MACRO sram_2_16_1_freepdk45
    CLASS RING ;
    ORIGIN 5.765 0.0 ;
    FOREIGN  sram 0.0 0.0 ;
    SIZE 19.165 BY 41.725 ;
    SYMMETRY X Y R90 ;
    PIN vdd 
        DIRECTION INOUT ; 
        USE POWER ; 
        SHAPE ABUTMENT ; 
        PORT             
        Layer metal1 ; 
        RECT  0.0 0.0 0.7 41.725 ;
        RECT  12.735 0.0 13.435 41.725 ;
        END             
    END vdd 
    PIN gnd 
        DIRECTION INOUT ; 
        USE GROUND ; 
        SHAPE ABUTMENT ; 
        PORT             
        Layer metal2 ; 
        RECT  8.89 0.0 9.59 41.725 ;
        END             
    END gnd 
    PIN DATA[0] 
        DIRECTION INOUT ; 
        PORT             
        Layer metal3 ; 
        RECT  11.4475 0.0 11.5175 3.22 ;
        RECT  11.4475 0.0 11.5175 0.135 ;
        END             
    END DATA[0] 
    PIN DATA[1] 
        DIRECTION INOUT ; 
        PORT             
        Layer metal3 ; 
        RECT  12.1525 0.0 12.2225 3.22 ;
        RECT  12.1525 0.0 12.2225 0.135 ;
        END             
    END DATA[1] 
    PIN ADDR[0] 
        DIRECTION INPUT ; 
        PORT             
        Layer metal3 ; 
        RECT  0.0 7.4525 0.9825 7.5225 ;
        END             
    END ADDR[0] 
    PIN ADDR[1] 
        DIRECTION INPUT ; 
        PORT             
        Layer metal3 ; 
        RECT  0.0 6.7475 0.9825 6.8175 ;
        END             
    END ADDR[1] 
    PIN ADDR[2] 
        DIRECTION INPUT ; 
        PORT             
        Layer metal3 ; 
        RECT  0.0 6.0425 0.9825 6.1125 ;
        END             
    END ADDR[2] 
    PIN ADDR[3] 
        DIRECTION INPUT ; 
        PORT             
        Layer metal3 ; 
        RECT  0.0 5.3375 0.9825 5.4075 ;
        END             
    END ADDR[3] 
    PIN CSb 
        DIRECTION INPUT ; 
        PORT             
        Layer metal3 ; 
        RECT  -5.4125 8.275 -5.3425 8.415 ;
        END             
    END CSb 
    PIN OEb 
        DIRECTION INPUT ; 
        PORT             
        Layer metal3 ; 
        RECT  -4.0025 8.275 -3.9325 8.415 ;
        END             
    END OEb 
    PIN WEb 
        DIRECTION INPUT ; 
        PORT             
        Layer metal3 ; 
        RECT  -4.7075 8.275 -4.6375 8.415 ;
        END             
    END WEb 
    PIN clk 
        DIRECTION INPUT ; 
        PORT             
        Layer metal3 ; 
        RECT  -2.0525 8.275 9.73 8.345 ;
        RECT  -2.085 8.275 -2.015 8.41 ;
        END             
    END clk 
    OBS 
        Layer  metal1 ; 
        RECT  -0.545 26.2325 0.0 26.2975 ;
        RECT  12.735 0.0 13.435 41.725 ;
        RECT  0.0 0.0 0.7 41.725 ;
        RECT  5.53 19.49 5.595 19.87 ;
        RECT  5.53 20.61 5.595 20.99 ;
        RECT  5.53 22.18 5.595 22.56 ;
        RECT  5.53 23.3 5.595 23.68 ;
        RECT  5.53 24.87 5.595 25.25 ;
        RECT  5.53 25.99 5.595 26.37 ;
        RECT  5.53 27.56 5.595 27.94 ;
        RECT  5.53 28.68 5.595 29.06 ;
        RECT  5.53 30.25 5.595 30.63 ;
        RECT  5.53 31.37 5.595 31.75 ;
        RECT  5.53 32.94 5.595 33.32 ;
        RECT  5.53 34.06 5.595 34.44 ;
        RECT  5.53 35.63 5.595 36.01 ;
        RECT  5.53 36.75 5.595 37.13 ;
        RECT  5.53 38.32 5.595 38.7 ;
        RECT  5.53 39.44 5.595 39.82 ;
        RECT  7.855 20.2075 11.13 20.2725 ;
        RECT  7.855 22.8975 11.13 22.9625 ;
        RECT  7.855 25.5875 11.13 25.6525 ;
        RECT  7.855 28.2775 11.13 28.3425 ;
        RECT  7.855 30.9675 11.13 31.0325 ;
        RECT  7.855 33.6575 11.13 33.7225 ;
        RECT  7.855 36.3475 11.13 36.4125 ;
        RECT  7.855 39.0375 11.13 39.1025 ;
        RECT  7.245 8.73 8.61 8.795 ;
        RECT  7.245 10.165 8.4 10.23 ;
        RECT  7.245 14.11 8.19 14.175 ;
        RECT  7.245 15.545 7.98 15.61 ;
        RECT  10.36 3.6 11.4825 3.665 ;
        RECT  9.94 1.415 11.5 1.48 ;
        RECT  10.15 2.9625 11.5 3.0275 ;
        RECT  10.36 41.1 11.13 41.165 ;
        RECT  10.57 10.1025 11.13 10.1675 ;
        RECT  10.78 14.1275 11.13 14.1925 ;
        RECT  11.13 20.2075 12.735 20.2725 ;
        RECT  11.13 22.8975 12.735 22.9625 ;
        RECT  11.13 25.5875 12.735 25.6525 ;
        RECT  11.13 28.2775 12.735 28.3425 ;
        RECT  11.13 30.9675 12.735 31.0325 ;
        RECT  11.13 33.6575 12.735 33.7225 ;
        RECT  11.13 36.3475 12.735 36.4125 ;
        RECT  11.13 39.0375 12.735 39.1025 ;
        RECT  11.13 41.66 12.735 41.725 ;
        RECT  11.13 18.7 12.735 18.765 ;
        RECT  11.13 10.2325 12.735 10.2975 ;
        RECT  11.13 9.565 12.735 9.63 ;
        RECT  11.5 1.545 12.735 1.61 ;
        RECT  12.17 1.545 12.735 1.61 ;
        RECT  0.0 20.2075 4.22 20.2725 ;
        RECT  0.0 22.8975 4.22 22.9625 ;
        RECT  0.0 25.5875 4.22 25.6525 ;
        RECT  0.0 28.2775 4.22 28.3425 ;
        RECT  0.0 30.9675 4.22 31.0325 ;
        RECT  0.0 33.6575 4.22 33.7225 ;
        RECT  0.0 36.3475 4.22 36.4125 ;
        RECT  0.0 39.0375 4.22 39.1025 ;
        RECT  0.0 12.1375 4.22 12.2025 ;
        RECT  0.0 17.5175 4.22 17.5825 ;
        RECT  8.89 40.545 12.54 40.61 ;
        RECT  9.385 0.355 12.54 0.42 ;
        RECT  4.22 13.4825 8.89 13.5475 ;
        RECT  4.22 18.8625 8.89 18.9275 ;
        RECT  7.35 7.8075 8.89 7.8725 ;
        RECT  7.35 6.3975 8.89 6.4625 ;
        RECT  7.35 6.3975 8.89 6.4625 ;
        RECT  7.35 4.9875 8.89 5.0525 ;
        RECT  11.8 20.0075 11.865 20.1425 ;
        RECT  11.615 20.0075 11.68 20.1425 ;
        RECT  11.1 20.0075 11.165 20.1425 ;
        RECT  11.285 20.0075 11.35 20.1425 ;
        RECT  11.615 19.5425 11.68 19.6775 ;
        RECT  11.8 19.5425 11.865 19.6775 ;
        RECT  11.285 19.5425 11.35 19.6775 ;
        RECT  11.1 19.5425 11.165 19.6775 ;
        RECT  11.72 19.1525 11.785 19.2875 ;
        RECT  11.535 19.1525 11.6 19.2875 ;
        RECT  11.365 19.1525 11.43 19.2875 ;
        RECT  11.18 19.1525 11.245 19.2875 ;
        RECT  11.8025 19.645 11.8675 19.78 ;
        RECT  11.8025 19.645 11.8675 19.78 ;
        RECT  11.8025 19.645 11.8675 19.78 ;
        RECT  11.8025 19.645 11.8675 19.78 ;
        RECT  11.8025 19.645 11.8675 19.78 ;
        RECT  11.8025 19.645 11.8675 19.78 ;
        RECT  11.41 20.2075 11.545 20.2725 ;
        RECT  11.0625 18.8625 11.1975 18.9275 ;
        RECT  11.7675 18.8625 11.9025 18.9275 ;
        RECT  11.3975 19.0025 11.5325 19.0675 ;
        RECT  11.8025 19.645 11.8675 19.78 ;
        RECT  11.8025 19.645 11.8675 19.78 ;
        RECT  11.8025 19.645 11.8675 19.78 ;
        RECT  11.8025 19.645 11.8675 19.78 ;
        RECT  11.3025 19.8925 11.4375 19.9575 ;
        RECT  11.3025 19.8925 11.4375 19.9575 ;
        RECT  11.5275 19.7425 11.6625 19.8075 ;
        RECT  11.5275 19.7425 11.6625 19.8075 ;
        RECT  11.8025 19.645 11.8675 19.78 ;
        RECT  11.8025 19.645 11.8675 19.78 ;
        RECT  11.8025 19.645 11.8675 19.78 ;
        RECT  11.8025 19.645 11.8675 19.78 ;
        RECT  11.3525 19.1525 11.4175 19.2875 ;
        RECT  11.0975 19.645 11.1625 19.78 ;
        RECT  11.0975 19.645 11.1625 19.78 ;
        RECT  11.0975 19.645 11.1625 19.78 ;
        RECT  11.0975 19.645 11.1625 19.78 ;
        RECT  11.0975 19.645 11.1625 19.78 ;
        RECT  11.0975 19.645 11.1625 19.78 ;
        RECT  11.8025 19.645 11.8675 19.78 ;
        RECT  11.8025 19.645 11.8675 19.78 ;
        RECT  11.8025 19.645 11.8675 19.78 ;
        RECT  11.8025 19.645 11.8675 19.78 ;
        RECT  11.5475 19.1525 11.6125 19.2875 ;
        RECT  11.415 18.8625 11.55 18.9275 ;
        RECT  11.415 18.8625 11.55 18.9275 ;
        RECT  11.7675 18.8625 11.9025 18.9275 ;
        RECT  11.41 20.2075 11.545 20.2725 ;
        RECT  11.7675 18.8625 11.9025 18.9275 ;
        RECT  11.7675 18.8625 11.9025 18.9275 ;
        RECT  11.8025 19.645 11.8675 19.78 ;
        RECT  11.8025 19.645 11.8675 19.78 ;
        RECT  11.8025 19.645 11.8675 19.78 ;
        RECT  11.8025 19.645 11.8675 19.78 ;
        RECT  11.8025 19.645 11.8675 19.78 ;
        RECT  11.8025 19.645 11.8675 19.78 ;
        RECT  11.0625 18.8625 11.1975 18.9275 ;
        RECT  11.4225 20.2075 11.5225 20.27 ;
        RECT  11.4225 20.21 11.5225 20.2725 ;
        RECT  11.75 19.005 11.8025 19.0675 ;
        RECT  11.4225 20.2075 11.5225 20.27 ;
        RECT  11.8 20.0075 11.87 20.2075 ;
        RECT  11.8 19.5425 11.87 19.6775 ;
        RECT  11.8 19.5425 11.87 19.6775 ;
        RECT  11.04 18.8625 11.925 18.9275 ;
        RECT  11.615 19.3775 11.79 19.4425 ;
        RECT  11.095 19.5425 11.165 19.6775 ;
        RECT  11.285 19.3775 11.35 20.1175 ;
        RECT  11.4225 20.21 11.5225 20.2725 ;
        RECT  11.045 19.005 11.0975 19.0675 ;
        RECT  11.8 19.5425 11.87 19.6775 ;
        RECT  11.04 20.2075 11.925 20.2725 ;
        RECT  11.615 19.3775 11.68 20.0075 ;
        RECT  11.8 19.5425 11.87 19.6775 ;
        RECT  11.8 19.5425 11.87 19.6775 ;
        RECT  11.18 19.1525 11.25 19.4425 ;
        RECT  11.095 19.5425 11.165 19.6775 ;
        RECT  11.04 19.0025 11.925 19.0675 ;
        RECT  11.8 19.5425 11.87 19.6775 ;
        RECT  11.8 20.0075 11.87 20.2075 ;
        RECT  11.095 20.0075 11.165 20.2075 ;
        RECT  11.72 19.1525 11.79 19.4425 ;
        RECT  11.18 19.3775 11.35 19.4425 ;
        RECT  11.8 20.3375 11.865 20.4725 ;
        RECT  11.615 20.3375 11.68 20.4725 ;
        RECT  11.1 20.3375 11.165 20.4725 ;
        RECT  11.285 20.3375 11.35 20.4725 ;
        RECT  11.615 20.8025 11.68 20.9375 ;
        RECT  11.8 20.8025 11.865 20.9375 ;
        RECT  11.285 20.8025 11.35 20.9375 ;
        RECT  11.1 20.8025 11.165 20.9375 ;
        RECT  11.72 21.1925 11.785 21.3275 ;
        RECT  11.535 21.1925 11.6 21.3275 ;
        RECT  11.365 21.1925 11.43 21.3275 ;
        RECT  11.18 21.1925 11.245 21.3275 ;
        RECT  11.8025 20.7 11.8675 20.835 ;
        RECT  11.8025 20.7 11.8675 20.835 ;
        RECT  11.8025 20.7 11.8675 20.835 ;
        RECT  11.8025 20.7 11.8675 20.835 ;
        RECT  11.8025 20.7 11.8675 20.835 ;
        RECT  11.8025 20.7 11.8675 20.835 ;
        RECT  11.41 20.2075 11.545 20.2725 ;
        RECT  11.0625 21.5525 11.1975 21.6175 ;
        RECT  11.7675 21.5525 11.9025 21.6175 ;
        RECT  11.3975 21.4125 11.5325 21.4775 ;
        RECT  11.8025 20.7 11.8675 20.835 ;
        RECT  11.8025 20.7 11.8675 20.835 ;
        RECT  11.8025 20.7 11.8675 20.835 ;
        RECT  11.8025 20.7 11.8675 20.835 ;
        RECT  11.3025 20.5225 11.4375 20.5875 ;
        RECT  11.3025 20.5225 11.4375 20.5875 ;
        RECT  11.5275 20.6725 11.6625 20.7375 ;
        RECT  11.5275 20.6725 11.6625 20.7375 ;
        RECT  11.8025 20.7 11.8675 20.835 ;
        RECT  11.8025 20.7 11.8675 20.835 ;
        RECT  11.8025 20.7 11.8675 20.835 ;
        RECT  11.8025 20.7 11.8675 20.835 ;
        RECT  11.3525 21.1925 11.4175 21.3275 ;
        RECT  11.0975 20.7 11.1625 20.835 ;
        RECT  11.0975 20.7 11.1625 20.835 ;
        RECT  11.0975 20.7 11.1625 20.835 ;
        RECT  11.0975 20.7 11.1625 20.835 ;
        RECT  11.0975 20.7 11.1625 20.835 ;
        RECT  11.0975 20.7 11.1625 20.835 ;
        RECT  11.8025 20.7 11.8675 20.835 ;
        RECT  11.8025 20.7 11.8675 20.835 ;
        RECT  11.8025 20.7 11.8675 20.835 ;
        RECT  11.8025 20.7 11.8675 20.835 ;
        RECT  11.5475 21.1925 11.6125 21.3275 ;
        RECT  11.415 21.5525 11.55 21.6175 ;
        RECT  11.415 21.5525 11.55 21.6175 ;
        RECT  11.7675 21.5525 11.9025 21.6175 ;
        RECT  11.41 20.2075 11.545 20.2725 ;
        RECT  11.7675 21.5525 11.9025 21.6175 ;
        RECT  11.7675 21.5525 11.9025 21.6175 ;
        RECT  11.8025 20.7 11.8675 20.835 ;
        RECT  11.8025 20.7 11.8675 20.835 ;
        RECT  11.8025 20.7 11.8675 20.835 ;
        RECT  11.8025 20.7 11.8675 20.835 ;
        RECT  11.8025 20.7 11.8675 20.835 ;
        RECT  11.8025 20.7 11.8675 20.835 ;
        RECT  11.0625 21.5525 11.1975 21.6175 ;
        RECT  11.4225 20.21 11.5225 20.2725 ;
        RECT  11.4225 20.2075 11.5225 20.27 ;
        RECT  11.75 21.4125 11.8025 21.475 ;
        RECT  11.4225 20.21 11.5225 20.2725 ;
        RECT  11.8 20.2725 11.87 20.4725 ;
        RECT  11.8 20.8025 11.87 20.9375 ;
        RECT  11.8 20.8025 11.87 20.9375 ;
        RECT  11.04 21.5525 11.925 21.6175 ;
        RECT  11.615 21.0375 11.79 21.1025 ;
        RECT  11.095 20.8025 11.165 20.9375 ;
        RECT  11.285 20.3625 11.35 21.1025 ;
        RECT  11.4225 20.2075 11.5225 20.27 ;
        RECT  11.045 21.4125 11.0975 21.475 ;
        RECT  11.8 20.8025 11.87 20.9375 ;
        RECT  11.04 20.2075 11.925 20.2725 ;
        RECT  11.615 20.4725 11.68 21.1025 ;
        RECT  11.8 20.8025 11.87 20.9375 ;
        RECT  11.8 20.8025 11.87 20.9375 ;
        RECT  11.18 21.0375 11.25 21.3275 ;
        RECT  11.095 20.8025 11.165 20.9375 ;
        RECT  11.04 21.4125 11.925 21.4775 ;
        RECT  11.8 20.8025 11.87 20.9375 ;
        RECT  11.8 20.2725 11.87 20.4725 ;
        RECT  11.095 20.2725 11.165 20.4725 ;
        RECT  11.72 21.0375 11.79 21.3275 ;
        RECT  11.18 21.0375 11.35 21.1025 ;
        RECT  11.8 22.6975 11.865 22.8325 ;
        RECT  11.615 22.6975 11.68 22.8325 ;
        RECT  11.1 22.6975 11.165 22.8325 ;
        RECT  11.285 22.6975 11.35 22.8325 ;
        RECT  11.615 22.2325 11.68 22.3675 ;
        RECT  11.8 22.2325 11.865 22.3675 ;
        RECT  11.285 22.2325 11.35 22.3675 ;
        RECT  11.1 22.2325 11.165 22.3675 ;
        RECT  11.72 21.8425 11.785 21.9775 ;
        RECT  11.535 21.8425 11.6 21.9775 ;
        RECT  11.365 21.8425 11.43 21.9775 ;
        RECT  11.18 21.8425 11.245 21.9775 ;
        RECT  11.8025 22.335 11.8675 22.47 ;
        RECT  11.8025 22.335 11.8675 22.47 ;
        RECT  11.8025 22.335 11.8675 22.47 ;
        RECT  11.8025 22.335 11.8675 22.47 ;
        RECT  11.8025 22.335 11.8675 22.47 ;
        RECT  11.8025 22.335 11.8675 22.47 ;
        RECT  11.41 22.8975 11.545 22.9625 ;
        RECT  11.0625 21.5525 11.1975 21.6175 ;
        RECT  11.7675 21.5525 11.9025 21.6175 ;
        RECT  11.3975 21.6925 11.5325 21.7575 ;
        RECT  11.8025 22.335 11.8675 22.47 ;
        RECT  11.8025 22.335 11.8675 22.47 ;
        RECT  11.8025 22.335 11.8675 22.47 ;
        RECT  11.8025 22.335 11.8675 22.47 ;
        RECT  11.3025 22.5825 11.4375 22.6475 ;
        RECT  11.3025 22.5825 11.4375 22.6475 ;
        RECT  11.5275 22.4325 11.6625 22.4975 ;
        RECT  11.5275 22.4325 11.6625 22.4975 ;
        RECT  11.8025 22.335 11.8675 22.47 ;
        RECT  11.8025 22.335 11.8675 22.47 ;
        RECT  11.8025 22.335 11.8675 22.47 ;
        RECT  11.8025 22.335 11.8675 22.47 ;
        RECT  11.3525 21.8425 11.4175 21.9775 ;
        RECT  11.0975 22.335 11.1625 22.47 ;
        RECT  11.0975 22.335 11.1625 22.47 ;
        RECT  11.0975 22.335 11.1625 22.47 ;
        RECT  11.0975 22.335 11.1625 22.47 ;
        RECT  11.0975 22.335 11.1625 22.47 ;
        RECT  11.0975 22.335 11.1625 22.47 ;
        RECT  11.8025 22.335 11.8675 22.47 ;
        RECT  11.8025 22.335 11.8675 22.47 ;
        RECT  11.8025 22.335 11.8675 22.47 ;
        RECT  11.8025 22.335 11.8675 22.47 ;
        RECT  11.5475 21.8425 11.6125 21.9775 ;
        RECT  11.415 21.5525 11.55 21.6175 ;
        RECT  11.415 21.5525 11.55 21.6175 ;
        RECT  11.7675 21.5525 11.9025 21.6175 ;
        RECT  11.41 22.8975 11.545 22.9625 ;
        RECT  11.7675 21.5525 11.9025 21.6175 ;
        RECT  11.7675 21.5525 11.9025 21.6175 ;
        RECT  11.8025 22.335 11.8675 22.47 ;
        RECT  11.8025 22.335 11.8675 22.47 ;
        RECT  11.8025 22.335 11.8675 22.47 ;
        RECT  11.8025 22.335 11.8675 22.47 ;
        RECT  11.8025 22.335 11.8675 22.47 ;
        RECT  11.8025 22.335 11.8675 22.47 ;
        RECT  11.0625 21.5525 11.1975 21.6175 ;
        RECT  11.4225 22.8975 11.5225 22.96 ;
        RECT  11.4225 22.9 11.5225 22.9625 ;
        RECT  11.75 21.695 11.8025 21.7575 ;
        RECT  11.4225 22.8975 11.5225 22.96 ;
        RECT  11.8 22.6975 11.87 22.8975 ;
        RECT  11.8 22.2325 11.87 22.3675 ;
        RECT  11.8 22.2325 11.87 22.3675 ;
        RECT  11.04 21.5525 11.925 21.6175 ;
        RECT  11.615 22.0675 11.79 22.1325 ;
        RECT  11.095 22.2325 11.165 22.3675 ;
        RECT  11.285 22.0675 11.35 22.8075 ;
        RECT  11.4225 22.9 11.5225 22.9625 ;
        RECT  11.045 21.695 11.0975 21.7575 ;
        RECT  11.8 22.2325 11.87 22.3675 ;
        RECT  11.04 22.8975 11.925 22.9625 ;
        RECT  11.615 22.0675 11.68 22.6975 ;
        RECT  11.8 22.2325 11.87 22.3675 ;
        RECT  11.8 22.2325 11.87 22.3675 ;
        RECT  11.18 21.8425 11.25 22.1325 ;
        RECT  11.095 22.2325 11.165 22.3675 ;
        RECT  11.04 21.6925 11.925 21.7575 ;
        RECT  11.8 22.2325 11.87 22.3675 ;
        RECT  11.8 22.6975 11.87 22.8975 ;
        RECT  11.095 22.6975 11.165 22.8975 ;
        RECT  11.72 21.8425 11.79 22.1325 ;
        RECT  11.18 22.0675 11.35 22.1325 ;
        RECT  11.8 23.0275 11.865 23.1625 ;
        RECT  11.615 23.0275 11.68 23.1625 ;
        RECT  11.1 23.0275 11.165 23.1625 ;
        RECT  11.285 23.0275 11.35 23.1625 ;
        RECT  11.615 23.4925 11.68 23.6275 ;
        RECT  11.8 23.4925 11.865 23.6275 ;
        RECT  11.285 23.4925 11.35 23.6275 ;
        RECT  11.1 23.4925 11.165 23.6275 ;
        RECT  11.72 23.8825 11.785 24.0175 ;
        RECT  11.535 23.8825 11.6 24.0175 ;
        RECT  11.365 23.8825 11.43 24.0175 ;
        RECT  11.18 23.8825 11.245 24.0175 ;
        RECT  11.8025 23.39 11.8675 23.525 ;
        RECT  11.8025 23.39 11.8675 23.525 ;
        RECT  11.8025 23.39 11.8675 23.525 ;
        RECT  11.8025 23.39 11.8675 23.525 ;
        RECT  11.8025 23.39 11.8675 23.525 ;
        RECT  11.8025 23.39 11.8675 23.525 ;
        RECT  11.41 22.8975 11.545 22.9625 ;
        RECT  11.0625 24.2425 11.1975 24.3075 ;
        RECT  11.7675 24.2425 11.9025 24.3075 ;
        RECT  11.3975 24.1025 11.5325 24.1675 ;
        RECT  11.8025 23.39 11.8675 23.525 ;
        RECT  11.8025 23.39 11.8675 23.525 ;
        RECT  11.8025 23.39 11.8675 23.525 ;
        RECT  11.8025 23.39 11.8675 23.525 ;
        RECT  11.3025 23.2125 11.4375 23.2775 ;
        RECT  11.3025 23.2125 11.4375 23.2775 ;
        RECT  11.5275 23.3625 11.6625 23.4275 ;
        RECT  11.5275 23.3625 11.6625 23.4275 ;
        RECT  11.8025 23.39 11.8675 23.525 ;
        RECT  11.8025 23.39 11.8675 23.525 ;
        RECT  11.8025 23.39 11.8675 23.525 ;
        RECT  11.8025 23.39 11.8675 23.525 ;
        RECT  11.3525 23.8825 11.4175 24.0175 ;
        RECT  11.0975 23.39 11.1625 23.525 ;
        RECT  11.0975 23.39 11.1625 23.525 ;
        RECT  11.0975 23.39 11.1625 23.525 ;
        RECT  11.0975 23.39 11.1625 23.525 ;
        RECT  11.0975 23.39 11.1625 23.525 ;
        RECT  11.0975 23.39 11.1625 23.525 ;
        RECT  11.8025 23.39 11.8675 23.525 ;
        RECT  11.8025 23.39 11.8675 23.525 ;
        RECT  11.8025 23.39 11.8675 23.525 ;
        RECT  11.8025 23.39 11.8675 23.525 ;
        RECT  11.5475 23.8825 11.6125 24.0175 ;
        RECT  11.415 24.2425 11.55 24.3075 ;
        RECT  11.415 24.2425 11.55 24.3075 ;
        RECT  11.7675 24.2425 11.9025 24.3075 ;
        RECT  11.41 22.8975 11.545 22.9625 ;
        RECT  11.7675 24.2425 11.9025 24.3075 ;
        RECT  11.7675 24.2425 11.9025 24.3075 ;
        RECT  11.8025 23.39 11.8675 23.525 ;
        RECT  11.8025 23.39 11.8675 23.525 ;
        RECT  11.8025 23.39 11.8675 23.525 ;
        RECT  11.8025 23.39 11.8675 23.525 ;
        RECT  11.8025 23.39 11.8675 23.525 ;
        RECT  11.8025 23.39 11.8675 23.525 ;
        RECT  11.0625 24.2425 11.1975 24.3075 ;
        RECT  11.4225 22.9 11.5225 22.9625 ;
        RECT  11.4225 22.8975 11.5225 22.96 ;
        RECT  11.75 24.1025 11.8025 24.165 ;
        RECT  11.4225 22.9 11.5225 22.9625 ;
        RECT  11.8 22.9625 11.87 23.1625 ;
        RECT  11.8 23.4925 11.87 23.6275 ;
        RECT  11.8 23.4925 11.87 23.6275 ;
        RECT  11.04 24.2425 11.925 24.3075 ;
        RECT  11.615 23.7275 11.79 23.7925 ;
        RECT  11.095 23.4925 11.165 23.6275 ;
        RECT  11.285 23.0525 11.35 23.7925 ;
        RECT  11.4225 22.8975 11.5225 22.96 ;
        RECT  11.045 24.1025 11.0975 24.165 ;
        RECT  11.8 23.4925 11.87 23.6275 ;
        RECT  11.04 22.8975 11.925 22.9625 ;
        RECT  11.615 23.1625 11.68 23.7925 ;
        RECT  11.8 23.4925 11.87 23.6275 ;
        RECT  11.8 23.4925 11.87 23.6275 ;
        RECT  11.18 23.7275 11.25 24.0175 ;
        RECT  11.095 23.4925 11.165 23.6275 ;
        RECT  11.04 24.1025 11.925 24.1675 ;
        RECT  11.8 23.4925 11.87 23.6275 ;
        RECT  11.8 22.9625 11.87 23.1625 ;
        RECT  11.095 22.9625 11.165 23.1625 ;
        RECT  11.72 23.7275 11.79 24.0175 ;
        RECT  11.18 23.7275 11.35 23.7925 ;
        RECT  11.8 25.3875 11.865 25.5225 ;
        RECT  11.615 25.3875 11.68 25.5225 ;
        RECT  11.1 25.3875 11.165 25.5225 ;
        RECT  11.285 25.3875 11.35 25.5225 ;
        RECT  11.615 24.9225 11.68 25.0575 ;
        RECT  11.8 24.9225 11.865 25.0575 ;
        RECT  11.285 24.9225 11.35 25.0575 ;
        RECT  11.1 24.9225 11.165 25.0575 ;
        RECT  11.72 24.5325 11.785 24.6675 ;
        RECT  11.535 24.5325 11.6 24.6675 ;
        RECT  11.365 24.5325 11.43 24.6675 ;
        RECT  11.18 24.5325 11.245 24.6675 ;
        RECT  11.8025 25.025 11.8675 25.16 ;
        RECT  11.8025 25.025 11.8675 25.16 ;
        RECT  11.8025 25.025 11.8675 25.16 ;
        RECT  11.8025 25.025 11.8675 25.16 ;
        RECT  11.8025 25.025 11.8675 25.16 ;
        RECT  11.8025 25.025 11.8675 25.16 ;
        RECT  11.41 25.5875 11.545 25.6525 ;
        RECT  11.0625 24.2425 11.1975 24.3075 ;
        RECT  11.7675 24.2425 11.9025 24.3075 ;
        RECT  11.3975 24.3825 11.5325 24.4475 ;
        RECT  11.8025 25.025 11.8675 25.16 ;
        RECT  11.8025 25.025 11.8675 25.16 ;
        RECT  11.8025 25.025 11.8675 25.16 ;
        RECT  11.8025 25.025 11.8675 25.16 ;
        RECT  11.3025 25.2725 11.4375 25.3375 ;
        RECT  11.3025 25.2725 11.4375 25.3375 ;
        RECT  11.5275 25.1225 11.6625 25.1875 ;
        RECT  11.5275 25.1225 11.6625 25.1875 ;
        RECT  11.8025 25.025 11.8675 25.16 ;
        RECT  11.8025 25.025 11.8675 25.16 ;
        RECT  11.8025 25.025 11.8675 25.16 ;
        RECT  11.8025 25.025 11.8675 25.16 ;
        RECT  11.3525 24.5325 11.4175 24.6675 ;
        RECT  11.0975 25.025 11.1625 25.16 ;
        RECT  11.0975 25.025 11.1625 25.16 ;
        RECT  11.0975 25.025 11.1625 25.16 ;
        RECT  11.0975 25.025 11.1625 25.16 ;
        RECT  11.0975 25.025 11.1625 25.16 ;
        RECT  11.0975 25.025 11.1625 25.16 ;
        RECT  11.8025 25.025 11.8675 25.16 ;
        RECT  11.8025 25.025 11.8675 25.16 ;
        RECT  11.8025 25.025 11.8675 25.16 ;
        RECT  11.8025 25.025 11.8675 25.16 ;
        RECT  11.5475 24.5325 11.6125 24.6675 ;
        RECT  11.415 24.2425 11.55 24.3075 ;
        RECT  11.415 24.2425 11.55 24.3075 ;
        RECT  11.7675 24.2425 11.9025 24.3075 ;
        RECT  11.41 25.5875 11.545 25.6525 ;
        RECT  11.7675 24.2425 11.9025 24.3075 ;
        RECT  11.7675 24.2425 11.9025 24.3075 ;
        RECT  11.8025 25.025 11.8675 25.16 ;
        RECT  11.8025 25.025 11.8675 25.16 ;
        RECT  11.8025 25.025 11.8675 25.16 ;
        RECT  11.8025 25.025 11.8675 25.16 ;
        RECT  11.8025 25.025 11.8675 25.16 ;
        RECT  11.8025 25.025 11.8675 25.16 ;
        RECT  11.0625 24.2425 11.1975 24.3075 ;
        RECT  11.4225 25.5875 11.5225 25.65 ;
        RECT  11.4225 25.59 11.5225 25.6525 ;
        RECT  11.75 24.385 11.8025 24.4475 ;
        RECT  11.4225 25.5875 11.5225 25.65 ;
        RECT  11.8 25.3875 11.87 25.5875 ;
        RECT  11.8 24.9225 11.87 25.0575 ;
        RECT  11.8 24.9225 11.87 25.0575 ;
        RECT  11.04 24.2425 11.925 24.3075 ;
        RECT  11.615 24.7575 11.79 24.8225 ;
        RECT  11.095 24.9225 11.165 25.0575 ;
        RECT  11.285 24.7575 11.35 25.4975 ;
        RECT  11.4225 25.59 11.5225 25.6525 ;
        RECT  11.045 24.385 11.0975 24.4475 ;
        RECT  11.8 24.9225 11.87 25.0575 ;
        RECT  11.04 25.5875 11.925 25.6525 ;
        RECT  11.615 24.7575 11.68 25.3875 ;
        RECT  11.8 24.9225 11.87 25.0575 ;
        RECT  11.8 24.9225 11.87 25.0575 ;
        RECT  11.18 24.5325 11.25 24.8225 ;
        RECT  11.095 24.9225 11.165 25.0575 ;
        RECT  11.04 24.3825 11.925 24.4475 ;
        RECT  11.8 24.9225 11.87 25.0575 ;
        RECT  11.8 25.3875 11.87 25.5875 ;
        RECT  11.095 25.3875 11.165 25.5875 ;
        RECT  11.72 24.5325 11.79 24.8225 ;
        RECT  11.18 24.7575 11.35 24.8225 ;
        RECT  11.8 25.7175 11.865 25.8525 ;
        RECT  11.615 25.7175 11.68 25.8525 ;
        RECT  11.1 25.7175 11.165 25.8525 ;
        RECT  11.285 25.7175 11.35 25.8525 ;
        RECT  11.615 26.1825 11.68 26.3175 ;
        RECT  11.8 26.1825 11.865 26.3175 ;
        RECT  11.285 26.1825 11.35 26.3175 ;
        RECT  11.1 26.1825 11.165 26.3175 ;
        RECT  11.72 26.5725 11.785 26.7075 ;
        RECT  11.535 26.5725 11.6 26.7075 ;
        RECT  11.365 26.5725 11.43 26.7075 ;
        RECT  11.18 26.5725 11.245 26.7075 ;
        RECT  11.8025 26.08 11.8675 26.215 ;
        RECT  11.8025 26.08 11.8675 26.215 ;
        RECT  11.8025 26.08 11.8675 26.215 ;
        RECT  11.8025 26.08 11.8675 26.215 ;
        RECT  11.8025 26.08 11.8675 26.215 ;
        RECT  11.8025 26.08 11.8675 26.215 ;
        RECT  11.41 25.5875 11.545 25.6525 ;
        RECT  11.0625 26.9325 11.1975 26.9975 ;
        RECT  11.7675 26.9325 11.9025 26.9975 ;
        RECT  11.3975 26.7925 11.5325 26.8575 ;
        RECT  11.8025 26.08 11.8675 26.215 ;
        RECT  11.8025 26.08 11.8675 26.215 ;
        RECT  11.8025 26.08 11.8675 26.215 ;
        RECT  11.8025 26.08 11.8675 26.215 ;
        RECT  11.3025 25.9025 11.4375 25.9675 ;
        RECT  11.3025 25.9025 11.4375 25.9675 ;
        RECT  11.5275 26.0525 11.6625 26.1175 ;
        RECT  11.5275 26.0525 11.6625 26.1175 ;
        RECT  11.8025 26.08 11.8675 26.215 ;
        RECT  11.8025 26.08 11.8675 26.215 ;
        RECT  11.8025 26.08 11.8675 26.215 ;
        RECT  11.8025 26.08 11.8675 26.215 ;
        RECT  11.3525 26.5725 11.4175 26.7075 ;
        RECT  11.0975 26.08 11.1625 26.215 ;
        RECT  11.0975 26.08 11.1625 26.215 ;
        RECT  11.0975 26.08 11.1625 26.215 ;
        RECT  11.0975 26.08 11.1625 26.215 ;
        RECT  11.0975 26.08 11.1625 26.215 ;
        RECT  11.0975 26.08 11.1625 26.215 ;
        RECT  11.8025 26.08 11.8675 26.215 ;
        RECT  11.8025 26.08 11.8675 26.215 ;
        RECT  11.8025 26.08 11.8675 26.215 ;
        RECT  11.8025 26.08 11.8675 26.215 ;
        RECT  11.5475 26.5725 11.6125 26.7075 ;
        RECT  11.415 26.9325 11.55 26.9975 ;
        RECT  11.415 26.9325 11.55 26.9975 ;
        RECT  11.7675 26.9325 11.9025 26.9975 ;
        RECT  11.41 25.5875 11.545 25.6525 ;
        RECT  11.7675 26.9325 11.9025 26.9975 ;
        RECT  11.7675 26.9325 11.9025 26.9975 ;
        RECT  11.8025 26.08 11.8675 26.215 ;
        RECT  11.8025 26.08 11.8675 26.215 ;
        RECT  11.8025 26.08 11.8675 26.215 ;
        RECT  11.8025 26.08 11.8675 26.215 ;
        RECT  11.8025 26.08 11.8675 26.215 ;
        RECT  11.8025 26.08 11.8675 26.215 ;
        RECT  11.0625 26.9325 11.1975 26.9975 ;
        RECT  11.4225 25.59 11.5225 25.6525 ;
        RECT  11.4225 25.5875 11.5225 25.65 ;
        RECT  11.75 26.7925 11.8025 26.855 ;
        RECT  11.4225 25.59 11.5225 25.6525 ;
        RECT  11.8 25.6525 11.87 25.8525 ;
        RECT  11.8 26.1825 11.87 26.3175 ;
        RECT  11.8 26.1825 11.87 26.3175 ;
        RECT  11.04 26.9325 11.925 26.9975 ;
        RECT  11.615 26.4175 11.79 26.4825 ;
        RECT  11.095 26.1825 11.165 26.3175 ;
        RECT  11.285 25.7425 11.35 26.4825 ;
        RECT  11.4225 25.5875 11.5225 25.65 ;
        RECT  11.045 26.7925 11.0975 26.855 ;
        RECT  11.8 26.1825 11.87 26.3175 ;
        RECT  11.04 25.5875 11.925 25.6525 ;
        RECT  11.615 25.8525 11.68 26.4825 ;
        RECT  11.8 26.1825 11.87 26.3175 ;
        RECT  11.8 26.1825 11.87 26.3175 ;
        RECT  11.18 26.4175 11.25 26.7075 ;
        RECT  11.095 26.1825 11.165 26.3175 ;
        RECT  11.04 26.7925 11.925 26.8575 ;
        RECT  11.8 26.1825 11.87 26.3175 ;
        RECT  11.8 25.6525 11.87 25.8525 ;
        RECT  11.095 25.6525 11.165 25.8525 ;
        RECT  11.72 26.4175 11.79 26.7075 ;
        RECT  11.18 26.4175 11.35 26.4825 ;
        RECT  11.8 28.0775 11.865 28.2125 ;
        RECT  11.615 28.0775 11.68 28.2125 ;
        RECT  11.1 28.0775 11.165 28.2125 ;
        RECT  11.285 28.0775 11.35 28.2125 ;
        RECT  11.615 27.6125 11.68 27.7475 ;
        RECT  11.8 27.6125 11.865 27.7475 ;
        RECT  11.285 27.6125 11.35 27.7475 ;
        RECT  11.1 27.6125 11.165 27.7475 ;
        RECT  11.72 27.2225 11.785 27.3575 ;
        RECT  11.535 27.2225 11.6 27.3575 ;
        RECT  11.365 27.2225 11.43 27.3575 ;
        RECT  11.18 27.2225 11.245 27.3575 ;
        RECT  11.8025 27.715 11.8675 27.85 ;
        RECT  11.8025 27.715 11.8675 27.85 ;
        RECT  11.8025 27.715 11.8675 27.85 ;
        RECT  11.8025 27.715 11.8675 27.85 ;
        RECT  11.8025 27.715 11.8675 27.85 ;
        RECT  11.8025 27.715 11.8675 27.85 ;
        RECT  11.41 28.2775 11.545 28.3425 ;
        RECT  11.0625 26.9325 11.1975 26.9975 ;
        RECT  11.7675 26.9325 11.9025 26.9975 ;
        RECT  11.3975 27.0725 11.5325 27.1375 ;
        RECT  11.8025 27.715 11.8675 27.85 ;
        RECT  11.8025 27.715 11.8675 27.85 ;
        RECT  11.8025 27.715 11.8675 27.85 ;
        RECT  11.8025 27.715 11.8675 27.85 ;
        RECT  11.3025 27.9625 11.4375 28.0275 ;
        RECT  11.3025 27.9625 11.4375 28.0275 ;
        RECT  11.5275 27.8125 11.6625 27.8775 ;
        RECT  11.5275 27.8125 11.6625 27.8775 ;
        RECT  11.8025 27.715 11.8675 27.85 ;
        RECT  11.8025 27.715 11.8675 27.85 ;
        RECT  11.8025 27.715 11.8675 27.85 ;
        RECT  11.8025 27.715 11.8675 27.85 ;
        RECT  11.3525 27.2225 11.4175 27.3575 ;
        RECT  11.0975 27.715 11.1625 27.85 ;
        RECT  11.0975 27.715 11.1625 27.85 ;
        RECT  11.0975 27.715 11.1625 27.85 ;
        RECT  11.0975 27.715 11.1625 27.85 ;
        RECT  11.0975 27.715 11.1625 27.85 ;
        RECT  11.0975 27.715 11.1625 27.85 ;
        RECT  11.8025 27.715 11.8675 27.85 ;
        RECT  11.8025 27.715 11.8675 27.85 ;
        RECT  11.8025 27.715 11.8675 27.85 ;
        RECT  11.8025 27.715 11.8675 27.85 ;
        RECT  11.5475 27.2225 11.6125 27.3575 ;
        RECT  11.415 26.9325 11.55 26.9975 ;
        RECT  11.415 26.9325 11.55 26.9975 ;
        RECT  11.7675 26.9325 11.9025 26.9975 ;
        RECT  11.41 28.2775 11.545 28.3425 ;
        RECT  11.7675 26.9325 11.9025 26.9975 ;
        RECT  11.7675 26.9325 11.9025 26.9975 ;
        RECT  11.8025 27.715 11.8675 27.85 ;
        RECT  11.8025 27.715 11.8675 27.85 ;
        RECT  11.8025 27.715 11.8675 27.85 ;
        RECT  11.8025 27.715 11.8675 27.85 ;
        RECT  11.8025 27.715 11.8675 27.85 ;
        RECT  11.8025 27.715 11.8675 27.85 ;
        RECT  11.0625 26.9325 11.1975 26.9975 ;
        RECT  11.4225 28.2775 11.5225 28.34 ;
        RECT  11.4225 28.28 11.5225 28.3425 ;
        RECT  11.75 27.075 11.8025 27.1375 ;
        RECT  11.4225 28.2775 11.5225 28.34 ;
        RECT  11.8 28.0775 11.87 28.2775 ;
        RECT  11.8 27.6125 11.87 27.7475 ;
        RECT  11.8 27.6125 11.87 27.7475 ;
        RECT  11.04 26.9325 11.925 26.9975 ;
        RECT  11.615 27.4475 11.79 27.5125 ;
        RECT  11.095 27.6125 11.165 27.7475 ;
        RECT  11.285 27.4475 11.35 28.1875 ;
        RECT  11.4225 28.28 11.5225 28.3425 ;
        RECT  11.045 27.075 11.0975 27.1375 ;
        RECT  11.8 27.6125 11.87 27.7475 ;
        RECT  11.04 28.2775 11.925 28.3425 ;
        RECT  11.615 27.4475 11.68 28.0775 ;
        RECT  11.8 27.6125 11.87 27.7475 ;
        RECT  11.8 27.6125 11.87 27.7475 ;
        RECT  11.18 27.2225 11.25 27.5125 ;
        RECT  11.095 27.6125 11.165 27.7475 ;
        RECT  11.04 27.0725 11.925 27.1375 ;
        RECT  11.8 27.6125 11.87 27.7475 ;
        RECT  11.8 28.0775 11.87 28.2775 ;
        RECT  11.095 28.0775 11.165 28.2775 ;
        RECT  11.72 27.2225 11.79 27.5125 ;
        RECT  11.18 27.4475 11.35 27.5125 ;
        RECT  11.8 28.4075 11.865 28.5425 ;
        RECT  11.615 28.4075 11.68 28.5425 ;
        RECT  11.1 28.4075 11.165 28.5425 ;
        RECT  11.285 28.4075 11.35 28.5425 ;
        RECT  11.615 28.8725 11.68 29.0075 ;
        RECT  11.8 28.8725 11.865 29.0075 ;
        RECT  11.285 28.8725 11.35 29.0075 ;
        RECT  11.1 28.8725 11.165 29.0075 ;
        RECT  11.72 29.2625 11.785 29.3975 ;
        RECT  11.535 29.2625 11.6 29.3975 ;
        RECT  11.365 29.2625 11.43 29.3975 ;
        RECT  11.18 29.2625 11.245 29.3975 ;
        RECT  11.8025 28.77 11.8675 28.905 ;
        RECT  11.8025 28.77 11.8675 28.905 ;
        RECT  11.8025 28.77 11.8675 28.905 ;
        RECT  11.8025 28.77 11.8675 28.905 ;
        RECT  11.8025 28.77 11.8675 28.905 ;
        RECT  11.8025 28.77 11.8675 28.905 ;
        RECT  11.41 28.2775 11.545 28.3425 ;
        RECT  11.0625 29.6225 11.1975 29.6875 ;
        RECT  11.7675 29.6225 11.9025 29.6875 ;
        RECT  11.3975 29.4825 11.5325 29.5475 ;
        RECT  11.8025 28.77 11.8675 28.905 ;
        RECT  11.8025 28.77 11.8675 28.905 ;
        RECT  11.8025 28.77 11.8675 28.905 ;
        RECT  11.8025 28.77 11.8675 28.905 ;
        RECT  11.3025 28.5925 11.4375 28.6575 ;
        RECT  11.3025 28.5925 11.4375 28.6575 ;
        RECT  11.5275 28.7425 11.6625 28.8075 ;
        RECT  11.5275 28.7425 11.6625 28.8075 ;
        RECT  11.8025 28.77 11.8675 28.905 ;
        RECT  11.8025 28.77 11.8675 28.905 ;
        RECT  11.8025 28.77 11.8675 28.905 ;
        RECT  11.8025 28.77 11.8675 28.905 ;
        RECT  11.3525 29.2625 11.4175 29.3975 ;
        RECT  11.0975 28.77 11.1625 28.905 ;
        RECT  11.0975 28.77 11.1625 28.905 ;
        RECT  11.0975 28.77 11.1625 28.905 ;
        RECT  11.0975 28.77 11.1625 28.905 ;
        RECT  11.0975 28.77 11.1625 28.905 ;
        RECT  11.0975 28.77 11.1625 28.905 ;
        RECT  11.8025 28.77 11.8675 28.905 ;
        RECT  11.8025 28.77 11.8675 28.905 ;
        RECT  11.8025 28.77 11.8675 28.905 ;
        RECT  11.8025 28.77 11.8675 28.905 ;
        RECT  11.5475 29.2625 11.6125 29.3975 ;
        RECT  11.415 29.6225 11.55 29.6875 ;
        RECT  11.415 29.6225 11.55 29.6875 ;
        RECT  11.7675 29.6225 11.9025 29.6875 ;
        RECT  11.41 28.2775 11.545 28.3425 ;
        RECT  11.7675 29.6225 11.9025 29.6875 ;
        RECT  11.7675 29.6225 11.9025 29.6875 ;
        RECT  11.8025 28.77 11.8675 28.905 ;
        RECT  11.8025 28.77 11.8675 28.905 ;
        RECT  11.8025 28.77 11.8675 28.905 ;
        RECT  11.8025 28.77 11.8675 28.905 ;
        RECT  11.8025 28.77 11.8675 28.905 ;
        RECT  11.8025 28.77 11.8675 28.905 ;
        RECT  11.0625 29.6225 11.1975 29.6875 ;
        RECT  11.4225 28.28 11.5225 28.3425 ;
        RECT  11.4225 28.2775 11.5225 28.34 ;
        RECT  11.75 29.4825 11.8025 29.545 ;
        RECT  11.4225 28.28 11.5225 28.3425 ;
        RECT  11.8 28.3425 11.87 28.5425 ;
        RECT  11.8 28.8725 11.87 29.0075 ;
        RECT  11.8 28.8725 11.87 29.0075 ;
        RECT  11.04 29.6225 11.925 29.6875 ;
        RECT  11.615 29.1075 11.79 29.1725 ;
        RECT  11.095 28.8725 11.165 29.0075 ;
        RECT  11.285 28.4325 11.35 29.1725 ;
        RECT  11.4225 28.2775 11.5225 28.34 ;
        RECT  11.045 29.4825 11.0975 29.545 ;
        RECT  11.8 28.8725 11.87 29.0075 ;
        RECT  11.04 28.2775 11.925 28.3425 ;
        RECT  11.615 28.5425 11.68 29.1725 ;
        RECT  11.8 28.8725 11.87 29.0075 ;
        RECT  11.8 28.8725 11.87 29.0075 ;
        RECT  11.18 29.1075 11.25 29.3975 ;
        RECT  11.095 28.8725 11.165 29.0075 ;
        RECT  11.04 29.4825 11.925 29.5475 ;
        RECT  11.8 28.8725 11.87 29.0075 ;
        RECT  11.8 28.3425 11.87 28.5425 ;
        RECT  11.095 28.3425 11.165 28.5425 ;
        RECT  11.72 29.1075 11.79 29.3975 ;
        RECT  11.18 29.1075 11.35 29.1725 ;
        RECT  11.8 30.7675 11.865 30.9025 ;
        RECT  11.615 30.7675 11.68 30.9025 ;
        RECT  11.1 30.7675 11.165 30.9025 ;
        RECT  11.285 30.7675 11.35 30.9025 ;
        RECT  11.615 30.3025 11.68 30.4375 ;
        RECT  11.8 30.3025 11.865 30.4375 ;
        RECT  11.285 30.3025 11.35 30.4375 ;
        RECT  11.1 30.3025 11.165 30.4375 ;
        RECT  11.72 29.9125 11.785 30.0475 ;
        RECT  11.535 29.9125 11.6 30.0475 ;
        RECT  11.365 29.9125 11.43 30.0475 ;
        RECT  11.18 29.9125 11.245 30.0475 ;
        RECT  11.8025 30.405 11.8675 30.54 ;
        RECT  11.8025 30.405 11.8675 30.54 ;
        RECT  11.8025 30.405 11.8675 30.54 ;
        RECT  11.8025 30.405 11.8675 30.54 ;
        RECT  11.8025 30.405 11.8675 30.54 ;
        RECT  11.8025 30.405 11.8675 30.54 ;
        RECT  11.41 30.9675 11.545 31.0325 ;
        RECT  11.0625 29.6225 11.1975 29.6875 ;
        RECT  11.7675 29.6225 11.9025 29.6875 ;
        RECT  11.3975 29.7625 11.5325 29.8275 ;
        RECT  11.8025 30.405 11.8675 30.54 ;
        RECT  11.8025 30.405 11.8675 30.54 ;
        RECT  11.8025 30.405 11.8675 30.54 ;
        RECT  11.8025 30.405 11.8675 30.54 ;
        RECT  11.3025 30.6525 11.4375 30.7175 ;
        RECT  11.3025 30.6525 11.4375 30.7175 ;
        RECT  11.5275 30.5025 11.6625 30.5675 ;
        RECT  11.5275 30.5025 11.6625 30.5675 ;
        RECT  11.8025 30.405 11.8675 30.54 ;
        RECT  11.8025 30.405 11.8675 30.54 ;
        RECT  11.8025 30.405 11.8675 30.54 ;
        RECT  11.8025 30.405 11.8675 30.54 ;
        RECT  11.3525 29.9125 11.4175 30.0475 ;
        RECT  11.0975 30.405 11.1625 30.54 ;
        RECT  11.0975 30.405 11.1625 30.54 ;
        RECT  11.0975 30.405 11.1625 30.54 ;
        RECT  11.0975 30.405 11.1625 30.54 ;
        RECT  11.0975 30.405 11.1625 30.54 ;
        RECT  11.0975 30.405 11.1625 30.54 ;
        RECT  11.8025 30.405 11.8675 30.54 ;
        RECT  11.8025 30.405 11.8675 30.54 ;
        RECT  11.8025 30.405 11.8675 30.54 ;
        RECT  11.8025 30.405 11.8675 30.54 ;
        RECT  11.5475 29.9125 11.6125 30.0475 ;
        RECT  11.415 29.6225 11.55 29.6875 ;
        RECT  11.415 29.6225 11.55 29.6875 ;
        RECT  11.7675 29.6225 11.9025 29.6875 ;
        RECT  11.41 30.9675 11.545 31.0325 ;
        RECT  11.7675 29.6225 11.9025 29.6875 ;
        RECT  11.7675 29.6225 11.9025 29.6875 ;
        RECT  11.8025 30.405 11.8675 30.54 ;
        RECT  11.8025 30.405 11.8675 30.54 ;
        RECT  11.8025 30.405 11.8675 30.54 ;
        RECT  11.8025 30.405 11.8675 30.54 ;
        RECT  11.8025 30.405 11.8675 30.54 ;
        RECT  11.8025 30.405 11.8675 30.54 ;
        RECT  11.0625 29.6225 11.1975 29.6875 ;
        RECT  11.4225 30.9675 11.5225 31.03 ;
        RECT  11.4225 30.97 11.5225 31.0325 ;
        RECT  11.75 29.765 11.8025 29.8275 ;
        RECT  11.4225 30.9675 11.5225 31.03 ;
        RECT  11.8 30.7675 11.87 30.9675 ;
        RECT  11.8 30.3025 11.87 30.4375 ;
        RECT  11.8 30.3025 11.87 30.4375 ;
        RECT  11.04 29.6225 11.925 29.6875 ;
        RECT  11.615 30.1375 11.79 30.2025 ;
        RECT  11.095 30.3025 11.165 30.4375 ;
        RECT  11.285 30.1375 11.35 30.8775 ;
        RECT  11.4225 30.97 11.5225 31.0325 ;
        RECT  11.045 29.765 11.0975 29.8275 ;
        RECT  11.8 30.3025 11.87 30.4375 ;
        RECT  11.04 30.9675 11.925 31.0325 ;
        RECT  11.615 30.1375 11.68 30.7675 ;
        RECT  11.8 30.3025 11.87 30.4375 ;
        RECT  11.8 30.3025 11.87 30.4375 ;
        RECT  11.18 29.9125 11.25 30.2025 ;
        RECT  11.095 30.3025 11.165 30.4375 ;
        RECT  11.04 29.7625 11.925 29.8275 ;
        RECT  11.8 30.3025 11.87 30.4375 ;
        RECT  11.8 30.7675 11.87 30.9675 ;
        RECT  11.095 30.7675 11.165 30.9675 ;
        RECT  11.72 29.9125 11.79 30.2025 ;
        RECT  11.18 30.1375 11.35 30.2025 ;
        RECT  11.8 31.0975 11.865 31.2325 ;
        RECT  11.615 31.0975 11.68 31.2325 ;
        RECT  11.1 31.0975 11.165 31.2325 ;
        RECT  11.285 31.0975 11.35 31.2325 ;
        RECT  11.615 31.5625 11.68 31.6975 ;
        RECT  11.8 31.5625 11.865 31.6975 ;
        RECT  11.285 31.5625 11.35 31.6975 ;
        RECT  11.1 31.5625 11.165 31.6975 ;
        RECT  11.72 31.9525 11.785 32.0875 ;
        RECT  11.535 31.9525 11.6 32.0875 ;
        RECT  11.365 31.9525 11.43 32.0875 ;
        RECT  11.18 31.9525 11.245 32.0875 ;
        RECT  11.8025 31.46 11.8675 31.595 ;
        RECT  11.8025 31.46 11.8675 31.595 ;
        RECT  11.8025 31.46 11.8675 31.595 ;
        RECT  11.8025 31.46 11.8675 31.595 ;
        RECT  11.8025 31.46 11.8675 31.595 ;
        RECT  11.8025 31.46 11.8675 31.595 ;
        RECT  11.41 30.9675 11.545 31.0325 ;
        RECT  11.0625 32.3125 11.1975 32.3775 ;
        RECT  11.7675 32.3125 11.9025 32.3775 ;
        RECT  11.3975 32.1725 11.5325 32.2375 ;
        RECT  11.8025 31.46 11.8675 31.595 ;
        RECT  11.8025 31.46 11.8675 31.595 ;
        RECT  11.8025 31.46 11.8675 31.595 ;
        RECT  11.8025 31.46 11.8675 31.595 ;
        RECT  11.3025 31.2825 11.4375 31.3475 ;
        RECT  11.3025 31.2825 11.4375 31.3475 ;
        RECT  11.5275 31.4325 11.6625 31.4975 ;
        RECT  11.5275 31.4325 11.6625 31.4975 ;
        RECT  11.8025 31.46 11.8675 31.595 ;
        RECT  11.8025 31.46 11.8675 31.595 ;
        RECT  11.8025 31.46 11.8675 31.595 ;
        RECT  11.8025 31.46 11.8675 31.595 ;
        RECT  11.3525 31.9525 11.4175 32.0875 ;
        RECT  11.0975 31.46 11.1625 31.595 ;
        RECT  11.0975 31.46 11.1625 31.595 ;
        RECT  11.0975 31.46 11.1625 31.595 ;
        RECT  11.0975 31.46 11.1625 31.595 ;
        RECT  11.0975 31.46 11.1625 31.595 ;
        RECT  11.0975 31.46 11.1625 31.595 ;
        RECT  11.8025 31.46 11.8675 31.595 ;
        RECT  11.8025 31.46 11.8675 31.595 ;
        RECT  11.8025 31.46 11.8675 31.595 ;
        RECT  11.8025 31.46 11.8675 31.595 ;
        RECT  11.5475 31.9525 11.6125 32.0875 ;
        RECT  11.415 32.3125 11.55 32.3775 ;
        RECT  11.415 32.3125 11.55 32.3775 ;
        RECT  11.7675 32.3125 11.9025 32.3775 ;
        RECT  11.41 30.9675 11.545 31.0325 ;
        RECT  11.7675 32.3125 11.9025 32.3775 ;
        RECT  11.7675 32.3125 11.9025 32.3775 ;
        RECT  11.8025 31.46 11.8675 31.595 ;
        RECT  11.8025 31.46 11.8675 31.595 ;
        RECT  11.8025 31.46 11.8675 31.595 ;
        RECT  11.8025 31.46 11.8675 31.595 ;
        RECT  11.8025 31.46 11.8675 31.595 ;
        RECT  11.8025 31.46 11.8675 31.595 ;
        RECT  11.0625 32.3125 11.1975 32.3775 ;
        RECT  11.4225 30.97 11.5225 31.0325 ;
        RECT  11.4225 30.9675 11.5225 31.03 ;
        RECT  11.75 32.1725 11.8025 32.235 ;
        RECT  11.4225 30.97 11.5225 31.0325 ;
        RECT  11.8 31.0325 11.87 31.2325 ;
        RECT  11.8 31.5625 11.87 31.6975 ;
        RECT  11.8 31.5625 11.87 31.6975 ;
        RECT  11.04 32.3125 11.925 32.3775 ;
        RECT  11.615 31.7975 11.79 31.8625 ;
        RECT  11.095 31.5625 11.165 31.6975 ;
        RECT  11.285 31.1225 11.35 31.8625 ;
        RECT  11.4225 30.9675 11.5225 31.03 ;
        RECT  11.045 32.1725 11.0975 32.235 ;
        RECT  11.8 31.5625 11.87 31.6975 ;
        RECT  11.04 30.9675 11.925 31.0325 ;
        RECT  11.615 31.2325 11.68 31.8625 ;
        RECT  11.8 31.5625 11.87 31.6975 ;
        RECT  11.8 31.5625 11.87 31.6975 ;
        RECT  11.18 31.7975 11.25 32.0875 ;
        RECT  11.095 31.5625 11.165 31.6975 ;
        RECT  11.04 32.1725 11.925 32.2375 ;
        RECT  11.8 31.5625 11.87 31.6975 ;
        RECT  11.8 31.0325 11.87 31.2325 ;
        RECT  11.095 31.0325 11.165 31.2325 ;
        RECT  11.72 31.7975 11.79 32.0875 ;
        RECT  11.18 31.7975 11.35 31.8625 ;
        RECT  11.8 33.4575 11.865 33.5925 ;
        RECT  11.615 33.4575 11.68 33.5925 ;
        RECT  11.1 33.4575 11.165 33.5925 ;
        RECT  11.285 33.4575 11.35 33.5925 ;
        RECT  11.615 32.9925 11.68 33.1275 ;
        RECT  11.8 32.9925 11.865 33.1275 ;
        RECT  11.285 32.9925 11.35 33.1275 ;
        RECT  11.1 32.9925 11.165 33.1275 ;
        RECT  11.72 32.6025 11.785 32.7375 ;
        RECT  11.535 32.6025 11.6 32.7375 ;
        RECT  11.365 32.6025 11.43 32.7375 ;
        RECT  11.18 32.6025 11.245 32.7375 ;
        RECT  11.8025 33.095 11.8675 33.23 ;
        RECT  11.8025 33.095 11.8675 33.23 ;
        RECT  11.8025 33.095 11.8675 33.23 ;
        RECT  11.8025 33.095 11.8675 33.23 ;
        RECT  11.8025 33.095 11.8675 33.23 ;
        RECT  11.8025 33.095 11.8675 33.23 ;
        RECT  11.41 33.6575 11.545 33.7225 ;
        RECT  11.0625 32.3125 11.1975 32.3775 ;
        RECT  11.7675 32.3125 11.9025 32.3775 ;
        RECT  11.3975 32.4525 11.5325 32.5175 ;
        RECT  11.8025 33.095 11.8675 33.23 ;
        RECT  11.8025 33.095 11.8675 33.23 ;
        RECT  11.8025 33.095 11.8675 33.23 ;
        RECT  11.8025 33.095 11.8675 33.23 ;
        RECT  11.3025 33.3425 11.4375 33.4075 ;
        RECT  11.3025 33.3425 11.4375 33.4075 ;
        RECT  11.5275 33.1925 11.6625 33.2575 ;
        RECT  11.5275 33.1925 11.6625 33.2575 ;
        RECT  11.8025 33.095 11.8675 33.23 ;
        RECT  11.8025 33.095 11.8675 33.23 ;
        RECT  11.8025 33.095 11.8675 33.23 ;
        RECT  11.8025 33.095 11.8675 33.23 ;
        RECT  11.3525 32.6025 11.4175 32.7375 ;
        RECT  11.0975 33.095 11.1625 33.23 ;
        RECT  11.0975 33.095 11.1625 33.23 ;
        RECT  11.0975 33.095 11.1625 33.23 ;
        RECT  11.0975 33.095 11.1625 33.23 ;
        RECT  11.0975 33.095 11.1625 33.23 ;
        RECT  11.0975 33.095 11.1625 33.23 ;
        RECT  11.8025 33.095 11.8675 33.23 ;
        RECT  11.8025 33.095 11.8675 33.23 ;
        RECT  11.8025 33.095 11.8675 33.23 ;
        RECT  11.8025 33.095 11.8675 33.23 ;
        RECT  11.5475 32.6025 11.6125 32.7375 ;
        RECT  11.415 32.3125 11.55 32.3775 ;
        RECT  11.415 32.3125 11.55 32.3775 ;
        RECT  11.7675 32.3125 11.9025 32.3775 ;
        RECT  11.41 33.6575 11.545 33.7225 ;
        RECT  11.7675 32.3125 11.9025 32.3775 ;
        RECT  11.7675 32.3125 11.9025 32.3775 ;
        RECT  11.8025 33.095 11.8675 33.23 ;
        RECT  11.8025 33.095 11.8675 33.23 ;
        RECT  11.8025 33.095 11.8675 33.23 ;
        RECT  11.8025 33.095 11.8675 33.23 ;
        RECT  11.8025 33.095 11.8675 33.23 ;
        RECT  11.8025 33.095 11.8675 33.23 ;
        RECT  11.0625 32.3125 11.1975 32.3775 ;
        RECT  11.4225 33.6575 11.5225 33.72 ;
        RECT  11.4225 33.66 11.5225 33.7225 ;
        RECT  11.75 32.455 11.8025 32.5175 ;
        RECT  11.4225 33.6575 11.5225 33.72 ;
        RECT  11.8 33.4575 11.87 33.6575 ;
        RECT  11.8 32.9925 11.87 33.1275 ;
        RECT  11.8 32.9925 11.87 33.1275 ;
        RECT  11.04 32.3125 11.925 32.3775 ;
        RECT  11.615 32.8275 11.79 32.8925 ;
        RECT  11.095 32.9925 11.165 33.1275 ;
        RECT  11.285 32.8275 11.35 33.5675 ;
        RECT  11.4225 33.66 11.5225 33.7225 ;
        RECT  11.045 32.455 11.0975 32.5175 ;
        RECT  11.8 32.9925 11.87 33.1275 ;
        RECT  11.04 33.6575 11.925 33.7225 ;
        RECT  11.615 32.8275 11.68 33.4575 ;
        RECT  11.8 32.9925 11.87 33.1275 ;
        RECT  11.8 32.9925 11.87 33.1275 ;
        RECT  11.18 32.6025 11.25 32.8925 ;
        RECT  11.095 32.9925 11.165 33.1275 ;
        RECT  11.04 32.4525 11.925 32.5175 ;
        RECT  11.8 32.9925 11.87 33.1275 ;
        RECT  11.8 33.4575 11.87 33.6575 ;
        RECT  11.095 33.4575 11.165 33.6575 ;
        RECT  11.72 32.6025 11.79 32.8925 ;
        RECT  11.18 32.8275 11.35 32.8925 ;
        RECT  11.8 33.7875 11.865 33.9225 ;
        RECT  11.615 33.7875 11.68 33.9225 ;
        RECT  11.1 33.7875 11.165 33.9225 ;
        RECT  11.285 33.7875 11.35 33.9225 ;
        RECT  11.615 34.2525 11.68 34.3875 ;
        RECT  11.8 34.2525 11.865 34.3875 ;
        RECT  11.285 34.2525 11.35 34.3875 ;
        RECT  11.1 34.2525 11.165 34.3875 ;
        RECT  11.72 34.6425 11.785 34.7775 ;
        RECT  11.535 34.6425 11.6 34.7775 ;
        RECT  11.365 34.6425 11.43 34.7775 ;
        RECT  11.18 34.6425 11.245 34.7775 ;
        RECT  11.8025 34.15 11.8675 34.285 ;
        RECT  11.8025 34.15 11.8675 34.285 ;
        RECT  11.8025 34.15 11.8675 34.285 ;
        RECT  11.8025 34.15 11.8675 34.285 ;
        RECT  11.8025 34.15 11.8675 34.285 ;
        RECT  11.8025 34.15 11.8675 34.285 ;
        RECT  11.41 33.6575 11.545 33.7225 ;
        RECT  11.0625 35.0025 11.1975 35.0675 ;
        RECT  11.7675 35.0025 11.9025 35.0675 ;
        RECT  11.3975 34.8625 11.5325 34.9275 ;
        RECT  11.8025 34.15 11.8675 34.285 ;
        RECT  11.8025 34.15 11.8675 34.285 ;
        RECT  11.8025 34.15 11.8675 34.285 ;
        RECT  11.8025 34.15 11.8675 34.285 ;
        RECT  11.3025 33.9725 11.4375 34.0375 ;
        RECT  11.3025 33.9725 11.4375 34.0375 ;
        RECT  11.5275 34.1225 11.6625 34.1875 ;
        RECT  11.5275 34.1225 11.6625 34.1875 ;
        RECT  11.8025 34.15 11.8675 34.285 ;
        RECT  11.8025 34.15 11.8675 34.285 ;
        RECT  11.8025 34.15 11.8675 34.285 ;
        RECT  11.8025 34.15 11.8675 34.285 ;
        RECT  11.3525 34.6425 11.4175 34.7775 ;
        RECT  11.0975 34.15 11.1625 34.285 ;
        RECT  11.0975 34.15 11.1625 34.285 ;
        RECT  11.0975 34.15 11.1625 34.285 ;
        RECT  11.0975 34.15 11.1625 34.285 ;
        RECT  11.0975 34.15 11.1625 34.285 ;
        RECT  11.0975 34.15 11.1625 34.285 ;
        RECT  11.8025 34.15 11.8675 34.285 ;
        RECT  11.8025 34.15 11.8675 34.285 ;
        RECT  11.8025 34.15 11.8675 34.285 ;
        RECT  11.8025 34.15 11.8675 34.285 ;
        RECT  11.5475 34.6425 11.6125 34.7775 ;
        RECT  11.415 35.0025 11.55 35.0675 ;
        RECT  11.415 35.0025 11.55 35.0675 ;
        RECT  11.7675 35.0025 11.9025 35.0675 ;
        RECT  11.41 33.6575 11.545 33.7225 ;
        RECT  11.7675 35.0025 11.9025 35.0675 ;
        RECT  11.7675 35.0025 11.9025 35.0675 ;
        RECT  11.8025 34.15 11.8675 34.285 ;
        RECT  11.8025 34.15 11.8675 34.285 ;
        RECT  11.8025 34.15 11.8675 34.285 ;
        RECT  11.8025 34.15 11.8675 34.285 ;
        RECT  11.8025 34.15 11.8675 34.285 ;
        RECT  11.8025 34.15 11.8675 34.285 ;
        RECT  11.0625 35.0025 11.1975 35.0675 ;
        RECT  11.4225 33.66 11.5225 33.7225 ;
        RECT  11.4225 33.6575 11.5225 33.72 ;
        RECT  11.75 34.8625 11.8025 34.925 ;
        RECT  11.4225 33.66 11.5225 33.7225 ;
        RECT  11.8 33.7225 11.87 33.9225 ;
        RECT  11.8 34.2525 11.87 34.3875 ;
        RECT  11.8 34.2525 11.87 34.3875 ;
        RECT  11.04 35.0025 11.925 35.0675 ;
        RECT  11.615 34.4875 11.79 34.5525 ;
        RECT  11.095 34.2525 11.165 34.3875 ;
        RECT  11.285 33.8125 11.35 34.5525 ;
        RECT  11.4225 33.6575 11.5225 33.72 ;
        RECT  11.045 34.8625 11.0975 34.925 ;
        RECT  11.8 34.2525 11.87 34.3875 ;
        RECT  11.04 33.6575 11.925 33.7225 ;
        RECT  11.615 33.9225 11.68 34.5525 ;
        RECT  11.8 34.2525 11.87 34.3875 ;
        RECT  11.8 34.2525 11.87 34.3875 ;
        RECT  11.18 34.4875 11.25 34.7775 ;
        RECT  11.095 34.2525 11.165 34.3875 ;
        RECT  11.04 34.8625 11.925 34.9275 ;
        RECT  11.8 34.2525 11.87 34.3875 ;
        RECT  11.8 33.7225 11.87 33.9225 ;
        RECT  11.095 33.7225 11.165 33.9225 ;
        RECT  11.72 34.4875 11.79 34.7775 ;
        RECT  11.18 34.4875 11.35 34.5525 ;
        RECT  11.8 36.1475 11.865 36.2825 ;
        RECT  11.615 36.1475 11.68 36.2825 ;
        RECT  11.1 36.1475 11.165 36.2825 ;
        RECT  11.285 36.1475 11.35 36.2825 ;
        RECT  11.615 35.6825 11.68 35.8175 ;
        RECT  11.8 35.6825 11.865 35.8175 ;
        RECT  11.285 35.6825 11.35 35.8175 ;
        RECT  11.1 35.6825 11.165 35.8175 ;
        RECT  11.72 35.2925 11.785 35.4275 ;
        RECT  11.535 35.2925 11.6 35.4275 ;
        RECT  11.365 35.2925 11.43 35.4275 ;
        RECT  11.18 35.2925 11.245 35.4275 ;
        RECT  11.8025 35.785 11.8675 35.92 ;
        RECT  11.8025 35.785 11.8675 35.92 ;
        RECT  11.8025 35.785 11.8675 35.92 ;
        RECT  11.8025 35.785 11.8675 35.92 ;
        RECT  11.8025 35.785 11.8675 35.92 ;
        RECT  11.8025 35.785 11.8675 35.92 ;
        RECT  11.41 36.3475 11.545 36.4125 ;
        RECT  11.0625 35.0025 11.1975 35.0675 ;
        RECT  11.7675 35.0025 11.9025 35.0675 ;
        RECT  11.3975 35.1425 11.5325 35.2075 ;
        RECT  11.8025 35.785 11.8675 35.92 ;
        RECT  11.8025 35.785 11.8675 35.92 ;
        RECT  11.8025 35.785 11.8675 35.92 ;
        RECT  11.8025 35.785 11.8675 35.92 ;
        RECT  11.3025 36.0325 11.4375 36.0975 ;
        RECT  11.3025 36.0325 11.4375 36.0975 ;
        RECT  11.5275 35.8825 11.6625 35.9475 ;
        RECT  11.5275 35.8825 11.6625 35.9475 ;
        RECT  11.8025 35.785 11.8675 35.92 ;
        RECT  11.8025 35.785 11.8675 35.92 ;
        RECT  11.8025 35.785 11.8675 35.92 ;
        RECT  11.8025 35.785 11.8675 35.92 ;
        RECT  11.3525 35.2925 11.4175 35.4275 ;
        RECT  11.0975 35.785 11.1625 35.92 ;
        RECT  11.0975 35.785 11.1625 35.92 ;
        RECT  11.0975 35.785 11.1625 35.92 ;
        RECT  11.0975 35.785 11.1625 35.92 ;
        RECT  11.0975 35.785 11.1625 35.92 ;
        RECT  11.0975 35.785 11.1625 35.92 ;
        RECT  11.8025 35.785 11.8675 35.92 ;
        RECT  11.8025 35.785 11.8675 35.92 ;
        RECT  11.8025 35.785 11.8675 35.92 ;
        RECT  11.8025 35.785 11.8675 35.92 ;
        RECT  11.5475 35.2925 11.6125 35.4275 ;
        RECT  11.415 35.0025 11.55 35.0675 ;
        RECT  11.415 35.0025 11.55 35.0675 ;
        RECT  11.7675 35.0025 11.9025 35.0675 ;
        RECT  11.41 36.3475 11.545 36.4125 ;
        RECT  11.7675 35.0025 11.9025 35.0675 ;
        RECT  11.7675 35.0025 11.9025 35.0675 ;
        RECT  11.8025 35.785 11.8675 35.92 ;
        RECT  11.8025 35.785 11.8675 35.92 ;
        RECT  11.8025 35.785 11.8675 35.92 ;
        RECT  11.8025 35.785 11.8675 35.92 ;
        RECT  11.8025 35.785 11.8675 35.92 ;
        RECT  11.8025 35.785 11.8675 35.92 ;
        RECT  11.0625 35.0025 11.1975 35.0675 ;
        RECT  11.4225 36.3475 11.5225 36.41 ;
        RECT  11.4225 36.35 11.5225 36.4125 ;
        RECT  11.75 35.145 11.8025 35.2075 ;
        RECT  11.4225 36.3475 11.5225 36.41 ;
        RECT  11.8 36.1475 11.87 36.3475 ;
        RECT  11.8 35.6825 11.87 35.8175 ;
        RECT  11.8 35.6825 11.87 35.8175 ;
        RECT  11.04 35.0025 11.925 35.0675 ;
        RECT  11.615 35.5175 11.79 35.5825 ;
        RECT  11.095 35.6825 11.165 35.8175 ;
        RECT  11.285 35.5175 11.35 36.2575 ;
        RECT  11.4225 36.35 11.5225 36.4125 ;
        RECT  11.045 35.145 11.0975 35.2075 ;
        RECT  11.8 35.6825 11.87 35.8175 ;
        RECT  11.04 36.3475 11.925 36.4125 ;
        RECT  11.615 35.5175 11.68 36.1475 ;
        RECT  11.8 35.6825 11.87 35.8175 ;
        RECT  11.8 35.6825 11.87 35.8175 ;
        RECT  11.18 35.2925 11.25 35.5825 ;
        RECT  11.095 35.6825 11.165 35.8175 ;
        RECT  11.04 35.1425 11.925 35.2075 ;
        RECT  11.8 35.6825 11.87 35.8175 ;
        RECT  11.8 36.1475 11.87 36.3475 ;
        RECT  11.095 36.1475 11.165 36.3475 ;
        RECT  11.72 35.2925 11.79 35.5825 ;
        RECT  11.18 35.5175 11.35 35.5825 ;
        RECT  11.8 36.4775 11.865 36.6125 ;
        RECT  11.615 36.4775 11.68 36.6125 ;
        RECT  11.1 36.4775 11.165 36.6125 ;
        RECT  11.285 36.4775 11.35 36.6125 ;
        RECT  11.615 36.9425 11.68 37.0775 ;
        RECT  11.8 36.9425 11.865 37.0775 ;
        RECT  11.285 36.9425 11.35 37.0775 ;
        RECT  11.1 36.9425 11.165 37.0775 ;
        RECT  11.72 37.3325 11.785 37.4675 ;
        RECT  11.535 37.3325 11.6 37.4675 ;
        RECT  11.365 37.3325 11.43 37.4675 ;
        RECT  11.18 37.3325 11.245 37.4675 ;
        RECT  11.8025 36.84 11.8675 36.975 ;
        RECT  11.8025 36.84 11.8675 36.975 ;
        RECT  11.8025 36.84 11.8675 36.975 ;
        RECT  11.8025 36.84 11.8675 36.975 ;
        RECT  11.8025 36.84 11.8675 36.975 ;
        RECT  11.8025 36.84 11.8675 36.975 ;
        RECT  11.41 36.3475 11.545 36.4125 ;
        RECT  11.0625 37.6925 11.1975 37.7575 ;
        RECT  11.7675 37.6925 11.9025 37.7575 ;
        RECT  11.3975 37.5525 11.5325 37.6175 ;
        RECT  11.8025 36.84 11.8675 36.975 ;
        RECT  11.8025 36.84 11.8675 36.975 ;
        RECT  11.8025 36.84 11.8675 36.975 ;
        RECT  11.8025 36.84 11.8675 36.975 ;
        RECT  11.3025 36.6625 11.4375 36.7275 ;
        RECT  11.3025 36.6625 11.4375 36.7275 ;
        RECT  11.5275 36.8125 11.6625 36.8775 ;
        RECT  11.5275 36.8125 11.6625 36.8775 ;
        RECT  11.8025 36.84 11.8675 36.975 ;
        RECT  11.8025 36.84 11.8675 36.975 ;
        RECT  11.8025 36.84 11.8675 36.975 ;
        RECT  11.8025 36.84 11.8675 36.975 ;
        RECT  11.3525 37.3325 11.4175 37.4675 ;
        RECT  11.0975 36.84 11.1625 36.975 ;
        RECT  11.0975 36.84 11.1625 36.975 ;
        RECT  11.0975 36.84 11.1625 36.975 ;
        RECT  11.0975 36.84 11.1625 36.975 ;
        RECT  11.0975 36.84 11.1625 36.975 ;
        RECT  11.0975 36.84 11.1625 36.975 ;
        RECT  11.8025 36.84 11.8675 36.975 ;
        RECT  11.8025 36.84 11.8675 36.975 ;
        RECT  11.8025 36.84 11.8675 36.975 ;
        RECT  11.8025 36.84 11.8675 36.975 ;
        RECT  11.5475 37.3325 11.6125 37.4675 ;
        RECT  11.415 37.6925 11.55 37.7575 ;
        RECT  11.415 37.6925 11.55 37.7575 ;
        RECT  11.7675 37.6925 11.9025 37.7575 ;
        RECT  11.41 36.3475 11.545 36.4125 ;
        RECT  11.7675 37.6925 11.9025 37.7575 ;
        RECT  11.7675 37.6925 11.9025 37.7575 ;
        RECT  11.8025 36.84 11.8675 36.975 ;
        RECT  11.8025 36.84 11.8675 36.975 ;
        RECT  11.8025 36.84 11.8675 36.975 ;
        RECT  11.8025 36.84 11.8675 36.975 ;
        RECT  11.8025 36.84 11.8675 36.975 ;
        RECT  11.8025 36.84 11.8675 36.975 ;
        RECT  11.0625 37.6925 11.1975 37.7575 ;
        RECT  11.4225 36.35 11.5225 36.4125 ;
        RECT  11.4225 36.3475 11.5225 36.41 ;
        RECT  11.75 37.5525 11.8025 37.615 ;
        RECT  11.4225 36.35 11.5225 36.4125 ;
        RECT  11.8 36.4125 11.87 36.6125 ;
        RECT  11.8 36.9425 11.87 37.0775 ;
        RECT  11.8 36.9425 11.87 37.0775 ;
        RECT  11.04 37.6925 11.925 37.7575 ;
        RECT  11.615 37.1775 11.79 37.2425 ;
        RECT  11.095 36.9425 11.165 37.0775 ;
        RECT  11.285 36.5025 11.35 37.2425 ;
        RECT  11.4225 36.3475 11.5225 36.41 ;
        RECT  11.045 37.5525 11.0975 37.615 ;
        RECT  11.8 36.9425 11.87 37.0775 ;
        RECT  11.04 36.3475 11.925 36.4125 ;
        RECT  11.615 36.6125 11.68 37.2425 ;
        RECT  11.8 36.9425 11.87 37.0775 ;
        RECT  11.8 36.9425 11.87 37.0775 ;
        RECT  11.18 37.1775 11.25 37.4675 ;
        RECT  11.095 36.9425 11.165 37.0775 ;
        RECT  11.04 37.5525 11.925 37.6175 ;
        RECT  11.8 36.9425 11.87 37.0775 ;
        RECT  11.8 36.4125 11.87 36.6125 ;
        RECT  11.095 36.4125 11.165 36.6125 ;
        RECT  11.72 37.1775 11.79 37.4675 ;
        RECT  11.18 37.1775 11.35 37.2425 ;
        RECT  11.8 38.8375 11.865 38.9725 ;
        RECT  11.615 38.8375 11.68 38.9725 ;
        RECT  11.1 38.8375 11.165 38.9725 ;
        RECT  11.285 38.8375 11.35 38.9725 ;
        RECT  11.615 38.3725 11.68 38.5075 ;
        RECT  11.8 38.3725 11.865 38.5075 ;
        RECT  11.285 38.3725 11.35 38.5075 ;
        RECT  11.1 38.3725 11.165 38.5075 ;
        RECT  11.72 37.9825 11.785 38.1175 ;
        RECT  11.535 37.9825 11.6 38.1175 ;
        RECT  11.365 37.9825 11.43 38.1175 ;
        RECT  11.18 37.9825 11.245 38.1175 ;
        RECT  11.8025 38.475 11.8675 38.61 ;
        RECT  11.8025 38.475 11.8675 38.61 ;
        RECT  11.8025 38.475 11.8675 38.61 ;
        RECT  11.8025 38.475 11.8675 38.61 ;
        RECT  11.8025 38.475 11.8675 38.61 ;
        RECT  11.8025 38.475 11.8675 38.61 ;
        RECT  11.41 39.0375 11.545 39.1025 ;
        RECT  11.0625 37.6925 11.1975 37.7575 ;
        RECT  11.7675 37.6925 11.9025 37.7575 ;
        RECT  11.3975 37.8325 11.5325 37.8975 ;
        RECT  11.8025 38.475 11.8675 38.61 ;
        RECT  11.8025 38.475 11.8675 38.61 ;
        RECT  11.8025 38.475 11.8675 38.61 ;
        RECT  11.8025 38.475 11.8675 38.61 ;
        RECT  11.3025 38.7225 11.4375 38.7875 ;
        RECT  11.3025 38.7225 11.4375 38.7875 ;
        RECT  11.5275 38.5725 11.6625 38.6375 ;
        RECT  11.5275 38.5725 11.6625 38.6375 ;
        RECT  11.8025 38.475 11.8675 38.61 ;
        RECT  11.8025 38.475 11.8675 38.61 ;
        RECT  11.8025 38.475 11.8675 38.61 ;
        RECT  11.8025 38.475 11.8675 38.61 ;
        RECT  11.3525 37.9825 11.4175 38.1175 ;
        RECT  11.0975 38.475 11.1625 38.61 ;
        RECT  11.0975 38.475 11.1625 38.61 ;
        RECT  11.0975 38.475 11.1625 38.61 ;
        RECT  11.0975 38.475 11.1625 38.61 ;
        RECT  11.0975 38.475 11.1625 38.61 ;
        RECT  11.0975 38.475 11.1625 38.61 ;
        RECT  11.8025 38.475 11.8675 38.61 ;
        RECT  11.8025 38.475 11.8675 38.61 ;
        RECT  11.8025 38.475 11.8675 38.61 ;
        RECT  11.8025 38.475 11.8675 38.61 ;
        RECT  11.5475 37.9825 11.6125 38.1175 ;
        RECT  11.415 37.6925 11.55 37.7575 ;
        RECT  11.415 37.6925 11.55 37.7575 ;
        RECT  11.7675 37.6925 11.9025 37.7575 ;
        RECT  11.41 39.0375 11.545 39.1025 ;
        RECT  11.7675 37.6925 11.9025 37.7575 ;
        RECT  11.7675 37.6925 11.9025 37.7575 ;
        RECT  11.8025 38.475 11.8675 38.61 ;
        RECT  11.8025 38.475 11.8675 38.61 ;
        RECT  11.8025 38.475 11.8675 38.61 ;
        RECT  11.8025 38.475 11.8675 38.61 ;
        RECT  11.8025 38.475 11.8675 38.61 ;
        RECT  11.8025 38.475 11.8675 38.61 ;
        RECT  11.0625 37.6925 11.1975 37.7575 ;
        RECT  11.4225 39.0375 11.5225 39.1 ;
        RECT  11.4225 39.04 11.5225 39.1025 ;
        RECT  11.75 37.835 11.8025 37.8975 ;
        RECT  11.4225 39.0375 11.5225 39.1 ;
        RECT  11.8 38.8375 11.87 39.0375 ;
        RECT  11.8 38.3725 11.87 38.5075 ;
        RECT  11.8 38.3725 11.87 38.5075 ;
        RECT  11.04 37.6925 11.925 37.7575 ;
        RECT  11.615 38.2075 11.79 38.2725 ;
        RECT  11.095 38.3725 11.165 38.5075 ;
        RECT  11.285 38.2075 11.35 38.9475 ;
        RECT  11.4225 39.04 11.5225 39.1025 ;
        RECT  11.045 37.835 11.0975 37.8975 ;
        RECT  11.8 38.3725 11.87 38.5075 ;
        RECT  11.04 39.0375 11.925 39.1025 ;
        RECT  11.615 38.2075 11.68 38.8375 ;
        RECT  11.8 38.3725 11.87 38.5075 ;
        RECT  11.8 38.3725 11.87 38.5075 ;
        RECT  11.18 37.9825 11.25 38.2725 ;
        RECT  11.095 38.3725 11.165 38.5075 ;
        RECT  11.04 37.8325 11.925 37.8975 ;
        RECT  11.8 38.3725 11.87 38.5075 ;
        RECT  11.8 38.8375 11.87 39.0375 ;
        RECT  11.095 38.8375 11.165 39.0375 ;
        RECT  11.72 37.9825 11.79 38.2725 ;
        RECT  11.18 38.2075 11.35 38.2725 ;
        RECT  11.8 39.1675 11.865 39.3025 ;
        RECT  11.615 39.1675 11.68 39.3025 ;
        RECT  11.1 39.1675 11.165 39.3025 ;
        RECT  11.285 39.1675 11.35 39.3025 ;
        RECT  11.615 39.6325 11.68 39.7675 ;
        RECT  11.8 39.6325 11.865 39.7675 ;
        RECT  11.285 39.6325 11.35 39.7675 ;
        RECT  11.1 39.6325 11.165 39.7675 ;
        RECT  11.72 40.0225 11.785 40.1575 ;
        RECT  11.535 40.0225 11.6 40.1575 ;
        RECT  11.365 40.0225 11.43 40.1575 ;
        RECT  11.18 40.0225 11.245 40.1575 ;
        RECT  11.8025 39.53 11.8675 39.665 ;
        RECT  11.8025 39.53 11.8675 39.665 ;
        RECT  11.8025 39.53 11.8675 39.665 ;
        RECT  11.8025 39.53 11.8675 39.665 ;
        RECT  11.8025 39.53 11.8675 39.665 ;
        RECT  11.8025 39.53 11.8675 39.665 ;
        RECT  11.41 39.0375 11.545 39.1025 ;
        RECT  11.0625 40.3825 11.1975 40.4475 ;
        RECT  11.7675 40.3825 11.9025 40.4475 ;
        RECT  11.3975 40.2425 11.5325 40.3075 ;
        RECT  11.8025 39.53 11.8675 39.665 ;
        RECT  11.8025 39.53 11.8675 39.665 ;
        RECT  11.8025 39.53 11.8675 39.665 ;
        RECT  11.8025 39.53 11.8675 39.665 ;
        RECT  11.3025 39.3525 11.4375 39.4175 ;
        RECT  11.3025 39.3525 11.4375 39.4175 ;
        RECT  11.5275 39.5025 11.6625 39.5675 ;
        RECT  11.5275 39.5025 11.6625 39.5675 ;
        RECT  11.8025 39.53 11.8675 39.665 ;
        RECT  11.8025 39.53 11.8675 39.665 ;
        RECT  11.8025 39.53 11.8675 39.665 ;
        RECT  11.8025 39.53 11.8675 39.665 ;
        RECT  11.3525 40.0225 11.4175 40.1575 ;
        RECT  11.0975 39.53 11.1625 39.665 ;
        RECT  11.0975 39.53 11.1625 39.665 ;
        RECT  11.0975 39.53 11.1625 39.665 ;
        RECT  11.0975 39.53 11.1625 39.665 ;
        RECT  11.0975 39.53 11.1625 39.665 ;
        RECT  11.0975 39.53 11.1625 39.665 ;
        RECT  11.8025 39.53 11.8675 39.665 ;
        RECT  11.8025 39.53 11.8675 39.665 ;
        RECT  11.8025 39.53 11.8675 39.665 ;
        RECT  11.8025 39.53 11.8675 39.665 ;
        RECT  11.5475 40.0225 11.6125 40.1575 ;
        RECT  11.415 40.3825 11.55 40.4475 ;
        RECT  11.415 40.3825 11.55 40.4475 ;
        RECT  11.7675 40.3825 11.9025 40.4475 ;
        RECT  11.41 39.0375 11.545 39.1025 ;
        RECT  11.7675 40.3825 11.9025 40.4475 ;
        RECT  11.7675 40.3825 11.9025 40.4475 ;
        RECT  11.8025 39.53 11.8675 39.665 ;
        RECT  11.8025 39.53 11.8675 39.665 ;
        RECT  11.8025 39.53 11.8675 39.665 ;
        RECT  11.8025 39.53 11.8675 39.665 ;
        RECT  11.8025 39.53 11.8675 39.665 ;
        RECT  11.8025 39.53 11.8675 39.665 ;
        RECT  11.0625 40.3825 11.1975 40.4475 ;
        RECT  11.4225 39.04 11.5225 39.1025 ;
        RECT  11.4225 39.0375 11.5225 39.1 ;
        RECT  11.75 40.2425 11.8025 40.305 ;
        RECT  11.4225 39.04 11.5225 39.1025 ;
        RECT  11.8 39.1025 11.87 39.3025 ;
        RECT  11.8 39.6325 11.87 39.7675 ;
        RECT  11.8 39.6325 11.87 39.7675 ;
        RECT  11.04 40.3825 11.925 40.4475 ;
        RECT  11.615 39.8675 11.79 39.9325 ;
        RECT  11.095 39.6325 11.165 39.7675 ;
        RECT  11.285 39.1925 11.35 39.9325 ;
        RECT  11.4225 39.0375 11.5225 39.1 ;
        RECT  11.045 40.2425 11.0975 40.305 ;
        RECT  11.8 39.6325 11.87 39.7675 ;
        RECT  11.04 39.0375 11.925 39.1025 ;
        RECT  11.615 39.3025 11.68 39.9325 ;
        RECT  11.8 39.6325 11.87 39.7675 ;
        RECT  11.8 39.6325 11.87 39.7675 ;
        RECT  11.18 39.8675 11.25 40.1575 ;
        RECT  11.095 39.6325 11.165 39.7675 ;
        RECT  11.04 40.2425 11.925 40.3075 ;
        RECT  11.8 39.6325 11.87 39.7675 ;
        RECT  11.8 39.1025 11.87 39.3025 ;
        RECT  11.095 39.1025 11.165 39.3025 ;
        RECT  11.72 39.8675 11.79 40.1575 ;
        RECT  11.18 39.8675 11.35 39.9325 ;
        RECT  12.505 20.0075 12.57 20.1425 ;
        RECT  12.32 20.0075 12.385 20.1425 ;
        RECT  11.805 20.0075 11.87 20.1425 ;
        RECT  11.99 20.0075 12.055 20.1425 ;
        RECT  12.32 19.5425 12.385 19.6775 ;
        RECT  12.505 19.5425 12.57 19.6775 ;
        RECT  11.99 19.5425 12.055 19.6775 ;
        RECT  11.805 19.5425 11.87 19.6775 ;
        RECT  12.425 19.1525 12.49 19.2875 ;
        RECT  12.24 19.1525 12.305 19.2875 ;
        RECT  12.07 19.1525 12.135 19.2875 ;
        RECT  11.885 19.1525 11.95 19.2875 ;
        RECT  12.5075 19.645 12.5725 19.78 ;
        RECT  12.5075 19.645 12.5725 19.78 ;
        RECT  12.5075 19.645 12.5725 19.78 ;
        RECT  12.5075 19.645 12.5725 19.78 ;
        RECT  12.5075 19.645 12.5725 19.78 ;
        RECT  12.5075 19.645 12.5725 19.78 ;
        RECT  12.115 20.2075 12.25 20.2725 ;
        RECT  11.7675 18.8625 11.9025 18.9275 ;
        RECT  12.4725 18.8625 12.6075 18.9275 ;
        RECT  12.1025 19.0025 12.2375 19.0675 ;
        RECT  12.5075 19.645 12.5725 19.78 ;
        RECT  12.5075 19.645 12.5725 19.78 ;
        RECT  12.5075 19.645 12.5725 19.78 ;
        RECT  12.5075 19.645 12.5725 19.78 ;
        RECT  12.0075 19.8925 12.1425 19.9575 ;
        RECT  12.0075 19.8925 12.1425 19.9575 ;
        RECT  12.2325 19.7425 12.3675 19.8075 ;
        RECT  12.2325 19.7425 12.3675 19.8075 ;
        RECT  12.5075 19.645 12.5725 19.78 ;
        RECT  12.5075 19.645 12.5725 19.78 ;
        RECT  12.5075 19.645 12.5725 19.78 ;
        RECT  12.5075 19.645 12.5725 19.78 ;
        RECT  12.0575 19.1525 12.1225 19.2875 ;
        RECT  11.8025 19.645 11.8675 19.78 ;
        RECT  11.8025 19.645 11.8675 19.78 ;
        RECT  11.8025 19.645 11.8675 19.78 ;
        RECT  11.8025 19.645 11.8675 19.78 ;
        RECT  11.8025 19.645 11.8675 19.78 ;
        RECT  11.8025 19.645 11.8675 19.78 ;
        RECT  12.5075 19.645 12.5725 19.78 ;
        RECT  12.5075 19.645 12.5725 19.78 ;
        RECT  12.5075 19.645 12.5725 19.78 ;
        RECT  12.5075 19.645 12.5725 19.78 ;
        RECT  12.2525 19.1525 12.3175 19.2875 ;
        RECT  12.12 18.8625 12.255 18.9275 ;
        RECT  12.12 18.8625 12.255 18.9275 ;
        RECT  12.4725 18.8625 12.6075 18.9275 ;
        RECT  12.115 20.2075 12.25 20.2725 ;
        RECT  12.4725 18.8625 12.6075 18.9275 ;
        RECT  12.4725 18.8625 12.6075 18.9275 ;
        RECT  12.5075 19.645 12.5725 19.78 ;
        RECT  12.5075 19.645 12.5725 19.78 ;
        RECT  12.5075 19.645 12.5725 19.78 ;
        RECT  12.5075 19.645 12.5725 19.78 ;
        RECT  12.5075 19.645 12.5725 19.78 ;
        RECT  12.5075 19.645 12.5725 19.78 ;
        RECT  11.7675 18.8625 11.9025 18.9275 ;
        RECT  12.1275 20.2075 12.2275 20.27 ;
        RECT  12.1275 20.21 12.2275 20.2725 ;
        RECT  12.455 19.005 12.5075 19.0675 ;
        RECT  12.1275 20.2075 12.2275 20.27 ;
        RECT  12.505 20.0075 12.575 20.2075 ;
        RECT  12.505 19.5425 12.575 19.6775 ;
        RECT  12.505 19.5425 12.575 19.6775 ;
        RECT  11.745 18.8625 12.63 18.9275 ;
        RECT  12.32 19.3775 12.495 19.4425 ;
        RECT  11.8 19.5425 11.87 19.6775 ;
        RECT  11.99 19.3775 12.055 20.1175 ;
        RECT  12.1275 20.21 12.2275 20.2725 ;
        RECT  11.75 19.005 11.8025 19.0675 ;
        RECT  12.505 19.5425 12.575 19.6775 ;
        RECT  11.745 20.2075 12.63 20.2725 ;
        RECT  12.32 19.3775 12.385 20.0075 ;
        RECT  12.505 19.5425 12.575 19.6775 ;
        RECT  12.505 19.5425 12.575 19.6775 ;
        RECT  11.885 19.1525 11.955 19.4425 ;
        RECT  11.8 19.5425 11.87 19.6775 ;
        RECT  11.745 19.0025 12.63 19.0675 ;
        RECT  12.505 19.5425 12.575 19.6775 ;
        RECT  12.505 20.0075 12.575 20.2075 ;
        RECT  11.8 20.0075 11.87 20.2075 ;
        RECT  12.425 19.1525 12.495 19.4425 ;
        RECT  11.885 19.3775 12.055 19.4425 ;
        RECT  12.505 20.3375 12.57 20.4725 ;
        RECT  12.32 20.3375 12.385 20.4725 ;
        RECT  11.805 20.3375 11.87 20.4725 ;
        RECT  11.99 20.3375 12.055 20.4725 ;
        RECT  12.32 20.8025 12.385 20.9375 ;
        RECT  12.505 20.8025 12.57 20.9375 ;
        RECT  11.99 20.8025 12.055 20.9375 ;
        RECT  11.805 20.8025 11.87 20.9375 ;
        RECT  12.425 21.1925 12.49 21.3275 ;
        RECT  12.24 21.1925 12.305 21.3275 ;
        RECT  12.07 21.1925 12.135 21.3275 ;
        RECT  11.885 21.1925 11.95 21.3275 ;
        RECT  12.5075 20.7 12.5725 20.835 ;
        RECT  12.5075 20.7 12.5725 20.835 ;
        RECT  12.5075 20.7 12.5725 20.835 ;
        RECT  12.5075 20.7 12.5725 20.835 ;
        RECT  12.5075 20.7 12.5725 20.835 ;
        RECT  12.5075 20.7 12.5725 20.835 ;
        RECT  12.115 20.2075 12.25 20.2725 ;
        RECT  11.7675 21.5525 11.9025 21.6175 ;
        RECT  12.4725 21.5525 12.6075 21.6175 ;
        RECT  12.1025 21.4125 12.2375 21.4775 ;
        RECT  12.5075 20.7 12.5725 20.835 ;
        RECT  12.5075 20.7 12.5725 20.835 ;
        RECT  12.5075 20.7 12.5725 20.835 ;
        RECT  12.5075 20.7 12.5725 20.835 ;
        RECT  12.0075 20.5225 12.1425 20.5875 ;
        RECT  12.0075 20.5225 12.1425 20.5875 ;
        RECT  12.2325 20.6725 12.3675 20.7375 ;
        RECT  12.2325 20.6725 12.3675 20.7375 ;
        RECT  12.5075 20.7 12.5725 20.835 ;
        RECT  12.5075 20.7 12.5725 20.835 ;
        RECT  12.5075 20.7 12.5725 20.835 ;
        RECT  12.5075 20.7 12.5725 20.835 ;
        RECT  12.0575 21.1925 12.1225 21.3275 ;
        RECT  11.8025 20.7 11.8675 20.835 ;
        RECT  11.8025 20.7 11.8675 20.835 ;
        RECT  11.8025 20.7 11.8675 20.835 ;
        RECT  11.8025 20.7 11.8675 20.835 ;
        RECT  11.8025 20.7 11.8675 20.835 ;
        RECT  11.8025 20.7 11.8675 20.835 ;
        RECT  12.5075 20.7 12.5725 20.835 ;
        RECT  12.5075 20.7 12.5725 20.835 ;
        RECT  12.5075 20.7 12.5725 20.835 ;
        RECT  12.5075 20.7 12.5725 20.835 ;
        RECT  12.2525 21.1925 12.3175 21.3275 ;
        RECT  12.12 21.5525 12.255 21.6175 ;
        RECT  12.12 21.5525 12.255 21.6175 ;
        RECT  12.4725 21.5525 12.6075 21.6175 ;
        RECT  12.115 20.2075 12.25 20.2725 ;
        RECT  12.4725 21.5525 12.6075 21.6175 ;
        RECT  12.4725 21.5525 12.6075 21.6175 ;
        RECT  12.5075 20.7 12.5725 20.835 ;
        RECT  12.5075 20.7 12.5725 20.835 ;
        RECT  12.5075 20.7 12.5725 20.835 ;
        RECT  12.5075 20.7 12.5725 20.835 ;
        RECT  12.5075 20.7 12.5725 20.835 ;
        RECT  12.5075 20.7 12.5725 20.835 ;
        RECT  11.7675 21.5525 11.9025 21.6175 ;
        RECT  12.1275 20.21 12.2275 20.2725 ;
        RECT  12.1275 20.2075 12.2275 20.27 ;
        RECT  12.455 21.4125 12.5075 21.475 ;
        RECT  12.1275 20.21 12.2275 20.2725 ;
        RECT  12.505 20.2725 12.575 20.4725 ;
        RECT  12.505 20.8025 12.575 20.9375 ;
        RECT  12.505 20.8025 12.575 20.9375 ;
        RECT  11.745 21.5525 12.63 21.6175 ;
        RECT  12.32 21.0375 12.495 21.1025 ;
        RECT  11.8 20.8025 11.87 20.9375 ;
        RECT  11.99 20.3625 12.055 21.1025 ;
        RECT  12.1275 20.2075 12.2275 20.27 ;
        RECT  11.75 21.4125 11.8025 21.475 ;
        RECT  12.505 20.8025 12.575 20.9375 ;
        RECT  11.745 20.2075 12.63 20.2725 ;
        RECT  12.32 20.4725 12.385 21.1025 ;
        RECT  12.505 20.8025 12.575 20.9375 ;
        RECT  12.505 20.8025 12.575 20.9375 ;
        RECT  11.885 21.0375 11.955 21.3275 ;
        RECT  11.8 20.8025 11.87 20.9375 ;
        RECT  11.745 21.4125 12.63 21.4775 ;
        RECT  12.505 20.8025 12.575 20.9375 ;
        RECT  12.505 20.2725 12.575 20.4725 ;
        RECT  11.8 20.2725 11.87 20.4725 ;
        RECT  12.425 21.0375 12.495 21.3275 ;
        RECT  11.885 21.0375 12.055 21.1025 ;
        RECT  12.505 22.6975 12.57 22.8325 ;
        RECT  12.32 22.6975 12.385 22.8325 ;
        RECT  11.805 22.6975 11.87 22.8325 ;
        RECT  11.99 22.6975 12.055 22.8325 ;
        RECT  12.32 22.2325 12.385 22.3675 ;
        RECT  12.505 22.2325 12.57 22.3675 ;
        RECT  11.99 22.2325 12.055 22.3675 ;
        RECT  11.805 22.2325 11.87 22.3675 ;
        RECT  12.425 21.8425 12.49 21.9775 ;
        RECT  12.24 21.8425 12.305 21.9775 ;
        RECT  12.07 21.8425 12.135 21.9775 ;
        RECT  11.885 21.8425 11.95 21.9775 ;
        RECT  12.5075 22.335 12.5725 22.47 ;
        RECT  12.5075 22.335 12.5725 22.47 ;
        RECT  12.5075 22.335 12.5725 22.47 ;
        RECT  12.5075 22.335 12.5725 22.47 ;
        RECT  12.5075 22.335 12.5725 22.47 ;
        RECT  12.5075 22.335 12.5725 22.47 ;
        RECT  12.115 22.8975 12.25 22.9625 ;
        RECT  11.7675 21.5525 11.9025 21.6175 ;
        RECT  12.4725 21.5525 12.6075 21.6175 ;
        RECT  12.1025 21.6925 12.2375 21.7575 ;
        RECT  12.5075 22.335 12.5725 22.47 ;
        RECT  12.5075 22.335 12.5725 22.47 ;
        RECT  12.5075 22.335 12.5725 22.47 ;
        RECT  12.5075 22.335 12.5725 22.47 ;
        RECT  12.0075 22.5825 12.1425 22.6475 ;
        RECT  12.0075 22.5825 12.1425 22.6475 ;
        RECT  12.2325 22.4325 12.3675 22.4975 ;
        RECT  12.2325 22.4325 12.3675 22.4975 ;
        RECT  12.5075 22.335 12.5725 22.47 ;
        RECT  12.5075 22.335 12.5725 22.47 ;
        RECT  12.5075 22.335 12.5725 22.47 ;
        RECT  12.5075 22.335 12.5725 22.47 ;
        RECT  12.0575 21.8425 12.1225 21.9775 ;
        RECT  11.8025 22.335 11.8675 22.47 ;
        RECT  11.8025 22.335 11.8675 22.47 ;
        RECT  11.8025 22.335 11.8675 22.47 ;
        RECT  11.8025 22.335 11.8675 22.47 ;
        RECT  11.8025 22.335 11.8675 22.47 ;
        RECT  11.8025 22.335 11.8675 22.47 ;
        RECT  12.5075 22.335 12.5725 22.47 ;
        RECT  12.5075 22.335 12.5725 22.47 ;
        RECT  12.5075 22.335 12.5725 22.47 ;
        RECT  12.5075 22.335 12.5725 22.47 ;
        RECT  12.2525 21.8425 12.3175 21.9775 ;
        RECT  12.12 21.5525 12.255 21.6175 ;
        RECT  12.12 21.5525 12.255 21.6175 ;
        RECT  12.4725 21.5525 12.6075 21.6175 ;
        RECT  12.115 22.8975 12.25 22.9625 ;
        RECT  12.4725 21.5525 12.6075 21.6175 ;
        RECT  12.4725 21.5525 12.6075 21.6175 ;
        RECT  12.5075 22.335 12.5725 22.47 ;
        RECT  12.5075 22.335 12.5725 22.47 ;
        RECT  12.5075 22.335 12.5725 22.47 ;
        RECT  12.5075 22.335 12.5725 22.47 ;
        RECT  12.5075 22.335 12.5725 22.47 ;
        RECT  12.5075 22.335 12.5725 22.47 ;
        RECT  11.7675 21.5525 11.9025 21.6175 ;
        RECT  12.1275 22.8975 12.2275 22.96 ;
        RECT  12.1275 22.9 12.2275 22.9625 ;
        RECT  12.455 21.695 12.5075 21.7575 ;
        RECT  12.1275 22.8975 12.2275 22.96 ;
        RECT  12.505 22.6975 12.575 22.8975 ;
        RECT  12.505 22.2325 12.575 22.3675 ;
        RECT  12.505 22.2325 12.575 22.3675 ;
        RECT  11.745 21.5525 12.63 21.6175 ;
        RECT  12.32 22.0675 12.495 22.1325 ;
        RECT  11.8 22.2325 11.87 22.3675 ;
        RECT  11.99 22.0675 12.055 22.8075 ;
        RECT  12.1275 22.9 12.2275 22.9625 ;
        RECT  11.75 21.695 11.8025 21.7575 ;
        RECT  12.505 22.2325 12.575 22.3675 ;
        RECT  11.745 22.8975 12.63 22.9625 ;
        RECT  12.32 22.0675 12.385 22.6975 ;
        RECT  12.505 22.2325 12.575 22.3675 ;
        RECT  12.505 22.2325 12.575 22.3675 ;
        RECT  11.885 21.8425 11.955 22.1325 ;
        RECT  11.8 22.2325 11.87 22.3675 ;
        RECT  11.745 21.6925 12.63 21.7575 ;
        RECT  12.505 22.2325 12.575 22.3675 ;
        RECT  12.505 22.6975 12.575 22.8975 ;
        RECT  11.8 22.6975 11.87 22.8975 ;
        RECT  12.425 21.8425 12.495 22.1325 ;
        RECT  11.885 22.0675 12.055 22.1325 ;
        RECT  12.505 23.0275 12.57 23.1625 ;
        RECT  12.32 23.0275 12.385 23.1625 ;
        RECT  11.805 23.0275 11.87 23.1625 ;
        RECT  11.99 23.0275 12.055 23.1625 ;
        RECT  12.32 23.4925 12.385 23.6275 ;
        RECT  12.505 23.4925 12.57 23.6275 ;
        RECT  11.99 23.4925 12.055 23.6275 ;
        RECT  11.805 23.4925 11.87 23.6275 ;
        RECT  12.425 23.8825 12.49 24.0175 ;
        RECT  12.24 23.8825 12.305 24.0175 ;
        RECT  12.07 23.8825 12.135 24.0175 ;
        RECT  11.885 23.8825 11.95 24.0175 ;
        RECT  12.5075 23.39 12.5725 23.525 ;
        RECT  12.5075 23.39 12.5725 23.525 ;
        RECT  12.5075 23.39 12.5725 23.525 ;
        RECT  12.5075 23.39 12.5725 23.525 ;
        RECT  12.5075 23.39 12.5725 23.525 ;
        RECT  12.5075 23.39 12.5725 23.525 ;
        RECT  12.115 22.8975 12.25 22.9625 ;
        RECT  11.7675 24.2425 11.9025 24.3075 ;
        RECT  12.4725 24.2425 12.6075 24.3075 ;
        RECT  12.1025 24.1025 12.2375 24.1675 ;
        RECT  12.5075 23.39 12.5725 23.525 ;
        RECT  12.5075 23.39 12.5725 23.525 ;
        RECT  12.5075 23.39 12.5725 23.525 ;
        RECT  12.5075 23.39 12.5725 23.525 ;
        RECT  12.0075 23.2125 12.1425 23.2775 ;
        RECT  12.0075 23.2125 12.1425 23.2775 ;
        RECT  12.2325 23.3625 12.3675 23.4275 ;
        RECT  12.2325 23.3625 12.3675 23.4275 ;
        RECT  12.5075 23.39 12.5725 23.525 ;
        RECT  12.5075 23.39 12.5725 23.525 ;
        RECT  12.5075 23.39 12.5725 23.525 ;
        RECT  12.5075 23.39 12.5725 23.525 ;
        RECT  12.0575 23.8825 12.1225 24.0175 ;
        RECT  11.8025 23.39 11.8675 23.525 ;
        RECT  11.8025 23.39 11.8675 23.525 ;
        RECT  11.8025 23.39 11.8675 23.525 ;
        RECT  11.8025 23.39 11.8675 23.525 ;
        RECT  11.8025 23.39 11.8675 23.525 ;
        RECT  11.8025 23.39 11.8675 23.525 ;
        RECT  12.5075 23.39 12.5725 23.525 ;
        RECT  12.5075 23.39 12.5725 23.525 ;
        RECT  12.5075 23.39 12.5725 23.525 ;
        RECT  12.5075 23.39 12.5725 23.525 ;
        RECT  12.2525 23.8825 12.3175 24.0175 ;
        RECT  12.12 24.2425 12.255 24.3075 ;
        RECT  12.12 24.2425 12.255 24.3075 ;
        RECT  12.4725 24.2425 12.6075 24.3075 ;
        RECT  12.115 22.8975 12.25 22.9625 ;
        RECT  12.4725 24.2425 12.6075 24.3075 ;
        RECT  12.4725 24.2425 12.6075 24.3075 ;
        RECT  12.5075 23.39 12.5725 23.525 ;
        RECT  12.5075 23.39 12.5725 23.525 ;
        RECT  12.5075 23.39 12.5725 23.525 ;
        RECT  12.5075 23.39 12.5725 23.525 ;
        RECT  12.5075 23.39 12.5725 23.525 ;
        RECT  12.5075 23.39 12.5725 23.525 ;
        RECT  11.7675 24.2425 11.9025 24.3075 ;
        RECT  12.1275 22.9 12.2275 22.9625 ;
        RECT  12.1275 22.8975 12.2275 22.96 ;
        RECT  12.455 24.1025 12.5075 24.165 ;
        RECT  12.1275 22.9 12.2275 22.9625 ;
        RECT  12.505 22.9625 12.575 23.1625 ;
        RECT  12.505 23.4925 12.575 23.6275 ;
        RECT  12.505 23.4925 12.575 23.6275 ;
        RECT  11.745 24.2425 12.63 24.3075 ;
        RECT  12.32 23.7275 12.495 23.7925 ;
        RECT  11.8 23.4925 11.87 23.6275 ;
        RECT  11.99 23.0525 12.055 23.7925 ;
        RECT  12.1275 22.8975 12.2275 22.96 ;
        RECT  11.75 24.1025 11.8025 24.165 ;
        RECT  12.505 23.4925 12.575 23.6275 ;
        RECT  11.745 22.8975 12.63 22.9625 ;
        RECT  12.32 23.1625 12.385 23.7925 ;
        RECT  12.505 23.4925 12.575 23.6275 ;
        RECT  12.505 23.4925 12.575 23.6275 ;
        RECT  11.885 23.7275 11.955 24.0175 ;
        RECT  11.8 23.4925 11.87 23.6275 ;
        RECT  11.745 24.1025 12.63 24.1675 ;
        RECT  12.505 23.4925 12.575 23.6275 ;
        RECT  12.505 22.9625 12.575 23.1625 ;
        RECT  11.8 22.9625 11.87 23.1625 ;
        RECT  12.425 23.7275 12.495 24.0175 ;
        RECT  11.885 23.7275 12.055 23.7925 ;
        RECT  12.505 25.3875 12.57 25.5225 ;
        RECT  12.32 25.3875 12.385 25.5225 ;
        RECT  11.805 25.3875 11.87 25.5225 ;
        RECT  11.99 25.3875 12.055 25.5225 ;
        RECT  12.32 24.9225 12.385 25.0575 ;
        RECT  12.505 24.9225 12.57 25.0575 ;
        RECT  11.99 24.9225 12.055 25.0575 ;
        RECT  11.805 24.9225 11.87 25.0575 ;
        RECT  12.425 24.5325 12.49 24.6675 ;
        RECT  12.24 24.5325 12.305 24.6675 ;
        RECT  12.07 24.5325 12.135 24.6675 ;
        RECT  11.885 24.5325 11.95 24.6675 ;
        RECT  12.5075 25.025 12.5725 25.16 ;
        RECT  12.5075 25.025 12.5725 25.16 ;
        RECT  12.5075 25.025 12.5725 25.16 ;
        RECT  12.5075 25.025 12.5725 25.16 ;
        RECT  12.5075 25.025 12.5725 25.16 ;
        RECT  12.5075 25.025 12.5725 25.16 ;
        RECT  12.115 25.5875 12.25 25.6525 ;
        RECT  11.7675 24.2425 11.9025 24.3075 ;
        RECT  12.4725 24.2425 12.6075 24.3075 ;
        RECT  12.1025 24.3825 12.2375 24.4475 ;
        RECT  12.5075 25.025 12.5725 25.16 ;
        RECT  12.5075 25.025 12.5725 25.16 ;
        RECT  12.5075 25.025 12.5725 25.16 ;
        RECT  12.5075 25.025 12.5725 25.16 ;
        RECT  12.0075 25.2725 12.1425 25.3375 ;
        RECT  12.0075 25.2725 12.1425 25.3375 ;
        RECT  12.2325 25.1225 12.3675 25.1875 ;
        RECT  12.2325 25.1225 12.3675 25.1875 ;
        RECT  12.5075 25.025 12.5725 25.16 ;
        RECT  12.5075 25.025 12.5725 25.16 ;
        RECT  12.5075 25.025 12.5725 25.16 ;
        RECT  12.5075 25.025 12.5725 25.16 ;
        RECT  12.0575 24.5325 12.1225 24.6675 ;
        RECT  11.8025 25.025 11.8675 25.16 ;
        RECT  11.8025 25.025 11.8675 25.16 ;
        RECT  11.8025 25.025 11.8675 25.16 ;
        RECT  11.8025 25.025 11.8675 25.16 ;
        RECT  11.8025 25.025 11.8675 25.16 ;
        RECT  11.8025 25.025 11.8675 25.16 ;
        RECT  12.5075 25.025 12.5725 25.16 ;
        RECT  12.5075 25.025 12.5725 25.16 ;
        RECT  12.5075 25.025 12.5725 25.16 ;
        RECT  12.5075 25.025 12.5725 25.16 ;
        RECT  12.2525 24.5325 12.3175 24.6675 ;
        RECT  12.12 24.2425 12.255 24.3075 ;
        RECT  12.12 24.2425 12.255 24.3075 ;
        RECT  12.4725 24.2425 12.6075 24.3075 ;
        RECT  12.115 25.5875 12.25 25.6525 ;
        RECT  12.4725 24.2425 12.6075 24.3075 ;
        RECT  12.4725 24.2425 12.6075 24.3075 ;
        RECT  12.5075 25.025 12.5725 25.16 ;
        RECT  12.5075 25.025 12.5725 25.16 ;
        RECT  12.5075 25.025 12.5725 25.16 ;
        RECT  12.5075 25.025 12.5725 25.16 ;
        RECT  12.5075 25.025 12.5725 25.16 ;
        RECT  12.5075 25.025 12.5725 25.16 ;
        RECT  11.7675 24.2425 11.9025 24.3075 ;
        RECT  12.1275 25.5875 12.2275 25.65 ;
        RECT  12.1275 25.59 12.2275 25.6525 ;
        RECT  12.455 24.385 12.5075 24.4475 ;
        RECT  12.1275 25.5875 12.2275 25.65 ;
        RECT  12.505 25.3875 12.575 25.5875 ;
        RECT  12.505 24.9225 12.575 25.0575 ;
        RECT  12.505 24.9225 12.575 25.0575 ;
        RECT  11.745 24.2425 12.63 24.3075 ;
        RECT  12.32 24.7575 12.495 24.8225 ;
        RECT  11.8 24.9225 11.87 25.0575 ;
        RECT  11.99 24.7575 12.055 25.4975 ;
        RECT  12.1275 25.59 12.2275 25.6525 ;
        RECT  11.75 24.385 11.8025 24.4475 ;
        RECT  12.505 24.9225 12.575 25.0575 ;
        RECT  11.745 25.5875 12.63 25.6525 ;
        RECT  12.32 24.7575 12.385 25.3875 ;
        RECT  12.505 24.9225 12.575 25.0575 ;
        RECT  12.505 24.9225 12.575 25.0575 ;
        RECT  11.885 24.5325 11.955 24.8225 ;
        RECT  11.8 24.9225 11.87 25.0575 ;
        RECT  11.745 24.3825 12.63 24.4475 ;
        RECT  12.505 24.9225 12.575 25.0575 ;
        RECT  12.505 25.3875 12.575 25.5875 ;
        RECT  11.8 25.3875 11.87 25.5875 ;
        RECT  12.425 24.5325 12.495 24.8225 ;
        RECT  11.885 24.7575 12.055 24.8225 ;
        RECT  12.505 25.7175 12.57 25.8525 ;
        RECT  12.32 25.7175 12.385 25.8525 ;
        RECT  11.805 25.7175 11.87 25.8525 ;
        RECT  11.99 25.7175 12.055 25.8525 ;
        RECT  12.32 26.1825 12.385 26.3175 ;
        RECT  12.505 26.1825 12.57 26.3175 ;
        RECT  11.99 26.1825 12.055 26.3175 ;
        RECT  11.805 26.1825 11.87 26.3175 ;
        RECT  12.425 26.5725 12.49 26.7075 ;
        RECT  12.24 26.5725 12.305 26.7075 ;
        RECT  12.07 26.5725 12.135 26.7075 ;
        RECT  11.885 26.5725 11.95 26.7075 ;
        RECT  12.5075 26.08 12.5725 26.215 ;
        RECT  12.5075 26.08 12.5725 26.215 ;
        RECT  12.5075 26.08 12.5725 26.215 ;
        RECT  12.5075 26.08 12.5725 26.215 ;
        RECT  12.5075 26.08 12.5725 26.215 ;
        RECT  12.5075 26.08 12.5725 26.215 ;
        RECT  12.115 25.5875 12.25 25.6525 ;
        RECT  11.7675 26.9325 11.9025 26.9975 ;
        RECT  12.4725 26.9325 12.6075 26.9975 ;
        RECT  12.1025 26.7925 12.2375 26.8575 ;
        RECT  12.5075 26.08 12.5725 26.215 ;
        RECT  12.5075 26.08 12.5725 26.215 ;
        RECT  12.5075 26.08 12.5725 26.215 ;
        RECT  12.5075 26.08 12.5725 26.215 ;
        RECT  12.0075 25.9025 12.1425 25.9675 ;
        RECT  12.0075 25.9025 12.1425 25.9675 ;
        RECT  12.2325 26.0525 12.3675 26.1175 ;
        RECT  12.2325 26.0525 12.3675 26.1175 ;
        RECT  12.5075 26.08 12.5725 26.215 ;
        RECT  12.5075 26.08 12.5725 26.215 ;
        RECT  12.5075 26.08 12.5725 26.215 ;
        RECT  12.5075 26.08 12.5725 26.215 ;
        RECT  12.0575 26.5725 12.1225 26.7075 ;
        RECT  11.8025 26.08 11.8675 26.215 ;
        RECT  11.8025 26.08 11.8675 26.215 ;
        RECT  11.8025 26.08 11.8675 26.215 ;
        RECT  11.8025 26.08 11.8675 26.215 ;
        RECT  11.8025 26.08 11.8675 26.215 ;
        RECT  11.8025 26.08 11.8675 26.215 ;
        RECT  12.5075 26.08 12.5725 26.215 ;
        RECT  12.5075 26.08 12.5725 26.215 ;
        RECT  12.5075 26.08 12.5725 26.215 ;
        RECT  12.5075 26.08 12.5725 26.215 ;
        RECT  12.2525 26.5725 12.3175 26.7075 ;
        RECT  12.12 26.9325 12.255 26.9975 ;
        RECT  12.12 26.9325 12.255 26.9975 ;
        RECT  12.4725 26.9325 12.6075 26.9975 ;
        RECT  12.115 25.5875 12.25 25.6525 ;
        RECT  12.4725 26.9325 12.6075 26.9975 ;
        RECT  12.4725 26.9325 12.6075 26.9975 ;
        RECT  12.5075 26.08 12.5725 26.215 ;
        RECT  12.5075 26.08 12.5725 26.215 ;
        RECT  12.5075 26.08 12.5725 26.215 ;
        RECT  12.5075 26.08 12.5725 26.215 ;
        RECT  12.5075 26.08 12.5725 26.215 ;
        RECT  12.5075 26.08 12.5725 26.215 ;
        RECT  11.7675 26.9325 11.9025 26.9975 ;
        RECT  12.1275 25.59 12.2275 25.6525 ;
        RECT  12.1275 25.5875 12.2275 25.65 ;
        RECT  12.455 26.7925 12.5075 26.855 ;
        RECT  12.1275 25.59 12.2275 25.6525 ;
        RECT  12.505 25.6525 12.575 25.8525 ;
        RECT  12.505 26.1825 12.575 26.3175 ;
        RECT  12.505 26.1825 12.575 26.3175 ;
        RECT  11.745 26.9325 12.63 26.9975 ;
        RECT  12.32 26.4175 12.495 26.4825 ;
        RECT  11.8 26.1825 11.87 26.3175 ;
        RECT  11.99 25.7425 12.055 26.4825 ;
        RECT  12.1275 25.5875 12.2275 25.65 ;
        RECT  11.75 26.7925 11.8025 26.855 ;
        RECT  12.505 26.1825 12.575 26.3175 ;
        RECT  11.745 25.5875 12.63 25.6525 ;
        RECT  12.32 25.8525 12.385 26.4825 ;
        RECT  12.505 26.1825 12.575 26.3175 ;
        RECT  12.505 26.1825 12.575 26.3175 ;
        RECT  11.885 26.4175 11.955 26.7075 ;
        RECT  11.8 26.1825 11.87 26.3175 ;
        RECT  11.745 26.7925 12.63 26.8575 ;
        RECT  12.505 26.1825 12.575 26.3175 ;
        RECT  12.505 25.6525 12.575 25.8525 ;
        RECT  11.8 25.6525 11.87 25.8525 ;
        RECT  12.425 26.4175 12.495 26.7075 ;
        RECT  11.885 26.4175 12.055 26.4825 ;
        RECT  12.505 28.0775 12.57 28.2125 ;
        RECT  12.32 28.0775 12.385 28.2125 ;
        RECT  11.805 28.0775 11.87 28.2125 ;
        RECT  11.99 28.0775 12.055 28.2125 ;
        RECT  12.32 27.6125 12.385 27.7475 ;
        RECT  12.505 27.6125 12.57 27.7475 ;
        RECT  11.99 27.6125 12.055 27.7475 ;
        RECT  11.805 27.6125 11.87 27.7475 ;
        RECT  12.425 27.2225 12.49 27.3575 ;
        RECT  12.24 27.2225 12.305 27.3575 ;
        RECT  12.07 27.2225 12.135 27.3575 ;
        RECT  11.885 27.2225 11.95 27.3575 ;
        RECT  12.5075 27.715 12.5725 27.85 ;
        RECT  12.5075 27.715 12.5725 27.85 ;
        RECT  12.5075 27.715 12.5725 27.85 ;
        RECT  12.5075 27.715 12.5725 27.85 ;
        RECT  12.5075 27.715 12.5725 27.85 ;
        RECT  12.5075 27.715 12.5725 27.85 ;
        RECT  12.115 28.2775 12.25 28.3425 ;
        RECT  11.7675 26.9325 11.9025 26.9975 ;
        RECT  12.4725 26.9325 12.6075 26.9975 ;
        RECT  12.1025 27.0725 12.2375 27.1375 ;
        RECT  12.5075 27.715 12.5725 27.85 ;
        RECT  12.5075 27.715 12.5725 27.85 ;
        RECT  12.5075 27.715 12.5725 27.85 ;
        RECT  12.5075 27.715 12.5725 27.85 ;
        RECT  12.0075 27.9625 12.1425 28.0275 ;
        RECT  12.0075 27.9625 12.1425 28.0275 ;
        RECT  12.2325 27.8125 12.3675 27.8775 ;
        RECT  12.2325 27.8125 12.3675 27.8775 ;
        RECT  12.5075 27.715 12.5725 27.85 ;
        RECT  12.5075 27.715 12.5725 27.85 ;
        RECT  12.5075 27.715 12.5725 27.85 ;
        RECT  12.5075 27.715 12.5725 27.85 ;
        RECT  12.0575 27.2225 12.1225 27.3575 ;
        RECT  11.8025 27.715 11.8675 27.85 ;
        RECT  11.8025 27.715 11.8675 27.85 ;
        RECT  11.8025 27.715 11.8675 27.85 ;
        RECT  11.8025 27.715 11.8675 27.85 ;
        RECT  11.8025 27.715 11.8675 27.85 ;
        RECT  11.8025 27.715 11.8675 27.85 ;
        RECT  12.5075 27.715 12.5725 27.85 ;
        RECT  12.5075 27.715 12.5725 27.85 ;
        RECT  12.5075 27.715 12.5725 27.85 ;
        RECT  12.5075 27.715 12.5725 27.85 ;
        RECT  12.2525 27.2225 12.3175 27.3575 ;
        RECT  12.12 26.9325 12.255 26.9975 ;
        RECT  12.12 26.9325 12.255 26.9975 ;
        RECT  12.4725 26.9325 12.6075 26.9975 ;
        RECT  12.115 28.2775 12.25 28.3425 ;
        RECT  12.4725 26.9325 12.6075 26.9975 ;
        RECT  12.4725 26.9325 12.6075 26.9975 ;
        RECT  12.5075 27.715 12.5725 27.85 ;
        RECT  12.5075 27.715 12.5725 27.85 ;
        RECT  12.5075 27.715 12.5725 27.85 ;
        RECT  12.5075 27.715 12.5725 27.85 ;
        RECT  12.5075 27.715 12.5725 27.85 ;
        RECT  12.5075 27.715 12.5725 27.85 ;
        RECT  11.7675 26.9325 11.9025 26.9975 ;
        RECT  12.1275 28.2775 12.2275 28.34 ;
        RECT  12.1275 28.28 12.2275 28.3425 ;
        RECT  12.455 27.075 12.5075 27.1375 ;
        RECT  12.1275 28.2775 12.2275 28.34 ;
        RECT  12.505 28.0775 12.575 28.2775 ;
        RECT  12.505 27.6125 12.575 27.7475 ;
        RECT  12.505 27.6125 12.575 27.7475 ;
        RECT  11.745 26.9325 12.63 26.9975 ;
        RECT  12.32 27.4475 12.495 27.5125 ;
        RECT  11.8 27.6125 11.87 27.7475 ;
        RECT  11.99 27.4475 12.055 28.1875 ;
        RECT  12.1275 28.28 12.2275 28.3425 ;
        RECT  11.75 27.075 11.8025 27.1375 ;
        RECT  12.505 27.6125 12.575 27.7475 ;
        RECT  11.745 28.2775 12.63 28.3425 ;
        RECT  12.32 27.4475 12.385 28.0775 ;
        RECT  12.505 27.6125 12.575 27.7475 ;
        RECT  12.505 27.6125 12.575 27.7475 ;
        RECT  11.885 27.2225 11.955 27.5125 ;
        RECT  11.8 27.6125 11.87 27.7475 ;
        RECT  11.745 27.0725 12.63 27.1375 ;
        RECT  12.505 27.6125 12.575 27.7475 ;
        RECT  12.505 28.0775 12.575 28.2775 ;
        RECT  11.8 28.0775 11.87 28.2775 ;
        RECT  12.425 27.2225 12.495 27.5125 ;
        RECT  11.885 27.4475 12.055 27.5125 ;
        RECT  12.505 28.4075 12.57 28.5425 ;
        RECT  12.32 28.4075 12.385 28.5425 ;
        RECT  11.805 28.4075 11.87 28.5425 ;
        RECT  11.99 28.4075 12.055 28.5425 ;
        RECT  12.32 28.8725 12.385 29.0075 ;
        RECT  12.505 28.8725 12.57 29.0075 ;
        RECT  11.99 28.8725 12.055 29.0075 ;
        RECT  11.805 28.8725 11.87 29.0075 ;
        RECT  12.425 29.2625 12.49 29.3975 ;
        RECT  12.24 29.2625 12.305 29.3975 ;
        RECT  12.07 29.2625 12.135 29.3975 ;
        RECT  11.885 29.2625 11.95 29.3975 ;
        RECT  12.5075 28.77 12.5725 28.905 ;
        RECT  12.5075 28.77 12.5725 28.905 ;
        RECT  12.5075 28.77 12.5725 28.905 ;
        RECT  12.5075 28.77 12.5725 28.905 ;
        RECT  12.5075 28.77 12.5725 28.905 ;
        RECT  12.5075 28.77 12.5725 28.905 ;
        RECT  12.115 28.2775 12.25 28.3425 ;
        RECT  11.7675 29.6225 11.9025 29.6875 ;
        RECT  12.4725 29.6225 12.6075 29.6875 ;
        RECT  12.1025 29.4825 12.2375 29.5475 ;
        RECT  12.5075 28.77 12.5725 28.905 ;
        RECT  12.5075 28.77 12.5725 28.905 ;
        RECT  12.5075 28.77 12.5725 28.905 ;
        RECT  12.5075 28.77 12.5725 28.905 ;
        RECT  12.0075 28.5925 12.1425 28.6575 ;
        RECT  12.0075 28.5925 12.1425 28.6575 ;
        RECT  12.2325 28.7425 12.3675 28.8075 ;
        RECT  12.2325 28.7425 12.3675 28.8075 ;
        RECT  12.5075 28.77 12.5725 28.905 ;
        RECT  12.5075 28.77 12.5725 28.905 ;
        RECT  12.5075 28.77 12.5725 28.905 ;
        RECT  12.5075 28.77 12.5725 28.905 ;
        RECT  12.0575 29.2625 12.1225 29.3975 ;
        RECT  11.8025 28.77 11.8675 28.905 ;
        RECT  11.8025 28.77 11.8675 28.905 ;
        RECT  11.8025 28.77 11.8675 28.905 ;
        RECT  11.8025 28.77 11.8675 28.905 ;
        RECT  11.8025 28.77 11.8675 28.905 ;
        RECT  11.8025 28.77 11.8675 28.905 ;
        RECT  12.5075 28.77 12.5725 28.905 ;
        RECT  12.5075 28.77 12.5725 28.905 ;
        RECT  12.5075 28.77 12.5725 28.905 ;
        RECT  12.5075 28.77 12.5725 28.905 ;
        RECT  12.2525 29.2625 12.3175 29.3975 ;
        RECT  12.12 29.6225 12.255 29.6875 ;
        RECT  12.12 29.6225 12.255 29.6875 ;
        RECT  12.4725 29.6225 12.6075 29.6875 ;
        RECT  12.115 28.2775 12.25 28.3425 ;
        RECT  12.4725 29.6225 12.6075 29.6875 ;
        RECT  12.4725 29.6225 12.6075 29.6875 ;
        RECT  12.5075 28.77 12.5725 28.905 ;
        RECT  12.5075 28.77 12.5725 28.905 ;
        RECT  12.5075 28.77 12.5725 28.905 ;
        RECT  12.5075 28.77 12.5725 28.905 ;
        RECT  12.5075 28.77 12.5725 28.905 ;
        RECT  12.5075 28.77 12.5725 28.905 ;
        RECT  11.7675 29.6225 11.9025 29.6875 ;
        RECT  12.1275 28.28 12.2275 28.3425 ;
        RECT  12.1275 28.2775 12.2275 28.34 ;
        RECT  12.455 29.4825 12.5075 29.545 ;
        RECT  12.1275 28.28 12.2275 28.3425 ;
        RECT  12.505 28.3425 12.575 28.5425 ;
        RECT  12.505 28.8725 12.575 29.0075 ;
        RECT  12.505 28.8725 12.575 29.0075 ;
        RECT  11.745 29.6225 12.63 29.6875 ;
        RECT  12.32 29.1075 12.495 29.1725 ;
        RECT  11.8 28.8725 11.87 29.0075 ;
        RECT  11.99 28.4325 12.055 29.1725 ;
        RECT  12.1275 28.2775 12.2275 28.34 ;
        RECT  11.75 29.4825 11.8025 29.545 ;
        RECT  12.505 28.8725 12.575 29.0075 ;
        RECT  11.745 28.2775 12.63 28.3425 ;
        RECT  12.32 28.5425 12.385 29.1725 ;
        RECT  12.505 28.8725 12.575 29.0075 ;
        RECT  12.505 28.8725 12.575 29.0075 ;
        RECT  11.885 29.1075 11.955 29.3975 ;
        RECT  11.8 28.8725 11.87 29.0075 ;
        RECT  11.745 29.4825 12.63 29.5475 ;
        RECT  12.505 28.8725 12.575 29.0075 ;
        RECT  12.505 28.3425 12.575 28.5425 ;
        RECT  11.8 28.3425 11.87 28.5425 ;
        RECT  12.425 29.1075 12.495 29.3975 ;
        RECT  11.885 29.1075 12.055 29.1725 ;
        RECT  12.505 30.7675 12.57 30.9025 ;
        RECT  12.32 30.7675 12.385 30.9025 ;
        RECT  11.805 30.7675 11.87 30.9025 ;
        RECT  11.99 30.7675 12.055 30.9025 ;
        RECT  12.32 30.3025 12.385 30.4375 ;
        RECT  12.505 30.3025 12.57 30.4375 ;
        RECT  11.99 30.3025 12.055 30.4375 ;
        RECT  11.805 30.3025 11.87 30.4375 ;
        RECT  12.425 29.9125 12.49 30.0475 ;
        RECT  12.24 29.9125 12.305 30.0475 ;
        RECT  12.07 29.9125 12.135 30.0475 ;
        RECT  11.885 29.9125 11.95 30.0475 ;
        RECT  12.5075 30.405 12.5725 30.54 ;
        RECT  12.5075 30.405 12.5725 30.54 ;
        RECT  12.5075 30.405 12.5725 30.54 ;
        RECT  12.5075 30.405 12.5725 30.54 ;
        RECT  12.5075 30.405 12.5725 30.54 ;
        RECT  12.5075 30.405 12.5725 30.54 ;
        RECT  12.115 30.9675 12.25 31.0325 ;
        RECT  11.7675 29.6225 11.9025 29.6875 ;
        RECT  12.4725 29.6225 12.6075 29.6875 ;
        RECT  12.1025 29.7625 12.2375 29.8275 ;
        RECT  12.5075 30.405 12.5725 30.54 ;
        RECT  12.5075 30.405 12.5725 30.54 ;
        RECT  12.5075 30.405 12.5725 30.54 ;
        RECT  12.5075 30.405 12.5725 30.54 ;
        RECT  12.0075 30.6525 12.1425 30.7175 ;
        RECT  12.0075 30.6525 12.1425 30.7175 ;
        RECT  12.2325 30.5025 12.3675 30.5675 ;
        RECT  12.2325 30.5025 12.3675 30.5675 ;
        RECT  12.5075 30.405 12.5725 30.54 ;
        RECT  12.5075 30.405 12.5725 30.54 ;
        RECT  12.5075 30.405 12.5725 30.54 ;
        RECT  12.5075 30.405 12.5725 30.54 ;
        RECT  12.0575 29.9125 12.1225 30.0475 ;
        RECT  11.8025 30.405 11.8675 30.54 ;
        RECT  11.8025 30.405 11.8675 30.54 ;
        RECT  11.8025 30.405 11.8675 30.54 ;
        RECT  11.8025 30.405 11.8675 30.54 ;
        RECT  11.8025 30.405 11.8675 30.54 ;
        RECT  11.8025 30.405 11.8675 30.54 ;
        RECT  12.5075 30.405 12.5725 30.54 ;
        RECT  12.5075 30.405 12.5725 30.54 ;
        RECT  12.5075 30.405 12.5725 30.54 ;
        RECT  12.5075 30.405 12.5725 30.54 ;
        RECT  12.2525 29.9125 12.3175 30.0475 ;
        RECT  12.12 29.6225 12.255 29.6875 ;
        RECT  12.12 29.6225 12.255 29.6875 ;
        RECT  12.4725 29.6225 12.6075 29.6875 ;
        RECT  12.115 30.9675 12.25 31.0325 ;
        RECT  12.4725 29.6225 12.6075 29.6875 ;
        RECT  12.4725 29.6225 12.6075 29.6875 ;
        RECT  12.5075 30.405 12.5725 30.54 ;
        RECT  12.5075 30.405 12.5725 30.54 ;
        RECT  12.5075 30.405 12.5725 30.54 ;
        RECT  12.5075 30.405 12.5725 30.54 ;
        RECT  12.5075 30.405 12.5725 30.54 ;
        RECT  12.5075 30.405 12.5725 30.54 ;
        RECT  11.7675 29.6225 11.9025 29.6875 ;
        RECT  12.1275 30.9675 12.2275 31.03 ;
        RECT  12.1275 30.97 12.2275 31.0325 ;
        RECT  12.455 29.765 12.5075 29.8275 ;
        RECT  12.1275 30.9675 12.2275 31.03 ;
        RECT  12.505 30.7675 12.575 30.9675 ;
        RECT  12.505 30.3025 12.575 30.4375 ;
        RECT  12.505 30.3025 12.575 30.4375 ;
        RECT  11.745 29.6225 12.63 29.6875 ;
        RECT  12.32 30.1375 12.495 30.2025 ;
        RECT  11.8 30.3025 11.87 30.4375 ;
        RECT  11.99 30.1375 12.055 30.8775 ;
        RECT  12.1275 30.97 12.2275 31.0325 ;
        RECT  11.75 29.765 11.8025 29.8275 ;
        RECT  12.505 30.3025 12.575 30.4375 ;
        RECT  11.745 30.9675 12.63 31.0325 ;
        RECT  12.32 30.1375 12.385 30.7675 ;
        RECT  12.505 30.3025 12.575 30.4375 ;
        RECT  12.505 30.3025 12.575 30.4375 ;
        RECT  11.885 29.9125 11.955 30.2025 ;
        RECT  11.8 30.3025 11.87 30.4375 ;
        RECT  11.745 29.7625 12.63 29.8275 ;
        RECT  12.505 30.3025 12.575 30.4375 ;
        RECT  12.505 30.7675 12.575 30.9675 ;
        RECT  11.8 30.7675 11.87 30.9675 ;
        RECT  12.425 29.9125 12.495 30.2025 ;
        RECT  11.885 30.1375 12.055 30.2025 ;
        RECT  12.505 31.0975 12.57 31.2325 ;
        RECT  12.32 31.0975 12.385 31.2325 ;
        RECT  11.805 31.0975 11.87 31.2325 ;
        RECT  11.99 31.0975 12.055 31.2325 ;
        RECT  12.32 31.5625 12.385 31.6975 ;
        RECT  12.505 31.5625 12.57 31.6975 ;
        RECT  11.99 31.5625 12.055 31.6975 ;
        RECT  11.805 31.5625 11.87 31.6975 ;
        RECT  12.425 31.9525 12.49 32.0875 ;
        RECT  12.24 31.9525 12.305 32.0875 ;
        RECT  12.07 31.9525 12.135 32.0875 ;
        RECT  11.885 31.9525 11.95 32.0875 ;
        RECT  12.5075 31.46 12.5725 31.595 ;
        RECT  12.5075 31.46 12.5725 31.595 ;
        RECT  12.5075 31.46 12.5725 31.595 ;
        RECT  12.5075 31.46 12.5725 31.595 ;
        RECT  12.5075 31.46 12.5725 31.595 ;
        RECT  12.5075 31.46 12.5725 31.595 ;
        RECT  12.115 30.9675 12.25 31.0325 ;
        RECT  11.7675 32.3125 11.9025 32.3775 ;
        RECT  12.4725 32.3125 12.6075 32.3775 ;
        RECT  12.1025 32.1725 12.2375 32.2375 ;
        RECT  12.5075 31.46 12.5725 31.595 ;
        RECT  12.5075 31.46 12.5725 31.595 ;
        RECT  12.5075 31.46 12.5725 31.595 ;
        RECT  12.5075 31.46 12.5725 31.595 ;
        RECT  12.0075 31.2825 12.1425 31.3475 ;
        RECT  12.0075 31.2825 12.1425 31.3475 ;
        RECT  12.2325 31.4325 12.3675 31.4975 ;
        RECT  12.2325 31.4325 12.3675 31.4975 ;
        RECT  12.5075 31.46 12.5725 31.595 ;
        RECT  12.5075 31.46 12.5725 31.595 ;
        RECT  12.5075 31.46 12.5725 31.595 ;
        RECT  12.5075 31.46 12.5725 31.595 ;
        RECT  12.0575 31.9525 12.1225 32.0875 ;
        RECT  11.8025 31.46 11.8675 31.595 ;
        RECT  11.8025 31.46 11.8675 31.595 ;
        RECT  11.8025 31.46 11.8675 31.595 ;
        RECT  11.8025 31.46 11.8675 31.595 ;
        RECT  11.8025 31.46 11.8675 31.595 ;
        RECT  11.8025 31.46 11.8675 31.595 ;
        RECT  12.5075 31.46 12.5725 31.595 ;
        RECT  12.5075 31.46 12.5725 31.595 ;
        RECT  12.5075 31.46 12.5725 31.595 ;
        RECT  12.5075 31.46 12.5725 31.595 ;
        RECT  12.2525 31.9525 12.3175 32.0875 ;
        RECT  12.12 32.3125 12.255 32.3775 ;
        RECT  12.12 32.3125 12.255 32.3775 ;
        RECT  12.4725 32.3125 12.6075 32.3775 ;
        RECT  12.115 30.9675 12.25 31.0325 ;
        RECT  12.4725 32.3125 12.6075 32.3775 ;
        RECT  12.4725 32.3125 12.6075 32.3775 ;
        RECT  12.5075 31.46 12.5725 31.595 ;
        RECT  12.5075 31.46 12.5725 31.595 ;
        RECT  12.5075 31.46 12.5725 31.595 ;
        RECT  12.5075 31.46 12.5725 31.595 ;
        RECT  12.5075 31.46 12.5725 31.595 ;
        RECT  12.5075 31.46 12.5725 31.595 ;
        RECT  11.7675 32.3125 11.9025 32.3775 ;
        RECT  12.1275 30.97 12.2275 31.0325 ;
        RECT  12.1275 30.9675 12.2275 31.03 ;
        RECT  12.455 32.1725 12.5075 32.235 ;
        RECT  12.1275 30.97 12.2275 31.0325 ;
        RECT  12.505 31.0325 12.575 31.2325 ;
        RECT  12.505 31.5625 12.575 31.6975 ;
        RECT  12.505 31.5625 12.575 31.6975 ;
        RECT  11.745 32.3125 12.63 32.3775 ;
        RECT  12.32 31.7975 12.495 31.8625 ;
        RECT  11.8 31.5625 11.87 31.6975 ;
        RECT  11.99 31.1225 12.055 31.8625 ;
        RECT  12.1275 30.9675 12.2275 31.03 ;
        RECT  11.75 32.1725 11.8025 32.235 ;
        RECT  12.505 31.5625 12.575 31.6975 ;
        RECT  11.745 30.9675 12.63 31.0325 ;
        RECT  12.32 31.2325 12.385 31.8625 ;
        RECT  12.505 31.5625 12.575 31.6975 ;
        RECT  12.505 31.5625 12.575 31.6975 ;
        RECT  11.885 31.7975 11.955 32.0875 ;
        RECT  11.8 31.5625 11.87 31.6975 ;
        RECT  11.745 32.1725 12.63 32.2375 ;
        RECT  12.505 31.5625 12.575 31.6975 ;
        RECT  12.505 31.0325 12.575 31.2325 ;
        RECT  11.8 31.0325 11.87 31.2325 ;
        RECT  12.425 31.7975 12.495 32.0875 ;
        RECT  11.885 31.7975 12.055 31.8625 ;
        RECT  12.505 33.4575 12.57 33.5925 ;
        RECT  12.32 33.4575 12.385 33.5925 ;
        RECT  11.805 33.4575 11.87 33.5925 ;
        RECT  11.99 33.4575 12.055 33.5925 ;
        RECT  12.32 32.9925 12.385 33.1275 ;
        RECT  12.505 32.9925 12.57 33.1275 ;
        RECT  11.99 32.9925 12.055 33.1275 ;
        RECT  11.805 32.9925 11.87 33.1275 ;
        RECT  12.425 32.6025 12.49 32.7375 ;
        RECT  12.24 32.6025 12.305 32.7375 ;
        RECT  12.07 32.6025 12.135 32.7375 ;
        RECT  11.885 32.6025 11.95 32.7375 ;
        RECT  12.5075 33.095 12.5725 33.23 ;
        RECT  12.5075 33.095 12.5725 33.23 ;
        RECT  12.5075 33.095 12.5725 33.23 ;
        RECT  12.5075 33.095 12.5725 33.23 ;
        RECT  12.5075 33.095 12.5725 33.23 ;
        RECT  12.5075 33.095 12.5725 33.23 ;
        RECT  12.115 33.6575 12.25 33.7225 ;
        RECT  11.7675 32.3125 11.9025 32.3775 ;
        RECT  12.4725 32.3125 12.6075 32.3775 ;
        RECT  12.1025 32.4525 12.2375 32.5175 ;
        RECT  12.5075 33.095 12.5725 33.23 ;
        RECT  12.5075 33.095 12.5725 33.23 ;
        RECT  12.5075 33.095 12.5725 33.23 ;
        RECT  12.5075 33.095 12.5725 33.23 ;
        RECT  12.0075 33.3425 12.1425 33.4075 ;
        RECT  12.0075 33.3425 12.1425 33.4075 ;
        RECT  12.2325 33.1925 12.3675 33.2575 ;
        RECT  12.2325 33.1925 12.3675 33.2575 ;
        RECT  12.5075 33.095 12.5725 33.23 ;
        RECT  12.5075 33.095 12.5725 33.23 ;
        RECT  12.5075 33.095 12.5725 33.23 ;
        RECT  12.5075 33.095 12.5725 33.23 ;
        RECT  12.0575 32.6025 12.1225 32.7375 ;
        RECT  11.8025 33.095 11.8675 33.23 ;
        RECT  11.8025 33.095 11.8675 33.23 ;
        RECT  11.8025 33.095 11.8675 33.23 ;
        RECT  11.8025 33.095 11.8675 33.23 ;
        RECT  11.8025 33.095 11.8675 33.23 ;
        RECT  11.8025 33.095 11.8675 33.23 ;
        RECT  12.5075 33.095 12.5725 33.23 ;
        RECT  12.5075 33.095 12.5725 33.23 ;
        RECT  12.5075 33.095 12.5725 33.23 ;
        RECT  12.5075 33.095 12.5725 33.23 ;
        RECT  12.2525 32.6025 12.3175 32.7375 ;
        RECT  12.12 32.3125 12.255 32.3775 ;
        RECT  12.12 32.3125 12.255 32.3775 ;
        RECT  12.4725 32.3125 12.6075 32.3775 ;
        RECT  12.115 33.6575 12.25 33.7225 ;
        RECT  12.4725 32.3125 12.6075 32.3775 ;
        RECT  12.4725 32.3125 12.6075 32.3775 ;
        RECT  12.5075 33.095 12.5725 33.23 ;
        RECT  12.5075 33.095 12.5725 33.23 ;
        RECT  12.5075 33.095 12.5725 33.23 ;
        RECT  12.5075 33.095 12.5725 33.23 ;
        RECT  12.5075 33.095 12.5725 33.23 ;
        RECT  12.5075 33.095 12.5725 33.23 ;
        RECT  11.7675 32.3125 11.9025 32.3775 ;
        RECT  12.1275 33.6575 12.2275 33.72 ;
        RECT  12.1275 33.66 12.2275 33.7225 ;
        RECT  12.455 32.455 12.5075 32.5175 ;
        RECT  12.1275 33.6575 12.2275 33.72 ;
        RECT  12.505 33.4575 12.575 33.6575 ;
        RECT  12.505 32.9925 12.575 33.1275 ;
        RECT  12.505 32.9925 12.575 33.1275 ;
        RECT  11.745 32.3125 12.63 32.3775 ;
        RECT  12.32 32.8275 12.495 32.8925 ;
        RECT  11.8 32.9925 11.87 33.1275 ;
        RECT  11.99 32.8275 12.055 33.5675 ;
        RECT  12.1275 33.66 12.2275 33.7225 ;
        RECT  11.75 32.455 11.8025 32.5175 ;
        RECT  12.505 32.9925 12.575 33.1275 ;
        RECT  11.745 33.6575 12.63 33.7225 ;
        RECT  12.32 32.8275 12.385 33.4575 ;
        RECT  12.505 32.9925 12.575 33.1275 ;
        RECT  12.505 32.9925 12.575 33.1275 ;
        RECT  11.885 32.6025 11.955 32.8925 ;
        RECT  11.8 32.9925 11.87 33.1275 ;
        RECT  11.745 32.4525 12.63 32.5175 ;
        RECT  12.505 32.9925 12.575 33.1275 ;
        RECT  12.505 33.4575 12.575 33.6575 ;
        RECT  11.8 33.4575 11.87 33.6575 ;
        RECT  12.425 32.6025 12.495 32.8925 ;
        RECT  11.885 32.8275 12.055 32.8925 ;
        RECT  12.505 33.7875 12.57 33.9225 ;
        RECT  12.32 33.7875 12.385 33.9225 ;
        RECT  11.805 33.7875 11.87 33.9225 ;
        RECT  11.99 33.7875 12.055 33.9225 ;
        RECT  12.32 34.2525 12.385 34.3875 ;
        RECT  12.505 34.2525 12.57 34.3875 ;
        RECT  11.99 34.2525 12.055 34.3875 ;
        RECT  11.805 34.2525 11.87 34.3875 ;
        RECT  12.425 34.6425 12.49 34.7775 ;
        RECT  12.24 34.6425 12.305 34.7775 ;
        RECT  12.07 34.6425 12.135 34.7775 ;
        RECT  11.885 34.6425 11.95 34.7775 ;
        RECT  12.5075 34.15 12.5725 34.285 ;
        RECT  12.5075 34.15 12.5725 34.285 ;
        RECT  12.5075 34.15 12.5725 34.285 ;
        RECT  12.5075 34.15 12.5725 34.285 ;
        RECT  12.5075 34.15 12.5725 34.285 ;
        RECT  12.5075 34.15 12.5725 34.285 ;
        RECT  12.115 33.6575 12.25 33.7225 ;
        RECT  11.7675 35.0025 11.9025 35.0675 ;
        RECT  12.4725 35.0025 12.6075 35.0675 ;
        RECT  12.1025 34.8625 12.2375 34.9275 ;
        RECT  12.5075 34.15 12.5725 34.285 ;
        RECT  12.5075 34.15 12.5725 34.285 ;
        RECT  12.5075 34.15 12.5725 34.285 ;
        RECT  12.5075 34.15 12.5725 34.285 ;
        RECT  12.0075 33.9725 12.1425 34.0375 ;
        RECT  12.0075 33.9725 12.1425 34.0375 ;
        RECT  12.2325 34.1225 12.3675 34.1875 ;
        RECT  12.2325 34.1225 12.3675 34.1875 ;
        RECT  12.5075 34.15 12.5725 34.285 ;
        RECT  12.5075 34.15 12.5725 34.285 ;
        RECT  12.5075 34.15 12.5725 34.285 ;
        RECT  12.5075 34.15 12.5725 34.285 ;
        RECT  12.0575 34.6425 12.1225 34.7775 ;
        RECT  11.8025 34.15 11.8675 34.285 ;
        RECT  11.8025 34.15 11.8675 34.285 ;
        RECT  11.8025 34.15 11.8675 34.285 ;
        RECT  11.8025 34.15 11.8675 34.285 ;
        RECT  11.8025 34.15 11.8675 34.285 ;
        RECT  11.8025 34.15 11.8675 34.285 ;
        RECT  12.5075 34.15 12.5725 34.285 ;
        RECT  12.5075 34.15 12.5725 34.285 ;
        RECT  12.5075 34.15 12.5725 34.285 ;
        RECT  12.5075 34.15 12.5725 34.285 ;
        RECT  12.2525 34.6425 12.3175 34.7775 ;
        RECT  12.12 35.0025 12.255 35.0675 ;
        RECT  12.12 35.0025 12.255 35.0675 ;
        RECT  12.4725 35.0025 12.6075 35.0675 ;
        RECT  12.115 33.6575 12.25 33.7225 ;
        RECT  12.4725 35.0025 12.6075 35.0675 ;
        RECT  12.4725 35.0025 12.6075 35.0675 ;
        RECT  12.5075 34.15 12.5725 34.285 ;
        RECT  12.5075 34.15 12.5725 34.285 ;
        RECT  12.5075 34.15 12.5725 34.285 ;
        RECT  12.5075 34.15 12.5725 34.285 ;
        RECT  12.5075 34.15 12.5725 34.285 ;
        RECT  12.5075 34.15 12.5725 34.285 ;
        RECT  11.7675 35.0025 11.9025 35.0675 ;
        RECT  12.1275 33.66 12.2275 33.7225 ;
        RECT  12.1275 33.6575 12.2275 33.72 ;
        RECT  12.455 34.8625 12.5075 34.925 ;
        RECT  12.1275 33.66 12.2275 33.7225 ;
        RECT  12.505 33.7225 12.575 33.9225 ;
        RECT  12.505 34.2525 12.575 34.3875 ;
        RECT  12.505 34.2525 12.575 34.3875 ;
        RECT  11.745 35.0025 12.63 35.0675 ;
        RECT  12.32 34.4875 12.495 34.5525 ;
        RECT  11.8 34.2525 11.87 34.3875 ;
        RECT  11.99 33.8125 12.055 34.5525 ;
        RECT  12.1275 33.6575 12.2275 33.72 ;
        RECT  11.75 34.8625 11.8025 34.925 ;
        RECT  12.505 34.2525 12.575 34.3875 ;
        RECT  11.745 33.6575 12.63 33.7225 ;
        RECT  12.32 33.9225 12.385 34.5525 ;
        RECT  12.505 34.2525 12.575 34.3875 ;
        RECT  12.505 34.2525 12.575 34.3875 ;
        RECT  11.885 34.4875 11.955 34.7775 ;
        RECT  11.8 34.2525 11.87 34.3875 ;
        RECT  11.745 34.8625 12.63 34.9275 ;
        RECT  12.505 34.2525 12.575 34.3875 ;
        RECT  12.505 33.7225 12.575 33.9225 ;
        RECT  11.8 33.7225 11.87 33.9225 ;
        RECT  12.425 34.4875 12.495 34.7775 ;
        RECT  11.885 34.4875 12.055 34.5525 ;
        RECT  12.505 36.1475 12.57 36.2825 ;
        RECT  12.32 36.1475 12.385 36.2825 ;
        RECT  11.805 36.1475 11.87 36.2825 ;
        RECT  11.99 36.1475 12.055 36.2825 ;
        RECT  12.32 35.6825 12.385 35.8175 ;
        RECT  12.505 35.6825 12.57 35.8175 ;
        RECT  11.99 35.6825 12.055 35.8175 ;
        RECT  11.805 35.6825 11.87 35.8175 ;
        RECT  12.425 35.2925 12.49 35.4275 ;
        RECT  12.24 35.2925 12.305 35.4275 ;
        RECT  12.07 35.2925 12.135 35.4275 ;
        RECT  11.885 35.2925 11.95 35.4275 ;
        RECT  12.5075 35.785 12.5725 35.92 ;
        RECT  12.5075 35.785 12.5725 35.92 ;
        RECT  12.5075 35.785 12.5725 35.92 ;
        RECT  12.5075 35.785 12.5725 35.92 ;
        RECT  12.5075 35.785 12.5725 35.92 ;
        RECT  12.5075 35.785 12.5725 35.92 ;
        RECT  12.115 36.3475 12.25 36.4125 ;
        RECT  11.7675 35.0025 11.9025 35.0675 ;
        RECT  12.4725 35.0025 12.6075 35.0675 ;
        RECT  12.1025 35.1425 12.2375 35.2075 ;
        RECT  12.5075 35.785 12.5725 35.92 ;
        RECT  12.5075 35.785 12.5725 35.92 ;
        RECT  12.5075 35.785 12.5725 35.92 ;
        RECT  12.5075 35.785 12.5725 35.92 ;
        RECT  12.0075 36.0325 12.1425 36.0975 ;
        RECT  12.0075 36.0325 12.1425 36.0975 ;
        RECT  12.2325 35.8825 12.3675 35.9475 ;
        RECT  12.2325 35.8825 12.3675 35.9475 ;
        RECT  12.5075 35.785 12.5725 35.92 ;
        RECT  12.5075 35.785 12.5725 35.92 ;
        RECT  12.5075 35.785 12.5725 35.92 ;
        RECT  12.5075 35.785 12.5725 35.92 ;
        RECT  12.0575 35.2925 12.1225 35.4275 ;
        RECT  11.8025 35.785 11.8675 35.92 ;
        RECT  11.8025 35.785 11.8675 35.92 ;
        RECT  11.8025 35.785 11.8675 35.92 ;
        RECT  11.8025 35.785 11.8675 35.92 ;
        RECT  11.8025 35.785 11.8675 35.92 ;
        RECT  11.8025 35.785 11.8675 35.92 ;
        RECT  12.5075 35.785 12.5725 35.92 ;
        RECT  12.5075 35.785 12.5725 35.92 ;
        RECT  12.5075 35.785 12.5725 35.92 ;
        RECT  12.5075 35.785 12.5725 35.92 ;
        RECT  12.2525 35.2925 12.3175 35.4275 ;
        RECT  12.12 35.0025 12.255 35.0675 ;
        RECT  12.12 35.0025 12.255 35.0675 ;
        RECT  12.4725 35.0025 12.6075 35.0675 ;
        RECT  12.115 36.3475 12.25 36.4125 ;
        RECT  12.4725 35.0025 12.6075 35.0675 ;
        RECT  12.4725 35.0025 12.6075 35.0675 ;
        RECT  12.5075 35.785 12.5725 35.92 ;
        RECT  12.5075 35.785 12.5725 35.92 ;
        RECT  12.5075 35.785 12.5725 35.92 ;
        RECT  12.5075 35.785 12.5725 35.92 ;
        RECT  12.5075 35.785 12.5725 35.92 ;
        RECT  12.5075 35.785 12.5725 35.92 ;
        RECT  11.7675 35.0025 11.9025 35.0675 ;
        RECT  12.1275 36.3475 12.2275 36.41 ;
        RECT  12.1275 36.35 12.2275 36.4125 ;
        RECT  12.455 35.145 12.5075 35.2075 ;
        RECT  12.1275 36.3475 12.2275 36.41 ;
        RECT  12.505 36.1475 12.575 36.3475 ;
        RECT  12.505 35.6825 12.575 35.8175 ;
        RECT  12.505 35.6825 12.575 35.8175 ;
        RECT  11.745 35.0025 12.63 35.0675 ;
        RECT  12.32 35.5175 12.495 35.5825 ;
        RECT  11.8 35.6825 11.87 35.8175 ;
        RECT  11.99 35.5175 12.055 36.2575 ;
        RECT  12.1275 36.35 12.2275 36.4125 ;
        RECT  11.75 35.145 11.8025 35.2075 ;
        RECT  12.505 35.6825 12.575 35.8175 ;
        RECT  11.745 36.3475 12.63 36.4125 ;
        RECT  12.32 35.5175 12.385 36.1475 ;
        RECT  12.505 35.6825 12.575 35.8175 ;
        RECT  12.505 35.6825 12.575 35.8175 ;
        RECT  11.885 35.2925 11.955 35.5825 ;
        RECT  11.8 35.6825 11.87 35.8175 ;
        RECT  11.745 35.1425 12.63 35.2075 ;
        RECT  12.505 35.6825 12.575 35.8175 ;
        RECT  12.505 36.1475 12.575 36.3475 ;
        RECT  11.8 36.1475 11.87 36.3475 ;
        RECT  12.425 35.2925 12.495 35.5825 ;
        RECT  11.885 35.5175 12.055 35.5825 ;
        RECT  12.505 36.4775 12.57 36.6125 ;
        RECT  12.32 36.4775 12.385 36.6125 ;
        RECT  11.805 36.4775 11.87 36.6125 ;
        RECT  11.99 36.4775 12.055 36.6125 ;
        RECT  12.32 36.9425 12.385 37.0775 ;
        RECT  12.505 36.9425 12.57 37.0775 ;
        RECT  11.99 36.9425 12.055 37.0775 ;
        RECT  11.805 36.9425 11.87 37.0775 ;
        RECT  12.425 37.3325 12.49 37.4675 ;
        RECT  12.24 37.3325 12.305 37.4675 ;
        RECT  12.07 37.3325 12.135 37.4675 ;
        RECT  11.885 37.3325 11.95 37.4675 ;
        RECT  12.5075 36.84 12.5725 36.975 ;
        RECT  12.5075 36.84 12.5725 36.975 ;
        RECT  12.5075 36.84 12.5725 36.975 ;
        RECT  12.5075 36.84 12.5725 36.975 ;
        RECT  12.5075 36.84 12.5725 36.975 ;
        RECT  12.5075 36.84 12.5725 36.975 ;
        RECT  12.115 36.3475 12.25 36.4125 ;
        RECT  11.7675 37.6925 11.9025 37.7575 ;
        RECT  12.4725 37.6925 12.6075 37.7575 ;
        RECT  12.1025 37.5525 12.2375 37.6175 ;
        RECT  12.5075 36.84 12.5725 36.975 ;
        RECT  12.5075 36.84 12.5725 36.975 ;
        RECT  12.5075 36.84 12.5725 36.975 ;
        RECT  12.5075 36.84 12.5725 36.975 ;
        RECT  12.0075 36.6625 12.1425 36.7275 ;
        RECT  12.0075 36.6625 12.1425 36.7275 ;
        RECT  12.2325 36.8125 12.3675 36.8775 ;
        RECT  12.2325 36.8125 12.3675 36.8775 ;
        RECT  12.5075 36.84 12.5725 36.975 ;
        RECT  12.5075 36.84 12.5725 36.975 ;
        RECT  12.5075 36.84 12.5725 36.975 ;
        RECT  12.5075 36.84 12.5725 36.975 ;
        RECT  12.0575 37.3325 12.1225 37.4675 ;
        RECT  11.8025 36.84 11.8675 36.975 ;
        RECT  11.8025 36.84 11.8675 36.975 ;
        RECT  11.8025 36.84 11.8675 36.975 ;
        RECT  11.8025 36.84 11.8675 36.975 ;
        RECT  11.8025 36.84 11.8675 36.975 ;
        RECT  11.8025 36.84 11.8675 36.975 ;
        RECT  12.5075 36.84 12.5725 36.975 ;
        RECT  12.5075 36.84 12.5725 36.975 ;
        RECT  12.5075 36.84 12.5725 36.975 ;
        RECT  12.5075 36.84 12.5725 36.975 ;
        RECT  12.2525 37.3325 12.3175 37.4675 ;
        RECT  12.12 37.6925 12.255 37.7575 ;
        RECT  12.12 37.6925 12.255 37.7575 ;
        RECT  12.4725 37.6925 12.6075 37.7575 ;
        RECT  12.115 36.3475 12.25 36.4125 ;
        RECT  12.4725 37.6925 12.6075 37.7575 ;
        RECT  12.4725 37.6925 12.6075 37.7575 ;
        RECT  12.5075 36.84 12.5725 36.975 ;
        RECT  12.5075 36.84 12.5725 36.975 ;
        RECT  12.5075 36.84 12.5725 36.975 ;
        RECT  12.5075 36.84 12.5725 36.975 ;
        RECT  12.5075 36.84 12.5725 36.975 ;
        RECT  12.5075 36.84 12.5725 36.975 ;
        RECT  11.7675 37.6925 11.9025 37.7575 ;
        RECT  12.1275 36.35 12.2275 36.4125 ;
        RECT  12.1275 36.3475 12.2275 36.41 ;
        RECT  12.455 37.5525 12.5075 37.615 ;
        RECT  12.1275 36.35 12.2275 36.4125 ;
        RECT  12.505 36.4125 12.575 36.6125 ;
        RECT  12.505 36.9425 12.575 37.0775 ;
        RECT  12.505 36.9425 12.575 37.0775 ;
        RECT  11.745 37.6925 12.63 37.7575 ;
        RECT  12.32 37.1775 12.495 37.2425 ;
        RECT  11.8 36.9425 11.87 37.0775 ;
        RECT  11.99 36.5025 12.055 37.2425 ;
        RECT  12.1275 36.3475 12.2275 36.41 ;
        RECT  11.75 37.5525 11.8025 37.615 ;
        RECT  12.505 36.9425 12.575 37.0775 ;
        RECT  11.745 36.3475 12.63 36.4125 ;
        RECT  12.32 36.6125 12.385 37.2425 ;
        RECT  12.505 36.9425 12.575 37.0775 ;
        RECT  12.505 36.9425 12.575 37.0775 ;
        RECT  11.885 37.1775 11.955 37.4675 ;
        RECT  11.8 36.9425 11.87 37.0775 ;
        RECT  11.745 37.5525 12.63 37.6175 ;
        RECT  12.505 36.9425 12.575 37.0775 ;
        RECT  12.505 36.4125 12.575 36.6125 ;
        RECT  11.8 36.4125 11.87 36.6125 ;
        RECT  12.425 37.1775 12.495 37.4675 ;
        RECT  11.885 37.1775 12.055 37.2425 ;
        RECT  12.505 38.8375 12.57 38.9725 ;
        RECT  12.32 38.8375 12.385 38.9725 ;
        RECT  11.805 38.8375 11.87 38.9725 ;
        RECT  11.99 38.8375 12.055 38.9725 ;
        RECT  12.32 38.3725 12.385 38.5075 ;
        RECT  12.505 38.3725 12.57 38.5075 ;
        RECT  11.99 38.3725 12.055 38.5075 ;
        RECT  11.805 38.3725 11.87 38.5075 ;
        RECT  12.425 37.9825 12.49 38.1175 ;
        RECT  12.24 37.9825 12.305 38.1175 ;
        RECT  12.07 37.9825 12.135 38.1175 ;
        RECT  11.885 37.9825 11.95 38.1175 ;
        RECT  12.5075 38.475 12.5725 38.61 ;
        RECT  12.5075 38.475 12.5725 38.61 ;
        RECT  12.5075 38.475 12.5725 38.61 ;
        RECT  12.5075 38.475 12.5725 38.61 ;
        RECT  12.5075 38.475 12.5725 38.61 ;
        RECT  12.5075 38.475 12.5725 38.61 ;
        RECT  12.115 39.0375 12.25 39.1025 ;
        RECT  11.7675 37.6925 11.9025 37.7575 ;
        RECT  12.4725 37.6925 12.6075 37.7575 ;
        RECT  12.1025 37.8325 12.2375 37.8975 ;
        RECT  12.5075 38.475 12.5725 38.61 ;
        RECT  12.5075 38.475 12.5725 38.61 ;
        RECT  12.5075 38.475 12.5725 38.61 ;
        RECT  12.5075 38.475 12.5725 38.61 ;
        RECT  12.0075 38.7225 12.1425 38.7875 ;
        RECT  12.0075 38.7225 12.1425 38.7875 ;
        RECT  12.2325 38.5725 12.3675 38.6375 ;
        RECT  12.2325 38.5725 12.3675 38.6375 ;
        RECT  12.5075 38.475 12.5725 38.61 ;
        RECT  12.5075 38.475 12.5725 38.61 ;
        RECT  12.5075 38.475 12.5725 38.61 ;
        RECT  12.5075 38.475 12.5725 38.61 ;
        RECT  12.0575 37.9825 12.1225 38.1175 ;
        RECT  11.8025 38.475 11.8675 38.61 ;
        RECT  11.8025 38.475 11.8675 38.61 ;
        RECT  11.8025 38.475 11.8675 38.61 ;
        RECT  11.8025 38.475 11.8675 38.61 ;
        RECT  11.8025 38.475 11.8675 38.61 ;
        RECT  11.8025 38.475 11.8675 38.61 ;
        RECT  12.5075 38.475 12.5725 38.61 ;
        RECT  12.5075 38.475 12.5725 38.61 ;
        RECT  12.5075 38.475 12.5725 38.61 ;
        RECT  12.5075 38.475 12.5725 38.61 ;
        RECT  12.2525 37.9825 12.3175 38.1175 ;
        RECT  12.12 37.6925 12.255 37.7575 ;
        RECT  12.12 37.6925 12.255 37.7575 ;
        RECT  12.4725 37.6925 12.6075 37.7575 ;
        RECT  12.115 39.0375 12.25 39.1025 ;
        RECT  12.4725 37.6925 12.6075 37.7575 ;
        RECT  12.4725 37.6925 12.6075 37.7575 ;
        RECT  12.5075 38.475 12.5725 38.61 ;
        RECT  12.5075 38.475 12.5725 38.61 ;
        RECT  12.5075 38.475 12.5725 38.61 ;
        RECT  12.5075 38.475 12.5725 38.61 ;
        RECT  12.5075 38.475 12.5725 38.61 ;
        RECT  12.5075 38.475 12.5725 38.61 ;
        RECT  11.7675 37.6925 11.9025 37.7575 ;
        RECT  12.1275 39.0375 12.2275 39.1 ;
        RECT  12.1275 39.04 12.2275 39.1025 ;
        RECT  12.455 37.835 12.5075 37.8975 ;
        RECT  12.1275 39.0375 12.2275 39.1 ;
        RECT  12.505 38.8375 12.575 39.0375 ;
        RECT  12.505 38.3725 12.575 38.5075 ;
        RECT  12.505 38.3725 12.575 38.5075 ;
        RECT  11.745 37.6925 12.63 37.7575 ;
        RECT  12.32 38.2075 12.495 38.2725 ;
        RECT  11.8 38.3725 11.87 38.5075 ;
        RECT  11.99 38.2075 12.055 38.9475 ;
        RECT  12.1275 39.04 12.2275 39.1025 ;
        RECT  11.75 37.835 11.8025 37.8975 ;
        RECT  12.505 38.3725 12.575 38.5075 ;
        RECT  11.745 39.0375 12.63 39.1025 ;
        RECT  12.32 38.2075 12.385 38.8375 ;
        RECT  12.505 38.3725 12.575 38.5075 ;
        RECT  12.505 38.3725 12.575 38.5075 ;
        RECT  11.885 37.9825 11.955 38.2725 ;
        RECT  11.8 38.3725 11.87 38.5075 ;
        RECT  11.745 37.8325 12.63 37.8975 ;
        RECT  12.505 38.3725 12.575 38.5075 ;
        RECT  12.505 38.8375 12.575 39.0375 ;
        RECT  11.8 38.8375 11.87 39.0375 ;
        RECT  12.425 37.9825 12.495 38.2725 ;
        RECT  11.885 38.2075 12.055 38.2725 ;
        RECT  12.505 39.1675 12.57 39.3025 ;
        RECT  12.32 39.1675 12.385 39.3025 ;
        RECT  11.805 39.1675 11.87 39.3025 ;
        RECT  11.99 39.1675 12.055 39.3025 ;
        RECT  12.32 39.6325 12.385 39.7675 ;
        RECT  12.505 39.6325 12.57 39.7675 ;
        RECT  11.99 39.6325 12.055 39.7675 ;
        RECT  11.805 39.6325 11.87 39.7675 ;
        RECT  12.425 40.0225 12.49 40.1575 ;
        RECT  12.24 40.0225 12.305 40.1575 ;
        RECT  12.07 40.0225 12.135 40.1575 ;
        RECT  11.885 40.0225 11.95 40.1575 ;
        RECT  12.5075 39.53 12.5725 39.665 ;
        RECT  12.5075 39.53 12.5725 39.665 ;
        RECT  12.5075 39.53 12.5725 39.665 ;
        RECT  12.5075 39.53 12.5725 39.665 ;
        RECT  12.5075 39.53 12.5725 39.665 ;
        RECT  12.5075 39.53 12.5725 39.665 ;
        RECT  12.115 39.0375 12.25 39.1025 ;
        RECT  11.7675 40.3825 11.9025 40.4475 ;
        RECT  12.4725 40.3825 12.6075 40.4475 ;
        RECT  12.1025 40.2425 12.2375 40.3075 ;
        RECT  12.5075 39.53 12.5725 39.665 ;
        RECT  12.5075 39.53 12.5725 39.665 ;
        RECT  12.5075 39.53 12.5725 39.665 ;
        RECT  12.5075 39.53 12.5725 39.665 ;
        RECT  12.0075 39.3525 12.1425 39.4175 ;
        RECT  12.0075 39.3525 12.1425 39.4175 ;
        RECT  12.2325 39.5025 12.3675 39.5675 ;
        RECT  12.2325 39.5025 12.3675 39.5675 ;
        RECT  12.5075 39.53 12.5725 39.665 ;
        RECT  12.5075 39.53 12.5725 39.665 ;
        RECT  12.5075 39.53 12.5725 39.665 ;
        RECT  12.5075 39.53 12.5725 39.665 ;
        RECT  12.0575 40.0225 12.1225 40.1575 ;
        RECT  11.8025 39.53 11.8675 39.665 ;
        RECT  11.8025 39.53 11.8675 39.665 ;
        RECT  11.8025 39.53 11.8675 39.665 ;
        RECT  11.8025 39.53 11.8675 39.665 ;
        RECT  11.8025 39.53 11.8675 39.665 ;
        RECT  11.8025 39.53 11.8675 39.665 ;
        RECT  12.5075 39.53 12.5725 39.665 ;
        RECT  12.5075 39.53 12.5725 39.665 ;
        RECT  12.5075 39.53 12.5725 39.665 ;
        RECT  12.5075 39.53 12.5725 39.665 ;
        RECT  12.2525 40.0225 12.3175 40.1575 ;
        RECT  12.12 40.3825 12.255 40.4475 ;
        RECT  12.12 40.3825 12.255 40.4475 ;
        RECT  12.4725 40.3825 12.6075 40.4475 ;
        RECT  12.115 39.0375 12.25 39.1025 ;
        RECT  12.4725 40.3825 12.6075 40.4475 ;
        RECT  12.4725 40.3825 12.6075 40.4475 ;
        RECT  12.5075 39.53 12.5725 39.665 ;
        RECT  12.5075 39.53 12.5725 39.665 ;
        RECT  12.5075 39.53 12.5725 39.665 ;
        RECT  12.5075 39.53 12.5725 39.665 ;
        RECT  12.5075 39.53 12.5725 39.665 ;
        RECT  12.5075 39.53 12.5725 39.665 ;
        RECT  11.7675 40.3825 11.9025 40.4475 ;
        RECT  12.1275 39.04 12.2275 39.1025 ;
        RECT  12.1275 39.0375 12.2275 39.1 ;
        RECT  12.455 40.2425 12.5075 40.305 ;
        RECT  12.1275 39.04 12.2275 39.1025 ;
        RECT  12.505 39.1025 12.575 39.3025 ;
        RECT  12.505 39.6325 12.575 39.7675 ;
        RECT  12.505 39.6325 12.575 39.7675 ;
        RECT  11.745 40.3825 12.63 40.4475 ;
        RECT  12.32 39.8675 12.495 39.9325 ;
        RECT  11.8 39.6325 11.87 39.7675 ;
        RECT  11.99 39.1925 12.055 39.9325 ;
        RECT  12.1275 39.0375 12.2275 39.1 ;
        RECT  11.75 40.2425 11.8025 40.305 ;
        RECT  12.505 39.6325 12.575 39.7675 ;
        RECT  11.745 39.0375 12.63 39.1025 ;
        RECT  12.32 39.3025 12.385 39.9325 ;
        RECT  12.505 39.6325 12.575 39.7675 ;
        RECT  12.505 39.6325 12.575 39.7675 ;
        RECT  11.885 39.8675 11.955 40.1575 ;
        RECT  11.8 39.6325 11.87 39.7675 ;
        RECT  11.745 40.2425 12.63 40.3075 ;
        RECT  12.505 39.6325 12.575 39.7675 ;
        RECT  12.505 39.1025 12.575 39.3025 ;
        RECT  11.8 39.1025 11.87 39.3025 ;
        RECT  12.425 39.8675 12.495 40.1575 ;
        RECT  11.885 39.8675 12.055 39.9325 ;
        RECT  11.13 41.66 12.54 41.725 ;
        RECT  11.13 41.1 12.54 41.165 ;
        RECT  11.13 41.1 11.835 41.165 ;
        RECT  11.13 41.66 11.835 41.725 ;
        RECT  11.515 41.3125 11.58 41.725 ;
        RECT  11.325 40.8625 11.39 40.9975 ;
        RECT  11.515 40.8625 11.58 40.9975 ;
        RECT  11.325 41.3125 11.39 41.4475 ;
        RECT  11.515 41.3125 11.58 41.4475 ;
        RECT  11.515 41.3125 11.58 41.4475 ;
        RECT  11.705 41.3125 11.77 41.4475 ;
        RECT  11.36 41.1 11.495 41.165 ;
        RECT  11.515 41.5575 11.58 41.6925 ;
        RECT  11.325 41.3125 11.39 41.4475 ;
        RECT  11.705 41.3125 11.77 41.4475 ;
        RECT  11.325 40.8625 11.39 40.9975 ;
        RECT  11.515 40.8625 11.58 40.9975 ;
        RECT  11.835 41.1 12.54 41.165 ;
        RECT  11.835 41.66 12.54 41.725 ;
        RECT  12.22 41.3125 12.285 41.725 ;
        RECT  12.03 40.8625 12.095 40.9975 ;
        RECT  12.22 40.8625 12.285 40.9975 ;
        RECT  12.03 41.3125 12.095 41.4475 ;
        RECT  12.22 41.3125 12.285 41.4475 ;
        RECT  12.22 41.3125 12.285 41.4475 ;
        RECT  12.41 41.3125 12.475 41.4475 ;
        RECT  12.065 41.1 12.2 41.165 ;
        RECT  12.22 41.5575 12.285 41.6925 ;
        RECT  12.03 41.3125 12.095 41.4475 ;
        RECT  12.41 41.3125 12.475 41.4475 ;
        RECT  12.03 40.8625 12.095 40.9975 ;
        RECT  12.22 40.8625 12.285 40.9975 ;
        RECT  11.13 18.7 12.54 18.765 ;
        RECT  11.13 14.2575 12.54 14.3225 ;
        RECT  11.13 14.1275 12.54 14.1925 ;
        RECT  11.6375 14.9225 11.7025 15.1975 ;
        RECT  11.4525 14.9225 11.5175 15.1975 ;
        RECT  11.4475 14.9225 11.5125 15.1975 ;
        RECT  11.2625 14.9225 11.3275 15.1975 ;
        RECT  11.5475 14.465 11.6125 14.74 ;
        RECT  11.3625 14.465 11.4275 14.74 ;
        RECT  11.4475 15.6675 11.5125 16.2225 ;
        RECT  11.2625 15.6675 11.3275 16.2225 ;
        RECT  11.6375 15.6675 11.7025 16.2225 ;
        RECT  11.4525 15.6675 11.5175 16.2225 ;
        RECT  11.4475 17.45 11.5125 18.145 ;
        RECT  11.2625 17.45 11.3275 18.145 ;
        RECT  11.6375 16.48 11.7025 17.175 ;
        RECT  11.4525 16.48 11.5175 17.175 ;
        RECT  11.445 18.4975 11.51 18.6325 ;
        RECT  11.42 14.1275 11.555 14.1925 ;
        RECT  11.8025 14.2575 11.8675 14.3925 ;
        RECT  11.0975 14.2575 11.1625 14.3925 ;
        RECT  11.64 17.04 11.705 17.175 ;
        RECT  11.7225 14.4875 11.7875 14.6225 ;
        RECT  11.2575 17.45 11.3225 17.585 ;
        RECT  11.415 18.3625 11.55 18.4275 ;
        RECT  11.45 18.2925 11.515 18.4275 ;
        RECT  11.45 16.15 11.515 16.285 ;
        RECT  11.3925 15.4625 11.4575 15.5975 ;
        RECT  11.5075 15.2625 11.5725 15.3975 ;
        RECT  11.4 14.2575 11.46 14.3225 ;
        RECT  11.36 14.1275 11.425 14.1925 ;
        RECT  11.7875 14.3225 11.8025 14.3925 ;
        RECT  11.1925 18.4275 11.26 18.765 ;
        RECT  11.1925 18.3625 11.55 18.4275 ;
        RECT  11.695 17.32 11.76 18.5675 ;
        RECT  11.1925 18.7 11.26 18.765 ;
        RECT  11.5475 14.3225 11.6125 14.475 ;
        RECT  11.7225 14.2575 11.7875 14.4875 ;
        RECT  11.4425 18.4975 11.76 18.5675 ;
        RECT  11.45 17.32 11.515 17.5175 ;
        RECT  11.2625 17.32 11.76 17.385 ;
        RECT  11.4525 16.35 11.5175 16.545 ;
        RECT  11.4525 16.35 11.7025 16.415 ;
        RECT  11.4125 14.6525 11.4825 14.98 ;
        RECT  11.095 14.2575 11.87 14.3225 ;
        RECT  11.6375 16.22 11.7025 16.415 ;
        RECT  11.2625 16.2225 11.3275 17.32 ;
        RECT  11.095 18.7 11.87 18.765 ;
        RECT  11.4125 15.4975 11.7025 15.5625 ;
        RECT  11.2625 15.2975 11.5525 15.3625 ;
        RECT  11.2625 15.1925 11.3275 16.06 ;
        RECT  11.6375 15.1975 11.7025 16.06 ;
        RECT  11.095 14.1275 11.87 14.1925 ;
        RECT  12.3425 14.9225 12.4075 15.1975 ;
        RECT  12.1575 14.9225 12.2225 15.1975 ;
        RECT  12.1525 14.9225 12.2175 15.1975 ;
        RECT  11.9675 14.9225 12.0325 15.1975 ;
        RECT  12.2525 14.465 12.3175 14.74 ;
        RECT  12.0675 14.465 12.1325 14.74 ;
        RECT  12.1525 15.6675 12.2175 16.2225 ;
        RECT  11.9675 15.6675 12.0325 16.2225 ;
        RECT  12.3425 15.6675 12.4075 16.2225 ;
        RECT  12.1575 15.6675 12.2225 16.2225 ;
        RECT  12.1525 17.45 12.2175 18.145 ;
        RECT  11.9675 17.45 12.0325 18.145 ;
        RECT  12.3425 16.48 12.4075 17.175 ;
        RECT  12.1575 16.48 12.2225 17.175 ;
        RECT  12.15 18.4975 12.215 18.6325 ;
        RECT  12.125 14.1275 12.26 14.1925 ;
        RECT  12.5075 14.2575 12.5725 14.3925 ;
        RECT  11.8025 14.2575 11.8675 14.3925 ;
        RECT  12.345 17.04 12.41 17.175 ;
        RECT  12.4275 14.4875 12.4925 14.6225 ;
        RECT  11.9625 17.45 12.0275 17.585 ;
        RECT  12.12 18.3625 12.255 18.4275 ;
        RECT  12.155 18.2925 12.22 18.4275 ;
        RECT  12.155 16.15 12.22 16.285 ;
        RECT  12.0975 15.4625 12.1625 15.5975 ;
        RECT  12.2125 15.2625 12.2775 15.3975 ;
        RECT  12.105 14.2575 12.165 14.3225 ;
        RECT  12.065 14.1275 12.13 14.1925 ;
        RECT  12.4925 14.3225 12.5075 14.3925 ;
        RECT  11.8975 18.4275 11.965 18.765 ;
        RECT  11.8975 18.3625 12.255 18.4275 ;
        RECT  12.4 17.32 12.465 18.5675 ;
        RECT  11.8975 18.7 11.965 18.765 ;
        RECT  12.2525 14.3225 12.3175 14.475 ;
        RECT  12.4275 14.2575 12.4925 14.4875 ;
        RECT  12.1475 18.4975 12.465 18.5675 ;
        RECT  12.155 17.32 12.22 17.5175 ;
        RECT  11.9675 17.32 12.465 17.385 ;
        RECT  12.1575 16.35 12.2225 16.545 ;
        RECT  12.1575 16.35 12.4075 16.415 ;
        RECT  12.1175 14.6525 12.1875 14.98 ;
        RECT  11.8 14.2575 12.575 14.3225 ;
        RECT  12.3425 16.22 12.4075 16.415 ;
        RECT  11.9675 16.2225 12.0325 17.32 ;
        RECT  11.8 18.7 12.575 18.765 ;
        RECT  12.1175 15.4975 12.4075 15.5625 ;
        RECT  11.9675 15.2975 12.2575 15.3625 ;
        RECT  11.9675 15.1925 12.0325 16.06 ;
        RECT  12.3425 15.1975 12.4075 16.06 ;
        RECT  11.8 14.1275 12.575 14.1925 ;
        RECT  11.13 10.1025 12.54 10.1675 ;
        RECT  11.13 10.2325 12.54 10.2975 ;
        RECT  11.13 11.035 12.54 11.1 ;
        RECT  11.55 13.4975 11.615 13.6325 ;
        RECT  11.175 13.4975 11.24 13.6325 ;
        RECT  11.175 11.57 11.24 11.705 ;
        RECT  11.55 11.57 11.615 11.705 ;
        RECT  11.55 12.7025 11.615 13.1175 ;
        RECT  11.175 12.7025 11.24 13.1175 ;
        RECT  11.175 12.085 11.24 12.5 ;
        RECT  11.55 12.085 11.615 12.5 ;
        RECT  11.36 10.515 11.425 10.93 ;
        RECT  11.175 10.515 11.24 10.93 ;
        RECT  11.515 10.515 11.58 10.93 ;
        RECT  11.7 10.515 11.765 10.93 ;
        RECT  11.36 11.205 11.425 11.34 ;
        RECT  11.175 11.205 11.24 11.34 ;
        RECT  11.515 11.205 11.58 11.34 ;
        RECT  11.7 11.205 11.765 11.34 ;
        RECT  11.3375 9.97 11.4725 10.035 ;
        RECT  11.4125 11.925 11.4775 12.06 ;
        RECT  11.8025 11.57 11.8675 11.705 ;
        RECT  11.715 11.57 11.78 11.705 ;
        RECT  11.0975 12.5325 11.1625 12.6675 ;
        RECT  11.8025 11.0 11.8675 11.135 ;
        RECT  11.0975 11.0 11.1625 11.135 ;
        RECT  11.5175 11.205 11.5825 11.34 ;
        RECT  11.8025 13.4975 11.8675 13.6325 ;
        RECT  11.7175 13.4975 11.7825 13.6325 ;
        RECT  11.5175 10.795 11.5825 10.93 ;
        RECT  11.3775 10.795 11.4425 10.93 ;
        RECT  11.4 10.3825 11.535 10.4475 ;
        RECT  11.2325 9.9725 11.3675 10.0375 ;
        RECT  11.5725 10.1025 11.7075 10.1675 ;
        RECT  11.8025 11.205 11.8675 11.34 ;
        RECT  11.0975 11.205 11.1625 11.34 ;
        RECT  11.235 10.2325 11.37 10.2975 ;
        RECT  11.3775 13.175 11.4425 13.31 ;
        RECT  11.5475 11.57 11.6125 11.705 ;
        RECT  11.2375 12.485 11.3025 12.62 ;
        RECT  11.3775 11.205 11.4425 11.34 ;
        RECT  11.315 13.175 11.38 13.31 ;
        RECT  11.0975 11.57 11.1625 11.705 ;
        RECT  11.5475 12.085 11.6125 12.22 ;
        RECT  11.2825 13.7075 11.3475 13.8425 ;
        RECT  11.0975 13.4975 11.1625 13.6325 ;
        RECT  11.7825 13.4975 11.8025 13.6325 ;
        RECT  11.78 11.57 11.8025 11.705 ;
        RECT  11.45 11.0375 11.5075 11.0975 ;
        RECT  11.425 10.1025 11.4975 10.1675 ;
        RECT  11.4275 10.2325 11.4975 10.2975 ;
        RECT  11.1575 13.4975 11.17 13.6325 ;
        RECT  11.1625 12.5325 11.305 12.6675 ;
        RECT  11.095 11.035 11.87 11.1 ;
        RECT  11.4325 10.2975 11.4975 10.4475 ;
        RECT  11.76 11.205 11.8025 11.34 ;
        RECT  11.7 10.2975 11.765 10.515 ;
        RECT  11.175 10.2975 11.24 10.515 ;
        RECT  11.095 10.2325 11.87 10.2975 ;
        RECT  11.095 10.1025 11.87 10.1675 ;
        RECT  11.1575 11.205 11.17 11.34 ;
        RECT  11.225 12.485 11.24 12.62 ;
        RECT  11.1575 11.57 11.17 11.705 ;
        RECT  11.175 12.5 11.24 12.7025 ;
        RECT  11.55 13.6325 11.615 13.7075 ;
        RECT  11.4125 11.4125 11.575 11.4775 ;
        RECT  11.165 13.4975 11.175 13.6325 ;
        RECT  11.165 11.57 11.175 11.705 ;
        RECT  11.51 11.2875 11.575 11.4125 ;
        RECT  11.4125 11.4125 11.4775 12.01 ;
        RECT  11.55 13.1175 11.615 13.4975 ;
        RECT  11.28 13.7075 11.615 13.7725 ;
        RECT  11.165 11.205 11.175 11.34 ;
        RECT  12.255 13.4975 12.32 13.6325 ;
        RECT  11.88 13.4975 11.945 13.6325 ;
        RECT  11.88 11.57 11.945 11.705 ;
        RECT  12.255 11.57 12.32 11.705 ;
        RECT  12.255 12.7025 12.32 13.1175 ;
        RECT  11.88 12.7025 11.945 13.1175 ;
        RECT  11.88 12.085 11.945 12.5 ;
        RECT  12.255 12.085 12.32 12.5 ;
        RECT  12.065 10.515 12.13 10.93 ;
        RECT  11.88 10.515 11.945 10.93 ;
        RECT  12.22 10.515 12.285 10.93 ;
        RECT  12.405 10.515 12.47 10.93 ;
        RECT  12.065 11.205 12.13 11.34 ;
        RECT  11.88 11.205 11.945 11.34 ;
        RECT  12.22 11.205 12.285 11.34 ;
        RECT  12.405 11.205 12.47 11.34 ;
        RECT  12.0425 9.97 12.1775 10.035 ;
        RECT  12.1175 11.925 12.1825 12.06 ;
        RECT  12.5075 11.57 12.5725 11.705 ;
        RECT  12.42 11.57 12.485 11.705 ;
        RECT  11.8025 12.5325 11.8675 12.6675 ;
        RECT  12.5075 11.0 12.5725 11.135 ;
        RECT  11.8025 11.0 11.8675 11.135 ;
        RECT  12.2225 11.205 12.2875 11.34 ;
        RECT  12.5075 13.4975 12.5725 13.6325 ;
        RECT  12.4225 13.4975 12.4875 13.6325 ;
        RECT  12.2225 10.795 12.2875 10.93 ;
        RECT  12.0825 10.795 12.1475 10.93 ;
        RECT  12.105 10.3825 12.24 10.4475 ;
        RECT  11.9375 9.9725 12.0725 10.0375 ;
        RECT  12.2775 10.1025 12.4125 10.1675 ;
        RECT  12.5075 11.205 12.5725 11.34 ;
        RECT  11.8025 11.205 11.8675 11.34 ;
        RECT  11.94 10.2325 12.075 10.2975 ;
        RECT  12.0825 13.175 12.1475 13.31 ;
        RECT  12.2525 11.57 12.3175 11.705 ;
        RECT  11.9425 12.485 12.0075 12.62 ;
        RECT  12.0825 11.205 12.1475 11.34 ;
        RECT  12.02 13.175 12.085 13.31 ;
        RECT  11.8025 11.57 11.8675 11.705 ;
        RECT  12.2525 12.085 12.3175 12.22 ;
        RECT  11.9875 13.7075 12.0525 13.8425 ;
        RECT  11.8025 13.4975 11.8675 13.6325 ;
        RECT  12.4875 13.4975 12.5075 13.6325 ;
        RECT  12.485 11.57 12.5075 11.705 ;
        RECT  12.155 11.0375 12.2125 11.0975 ;
        RECT  12.13 10.1025 12.2025 10.1675 ;
        RECT  12.1325 10.2325 12.2025 10.2975 ;
        RECT  11.8625 13.4975 11.875 13.6325 ;
        RECT  11.8675 12.5325 12.01 12.6675 ;
        RECT  11.8 11.035 12.575 11.1 ;
        RECT  12.1375 10.2975 12.2025 10.4475 ;
        RECT  12.465 11.205 12.5075 11.34 ;
        RECT  12.405 10.2975 12.47 10.515 ;
        RECT  11.88 10.2975 11.945 10.515 ;
        RECT  11.8 10.2325 12.575 10.2975 ;
        RECT  11.8 10.1025 12.575 10.1675 ;
        RECT  11.8625 11.205 11.875 11.34 ;
        RECT  11.93 12.485 11.945 12.62 ;
        RECT  11.8625 11.57 11.875 11.705 ;
        RECT  11.88 12.5 11.945 12.7025 ;
        RECT  12.255 13.6325 12.32 13.7075 ;
        RECT  12.1175 11.4125 12.28 11.4775 ;
        RECT  11.87 13.4975 11.88 13.6325 ;
        RECT  11.87 11.57 11.88 11.705 ;
        RECT  12.215 11.2875 12.28 11.4125 ;
        RECT  12.1175 11.4125 12.1825 12.01 ;
        RECT  12.255 13.1175 12.32 13.4975 ;
        RECT  11.985 13.7075 12.32 13.7725 ;
        RECT  11.87 11.205 11.88 11.34 ;
        RECT  11.13 3.5675 12.54 3.6325 ;
        RECT  11.13 9.565 12.54 9.63 ;
        RECT  11.67 6.085 11.735 6.22 ;
        RECT  11.485 6.085 11.55 6.22 ;
        RECT  11.67 4.85 11.735 4.985 ;
        RECT  11.485 4.85 11.55 4.985 ;
        RECT  11.48 6.085 11.545 6.22 ;
        RECT  11.295 6.085 11.36 6.22 ;
        RECT  11.48 9.045 11.545 9.18 ;
        RECT  11.295 9.045 11.36 9.18 ;
        RECT  11.48 4.85 11.545 4.985 ;
        RECT  11.295 4.85 11.36 4.985 ;
        RECT  11.67 9.045 11.735 9.18 ;
        RECT  11.485 9.045 11.55 9.18 ;
        RECT  11.48 4.315 11.545 4.45 ;
        RECT  11.295 4.315 11.36 4.45 ;
        RECT  11.62 7.275 11.685 7.41 ;
        RECT  11.435 7.275 11.5 7.41 ;
        RECT  11.67 7.81 11.735 7.945 ;
        RECT  11.485 7.81 11.55 7.945 ;
        RECT  11.48 7.81 11.545 7.945 ;
        RECT  11.295 7.81 11.36 7.945 ;
        RECT  11.67 8.235 11.735 8.37 ;
        RECT  11.485 8.235 11.55 8.37 ;
        RECT  11.67 5.275 11.735 5.41 ;
        RECT  11.485 5.275 11.55 5.41 ;
        RECT  11.67 8.62 11.735 8.755 ;
        RECT  11.485 8.62 11.55 8.755 ;
        RECT  11.48 8.62 11.545 8.755 ;
        RECT  11.295 8.62 11.36 8.755 ;
        RECT  11.48 5.275 11.545 5.41 ;
        RECT  11.295 5.275 11.36 5.41 ;
        RECT  11.48 8.235 11.545 8.37 ;
        RECT  11.295 8.235 11.36 8.37 ;
        RECT  11.48 5.66 11.545 5.795 ;
        RECT  11.295 5.66 11.36 5.795 ;
        RECT  11.67 5.66 11.735 5.795 ;
        RECT  11.485 5.66 11.55 5.795 ;
        RECT  11.48 3.89 11.545 4.025 ;
        RECT  11.295 3.89 11.36 4.025 ;
        RECT  11.555 6.865 11.62 7.0 ;
        RECT  11.37 6.865 11.435 7.0 ;
        RECT  11.3575 3.6 11.4925 3.665 ;
        RECT  11.295 9.0975 11.36 9.2325 ;
        RECT  11.185 7.2825 11.25 7.4175 ;
        RECT  11.295 6.3825 11.36 6.5175 ;
        RECT  11.7175 6.8575 11.7825 6.9925 ;
        RECT  11.295 9.4625 11.36 9.5975 ;
        RECT  11.8025 3.92 11.8675 4.055 ;
        RECT  11.66 8.0025 11.725 8.1375 ;
        RECT  11.6625 6.395 11.7275 6.53 ;
        RECT  11.6625 4.9975 11.7275 5.1325 ;
        RECT  11.0975 3.78 11.1625 3.915 ;
        RECT  11.6725 3.8975 11.7375 4.0325 ;
        RECT  11.6725 5.5075 11.8075 5.5725 ;
        RECT  11.7125 4.4225 11.7775 4.5575 ;
        RECT  11.6725 8.4675 11.8075 8.5325 ;
        RECT  11.62 9.355 11.685 9.49 ;
        RECT  11.54 5.885 11.605 6.02 ;
        RECT  11.53 8.845 11.595 8.98 ;
        RECT  11.2975 7.155 11.4325 7.22 ;
        RECT  11.8025 6.8575 11.8675 6.9925 ;
        RECT  11.1875 4.15 11.3225 4.215 ;
        RECT  11.2975 5.6625 11.3625 5.7975 ;
        RECT  11.6625 9.355 11.7275 9.49 ;
        RECT  11.485 8.845 11.55 8.98 ;
        RECT  11.8025 8.4325 11.8675 8.5675 ;
        RECT  11.8025 3.73 11.8675 3.865 ;
        RECT  11.6625 6.395 11.7275 6.53 ;
        RECT  11.8025 5.4725 11.8675 5.6075 ;
        RECT  11.2975 5.2725 11.3625 5.4075 ;
        RECT  11.485 5.2725 11.55 5.4075 ;
        RECT  11.485 5.885 11.55 6.02 ;
        RECT  11.295 8.2325 11.36 8.3675 ;
        RECT  11.485 8.2325 11.55 8.3675 ;
        RECT  11.095 3.6 11.87 3.665 ;
        RECT  11.165 6.67 11.23 9.565 ;
        RECT  11.67 9.18 11.735 9.49 ;
        RECT  11.295 8.755 11.36 9.045 ;
        RECT  11.295 7.945 11.36 8.235 ;
        RECT  11.435 9.5675 11.5075 9.63 ;
        RECT  11.48 9.18 11.55 9.565 ;
        RECT  11.48 7.945 11.55 8.235 ;
        RECT  11.48 8.465 11.55 8.6225 ;
        RECT  11.67 8.755 11.735 9.045 ;
        RECT  11.67 7.945 11.735 8.235 ;
        RECT  11.48 8.465 11.865 8.535 ;
        RECT  11.095 9.565 11.87 9.63 ;
        RECT  11.095 7.575 11.87 7.64 ;
        RECT  11.165 4.68 11.23 6.605 ;
        RECT  11.67 6.22 11.735 6.53 ;
        RECT  11.295 5.795 11.36 6.085 ;
        RECT  11.37 6.96 11.435 7.41 ;
        RECT  11.48 6.22 11.55 6.605 ;
        RECT  11.48 5.505 11.55 5.6625 ;
        RECT  11.295 6.5175 11.36 6.605 ;
        RECT  11.67 5.795 11.735 6.085 ;
        RECT  11.555 6.735 11.8 6.8 ;
        RECT  11.7175 6.735 11.8 6.8575 ;
        RECT  11.7375 6.8575 11.805 6.9925 ;
        RECT  11.095 6.605 11.87 6.67 ;
        RECT  11.295 4.985 11.36 5.275 ;
        RECT  11.48 4.4475 11.545 4.615 ;
        RECT  11.545 3.955 11.8025 4.025 ;
        RECT  11.295 3.89 11.36 4.315 ;
        RECT  11.48 4.985 11.55 5.275 ;
        RECT  11.1875 4.145 11.36 4.22 ;
        RECT  11.67 4.985 11.735 5.275 ;
        RECT  11.6725 3.825 11.7375 3.8975 ;
        RECT  11.48 5.505 11.865 5.575 ;
        RECT  11.7125 4.535 11.7775 4.65 ;
        RECT  11.095 3.76 11.87 3.825 ;
        RECT  11.095 4.615 11.87 4.68 ;
        RECT  11.235 3.605 11.3 3.6625 ;
        RECT  11.8025 3.845 11.8675 3.9675 ;
        RECT  11.62 7.4075 11.685 7.575 ;
        RECT  11.555 6.8 11.6225 6.9025 ;
        RECT  11.935 6.085 12.0 6.22 ;
        RECT  12.12 6.085 12.185 6.22 ;
        RECT  11.935 4.85 12.0 4.985 ;
        RECT  12.12 4.85 12.185 4.985 ;
        RECT  12.125 6.085 12.19 6.22 ;
        RECT  12.31 6.085 12.375 6.22 ;
        RECT  12.125 9.045 12.19 9.18 ;
        RECT  12.31 9.045 12.375 9.18 ;
        RECT  12.125 4.85 12.19 4.985 ;
        RECT  12.31 4.85 12.375 4.985 ;
        RECT  11.935 9.045 12.0 9.18 ;
        RECT  12.12 9.045 12.185 9.18 ;
        RECT  12.125 4.315 12.19 4.45 ;
        RECT  12.31 4.315 12.375 4.45 ;
        RECT  11.985 7.275 12.05 7.41 ;
        RECT  12.17 7.275 12.235 7.41 ;
        RECT  11.935 7.81 12.0 7.945 ;
        RECT  12.12 7.81 12.185 7.945 ;
        RECT  12.125 7.81 12.19 7.945 ;
        RECT  12.31 7.81 12.375 7.945 ;
        RECT  11.935 8.235 12.0 8.37 ;
        RECT  12.12 8.235 12.185 8.37 ;
        RECT  11.935 5.275 12.0 5.41 ;
        RECT  12.12 5.275 12.185 5.41 ;
        RECT  11.935 8.62 12.0 8.755 ;
        RECT  12.12 8.62 12.185 8.755 ;
        RECT  12.125 8.62 12.19 8.755 ;
        RECT  12.31 8.62 12.375 8.755 ;
        RECT  12.125 5.275 12.19 5.41 ;
        RECT  12.31 5.275 12.375 5.41 ;
        RECT  12.125 8.235 12.19 8.37 ;
        RECT  12.31 8.235 12.375 8.37 ;
        RECT  12.125 5.66 12.19 5.795 ;
        RECT  12.31 5.66 12.375 5.795 ;
        RECT  11.935 5.66 12.0 5.795 ;
        RECT  12.12 5.66 12.185 5.795 ;
        RECT  12.125 3.89 12.19 4.025 ;
        RECT  12.31 3.89 12.375 4.025 ;
        RECT  12.05 6.865 12.115 7.0 ;
        RECT  12.235 6.865 12.3 7.0 ;
        RECT  12.1775 3.6 12.3125 3.665 ;
        RECT  12.31 9.0975 12.375 9.2325 ;
        RECT  12.42 7.2825 12.485 7.4175 ;
        RECT  12.31 6.3825 12.375 6.5175 ;
        RECT  11.8875 6.8575 11.9525 6.9925 ;
        RECT  12.31 9.4625 12.375 9.5975 ;
        RECT  11.8025 3.92 11.8675 4.055 ;
        RECT  11.945 8.0025 12.01 8.1375 ;
        RECT  11.9425 6.395 12.0075 6.53 ;
        RECT  11.9425 4.9975 12.0075 5.1325 ;
        RECT  12.5075 3.78 12.5725 3.915 ;
        RECT  11.9325 3.8975 11.9975 4.0325 ;
        RECT  11.8625 5.5075 11.9975 5.5725 ;
        RECT  11.8925 4.4225 11.9575 4.5575 ;
        RECT  11.8625 8.4675 11.9975 8.5325 ;
        RECT  11.985 9.355 12.05 9.49 ;
        RECT  12.065 5.885 12.13 6.02 ;
        RECT  12.075 8.845 12.14 8.98 ;
        RECT  12.2375 7.155 12.3725 7.22 ;
        RECT  11.8025 6.8575 11.8675 6.9925 ;
        RECT  12.3475 4.15 12.4825 4.215 ;
        RECT  12.3075 5.6625 12.3725 5.7975 ;
        RECT  11.9425 9.355 12.0075 9.49 ;
        RECT  12.12 8.845 12.185 8.98 ;
        RECT  11.8025 8.4325 11.8675 8.5675 ;
        RECT  11.8025 3.73 11.8675 3.865 ;
        RECT  11.9425 6.395 12.0075 6.53 ;
        RECT  11.8025 5.4725 11.8675 5.6075 ;
        RECT  12.3075 5.2725 12.3725 5.4075 ;
        RECT  12.12 5.2725 12.185 5.4075 ;
        RECT  12.12 5.885 12.185 6.02 ;
        RECT  12.31 8.2325 12.375 8.3675 ;
        RECT  12.12 8.2325 12.185 8.3675 ;
        RECT  11.8 3.6 12.575 3.665 ;
        RECT  12.44 6.67 12.505 9.565 ;
        RECT  11.935 9.18 12.0 9.49 ;
        RECT  12.31 8.755 12.375 9.045 ;
        RECT  12.31 7.945 12.375 8.235 ;
        RECT  12.1625 9.5675 12.235 9.63 ;
        RECT  12.12 9.18 12.19 9.565 ;
        RECT  12.12 7.945 12.19 8.235 ;
        RECT  12.12 8.465 12.19 8.6225 ;
        RECT  11.935 8.755 12.0 9.045 ;
        RECT  11.935 7.945 12.0 8.235 ;
        RECT  11.805 8.465 12.19 8.535 ;
        RECT  11.8 9.565 12.575 9.63 ;
        RECT  11.8 7.575 12.575 7.64 ;
        RECT  12.44 4.68 12.505 6.605 ;
        RECT  11.935 6.22 12.0 6.53 ;
        RECT  12.31 5.795 12.375 6.085 ;
        RECT  12.235 6.96 12.3 7.41 ;
        RECT  12.12 6.22 12.19 6.605 ;
        RECT  12.12 5.505 12.19 5.6625 ;
        RECT  12.31 6.5175 12.375 6.605 ;
        RECT  11.935 5.795 12.0 6.085 ;
        RECT  11.87 6.735 12.115 6.8 ;
        RECT  11.87 6.735 11.9525 6.8575 ;
        RECT  11.865 6.8575 11.9325 6.9925 ;
        RECT  11.8 6.605 12.575 6.67 ;
        RECT  12.31 4.985 12.375 5.275 ;
        RECT  12.125 4.4475 12.19 4.615 ;
        RECT  11.8675 3.955 12.125 4.025 ;
        RECT  12.31 3.89 12.375 4.315 ;
        RECT  12.12 4.985 12.19 5.275 ;
        RECT  12.31 4.145 12.4825 4.22 ;
        RECT  11.935 4.985 12.0 5.275 ;
        RECT  11.9325 3.825 11.9975 3.8975 ;
        RECT  11.805 5.505 12.19 5.575 ;
        RECT  11.8925 4.535 11.9575 4.65 ;
        RECT  11.8 3.76 12.575 3.825 ;
        RECT  11.8 4.615 12.575 4.68 ;
        RECT  12.37 3.605 12.435 3.6625 ;
        RECT  11.8025 3.845 11.8675 3.9675 ;
        RECT  11.985 7.4075 12.05 7.575 ;
        RECT  12.0475 6.8 12.115 6.9025 ;
        RECT  11.13 2.9625 12.54 3.0275 ;
        RECT  11.13 1.415 12.54 1.48 ;
        RECT  11.13 1.545 12.54 1.61 ;
        RECT  11.485 5.44 11.55 5.575 ;
        RECT  11.3 5.44 11.365 5.575 ;
        RECT  11.485 5.955 11.55 6.09 ;
        RECT  11.3 5.955 11.365 6.09 ;
        RECT  11.6125 4.045 11.6775 4.18 ;
        RECT  11.2375 4.045 11.3025 4.18 ;
        RECT  11.6125 4.6725 11.6775 5.0875 ;
        RECT  11.2375 4.6725 11.3025 5.0875 ;
        RECT  11.6275 4.3125 11.7625 4.3775 ;
        RECT  11.65 5.9625 11.715 6.0975 ;
        RECT  11.415 5.18 11.55 5.245 ;
        RECT  11.57 3.8925 11.705 3.9575 ;
        RECT  11.8025 3.8925 11.8675 4.0275 ;
        RECT  11.1875 5.31 11.3225 5.375 ;
        RECT  11.2925 3.7625 11.4275 3.8275 ;
        RECT  11.5475 5.82 11.6825 5.885 ;
        RECT  11.8025 5.9525 11.8675 6.0875 ;
        RECT  11.5475 5.78 11.6825 5.845 ;
        RECT  11.57 5.18 11.705 5.245 ;
        RECT  11.275 5.7625 11.34 5.8975 ;
        RECT  11.4825 5.485 11.5475 5.62 ;
        RECT  11.455 3.7625 11.5125 3.8275 ;
        RECT  11.4075 5.31 11.47 5.375 ;
        RECT  11.3 5.57 11.365 6.09 ;
        RECT  11.2375 4.1575 11.3025 4.6725 ;
        RECT  11.5475 4.3125 11.6825 4.3775 ;
        RECT  11.13 3.7625 11.87 3.8275 ;
        RECT  11.13 3.8925 11.87 3.9575 ;
        RECT  11.6125 3.9575 11.6775 4.045 ;
        RECT  11.505 5.9525 11.8025 6.0875 ;
        RECT  11.13 5.31 11.87 5.375 ;
        RECT  11.13 5.18 11.87 5.245 ;
        RECT  11.6125 5.0875 11.6775 5.18 ;
        RECT  11.2725 5.18 11.3375 5.245 ;
        RECT  11.2375 4.045 11.3025 4.18 ;
        RECT  12.12 5.44 12.185 5.575 ;
        RECT  12.305 5.44 12.37 5.575 ;
        RECT  12.12 5.955 12.185 6.09 ;
        RECT  12.305 5.955 12.37 6.09 ;
        RECT  11.9925 4.045 12.0575 4.18 ;
        RECT  12.3675 4.045 12.4325 4.18 ;
        RECT  11.9925 4.6725 12.0575 5.0875 ;
        RECT  12.3675 4.6725 12.4325 5.0875 ;
        RECT  11.9075 4.3125 12.0425 4.3775 ;
        RECT  11.955 5.9625 12.02 6.0975 ;
        RECT  12.12 5.18 12.255 5.245 ;
        RECT  11.965 3.8925 12.1 3.9575 ;
        RECT  11.8025 3.8925 11.8675 4.0275 ;
        RECT  12.3475 5.31 12.4825 5.375 ;
        RECT  12.2425 3.7625 12.3775 3.8275 ;
        RECT  11.9875 5.82 12.1225 5.885 ;
        RECT  11.8025 5.9525 11.8675 6.0875 ;
        RECT  11.9875 5.78 12.1225 5.845 ;
        RECT  11.965 5.18 12.1 5.245 ;
        RECT  12.33 5.7625 12.395 5.8975 ;
        RECT  12.1225 5.485 12.1875 5.62 ;
        RECT  12.1575 3.7625 12.215 3.8275 ;
        RECT  12.2 5.31 12.2625 5.375 ;
        RECT  12.305 5.57 12.37 6.09 ;
        RECT  12.3675 4.1575 12.4325 4.6725 ;
        RECT  11.9875 4.3125 12.1225 4.3775 ;
        RECT  11.8 3.7625 12.54 3.8275 ;
        RECT  11.8 3.8925 12.54 3.9575 ;
        RECT  11.9925 3.9575 12.0575 4.045 ;
        RECT  11.8675 5.9525 12.165 6.0875 ;
        RECT  11.8 5.31 12.54 5.375 ;
        RECT  11.8 5.18 12.54 5.245 ;
        RECT  11.9925 5.0875 12.0575 5.18 ;
        RECT  12.3325 5.18 12.3975 5.245 ;
        RECT  12.3675 4.045 12.4325 4.18 ;
        RECT  4.97 19.4925 5.035 19.5575 ;
        RECT  4.97 20.9225 5.035 20.9875 ;
        RECT  4.97 22.1825 5.035 22.2475 ;
        RECT  4.97 23.6125 5.035 23.6775 ;
        RECT  4.97 24.8725 5.035 24.9375 ;
        RECT  4.97 26.3025 5.035 26.3675 ;
        RECT  4.97 27.5625 5.035 27.6275 ;
        RECT  4.97 28.9925 5.035 29.0575 ;
        RECT  4.97 30.2525 5.035 30.3175 ;
        RECT  4.97 31.6825 5.035 31.7475 ;
        RECT  4.97 32.9425 5.035 33.0075 ;
        RECT  4.97 34.3725 5.035 34.4375 ;
        RECT  4.97 35.6325 5.035 35.6975 ;
        RECT  4.97 37.0625 5.035 37.1275 ;
        RECT  4.97 38.3225 5.035 38.3875 ;
        RECT  4.97 39.7525 5.035 39.8175 ;
        RECT  2.82 8.73 4.22 8.795 ;
        RECT  2.995 10.165 4.22 10.23 ;
        RECT  3.17 11.42 4.22 11.485 ;
        RECT  3.345 12.855 4.22 12.92 ;
        RECT  3.52 14.11 4.22 14.175 ;
        RECT  3.695 15.545 4.22 15.61 ;
        RECT  3.87 16.8 4.22 16.865 ;
        RECT  4.045 18.235 4.22 18.3 ;
        RECT  2.82 19.805 4.22 19.87 ;
        RECT  3.52 19.275 4.22 19.34 ;
        RECT  2.82 20.61 4.22 20.675 ;
        RECT  3.695 21.14 4.22 21.205 ;
        RECT  2.82 22.495 4.22 22.56 ;
        RECT  3.87 21.965 4.22 22.03 ;
        RECT  2.82 23.3 4.22 23.365 ;
        RECT  4.045 23.83 4.22 23.895 ;
        RECT  2.995 25.185 4.22 25.25 ;
        RECT  3.52 24.655 4.22 24.72 ;
        RECT  2.995 25.99 4.22 26.055 ;
        RECT  3.695 26.52 4.22 26.585 ;
        RECT  2.995 27.875 4.22 27.94 ;
        RECT  3.87 27.345 4.22 27.41 ;
        RECT  2.995 28.68 4.22 28.745 ;
        RECT  4.045 29.21 4.22 29.275 ;
        RECT  3.17 30.565 4.22 30.63 ;
        RECT  3.52 30.035 4.22 30.1 ;
        RECT  3.17 31.37 4.22 31.435 ;
        RECT  3.695 31.9 4.22 31.965 ;
        RECT  3.17 33.255 4.22 33.32 ;
        RECT  3.87 32.725 4.22 32.79 ;
        RECT  3.17 34.06 4.22 34.125 ;
        RECT  4.045 34.59 4.22 34.655 ;
        RECT  3.345 35.945 4.22 36.01 ;
        RECT  3.52 35.415 4.22 35.48 ;
        RECT  3.345 36.75 4.22 36.815 ;
        RECT  3.695 37.28 4.22 37.345 ;
        RECT  3.345 38.635 4.22 38.7 ;
        RECT  3.87 38.105 4.22 38.17 ;
        RECT  3.345 39.44 4.22 39.505 ;
        RECT  4.045 39.97 4.22 40.035 ;
        RECT  4.715 8.7325 4.78 8.7975 ;
        RECT  4.715 10.1625 4.78 10.2275 ;
        RECT  4.715 11.4225 4.78 11.4875 ;
        RECT  4.715 12.8525 4.78 12.9175 ;
        RECT  6.62 8.73 6.685 9.3175 ;
        RECT  6.16 9.2525 6.685 9.3175 ;
        RECT  7.175 8.73 7.595 8.795 ;
        RECT  6.51 9.4475 7.245 9.5125 ;
        RECT  6.335 8.1025 7.245 8.1675 ;
        RECT  6.62 9.6425 6.685 10.23 ;
        RECT  5.985 9.6425 6.685 9.7075 ;
        RECT  7.175 10.165 7.42 10.23 ;
        RECT  6.51 9.4475 7.245 9.5125 ;
        RECT  6.335 10.7925 7.245 10.8575 ;
        RECT  5.53 9.045 6.23 9.11 ;
        RECT  5.53 8.515 6.055 8.58 ;
        RECT  5.53 9.85 5.88 9.915 ;
        RECT  5.53 10.38 6.055 10.445 ;
        RECT  5.53 11.735 6.23 11.8 ;
        RECT  5.53 11.205 5.705 11.27 ;
        RECT  5.53 12.54 5.88 12.605 ;
        RECT  5.53 12.54 7.595 12.605 ;
        RECT  5.53 13.07 5.705 13.135 ;
        RECT  5.53 13.07 7.42 13.135 ;
        RECT  5.53 8.1025 6.405 8.1675 ;
        RECT  5.53 9.4475 6.58 9.5125 ;
        RECT  5.53 10.7925 6.405 10.8575 ;
        RECT  5.53 12.1375 6.58 12.2025 ;
        RECT  5.53 13.4825 6.405 13.5475 ;
        RECT  6.34 13.305 6.405 13.4825 ;
        RECT  6.685 8.1025 7.245 8.1675 ;
        RECT  6.685 6.7575 7.245 6.8225 ;
        RECT  6.7525 6.8225 6.8175 7.0725 ;
        RECT  6.7525 7.9675 6.8175 8.1025 ;
        RECT  7.1125 8.0325 7.1775 8.1025 ;
        RECT  7.1125 6.8225 7.1775 6.9375 ;
        RECT  6.9225 6.9375 6.9875 8.0 ;
        RECT  7.21 7.475 7.245 7.54 ;
        RECT  6.685 7.475 6.9225 7.54 ;
        RECT  7.1125 7.7625 7.1775 7.8975 ;
        RECT  6.9225 7.7625 6.9875 7.8975 ;
        RECT  7.1125 6.9375 7.1775 7.0725 ;
        RECT  6.9225 6.9375 6.9875 7.0725 ;
        RECT  6.7525 6.9375 6.8175 7.0725 ;
        RECT  6.7525 7.8975 6.8175 8.0325 ;
        RECT  7.075 7.475 7.21 7.54 ;
        RECT  6.685 10.7925 7.245 10.8575 ;
        RECT  6.685 12.1375 7.245 12.2025 ;
        RECT  6.7525 11.8875 6.8175 12.1375 ;
        RECT  6.7525 10.8575 6.8175 10.9925 ;
        RECT  7.1125 10.8575 7.1775 10.9275 ;
        RECT  7.1125 12.0225 7.1775 12.1375 ;
        RECT  6.9225 10.96 6.9875 12.0225 ;
        RECT  7.21 11.42 7.245 11.485 ;
        RECT  6.685 11.42 6.9225 11.485 ;
        RECT  7.1125 10.9925 7.1775 11.1275 ;
        RECT  6.9225 10.9925 6.9875 11.1275 ;
        RECT  7.1125 11.5975 7.1775 11.7325 ;
        RECT  6.9225 11.5975 6.9875 11.7325 ;
        RECT  6.7525 11.7525 6.8175 11.8875 ;
        RECT  6.7525 10.7925 6.8175 10.9275 ;
        RECT  7.075 11.345 7.21 11.41 ;
        RECT  4.22 8.1025 4.78 8.1675 ;
        RECT  4.22 6.7575 4.78 6.8225 ;
        RECT  4.2875 6.8225 4.3525 7.0725 ;
        RECT  4.2875 7.9675 4.3525 8.1025 ;
        RECT  4.6475 8.0325 4.7125 8.1025 ;
        RECT  4.6475 6.8225 4.7125 6.9375 ;
        RECT  4.4575 6.9375 4.5225 8.0 ;
        RECT  4.745 7.475 4.78 7.54 ;
        RECT  4.22 7.475 4.4575 7.54 ;
        RECT  4.6475 7.7625 4.7125 7.8975 ;
        RECT  4.4575 7.7625 4.5225 7.8975 ;
        RECT  4.6475 6.9375 4.7125 7.0725 ;
        RECT  4.4575 6.9375 4.5225 7.0725 ;
        RECT  4.2875 6.9375 4.3525 7.0725 ;
        RECT  4.2875 7.8975 4.3525 8.0325 ;
        RECT  4.61 7.475 4.745 7.54 ;
        RECT  4.22 10.7925 4.78 10.8575 ;
        RECT  4.22 12.1375 4.78 12.2025 ;
        RECT  4.2875 11.8875 4.3525 12.1375 ;
        RECT  4.2875 10.8575 4.3525 10.9925 ;
        RECT  4.6475 10.8575 4.7125 10.9275 ;
        RECT  4.6475 12.0225 4.7125 12.1375 ;
        RECT  4.4575 10.96 4.5225 12.0225 ;
        RECT  4.745 11.42 4.78 11.485 ;
        RECT  4.22 11.42 4.4575 11.485 ;
        RECT  4.6475 10.9925 4.7125 11.1275 ;
        RECT  4.4575 10.9925 4.5225 11.1275 ;
        RECT  4.6475 11.5975 4.7125 11.7325 ;
        RECT  4.4575 11.5975 4.5225 11.7325 ;
        RECT  4.2875 11.7525 4.3525 11.8875 ;
        RECT  4.2875 10.7925 4.3525 10.9275 ;
        RECT  4.61 11.345 4.745 11.41 ;
        RECT  4.22 10.7925 4.78 10.8575 ;
        RECT  4.22 9.4475 4.78 9.5125 ;
        RECT  4.2875 9.5125 4.3525 9.7625 ;
        RECT  4.2875 10.6575 4.3525 10.7925 ;
        RECT  4.6475 10.7225 4.7125 10.7925 ;
        RECT  4.6475 9.5125 4.7125 9.6275 ;
        RECT  4.4575 9.6275 4.5225 10.69 ;
        RECT  4.745 10.165 4.78 10.23 ;
        RECT  4.22 10.165 4.4575 10.23 ;
        RECT  4.6475 10.4525 4.7125 10.5875 ;
        RECT  4.4575 10.4525 4.5225 10.5875 ;
        RECT  4.6475 9.6275 4.7125 9.7625 ;
        RECT  4.4575 9.6275 4.5225 9.7625 ;
        RECT  4.2875 9.6275 4.3525 9.7625 ;
        RECT  4.2875 10.5875 4.3525 10.7225 ;
        RECT  4.61 10.165 4.745 10.23 ;
        RECT  4.22 13.4825 4.78 13.5475 ;
        RECT  4.22 14.8275 4.78 14.8925 ;
        RECT  4.2875 14.5775 4.3525 14.8275 ;
        RECT  4.2875 13.5475 4.3525 13.6825 ;
        RECT  4.6475 13.5475 4.7125 13.6175 ;
        RECT  4.6475 14.7125 4.7125 14.8275 ;
        RECT  4.4575 13.65 4.5225 14.7125 ;
        RECT  4.745 14.11 4.78 14.175 ;
        RECT  4.22 14.11 4.4575 14.175 ;
        RECT  4.6475 13.6825 4.7125 13.8175 ;
        RECT  4.4575 13.6825 4.5225 13.8175 ;
        RECT  4.6475 14.2875 4.7125 14.4225 ;
        RECT  4.4575 14.2875 4.5225 14.4225 ;
        RECT  4.2875 14.4425 4.3525 14.5775 ;
        RECT  4.2875 13.4825 4.3525 13.6175 ;
        RECT  4.61 14.035 4.745 14.1 ;
        RECT  4.78 8.1025 5.53 8.1675 ;
        RECT  4.78 6.7575 5.53 6.8225 ;
        RECT  4.8475 6.79 4.9125 7.0725 ;
        RECT  4.8475 7.955 4.9125 8.135 ;
        RECT  5.3975 6.79 5.4625 7.0725 ;
        RECT  5.0175 6.79 5.0825 7.0725 ;
        RECT  5.3975 7.8525 5.4625 8.135 ;
        RECT  5.495 7.16 5.53 7.225 ;
        RECT  5.255 7.69 5.53 7.755 ;
        RECT  4.78 7.4725 5.0175 7.5375 ;
        RECT  5.3975 7.7175 5.4625 7.8525 ;
        RECT  5.2075 7.7175 5.2725 7.8525 ;
        RECT  5.2075 7.7175 5.2725 7.8525 ;
        RECT  5.0175 7.7175 5.0825 7.8525 ;
        RECT  5.3975 6.9375 5.4625 7.0725 ;
        RECT  5.2075 6.9375 5.2725 7.0725 ;
        RECT  5.2075 6.9375 5.2725 7.0725 ;
        RECT  5.0175 6.9375 5.0825 7.0725 ;
        RECT  4.8475 6.9375 4.9125 7.0725 ;
        RECT  4.8475 7.8525 4.9125 7.9875 ;
        RECT  4.985 7.175 5.05 7.24 ;
        RECT  5.2075 7.175 5.2725 7.24 ;
        RECT  4.985 7.2075 5.05 7.9875 ;
        RECT  5.0175 7.175 5.24 7.24 ;
        RECT  5.2075 7.0725 5.2725 7.2075 ;
        RECT  5.36 7.16 5.495 7.225 ;
        RECT  5.12 7.69 5.255 7.755 ;
        RECT  4.78 10.7925 5.53 10.8575 ;
        RECT  4.78 12.1375 5.53 12.2025 ;
        RECT  4.8475 11.8875 4.9125 12.17 ;
        RECT  4.8475 10.825 4.9125 11.005 ;
        RECT  5.3975 11.8875 5.4625 12.17 ;
        RECT  5.0175 11.8875 5.0825 12.17 ;
        RECT  5.3975 10.825 5.4625 11.1075 ;
        RECT  5.495 11.735 5.53 11.8 ;
        RECT  5.255 11.205 5.53 11.27 ;
        RECT  4.78 11.4225 5.0175 11.4875 ;
        RECT  5.3975 11.1275 5.4625 11.2625 ;
        RECT  5.2075 11.1275 5.2725 11.2625 ;
        RECT  5.2075 11.1275 5.2725 11.2625 ;
        RECT  5.0175 11.1275 5.0825 11.2625 ;
        RECT  5.3975 11.5975 5.4625 11.7325 ;
        RECT  5.2075 11.5975 5.2725 11.7325 ;
        RECT  5.2075 11.5975 5.2725 11.7325 ;
        RECT  5.0175 11.5975 5.0825 11.7325 ;
        RECT  4.8475 11.7525 4.9125 11.8875 ;
        RECT  4.8475 10.8375 4.9125 10.9725 ;
        RECT  4.985 10.16 5.05 10.225 ;
        RECT  5.2075 10.16 5.2725 10.225 ;
        RECT  4.985 10.1925 5.05 10.9725 ;
        RECT  5.0175 10.16 5.24 10.225 ;
        RECT  5.2075 10.0575 5.2725 10.1925 ;
        RECT  5.36 11.66 5.495 11.725 ;
        RECT  5.12 11.13 5.255 11.195 ;
        RECT  4.78 10.7925 5.53 10.8575 ;
        RECT  4.78 9.4475 5.53 9.5125 ;
        RECT  4.8475 9.48 4.9125 9.7625 ;
        RECT  4.8475 10.645 4.9125 10.825 ;
        RECT  5.3975 9.48 5.4625 9.7625 ;
        RECT  5.0175 9.48 5.0825 9.7625 ;
        RECT  5.3975 10.5425 5.4625 10.825 ;
        RECT  5.495 9.85 5.53 9.915 ;
        RECT  5.255 10.38 5.53 10.445 ;
        RECT  4.78 10.1625 5.0175 10.2275 ;
        RECT  5.3975 10.4075 5.4625 10.5425 ;
        RECT  5.2075 10.4075 5.2725 10.5425 ;
        RECT  5.2075 10.4075 5.2725 10.5425 ;
        RECT  5.0175 10.4075 5.0825 10.5425 ;
        RECT  5.3975 9.6275 5.4625 9.7625 ;
        RECT  5.2075 9.6275 5.2725 9.7625 ;
        RECT  5.2075 9.6275 5.2725 9.7625 ;
        RECT  5.0175 9.6275 5.0825 9.7625 ;
        RECT  4.8475 9.6275 4.9125 9.7625 ;
        RECT  4.8475 10.5425 4.9125 10.6775 ;
        RECT  4.985 9.865 5.05 9.93 ;
        RECT  5.2075 9.865 5.2725 9.93 ;
        RECT  4.985 9.8975 5.05 10.6775 ;
        RECT  5.0175 9.865 5.24 9.93 ;
        RECT  5.2075 9.7625 5.2725 9.8975 ;
        RECT  5.36 9.85 5.495 9.915 ;
        RECT  5.12 10.38 5.255 10.445 ;
        RECT  4.78 13.4825 5.53 13.5475 ;
        RECT  4.78 14.8275 5.53 14.8925 ;
        RECT  4.8475 14.5775 4.9125 14.86 ;
        RECT  4.8475 13.515 4.9125 13.695 ;
        RECT  5.3975 14.5775 5.4625 14.86 ;
        RECT  5.0175 14.5775 5.0825 14.86 ;
        RECT  5.3975 13.515 5.4625 13.7975 ;
        RECT  5.495 14.425 5.53 14.49 ;
        RECT  5.255 13.895 5.53 13.96 ;
        RECT  4.78 14.1125 5.0175 14.1775 ;
        RECT  5.3975 13.8175 5.4625 13.9525 ;
        RECT  5.2075 13.8175 5.2725 13.9525 ;
        RECT  5.2075 13.8175 5.2725 13.9525 ;
        RECT  5.0175 13.8175 5.0825 13.9525 ;
        RECT  5.3975 14.2875 5.4625 14.4225 ;
        RECT  5.2075 14.2875 5.2725 14.4225 ;
        RECT  5.2075 14.2875 5.2725 14.4225 ;
        RECT  5.0175 14.2875 5.0825 14.4225 ;
        RECT  4.8475 14.4425 4.9125 14.5775 ;
        RECT  4.8475 13.5275 4.9125 13.6625 ;
        RECT  4.985 12.85 5.05 12.915 ;
        RECT  5.2075 12.85 5.2725 12.915 ;
        RECT  4.985 12.8825 5.05 13.6625 ;
        RECT  5.0175 12.85 5.24 12.915 ;
        RECT  5.2075 12.7475 5.2725 12.8825 ;
        RECT  5.36 14.35 5.495 14.415 ;
        RECT  5.12 13.82 5.255 13.885 ;
        RECT  6.125 9.1825 6.26 9.2475 ;
        RECT  7.49 8.66 7.625 8.725 ;
        RECT  5.95 9.5725 6.085 9.6375 ;
        RECT  7.315 10.095 7.45 10.16 ;
        RECT  6.125 8.975 6.26 9.04 ;
        RECT  5.95 8.445 6.085 8.51 ;
        RECT  5.775 9.78 5.91 9.845 ;
        RECT  5.95 10.31 6.085 10.375 ;
        RECT  6.125 11.665 6.26 11.73 ;
        RECT  5.6 11.135 5.735 11.2 ;
        RECT  5.775 12.47 5.91 12.535 ;
        RECT  7.49 12.47 7.625 12.535 ;
        RECT  5.6 13.0 5.735 13.065 ;
        RECT  7.315 13.0 7.45 13.065 ;
        RECT  6.3 8.0325 6.435 8.0975 ;
        RECT  6.475 9.3775 6.61 9.4425 ;
        RECT  6.3 10.7225 6.435 10.7875 ;
        RECT  6.475 12.0675 6.61 12.1325 ;
        RECT  6.3 13.235 6.435 13.3 ;
        RECT  4.715 14.1125 4.78 14.1775 ;
        RECT  4.715 15.5425 4.78 15.6075 ;
        RECT  4.715 16.8025 4.78 16.8675 ;
        RECT  4.715 18.2325 4.78 18.2975 ;
        RECT  6.62 14.11 6.685 14.6975 ;
        RECT  6.16 14.6325 6.685 14.6975 ;
        RECT  7.175 14.11 7.595 14.175 ;
        RECT  6.51 14.8275 7.245 14.8925 ;
        RECT  6.335 13.4825 7.245 13.5475 ;
        RECT  6.62 15.0225 6.685 15.61 ;
        RECT  5.985 15.0225 6.685 15.0875 ;
        RECT  7.175 15.545 7.42 15.61 ;
        RECT  6.51 14.8275 7.245 14.8925 ;
        RECT  6.335 16.1725 7.245 16.2375 ;
        RECT  5.53 14.425 6.23 14.49 ;
        RECT  5.53 13.895 6.055 13.96 ;
        RECT  5.53 15.23 5.88 15.295 ;
        RECT  5.53 15.76 6.055 15.825 ;
        RECT  5.53 17.115 6.23 17.18 ;
        RECT  5.53 16.585 5.705 16.65 ;
        RECT  5.53 17.92 5.88 17.985 ;
        RECT  5.53 17.92 7.595 17.985 ;
        RECT  5.53 18.45 5.705 18.515 ;
        RECT  5.53 18.45 7.42 18.515 ;
        RECT  5.53 13.4825 6.405 13.5475 ;
        RECT  5.53 14.8275 6.58 14.8925 ;
        RECT  5.53 16.1725 6.405 16.2375 ;
        RECT  5.53 17.5175 6.58 17.5825 ;
        RECT  5.53 18.8625 6.405 18.9275 ;
        RECT  6.34 18.685 6.405 18.8625 ;
        RECT  6.685 13.4825 7.245 13.5475 ;
        RECT  6.685 12.1375 7.245 12.2025 ;
        RECT  6.7525 12.2025 6.8175 12.4525 ;
        RECT  6.7525 13.3475 6.8175 13.4825 ;
        RECT  7.1125 13.4125 7.1775 13.4825 ;
        RECT  7.1125 12.2025 7.1775 12.3175 ;
        RECT  6.9225 12.3175 6.9875 13.38 ;
        RECT  7.21 12.855 7.245 12.92 ;
        RECT  6.685 12.855 6.9225 12.92 ;
        RECT  7.1125 13.1425 7.1775 13.2775 ;
        RECT  6.9225 13.1425 6.9875 13.2775 ;
        RECT  7.1125 12.3175 7.1775 12.4525 ;
        RECT  6.9225 12.3175 6.9875 12.4525 ;
        RECT  6.7525 12.3175 6.8175 12.4525 ;
        RECT  6.7525 13.2775 6.8175 13.4125 ;
        RECT  7.075 12.855 7.21 12.92 ;
        RECT  6.685 16.1725 7.245 16.2375 ;
        RECT  6.685 17.5175 7.245 17.5825 ;
        RECT  6.7525 17.2675 6.8175 17.5175 ;
        RECT  6.7525 16.2375 6.8175 16.3725 ;
        RECT  7.1125 16.2375 7.1775 16.3075 ;
        RECT  7.1125 17.4025 7.1775 17.5175 ;
        RECT  6.9225 16.34 6.9875 17.4025 ;
        RECT  7.21 16.8 7.245 16.865 ;
        RECT  6.685 16.8 6.9225 16.865 ;
        RECT  7.1125 16.3725 7.1775 16.5075 ;
        RECT  6.9225 16.3725 6.9875 16.5075 ;
        RECT  7.1125 16.9775 7.1775 17.1125 ;
        RECT  6.9225 16.9775 6.9875 17.1125 ;
        RECT  6.7525 17.1325 6.8175 17.2675 ;
        RECT  6.7525 16.1725 6.8175 16.3075 ;
        RECT  7.075 16.725 7.21 16.79 ;
        RECT  4.22 13.4825 4.78 13.5475 ;
        RECT  4.22 12.1375 4.78 12.2025 ;
        RECT  4.2875 12.2025 4.3525 12.4525 ;
        RECT  4.2875 13.3475 4.3525 13.4825 ;
        RECT  4.6475 13.4125 4.7125 13.4825 ;
        RECT  4.6475 12.2025 4.7125 12.3175 ;
        RECT  4.4575 12.3175 4.5225 13.38 ;
        RECT  4.745 12.855 4.78 12.92 ;
        RECT  4.22 12.855 4.4575 12.92 ;
        RECT  4.6475 13.1425 4.7125 13.2775 ;
        RECT  4.4575 13.1425 4.5225 13.2775 ;
        RECT  4.6475 12.3175 4.7125 12.4525 ;
        RECT  4.4575 12.3175 4.5225 12.4525 ;
        RECT  4.2875 12.3175 4.3525 12.4525 ;
        RECT  4.2875 13.2775 4.3525 13.4125 ;
        RECT  4.61 12.855 4.745 12.92 ;
        RECT  4.22 16.1725 4.78 16.2375 ;
        RECT  4.22 17.5175 4.78 17.5825 ;
        RECT  4.2875 17.2675 4.3525 17.5175 ;
        RECT  4.2875 16.2375 4.3525 16.3725 ;
        RECT  4.6475 16.2375 4.7125 16.3075 ;
        RECT  4.6475 17.4025 4.7125 17.5175 ;
        RECT  4.4575 16.34 4.5225 17.4025 ;
        RECT  4.745 16.8 4.78 16.865 ;
        RECT  4.22 16.8 4.4575 16.865 ;
        RECT  4.6475 16.3725 4.7125 16.5075 ;
        RECT  4.4575 16.3725 4.5225 16.5075 ;
        RECT  4.6475 16.9775 4.7125 17.1125 ;
        RECT  4.4575 16.9775 4.5225 17.1125 ;
        RECT  4.2875 17.1325 4.3525 17.2675 ;
        RECT  4.2875 16.1725 4.3525 16.3075 ;
        RECT  4.61 16.725 4.745 16.79 ;
        RECT  4.22 16.1725 4.78 16.2375 ;
        RECT  4.22 14.8275 4.78 14.8925 ;
        RECT  4.2875 14.8925 4.3525 15.1425 ;
        RECT  4.2875 16.0375 4.3525 16.1725 ;
        RECT  4.6475 16.1025 4.7125 16.1725 ;
        RECT  4.6475 14.8925 4.7125 15.0075 ;
        RECT  4.4575 15.0075 4.5225 16.07 ;
        RECT  4.745 15.545 4.78 15.61 ;
        RECT  4.22 15.545 4.4575 15.61 ;
        RECT  4.6475 15.8325 4.7125 15.9675 ;
        RECT  4.4575 15.8325 4.5225 15.9675 ;
        RECT  4.6475 15.0075 4.7125 15.1425 ;
        RECT  4.4575 15.0075 4.5225 15.1425 ;
        RECT  4.2875 15.0075 4.3525 15.1425 ;
        RECT  4.2875 15.9675 4.3525 16.1025 ;
        RECT  4.61 15.545 4.745 15.61 ;
        RECT  4.22 18.8625 4.78 18.9275 ;
        RECT  4.22 20.2075 4.78 20.2725 ;
        RECT  4.2875 19.9575 4.3525 20.2075 ;
        RECT  4.2875 18.9275 4.3525 19.0625 ;
        RECT  4.6475 18.9275 4.7125 18.9975 ;
        RECT  4.6475 20.0925 4.7125 20.2075 ;
        RECT  4.4575 19.03 4.5225 20.0925 ;
        RECT  4.745 19.49 4.78 19.555 ;
        RECT  4.22 19.49 4.4575 19.555 ;
        RECT  4.6475 19.0625 4.7125 19.1975 ;
        RECT  4.4575 19.0625 4.5225 19.1975 ;
        RECT  4.6475 19.6675 4.7125 19.8025 ;
        RECT  4.4575 19.6675 4.5225 19.8025 ;
        RECT  4.2875 19.8225 4.3525 19.9575 ;
        RECT  4.2875 18.8625 4.3525 18.9975 ;
        RECT  4.61 19.415 4.745 19.48 ;
        RECT  4.78 13.4825 5.53 13.5475 ;
        RECT  4.78 12.1375 5.53 12.2025 ;
        RECT  4.8475 12.17 4.9125 12.4525 ;
        RECT  4.8475 13.335 4.9125 13.515 ;
        RECT  5.3975 12.17 5.4625 12.4525 ;
        RECT  5.0175 12.17 5.0825 12.4525 ;
        RECT  5.3975 13.2325 5.4625 13.515 ;
        RECT  5.495 12.54 5.53 12.605 ;
        RECT  5.255 13.07 5.53 13.135 ;
        RECT  4.78 12.8525 5.0175 12.9175 ;
        RECT  5.3975 13.0975 5.4625 13.2325 ;
        RECT  5.2075 13.0975 5.2725 13.2325 ;
        RECT  5.2075 13.0975 5.2725 13.2325 ;
        RECT  5.0175 13.0975 5.0825 13.2325 ;
        RECT  5.3975 12.3175 5.4625 12.4525 ;
        RECT  5.2075 12.3175 5.2725 12.4525 ;
        RECT  5.2075 12.3175 5.2725 12.4525 ;
        RECT  5.0175 12.3175 5.0825 12.4525 ;
        RECT  4.8475 12.3175 4.9125 12.4525 ;
        RECT  4.8475 13.2325 4.9125 13.3675 ;
        RECT  4.985 12.555 5.05 12.62 ;
        RECT  5.2075 12.555 5.2725 12.62 ;
        RECT  4.985 12.5875 5.05 13.3675 ;
        RECT  5.0175 12.555 5.24 12.62 ;
        RECT  5.2075 12.4525 5.2725 12.5875 ;
        RECT  5.36 12.54 5.495 12.605 ;
        RECT  5.12 13.07 5.255 13.135 ;
        RECT  4.78 16.1725 5.53 16.2375 ;
        RECT  4.78 17.5175 5.53 17.5825 ;
        RECT  4.8475 17.2675 4.9125 17.55 ;
        RECT  4.8475 16.205 4.9125 16.385 ;
        RECT  5.3975 17.2675 5.4625 17.55 ;
        RECT  5.0175 17.2675 5.0825 17.55 ;
        RECT  5.3975 16.205 5.4625 16.4875 ;
        RECT  5.495 17.115 5.53 17.18 ;
        RECT  5.255 16.585 5.53 16.65 ;
        RECT  4.78 16.8025 5.0175 16.8675 ;
        RECT  5.3975 16.5075 5.4625 16.6425 ;
        RECT  5.2075 16.5075 5.2725 16.6425 ;
        RECT  5.2075 16.5075 5.2725 16.6425 ;
        RECT  5.0175 16.5075 5.0825 16.6425 ;
        RECT  5.3975 16.9775 5.4625 17.1125 ;
        RECT  5.2075 16.9775 5.2725 17.1125 ;
        RECT  5.2075 16.9775 5.2725 17.1125 ;
        RECT  5.0175 16.9775 5.0825 17.1125 ;
        RECT  4.8475 17.1325 4.9125 17.2675 ;
        RECT  4.8475 16.2175 4.9125 16.3525 ;
        RECT  4.985 15.54 5.05 15.605 ;
        RECT  5.2075 15.54 5.2725 15.605 ;
        RECT  4.985 15.5725 5.05 16.3525 ;
        RECT  5.0175 15.54 5.24 15.605 ;
        RECT  5.2075 15.4375 5.2725 15.5725 ;
        RECT  5.36 17.04 5.495 17.105 ;
        RECT  5.12 16.51 5.255 16.575 ;
        RECT  4.78 16.1725 5.53 16.2375 ;
        RECT  4.78 14.8275 5.53 14.8925 ;
        RECT  4.8475 14.86 4.9125 15.1425 ;
        RECT  4.8475 16.025 4.9125 16.205 ;
        RECT  5.3975 14.86 5.4625 15.1425 ;
        RECT  5.0175 14.86 5.0825 15.1425 ;
        RECT  5.3975 15.9225 5.4625 16.205 ;
        RECT  5.495 15.23 5.53 15.295 ;
        RECT  5.255 15.76 5.53 15.825 ;
        RECT  4.78 15.5425 5.0175 15.6075 ;
        RECT  5.3975 15.7875 5.4625 15.9225 ;
        RECT  5.2075 15.7875 5.2725 15.9225 ;
        RECT  5.2075 15.7875 5.2725 15.9225 ;
        RECT  5.0175 15.7875 5.0825 15.9225 ;
        RECT  5.3975 15.0075 5.4625 15.1425 ;
        RECT  5.2075 15.0075 5.2725 15.1425 ;
        RECT  5.2075 15.0075 5.2725 15.1425 ;
        RECT  5.0175 15.0075 5.0825 15.1425 ;
        RECT  4.8475 15.0075 4.9125 15.1425 ;
        RECT  4.8475 15.9225 4.9125 16.0575 ;
        RECT  4.985 15.245 5.05 15.31 ;
        RECT  5.2075 15.245 5.2725 15.31 ;
        RECT  4.985 15.2775 5.05 16.0575 ;
        RECT  5.0175 15.245 5.24 15.31 ;
        RECT  5.2075 15.1425 5.2725 15.2775 ;
        RECT  5.36 15.23 5.495 15.295 ;
        RECT  5.12 15.76 5.255 15.825 ;
        RECT  4.78 18.8625 5.53 18.9275 ;
        RECT  4.78 20.2075 5.53 20.2725 ;
        RECT  4.8475 19.9575 4.9125 20.24 ;
        RECT  4.8475 18.895 4.9125 19.075 ;
        RECT  5.3975 19.9575 5.4625 20.24 ;
        RECT  5.0175 19.9575 5.0825 20.24 ;
        RECT  5.3975 18.895 5.4625 19.1775 ;
        RECT  5.495 19.805 5.53 19.87 ;
        RECT  5.255 19.275 5.53 19.34 ;
        RECT  4.78 19.4925 5.0175 19.5575 ;
        RECT  5.3975 19.1975 5.4625 19.3325 ;
        RECT  5.2075 19.1975 5.2725 19.3325 ;
        RECT  5.2075 19.1975 5.2725 19.3325 ;
        RECT  5.0175 19.1975 5.0825 19.3325 ;
        RECT  5.3975 19.6675 5.4625 19.8025 ;
        RECT  5.2075 19.6675 5.2725 19.8025 ;
        RECT  5.2075 19.6675 5.2725 19.8025 ;
        RECT  5.0175 19.6675 5.0825 19.8025 ;
        RECT  4.8475 19.8225 4.9125 19.9575 ;
        RECT  4.8475 18.9075 4.9125 19.0425 ;
        RECT  4.985 18.23 5.05 18.295 ;
        RECT  5.2075 18.23 5.2725 18.295 ;
        RECT  4.985 18.2625 5.05 19.0425 ;
        RECT  5.0175 18.23 5.24 18.295 ;
        RECT  5.2075 18.1275 5.2725 18.2625 ;
        RECT  5.36 19.73 5.495 19.795 ;
        RECT  5.12 19.2 5.255 19.265 ;
        RECT  6.125 14.5625 6.26 14.6275 ;
        RECT  7.49 14.04 7.625 14.105 ;
        RECT  5.95 14.9525 6.085 15.0175 ;
        RECT  7.315 15.475 7.45 15.54 ;
        RECT  6.125 14.355 6.26 14.42 ;
        RECT  5.95 13.825 6.085 13.89 ;
        RECT  5.775 15.16 5.91 15.225 ;
        RECT  5.95 15.69 6.085 15.755 ;
        RECT  6.125 17.045 6.26 17.11 ;
        RECT  5.6 16.515 5.735 16.58 ;
        RECT  5.775 17.85 5.91 17.915 ;
        RECT  7.49 17.85 7.625 17.915 ;
        RECT  5.6 18.38 5.735 18.445 ;
        RECT  7.315 18.38 7.45 18.445 ;
        RECT  6.3 13.4125 6.435 13.4775 ;
        RECT  6.475 14.7575 6.61 14.8225 ;
        RECT  6.3 16.1025 6.435 16.1675 ;
        RECT  6.475 17.4475 6.61 17.5125 ;
        RECT  6.3 18.615 6.435 18.68 ;
        RECT  4.22 18.8625 4.97 18.9275 ;
        RECT  4.22 20.2075 4.97 20.2725 ;
        RECT  4.8375 19.9575 4.9025 20.24 ;
        RECT  4.8375 18.895 4.9025 19.075 ;
        RECT  4.2875 19.9575 4.3525 20.24 ;
        RECT  4.6675 19.9575 4.7325 20.24 ;
        RECT  4.2875 18.895 4.3525 19.1775 ;
        RECT  4.22 19.805 4.255 19.87 ;
        RECT  4.22 19.275 4.495 19.34 ;
        RECT  4.7325 19.4925 4.97 19.5575 ;
        RECT  4.2875 19.1775 4.3525 19.3125 ;
        RECT  4.4775 19.1775 4.5425 19.3125 ;
        RECT  4.4775 19.1775 4.5425 19.3125 ;
        RECT  4.6675 19.1775 4.7325 19.3125 ;
        RECT  4.2875 19.9575 4.3525 20.0925 ;
        RECT  4.4775 19.9575 4.5425 20.0925 ;
        RECT  4.4775 19.9575 4.5425 20.0925 ;
        RECT  4.6675 19.9575 4.7325 20.0925 ;
        RECT  4.8375 19.9575 4.9025 20.0925 ;
        RECT  4.8375 19.0425 4.9025 19.1775 ;
        RECT  4.7 19.79 4.765 19.855 ;
        RECT  4.4775 19.79 4.5425 19.855 ;
        RECT  4.7 19.0425 4.765 19.8225 ;
        RECT  4.51 19.79 4.7325 19.855 ;
        RECT  4.4775 19.8225 4.5425 19.9575 ;
        RECT  4.255 19.805 4.39 19.87 ;
        RECT  4.495 19.275 4.63 19.34 ;
        RECT  4.22 21.5525 4.97 21.6175 ;
        RECT  4.22 20.2075 4.97 20.2725 ;
        RECT  4.8375 20.24 4.9025 20.5225 ;
        RECT  4.8375 21.405 4.9025 21.585 ;
        RECT  4.2875 20.24 4.3525 20.5225 ;
        RECT  4.6675 20.24 4.7325 20.5225 ;
        RECT  4.2875 21.3025 4.3525 21.585 ;
        RECT  4.22 20.61 4.255 20.675 ;
        RECT  4.22 21.14 4.495 21.205 ;
        RECT  4.7325 20.9225 4.97 20.9875 ;
        RECT  4.2875 21.1475 4.3525 21.2825 ;
        RECT  4.4775 21.1475 4.5425 21.2825 ;
        RECT  4.4775 21.1475 4.5425 21.2825 ;
        RECT  4.6675 21.1475 4.7325 21.2825 ;
        RECT  4.2875 20.6775 4.3525 20.8125 ;
        RECT  4.4775 20.6775 4.5425 20.8125 ;
        RECT  4.4775 20.6775 4.5425 20.8125 ;
        RECT  4.6675 20.6775 4.7325 20.8125 ;
        RECT  4.8375 20.5225 4.9025 20.6575 ;
        RECT  4.8375 21.4375 4.9025 21.5725 ;
        RECT  4.7 22.185 4.765 22.25 ;
        RECT  4.4775 22.185 4.5425 22.25 ;
        RECT  4.7 21.4375 4.765 22.2175 ;
        RECT  4.51 22.185 4.7325 22.25 ;
        RECT  4.4775 22.2175 4.5425 22.3525 ;
        RECT  4.255 20.685 4.39 20.75 ;
        RECT  4.495 21.215 4.63 21.28 ;
        RECT  4.22 21.5525 4.97 21.6175 ;
        RECT  4.22 22.8975 4.97 22.9625 ;
        RECT  4.8375 22.6475 4.9025 22.93 ;
        RECT  4.8375 21.585 4.9025 21.765 ;
        RECT  4.2875 22.6475 4.3525 22.93 ;
        RECT  4.6675 22.6475 4.7325 22.93 ;
        RECT  4.2875 21.585 4.3525 21.8675 ;
        RECT  4.22 22.495 4.255 22.56 ;
        RECT  4.22 21.965 4.495 22.03 ;
        RECT  4.7325 22.1825 4.97 22.2475 ;
        RECT  4.2875 21.8675 4.3525 22.0025 ;
        RECT  4.4775 21.8675 4.5425 22.0025 ;
        RECT  4.4775 21.8675 4.5425 22.0025 ;
        RECT  4.6675 21.8675 4.7325 22.0025 ;
        RECT  4.2875 22.6475 4.3525 22.7825 ;
        RECT  4.4775 22.6475 4.5425 22.7825 ;
        RECT  4.4775 22.6475 4.5425 22.7825 ;
        RECT  4.6675 22.6475 4.7325 22.7825 ;
        RECT  4.8375 22.6475 4.9025 22.7825 ;
        RECT  4.8375 21.7325 4.9025 21.8675 ;
        RECT  4.7 22.48 4.765 22.545 ;
        RECT  4.4775 22.48 4.5425 22.545 ;
        RECT  4.7 21.7325 4.765 22.5125 ;
        RECT  4.51 22.48 4.7325 22.545 ;
        RECT  4.4775 22.5125 4.5425 22.6475 ;
        RECT  4.255 22.495 4.39 22.56 ;
        RECT  4.495 21.965 4.63 22.03 ;
        RECT  4.22 24.2425 4.97 24.3075 ;
        RECT  4.22 22.8975 4.97 22.9625 ;
        RECT  4.8375 22.93 4.9025 23.2125 ;
        RECT  4.8375 24.095 4.9025 24.275 ;
        RECT  4.2875 22.93 4.3525 23.2125 ;
        RECT  4.6675 22.93 4.7325 23.2125 ;
        RECT  4.2875 23.9925 4.3525 24.275 ;
        RECT  4.22 23.3 4.255 23.365 ;
        RECT  4.22 23.83 4.495 23.895 ;
        RECT  4.7325 23.6125 4.97 23.6775 ;
        RECT  4.2875 23.8375 4.3525 23.9725 ;
        RECT  4.4775 23.8375 4.5425 23.9725 ;
        RECT  4.4775 23.8375 4.5425 23.9725 ;
        RECT  4.6675 23.8375 4.7325 23.9725 ;
        RECT  4.2875 23.3675 4.3525 23.5025 ;
        RECT  4.4775 23.3675 4.5425 23.5025 ;
        RECT  4.4775 23.3675 4.5425 23.5025 ;
        RECT  4.6675 23.3675 4.7325 23.5025 ;
        RECT  4.8375 23.2125 4.9025 23.3475 ;
        RECT  4.8375 24.1275 4.9025 24.2625 ;
        RECT  4.7 24.875 4.765 24.94 ;
        RECT  4.4775 24.875 4.5425 24.94 ;
        RECT  4.7 24.1275 4.765 24.9075 ;
        RECT  4.51 24.875 4.7325 24.94 ;
        RECT  4.4775 24.9075 4.5425 25.0425 ;
        RECT  4.255 23.375 4.39 23.44 ;
        RECT  4.495 23.905 4.63 23.97 ;
        RECT  4.22 24.2425 4.97 24.3075 ;
        RECT  4.22 25.5875 4.97 25.6525 ;
        RECT  4.8375 25.3375 4.9025 25.62 ;
        RECT  4.8375 24.275 4.9025 24.455 ;
        RECT  4.2875 25.3375 4.3525 25.62 ;
        RECT  4.6675 25.3375 4.7325 25.62 ;
        RECT  4.2875 24.275 4.3525 24.5575 ;
        RECT  4.22 25.185 4.255 25.25 ;
        RECT  4.22 24.655 4.495 24.72 ;
        RECT  4.7325 24.8725 4.97 24.9375 ;
        RECT  4.2875 24.5575 4.3525 24.6925 ;
        RECT  4.4775 24.5575 4.5425 24.6925 ;
        RECT  4.4775 24.5575 4.5425 24.6925 ;
        RECT  4.6675 24.5575 4.7325 24.6925 ;
        RECT  4.2875 25.3375 4.3525 25.4725 ;
        RECT  4.4775 25.3375 4.5425 25.4725 ;
        RECT  4.4775 25.3375 4.5425 25.4725 ;
        RECT  4.6675 25.3375 4.7325 25.4725 ;
        RECT  4.8375 25.3375 4.9025 25.4725 ;
        RECT  4.8375 24.4225 4.9025 24.5575 ;
        RECT  4.7 25.17 4.765 25.235 ;
        RECT  4.4775 25.17 4.5425 25.235 ;
        RECT  4.7 24.4225 4.765 25.2025 ;
        RECT  4.51 25.17 4.7325 25.235 ;
        RECT  4.4775 25.2025 4.5425 25.3375 ;
        RECT  4.255 25.185 4.39 25.25 ;
        RECT  4.495 24.655 4.63 24.72 ;
        RECT  4.22 26.9325 4.97 26.9975 ;
        RECT  4.22 25.5875 4.97 25.6525 ;
        RECT  4.8375 25.62 4.9025 25.9025 ;
        RECT  4.8375 26.785 4.9025 26.965 ;
        RECT  4.2875 25.62 4.3525 25.9025 ;
        RECT  4.6675 25.62 4.7325 25.9025 ;
        RECT  4.2875 26.6825 4.3525 26.965 ;
        RECT  4.22 25.99 4.255 26.055 ;
        RECT  4.22 26.52 4.495 26.585 ;
        RECT  4.7325 26.3025 4.97 26.3675 ;
        RECT  4.2875 26.5275 4.3525 26.6625 ;
        RECT  4.4775 26.5275 4.5425 26.6625 ;
        RECT  4.4775 26.5275 4.5425 26.6625 ;
        RECT  4.6675 26.5275 4.7325 26.6625 ;
        RECT  4.2875 26.0575 4.3525 26.1925 ;
        RECT  4.4775 26.0575 4.5425 26.1925 ;
        RECT  4.4775 26.0575 4.5425 26.1925 ;
        RECT  4.6675 26.0575 4.7325 26.1925 ;
        RECT  4.8375 25.9025 4.9025 26.0375 ;
        RECT  4.8375 26.8175 4.9025 26.9525 ;
        RECT  4.7 27.565 4.765 27.63 ;
        RECT  4.4775 27.565 4.5425 27.63 ;
        RECT  4.7 26.8175 4.765 27.5975 ;
        RECT  4.51 27.565 4.7325 27.63 ;
        RECT  4.4775 27.5975 4.5425 27.7325 ;
        RECT  4.255 26.065 4.39 26.13 ;
        RECT  4.495 26.595 4.63 26.66 ;
        RECT  4.22 26.9325 4.97 26.9975 ;
        RECT  4.22 28.2775 4.97 28.3425 ;
        RECT  4.8375 28.0275 4.9025 28.31 ;
        RECT  4.8375 26.965 4.9025 27.145 ;
        RECT  4.2875 28.0275 4.3525 28.31 ;
        RECT  4.6675 28.0275 4.7325 28.31 ;
        RECT  4.2875 26.965 4.3525 27.2475 ;
        RECT  4.22 27.875 4.255 27.94 ;
        RECT  4.22 27.345 4.495 27.41 ;
        RECT  4.7325 27.5625 4.97 27.6275 ;
        RECT  4.2875 27.2475 4.3525 27.3825 ;
        RECT  4.4775 27.2475 4.5425 27.3825 ;
        RECT  4.4775 27.2475 4.5425 27.3825 ;
        RECT  4.6675 27.2475 4.7325 27.3825 ;
        RECT  4.2875 28.0275 4.3525 28.1625 ;
        RECT  4.4775 28.0275 4.5425 28.1625 ;
        RECT  4.4775 28.0275 4.5425 28.1625 ;
        RECT  4.6675 28.0275 4.7325 28.1625 ;
        RECT  4.8375 28.0275 4.9025 28.1625 ;
        RECT  4.8375 27.1125 4.9025 27.2475 ;
        RECT  4.7 27.86 4.765 27.925 ;
        RECT  4.4775 27.86 4.5425 27.925 ;
        RECT  4.7 27.1125 4.765 27.8925 ;
        RECT  4.51 27.86 4.7325 27.925 ;
        RECT  4.4775 27.8925 4.5425 28.0275 ;
        RECT  4.255 27.875 4.39 27.94 ;
        RECT  4.495 27.345 4.63 27.41 ;
        RECT  4.22 29.6225 4.97 29.6875 ;
        RECT  4.22 28.2775 4.97 28.3425 ;
        RECT  4.8375 28.31 4.9025 28.5925 ;
        RECT  4.8375 29.475 4.9025 29.655 ;
        RECT  4.2875 28.31 4.3525 28.5925 ;
        RECT  4.6675 28.31 4.7325 28.5925 ;
        RECT  4.2875 29.3725 4.3525 29.655 ;
        RECT  4.22 28.68 4.255 28.745 ;
        RECT  4.22 29.21 4.495 29.275 ;
        RECT  4.7325 28.9925 4.97 29.0575 ;
        RECT  4.2875 29.2175 4.3525 29.3525 ;
        RECT  4.4775 29.2175 4.5425 29.3525 ;
        RECT  4.4775 29.2175 4.5425 29.3525 ;
        RECT  4.6675 29.2175 4.7325 29.3525 ;
        RECT  4.2875 28.7475 4.3525 28.8825 ;
        RECT  4.4775 28.7475 4.5425 28.8825 ;
        RECT  4.4775 28.7475 4.5425 28.8825 ;
        RECT  4.6675 28.7475 4.7325 28.8825 ;
        RECT  4.8375 28.5925 4.9025 28.7275 ;
        RECT  4.8375 29.5075 4.9025 29.6425 ;
        RECT  4.7 30.255 4.765 30.32 ;
        RECT  4.4775 30.255 4.5425 30.32 ;
        RECT  4.7 29.5075 4.765 30.2875 ;
        RECT  4.51 30.255 4.7325 30.32 ;
        RECT  4.4775 30.2875 4.5425 30.4225 ;
        RECT  4.255 28.755 4.39 28.82 ;
        RECT  4.495 29.285 4.63 29.35 ;
        RECT  4.22 29.6225 4.97 29.6875 ;
        RECT  4.22 30.9675 4.97 31.0325 ;
        RECT  4.8375 30.7175 4.9025 31.0 ;
        RECT  4.8375 29.655 4.9025 29.835 ;
        RECT  4.2875 30.7175 4.3525 31.0 ;
        RECT  4.6675 30.7175 4.7325 31.0 ;
        RECT  4.2875 29.655 4.3525 29.9375 ;
        RECT  4.22 30.565 4.255 30.63 ;
        RECT  4.22 30.035 4.495 30.1 ;
        RECT  4.7325 30.2525 4.97 30.3175 ;
        RECT  4.2875 29.9375 4.3525 30.0725 ;
        RECT  4.4775 29.9375 4.5425 30.0725 ;
        RECT  4.4775 29.9375 4.5425 30.0725 ;
        RECT  4.6675 29.9375 4.7325 30.0725 ;
        RECT  4.2875 30.7175 4.3525 30.8525 ;
        RECT  4.4775 30.7175 4.5425 30.8525 ;
        RECT  4.4775 30.7175 4.5425 30.8525 ;
        RECT  4.6675 30.7175 4.7325 30.8525 ;
        RECT  4.8375 30.7175 4.9025 30.8525 ;
        RECT  4.8375 29.8025 4.9025 29.9375 ;
        RECT  4.7 30.55 4.765 30.615 ;
        RECT  4.4775 30.55 4.5425 30.615 ;
        RECT  4.7 29.8025 4.765 30.5825 ;
        RECT  4.51 30.55 4.7325 30.615 ;
        RECT  4.4775 30.5825 4.5425 30.7175 ;
        RECT  4.255 30.565 4.39 30.63 ;
        RECT  4.495 30.035 4.63 30.1 ;
        RECT  4.22 32.3125 4.97 32.3775 ;
        RECT  4.22 30.9675 4.97 31.0325 ;
        RECT  4.8375 31.0 4.9025 31.2825 ;
        RECT  4.8375 32.165 4.9025 32.345 ;
        RECT  4.2875 31.0 4.3525 31.2825 ;
        RECT  4.6675 31.0 4.7325 31.2825 ;
        RECT  4.2875 32.0625 4.3525 32.345 ;
        RECT  4.22 31.37 4.255 31.435 ;
        RECT  4.22 31.9 4.495 31.965 ;
        RECT  4.7325 31.6825 4.97 31.7475 ;
        RECT  4.2875 31.9075 4.3525 32.0425 ;
        RECT  4.4775 31.9075 4.5425 32.0425 ;
        RECT  4.4775 31.9075 4.5425 32.0425 ;
        RECT  4.6675 31.9075 4.7325 32.0425 ;
        RECT  4.2875 31.4375 4.3525 31.5725 ;
        RECT  4.4775 31.4375 4.5425 31.5725 ;
        RECT  4.4775 31.4375 4.5425 31.5725 ;
        RECT  4.6675 31.4375 4.7325 31.5725 ;
        RECT  4.8375 31.2825 4.9025 31.4175 ;
        RECT  4.8375 32.1975 4.9025 32.3325 ;
        RECT  4.7 32.945 4.765 33.01 ;
        RECT  4.4775 32.945 4.5425 33.01 ;
        RECT  4.7 32.1975 4.765 32.9775 ;
        RECT  4.51 32.945 4.7325 33.01 ;
        RECT  4.4775 32.9775 4.5425 33.1125 ;
        RECT  4.255 31.445 4.39 31.51 ;
        RECT  4.495 31.975 4.63 32.04 ;
        RECT  4.22 32.3125 4.97 32.3775 ;
        RECT  4.22 33.6575 4.97 33.7225 ;
        RECT  4.8375 33.4075 4.9025 33.69 ;
        RECT  4.8375 32.345 4.9025 32.525 ;
        RECT  4.2875 33.4075 4.3525 33.69 ;
        RECT  4.6675 33.4075 4.7325 33.69 ;
        RECT  4.2875 32.345 4.3525 32.6275 ;
        RECT  4.22 33.255 4.255 33.32 ;
        RECT  4.22 32.725 4.495 32.79 ;
        RECT  4.7325 32.9425 4.97 33.0075 ;
        RECT  4.2875 32.6275 4.3525 32.7625 ;
        RECT  4.4775 32.6275 4.5425 32.7625 ;
        RECT  4.4775 32.6275 4.5425 32.7625 ;
        RECT  4.6675 32.6275 4.7325 32.7625 ;
        RECT  4.2875 33.4075 4.3525 33.5425 ;
        RECT  4.4775 33.4075 4.5425 33.5425 ;
        RECT  4.4775 33.4075 4.5425 33.5425 ;
        RECT  4.6675 33.4075 4.7325 33.5425 ;
        RECT  4.8375 33.4075 4.9025 33.5425 ;
        RECT  4.8375 32.4925 4.9025 32.6275 ;
        RECT  4.7 33.24 4.765 33.305 ;
        RECT  4.4775 33.24 4.5425 33.305 ;
        RECT  4.7 32.4925 4.765 33.2725 ;
        RECT  4.51 33.24 4.7325 33.305 ;
        RECT  4.4775 33.2725 4.5425 33.4075 ;
        RECT  4.255 33.255 4.39 33.32 ;
        RECT  4.495 32.725 4.63 32.79 ;
        RECT  4.22 35.0025 4.97 35.0675 ;
        RECT  4.22 33.6575 4.97 33.7225 ;
        RECT  4.8375 33.69 4.9025 33.9725 ;
        RECT  4.8375 34.855 4.9025 35.035 ;
        RECT  4.2875 33.69 4.3525 33.9725 ;
        RECT  4.6675 33.69 4.7325 33.9725 ;
        RECT  4.2875 34.7525 4.3525 35.035 ;
        RECT  4.22 34.06 4.255 34.125 ;
        RECT  4.22 34.59 4.495 34.655 ;
        RECT  4.7325 34.3725 4.97 34.4375 ;
        RECT  4.2875 34.5975 4.3525 34.7325 ;
        RECT  4.4775 34.5975 4.5425 34.7325 ;
        RECT  4.4775 34.5975 4.5425 34.7325 ;
        RECT  4.6675 34.5975 4.7325 34.7325 ;
        RECT  4.2875 34.1275 4.3525 34.2625 ;
        RECT  4.4775 34.1275 4.5425 34.2625 ;
        RECT  4.4775 34.1275 4.5425 34.2625 ;
        RECT  4.6675 34.1275 4.7325 34.2625 ;
        RECT  4.8375 33.9725 4.9025 34.1075 ;
        RECT  4.8375 34.8875 4.9025 35.0225 ;
        RECT  4.7 35.635 4.765 35.7 ;
        RECT  4.4775 35.635 4.5425 35.7 ;
        RECT  4.7 34.8875 4.765 35.6675 ;
        RECT  4.51 35.635 4.7325 35.7 ;
        RECT  4.4775 35.6675 4.5425 35.8025 ;
        RECT  4.255 34.135 4.39 34.2 ;
        RECT  4.495 34.665 4.63 34.73 ;
        RECT  4.22 35.0025 4.97 35.0675 ;
        RECT  4.22 36.3475 4.97 36.4125 ;
        RECT  4.8375 36.0975 4.9025 36.38 ;
        RECT  4.8375 35.035 4.9025 35.215 ;
        RECT  4.2875 36.0975 4.3525 36.38 ;
        RECT  4.6675 36.0975 4.7325 36.38 ;
        RECT  4.2875 35.035 4.3525 35.3175 ;
        RECT  4.22 35.945 4.255 36.01 ;
        RECT  4.22 35.415 4.495 35.48 ;
        RECT  4.7325 35.6325 4.97 35.6975 ;
        RECT  4.2875 35.3175 4.3525 35.4525 ;
        RECT  4.4775 35.3175 4.5425 35.4525 ;
        RECT  4.4775 35.3175 4.5425 35.4525 ;
        RECT  4.6675 35.3175 4.7325 35.4525 ;
        RECT  4.2875 36.0975 4.3525 36.2325 ;
        RECT  4.4775 36.0975 4.5425 36.2325 ;
        RECT  4.4775 36.0975 4.5425 36.2325 ;
        RECT  4.6675 36.0975 4.7325 36.2325 ;
        RECT  4.8375 36.0975 4.9025 36.2325 ;
        RECT  4.8375 35.1825 4.9025 35.3175 ;
        RECT  4.7 35.93 4.765 35.995 ;
        RECT  4.4775 35.93 4.5425 35.995 ;
        RECT  4.7 35.1825 4.765 35.9625 ;
        RECT  4.51 35.93 4.7325 35.995 ;
        RECT  4.4775 35.9625 4.5425 36.0975 ;
        RECT  4.255 35.945 4.39 36.01 ;
        RECT  4.495 35.415 4.63 35.48 ;
        RECT  4.22 37.6925 4.97 37.7575 ;
        RECT  4.22 36.3475 4.97 36.4125 ;
        RECT  4.8375 36.38 4.9025 36.6625 ;
        RECT  4.8375 37.545 4.9025 37.725 ;
        RECT  4.2875 36.38 4.3525 36.6625 ;
        RECT  4.6675 36.38 4.7325 36.6625 ;
        RECT  4.2875 37.4425 4.3525 37.725 ;
        RECT  4.22 36.75 4.255 36.815 ;
        RECT  4.22 37.28 4.495 37.345 ;
        RECT  4.7325 37.0625 4.97 37.1275 ;
        RECT  4.2875 37.2875 4.3525 37.4225 ;
        RECT  4.4775 37.2875 4.5425 37.4225 ;
        RECT  4.4775 37.2875 4.5425 37.4225 ;
        RECT  4.6675 37.2875 4.7325 37.4225 ;
        RECT  4.2875 36.8175 4.3525 36.9525 ;
        RECT  4.4775 36.8175 4.5425 36.9525 ;
        RECT  4.4775 36.8175 4.5425 36.9525 ;
        RECT  4.6675 36.8175 4.7325 36.9525 ;
        RECT  4.8375 36.6625 4.9025 36.7975 ;
        RECT  4.8375 37.5775 4.9025 37.7125 ;
        RECT  4.7 38.325 4.765 38.39 ;
        RECT  4.4775 38.325 4.5425 38.39 ;
        RECT  4.7 37.5775 4.765 38.3575 ;
        RECT  4.51 38.325 4.7325 38.39 ;
        RECT  4.4775 38.3575 4.5425 38.4925 ;
        RECT  4.255 36.825 4.39 36.89 ;
        RECT  4.495 37.355 4.63 37.42 ;
        RECT  4.22 37.6925 4.97 37.7575 ;
        RECT  4.22 39.0375 4.97 39.1025 ;
        RECT  4.8375 38.7875 4.9025 39.07 ;
        RECT  4.8375 37.725 4.9025 37.905 ;
        RECT  4.2875 38.7875 4.3525 39.07 ;
        RECT  4.6675 38.7875 4.7325 39.07 ;
        RECT  4.2875 37.725 4.3525 38.0075 ;
        RECT  4.22 38.635 4.255 38.7 ;
        RECT  4.22 38.105 4.495 38.17 ;
        RECT  4.7325 38.3225 4.97 38.3875 ;
        RECT  4.2875 38.0075 4.3525 38.1425 ;
        RECT  4.4775 38.0075 4.5425 38.1425 ;
        RECT  4.4775 38.0075 4.5425 38.1425 ;
        RECT  4.6675 38.0075 4.7325 38.1425 ;
        RECT  4.2875 38.7875 4.3525 38.9225 ;
        RECT  4.4775 38.7875 4.5425 38.9225 ;
        RECT  4.4775 38.7875 4.5425 38.9225 ;
        RECT  4.6675 38.7875 4.7325 38.9225 ;
        RECT  4.8375 38.7875 4.9025 38.9225 ;
        RECT  4.8375 37.8725 4.9025 38.0075 ;
        RECT  4.7 38.62 4.765 38.685 ;
        RECT  4.4775 38.62 4.5425 38.685 ;
        RECT  4.7 37.8725 4.765 38.6525 ;
        RECT  4.51 38.62 4.7325 38.685 ;
        RECT  4.4775 38.6525 4.5425 38.7875 ;
        RECT  4.255 38.635 4.39 38.7 ;
        RECT  4.495 38.105 4.63 38.17 ;
        RECT  4.22 40.3825 4.97 40.4475 ;
        RECT  4.22 39.0375 4.97 39.1025 ;
        RECT  4.8375 39.07 4.9025 39.3525 ;
        RECT  4.8375 40.235 4.9025 40.415 ;
        RECT  4.2875 39.07 4.3525 39.3525 ;
        RECT  4.6675 39.07 4.7325 39.3525 ;
        RECT  4.2875 40.1325 4.3525 40.415 ;
        RECT  4.22 39.44 4.255 39.505 ;
        RECT  4.22 39.97 4.495 40.035 ;
        RECT  4.7325 39.7525 4.97 39.8175 ;
        RECT  4.2875 39.9775 4.3525 40.1125 ;
        RECT  4.4775 39.9775 4.5425 40.1125 ;
        RECT  4.4775 39.9775 4.5425 40.1125 ;
        RECT  4.6675 39.9775 4.7325 40.1125 ;
        RECT  4.2875 39.5075 4.3525 39.6425 ;
        RECT  4.4775 39.5075 4.5425 39.6425 ;
        RECT  4.4775 39.5075 4.5425 39.6425 ;
        RECT  4.6675 39.5075 4.7325 39.6425 ;
        RECT  4.8375 39.3525 4.9025 39.4875 ;
        RECT  4.8375 40.2675 4.9025 40.4025 ;
        RECT  4.7 41.015 4.765 41.08 ;
        RECT  4.4775 41.015 4.5425 41.08 ;
        RECT  4.7 40.2675 4.765 41.0475 ;
        RECT  4.51 41.015 4.7325 41.08 ;
        RECT  4.4775 41.0475 4.5425 41.1825 ;
        RECT  4.255 39.515 4.39 39.58 ;
        RECT  4.495 40.045 4.63 40.11 ;
        RECT  4.97 18.8625 5.53 18.9275 ;
        RECT  4.97 20.2075 5.53 20.2725 ;
        RECT  5.3975 19.9575 5.4625 20.2075 ;
        RECT  5.3975 18.9275 5.4625 19.0625 ;
        RECT  5.0375 18.9275 5.1025 18.9975 ;
        RECT  5.0375 20.0925 5.1025 20.2075 ;
        RECT  5.2275 19.03 5.2925 20.0925 ;
        RECT  4.97 19.49 5.005 19.555 ;
        RECT  5.2925 19.49 5.53 19.555 ;
        RECT  5.0375 19.1325 5.1025 19.2675 ;
        RECT  5.2275 19.1325 5.2925 19.2675 ;
        RECT  5.0375 19.9575 5.1025 20.0925 ;
        RECT  5.2275 19.9575 5.2925 20.0925 ;
        RECT  5.3975 19.9575 5.4625 20.0925 ;
        RECT  5.3975 18.9975 5.4625 19.1325 ;
        RECT  5.005 19.49 5.14 19.555 ;
        RECT  4.97 21.5525 5.53 21.6175 ;
        RECT  4.97 20.2075 5.53 20.2725 ;
        RECT  5.3975 20.2725 5.4625 20.5225 ;
        RECT  5.3975 21.4175 5.4625 21.5525 ;
        RECT  5.0375 21.4825 5.1025 21.5525 ;
        RECT  5.0375 20.2725 5.1025 20.3875 ;
        RECT  5.2275 20.3875 5.2925 21.45 ;
        RECT  4.97 20.925 5.005 20.99 ;
        RECT  5.2925 20.925 5.53 20.99 ;
        RECT  5.0375 21.2825 5.1025 21.4175 ;
        RECT  5.2275 21.2825 5.2925 21.4175 ;
        RECT  5.0375 20.6775 5.1025 20.8125 ;
        RECT  5.2275 20.6775 5.2925 20.8125 ;
        RECT  5.3975 20.5225 5.4625 20.6575 ;
        RECT  5.3975 21.4825 5.4625 21.6175 ;
        RECT  5.005 21.0 5.14 21.065 ;
        RECT  4.97 21.5525 5.53 21.6175 ;
        RECT  4.97 22.8975 5.53 22.9625 ;
        RECT  5.3975 22.6475 5.4625 22.8975 ;
        RECT  5.3975 21.6175 5.4625 21.7525 ;
        RECT  5.0375 21.6175 5.1025 21.6875 ;
        RECT  5.0375 22.7825 5.1025 22.8975 ;
        RECT  5.2275 21.72 5.2925 22.7825 ;
        RECT  4.97 22.18 5.005 22.245 ;
        RECT  5.2925 22.18 5.53 22.245 ;
        RECT  5.0375 21.8225 5.1025 21.9575 ;
        RECT  5.2275 21.8225 5.2925 21.9575 ;
        RECT  5.0375 22.6475 5.1025 22.7825 ;
        RECT  5.2275 22.6475 5.2925 22.7825 ;
        RECT  5.3975 22.6475 5.4625 22.7825 ;
        RECT  5.3975 21.6875 5.4625 21.8225 ;
        RECT  5.005 22.18 5.14 22.245 ;
        RECT  4.97 24.2425 5.53 24.3075 ;
        RECT  4.97 22.8975 5.53 22.9625 ;
        RECT  5.3975 22.9625 5.4625 23.2125 ;
        RECT  5.3975 24.1075 5.4625 24.2425 ;
        RECT  5.0375 24.1725 5.1025 24.2425 ;
        RECT  5.0375 22.9625 5.1025 23.0775 ;
        RECT  5.2275 23.0775 5.2925 24.14 ;
        RECT  4.97 23.615 5.005 23.68 ;
        RECT  5.2925 23.615 5.53 23.68 ;
        RECT  5.0375 23.9725 5.1025 24.1075 ;
        RECT  5.2275 23.9725 5.2925 24.1075 ;
        RECT  5.0375 23.3675 5.1025 23.5025 ;
        RECT  5.2275 23.3675 5.2925 23.5025 ;
        RECT  5.3975 23.2125 5.4625 23.3475 ;
        RECT  5.3975 24.1725 5.4625 24.3075 ;
        RECT  5.005 23.69 5.14 23.755 ;
        RECT  4.97 24.2425 5.53 24.3075 ;
        RECT  4.97 25.5875 5.53 25.6525 ;
        RECT  5.3975 25.3375 5.4625 25.5875 ;
        RECT  5.3975 24.3075 5.4625 24.4425 ;
        RECT  5.0375 24.3075 5.1025 24.3775 ;
        RECT  5.0375 25.4725 5.1025 25.5875 ;
        RECT  5.2275 24.41 5.2925 25.4725 ;
        RECT  4.97 24.87 5.005 24.935 ;
        RECT  5.2925 24.87 5.53 24.935 ;
        RECT  5.0375 24.5125 5.1025 24.6475 ;
        RECT  5.2275 24.5125 5.2925 24.6475 ;
        RECT  5.0375 25.3375 5.1025 25.4725 ;
        RECT  5.2275 25.3375 5.2925 25.4725 ;
        RECT  5.3975 25.3375 5.4625 25.4725 ;
        RECT  5.3975 24.3775 5.4625 24.5125 ;
        RECT  5.005 24.87 5.14 24.935 ;
        RECT  4.97 26.9325 5.53 26.9975 ;
        RECT  4.97 25.5875 5.53 25.6525 ;
        RECT  5.3975 25.6525 5.4625 25.9025 ;
        RECT  5.3975 26.7975 5.4625 26.9325 ;
        RECT  5.0375 26.8625 5.1025 26.9325 ;
        RECT  5.0375 25.6525 5.1025 25.7675 ;
        RECT  5.2275 25.7675 5.2925 26.83 ;
        RECT  4.97 26.305 5.005 26.37 ;
        RECT  5.2925 26.305 5.53 26.37 ;
        RECT  5.0375 26.6625 5.1025 26.7975 ;
        RECT  5.2275 26.6625 5.2925 26.7975 ;
        RECT  5.0375 26.0575 5.1025 26.1925 ;
        RECT  5.2275 26.0575 5.2925 26.1925 ;
        RECT  5.3975 25.9025 5.4625 26.0375 ;
        RECT  5.3975 26.8625 5.4625 26.9975 ;
        RECT  5.005 26.38 5.14 26.445 ;
        RECT  4.97 26.9325 5.53 26.9975 ;
        RECT  4.97 28.2775 5.53 28.3425 ;
        RECT  5.3975 28.0275 5.4625 28.2775 ;
        RECT  5.3975 26.9975 5.4625 27.1325 ;
        RECT  5.0375 26.9975 5.1025 27.0675 ;
        RECT  5.0375 28.1625 5.1025 28.2775 ;
        RECT  5.2275 27.1 5.2925 28.1625 ;
        RECT  4.97 27.56 5.005 27.625 ;
        RECT  5.2925 27.56 5.53 27.625 ;
        RECT  5.0375 27.2025 5.1025 27.3375 ;
        RECT  5.2275 27.2025 5.2925 27.3375 ;
        RECT  5.0375 28.0275 5.1025 28.1625 ;
        RECT  5.2275 28.0275 5.2925 28.1625 ;
        RECT  5.3975 28.0275 5.4625 28.1625 ;
        RECT  5.3975 27.0675 5.4625 27.2025 ;
        RECT  5.005 27.56 5.14 27.625 ;
        RECT  4.97 29.6225 5.53 29.6875 ;
        RECT  4.97 28.2775 5.53 28.3425 ;
        RECT  5.3975 28.3425 5.4625 28.5925 ;
        RECT  5.3975 29.4875 5.4625 29.6225 ;
        RECT  5.0375 29.5525 5.1025 29.6225 ;
        RECT  5.0375 28.3425 5.1025 28.4575 ;
        RECT  5.2275 28.4575 5.2925 29.52 ;
        RECT  4.97 28.995 5.005 29.06 ;
        RECT  5.2925 28.995 5.53 29.06 ;
        RECT  5.0375 29.3525 5.1025 29.4875 ;
        RECT  5.2275 29.3525 5.2925 29.4875 ;
        RECT  5.0375 28.7475 5.1025 28.8825 ;
        RECT  5.2275 28.7475 5.2925 28.8825 ;
        RECT  5.3975 28.5925 5.4625 28.7275 ;
        RECT  5.3975 29.5525 5.4625 29.6875 ;
        RECT  5.005 29.07 5.14 29.135 ;
        RECT  4.97 29.6225 5.53 29.6875 ;
        RECT  4.97 30.9675 5.53 31.0325 ;
        RECT  5.3975 30.7175 5.4625 30.9675 ;
        RECT  5.3975 29.6875 5.4625 29.8225 ;
        RECT  5.0375 29.6875 5.1025 29.7575 ;
        RECT  5.0375 30.8525 5.1025 30.9675 ;
        RECT  5.2275 29.79 5.2925 30.8525 ;
        RECT  4.97 30.25 5.005 30.315 ;
        RECT  5.2925 30.25 5.53 30.315 ;
        RECT  5.0375 29.8925 5.1025 30.0275 ;
        RECT  5.2275 29.8925 5.2925 30.0275 ;
        RECT  5.0375 30.7175 5.1025 30.8525 ;
        RECT  5.2275 30.7175 5.2925 30.8525 ;
        RECT  5.3975 30.7175 5.4625 30.8525 ;
        RECT  5.3975 29.7575 5.4625 29.8925 ;
        RECT  5.005 30.25 5.14 30.315 ;
        RECT  4.97 32.3125 5.53 32.3775 ;
        RECT  4.97 30.9675 5.53 31.0325 ;
        RECT  5.3975 31.0325 5.4625 31.2825 ;
        RECT  5.3975 32.1775 5.4625 32.3125 ;
        RECT  5.0375 32.2425 5.1025 32.3125 ;
        RECT  5.0375 31.0325 5.1025 31.1475 ;
        RECT  5.2275 31.1475 5.2925 32.21 ;
        RECT  4.97 31.685 5.005 31.75 ;
        RECT  5.2925 31.685 5.53 31.75 ;
        RECT  5.0375 32.0425 5.1025 32.1775 ;
        RECT  5.2275 32.0425 5.2925 32.1775 ;
        RECT  5.0375 31.4375 5.1025 31.5725 ;
        RECT  5.2275 31.4375 5.2925 31.5725 ;
        RECT  5.3975 31.2825 5.4625 31.4175 ;
        RECT  5.3975 32.2425 5.4625 32.3775 ;
        RECT  5.005 31.76 5.14 31.825 ;
        RECT  4.97 32.3125 5.53 32.3775 ;
        RECT  4.97 33.6575 5.53 33.7225 ;
        RECT  5.3975 33.4075 5.4625 33.6575 ;
        RECT  5.3975 32.3775 5.4625 32.5125 ;
        RECT  5.0375 32.3775 5.1025 32.4475 ;
        RECT  5.0375 33.5425 5.1025 33.6575 ;
        RECT  5.2275 32.48 5.2925 33.5425 ;
        RECT  4.97 32.94 5.005 33.005 ;
        RECT  5.2925 32.94 5.53 33.005 ;
        RECT  5.0375 32.5825 5.1025 32.7175 ;
        RECT  5.2275 32.5825 5.2925 32.7175 ;
        RECT  5.0375 33.4075 5.1025 33.5425 ;
        RECT  5.2275 33.4075 5.2925 33.5425 ;
        RECT  5.3975 33.4075 5.4625 33.5425 ;
        RECT  5.3975 32.4475 5.4625 32.5825 ;
        RECT  5.005 32.94 5.14 33.005 ;
        RECT  4.97 35.0025 5.53 35.0675 ;
        RECT  4.97 33.6575 5.53 33.7225 ;
        RECT  5.3975 33.7225 5.4625 33.9725 ;
        RECT  5.3975 34.8675 5.4625 35.0025 ;
        RECT  5.0375 34.9325 5.1025 35.0025 ;
        RECT  5.0375 33.7225 5.1025 33.8375 ;
        RECT  5.2275 33.8375 5.2925 34.9 ;
        RECT  4.97 34.375 5.005 34.44 ;
        RECT  5.2925 34.375 5.53 34.44 ;
        RECT  5.0375 34.7325 5.1025 34.8675 ;
        RECT  5.2275 34.7325 5.2925 34.8675 ;
        RECT  5.0375 34.1275 5.1025 34.2625 ;
        RECT  5.2275 34.1275 5.2925 34.2625 ;
        RECT  5.3975 33.9725 5.4625 34.1075 ;
        RECT  5.3975 34.9325 5.4625 35.0675 ;
        RECT  5.005 34.45 5.14 34.515 ;
        RECT  4.97 35.0025 5.53 35.0675 ;
        RECT  4.97 36.3475 5.53 36.4125 ;
        RECT  5.3975 36.0975 5.4625 36.3475 ;
        RECT  5.3975 35.0675 5.4625 35.2025 ;
        RECT  5.0375 35.0675 5.1025 35.1375 ;
        RECT  5.0375 36.2325 5.1025 36.3475 ;
        RECT  5.2275 35.17 5.2925 36.2325 ;
        RECT  4.97 35.63 5.005 35.695 ;
        RECT  5.2925 35.63 5.53 35.695 ;
        RECT  5.0375 35.2725 5.1025 35.4075 ;
        RECT  5.2275 35.2725 5.2925 35.4075 ;
        RECT  5.0375 36.0975 5.1025 36.2325 ;
        RECT  5.2275 36.0975 5.2925 36.2325 ;
        RECT  5.3975 36.0975 5.4625 36.2325 ;
        RECT  5.3975 35.1375 5.4625 35.2725 ;
        RECT  5.005 35.63 5.14 35.695 ;
        RECT  4.97 37.6925 5.53 37.7575 ;
        RECT  4.97 36.3475 5.53 36.4125 ;
        RECT  5.3975 36.4125 5.4625 36.6625 ;
        RECT  5.3975 37.5575 5.4625 37.6925 ;
        RECT  5.0375 37.6225 5.1025 37.6925 ;
        RECT  5.0375 36.4125 5.1025 36.5275 ;
        RECT  5.2275 36.5275 5.2925 37.59 ;
        RECT  4.97 37.065 5.005 37.13 ;
        RECT  5.2925 37.065 5.53 37.13 ;
        RECT  5.0375 37.4225 5.1025 37.5575 ;
        RECT  5.2275 37.4225 5.2925 37.5575 ;
        RECT  5.0375 36.8175 5.1025 36.9525 ;
        RECT  5.2275 36.8175 5.2925 36.9525 ;
        RECT  5.3975 36.6625 5.4625 36.7975 ;
        RECT  5.3975 37.6225 5.4625 37.7575 ;
        RECT  5.005 37.14 5.14 37.205 ;
        RECT  4.97 37.6925 5.53 37.7575 ;
        RECT  4.97 39.0375 5.53 39.1025 ;
        RECT  5.3975 38.7875 5.4625 39.0375 ;
        RECT  5.3975 37.7575 5.4625 37.8925 ;
        RECT  5.0375 37.7575 5.1025 37.8275 ;
        RECT  5.0375 38.9225 5.1025 39.0375 ;
        RECT  5.2275 37.86 5.2925 38.9225 ;
        RECT  4.97 38.32 5.005 38.385 ;
        RECT  5.2925 38.32 5.53 38.385 ;
        RECT  5.0375 37.9625 5.1025 38.0975 ;
        RECT  5.2275 37.9625 5.2925 38.0975 ;
        RECT  5.0375 38.7875 5.1025 38.9225 ;
        RECT  5.2275 38.7875 5.2925 38.9225 ;
        RECT  5.3975 38.7875 5.4625 38.9225 ;
        RECT  5.3975 37.8275 5.4625 37.9625 ;
        RECT  5.005 38.32 5.14 38.385 ;
        RECT  4.97 40.3825 5.53 40.4475 ;
        RECT  4.97 39.0375 5.53 39.1025 ;
        RECT  5.3975 39.1025 5.4625 39.3525 ;
        RECT  5.3975 40.2475 5.4625 40.3825 ;
        RECT  5.0375 40.3125 5.1025 40.3825 ;
        RECT  5.0375 39.1025 5.1025 39.2175 ;
        RECT  5.2275 39.2175 5.2925 40.28 ;
        RECT  4.97 39.755 5.005 39.82 ;
        RECT  5.2925 39.755 5.53 39.82 ;
        RECT  5.0375 40.1125 5.1025 40.2475 ;
        RECT  5.2275 40.1125 5.2925 40.2475 ;
        RECT  5.0375 39.5075 5.1025 39.6425 ;
        RECT  5.2275 39.5075 5.2925 39.6425 ;
        RECT  5.3975 39.3525 5.4625 39.4875 ;
        RECT  5.3975 40.3125 5.4625 40.4475 ;
        RECT  5.005 39.83 5.14 39.895 ;
        RECT  2.79 8.73 2.925 8.795 ;
        RECT  2.965 10.165 3.1 10.23 ;
        RECT  3.14 11.42 3.275 11.485 ;
        RECT  3.315 12.855 3.45 12.92 ;
        RECT  3.49 14.11 3.625 14.175 ;
        RECT  3.665 15.545 3.8 15.61 ;
        RECT  3.84 16.8 3.975 16.865 ;
        RECT  4.015 18.235 4.15 18.3 ;
        RECT  2.79 19.805 2.925 19.87 ;
        RECT  3.49 19.275 3.625 19.34 ;
        RECT  2.79 20.61 2.925 20.675 ;
        RECT  3.665 21.14 3.8 21.205 ;
        RECT  2.79 22.495 2.925 22.56 ;
        RECT  3.84 21.965 3.975 22.03 ;
        RECT  2.79 23.3 2.925 23.365 ;
        RECT  4.015 23.83 4.15 23.895 ;
        RECT  2.965 25.185 3.1 25.25 ;
        RECT  3.49 24.655 3.625 24.72 ;
        RECT  2.965 25.99 3.1 26.055 ;
        RECT  3.665 26.52 3.8 26.585 ;
        RECT  2.965 27.875 3.1 27.94 ;
        RECT  3.84 27.345 3.975 27.41 ;
        RECT  2.965 28.68 3.1 28.745 ;
        RECT  4.015 29.21 4.15 29.275 ;
        RECT  3.14 30.565 3.275 30.63 ;
        RECT  3.49 30.035 3.625 30.1 ;
        RECT  3.14 31.37 3.275 31.435 ;
        RECT  3.665 31.9 3.8 31.965 ;
        RECT  3.14 33.255 3.275 33.32 ;
        RECT  3.84 32.725 3.975 32.79 ;
        RECT  3.14 34.06 3.275 34.125 ;
        RECT  4.015 34.59 4.15 34.655 ;
        RECT  3.315 35.945 3.45 36.01 ;
        RECT  3.49 35.415 3.625 35.48 ;
        RECT  3.315 36.75 3.45 36.815 ;
        RECT  3.665 37.28 3.8 37.345 ;
        RECT  3.315 38.635 3.45 38.7 ;
        RECT  3.84 38.105 3.975 38.17 ;
        RECT  3.315 39.44 3.45 39.505 ;
        RECT  4.015 39.97 4.15 40.035 ;
        RECT  5.725 19.025 5.79 40.805 ;
        RECT  5.725 19.445 6.05 19.51 ;
        RECT  6.48 19.275 6.545 19.51 ;
        RECT  7.295 19.4925 7.36 19.5575 ;
        RECT  7.855 19.445 7.92 19.51 ;
        RECT  5.725 20.97 6.05 21.035 ;
        RECT  6.48 20.97 6.545 21.205 ;
        RECT  7.295 20.9225 7.36 20.9875 ;
        RECT  7.79 20.97 7.855 21.035 ;
        RECT  5.725 22.135 6.05 22.2 ;
        RECT  6.48 21.965 6.545 22.2 ;
        RECT  7.295 22.1825 7.36 22.2475 ;
        RECT  7.855 22.135 7.92 22.2 ;
        RECT  5.725 23.66 6.05 23.725 ;
        RECT  6.48 23.66 6.545 23.895 ;
        RECT  7.295 23.6125 7.36 23.6775 ;
        RECT  7.79 23.66 7.855 23.725 ;
        RECT  5.725 24.825 6.05 24.89 ;
        RECT  6.48 24.655 6.545 24.89 ;
        RECT  7.295 24.8725 7.36 24.9375 ;
        RECT  7.855 24.825 7.92 24.89 ;
        RECT  5.725 26.35 6.05 26.415 ;
        RECT  6.48 26.35 6.545 26.585 ;
        RECT  7.295 26.3025 7.36 26.3675 ;
        RECT  7.79 26.35 7.855 26.415 ;
        RECT  5.725 27.515 6.05 27.58 ;
        RECT  6.48 27.345 6.545 27.58 ;
        RECT  7.295 27.5625 7.36 27.6275 ;
        RECT  7.855 27.515 7.92 27.58 ;
        RECT  5.725 29.04 6.05 29.105 ;
        RECT  6.48 29.04 6.545 29.275 ;
        RECT  7.295 28.9925 7.36 29.0575 ;
        RECT  7.79 29.04 7.855 29.105 ;
        RECT  5.725 30.205 6.05 30.27 ;
        RECT  6.48 30.035 6.545 30.27 ;
        RECT  7.295 30.2525 7.36 30.3175 ;
        RECT  7.855 30.205 7.92 30.27 ;
        RECT  5.725 31.73 6.05 31.795 ;
        RECT  6.48 31.73 6.545 31.965 ;
        RECT  7.295 31.6825 7.36 31.7475 ;
        RECT  7.79 31.73 7.855 31.795 ;
        RECT  5.725 32.895 6.05 32.96 ;
        RECT  6.48 32.725 6.545 32.96 ;
        RECT  7.295 32.9425 7.36 33.0075 ;
        RECT  7.855 32.895 7.92 32.96 ;
        RECT  5.725 34.42 6.05 34.485 ;
        RECT  6.48 34.42 6.545 34.655 ;
        RECT  7.295 34.3725 7.36 34.4375 ;
        RECT  7.79 34.42 7.855 34.485 ;
        RECT  5.725 35.585 6.05 35.65 ;
        RECT  6.48 35.415 6.545 35.65 ;
        RECT  7.295 35.6325 7.36 35.6975 ;
        RECT  7.855 35.585 7.92 35.65 ;
        RECT  5.725 37.11 6.05 37.175 ;
        RECT  6.48 37.11 6.545 37.345 ;
        RECT  7.295 37.0625 7.36 37.1275 ;
        RECT  7.79 37.11 7.855 37.175 ;
        RECT  5.725 38.275 6.05 38.34 ;
        RECT  6.48 38.105 6.545 38.34 ;
        RECT  7.295 38.3225 7.36 38.3875 ;
        RECT  7.855 38.275 7.92 38.34 ;
        RECT  5.725 39.8 6.05 39.865 ;
        RECT  6.48 39.8 6.545 40.035 ;
        RECT  7.295 39.7525 7.36 39.8175 ;
        RECT  7.79 39.8 7.855 39.865 ;
        RECT  5.46 20.2075 5.595 20.2725 ;
        RECT  5.915 20.2075 6.05 20.2725 ;
        RECT  5.985 18.8625 6.545 18.9275 ;
        RECT  5.985 20.2075 6.545 20.2725 ;
        RECT  6.4125 19.9575 6.4775 20.2075 ;
        RECT  6.4125 18.9275 6.4775 19.0625 ;
        RECT  6.0525 18.9275 6.1175 18.9975 ;
        RECT  6.0525 20.0925 6.1175 20.2075 ;
        RECT  6.2425 19.03 6.3075 20.0925 ;
        RECT  5.985 19.49 6.02 19.555 ;
        RECT  6.3075 19.49 6.545 19.555 ;
        RECT  6.0525 19.1325 6.1175 19.2675 ;
        RECT  6.2425 19.1325 6.3075 19.2675 ;
        RECT  6.0525 19.9575 6.1175 20.0925 ;
        RECT  6.2425 19.9575 6.3075 20.0925 ;
        RECT  6.4125 19.9575 6.4775 20.0925 ;
        RECT  6.4125 18.9975 6.4775 19.1325 ;
        RECT  6.02 19.49 6.155 19.555 ;
        RECT  6.545 18.8625 7.295 18.9275 ;
        RECT  6.545 20.2075 7.295 20.2725 ;
        RECT  7.1625 19.9575 7.2275 20.24 ;
        RECT  7.1625 18.895 7.2275 19.075 ;
        RECT  6.6125 19.9575 6.6775 20.24 ;
        RECT  6.9925 19.9575 7.0575 20.24 ;
        RECT  6.6125 18.895 6.6775 19.1775 ;
        RECT  6.545 19.805 6.58 19.87 ;
        RECT  6.545 19.275 6.82 19.34 ;
        RECT  7.0575 19.4925 7.295 19.5575 ;
        RECT  6.6125 19.1775 6.6775 19.3125 ;
        RECT  6.8025 19.1775 6.8675 19.3125 ;
        RECT  6.8025 19.1775 6.8675 19.3125 ;
        RECT  6.9925 19.1775 7.0575 19.3125 ;
        RECT  6.6125 19.9575 6.6775 20.0925 ;
        RECT  6.8025 19.9575 6.8675 20.0925 ;
        RECT  6.8025 19.9575 6.8675 20.0925 ;
        RECT  6.9925 19.9575 7.0575 20.0925 ;
        RECT  7.1625 19.9575 7.2275 20.0925 ;
        RECT  7.1625 19.0425 7.2275 19.1775 ;
        RECT  7.025 19.79 7.09 19.855 ;
        RECT  6.8025 19.79 6.8675 19.855 ;
        RECT  7.025 19.0425 7.09 19.8225 ;
        RECT  6.835 19.79 7.0575 19.855 ;
        RECT  6.8025 19.8225 6.8675 19.9575 ;
        RECT  6.58 19.805 6.715 19.87 ;
        RECT  6.82 19.275 6.955 19.34 ;
        RECT  7.295 18.8625 7.855 18.9275 ;
        RECT  7.295 20.2075 7.855 20.2725 ;
        RECT  7.7225 19.9575 7.7875 20.2075 ;
        RECT  7.7225 18.9275 7.7875 19.0625 ;
        RECT  7.3625 18.9275 7.4275 18.9975 ;
        RECT  7.3625 20.0925 7.4275 20.2075 ;
        RECT  7.5525 19.03 7.6175 20.0925 ;
        RECT  7.295 19.49 7.33 19.555 ;
        RECT  7.6175 19.49 7.855 19.555 ;
        RECT  7.3625 19.1325 7.4275 19.2675 ;
        RECT  7.5525 19.1325 7.6175 19.2675 ;
        RECT  7.3625 19.9575 7.4275 20.0925 ;
        RECT  7.5525 19.9575 7.6175 20.0925 ;
        RECT  7.7225 19.9575 7.7875 20.0925 ;
        RECT  7.7225 18.9975 7.7875 19.1325 ;
        RECT  7.33 19.49 7.465 19.555 ;
        RECT  6.545 19.8075 6.68 19.8725 ;
        RECT  5.5325 19.805 5.5975 19.94 ;
        RECT  5.46 21.5525 5.595 21.6175 ;
        RECT  5.915 21.5525 6.05 21.6175 ;
        RECT  5.985 21.5525 6.545 21.6175 ;
        RECT  5.985 20.2075 6.545 20.2725 ;
        RECT  6.4125 20.2725 6.4775 20.5225 ;
        RECT  6.4125 21.4175 6.4775 21.5525 ;
        RECT  6.0525 21.4825 6.1175 21.5525 ;
        RECT  6.0525 20.2725 6.1175 20.3875 ;
        RECT  6.2425 20.3875 6.3075 21.45 ;
        RECT  5.985 20.925 6.02 20.99 ;
        RECT  6.3075 20.925 6.545 20.99 ;
        RECT  6.0525 21.2825 6.1175 21.4175 ;
        RECT  6.2425 21.2825 6.3075 21.4175 ;
        RECT  6.0525 20.6775 6.1175 20.8125 ;
        RECT  6.2425 20.6775 6.3075 20.8125 ;
        RECT  6.4125 20.5225 6.4775 20.6575 ;
        RECT  6.4125 21.4825 6.4775 21.6175 ;
        RECT  6.02 21.0 6.155 21.065 ;
        RECT  6.545 21.5525 7.295 21.6175 ;
        RECT  6.545 20.2075 7.295 20.2725 ;
        RECT  7.1625 20.24 7.2275 20.5225 ;
        RECT  7.1625 21.405 7.2275 21.585 ;
        RECT  6.6125 20.24 6.6775 20.5225 ;
        RECT  6.9925 20.24 7.0575 20.5225 ;
        RECT  6.6125 21.3025 6.6775 21.585 ;
        RECT  6.545 20.61 6.58 20.675 ;
        RECT  6.545 21.14 6.82 21.205 ;
        RECT  7.0575 20.9225 7.295 20.9875 ;
        RECT  6.6125 21.1475 6.6775 21.2825 ;
        RECT  6.8025 21.1475 6.8675 21.2825 ;
        RECT  6.8025 21.1475 6.8675 21.2825 ;
        RECT  6.9925 21.1475 7.0575 21.2825 ;
        RECT  6.6125 20.6775 6.6775 20.8125 ;
        RECT  6.8025 20.6775 6.8675 20.8125 ;
        RECT  6.8025 20.6775 6.8675 20.8125 ;
        RECT  6.9925 20.6775 7.0575 20.8125 ;
        RECT  7.1625 20.5225 7.2275 20.6575 ;
        RECT  7.1625 21.4375 7.2275 21.5725 ;
        RECT  7.025 22.185 7.09 22.25 ;
        RECT  6.8025 22.185 6.8675 22.25 ;
        RECT  7.025 21.4375 7.09 22.2175 ;
        RECT  6.835 22.185 7.0575 22.25 ;
        RECT  6.8025 22.2175 6.8675 22.3525 ;
        RECT  6.58 20.685 6.715 20.75 ;
        RECT  6.82 21.215 6.955 21.28 ;
        RECT  7.295 21.5525 7.855 21.6175 ;
        RECT  7.295 20.2075 7.855 20.2725 ;
        RECT  7.7225 20.2725 7.7875 20.5225 ;
        RECT  7.7225 21.4175 7.7875 21.5525 ;
        RECT  7.3625 21.4825 7.4275 21.5525 ;
        RECT  7.3625 20.2725 7.4275 20.3875 ;
        RECT  7.5525 20.3875 7.6175 21.45 ;
        RECT  7.295 20.925 7.33 20.99 ;
        RECT  7.6175 20.925 7.855 20.99 ;
        RECT  7.3625 21.2825 7.4275 21.4175 ;
        RECT  7.5525 21.2825 7.6175 21.4175 ;
        RECT  7.3625 20.6775 7.4275 20.8125 ;
        RECT  7.5525 20.6775 7.6175 20.8125 ;
        RECT  7.7225 20.5225 7.7875 20.6575 ;
        RECT  7.7225 21.4825 7.7875 21.6175 ;
        RECT  7.33 21.0 7.465 21.065 ;
        RECT  6.545 20.6075 6.68 20.6725 ;
        RECT  5.5325 20.54 5.5975 20.675 ;
        RECT  5.46 22.8975 5.595 22.9625 ;
        RECT  5.915 22.8975 6.05 22.9625 ;
        RECT  5.985 21.5525 6.545 21.6175 ;
        RECT  5.985 22.8975 6.545 22.9625 ;
        RECT  6.4125 22.6475 6.4775 22.8975 ;
        RECT  6.4125 21.6175 6.4775 21.7525 ;
        RECT  6.0525 21.6175 6.1175 21.6875 ;
        RECT  6.0525 22.7825 6.1175 22.8975 ;
        RECT  6.2425 21.72 6.3075 22.7825 ;
        RECT  5.985 22.18 6.02 22.245 ;
        RECT  6.3075 22.18 6.545 22.245 ;
        RECT  6.0525 21.8225 6.1175 21.9575 ;
        RECT  6.2425 21.8225 6.3075 21.9575 ;
        RECT  6.0525 22.6475 6.1175 22.7825 ;
        RECT  6.2425 22.6475 6.3075 22.7825 ;
        RECT  6.4125 22.6475 6.4775 22.7825 ;
        RECT  6.4125 21.6875 6.4775 21.8225 ;
        RECT  6.02 22.18 6.155 22.245 ;
        RECT  6.545 21.5525 7.295 21.6175 ;
        RECT  6.545 22.8975 7.295 22.9625 ;
        RECT  7.1625 22.6475 7.2275 22.93 ;
        RECT  7.1625 21.585 7.2275 21.765 ;
        RECT  6.6125 22.6475 6.6775 22.93 ;
        RECT  6.9925 22.6475 7.0575 22.93 ;
        RECT  6.6125 21.585 6.6775 21.8675 ;
        RECT  6.545 22.495 6.58 22.56 ;
        RECT  6.545 21.965 6.82 22.03 ;
        RECT  7.0575 22.1825 7.295 22.2475 ;
        RECT  6.6125 21.8675 6.6775 22.0025 ;
        RECT  6.8025 21.8675 6.8675 22.0025 ;
        RECT  6.8025 21.8675 6.8675 22.0025 ;
        RECT  6.9925 21.8675 7.0575 22.0025 ;
        RECT  6.6125 22.6475 6.6775 22.7825 ;
        RECT  6.8025 22.6475 6.8675 22.7825 ;
        RECT  6.8025 22.6475 6.8675 22.7825 ;
        RECT  6.9925 22.6475 7.0575 22.7825 ;
        RECT  7.1625 22.6475 7.2275 22.7825 ;
        RECT  7.1625 21.7325 7.2275 21.8675 ;
        RECT  7.025 22.48 7.09 22.545 ;
        RECT  6.8025 22.48 6.8675 22.545 ;
        RECT  7.025 21.7325 7.09 22.5125 ;
        RECT  6.835 22.48 7.0575 22.545 ;
        RECT  6.8025 22.5125 6.8675 22.6475 ;
        RECT  6.58 22.495 6.715 22.56 ;
        RECT  6.82 21.965 6.955 22.03 ;
        RECT  7.295 21.5525 7.855 21.6175 ;
        RECT  7.295 22.8975 7.855 22.9625 ;
        RECT  7.7225 22.6475 7.7875 22.8975 ;
        RECT  7.7225 21.6175 7.7875 21.7525 ;
        RECT  7.3625 21.6175 7.4275 21.6875 ;
        RECT  7.3625 22.7825 7.4275 22.8975 ;
        RECT  7.5525 21.72 7.6175 22.7825 ;
        RECT  7.295 22.18 7.33 22.245 ;
        RECT  7.6175 22.18 7.855 22.245 ;
        RECT  7.3625 21.8225 7.4275 21.9575 ;
        RECT  7.5525 21.8225 7.6175 21.9575 ;
        RECT  7.3625 22.6475 7.4275 22.7825 ;
        RECT  7.5525 22.6475 7.6175 22.7825 ;
        RECT  7.7225 22.6475 7.7875 22.7825 ;
        RECT  7.7225 21.6875 7.7875 21.8225 ;
        RECT  7.33 22.18 7.465 22.245 ;
        RECT  6.545 22.4975 6.68 22.5625 ;
        RECT  5.5325 22.495 5.5975 22.63 ;
        RECT  5.46 24.2425 5.595 24.3075 ;
        RECT  5.915 24.2425 6.05 24.3075 ;
        RECT  5.985 24.2425 6.545 24.3075 ;
        RECT  5.985 22.8975 6.545 22.9625 ;
        RECT  6.4125 22.9625 6.4775 23.2125 ;
        RECT  6.4125 24.1075 6.4775 24.2425 ;
        RECT  6.0525 24.1725 6.1175 24.2425 ;
        RECT  6.0525 22.9625 6.1175 23.0775 ;
        RECT  6.2425 23.0775 6.3075 24.14 ;
        RECT  5.985 23.615 6.02 23.68 ;
        RECT  6.3075 23.615 6.545 23.68 ;
        RECT  6.0525 23.9725 6.1175 24.1075 ;
        RECT  6.2425 23.9725 6.3075 24.1075 ;
        RECT  6.0525 23.3675 6.1175 23.5025 ;
        RECT  6.2425 23.3675 6.3075 23.5025 ;
        RECT  6.4125 23.2125 6.4775 23.3475 ;
        RECT  6.4125 24.1725 6.4775 24.3075 ;
        RECT  6.02 23.69 6.155 23.755 ;
        RECT  6.545 24.2425 7.295 24.3075 ;
        RECT  6.545 22.8975 7.295 22.9625 ;
        RECT  7.1625 22.93 7.2275 23.2125 ;
        RECT  7.1625 24.095 7.2275 24.275 ;
        RECT  6.6125 22.93 6.6775 23.2125 ;
        RECT  6.9925 22.93 7.0575 23.2125 ;
        RECT  6.6125 23.9925 6.6775 24.275 ;
        RECT  6.545 23.3 6.58 23.365 ;
        RECT  6.545 23.83 6.82 23.895 ;
        RECT  7.0575 23.6125 7.295 23.6775 ;
        RECT  6.6125 23.8375 6.6775 23.9725 ;
        RECT  6.8025 23.8375 6.8675 23.9725 ;
        RECT  6.8025 23.8375 6.8675 23.9725 ;
        RECT  6.9925 23.8375 7.0575 23.9725 ;
        RECT  6.6125 23.3675 6.6775 23.5025 ;
        RECT  6.8025 23.3675 6.8675 23.5025 ;
        RECT  6.8025 23.3675 6.8675 23.5025 ;
        RECT  6.9925 23.3675 7.0575 23.5025 ;
        RECT  7.1625 23.2125 7.2275 23.3475 ;
        RECT  7.1625 24.1275 7.2275 24.2625 ;
        RECT  7.025 24.875 7.09 24.94 ;
        RECT  6.8025 24.875 6.8675 24.94 ;
        RECT  7.025 24.1275 7.09 24.9075 ;
        RECT  6.835 24.875 7.0575 24.94 ;
        RECT  6.8025 24.9075 6.8675 25.0425 ;
        RECT  6.58 23.375 6.715 23.44 ;
        RECT  6.82 23.905 6.955 23.97 ;
        RECT  7.295 24.2425 7.855 24.3075 ;
        RECT  7.295 22.8975 7.855 22.9625 ;
        RECT  7.7225 22.9625 7.7875 23.2125 ;
        RECT  7.7225 24.1075 7.7875 24.2425 ;
        RECT  7.3625 24.1725 7.4275 24.2425 ;
        RECT  7.3625 22.9625 7.4275 23.0775 ;
        RECT  7.5525 23.0775 7.6175 24.14 ;
        RECT  7.295 23.615 7.33 23.68 ;
        RECT  7.6175 23.615 7.855 23.68 ;
        RECT  7.3625 23.9725 7.4275 24.1075 ;
        RECT  7.5525 23.9725 7.6175 24.1075 ;
        RECT  7.3625 23.3675 7.4275 23.5025 ;
        RECT  7.5525 23.3675 7.6175 23.5025 ;
        RECT  7.7225 23.2125 7.7875 23.3475 ;
        RECT  7.7225 24.1725 7.7875 24.3075 ;
        RECT  7.33 23.69 7.465 23.755 ;
        RECT  6.545 23.2975 6.68 23.3625 ;
        RECT  5.5325 23.23 5.5975 23.365 ;
        RECT  5.46 25.5875 5.595 25.6525 ;
        RECT  5.915 25.5875 6.05 25.6525 ;
        RECT  5.985 24.2425 6.545 24.3075 ;
        RECT  5.985 25.5875 6.545 25.6525 ;
        RECT  6.4125 25.3375 6.4775 25.5875 ;
        RECT  6.4125 24.3075 6.4775 24.4425 ;
        RECT  6.0525 24.3075 6.1175 24.3775 ;
        RECT  6.0525 25.4725 6.1175 25.5875 ;
        RECT  6.2425 24.41 6.3075 25.4725 ;
        RECT  5.985 24.87 6.02 24.935 ;
        RECT  6.3075 24.87 6.545 24.935 ;
        RECT  6.0525 24.5125 6.1175 24.6475 ;
        RECT  6.2425 24.5125 6.3075 24.6475 ;
        RECT  6.0525 25.3375 6.1175 25.4725 ;
        RECT  6.2425 25.3375 6.3075 25.4725 ;
        RECT  6.4125 25.3375 6.4775 25.4725 ;
        RECT  6.4125 24.3775 6.4775 24.5125 ;
        RECT  6.02 24.87 6.155 24.935 ;
        RECT  6.545 24.2425 7.295 24.3075 ;
        RECT  6.545 25.5875 7.295 25.6525 ;
        RECT  7.1625 25.3375 7.2275 25.62 ;
        RECT  7.1625 24.275 7.2275 24.455 ;
        RECT  6.6125 25.3375 6.6775 25.62 ;
        RECT  6.9925 25.3375 7.0575 25.62 ;
        RECT  6.6125 24.275 6.6775 24.5575 ;
        RECT  6.545 25.185 6.58 25.25 ;
        RECT  6.545 24.655 6.82 24.72 ;
        RECT  7.0575 24.8725 7.295 24.9375 ;
        RECT  6.6125 24.5575 6.6775 24.6925 ;
        RECT  6.8025 24.5575 6.8675 24.6925 ;
        RECT  6.8025 24.5575 6.8675 24.6925 ;
        RECT  6.9925 24.5575 7.0575 24.6925 ;
        RECT  6.6125 25.3375 6.6775 25.4725 ;
        RECT  6.8025 25.3375 6.8675 25.4725 ;
        RECT  6.8025 25.3375 6.8675 25.4725 ;
        RECT  6.9925 25.3375 7.0575 25.4725 ;
        RECT  7.1625 25.3375 7.2275 25.4725 ;
        RECT  7.1625 24.4225 7.2275 24.5575 ;
        RECT  7.025 25.17 7.09 25.235 ;
        RECT  6.8025 25.17 6.8675 25.235 ;
        RECT  7.025 24.4225 7.09 25.2025 ;
        RECT  6.835 25.17 7.0575 25.235 ;
        RECT  6.8025 25.2025 6.8675 25.3375 ;
        RECT  6.58 25.185 6.715 25.25 ;
        RECT  6.82 24.655 6.955 24.72 ;
        RECT  7.295 24.2425 7.855 24.3075 ;
        RECT  7.295 25.5875 7.855 25.6525 ;
        RECT  7.7225 25.3375 7.7875 25.5875 ;
        RECT  7.7225 24.3075 7.7875 24.4425 ;
        RECT  7.3625 24.3075 7.4275 24.3775 ;
        RECT  7.3625 25.4725 7.4275 25.5875 ;
        RECT  7.5525 24.41 7.6175 25.4725 ;
        RECT  7.295 24.87 7.33 24.935 ;
        RECT  7.6175 24.87 7.855 24.935 ;
        RECT  7.3625 24.5125 7.4275 24.6475 ;
        RECT  7.5525 24.5125 7.6175 24.6475 ;
        RECT  7.3625 25.3375 7.4275 25.4725 ;
        RECT  7.5525 25.3375 7.6175 25.4725 ;
        RECT  7.7225 25.3375 7.7875 25.4725 ;
        RECT  7.7225 24.3775 7.7875 24.5125 ;
        RECT  7.33 24.87 7.465 24.935 ;
        RECT  6.545 25.1875 6.68 25.2525 ;
        RECT  5.5325 25.185 5.5975 25.32 ;
        RECT  5.46 26.9325 5.595 26.9975 ;
        RECT  5.915 26.9325 6.05 26.9975 ;
        RECT  5.985 26.9325 6.545 26.9975 ;
        RECT  5.985 25.5875 6.545 25.6525 ;
        RECT  6.4125 25.6525 6.4775 25.9025 ;
        RECT  6.4125 26.7975 6.4775 26.9325 ;
        RECT  6.0525 26.8625 6.1175 26.9325 ;
        RECT  6.0525 25.6525 6.1175 25.7675 ;
        RECT  6.2425 25.7675 6.3075 26.83 ;
        RECT  5.985 26.305 6.02 26.37 ;
        RECT  6.3075 26.305 6.545 26.37 ;
        RECT  6.0525 26.6625 6.1175 26.7975 ;
        RECT  6.2425 26.6625 6.3075 26.7975 ;
        RECT  6.0525 26.0575 6.1175 26.1925 ;
        RECT  6.2425 26.0575 6.3075 26.1925 ;
        RECT  6.4125 25.9025 6.4775 26.0375 ;
        RECT  6.4125 26.8625 6.4775 26.9975 ;
        RECT  6.02 26.38 6.155 26.445 ;
        RECT  6.545 26.9325 7.295 26.9975 ;
        RECT  6.545 25.5875 7.295 25.6525 ;
        RECT  7.1625 25.62 7.2275 25.9025 ;
        RECT  7.1625 26.785 7.2275 26.965 ;
        RECT  6.6125 25.62 6.6775 25.9025 ;
        RECT  6.9925 25.62 7.0575 25.9025 ;
        RECT  6.6125 26.6825 6.6775 26.965 ;
        RECT  6.545 25.99 6.58 26.055 ;
        RECT  6.545 26.52 6.82 26.585 ;
        RECT  7.0575 26.3025 7.295 26.3675 ;
        RECT  6.6125 26.5275 6.6775 26.6625 ;
        RECT  6.8025 26.5275 6.8675 26.6625 ;
        RECT  6.8025 26.5275 6.8675 26.6625 ;
        RECT  6.9925 26.5275 7.0575 26.6625 ;
        RECT  6.6125 26.0575 6.6775 26.1925 ;
        RECT  6.8025 26.0575 6.8675 26.1925 ;
        RECT  6.8025 26.0575 6.8675 26.1925 ;
        RECT  6.9925 26.0575 7.0575 26.1925 ;
        RECT  7.1625 25.9025 7.2275 26.0375 ;
        RECT  7.1625 26.8175 7.2275 26.9525 ;
        RECT  7.025 27.565 7.09 27.63 ;
        RECT  6.8025 27.565 6.8675 27.63 ;
        RECT  7.025 26.8175 7.09 27.5975 ;
        RECT  6.835 27.565 7.0575 27.63 ;
        RECT  6.8025 27.5975 6.8675 27.7325 ;
        RECT  6.58 26.065 6.715 26.13 ;
        RECT  6.82 26.595 6.955 26.66 ;
        RECT  7.295 26.9325 7.855 26.9975 ;
        RECT  7.295 25.5875 7.855 25.6525 ;
        RECT  7.7225 25.6525 7.7875 25.9025 ;
        RECT  7.7225 26.7975 7.7875 26.9325 ;
        RECT  7.3625 26.8625 7.4275 26.9325 ;
        RECT  7.3625 25.6525 7.4275 25.7675 ;
        RECT  7.5525 25.7675 7.6175 26.83 ;
        RECT  7.295 26.305 7.33 26.37 ;
        RECT  7.6175 26.305 7.855 26.37 ;
        RECT  7.3625 26.6625 7.4275 26.7975 ;
        RECT  7.5525 26.6625 7.6175 26.7975 ;
        RECT  7.3625 26.0575 7.4275 26.1925 ;
        RECT  7.5525 26.0575 7.6175 26.1925 ;
        RECT  7.7225 25.9025 7.7875 26.0375 ;
        RECT  7.7225 26.8625 7.7875 26.9975 ;
        RECT  7.33 26.38 7.465 26.445 ;
        RECT  6.545 25.9875 6.68 26.0525 ;
        RECT  5.5325 25.92 5.5975 26.055 ;
        RECT  5.46 28.2775 5.595 28.3425 ;
        RECT  5.915 28.2775 6.05 28.3425 ;
        RECT  5.985 26.9325 6.545 26.9975 ;
        RECT  5.985 28.2775 6.545 28.3425 ;
        RECT  6.4125 28.0275 6.4775 28.2775 ;
        RECT  6.4125 26.9975 6.4775 27.1325 ;
        RECT  6.0525 26.9975 6.1175 27.0675 ;
        RECT  6.0525 28.1625 6.1175 28.2775 ;
        RECT  6.2425 27.1 6.3075 28.1625 ;
        RECT  5.985 27.56 6.02 27.625 ;
        RECT  6.3075 27.56 6.545 27.625 ;
        RECT  6.0525 27.2025 6.1175 27.3375 ;
        RECT  6.2425 27.2025 6.3075 27.3375 ;
        RECT  6.0525 28.0275 6.1175 28.1625 ;
        RECT  6.2425 28.0275 6.3075 28.1625 ;
        RECT  6.4125 28.0275 6.4775 28.1625 ;
        RECT  6.4125 27.0675 6.4775 27.2025 ;
        RECT  6.02 27.56 6.155 27.625 ;
        RECT  6.545 26.9325 7.295 26.9975 ;
        RECT  6.545 28.2775 7.295 28.3425 ;
        RECT  7.1625 28.0275 7.2275 28.31 ;
        RECT  7.1625 26.965 7.2275 27.145 ;
        RECT  6.6125 28.0275 6.6775 28.31 ;
        RECT  6.9925 28.0275 7.0575 28.31 ;
        RECT  6.6125 26.965 6.6775 27.2475 ;
        RECT  6.545 27.875 6.58 27.94 ;
        RECT  6.545 27.345 6.82 27.41 ;
        RECT  7.0575 27.5625 7.295 27.6275 ;
        RECT  6.6125 27.2475 6.6775 27.3825 ;
        RECT  6.8025 27.2475 6.8675 27.3825 ;
        RECT  6.8025 27.2475 6.8675 27.3825 ;
        RECT  6.9925 27.2475 7.0575 27.3825 ;
        RECT  6.6125 28.0275 6.6775 28.1625 ;
        RECT  6.8025 28.0275 6.8675 28.1625 ;
        RECT  6.8025 28.0275 6.8675 28.1625 ;
        RECT  6.9925 28.0275 7.0575 28.1625 ;
        RECT  7.1625 28.0275 7.2275 28.1625 ;
        RECT  7.1625 27.1125 7.2275 27.2475 ;
        RECT  7.025 27.86 7.09 27.925 ;
        RECT  6.8025 27.86 6.8675 27.925 ;
        RECT  7.025 27.1125 7.09 27.8925 ;
        RECT  6.835 27.86 7.0575 27.925 ;
        RECT  6.8025 27.8925 6.8675 28.0275 ;
        RECT  6.58 27.875 6.715 27.94 ;
        RECT  6.82 27.345 6.955 27.41 ;
        RECT  7.295 26.9325 7.855 26.9975 ;
        RECT  7.295 28.2775 7.855 28.3425 ;
        RECT  7.7225 28.0275 7.7875 28.2775 ;
        RECT  7.7225 26.9975 7.7875 27.1325 ;
        RECT  7.3625 26.9975 7.4275 27.0675 ;
        RECT  7.3625 28.1625 7.4275 28.2775 ;
        RECT  7.5525 27.1 7.6175 28.1625 ;
        RECT  7.295 27.56 7.33 27.625 ;
        RECT  7.6175 27.56 7.855 27.625 ;
        RECT  7.3625 27.2025 7.4275 27.3375 ;
        RECT  7.5525 27.2025 7.6175 27.3375 ;
        RECT  7.3625 28.0275 7.4275 28.1625 ;
        RECT  7.5525 28.0275 7.6175 28.1625 ;
        RECT  7.7225 28.0275 7.7875 28.1625 ;
        RECT  7.7225 27.0675 7.7875 27.2025 ;
        RECT  7.33 27.56 7.465 27.625 ;
        RECT  6.545 27.8775 6.68 27.9425 ;
        RECT  5.5325 27.875 5.5975 28.01 ;
        RECT  5.46 29.6225 5.595 29.6875 ;
        RECT  5.915 29.6225 6.05 29.6875 ;
        RECT  5.985 29.6225 6.545 29.6875 ;
        RECT  5.985 28.2775 6.545 28.3425 ;
        RECT  6.4125 28.3425 6.4775 28.5925 ;
        RECT  6.4125 29.4875 6.4775 29.6225 ;
        RECT  6.0525 29.5525 6.1175 29.6225 ;
        RECT  6.0525 28.3425 6.1175 28.4575 ;
        RECT  6.2425 28.4575 6.3075 29.52 ;
        RECT  5.985 28.995 6.02 29.06 ;
        RECT  6.3075 28.995 6.545 29.06 ;
        RECT  6.0525 29.3525 6.1175 29.4875 ;
        RECT  6.2425 29.3525 6.3075 29.4875 ;
        RECT  6.0525 28.7475 6.1175 28.8825 ;
        RECT  6.2425 28.7475 6.3075 28.8825 ;
        RECT  6.4125 28.5925 6.4775 28.7275 ;
        RECT  6.4125 29.5525 6.4775 29.6875 ;
        RECT  6.02 29.07 6.155 29.135 ;
        RECT  6.545 29.6225 7.295 29.6875 ;
        RECT  6.545 28.2775 7.295 28.3425 ;
        RECT  7.1625 28.31 7.2275 28.5925 ;
        RECT  7.1625 29.475 7.2275 29.655 ;
        RECT  6.6125 28.31 6.6775 28.5925 ;
        RECT  6.9925 28.31 7.0575 28.5925 ;
        RECT  6.6125 29.3725 6.6775 29.655 ;
        RECT  6.545 28.68 6.58 28.745 ;
        RECT  6.545 29.21 6.82 29.275 ;
        RECT  7.0575 28.9925 7.295 29.0575 ;
        RECT  6.6125 29.2175 6.6775 29.3525 ;
        RECT  6.8025 29.2175 6.8675 29.3525 ;
        RECT  6.8025 29.2175 6.8675 29.3525 ;
        RECT  6.9925 29.2175 7.0575 29.3525 ;
        RECT  6.6125 28.7475 6.6775 28.8825 ;
        RECT  6.8025 28.7475 6.8675 28.8825 ;
        RECT  6.8025 28.7475 6.8675 28.8825 ;
        RECT  6.9925 28.7475 7.0575 28.8825 ;
        RECT  7.1625 28.5925 7.2275 28.7275 ;
        RECT  7.1625 29.5075 7.2275 29.6425 ;
        RECT  7.025 30.255 7.09 30.32 ;
        RECT  6.8025 30.255 6.8675 30.32 ;
        RECT  7.025 29.5075 7.09 30.2875 ;
        RECT  6.835 30.255 7.0575 30.32 ;
        RECT  6.8025 30.2875 6.8675 30.4225 ;
        RECT  6.58 28.755 6.715 28.82 ;
        RECT  6.82 29.285 6.955 29.35 ;
        RECT  7.295 29.6225 7.855 29.6875 ;
        RECT  7.295 28.2775 7.855 28.3425 ;
        RECT  7.7225 28.3425 7.7875 28.5925 ;
        RECT  7.7225 29.4875 7.7875 29.6225 ;
        RECT  7.3625 29.5525 7.4275 29.6225 ;
        RECT  7.3625 28.3425 7.4275 28.4575 ;
        RECT  7.5525 28.4575 7.6175 29.52 ;
        RECT  7.295 28.995 7.33 29.06 ;
        RECT  7.6175 28.995 7.855 29.06 ;
        RECT  7.3625 29.3525 7.4275 29.4875 ;
        RECT  7.5525 29.3525 7.6175 29.4875 ;
        RECT  7.3625 28.7475 7.4275 28.8825 ;
        RECT  7.5525 28.7475 7.6175 28.8825 ;
        RECT  7.7225 28.5925 7.7875 28.7275 ;
        RECT  7.7225 29.5525 7.7875 29.6875 ;
        RECT  7.33 29.07 7.465 29.135 ;
        RECT  6.545 28.6775 6.68 28.7425 ;
        RECT  5.5325 28.61 5.5975 28.745 ;
        RECT  5.46 30.9675 5.595 31.0325 ;
        RECT  5.915 30.9675 6.05 31.0325 ;
        RECT  5.985 29.6225 6.545 29.6875 ;
        RECT  5.985 30.9675 6.545 31.0325 ;
        RECT  6.4125 30.7175 6.4775 30.9675 ;
        RECT  6.4125 29.6875 6.4775 29.8225 ;
        RECT  6.0525 29.6875 6.1175 29.7575 ;
        RECT  6.0525 30.8525 6.1175 30.9675 ;
        RECT  6.2425 29.79 6.3075 30.8525 ;
        RECT  5.985 30.25 6.02 30.315 ;
        RECT  6.3075 30.25 6.545 30.315 ;
        RECT  6.0525 29.8925 6.1175 30.0275 ;
        RECT  6.2425 29.8925 6.3075 30.0275 ;
        RECT  6.0525 30.7175 6.1175 30.8525 ;
        RECT  6.2425 30.7175 6.3075 30.8525 ;
        RECT  6.4125 30.7175 6.4775 30.8525 ;
        RECT  6.4125 29.7575 6.4775 29.8925 ;
        RECT  6.02 30.25 6.155 30.315 ;
        RECT  6.545 29.6225 7.295 29.6875 ;
        RECT  6.545 30.9675 7.295 31.0325 ;
        RECT  7.1625 30.7175 7.2275 31.0 ;
        RECT  7.1625 29.655 7.2275 29.835 ;
        RECT  6.6125 30.7175 6.6775 31.0 ;
        RECT  6.9925 30.7175 7.0575 31.0 ;
        RECT  6.6125 29.655 6.6775 29.9375 ;
        RECT  6.545 30.565 6.58 30.63 ;
        RECT  6.545 30.035 6.82 30.1 ;
        RECT  7.0575 30.2525 7.295 30.3175 ;
        RECT  6.6125 29.9375 6.6775 30.0725 ;
        RECT  6.8025 29.9375 6.8675 30.0725 ;
        RECT  6.8025 29.9375 6.8675 30.0725 ;
        RECT  6.9925 29.9375 7.0575 30.0725 ;
        RECT  6.6125 30.7175 6.6775 30.8525 ;
        RECT  6.8025 30.7175 6.8675 30.8525 ;
        RECT  6.8025 30.7175 6.8675 30.8525 ;
        RECT  6.9925 30.7175 7.0575 30.8525 ;
        RECT  7.1625 30.7175 7.2275 30.8525 ;
        RECT  7.1625 29.8025 7.2275 29.9375 ;
        RECT  7.025 30.55 7.09 30.615 ;
        RECT  6.8025 30.55 6.8675 30.615 ;
        RECT  7.025 29.8025 7.09 30.5825 ;
        RECT  6.835 30.55 7.0575 30.615 ;
        RECT  6.8025 30.5825 6.8675 30.7175 ;
        RECT  6.58 30.565 6.715 30.63 ;
        RECT  6.82 30.035 6.955 30.1 ;
        RECT  7.295 29.6225 7.855 29.6875 ;
        RECT  7.295 30.9675 7.855 31.0325 ;
        RECT  7.7225 30.7175 7.7875 30.9675 ;
        RECT  7.7225 29.6875 7.7875 29.8225 ;
        RECT  7.3625 29.6875 7.4275 29.7575 ;
        RECT  7.3625 30.8525 7.4275 30.9675 ;
        RECT  7.5525 29.79 7.6175 30.8525 ;
        RECT  7.295 30.25 7.33 30.315 ;
        RECT  7.6175 30.25 7.855 30.315 ;
        RECT  7.3625 29.8925 7.4275 30.0275 ;
        RECT  7.5525 29.8925 7.6175 30.0275 ;
        RECT  7.3625 30.7175 7.4275 30.8525 ;
        RECT  7.5525 30.7175 7.6175 30.8525 ;
        RECT  7.7225 30.7175 7.7875 30.8525 ;
        RECT  7.7225 29.7575 7.7875 29.8925 ;
        RECT  7.33 30.25 7.465 30.315 ;
        RECT  6.545 30.5675 6.68 30.6325 ;
        RECT  5.5325 30.565 5.5975 30.7 ;
        RECT  5.46 32.3125 5.595 32.3775 ;
        RECT  5.915 32.3125 6.05 32.3775 ;
        RECT  5.985 32.3125 6.545 32.3775 ;
        RECT  5.985 30.9675 6.545 31.0325 ;
        RECT  6.4125 31.0325 6.4775 31.2825 ;
        RECT  6.4125 32.1775 6.4775 32.3125 ;
        RECT  6.0525 32.2425 6.1175 32.3125 ;
        RECT  6.0525 31.0325 6.1175 31.1475 ;
        RECT  6.2425 31.1475 6.3075 32.21 ;
        RECT  5.985 31.685 6.02 31.75 ;
        RECT  6.3075 31.685 6.545 31.75 ;
        RECT  6.0525 32.0425 6.1175 32.1775 ;
        RECT  6.2425 32.0425 6.3075 32.1775 ;
        RECT  6.0525 31.4375 6.1175 31.5725 ;
        RECT  6.2425 31.4375 6.3075 31.5725 ;
        RECT  6.4125 31.2825 6.4775 31.4175 ;
        RECT  6.4125 32.2425 6.4775 32.3775 ;
        RECT  6.02 31.76 6.155 31.825 ;
        RECT  6.545 32.3125 7.295 32.3775 ;
        RECT  6.545 30.9675 7.295 31.0325 ;
        RECT  7.1625 31.0 7.2275 31.2825 ;
        RECT  7.1625 32.165 7.2275 32.345 ;
        RECT  6.6125 31.0 6.6775 31.2825 ;
        RECT  6.9925 31.0 7.0575 31.2825 ;
        RECT  6.6125 32.0625 6.6775 32.345 ;
        RECT  6.545 31.37 6.58 31.435 ;
        RECT  6.545 31.9 6.82 31.965 ;
        RECT  7.0575 31.6825 7.295 31.7475 ;
        RECT  6.6125 31.9075 6.6775 32.0425 ;
        RECT  6.8025 31.9075 6.8675 32.0425 ;
        RECT  6.8025 31.9075 6.8675 32.0425 ;
        RECT  6.9925 31.9075 7.0575 32.0425 ;
        RECT  6.6125 31.4375 6.6775 31.5725 ;
        RECT  6.8025 31.4375 6.8675 31.5725 ;
        RECT  6.8025 31.4375 6.8675 31.5725 ;
        RECT  6.9925 31.4375 7.0575 31.5725 ;
        RECT  7.1625 31.2825 7.2275 31.4175 ;
        RECT  7.1625 32.1975 7.2275 32.3325 ;
        RECT  7.025 32.945 7.09 33.01 ;
        RECT  6.8025 32.945 6.8675 33.01 ;
        RECT  7.025 32.1975 7.09 32.9775 ;
        RECT  6.835 32.945 7.0575 33.01 ;
        RECT  6.8025 32.9775 6.8675 33.1125 ;
        RECT  6.58 31.445 6.715 31.51 ;
        RECT  6.82 31.975 6.955 32.04 ;
        RECT  7.295 32.3125 7.855 32.3775 ;
        RECT  7.295 30.9675 7.855 31.0325 ;
        RECT  7.7225 31.0325 7.7875 31.2825 ;
        RECT  7.7225 32.1775 7.7875 32.3125 ;
        RECT  7.3625 32.2425 7.4275 32.3125 ;
        RECT  7.3625 31.0325 7.4275 31.1475 ;
        RECT  7.5525 31.1475 7.6175 32.21 ;
        RECT  7.295 31.685 7.33 31.75 ;
        RECT  7.6175 31.685 7.855 31.75 ;
        RECT  7.3625 32.0425 7.4275 32.1775 ;
        RECT  7.5525 32.0425 7.6175 32.1775 ;
        RECT  7.3625 31.4375 7.4275 31.5725 ;
        RECT  7.5525 31.4375 7.6175 31.5725 ;
        RECT  7.7225 31.2825 7.7875 31.4175 ;
        RECT  7.7225 32.2425 7.7875 32.3775 ;
        RECT  7.33 31.76 7.465 31.825 ;
        RECT  6.545 31.3675 6.68 31.4325 ;
        RECT  5.5325 31.3 5.5975 31.435 ;
        RECT  5.46 33.6575 5.595 33.7225 ;
        RECT  5.915 33.6575 6.05 33.7225 ;
        RECT  5.985 32.3125 6.545 32.3775 ;
        RECT  5.985 33.6575 6.545 33.7225 ;
        RECT  6.4125 33.4075 6.4775 33.6575 ;
        RECT  6.4125 32.3775 6.4775 32.5125 ;
        RECT  6.0525 32.3775 6.1175 32.4475 ;
        RECT  6.0525 33.5425 6.1175 33.6575 ;
        RECT  6.2425 32.48 6.3075 33.5425 ;
        RECT  5.985 32.94 6.02 33.005 ;
        RECT  6.3075 32.94 6.545 33.005 ;
        RECT  6.0525 32.5825 6.1175 32.7175 ;
        RECT  6.2425 32.5825 6.3075 32.7175 ;
        RECT  6.0525 33.4075 6.1175 33.5425 ;
        RECT  6.2425 33.4075 6.3075 33.5425 ;
        RECT  6.4125 33.4075 6.4775 33.5425 ;
        RECT  6.4125 32.4475 6.4775 32.5825 ;
        RECT  6.02 32.94 6.155 33.005 ;
        RECT  6.545 32.3125 7.295 32.3775 ;
        RECT  6.545 33.6575 7.295 33.7225 ;
        RECT  7.1625 33.4075 7.2275 33.69 ;
        RECT  7.1625 32.345 7.2275 32.525 ;
        RECT  6.6125 33.4075 6.6775 33.69 ;
        RECT  6.9925 33.4075 7.0575 33.69 ;
        RECT  6.6125 32.345 6.6775 32.6275 ;
        RECT  6.545 33.255 6.58 33.32 ;
        RECT  6.545 32.725 6.82 32.79 ;
        RECT  7.0575 32.9425 7.295 33.0075 ;
        RECT  6.6125 32.6275 6.6775 32.7625 ;
        RECT  6.8025 32.6275 6.8675 32.7625 ;
        RECT  6.8025 32.6275 6.8675 32.7625 ;
        RECT  6.9925 32.6275 7.0575 32.7625 ;
        RECT  6.6125 33.4075 6.6775 33.5425 ;
        RECT  6.8025 33.4075 6.8675 33.5425 ;
        RECT  6.8025 33.4075 6.8675 33.5425 ;
        RECT  6.9925 33.4075 7.0575 33.5425 ;
        RECT  7.1625 33.4075 7.2275 33.5425 ;
        RECT  7.1625 32.4925 7.2275 32.6275 ;
        RECT  7.025 33.24 7.09 33.305 ;
        RECT  6.8025 33.24 6.8675 33.305 ;
        RECT  7.025 32.4925 7.09 33.2725 ;
        RECT  6.835 33.24 7.0575 33.305 ;
        RECT  6.8025 33.2725 6.8675 33.4075 ;
        RECT  6.58 33.255 6.715 33.32 ;
        RECT  6.82 32.725 6.955 32.79 ;
        RECT  7.295 32.3125 7.855 32.3775 ;
        RECT  7.295 33.6575 7.855 33.7225 ;
        RECT  7.7225 33.4075 7.7875 33.6575 ;
        RECT  7.7225 32.3775 7.7875 32.5125 ;
        RECT  7.3625 32.3775 7.4275 32.4475 ;
        RECT  7.3625 33.5425 7.4275 33.6575 ;
        RECT  7.5525 32.48 7.6175 33.5425 ;
        RECT  7.295 32.94 7.33 33.005 ;
        RECT  7.6175 32.94 7.855 33.005 ;
        RECT  7.3625 32.5825 7.4275 32.7175 ;
        RECT  7.5525 32.5825 7.6175 32.7175 ;
        RECT  7.3625 33.4075 7.4275 33.5425 ;
        RECT  7.5525 33.4075 7.6175 33.5425 ;
        RECT  7.7225 33.4075 7.7875 33.5425 ;
        RECT  7.7225 32.4475 7.7875 32.5825 ;
        RECT  7.33 32.94 7.465 33.005 ;
        RECT  6.545 33.2575 6.68 33.3225 ;
        RECT  5.5325 33.255 5.5975 33.39 ;
        RECT  5.46 35.0025 5.595 35.0675 ;
        RECT  5.915 35.0025 6.05 35.0675 ;
        RECT  5.985 35.0025 6.545 35.0675 ;
        RECT  5.985 33.6575 6.545 33.7225 ;
        RECT  6.4125 33.7225 6.4775 33.9725 ;
        RECT  6.4125 34.8675 6.4775 35.0025 ;
        RECT  6.0525 34.9325 6.1175 35.0025 ;
        RECT  6.0525 33.7225 6.1175 33.8375 ;
        RECT  6.2425 33.8375 6.3075 34.9 ;
        RECT  5.985 34.375 6.02 34.44 ;
        RECT  6.3075 34.375 6.545 34.44 ;
        RECT  6.0525 34.7325 6.1175 34.8675 ;
        RECT  6.2425 34.7325 6.3075 34.8675 ;
        RECT  6.0525 34.1275 6.1175 34.2625 ;
        RECT  6.2425 34.1275 6.3075 34.2625 ;
        RECT  6.4125 33.9725 6.4775 34.1075 ;
        RECT  6.4125 34.9325 6.4775 35.0675 ;
        RECT  6.02 34.45 6.155 34.515 ;
        RECT  6.545 35.0025 7.295 35.0675 ;
        RECT  6.545 33.6575 7.295 33.7225 ;
        RECT  7.1625 33.69 7.2275 33.9725 ;
        RECT  7.1625 34.855 7.2275 35.035 ;
        RECT  6.6125 33.69 6.6775 33.9725 ;
        RECT  6.9925 33.69 7.0575 33.9725 ;
        RECT  6.6125 34.7525 6.6775 35.035 ;
        RECT  6.545 34.06 6.58 34.125 ;
        RECT  6.545 34.59 6.82 34.655 ;
        RECT  7.0575 34.3725 7.295 34.4375 ;
        RECT  6.6125 34.5975 6.6775 34.7325 ;
        RECT  6.8025 34.5975 6.8675 34.7325 ;
        RECT  6.8025 34.5975 6.8675 34.7325 ;
        RECT  6.9925 34.5975 7.0575 34.7325 ;
        RECT  6.6125 34.1275 6.6775 34.2625 ;
        RECT  6.8025 34.1275 6.8675 34.2625 ;
        RECT  6.8025 34.1275 6.8675 34.2625 ;
        RECT  6.9925 34.1275 7.0575 34.2625 ;
        RECT  7.1625 33.9725 7.2275 34.1075 ;
        RECT  7.1625 34.8875 7.2275 35.0225 ;
        RECT  7.025 35.635 7.09 35.7 ;
        RECT  6.8025 35.635 6.8675 35.7 ;
        RECT  7.025 34.8875 7.09 35.6675 ;
        RECT  6.835 35.635 7.0575 35.7 ;
        RECT  6.8025 35.6675 6.8675 35.8025 ;
        RECT  6.58 34.135 6.715 34.2 ;
        RECT  6.82 34.665 6.955 34.73 ;
        RECT  7.295 35.0025 7.855 35.0675 ;
        RECT  7.295 33.6575 7.855 33.7225 ;
        RECT  7.7225 33.7225 7.7875 33.9725 ;
        RECT  7.7225 34.8675 7.7875 35.0025 ;
        RECT  7.3625 34.9325 7.4275 35.0025 ;
        RECT  7.3625 33.7225 7.4275 33.8375 ;
        RECT  7.5525 33.8375 7.6175 34.9 ;
        RECT  7.295 34.375 7.33 34.44 ;
        RECT  7.6175 34.375 7.855 34.44 ;
        RECT  7.3625 34.7325 7.4275 34.8675 ;
        RECT  7.5525 34.7325 7.6175 34.8675 ;
        RECT  7.3625 34.1275 7.4275 34.2625 ;
        RECT  7.5525 34.1275 7.6175 34.2625 ;
        RECT  7.7225 33.9725 7.7875 34.1075 ;
        RECT  7.7225 34.9325 7.7875 35.0675 ;
        RECT  7.33 34.45 7.465 34.515 ;
        RECT  6.545 34.0575 6.68 34.1225 ;
        RECT  5.5325 33.99 5.5975 34.125 ;
        RECT  5.46 36.3475 5.595 36.4125 ;
        RECT  5.915 36.3475 6.05 36.4125 ;
        RECT  5.985 35.0025 6.545 35.0675 ;
        RECT  5.985 36.3475 6.545 36.4125 ;
        RECT  6.4125 36.0975 6.4775 36.3475 ;
        RECT  6.4125 35.0675 6.4775 35.2025 ;
        RECT  6.0525 35.0675 6.1175 35.1375 ;
        RECT  6.0525 36.2325 6.1175 36.3475 ;
        RECT  6.2425 35.17 6.3075 36.2325 ;
        RECT  5.985 35.63 6.02 35.695 ;
        RECT  6.3075 35.63 6.545 35.695 ;
        RECT  6.0525 35.2725 6.1175 35.4075 ;
        RECT  6.2425 35.2725 6.3075 35.4075 ;
        RECT  6.0525 36.0975 6.1175 36.2325 ;
        RECT  6.2425 36.0975 6.3075 36.2325 ;
        RECT  6.4125 36.0975 6.4775 36.2325 ;
        RECT  6.4125 35.1375 6.4775 35.2725 ;
        RECT  6.02 35.63 6.155 35.695 ;
        RECT  6.545 35.0025 7.295 35.0675 ;
        RECT  6.545 36.3475 7.295 36.4125 ;
        RECT  7.1625 36.0975 7.2275 36.38 ;
        RECT  7.1625 35.035 7.2275 35.215 ;
        RECT  6.6125 36.0975 6.6775 36.38 ;
        RECT  6.9925 36.0975 7.0575 36.38 ;
        RECT  6.6125 35.035 6.6775 35.3175 ;
        RECT  6.545 35.945 6.58 36.01 ;
        RECT  6.545 35.415 6.82 35.48 ;
        RECT  7.0575 35.6325 7.295 35.6975 ;
        RECT  6.6125 35.3175 6.6775 35.4525 ;
        RECT  6.8025 35.3175 6.8675 35.4525 ;
        RECT  6.8025 35.3175 6.8675 35.4525 ;
        RECT  6.9925 35.3175 7.0575 35.4525 ;
        RECT  6.6125 36.0975 6.6775 36.2325 ;
        RECT  6.8025 36.0975 6.8675 36.2325 ;
        RECT  6.8025 36.0975 6.8675 36.2325 ;
        RECT  6.9925 36.0975 7.0575 36.2325 ;
        RECT  7.1625 36.0975 7.2275 36.2325 ;
        RECT  7.1625 35.1825 7.2275 35.3175 ;
        RECT  7.025 35.93 7.09 35.995 ;
        RECT  6.8025 35.93 6.8675 35.995 ;
        RECT  7.025 35.1825 7.09 35.9625 ;
        RECT  6.835 35.93 7.0575 35.995 ;
        RECT  6.8025 35.9625 6.8675 36.0975 ;
        RECT  6.58 35.945 6.715 36.01 ;
        RECT  6.82 35.415 6.955 35.48 ;
        RECT  7.295 35.0025 7.855 35.0675 ;
        RECT  7.295 36.3475 7.855 36.4125 ;
        RECT  7.7225 36.0975 7.7875 36.3475 ;
        RECT  7.7225 35.0675 7.7875 35.2025 ;
        RECT  7.3625 35.0675 7.4275 35.1375 ;
        RECT  7.3625 36.2325 7.4275 36.3475 ;
        RECT  7.5525 35.17 7.6175 36.2325 ;
        RECT  7.295 35.63 7.33 35.695 ;
        RECT  7.6175 35.63 7.855 35.695 ;
        RECT  7.3625 35.2725 7.4275 35.4075 ;
        RECT  7.5525 35.2725 7.6175 35.4075 ;
        RECT  7.3625 36.0975 7.4275 36.2325 ;
        RECT  7.5525 36.0975 7.6175 36.2325 ;
        RECT  7.7225 36.0975 7.7875 36.2325 ;
        RECT  7.7225 35.1375 7.7875 35.2725 ;
        RECT  7.33 35.63 7.465 35.695 ;
        RECT  6.545 35.9475 6.68 36.0125 ;
        RECT  5.5325 35.945 5.5975 36.08 ;
        RECT  5.46 37.6925 5.595 37.7575 ;
        RECT  5.915 37.6925 6.05 37.7575 ;
        RECT  5.985 37.6925 6.545 37.7575 ;
        RECT  5.985 36.3475 6.545 36.4125 ;
        RECT  6.4125 36.4125 6.4775 36.6625 ;
        RECT  6.4125 37.5575 6.4775 37.6925 ;
        RECT  6.0525 37.6225 6.1175 37.6925 ;
        RECT  6.0525 36.4125 6.1175 36.5275 ;
        RECT  6.2425 36.5275 6.3075 37.59 ;
        RECT  5.985 37.065 6.02 37.13 ;
        RECT  6.3075 37.065 6.545 37.13 ;
        RECT  6.0525 37.4225 6.1175 37.5575 ;
        RECT  6.2425 37.4225 6.3075 37.5575 ;
        RECT  6.0525 36.8175 6.1175 36.9525 ;
        RECT  6.2425 36.8175 6.3075 36.9525 ;
        RECT  6.4125 36.6625 6.4775 36.7975 ;
        RECT  6.4125 37.6225 6.4775 37.7575 ;
        RECT  6.02 37.14 6.155 37.205 ;
        RECT  6.545 37.6925 7.295 37.7575 ;
        RECT  6.545 36.3475 7.295 36.4125 ;
        RECT  7.1625 36.38 7.2275 36.6625 ;
        RECT  7.1625 37.545 7.2275 37.725 ;
        RECT  6.6125 36.38 6.6775 36.6625 ;
        RECT  6.9925 36.38 7.0575 36.6625 ;
        RECT  6.6125 37.4425 6.6775 37.725 ;
        RECT  6.545 36.75 6.58 36.815 ;
        RECT  6.545 37.28 6.82 37.345 ;
        RECT  7.0575 37.0625 7.295 37.1275 ;
        RECT  6.6125 37.2875 6.6775 37.4225 ;
        RECT  6.8025 37.2875 6.8675 37.4225 ;
        RECT  6.8025 37.2875 6.8675 37.4225 ;
        RECT  6.9925 37.2875 7.0575 37.4225 ;
        RECT  6.6125 36.8175 6.6775 36.9525 ;
        RECT  6.8025 36.8175 6.8675 36.9525 ;
        RECT  6.8025 36.8175 6.8675 36.9525 ;
        RECT  6.9925 36.8175 7.0575 36.9525 ;
        RECT  7.1625 36.6625 7.2275 36.7975 ;
        RECT  7.1625 37.5775 7.2275 37.7125 ;
        RECT  7.025 38.325 7.09 38.39 ;
        RECT  6.8025 38.325 6.8675 38.39 ;
        RECT  7.025 37.5775 7.09 38.3575 ;
        RECT  6.835 38.325 7.0575 38.39 ;
        RECT  6.8025 38.3575 6.8675 38.4925 ;
        RECT  6.58 36.825 6.715 36.89 ;
        RECT  6.82 37.355 6.955 37.42 ;
        RECT  7.295 37.6925 7.855 37.7575 ;
        RECT  7.295 36.3475 7.855 36.4125 ;
        RECT  7.7225 36.4125 7.7875 36.6625 ;
        RECT  7.7225 37.5575 7.7875 37.6925 ;
        RECT  7.3625 37.6225 7.4275 37.6925 ;
        RECT  7.3625 36.4125 7.4275 36.5275 ;
        RECT  7.5525 36.5275 7.6175 37.59 ;
        RECT  7.295 37.065 7.33 37.13 ;
        RECT  7.6175 37.065 7.855 37.13 ;
        RECT  7.3625 37.4225 7.4275 37.5575 ;
        RECT  7.5525 37.4225 7.6175 37.5575 ;
        RECT  7.3625 36.8175 7.4275 36.9525 ;
        RECT  7.5525 36.8175 7.6175 36.9525 ;
        RECT  7.7225 36.6625 7.7875 36.7975 ;
        RECT  7.7225 37.6225 7.7875 37.7575 ;
        RECT  7.33 37.14 7.465 37.205 ;
        RECT  6.545 36.7475 6.68 36.8125 ;
        RECT  5.5325 36.68 5.5975 36.815 ;
        RECT  5.46 39.0375 5.595 39.1025 ;
        RECT  5.915 39.0375 6.05 39.1025 ;
        RECT  5.985 37.6925 6.545 37.7575 ;
        RECT  5.985 39.0375 6.545 39.1025 ;
        RECT  6.4125 38.7875 6.4775 39.0375 ;
        RECT  6.4125 37.7575 6.4775 37.8925 ;
        RECT  6.0525 37.7575 6.1175 37.8275 ;
        RECT  6.0525 38.9225 6.1175 39.0375 ;
        RECT  6.2425 37.86 6.3075 38.9225 ;
        RECT  5.985 38.32 6.02 38.385 ;
        RECT  6.3075 38.32 6.545 38.385 ;
        RECT  6.0525 37.9625 6.1175 38.0975 ;
        RECT  6.2425 37.9625 6.3075 38.0975 ;
        RECT  6.0525 38.7875 6.1175 38.9225 ;
        RECT  6.2425 38.7875 6.3075 38.9225 ;
        RECT  6.4125 38.7875 6.4775 38.9225 ;
        RECT  6.4125 37.8275 6.4775 37.9625 ;
        RECT  6.02 38.32 6.155 38.385 ;
        RECT  6.545 37.6925 7.295 37.7575 ;
        RECT  6.545 39.0375 7.295 39.1025 ;
        RECT  7.1625 38.7875 7.2275 39.07 ;
        RECT  7.1625 37.725 7.2275 37.905 ;
        RECT  6.6125 38.7875 6.6775 39.07 ;
        RECT  6.9925 38.7875 7.0575 39.07 ;
        RECT  6.6125 37.725 6.6775 38.0075 ;
        RECT  6.545 38.635 6.58 38.7 ;
        RECT  6.545 38.105 6.82 38.17 ;
        RECT  7.0575 38.3225 7.295 38.3875 ;
        RECT  6.6125 38.0075 6.6775 38.1425 ;
        RECT  6.8025 38.0075 6.8675 38.1425 ;
        RECT  6.8025 38.0075 6.8675 38.1425 ;
        RECT  6.9925 38.0075 7.0575 38.1425 ;
        RECT  6.6125 38.7875 6.6775 38.9225 ;
        RECT  6.8025 38.7875 6.8675 38.9225 ;
        RECT  6.8025 38.7875 6.8675 38.9225 ;
        RECT  6.9925 38.7875 7.0575 38.9225 ;
        RECT  7.1625 38.7875 7.2275 38.9225 ;
        RECT  7.1625 37.8725 7.2275 38.0075 ;
        RECT  7.025 38.62 7.09 38.685 ;
        RECT  6.8025 38.62 6.8675 38.685 ;
        RECT  7.025 37.8725 7.09 38.6525 ;
        RECT  6.835 38.62 7.0575 38.685 ;
        RECT  6.8025 38.6525 6.8675 38.7875 ;
        RECT  6.58 38.635 6.715 38.7 ;
        RECT  6.82 38.105 6.955 38.17 ;
        RECT  7.295 37.6925 7.855 37.7575 ;
        RECT  7.295 39.0375 7.855 39.1025 ;
        RECT  7.7225 38.7875 7.7875 39.0375 ;
        RECT  7.7225 37.7575 7.7875 37.8925 ;
        RECT  7.3625 37.7575 7.4275 37.8275 ;
        RECT  7.3625 38.9225 7.4275 39.0375 ;
        RECT  7.5525 37.86 7.6175 38.9225 ;
        RECT  7.295 38.32 7.33 38.385 ;
        RECT  7.6175 38.32 7.855 38.385 ;
        RECT  7.3625 37.9625 7.4275 38.0975 ;
        RECT  7.5525 37.9625 7.6175 38.0975 ;
        RECT  7.3625 38.7875 7.4275 38.9225 ;
        RECT  7.5525 38.7875 7.6175 38.9225 ;
        RECT  7.7225 38.7875 7.7875 38.9225 ;
        RECT  7.7225 37.8275 7.7875 37.9625 ;
        RECT  7.33 38.32 7.465 38.385 ;
        RECT  6.545 38.6375 6.68 38.7025 ;
        RECT  5.5325 38.635 5.5975 38.77 ;
        RECT  5.46 40.3825 5.595 40.4475 ;
        RECT  5.915 40.3825 6.05 40.4475 ;
        RECT  5.985 40.3825 6.545 40.4475 ;
        RECT  5.985 39.0375 6.545 39.1025 ;
        RECT  6.4125 39.1025 6.4775 39.3525 ;
        RECT  6.4125 40.2475 6.4775 40.3825 ;
        RECT  6.0525 40.3125 6.1175 40.3825 ;
        RECT  6.0525 39.1025 6.1175 39.2175 ;
        RECT  6.2425 39.2175 6.3075 40.28 ;
        RECT  5.985 39.755 6.02 39.82 ;
        RECT  6.3075 39.755 6.545 39.82 ;
        RECT  6.0525 40.1125 6.1175 40.2475 ;
        RECT  6.2425 40.1125 6.3075 40.2475 ;
        RECT  6.0525 39.5075 6.1175 39.6425 ;
        RECT  6.2425 39.5075 6.3075 39.6425 ;
        RECT  6.4125 39.3525 6.4775 39.4875 ;
        RECT  6.4125 40.3125 6.4775 40.4475 ;
        RECT  6.02 39.83 6.155 39.895 ;
        RECT  6.545 40.3825 7.295 40.4475 ;
        RECT  6.545 39.0375 7.295 39.1025 ;
        RECT  7.1625 39.07 7.2275 39.3525 ;
        RECT  7.1625 40.235 7.2275 40.415 ;
        RECT  6.6125 39.07 6.6775 39.3525 ;
        RECT  6.9925 39.07 7.0575 39.3525 ;
        RECT  6.6125 40.1325 6.6775 40.415 ;
        RECT  6.545 39.44 6.58 39.505 ;
        RECT  6.545 39.97 6.82 40.035 ;
        RECT  7.0575 39.7525 7.295 39.8175 ;
        RECT  6.6125 39.9775 6.6775 40.1125 ;
        RECT  6.8025 39.9775 6.8675 40.1125 ;
        RECT  6.8025 39.9775 6.8675 40.1125 ;
        RECT  6.9925 39.9775 7.0575 40.1125 ;
        RECT  6.6125 39.5075 6.6775 39.6425 ;
        RECT  6.8025 39.5075 6.8675 39.6425 ;
        RECT  6.8025 39.5075 6.8675 39.6425 ;
        RECT  6.9925 39.5075 7.0575 39.6425 ;
        RECT  7.1625 39.3525 7.2275 39.4875 ;
        RECT  7.1625 40.2675 7.2275 40.4025 ;
        RECT  7.025 41.015 7.09 41.08 ;
        RECT  6.8025 41.015 6.8675 41.08 ;
        RECT  7.025 40.2675 7.09 41.0475 ;
        RECT  6.835 41.015 7.0575 41.08 ;
        RECT  6.8025 41.0475 6.8675 41.1825 ;
        RECT  6.58 39.515 6.715 39.58 ;
        RECT  6.82 40.045 6.955 40.11 ;
        RECT  7.295 40.3825 7.855 40.4475 ;
        RECT  7.295 39.0375 7.855 39.1025 ;
        RECT  7.7225 39.1025 7.7875 39.3525 ;
        RECT  7.7225 40.2475 7.7875 40.3825 ;
        RECT  7.3625 40.3125 7.4275 40.3825 ;
        RECT  7.3625 39.1025 7.4275 39.2175 ;
        RECT  7.5525 39.2175 7.6175 40.28 ;
        RECT  7.295 39.755 7.33 39.82 ;
        RECT  7.6175 39.755 7.855 39.82 ;
        RECT  7.3625 40.1125 7.4275 40.2475 ;
        RECT  7.5525 40.1125 7.6175 40.2475 ;
        RECT  7.3625 39.5075 7.4275 39.6425 ;
        RECT  7.5525 39.5075 7.6175 39.6425 ;
        RECT  7.7225 39.3525 7.7875 39.4875 ;
        RECT  7.7225 40.3125 7.7875 40.4475 ;
        RECT  7.33 39.83 7.465 39.895 ;
        RECT  6.545 39.4375 6.68 39.5025 ;
        RECT  5.5325 39.37 5.5975 39.505 ;
        RECT  1.0825 5.02 1.1475 7.84 ;
        RECT  7.08 5.02 7.145 7.84 ;
        RECT  3.6 7.235 3.735 7.3 ;
        RECT  3.6 7.42 3.735 7.485 ;
        RECT  2.365 7.235 2.5 7.3 ;
        RECT  2.365 7.42 2.5 7.485 ;
        RECT  3.6 7.425 3.735 7.49 ;
        RECT  3.6 7.61 3.735 7.675 ;
        RECT  6.56 7.425 6.695 7.49 ;
        RECT  6.56 7.61 6.695 7.675 ;
        RECT  2.365 7.425 2.5 7.49 ;
        RECT  2.365 7.61 2.5 7.675 ;
        RECT  6.56 7.235 6.695 7.3 ;
        RECT  6.56 7.42 6.695 7.485 ;
        RECT  1.83 7.425 1.965 7.49 ;
        RECT  1.83 7.61 1.965 7.675 ;
        RECT  4.79 7.285 4.925 7.35 ;
        RECT  4.79 7.47 4.925 7.535 ;
        RECT  5.325 7.235 5.46 7.3 ;
        RECT  5.325 7.42 5.46 7.485 ;
        RECT  5.325 7.425 5.46 7.49 ;
        RECT  5.325 7.61 5.46 7.675 ;
        RECT  5.75 7.235 5.885 7.3 ;
        RECT  5.75 7.42 5.885 7.485 ;
        RECT  2.79 7.235 2.925 7.3 ;
        RECT  2.79 7.42 2.925 7.485 ;
        RECT  6.135 7.235 6.27 7.3 ;
        RECT  6.135 7.42 6.27 7.485 ;
        RECT  6.135 7.425 6.27 7.49 ;
        RECT  6.135 7.61 6.27 7.675 ;
        RECT  2.79 7.425 2.925 7.49 ;
        RECT  2.79 7.61 2.925 7.675 ;
        RECT  5.75 7.425 5.885 7.49 ;
        RECT  5.75 7.61 5.885 7.675 ;
        RECT  3.175 7.425 3.31 7.49 ;
        RECT  3.175 7.61 3.31 7.675 ;
        RECT  3.175 7.235 3.31 7.3 ;
        RECT  3.175 7.42 3.31 7.485 ;
        RECT  1.405 7.425 1.54 7.49 ;
        RECT  1.405 7.61 1.54 7.675 ;
        RECT  4.38 7.35 4.515 7.415 ;
        RECT  4.38 7.535 4.515 7.6 ;
        RECT  1.115 7.4775 1.18 7.6125 ;
        RECT  6.6125 7.61 6.7475 7.675 ;
        RECT  4.7975 7.72 4.9325 7.785 ;
        RECT  3.8975 7.61 4.0325 7.675 ;
        RECT  4.3725 7.1875 4.5075 7.2525 ;
        RECT  6.9775 7.61 7.1125 7.675 ;
        RECT  1.435 7.1025 1.57 7.1675 ;
        RECT  5.5175 7.245 5.6525 7.31 ;
        RECT  3.91 7.2425 4.045 7.3075 ;
        RECT  2.5125 7.2425 2.6475 7.3075 ;
        RECT  1.295 7.8075 1.43 7.8725 ;
        RECT  1.4125 7.2325 1.5475 7.2975 ;
        RECT  3.0225 7.1625 3.0875 7.2975 ;
        RECT  1.9375 7.1925 2.0725 7.2575 ;
        RECT  5.9825 7.1625 6.0475 7.2975 ;
        RECT  6.87 7.285 7.005 7.35 ;
        RECT  3.4 7.365 3.535 7.43 ;
        RECT  6.36 7.375 6.495 7.44 ;
        RECT  4.67 7.5375 4.735 7.6725 ;
        RECT  4.3725 7.1025 4.5075 7.1675 ;
        RECT  1.665 7.6475 1.73 7.7825 ;
        RECT  3.1775 7.6075 3.3125 7.6725 ;
        RECT  6.87 7.2425 7.005 7.3075 ;
        RECT  6.36 7.42 6.495 7.485 ;
        RECT  5.9475 7.1025 6.0825 7.1675 ;
        RECT  1.245 7.1025 1.38 7.1675 ;
        RECT  3.91 7.2425 4.045 7.3075 ;
        RECT  2.9875 7.1025 3.1225 7.1675 ;
        RECT  2.7875 7.6075 2.9225 7.6725 ;
        RECT  2.7875 7.42 2.9225 7.485 ;
        RECT  3.4 7.42 3.535 7.485 ;
        RECT  5.7475 7.61 5.8825 7.675 ;
        RECT  5.7475 7.42 5.8825 7.485 ;
        RECT  1.115 7.1 1.18 7.875 ;
        RECT  4.185 7.74 7.08 7.805 ;
        RECT  6.695 7.235 7.005 7.3 ;
        RECT  6.27 7.61 6.56 7.675 ;
        RECT  5.46 7.61 5.75 7.675 ;
        RECT  7.0825 7.4625 7.145 7.535 ;
        RECT  6.695 7.42 7.08 7.49 ;
        RECT  5.46 7.42 5.75 7.49 ;
        RECT  5.98 7.42 6.1375 7.49 ;
        RECT  6.27 7.235 6.56 7.3 ;
        RECT  5.46 7.235 5.75 7.3 ;
        RECT  5.98 7.105 6.05 7.49 ;
        RECT  7.08 7.1 7.145 7.875 ;
        RECT  5.09 7.1 5.155 7.875 ;
        RECT  2.195 7.74 4.12 7.805 ;
        RECT  3.735 7.235 4.045 7.3 ;
        RECT  3.31 7.61 3.6 7.675 ;
        RECT  4.475 7.535 4.925 7.6 ;
        RECT  3.735 7.42 4.12 7.49 ;
        RECT  3.02 7.42 3.1775 7.49 ;
        RECT  4.0325 7.61 4.12 7.675 ;
        RECT  3.31 7.235 3.6 7.3 ;
        RECT  4.25 7.17 4.315 7.415 ;
        RECT  4.25 7.17 4.3725 7.2525 ;
        RECT  4.3725 7.165 4.5075 7.2325 ;
        RECT  4.12 7.1 4.185 7.875 ;
        RECT  2.5 7.61 2.79 7.675 ;
        RECT  1.9625 7.425 2.13 7.49 ;
        RECT  1.47 7.1675 1.54 7.425 ;
        RECT  1.405 7.61 1.83 7.675 ;
        RECT  2.5 7.42 2.79 7.49 ;
        RECT  1.66 7.61 1.735 7.7825 ;
        RECT  2.5 7.235 2.79 7.3 ;
        RECT  1.34 7.2325 1.4125 7.2975 ;
        RECT  3.02 7.105 3.09 7.49 ;
        RECT  2.05 7.1925 2.165 7.2575 ;
        RECT  1.275 7.1 1.34 7.875 ;
        RECT  2.13 7.1 2.195 7.875 ;
        RECT  1.12 7.67 1.1775 7.735 ;
        RECT  1.36 7.1025 1.4825 7.1675 ;
        RECT  4.9225 7.285 5.09 7.35 ;
        RECT  4.315 7.3475 4.4175 7.415 ;
        RECT  3.6 6.97 3.735 7.035 ;
        RECT  3.6 6.785 3.735 6.85 ;
        RECT  2.365 6.97 2.5 7.035 ;
        RECT  2.365 6.785 2.5 6.85 ;
        RECT  3.6 6.78 3.735 6.845 ;
        RECT  3.6 6.595 3.735 6.66 ;
        RECT  6.56 6.78 6.695 6.845 ;
        RECT  6.56 6.595 6.695 6.66 ;
        RECT  2.365 6.78 2.5 6.845 ;
        RECT  2.365 6.595 2.5 6.66 ;
        RECT  6.56 6.97 6.695 7.035 ;
        RECT  6.56 6.785 6.695 6.85 ;
        RECT  1.83 6.78 1.965 6.845 ;
        RECT  1.83 6.595 1.965 6.66 ;
        RECT  4.79 6.92 4.925 6.985 ;
        RECT  4.79 6.735 4.925 6.8 ;
        RECT  5.325 6.97 5.46 7.035 ;
        RECT  5.325 6.785 5.46 6.85 ;
        RECT  5.325 6.78 5.46 6.845 ;
        RECT  5.325 6.595 5.46 6.66 ;
        RECT  5.75 6.97 5.885 7.035 ;
        RECT  5.75 6.785 5.885 6.85 ;
        RECT  2.79 6.97 2.925 7.035 ;
        RECT  2.79 6.785 2.925 6.85 ;
        RECT  6.135 6.97 6.27 7.035 ;
        RECT  6.135 6.785 6.27 6.85 ;
        RECT  6.135 6.78 6.27 6.845 ;
        RECT  6.135 6.595 6.27 6.66 ;
        RECT  2.79 6.78 2.925 6.845 ;
        RECT  2.79 6.595 2.925 6.66 ;
        RECT  5.75 6.78 5.885 6.845 ;
        RECT  5.75 6.595 5.885 6.66 ;
        RECT  3.175 6.78 3.31 6.845 ;
        RECT  3.175 6.595 3.31 6.66 ;
        RECT  3.175 6.97 3.31 7.035 ;
        RECT  3.175 6.785 3.31 6.85 ;
        RECT  1.405 6.78 1.54 6.845 ;
        RECT  1.405 6.595 1.54 6.66 ;
        RECT  4.38 6.855 4.515 6.92 ;
        RECT  4.38 6.67 4.515 6.735 ;
        RECT  1.115 6.6575 1.18 6.7925 ;
        RECT  6.6125 6.595 6.7475 6.66 ;
        RECT  4.7975 6.485 4.9325 6.55 ;
        RECT  3.8975 6.595 4.0325 6.66 ;
        RECT  4.3725 7.0175 4.5075 7.0825 ;
        RECT  6.9775 6.595 7.1125 6.66 ;
        RECT  1.435 7.1025 1.57 7.1675 ;
        RECT  5.5175 6.96 5.6525 7.025 ;
        RECT  3.91 6.9625 4.045 7.0275 ;
        RECT  2.5125 6.9625 2.6475 7.0275 ;
        RECT  1.295 6.3975 1.43 6.4625 ;
        RECT  1.4125 6.9725 1.5475 7.0375 ;
        RECT  3.0225 6.9725 3.0875 7.1075 ;
        RECT  1.9375 7.0125 2.0725 7.0775 ;
        RECT  5.9825 6.9725 6.0475 7.1075 ;
        RECT  6.87 6.92 7.005 6.985 ;
        RECT  3.4 6.84 3.535 6.905 ;
        RECT  6.36 6.83 6.495 6.895 ;
        RECT  4.67 6.5975 4.735 6.7325 ;
        RECT  4.3725 7.1025 4.5075 7.1675 ;
        RECT  1.665 6.4875 1.73 6.6225 ;
        RECT  3.1775 6.5975 3.3125 6.6625 ;
        RECT  6.87 6.9625 7.005 7.0275 ;
        RECT  6.36 6.785 6.495 6.85 ;
        RECT  5.9475 7.1025 6.0825 7.1675 ;
        RECT  1.245 7.1025 1.38 7.1675 ;
        RECT  3.91 6.9625 4.045 7.0275 ;
        RECT  2.9875 7.1025 3.1225 7.1675 ;
        RECT  2.7875 6.5975 2.9225 6.6625 ;
        RECT  2.7875 6.785 2.9225 6.85 ;
        RECT  3.4 6.785 3.535 6.85 ;
        RECT  5.7475 6.595 5.8825 6.66 ;
        RECT  5.7475 6.785 5.8825 6.85 ;
        RECT  1.115 6.395 1.18 7.17 ;
        RECT  4.185 6.465 7.08 6.53 ;
        RECT  6.695 6.97 7.005 7.035 ;
        RECT  6.27 6.595 6.56 6.66 ;
        RECT  5.46 6.595 5.75 6.66 ;
        RECT  7.0825 6.735 7.145 6.8075 ;
        RECT  6.695 6.78 7.08 6.85 ;
        RECT  5.46 6.78 5.75 6.85 ;
        RECT  5.98 6.78 6.1375 6.85 ;
        RECT  6.27 6.97 6.56 7.035 ;
        RECT  5.46 6.97 5.75 7.035 ;
        RECT  5.98 6.78 6.05 7.165 ;
        RECT  7.08 6.395 7.145 7.17 ;
        RECT  5.09 6.395 5.155 7.17 ;
        RECT  2.195 6.465 4.12 6.53 ;
        RECT  3.735 6.97 4.045 7.035 ;
        RECT  3.31 6.595 3.6 6.66 ;
        RECT  4.475 6.67 4.925 6.735 ;
        RECT  3.735 6.78 4.12 6.85 ;
        RECT  3.02 6.78 3.1775 6.85 ;
        RECT  4.0325 6.595 4.12 6.66 ;
        RECT  3.31 6.97 3.6 7.035 ;
        RECT  4.25 6.855 4.315 7.1 ;
        RECT  4.25 7.0175 4.3725 7.1 ;
        RECT  4.3725 7.0375 4.5075 7.105 ;
        RECT  4.12 6.395 4.185 7.17 ;
        RECT  2.5 6.595 2.79 6.66 ;
        RECT  1.9625 6.78 2.13 6.845 ;
        RECT  1.47 6.845 1.54 7.1025 ;
        RECT  1.405 6.595 1.83 6.66 ;
        RECT  2.5 6.78 2.79 6.85 ;
        RECT  1.66 6.4875 1.735 6.66 ;
        RECT  2.5 6.97 2.79 7.035 ;
        RECT  1.34 6.9725 1.4125 7.0375 ;
        RECT  3.02 6.78 3.09 7.165 ;
        RECT  2.05 7.0125 2.165 7.0775 ;
        RECT  1.275 6.395 1.34 7.17 ;
        RECT  2.13 6.395 2.195 7.17 ;
        RECT  1.12 6.535 1.1775 6.6 ;
        RECT  1.36 7.1025 1.4825 7.1675 ;
        RECT  4.9225 6.92 5.09 6.985 ;
        RECT  4.315 6.855 4.4175 6.9225 ;
        RECT  3.6 5.825 3.735 5.89 ;
        RECT  3.6 6.01 3.735 6.075 ;
        RECT  2.365 5.825 2.5 5.89 ;
        RECT  2.365 6.01 2.5 6.075 ;
        RECT  3.6 6.015 3.735 6.08 ;
        RECT  3.6 6.2 3.735 6.265 ;
        RECT  6.56 6.015 6.695 6.08 ;
        RECT  6.56 6.2 6.695 6.265 ;
        RECT  2.365 6.015 2.5 6.08 ;
        RECT  2.365 6.2 2.5 6.265 ;
        RECT  6.56 5.825 6.695 5.89 ;
        RECT  6.56 6.01 6.695 6.075 ;
        RECT  1.83 6.015 1.965 6.08 ;
        RECT  1.83 6.2 1.965 6.265 ;
        RECT  4.79 5.875 4.925 5.94 ;
        RECT  4.79 6.06 4.925 6.125 ;
        RECT  5.325 5.825 5.46 5.89 ;
        RECT  5.325 6.01 5.46 6.075 ;
        RECT  5.325 6.015 5.46 6.08 ;
        RECT  5.325 6.2 5.46 6.265 ;
        RECT  5.75 5.825 5.885 5.89 ;
        RECT  5.75 6.01 5.885 6.075 ;
        RECT  2.79 5.825 2.925 5.89 ;
        RECT  2.79 6.01 2.925 6.075 ;
        RECT  6.135 5.825 6.27 5.89 ;
        RECT  6.135 6.01 6.27 6.075 ;
        RECT  6.135 6.015 6.27 6.08 ;
        RECT  6.135 6.2 6.27 6.265 ;
        RECT  2.79 6.015 2.925 6.08 ;
        RECT  2.79 6.2 2.925 6.265 ;
        RECT  5.75 6.015 5.885 6.08 ;
        RECT  5.75 6.2 5.885 6.265 ;
        RECT  3.175 6.015 3.31 6.08 ;
        RECT  3.175 6.2 3.31 6.265 ;
        RECT  3.175 5.825 3.31 5.89 ;
        RECT  3.175 6.01 3.31 6.075 ;
        RECT  1.405 6.015 1.54 6.08 ;
        RECT  1.405 6.2 1.54 6.265 ;
        RECT  4.38 5.94 4.515 6.005 ;
        RECT  4.38 6.125 4.515 6.19 ;
        RECT  1.115 6.0675 1.18 6.2025 ;
        RECT  6.6125 6.2 6.7475 6.265 ;
        RECT  4.7975 6.31 4.9325 6.375 ;
        RECT  3.8975 6.2 4.0325 6.265 ;
        RECT  4.3725 5.7775 4.5075 5.8425 ;
        RECT  6.9775 6.2 7.1125 6.265 ;
        RECT  1.435 5.6925 1.57 5.7575 ;
        RECT  5.5175 5.835 5.6525 5.9 ;
        RECT  3.91 5.8325 4.045 5.8975 ;
        RECT  2.5125 5.8325 2.6475 5.8975 ;
        RECT  1.295 6.3975 1.43 6.4625 ;
        RECT  1.4125 5.8225 1.5475 5.8875 ;
        RECT  3.0225 5.7525 3.0875 5.8875 ;
        RECT  1.9375 5.7825 2.0725 5.8475 ;
        RECT  5.9825 5.7525 6.0475 5.8875 ;
        RECT  6.87 5.875 7.005 5.94 ;
        RECT  3.4 5.955 3.535 6.02 ;
        RECT  6.36 5.965 6.495 6.03 ;
        RECT  4.67 6.1275 4.735 6.2625 ;
        RECT  4.3725 5.6925 4.5075 5.7575 ;
        RECT  1.665 6.2375 1.73 6.3725 ;
        RECT  3.1775 6.1975 3.3125 6.2625 ;
        RECT  6.87 5.8325 7.005 5.8975 ;
        RECT  6.36 6.01 6.495 6.075 ;
        RECT  5.9475 5.6925 6.0825 5.7575 ;
        RECT  1.245 5.6925 1.38 5.7575 ;
        RECT  3.91 5.8325 4.045 5.8975 ;
        RECT  2.9875 5.6925 3.1225 5.7575 ;
        RECT  2.7875 6.1975 2.9225 6.2625 ;
        RECT  2.7875 6.01 2.9225 6.075 ;
        RECT  3.4 6.01 3.535 6.075 ;
        RECT  5.7475 6.2 5.8825 6.265 ;
        RECT  5.7475 6.01 5.8825 6.075 ;
        RECT  1.115 5.69 1.18 6.465 ;
        RECT  4.185 6.33 7.08 6.395 ;
        RECT  6.695 5.825 7.005 5.89 ;
        RECT  6.27 6.2 6.56 6.265 ;
        RECT  5.46 6.2 5.75 6.265 ;
        RECT  7.0825 6.0525 7.145 6.125 ;
        RECT  6.695 6.01 7.08 6.08 ;
        RECT  5.46 6.01 5.75 6.08 ;
        RECT  5.98 6.01 6.1375 6.08 ;
        RECT  6.27 5.825 6.56 5.89 ;
        RECT  5.46 5.825 5.75 5.89 ;
        RECT  5.98 5.695 6.05 6.08 ;
        RECT  7.08 5.69 7.145 6.465 ;
        RECT  5.09 5.69 5.155 6.465 ;
        RECT  2.195 6.33 4.12 6.395 ;
        RECT  3.735 5.825 4.045 5.89 ;
        RECT  3.31 6.2 3.6 6.265 ;
        RECT  4.475 6.125 4.925 6.19 ;
        RECT  3.735 6.01 4.12 6.08 ;
        RECT  3.02 6.01 3.1775 6.08 ;
        RECT  4.0325 6.2 4.12 6.265 ;
        RECT  3.31 5.825 3.6 5.89 ;
        RECT  4.25 5.76 4.315 6.005 ;
        RECT  4.25 5.76 4.3725 5.8425 ;
        RECT  4.3725 5.755 4.5075 5.8225 ;
        RECT  4.12 5.69 4.185 6.465 ;
        RECT  2.5 6.2 2.79 6.265 ;
        RECT  1.9625 6.015 2.13 6.08 ;
        RECT  1.47 5.7575 1.54 6.015 ;
        RECT  1.405 6.2 1.83 6.265 ;
        RECT  2.5 6.01 2.79 6.08 ;
        RECT  1.66 6.2 1.735 6.3725 ;
        RECT  2.5 5.825 2.79 5.89 ;
        RECT  1.34 5.8225 1.4125 5.8875 ;
        RECT  3.02 5.695 3.09 6.08 ;
        RECT  2.05 5.7825 2.165 5.8475 ;
        RECT  1.275 5.69 1.34 6.465 ;
        RECT  2.13 5.69 2.195 6.465 ;
        RECT  1.12 6.26 1.1775 6.325 ;
        RECT  1.36 5.6925 1.4825 5.7575 ;
        RECT  4.9225 5.875 5.09 5.94 ;
        RECT  4.315 5.9375 4.4175 6.005 ;
        RECT  3.6 5.56 3.735 5.625 ;
        RECT  3.6 5.375 3.735 5.44 ;
        RECT  2.365 5.56 2.5 5.625 ;
        RECT  2.365 5.375 2.5 5.44 ;
        RECT  3.6 5.37 3.735 5.435 ;
        RECT  3.6 5.185 3.735 5.25 ;
        RECT  6.56 5.37 6.695 5.435 ;
        RECT  6.56 5.185 6.695 5.25 ;
        RECT  2.365 5.37 2.5 5.435 ;
        RECT  2.365 5.185 2.5 5.25 ;
        RECT  6.56 5.56 6.695 5.625 ;
        RECT  6.56 5.375 6.695 5.44 ;
        RECT  1.83 5.37 1.965 5.435 ;
        RECT  1.83 5.185 1.965 5.25 ;
        RECT  4.79 5.51 4.925 5.575 ;
        RECT  4.79 5.325 4.925 5.39 ;
        RECT  5.325 5.56 5.46 5.625 ;
        RECT  5.325 5.375 5.46 5.44 ;
        RECT  5.325 5.37 5.46 5.435 ;
        RECT  5.325 5.185 5.46 5.25 ;
        RECT  5.75 5.56 5.885 5.625 ;
        RECT  5.75 5.375 5.885 5.44 ;
        RECT  2.79 5.56 2.925 5.625 ;
        RECT  2.79 5.375 2.925 5.44 ;
        RECT  6.135 5.56 6.27 5.625 ;
        RECT  6.135 5.375 6.27 5.44 ;
        RECT  6.135 5.37 6.27 5.435 ;
        RECT  6.135 5.185 6.27 5.25 ;
        RECT  2.79 5.37 2.925 5.435 ;
        RECT  2.79 5.185 2.925 5.25 ;
        RECT  5.75 5.37 5.885 5.435 ;
        RECT  5.75 5.185 5.885 5.25 ;
        RECT  3.175 5.37 3.31 5.435 ;
        RECT  3.175 5.185 3.31 5.25 ;
        RECT  3.175 5.56 3.31 5.625 ;
        RECT  3.175 5.375 3.31 5.44 ;
        RECT  1.405 5.37 1.54 5.435 ;
        RECT  1.405 5.185 1.54 5.25 ;
        RECT  4.38 5.445 4.515 5.51 ;
        RECT  4.38 5.26 4.515 5.325 ;
        RECT  1.115 5.2475 1.18 5.3825 ;
        RECT  6.6125 5.185 6.7475 5.25 ;
        RECT  4.7975 5.075 4.9325 5.14 ;
        RECT  3.8975 5.185 4.0325 5.25 ;
        RECT  4.3725 5.6075 4.5075 5.6725 ;
        RECT  6.9775 5.185 7.1125 5.25 ;
        RECT  1.435 5.6925 1.57 5.7575 ;
        RECT  5.5175 5.55 5.6525 5.615 ;
        RECT  3.91 5.5525 4.045 5.6175 ;
        RECT  2.5125 5.5525 2.6475 5.6175 ;
        RECT  1.295 4.9875 1.43 5.0525 ;
        RECT  1.4125 5.5625 1.5475 5.6275 ;
        RECT  3.0225 5.5625 3.0875 5.6975 ;
        RECT  1.9375 5.6025 2.0725 5.6675 ;
        RECT  5.9825 5.5625 6.0475 5.6975 ;
        RECT  6.87 5.51 7.005 5.575 ;
        RECT  3.4 5.43 3.535 5.495 ;
        RECT  6.36 5.42 6.495 5.485 ;
        RECT  4.67 5.1875 4.735 5.3225 ;
        RECT  4.3725 5.6925 4.5075 5.7575 ;
        RECT  1.665 5.0775 1.73 5.2125 ;
        RECT  3.1775 5.1875 3.3125 5.2525 ;
        RECT  6.87 5.5525 7.005 5.6175 ;
        RECT  6.36 5.375 6.495 5.44 ;
        RECT  5.9475 5.6925 6.0825 5.7575 ;
        RECT  1.245 5.6925 1.38 5.7575 ;
        RECT  3.91 5.5525 4.045 5.6175 ;
        RECT  2.9875 5.6925 3.1225 5.7575 ;
        RECT  2.7875 5.1875 2.9225 5.2525 ;
        RECT  2.7875 5.375 2.9225 5.44 ;
        RECT  3.4 5.375 3.535 5.44 ;
        RECT  5.7475 5.185 5.8825 5.25 ;
        RECT  5.7475 5.375 5.8825 5.44 ;
        RECT  1.115 4.985 1.18 5.76 ;
        RECT  4.185 5.055 7.08 5.12 ;
        RECT  6.695 5.56 7.005 5.625 ;
        RECT  6.27 5.185 6.56 5.25 ;
        RECT  5.46 5.185 5.75 5.25 ;
        RECT  7.0825 5.325 7.145 5.3975 ;
        RECT  6.695 5.37 7.08 5.44 ;
        RECT  5.46 5.37 5.75 5.44 ;
        RECT  5.98 5.37 6.1375 5.44 ;
        RECT  6.27 5.56 6.56 5.625 ;
        RECT  5.46 5.56 5.75 5.625 ;
        RECT  5.98 5.37 6.05 5.755 ;
        RECT  7.08 4.985 7.145 5.76 ;
        RECT  5.09 4.985 5.155 5.76 ;
        RECT  2.195 5.055 4.12 5.12 ;
        RECT  3.735 5.56 4.045 5.625 ;
        RECT  3.31 5.185 3.6 5.25 ;
        RECT  4.475 5.26 4.925 5.325 ;
        RECT  3.735 5.37 4.12 5.44 ;
        RECT  3.02 5.37 3.1775 5.44 ;
        RECT  4.0325 5.185 4.12 5.25 ;
        RECT  3.31 5.56 3.6 5.625 ;
        RECT  4.25 5.445 4.315 5.69 ;
        RECT  4.25 5.6075 4.3725 5.69 ;
        RECT  4.3725 5.6275 4.5075 5.695 ;
        RECT  4.12 4.985 4.185 5.76 ;
        RECT  2.5 5.185 2.79 5.25 ;
        RECT  1.9625 5.37 2.13 5.435 ;
        RECT  1.47 5.435 1.54 5.6925 ;
        RECT  1.405 5.185 1.83 5.25 ;
        RECT  2.5 5.37 2.79 5.44 ;
        RECT  1.66 5.0775 1.735 5.25 ;
        RECT  2.5 5.56 2.79 5.625 ;
        RECT  1.34 5.5625 1.4125 5.6275 ;
        RECT  3.02 5.37 3.09 5.755 ;
        RECT  2.05 5.6025 2.165 5.6675 ;
        RECT  1.275 4.985 1.34 5.76 ;
        RECT  2.13 4.985 2.195 5.76 ;
        RECT  1.12 5.125 1.1775 5.19 ;
        RECT  1.36 5.6925 1.4825 5.7575 ;
        RECT  4.9225 5.51 5.09 5.575 ;
        RECT  4.315 5.445 4.4175 5.5125 ;
        RECT  7.855 19.0025 7.92 19.0675 ;
        RECT  7.8875 19.0025 11.1625 19.0675 ;
        RECT  7.855 19.035 7.92 19.575 ;
        RECT  7.855 21.4125 7.92 21.4775 ;
        RECT  7.8875 21.4125 11.1625 21.4775 ;
        RECT  7.855 20.905 7.92 21.445 ;
        RECT  7.855 21.6925 7.92 21.7575 ;
        RECT  7.8875 21.6925 11.1625 21.7575 ;
        RECT  7.855 21.725 7.92 22.265 ;
        RECT  7.855 24.1025 7.92 24.1675 ;
        RECT  7.8875 24.1025 11.1625 24.1675 ;
        RECT  7.855 23.595 7.92 24.135 ;
        RECT  7.855 24.3825 7.92 24.4475 ;
        RECT  7.8875 24.3825 11.1625 24.4475 ;
        RECT  7.855 24.415 7.92 24.955 ;
        RECT  7.855 26.7925 7.92 26.8575 ;
        RECT  7.8875 26.7925 11.1625 26.8575 ;
        RECT  7.855 26.285 7.92 26.825 ;
        RECT  7.855 27.0725 7.92 27.1375 ;
        RECT  7.8875 27.0725 11.1625 27.1375 ;
        RECT  7.855 27.105 7.92 27.645 ;
        RECT  7.855 29.4825 7.92 29.5475 ;
        RECT  7.8875 29.4825 11.1625 29.5475 ;
        RECT  7.855 28.975 7.92 29.515 ;
        RECT  7.855 29.7625 7.92 29.8275 ;
        RECT  7.8875 29.7625 11.1625 29.8275 ;
        RECT  7.855 29.795 7.92 30.335 ;
        RECT  7.855 32.1725 7.92 32.2375 ;
        RECT  7.8875 32.1725 11.1625 32.2375 ;
        RECT  7.855 31.665 7.92 32.205 ;
        RECT  7.855 32.4525 7.92 32.5175 ;
        RECT  7.8875 32.4525 11.1625 32.5175 ;
        RECT  7.855 32.485 7.92 33.025 ;
        RECT  7.855 34.8625 7.92 34.9275 ;
        RECT  7.8875 34.8625 11.1625 34.9275 ;
        RECT  7.855 34.355 7.92 34.895 ;
        RECT  7.855 35.1425 7.92 35.2075 ;
        RECT  7.8875 35.1425 11.1625 35.2075 ;
        RECT  7.855 35.175 7.92 35.715 ;
        RECT  7.855 37.5525 7.92 37.6175 ;
        RECT  7.8875 37.5525 11.1625 37.6175 ;
        RECT  7.855 37.045 7.92 37.585 ;
        RECT  7.855 37.8325 7.92 37.8975 ;
        RECT  7.8875 37.8325 11.1625 37.8975 ;
        RECT  7.855 37.865 7.92 38.405 ;
        RECT  7.855 40.2425 7.92 40.3075 ;
        RECT  7.8875 40.2425 11.1625 40.3075 ;
        RECT  7.855 39.735 7.92 40.275 ;
        RECT  8.5425 8.73 8.6075 8.865 ;
        RECT  8.3325 10.165 8.3975 10.3 ;
        RECT  8.1225 14.11 8.1875 14.245 ;
        RECT  7.9125 15.545 7.9775 15.68 ;
        RECT  10.3625 3.6 10.4275 3.735 ;
        RECT  9.9425 1.415 10.0075 1.55 ;
        RECT  10.1525 2.9625 10.2175 3.0975 ;
        RECT  10.3625 41.1 10.4275 41.235 ;
        RECT  10.5725 10.1025 10.6375 10.2375 ;
        RECT  10.7825 14.1275 10.8475 14.2625 ;
        RECT  0.98 7.63 1.115 7.695 ;
        RECT  5.725 41.53 5.79 41.595 ;
        RECT  5.725 40.415 5.79 41.5625 ;
        RECT  5.7575 41.53 9.8275 41.595 ;
        RECT  9.7325 41.53 9.7975 41.665 ;
        RECT  7.08 4.7925 7.145 4.8575 ;
        RECT  0.0 4.7925 7.1125 4.8575 ;
        RECT  7.08 4.825 7.145 5.02 ;
        RECT  8.89 40.545 9.095 40.68 ;
        RECT  11.77 40.5475 11.905 40.6125 ;
        RECT  12.475 40.5475 12.61 40.6125 ;
        RECT  10.995 40.5475 11.13 40.6125 ;
        RECT  9.385 0.355 9.59 0.49 ;
        RECT  11.8025 0.355 11.8675 0.49 ;
        RECT  11.8025 0.355 11.8675 0.49 ;
        RECT  7.755 21.555 7.89 21.62 ;
        RECT  7.755 24.245 7.89 24.31 ;
        RECT  7.755 26.935 7.89 27.0 ;
        RECT  7.755 29.625 7.89 29.69 ;
        RECT  7.755 32.315 7.89 32.38 ;
        RECT  7.755 35.005 7.89 35.07 ;
        RECT  7.755 37.695 7.89 37.76 ;
        RECT  7.755 40.385 7.89 40.45 ;
        RECT  8.89 13.4125 9.095 13.5475 ;
        RECT  8.89 18.7925 9.095 18.9275 ;
        RECT  7.28 7.81 7.415 7.875 ;
        RECT  8.89 7.8075 9.095 7.9425 ;
        RECT  7.28 6.4 7.415 6.465 ;
        RECT  8.89 6.3975 9.095 6.5325 ;
        RECT  7.28 6.4 7.415 6.465 ;
        RECT  8.89 6.3975 9.095 6.5325 ;
        RECT  7.28 4.99 7.415 5.055 ;
        RECT  8.89 4.9875 9.095 5.1225 ;
        RECT  -2.49 17.335 -2.3225 17.4 ;
        RECT  -3.7575 17.335 -3.59 17.4 ;
        RECT  -3.9975 14.715 -3.9325 15.205 ;
        RECT  -4.1525 14.715 -4.0875 15.415 ;
        RECT  -5.5625 14.715 -5.4975 15.625 ;
        RECT  -4.5475 14.715 -4.4825 15.835 ;
        RECT  -1.325 15.345 -1.26 16.185 ;
        RECT  -0.795 15.975 -0.73 16.185 ;
        RECT  -2.12 15.975 -2.055 16.185 ;
        RECT  -2.6425 15.345 -2.5775 16.185 ;
        RECT  -2.7825 15.555 -2.7175 16.185 ;
        RECT  -4.025 15.975 -3.96 16.185 ;
        RECT  -3.5025 15.765 -3.4375 16.185 ;
        RECT  -3.3625 15.555 -3.2975 16.185 ;
        RECT  -2.49 17.895 -2.425 19.505 ;
        RECT  -3.655 19.015 -3.59 19.295 ;
        RECT  -0.965 18.455 -0.9 19.715 ;
        RECT  -0.3825 23.7575 -0.14 23.8225 ;
        RECT  -1.7275 8.415 -1.6625 20.065 ;
        RECT  -4.4175 17.335 -4.3525 19.925 ;
        RECT  -5.73 14.4425 -1.6625 14.5075 ;
        RECT  -0.3825 8.415 -0.3175 20.835 ;
        RECT  -3.0725 17.335 -3.0075 20.695 ;
        RECT  -5.3775 8.4775 -2.0525 8.5425 ;
        RECT  -5.73 8.4475 -3.615 8.5125 ;
        RECT  -5.73 14.445 -3.615 14.51 ;
        RECT  -5.19 10.965 -5.125 11.1 ;
        RECT  -5.375 10.965 -5.31 11.1 ;
        RECT  -5.19 9.73 -5.125 9.865 ;
        RECT  -5.375 9.73 -5.31 9.865 ;
        RECT  -5.38 10.965 -5.315 11.1 ;
        RECT  -5.565 10.965 -5.5 11.1 ;
        RECT  -5.38 13.925 -5.315 14.06 ;
        RECT  -5.565 13.925 -5.5 14.06 ;
        RECT  -5.38 9.73 -5.315 9.865 ;
        RECT  -5.565 9.73 -5.5 9.865 ;
        RECT  -5.19 13.925 -5.125 14.06 ;
        RECT  -5.375 13.925 -5.31 14.06 ;
        RECT  -5.38 9.195 -5.315 9.33 ;
        RECT  -5.565 9.195 -5.5 9.33 ;
        RECT  -5.24 12.155 -5.175 12.29 ;
        RECT  -5.425 12.155 -5.36 12.29 ;
        RECT  -5.19 12.69 -5.125 12.825 ;
        RECT  -5.375 12.69 -5.31 12.825 ;
        RECT  -5.38 12.69 -5.315 12.825 ;
        RECT  -5.565 12.69 -5.5 12.825 ;
        RECT  -5.19 13.115 -5.125 13.25 ;
        RECT  -5.375 13.115 -5.31 13.25 ;
        RECT  -5.19 10.155 -5.125 10.29 ;
        RECT  -5.375 10.155 -5.31 10.29 ;
        RECT  -5.19 13.5 -5.125 13.635 ;
        RECT  -5.375 13.5 -5.31 13.635 ;
        RECT  -5.38 13.5 -5.315 13.635 ;
        RECT  -5.565 13.5 -5.5 13.635 ;
        RECT  -5.38 10.155 -5.315 10.29 ;
        RECT  -5.565 10.155 -5.5 10.29 ;
        RECT  -5.38 13.115 -5.315 13.25 ;
        RECT  -5.565 13.115 -5.5 13.25 ;
        RECT  -5.38 10.54 -5.315 10.675 ;
        RECT  -5.565 10.54 -5.5 10.675 ;
        RECT  -5.19 10.54 -5.125 10.675 ;
        RECT  -5.375 10.54 -5.31 10.675 ;
        RECT  -5.38 8.77 -5.315 8.905 ;
        RECT  -5.565 8.77 -5.5 8.905 ;
        RECT  -5.305 11.745 -5.24 11.88 ;
        RECT  -5.49 11.745 -5.425 11.88 ;
        RECT  -5.5025 8.48 -5.3675 8.545 ;
        RECT  -5.565 13.9775 -5.5 14.1125 ;
        RECT  -5.675 12.1625 -5.61 12.2975 ;
        RECT  -5.565 11.2625 -5.5 11.3975 ;
        RECT  -5.1425 11.7375 -5.0775 11.8725 ;
        RECT  -5.565 14.3425 -5.5 14.4775 ;
        RECT  -5.0575 8.8 -4.9925 8.935 ;
        RECT  -5.2 12.8825 -5.135 13.0175 ;
        RECT  -5.1975 11.275 -5.1325 11.41 ;
        RECT  -5.1975 9.8775 -5.1325 10.0125 ;
        RECT  -5.7625 8.66 -5.6975 8.795 ;
        RECT  -5.1875 8.7775 -5.1225 8.9125 ;
        RECT  -5.1875 10.3875 -5.0525 10.4525 ;
        RECT  -5.1475 9.3025 -5.0825 9.4375 ;
        RECT  -5.1875 13.3475 -5.0525 13.4125 ;
        RECT  -5.24 14.235 -5.175 14.37 ;
        RECT  -5.32 10.765 -5.255 10.9 ;
        RECT  -5.33 13.725 -5.265 13.86 ;
        RECT  -5.5625 12.035 -5.4275 12.1 ;
        RECT  -5.0575 11.7375 -4.9925 11.8725 ;
        RECT  -5.6725 9.03 -5.5375 9.095 ;
        RECT  -5.5625 10.5425 -5.4975 10.6775 ;
        RECT  -5.1975 14.235 -5.1325 14.37 ;
        RECT  -5.375 13.725 -5.31 13.86 ;
        RECT  -5.0575 13.3125 -4.9925 13.4475 ;
        RECT  -5.0575 8.61 -4.9925 8.745 ;
        RECT  -5.1975 11.275 -5.1325 11.41 ;
        RECT  -5.0575 10.3525 -4.9925 10.4875 ;
        RECT  -5.5625 10.1525 -5.4975 10.2875 ;
        RECT  -5.375 10.1525 -5.31 10.2875 ;
        RECT  -5.375 10.765 -5.31 10.9 ;
        RECT  -5.565 13.1125 -5.5 13.2475 ;
        RECT  -5.375 13.1125 -5.31 13.2475 ;
        RECT  -5.765 8.48 -4.99 8.545 ;
        RECT  -5.695 11.55 -5.63 14.445 ;
        RECT  -5.19 14.06 -5.125 14.37 ;
        RECT  -5.565 13.635 -5.5 13.925 ;
        RECT  -5.565 12.825 -5.5 13.115 ;
        RECT  -5.425 14.4475 -5.3525 14.51 ;
        RECT  -5.38 14.06 -5.31 14.445 ;
        RECT  -5.38 12.825 -5.31 13.115 ;
        RECT  -5.38 13.345 -5.31 13.5025 ;
        RECT  -5.19 13.635 -5.125 13.925 ;
        RECT  -5.19 12.825 -5.125 13.115 ;
        RECT  -5.38 13.345 -4.995 13.415 ;
        RECT  -5.765 14.445 -4.99 14.51 ;
        RECT  -5.765 12.455 -4.99 12.52 ;
        RECT  -5.695 9.56 -5.63 11.485 ;
        RECT  -5.19 11.1 -5.125 11.41 ;
        RECT  -5.565 10.675 -5.5 10.965 ;
        RECT  -5.49 11.84 -5.425 12.29 ;
        RECT  -5.38 11.1 -5.31 11.485 ;
        RECT  -5.38 10.385 -5.31 10.5425 ;
        RECT  -5.565 11.3975 -5.5 11.485 ;
        RECT  -5.19 10.675 -5.125 10.965 ;
        RECT  -5.305 11.615 -5.06 11.68 ;
        RECT  -5.1425 11.615 -5.06 11.7375 ;
        RECT  -5.1225 11.7375 -5.055 11.8725 ;
        RECT  -5.765 11.485 -4.99 11.55 ;
        RECT  -5.565 9.865 -5.5 10.155 ;
        RECT  -5.38 9.3275 -5.315 9.495 ;
        RECT  -5.315 8.835 -5.0575 8.905 ;
        RECT  -5.565 8.77 -5.5 9.195 ;
        RECT  -5.38 9.865 -5.31 10.155 ;
        RECT  -5.6725 9.025 -5.5 9.1 ;
        RECT  -5.19 9.865 -5.125 10.155 ;
        RECT  -5.1875 8.705 -5.1225 8.7775 ;
        RECT  -5.38 10.385 -4.995 10.455 ;
        RECT  -5.1475 9.415 -5.0825 9.53 ;
        RECT  -5.765 8.64 -4.99 8.705 ;
        RECT  -5.765 9.495 -4.99 9.56 ;
        RECT  -5.625 8.485 -5.56 8.5425 ;
        RECT  -5.0575 8.725 -4.9925 8.8475 ;
        RECT  -5.24 12.2875 -5.175 12.455 ;
        RECT  -5.305 11.68 -5.2375 11.7825 ;
        RECT  -4.925 10.965 -4.86 11.1 ;
        RECT  -4.74 10.965 -4.675 11.1 ;
        RECT  -4.925 9.73 -4.86 9.865 ;
        RECT  -4.74 9.73 -4.675 9.865 ;
        RECT  -4.735 10.965 -4.67 11.1 ;
        RECT  -4.55 10.965 -4.485 11.1 ;
        RECT  -4.735 13.925 -4.67 14.06 ;
        RECT  -4.55 13.925 -4.485 14.06 ;
        RECT  -4.735 9.73 -4.67 9.865 ;
        RECT  -4.55 9.73 -4.485 9.865 ;
        RECT  -4.925 13.925 -4.86 14.06 ;
        RECT  -4.74 13.925 -4.675 14.06 ;
        RECT  -4.735 9.195 -4.67 9.33 ;
        RECT  -4.55 9.195 -4.485 9.33 ;
        RECT  -4.875 12.155 -4.81 12.29 ;
        RECT  -4.69 12.155 -4.625 12.29 ;
        RECT  -4.925 12.69 -4.86 12.825 ;
        RECT  -4.74 12.69 -4.675 12.825 ;
        RECT  -4.735 12.69 -4.67 12.825 ;
        RECT  -4.55 12.69 -4.485 12.825 ;
        RECT  -4.925 13.115 -4.86 13.25 ;
        RECT  -4.74 13.115 -4.675 13.25 ;
        RECT  -4.925 10.155 -4.86 10.29 ;
        RECT  -4.74 10.155 -4.675 10.29 ;
        RECT  -4.925 13.5 -4.86 13.635 ;
        RECT  -4.74 13.5 -4.675 13.635 ;
        RECT  -4.735 13.5 -4.67 13.635 ;
        RECT  -4.55 13.5 -4.485 13.635 ;
        RECT  -4.735 10.155 -4.67 10.29 ;
        RECT  -4.55 10.155 -4.485 10.29 ;
        RECT  -4.735 13.115 -4.67 13.25 ;
        RECT  -4.55 13.115 -4.485 13.25 ;
        RECT  -4.735 10.54 -4.67 10.675 ;
        RECT  -4.55 10.54 -4.485 10.675 ;
        RECT  -4.925 10.54 -4.86 10.675 ;
        RECT  -4.74 10.54 -4.675 10.675 ;
        RECT  -4.735 8.77 -4.67 8.905 ;
        RECT  -4.55 8.77 -4.485 8.905 ;
        RECT  -4.81 11.745 -4.745 11.88 ;
        RECT  -4.625 11.745 -4.56 11.88 ;
        RECT  -4.6825 8.48 -4.5475 8.545 ;
        RECT  -4.55 13.9775 -4.485 14.1125 ;
        RECT  -4.44 12.1625 -4.375 12.2975 ;
        RECT  -4.55 11.2625 -4.485 11.3975 ;
        RECT  -4.9725 11.7375 -4.9075 11.8725 ;
        RECT  -4.55 14.3425 -4.485 14.4775 ;
        RECT  -5.0575 8.8 -4.9925 8.935 ;
        RECT  -4.915 12.8825 -4.85 13.0175 ;
        RECT  -4.9175 11.275 -4.8525 11.41 ;
        RECT  -4.9175 9.8775 -4.8525 10.0125 ;
        RECT  -4.3525 8.66 -4.2875 8.795 ;
        RECT  -4.9275 8.7775 -4.8625 8.9125 ;
        RECT  -4.9975 10.3875 -4.8625 10.4525 ;
        RECT  -4.9675 9.3025 -4.9025 9.4375 ;
        RECT  -4.9975 13.3475 -4.8625 13.4125 ;
        RECT  -4.875 14.235 -4.81 14.37 ;
        RECT  -4.795 10.765 -4.73 10.9 ;
        RECT  -4.785 13.725 -4.72 13.86 ;
        RECT  -4.6225 12.035 -4.4875 12.1 ;
        RECT  -5.0575 11.7375 -4.9925 11.8725 ;
        RECT  -4.5125 9.03 -4.3775 9.095 ;
        RECT  -4.5525 10.5425 -4.4875 10.6775 ;
        RECT  -4.9175 14.235 -4.8525 14.37 ;
        RECT  -4.74 13.725 -4.675 13.86 ;
        RECT  -5.0575 13.3125 -4.9925 13.4475 ;
        RECT  -5.0575 8.61 -4.9925 8.745 ;
        RECT  -4.9175 11.275 -4.8525 11.41 ;
        RECT  -5.0575 10.3525 -4.9925 10.4875 ;
        RECT  -4.5525 10.1525 -4.4875 10.2875 ;
        RECT  -4.74 10.1525 -4.675 10.2875 ;
        RECT  -4.74 10.765 -4.675 10.9 ;
        RECT  -4.55 13.1125 -4.485 13.2475 ;
        RECT  -4.74 13.1125 -4.675 13.2475 ;
        RECT  -5.06 8.48 -4.285 8.545 ;
        RECT  -4.42 11.55 -4.355 14.445 ;
        RECT  -4.925 14.06 -4.86 14.37 ;
        RECT  -4.55 13.635 -4.485 13.925 ;
        RECT  -4.55 12.825 -4.485 13.115 ;
        RECT  -4.6975 14.4475 -4.625 14.51 ;
        RECT  -4.74 14.06 -4.67 14.445 ;
        RECT  -4.74 12.825 -4.67 13.115 ;
        RECT  -4.74 13.345 -4.67 13.5025 ;
        RECT  -4.925 13.635 -4.86 13.925 ;
        RECT  -4.925 12.825 -4.86 13.115 ;
        RECT  -5.055 13.345 -4.67 13.415 ;
        RECT  -5.06 14.445 -4.285 14.51 ;
        RECT  -5.06 12.455 -4.285 12.52 ;
        RECT  -4.42 9.56 -4.355 11.485 ;
        RECT  -4.925 11.1 -4.86 11.41 ;
        RECT  -4.55 10.675 -4.485 10.965 ;
        RECT  -4.625 11.84 -4.56 12.29 ;
        RECT  -4.74 11.1 -4.67 11.485 ;
        RECT  -4.74 10.385 -4.67 10.5425 ;
        RECT  -4.55 11.3975 -4.485 11.485 ;
        RECT  -4.925 10.675 -4.86 10.965 ;
        RECT  -4.99 11.615 -4.745 11.68 ;
        RECT  -4.99 11.615 -4.9075 11.7375 ;
        RECT  -4.995 11.7375 -4.9275 11.8725 ;
        RECT  -5.06 11.485 -4.285 11.55 ;
        RECT  -4.55 9.865 -4.485 10.155 ;
        RECT  -4.735 9.3275 -4.67 9.495 ;
        RECT  -4.9925 8.835 -4.735 8.905 ;
        RECT  -4.55 8.77 -4.485 9.195 ;
        RECT  -4.74 9.865 -4.67 10.155 ;
        RECT  -4.55 9.025 -4.3775 9.1 ;
        RECT  -4.925 9.865 -4.86 10.155 ;
        RECT  -4.9275 8.705 -4.8625 8.7775 ;
        RECT  -5.055 10.385 -4.67 10.455 ;
        RECT  -4.9675 9.415 -4.9025 9.53 ;
        RECT  -5.06 8.64 -4.285 8.705 ;
        RECT  -5.06 9.495 -4.285 9.56 ;
        RECT  -4.49 8.485 -4.425 8.5425 ;
        RECT  -5.0575 8.725 -4.9925 8.8475 ;
        RECT  -4.875 12.2875 -4.81 12.455 ;
        RECT  -4.8125 11.68 -4.745 11.7825 ;
        RECT  -3.78 10.965 -3.715 11.1 ;
        RECT  -3.965 10.965 -3.9 11.1 ;
        RECT  -3.78 9.73 -3.715 9.865 ;
        RECT  -3.965 9.73 -3.9 9.865 ;
        RECT  -3.97 10.965 -3.905 11.1 ;
        RECT  -4.155 10.965 -4.09 11.1 ;
        RECT  -3.97 13.925 -3.905 14.06 ;
        RECT  -4.155 13.925 -4.09 14.06 ;
        RECT  -3.97 9.73 -3.905 9.865 ;
        RECT  -4.155 9.73 -4.09 9.865 ;
        RECT  -3.78 13.925 -3.715 14.06 ;
        RECT  -3.965 13.925 -3.9 14.06 ;
        RECT  -3.97 9.195 -3.905 9.33 ;
        RECT  -4.155 9.195 -4.09 9.33 ;
        RECT  -3.83 12.155 -3.765 12.29 ;
        RECT  -4.015 12.155 -3.95 12.29 ;
        RECT  -3.78 12.69 -3.715 12.825 ;
        RECT  -3.965 12.69 -3.9 12.825 ;
        RECT  -3.97 12.69 -3.905 12.825 ;
        RECT  -4.155 12.69 -4.09 12.825 ;
        RECT  -3.78 13.115 -3.715 13.25 ;
        RECT  -3.965 13.115 -3.9 13.25 ;
        RECT  -3.78 10.155 -3.715 10.29 ;
        RECT  -3.965 10.155 -3.9 10.29 ;
        RECT  -3.78 13.5 -3.715 13.635 ;
        RECT  -3.965 13.5 -3.9 13.635 ;
        RECT  -3.97 13.5 -3.905 13.635 ;
        RECT  -4.155 13.5 -4.09 13.635 ;
        RECT  -3.97 10.155 -3.905 10.29 ;
        RECT  -4.155 10.155 -4.09 10.29 ;
        RECT  -3.97 13.115 -3.905 13.25 ;
        RECT  -4.155 13.115 -4.09 13.25 ;
        RECT  -3.97 10.54 -3.905 10.675 ;
        RECT  -4.155 10.54 -4.09 10.675 ;
        RECT  -3.78 10.54 -3.715 10.675 ;
        RECT  -3.965 10.54 -3.9 10.675 ;
        RECT  -3.97 8.77 -3.905 8.905 ;
        RECT  -4.155 8.77 -4.09 8.905 ;
        RECT  -3.895 11.745 -3.83 11.88 ;
        RECT  -4.08 11.745 -4.015 11.88 ;
        RECT  -4.0925 8.48 -3.9575 8.545 ;
        RECT  -4.155 13.9775 -4.09 14.1125 ;
        RECT  -4.265 12.1625 -4.2 12.2975 ;
        RECT  -4.155 11.2625 -4.09 11.3975 ;
        RECT  -3.7325 11.7375 -3.6675 11.8725 ;
        RECT  -4.155 14.3425 -4.09 14.4775 ;
        RECT  -3.6475 8.8 -3.5825 8.935 ;
        RECT  -3.79 12.8825 -3.725 13.0175 ;
        RECT  -3.7875 11.275 -3.7225 11.41 ;
        RECT  -3.7875 9.8775 -3.7225 10.0125 ;
        RECT  -4.3525 8.66 -4.2875 8.795 ;
        RECT  -3.7775 8.7775 -3.7125 8.9125 ;
        RECT  -3.7775 10.3875 -3.6425 10.4525 ;
        RECT  -3.7375 9.3025 -3.6725 9.4375 ;
        RECT  -3.7775 13.3475 -3.6425 13.4125 ;
        RECT  -3.83 14.235 -3.765 14.37 ;
        RECT  -3.91 10.765 -3.845 10.9 ;
        RECT  -3.92 13.725 -3.855 13.86 ;
        RECT  -4.1525 12.035 -4.0175 12.1 ;
        RECT  -3.6475 11.7375 -3.5825 11.8725 ;
        RECT  -4.2625 9.03 -4.1275 9.095 ;
        RECT  -4.1525 10.5425 -4.0875 10.6775 ;
        RECT  -3.7875 14.235 -3.7225 14.37 ;
        RECT  -3.965 13.725 -3.9 13.86 ;
        RECT  -3.6475 13.3125 -3.5825 13.4475 ;
        RECT  -3.6475 8.61 -3.5825 8.745 ;
        RECT  -3.7875 11.275 -3.7225 11.41 ;
        RECT  -3.6475 10.3525 -3.5825 10.4875 ;
        RECT  -4.1525 10.1525 -4.0875 10.2875 ;
        RECT  -3.965 10.1525 -3.9 10.2875 ;
        RECT  -3.965 10.765 -3.9 10.9 ;
        RECT  -4.155 13.1125 -4.09 13.2475 ;
        RECT  -3.965 13.1125 -3.9 13.2475 ;
        RECT  -4.355 8.48 -3.58 8.545 ;
        RECT  -4.285 11.55 -4.22 14.445 ;
        RECT  -3.78 14.06 -3.715 14.37 ;
        RECT  -4.155 13.635 -4.09 13.925 ;
        RECT  -4.155 12.825 -4.09 13.115 ;
        RECT  -4.015 14.4475 -3.9425 14.51 ;
        RECT  -3.97 14.06 -3.9 14.445 ;
        RECT  -3.97 12.825 -3.9 13.115 ;
        RECT  -3.97 13.345 -3.9 13.5025 ;
        RECT  -3.78 13.635 -3.715 13.925 ;
        RECT  -3.78 12.825 -3.715 13.115 ;
        RECT  -3.97 13.345 -3.585 13.415 ;
        RECT  -4.355 14.445 -3.58 14.51 ;
        RECT  -4.355 12.455 -3.58 12.52 ;
        RECT  -4.285 9.56 -4.22 11.485 ;
        RECT  -3.78 11.1 -3.715 11.41 ;
        RECT  -4.155 10.675 -4.09 10.965 ;
        RECT  -4.08 11.84 -4.015 12.29 ;
        RECT  -3.97 11.1 -3.9 11.485 ;
        RECT  -3.97 10.385 -3.9 10.5425 ;
        RECT  -4.155 11.3975 -4.09 11.485 ;
        RECT  -3.78 10.675 -3.715 10.965 ;
        RECT  -3.895 11.615 -3.65 11.68 ;
        RECT  -3.7325 11.615 -3.65 11.7375 ;
        RECT  -3.7125 11.7375 -3.645 11.8725 ;
        RECT  -4.355 11.485 -3.58 11.55 ;
        RECT  -4.155 9.865 -4.09 10.155 ;
        RECT  -3.97 9.3275 -3.905 9.495 ;
        RECT  -3.905 8.835 -3.6475 8.905 ;
        RECT  -4.155 8.77 -4.09 9.195 ;
        RECT  -3.97 9.865 -3.9 10.155 ;
        RECT  -4.2625 9.025 -4.09 9.1 ;
        RECT  -3.78 9.865 -3.715 10.155 ;
        RECT  -3.7775 8.705 -3.7125 8.7775 ;
        RECT  -3.97 10.385 -3.585 10.455 ;
        RECT  -3.7375 9.415 -3.6725 9.53 ;
        RECT  -4.355 8.64 -3.58 8.705 ;
        RECT  -4.355 9.495 -3.58 9.56 ;
        RECT  -4.215 8.485 -4.15 8.5425 ;
        RECT  -3.6475 8.725 -3.5825 8.8475 ;
        RECT  -3.83 12.2875 -3.765 12.455 ;
        RECT  -3.895 11.68 -3.8275 11.7825 ;
        RECT  -0.3825 13.585 -0.3175 14.715 ;
        RECT  -1.7275 13.585 -1.6625 14.715 ;
        RECT  -1.6625 14.5825 -1.2975 14.6475 ;
        RECT  -0.5175 14.5825 -0.3825 14.6475 ;
        RECT  -1.4325 13.8425 -0.485 13.9075 ;
        RECT  -1.4325 14.2225 -0.485 14.2875 ;
        RECT  -0.965 13.585 -0.9 13.62 ;
        RECT  -0.965 14.2875 -0.9 14.715 ;
        RECT  -0.7225 13.6525 -0.5875 13.7175 ;
        RECT  -0.7225 13.8425 -0.5875 13.9075 ;
        RECT  -0.7225 14.0325 -0.5875 14.0975 ;
        RECT  -0.7225 14.2225 -0.5875 14.2875 ;
        RECT  -0.7225 14.4125 -0.5875 14.4775 ;
        RECT  -0.855 13.6525 -0.79 13.7175 ;
        RECT  -0.855 14.0325 -0.79 14.0975 ;
        RECT  -0.855 14.0325 -0.79 14.0975 ;
        RECT  -0.855 14.4125 -0.79 14.4775 ;
        RECT  -0.7875 13.6525 -0.5875 13.7175 ;
        RECT  -0.8225 13.6525 -0.7875 13.7175 ;
        RECT  -0.855 13.685 -0.79 14.065 ;
        RECT  -0.8225 14.0325 -0.5875 14.0975 ;
        RECT  -0.7875 14.0325 -0.5875 14.0975 ;
        RECT  -0.8225 14.0325 -0.7875 14.0975 ;
        RECT  -0.855 14.065 -0.79 14.445 ;
        RECT  -0.8225 14.4125 -0.5875 14.4775 ;
        RECT  -0.5225 13.8425 -0.4575 13.9075 ;
        RECT  -0.5225 14.2225 -0.4575 14.2875 ;
        RECT  -0.5875 13.8425 -0.5225 13.9075 ;
        RECT  -0.5225 13.8425 -0.49 13.9075 ;
        RECT  -0.5225 13.875 -0.4575 14.255 ;
        RECT  -0.5875 14.2225 -0.49 14.2875 ;
        RECT  -1.5725 13.6525 -1.2975 13.7175 ;
        RECT  -1.5725 13.8425 -1.2975 13.9075 ;
        RECT  -1.5725 14.0325 -1.2975 14.0975 ;
        RECT  -1.5725 14.2225 -1.2975 14.2875 ;
        RECT  -1.5725 14.4125 -1.2975 14.4775 ;
        RECT  -1.705 13.6525 -1.64 13.7175 ;
        RECT  -1.705 14.0325 -1.64 14.0975 ;
        RECT  -1.705 14.0325 -1.64 14.0975 ;
        RECT  -1.705 14.4125 -1.64 14.4775 ;
        RECT  -1.6375 13.6525 -1.3675 13.7175 ;
        RECT  -1.6725 13.6525 -1.6375 13.7175 ;
        RECT  -1.705 13.685 -1.64 14.065 ;
        RECT  -1.6725 14.0325 -1.3675 14.0975 ;
        RECT  -1.6375 14.0325 -1.3675 14.0975 ;
        RECT  -1.6725 14.0325 -1.6375 14.0975 ;
        RECT  -1.705 14.065 -1.64 14.445 ;
        RECT  -1.6725 14.4125 -1.3675 14.4775 ;
        RECT  -1.2325 13.8425 -1.1675 13.9075 ;
        RECT  -1.2325 14.2225 -1.1675 14.2875 ;
        RECT  -1.3675 13.8425 -1.2325 13.9075 ;
        RECT  -1.2325 13.8425 -1.2 13.9075 ;
        RECT  -1.2325 13.875 -1.1675 14.255 ;
        RECT  -1.3675 14.2225 -1.2 14.2875 ;
        RECT  -1.5725 14.5825 -1.2975 14.6475 ;
        RECT  -0.5875 14.5825 -0.4525 14.6475 ;
        RECT  -0.965 13.62 -0.9 13.755 ;
        RECT  -0.3825 8.415 -0.3175 9.745 ;
        RECT  -1.7275 8.415 -1.6625 9.745 ;
        RECT  -0.8675 9.575 -0.8025 9.745 ;
        RECT  -0.9975 8.995 -0.9325 9.745 ;
        RECT  -1.695 8.4825 -1.4125 8.5475 ;
        RECT  -0.4525 9.0625 -0.35 9.1275 ;
        RECT  -1.6625 9.6125 -1.4125 9.6775 ;
        RECT  -1.6625 9.2325 -1.4125 9.2975 ;
        RECT  -0.4525 9.6125 -0.3175 9.6775 ;
        RECT  -0.4525 9.2325 -0.3175 9.2975 ;
        RECT  -0.6525 9.6125 -0.5175 9.6775 ;
        RECT  -0.6525 9.4225 -0.5175 9.4875 ;
        RECT  -0.6525 9.4225 -0.5175 9.4875 ;
        RECT  -0.6525 9.2325 -0.5175 9.2975 ;
        RECT  -1.2575 9.6125 -1.1225 9.6775 ;
        RECT  -1.2575 9.4225 -1.1225 9.4875 ;
        RECT  -1.2575 9.2325 -1.1225 9.2975 ;
        RECT  -1.2575 9.0325 -1.1225 9.0975 ;
        RECT  -1.2575 8.8425 -1.1225 8.9075 ;
        RECT  -1.2575 8.6525 -1.1225 8.7175 ;
        RECT  -1.4125 8.4825 -1.2775 8.5475 ;
        RECT  -0.4525 9.0625 -0.3175 9.1275 ;
        RECT  -0.7925 9.575 -0.7275 9.71 ;
        RECT  -0.9225 8.995 -0.8575 9.13 ;
        RECT  -0.8675 9.4225 -0.8025 9.4875 ;
        RECT  -0.8675 8.415 -0.8025 9.455 ;
        RECT  -1.2175 9.4225 -0.835 9.4875 ;
        RECT  -1.4125 8.8425 -1.2775 8.9075 ;
        RECT  -0.8675 8.84 -0.8025 8.91 ;
        RECT  -0.8675 8.415 -0.8025 8.875 ;
        RECT  -0.8675 8.8075 -0.8025 8.9425 ;
        RECT  -1.7625 9.4225 -1.6975 9.4875 ;
        RECT  -1.73 9.4225 -1.4125 9.4875 ;
        RECT  -1.7625 9.165 -1.6975 9.455 ;
        RECT  -1.7625 9.0325 -1.6975 9.0975 ;
        RECT  -1.73 9.0325 -1.4125 9.0975 ;
        RECT  -1.7625 9.065 -1.6975 9.165 ;
        RECT  -1.7625 8.6525 -1.6975 8.7175 ;
        RECT  -1.73 8.6525 -1.4125 8.7175 ;
        RECT  -1.7625 8.685 -1.6975 9.165 ;
        RECT  -0.3825 16.185 -0.3175 16.935 ;
        RECT  -1.7275 16.185 -1.6625 16.935 ;
        RECT  -1.695 16.8025 -1.4125 16.8675 ;
        RECT  -0.53 16.8025 -0.35 16.8675 ;
        RECT  -1.695 16.2525 -1.4125 16.3175 ;
        RECT  -1.695 16.6325 -1.4125 16.6975 ;
        RECT  -0.6325 16.2525 -0.35 16.3175 ;
        RECT  -1.325 16.185 -1.26 16.22 ;
        RECT  -0.795 16.185 -0.73 16.46 ;
        RECT  -1.0125 16.6975 -0.9475 16.935 ;
        RECT  -0.7675 16.2525 -0.6325 16.3175 ;
        RECT  -0.7675 16.4425 -0.6325 16.5075 ;
        RECT  -0.7675 16.4425 -0.6325 16.5075 ;
        RECT  -0.7675 16.6325 -0.6325 16.6975 ;
        RECT  -1.5475 16.2525 -1.4125 16.3175 ;
        RECT  -1.5475 16.4425 -1.4125 16.5075 ;
        RECT  -1.5475 16.4425 -1.4125 16.5075 ;
        RECT  -1.5475 16.6325 -1.4125 16.6975 ;
        RECT  -1.5475 16.8025 -1.4125 16.8675 ;
        RECT  -0.6325 16.8025 -0.4975 16.8675 ;
        RECT  -1.31 16.665 -1.245 16.73 ;
        RECT  -1.31 16.4425 -1.245 16.5075 ;
        RECT  -1.2775 16.665 -0.4975 16.73 ;
        RECT  -1.31 16.475 -1.245 16.6975 ;
        RECT  -1.4125 16.4425 -1.2775 16.5075 ;
        RECT  -1.325 16.22 -1.26 16.355 ;
        RECT  -0.795 16.46 -0.73 16.595 ;
        RECT  -1.9775 21.245 -1.9075 21.38 ;
        RECT  -2.135 21.1325 -2.07 21.1975 ;
        RECT  -4.1925 22.5675 -3.96 22.6325 ;
        RECT  -4.9025 26.2325 -0.3825 26.2975 ;
        RECT  -0.415 24.07 -0.35 25.19 ;
        RECT  -3.105 24.07 -3.04 25.19 ;
        RECT  -1.9075 20.6625 -1.3475 20.7275 ;
        RECT  -1.9075 19.3175 -1.3475 19.3825 ;
        RECT  -1.84 19.3825 -1.775 19.7475 ;
        RECT  -1.84 20.5275 -1.775 20.6625 ;
        RECT  -1.48 20.5925 -1.415 20.6625 ;
        RECT  -1.48 19.3825 -1.415 19.4725 ;
        RECT  -1.67 19.6125 -1.605 20.56 ;
        RECT  -1.3825 20.08 -1.3475 20.145 ;
        RECT  -1.9075 20.08 -1.67 20.145 ;
        RECT  -1.48 20.3225 -1.415 20.4575 ;
        RECT  -1.67 20.3225 -1.605 20.4575 ;
        RECT  -1.48 19.4725 -1.415 19.7475 ;
        RECT  -1.67 19.4725 -1.605 19.7475 ;
        RECT  -1.84 19.4725 -1.775 19.7475 ;
        RECT  -1.84 20.4575 -1.775 20.5925 ;
        RECT  -1.5175 20.08 -1.3825 20.145 ;
        RECT  -0.94 21.235 -0.805 21.3 ;
        RECT  -0.94 21.045 -0.805 21.11 ;
        RECT  -1.0 23.795 -0.935 23.93 ;
        RECT  -0.415 23.37 -0.35 23.93 ;
        RECT  -1.76 23.37 -1.695 23.93 ;
        RECT  -1.695 23.4375 -1.33 23.5025 ;
        RECT  -0.55 23.4375 -0.415 23.5025 ;
        RECT  -0.485 23.7975 -0.415 23.8625 ;
        RECT  -1.695 23.7975 -1.605 23.8625 ;
        RECT  -1.465 23.6075 -0.5175 23.6725 ;
        RECT  -0.9975 23.895 -0.9325 23.93 ;
        RECT  -0.685 23.7975 -0.55 23.8625 ;
        RECT  -0.685 23.6075 -0.55 23.6725 ;
        RECT  -1.225 23.7975 -0.95 23.8625 ;
        RECT  -1.225 23.6075 -0.95 23.6725 ;
        RECT  -1.33 23.4375 -1.055 23.5025 ;
        RECT  -0.485 23.4375 -0.35 23.5025 ;
        RECT  -0.9225 23.76 -0.8575 23.895 ;
        RECT  -1.0 23.235 -0.935 23.37 ;
        RECT  -0.415 22.81 -0.35 23.37 ;
        RECT  -1.76 22.81 -1.695 23.37 ;
        RECT  -1.695 22.8775 -1.33 22.9425 ;
        RECT  -0.55 22.8775 -0.415 22.9425 ;
        RECT  -0.485 23.2375 -0.415 23.3025 ;
        RECT  -1.695 23.2375 -1.605 23.3025 ;
        RECT  -1.465 23.0475 -0.5175 23.1125 ;
        RECT  -0.9975 23.335 -0.9325 23.37 ;
        RECT  -0.685 23.2375 -0.55 23.3025 ;
        RECT  -0.685 23.0475 -0.55 23.1125 ;
        RECT  -1.225 23.2375 -0.95 23.3025 ;
        RECT  -1.225 23.0475 -0.95 23.1125 ;
        RECT  -1.33 22.8775 -1.055 22.9425 ;
        RECT  -0.485 22.8775 -0.35 22.9425 ;
        RECT  -0.9225 23.2 -0.8575 23.335 ;
        RECT  -2.52 22.81 -2.455 22.945 ;
        RECT  -3.105 22.81 -3.04 23.37 ;
        RECT  -1.76 22.81 -1.695 23.37 ;
        RECT  -2.125 23.2375 -1.76 23.3025 ;
        RECT  -3.04 23.2375 -2.905 23.3025 ;
        RECT  -3.04 22.8775 -2.97 22.9425 ;
        RECT  -1.85 22.8775 -1.76 22.9425 ;
        RECT  -2.9375 23.0675 -1.99 23.1325 ;
        RECT  -2.5225 22.81 -2.4575 22.845 ;
        RECT  -2.905 22.8775 -2.77 22.9425 ;
        RECT  -2.905 23.0675 -2.77 23.1325 ;
        RECT  -2.505 22.8775 -2.23 22.9425 ;
        RECT  -2.505 23.0675 -2.23 23.1325 ;
        RECT  -2.4 23.2375 -2.125 23.3025 ;
        RECT  -3.105 23.2375 -2.97 23.3025 ;
        RECT  -2.5975 22.845 -2.5325 22.98 ;
        RECT  -2.52 23.37 -2.455 23.505 ;
        RECT  -3.105 23.37 -3.04 23.93 ;
        RECT  -1.76 23.37 -1.695 23.93 ;
        RECT  -2.125 23.7975 -1.76 23.8625 ;
        RECT  -3.04 23.7975 -2.905 23.8625 ;
        RECT  -3.04 23.4375 -2.97 23.5025 ;
        RECT  -1.85 23.4375 -1.76 23.5025 ;
        RECT  -2.9375 23.6275 -1.99 23.6925 ;
        RECT  -2.5225 23.37 -2.4575 23.405 ;
        RECT  -2.905 23.4375 -2.77 23.5025 ;
        RECT  -2.905 23.6275 -2.77 23.6925 ;
        RECT  -2.505 23.4375 -2.23 23.5025 ;
        RECT  -2.505 23.6275 -2.23 23.6925 ;
        RECT  -2.4 23.7975 -2.125 23.8625 ;
        RECT  -3.105 23.7975 -2.97 23.8625 ;
        RECT  -2.5975 23.405 -2.5325 23.54 ;
        RECT  -1.0 23.4725 -0.935 23.6075 ;
        RECT  -1.0 22.9125 -0.935 23.0475 ;
        RECT  -2.52 23.1325 -2.455 23.2675 ;
        RECT  -4.8475 22.9975 -4.7825 23.1325 ;
        RECT  -4.6625 22.9975 -4.5975 23.1325 ;
        RECT  -4.4925 23.0025 -4.4275 23.1375 ;
        RECT  -4.3075 23.0025 -4.2425 23.1375 ;
        RECT  -4.9275 23.3875 -4.8625 23.5225 ;
        RECT  -4.7425 23.3875 -4.6775 23.5225 ;
        RECT  -4.4125 23.3875 -4.3475 23.5225 ;
        RECT  -4.2275 23.3875 -4.1625 23.5225 ;
        RECT  -4.9275 23.8525 -4.8625 23.9875 ;
        RECT  -4.7425 23.8525 -4.6775 23.9875 ;
        RECT  -4.4125 23.8525 -4.3475 23.9875 ;
        RECT  -4.2275 23.8525 -4.1625 23.9875 ;
        RECT  -4.225 23.0025 -4.16 23.1375 ;
        RECT  -4.93 23.4775 -4.865 23.6125 ;
        RECT  -4.225 23.4775 -4.16 23.6125 ;
        RECT  -4.6775 22.9975 -4.6125 23.1325 ;
        RECT  -4.4775 23.0025 -4.4125 23.1375 ;
        RECT  -4.725 23.5925 -4.59 23.6575 ;
        RECT  -4.5 23.7425 -4.365 23.8075 ;
        RECT  -4.6025 22.8475 -4.4675 22.9125 ;
        RECT  -4.61 24.0525 -4.475 24.1175 ;
        RECT  -4.6075 22.7075 -4.4725 22.7725 ;
        RECT  -4.965 22.7075 -4.83 22.7725 ;
        RECT  -4.245 23.0025 -4.1925 23.1375 ;
        RECT  -4.26 22.7075 -4.125 22.7725 ;
        RECT  -4.575 24.0525 -4.51 24.1175 ;
        RECT  -4.2275 22.8475 -4.1575 22.9125 ;
        RECT  -4.7825 23.2225 -4.6775 23.2875 ;
        RECT  -4.7425 23.2875 -4.6775 23.3875 ;
        RECT  -4.8475 23.1325 -4.7825 23.2875 ;
        RECT  -4.4125 23.2225 -4.3075 23.2875 ;
        RECT  -4.4125 23.2875 -4.3475 23.3875 ;
        RECT  -4.3075 23.1375 -4.2425 23.2875 ;
        RECT  -4.9275 23.9875 -4.8625 24.0525 ;
        RECT  -4.2275 23.9875 -4.1625 24.0525 ;
        RECT  -4.7425 23.3875 -4.6775 23.8775 ;
        RECT  -4.4125 23.3875 -4.3475 23.8775 ;
        RECT  -4.9875 22.8475 -4.1025 22.9125 ;
        RECT  -4.9875 24.0525 -4.1025 24.1175 ;
        RECT  -4.9875 22.7075 -4.1025 22.7725 ;
        RECT  -4.9275 21.4925 -4.8625 21.6275 ;
        RECT  -4.7425 21.4925 -4.6775 21.6275 ;
        RECT  -4.2275 21.4925 -4.1625 21.6275 ;
        RECT  -4.4125 21.4925 -4.3475 21.6275 ;
        RECT  -4.7425 21.9575 -4.6775 22.0925 ;
        RECT  -4.9275 21.9575 -4.8625 22.0925 ;
        RECT  -4.4125 21.9575 -4.3475 22.0925 ;
        RECT  -4.2275 21.9575 -4.1625 22.0925 ;
        RECT  -4.8475 22.3475 -4.7825 22.4825 ;
        RECT  -4.6625 22.3475 -4.5975 22.4825 ;
        RECT  -4.4925 22.3475 -4.4275 22.4825 ;
        RECT  -4.3075 22.3475 -4.2425 22.4825 ;
        RECT  -4.93 21.855 -4.865 21.99 ;
        RECT  -4.93 21.855 -4.865 21.99 ;
        RECT  -4.93 21.855 -4.865 21.99 ;
        RECT  -4.93 21.855 -4.865 21.99 ;
        RECT  -4.93 21.855 -4.865 21.99 ;
        RECT  -4.93 21.855 -4.865 21.99 ;
        RECT  -4.6075 21.3625 -4.4725 21.4275 ;
        RECT  -4.26 22.7075 -4.125 22.7725 ;
        RECT  -4.965 22.7075 -4.83 22.7725 ;
        RECT  -4.595 22.5675 -4.46 22.6325 ;
        RECT  -4.93 21.855 -4.865 21.99 ;
        RECT  -4.93 21.855 -4.865 21.99 ;
        RECT  -4.93 21.855 -4.865 21.99 ;
        RECT  -4.93 21.855 -4.865 21.99 ;
        RECT  -4.5 21.6775 -4.365 21.7425 ;
        RECT  -4.5 21.6775 -4.365 21.7425 ;
        RECT  -4.725 21.8275 -4.59 21.8925 ;
        RECT  -4.725 21.8275 -4.59 21.8925 ;
        RECT  -4.93 21.855 -4.865 21.99 ;
        RECT  -4.93 21.855 -4.865 21.99 ;
        RECT  -4.93 21.855 -4.865 21.99 ;
        RECT  -4.93 21.855 -4.865 21.99 ;
        RECT  -4.48 22.3475 -4.415 22.4825 ;
        RECT  -4.225 21.855 -4.16 21.99 ;
        RECT  -4.225 21.855 -4.16 21.99 ;
        RECT  -4.225 21.855 -4.16 21.99 ;
        RECT  -4.225 21.855 -4.16 21.99 ;
        RECT  -4.225 21.855 -4.16 21.99 ;
        RECT  -4.225 21.855 -4.16 21.99 ;
        RECT  -4.93 21.855 -4.865 21.99 ;
        RECT  -4.93 21.855 -4.865 21.99 ;
        RECT  -4.93 21.855 -4.865 21.99 ;
        RECT  -4.93 21.855 -4.865 21.99 ;
        RECT  -4.675 22.3475 -4.61 22.4825 ;
        RECT  -4.6125 22.7075 -4.4775 22.7725 ;
        RECT  -4.6125 22.7075 -4.4775 22.7725 ;
        RECT  -4.965 22.7075 -4.83 22.7725 ;
        RECT  -4.6075 21.3625 -4.4725 21.4275 ;
        RECT  -4.965 22.7075 -4.83 22.7725 ;
        RECT  -4.965 22.7075 -4.83 22.7725 ;
        RECT  -4.93 21.855 -4.865 21.99 ;
        RECT  -4.93 21.855 -4.865 21.99 ;
        RECT  -4.93 21.855 -4.865 21.99 ;
        RECT  -4.93 21.855 -4.865 21.99 ;
        RECT  -4.93 21.855 -4.865 21.99 ;
        RECT  -4.93 21.855 -4.865 21.99 ;
        RECT  -4.26 22.7075 -4.125 22.7725 ;
        RECT  -4.585 21.365 -4.485 21.4275 ;
        RECT  -4.585 21.3625 -4.485 21.425 ;
        RECT  -4.865 22.5675 -4.8125 22.63 ;
        RECT  -4.585 21.365 -4.485 21.4275 ;
        RECT  -4.9325 21.4275 -4.8625 21.6275 ;
        RECT  -4.9325 21.9575 -4.8625 22.0925 ;
        RECT  -4.9325 21.9575 -4.8625 22.0925 ;
        RECT  -4.9875 22.7075 -4.1025 22.7725 ;
        RECT  -4.8525 22.1925 -4.6775 22.2575 ;
        RECT  -4.2275 21.9575 -4.1575 22.0925 ;
        RECT  -4.4125 21.5175 -4.3475 22.2575 ;
        RECT  -4.585 21.3625 -4.485 21.425 ;
        RECT  -4.16 22.5675 -4.1075 22.63 ;
        RECT  -4.9325 21.9575 -4.8625 22.0925 ;
        RECT  -4.9875 21.3625 -4.1025 21.4275 ;
        RECT  -4.7425 21.6275 -4.6775 22.2575 ;
        RECT  -4.9325 21.9575 -4.8625 22.0925 ;
        RECT  -4.9325 21.9575 -4.8625 22.0925 ;
        RECT  -4.3125 22.1925 -4.2425 22.4825 ;
        RECT  -4.2275 21.9575 -4.1575 22.0925 ;
        RECT  -4.9875 22.5675 -4.1025 22.6325 ;
        RECT  -4.9325 21.9575 -4.8625 22.0925 ;
        RECT  -4.9325 21.4275 -4.8625 21.6275 ;
        RECT  -4.2275 21.4275 -4.1575 21.6275 ;
        RECT  -4.8525 22.1925 -4.7825 22.4825 ;
        RECT  -4.4125 22.1925 -4.2425 22.2575 ;
        RECT  -4.9275 21.1625 -4.8625 21.2975 ;
        RECT  -4.7425 21.1625 -4.6775 21.2975 ;
        RECT  -4.2275 21.1625 -4.1625 21.2975 ;
        RECT  -4.4125 21.1625 -4.3475 21.2975 ;
        RECT  -4.7425 20.6975 -4.6775 20.8325 ;
        RECT  -4.9275 20.6975 -4.8625 20.8325 ;
        RECT  -4.4125 20.6975 -4.3475 20.8325 ;
        RECT  -4.2275 20.6975 -4.1625 20.8325 ;
        RECT  -4.8475 20.3075 -4.7825 20.4425 ;
        RECT  -4.6625 20.3075 -4.5975 20.4425 ;
        RECT  -4.4925 20.3075 -4.4275 20.4425 ;
        RECT  -4.3075 20.3075 -4.2425 20.4425 ;
        RECT  -4.93 20.8 -4.865 20.935 ;
        RECT  -4.93 20.8 -4.865 20.935 ;
        RECT  -4.93 20.8 -4.865 20.935 ;
        RECT  -4.93 20.8 -4.865 20.935 ;
        RECT  -4.93 20.8 -4.865 20.935 ;
        RECT  -4.93 20.8 -4.865 20.935 ;
        RECT  -4.6075 21.3625 -4.4725 21.4275 ;
        RECT  -4.26 20.0175 -4.125 20.0825 ;
        RECT  -4.965 20.0175 -4.83 20.0825 ;
        RECT  -4.595 20.1575 -4.46 20.2225 ;
        RECT  -4.93 20.8 -4.865 20.935 ;
        RECT  -4.93 20.8 -4.865 20.935 ;
        RECT  -4.93 20.8 -4.865 20.935 ;
        RECT  -4.93 20.8 -4.865 20.935 ;
        RECT  -4.5 21.0475 -4.365 21.1125 ;
        RECT  -4.5 21.0475 -4.365 21.1125 ;
        RECT  -4.725 20.8975 -4.59 20.9625 ;
        RECT  -4.725 20.8975 -4.59 20.9625 ;
        RECT  -4.93 20.8 -4.865 20.935 ;
        RECT  -4.93 20.8 -4.865 20.935 ;
        RECT  -4.93 20.8 -4.865 20.935 ;
        RECT  -4.93 20.8 -4.865 20.935 ;
        RECT  -4.48 20.3075 -4.415 20.4425 ;
        RECT  -4.225 20.8 -4.16 20.935 ;
        RECT  -4.225 20.8 -4.16 20.935 ;
        RECT  -4.225 20.8 -4.16 20.935 ;
        RECT  -4.225 20.8 -4.16 20.935 ;
        RECT  -4.225 20.8 -4.16 20.935 ;
        RECT  -4.225 20.8 -4.16 20.935 ;
        RECT  -4.93 20.8 -4.865 20.935 ;
        RECT  -4.93 20.8 -4.865 20.935 ;
        RECT  -4.93 20.8 -4.865 20.935 ;
        RECT  -4.93 20.8 -4.865 20.935 ;
        RECT  -4.675 20.3075 -4.61 20.4425 ;
        RECT  -4.6125 20.0175 -4.4775 20.0825 ;
        RECT  -4.6125 20.0175 -4.4775 20.0825 ;
        RECT  -4.965 20.0175 -4.83 20.0825 ;
        RECT  -4.6075 21.3625 -4.4725 21.4275 ;
        RECT  -4.965 20.0175 -4.83 20.0825 ;
        RECT  -4.965 20.0175 -4.83 20.0825 ;
        RECT  -4.93 20.8 -4.865 20.935 ;
        RECT  -4.93 20.8 -4.865 20.935 ;
        RECT  -4.93 20.8 -4.865 20.935 ;
        RECT  -4.93 20.8 -4.865 20.935 ;
        RECT  -4.93 20.8 -4.865 20.935 ;
        RECT  -4.93 20.8 -4.865 20.935 ;
        RECT  -4.26 20.0175 -4.125 20.0825 ;
        RECT  -4.585 21.3625 -4.485 21.425 ;
        RECT  -4.585 21.365 -4.485 21.4275 ;
        RECT  -4.865 20.16 -4.8125 20.2225 ;
        RECT  -4.585 21.3625 -4.485 21.425 ;
        RECT  -4.9325 21.1625 -4.8625 21.3625 ;
        RECT  -4.9325 20.6975 -4.8625 20.8325 ;
        RECT  -4.9325 20.6975 -4.8625 20.8325 ;
        RECT  -4.9875 20.0175 -4.1025 20.0825 ;
        RECT  -4.8525 20.5325 -4.6775 20.5975 ;
        RECT  -4.2275 20.6975 -4.1575 20.8325 ;
        RECT  -4.4125 20.5325 -4.3475 21.2725 ;
        RECT  -4.585 21.365 -4.485 21.4275 ;
        RECT  -4.16 20.16 -4.1075 20.2225 ;
        RECT  -4.9325 20.6975 -4.8625 20.8325 ;
        RECT  -4.9875 21.3625 -4.1025 21.4275 ;
        RECT  -4.7425 20.5325 -4.6775 21.1625 ;
        RECT  -4.9325 20.6975 -4.8625 20.8325 ;
        RECT  -4.9325 20.6975 -4.8625 20.8325 ;
        RECT  -4.3125 20.3075 -4.2425 20.5975 ;
        RECT  -4.2275 20.6975 -4.1575 20.8325 ;
        RECT  -4.9875 20.1575 -4.1025 20.2225 ;
        RECT  -4.9325 20.6975 -4.8625 20.8325 ;
        RECT  -4.9325 21.1625 -4.8625 21.3625 ;
        RECT  -4.2275 21.1625 -4.1575 21.3625 ;
        RECT  -4.8525 20.3075 -4.7825 20.5975 ;
        RECT  -4.4125 20.5325 -4.2425 20.5975 ;
        RECT  -1.975 21.1425 -1.91 21.2775 ;
        RECT  -0.9975 23.7575 -0.9325 23.8225 ;
        RECT  -0.965 23.7575 -0.3825 23.8225 ;
        RECT  -0.9975 23.65 -0.9325 23.79 ;
        RECT  -1.38 21.3825 -1.315 21.4525 ;
        RECT  -2.135 21.3825 -2.07 21.4525 ;
        RECT  -1.38 21.2775 -1.315 21.4175 ;
        RECT  -2.135 21.39 -2.07 21.4175 ;
        RECT  -1.415 21.385 -1.28 21.45 ;
        RECT  -2.17 21.385 -2.035 21.45 ;
        RECT  -4.4125 24.28 -4.3425 24.345 ;
        RECT  -4.3775 24.2825 -2.1025 24.3475 ;
        RECT  -4.445 24.28 -4.31 24.345 ;
        RECT  -0.6525 21.36 -0.5875 21.495 ;
        RECT  -0.65 19.52 -0.58 19.585 ;
        RECT  -2.5575 19.5225 -2.4875 19.5875 ;
        RECT  -2.5225 19.5225 -0.615 19.5875 ;
        RECT  -0.6825 19.52 -0.5475 19.585 ;
        RECT  -2.59 19.5225 -2.455 19.5875 ;
        RECT  -2.59 24.1675 -2.525 24.3025 ;
        RECT  -0.6475 21.33 -0.5825 21.465 ;
        RECT  -4.025 22.3975 -3.96 22.5325 ;
        RECT  -0.94 21.2425 -0.875 21.3075 ;
        RECT  -0.94 21.275 -0.875 21.6575 ;
        RECT  -1.3475 21.2425 -0.9075 21.3075 ;
        RECT  -3.7375 22.0075 -3.6675 22.0725 ;
        RECT  -3.7025 22.0075 -1.3475 22.0725 ;
        RECT  -3.77 22.0075 -3.635 22.0725 ;
        RECT  -0.94 21.625 -0.875 21.69 ;
        RECT  -0.94 21.4675 -0.875 21.6575 ;
        RECT  -1.3475 21.625 -0.9075 21.69 ;
        RECT  -1.76 24.0275 -1.695 24.0925 ;
        RECT  -1.76 23.93 -1.695 24.06 ;
        RECT  -3.7025 24.0275 -1.7275 24.0925 ;
        RECT  -3.7375 23.7675 -3.6675 23.8325 ;
        RECT  -3.7025 23.7675 -1.7275 23.8325 ;
        RECT  -3.77 23.7675 -3.635 23.8325 ;
        RECT  -0.4175 20.6625 -0.3475 20.7275 ;
        RECT  -0.4175 16.165 -0.3475 16.23 ;
        RECT  -3.1075 16.1675 -3.0375 16.2325 ;
        RECT  -1.3475 20.6625 -0.3825 20.7275 ;
        RECT  -3.0725 16.1675 -0.3825 16.2325 ;
        RECT  -0.45 20.6625 -0.315 20.7275 ;
        RECT  -0.45 16.165 -0.315 16.23 ;
        RECT  -3.14 16.1675 -3.005 16.2325 ;
        RECT  -3.77 26.2325 -3.705 26.3675 ;
        RECT  -3.5275 23.93 -3.4575 23.995 ;
        RECT  -3.5275 25.01 -3.4575 25.075 ;
        RECT  -3.4925 23.93 -3.04 23.995 ;
        RECT  -4.1925 25.0125 -3.4925 25.0775 ;
        RECT  -3.56 23.93 -3.425 23.995 ;
        RECT  -3.56 25.01 -3.425 25.075 ;
        RECT  -3.7375 28.345 -3.6675 28.41 ;
        RECT  -4.1925 28.3475 -3.7025 28.4125 ;
        RECT  -3.77 28.345 -3.635 28.41 ;
        RECT  -3.5275 23.93 -3.4575 23.995 ;
        RECT  -3.5275 22.6 -3.4575 22.665 ;
        RECT  -3.4925 23.93 -3.04 23.995 ;
        RECT  -4.1925 22.6025 -3.4925 22.6675 ;
        RECT  -3.56 23.93 -3.425 23.995 ;
        RECT  -3.56 22.6 -3.425 22.665 ;
        RECT  -3.7375 31.035 -3.6675 31.1 ;
        RECT  -4.545 31.0375 -3.7025 31.1025 ;
        RECT  -3.77 31.035 -3.635 31.1 ;
        RECT  -4.9325 20.6625 -4.8625 20.7275 ;
        RECT  -4.8975 20.6625 -0.7875 20.7275 ;
        RECT  -4.965 20.6625 -4.83 20.7275 ;
        RECT  -4.2275 20.6625 -4.1575 20.7275 ;
        RECT  -4.1925 20.6625 -0.7875 20.7275 ;
        RECT  -4.26 20.6625 -4.125 20.7275 ;
        RECT  -0.3825 17.335 -0.3175 17.895 ;
        RECT  -1.7275 17.335 -1.6625 17.895 ;
        RECT  -1.6625 17.4025 -1.2975 17.4675 ;
        RECT  -0.5175 17.4025 -0.3825 17.4675 ;
        RECT  -0.4525 17.7625 -0.3825 17.8275 ;
        RECT  -1.6625 17.7625 -1.5725 17.8275 ;
        RECT  -1.4325 17.5725 -0.485 17.6375 ;
        RECT  -0.965 17.86 -0.9 17.895 ;
        RECT  -0.965 17.335 -0.9 17.5725 ;
        RECT  -0.6525 17.7625 -0.5175 17.8275 ;
        RECT  -0.6525 17.5725 -0.5175 17.6375 ;
        RECT  -1.1925 17.7625 -0.9175 17.8275 ;
        RECT  -1.1925 17.5725 -0.9175 17.6375 ;
        RECT  -1.2975 17.4025 -1.0225 17.4675 ;
        RECT  -0.4525 17.4025 -0.3175 17.4675 ;
        RECT  -0.89 17.725 -0.825 17.86 ;
        RECT  -0.3825 17.895 -0.3175 18.455 ;
        RECT  -1.7275 17.895 -1.6625 18.455 ;
        RECT  -1.6625 17.9625 -1.2975 18.0275 ;
        RECT  -0.5175 17.9625 -0.3825 18.0275 ;
        RECT  -0.4525 18.3225 -0.3825 18.3875 ;
        RECT  -1.6625 18.3225 -1.5725 18.3875 ;
        RECT  -1.4325 18.1325 -0.485 18.1975 ;
        RECT  -0.965 18.42 -0.9 18.455 ;
        RECT  -0.965 17.895 -0.9 18.1325 ;
        RECT  -0.6525 18.3225 -0.5175 18.3875 ;
        RECT  -0.6525 18.1325 -0.5175 18.1975 ;
        RECT  -1.1925 18.3225 -0.9175 18.3875 ;
        RECT  -1.1925 18.1325 -0.9175 18.1975 ;
        RECT  -1.2975 17.9625 -1.0225 18.0275 ;
        RECT  -0.4525 17.9625 -0.3175 18.0275 ;
        RECT  -0.89 18.285 -0.825 18.42 ;
        RECT  -3.0725 16.185 -3.0075 17.335 ;
        RECT  -1.7275 16.185 -1.6625 17.335 ;
        RECT  -2.91 17.02 -1.825 17.085 ;
        RECT  -1.9775 17.1575 -1.695 17.2225 ;
        RECT  -3.04 17.1575 -2.77 17.2225 ;
        RECT  -1.9775 16.4175 -1.695 16.4825 ;
        RECT  -1.9775 16.7975 -1.695 16.8625 ;
        RECT  -3.04 16.4175 -2.7575 16.4825 ;
        RECT  -2.12 16.185 -2.055 16.495 ;
        RECT  -2.6425 16.185 -2.5775 16.35 ;
        RECT  -2.7825 16.185 -2.7175 16.35 ;
        RECT  -2.3875 17.02 -2.3225 17.335 ;
        RECT  -2.8125 16.4175 -2.5375 16.4825 ;
        RECT  -2.8125 16.6075 -2.5375 16.6725 ;
        RECT  -2.8125 16.6075 -2.5375 16.6725 ;
        RECT  -2.8125 16.7975 -2.5375 16.8625 ;
        RECT  -2.8125 16.7975 -2.5375 16.8625 ;
        RECT  -2.8125 16.9875 -2.5375 17.0525 ;
        RECT  -2.2675 16.4175 -2.1325 16.4825 ;
        RECT  -2.2675 16.6075 -2.1325 16.6725 ;
        RECT  -2.2675 16.6075 -2.1325 16.6725 ;
        RECT  -2.2675 16.7975 -2.1325 16.8625 ;
        RECT  -2.2675 16.7975 -2.1325 16.8625 ;
        RECT  -2.2675 16.9875 -2.1325 17.0525 ;
        RECT  -2.1125 17.1575 -1.9775 17.2225 ;
        RECT  -3.1925 17.1575 -2.9175 17.2225 ;
        RECT  -2.1125 16.6075 -1.9775 16.6725 ;
        RECT  -2.1125 16.9875 -1.9775 17.0525 ;
        RECT  -2.2 16.36 -2.135 16.495 ;
        RECT  -2.7125 16.665 -2.5775 16.73 ;
        RECT  -2.7125 16.6625 -2.5775 16.7275 ;
        RECT  -2.715 16.215 -2.65 16.35 ;
        RECT  -2.7125 16.855 -2.5775 16.92 ;
        RECT  -2.7125 16.8525 -2.5775 16.9175 ;
        RECT  -2.855 16.215 -2.79 16.35 ;
        RECT  -3.0725 16.185 -3.0075 17.335 ;
        RECT  -4.4175 16.185 -4.3525 17.335 ;
        RECT  -4.255 17.02 -3.17 17.085 ;
        RECT  -4.385 17.1575 -4.1025 17.2225 ;
        RECT  -3.31 17.1575 -3.04 17.2225 ;
        RECT  -4.385 16.4175 -4.1025 16.4825 ;
        RECT  -4.385 16.7975 -4.1025 16.8625 ;
        RECT  -3.3225 16.4175 -3.04 16.4825 ;
        RECT  -4.025 16.185 -3.96 16.495 ;
        RECT  -3.5025 16.185 -3.4375 16.35 ;
        RECT  -3.3625 16.185 -3.2975 16.35 ;
        RECT  -3.7575 17.02 -3.6925 17.335 ;
        RECT  -3.7125 16.4175 -3.4375 16.4825 ;
        RECT  -3.7125 16.6075 -3.4375 16.6725 ;
        RECT  -3.7125 16.6075 -3.4375 16.6725 ;
        RECT  -3.7125 16.7975 -3.4375 16.8625 ;
        RECT  -3.7125 16.7975 -3.4375 16.8625 ;
        RECT  -3.7125 16.9875 -3.4375 17.0525 ;
        RECT  -4.2375 16.4175 -4.1025 16.4825 ;
        RECT  -4.2375 16.6075 -4.1025 16.6725 ;
        RECT  -4.2375 16.6075 -4.1025 16.6725 ;
        RECT  -4.2375 16.7975 -4.1025 16.8625 ;
        RECT  -4.2375 16.7975 -4.1025 16.8625 ;
        RECT  -4.2375 16.9875 -4.1025 17.0525 ;
        RECT  -4.2375 17.1575 -4.1025 17.2225 ;
        RECT  -3.4375 17.1575 -3.1625 17.2225 ;
        RECT  -4.2375 16.6075 -4.1025 16.6725 ;
        RECT  -4.2375 16.9875 -4.1025 17.0525 ;
        RECT  -4.02 16.36 -3.955 16.495 ;
        RECT  -3.6375 16.665 -3.5025 16.73 ;
        RECT  -3.6375 16.6625 -3.5025 16.7275 ;
        RECT  -3.5 16.215 -3.435 16.35 ;
        RECT  -3.6375 16.855 -3.5025 16.92 ;
        RECT  -3.6375 16.8525 -3.5025 16.9175 ;
        RECT  -3.36 16.215 -3.295 16.35 ;
        RECT  -3.0725 17.335 -3.0075 17.895 ;
        RECT  -1.7275 17.335 -1.6625 17.895 ;
        RECT  -2.0925 17.7625 -1.7275 17.8275 ;
        RECT  -3.0075 17.7625 -2.8725 17.8275 ;
        RECT  -3.0075 17.4025 -2.9375 17.4675 ;
        RECT  -1.8175 17.4025 -1.7275 17.4675 ;
        RECT  -2.905 17.5925 -1.9575 17.6575 ;
        RECT  -2.49 17.335 -2.425 17.37 ;
        RECT  -2.49 17.6575 -2.425 17.895 ;
        RECT  -2.8725 17.4025 -2.7375 17.4675 ;
        RECT  -2.8725 17.5925 -2.7375 17.6575 ;
        RECT  -2.4725 17.4025 -2.1975 17.4675 ;
        RECT  -2.4725 17.5925 -2.1975 17.6575 ;
        RECT  -2.3675 17.7625 -2.0925 17.8275 ;
        RECT  -3.0725 17.7625 -2.9375 17.8275 ;
        RECT  -2.565 17.37 -2.5 17.505 ;
        RECT  -3.0725 17.335 -3.0075 17.895 ;
        RECT  -4.4175 17.335 -4.3525 17.895 ;
        RECT  -4.3525 17.7625 -3.9875 17.8275 ;
        RECT  -3.2075 17.7625 -3.0725 17.8275 ;
        RECT  -3.1425 17.4025 -3.0725 17.4675 ;
        RECT  -4.3525 17.4025 -4.2625 17.4675 ;
        RECT  -4.1225 17.5925 -3.175 17.6575 ;
        RECT  -3.655 17.335 -3.59 17.37 ;
        RECT  -3.655 17.6575 -3.59 17.895 ;
        RECT  -3.4125 17.4025 -3.2775 17.4675 ;
        RECT  -3.4125 17.5925 -3.2775 17.6575 ;
        RECT  -4.2625 17.4025 -3.9875 17.4675 ;
        RECT  -4.2625 17.5925 -3.9875 17.6575 ;
        RECT  -4.2625 17.7625 -3.9875 17.8275 ;
        RECT  -3.2775 17.7625 -3.1425 17.8275 ;
        RECT  -3.655 17.37 -3.59 17.505 ;
        RECT  -3.0725 17.895 -3.0075 18.455 ;
        RECT  -4.4175 17.895 -4.3525 18.455 ;
        RECT  -4.3525 18.3225 -3.9875 18.3875 ;
        RECT  -3.2075 18.3225 -3.0725 18.3875 ;
        RECT  -3.1425 17.9625 -3.0725 18.0275 ;
        RECT  -4.3525 17.9625 -4.2625 18.0275 ;
        RECT  -4.1225 18.1525 -3.175 18.2175 ;
        RECT  -3.655 17.895 -3.59 17.93 ;
        RECT  -3.655 18.2175 -3.59 18.455 ;
        RECT  -3.4125 17.9625 -3.2775 18.0275 ;
        RECT  -3.4125 18.1525 -3.2775 18.2175 ;
        RECT  -4.2625 17.9625 -3.9875 18.0275 ;
        RECT  -4.2625 18.1525 -3.9875 18.2175 ;
        RECT  -4.2625 18.3225 -3.9875 18.3875 ;
        RECT  -3.2775 18.3225 -3.1425 18.3875 ;
        RECT  -3.655 17.93 -3.59 18.065 ;
        RECT  -3.0725 18.455 -3.0075 19.015 ;
        RECT  -4.4175 18.455 -4.3525 19.015 ;
        RECT  -4.3525 18.8825 -3.9875 18.9475 ;
        RECT  -3.2075 18.8825 -3.0725 18.9475 ;
        RECT  -3.1425 18.5225 -3.0725 18.5875 ;
        RECT  -4.3525 18.5225 -4.2625 18.5875 ;
        RECT  -4.1225 18.7125 -3.175 18.7775 ;
        RECT  -3.655 18.455 -3.59 18.49 ;
        RECT  -3.655 18.7775 -3.59 19.015 ;
        RECT  -3.4125 18.5225 -3.2775 18.5875 ;
        RECT  -3.4125 18.7125 -3.2775 18.7775 ;
        RECT  -4.2625 18.5225 -3.9875 18.5875 ;
        RECT  -4.2625 18.7125 -3.9875 18.7775 ;
        RECT  -4.2625 18.8825 -3.9875 18.9475 ;
        RECT  -3.2775 18.8825 -3.1425 18.9475 ;
        RECT  -3.655 18.49 -3.59 18.625 ;
        RECT  -3.9975 14.615 -3.9325 14.75 ;
        RECT  -3.9975 15.105 -3.9325 15.24 ;
        RECT  -4.1525 14.615 -4.0875 14.75 ;
        RECT  -4.1525 15.315 -4.0875 15.45 ;
        RECT  -5.5625 14.615 -5.4975 14.75 ;
        RECT  -5.5625 15.525 -5.4975 15.66 ;
        RECT  -4.5475 14.615 -4.4825 14.75 ;
        RECT  -4.5475 15.735 -4.4825 15.87 ;
        RECT  -1.325 15.315 -1.26 15.45 ;
        RECT  -0.795 15.945 -0.73 16.08 ;
        RECT  -2.12 15.945 -2.055 16.08 ;
        RECT  -2.6425 15.315 -2.5775 15.45 ;
        RECT  -2.7825 15.525 -2.7175 15.66 ;
        RECT  -4.025 15.945 -3.96 16.08 ;
        RECT  -3.5025 15.735 -3.4375 15.87 ;
        RECT  -3.3625 15.525 -3.2975 15.66 ;
        RECT  -0.9975 9.85 -0.9325 9.92 ;
        RECT  -0.2225 9.85 -0.1575 9.92 ;
        RECT  -0.22 15.135 -0.155 15.205 ;
        RECT  -0.9975 9.745 -0.9325 9.885 ;
        RECT  -0.22 9.885 -0.155 15.17 ;
        RECT  -0.9975 9.8175 -0.9325 9.9525 ;
        RECT  -0.2225 9.8175 -0.1575 9.9525 ;
        RECT  -0.22 15.1025 -0.155 15.2375 ;
        RECT  -0.965 14.7525 -0.9 14.8175 ;
        RECT  -0.795 14.7525 -0.73 14.8175 ;
        RECT  -0.965 14.715 -0.9 14.785 ;
        RECT  -0.9325 14.7525 -0.7625 14.8175 ;
        RECT  -0.795 14.785 -0.73 16.185 ;
        RECT  -2.49 19.405 -2.425 19.54 ;
        RECT  -3.655 19.195 -3.59 19.33 ;
        RECT  -0.965 19.615 -0.9 19.75 ;
        RECT  -0.2075 19.435 -0.1425 19.505 ;
        RECT  -0.205 19.47 -0.14 23.79 ;
        RECT  -0.2075 19.4025 -0.1425 19.5375 ;
        RECT  -1.7275 19.825 -1.6625 19.96 ;
        RECT  -4.4175 19.825 -4.3525 19.96 ;
        RECT  -0.3825 14.895 -0.3175 15.03 ;
        RECT  -0.965 13.41 -0.9 13.48 ;
        RECT  -2.0875 13.41 -2.0225 13.48 ;
        RECT  -0.965 13.445 -0.9 13.585 ;
        RECT  -2.085 8.275 -2.02 13.445 ;
        RECT  -0.965 13.3775 -0.9 13.5125 ;
        RECT  -2.0875 13.3775 -2.0225 13.5125 ;
        RECT  -0.965 13.2025 -0.9 13.2675 ;
        RECT  -0.8675 13.2025 -0.8025 13.2675 ;
        RECT  -0.965 13.235 -0.9 13.445 ;
        RECT  -0.9325 13.2025 -0.835 13.2675 ;
        RECT  -0.8675 9.745 -0.8025 13.235 ;
        RECT  -2.0825 8.275 -2.0175 8.41 ;
        RECT  -0.865 8.415 -0.8 8.55 ;
        RECT  -1.0825 16.8675 -0.9475 16.9325 ;
        RECT  -1.035 17.3375 -0.9 17.4025 ;
        RECT  0.0 19.855 0.205 19.99 ;
        Layer  via1 ; 
        RECT  11.8025 19.68 11.8675 19.745 ;
        RECT  11.8025 19.68 11.8675 19.745 ;
        RECT  11.8025 19.68 11.8675 19.745 ;
        RECT  11.8025 19.68 11.8675 19.745 ;
        RECT  11.8025 19.68 11.8675 19.745 ;
        RECT  11.8025 19.68 11.8675 19.745 ;
        RECT  11.0975 18.8625 11.1625 18.9275 ;
        RECT  11.8025 18.8625 11.8675 18.9275 ;
        RECT  11.8025 19.68 11.8675 19.745 ;
        RECT  11.8025 19.68 11.8675 19.745 ;
        RECT  11.8025 19.68 11.8675 19.745 ;
        RECT  11.8025 19.68 11.8675 19.745 ;
        RECT  11.8025 19.68 11.8675 19.745 ;
        RECT  11.8025 19.68 11.8675 19.745 ;
        RECT  11.8025 19.68 11.8675 19.745 ;
        RECT  11.8025 19.68 11.8675 19.745 ;
        RECT  11.3525 19.1875 11.4175 19.2525 ;
        RECT  11.0975 19.68 11.1625 19.745 ;
        RECT  11.0975 19.68 11.1625 19.745 ;
        RECT  11.0975 19.68 11.1625 19.745 ;
        RECT  11.0975 19.68 11.1625 19.745 ;
        RECT  11.0975 19.68 11.1625 19.745 ;
        RECT  11.0975 19.68 11.1625 19.745 ;
        RECT  11.8025 19.68 11.8675 19.745 ;
        RECT  11.8025 19.68 11.8675 19.745 ;
        RECT  11.8025 19.68 11.8675 19.745 ;
        RECT  11.8025 19.68 11.8675 19.745 ;
        RECT  11.5475 19.1875 11.6125 19.2525 ;
        RECT  11.8025 18.8625 11.8675 18.9275 ;
        RECT  11.8025 18.8625 11.8675 18.9275 ;
        RECT  11.8025 18.8625 11.8675 18.9275 ;
        RECT  11.8025 19.68 11.8675 19.745 ;
        RECT  11.8025 19.68 11.8675 19.745 ;
        RECT  11.8025 19.68 11.8675 19.745 ;
        RECT  11.8025 19.68 11.8675 19.745 ;
        RECT  11.8025 19.68 11.8675 19.745 ;
        RECT  11.8025 19.68 11.8675 19.745 ;
        RECT  11.0975 18.8625 11.1625 18.9275 ;
        RECT  11.8025 20.735 11.8675 20.8 ;
        RECT  11.8025 20.735 11.8675 20.8 ;
        RECT  11.8025 20.735 11.8675 20.8 ;
        RECT  11.8025 20.735 11.8675 20.8 ;
        RECT  11.8025 20.735 11.8675 20.8 ;
        RECT  11.8025 20.735 11.8675 20.8 ;
        RECT  11.0975 21.5525 11.1625 21.6175 ;
        RECT  11.8025 21.5525 11.8675 21.6175 ;
        RECT  11.8025 20.735 11.8675 20.8 ;
        RECT  11.8025 20.735 11.8675 20.8 ;
        RECT  11.8025 20.735 11.8675 20.8 ;
        RECT  11.8025 20.735 11.8675 20.8 ;
        RECT  11.8025 20.735 11.8675 20.8 ;
        RECT  11.8025 20.735 11.8675 20.8 ;
        RECT  11.8025 20.735 11.8675 20.8 ;
        RECT  11.8025 20.735 11.8675 20.8 ;
        RECT  11.3525 21.2275 11.4175 21.2925 ;
        RECT  11.0975 20.735 11.1625 20.8 ;
        RECT  11.0975 20.735 11.1625 20.8 ;
        RECT  11.0975 20.735 11.1625 20.8 ;
        RECT  11.0975 20.735 11.1625 20.8 ;
        RECT  11.0975 20.735 11.1625 20.8 ;
        RECT  11.0975 20.735 11.1625 20.8 ;
        RECT  11.8025 20.735 11.8675 20.8 ;
        RECT  11.8025 20.735 11.8675 20.8 ;
        RECT  11.8025 20.735 11.8675 20.8 ;
        RECT  11.8025 20.735 11.8675 20.8 ;
        RECT  11.5475 21.2275 11.6125 21.2925 ;
        RECT  11.8025 21.5525 11.8675 21.6175 ;
        RECT  11.8025 21.5525 11.8675 21.6175 ;
        RECT  11.8025 21.5525 11.8675 21.6175 ;
        RECT  11.8025 20.735 11.8675 20.8 ;
        RECT  11.8025 20.735 11.8675 20.8 ;
        RECT  11.8025 20.735 11.8675 20.8 ;
        RECT  11.8025 20.735 11.8675 20.8 ;
        RECT  11.8025 20.735 11.8675 20.8 ;
        RECT  11.8025 20.735 11.8675 20.8 ;
        RECT  11.0975 21.5525 11.1625 21.6175 ;
        RECT  11.8025 22.37 11.8675 22.435 ;
        RECT  11.8025 22.37 11.8675 22.435 ;
        RECT  11.8025 22.37 11.8675 22.435 ;
        RECT  11.8025 22.37 11.8675 22.435 ;
        RECT  11.8025 22.37 11.8675 22.435 ;
        RECT  11.8025 22.37 11.8675 22.435 ;
        RECT  11.0975 21.5525 11.1625 21.6175 ;
        RECT  11.8025 21.5525 11.8675 21.6175 ;
        RECT  11.8025 22.37 11.8675 22.435 ;
        RECT  11.8025 22.37 11.8675 22.435 ;
        RECT  11.8025 22.37 11.8675 22.435 ;
        RECT  11.8025 22.37 11.8675 22.435 ;
        RECT  11.8025 22.37 11.8675 22.435 ;
        RECT  11.8025 22.37 11.8675 22.435 ;
        RECT  11.8025 22.37 11.8675 22.435 ;
        RECT  11.8025 22.37 11.8675 22.435 ;
        RECT  11.3525 21.8775 11.4175 21.9425 ;
        RECT  11.0975 22.37 11.1625 22.435 ;
        RECT  11.0975 22.37 11.1625 22.435 ;
        RECT  11.0975 22.37 11.1625 22.435 ;
        RECT  11.0975 22.37 11.1625 22.435 ;
        RECT  11.0975 22.37 11.1625 22.435 ;
        RECT  11.0975 22.37 11.1625 22.435 ;
        RECT  11.8025 22.37 11.8675 22.435 ;
        RECT  11.8025 22.37 11.8675 22.435 ;
        RECT  11.8025 22.37 11.8675 22.435 ;
        RECT  11.8025 22.37 11.8675 22.435 ;
        RECT  11.5475 21.8775 11.6125 21.9425 ;
        RECT  11.8025 21.5525 11.8675 21.6175 ;
        RECT  11.8025 21.5525 11.8675 21.6175 ;
        RECT  11.8025 21.5525 11.8675 21.6175 ;
        RECT  11.8025 22.37 11.8675 22.435 ;
        RECT  11.8025 22.37 11.8675 22.435 ;
        RECT  11.8025 22.37 11.8675 22.435 ;
        RECT  11.8025 22.37 11.8675 22.435 ;
        RECT  11.8025 22.37 11.8675 22.435 ;
        RECT  11.8025 22.37 11.8675 22.435 ;
        RECT  11.0975 21.5525 11.1625 21.6175 ;
        RECT  11.8025 23.425 11.8675 23.49 ;
        RECT  11.8025 23.425 11.8675 23.49 ;
        RECT  11.8025 23.425 11.8675 23.49 ;
        RECT  11.8025 23.425 11.8675 23.49 ;
        RECT  11.8025 23.425 11.8675 23.49 ;
        RECT  11.8025 23.425 11.8675 23.49 ;
        RECT  11.0975 24.2425 11.1625 24.3075 ;
        RECT  11.8025 24.2425 11.8675 24.3075 ;
        RECT  11.8025 23.425 11.8675 23.49 ;
        RECT  11.8025 23.425 11.8675 23.49 ;
        RECT  11.8025 23.425 11.8675 23.49 ;
        RECT  11.8025 23.425 11.8675 23.49 ;
        RECT  11.8025 23.425 11.8675 23.49 ;
        RECT  11.8025 23.425 11.8675 23.49 ;
        RECT  11.8025 23.425 11.8675 23.49 ;
        RECT  11.8025 23.425 11.8675 23.49 ;
        RECT  11.3525 23.9175 11.4175 23.9825 ;
        RECT  11.0975 23.425 11.1625 23.49 ;
        RECT  11.0975 23.425 11.1625 23.49 ;
        RECT  11.0975 23.425 11.1625 23.49 ;
        RECT  11.0975 23.425 11.1625 23.49 ;
        RECT  11.0975 23.425 11.1625 23.49 ;
        RECT  11.0975 23.425 11.1625 23.49 ;
        RECT  11.8025 23.425 11.8675 23.49 ;
        RECT  11.8025 23.425 11.8675 23.49 ;
        RECT  11.8025 23.425 11.8675 23.49 ;
        RECT  11.8025 23.425 11.8675 23.49 ;
        RECT  11.5475 23.9175 11.6125 23.9825 ;
        RECT  11.8025 24.2425 11.8675 24.3075 ;
        RECT  11.8025 24.2425 11.8675 24.3075 ;
        RECT  11.8025 24.2425 11.8675 24.3075 ;
        RECT  11.8025 23.425 11.8675 23.49 ;
        RECT  11.8025 23.425 11.8675 23.49 ;
        RECT  11.8025 23.425 11.8675 23.49 ;
        RECT  11.8025 23.425 11.8675 23.49 ;
        RECT  11.8025 23.425 11.8675 23.49 ;
        RECT  11.8025 23.425 11.8675 23.49 ;
        RECT  11.0975 24.2425 11.1625 24.3075 ;
        RECT  11.8025 25.06 11.8675 25.125 ;
        RECT  11.8025 25.06 11.8675 25.125 ;
        RECT  11.8025 25.06 11.8675 25.125 ;
        RECT  11.8025 25.06 11.8675 25.125 ;
        RECT  11.8025 25.06 11.8675 25.125 ;
        RECT  11.8025 25.06 11.8675 25.125 ;
        RECT  11.0975 24.2425 11.1625 24.3075 ;
        RECT  11.8025 24.2425 11.8675 24.3075 ;
        RECT  11.8025 25.06 11.8675 25.125 ;
        RECT  11.8025 25.06 11.8675 25.125 ;
        RECT  11.8025 25.06 11.8675 25.125 ;
        RECT  11.8025 25.06 11.8675 25.125 ;
        RECT  11.8025 25.06 11.8675 25.125 ;
        RECT  11.8025 25.06 11.8675 25.125 ;
        RECT  11.8025 25.06 11.8675 25.125 ;
        RECT  11.8025 25.06 11.8675 25.125 ;
        RECT  11.3525 24.5675 11.4175 24.6325 ;
        RECT  11.0975 25.06 11.1625 25.125 ;
        RECT  11.0975 25.06 11.1625 25.125 ;
        RECT  11.0975 25.06 11.1625 25.125 ;
        RECT  11.0975 25.06 11.1625 25.125 ;
        RECT  11.0975 25.06 11.1625 25.125 ;
        RECT  11.0975 25.06 11.1625 25.125 ;
        RECT  11.8025 25.06 11.8675 25.125 ;
        RECT  11.8025 25.06 11.8675 25.125 ;
        RECT  11.8025 25.06 11.8675 25.125 ;
        RECT  11.8025 25.06 11.8675 25.125 ;
        RECT  11.5475 24.5675 11.6125 24.6325 ;
        RECT  11.8025 24.2425 11.8675 24.3075 ;
        RECT  11.8025 24.2425 11.8675 24.3075 ;
        RECT  11.8025 24.2425 11.8675 24.3075 ;
        RECT  11.8025 25.06 11.8675 25.125 ;
        RECT  11.8025 25.06 11.8675 25.125 ;
        RECT  11.8025 25.06 11.8675 25.125 ;
        RECT  11.8025 25.06 11.8675 25.125 ;
        RECT  11.8025 25.06 11.8675 25.125 ;
        RECT  11.8025 25.06 11.8675 25.125 ;
        RECT  11.0975 24.2425 11.1625 24.3075 ;
        RECT  11.8025 26.115 11.8675 26.18 ;
        RECT  11.8025 26.115 11.8675 26.18 ;
        RECT  11.8025 26.115 11.8675 26.18 ;
        RECT  11.8025 26.115 11.8675 26.18 ;
        RECT  11.8025 26.115 11.8675 26.18 ;
        RECT  11.8025 26.115 11.8675 26.18 ;
        RECT  11.0975 26.9325 11.1625 26.9975 ;
        RECT  11.8025 26.9325 11.8675 26.9975 ;
        RECT  11.8025 26.115 11.8675 26.18 ;
        RECT  11.8025 26.115 11.8675 26.18 ;
        RECT  11.8025 26.115 11.8675 26.18 ;
        RECT  11.8025 26.115 11.8675 26.18 ;
        RECT  11.8025 26.115 11.8675 26.18 ;
        RECT  11.8025 26.115 11.8675 26.18 ;
        RECT  11.8025 26.115 11.8675 26.18 ;
        RECT  11.8025 26.115 11.8675 26.18 ;
        RECT  11.3525 26.6075 11.4175 26.6725 ;
        RECT  11.0975 26.115 11.1625 26.18 ;
        RECT  11.0975 26.115 11.1625 26.18 ;
        RECT  11.0975 26.115 11.1625 26.18 ;
        RECT  11.0975 26.115 11.1625 26.18 ;
        RECT  11.0975 26.115 11.1625 26.18 ;
        RECT  11.0975 26.115 11.1625 26.18 ;
        RECT  11.8025 26.115 11.8675 26.18 ;
        RECT  11.8025 26.115 11.8675 26.18 ;
        RECT  11.8025 26.115 11.8675 26.18 ;
        RECT  11.8025 26.115 11.8675 26.18 ;
        RECT  11.5475 26.6075 11.6125 26.6725 ;
        RECT  11.8025 26.9325 11.8675 26.9975 ;
        RECT  11.8025 26.9325 11.8675 26.9975 ;
        RECT  11.8025 26.9325 11.8675 26.9975 ;
        RECT  11.8025 26.115 11.8675 26.18 ;
        RECT  11.8025 26.115 11.8675 26.18 ;
        RECT  11.8025 26.115 11.8675 26.18 ;
        RECT  11.8025 26.115 11.8675 26.18 ;
        RECT  11.8025 26.115 11.8675 26.18 ;
        RECT  11.8025 26.115 11.8675 26.18 ;
        RECT  11.0975 26.9325 11.1625 26.9975 ;
        RECT  11.8025 27.75 11.8675 27.815 ;
        RECT  11.8025 27.75 11.8675 27.815 ;
        RECT  11.8025 27.75 11.8675 27.815 ;
        RECT  11.8025 27.75 11.8675 27.815 ;
        RECT  11.8025 27.75 11.8675 27.815 ;
        RECT  11.8025 27.75 11.8675 27.815 ;
        RECT  11.0975 26.9325 11.1625 26.9975 ;
        RECT  11.8025 26.9325 11.8675 26.9975 ;
        RECT  11.8025 27.75 11.8675 27.815 ;
        RECT  11.8025 27.75 11.8675 27.815 ;
        RECT  11.8025 27.75 11.8675 27.815 ;
        RECT  11.8025 27.75 11.8675 27.815 ;
        RECT  11.8025 27.75 11.8675 27.815 ;
        RECT  11.8025 27.75 11.8675 27.815 ;
        RECT  11.8025 27.75 11.8675 27.815 ;
        RECT  11.8025 27.75 11.8675 27.815 ;
        RECT  11.3525 27.2575 11.4175 27.3225 ;
        RECT  11.0975 27.75 11.1625 27.815 ;
        RECT  11.0975 27.75 11.1625 27.815 ;
        RECT  11.0975 27.75 11.1625 27.815 ;
        RECT  11.0975 27.75 11.1625 27.815 ;
        RECT  11.0975 27.75 11.1625 27.815 ;
        RECT  11.0975 27.75 11.1625 27.815 ;
        RECT  11.8025 27.75 11.8675 27.815 ;
        RECT  11.8025 27.75 11.8675 27.815 ;
        RECT  11.8025 27.75 11.8675 27.815 ;
        RECT  11.8025 27.75 11.8675 27.815 ;
        RECT  11.5475 27.2575 11.6125 27.3225 ;
        RECT  11.8025 26.9325 11.8675 26.9975 ;
        RECT  11.8025 26.9325 11.8675 26.9975 ;
        RECT  11.8025 26.9325 11.8675 26.9975 ;
        RECT  11.8025 27.75 11.8675 27.815 ;
        RECT  11.8025 27.75 11.8675 27.815 ;
        RECT  11.8025 27.75 11.8675 27.815 ;
        RECT  11.8025 27.75 11.8675 27.815 ;
        RECT  11.8025 27.75 11.8675 27.815 ;
        RECT  11.8025 27.75 11.8675 27.815 ;
        RECT  11.0975 26.9325 11.1625 26.9975 ;
        RECT  11.8025 28.805 11.8675 28.87 ;
        RECT  11.8025 28.805 11.8675 28.87 ;
        RECT  11.8025 28.805 11.8675 28.87 ;
        RECT  11.8025 28.805 11.8675 28.87 ;
        RECT  11.8025 28.805 11.8675 28.87 ;
        RECT  11.8025 28.805 11.8675 28.87 ;
        RECT  11.0975 29.6225 11.1625 29.6875 ;
        RECT  11.8025 29.6225 11.8675 29.6875 ;
        RECT  11.8025 28.805 11.8675 28.87 ;
        RECT  11.8025 28.805 11.8675 28.87 ;
        RECT  11.8025 28.805 11.8675 28.87 ;
        RECT  11.8025 28.805 11.8675 28.87 ;
        RECT  11.8025 28.805 11.8675 28.87 ;
        RECT  11.8025 28.805 11.8675 28.87 ;
        RECT  11.8025 28.805 11.8675 28.87 ;
        RECT  11.8025 28.805 11.8675 28.87 ;
        RECT  11.3525 29.2975 11.4175 29.3625 ;
        RECT  11.0975 28.805 11.1625 28.87 ;
        RECT  11.0975 28.805 11.1625 28.87 ;
        RECT  11.0975 28.805 11.1625 28.87 ;
        RECT  11.0975 28.805 11.1625 28.87 ;
        RECT  11.0975 28.805 11.1625 28.87 ;
        RECT  11.0975 28.805 11.1625 28.87 ;
        RECT  11.8025 28.805 11.8675 28.87 ;
        RECT  11.8025 28.805 11.8675 28.87 ;
        RECT  11.8025 28.805 11.8675 28.87 ;
        RECT  11.8025 28.805 11.8675 28.87 ;
        RECT  11.5475 29.2975 11.6125 29.3625 ;
        RECT  11.8025 29.6225 11.8675 29.6875 ;
        RECT  11.8025 29.6225 11.8675 29.6875 ;
        RECT  11.8025 29.6225 11.8675 29.6875 ;
        RECT  11.8025 28.805 11.8675 28.87 ;
        RECT  11.8025 28.805 11.8675 28.87 ;
        RECT  11.8025 28.805 11.8675 28.87 ;
        RECT  11.8025 28.805 11.8675 28.87 ;
        RECT  11.8025 28.805 11.8675 28.87 ;
        RECT  11.8025 28.805 11.8675 28.87 ;
        RECT  11.0975 29.6225 11.1625 29.6875 ;
        RECT  11.8025 30.44 11.8675 30.505 ;
        RECT  11.8025 30.44 11.8675 30.505 ;
        RECT  11.8025 30.44 11.8675 30.505 ;
        RECT  11.8025 30.44 11.8675 30.505 ;
        RECT  11.8025 30.44 11.8675 30.505 ;
        RECT  11.8025 30.44 11.8675 30.505 ;
        RECT  11.0975 29.6225 11.1625 29.6875 ;
        RECT  11.8025 29.6225 11.8675 29.6875 ;
        RECT  11.8025 30.44 11.8675 30.505 ;
        RECT  11.8025 30.44 11.8675 30.505 ;
        RECT  11.8025 30.44 11.8675 30.505 ;
        RECT  11.8025 30.44 11.8675 30.505 ;
        RECT  11.8025 30.44 11.8675 30.505 ;
        RECT  11.8025 30.44 11.8675 30.505 ;
        RECT  11.8025 30.44 11.8675 30.505 ;
        RECT  11.8025 30.44 11.8675 30.505 ;
        RECT  11.3525 29.9475 11.4175 30.0125 ;
        RECT  11.0975 30.44 11.1625 30.505 ;
        RECT  11.0975 30.44 11.1625 30.505 ;
        RECT  11.0975 30.44 11.1625 30.505 ;
        RECT  11.0975 30.44 11.1625 30.505 ;
        RECT  11.0975 30.44 11.1625 30.505 ;
        RECT  11.0975 30.44 11.1625 30.505 ;
        RECT  11.8025 30.44 11.8675 30.505 ;
        RECT  11.8025 30.44 11.8675 30.505 ;
        RECT  11.8025 30.44 11.8675 30.505 ;
        RECT  11.8025 30.44 11.8675 30.505 ;
        RECT  11.5475 29.9475 11.6125 30.0125 ;
        RECT  11.8025 29.6225 11.8675 29.6875 ;
        RECT  11.8025 29.6225 11.8675 29.6875 ;
        RECT  11.8025 29.6225 11.8675 29.6875 ;
        RECT  11.8025 30.44 11.8675 30.505 ;
        RECT  11.8025 30.44 11.8675 30.505 ;
        RECT  11.8025 30.44 11.8675 30.505 ;
        RECT  11.8025 30.44 11.8675 30.505 ;
        RECT  11.8025 30.44 11.8675 30.505 ;
        RECT  11.8025 30.44 11.8675 30.505 ;
        RECT  11.0975 29.6225 11.1625 29.6875 ;
        RECT  11.8025 31.495 11.8675 31.56 ;
        RECT  11.8025 31.495 11.8675 31.56 ;
        RECT  11.8025 31.495 11.8675 31.56 ;
        RECT  11.8025 31.495 11.8675 31.56 ;
        RECT  11.8025 31.495 11.8675 31.56 ;
        RECT  11.8025 31.495 11.8675 31.56 ;
        RECT  11.0975 32.3125 11.1625 32.3775 ;
        RECT  11.8025 32.3125 11.8675 32.3775 ;
        RECT  11.8025 31.495 11.8675 31.56 ;
        RECT  11.8025 31.495 11.8675 31.56 ;
        RECT  11.8025 31.495 11.8675 31.56 ;
        RECT  11.8025 31.495 11.8675 31.56 ;
        RECT  11.8025 31.495 11.8675 31.56 ;
        RECT  11.8025 31.495 11.8675 31.56 ;
        RECT  11.8025 31.495 11.8675 31.56 ;
        RECT  11.8025 31.495 11.8675 31.56 ;
        RECT  11.3525 31.9875 11.4175 32.0525 ;
        RECT  11.0975 31.495 11.1625 31.56 ;
        RECT  11.0975 31.495 11.1625 31.56 ;
        RECT  11.0975 31.495 11.1625 31.56 ;
        RECT  11.0975 31.495 11.1625 31.56 ;
        RECT  11.0975 31.495 11.1625 31.56 ;
        RECT  11.0975 31.495 11.1625 31.56 ;
        RECT  11.8025 31.495 11.8675 31.56 ;
        RECT  11.8025 31.495 11.8675 31.56 ;
        RECT  11.8025 31.495 11.8675 31.56 ;
        RECT  11.8025 31.495 11.8675 31.56 ;
        RECT  11.5475 31.9875 11.6125 32.0525 ;
        RECT  11.8025 32.3125 11.8675 32.3775 ;
        RECT  11.8025 32.3125 11.8675 32.3775 ;
        RECT  11.8025 32.3125 11.8675 32.3775 ;
        RECT  11.8025 31.495 11.8675 31.56 ;
        RECT  11.8025 31.495 11.8675 31.56 ;
        RECT  11.8025 31.495 11.8675 31.56 ;
        RECT  11.8025 31.495 11.8675 31.56 ;
        RECT  11.8025 31.495 11.8675 31.56 ;
        RECT  11.8025 31.495 11.8675 31.56 ;
        RECT  11.0975 32.3125 11.1625 32.3775 ;
        RECT  11.8025 33.13 11.8675 33.195 ;
        RECT  11.8025 33.13 11.8675 33.195 ;
        RECT  11.8025 33.13 11.8675 33.195 ;
        RECT  11.8025 33.13 11.8675 33.195 ;
        RECT  11.8025 33.13 11.8675 33.195 ;
        RECT  11.8025 33.13 11.8675 33.195 ;
        RECT  11.0975 32.3125 11.1625 32.3775 ;
        RECT  11.8025 32.3125 11.8675 32.3775 ;
        RECT  11.8025 33.13 11.8675 33.195 ;
        RECT  11.8025 33.13 11.8675 33.195 ;
        RECT  11.8025 33.13 11.8675 33.195 ;
        RECT  11.8025 33.13 11.8675 33.195 ;
        RECT  11.8025 33.13 11.8675 33.195 ;
        RECT  11.8025 33.13 11.8675 33.195 ;
        RECT  11.8025 33.13 11.8675 33.195 ;
        RECT  11.8025 33.13 11.8675 33.195 ;
        RECT  11.3525 32.6375 11.4175 32.7025 ;
        RECT  11.0975 33.13 11.1625 33.195 ;
        RECT  11.0975 33.13 11.1625 33.195 ;
        RECT  11.0975 33.13 11.1625 33.195 ;
        RECT  11.0975 33.13 11.1625 33.195 ;
        RECT  11.0975 33.13 11.1625 33.195 ;
        RECT  11.0975 33.13 11.1625 33.195 ;
        RECT  11.8025 33.13 11.8675 33.195 ;
        RECT  11.8025 33.13 11.8675 33.195 ;
        RECT  11.8025 33.13 11.8675 33.195 ;
        RECT  11.8025 33.13 11.8675 33.195 ;
        RECT  11.5475 32.6375 11.6125 32.7025 ;
        RECT  11.8025 32.3125 11.8675 32.3775 ;
        RECT  11.8025 32.3125 11.8675 32.3775 ;
        RECT  11.8025 32.3125 11.8675 32.3775 ;
        RECT  11.8025 33.13 11.8675 33.195 ;
        RECT  11.8025 33.13 11.8675 33.195 ;
        RECT  11.8025 33.13 11.8675 33.195 ;
        RECT  11.8025 33.13 11.8675 33.195 ;
        RECT  11.8025 33.13 11.8675 33.195 ;
        RECT  11.8025 33.13 11.8675 33.195 ;
        RECT  11.0975 32.3125 11.1625 32.3775 ;
        RECT  11.8025 34.185 11.8675 34.25 ;
        RECT  11.8025 34.185 11.8675 34.25 ;
        RECT  11.8025 34.185 11.8675 34.25 ;
        RECT  11.8025 34.185 11.8675 34.25 ;
        RECT  11.8025 34.185 11.8675 34.25 ;
        RECT  11.8025 34.185 11.8675 34.25 ;
        RECT  11.0975 35.0025 11.1625 35.0675 ;
        RECT  11.8025 35.0025 11.8675 35.0675 ;
        RECT  11.8025 34.185 11.8675 34.25 ;
        RECT  11.8025 34.185 11.8675 34.25 ;
        RECT  11.8025 34.185 11.8675 34.25 ;
        RECT  11.8025 34.185 11.8675 34.25 ;
        RECT  11.8025 34.185 11.8675 34.25 ;
        RECT  11.8025 34.185 11.8675 34.25 ;
        RECT  11.8025 34.185 11.8675 34.25 ;
        RECT  11.8025 34.185 11.8675 34.25 ;
        RECT  11.3525 34.6775 11.4175 34.7425 ;
        RECT  11.0975 34.185 11.1625 34.25 ;
        RECT  11.0975 34.185 11.1625 34.25 ;
        RECT  11.0975 34.185 11.1625 34.25 ;
        RECT  11.0975 34.185 11.1625 34.25 ;
        RECT  11.0975 34.185 11.1625 34.25 ;
        RECT  11.0975 34.185 11.1625 34.25 ;
        RECT  11.8025 34.185 11.8675 34.25 ;
        RECT  11.8025 34.185 11.8675 34.25 ;
        RECT  11.8025 34.185 11.8675 34.25 ;
        RECT  11.8025 34.185 11.8675 34.25 ;
        RECT  11.5475 34.6775 11.6125 34.7425 ;
        RECT  11.8025 35.0025 11.8675 35.0675 ;
        RECT  11.8025 35.0025 11.8675 35.0675 ;
        RECT  11.8025 35.0025 11.8675 35.0675 ;
        RECT  11.8025 34.185 11.8675 34.25 ;
        RECT  11.8025 34.185 11.8675 34.25 ;
        RECT  11.8025 34.185 11.8675 34.25 ;
        RECT  11.8025 34.185 11.8675 34.25 ;
        RECT  11.8025 34.185 11.8675 34.25 ;
        RECT  11.8025 34.185 11.8675 34.25 ;
        RECT  11.0975 35.0025 11.1625 35.0675 ;
        RECT  11.8025 35.82 11.8675 35.885 ;
        RECT  11.8025 35.82 11.8675 35.885 ;
        RECT  11.8025 35.82 11.8675 35.885 ;
        RECT  11.8025 35.82 11.8675 35.885 ;
        RECT  11.8025 35.82 11.8675 35.885 ;
        RECT  11.8025 35.82 11.8675 35.885 ;
        RECT  11.0975 35.0025 11.1625 35.0675 ;
        RECT  11.8025 35.0025 11.8675 35.0675 ;
        RECT  11.8025 35.82 11.8675 35.885 ;
        RECT  11.8025 35.82 11.8675 35.885 ;
        RECT  11.8025 35.82 11.8675 35.885 ;
        RECT  11.8025 35.82 11.8675 35.885 ;
        RECT  11.8025 35.82 11.8675 35.885 ;
        RECT  11.8025 35.82 11.8675 35.885 ;
        RECT  11.8025 35.82 11.8675 35.885 ;
        RECT  11.8025 35.82 11.8675 35.885 ;
        RECT  11.3525 35.3275 11.4175 35.3925 ;
        RECT  11.0975 35.82 11.1625 35.885 ;
        RECT  11.0975 35.82 11.1625 35.885 ;
        RECT  11.0975 35.82 11.1625 35.885 ;
        RECT  11.0975 35.82 11.1625 35.885 ;
        RECT  11.0975 35.82 11.1625 35.885 ;
        RECT  11.0975 35.82 11.1625 35.885 ;
        RECT  11.8025 35.82 11.8675 35.885 ;
        RECT  11.8025 35.82 11.8675 35.885 ;
        RECT  11.8025 35.82 11.8675 35.885 ;
        RECT  11.8025 35.82 11.8675 35.885 ;
        RECT  11.5475 35.3275 11.6125 35.3925 ;
        RECT  11.8025 35.0025 11.8675 35.0675 ;
        RECT  11.8025 35.0025 11.8675 35.0675 ;
        RECT  11.8025 35.0025 11.8675 35.0675 ;
        RECT  11.8025 35.82 11.8675 35.885 ;
        RECT  11.8025 35.82 11.8675 35.885 ;
        RECT  11.8025 35.82 11.8675 35.885 ;
        RECT  11.8025 35.82 11.8675 35.885 ;
        RECT  11.8025 35.82 11.8675 35.885 ;
        RECT  11.8025 35.82 11.8675 35.885 ;
        RECT  11.0975 35.0025 11.1625 35.0675 ;
        RECT  11.8025 36.875 11.8675 36.94 ;
        RECT  11.8025 36.875 11.8675 36.94 ;
        RECT  11.8025 36.875 11.8675 36.94 ;
        RECT  11.8025 36.875 11.8675 36.94 ;
        RECT  11.8025 36.875 11.8675 36.94 ;
        RECT  11.8025 36.875 11.8675 36.94 ;
        RECT  11.0975 37.6925 11.1625 37.7575 ;
        RECT  11.8025 37.6925 11.8675 37.7575 ;
        RECT  11.8025 36.875 11.8675 36.94 ;
        RECT  11.8025 36.875 11.8675 36.94 ;
        RECT  11.8025 36.875 11.8675 36.94 ;
        RECT  11.8025 36.875 11.8675 36.94 ;
        RECT  11.8025 36.875 11.8675 36.94 ;
        RECT  11.8025 36.875 11.8675 36.94 ;
        RECT  11.8025 36.875 11.8675 36.94 ;
        RECT  11.8025 36.875 11.8675 36.94 ;
        RECT  11.3525 37.3675 11.4175 37.4325 ;
        RECT  11.0975 36.875 11.1625 36.94 ;
        RECT  11.0975 36.875 11.1625 36.94 ;
        RECT  11.0975 36.875 11.1625 36.94 ;
        RECT  11.0975 36.875 11.1625 36.94 ;
        RECT  11.0975 36.875 11.1625 36.94 ;
        RECT  11.0975 36.875 11.1625 36.94 ;
        RECT  11.8025 36.875 11.8675 36.94 ;
        RECT  11.8025 36.875 11.8675 36.94 ;
        RECT  11.8025 36.875 11.8675 36.94 ;
        RECT  11.8025 36.875 11.8675 36.94 ;
        RECT  11.5475 37.3675 11.6125 37.4325 ;
        RECT  11.8025 37.6925 11.8675 37.7575 ;
        RECT  11.8025 37.6925 11.8675 37.7575 ;
        RECT  11.8025 37.6925 11.8675 37.7575 ;
        RECT  11.8025 36.875 11.8675 36.94 ;
        RECT  11.8025 36.875 11.8675 36.94 ;
        RECT  11.8025 36.875 11.8675 36.94 ;
        RECT  11.8025 36.875 11.8675 36.94 ;
        RECT  11.8025 36.875 11.8675 36.94 ;
        RECT  11.8025 36.875 11.8675 36.94 ;
        RECT  11.0975 37.6925 11.1625 37.7575 ;
        RECT  11.8025 38.51 11.8675 38.575 ;
        RECT  11.8025 38.51 11.8675 38.575 ;
        RECT  11.8025 38.51 11.8675 38.575 ;
        RECT  11.8025 38.51 11.8675 38.575 ;
        RECT  11.8025 38.51 11.8675 38.575 ;
        RECT  11.8025 38.51 11.8675 38.575 ;
        RECT  11.0975 37.6925 11.1625 37.7575 ;
        RECT  11.8025 37.6925 11.8675 37.7575 ;
        RECT  11.8025 38.51 11.8675 38.575 ;
        RECT  11.8025 38.51 11.8675 38.575 ;
        RECT  11.8025 38.51 11.8675 38.575 ;
        RECT  11.8025 38.51 11.8675 38.575 ;
        RECT  11.8025 38.51 11.8675 38.575 ;
        RECT  11.8025 38.51 11.8675 38.575 ;
        RECT  11.8025 38.51 11.8675 38.575 ;
        RECT  11.8025 38.51 11.8675 38.575 ;
        RECT  11.3525 38.0175 11.4175 38.0825 ;
        RECT  11.0975 38.51 11.1625 38.575 ;
        RECT  11.0975 38.51 11.1625 38.575 ;
        RECT  11.0975 38.51 11.1625 38.575 ;
        RECT  11.0975 38.51 11.1625 38.575 ;
        RECT  11.0975 38.51 11.1625 38.575 ;
        RECT  11.0975 38.51 11.1625 38.575 ;
        RECT  11.8025 38.51 11.8675 38.575 ;
        RECT  11.8025 38.51 11.8675 38.575 ;
        RECT  11.8025 38.51 11.8675 38.575 ;
        RECT  11.8025 38.51 11.8675 38.575 ;
        RECT  11.5475 38.0175 11.6125 38.0825 ;
        RECT  11.8025 37.6925 11.8675 37.7575 ;
        RECT  11.8025 37.6925 11.8675 37.7575 ;
        RECT  11.8025 37.6925 11.8675 37.7575 ;
        RECT  11.8025 38.51 11.8675 38.575 ;
        RECT  11.8025 38.51 11.8675 38.575 ;
        RECT  11.8025 38.51 11.8675 38.575 ;
        RECT  11.8025 38.51 11.8675 38.575 ;
        RECT  11.8025 38.51 11.8675 38.575 ;
        RECT  11.8025 38.51 11.8675 38.575 ;
        RECT  11.0975 37.6925 11.1625 37.7575 ;
        RECT  11.8025 39.565 11.8675 39.63 ;
        RECT  11.8025 39.565 11.8675 39.63 ;
        RECT  11.8025 39.565 11.8675 39.63 ;
        RECT  11.8025 39.565 11.8675 39.63 ;
        RECT  11.8025 39.565 11.8675 39.63 ;
        RECT  11.8025 39.565 11.8675 39.63 ;
        RECT  11.0975 40.3825 11.1625 40.4475 ;
        RECT  11.8025 40.3825 11.8675 40.4475 ;
        RECT  11.8025 39.565 11.8675 39.63 ;
        RECT  11.8025 39.565 11.8675 39.63 ;
        RECT  11.8025 39.565 11.8675 39.63 ;
        RECT  11.8025 39.565 11.8675 39.63 ;
        RECT  11.8025 39.565 11.8675 39.63 ;
        RECT  11.8025 39.565 11.8675 39.63 ;
        RECT  11.8025 39.565 11.8675 39.63 ;
        RECT  11.8025 39.565 11.8675 39.63 ;
        RECT  11.3525 40.0575 11.4175 40.1225 ;
        RECT  11.0975 39.565 11.1625 39.63 ;
        RECT  11.0975 39.565 11.1625 39.63 ;
        RECT  11.0975 39.565 11.1625 39.63 ;
        RECT  11.0975 39.565 11.1625 39.63 ;
        RECT  11.0975 39.565 11.1625 39.63 ;
        RECT  11.0975 39.565 11.1625 39.63 ;
        RECT  11.8025 39.565 11.8675 39.63 ;
        RECT  11.8025 39.565 11.8675 39.63 ;
        RECT  11.8025 39.565 11.8675 39.63 ;
        RECT  11.8025 39.565 11.8675 39.63 ;
        RECT  11.5475 40.0575 11.6125 40.1225 ;
        RECT  11.8025 40.3825 11.8675 40.4475 ;
        RECT  11.8025 40.3825 11.8675 40.4475 ;
        RECT  11.8025 40.3825 11.8675 40.4475 ;
        RECT  11.8025 39.565 11.8675 39.63 ;
        RECT  11.8025 39.565 11.8675 39.63 ;
        RECT  11.8025 39.565 11.8675 39.63 ;
        RECT  11.8025 39.565 11.8675 39.63 ;
        RECT  11.8025 39.565 11.8675 39.63 ;
        RECT  11.8025 39.565 11.8675 39.63 ;
        RECT  11.0975 40.3825 11.1625 40.4475 ;
        RECT  12.5075 19.68 12.5725 19.745 ;
        RECT  12.5075 19.68 12.5725 19.745 ;
        RECT  12.5075 19.68 12.5725 19.745 ;
        RECT  12.5075 19.68 12.5725 19.745 ;
        RECT  12.5075 19.68 12.5725 19.745 ;
        RECT  12.5075 19.68 12.5725 19.745 ;
        RECT  11.8025 18.8625 11.8675 18.9275 ;
        RECT  12.5075 18.8625 12.5725 18.9275 ;
        RECT  12.5075 19.68 12.5725 19.745 ;
        RECT  12.5075 19.68 12.5725 19.745 ;
        RECT  12.5075 19.68 12.5725 19.745 ;
        RECT  12.5075 19.68 12.5725 19.745 ;
        RECT  12.5075 19.68 12.5725 19.745 ;
        RECT  12.5075 19.68 12.5725 19.745 ;
        RECT  12.5075 19.68 12.5725 19.745 ;
        RECT  12.5075 19.68 12.5725 19.745 ;
        RECT  12.0575 19.1875 12.1225 19.2525 ;
        RECT  11.8025 19.68 11.8675 19.745 ;
        RECT  11.8025 19.68 11.8675 19.745 ;
        RECT  11.8025 19.68 11.8675 19.745 ;
        RECT  11.8025 19.68 11.8675 19.745 ;
        RECT  11.8025 19.68 11.8675 19.745 ;
        RECT  11.8025 19.68 11.8675 19.745 ;
        RECT  12.5075 19.68 12.5725 19.745 ;
        RECT  12.5075 19.68 12.5725 19.745 ;
        RECT  12.5075 19.68 12.5725 19.745 ;
        RECT  12.5075 19.68 12.5725 19.745 ;
        RECT  12.2525 19.1875 12.3175 19.2525 ;
        RECT  12.5075 18.8625 12.5725 18.9275 ;
        RECT  12.5075 18.8625 12.5725 18.9275 ;
        RECT  12.5075 18.8625 12.5725 18.9275 ;
        RECT  12.5075 19.68 12.5725 19.745 ;
        RECT  12.5075 19.68 12.5725 19.745 ;
        RECT  12.5075 19.68 12.5725 19.745 ;
        RECT  12.5075 19.68 12.5725 19.745 ;
        RECT  12.5075 19.68 12.5725 19.745 ;
        RECT  12.5075 19.68 12.5725 19.745 ;
        RECT  11.8025 18.8625 11.8675 18.9275 ;
        RECT  12.5075 20.735 12.5725 20.8 ;
        RECT  12.5075 20.735 12.5725 20.8 ;
        RECT  12.5075 20.735 12.5725 20.8 ;
        RECT  12.5075 20.735 12.5725 20.8 ;
        RECT  12.5075 20.735 12.5725 20.8 ;
        RECT  12.5075 20.735 12.5725 20.8 ;
        RECT  11.8025 21.5525 11.8675 21.6175 ;
        RECT  12.5075 21.5525 12.5725 21.6175 ;
        RECT  12.5075 20.735 12.5725 20.8 ;
        RECT  12.5075 20.735 12.5725 20.8 ;
        RECT  12.5075 20.735 12.5725 20.8 ;
        RECT  12.5075 20.735 12.5725 20.8 ;
        RECT  12.5075 20.735 12.5725 20.8 ;
        RECT  12.5075 20.735 12.5725 20.8 ;
        RECT  12.5075 20.735 12.5725 20.8 ;
        RECT  12.5075 20.735 12.5725 20.8 ;
        RECT  12.0575 21.2275 12.1225 21.2925 ;
        RECT  11.8025 20.735 11.8675 20.8 ;
        RECT  11.8025 20.735 11.8675 20.8 ;
        RECT  11.8025 20.735 11.8675 20.8 ;
        RECT  11.8025 20.735 11.8675 20.8 ;
        RECT  11.8025 20.735 11.8675 20.8 ;
        RECT  11.8025 20.735 11.8675 20.8 ;
        RECT  12.5075 20.735 12.5725 20.8 ;
        RECT  12.5075 20.735 12.5725 20.8 ;
        RECT  12.5075 20.735 12.5725 20.8 ;
        RECT  12.5075 20.735 12.5725 20.8 ;
        RECT  12.2525 21.2275 12.3175 21.2925 ;
        RECT  12.5075 21.5525 12.5725 21.6175 ;
        RECT  12.5075 21.5525 12.5725 21.6175 ;
        RECT  12.5075 21.5525 12.5725 21.6175 ;
        RECT  12.5075 20.735 12.5725 20.8 ;
        RECT  12.5075 20.735 12.5725 20.8 ;
        RECT  12.5075 20.735 12.5725 20.8 ;
        RECT  12.5075 20.735 12.5725 20.8 ;
        RECT  12.5075 20.735 12.5725 20.8 ;
        RECT  12.5075 20.735 12.5725 20.8 ;
        RECT  11.8025 21.5525 11.8675 21.6175 ;
        RECT  12.5075 22.37 12.5725 22.435 ;
        RECT  12.5075 22.37 12.5725 22.435 ;
        RECT  12.5075 22.37 12.5725 22.435 ;
        RECT  12.5075 22.37 12.5725 22.435 ;
        RECT  12.5075 22.37 12.5725 22.435 ;
        RECT  12.5075 22.37 12.5725 22.435 ;
        RECT  11.8025 21.5525 11.8675 21.6175 ;
        RECT  12.5075 21.5525 12.5725 21.6175 ;
        RECT  12.5075 22.37 12.5725 22.435 ;
        RECT  12.5075 22.37 12.5725 22.435 ;
        RECT  12.5075 22.37 12.5725 22.435 ;
        RECT  12.5075 22.37 12.5725 22.435 ;
        RECT  12.5075 22.37 12.5725 22.435 ;
        RECT  12.5075 22.37 12.5725 22.435 ;
        RECT  12.5075 22.37 12.5725 22.435 ;
        RECT  12.5075 22.37 12.5725 22.435 ;
        RECT  12.0575 21.8775 12.1225 21.9425 ;
        RECT  11.8025 22.37 11.8675 22.435 ;
        RECT  11.8025 22.37 11.8675 22.435 ;
        RECT  11.8025 22.37 11.8675 22.435 ;
        RECT  11.8025 22.37 11.8675 22.435 ;
        RECT  11.8025 22.37 11.8675 22.435 ;
        RECT  11.8025 22.37 11.8675 22.435 ;
        RECT  12.5075 22.37 12.5725 22.435 ;
        RECT  12.5075 22.37 12.5725 22.435 ;
        RECT  12.5075 22.37 12.5725 22.435 ;
        RECT  12.5075 22.37 12.5725 22.435 ;
        RECT  12.2525 21.8775 12.3175 21.9425 ;
        RECT  12.5075 21.5525 12.5725 21.6175 ;
        RECT  12.5075 21.5525 12.5725 21.6175 ;
        RECT  12.5075 21.5525 12.5725 21.6175 ;
        RECT  12.5075 22.37 12.5725 22.435 ;
        RECT  12.5075 22.37 12.5725 22.435 ;
        RECT  12.5075 22.37 12.5725 22.435 ;
        RECT  12.5075 22.37 12.5725 22.435 ;
        RECT  12.5075 22.37 12.5725 22.435 ;
        RECT  12.5075 22.37 12.5725 22.435 ;
        RECT  11.8025 21.5525 11.8675 21.6175 ;
        RECT  12.5075 23.425 12.5725 23.49 ;
        RECT  12.5075 23.425 12.5725 23.49 ;
        RECT  12.5075 23.425 12.5725 23.49 ;
        RECT  12.5075 23.425 12.5725 23.49 ;
        RECT  12.5075 23.425 12.5725 23.49 ;
        RECT  12.5075 23.425 12.5725 23.49 ;
        RECT  11.8025 24.2425 11.8675 24.3075 ;
        RECT  12.5075 24.2425 12.5725 24.3075 ;
        RECT  12.5075 23.425 12.5725 23.49 ;
        RECT  12.5075 23.425 12.5725 23.49 ;
        RECT  12.5075 23.425 12.5725 23.49 ;
        RECT  12.5075 23.425 12.5725 23.49 ;
        RECT  12.5075 23.425 12.5725 23.49 ;
        RECT  12.5075 23.425 12.5725 23.49 ;
        RECT  12.5075 23.425 12.5725 23.49 ;
        RECT  12.5075 23.425 12.5725 23.49 ;
        RECT  12.0575 23.9175 12.1225 23.9825 ;
        RECT  11.8025 23.425 11.8675 23.49 ;
        RECT  11.8025 23.425 11.8675 23.49 ;
        RECT  11.8025 23.425 11.8675 23.49 ;
        RECT  11.8025 23.425 11.8675 23.49 ;
        RECT  11.8025 23.425 11.8675 23.49 ;
        RECT  11.8025 23.425 11.8675 23.49 ;
        RECT  12.5075 23.425 12.5725 23.49 ;
        RECT  12.5075 23.425 12.5725 23.49 ;
        RECT  12.5075 23.425 12.5725 23.49 ;
        RECT  12.5075 23.425 12.5725 23.49 ;
        RECT  12.2525 23.9175 12.3175 23.9825 ;
        RECT  12.5075 24.2425 12.5725 24.3075 ;
        RECT  12.5075 24.2425 12.5725 24.3075 ;
        RECT  12.5075 24.2425 12.5725 24.3075 ;
        RECT  12.5075 23.425 12.5725 23.49 ;
        RECT  12.5075 23.425 12.5725 23.49 ;
        RECT  12.5075 23.425 12.5725 23.49 ;
        RECT  12.5075 23.425 12.5725 23.49 ;
        RECT  12.5075 23.425 12.5725 23.49 ;
        RECT  12.5075 23.425 12.5725 23.49 ;
        RECT  11.8025 24.2425 11.8675 24.3075 ;
        RECT  12.5075 25.06 12.5725 25.125 ;
        RECT  12.5075 25.06 12.5725 25.125 ;
        RECT  12.5075 25.06 12.5725 25.125 ;
        RECT  12.5075 25.06 12.5725 25.125 ;
        RECT  12.5075 25.06 12.5725 25.125 ;
        RECT  12.5075 25.06 12.5725 25.125 ;
        RECT  11.8025 24.2425 11.8675 24.3075 ;
        RECT  12.5075 24.2425 12.5725 24.3075 ;
        RECT  12.5075 25.06 12.5725 25.125 ;
        RECT  12.5075 25.06 12.5725 25.125 ;
        RECT  12.5075 25.06 12.5725 25.125 ;
        RECT  12.5075 25.06 12.5725 25.125 ;
        RECT  12.5075 25.06 12.5725 25.125 ;
        RECT  12.5075 25.06 12.5725 25.125 ;
        RECT  12.5075 25.06 12.5725 25.125 ;
        RECT  12.5075 25.06 12.5725 25.125 ;
        RECT  12.0575 24.5675 12.1225 24.6325 ;
        RECT  11.8025 25.06 11.8675 25.125 ;
        RECT  11.8025 25.06 11.8675 25.125 ;
        RECT  11.8025 25.06 11.8675 25.125 ;
        RECT  11.8025 25.06 11.8675 25.125 ;
        RECT  11.8025 25.06 11.8675 25.125 ;
        RECT  11.8025 25.06 11.8675 25.125 ;
        RECT  12.5075 25.06 12.5725 25.125 ;
        RECT  12.5075 25.06 12.5725 25.125 ;
        RECT  12.5075 25.06 12.5725 25.125 ;
        RECT  12.5075 25.06 12.5725 25.125 ;
        RECT  12.2525 24.5675 12.3175 24.6325 ;
        RECT  12.5075 24.2425 12.5725 24.3075 ;
        RECT  12.5075 24.2425 12.5725 24.3075 ;
        RECT  12.5075 24.2425 12.5725 24.3075 ;
        RECT  12.5075 25.06 12.5725 25.125 ;
        RECT  12.5075 25.06 12.5725 25.125 ;
        RECT  12.5075 25.06 12.5725 25.125 ;
        RECT  12.5075 25.06 12.5725 25.125 ;
        RECT  12.5075 25.06 12.5725 25.125 ;
        RECT  12.5075 25.06 12.5725 25.125 ;
        RECT  11.8025 24.2425 11.8675 24.3075 ;
        RECT  12.5075 26.115 12.5725 26.18 ;
        RECT  12.5075 26.115 12.5725 26.18 ;
        RECT  12.5075 26.115 12.5725 26.18 ;
        RECT  12.5075 26.115 12.5725 26.18 ;
        RECT  12.5075 26.115 12.5725 26.18 ;
        RECT  12.5075 26.115 12.5725 26.18 ;
        RECT  11.8025 26.9325 11.8675 26.9975 ;
        RECT  12.5075 26.9325 12.5725 26.9975 ;
        RECT  12.5075 26.115 12.5725 26.18 ;
        RECT  12.5075 26.115 12.5725 26.18 ;
        RECT  12.5075 26.115 12.5725 26.18 ;
        RECT  12.5075 26.115 12.5725 26.18 ;
        RECT  12.5075 26.115 12.5725 26.18 ;
        RECT  12.5075 26.115 12.5725 26.18 ;
        RECT  12.5075 26.115 12.5725 26.18 ;
        RECT  12.5075 26.115 12.5725 26.18 ;
        RECT  12.0575 26.6075 12.1225 26.6725 ;
        RECT  11.8025 26.115 11.8675 26.18 ;
        RECT  11.8025 26.115 11.8675 26.18 ;
        RECT  11.8025 26.115 11.8675 26.18 ;
        RECT  11.8025 26.115 11.8675 26.18 ;
        RECT  11.8025 26.115 11.8675 26.18 ;
        RECT  11.8025 26.115 11.8675 26.18 ;
        RECT  12.5075 26.115 12.5725 26.18 ;
        RECT  12.5075 26.115 12.5725 26.18 ;
        RECT  12.5075 26.115 12.5725 26.18 ;
        RECT  12.5075 26.115 12.5725 26.18 ;
        RECT  12.2525 26.6075 12.3175 26.6725 ;
        RECT  12.5075 26.9325 12.5725 26.9975 ;
        RECT  12.5075 26.9325 12.5725 26.9975 ;
        RECT  12.5075 26.9325 12.5725 26.9975 ;
        RECT  12.5075 26.115 12.5725 26.18 ;
        RECT  12.5075 26.115 12.5725 26.18 ;
        RECT  12.5075 26.115 12.5725 26.18 ;
        RECT  12.5075 26.115 12.5725 26.18 ;
        RECT  12.5075 26.115 12.5725 26.18 ;
        RECT  12.5075 26.115 12.5725 26.18 ;
        RECT  11.8025 26.9325 11.8675 26.9975 ;
        RECT  12.5075 27.75 12.5725 27.815 ;
        RECT  12.5075 27.75 12.5725 27.815 ;
        RECT  12.5075 27.75 12.5725 27.815 ;
        RECT  12.5075 27.75 12.5725 27.815 ;
        RECT  12.5075 27.75 12.5725 27.815 ;
        RECT  12.5075 27.75 12.5725 27.815 ;
        RECT  11.8025 26.9325 11.8675 26.9975 ;
        RECT  12.5075 26.9325 12.5725 26.9975 ;
        RECT  12.5075 27.75 12.5725 27.815 ;
        RECT  12.5075 27.75 12.5725 27.815 ;
        RECT  12.5075 27.75 12.5725 27.815 ;
        RECT  12.5075 27.75 12.5725 27.815 ;
        RECT  12.5075 27.75 12.5725 27.815 ;
        RECT  12.5075 27.75 12.5725 27.815 ;
        RECT  12.5075 27.75 12.5725 27.815 ;
        RECT  12.5075 27.75 12.5725 27.815 ;
        RECT  12.0575 27.2575 12.1225 27.3225 ;
        RECT  11.8025 27.75 11.8675 27.815 ;
        RECT  11.8025 27.75 11.8675 27.815 ;
        RECT  11.8025 27.75 11.8675 27.815 ;
        RECT  11.8025 27.75 11.8675 27.815 ;
        RECT  11.8025 27.75 11.8675 27.815 ;
        RECT  11.8025 27.75 11.8675 27.815 ;
        RECT  12.5075 27.75 12.5725 27.815 ;
        RECT  12.5075 27.75 12.5725 27.815 ;
        RECT  12.5075 27.75 12.5725 27.815 ;
        RECT  12.5075 27.75 12.5725 27.815 ;
        RECT  12.2525 27.2575 12.3175 27.3225 ;
        RECT  12.5075 26.9325 12.5725 26.9975 ;
        RECT  12.5075 26.9325 12.5725 26.9975 ;
        RECT  12.5075 26.9325 12.5725 26.9975 ;
        RECT  12.5075 27.75 12.5725 27.815 ;
        RECT  12.5075 27.75 12.5725 27.815 ;
        RECT  12.5075 27.75 12.5725 27.815 ;
        RECT  12.5075 27.75 12.5725 27.815 ;
        RECT  12.5075 27.75 12.5725 27.815 ;
        RECT  12.5075 27.75 12.5725 27.815 ;
        RECT  11.8025 26.9325 11.8675 26.9975 ;
        RECT  12.5075 28.805 12.5725 28.87 ;
        RECT  12.5075 28.805 12.5725 28.87 ;
        RECT  12.5075 28.805 12.5725 28.87 ;
        RECT  12.5075 28.805 12.5725 28.87 ;
        RECT  12.5075 28.805 12.5725 28.87 ;
        RECT  12.5075 28.805 12.5725 28.87 ;
        RECT  11.8025 29.6225 11.8675 29.6875 ;
        RECT  12.5075 29.6225 12.5725 29.6875 ;
        RECT  12.5075 28.805 12.5725 28.87 ;
        RECT  12.5075 28.805 12.5725 28.87 ;
        RECT  12.5075 28.805 12.5725 28.87 ;
        RECT  12.5075 28.805 12.5725 28.87 ;
        RECT  12.5075 28.805 12.5725 28.87 ;
        RECT  12.5075 28.805 12.5725 28.87 ;
        RECT  12.5075 28.805 12.5725 28.87 ;
        RECT  12.5075 28.805 12.5725 28.87 ;
        RECT  12.0575 29.2975 12.1225 29.3625 ;
        RECT  11.8025 28.805 11.8675 28.87 ;
        RECT  11.8025 28.805 11.8675 28.87 ;
        RECT  11.8025 28.805 11.8675 28.87 ;
        RECT  11.8025 28.805 11.8675 28.87 ;
        RECT  11.8025 28.805 11.8675 28.87 ;
        RECT  11.8025 28.805 11.8675 28.87 ;
        RECT  12.5075 28.805 12.5725 28.87 ;
        RECT  12.5075 28.805 12.5725 28.87 ;
        RECT  12.5075 28.805 12.5725 28.87 ;
        RECT  12.5075 28.805 12.5725 28.87 ;
        RECT  12.2525 29.2975 12.3175 29.3625 ;
        RECT  12.5075 29.6225 12.5725 29.6875 ;
        RECT  12.5075 29.6225 12.5725 29.6875 ;
        RECT  12.5075 29.6225 12.5725 29.6875 ;
        RECT  12.5075 28.805 12.5725 28.87 ;
        RECT  12.5075 28.805 12.5725 28.87 ;
        RECT  12.5075 28.805 12.5725 28.87 ;
        RECT  12.5075 28.805 12.5725 28.87 ;
        RECT  12.5075 28.805 12.5725 28.87 ;
        RECT  12.5075 28.805 12.5725 28.87 ;
        RECT  11.8025 29.6225 11.8675 29.6875 ;
        RECT  12.5075 30.44 12.5725 30.505 ;
        RECT  12.5075 30.44 12.5725 30.505 ;
        RECT  12.5075 30.44 12.5725 30.505 ;
        RECT  12.5075 30.44 12.5725 30.505 ;
        RECT  12.5075 30.44 12.5725 30.505 ;
        RECT  12.5075 30.44 12.5725 30.505 ;
        RECT  11.8025 29.6225 11.8675 29.6875 ;
        RECT  12.5075 29.6225 12.5725 29.6875 ;
        RECT  12.5075 30.44 12.5725 30.505 ;
        RECT  12.5075 30.44 12.5725 30.505 ;
        RECT  12.5075 30.44 12.5725 30.505 ;
        RECT  12.5075 30.44 12.5725 30.505 ;
        RECT  12.5075 30.44 12.5725 30.505 ;
        RECT  12.5075 30.44 12.5725 30.505 ;
        RECT  12.5075 30.44 12.5725 30.505 ;
        RECT  12.5075 30.44 12.5725 30.505 ;
        RECT  12.0575 29.9475 12.1225 30.0125 ;
        RECT  11.8025 30.44 11.8675 30.505 ;
        RECT  11.8025 30.44 11.8675 30.505 ;
        RECT  11.8025 30.44 11.8675 30.505 ;
        RECT  11.8025 30.44 11.8675 30.505 ;
        RECT  11.8025 30.44 11.8675 30.505 ;
        RECT  11.8025 30.44 11.8675 30.505 ;
        RECT  12.5075 30.44 12.5725 30.505 ;
        RECT  12.5075 30.44 12.5725 30.505 ;
        RECT  12.5075 30.44 12.5725 30.505 ;
        RECT  12.5075 30.44 12.5725 30.505 ;
        RECT  12.2525 29.9475 12.3175 30.0125 ;
        RECT  12.5075 29.6225 12.5725 29.6875 ;
        RECT  12.5075 29.6225 12.5725 29.6875 ;
        RECT  12.5075 29.6225 12.5725 29.6875 ;
        RECT  12.5075 30.44 12.5725 30.505 ;
        RECT  12.5075 30.44 12.5725 30.505 ;
        RECT  12.5075 30.44 12.5725 30.505 ;
        RECT  12.5075 30.44 12.5725 30.505 ;
        RECT  12.5075 30.44 12.5725 30.505 ;
        RECT  12.5075 30.44 12.5725 30.505 ;
        RECT  11.8025 29.6225 11.8675 29.6875 ;
        RECT  12.5075 31.495 12.5725 31.56 ;
        RECT  12.5075 31.495 12.5725 31.56 ;
        RECT  12.5075 31.495 12.5725 31.56 ;
        RECT  12.5075 31.495 12.5725 31.56 ;
        RECT  12.5075 31.495 12.5725 31.56 ;
        RECT  12.5075 31.495 12.5725 31.56 ;
        RECT  11.8025 32.3125 11.8675 32.3775 ;
        RECT  12.5075 32.3125 12.5725 32.3775 ;
        RECT  12.5075 31.495 12.5725 31.56 ;
        RECT  12.5075 31.495 12.5725 31.56 ;
        RECT  12.5075 31.495 12.5725 31.56 ;
        RECT  12.5075 31.495 12.5725 31.56 ;
        RECT  12.5075 31.495 12.5725 31.56 ;
        RECT  12.5075 31.495 12.5725 31.56 ;
        RECT  12.5075 31.495 12.5725 31.56 ;
        RECT  12.5075 31.495 12.5725 31.56 ;
        RECT  12.0575 31.9875 12.1225 32.0525 ;
        RECT  11.8025 31.495 11.8675 31.56 ;
        RECT  11.8025 31.495 11.8675 31.56 ;
        RECT  11.8025 31.495 11.8675 31.56 ;
        RECT  11.8025 31.495 11.8675 31.56 ;
        RECT  11.8025 31.495 11.8675 31.56 ;
        RECT  11.8025 31.495 11.8675 31.56 ;
        RECT  12.5075 31.495 12.5725 31.56 ;
        RECT  12.5075 31.495 12.5725 31.56 ;
        RECT  12.5075 31.495 12.5725 31.56 ;
        RECT  12.5075 31.495 12.5725 31.56 ;
        RECT  12.2525 31.9875 12.3175 32.0525 ;
        RECT  12.5075 32.3125 12.5725 32.3775 ;
        RECT  12.5075 32.3125 12.5725 32.3775 ;
        RECT  12.5075 32.3125 12.5725 32.3775 ;
        RECT  12.5075 31.495 12.5725 31.56 ;
        RECT  12.5075 31.495 12.5725 31.56 ;
        RECT  12.5075 31.495 12.5725 31.56 ;
        RECT  12.5075 31.495 12.5725 31.56 ;
        RECT  12.5075 31.495 12.5725 31.56 ;
        RECT  12.5075 31.495 12.5725 31.56 ;
        RECT  11.8025 32.3125 11.8675 32.3775 ;
        RECT  12.5075 33.13 12.5725 33.195 ;
        RECT  12.5075 33.13 12.5725 33.195 ;
        RECT  12.5075 33.13 12.5725 33.195 ;
        RECT  12.5075 33.13 12.5725 33.195 ;
        RECT  12.5075 33.13 12.5725 33.195 ;
        RECT  12.5075 33.13 12.5725 33.195 ;
        RECT  11.8025 32.3125 11.8675 32.3775 ;
        RECT  12.5075 32.3125 12.5725 32.3775 ;
        RECT  12.5075 33.13 12.5725 33.195 ;
        RECT  12.5075 33.13 12.5725 33.195 ;
        RECT  12.5075 33.13 12.5725 33.195 ;
        RECT  12.5075 33.13 12.5725 33.195 ;
        RECT  12.5075 33.13 12.5725 33.195 ;
        RECT  12.5075 33.13 12.5725 33.195 ;
        RECT  12.5075 33.13 12.5725 33.195 ;
        RECT  12.5075 33.13 12.5725 33.195 ;
        RECT  12.0575 32.6375 12.1225 32.7025 ;
        RECT  11.8025 33.13 11.8675 33.195 ;
        RECT  11.8025 33.13 11.8675 33.195 ;
        RECT  11.8025 33.13 11.8675 33.195 ;
        RECT  11.8025 33.13 11.8675 33.195 ;
        RECT  11.8025 33.13 11.8675 33.195 ;
        RECT  11.8025 33.13 11.8675 33.195 ;
        RECT  12.5075 33.13 12.5725 33.195 ;
        RECT  12.5075 33.13 12.5725 33.195 ;
        RECT  12.5075 33.13 12.5725 33.195 ;
        RECT  12.5075 33.13 12.5725 33.195 ;
        RECT  12.2525 32.6375 12.3175 32.7025 ;
        RECT  12.5075 32.3125 12.5725 32.3775 ;
        RECT  12.5075 32.3125 12.5725 32.3775 ;
        RECT  12.5075 32.3125 12.5725 32.3775 ;
        RECT  12.5075 33.13 12.5725 33.195 ;
        RECT  12.5075 33.13 12.5725 33.195 ;
        RECT  12.5075 33.13 12.5725 33.195 ;
        RECT  12.5075 33.13 12.5725 33.195 ;
        RECT  12.5075 33.13 12.5725 33.195 ;
        RECT  12.5075 33.13 12.5725 33.195 ;
        RECT  11.8025 32.3125 11.8675 32.3775 ;
        RECT  12.5075 34.185 12.5725 34.25 ;
        RECT  12.5075 34.185 12.5725 34.25 ;
        RECT  12.5075 34.185 12.5725 34.25 ;
        RECT  12.5075 34.185 12.5725 34.25 ;
        RECT  12.5075 34.185 12.5725 34.25 ;
        RECT  12.5075 34.185 12.5725 34.25 ;
        RECT  11.8025 35.0025 11.8675 35.0675 ;
        RECT  12.5075 35.0025 12.5725 35.0675 ;
        RECT  12.5075 34.185 12.5725 34.25 ;
        RECT  12.5075 34.185 12.5725 34.25 ;
        RECT  12.5075 34.185 12.5725 34.25 ;
        RECT  12.5075 34.185 12.5725 34.25 ;
        RECT  12.5075 34.185 12.5725 34.25 ;
        RECT  12.5075 34.185 12.5725 34.25 ;
        RECT  12.5075 34.185 12.5725 34.25 ;
        RECT  12.5075 34.185 12.5725 34.25 ;
        RECT  12.0575 34.6775 12.1225 34.7425 ;
        RECT  11.8025 34.185 11.8675 34.25 ;
        RECT  11.8025 34.185 11.8675 34.25 ;
        RECT  11.8025 34.185 11.8675 34.25 ;
        RECT  11.8025 34.185 11.8675 34.25 ;
        RECT  11.8025 34.185 11.8675 34.25 ;
        RECT  11.8025 34.185 11.8675 34.25 ;
        RECT  12.5075 34.185 12.5725 34.25 ;
        RECT  12.5075 34.185 12.5725 34.25 ;
        RECT  12.5075 34.185 12.5725 34.25 ;
        RECT  12.5075 34.185 12.5725 34.25 ;
        RECT  12.2525 34.6775 12.3175 34.7425 ;
        RECT  12.5075 35.0025 12.5725 35.0675 ;
        RECT  12.5075 35.0025 12.5725 35.0675 ;
        RECT  12.5075 35.0025 12.5725 35.0675 ;
        RECT  12.5075 34.185 12.5725 34.25 ;
        RECT  12.5075 34.185 12.5725 34.25 ;
        RECT  12.5075 34.185 12.5725 34.25 ;
        RECT  12.5075 34.185 12.5725 34.25 ;
        RECT  12.5075 34.185 12.5725 34.25 ;
        RECT  12.5075 34.185 12.5725 34.25 ;
        RECT  11.8025 35.0025 11.8675 35.0675 ;
        RECT  12.5075 35.82 12.5725 35.885 ;
        RECT  12.5075 35.82 12.5725 35.885 ;
        RECT  12.5075 35.82 12.5725 35.885 ;
        RECT  12.5075 35.82 12.5725 35.885 ;
        RECT  12.5075 35.82 12.5725 35.885 ;
        RECT  12.5075 35.82 12.5725 35.885 ;
        RECT  11.8025 35.0025 11.8675 35.0675 ;
        RECT  12.5075 35.0025 12.5725 35.0675 ;
        RECT  12.5075 35.82 12.5725 35.885 ;
        RECT  12.5075 35.82 12.5725 35.885 ;
        RECT  12.5075 35.82 12.5725 35.885 ;
        RECT  12.5075 35.82 12.5725 35.885 ;
        RECT  12.5075 35.82 12.5725 35.885 ;
        RECT  12.5075 35.82 12.5725 35.885 ;
        RECT  12.5075 35.82 12.5725 35.885 ;
        RECT  12.5075 35.82 12.5725 35.885 ;
        RECT  12.0575 35.3275 12.1225 35.3925 ;
        RECT  11.8025 35.82 11.8675 35.885 ;
        RECT  11.8025 35.82 11.8675 35.885 ;
        RECT  11.8025 35.82 11.8675 35.885 ;
        RECT  11.8025 35.82 11.8675 35.885 ;
        RECT  11.8025 35.82 11.8675 35.885 ;
        RECT  11.8025 35.82 11.8675 35.885 ;
        RECT  12.5075 35.82 12.5725 35.885 ;
        RECT  12.5075 35.82 12.5725 35.885 ;
        RECT  12.5075 35.82 12.5725 35.885 ;
        RECT  12.5075 35.82 12.5725 35.885 ;
        RECT  12.2525 35.3275 12.3175 35.3925 ;
        RECT  12.5075 35.0025 12.5725 35.0675 ;
        RECT  12.5075 35.0025 12.5725 35.0675 ;
        RECT  12.5075 35.0025 12.5725 35.0675 ;
        RECT  12.5075 35.82 12.5725 35.885 ;
        RECT  12.5075 35.82 12.5725 35.885 ;
        RECT  12.5075 35.82 12.5725 35.885 ;
        RECT  12.5075 35.82 12.5725 35.885 ;
        RECT  12.5075 35.82 12.5725 35.885 ;
        RECT  12.5075 35.82 12.5725 35.885 ;
        RECT  11.8025 35.0025 11.8675 35.0675 ;
        RECT  12.5075 36.875 12.5725 36.94 ;
        RECT  12.5075 36.875 12.5725 36.94 ;
        RECT  12.5075 36.875 12.5725 36.94 ;
        RECT  12.5075 36.875 12.5725 36.94 ;
        RECT  12.5075 36.875 12.5725 36.94 ;
        RECT  12.5075 36.875 12.5725 36.94 ;
        RECT  11.8025 37.6925 11.8675 37.7575 ;
        RECT  12.5075 37.6925 12.5725 37.7575 ;
        RECT  12.5075 36.875 12.5725 36.94 ;
        RECT  12.5075 36.875 12.5725 36.94 ;
        RECT  12.5075 36.875 12.5725 36.94 ;
        RECT  12.5075 36.875 12.5725 36.94 ;
        RECT  12.5075 36.875 12.5725 36.94 ;
        RECT  12.5075 36.875 12.5725 36.94 ;
        RECT  12.5075 36.875 12.5725 36.94 ;
        RECT  12.5075 36.875 12.5725 36.94 ;
        RECT  12.0575 37.3675 12.1225 37.4325 ;
        RECT  11.8025 36.875 11.8675 36.94 ;
        RECT  11.8025 36.875 11.8675 36.94 ;
        RECT  11.8025 36.875 11.8675 36.94 ;
        RECT  11.8025 36.875 11.8675 36.94 ;
        RECT  11.8025 36.875 11.8675 36.94 ;
        RECT  11.8025 36.875 11.8675 36.94 ;
        RECT  12.5075 36.875 12.5725 36.94 ;
        RECT  12.5075 36.875 12.5725 36.94 ;
        RECT  12.5075 36.875 12.5725 36.94 ;
        RECT  12.5075 36.875 12.5725 36.94 ;
        RECT  12.2525 37.3675 12.3175 37.4325 ;
        RECT  12.5075 37.6925 12.5725 37.7575 ;
        RECT  12.5075 37.6925 12.5725 37.7575 ;
        RECT  12.5075 37.6925 12.5725 37.7575 ;
        RECT  12.5075 36.875 12.5725 36.94 ;
        RECT  12.5075 36.875 12.5725 36.94 ;
        RECT  12.5075 36.875 12.5725 36.94 ;
        RECT  12.5075 36.875 12.5725 36.94 ;
        RECT  12.5075 36.875 12.5725 36.94 ;
        RECT  12.5075 36.875 12.5725 36.94 ;
        RECT  11.8025 37.6925 11.8675 37.7575 ;
        RECT  12.5075 38.51 12.5725 38.575 ;
        RECT  12.5075 38.51 12.5725 38.575 ;
        RECT  12.5075 38.51 12.5725 38.575 ;
        RECT  12.5075 38.51 12.5725 38.575 ;
        RECT  12.5075 38.51 12.5725 38.575 ;
        RECT  12.5075 38.51 12.5725 38.575 ;
        RECT  11.8025 37.6925 11.8675 37.7575 ;
        RECT  12.5075 37.6925 12.5725 37.7575 ;
        RECT  12.5075 38.51 12.5725 38.575 ;
        RECT  12.5075 38.51 12.5725 38.575 ;
        RECT  12.5075 38.51 12.5725 38.575 ;
        RECT  12.5075 38.51 12.5725 38.575 ;
        RECT  12.5075 38.51 12.5725 38.575 ;
        RECT  12.5075 38.51 12.5725 38.575 ;
        RECT  12.5075 38.51 12.5725 38.575 ;
        RECT  12.5075 38.51 12.5725 38.575 ;
        RECT  12.0575 38.0175 12.1225 38.0825 ;
        RECT  11.8025 38.51 11.8675 38.575 ;
        RECT  11.8025 38.51 11.8675 38.575 ;
        RECT  11.8025 38.51 11.8675 38.575 ;
        RECT  11.8025 38.51 11.8675 38.575 ;
        RECT  11.8025 38.51 11.8675 38.575 ;
        RECT  11.8025 38.51 11.8675 38.575 ;
        RECT  12.5075 38.51 12.5725 38.575 ;
        RECT  12.5075 38.51 12.5725 38.575 ;
        RECT  12.5075 38.51 12.5725 38.575 ;
        RECT  12.5075 38.51 12.5725 38.575 ;
        RECT  12.2525 38.0175 12.3175 38.0825 ;
        RECT  12.5075 37.6925 12.5725 37.7575 ;
        RECT  12.5075 37.6925 12.5725 37.7575 ;
        RECT  12.5075 37.6925 12.5725 37.7575 ;
        RECT  12.5075 38.51 12.5725 38.575 ;
        RECT  12.5075 38.51 12.5725 38.575 ;
        RECT  12.5075 38.51 12.5725 38.575 ;
        RECT  12.5075 38.51 12.5725 38.575 ;
        RECT  12.5075 38.51 12.5725 38.575 ;
        RECT  12.5075 38.51 12.5725 38.575 ;
        RECT  11.8025 37.6925 11.8675 37.7575 ;
        RECT  12.5075 39.565 12.5725 39.63 ;
        RECT  12.5075 39.565 12.5725 39.63 ;
        RECT  12.5075 39.565 12.5725 39.63 ;
        RECT  12.5075 39.565 12.5725 39.63 ;
        RECT  12.5075 39.565 12.5725 39.63 ;
        RECT  12.5075 39.565 12.5725 39.63 ;
        RECT  11.8025 40.3825 11.8675 40.4475 ;
        RECT  12.5075 40.3825 12.5725 40.4475 ;
        RECT  12.5075 39.565 12.5725 39.63 ;
        RECT  12.5075 39.565 12.5725 39.63 ;
        RECT  12.5075 39.565 12.5725 39.63 ;
        RECT  12.5075 39.565 12.5725 39.63 ;
        RECT  12.5075 39.565 12.5725 39.63 ;
        RECT  12.5075 39.565 12.5725 39.63 ;
        RECT  12.5075 39.565 12.5725 39.63 ;
        RECT  12.5075 39.565 12.5725 39.63 ;
        RECT  12.0575 40.0575 12.1225 40.1225 ;
        RECT  11.8025 39.565 11.8675 39.63 ;
        RECT  11.8025 39.565 11.8675 39.63 ;
        RECT  11.8025 39.565 11.8675 39.63 ;
        RECT  11.8025 39.565 11.8675 39.63 ;
        RECT  11.8025 39.565 11.8675 39.63 ;
        RECT  11.8025 39.565 11.8675 39.63 ;
        RECT  12.5075 39.565 12.5725 39.63 ;
        RECT  12.5075 39.565 12.5725 39.63 ;
        RECT  12.5075 39.565 12.5725 39.63 ;
        RECT  12.5075 39.565 12.5725 39.63 ;
        RECT  12.2525 40.0575 12.3175 40.1225 ;
        RECT  12.5075 40.3825 12.5725 40.4475 ;
        RECT  12.5075 40.3825 12.5725 40.4475 ;
        RECT  12.5075 40.3825 12.5725 40.4475 ;
        RECT  12.5075 39.565 12.5725 39.63 ;
        RECT  12.5075 39.565 12.5725 39.63 ;
        RECT  12.5075 39.565 12.5725 39.63 ;
        RECT  12.5075 39.565 12.5725 39.63 ;
        RECT  12.5075 39.565 12.5725 39.63 ;
        RECT  12.5075 39.565 12.5725 39.63 ;
        RECT  11.8025 40.3825 11.8675 40.4475 ;
        RECT  11.325 41.3475 11.39 41.4125 ;
        RECT  11.705 41.3475 11.77 41.4125 ;
        RECT  11.325 40.8975 11.39 40.9625 ;
        RECT  11.515 40.8975 11.58 40.9625 ;
        RECT  12.03 41.3475 12.095 41.4125 ;
        RECT  12.41 41.3475 12.475 41.4125 ;
        RECT  12.03 40.8975 12.095 40.9625 ;
        RECT  12.22 40.8975 12.285 40.9625 ;
        RECT  11.445 18.5325 11.51 18.5975 ;
        RECT  11.8025 14.2925 11.8675 14.3575 ;
        RECT  11.0975 14.2925 11.1625 14.3575 ;
        RECT  11.64 17.075 11.705 17.14 ;
        RECT  11.2575 17.485 11.3225 17.55 ;
        RECT  11.45 18.3275 11.515 18.3925 ;
        RECT  11.45 16.185 11.515 16.25 ;
        RECT  12.15 18.5325 12.215 18.5975 ;
        RECT  12.5075 14.2925 12.5725 14.3575 ;
        RECT  11.8025 14.2925 11.8675 14.3575 ;
        RECT  12.345 17.075 12.41 17.14 ;
        RECT  11.9625 17.485 12.0275 17.55 ;
        RECT  12.155 18.3275 12.22 18.3925 ;
        RECT  12.155 16.185 12.22 16.25 ;
        RECT  11.3725 9.97 11.4375 10.035 ;
        RECT  11.8025 11.605 11.8675 11.67 ;
        RECT  11.8025 11.035 11.8675 11.1 ;
        RECT  11.0975 11.035 11.1625 11.1 ;
        RECT  11.5175 11.24 11.5825 11.305 ;
        RECT  11.8025 13.5325 11.8675 13.5975 ;
        RECT  11.5175 10.83 11.5825 10.895 ;
        RECT  11.3775 10.83 11.4425 10.895 ;
        RECT  11.8025 11.24 11.8675 11.305 ;
        RECT  11.0975 11.24 11.1625 11.305 ;
        RECT  11.27 10.2325 11.335 10.2975 ;
        RECT  11.3775 13.21 11.4425 13.275 ;
        RECT  11.5475 11.605 11.6125 11.67 ;
        RECT  11.2375 12.52 11.3025 12.585 ;
        RECT  11.3775 11.24 11.4425 11.305 ;
        RECT  11.0975 11.605 11.1625 11.67 ;
        RECT  11.5475 12.12 11.6125 12.185 ;
        RECT  11.2825 13.7425 11.3475 13.8075 ;
        RECT  11.0975 13.5325 11.1625 13.5975 ;
        RECT  12.0775 9.97 12.1425 10.035 ;
        RECT  12.5075 11.605 12.5725 11.67 ;
        RECT  12.5075 11.035 12.5725 11.1 ;
        RECT  11.8025 11.035 11.8675 11.1 ;
        RECT  12.2225 11.24 12.2875 11.305 ;
        RECT  12.5075 13.5325 12.5725 13.5975 ;
        RECT  12.2225 10.83 12.2875 10.895 ;
        RECT  12.0825 10.83 12.1475 10.895 ;
        RECT  12.5075 11.24 12.5725 11.305 ;
        RECT  11.8025 11.24 11.8675 11.305 ;
        RECT  11.975 10.2325 12.04 10.2975 ;
        RECT  12.0825 13.21 12.1475 13.275 ;
        RECT  12.2525 11.605 12.3175 11.67 ;
        RECT  11.9425 12.52 12.0075 12.585 ;
        RECT  12.0825 11.24 12.1475 11.305 ;
        RECT  11.8025 11.605 11.8675 11.67 ;
        RECT  12.2525 12.12 12.3175 12.185 ;
        RECT  11.9875 13.7425 12.0525 13.8075 ;
        RECT  11.8025 13.5325 11.8675 13.5975 ;
        RECT  11.295 9.1325 11.36 9.1975 ;
        RECT  11.8025 3.955 11.8675 4.02 ;
        RECT  11.66 8.0375 11.725 8.1025 ;
        RECT  11.6625 6.43 11.7275 6.495 ;
        RECT  11.6625 5.0325 11.7275 5.0975 ;
        RECT  11.0975 3.815 11.1625 3.88 ;
        RECT  11.8025 6.8925 11.8675 6.9575 ;
        RECT  11.2975 5.6975 11.3625 5.7625 ;
        RECT  11.6625 9.39 11.7275 9.455 ;
        RECT  11.485 8.88 11.55 8.945 ;
        RECT  11.8025 8.4675 11.8675 8.5325 ;
        RECT  11.8025 3.765 11.8675 3.83 ;
        RECT  11.8025 5.5075 11.8675 5.5725 ;
        RECT  11.2975 5.3075 11.3625 5.3725 ;
        RECT  11.485 5.3075 11.55 5.3725 ;
        RECT  11.485 5.92 11.55 5.985 ;
        RECT  11.295 8.2675 11.36 8.3325 ;
        RECT  11.485 8.2675 11.55 8.3325 ;
        RECT  12.31 9.1325 12.375 9.1975 ;
        RECT  11.8025 3.955 11.8675 4.02 ;
        RECT  11.945 8.0375 12.01 8.1025 ;
        RECT  11.9425 6.43 12.0075 6.495 ;
        RECT  11.9425 5.0325 12.0075 5.0975 ;
        RECT  12.5075 3.815 12.5725 3.88 ;
        RECT  11.8025 6.8925 11.8675 6.9575 ;
        RECT  12.3075 5.6975 12.3725 5.7625 ;
        RECT  11.9425 9.39 12.0075 9.455 ;
        RECT  12.12 8.88 12.185 8.945 ;
        RECT  11.8025 8.4675 11.8675 8.5325 ;
        RECT  11.8025 3.765 11.8675 3.83 ;
        RECT  11.8025 5.5075 11.8675 5.5725 ;
        RECT  12.3075 5.3075 12.3725 5.3725 ;
        RECT  12.12 5.3075 12.185 5.3725 ;
        RECT  12.12 5.92 12.185 5.985 ;
        RECT  12.31 8.2675 12.375 8.3325 ;
        RECT  12.12 8.2675 12.185 8.3325 ;
        RECT  11.45 5.18 11.515 5.245 ;
        RECT  11.8025 3.9275 11.8675 3.9925 ;
        RECT  11.5825 5.82 11.6475 5.885 ;
        RECT  11.8025 5.9875 11.8675 6.0525 ;
        RECT  11.275 5.7975 11.34 5.8625 ;
        RECT  11.4825 5.52 11.5475 5.585 ;
        RECT  11.5825 4.3125 11.6475 4.3775 ;
        RECT  11.2375 4.08 11.3025 4.145 ;
        RECT  12.155 5.18 12.22 5.245 ;
        RECT  11.8025 3.9275 11.8675 3.9925 ;
        RECT  12.0225 5.82 12.0875 5.885 ;
        RECT  11.8025 5.9875 11.8675 6.0525 ;
        RECT  12.33 5.7975 12.395 5.8625 ;
        RECT  12.1225 5.52 12.1875 5.585 ;
        RECT  12.0225 4.3125 12.0875 4.3775 ;
        RECT  12.3675 4.08 12.4325 4.145 ;
        RECT  6.16 9.1825 6.225 9.2475 ;
        RECT  7.525 8.66 7.59 8.725 ;
        RECT  5.985 9.5725 6.05 9.6375 ;
        RECT  7.35 10.095 7.415 10.16 ;
        RECT  6.16 8.975 6.225 9.04 ;
        RECT  5.985 8.445 6.05 8.51 ;
        RECT  5.81 9.78 5.875 9.845 ;
        RECT  5.985 10.31 6.05 10.375 ;
        RECT  6.16 11.665 6.225 11.73 ;
        RECT  5.635 11.135 5.7 11.2 ;
        RECT  5.81 12.47 5.875 12.535 ;
        RECT  7.525 12.47 7.59 12.535 ;
        RECT  5.635 13.0 5.7 13.065 ;
        RECT  7.35 13.0 7.415 13.065 ;
        RECT  6.335 8.0325 6.4 8.0975 ;
        RECT  6.51 9.3775 6.575 9.4425 ;
        RECT  6.335 10.7225 6.4 10.7875 ;
        RECT  6.51 12.0675 6.575 12.1325 ;
        RECT  6.335 13.235 6.4 13.3 ;
        RECT  6.16 14.5625 6.225 14.6275 ;
        RECT  7.525 14.04 7.59 14.105 ;
        RECT  5.985 14.9525 6.05 15.0175 ;
        RECT  7.35 15.475 7.415 15.54 ;
        RECT  6.16 14.355 6.225 14.42 ;
        RECT  5.985 13.825 6.05 13.89 ;
        RECT  5.81 15.16 5.875 15.225 ;
        RECT  5.985 15.69 6.05 15.755 ;
        RECT  6.16 17.045 6.225 17.11 ;
        RECT  5.635 16.515 5.7 16.58 ;
        RECT  5.81 17.85 5.875 17.915 ;
        RECT  7.525 17.85 7.59 17.915 ;
        RECT  5.635 18.38 5.7 18.445 ;
        RECT  7.35 18.38 7.415 18.445 ;
        RECT  6.335 13.4125 6.4 13.4775 ;
        RECT  6.51 14.7575 6.575 14.8225 ;
        RECT  6.335 16.1025 6.4 16.1675 ;
        RECT  6.51 17.4475 6.575 17.5125 ;
        RECT  6.335 18.615 6.4 18.68 ;
        RECT  2.825 8.73 2.89 8.795 ;
        RECT  3.0 10.165 3.065 10.23 ;
        RECT  3.175 11.42 3.24 11.485 ;
        RECT  3.35 12.855 3.415 12.92 ;
        RECT  3.525 14.11 3.59 14.175 ;
        RECT  3.7 15.545 3.765 15.61 ;
        RECT  3.875 16.8 3.94 16.865 ;
        RECT  4.05 18.235 4.115 18.3 ;
        RECT  2.825 19.805 2.89 19.87 ;
        RECT  3.525 19.275 3.59 19.34 ;
        RECT  2.825 20.61 2.89 20.675 ;
        RECT  3.7 21.14 3.765 21.205 ;
        RECT  2.825 22.495 2.89 22.56 ;
        RECT  3.875 21.965 3.94 22.03 ;
        RECT  2.825 23.3 2.89 23.365 ;
        RECT  4.05 23.83 4.115 23.895 ;
        RECT  3.0 25.185 3.065 25.25 ;
        RECT  3.525 24.655 3.59 24.72 ;
        RECT  3.0 25.99 3.065 26.055 ;
        RECT  3.7 26.52 3.765 26.585 ;
        RECT  3.0 27.875 3.065 27.94 ;
        RECT  3.875 27.345 3.94 27.41 ;
        RECT  3.0 28.68 3.065 28.745 ;
        RECT  4.05 29.21 4.115 29.275 ;
        RECT  3.175 30.565 3.24 30.63 ;
        RECT  3.525 30.035 3.59 30.1 ;
        RECT  3.175 31.37 3.24 31.435 ;
        RECT  3.7 31.9 3.765 31.965 ;
        RECT  3.175 33.255 3.24 33.32 ;
        RECT  3.875 32.725 3.94 32.79 ;
        RECT  3.175 34.06 3.24 34.125 ;
        RECT  4.05 34.59 4.115 34.655 ;
        RECT  3.35 35.945 3.415 36.01 ;
        RECT  3.525 35.415 3.59 35.48 ;
        RECT  3.35 36.75 3.415 36.815 ;
        RECT  3.7 37.28 3.765 37.345 ;
        RECT  3.35 38.635 3.415 38.7 ;
        RECT  3.875 38.105 3.94 38.17 ;
        RECT  3.35 39.44 3.415 39.505 ;
        RECT  4.05 39.97 4.115 40.035 ;
        RECT  5.495 20.2075 5.56 20.2725 ;
        RECT  5.95 20.2075 6.015 20.2725 ;
        RECT  6.58 19.8075 6.645 19.8725 ;
        RECT  5.5325 19.84 5.5975 19.905 ;
        RECT  5.495 21.5525 5.56 21.6175 ;
        RECT  5.95 21.5525 6.015 21.6175 ;
        RECT  6.58 20.6075 6.645 20.6725 ;
        RECT  5.5325 20.575 5.5975 20.64 ;
        RECT  5.495 22.8975 5.56 22.9625 ;
        RECT  5.95 22.8975 6.015 22.9625 ;
        RECT  6.58 22.4975 6.645 22.5625 ;
        RECT  5.5325 22.53 5.5975 22.595 ;
        RECT  5.495 24.2425 5.56 24.3075 ;
        RECT  5.95 24.2425 6.015 24.3075 ;
        RECT  6.58 23.2975 6.645 23.3625 ;
        RECT  5.5325 23.265 5.5975 23.33 ;
        RECT  5.495 25.5875 5.56 25.6525 ;
        RECT  5.95 25.5875 6.015 25.6525 ;
        RECT  6.58 25.1875 6.645 25.2525 ;
        RECT  5.5325 25.22 5.5975 25.285 ;
        RECT  5.495 26.9325 5.56 26.9975 ;
        RECT  5.95 26.9325 6.015 26.9975 ;
        RECT  6.58 25.9875 6.645 26.0525 ;
        RECT  5.5325 25.955 5.5975 26.02 ;
        RECT  5.495 28.2775 5.56 28.3425 ;
        RECT  5.95 28.2775 6.015 28.3425 ;
        RECT  6.58 27.8775 6.645 27.9425 ;
        RECT  5.5325 27.91 5.5975 27.975 ;
        RECT  5.495 29.6225 5.56 29.6875 ;
        RECT  5.95 29.6225 6.015 29.6875 ;
        RECT  6.58 28.6775 6.645 28.7425 ;
        RECT  5.5325 28.645 5.5975 28.71 ;
        RECT  5.495 30.9675 5.56 31.0325 ;
        RECT  5.95 30.9675 6.015 31.0325 ;
        RECT  6.58 30.5675 6.645 30.6325 ;
        RECT  5.5325 30.6 5.5975 30.665 ;
        RECT  5.495 32.3125 5.56 32.3775 ;
        RECT  5.95 32.3125 6.015 32.3775 ;
        RECT  6.58 31.3675 6.645 31.4325 ;
        RECT  5.5325 31.335 5.5975 31.4 ;
        RECT  5.495 33.6575 5.56 33.7225 ;
        RECT  5.95 33.6575 6.015 33.7225 ;
        RECT  6.58 33.2575 6.645 33.3225 ;
        RECT  5.5325 33.29 5.5975 33.355 ;
        RECT  5.495 35.0025 5.56 35.0675 ;
        RECT  5.95 35.0025 6.015 35.0675 ;
        RECT  6.58 34.0575 6.645 34.1225 ;
        RECT  5.5325 34.025 5.5975 34.09 ;
        RECT  5.495 36.3475 5.56 36.4125 ;
        RECT  5.95 36.3475 6.015 36.4125 ;
        RECT  6.58 35.9475 6.645 36.0125 ;
        RECT  5.5325 35.98 5.5975 36.045 ;
        RECT  5.495 37.6925 5.56 37.7575 ;
        RECT  5.95 37.6925 6.015 37.7575 ;
        RECT  6.58 36.7475 6.645 36.8125 ;
        RECT  5.5325 36.715 5.5975 36.78 ;
        RECT  5.495 39.0375 5.56 39.1025 ;
        RECT  5.95 39.0375 6.015 39.1025 ;
        RECT  6.58 38.6375 6.645 38.7025 ;
        RECT  5.5325 38.67 5.5975 38.735 ;
        RECT  5.495 40.3825 5.56 40.4475 ;
        RECT  5.95 40.3825 6.015 40.4475 ;
        RECT  6.58 39.4375 6.645 39.5025 ;
        RECT  5.5325 39.405 5.5975 39.47 ;
        RECT  6.6475 7.61 6.7125 7.675 ;
        RECT  1.47 7.1025 1.535 7.1675 ;
        RECT  5.5525 7.245 5.6175 7.31 ;
        RECT  3.945 7.2425 4.01 7.3075 ;
        RECT  2.5475 7.2425 2.6125 7.3075 ;
        RECT  1.33 7.8075 1.395 7.8725 ;
        RECT  4.4075 7.1025 4.4725 7.1675 ;
        RECT  3.2125 7.6075 3.2775 7.6725 ;
        RECT  6.905 7.2425 6.97 7.3075 ;
        RECT  6.395 7.42 6.46 7.485 ;
        RECT  5.9825 7.1025 6.0475 7.1675 ;
        RECT  1.28 7.1025 1.345 7.1675 ;
        RECT  3.0225 7.1025 3.0875 7.1675 ;
        RECT  2.8225 7.6075 2.8875 7.6725 ;
        RECT  2.8225 7.42 2.8875 7.485 ;
        RECT  3.435 7.42 3.5 7.485 ;
        RECT  5.7825 7.61 5.8475 7.675 ;
        RECT  5.7825 7.42 5.8475 7.485 ;
        RECT  6.6475 6.595 6.7125 6.66 ;
        RECT  1.47 7.1025 1.535 7.1675 ;
        RECT  5.5525 6.96 5.6175 7.025 ;
        RECT  3.945 6.9625 4.01 7.0275 ;
        RECT  2.5475 6.9625 2.6125 7.0275 ;
        RECT  1.33 6.3975 1.395 6.4625 ;
        RECT  4.4075 7.1025 4.4725 7.1675 ;
        RECT  3.2125 6.5975 3.2775 6.6625 ;
        RECT  6.905 6.9625 6.97 7.0275 ;
        RECT  6.395 6.785 6.46 6.85 ;
        RECT  5.9825 7.1025 6.0475 7.1675 ;
        RECT  1.28 7.1025 1.345 7.1675 ;
        RECT  3.0225 7.1025 3.0875 7.1675 ;
        RECT  2.8225 6.5975 2.8875 6.6625 ;
        RECT  2.8225 6.785 2.8875 6.85 ;
        RECT  3.435 6.785 3.5 6.85 ;
        RECT  5.7825 6.595 5.8475 6.66 ;
        RECT  5.7825 6.785 5.8475 6.85 ;
        RECT  6.6475 6.2 6.7125 6.265 ;
        RECT  1.47 5.6925 1.535 5.7575 ;
        RECT  5.5525 5.835 5.6175 5.9 ;
        RECT  3.945 5.8325 4.01 5.8975 ;
        RECT  2.5475 5.8325 2.6125 5.8975 ;
        RECT  1.33 6.3975 1.395 6.4625 ;
        RECT  4.4075 5.6925 4.4725 5.7575 ;
        RECT  3.2125 6.1975 3.2775 6.2625 ;
        RECT  6.905 5.8325 6.97 5.8975 ;
        RECT  6.395 6.01 6.46 6.075 ;
        RECT  5.9825 5.6925 6.0475 5.7575 ;
        RECT  1.28 5.6925 1.345 5.7575 ;
        RECT  3.0225 5.6925 3.0875 5.7575 ;
        RECT  2.8225 6.1975 2.8875 6.2625 ;
        RECT  2.8225 6.01 2.8875 6.075 ;
        RECT  3.435 6.01 3.5 6.075 ;
        RECT  5.7825 6.2 5.8475 6.265 ;
        RECT  5.7825 6.01 5.8475 6.075 ;
        RECT  6.6475 5.185 6.7125 5.25 ;
        RECT  1.47 5.6925 1.535 5.7575 ;
        RECT  5.5525 5.55 5.6175 5.615 ;
        RECT  3.945 5.5525 4.01 5.6175 ;
        RECT  2.5475 5.5525 2.6125 5.6175 ;
        RECT  1.33 4.9875 1.395 5.0525 ;
        RECT  4.4075 5.6925 4.4725 5.7575 ;
        RECT  3.2125 5.1875 3.2775 5.2525 ;
        RECT  6.905 5.5525 6.97 5.6175 ;
        RECT  6.395 5.375 6.46 5.44 ;
        RECT  5.9825 5.6925 6.0475 5.7575 ;
        RECT  1.28 5.6925 1.345 5.7575 ;
        RECT  3.0225 5.6925 3.0875 5.7575 ;
        RECT  2.8225 5.1875 2.8875 5.2525 ;
        RECT  2.8225 5.375 2.8875 5.44 ;
        RECT  3.435 5.375 3.5 5.44 ;
        RECT  5.7825 5.185 5.8475 5.25 ;
        RECT  5.7825 5.375 5.8475 5.44 ;
        RECT  8.5425 8.765 8.6075 8.83 ;
        RECT  8.3325 10.2 8.3975 10.265 ;
        RECT  8.1225 14.145 8.1875 14.21 ;
        RECT  7.9125 15.58 7.9775 15.645 ;
        RECT  10.3625 3.635 10.4275 3.7 ;
        RECT  9.9425 1.45 10.0075 1.515 ;
        RECT  10.1525 2.9975 10.2175 3.0625 ;
        RECT  10.3625 41.135 10.4275 41.2 ;
        RECT  10.5725 10.1375 10.6375 10.2025 ;
        RECT  10.7825 14.1625 10.8475 14.2275 ;
        RECT  1.015 7.63 1.08 7.695 ;
        RECT  9.7325 41.565 9.7975 41.63 ;
        RECT  8.89 40.58 8.955 40.645 ;
        RECT  9.03 40.58 9.095 40.645 ;
        RECT  11.805 40.5475 11.87 40.6125 ;
        RECT  12.51 40.5475 12.575 40.6125 ;
        RECT  11.03 40.5475 11.095 40.6125 ;
        RECT  9.385 0.39 9.45 0.455 ;
        RECT  9.525 0.39 9.59 0.455 ;
        RECT  11.8025 0.39 11.8675 0.455 ;
        RECT  11.8025 0.39 11.8675 0.455 ;
        RECT  7.79 21.555 7.855 21.62 ;
        RECT  7.79 24.245 7.855 24.31 ;
        RECT  7.79 26.935 7.855 27.0 ;
        RECT  7.79 29.625 7.855 29.69 ;
        RECT  7.79 32.315 7.855 32.38 ;
        RECT  7.79 35.005 7.855 35.07 ;
        RECT  7.79 37.695 7.855 37.76 ;
        RECT  7.79 40.385 7.855 40.45 ;
        RECT  8.89 13.4475 8.955 13.5125 ;
        RECT  9.03 13.4475 9.095 13.5125 ;
        RECT  8.89 18.8275 8.955 18.8925 ;
        RECT  9.03 18.8275 9.095 18.8925 ;
        RECT  7.315 7.81 7.38 7.875 ;
        RECT  8.89 7.8425 8.955 7.9075 ;
        RECT  9.03 7.8425 9.095 7.9075 ;
        RECT  7.315 6.4 7.38 6.465 ;
        RECT  8.89 6.4325 8.955 6.4975 ;
        RECT  9.03 6.4325 9.095 6.4975 ;
        RECT  7.315 6.4 7.38 6.465 ;
        RECT  8.89 6.4325 8.955 6.4975 ;
        RECT  9.03 6.4325 9.095 6.4975 ;
        RECT  7.315 4.99 7.38 5.055 ;
        RECT  8.89 5.0225 8.955 5.0875 ;
        RECT  9.03 5.0225 9.095 5.0875 ;
        RECT  -5.565 14.0125 -5.5 14.0775 ;
        RECT  -5.0575 8.835 -4.9925 8.9 ;
        RECT  -5.2 12.9175 -5.135 12.9825 ;
        RECT  -5.1975 11.31 -5.1325 11.375 ;
        RECT  -5.1975 9.9125 -5.1325 9.9775 ;
        RECT  -5.7625 8.695 -5.6975 8.76 ;
        RECT  -5.0575 11.7725 -4.9925 11.8375 ;
        RECT  -5.5625 10.5775 -5.4975 10.6425 ;
        RECT  -5.1975 14.27 -5.1325 14.335 ;
        RECT  -5.375 13.76 -5.31 13.825 ;
        RECT  -5.0575 13.3475 -4.9925 13.4125 ;
        RECT  -5.0575 8.645 -4.9925 8.71 ;
        RECT  -5.0575 10.3875 -4.9925 10.4525 ;
        RECT  -5.5625 10.1875 -5.4975 10.2525 ;
        RECT  -5.375 10.1875 -5.31 10.2525 ;
        RECT  -5.375 10.8 -5.31 10.865 ;
        RECT  -5.565 13.1475 -5.5 13.2125 ;
        RECT  -5.375 13.1475 -5.31 13.2125 ;
        RECT  -4.55 14.0125 -4.485 14.0775 ;
        RECT  -5.0575 8.835 -4.9925 8.9 ;
        RECT  -4.915 12.9175 -4.85 12.9825 ;
        RECT  -4.9175 11.31 -4.8525 11.375 ;
        RECT  -4.9175 9.9125 -4.8525 9.9775 ;
        RECT  -4.3525 8.695 -4.2875 8.76 ;
        RECT  -5.0575 11.7725 -4.9925 11.8375 ;
        RECT  -4.5525 10.5775 -4.4875 10.6425 ;
        RECT  -4.9175 14.27 -4.8525 14.335 ;
        RECT  -4.74 13.76 -4.675 13.825 ;
        RECT  -5.0575 13.3475 -4.9925 13.4125 ;
        RECT  -5.0575 8.645 -4.9925 8.71 ;
        RECT  -5.0575 10.3875 -4.9925 10.4525 ;
        RECT  -4.5525 10.1875 -4.4875 10.2525 ;
        RECT  -4.74 10.1875 -4.675 10.2525 ;
        RECT  -4.74 10.8 -4.675 10.865 ;
        RECT  -4.55 13.1475 -4.485 13.2125 ;
        RECT  -4.74 13.1475 -4.675 13.2125 ;
        RECT  -4.155 14.0125 -4.09 14.0775 ;
        RECT  -3.6475 8.835 -3.5825 8.9 ;
        RECT  -3.79 12.9175 -3.725 12.9825 ;
        RECT  -3.7875 11.31 -3.7225 11.375 ;
        RECT  -3.7875 9.9125 -3.7225 9.9775 ;
        RECT  -4.3525 8.695 -4.2875 8.76 ;
        RECT  -3.6475 11.7725 -3.5825 11.8375 ;
        RECT  -4.1525 10.5775 -4.0875 10.6425 ;
        RECT  -3.7875 14.27 -3.7225 14.335 ;
        RECT  -3.965 13.76 -3.9 13.825 ;
        RECT  -3.6475 13.3475 -3.5825 13.4125 ;
        RECT  -3.6475 8.645 -3.5825 8.71 ;
        RECT  -3.6475 10.3875 -3.5825 10.4525 ;
        RECT  -4.1525 10.1875 -4.0875 10.2525 ;
        RECT  -3.965 10.1875 -3.9 10.2525 ;
        RECT  -3.965 10.8 -3.9 10.865 ;
        RECT  -4.155 13.1475 -4.09 13.2125 ;
        RECT  -3.965 13.1475 -3.9 13.2125 ;
        RECT  -1.3775 8.8425 -1.3125 8.9075 ;
        RECT  -0.8675 8.8425 -0.8025 8.9075 ;
        RECT  -1.0 23.83 -0.935 23.895 ;
        RECT  -1.0 23.27 -0.935 23.335 ;
        RECT  -2.52 22.845 -2.455 22.91 ;
        RECT  -2.52 23.405 -2.455 23.47 ;
        RECT  -1.0 23.5075 -0.935 23.5725 ;
        RECT  -1.0 22.9475 -0.935 23.0125 ;
        RECT  -2.52 23.1675 -2.455 23.2325 ;
        RECT  -4.225 23.0375 -4.16 23.1025 ;
        RECT  -4.93 23.5125 -4.865 23.5775 ;
        RECT  -4.225 23.5125 -4.16 23.5775 ;
        RECT  -4.6775 23.0325 -4.6125 23.0975 ;
        RECT  -4.4775 23.0375 -4.4125 23.1025 ;
        RECT  -4.93 22.7075 -4.865 22.7725 ;
        RECT  -4.225 22.7075 -4.16 22.7725 ;
        RECT  -4.93 21.89 -4.865 21.955 ;
        RECT  -4.93 21.89 -4.865 21.955 ;
        RECT  -4.93 21.89 -4.865 21.955 ;
        RECT  -4.93 21.89 -4.865 21.955 ;
        RECT  -4.93 21.89 -4.865 21.955 ;
        RECT  -4.93 21.89 -4.865 21.955 ;
        RECT  -4.225 22.7075 -4.16 22.7725 ;
        RECT  -4.93 22.7075 -4.865 22.7725 ;
        RECT  -4.93 21.89 -4.865 21.955 ;
        RECT  -4.93 21.89 -4.865 21.955 ;
        RECT  -4.93 21.89 -4.865 21.955 ;
        RECT  -4.93 21.89 -4.865 21.955 ;
        RECT  -4.93 21.89 -4.865 21.955 ;
        RECT  -4.93 21.89 -4.865 21.955 ;
        RECT  -4.93 21.89 -4.865 21.955 ;
        RECT  -4.93 21.89 -4.865 21.955 ;
        RECT  -4.48 22.3825 -4.415 22.4475 ;
        RECT  -4.225 21.89 -4.16 21.955 ;
        RECT  -4.225 21.89 -4.16 21.955 ;
        RECT  -4.225 21.89 -4.16 21.955 ;
        RECT  -4.225 21.89 -4.16 21.955 ;
        RECT  -4.225 21.89 -4.16 21.955 ;
        RECT  -4.225 21.89 -4.16 21.955 ;
        RECT  -4.93 21.89 -4.865 21.955 ;
        RECT  -4.93 21.89 -4.865 21.955 ;
        RECT  -4.93 21.89 -4.865 21.955 ;
        RECT  -4.93 21.89 -4.865 21.955 ;
        RECT  -4.675 22.3825 -4.61 22.4475 ;
        RECT  -4.93 22.7075 -4.865 22.7725 ;
        RECT  -4.93 22.7075 -4.865 22.7725 ;
        RECT  -4.93 22.7075 -4.865 22.7725 ;
        RECT  -4.93 21.89 -4.865 21.955 ;
        RECT  -4.93 21.89 -4.865 21.955 ;
        RECT  -4.93 21.89 -4.865 21.955 ;
        RECT  -4.93 21.89 -4.865 21.955 ;
        RECT  -4.93 21.89 -4.865 21.955 ;
        RECT  -4.93 21.89 -4.865 21.955 ;
        RECT  -4.225 22.7075 -4.16 22.7725 ;
        RECT  -4.93 20.835 -4.865 20.9 ;
        RECT  -4.93 20.835 -4.865 20.9 ;
        RECT  -4.93 20.835 -4.865 20.9 ;
        RECT  -4.93 20.835 -4.865 20.9 ;
        RECT  -4.93 20.835 -4.865 20.9 ;
        RECT  -4.93 20.835 -4.865 20.9 ;
        RECT  -4.225 20.0175 -4.16 20.0825 ;
        RECT  -4.93 20.0175 -4.865 20.0825 ;
        RECT  -4.93 20.835 -4.865 20.9 ;
        RECT  -4.93 20.835 -4.865 20.9 ;
        RECT  -4.93 20.835 -4.865 20.9 ;
        RECT  -4.93 20.835 -4.865 20.9 ;
        RECT  -4.93 20.835 -4.865 20.9 ;
        RECT  -4.93 20.835 -4.865 20.9 ;
        RECT  -4.93 20.835 -4.865 20.9 ;
        RECT  -4.93 20.835 -4.865 20.9 ;
        RECT  -4.48 20.3425 -4.415 20.4075 ;
        RECT  -4.225 20.835 -4.16 20.9 ;
        RECT  -4.225 20.835 -4.16 20.9 ;
        RECT  -4.225 20.835 -4.16 20.9 ;
        RECT  -4.225 20.835 -4.16 20.9 ;
        RECT  -4.225 20.835 -4.16 20.9 ;
        RECT  -4.225 20.835 -4.16 20.9 ;
        RECT  -4.93 20.835 -4.865 20.9 ;
        RECT  -4.93 20.835 -4.865 20.9 ;
        RECT  -4.93 20.835 -4.865 20.9 ;
        RECT  -4.93 20.835 -4.865 20.9 ;
        RECT  -4.675 20.3425 -4.61 20.4075 ;
        RECT  -4.93 20.0175 -4.865 20.0825 ;
        RECT  -4.93 20.0175 -4.865 20.0825 ;
        RECT  -4.93 20.0175 -4.865 20.0825 ;
        RECT  -4.93 20.835 -4.865 20.9 ;
        RECT  -4.93 20.835 -4.865 20.9 ;
        RECT  -4.93 20.835 -4.865 20.9 ;
        RECT  -4.93 20.835 -4.865 20.9 ;
        RECT  -4.93 20.835 -4.865 20.9 ;
        RECT  -4.93 20.835 -4.865 20.9 ;
        RECT  -4.225 20.0175 -4.16 20.0825 ;
        RECT  -1.975 21.1775 -1.91 21.2425 ;
        RECT  -1.38 21.385 -1.315 21.45 ;
        RECT  -2.135 21.385 -2.07 21.45 ;
        RECT  -4.41 24.28 -4.345 24.345 ;
        RECT  -0.6475 19.52 -0.5825 19.585 ;
        RECT  -2.555 19.5225 -2.49 19.5875 ;
        RECT  -2.59 24.2025 -2.525 24.2675 ;
        RECT  -0.6475 21.365 -0.5825 21.43 ;
        RECT  -4.025 22.4325 -3.96 22.4975 ;
        RECT  -3.735 22.0075 -3.67 22.0725 ;
        RECT  -3.735 23.7675 -3.67 23.8325 ;
        RECT  -0.415 20.6625 -0.35 20.7275 ;
        RECT  -0.415 16.165 -0.35 16.23 ;
        RECT  -3.105 16.1675 -3.04 16.2325 ;
        RECT  -3.77 26.2675 -3.705 26.3325 ;
        RECT  -3.525 23.93 -3.46 23.995 ;
        RECT  -3.525 25.01 -3.46 25.075 ;
        RECT  -3.735 28.345 -3.67 28.41 ;
        RECT  -3.525 23.93 -3.46 23.995 ;
        RECT  -3.525 22.6 -3.46 22.665 ;
        RECT  -3.735 31.035 -3.67 31.1 ;
        RECT  -4.93 20.6625 -4.865 20.7275 ;
        RECT  -4.225 20.6625 -4.16 20.7275 ;
        RECT  -2.0775 16.6075 -2.0125 16.6725 ;
        RECT  -2.0775 16.9875 -2.0125 17.0525 ;
        RECT  -2.6775 16.6625 -2.6125 16.7275 ;
        RECT  -2.715 16.25 -2.65 16.315 ;
        RECT  -2.6775 16.8525 -2.6125 16.9175 ;
        RECT  -2.855 16.25 -2.79 16.315 ;
        RECT  -4.2025 16.6075 -4.1375 16.6725 ;
        RECT  -4.2025 16.9875 -4.1375 17.0525 ;
        RECT  -3.6025 16.6625 -3.5375 16.7275 ;
        RECT  -3.5 16.25 -3.435 16.315 ;
        RECT  -3.6025 16.8525 -3.5375 16.9175 ;
        RECT  -3.36 16.25 -3.295 16.315 ;
        RECT  -3.9975 14.65 -3.9325 14.715 ;
        RECT  -3.9975 15.14 -3.9325 15.205 ;
        RECT  -4.1525 14.65 -4.0875 14.715 ;
        RECT  -4.1525 15.35 -4.0875 15.415 ;
        RECT  -5.5625 14.65 -5.4975 14.715 ;
        RECT  -5.5625 15.56 -5.4975 15.625 ;
        RECT  -4.5475 14.65 -4.4825 14.715 ;
        RECT  -4.5475 15.77 -4.4825 15.835 ;
        RECT  -1.325 15.35 -1.26 15.415 ;
        RECT  -0.795 15.98 -0.73 16.045 ;
        RECT  -2.12 15.98 -2.055 16.045 ;
        RECT  -2.6425 15.35 -2.5775 15.415 ;
        RECT  -2.7825 15.56 -2.7175 15.625 ;
        RECT  -4.025 15.98 -3.96 16.045 ;
        RECT  -3.5025 15.77 -3.4375 15.835 ;
        RECT  -3.3625 15.56 -3.2975 15.625 ;
        RECT  -0.9975 9.8525 -0.9325 9.9175 ;
        RECT  -0.2225 9.8525 -0.1575 9.9175 ;
        RECT  -0.22 15.1375 -0.155 15.2025 ;
        RECT  -2.49 19.44 -2.425 19.505 ;
        RECT  -3.655 19.23 -3.59 19.295 ;
        RECT  -0.965 19.65 -0.9 19.715 ;
        RECT  -0.2075 19.4375 -0.1425 19.5025 ;
        RECT  -1.7275 19.86 -1.6625 19.925 ;
        RECT  -4.4175 19.86 -4.3525 19.925 ;
        RECT  -0.3825 14.93 -0.3175 14.995 ;
        RECT  -0.965 13.4125 -0.9 13.4775 ;
        RECT  -2.0875 13.4125 -2.0225 13.4775 ;
        RECT  -2.0825 8.31 -2.0175 8.375 ;
        RECT  -0.865 8.45 -0.8 8.515 ;
        RECT  -1.0475 16.8675 -0.9825 16.9325 ;
        RECT  -1.0 17.3375 -0.935 17.4025 ;
        RECT  0.0 19.89 0.065 19.955 ;
        RECT  0.14 19.89 0.205 19.955 ;
        Layer  metal2 ; 
        RECT  -0.35 19.855 0.0 19.925 ;
        RECT  8.89 0.0 9.59 41.725 ;
        RECT  10.78 0.0 10.85 41.725 ;
        RECT  10.57 0.0 10.64 41.725 ;
        RECT  10.36 0.0 10.43 41.725 ;
        RECT  10.15 0.0 10.22 41.725 ;
        RECT  9.94 0.0 10.01 41.725 ;
        RECT  9.73 0.0 9.8 41.725 ;
        RECT  8.54 5.02 8.61 18.615 ;
        RECT  8.33 5.02 8.4 18.615 ;
        RECT  8.12 5.02 8.19 18.615 ;
        RECT  7.91 5.02 7.98 18.615 ;
        RECT  11.28 40.415 11.35 40.765 ;
        RECT  11.615 40.415 11.685 40.765 ;
        RECT  11.985 40.415 12.055 40.765 ;
        RECT  12.32 40.415 12.39 40.765 ;
        RECT  10.36 18.895 10.43 41.24 ;
        RECT  11.8 40.415 11.87 40.61 ;
        RECT  12.505 40.415 12.575 40.61 ;
        RECT  11.06 18.895 11.13 40.61 ;
        RECT  7.855 21.5525 8.89 21.6225 ;
        RECT  7.855 24.2425 8.89 24.3125 ;
        RECT  7.855 26.9325 8.89 27.0025 ;
        RECT  7.855 29.6225 8.89 29.6925 ;
        RECT  7.855 32.3125 8.89 32.3825 ;
        RECT  7.855 35.0025 8.89 35.0725 ;
        RECT  7.855 37.6925 8.89 37.7625 ;
        RECT  7.855 40.3825 8.89 40.4525 ;
        RECT  11.8 19.645 11.87 19.78 ;
        RECT  11.8 19.645 11.87 19.78 ;
        RECT  11.8 19.645 11.87 19.78 ;
        RECT  11.8 19.645 11.87 19.78 ;
        RECT  11.8 19.645 11.87 19.78 ;
        RECT  11.8 19.645 11.87 19.78 ;
        RECT  11.0625 18.86 11.1975 18.93 ;
        RECT  11.7675 18.86 11.9025 18.93 ;
        RECT  11.8 19.645 11.87 19.78 ;
        RECT  11.8 19.645 11.87 19.78 ;
        RECT  11.8 19.645 11.87 19.78 ;
        RECT  11.8 19.645 11.87 19.78 ;
        RECT  11.8 19.645 11.87 19.78 ;
        RECT  11.8 19.645 11.87 19.78 ;
        RECT  11.8 19.645 11.87 19.78 ;
        RECT  11.8 19.645 11.87 19.78 ;
        RECT  11.35 19.1525 11.42 19.2875 ;
        RECT  11.095 19.645 11.165 19.78 ;
        RECT  11.095 19.645 11.165 19.78 ;
        RECT  11.095 19.645 11.165 19.78 ;
        RECT  11.095 19.645 11.165 19.78 ;
        RECT  11.095 19.645 11.165 19.78 ;
        RECT  11.095 19.645 11.165 19.78 ;
        RECT  11.8 19.645 11.87 19.78 ;
        RECT  11.8 19.645 11.87 19.78 ;
        RECT  11.8 19.645 11.87 19.78 ;
        RECT  11.8 19.645 11.87 19.78 ;
        RECT  11.545 19.1525 11.615 19.2875 ;
        RECT  11.7675 18.86 11.9025 18.93 ;
        RECT  11.7675 18.86 11.9025 18.93 ;
        RECT  11.7675 18.86 11.9025 18.93 ;
        RECT  11.8 19.645 11.87 19.78 ;
        RECT  11.8 19.645 11.87 19.78 ;
        RECT  11.8 19.645 11.87 19.78 ;
        RECT  11.8 19.645 11.87 19.78 ;
        RECT  11.8 19.645 11.87 19.78 ;
        RECT  11.8 19.645 11.87 19.78 ;
        RECT  11.0625 18.86 11.1975 18.93 ;
        RECT  11.8 18.8625 11.87 20.2725 ;
        RECT  11.1 18.865 11.16 18.9225 ;
        RECT  11.2875 18.87 11.3425 18.9225 ;
        RECT  11.6225 18.8625 11.68 18.9225 ;
        RECT  11.805 18.87 11.865 18.9275 ;
        RECT  11.615 18.795 11.685 20.34 ;
        RECT  11.28 18.795 11.35 20.34 ;
        RECT  11.095 18.795 11.165 20.34 ;
        RECT  11.8 18.795 11.87 20.34 ;
        RECT  11.8 20.7 11.87 20.835 ;
        RECT  11.8 20.7 11.87 20.835 ;
        RECT  11.8 20.7 11.87 20.835 ;
        RECT  11.8 20.7 11.87 20.835 ;
        RECT  11.8 20.7 11.87 20.835 ;
        RECT  11.8 20.7 11.87 20.835 ;
        RECT  11.0625 21.55 11.1975 21.62 ;
        RECT  11.7675 21.55 11.9025 21.62 ;
        RECT  11.8 20.7 11.87 20.835 ;
        RECT  11.8 20.7 11.87 20.835 ;
        RECT  11.8 20.7 11.87 20.835 ;
        RECT  11.8 20.7 11.87 20.835 ;
        RECT  11.8 20.7 11.87 20.835 ;
        RECT  11.8 20.7 11.87 20.835 ;
        RECT  11.8 20.7 11.87 20.835 ;
        RECT  11.8 20.7 11.87 20.835 ;
        RECT  11.35 21.1925 11.42 21.3275 ;
        RECT  11.095 20.7 11.165 20.835 ;
        RECT  11.095 20.7 11.165 20.835 ;
        RECT  11.095 20.7 11.165 20.835 ;
        RECT  11.095 20.7 11.165 20.835 ;
        RECT  11.095 20.7 11.165 20.835 ;
        RECT  11.095 20.7 11.165 20.835 ;
        RECT  11.8 20.7 11.87 20.835 ;
        RECT  11.8 20.7 11.87 20.835 ;
        RECT  11.8 20.7 11.87 20.835 ;
        RECT  11.8 20.7 11.87 20.835 ;
        RECT  11.545 21.1925 11.615 21.3275 ;
        RECT  11.7675 21.55 11.9025 21.62 ;
        RECT  11.7675 21.55 11.9025 21.62 ;
        RECT  11.7675 21.55 11.9025 21.62 ;
        RECT  11.8 20.7 11.87 20.835 ;
        RECT  11.8 20.7 11.87 20.835 ;
        RECT  11.8 20.7 11.87 20.835 ;
        RECT  11.8 20.7 11.87 20.835 ;
        RECT  11.8 20.7 11.87 20.835 ;
        RECT  11.8 20.7 11.87 20.835 ;
        RECT  11.0625 21.55 11.1975 21.62 ;
        RECT  11.8 20.2075 11.87 21.6175 ;
        RECT  11.1 21.5575 11.16 21.615 ;
        RECT  11.2875 21.5575 11.3425 21.61 ;
        RECT  11.6225 21.5575 11.68 21.6175 ;
        RECT  11.805 21.5525 11.865 21.61 ;
        RECT  11.615 20.14 11.685 21.685 ;
        RECT  11.28 20.14 11.35 21.685 ;
        RECT  11.095 20.14 11.165 21.685 ;
        RECT  11.8 20.14 11.87 21.685 ;
        RECT  11.8 22.335 11.87 22.47 ;
        RECT  11.8 22.335 11.87 22.47 ;
        RECT  11.8 22.335 11.87 22.47 ;
        RECT  11.8 22.335 11.87 22.47 ;
        RECT  11.8 22.335 11.87 22.47 ;
        RECT  11.8 22.335 11.87 22.47 ;
        RECT  11.0625 21.55 11.1975 21.62 ;
        RECT  11.7675 21.55 11.9025 21.62 ;
        RECT  11.8 22.335 11.87 22.47 ;
        RECT  11.8 22.335 11.87 22.47 ;
        RECT  11.8 22.335 11.87 22.47 ;
        RECT  11.8 22.335 11.87 22.47 ;
        RECT  11.8 22.335 11.87 22.47 ;
        RECT  11.8 22.335 11.87 22.47 ;
        RECT  11.8 22.335 11.87 22.47 ;
        RECT  11.8 22.335 11.87 22.47 ;
        RECT  11.35 21.8425 11.42 21.9775 ;
        RECT  11.095 22.335 11.165 22.47 ;
        RECT  11.095 22.335 11.165 22.47 ;
        RECT  11.095 22.335 11.165 22.47 ;
        RECT  11.095 22.335 11.165 22.47 ;
        RECT  11.095 22.335 11.165 22.47 ;
        RECT  11.095 22.335 11.165 22.47 ;
        RECT  11.8 22.335 11.87 22.47 ;
        RECT  11.8 22.335 11.87 22.47 ;
        RECT  11.8 22.335 11.87 22.47 ;
        RECT  11.8 22.335 11.87 22.47 ;
        RECT  11.545 21.8425 11.615 21.9775 ;
        RECT  11.7675 21.55 11.9025 21.62 ;
        RECT  11.7675 21.55 11.9025 21.62 ;
        RECT  11.7675 21.55 11.9025 21.62 ;
        RECT  11.8 22.335 11.87 22.47 ;
        RECT  11.8 22.335 11.87 22.47 ;
        RECT  11.8 22.335 11.87 22.47 ;
        RECT  11.8 22.335 11.87 22.47 ;
        RECT  11.8 22.335 11.87 22.47 ;
        RECT  11.8 22.335 11.87 22.47 ;
        RECT  11.0625 21.55 11.1975 21.62 ;
        RECT  11.8 21.5525 11.87 22.9625 ;
        RECT  11.1 21.555 11.16 21.6125 ;
        RECT  11.2875 21.56 11.3425 21.6125 ;
        RECT  11.6225 21.5525 11.68 21.6125 ;
        RECT  11.805 21.56 11.865 21.6175 ;
        RECT  11.615 21.485 11.685 23.03 ;
        RECT  11.28 21.485 11.35 23.03 ;
        RECT  11.095 21.485 11.165 23.03 ;
        RECT  11.8 21.485 11.87 23.03 ;
        RECT  11.8 23.39 11.87 23.525 ;
        RECT  11.8 23.39 11.87 23.525 ;
        RECT  11.8 23.39 11.87 23.525 ;
        RECT  11.8 23.39 11.87 23.525 ;
        RECT  11.8 23.39 11.87 23.525 ;
        RECT  11.8 23.39 11.87 23.525 ;
        RECT  11.0625 24.24 11.1975 24.31 ;
        RECT  11.7675 24.24 11.9025 24.31 ;
        RECT  11.8 23.39 11.87 23.525 ;
        RECT  11.8 23.39 11.87 23.525 ;
        RECT  11.8 23.39 11.87 23.525 ;
        RECT  11.8 23.39 11.87 23.525 ;
        RECT  11.8 23.39 11.87 23.525 ;
        RECT  11.8 23.39 11.87 23.525 ;
        RECT  11.8 23.39 11.87 23.525 ;
        RECT  11.8 23.39 11.87 23.525 ;
        RECT  11.35 23.8825 11.42 24.0175 ;
        RECT  11.095 23.39 11.165 23.525 ;
        RECT  11.095 23.39 11.165 23.525 ;
        RECT  11.095 23.39 11.165 23.525 ;
        RECT  11.095 23.39 11.165 23.525 ;
        RECT  11.095 23.39 11.165 23.525 ;
        RECT  11.095 23.39 11.165 23.525 ;
        RECT  11.8 23.39 11.87 23.525 ;
        RECT  11.8 23.39 11.87 23.525 ;
        RECT  11.8 23.39 11.87 23.525 ;
        RECT  11.8 23.39 11.87 23.525 ;
        RECT  11.545 23.8825 11.615 24.0175 ;
        RECT  11.7675 24.24 11.9025 24.31 ;
        RECT  11.7675 24.24 11.9025 24.31 ;
        RECT  11.7675 24.24 11.9025 24.31 ;
        RECT  11.8 23.39 11.87 23.525 ;
        RECT  11.8 23.39 11.87 23.525 ;
        RECT  11.8 23.39 11.87 23.525 ;
        RECT  11.8 23.39 11.87 23.525 ;
        RECT  11.8 23.39 11.87 23.525 ;
        RECT  11.8 23.39 11.87 23.525 ;
        RECT  11.0625 24.24 11.1975 24.31 ;
        RECT  11.8 22.8975 11.87 24.3075 ;
        RECT  11.1 24.2475 11.16 24.305 ;
        RECT  11.2875 24.2475 11.3425 24.3 ;
        RECT  11.6225 24.2475 11.68 24.3075 ;
        RECT  11.805 24.2425 11.865 24.3 ;
        RECT  11.615 22.83 11.685 24.375 ;
        RECT  11.28 22.83 11.35 24.375 ;
        RECT  11.095 22.83 11.165 24.375 ;
        RECT  11.8 22.83 11.87 24.375 ;
        RECT  11.8 25.025 11.87 25.16 ;
        RECT  11.8 25.025 11.87 25.16 ;
        RECT  11.8 25.025 11.87 25.16 ;
        RECT  11.8 25.025 11.87 25.16 ;
        RECT  11.8 25.025 11.87 25.16 ;
        RECT  11.8 25.025 11.87 25.16 ;
        RECT  11.0625 24.24 11.1975 24.31 ;
        RECT  11.7675 24.24 11.9025 24.31 ;
        RECT  11.8 25.025 11.87 25.16 ;
        RECT  11.8 25.025 11.87 25.16 ;
        RECT  11.8 25.025 11.87 25.16 ;
        RECT  11.8 25.025 11.87 25.16 ;
        RECT  11.8 25.025 11.87 25.16 ;
        RECT  11.8 25.025 11.87 25.16 ;
        RECT  11.8 25.025 11.87 25.16 ;
        RECT  11.8 25.025 11.87 25.16 ;
        RECT  11.35 24.5325 11.42 24.6675 ;
        RECT  11.095 25.025 11.165 25.16 ;
        RECT  11.095 25.025 11.165 25.16 ;
        RECT  11.095 25.025 11.165 25.16 ;
        RECT  11.095 25.025 11.165 25.16 ;
        RECT  11.095 25.025 11.165 25.16 ;
        RECT  11.095 25.025 11.165 25.16 ;
        RECT  11.8 25.025 11.87 25.16 ;
        RECT  11.8 25.025 11.87 25.16 ;
        RECT  11.8 25.025 11.87 25.16 ;
        RECT  11.8 25.025 11.87 25.16 ;
        RECT  11.545 24.5325 11.615 24.6675 ;
        RECT  11.7675 24.24 11.9025 24.31 ;
        RECT  11.7675 24.24 11.9025 24.31 ;
        RECT  11.7675 24.24 11.9025 24.31 ;
        RECT  11.8 25.025 11.87 25.16 ;
        RECT  11.8 25.025 11.87 25.16 ;
        RECT  11.8 25.025 11.87 25.16 ;
        RECT  11.8 25.025 11.87 25.16 ;
        RECT  11.8 25.025 11.87 25.16 ;
        RECT  11.8 25.025 11.87 25.16 ;
        RECT  11.0625 24.24 11.1975 24.31 ;
        RECT  11.8 24.2425 11.87 25.6525 ;
        RECT  11.1 24.245 11.16 24.3025 ;
        RECT  11.2875 24.25 11.3425 24.3025 ;
        RECT  11.6225 24.2425 11.68 24.3025 ;
        RECT  11.805 24.25 11.865 24.3075 ;
        RECT  11.615 24.175 11.685 25.72 ;
        RECT  11.28 24.175 11.35 25.72 ;
        RECT  11.095 24.175 11.165 25.72 ;
        RECT  11.8 24.175 11.87 25.72 ;
        RECT  11.8 26.08 11.87 26.215 ;
        RECT  11.8 26.08 11.87 26.215 ;
        RECT  11.8 26.08 11.87 26.215 ;
        RECT  11.8 26.08 11.87 26.215 ;
        RECT  11.8 26.08 11.87 26.215 ;
        RECT  11.8 26.08 11.87 26.215 ;
        RECT  11.0625 26.93 11.1975 27.0 ;
        RECT  11.7675 26.93 11.9025 27.0 ;
        RECT  11.8 26.08 11.87 26.215 ;
        RECT  11.8 26.08 11.87 26.215 ;
        RECT  11.8 26.08 11.87 26.215 ;
        RECT  11.8 26.08 11.87 26.215 ;
        RECT  11.8 26.08 11.87 26.215 ;
        RECT  11.8 26.08 11.87 26.215 ;
        RECT  11.8 26.08 11.87 26.215 ;
        RECT  11.8 26.08 11.87 26.215 ;
        RECT  11.35 26.5725 11.42 26.7075 ;
        RECT  11.095 26.08 11.165 26.215 ;
        RECT  11.095 26.08 11.165 26.215 ;
        RECT  11.095 26.08 11.165 26.215 ;
        RECT  11.095 26.08 11.165 26.215 ;
        RECT  11.095 26.08 11.165 26.215 ;
        RECT  11.095 26.08 11.165 26.215 ;
        RECT  11.8 26.08 11.87 26.215 ;
        RECT  11.8 26.08 11.87 26.215 ;
        RECT  11.8 26.08 11.87 26.215 ;
        RECT  11.8 26.08 11.87 26.215 ;
        RECT  11.545 26.5725 11.615 26.7075 ;
        RECT  11.7675 26.93 11.9025 27.0 ;
        RECT  11.7675 26.93 11.9025 27.0 ;
        RECT  11.7675 26.93 11.9025 27.0 ;
        RECT  11.8 26.08 11.87 26.215 ;
        RECT  11.8 26.08 11.87 26.215 ;
        RECT  11.8 26.08 11.87 26.215 ;
        RECT  11.8 26.08 11.87 26.215 ;
        RECT  11.8 26.08 11.87 26.215 ;
        RECT  11.8 26.08 11.87 26.215 ;
        RECT  11.0625 26.93 11.1975 27.0 ;
        RECT  11.8 25.5875 11.87 26.9975 ;
        RECT  11.1 26.9375 11.16 26.995 ;
        RECT  11.2875 26.9375 11.3425 26.99 ;
        RECT  11.6225 26.9375 11.68 26.9975 ;
        RECT  11.805 26.9325 11.865 26.99 ;
        RECT  11.615 25.52 11.685 27.065 ;
        RECT  11.28 25.52 11.35 27.065 ;
        RECT  11.095 25.52 11.165 27.065 ;
        RECT  11.8 25.52 11.87 27.065 ;
        RECT  11.8 27.715 11.87 27.85 ;
        RECT  11.8 27.715 11.87 27.85 ;
        RECT  11.8 27.715 11.87 27.85 ;
        RECT  11.8 27.715 11.87 27.85 ;
        RECT  11.8 27.715 11.87 27.85 ;
        RECT  11.8 27.715 11.87 27.85 ;
        RECT  11.0625 26.93 11.1975 27.0 ;
        RECT  11.7675 26.93 11.9025 27.0 ;
        RECT  11.8 27.715 11.87 27.85 ;
        RECT  11.8 27.715 11.87 27.85 ;
        RECT  11.8 27.715 11.87 27.85 ;
        RECT  11.8 27.715 11.87 27.85 ;
        RECT  11.8 27.715 11.87 27.85 ;
        RECT  11.8 27.715 11.87 27.85 ;
        RECT  11.8 27.715 11.87 27.85 ;
        RECT  11.8 27.715 11.87 27.85 ;
        RECT  11.35 27.2225 11.42 27.3575 ;
        RECT  11.095 27.715 11.165 27.85 ;
        RECT  11.095 27.715 11.165 27.85 ;
        RECT  11.095 27.715 11.165 27.85 ;
        RECT  11.095 27.715 11.165 27.85 ;
        RECT  11.095 27.715 11.165 27.85 ;
        RECT  11.095 27.715 11.165 27.85 ;
        RECT  11.8 27.715 11.87 27.85 ;
        RECT  11.8 27.715 11.87 27.85 ;
        RECT  11.8 27.715 11.87 27.85 ;
        RECT  11.8 27.715 11.87 27.85 ;
        RECT  11.545 27.2225 11.615 27.3575 ;
        RECT  11.7675 26.93 11.9025 27.0 ;
        RECT  11.7675 26.93 11.9025 27.0 ;
        RECT  11.7675 26.93 11.9025 27.0 ;
        RECT  11.8 27.715 11.87 27.85 ;
        RECT  11.8 27.715 11.87 27.85 ;
        RECT  11.8 27.715 11.87 27.85 ;
        RECT  11.8 27.715 11.87 27.85 ;
        RECT  11.8 27.715 11.87 27.85 ;
        RECT  11.8 27.715 11.87 27.85 ;
        RECT  11.0625 26.93 11.1975 27.0 ;
        RECT  11.8 26.9325 11.87 28.3425 ;
        RECT  11.1 26.935 11.16 26.9925 ;
        RECT  11.2875 26.94 11.3425 26.9925 ;
        RECT  11.6225 26.9325 11.68 26.9925 ;
        RECT  11.805 26.94 11.865 26.9975 ;
        RECT  11.615 26.865 11.685 28.41 ;
        RECT  11.28 26.865 11.35 28.41 ;
        RECT  11.095 26.865 11.165 28.41 ;
        RECT  11.8 26.865 11.87 28.41 ;
        RECT  11.8 28.77 11.87 28.905 ;
        RECT  11.8 28.77 11.87 28.905 ;
        RECT  11.8 28.77 11.87 28.905 ;
        RECT  11.8 28.77 11.87 28.905 ;
        RECT  11.8 28.77 11.87 28.905 ;
        RECT  11.8 28.77 11.87 28.905 ;
        RECT  11.0625 29.62 11.1975 29.69 ;
        RECT  11.7675 29.62 11.9025 29.69 ;
        RECT  11.8 28.77 11.87 28.905 ;
        RECT  11.8 28.77 11.87 28.905 ;
        RECT  11.8 28.77 11.87 28.905 ;
        RECT  11.8 28.77 11.87 28.905 ;
        RECT  11.8 28.77 11.87 28.905 ;
        RECT  11.8 28.77 11.87 28.905 ;
        RECT  11.8 28.77 11.87 28.905 ;
        RECT  11.8 28.77 11.87 28.905 ;
        RECT  11.35 29.2625 11.42 29.3975 ;
        RECT  11.095 28.77 11.165 28.905 ;
        RECT  11.095 28.77 11.165 28.905 ;
        RECT  11.095 28.77 11.165 28.905 ;
        RECT  11.095 28.77 11.165 28.905 ;
        RECT  11.095 28.77 11.165 28.905 ;
        RECT  11.095 28.77 11.165 28.905 ;
        RECT  11.8 28.77 11.87 28.905 ;
        RECT  11.8 28.77 11.87 28.905 ;
        RECT  11.8 28.77 11.87 28.905 ;
        RECT  11.8 28.77 11.87 28.905 ;
        RECT  11.545 29.2625 11.615 29.3975 ;
        RECT  11.7675 29.62 11.9025 29.69 ;
        RECT  11.7675 29.62 11.9025 29.69 ;
        RECT  11.7675 29.62 11.9025 29.69 ;
        RECT  11.8 28.77 11.87 28.905 ;
        RECT  11.8 28.77 11.87 28.905 ;
        RECT  11.8 28.77 11.87 28.905 ;
        RECT  11.8 28.77 11.87 28.905 ;
        RECT  11.8 28.77 11.87 28.905 ;
        RECT  11.8 28.77 11.87 28.905 ;
        RECT  11.0625 29.62 11.1975 29.69 ;
        RECT  11.8 28.2775 11.87 29.6875 ;
        RECT  11.1 29.6275 11.16 29.685 ;
        RECT  11.2875 29.6275 11.3425 29.68 ;
        RECT  11.6225 29.6275 11.68 29.6875 ;
        RECT  11.805 29.6225 11.865 29.68 ;
        RECT  11.615 28.21 11.685 29.755 ;
        RECT  11.28 28.21 11.35 29.755 ;
        RECT  11.095 28.21 11.165 29.755 ;
        RECT  11.8 28.21 11.87 29.755 ;
        RECT  11.8 30.405 11.87 30.54 ;
        RECT  11.8 30.405 11.87 30.54 ;
        RECT  11.8 30.405 11.87 30.54 ;
        RECT  11.8 30.405 11.87 30.54 ;
        RECT  11.8 30.405 11.87 30.54 ;
        RECT  11.8 30.405 11.87 30.54 ;
        RECT  11.0625 29.62 11.1975 29.69 ;
        RECT  11.7675 29.62 11.9025 29.69 ;
        RECT  11.8 30.405 11.87 30.54 ;
        RECT  11.8 30.405 11.87 30.54 ;
        RECT  11.8 30.405 11.87 30.54 ;
        RECT  11.8 30.405 11.87 30.54 ;
        RECT  11.8 30.405 11.87 30.54 ;
        RECT  11.8 30.405 11.87 30.54 ;
        RECT  11.8 30.405 11.87 30.54 ;
        RECT  11.8 30.405 11.87 30.54 ;
        RECT  11.35 29.9125 11.42 30.0475 ;
        RECT  11.095 30.405 11.165 30.54 ;
        RECT  11.095 30.405 11.165 30.54 ;
        RECT  11.095 30.405 11.165 30.54 ;
        RECT  11.095 30.405 11.165 30.54 ;
        RECT  11.095 30.405 11.165 30.54 ;
        RECT  11.095 30.405 11.165 30.54 ;
        RECT  11.8 30.405 11.87 30.54 ;
        RECT  11.8 30.405 11.87 30.54 ;
        RECT  11.8 30.405 11.87 30.54 ;
        RECT  11.8 30.405 11.87 30.54 ;
        RECT  11.545 29.9125 11.615 30.0475 ;
        RECT  11.7675 29.62 11.9025 29.69 ;
        RECT  11.7675 29.62 11.9025 29.69 ;
        RECT  11.7675 29.62 11.9025 29.69 ;
        RECT  11.8 30.405 11.87 30.54 ;
        RECT  11.8 30.405 11.87 30.54 ;
        RECT  11.8 30.405 11.87 30.54 ;
        RECT  11.8 30.405 11.87 30.54 ;
        RECT  11.8 30.405 11.87 30.54 ;
        RECT  11.8 30.405 11.87 30.54 ;
        RECT  11.0625 29.62 11.1975 29.69 ;
        RECT  11.8 29.6225 11.87 31.0325 ;
        RECT  11.1 29.625 11.16 29.6825 ;
        RECT  11.2875 29.63 11.3425 29.6825 ;
        RECT  11.6225 29.6225 11.68 29.6825 ;
        RECT  11.805 29.63 11.865 29.6875 ;
        RECT  11.615 29.555 11.685 31.1 ;
        RECT  11.28 29.555 11.35 31.1 ;
        RECT  11.095 29.555 11.165 31.1 ;
        RECT  11.8 29.555 11.87 31.1 ;
        RECT  11.8 31.46 11.87 31.595 ;
        RECT  11.8 31.46 11.87 31.595 ;
        RECT  11.8 31.46 11.87 31.595 ;
        RECT  11.8 31.46 11.87 31.595 ;
        RECT  11.8 31.46 11.87 31.595 ;
        RECT  11.8 31.46 11.87 31.595 ;
        RECT  11.0625 32.31 11.1975 32.38 ;
        RECT  11.7675 32.31 11.9025 32.38 ;
        RECT  11.8 31.46 11.87 31.595 ;
        RECT  11.8 31.46 11.87 31.595 ;
        RECT  11.8 31.46 11.87 31.595 ;
        RECT  11.8 31.46 11.87 31.595 ;
        RECT  11.8 31.46 11.87 31.595 ;
        RECT  11.8 31.46 11.87 31.595 ;
        RECT  11.8 31.46 11.87 31.595 ;
        RECT  11.8 31.46 11.87 31.595 ;
        RECT  11.35 31.9525 11.42 32.0875 ;
        RECT  11.095 31.46 11.165 31.595 ;
        RECT  11.095 31.46 11.165 31.595 ;
        RECT  11.095 31.46 11.165 31.595 ;
        RECT  11.095 31.46 11.165 31.595 ;
        RECT  11.095 31.46 11.165 31.595 ;
        RECT  11.095 31.46 11.165 31.595 ;
        RECT  11.8 31.46 11.87 31.595 ;
        RECT  11.8 31.46 11.87 31.595 ;
        RECT  11.8 31.46 11.87 31.595 ;
        RECT  11.8 31.46 11.87 31.595 ;
        RECT  11.545 31.9525 11.615 32.0875 ;
        RECT  11.7675 32.31 11.9025 32.38 ;
        RECT  11.7675 32.31 11.9025 32.38 ;
        RECT  11.7675 32.31 11.9025 32.38 ;
        RECT  11.8 31.46 11.87 31.595 ;
        RECT  11.8 31.46 11.87 31.595 ;
        RECT  11.8 31.46 11.87 31.595 ;
        RECT  11.8 31.46 11.87 31.595 ;
        RECT  11.8 31.46 11.87 31.595 ;
        RECT  11.8 31.46 11.87 31.595 ;
        RECT  11.0625 32.31 11.1975 32.38 ;
        RECT  11.8 30.9675 11.87 32.3775 ;
        RECT  11.1 32.3175 11.16 32.375 ;
        RECT  11.2875 32.3175 11.3425 32.37 ;
        RECT  11.6225 32.3175 11.68 32.3775 ;
        RECT  11.805 32.3125 11.865 32.37 ;
        RECT  11.615 30.9 11.685 32.445 ;
        RECT  11.28 30.9 11.35 32.445 ;
        RECT  11.095 30.9 11.165 32.445 ;
        RECT  11.8 30.9 11.87 32.445 ;
        RECT  11.8 33.095 11.87 33.23 ;
        RECT  11.8 33.095 11.87 33.23 ;
        RECT  11.8 33.095 11.87 33.23 ;
        RECT  11.8 33.095 11.87 33.23 ;
        RECT  11.8 33.095 11.87 33.23 ;
        RECT  11.8 33.095 11.87 33.23 ;
        RECT  11.0625 32.31 11.1975 32.38 ;
        RECT  11.7675 32.31 11.9025 32.38 ;
        RECT  11.8 33.095 11.87 33.23 ;
        RECT  11.8 33.095 11.87 33.23 ;
        RECT  11.8 33.095 11.87 33.23 ;
        RECT  11.8 33.095 11.87 33.23 ;
        RECT  11.8 33.095 11.87 33.23 ;
        RECT  11.8 33.095 11.87 33.23 ;
        RECT  11.8 33.095 11.87 33.23 ;
        RECT  11.8 33.095 11.87 33.23 ;
        RECT  11.35 32.6025 11.42 32.7375 ;
        RECT  11.095 33.095 11.165 33.23 ;
        RECT  11.095 33.095 11.165 33.23 ;
        RECT  11.095 33.095 11.165 33.23 ;
        RECT  11.095 33.095 11.165 33.23 ;
        RECT  11.095 33.095 11.165 33.23 ;
        RECT  11.095 33.095 11.165 33.23 ;
        RECT  11.8 33.095 11.87 33.23 ;
        RECT  11.8 33.095 11.87 33.23 ;
        RECT  11.8 33.095 11.87 33.23 ;
        RECT  11.8 33.095 11.87 33.23 ;
        RECT  11.545 32.6025 11.615 32.7375 ;
        RECT  11.7675 32.31 11.9025 32.38 ;
        RECT  11.7675 32.31 11.9025 32.38 ;
        RECT  11.7675 32.31 11.9025 32.38 ;
        RECT  11.8 33.095 11.87 33.23 ;
        RECT  11.8 33.095 11.87 33.23 ;
        RECT  11.8 33.095 11.87 33.23 ;
        RECT  11.8 33.095 11.87 33.23 ;
        RECT  11.8 33.095 11.87 33.23 ;
        RECT  11.8 33.095 11.87 33.23 ;
        RECT  11.0625 32.31 11.1975 32.38 ;
        RECT  11.8 32.3125 11.87 33.7225 ;
        RECT  11.1 32.315 11.16 32.3725 ;
        RECT  11.2875 32.32 11.3425 32.3725 ;
        RECT  11.6225 32.3125 11.68 32.3725 ;
        RECT  11.805 32.32 11.865 32.3775 ;
        RECT  11.615 32.245 11.685 33.79 ;
        RECT  11.28 32.245 11.35 33.79 ;
        RECT  11.095 32.245 11.165 33.79 ;
        RECT  11.8 32.245 11.87 33.79 ;
        RECT  11.8 34.15 11.87 34.285 ;
        RECT  11.8 34.15 11.87 34.285 ;
        RECT  11.8 34.15 11.87 34.285 ;
        RECT  11.8 34.15 11.87 34.285 ;
        RECT  11.8 34.15 11.87 34.285 ;
        RECT  11.8 34.15 11.87 34.285 ;
        RECT  11.0625 35.0 11.1975 35.07 ;
        RECT  11.7675 35.0 11.9025 35.07 ;
        RECT  11.8 34.15 11.87 34.285 ;
        RECT  11.8 34.15 11.87 34.285 ;
        RECT  11.8 34.15 11.87 34.285 ;
        RECT  11.8 34.15 11.87 34.285 ;
        RECT  11.8 34.15 11.87 34.285 ;
        RECT  11.8 34.15 11.87 34.285 ;
        RECT  11.8 34.15 11.87 34.285 ;
        RECT  11.8 34.15 11.87 34.285 ;
        RECT  11.35 34.6425 11.42 34.7775 ;
        RECT  11.095 34.15 11.165 34.285 ;
        RECT  11.095 34.15 11.165 34.285 ;
        RECT  11.095 34.15 11.165 34.285 ;
        RECT  11.095 34.15 11.165 34.285 ;
        RECT  11.095 34.15 11.165 34.285 ;
        RECT  11.095 34.15 11.165 34.285 ;
        RECT  11.8 34.15 11.87 34.285 ;
        RECT  11.8 34.15 11.87 34.285 ;
        RECT  11.8 34.15 11.87 34.285 ;
        RECT  11.8 34.15 11.87 34.285 ;
        RECT  11.545 34.6425 11.615 34.7775 ;
        RECT  11.7675 35.0 11.9025 35.07 ;
        RECT  11.7675 35.0 11.9025 35.07 ;
        RECT  11.7675 35.0 11.9025 35.07 ;
        RECT  11.8 34.15 11.87 34.285 ;
        RECT  11.8 34.15 11.87 34.285 ;
        RECT  11.8 34.15 11.87 34.285 ;
        RECT  11.8 34.15 11.87 34.285 ;
        RECT  11.8 34.15 11.87 34.285 ;
        RECT  11.8 34.15 11.87 34.285 ;
        RECT  11.0625 35.0 11.1975 35.07 ;
        RECT  11.8 33.6575 11.87 35.0675 ;
        RECT  11.1 35.0075 11.16 35.065 ;
        RECT  11.2875 35.0075 11.3425 35.06 ;
        RECT  11.6225 35.0075 11.68 35.0675 ;
        RECT  11.805 35.0025 11.865 35.06 ;
        RECT  11.615 33.59 11.685 35.135 ;
        RECT  11.28 33.59 11.35 35.135 ;
        RECT  11.095 33.59 11.165 35.135 ;
        RECT  11.8 33.59 11.87 35.135 ;
        RECT  11.8 35.785 11.87 35.92 ;
        RECT  11.8 35.785 11.87 35.92 ;
        RECT  11.8 35.785 11.87 35.92 ;
        RECT  11.8 35.785 11.87 35.92 ;
        RECT  11.8 35.785 11.87 35.92 ;
        RECT  11.8 35.785 11.87 35.92 ;
        RECT  11.0625 35.0 11.1975 35.07 ;
        RECT  11.7675 35.0 11.9025 35.07 ;
        RECT  11.8 35.785 11.87 35.92 ;
        RECT  11.8 35.785 11.87 35.92 ;
        RECT  11.8 35.785 11.87 35.92 ;
        RECT  11.8 35.785 11.87 35.92 ;
        RECT  11.8 35.785 11.87 35.92 ;
        RECT  11.8 35.785 11.87 35.92 ;
        RECT  11.8 35.785 11.87 35.92 ;
        RECT  11.8 35.785 11.87 35.92 ;
        RECT  11.35 35.2925 11.42 35.4275 ;
        RECT  11.095 35.785 11.165 35.92 ;
        RECT  11.095 35.785 11.165 35.92 ;
        RECT  11.095 35.785 11.165 35.92 ;
        RECT  11.095 35.785 11.165 35.92 ;
        RECT  11.095 35.785 11.165 35.92 ;
        RECT  11.095 35.785 11.165 35.92 ;
        RECT  11.8 35.785 11.87 35.92 ;
        RECT  11.8 35.785 11.87 35.92 ;
        RECT  11.8 35.785 11.87 35.92 ;
        RECT  11.8 35.785 11.87 35.92 ;
        RECT  11.545 35.2925 11.615 35.4275 ;
        RECT  11.7675 35.0 11.9025 35.07 ;
        RECT  11.7675 35.0 11.9025 35.07 ;
        RECT  11.7675 35.0 11.9025 35.07 ;
        RECT  11.8 35.785 11.87 35.92 ;
        RECT  11.8 35.785 11.87 35.92 ;
        RECT  11.8 35.785 11.87 35.92 ;
        RECT  11.8 35.785 11.87 35.92 ;
        RECT  11.8 35.785 11.87 35.92 ;
        RECT  11.8 35.785 11.87 35.92 ;
        RECT  11.0625 35.0 11.1975 35.07 ;
        RECT  11.8 35.0025 11.87 36.4125 ;
        RECT  11.1 35.005 11.16 35.0625 ;
        RECT  11.2875 35.01 11.3425 35.0625 ;
        RECT  11.6225 35.0025 11.68 35.0625 ;
        RECT  11.805 35.01 11.865 35.0675 ;
        RECT  11.615 34.935 11.685 36.48 ;
        RECT  11.28 34.935 11.35 36.48 ;
        RECT  11.095 34.935 11.165 36.48 ;
        RECT  11.8 34.935 11.87 36.48 ;
        RECT  11.8 36.84 11.87 36.975 ;
        RECT  11.8 36.84 11.87 36.975 ;
        RECT  11.8 36.84 11.87 36.975 ;
        RECT  11.8 36.84 11.87 36.975 ;
        RECT  11.8 36.84 11.87 36.975 ;
        RECT  11.8 36.84 11.87 36.975 ;
        RECT  11.0625 37.69 11.1975 37.76 ;
        RECT  11.7675 37.69 11.9025 37.76 ;
        RECT  11.8 36.84 11.87 36.975 ;
        RECT  11.8 36.84 11.87 36.975 ;
        RECT  11.8 36.84 11.87 36.975 ;
        RECT  11.8 36.84 11.87 36.975 ;
        RECT  11.8 36.84 11.87 36.975 ;
        RECT  11.8 36.84 11.87 36.975 ;
        RECT  11.8 36.84 11.87 36.975 ;
        RECT  11.8 36.84 11.87 36.975 ;
        RECT  11.35 37.3325 11.42 37.4675 ;
        RECT  11.095 36.84 11.165 36.975 ;
        RECT  11.095 36.84 11.165 36.975 ;
        RECT  11.095 36.84 11.165 36.975 ;
        RECT  11.095 36.84 11.165 36.975 ;
        RECT  11.095 36.84 11.165 36.975 ;
        RECT  11.095 36.84 11.165 36.975 ;
        RECT  11.8 36.84 11.87 36.975 ;
        RECT  11.8 36.84 11.87 36.975 ;
        RECT  11.8 36.84 11.87 36.975 ;
        RECT  11.8 36.84 11.87 36.975 ;
        RECT  11.545 37.3325 11.615 37.4675 ;
        RECT  11.7675 37.69 11.9025 37.76 ;
        RECT  11.7675 37.69 11.9025 37.76 ;
        RECT  11.7675 37.69 11.9025 37.76 ;
        RECT  11.8 36.84 11.87 36.975 ;
        RECT  11.8 36.84 11.87 36.975 ;
        RECT  11.8 36.84 11.87 36.975 ;
        RECT  11.8 36.84 11.87 36.975 ;
        RECT  11.8 36.84 11.87 36.975 ;
        RECT  11.8 36.84 11.87 36.975 ;
        RECT  11.0625 37.69 11.1975 37.76 ;
        RECT  11.8 36.3475 11.87 37.7575 ;
        RECT  11.1 37.6975 11.16 37.755 ;
        RECT  11.2875 37.6975 11.3425 37.75 ;
        RECT  11.6225 37.6975 11.68 37.7575 ;
        RECT  11.805 37.6925 11.865 37.75 ;
        RECT  11.615 36.28 11.685 37.825 ;
        RECT  11.28 36.28 11.35 37.825 ;
        RECT  11.095 36.28 11.165 37.825 ;
        RECT  11.8 36.28 11.87 37.825 ;
        RECT  11.8 38.475 11.87 38.61 ;
        RECT  11.8 38.475 11.87 38.61 ;
        RECT  11.8 38.475 11.87 38.61 ;
        RECT  11.8 38.475 11.87 38.61 ;
        RECT  11.8 38.475 11.87 38.61 ;
        RECT  11.8 38.475 11.87 38.61 ;
        RECT  11.0625 37.69 11.1975 37.76 ;
        RECT  11.7675 37.69 11.9025 37.76 ;
        RECT  11.8 38.475 11.87 38.61 ;
        RECT  11.8 38.475 11.87 38.61 ;
        RECT  11.8 38.475 11.87 38.61 ;
        RECT  11.8 38.475 11.87 38.61 ;
        RECT  11.8 38.475 11.87 38.61 ;
        RECT  11.8 38.475 11.87 38.61 ;
        RECT  11.8 38.475 11.87 38.61 ;
        RECT  11.8 38.475 11.87 38.61 ;
        RECT  11.35 37.9825 11.42 38.1175 ;
        RECT  11.095 38.475 11.165 38.61 ;
        RECT  11.095 38.475 11.165 38.61 ;
        RECT  11.095 38.475 11.165 38.61 ;
        RECT  11.095 38.475 11.165 38.61 ;
        RECT  11.095 38.475 11.165 38.61 ;
        RECT  11.095 38.475 11.165 38.61 ;
        RECT  11.8 38.475 11.87 38.61 ;
        RECT  11.8 38.475 11.87 38.61 ;
        RECT  11.8 38.475 11.87 38.61 ;
        RECT  11.8 38.475 11.87 38.61 ;
        RECT  11.545 37.9825 11.615 38.1175 ;
        RECT  11.7675 37.69 11.9025 37.76 ;
        RECT  11.7675 37.69 11.9025 37.76 ;
        RECT  11.7675 37.69 11.9025 37.76 ;
        RECT  11.8 38.475 11.87 38.61 ;
        RECT  11.8 38.475 11.87 38.61 ;
        RECT  11.8 38.475 11.87 38.61 ;
        RECT  11.8 38.475 11.87 38.61 ;
        RECT  11.8 38.475 11.87 38.61 ;
        RECT  11.8 38.475 11.87 38.61 ;
        RECT  11.0625 37.69 11.1975 37.76 ;
        RECT  11.8 37.6925 11.87 39.1025 ;
        RECT  11.1 37.695 11.16 37.7525 ;
        RECT  11.2875 37.7 11.3425 37.7525 ;
        RECT  11.6225 37.6925 11.68 37.7525 ;
        RECT  11.805 37.7 11.865 37.7575 ;
        RECT  11.615 37.625 11.685 39.17 ;
        RECT  11.28 37.625 11.35 39.17 ;
        RECT  11.095 37.625 11.165 39.17 ;
        RECT  11.8 37.625 11.87 39.17 ;
        RECT  11.8 39.53 11.87 39.665 ;
        RECT  11.8 39.53 11.87 39.665 ;
        RECT  11.8 39.53 11.87 39.665 ;
        RECT  11.8 39.53 11.87 39.665 ;
        RECT  11.8 39.53 11.87 39.665 ;
        RECT  11.8 39.53 11.87 39.665 ;
        RECT  11.0625 40.38 11.1975 40.45 ;
        RECT  11.7675 40.38 11.9025 40.45 ;
        RECT  11.8 39.53 11.87 39.665 ;
        RECT  11.8 39.53 11.87 39.665 ;
        RECT  11.8 39.53 11.87 39.665 ;
        RECT  11.8 39.53 11.87 39.665 ;
        RECT  11.8 39.53 11.87 39.665 ;
        RECT  11.8 39.53 11.87 39.665 ;
        RECT  11.8 39.53 11.87 39.665 ;
        RECT  11.8 39.53 11.87 39.665 ;
        RECT  11.35 40.0225 11.42 40.1575 ;
        RECT  11.095 39.53 11.165 39.665 ;
        RECT  11.095 39.53 11.165 39.665 ;
        RECT  11.095 39.53 11.165 39.665 ;
        RECT  11.095 39.53 11.165 39.665 ;
        RECT  11.095 39.53 11.165 39.665 ;
        RECT  11.095 39.53 11.165 39.665 ;
        RECT  11.8 39.53 11.87 39.665 ;
        RECT  11.8 39.53 11.87 39.665 ;
        RECT  11.8 39.53 11.87 39.665 ;
        RECT  11.8 39.53 11.87 39.665 ;
        RECT  11.545 40.0225 11.615 40.1575 ;
        RECT  11.7675 40.38 11.9025 40.45 ;
        RECT  11.7675 40.38 11.9025 40.45 ;
        RECT  11.7675 40.38 11.9025 40.45 ;
        RECT  11.8 39.53 11.87 39.665 ;
        RECT  11.8 39.53 11.87 39.665 ;
        RECT  11.8 39.53 11.87 39.665 ;
        RECT  11.8 39.53 11.87 39.665 ;
        RECT  11.8 39.53 11.87 39.665 ;
        RECT  11.8 39.53 11.87 39.665 ;
        RECT  11.0625 40.38 11.1975 40.45 ;
        RECT  11.8 39.0375 11.87 40.4475 ;
        RECT  11.1 40.3875 11.16 40.445 ;
        RECT  11.2875 40.3875 11.3425 40.44 ;
        RECT  11.6225 40.3875 11.68 40.4475 ;
        RECT  11.805 40.3825 11.865 40.44 ;
        RECT  11.615 38.97 11.685 40.515 ;
        RECT  11.28 38.97 11.35 40.515 ;
        RECT  11.095 38.97 11.165 40.515 ;
        RECT  11.8 38.97 11.87 40.515 ;
        RECT  12.505 19.645 12.575 19.78 ;
        RECT  12.505 19.645 12.575 19.78 ;
        RECT  12.505 19.645 12.575 19.78 ;
        RECT  12.505 19.645 12.575 19.78 ;
        RECT  12.505 19.645 12.575 19.78 ;
        RECT  12.505 19.645 12.575 19.78 ;
        RECT  11.7675 18.86 11.9025 18.93 ;
        RECT  12.4725 18.86 12.6075 18.93 ;
        RECT  12.505 19.645 12.575 19.78 ;
        RECT  12.505 19.645 12.575 19.78 ;
        RECT  12.505 19.645 12.575 19.78 ;
        RECT  12.505 19.645 12.575 19.78 ;
        RECT  12.505 19.645 12.575 19.78 ;
        RECT  12.505 19.645 12.575 19.78 ;
        RECT  12.505 19.645 12.575 19.78 ;
        RECT  12.505 19.645 12.575 19.78 ;
        RECT  12.055 19.1525 12.125 19.2875 ;
        RECT  11.8 19.645 11.87 19.78 ;
        RECT  11.8 19.645 11.87 19.78 ;
        RECT  11.8 19.645 11.87 19.78 ;
        RECT  11.8 19.645 11.87 19.78 ;
        RECT  11.8 19.645 11.87 19.78 ;
        RECT  11.8 19.645 11.87 19.78 ;
        RECT  12.505 19.645 12.575 19.78 ;
        RECT  12.505 19.645 12.575 19.78 ;
        RECT  12.505 19.645 12.575 19.78 ;
        RECT  12.505 19.645 12.575 19.78 ;
        RECT  12.25 19.1525 12.32 19.2875 ;
        RECT  12.4725 18.86 12.6075 18.93 ;
        RECT  12.4725 18.86 12.6075 18.93 ;
        RECT  12.4725 18.86 12.6075 18.93 ;
        RECT  12.505 19.645 12.575 19.78 ;
        RECT  12.505 19.645 12.575 19.78 ;
        RECT  12.505 19.645 12.575 19.78 ;
        RECT  12.505 19.645 12.575 19.78 ;
        RECT  12.505 19.645 12.575 19.78 ;
        RECT  12.505 19.645 12.575 19.78 ;
        RECT  11.7675 18.86 11.9025 18.93 ;
        RECT  12.505 18.8625 12.575 20.2725 ;
        RECT  11.805 18.865 11.865 18.9225 ;
        RECT  11.9925 18.87 12.0475 18.9225 ;
        RECT  12.3275 18.8625 12.385 18.9225 ;
        RECT  12.51 18.87 12.57 18.9275 ;
        RECT  12.32 18.795 12.39 20.34 ;
        RECT  11.985 18.795 12.055 20.34 ;
        RECT  11.8 18.795 11.87 20.34 ;
        RECT  12.505 18.795 12.575 20.34 ;
        RECT  12.505 20.7 12.575 20.835 ;
        RECT  12.505 20.7 12.575 20.835 ;
        RECT  12.505 20.7 12.575 20.835 ;
        RECT  12.505 20.7 12.575 20.835 ;
        RECT  12.505 20.7 12.575 20.835 ;
        RECT  12.505 20.7 12.575 20.835 ;
        RECT  11.7675 21.55 11.9025 21.62 ;
        RECT  12.4725 21.55 12.6075 21.62 ;
        RECT  12.505 20.7 12.575 20.835 ;
        RECT  12.505 20.7 12.575 20.835 ;
        RECT  12.505 20.7 12.575 20.835 ;
        RECT  12.505 20.7 12.575 20.835 ;
        RECT  12.505 20.7 12.575 20.835 ;
        RECT  12.505 20.7 12.575 20.835 ;
        RECT  12.505 20.7 12.575 20.835 ;
        RECT  12.505 20.7 12.575 20.835 ;
        RECT  12.055 21.1925 12.125 21.3275 ;
        RECT  11.8 20.7 11.87 20.835 ;
        RECT  11.8 20.7 11.87 20.835 ;
        RECT  11.8 20.7 11.87 20.835 ;
        RECT  11.8 20.7 11.87 20.835 ;
        RECT  11.8 20.7 11.87 20.835 ;
        RECT  11.8 20.7 11.87 20.835 ;
        RECT  12.505 20.7 12.575 20.835 ;
        RECT  12.505 20.7 12.575 20.835 ;
        RECT  12.505 20.7 12.575 20.835 ;
        RECT  12.505 20.7 12.575 20.835 ;
        RECT  12.25 21.1925 12.32 21.3275 ;
        RECT  12.4725 21.55 12.6075 21.62 ;
        RECT  12.4725 21.55 12.6075 21.62 ;
        RECT  12.4725 21.55 12.6075 21.62 ;
        RECT  12.505 20.7 12.575 20.835 ;
        RECT  12.505 20.7 12.575 20.835 ;
        RECT  12.505 20.7 12.575 20.835 ;
        RECT  12.505 20.7 12.575 20.835 ;
        RECT  12.505 20.7 12.575 20.835 ;
        RECT  12.505 20.7 12.575 20.835 ;
        RECT  11.7675 21.55 11.9025 21.62 ;
        RECT  12.505 20.2075 12.575 21.6175 ;
        RECT  11.805 21.5575 11.865 21.615 ;
        RECT  11.9925 21.5575 12.0475 21.61 ;
        RECT  12.3275 21.5575 12.385 21.6175 ;
        RECT  12.51 21.5525 12.57 21.61 ;
        RECT  12.32 20.14 12.39 21.685 ;
        RECT  11.985 20.14 12.055 21.685 ;
        RECT  11.8 20.14 11.87 21.685 ;
        RECT  12.505 20.14 12.575 21.685 ;
        RECT  12.505 22.335 12.575 22.47 ;
        RECT  12.505 22.335 12.575 22.47 ;
        RECT  12.505 22.335 12.575 22.47 ;
        RECT  12.505 22.335 12.575 22.47 ;
        RECT  12.505 22.335 12.575 22.47 ;
        RECT  12.505 22.335 12.575 22.47 ;
        RECT  11.7675 21.55 11.9025 21.62 ;
        RECT  12.4725 21.55 12.6075 21.62 ;
        RECT  12.505 22.335 12.575 22.47 ;
        RECT  12.505 22.335 12.575 22.47 ;
        RECT  12.505 22.335 12.575 22.47 ;
        RECT  12.505 22.335 12.575 22.47 ;
        RECT  12.505 22.335 12.575 22.47 ;
        RECT  12.505 22.335 12.575 22.47 ;
        RECT  12.505 22.335 12.575 22.47 ;
        RECT  12.505 22.335 12.575 22.47 ;
        RECT  12.055 21.8425 12.125 21.9775 ;
        RECT  11.8 22.335 11.87 22.47 ;
        RECT  11.8 22.335 11.87 22.47 ;
        RECT  11.8 22.335 11.87 22.47 ;
        RECT  11.8 22.335 11.87 22.47 ;
        RECT  11.8 22.335 11.87 22.47 ;
        RECT  11.8 22.335 11.87 22.47 ;
        RECT  12.505 22.335 12.575 22.47 ;
        RECT  12.505 22.335 12.575 22.47 ;
        RECT  12.505 22.335 12.575 22.47 ;
        RECT  12.505 22.335 12.575 22.47 ;
        RECT  12.25 21.8425 12.32 21.9775 ;
        RECT  12.4725 21.55 12.6075 21.62 ;
        RECT  12.4725 21.55 12.6075 21.62 ;
        RECT  12.4725 21.55 12.6075 21.62 ;
        RECT  12.505 22.335 12.575 22.47 ;
        RECT  12.505 22.335 12.575 22.47 ;
        RECT  12.505 22.335 12.575 22.47 ;
        RECT  12.505 22.335 12.575 22.47 ;
        RECT  12.505 22.335 12.575 22.47 ;
        RECT  12.505 22.335 12.575 22.47 ;
        RECT  11.7675 21.55 11.9025 21.62 ;
        RECT  12.505 21.5525 12.575 22.9625 ;
        RECT  11.805 21.555 11.865 21.6125 ;
        RECT  11.9925 21.56 12.0475 21.6125 ;
        RECT  12.3275 21.5525 12.385 21.6125 ;
        RECT  12.51 21.56 12.57 21.6175 ;
        RECT  12.32 21.485 12.39 23.03 ;
        RECT  11.985 21.485 12.055 23.03 ;
        RECT  11.8 21.485 11.87 23.03 ;
        RECT  12.505 21.485 12.575 23.03 ;
        RECT  12.505 23.39 12.575 23.525 ;
        RECT  12.505 23.39 12.575 23.525 ;
        RECT  12.505 23.39 12.575 23.525 ;
        RECT  12.505 23.39 12.575 23.525 ;
        RECT  12.505 23.39 12.575 23.525 ;
        RECT  12.505 23.39 12.575 23.525 ;
        RECT  11.7675 24.24 11.9025 24.31 ;
        RECT  12.4725 24.24 12.6075 24.31 ;
        RECT  12.505 23.39 12.575 23.525 ;
        RECT  12.505 23.39 12.575 23.525 ;
        RECT  12.505 23.39 12.575 23.525 ;
        RECT  12.505 23.39 12.575 23.525 ;
        RECT  12.505 23.39 12.575 23.525 ;
        RECT  12.505 23.39 12.575 23.525 ;
        RECT  12.505 23.39 12.575 23.525 ;
        RECT  12.505 23.39 12.575 23.525 ;
        RECT  12.055 23.8825 12.125 24.0175 ;
        RECT  11.8 23.39 11.87 23.525 ;
        RECT  11.8 23.39 11.87 23.525 ;
        RECT  11.8 23.39 11.87 23.525 ;
        RECT  11.8 23.39 11.87 23.525 ;
        RECT  11.8 23.39 11.87 23.525 ;
        RECT  11.8 23.39 11.87 23.525 ;
        RECT  12.505 23.39 12.575 23.525 ;
        RECT  12.505 23.39 12.575 23.525 ;
        RECT  12.505 23.39 12.575 23.525 ;
        RECT  12.505 23.39 12.575 23.525 ;
        RECT  12.25 23.8825 12.32 24.0175 ;
        RECT  12.4725 24.24 12.6075 24.31 ;
        RECT  12.4725 24.24 12.6075 24.31 ;
        RECT  12.4725 24.24 12.6075 24.31 ;
        RECT  12.505 23.39 12.575 23.525 ;
        RECT  12.505 23.39 12.575 23.525 ;
        RECT  12.505 23.39 12.575 23.525 ;
        RECT  12.505 23.39 12.575 23.525 ;
        RECT  12.505 23.39 12.575 23.525 ;
        RECT  12.505 23.39 12.575 23.525 ;
        RECT  11.7675 24.24 11.9025 24.31 ;
        RECT  12.505 22.8975 12.575 24.3075 ;
        RECT  11.805 24.2475 11.865 24.305 ;
        RECT  11.9925 24.2475 12.0475 24.3 ;
        RECT  12.3275 24.2475 12.385 24.3075 ;
        RECT  12.51 24.2425 12.57 24.3 ;
        RECT  12.32 22.83 12.39 24.375 ;
        RECT  11.985 22.83 12.055 24.375 ;
        RECT  11.8 22.83 11.87 24.375 ;
        RECT  12.505 22.83 12.575 24.375 ;
        RECT  12.505 25.025 12.575 25.16 ;
        RECT  12.505 25.025 12.575 25.16 ;
        RECT  12.505 25.025 12.575 25.16 ;
        RECT  12.505 25.025 12.575 25.16 ;
        RECT  12.505 25.025 12.575 25.16 ;
        RECT  12.505 25.025 12.575 25.16 ;
        RECT  11.7675 24.24 11.9025 24.31 ;
        RECT  12.4725 24.24 12.6075 24.31 ;
        RECT  12.505 25.025 12.575 25.16 ;
        RECT  12.505 25.025 12.575 25.16 ;
        RECT  12.505 25.025 12.575 25.16 ;
        RECT  12.505 25.025 12.575 25.16 ;
        RECT  12.505 25.025 12.575 25.16 ;
        RECT  12.505 25.025 12.575 25.16 ;
        RECT  12.505 25.025 12.575 25.16 ;
        RECT  12.505 25.025 12.575 25.16 ;
        RECT  12.055 24.5325 12.125 24.6675 ;
        RECT  11.8 25.025 11.87 25.16 ;
        RECT  11.8 25.025 11.87 25.16 ;
        RECT  11.8 25.025 11.87 25.16 ;
        RECT  11.8 25.025 11.87 25.16 ;
        RECT  11.8 25.025 11.87 25.16 ;
        RECT  11.8 25.025 11.87 25.16 ;
        RECT  12.505 25.025 12.575 25.16 ;
        RECT  12.505 25.025 12.575 25.16 ;
        RECT  12.505 25.025 12.575 25.16 ;
        RECT  12.505 25.025 12.575 25.16 ;
        RECT  12.25 24.5325 12.32 24.6675 ;
        RECT  12.4725 24.24 12.6075 24.31 ;
        RECT  12.4725 24.24 12.6075 24.31 ;
        RECT  12.4725 24.24 12.6075 24.31 ;
        RECT  12.505 25.025 12.575 25.16 ;
        RECT  12.505 25.025 12.575 25.16 ;
        RECT  12.505 25.025 12.575 25.16 ;
        RECT  12.505 25.025 12.575 25.16 ;
        RECT  12.505 25.025 12.575 25.16 ;
        RECT  12.505 25.025 12.575 25.16 ;
        RECT  11.7675 24.24 11.9025 24.31 ;
        RECT  12.505 24.2425 12.575 25.6525 ;
        RECT  11.805 24.245 11.865 24.3025 ;
        RECT  11.9925 24.25 12.0475 24.3025 ;
        RECT  12.3275 24.2425 12.385 24.3025 ;
        RECT  12.51 24.25 12.57 24.3075 ;
        RECT  12.32 24.175 12.39 25.72 ;
        RECT  11.985 24.175 12.055 25.72 ;
        RECT  11.8 24.175 11.87 25.72 ;
        RECT  12.505 24.175 12.575 25.72 ;
        RECT  12.505 26.08 12.575 26.215 ;
        RECT  12.505 26.08 12.575 26.215 ;
        RECT  12.505 26.08 12.575 26.215 ;
        RECT  12.505 26.08 12.575 26.215 ;
        RECT  12.505 26.08 12.575 26.215 ;
        RECT  12.505 26.08 12.575 26.215 ;
        RECT  11.7675 26.93 11.9025 27.0 ;
        RECT  12.4725 26.93 12.6075 27.0 ;
        RECT  12.505 26.08 12.575 26.215 ;
        RECT  12.505 26.08 12.575 26.215 ;
        RECT  12.505 26.08 12.575 26.215 ;
        RECT  12.505 26.08 12.575 26.215 ;
        RECT  12.505 26.08 12.575 26.215 ;
        RECT  12.505 26.08 12.575 26.215 ;
        RECT  12.505 26.08 12.575 26.215 ;
        RECT  12.505 26.08 12.575 26.215 ;
        RECT  12.055 26.5725 12.125 26.7075 ;
        RECT  11.8 26.08 11.87 26.215 ;
        RECT  11.8 26.08 11.87 26.215 ;
        RECT  11.8 26.08 11.87 26.215 ;
        RECT  11.8 26.08 11.87 26.215 ;
        RECT  11.8 26.08 11.87 26.215 ;
        RECT  11.8 26.08 11.87 26.215 ;
        RECT  12.505 26.08 12.575 26.215 ;
        RECT  12.505 26.08 12.575 26.215 ;
        RECT  12.505 26.08 12.575 26.215 ;
        RECT  12.505 26.08 12.575 26.215 ;
        RECT  12.25 26.5725 12.32 26.7075 ;
        RECT  12.4725 26.93 12.6075 27.0 ;
        RECT  12.4725 26.93 12.6075 27.0 ;
        RECT  12.4725 26.93 12.6075 27.0 ;
        RECT  12.505 26.08 12.575 26.215 ;
        RECT  12.505 26.08 12.575 26.215 ;
        RECT  12.505 26.08 12.575 26.215 ;
        RECT  12.505 26.08 12.575 26.215 ;
        RECT  12.505 26.08 12.575 26.215 ;
        RECT  12.505 26.08 12.575 26.215 ;
        RECT  11.7675 26.93 11.9025 27.0 ;
        RECT  12.505 25.5875 12.575 26.9975 ;
        RECT  11.805 26.9375 11.865 26.995 ;
        RECT  11.9925 26.9375 12.0475 26.99 ;
        RECT  12.3275 26.9375 12.385 26.9975 ;
        RECT  12.51 26.9325 12.57 26.99 ;
        RECT  12.32 25.52 12.39 27.065 ;
        RECT  11.985 25.52 12.055 27.065 ;
        RECT  11.8 25.52 11.87 27.065 ;
        RECT  12.505 25.52 12.575 27.065 ;
        RECT  12.505 27.715 12.575 27.85 ;
        RECT  12.505 27.715 12.575 27.85 ;
        RECT  12.505 27.715 12.575 27.85 ;
        RECT  12.505 27.715 12.575 27.85 ;
        RECT  12.505 27.715 12.575 27.85 ;
        RECT  12.505 27.715 12.575 27.85 ;
        RECT  11.7675 26.93 11.9025 27.0 ;
        RECT  12.4725 26.93 12.6075 27.0 ;
        RECT  12.505 27.715 12.575 27.85 ;
        RECT  12.505 27.715 12.575 27.85 ;
        RECT  12.505 27.715 12.575 27.85 ;
        RECT  12.505 27.715 12.575 27.85 ;
        RECT  12.505 27.715 12.575 27.85 ;
        RECT  12.505 27.715 12.575 27.85 ;
        RECT  12.505 27.715 12.575 27.85 ;
        RECT  12.505 27.715 12.575 27.85 ;
        RECT  12.055 27.2225 12.125 27.3575 ;
        RECT  11.8 27.715 11.87 27.85 ;
        RECT  11.8 27.715 11.87 27.85 ;
        RECT  11.8 27.715 11.87 27.85 ;
        RECT  11.8 27.715 11.87 27.85 ;
        RECT  11.8 27.715 11.87 27.85 ;
        RECT  11.8 27.715 11.87 27.85 ;
        RECT  12.505 27.715 12.575 27.85 ;
        RECT  12.505 27.715 12.575 27.85 ;
        RECT  12.505 27.715 12.575 27.85 ;
        RECT  12.505 27.715 12.575 27.85 ;
        RECT  12.25 27.2225 12.32 27.3575 ;
        RECT  12.4725 26.93 12.6075 27.0 ;
        RECT  12.4725 26.93 12.6075 27.0 ;
        RECT  12.4725 26.93 12.6075 27.0 ;
        RECT  12.505 27.715 12.575 27.85 ;
        RECT  12.505 27.715 12.575 27.85 ;
        RECT  12.505 27.715 12.575 27.85 ;
        RECT  12.505 27.715 12.575 27.85 ;
        RECT  12.505 27.715 12.575 27.85 ;
        RECT  12.505 27.715 12.575 27.85 ;
        RECT  11.7675 26.93 11.9025 27.0 ;
        RECT  12.505 26.9325 12.575 28.3425 ;
        RECT  11.805 26.935 11.865 26.9925 ;
        RECT  11.9925 26.94 12.0475 26.9925 ;
        RECT  12.3275 26.9325 12.385 26.9925 ;
        RECT  12.51 26.94 12.57 26.9975 ;
        RECT  12.32 26.865 12.39 28.41 ;
        RECT  11.985 26.865 12.055 28.41 ;
        RECT  11.8 26.865 11.87 28.41 ;
        RECT  12.505 26.865 12.575 28.41 ;
        RECT  12.505 28.77 12.575 28.905 ;
        RECT  12.505 28.77 12.575 28.905 ;
        RECT  12.505 28.77 12.575 28.905 ;
        RECT  12.505 28.77 12.575 28.905 ;
        RECT  12.505 28.77 12.575 28.905 ;
        RECT  12.505 28.77 12.575 28.905 ;
        RECT  11.7675 29.62 11.9025 29.69 ;
        RECT  12.4725 29.62 12.6075 29.69 ;
        RECT  12.505 28.77 12.575 28.905 ;
        RECT  12.505 28.77 12.575 28.905 ;
        RECT  12.505 28.77 12.575 28.905 ;
        RECT  12.505 28.77 12.575 28.905 ;
        RECT  12.505 28.77 12.575 28.905 ;
        RECT  12.505 28.77 12.575 28.905 ;
        RECT  12.505 28.77 12.575 28.905 ;
        RECT  12.505 28.77 12.575 28.905 ;
        RECT  12.055 29.2625 12.125 29.3975 ;
        RECT  11.8 28.77 11.87 28.905 ;
        RECT  11.8 28.77 11.87 28.905 ;
        RECT  11.8 28.77 11.87 28.905 ;
        RECT  11.8 28.77 11.87 28.905 ;
        RECT  11.8 28.77 11.87 28.905 ;
        RECT  11.8 28.77 11.87 28.905 ;
        RECT  12.505 28.77 12.575 28.905 ;
        RECT  12.505 28.77 12.575 28.905 ;
        RECT  12.505 28.77 12.575 28.905 ;
        RECT  12.505 28.77 12.575 28.905 ;
        RECT  12.25 29.2625 12.32 29.3975 ;
        RECT  12.4725 29.62 12.6075 29.69 ;
        RECT  12.4725 29.62 12.6075 29.69 ;
        RECT  12.4725 29.62 12.6075 29.69 ;
        RECT  12.505 28.77 12.575 28.905 ;
        RECT  12.505 28.77 12.575 28.905 ;
        RECT  12.505 28.77 12.575 28.905 ;
        RECT  12.505 28.77 12.575 28.905 ;
        RECT  12.505 28.77 12.575 28.905 ;
        RECT  12.505 28.77 12.575 28.905 ;
        RECT  11.7675 29.62 11.9025 29.69 ;
        RECT  12.505 28.2775 12.575 29.6875 ;
        RECT  11.805 29.6275 11.865 29.685 ;
        RECT  11.9925 29.6275 12.0475 29.68 ;
        RECT  12.3275 29.6275 12.385 29.6875 ;
        RECT  12.51 29.6225 12.57 29.68 ;
        RECT  12.32 28.21 12.39 29.755 ;
        RECT  11.985 28.21 12.055 29.755 ;
        RECT  11.8 28.21 11.87 29.755 ;
        RECT  12.505 28.21 12.575 29.755 ;
        RECT  12.505 30.405 12.575 30.54 ;
        RECT  12.505 30.405 12.575 30.54 ;
        RECT  12.505 30.405 12.575 30.54 ;
        RECT  12.505 30.405 12.575 30.54 ;
        RECT  12.505 30.405 12.575 30.54 ;
        RECT  12.505 30.405 12.575 30.54 ;
        RECT  11.7675 29.62 11.9025 29.69 ;
        RECT  12.4725 29.62 12.6075 29.69 ;
        RECT  12.505 30.405 12.575 30.54 ;
        RECT  12.505 30.405 12.575 30.54 ;
        RECT  12.505 30.405 12.575 30.54 ;
        RECT  12.505 30.405 12.575 30.54 ;
        RECT  12.505 30.405 12.575 30.54 ;
        RECT  12.505 30.405 12.575 30.54 ;
        RECT  12.505 30.405 12.575 30.54 ;
        RECT  12.505 30.405 12.575 30.54 ;
        RECT  12.055 29.9125 12.125 30.0475 ;
        RECT  11.8 30.405 11.87 30.54 ;
        RECT  11.8 30.405 11.87 30.54 ;
        RECT  11.8 30.405 11.87 30.54 ;
        RECT  11.8 30.405 11.87 30.54 ;
        RECT  11.8 30.405 11.87 30.54 ;
        RECT  11.8 30.405 11.87 30.54 ;
        RECT  12.505 30.405 12.575 30.54 ;
        RECT  12.505 30.405 12.575 30.54 ;
        RECT  12.505 30.405 12.575 30.54 ;
        RECT  12.505 30.405 12.575 30.54 ;
        RECT  12.25 29.9125 12.32 30.0475 ;
        RECT  12.4725 29.62 12.6075 29.69 ;
        RECT  12.4725 29.62 12.6075 29.69 ;
        RECT  12.4725 29.62 12.6075 29.69 ;
        RECT  12.505 30.405 12.575 30.54 ;
        RECT  12.505 30.405 12.575 30.54 ;
        RECT  12.505 30.405 12.575 30.54 ;
        RECT  12.505 30.405 12.575 30.54 ;
        RECT  12.505 30.405 12.575 30.54 ;
        RECT  12.505 30.405 12.575 30.54 ;
        RECT  11.7675 29.62 11.9025 29.69 ;
        RECT  12.505 29.6225 12.575 31.0325 ;
        RECT  11.805 29.625 11.865 29.6825 ;
        RECT  11.9925 29.63 12.0475 29.6825 ;
        RECT  12.3275 29.6225 12.385 29.6825 ;
        RECT  12.51 29.63 12.57 29.6875 ;
        RECT  12.32 29.555 12.39 31.1 ;
        RECT  11.985 29.555 12.055 31.1 ;
        RECT  11.8 29.555 11.87 31.1 ;
        RECT  12.505 29.555 12.575 31.1 ;
        RECT  12.505 31.46 12.575 31.595 ;
        RECT  12.505 31.46 12.575 31.595 ;
        RECT  12.505 31.46 12.575 31.595 ;
        RECT  12.505 31.46 12.575 31.595 ;
        RECT  12.505 31.46 12.575 31.595 ;
        RECT  12.505 31.46 12.575 31.595 ;
        RECT  11.7675 32.31 11.9025 32.38 ;
        RECT  12.4725 32.31 12.6075 32.38 ;
        RECT  12.505 31.46 12.575 31.595 ;
        RECT  12.505 31.46 12.575 31.595 ;
        RECT  12.505 31.46 12.575 31.595 ;
        RECT  12.505 31.46 12.575 31.595 ;
        RECT  12.505 31.46 12.575 31.595 ;
        RECT  12.505 31.46 12.575 31.595 ;
        RECT  12.505 31.46 12.575 31.595 ;
        RECT  12.505 31.46 12.575 31.595 ;
        RECT  12.055 31.9525 12.125 32.0875 ;
        RECT  11.8 31.46 11.87 31.595 ;
        RECT  11.8 31.46 11.87 31.595 ;
        RECT  11.8 31.46 11.87 31.595 ;
        RECT  11.8 31.46 11.87 31.595 ;
        RECT  11.8 31.46 11.87 31.595 ;
        RECT  11.8 31.46 11.87 31.595 ;
        RECT  12.505 31.46 12.575 31.595 ;
        RECT  12.505 31.46 12.575 31.595 ;
        RECT  12.505 31.46 12.575 31.595 ;
        RECT  12.505 31.46 12.575 31.595 ;
        RECT  12.25 31.9525 12.32 32.0875 ;
        RECT  12.4725 32.31 12.6075 32.38 ;
        RECT  12.4725 32.31 12.6075 32.38 ;
        RECT  12.4725 32.31 12.6075 32.38 ;
        RECT  12.505 31.46 12.575 31.595 ;
        RECT  12.505 31.46 12.575 31.595 ;
        RECT  12.505 31.46 12.575 31.595 ;
        RECT  12.505 31.46 12.575 31.595 ;
        RECT  12.505 31.46 12.575 31.595 ;
        RECT  12.505 31.46 12.575 31.595 ;
        RECT  11.7675 32.31 11.9025 32.38 ;
        RECT  12.505 30.9675 12.575 32.3775 ;
        RECT  11.805 32.3175 11.865 32.375 ;
        RECT  11.9925 32.3175 12.0475 32.37 ;
        RECT  12.3275 32.3175 12.385 32.3775 ;
        RECT  12.51 32.3125 12.57 32.37 ;
        RECT  12.32 30.9 12.39 32.445 ;
        RECT  11.985 30.9 12.055 32.445 ;
        RECT  11.8 30.9 11.87 32.445 ;
        RECT  12.505 30.9 12.575 32.445 ;
        RECT  12.505 33.095 12.575 33.23 ;
        RECT  12.505 33.095 12.575 33.23 ;
        RECT  12.505 33.095 12.575 33.23 ;
        RECT  12.505 33.095 12.575 33.23 ;
        RECT  12.505 33.095 12.575 33.23 ;
        RECT  12.505 33.095 12.575 33.23 ;
        RECT  11.7675 32.31 11.9025 32.38 ;
        RECT  12.4725 32.31 12.6075 32.38 ;
        RECT  12.505 33.095 12.575 33.23 ;
        RECT  12.505 33.095 12.575 33.23 ;
        RECT  12.505 33.095 12.575 33.23 ;
        RECT  12.505 33.095 12.575 33.23 ;
        RECT  12.505 33.095 12.575 33.23 ;
        RECT  12.505 33.095 12.575 33.23 ;
        RECT  12.505 33.095 12.575 33.23 ;
        RECT  12.505 33.095 12.575 33.23 ;
        RECT  12.055 32.6025 12.125 32.7375 ;
        RECT  11.8 33.095 11.87 33.23 ;
        RECT  11.8 33.095 11.87 33.23 ;
        RECT  11.8 33.095 11.87 33.23 ;
        RECT  11.8 33.095 11.87 33.23 ;
        RECT  11.8 33.095 11.87 33.23 ;
        RECT  11.8 33.095 11.87 33.23 ;
        RECT  12.505 33.095 12.575 33.23 ;
        RECT  12.505 33.095 12.575 33.23 ;
        RECT  12.505 33.095 12.575 33.23 ;
        RECT  12.505 33.095 12.575 33.23 ;
        RECT  12.25 32.6025 12.32 32.7375 ;
        RECT  12.4725 32.31 12.6075 32.38 ;
        RECT  12.4725 32.31 12.6075 32.38 ;
        RECT  12.4725 32.31 12.6075 32.38 ;
        RECT  12.505 33.095 12.575 33.23 ;
        RECT  12.505 33.095 12.575 33.23 ;
        RECT  12.505 33.095 12.575 33.23 ;
        RECT  12.505 33.095 12.575 33.23 ;
        RECT  12.505 33.095 12.575 33.23 ;
        RECT  12.505 33.095 12.575 33.23 ;
        RECT  11.7675 32.31 11.9025 32.38 ;
        RECT  12.505 32.3125 12.575 33.7225 ;
        RECT  11.805 32.315 11.865 32.3725 ;
        RECT  11.9925 32.32 12.0475 32.3725 ;
        RECT  12.3275 32.3125 12.385 32.3725 ;
        RECT  12.51 32.32 12.57 32.3775 ;
        RECT  12.32 32.245 12.39 33.79 ;
        RECT  11.985 32.245 12.055 33.79 ;
        RECT  11.8 32.245 11.87 33.79 ;
        RECT  12.505 32.245 12.575 33.79 ;
        RECT  12.505 34.15 12.575 34.285 ;
        RECT  12.505 34.15 12.575 34.285 ;
        RECT  12.505 34.15 12.575 34.285 ;
        RECT  12.505 34.15 12.575 34.285 ;
        RECT  12.505 34.15 12.575 34.285 ;
        RECT  12.505 34.15 12.575 34.285 ;
        RECT  11.7675 35.0 11.9025 35.07 ;
        RECT  12.4725 35.0 12.6075 35.07 ;
        RECT  12.505 34.15 12.575 34.285 ;
        RECT  12.505 34.15 12.575 34.285 ;
        RECT  12.505 34.15 12.575 34.285 ;
        RECT  12.505 34.15 12.575 34.285 ;
        RECT  12.505 34.15 12.575 34.285 ;
        RECT  12.505 34.15 12.575 34.285 ;
        RECT  12.505 34.15 12.575 34.285 ;
        RECT  12.505 34.15 12.575 34.285 ;
        RECT  12.055 34.6425 12.125 34.7775 ;
        RECT  11.8 34.15 11.87 34.285 ;
        RECT  11.8 34.15 11.87 34.285 ;
        RECT  11.8 34.15 11.87 34.285 ;
        RECT  11.8 34.15 11.87 34.285 ;
        RECT  11.8 34.15 11.87 34.285 ;
        RECT  11.8 34.15 11.87 34.285 ;
        RECT  12.505 34.15 12.575 34.285 ;
        RECT  12.505 34.15 12.575 34.285 ;
        RECT  12.505 34.15 12.575 34.285 ;
        RECT  12.505 34.15 12.575 34.285 ;
        RECT  12.25 34.6425 12.32 34.7775 ;
        RECT  12.4725 35.0 12.6075 35.07 ;
        RECT  12.4725 35.0 12.6075 35.07 ;
        RECT  12.4725 35.0 12.6075 35.07 ;
        RECT  12.505 34.15 12.575 34.285 ;
        RECT  12.505 34.15 12.575 34.285 ;
        RECT  12.505 34.15 12.575 34.285 ;
        RECT  12.505 34.15 12.575 34.285 ;
        RECT  12.505 34.15 12.575 34.285 ;
        RECT  12.505 34.15 12.575 34.285 ;
        RECT  11.7675 35.0 11.9025 35.07 ;
        RECT  12.505 33.6575 12.575 35.0675 ;
        RECT  11.805 35.0075 11.865 35.065 ;
        RECT  11.9925 35.0075 12.0475 35.06 ;
        RECT  12.3275 35.0075 12.385 35.0675 ;
        RECT  12.51 35.0025 12.57 35.06 ;
        RECT  12.32 33.59 12.39 35.135 ;
        RECT  11.985 33.59 12.055 35.135 ;
        RECT  11.8 33.59 11.87 35.135 ;
        RECT  12.505 33.59 12.575 35.135 ;
        RECT  12.505 35.785 12.575 35.92 ;
        RECT  12.505 35.785 12.575 35.92 ;
        RECT  12.505 35.785 12.575 35.92 ;
        RECT  12.505 35.785 12.575 35.92 ;
        RECT  12.505 35.785 12.575 35.92 ;
        RECT  12.505 35.785 12.575 35.92 ;
        RECT  11.7675 35.0 11.9025 35.07 ;
        RECT  12.4725 35.0 12.6075 35.07 ;
        RECT  12.505 35.785 12.575 35.92 ;
        RECT  12.505 35.785 12.575 35.92 ;
        RECT  12.505 35.785 12.575 35.92 ;
        RECT  12.505 35.785 12.575 35.92 ;
        RECT  12.505 35.785 12.575 35.92 ;
        RECT  12.505 35.785 12.575 35.92 ;
        RECT  12.505 35.785 12.575 35.92 ;
        RECT  12.505 35.785 12.575 35.92 ;
        RECT  12.055 35.2925 12.125 35.4275 ;
        RECT  11.8 35.785 11.87 35.92 ;
        RECT  11.8 35.785 11.87 35.92 ;
        RECT  11.8 35.785 11.87 35.92 ;
        RECT  11.8 35.785 11.87 35.92 ;
        RECT  11.8 35.785 11.87 35.92 ;
        RECT  11.8 35.785 11.87 35.92 ;
        RECT  12.505 35.785 12.575 35.92 ;
        RECT  12.505 35.785 12.575 35.92 ;
        RECT  12.505 35.785 12.575 35.92 ;
        RECT  12.505 35.785 12.575 35.92 ;
        RECT  12.25 35.2925 12.32 35.4275 ;
        RECT  12.4725 35.0 12.6075 35.07 ;
        RECT  12.4725 35.0 12.6075 35.07 ;
        RECT  12.4725 35.0 12.6075 35.07 ;
        RECT  12.505 35.785 12.575 35.92 ;
        RECT  12.505 35.785 12.575 35.92 ;
        RECT  12.505 35.785 12.575 35.92 ;
        RECT  12.505 35.785 12.575 35.92 ;
        RECT  12.505 35.785 12.575 35.92 ;
        RECT  12.505 35.785 12.575 35.92 ;
        RECT  11.7675 35.0 11.9025 35.07 ;
        RECT  12.505 35.0025 12.575 36.4125 ;
        RECT  11.805 35.005 11.865 35.0625 ;
        RECT  11.9925 35.01 12.0475 35.0625 ;
        RECT  12.3275 35.0025 12.385 35.0625 ;
        RECT  12.51 35.01 12.57 35.0675 ;
        RECT  12.32 34.935 12.39 36.48 ;
        RECT  11.985 34.935 12.055 36.48 ;
        RECT  11.8 34.935 11.87 36.48 ;
        RECT  12.505 34.935 12.575 36.48 ;
        RECT  12.505 36.84 12.575 36.975 ;
        RECT  12.505 36.84 12.575 36.975 ;
        RECT  12.505 36.84 12.575 36.975 ;
        RECT  12.505 36.84 12.575 36.975 ;
        RECT  12.505 36.84 12.575 36.975 ;
        RECT  12.505 36.84 12.575 36.975 ;
        RECT  11.7675 37.69 11.9025 37.76 ;
        RECT  12.4725 37.69 12.6075 37.76 ;
        RECT  12.505 36.84 12.575 36.975 ;
        RECT  12.505 36.84 12.575 36.975 ;
        RECT  12.505 36.84 12.575 36.975 ;
        RECT  12.505 36.84 12.575 36.975 ;
        RECT  12.505 36.84 12.575 36.975 ;
        RECT  12.505 36.84 12.575 36.975 ;
        RECT  12.505 36.84 12.575 36.975 ;
        RECT  12.505 36.84 12.575 36.975 ;
        RECT  12.055 37.3325 12.125 37.4675 ;
        RECT  11.8 36.84 11.87 36.975 ;
        RECT  11.8 36.84 11.87 36.975 ;
        RECT  11.8 36.84 11.87 36.975 ;
        RECT  11.8 36.84 11.87 36.975 ;
        RECT  11.8 36.84 11.87 36.975 ;
        RECT  11.8 36.84 11.87 36.975 ;
        RECT  12.505 36.84 12.575 36.975 ;
        RECT  12.505 36.84 12.575 36.975 ;
        RECT  12.505 36.84 12.575 36.975 ;
        RECT  12.505 36.84 12.575 36.975 ;
        RECT  12.25 37.3325 12.32 37.4675 ;
        RECT  12.4725 37.69 12.6075 37.76 ;
        RECT  12.4725 37.69 12.6075 37.76 ;
        RECT  12.4725 37.69 12.6075 37.76 ;
        RECT  12.505 36.84 12.575 36.975 ;
        RECT  12.505 36.84 12.575 36.975 ;
        RECT  12.505 36.84 12.575 36.975 ;
        RECT  12.505 36.84 12.575 36.975 ;
        RECT  12.505 36.84 12.575 36.975 ;
        RECT  12.505 36.84 12.575 36.975 ;
        RECT  11.7675 37.69 11.9025 37.76 ;
        RECT  12.505 36.3475 12.575 37.7575 ;
        RECT  11.805 37.6975 11.865 37.755 ;
        RECT  11.9925 37.6975 12.0475 37.75 ;
        RECT  12.3275 37.6975 12.385 37.7575 ;
        RECT  12.51 37.6925 12.57 37.75 ;
        RECT  12.32 36.28 12.39 37.825 ;
        RECT  11.985 36.28 12.055 37.825 ;
        RECT  11.8 36.28 11.87 37.825 ;
        RECT  12.505 36.28 12.575 37.825 ;
        RECT  12.505 38.475 12.575 38.61 ;
        RECT  12.505 38.475 12.575 38.61 ;
        RECT  12.505 38.475 12.575 38.61 ;
        RECT  12.505 38.475 12.575 38.61 ;
        RECT  12.505 38.475 12.575 38.61 ;
        RECT  12.505 38.475 12.575 38.61 ;
        RECT  11.7675 37.69 11.9025 37.76 ;
        RECT  12.4725 37.69 12.6075 37.76 ;
        RECT  12.505 38.475 12.575 38.61 ;
        RECT  12.505 38.475 12.575 38.61 ;
        RECT  12.505 38.475 12.575 38.61 ;
        RECT  12.505 38.475 12.575 38.61 ;
        RECT  12.505 38.475 12.575 38.61 ;
        RECT  12.505 38.475 12.575 38.61 ;
        RECT  12.505 38.475 12.575 38.61 ;
        RECT  12.505 38.475 12.575 38.61 ;
        RECT  12.055 37.9825 12.125 38.1175 ;
        RECT  11.8 38.475 11.87 38.61 ;
        RECT  11.8 38.475 11.87 38.61 ;
        RECT  11.8 38.475 11.87 38.61 ;
        RECT  11.8 38.475 11.87 38.61 ;
        RECT  11.8 38.475 11.87 38.61 ;
        RECT  11.8 38.475 11.87 38.61 ;
        RECT  12.505 38.475 12.575 38.61 ;
        RECT  12.505 38.475 12.575 38.61 ;
        RECT  12.505 38.475 12.575 38.61 ;
        RECT  12.505 38.475 12.575 38.61 ;
        RECT  12.25 37.9825 12.32 38.1175 ;
        RECT  12.4725 37.69 12.6075 37.76 ;
        RECT  12.4725 37.69 12.6075 37.76 ;
        RECT  12.4725 37.69 12.6075 37.76 ;
        RECT  12.505 38.475 12.575 38.61 ;
        RECT  12.505 38.475 12.575 38.61 ;
        RECT  12.505 38.475 12.575 38.61 ;
        RECT  12.505 38.475 12.575 38.61 ;
        RECT  12.505 38.475 12.575 38.61 ;
        RECT  12.505 38.475 12.575 38.61 ;
        RECT  11.7675 37.69 11.9025 37.76 ;
        RECT  12.505 37.6925 12.575 39.1025 ;
        RECT  11.805 37.695 11.865 37.7525 ;
        RECT  11.9925 37.7 12.0475 37.7525 ;
        RECT  12.3275 37.6925 12.385 37.7525 ;
        RECT  12.51 37.7 12.57 37.7575 ;
        RECT  12.32 37.625 12.39 39.17 ;
        RECT  11.985 37.625 12.055 39.17 ;
        RECT  11.8 37.625 11.87 39.17 ;
        RECT  12.505 37.625 12.575 39.17 ;
        RECT  12.505 39.53 12.575 39.665 ;
        RECT  12.505 39.53 12.575 39.665 ;
        RECT  12.505 39.53 12.575 39.665 ;
        RECT  12.505 39.53 12.575 39.665 ;
        RECT  12.505 39.53 12.575 39.665 ;
        RECT  12.505 39.53 12.575 39.665 ;
        RECT  11.7675 40.38 11.9025 40.45 ;
        RECT  12.4725 40.38 12.6075 40.45 ;
        RECT  12.505 39.53 12.575 39.665 ;
        RECT  12.505 39.53 12.575 39.665 ;
        RECT  12.505 39.53 12.575 39.665 ;
        RECT  12.505 39.53 12.575 39.665 ;
        RECT  12.505 39.53 12.575 39.665 ;
        RECT  12.505 39.53 12.575 39.665 ;
        RECT  12.505 39.53 12.575 39.665 ;
        RECT  12.505 39.53 12.575 39.665 ;
        RECT  12.055 40.0225 12.125 40.1575 ;
        RECT  11.8 39.53 11.87 39.665 ;
        RECT  11.8 39.53 11.87 39.665 ;
        RECT  11.8 39.53 11.87 39.665 ;
        RECT  11.8 39.53 11.87 39.665 ;
        RECT  11.8 39.53 11.87 39.665 ;
        RECT  11.8 39.53 11.87 39.665 ;
        RECT  12.505 39.53 12.575 39.665 ;
        RECT  12.505 39.53 12.575 39.665 ;
        RECT  12.505 39.53 12.575 39.665 ;
        RECT  12.505 39.53 12.575 39.665 ;
        RECT  12.25 40.0225 12.32 40.1575 ;
        RECT  12.4725 40.38 12.6075 40.45 ;
        RECT  12.4725 40.38 12.6075 40.45 ;
        RECT  12.4725 40.38 12.6075 40.45 ;
        RECT  12.505 39.53 12.575 39.665 ;
        RECT  12.505 39.53 12.575 39.665 ;
        RECT  12.505 39.53 12.575 39.665 ;
        RECT  12.505 39.53 12.575 39.665 ;
        RECT  12.505 39.53 12.575 39.665 ;
        RECT  12.505 39.53 12.575 39.665 ;
        RECT  11.7675 40.38 11.9025 40.45 ;
        RECT  12.505 39.0375 12.575 40.4475 ;
        RECT  11.805 40.3875 11.865 40.445 ;
        RECT  11.9925 40.3875 12.0475 40.44 ;
        RECT  12.3275 40.3875 12.385 40.4475 ;
        RECT  12.51 40.3825 12.57 40.44 ;
        RECT  12.32 38.97 12.39 40.515 ;
        RECT  11.985 38.97 12.055 40.515 ;
        RECT  11.8 38.97 11.87 40.515 ;
        RECT  12.505 38.97 12.575 40.515 ;
        RECT  11.28 40.765 11.35 41.725 ;
        RECT  11.615 40.765 11.685 41.725 ;
        RECT  11.315 41.3125 11.3575 41.4475 ;
        RECT  11.615 41.3125 11.7025 41.4475 ;
        RECT  11.315 40.8625 11.36 40.9975 ;
        RECT  11.515 40.8625 11.615 40.9975 ;
        RECT  11.3225 41.3125 11.3925 41.4475 ;
        RECT  11.7025 41.3125 11.7725 41.4475 ;
        RECT  11.3225 40.8625 11.3925 40.9975 ;
        RECT  11.5125 40.8625 11.5825 40.9975 ;
        RECT  11.985 40.765 12.055 41.725 ;
        RECT  12.32 40.765 12.39 41.725 ;
        RECT  12.02 41.3125 12.0625 41.4475 ;
        RECT  12.32 41.3125 12.4075 41.4475 ;
        RECT  12.02 40.8625 12.065 40.9975 ;
        RECT  12.22 40.8625 12.32 40.9975 ;
        RECT  12.0275 41.3125 12.0975 41.4475 ;
        RECT  12.4075 41.3125 12.4775 41.4475 ;
        RECT  12.0275 40.8625 12.0975 40.9975 ;
        RECT  12.2175 40.8625 12.2875 40.9975 ;
        RECT  11.4425 18.755 11.5125 18.895 ;
        RECT  11.4425 18.4975 11.5125 18.6325 ;
        RECT  11.8 14.2575 11.87 14.3925 ;
        RECT  11.095 14.2575 11.165 14.3925 ;
        RECT  11.6375 17.04 11.7075 17.175 ;
        RECT  11.255 17.45 11.325 17.585 ;
        RECT  11.4475 18.2925 11.5175 18.4275 ;
        RECT  11.4475 16.15 11.5175 16.285 ;
        RECT  11.4425 18.4975 11.5125 18.895 ;
        RECT  11.4425 18.84 11.5125 18.895 ;
        RECT  11.28 18.835 11.35 18.895 ;
        RECT  11.62 18.845 11.68 18.895 ;
        RECT  11.8 14.01 11.87 18.895 ;
        RECT  11.615 14.81 11.685 18.895 ;
        RECT  11.4475 16.285 11.5175 18.295 ;
        RECT  11.615 14.01 11.685 17.555 ;
        RECT  11.28 14.01 11.35 18.895 ;
        RECT  11.095 14.01 11.165 18.895 ;
        RECT  12.1475 18.755 12.2175 18.895 ;
        RECT  12.1475 18.4975 12.2175 18.6325 ;
        RECT  12.505 14.2575 12.575 14.3925 ;
        RECT  11.8 14.2575 11.87 14.3925 ;
        RECT  12.3425 17.04 12.4125 17.175 ;
        RECT  11.96 17.45 12.03 17.585 ;
        RECT  12.1525 18.2925 12.2225 18.4275 ;
        RECT  12.1525 16.15 12.2225 16.285 ;
        RECT  12.1475 18.4975 12.2175 18.895 ;
        RECT  12.1475 18.84 12.2175 18.895 ;
        RECT  11.985 18.835 12.055 18.895 ;
        RECT  12.325 18.845 12.385 18.895 ;
        RECT  12.505 14.01 12.575 18.895 ;
        RECT  12.32 14.81 12.39 18.895 ;
        RECT  12.1525 16.285 12.2225 18.295 ;
        RECT  12.32 14.01 12.39 17.555 ;
        RECT  11.985 14.01 12.055 18.895 ;
        RECT  11.8 14.01 11.87 18.895 ;
        RECT  11.3375 9.9675 11.4725 10.0375 ;
        RECT  11.4475 9.835 11.5175 9.975 ;
        RECT  11.8 11.57 11.87 11.705 ;
        RECT  11.8 11.0 11.87 11.135 ;
        RECT  11.095 11.0 11.165 11.135 ;
        RECT  11.515 11.205 11.585 11.34 ;
        RECT  11.8 13.4975 11.87 13.6325 ;
        RECT  11.515 10.795 11.585 10.93 ;
        RECT  11.375 10.795 11.445 10.93 ;
        RECT  11.8 11.205 11.87 11.34 ;
        RECT  11.095 11.205 11.165 11.34 ;
        RECT  11.235 10.23 11.37 10.3 ;
        RECT  11.375 13.175 11.445 13.31 ;
        RECT  11.545 11.57 11.615 11.705 ;
        RECT  11.235 12.485 11.305 12.62 ;
        RECT  11.375 11.205 11.445 11.34 ;
        RECT  11.095 11.57 11.165 11.705 ;
        RECT  11.545 12.085 11.615 12.22 ;
        RECT  11.28 13.7075 11.35 13.8425 ;
        RECT  11.095 13.4975 11.165 13.6325 ;
        RECT  11.28 13.71 11.35 14.01 ;
        RECT  11.28 13.945 11.35 14.01 ;
        RECT  11.6175 13.95 11.6825 14.01 ;
        RECT  11.45 9.84 11.515 9.9025 ;
        RECT  11.8 9.835 11.87 14.01 ;
        RECT  11.095 9.835 11.165 14.01 ;
        RECT  11.615 11.57 11.685 14.01 ;
        RECT  11.325 9.9675 11.5175 10.0375 ;
        RECT  11.515 10.93 11.585 11.205 ;
        RECT  11.235 10.3 11.305 12.62 ;
        RECT  11.375 10.93 11.445 11.205 ;
        RECT  11.375 11.205 11.445 13.3025 ;
        RECT  12.0425 9.9675 12.1775 10.0375 ;
        RECT  12.1525 9.835 12.2225 9.975 ;
        RECT  12.505 11.57 12.575 11.705 ;
        RECT  12.505 11.0 12.575 11.135 ;
        RECT  11.8 11.0 11.87 11.135 ;
        RECT  12.22 11.205 12.29 11.34 ;
        RECT  12.505 13.4975 12.575 13.6325 ;
        RECT  12.22 10.795 12.29 10.93 ;
        RECT  12.08 10.795 12.15 10.93 ;
        RECT  12.505 11.205 12.575 11.34 ;
        RECT  11.8 11.205 11.87 11.34 ;
        RECT  11.94 10.23 12.075 10.3 ;
        RECT  12.08 13.175 12.15 13.31 ;
        RECT  12.25 11.57 12.32 11.705 ;
        RECT  11.94 12.485 12.01 12.62 ;
        RECT  12.08 11.205 12.15 11.34 ;
        RECT  11.8 11.57 11.87 11.705 ;
        RECT  12.25 12.085 12.32 12.22 ;
        RECT  11.985 13.7075 12.055 13.8425 ;
        RECT  11.8 13.4975 11.87 13.6325 ;
        RECT  11.985 13.71 12.055 14.01 ;
        RECT  11.985 13.945 12.055 14.01 ;
        RECT  12.3225 13.95 12.3875 14.01 ;
        RECT  12.155 9.84 12.22 9.9025 ;
        RECT  12.505 9.835 12.575 14.01 ;
        RECT  11.8 9.835 11.87 14.01 ;
        RECT  12.32 11.57 12.39 14.01 ;
        RECT  12.03 9.9675 12.2225 10.0375 ;
        RECT  12.22 10.93 12.29 11.205 ;
        RECT  11.94 10.3 12.01 12.62 ;
        RECT  12.08 10.93 12.15 11.205 ;
        RECT  12.08 11.205 12.15 13.3025 ;
        RECT  11.2925 9.0975 11.3625 9.2325 ;
        RECT  11.8 3.92 11.87 4.055 ;
        RECT  11.6575 8.0025 11.7275 8.1375 ;
        RECT  11.66 6.395 11.73 6.53 ;
        RECT  11.66 4.9975 11.73 5.1325 ;
        RECT  11.095 3.78 11.165 3.915 ;
        RECT  11.4475 3.395 11.5175 3.535 ;
        RECT  11.8 6.8575 11.87 6.9925 ;
        RECT  11.295 5.6625 11.365 5.7975 ;
        RECT  11.66 9.355 11.73 9.49 ;
        RECT  11.4825 8.845 11.5525 8.98 ;
        RECT  11.8 8.4325 11.87 8.5675 ;
        RECT  11.8 3.73 11.87 3.865 ;
        RECT  11.8 5.4725 11.87 5.6075 ;
        RECT  11.295 5.2725 11.365 5.4075 ;
        RECT  11.4825 5.2725 11.5525 5.4075 ;
        RECT  11.4825 5.885 11.5525 6.02 ;
        RECT  11.2925 8.2325 11.3625 8.3675 ;
        RECT  11.4825 8.2325 11.5525 8.3675 ;
        RECT  11.5175 9.565 11.66 9.635 ;
        RECT  11.4475 3.395 11.5175 3.54 ;
        RECT  11.5125 3.47 11.66 3.54 ;
        RECT  11.4475 9.565 11.5175 9.835 ;
        RECT  11.0975 9.3575 11.16 9.4175 ;
        RECT  11.095 3.395 11.165 9.835 ;
        RECT  11.45 9.77 11.515 9.83 ;
        RECT  11.66 9.355 11.73 9.635 ;
        RECT  11.66 3.47 11.73 5.1325 ;
        RECT  11.2925 9.1475 11.3625 9.835 ;
        RECT  11.66 6.53 11.73 8.1375 ;
        RECT  11.4825 8.2325 11.5525 8.95 ;
        RECT  11.295 5.2725 11.365 5.7975 ;
        RECT  11.2975 9.6975 11.36 9.7575 ;
        RECT  11.2925 8.2325 11.3625 9.1725 ;
        RECT  11.4475 3.4 11.515 3.465 ;
        RECT  11.8 3.395 11.87 9.835 ;
        RECT  11.4825 5.2725 11.5525 5.99 ;
        RECT  12.3075 9.0975 12.3775 9.2325 ;
        RECT  11.8 3.92 11.87 4.055 ;
        RECT  11.9425 8.0025 12.0125 8.1375 ;
        RECT  11.94 6.395 12.01 6.53 ;
        RECT  11.94 4.9975 12.01 5.1325 ;
        RECT  12.505 3.78 12.575 3.915 ;
        RECT  12.1525 3.395 12.2225 3.535 ;
        RECT  11.8 6.8575 11.87 6.9925 ;
        RECT  12.305 5.6625 12.375 5.7975 ;
        RECT  11.94 9.355 12.01 9.49 ;
        RECT  12.1175 8.845 12.1875 8.98 ;
        RECT  11.8 8.4325 11.87 8.5675 ;
        RECT  11.8 3.73 11.87 3.865 ;
        RECT  11.8 5.4725 11.87 5.6075 ;
        RECT  12.305 5.2725 12.375 5.4075 ;
        RECT  12.1175 5.2725 12.1875 5.4075 ;
        RECT  12.1175 5.885 12.1875 6.02 ;
        RECT  12.3075 8.2325 12.3775 8.3675 ;
        RECT  12.1175 8.2325 12.1875 8.3675 ;
        RECT  12.01 9.565 12.1525 9.635 ;
        RECT  12.1525 3.395 12.2225 3.54 ;
        RECT  12.01 3.47 12.1575 3.54 ;
        RECT  12.1525 9.565 12.2225 9.835 ;
        RECT  12.51 9.3575 12.5725 9.4175 ;
        RECT  12.505 3.395 12.575 9.835 ;
        RECT  12.155 9.77 12.22 9.83 ;
        RECT  11.94 9.355 12.01 9.635 ;
        RECT  11.94 3.47 12.01 5.1325 ;
        RECT  12.3075 9.1475 12.3775 9.835 ;
        RECT  11.94 6.53 12.01 8.1375 ;
        RECT  12.1175 8.2325 12.1875 8.95 ;
        RECT  12.305 5.2725 12.375 5.7975 ;
        RECT  12.31 9.6975 12.3725 9.7575 ;
        RECT  12.3075 8.2325 12.3775 9.1725 ;
        RECT  12.155 3.4 12.2225 3.465 ;
        RECT  11.8 3.395 11.87 9.835 ;
        RECT  12.1175 5.2725 12.1875 5.99 ;
        RECT  11.415 5.1775 11.55 5.2475 ;
        RECT  11.8 3.8925 11.87 4.0275 ;
        RECT  11.4475 3.5475 11.5175 3.6875 ;
        RECT  11.5475 5.8175 11.6825 5.8875 ;
        RECT  11.8 5.9525 11.87 6.0875 ;
        RECT  11.2725 5.7625 11.3425 5.8975 ;
        RECT  11.48 5.485 11.55 5.62 ;
        RECT  11.235 3.675 11.4475 3.745 ;
        RECT  11.4475 3.395 11.5175 3.745 ;
        RECT  11.5175 6.13 11.62 6.2 ;
        RECT  11.4475 6.13 11.5175 6.37 ;
        RECT  11.4475 6.3125 11.5175 6.365 ;
        RECT  11.4475 3.55 11.5175 3.6125 ;
        RECT  11.2375 4.31 11.3075 5.8975 ;
        RECT  11.62 5.8175 11.69 6.2 ;
        RECT  11.48 5.2475 11.55 5.485 ;
        RECT  11.8 3.395 11.87 6.37 ;
        RECT  11.8 3.9675 11.87 4.025 ;
        RECT  11.5475 4.31 11.6825 4.38 ;
        RECT  11.3075 4.31 11.5475 4.38 ;
        RECT  11.235 3.675 11.305 4.045 ;
        RECT  11.235 4.045 11.305 4.18 ;
        RECT  12.12 5.1775 12.255 5.2475 ;
        RECT  11.8 3.8925 11.87 4.0275 ;
        RECT  12.1525 3.5475 12.2225 3.6875 ;
        RECT  11.9875 5.8175 12.1225 5.8875 ;
        RECT  11.8 5.9525 11.87 6.0875 ;
        RECT  12.3275 5.7625 12.3975 5.8975 ;
        RECT  12.12 5.485 12.19 5.62 ;
        RECT  12.2225 3.675 12.435 3.745 ;
        RECT  12.1525 3.395 12.2225 3.745 ;
        RECT  12.05 6.13 12.1525 6.2 ;
        RECT  12.1525 6.13 12.2225 6.37 ;
        RECT  12.1525 6.3125 12.2225 6.365 ;
        RECT  12.1525 3.55 12.2225 3.6125 ;
        RECT  12.3625 4.31 12.4325 5.8975 ;
        RECT  11.98 5.8175 12.05 6.2 ;
        RECT  12.12 5.2475 12.19 5.485 ;
        RECT  11.8 3.395 11.87 6.37 ;
        RECT  11.8 3.9675 11.87 4.025 ;
        RECT  11.9875 4.31 12.1225 4.38 ;
        RECT  12.1225 4.31 12.3625 4.38 ;
        RECT  12.365 3.675 12.435 4.045 ;
        RECT  12.365 4.045 12.435 4.18 ;
        RECT  4.045 8.135 4.115 40.415 ;
        RECT  3.87 8.135 3.94 40.415 ;
        RECT  3.695 8.135 3.765 40.415 ;
        RECT  3.52 8.135 3.59 40.415 ;
        RECT  3.345 8.135 3.415 40.415 ;
        RECT  3.17 8.135 3.24 40.415 ;
        RECT  2.995 8.135 3.065 40.415 ;
        RECT  2.82 8.135 2.89 40.415 ;
        RECT  7.525 8.135 7.595 13.305 ;
        RECT  7.35 8.135 7.42 13.305 ;
        RECT  6.51 8.135 6.58 13.305 ;
        RECT  6.335 8.135 6.405 13.305 ;
        RECT  6.16 8.135 6.23 13.305 ;
        RECT  5.985 8.135 6.055 13.305 ;
        RECT  5.81 8.135 5.88 13.305 ;
        RECT  5.635 8.135 5.705 13.305 ;
        RECT  6.125 9.18 6.26 9.25 ;
        RECT  7.49 8.6575 7.625 8.7275 ;
        RECT  5.95 9.57 6.085 9.64 ;
        RECT  7.315 10.0925 7.45 10.1625 ;
        RECT  6.125 8.9725 6.26 9.0425 ;
        RECT  5.95 8.4425 6.085 8.5125 ;
        RECT  5.775 9.7775 5.91 9.8475 ;
        RECT  5.95 10.3075 6.085 10.3775 ;
        RECT  6.125 11.6625 6.26 11.7325 ;
        RECT  5.6 11.1325 5.735 11.2025 ;
        RECT  5.775 12.4675 5.91 12.5375 ;
        RECT  7.49 12.4675 7.625 12.5375 ;
        RECT  5.6 12.9975 5.735 13.0675 ;
        RECT  7.315 12.9975 7.45 13.0675 ;
        RECT  6.3 8.03 6.435 8.1 ;
        RECT  6.475 9.375 6.61 9.445 ;
        RECT  6.3 10.72 6.435 10.79 ;
        RECT  6.475 12.065 6.61 12.135 ;
        RECT  6.3 13.2325 6.435 13.3025 ;
        RECT  7.525 13.515 7.595 18.685 ;
        RECT  7.35 13.515 7.42 18.685 ;
        RECT  6.51 13.515 6.58 18.685 ;
        RECT  6.335 13.515 6.405 18.685 ;
        RECT  6.16 13.515 6.23 18.685 ;
        RECT  5.985 13.515 6.055 18.685 ;
        RECT  5.81 13.515 5.88 18.685 ;
        RECT  5.635 13.515 5.705 18.685 ;
        RECT  6.125 14.56 6.26 14.63 ;
        RECT  7.49 14.0375 7.625 14.1075 ;
        RECT  5.95 14.95 6.085 15.02 ;
        RECT  7.315 15.4725 7.45 15.5425 ;
        RECT  6.125 14.3525 6.26 14.4225 ;
        RECT  5.95 13.8225 6.085 13.8925 ;
        RECT  5.775 15.1575 5.91 15.2275 ;
        RECT  5.95 15.6875 6.085 15.7575 ;
        RECT  6.125 17.0425 6.26 17.1125 ;
        RECT  5.6 16.5125 5.735 16.5825 ;
        RECT  5.775 17.8475 5.91 17.9175 ;
        RECT  7.49 17.8475 7.625 17.9175 ;
        RECT  5.6 18.3775 5.735 18.4475 ;
        RECT  7.315 18.3775 7.45 18.4475 ;
        RECT  6.3 13.41 6.435 13.48 ;
        RECT  6.475 14.755 6.61 14.825 ;
        RECT  6.3 16.1 6.435 16.17 ;
        RECT  6.475 17.445 6.61 17.515 ;
        RECT  6.3 18.6125 6.435 18.6825 ;
        RECT  2.79 8.7275 2.925 8.7975 ;
        RECT  2.965 10.1625 3.1 10.2325 ;
        RECT  3.14 11.4175 3.275 11.4875 ;
        RECT  3.315 12.8525 3.45 12.9225 ;
        RECT  3.49 14.1075 3.625 14.1775 ;
        RECT  3.665 15.5425 3.8 15.6125 ;
        RECT  3.84 16.7975 3.975 16.8675 ;
        RECT  4.015 18.2325 4.15 18.3025 ;
        RECT  2.79 19.8025 2.925 19.8725 ;
        RECT  3.49 19.2725 3.625 19.3425 ;
        RECT  2.79 20.6075 2.925 20.6775 ;
        RECT  3.665 21.1375 3.8 21.2075 ;
        RECT  2.79 22.4925 2.925 22.5625 ;
        RECT  3.84 21.9625 3.975 22.0325 ;
        RECT  2.79 23.2975 2.925 23.3675 ;
        RECT  4.015 23.8275 4.15 23.8975 ;
        RECT  2.965 25.1825 3.1 25.2525 ;
        RECT  3.49 24.6525 3.625 24.7225 ;
        RECT  2.965 25.9875 3.1 26.0575 ;
        RECT  3.665 26.5175 3.8 26.5875 ;
        RECT  2.965 27.8725 3.1 27.9425 ;
        RECT  3.84 27.3425 3.975 27.4125 ;
        RECT  2.965 28.6775 3.1 28.7475 ;
        RECT  4.015 29.2075 4.15 29.2775 ;
        RECT  3.14 30.5625 3.275 30.6325 ;
        RECT  3.49 30.0325 3.625 30.1025 ;
        RECT  3.14 31.3675 3.275 31.4375 ;
        RECT  3.665 31.8975 3.8 31.9675 ;
        RECT  3.14 33.2525 3.275 33.3225 ;
        RECT  3.84 32.7225 3.975 32.7925 ;
        RECT  3.14 34.0575 3.275 34.1275 ;
        RECT  4.015 34.5875 4.15 34.6575 ;
        RECT  3.315 35.9425 3.45 36.0125 ;
        RECT  3.49 35.4125 3.625 35.4825 ;
        RECT  3.315 36.7475 3.45 36.8175 ;
        RECT  3.665 37.2775 3.8 37.3475 ;
        RECT  3.315 38.6325 3.45 38.7025 ;
        RECT  3.84 38.1025 3.975 38.1725 ;
        RECT  3.315 39.4375 3.45 39.5075 ;
        RECT  4.015 39.9675 4.15 40.0375 ;
        RECT  5.53 20.205 5.985 20.275 ;
        RECT  5.53 19.805 6.545 19.875 ;
        RECT  5.53 21.55 5.985 21.62 ;
        RECT  5.53 20.605 6.545 20.675 ;
        RECT  5.53 22.895 5.985 22.965 ;
        RECT  5.53 22.495 6.545 22.565 ;
        RECT  5.53 24.24 5.985 24.31 ;
        RECT  5.53 23.295 6.545 23.365 ;
        RECT  5.53 25.585 5.985 25.655 ;
        RECT  5.53 25.185 6.545 25.255 ;
        RECT  5.53 26.93 5.985 27.0 ;
        RECT  5.53 25.985 6.545 26.055 ;
        RECT  5.53 28.275 5.985 28.345 ;
        RECT  5.53 27.875 6.545 27.945 ;
        RECT  5.53 29.62 5.985 29.69 ;
        RECT  5.53 28.675 6.545 28.745 ;
        RECT  5.53 30.965 5.985 31.035 ;
        RECT  5.53 30.565 6.545 30.635 ;
        RECT  5.53 32.31 5.985 32.38 ;
        RECT  5.53 31.365 6.545 31.435 ;
        RECT  5.53 33.655 5.985 33.725 ;
        RECT  5.53 33.255 6.545 33.325 ;
        RECT  5.53 35.0 5.985 35.07 ;
        RECT  5.53 34.055 6.545 34.125 ;
        RECT  5.53 36.345 5.985 36.415 ;
        RECT  5.53 35.945 6.545 36.015 ;
        RECT  5.53 37.69 5.985 37.76 ;
        RECT  5.53 36.745 6.545 36.815 ;
        RECT  5.53 39.035 5.985 39.105 ;
        RECT  5.53 38.635 6.545 38.705 ;
        RECT  5.53 40.38 5.985 40.45 ;
        RECT  5.53 39.435 6.545 39.505 ;
        RECT  5.46 20.205 5.595 20.275 ;
        RECT  5.915 20.205 6.05 20.275 ;
        RECT  6.545 19.805 6.68 19.875 ;
        RECT  5.53 19.805 5.6 19.94 ;
        RECT  5.46 21.55 5.595 21.62 ;
        RECT  5.915 21.55 6.05 21.62 ;
        RECT  6.545 20.605 6.68 20.675 ;
        RECT  5.53 20.54 5.6 20.675 ;
        RECT  5.46 22.895 5.595 22.965 ;
        RECT  5.915 22.895 6.05 22.965 ;
        RECT  6.545 22.495 6.68 22.565 ;
        RECT  5.53 22.495 5.6 22.63 ;
        RECT  5.46 24.24 5.595 24.31 ;
        RECT  5.915 24.24 6.05 24.31 ;
        RECT  6.545 23.295 6.68 23.365 ;
        RECT  5.53 23.23 5.6 23.365 ;
        RECT  5.46 25.585 5.595 25.655 ;
        RECT  5.915 25.585 6.05 25.655 ;
        RECT  6.545 25.185 6.68 25.255 ;
        RECT  5.53 25.185 5.6 25.32 ;
        RECT  5.46 26.93 5.595 27.0 ;
        RECT  5.915 26.93 6.05 27.0 ;
        RECT  6.545 25.985 6.68 26.055 ;
        RECT  5.53 25.92 5.6 26.055 ;
        RECT  5.46 28.275 5.595 28.345 ;
        RECT  5.915 28.275 6.05 28.345 ;
        RECT  6.545 27.875 6.68 27.945 ;
        RECT  5.53 27.875 5.6 28.01 ;
        RECT  5.46 29.62 5.595 29.69 ;
        RECT  5.915 29.62 6.05 29.69 ;
        RECT  6.545 28.675 6.68 28.745 ;
        RECT  5.53 28.61 5.6 28.745 ;
        RECT  5.46 30.965 5.595 31.035 ;
        RECT  5.915 30.965 6.05 31.035 ;
        RECT  6.545 30.565 6.68 30.635 ;
        RECT  5.53 30.565 5.6 30.7 ;
        RECT  5.46 32.31 5.595 32.38 ;
        RECT  5.915 32.31 6.05 32.38 ;
        RECT  6.545 31.365 6.68 31.435 ;
        RECT  5.53 31.3 5.6 31.435 ;
        RECT  5.46 33.655 5.595 33.725 ;
        RECT  5.915 33.655 6.05 33.725 ;
        RECT  6.545 33.255 6.68 33.325 ;
        RECT  5.53 33.255 5.6 33.39 ;
        RECT  5.46 35.0 5.595 35.07 ;
        RECT  5.915 35.0 6.05 35.07 ;
        RECT  6.545 34.055 6.68 34.125 ;
        RECT  5.53 33.99 5.6 34.125 ;
        RECT  5.46 36.345 5.595 36.415 ;
        RECT  5.915 36.345 6.05 36.415 ;
        RECT  6.545 35.945 6.68 36.015 ;
        RECT  5.53 35.945 5.6 36.08 ;
        RECT  5.46 37.69 5.595 37.76 ;
        RECT  5.915 37.69 6.05 37.76 ;
        RECT  6.545 36.745 6.68 36.815 ;
        RECT  5.53 36.68 5.6 36.815 ;
        RECT  5.46 39.035 5.595 39.105 ;
        RECT  5.915 39.035 6.05 39.105 ;
        RECT  6.545 38.635 6.68 38.705 ;
        RECT  5.53 38.635 5.6 38.77 ;
        RECT  5.46 40.38 5.595 40.45 ;
        RECT  5.915 40.38 6.05 40.45 ;
        RECT  6.545 39.435 6.68 39.505 ;
        RECT  5.53 39.37 5.6 39.505 ;
        RECT  6.6125 7.6075 6.7475 7.6775 ;
        RECT  1.435 7.1 1.57 7.17 ;
        RECT  5.5175 7.2425 5.6525 7.3125 ;
        RECT  3.91 7.24 4.045 7.31 ;
        RECT  2.5125 7.24 2.6475 7.31 ;
        RECT  1.295 7.805 1.43 7.875 ;
        RECT  0.91 7.4525 1.05 7.5225 ;
        RECT  4.3725 7.1 4.5075 7.17 ;
        RECT  3.1775 7.605 3.3125 7.675 ;
        RECT  6.87 7.24 7.005 7.31 ;
        RECT  6.36 7.4175 6.495 7.4875 ;
        RECT  5.9475 7.1 6.0825 7.17 ;
        RECT  1.245 7.1 1.38 7.17 ;
        RECT  2.9875 7.1 3.1225 7.17 ;
        RECT  2.7875 7.605 2.9225 7.675 ;
        RECT  2.7875 7.4175 2.9225 7.4875 ;
        RECT  3.4 7.4175 3.535 7.4875 ;
        RECT  5.7475 7.6075 5.8825 7.6775 ;
        RECT  5.7475 7.4175 5.8825 7.4875 ;
        RECT  7.08 7.31 7.15 7.4525 ;
        RECT  0.91 7.4525 1.055 7.5225 ;
        RECT  0.985 7.31 1.055 7.4575 ;
        RECT  7.08 7.4525 7.35 7.5225 ;
        RECT  6.8725 7.81 6.9325 7.8725 ;
        RECT  0.91 7.805 7.35 7.875 ;
        RECT  7.285 7.455 7.345 7.52 ;
        RECT  6.87 7.24 7.15 7.31 ;
        RECT  0.985 7.24 2.6475 7.31 ;
        RECT  6.6625 7.6075 7.35 7.6775 ;
        RECT  4.045 7.24 5.6525 7.31 ;
        RECT  5.7475 7.4175 6.465 7.4875 ;
        RECT  2.7875 7.605 3.3125 7.675 ;
        RECT  7.2125 7.61 7.2725 7.6725 ;
        RECT  5.7475 7.6075 6.6875 7.6775 ;
        RECT  0.915 7.455 0.98 7.5225 ;
        RECT  0.91 7.1 7.35 7.17 ;
        RECT  2.7875 7.4175 3.505 7.4875 ;
        RECT  6.6125 6.5925 6.7475 6.6625 ;
        RECT  1.435 7.1 1.57 7.17 ;
        RECT  5.5175 6.9575 5.6525 7.0275 ;
        RECT  3.91 6.96 4.045 7.03 ;
        RECT  2.5125 6.96 2.6475 7.03 ;
        RECT  1.295 6.395 1.43 6.465 ;
        RECT  0.91 6.7475 1.05 6.8175 ;
        RECT  4.3725 7.1 4.5075 7.17 ;
        RECT  3.1775 6.595 3.3125 6.665 ;
        RECT  6.87 6.96 7.005 7.03 ;
        RECT  6.36 6.7825 6.495 6.8525 ;
        RECT  5.9475 7.1 6.0825 7.17 ;
        RECT  1.245 7.1 1.38 7.17 ;
        RECT  2.9875 7.1 3.1225 7.17 ;
        RECT  2.7875 6.595 2.9225 6.665 ;
        RECT  2.7875 6.7825 2.9225 6.8525 ;
        RECT  3.4 6.7825 3.535 6.8525 ;
        RECT  5.7475 6.5925 5.8825 6.6625 ;
        RECT  5.7475 6.7825 5.8825 6.8525 ;
        RECT  7.08 6.8175 7.15 6.96 ;
        RECT  0.91 6.7475 1.055 6.8175 ;
        RECT  0.985 6.8125 1.055 6.96 ;
        RECT  7.08 6.7475 7.35 6.8175 ;
        RECT  6.8725 6.3975 6.9325 6.46 ;
        RECT  0.91 6.395 7.35 6.465 ;
        RECT  7.285 6.75 7.345 6.815 ;
        RECT  6.87 6.96 7.15 7.03 ;
        RECT  0.985 6.96 2.6475 7.03 ;
        RECT  6.6625 6.5925 7.35 6.6625 ;
        RECT  4.045 6.96 5.6525 7.03 ;
        RECT  5.7475 6.7825 6.465 6.8525 ;
        RECT  2.7875 6.595 3.3125 6.665 ;
        RECT  7.2125 6.5975 7.2725 6.66 ;
        RECT  5.7475 6.5925 6.6875 6.6625 ;
        RECT  0.915 6.7475 0.98 6.815 ;
        RECT  0.91 7.1 7.35 7.17 ;
        RECT  2.7875 6.7825 3.505 6.8525 ;
        RECT  6.6125 6.1975 6.7475 6.2675 ;
        RECT  1.435 5.69 1.57 5.76 ;
        RECT  5.5175 5.8325 5.6525 5.9025 ;
        RECT  3.91 5.83 4.045 5.9 ;
        RECT  2.5125 5.83 2.6475 5.9 ;
        RECT  1.295 6.395 1.43 6.465 ;
        RECT  0.91 6.0425 1.05 6.1125 ;
        RECT  4.3725 5.69 4.5075 5.76 ;
        RECT  3.1775 6.195 3.3125 6.265 ;
        RECT  6.87 5.83 7.005 5.9 ;
        RECT  6.36 6.0075 6.495 6.0775 ;
        RECT  5.9475 5.69 6.0825 5.76 ;
        RECT  1.245 5.69 1.38 5.76 ;
        RECT  2.9875 5.69 3.1225 5.76 ;
        RECT  2.7875 6.195 2.9225 6.265 ;
        RECT  2.7875 6.0075 2.9225 6.0775 ;
        RECT  3.4 6.0075 3.535 6.0775 ;
        RECT  5.7475 6.1975 5.8825 6.2675 ;
        RECT  5.7475 6.0075 5.8825 6.0775 ;
        RECT  7.08 5.9 7.15 6.0425 ;
        RECT  0.91 6.0425 1.055 6.1125 ;
        RECT  0.985 5.9 1.055 6.0475 ;
        RECT  7.08 6.0425 7.35 6.1125 ;
        RECT  6.8725 6.4 6.9325 6.4625 ;
        RECT  0.91 6.395 7.35 6.465 ;
        RECT  7.285 6.045 7.345 6.11 ;
        RECT  6.87 5.83 7.15 5.9 ;
        RECT  0.985 5.83 2.6475 5.9 ;
        RECT  6.6625 6.1975 7.35 6.2675 ;
        RECT  4.045 5.83 5.6525 5.9 ;
        RECT  5.7475 6.0075 6.465 6.0775 ;
        RECT  2.7875 6.195 3.3125 6.265 ;
        RECT  7.2125 6.2 7.2725 6.2625 ;
        RECT  5.7475 6.1975 6.6875 6.2675 ;
        RECT  0.915 6.045 0.98 6.1125 ;
        RECT  0.91 5.69 7.35 5.76 ;
        RECT  2.7875 6.0075 3.505 6.0775 ;
        RECT  6.6125 5.1825 6.7475 5.2525 ;
        RECT  1.435 5.69 1.57 5.76 ;
        RECT  5.5175 5.5475 5.6525 5.6175 ;
        RECT  3.91 5.55 4.045 5.62 ;
        RECT  2.5125 5.55 2.6475 5.62 ;
        RECT  1.295 4.985 1.43 5.055 ;
        RECT  0.91 5.3375 1.05 5.4075 ;
        RECT  4.3725 5.69 4.5075 5.76 ;
        RECT  3.1775 5.185 3.3125 5.255 ;
        RECT  6.87 5.55 7.005 5.62 ;
        RECT  6.36 5.3725 6.495 5.4425 ;
        RECT  5.9475 5.69 6.0825 5.76 ;
        RECT  1.245 5.69 1.38 5.76 ;
        RECT  2.9875 5.69 3.1225 5.76 ;
        RECT  2.7875 5.185 2.9225 5.255 ;
        RECT  2.7875 5.3725 2.9225 5.4425 ;
        RECT  3.4 5.3725 3.535 5.4425 ;
        RECT  5.7475 5.1825 5.8825 5.2525 ;
        RECT  5.7475 5.3725 5.8825 5.4425 ;
        RECT  7.08 5.4075 7.15 5.55 ;
        RECT  0.91 5.3375 1.055 5.4075 ;
        RECT  0.985 5.4025 1.055 5.55 ;
        RECT  7.08 5.3375 7.35 5.4075 ;
        RECT  6.8725 4.9875 6.9325 5.05 ;
        RECT  0.91 4.985 7.35 5.055 ;
        RECT  7.285 5.34 7.345 5.405 ;
        RECT  6.87 5.55 7.15 5.62 ;
        RECT  0.985 5.55 2.6475 5.62 ;
        RECT  6.6625 5.1825 7.35 5.2525 ;
        RECT  4.045 5.55 5.6525 5.62 ;
        RECT  5.7475 5.3725 6.465 5.4425 ;
        RECT  2.7875 5.185 3.3125 5.255 ;
        RECT  7.2125 5.1875 7.2725 5.25 ;
        RECT  5.7475 5.1825 6.6875 5.2525 ;
        RECT  0.915 5.3375 0.98 5.405 ;
        RECT  0.91 5.69 7.35 5.76 ;
        RECT  2.7875 5.3725 3.505 5.4425 ;
        RECT  11.4475 0.2775 11.5175 0.3475 ;
        RECT  11.2725 0.2775 11.4825 0.3475 ;
        RECT  11.4475 0.3125 11.5175 0.54 ;
        RECT  11.2375 0.2775 11.3075 0.4125 ;
        RECT  12.1525 0.2775 12.2225 0.3475 ;
        RECT  11.9775 0.2775 12.1875 0.3475 ;
        RECT  12.1525 0.3125 12.2225 0.54 ;
        RECT  11.9425 0.2775 12.0125 0.4125 ;
        RECT  11.4475 0.0 11.5175 0.135 ;
        RECT  12.1525 0.0 12.2225 0.135 ;
        RECT  8.54 8.73 8.61 8.865 ;
        RECT  8.54 7.4525 8.61 7.5875 ;
        RECT  7.08 7.4525 7.215 7.5225 ;
        RECT  8.33 10.165 8.4 10.3 ;
        RECT  8.33 6.7475 8.4 6.8825 ;
        RECT  7.08 6.7475 7.215 6.8175 ;
        RECT  8.12 14.11 8.19 14.245 ;
        RECT  8.12 6.0425 8.19 6.1775 ;
        RECT  7.08 6.0425 7.215 6.1125 ;
        RECT  7.91 15.545 7.98 15.68 ;
        RECT  7.91 5.3375 7.98 5.4725 ;
        RECT  7.08 5.3375 7.215 5.4075 ;
        RECT  10.36 3.6 10.43 3.735 ;
        RECT  9.94 1.415 10.01 1.55 ;
        RECT  10.15 2.9625 10.22 3.0975 ;
        RECT  10.36 41.1 10.43 41.235 ;
        RECT  10.57 10.1025 10.64 10.2375 ;
        RECT  10.78 14.1275 10.85 14.2625 ;
        RECT  0.98 7.6275 1.115 7.6975 ;
        RECT  0.98 7.6275 1.115 7.6975 ;
        RECT  9.73 7.98 9.8 8.115 ;
        RECT  9.73 41.53 9.8 41.665 ;
        RECT  8.89 40.545 9.095 40.68 ;
        RECT  11.77 40.545 11.905 40.615 ;
        RECT  12.475 40.545 12.61 40.615 ;
        RECT  10.995 40.545 11.13 40.615 ;
        RECT  9.385 0.355 9.59 0.49 ;
        RECT  11.8 0.355 11.87 0.49 ;
        RECT  11.8 0.355 11.87 0.49 ;
        RECT  7.755 21.5525 7.89 21.6225 ;
        RECT  7.755 24.2425 7.89 24.3125 ;
        RECT  7.755 26.9325 7.89 27.0025 ;
        RECT  7.755 29.6225 7.89 29.6925 ;
        RECT  7.755 32.3125 7.89 32.3825 ;
        RECT  7.755 35.0025 7.89 35.0725 ;
        RECT  7.755 37.6925 7.89 37.7625 ;
        RECT  7.755 40.3825 7.89 40.4525 ;
        RECT  8.89 13.4125 9.095 13.5475 ;
        RECT  8.89 18.7925 9.095 18.9275 ;
        RECT  7.28 7.8075 7.415 7.8775 ;
        RECT  8.89 7.8075 9.095 7.9425 ;
        RECT  7.28 6.3975 7.415 6.4675 ;
        RECT  8.89 6.3975 9.095 6.5325 ;
        RECT  7.28 6.3975 7.415 6.4675 ;
        RECT  8.89 6.3975 9.095 6.5325 ;
        RECT  7.28 4.9875 7.415 5.0575 ;
        RECT  8.89 4.9875 9.095 5.1225 ;
        RECT  -5.73 14.925 -0.35 14.995 ;
        RECT  -5.73 15.135 -0.35 15.205 ;
        RECT  -5.73 15.345 -0.35 15.415 ;
        RECT  -5.73 15.555 -0.35 15.625 ;
        RECT  -5.73 15.765 -0.35 15.835 ;
        RECT  -5.73 15.975 -0.35 16.045 ;
        RECT  -5.73 19.225 -0.35 19.295 ;
        RECT  -5.73 19.435 -0.35 19.505 ;
        RECT  -5.73 19.645 -0.35 19.715 ;
        RECT  -5.73 19.855 -0.35 19.925 ;
        RECT  -5.765 14.715 -5.695 14.995 ;
        RECT  -4.355 14.715 -4.285 14.995 ;
        RECT  -4.355 14.715 -4.285 14.995 ;
        RECT  -0.35 15.975 -0.14 16.045 ;
        RECT  -0.8675 8.415 -0.14 8.485 ;
        RECT  -1.0125 16.865 -0.14 16.935 ;
        RECT  -0.35 19.225 -0.14 19.295 ;
        RECT  -0.965 17.335 -0.14 17.405 ;
        RECT  -5.5675 13.9775 -5.4975 14.1125 ;
        RECT  -5.06 8.8 -4.99 8.935 ;
        RECT  -5.2025 12.8825 -5.1325 13.0175 ;
        RECT  -5.2 11.275 -5.13 11.41 ;
        RECT  -5.2 9.8775 -5.13 10.0125 ;
        RECT  -5.765 8.66 -5.695 8.795 ;
        RECT  -5.4125 8.275 -5.3425 8.415 ;
        RECT  -5.06 11.7375 -4.99 11.8725 ;
        RECT  -5.565 10.5425 -5.495 10.6775 ;
        RECT  -5.2 14.235 -5.13 14.37 ;
        RECT  -5.3775 13.725 -5.3075 13.86 ;
        RECT  -5.06 13.3125 -4.99 13.4475 ;
        RECT  -5.06 8.61 -4.99 8.745 ;
        RECT  -5.06 10.3525 -4.99 10.4875 ;
        RECT  -5.565 10.1525 -5.495 10.2875 ;
        RECT  -5.3775 10.1525 -5.3075 10.2875 ;
        RECT  -5.3775 10.765 -5.3075 10.9 ;
        RECT  -5.5675 13.1125 -5.4975 13.2475 ;
        RECT  -5.3775 13.1125 -5.3075 13.2475 ;
        RECT  -5.3425 14.445 -5.2 14.515 ;
        RECT  -5.4125 8.275 -5.3425 8.42 ;
        RECT  -5.3475 8.35 -5.2 8.42 ;
        RECT  -5.4125 14.445 -5.3425 14.715 ;
        RECT  -5.7625 14.2375 -5.7 14.2975 ;
        RECT  -5.765 8.275 -5.695 14.715 ;
        RECT  -5.41 14.65 -5.345 14.71 ;
        RECT  -5.2 14.235 -5.13 14.515 ;
        RECT  -5.2 8.35 -5.13 10.0125 ;
        RECT  -5.5675 14.0275 -5.4975 14.715 ;
        RECT  -5.2 11.41 -5.13 13.0175 ;
        RECT  -5.3775 13.1125 -5.3075 13.83 ;
        RECT  -5.565 10.1525 -5.495 10.6775 ;
        RECT  -5.5625 14.5775 -5.5 14.6375 ;
        RECT  -5.5675 13.1125 -5.4975 14.0525 ;
        RECT  -5.4125 8.28 -5.345 8.345 ;
        RECT  -5.06 8.275 -4.99 14.715 ;
        RECT  -5.3775 10.1525 -5.3075 10.87 ;
        RECT  -4.5525 13.9775 -4.4825 14.1125 ;
        RECT  -5.06 8.8 -4.99 8.935 ;
        RECT  -4.9175 12.8825 -4.8475 13.0175 ;
        RECT  -4.92 11.275 -4.85 11.41 ;
        RECT  -4.92 9.8775 -4.85 10.0125 ;
        RECT  -4.355 8.66 -4.285 8.795 ;
        RECT  -4.7075 8.275 -4.6375 8.415 ;
        RECT  -5.06 11.7375 -4.99 11.8725 ;
        RECT  -4.555 10.5425 -4.485 10.6775 ;
        RECT  -4.92 14.235 -4.85 14.37 ;
        RECT  -4.7425 13.725 -4.6725 13.86 ;
        RECT  -5.06 13.3125 -4.99 13.4475 ;
        RECT  -5.06 8.61 -4.99 8.745 ;
        RECT  -5.06 10.3525 -4.99 10.4875 ;
        RECT  -4.555 10.1525 -4.485 10.2875 ;
        RECT  -4.7425 10.1525 -4.6725 10.2875 ;
        RECT  -4.7425 10.765 -4.6725 10.9 ;
        RECT  -4.5525 13.1125 -4.4825 13.2475 ;
        RECT  -4.7425 13.1125 -4.6725 13.2475 ;
        RECT  -4.85 14.445 -4.7075 14.515 ;
        RECT  -4.7075 8.275 -4.6375 8.42 ;
        RECT  -4.85 8.35 -4.7025 8.42 ;
        RECT  -4.7075 14.445 -4.6375 14.715 ;
        RECT  -4.35 14.2375 -4.2875 14.2975 ;
        RECT  -4.355 8.275 -4.285 14.715 ;
        RECT  -4.705 14.65 -4.64 14.71 ;
        RECT  -4.92 14.235 -4.85 14.515 ;
        RECT  -4.92 8.35 -4.85 10.0125 ;
        RECT  -4.5525 14.0275 -4.4825 14.715 ;
        RECT  -4.92 11.41 -4.85 13.0175 ;
        RECT  -4.7425 13.1125 -4.6725 13.83 ;
        RECT  -4.555 10.1525 -4.485 10.6775 ;
        RECT  -4.55 14.5775 -4.4875 14.6375 ;
        RECT  -4.5525 13.1125 -4.4825 14.0525 ;
        RECT  -4.705 8.28 -4.6375 8.345 ;
        RECT  -5.06 8.275 -4.99 14.715 ;
        RECT  -4.7425 10.1525 -4.6725 10.87 ;
        RECT  -4.1575 13.9775 -4.0875 14.1125 ;
        RECT  -3.65 8.8 -3.58 8.935 ;
        RECT  -3.7925 12.8825 -3.7225 13.0175 ;
        RECT  -3.79 11.275 -3.72 11.41 ;
        RECT  -3.79 9.8775 -3.72 10.0125 ;
        RECT  -4.355 8.66 -4.285 8.795 ;
        RECT  -4.0025 8.275 -3.9325 8.415 ;
        RECT  -3.65 11.7375 -3.58 11.8725 ;
        RECT  -4.155 10.5425 -4.085 10.6775 ;
        RECT  -3.79 14.235 -3.72 14.37 ;
        RECT  -3.9675 13.725 -3.8975 13.86 ;
        RECT  -3.65 13.3125 -3.58 13.4475 ;
        RECT  -3.65 8.61 -3.58 8.745 ;
        RECT  -3.65 10.3525 -3.58 10.4875 ;
        RECT  -4.155 10.1525 -4.085 10.2875 ;
        RECT  -3.9675 10.1525 -3.8975 10.2875 ;
        RECT  -3.9675 10.765 -3.8975 10.9 ;
        RECT  -4.1575 13.1125 -4.0875 13.2475 ;
        RECT  -3.9675 13.1125 -3.8975 13.2475 ;
        RECT  -3.9325 14.445 -3.79 14.515 ;
        RECT  -4.0025 8.275 -3.9325 8.42 ;
        RECT  -3.9375 8.35 -3.79 8.42 ;
        RECT  -4.0025 14.445 -3.9325 14.715 ;
        RECT  -4.3525 14.2375 -4.29 14.2975 ;
        RECT  -4.355 8.275 -4.285 14.715 ;
        RECT  -4.0 14.65 -3.935 14.71 ;
        RECT  -3.79 14.235 -3.72 14.515 ;
        RECT  -3.79 8.35 -3.72 10.0125 ;
        RECT  -4.1575 14.0275 -4.0875 14.715 ;
        RECT  -3.79 11.41 -3.72 13.0175 ;
        RECT  -3.9675 13.1125 -3.8975 13.83 ;
        RECT  -4.155 10.1525 -4.085 10.6775 ;
        RECT  -4.1525 14.5775 -4.09 14.6375 ;
        RECT  -4.1575 13.1125 -4.0875 14.0525 ;
        RECT  -4.0025 8.28 -3.935 8.345 ;
        RECT  -3.65 8.275 -3.58 14.715 ;
        RECT  -3.9675 10.1525 -3.8975 10.87 ;
        RECT  -1.4125 8.84 -1.2775 8.91 ;
        RECT  -0.8675 8.84 -0.8025 8.91 ;
        RECT  -0.835 8.84 -0.2575 8.91 ;
        RECT  -0.87 8.8075 -0.8 8.9425 ;
        RECT  -1.9775 21.245 -1.9075 21.38 ;
        RECT  -1.0025 23.795 -0.9325 23.93 ;
        RECT  -1.0025 23.235 -0.9325 23.37 ;
        RECT  -2.5225 22.81 -2.4525 22.945 ;
        RECT  -2.5225 23.37 -2.4525 23.505 ;
        RECT  -1.0025 23.4725 -0.9325 23.6075 ;
        RECT  -1.0025 23.37 -0.9325 23.6075 ;
        RECT  -1.0025 22.9125 -0.9325 23.0475 ;
        RECT  -1.0025 22.81 -0.9325 22.88 ;
        RECT  -2.5225 22.81 -2.4525 22.88 ;
        RECT  -1.0025 22.845 -0.9325 23.0475 ;
        RECT  -2.5225 22.81 -2.4525 22.845 ;
        RECT  -1.0025 22.7775 -0.9325 22.9125 ;
        RECT  -2.5225 22.7775 -2.4525 22.9125 ;
        RECT  -2.5225 23.1325 -2.4525 23.2675 ;
        RECT  -2.5225 23.1325 -2.4525 23.37 ;
        RECT  -4.2275 23.0025 -4.1575 23.1375 ;
        RECT  -4.9325 23.4775 -4.8625 23.6125 ;
        RECT  -4.2275 23.4775 -4.1575 23.6125 ;
        RECT  -4.68 22.9975 -4.61 23.1325 ;
        RECT  -4.48 23.0025 -4.41 23.1375 ;
        RECT  -4.965 22.705 -4.83 22.775 ;
        RECT  -4.26 22.705 -4.125 22.775 ;
        RECT  -4.7475 22.7075 -4.6775 22.7725 ;
        RECT  -4.4125 22.7075 -4.3425 22.7725 ;
        RECT  -4.2275 22.705 -4.1575 22.775 ;
        RECT  -4.4125 22.64 -4.3425 24.1975 ;
        RECT  -4.7475 22.64 -4.6775 24.205 ;
        RECT  -4.9325 22.64 -4.8625 24.2075 ;
        RECT  -4.2275 22.64 -4.1575 24.185 ;
        RECT  -4.9325 21.855 -4.8625 21.99 ;
        RECT  -4.9325 21.855 -4.8625 21.99 ;
        RECT  -4.9325 21.855 -4.8625 21.99 ;
        RECT  -4.9325 21.855 -4.8625 21.99 ;
        RECT  -4.9325 21.855 -4.8625 21.99 ;
        RECT  -4.9325 21.855 -4.8625 21.99 ;
        RECT  -4.26 22.705 -4.125 22.775 ;
        RECT  -4.965 22.705 -4.83 22.775 ;
        RECT  -4.9325 21.855 -4.8625 21.99 ;
        RECT  -4.9325 21.855 -4.8625 21.99 ;
        RECT  -4.9325 21.855 -4.8625 21.99 ;
        RECT  -4.9325 21.855 -4.8625 21.99 ;
        RECT  -4.9325 21.855 -4.8625 21.99 ;
        RECT  -4.9325 21.855 -4.8625 21.99 ;
        RECT  -4.9325 21.855 -4.8625 21.99 ;
        RECT  -4.9325 21.855 -4.8625 21.99 ;
        RECT  -4.4825 22.3475 -4.4125 22.4825 ;
        RECT  -4.2275 21.855 -4.1575 21.99 ;
        RECT  -4.2275 21.855 -4.1575 21.99 ;
        RECT  -4.2275 21.855 -4.1575 21.99 ;
        RECT  -4.2275 21.855 -4.1575 21.99 ;
        RECT  -4.2275 21.855 -4.1575 21.99 ;
        RECT  -4.2275 21.855 -4.1575 21.99 ;
        RECT  -4.9325 21.855 -4.8625 21.99 ;
        RECT  -4.9325 21.855 -4.8625 21.99 ;
        RECT  -4.9325 21.855 -4.8625 21.99 ;
        RECT  -4.9325 21.855 -4.8625 21.99 ;
        RECT  -4.6775 22.3475 -4.6075 22.4825 ;
        RECT  -4.965 22.705 -4.83 22.775 ;
        RECT  -4.965 22.705 -4.83 22.775 ;
        RECT  -4.965 22.705 -4.83 22.775 ;
        RECT  -4.9325 21.855 -4.8625 21.99 ;
        RECT  -4.9325 21.855 -4.8625 21.99 ;
        RECT  -4.9325 21.855 -4.8625 21.99 ;
        RECT  -4.9325 21.855 -4.8625 21.99 ;
        RECT  -4.9325 21.855 -4.8625 21.99 ;
        RECT  -4.9325 21.855 -4.8625 21.99 ;
        RECT  -4.26 22.705 -4.125 22.775 ;
        RECT  -4.9325 21.3625 -4.8625 22.7725 ;
        RECT  -4.2225 22.7125 -4.1625 22.77 ;
        RECT  -4.405 22.7125 -4.35 22.765 ;
        RECT  -4.7425 22.7125 -4.685 22.7725 ;
        RECT  -4.9275 22.7075 -4.8675 22.765 ;
        RECT  -4.7475 21.295 -4.6775 22.84 ;
        RECT  -4.4125 21.295 -4.3425 22.84 ;
        RECT  -4.2275 21.295 -4.1575 22.84 ;
        RECT  -4.9325 21.295 -4.8625 22.84 ;
        RECT  -4.9325 20.8 -4.8625 20.935 ;
        RECT  -4.9325 20.8 -4.8625 20.935 ;
        RECT  -4.9325 20.8 -4.8625 20.935 ;
        RECT  -4.9325 20.8 -4.8625 20.935 ;
        RECT  -4.9325 20.8 -4.8625 20.935 ;
        RECT  -4.9325 20.8 -4.8625 20.935 ;
        RECT  -4.26 20.015 -4.125 20.085 ;
        RECT  -4.965 20.015 -4.83 20.085 ;
        RECT  -4.9325 20.8 -4.8625 20.935 ;
        RECT  -4.9325 20.8 -4.8625 20.935 ;
        RECT  -4.9325 20.8 -4.8625 20.935 ;
        RECT  -4.9325 20.8 -4.8625 20.935 ;
        RECT  -4.9325 20.8 -4.8625 20.935 ;
        RECT  -4.9325 20.8 -4.8625 20.935 ;
        RECT  -4.9325 20.8 -4.8625 20.935 ;
        RECT  -4.9325 20.8 -4.8625 20.935 ;
        RECT  -4.4825 20.3075 -4.4125 20.4425 ;
        RECT  -4.2275 20.8 -4.1575 20.935 ;
        RECT  -4.2275 20.8 -4.1575 20.935 ;
        RECT  -4.2275 20.8 -4.1575 20.935 ;
        RECT  -4.2275 20.8 -4.1575 20.935 ;
        RECT  -4.2275 20.8 -4.1575 20.935 ;
        RECT  -4.2275 20.8 -4.1575 20.935 ;
        RECT  -4.9325 20.8 -4.8625 20.935 ;
        RECT  -4.9325 20.8 -4.8625 20.935 ;
        RECT  -4.9325 20.8 -4.8625 20.935 ;
        RECT  -4.9325 20.8 -4.8625 20.935 ;
        RECT  -4.6775 20.3075 -4.6075 20.4425 ;
        RECT  -4.965 20.015 -4.83 20.085 ;
        RECT  -4.965 20.015 -4.83 20.085 ;
        RECT  -4.965 20.015 -4.83 20.085 ;
        RECT  -4.9325 20.8 -4.8625 20.935 ;
        RECT  -4.9325 20.8 -4.8625 20.935 ;
        RECT  -4.9325 20.8 -4.8625 20.935 ;
        RECT  -4.9325 20.8 -4.8625 20.935 ;
        RECT  -4.9325 20.8 -4.8625 20.935 ;
        RECT  -4.9325 20.8 -4.8625 20.935 ;
        RECT  -4.26 20.015 -4.125 20.085 ;
        RECT  -4.9325 20.0175 -4.8625 21.4275 ;
        RECT  -4.2225 20.02 -4.1625 20.0775 ;
        RECT  -4.405 20.025 -4.35 20.0775 ;
        RECT  -4.7425 20.0175 -4.685 20.0775 ;
        RECT  -4.9275 20.025 -4.8675 20.0825 ;
        RECT  -4.7475 19.95 -4.6775 21.495 ;
        RECT  -4.4125 19.95 -4.3425 21.495 ;
        RECT  -4.2275 19.95 -4.1575 21.495 ;
        RECT  -4.9325 19.95 -4.8625 21.495 ;
        RECT  -1.9775 21.1425 -1.9075 21.2775 ;
        RECT  -1.38 21.3825 -1.315 21.4525 ;
        RECT  -2.135 21.3825 -2.07 21.4525 ;
        RECT  -2.1025 21.3825 -1.3475 21.4525 ;
        RECT  -1.415 21.3825 -1.28 21.4525 ;
        RECT  -2.17 21.3825 -2.035 21.4525 ;
        RECT  -4.4125 24.28 -4.3425 24.345 ;
        RECT  -4.4125 22.74 -4.3425 24.315 ;
        RECT  -4.445 24.2775 -4.31 24.3475 ;
        RECT  -0.65 19.52 -0.58 19.585 ;
        RECT  -2.5575 19.5225 -2.4875 19.5875 ;
        RECT  -0.65 19.555 -0.58 21.5325 ;
        RECT  -2.5575 18.8975 -2.4875 19.555 ;
        RECT  -0.6825 19.5175 -0.5475 19.5875 ;
        RECT  -2.59 19.52 -2.455 19.59 ;
        RECT  -2.5925 24.1675 -2.5225 24.3025 ;
        RECT  -0.65 21.33 -0.58 21.465 ;
        RECT  -0.65 22.335 -0.58 22.405 ;
        RECT  -4.0275 22.335 -3.9575 22.405 ;
        RECT  -0.65 21.5325 -0.58 22.37 ;
        RECT  -2.1025 22.335 -0.615 22.405 ;
        RECT  -3.9925 22.335 -2.1025 22.405 ;
        RECT  -4.0275 20.465 -3.9575 22.37 ;
        RECT  -4.0275 22.3975 -3.9575 22.5325 ;
        RECT  -3.7375 22.0075 -3.6675 22.0725 ;
        RECT  -3.7375 17.8475 -3.6675 22.04 ;
        RECT  -3.77 22.005 -3.635 22.075 ;
        RECT  -3.7375 23.7675 -3.6675 23.8325 ;
        RECT  -3.7375 21.3675 -3.6675 23.8 ;
        RECT  -3.77 23.765 -3.635 23.835 ;
        RECT  -0.4175 20.6625 -0.3475 20.7275 ;
        RECT  -0.4175 16.165 -0.3475 16.23 ;
        RECT  -3.1075 16.1675 -3.0375 16.2325 ;
        RECT  -0.4175 16.2 -0.3475 20.695 ;
        RECT  -3.1075 16.2 -3.0375 17.46 ;
        RECT  -0.45 20.66 -0.315 20.73 ;
        RECT  -0.45 16.1625 -0.315 16.2325 ;
        RECT  -3.14 16.165 -3.005 16.235 ;
        RECT  -3.7725 26.2325 -3.7025 26.3675 ;
        RECT  -3.5275 23.93 -3.4575 23.995 ;
        RECT  -3.5275 25.01 -3.4575 25.075 ;
        RECT  -3.5275 23.9625 -3.4575 25.045 ;
        RECT  -3.56 23.9275 -3.425 23.9975 ;
        RECT  -3.56 25.0075 -3.425 25.0775 ;
        RECT  -3.7375 28.345 -3.6675 28.41 ;
        RECT  -3.7375 26.2325 -3.6675 28.38 ;
        RECT  -3.77 28.3425 -3.635 28.4125 ;
        RECT  -3.5275 23.93 -3.4575 23.995 ;
        RECT  -3.5275 22.6 -3.4575 22.665 ;
        RECT  -3.5275 22.635 -3.4575 23.9625 ;
        RECT  -3.56 23.9275 -3.425 23.9975 ;
        RECT  -3.56 22.5975 -3.425 22.6675 ;
        RECT  -3.7375 31.035 -3.6675 31.1 ;
        RECT  -3.7375 26.2325 -3.6675 31.07 ;
        RECT  -3.77 31.0325 -3.635 31.1025 ;
        RECT  -4.9325 20.6625 -4.8625 20.7275 ;
        RECT  -4.9325 15.96 -4.8625 20.695 ;
        RECT  -4.965 20.66 -4.83 20.73 ;
        RECT  -4.2275 20.6625 -4.1575 20.7275 ;
        RECT  -4.2275 15.96 -4.1575 20.695 ;
        RECT  -4.26 20.66 -4.125 20.73 ;
        RECT  -1.9775 16.605 -1.9075 17.055 ;
        RECT  -2.6475 16.255 -2.5775 16.73 ;
        RECT  -2.7875 16.255 -2.7175 16.92 ;
        RECT  -2.7175 16.85 -2.5775 16.92 ;
        RECT  -2.1125 16.605 -1.9775 16.675 ;
        RECT  -2.1125 16.985 -1.9775 17.055 ;
        RECT  -2.7125 16.66 -2.5775 16.73 ;
        RECT  -2.7175 16.215 -2.6475 16.35 ;
        RECT  -2.7125 16.85 -2.5775 16.92 ;
        RECT  -2.8575 16.215 -2.7875 16.35 ;
        RECT  -4.1725 16.605 -4.1025 17.055 ;
        RECT  -3.5025 16.255 -3.4325 16.73 ;
        RECT  -3.3625 16.255 -3.2925 16.92 ;
        RECT  -3.5025 16.85 -3.3625 16.92 ;
        RECT  -4.2375 16.605 -4.1025 16.675 ;
        RECT  -4.2375 16.985 -4.1025 17.055 ;
        RECT  -3.6375 16.66 -3.5025 16.73 ;
        RECT  -3.5025 16.215 -3.4325 16.35 ;
        RECT  -3.6375 16.85 -3.5025 16.92 ;
        RECT  -3.3625 16.215 -3.2925 16.35 ;
        RECT  -4.0 14.615 -3.93 14.75 ;
        RECT  -4.0 15.105 -3.93 15.24 ;
        RECT  -4.155 14.615 -4.085 14.75 ;
        RECT  -4.155 15.315 -4.085 15.45 ;
        RECT  -5.565 14.615 -5.495 14.75 ;
        RECT  -5.565 15.525 -5.495 15.66 ;
        RECT  -4.55 14.615 -4.48 14.75 ;
        RECT  -4.55 15.735 -4.48 15.87 ;
        RECT  -1.3275 15.315 -1.2575 15.45 ;
        RECT  -0.7975 15.945 -0.7275 16.08 ;
        RECT  -2.1225 15.945 -2.0525 16.08 ;
        RECT  -2.645 15.315 -2.575 15.45 ;
        RECT  -2.785 15.525 -2.715 15.66 ;
        RECT  -4.0275 15.945 -3.9575 16.08 ;
        RECT  -3.505 15.735 -3.435 15.87 ;
        RECT  -3.365 15.525 -3.295 15.66 ;
        RECT  -0.9975 9.85 -0.9325 9.92 ;
        RECT  -0.2225 9.85 -0.1575 9.92 ;
        RECT  -0.22 15.135 -0.155 15.205 ;
        RECT  -0.965 9.85 -0.1875 9.92 ;
        RECT  -0.35 15.135 -0.1875 15.205 ;
        RECT  -1.0 9.8175 -0.93 9.9525 ;
        RECT  -0.225 9.8175 -0.155 9.9525 ;
        RECT  -0.2225 15.1025 -0.1525 15.2375 ;
        RECT  -2.4925 19.405 -2.4225 19.54 ;
        RECT  -3.6575 19.195 -3.5875 19.33 ;
        RECT  -0.9675 19.615 -0.8975 19.75 ;
        RECT  -0.2075 19.435 -0.1425 19.505 ;
        RECT  -0.35 19.435 -0.1725 19.505 ;
        RECT  -0.21 19.4025 -0.14 19.5375 ;
        RECT  -2.0425 19.645 -1.9075 19.715 ;
        RECT  -2.0425 21.245 -1.9075 21.315 ;
        RECT  -1.73 19.825 -1.66 19.96 ;
        RECT  -4.42 19.825 -4.35 19.96 ;
        RECT  -0.385 14.895 -0.315 15.03 ;
        RECT  -0.965 13.41 -0.9 13.48 ;
        RECT  -2.0875 13.41 -2.0225 13.48 ;
        RECT  -2.0525 13.41 -0.9325 13.48 ;
        RECT  -0.9675 13.3775 -0.8975 13.5125 ;
        RECT  -2.09 13.3775 -2.02 13.5125 ;
        RECT  -2.085 8.275 -2.015 8.41 ;
        RECT  -2.085 8.275 -2.015 8.41 ;
        RECT  -0.275 15.975 -0.14 16.045 ;
        RECT  -0.8675 8.415 -0.7975 8.55 ;
        RECT  -0.275 8.415 -0.14 8.485 ;
        RECT  -1.0825 16.865 -0.9475 16.935 ;
        RECT  -0.275 16.865 -0.14 16.935 ;
        RECT  -0.275 19.225 -0.14 19.295 ;
        RECT  -1.035 17.335 -0.9 17.405 ;
        RECT  -0.275 17.335 -0.14 17.405 ;
        RECT  9.665 8.275 9.8 8.345 ;
        RECT  10.295 15.975 10.43 16.045 ;
        RECT  10.085 8.415 10.22 8.485 ;
        RECT  9.875 16.865 10.01 16.935 ;
        RECT  10.505 19.225 10.64 19.295 ;
        RECT  10.715 17.335 10.85 17.405 ;
        RECT  0.0 19.855 0.205 19.99 ;
        RECT  8.89 20.695 9.095 20.83 ;
        RECT  -0.415 20.695 -0.28 20.765 ;
        Layer  via2 ; 
        RECT  11.4425 18.79 11.5125 18.86 ;
        RECT  12.1475 18.79 12.2175 18.86 ;
        RECT  11.4475 9.87 11.5175 9.94 ;
        RECT  12.1525 9.87 12.2225 9.94 ;
        RECT  11.4475 3.43 11.5175 3.5 ;
        RECT  12.1525 3.43 12.2225 3.5 ;
        RECT  11.4475 3.5825 11.5175 3.6525 ;
        RECT  12.1525 3.5825 12.2225 3.6525 ;
        RECT  0.945 7.4525 1.015 7.5225 ;
        RECT  0.945 6.7475 1.015 6.8175 ;
        RECT  0.945 6.0425 1.015 6.1125 ;
        RECT  0.945 5.3375 1.015 5.4075 ;
        RECT  11.24 0.3125 11.305 0.3775 ;
        RECT  11.945 0.3125 12.01 0.3775 ;
        RECT  11.45 0.035 11.515 0.1 ;
        RECT  12.155 0.035 12.22 0.1 ;
        RECT  8.5425 7.4875 8.6075 7.5525 ;
        RECT  7.115 7.455 7.18 7.52 ;
        RECT  8.3325 6.7825 8.3975 6.8475 ;
        RECT  7.115 6.75 7.18 6.815 ;
        RECT  8.1225 6.0775 8.1875 6.1425 ;
        RECT  7.115 6.045 7.18 6.11 ;
        RECT  7.9125 5.3725 7.9775 5.4375 ;
        RECT  7.115 5.34 7.18 5.405 ;
        RECT  1.015 7.63 1.08 7.695 ;
        RECT  9.7325 8.015 9.7975 8.08 ;
        RECT  -5.4125 8.31 -5.3425 8.38 ;
        RECT  -4.7075 8.31 -4.6375 8.38 ;
        RECT  -4.0025 8.31 -3.9325 8.38 ;
        RECT  -1.0 22.8125 -0.935 22.8775 ;
        RECT  -2.52 22.8125 -2.455 22.8775 ;
        RECT  -2.0075 19.6475 -1.9425 19.7125 ;
        RECT  -2.0075 21.2475 -1.9425 21.3125 ;
        RECT  -2.0825 8.31 -2.0175 8.375 ;
        RECT  -0.24 15.9775 -0.175 16.0425 ;
        RECT  -0.24 8.4175 -0.175 8.4825 ;
        RECT  -0.24 16.8675 -0.175 16.9325 ;
        RECT  -0.24 19.2275 -0.175 19.2925 ;
        RECT  -0.24 17.3375 -0.175 17.4025 ;
        RECT  9.7 8.2775 9.765 8.3425 ;
        RECT  10.33 15.9775 10.395 16.0425 ;
        RECT  10.12 8.4175 10.185 8.4825 ;
        RECT  9.91 16.8675 9.975 16.9325 ;
        RECT  10.54 19.2275 10.605 19.2925 ;
        RECT  10.75 17.3375 10.815 17.4025 ;
        RECT  8.89 20.73 8.955 20.795 ;
        RECT  9.03 20.73 9.095 20.795 ;
        RECT  -0.38 20.6975 -0.315 20.7625 ;
        Layer  metal3 ; 
        RECT  -2.0525 8.275 9.73 8.345 ;
        RECT  -0.14 15.975 10.36 16.045 ;
        RECT  -0.14 8.415 10.15 8.485 ;
        RECT  -0.14 16.865 9.94 16.935 ;
        RECT  -0.14 19.225 10.57 19.295 ;
        RECT  -0.14 17.335 10.78 17.405 ;
        RECT  -0.28 20.695 8.89 20.765 ;
        RECT  11.4475 0.0 11.5175 3.22 ;
        RECT  12.1525 0.0 12.2225 3.22 ;
        RECT  7.215 7.4525 8.61 7.5225 ;
        RECT  7.215 6.7475 8.4 6.8175 ;
        RECT  7.215 6.0425 8.19 6.1125 ;
        RECT  7.215 5.3375 7.98 5.4075 ;
        RECT  0.0 7.4525 0.9825 7.5225 ;
        RECT  0.0 6.7475 0.9825 6.8175 ;
        RECT  0.0 6.0425 0.9825 6.1125 ;
        RECT  0.0 5.3375 0.9825 5.4075 ;
        RECT  11.4425 18.755 11.5125 18.895 ;
        RECT  12.1475 18.755 12.2175 18.895 ;
        RECT  11.4475 9.835 11.5175 9.975 ;
        RECT  12.1525 9.835 12.2225 9.975 ;
        RECT  11.4475 3.395 11.5175 3.535 ;
        RECT  12.1525 3.395 12.2225 3.535 ;
        RECT  11.4475 3.5475 11.5175 3.6875 ;
        RECT  12.1525 3.5475 12.2225 3.6875 ;
        RECT  0.91 7.4525 1.05 7.5225 ;
        RECT  0.91 6.7475 1.05 6.8175 ;
        RECT  0.91 6.0425 1.05 6.1125 ;
        RECT  0.91 5.3375 1.05 5.4075 ;
        RECT  11.2375 18.7325 11.3075 18.8025 ;
        RECT  11.2375 0.3125 11.3075 18.7675 ;
        RECT  11.2725 18.7325 11.5125 18.8025 ;
        RECT  11.2375 0.2775 11.3075 0.4125 ;
        RECT  11.9425 18.7325 12.0125 18.8025 ;
        RECT  11.9425 0.3125 12.0125 18.7675 ;
        RECT  11.9775 18.7325 12.2175 18.8025 ;
        RECT  11.9425 0.2775 12.0125 0.4125 ;
        RECT  11.4475 0.0 11.5175 0.135 ;
        RECT  12.1525 0.0 12.2225 0.135 ;
        RECT  8.54 7.4525 8.61 7.5875 ;
        RECT  7.08 7.4525 7.215 7.5225 ;
        RECT  8.33 6.7475 8.4 6.8825 ;
        RECT  7.08 6.7475 7.215 6.8175 ;
        RECT  8.12 6.0425 8.19 6.1775 ;
        RECT  7.08 6.0425 7.215 6.1125 ;
        RECT  7.91 5.3375 7.98 5.4725 ;
        RECT  7.08 5.3375 7.215 5.4075 ;
        RECT  0.98 7.6275 1.115 7.6975 ;
        RECT  1.08 7.98 1.15 8.05 ;
        RECT  1.08 7.6275 1.15 8.015 ;
        RECT  1.115 7.98 9.7325 8.05 ;
        RECT  9.73 7.98 9.8 8.115 ;
        RECT  -1.9775 19.645 -1.9075 21.2775 ;
        RECT  -5.4125 8.275 -5.3425 8.415 ;
        RECT  -4.7075 8.275 -4.6375 8.415 ;
        RECT  -4.0025 8.275 -3.9325 8.415 ;
        RECT  -1.0025 22.81 -0.9325 22.88 ;
        RECT  -2.5225 22.81 -2.4525 22.88 ;
        RECT  -2.4875 22.81 -0.9675 22.88 ;
        RECT  -1.0025 22.7775 -0.9325 22.9125 ;
        RECT  -2.5225 22.7775 -2.4525 22.9125 ;
        RECT  -2.0425 19.645 -1.9075 19.715 ;
        RECT  -2.0425 21.245 -1.9075 21.315 ;
        RECT  -2.085 8.275 -2.015 8.41 ;
        RECT  -0.275 15.975 -0.14 16.045 ;
        RECT  -0.275 8.415 -0.14 8.485 ;
        RECT  -0.275 16.865 -0.14 16.935 ;
        RECT  -0.275 19.225 -0.14 19.295 ;
        RECT  -0.275 17.335 -0.14 17.405 ;
        RECT  9.665 8.275 9.8 8.345 ;
        RECT  10.295 15.975 10.43 16.045 ;
        RECT  10.085 8.415 10.22 8.485 ;
        RECT  9.875 16.865 10.01 16.935 ;
        RECT  10.505 19.225 10.64 19.295 ;
        RECT  10.715 17.335 10.85 17.405 ;
        RECT  8.89 20.695 9.095 20.83 ;
        RECT  -0.415 20.695 -0.28 20.765 ;
    END 
END    sram_2_16_1_freepdk45 
END    LIBRARY 
