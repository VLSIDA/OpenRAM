magic
tech scmos
timestamp 1539900829
<< nwell >>
rect -18 -1 32 26
<< pwell >>
rect -18 -51 32 -6
<< ntransistor >>
rect -6 -18 -4 -12
rect 2 -24 4 -12
rect 10 -24 12 -12
rect 18 -18 20 -12
rect -6 -36 -4 -28
rect 2 -36 4 -28
rect 10 -36 12 -28
rect 18 -36 20 -28
<< ptransistor >>
rect 2 5 4 9
rect 10 5 12 9
<< ndiffusion >>
rect -11 -14 -6 -12
rect -7 -18 -6 -14
rect -4 -18 -3 -12
rect 1 -20 2 -12
rect -3 -24 2 -20
rect 4 -24 5 -12
rect 9 -24 10 -12
rect 12 -20 13 -12
rect 17 -18 18 -12
rect 20 -14 25 -12
rect 20 -18 21 -14
rect 12 -24 17 -20
rect -11 -30 -6 -28
rect -7 -34 -6 -30
rect -11 -36 -6 -34
rect -4 -36 2 -28
rect 4 -36 5 -28
rect 9 -36 10 -28
rect 12 -36 18 -28
rect 20 -30 25 -28
rect 20 -34 21 -30
rect 20 -36 25 -34
<< pdiffusion >>
rect 1 5 2 9
rect 4 5 5 9
rect 9 5 10 9
rect 12 5 13 9
<< ndcontact >>
rect -11 -18 -7 -14
rect -3 -20 1 -12
rect 5 -24 9 -12
rect 13 -20 17 -12
rect 21 -18 25 -14
rect -11 -34 -7 -30
rect 5 -36 9 -28
rect 21 -34 25 -30
<< pdcontact >>
rect -3 5 1 9
rect 5 5 9 9
rect 13 5 17 9
<< psubstratepcontact >>
rect 5 -44 9 -40
<< nsubstratencontact >>
rect 5 19 9 23
<< polysilicon >>
rect 2 9 4 11
rect 10 9 12 11
rect 2 -5 4 5
rect 10 2 12 5
rect 11 -2 12 2
rect -6 -12 -4 -7
rect 2 -9 3 -5
rect 2 -12 4 -9
rect 10 -12 12 -2
rect 18 -12 20 -7
rect -6 -20 -4 -18
rect 18 -20 20 -18
rect -6 -28 -4 -27
rect 2 -28 4 -24
rect 10 -28 12 -24
rect 18 -28 20 -27
rect -6 -38 -4 -36
rect 2 -38 4 -36
rect 10 -38 12 -36
rect 18 -38 20 -36
<< polycontact >>
rect 7 -2 11 2
rect -10 -11 -6 -7
rect 3 -9 7 -5
rect 20 -11 24 -7
rect -8 -27 -4 -23
rect 18 -27 22 -23
<< metal1 >>
rect -18 19 5 23
rect 9 19 32 23
rect -18 12 32 16
rect -10 -7 -6 12
rect -3 2 0 5
rect -3 -2 7 2
rect -3 -12 0 -2
rect 14 -5 17 5
rect 7 -9 17 -5
rect 14 -12 17 -9
rect 20 -7 24 12
rect -14 -18 -11 -14
rect 25 -18 28 -14
rect 5 -28 9 -24
rect 5 -40 9 -36
rect -17 -44 5 -40
rect 9 -44 31 -40
rect -17 -51 -4 -47
rect 0 -51 14 -47
rect 18 -51 31 -47
<< m2contact >>
rect 5 19 9 23
rect 5 5 9 9
rect -18 -18 -14 -14
rect -4 -27 0 -23
rect 28 -18 32 -14
rect 14 -27 18 -23
rect -11 -34 -7 -30
rect 21 -34 25 -30
rect -4 -51 0 -47
rect 14 -51 18 -47
<< metal2 >>
rect -18 -14 -14 23
rect -18 -51 -14 -18
rect -11 -30 -7 23
rect 5 9 9 19
rect -11 -51 -7 -34
rect -4 -47 0 -27
rect 14 -47 18 -27
rect 21 -30 25 23
rect 21 -51 25 -34
rect 28 -14 32 23
rect 28 -51 32 -18
<< labels >>
rlabel metal1 7 -49 7 -49 1 wl1
rlabel psubstratepcontact 7 -42 7 -42 1 gnd
rlabel m2contact 7 21 7 21 5 vdd
rlabel metal1 -1 14 -1 14 1 wl0
rlabel metal2 -16 -46 -16 -46 2 bl0
rlabel metal2 -9 -46 -9 -46 1 bl1
rlabel metal2 23 -46 23 -46 1 br1
rlabel metal2 30 -46 30 -46 8 br0
<< end >>
