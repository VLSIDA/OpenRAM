magic
tech scmos
timestamp 1680718477
<< nwell >>
rect 0 28 40 153
<< pwell >>
rect 0 153 40 214
rect 0 0 40 28
<< ntransistor >>
rect 21 181 23 190
rect 12 159 14 168
rect 20 159 22 168
rect 13 10 15 22
rect 21 18 23 22
<< ptransistor >>
rect 12 129 14 147
rect 20 129 22 147
rect 11 71 13 95
rect 27 71 29 95
rect 13 34 15 58
rect 21 34 23 42
<< ndiffusion >>
rect 20 181 21 190
rect 23 181 24 190
rect 11 159 12 168
rect 14 159 15 168
rect 19 159 20 168
rect 22 159 23 168
rect 12 10 13 22
rect 15 10 16 22
rect 20 18 21 22
rect 23 18 24 22
<< pdiffusion >>
rect 7 145 12 147
rect 11 131 12 145
rect 7 129 12 131
rect 14 145 20 147
rect 14 131 15 145
rect 19 131 20 145
rect 14 129 20 131
rect 22 145 27 147
rect 22 131 23 145
rect 22 129 27 131
rect 10 71 11 95
rect 13 71 14 95
rect 26 71 27 95
rect 29 71 30 95
rect 12 34 13 58
rect 15 34 16 58
rect 20 34 21 42
rect 23 34 24 42
<< ndcontact >>
rect 16 181 20 190
rect 24 181 28 190
rect 7 159 11 168
rect 15 159 19 168
rect 23 159 27 168
rect 8 10 12 22
rect 16 10 20 22
rect 24 18 28 22
<< pdcontact >>
rect 7 131 11 145
rect 15 131 19 145
rect 23 131 27 145
rect 6 71 10 95
rect 14 71 18 95
rect 22 71 26 95
rect 30 71 34 95
rect 8 34 12 58
rect 16 34 20 58
rect 24 34 28 42
<< psubstratepcontact >>
rect 32 188 36 192
rect 28 4 32 8
<< nsubstratencontact >>
rect 27 121 31 125
rect 27 55 31 59
<< polysilicon >>
rect 21 190 23 200
rect 21 180 23 181
rect 3 178 23 180
rect 3 98 5 178
rect 12 173 34 175
rect 12 168 14 173
rect 20 168 22 170
rect 12 147 14 159
rect 20 147 22 159
rect 32 156 34 173
rect 30 152 34 156
rect 12 127 14 129
rect 20 120 22 129
rect 13 118 22 120
rect 9 106 11 116
rect 32 106 34 152
rect 33 102 34 106
rect 3 96 13 98
rect 11 95 13 96
rect 27 95 29 97
rect 11 70 13 71
rect 27 70 29 71
rect 11 68 29 70
rect 7 63 23 65
rect 13 58 15 60
rect 21 42 23 63
rect 13 31 15 34
rect 13 27 14 31
rect 13 22 15 27
rect 21 22 23 34
rect 21 16 23 18
rect 13 8 15 10
<< polycontact >>
rect 20 200 24 204
rect 26 152 30 156
rect 9 116 13 120
rect 9 102 13 106
rect 29 102 33 106
rect 3 63 7 67
rect 14 27 18 31
<< metal1 >>
rect -2 200 20 204
rect 24 200 36 204
rect 28 184 32 188
rect 16 168 19 181
rect 7 145 11 159
rect 23 156 27 159
rect 23 152 26 156
rect 7 120 11 131
rect 15 145 19 147
rect 15 129 19 131
rect 23 145 27 152
rect 23 129 27 131
rect 15 126 18 129
rect 15 125 31 126
rect 15 123 27 125
rect 7 116 9 120
rect 6 95 9 105
rect 33 102 34 106
rect 31 95 34 102
rect 3 71 6 74
rect 3 67 7 71
rect 20 55 27 58
rect 8 22 11 34
rect 24 30 28 34
rect 18 27 28 30
rect 24 22 28 27
rect 3 10 8 13
rect 3 9 10 10
rect 3 8 7 9
rect 16 7 20 10
rect 16 4 28 7
<< m2contact >>
rect 32 184 36 188
rect 27 117 31 121
rect 13 95 17 99
rect 22 95 26 99
rect 27 51 31 55
rect 3 4 7 8
rect 28 8 32 12
<< metal2 >>
rect 10 99 14 214
rect 20 99 24 214
rect 32 180 36 184
rect 27 113 31 117
rect 10 95 13 99
rect 20 95 22 99
rect 3 0 7 4
rect 10 0 14 95
rect 20 0 24 95
rect 27 47 31 51
rect 28 12 32 16
<< bb >>
rect 0 0 34 214
<< labels >>
rlabel metal2 5 2 5 2 1 dout
rlabel metal2 30 14 30 14 1 gnd
rlabel metal2 29 49 29 49 1 vdd
rlabel metal2 22 212 22 212 5 br
rlabel metal2 12 212 12 212 5 bl
rlabel metal2 29 115 29 115 1 vdd
rlabel metal2 34 182 34 182 1 gnd
flabel metal1 0 200 0 200 4 FreeSans 26 0 0 0 en
<< properties >>
string path 270.000 468.000 270.000 486.000 288.000 486.000 288.000 468.000 270.000 468.000 
<< end >>
