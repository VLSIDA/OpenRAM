
.SUBCKT row_cap_cell_1rw_1r wl0 wl1 gnd

.ENDS
