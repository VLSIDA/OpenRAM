magic
tech sky130A
magscale 1 2
timestamp 1595931502
<< checkpaint >>
rect -1319 -1316 1685 1714
<< nwell >>
rect -54 -54 420 454
<< scpmos >>
rect 60 0 90 400
rect 168 0 198 400
rect 276 0 306 400
<< pdiff >>
rect 0 0 60 400
rect 90 0 168 400
rect 198 0 276 400
rect 306 0 366 400
<< poly >>
rect 60 400 90 426
rect 168 400 198 426
rect 276 400 306 426
rect 60 -26 90 0
rect 168 -26 198 0
rect 276 -26 306 0
rect 60 -56 306 -26
<< locali >>
rect 8 167 42 233
rect 112 133 146 200
rect 220 167 254 233
rect 324 133 358 200
rect 112 99 358 133
use contact_11  contact_11_3
timestamp 1595931502
transform 1 0 0 0 1 167
box -59 -51 109 117
use contact_11  contact_11_2
timestamp 1595931502
transform 1 0 104 0 1 167
box -59 -51 109 117
use contact_11  contact_11_1
timestamp 1595931502
transform 1 0 212 0 1 167
box -59 -51 109 117
use contact_11  contact_11_0
timestamp 1595931502
transform 1 0 316 0 1 167
box -59 -51 109 117
<< labels >>
rlabel poly s 183 -41 183 -41 4 G
rlabel corelocali s 25 200 25 200 4 S
rlabel corelocali s 237 200 237 200 4 S
rlabel corelocali s 235 116 235 116 4 D
<< properties >>
string FIXED_BBOX -54 -54 420 454
<< end >>
