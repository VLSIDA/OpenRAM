VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO sram_1rw1r_2_16_sky130
   CLASS BLOCK ;
   SIZE 152.02 BY 140.435 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  34.45 0.125 34.75 0.425 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  40.29 0.125 40.59 0.425 ;
      END
   END din0[1]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER m3 ;
         RECT  0.53 111.505 0.83 111.805 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER m3 ;
         RECT  0.53 120.005 0.83 120.305 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER m3 ;
         RECT  0.53 125.645 0.83 125.945 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER m3 ;
         RECT  0.53 134.145 0.83 134.445 ;
      END
   END addr0[3]
   PIN addr1[0]
      DIRECTION INPUT ;
      PORT
         LAYER m3 ;
         RECT  151.82 42.965 152.12 43.265 ;
      END
   END addr1[0]
   PIN addr1[1]
      DIRECTION INPUT ;
      PORT
         LAYER m3 ;
         RECT  151.82 34.465 152.12 34.765 ;
      END
   END addr1[1]
   PIN addr1[2]
      DIRECTION INPUT ;
      PORT
         LAYER m3 ;
         RECT  151.82 28.825 152.12 29.125 ;
      END
   END addr1[2]
   PIN addr1[3]
      DIRECTION INPUT ;
      PORT
         LAYER m3 ;
         RECT  151.82 20.325 152.12 20.625 ;
      END
   END addr1[3]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER m3 ;
         RECT  0.53 2.945 0.83 3.245 ;
      END
   END csb0
   PIN csb1
      DIRECTION INPUT ;
      PORT
         LAYER m3 ;
         RECT  151.82 137.385 152.12 137.685 ;
      END
   END csb1
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER m3 ;
         RECT  0.53 11.445 0.83 11.745 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  16.035 0.125 16.335 0.425 ;
      END
   END clk0
   PIN clk1
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  136.735 140.205 137.035 140.505 ;
      END
   END clk1
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER m4 ;
         RECT  35.07 0.125 35.37 0.425 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER m4 ;
         RECT  40.91 0.125 41.21 0.425 ;
      END
   END dout0[1]
   PIN dout1[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER m4 ;
         RECT  74.245 140.205 74.545 140.505 ;
      END
   END dout1[0]
   PIN dout1[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER m4 ;
         RECT  78.595 140.205 78.895 140.505 ;
      END
   END dout1[1]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER m3 ;
         RECT  0.0 25.16 26.22 25.54 ;
         LAYER m4 ;
         RECT  133.96 0.0 134.34 139.78 ;
         LAYER m3 ;
         RECT  0.0 108.12 23.5 108.5 ;
         LAYER m3 ;
         RECT  24.745 115.66 25.235 116.15 ;
         LAYER m3 ;
         RECT  0.0 127.16 152.02 127.54 ;
         LAYER m4 ;
         RECT  51.0 0.0 51.38 139.78 ;
         LAYER m4 ;
         RECT  105.4 0.0 105.78 139.78 ;
         LAYER m3 ;
         RECT  7.48 79.56 37.78 79.94 ;
         LAYER m3 ;
         RECT  86.36 64.6 152.02 64.98 ;
         LAYER m3 ;
         RECT  105.4 80.92 152.02 81.3 ;
         LAYER m3 ;
         RECT  78.79 55.58 79.28 56.07 ;
         LAYER m3 ;
         RECT  98.045 63.46 98.535 63.95 ;
         LAYER m3 ;
         RECT  109.115 63.46 109.605 63.95 ;
         LAYER m3 ;
         RECT  101.3 69.545 101.79 70.035 ;
         LAYER m3 ;
         RECT  86.36 70.04 98.3 70.42 ;
         LAYER m3 ;
         RECT  101.32 72.76 152.02 73.14 ;
         LAYER m3 ;
         RECT  28.56 42.84 123.46 43.22 ;
         LAYER m3 ;
         RECT  151.725 133.04 152.215 133.53 ;
         LAYER m3 ;
         RECT  86.36 86.36 144.54 86.74 ;
         LAYER m4 ;
         RECT  135.32 0.0 135.7 139.78 ;
         LAYER m3 ;
         RECT  25.84 136.68 135.02 137.06 ;
         LAYER m3 ;
         RECT  0.0 30.6 152.02 30.98 ;
         LAYER m4 ;
         RECT  113.56 0.0 113.94 139.78 ;
         LAYER m4 ;
         RECT  102.68 0.0 103.06 139.78 ;
         LAYER m3 ;
         RECT  80.72 98.7 81.21 99.19 ;
         LAYER m3 ;
         RECT  118.985 75.31 119.475 75.8 ;
         LAYER m3 ;
         RECT  55.76 67.32 98.3 67.7 ;
         LAYER m3 ;
         RECT  80.24 113.56 152.02 113.94 ;
         LAYER m3 ;
         RECT  55.225 63.46 55.715 63.95 ;
         LAYER m4 ;
         RECT  48.28 0.0 48.66 139.78 ;
         LAYER m3 ;
         RECT  98.045 85.185 98.535 85.675 ;
         LAYER m3 ;
         RECT  86.36 63.24 98.3 63.62 ;
         LAYER m4 ;
         RECT  72.76 0.0 73.14 139.78 ;
         LAYER m4 ;
         RECT  139.4 0.0 139.78 139.78 ;
         LAYER m3 ;
         RECT  9.52 71.4 48.66 71.78 ;
         LAYER m3 ;
         RECT  0.0 121.72 152.02 122.1 ;
         LAYER m3 ;
         RECT  145.805 91.29 146.295 91.78 ;
         LAYER m3 ;
         RECT  0.0 44.2 124.14 44.58 ;
         LAYER m3 ;
         RECT  17.0 3.4 152.02 3.78 ;
         LAYER m3 ;
         RECT  70.04 65.96 83.34 66.34 ;
         LAYER m4 ;
         RECT  64.6 0.0 64.98 139.78 ;
         LAYER m3 ;
         RECT  51.97 63.495 52.46 63.985 ;
         LAYER m3 ;
         RECT  55.76 65.96 67.02 66.34 ;
         LAYER m3 ;
         RECT  140.08 139.4 152.02 139.78 ;
         LAYER m3 ;
         RECT  78.88 40.12 152.02 40.5 ;
         LAYER m3 ;
         RECT  51.97 73.495 52.46 73.985 ;
         LAYER m3 ;
         RECT  44.155 67.41 44.645 67.9 ;
         LAYER m3 ;
         RECT  0.0 51.0 62.94 51.38 ;
         LAYER m3 ;
         RECT  9.52 65.96 48.66 66.34 ;
         LAYER m4 ;
         RECT  91.8 0.0 92.18 139.78 ;
         LAYER m3 ;
         RECT  67.32 38.76 152.02 39.14 ;
         LAYER m3 ;
         RECT  98.045 71.36 98.535 71.85 ;
         LAYER m4 ;
         RECT  74.12 0.0 74.5 112.58 ;
         LAYER m3 ;
         RECT  55.225 69.385 55.715 69.875 ;
         LAYER m3 ;
         RECT  140.76 123.08 152.02 123.46 ;
         LAYER m4 ;
         RECT  38.76 0.0 39.14 139.78 ;
         LAYER m3 ;
         RECT  0.0 75.48 31.66 75.86 ;
         LAYER m3 ;
         RECT  75.42 112.31 75.91 112.8 ;
         LAYER m3 ;
         RECT  55.76 63.24 67.02 63.62 ;
         LAYER m3 ;
         RECT  55.76 79.56 67.02 79.94 ;
         LAYER m3 ;
         RECT  55.76 89.08 67.02 89.46 ;
         LAYER m3 ;
         RECT  2.675 85.39 3.165 85.88 ;
         LAYER m3 ;
         RECT  0.0 132.6 129.58 132.98 ;
         LAYER m3 ;
         RECT  55.225 71.36 55.715 71.85 ;
         LAYER m3 ;
         RECT  71.955 58.535 72.445 59.025 ;
         LAYER m4 ;
         RECT  87.72 0.0 88.1 139.78 ;
         LAYER m4 ;
         RECT  36.04 0.0 36.42 139.78 ;
         LAYER m3 ;
         RECT  0.0 64.6 67.02 64.98 ;
         LAYER m3 ;
         RECT  0.0 95.88 141.82 96.26 ;
         LAYER m3 ;
         RECT  0.0 21.08 122.1 21.46 ;
         LAYER m3 ;
         RECT  98.045 79.26 98.535 79.75 ;
         LAYER m3 ;
         RECT  78.29 58.63 78.59 58.93 ;
         LAYER m3 ;
         RECT  86.36 89.08 98.3 89.46 ;
         LAYER m3 ;
         RECT  70.04 61.88 83.34 62.26 ;
         LAYER m3 ;
         RECT  105.4 83.64 142.5 84.02 ;
         LAYER m3 ;
         RECT  127.84 27.88 152.02 28.26 ;
         LAYER m3 ;
         RECT  9.52 60.52 67.02 60.9 ;
         LAYER m4 ;
         RECT  29.24 0.0 29.62 139.78 ;
         LAYER m3 ;
         RECT  0.0 128.52 132.98 128.9 ;
         LAYER m3 ;
         RECT  0.0 6.12 152.02 6.5 ;
         LAYER m4 ;
         RECT  142.12 0.0 142.5 139.78 ;
         LAYER m3 ;
         RECT  0.0 36.04 73.82 36.42 ;
         LAYER m3 ;
         RECT  127.84 114.92 152.02 115.3 ;
         LAYER m3 ;
         RECT  0.0 131.24 152.02 131.62 ;
         LAYER m3 ;
         RECT  77.29 46.16 77.78 46.65 ;
         LAYER m3 ;
         RECT  19.72 11.56 152.02 11.94 ;
         LAYER m4 ;
         RECT  8.84 0.0 9.22 139.78 ;
         LAYER m3 ;
         RECT  70.04 94.52 83.34 94.9 ;
         LAYER m3 ;
         RECT  55.225 67.41 55.715 67.9 ;
         LAYER m3 ;
         RECT  59.58 77.06 60.07 77.55 ;
         LAYER m3 ;
         RECT  10.2 59.16 152.02 59.54 ;
         LAYER m3 ;
         RECT  105.4 71.4 142.5 71.78 ;
         LAYER m4 ;
         RECT  55.08 0.0 55.46 139.78 ;
         LAYER m4 ;
         RECT  98.6 0.0 98.98 139.78 ;
         LAYER m3 ;
         RECT  9.52 76.84 48.66 77.22 ;
         LAYER m3 ;
         RECT  0.0 45.56 127.54 45.94 ;
         LAYER m3 ;
         RECT  86.36 60.52 142.5 60.9 ;
         LAYER m3 ;
         RECT  0.0 112.2 26.22 112.58 ;
         LAYER m4 ;
         RECT  11.56 0.0 11.94 139.78 ;
         LAYER m3 ;
         RECT  112.37 75.345 112.86 75.835 ;
         LAYER m3 ;
         RECT  101.32 90.44 152.02 90.82 ;
         LAYER m3 ;
         RECT  101.3 67.445 101.79 67.935 ;
         LAYER m3 ;
         RECT  7.48 68.68 67.02 69.06 ;
         LAYER m4 ;
         RECT  114.92 0.0 115.3 139.78 ;
         LAYER m3 ;
         RECT  0.0 63.24 31.66 63.62 ;
         LAYER m3 ;
         RECT  77.23 112.31 77.72 112.8 ;
         LAYER m3 ;
         RECT  68.0 25.16 152.02 25.54 ;
         LAYER m3 ;
         RECT  105.4 70.04 152.02 70.42 ;
         LAYER m4 ;
         RECT  136.68 0.0 137.06 135.7 ;
         LAYER m3 ;
         RECT  0.0 40.12 73.82 40.5 ;
         LAYER m3 ;
         RECT  86.36 82.28 152.02 82.66 ;
         LAYER m4 ;
         RECT  59.16 0.0 59.54 139.78 ;
         LAYER m3 ;
         RECT  118.985 63.46 119.475 63.95 ;
         LAYER m3 ;
         RECT  112.37 63.495 112.86 63.985 ;
         LAYER m3 ;
         RECT  149.485 46.49 149.975 46.98 ;
         LAYER m3 ;
         RECT  105.4 65.96 142.5 66.34 ;
         LAYER m4 ;
         RECT  151.64 0.0 152.02 139.78 ;
         LAYER m3 ;
         RECT  0.0 80.92 48.66 81.3 ;
         LAYER m3 ;
         RECT  51.97 91.145 52.46 91.635 ;
         LAYER m3 ;
         RECT  130.56 31.96 152.02 32.34 ;
         LAYER m3 ;
         RECT  0.0 117.64 152.02 118.02 ;
         LAYER m3 ;
         RECT  86.36 87.72 98.3 88.1 ;
         LAYER m3 ;
         RECT  79.56 36.04 152.02 36.42 ;
         LAYER m3 ;
         RECT  101.3 87.195 101.79 87.685 ;
         LAYER m3 ;
         RECT  17.68 42.84 26.22 43.22 ;
         LAYER m3 ;
         RECT  9.52 82.28 67.02 82.66 ;
         LAYER m3 ;
         RECT  127.84 108.12 152.02 108.5 ;
         LAYER m3 ;
         RECT  44.2 12.92 152.02 13.3 ;
         LAYER m4 ;
         RECT  40.12 17.0 40.5 139.78 ;
         LAYER m3 ;
         RECT  0.0 12.92 35.06 13.3 ;
         LAYER m3 ;
         RECT  0.0 61.88 67.02 62.26 ;
         LAYER m4 ;
         RECT  86.36 0.0 86.74 139.78 ;
         LAYER m3 ;
         RECT  46.92 14.28 152.02 14.66 ;
         LAYER m3 ;
         RECT  25.84 123.08 131.62 123.46 ;
         LAYER m4 ;
         RECT  23.8 0.0 24.18 139.78 ;
         LAYER m3 ;
         RECT  86.36 75.48 98.3 75.86 ;
         LAYER m3 ;
         RECT  116.28 79.56 152.02 79.94 ;
         LAYER m3 ;
         RECT  30.6 119.0 152.02 119.38 ;
         LAYER m3 ;
         RECT  70.04 82.28 83.34 82.66 ;
         LAYER m3 ;
         RECT  7.48 57.8 152.02 58.18 ;
         LAYER m3 ;
         RECT  0.0 85.0 48.66 85.38 ;
         LAYER m3 ;
         RECT  42.265 19.965 42.755 20.455 ;
         LAYER m4 ;
         RECT  104.04 0.0 104.42 139.78 ;
         LAYER m3 ;
         RECT  101.3 85.345 101.79 85.835 ;
         LAYER m3 ;
         RECT  0.0 129.88 152.02 130.26 ;
         LAYER m3 ;
         RECT  44.155 79.26 44.645 79.75 ;
         LAYER m3 ;
         RECT  101.3 65.595 101.79 66.085 ;
         LAYER m3 ;
         RECT  0.0 7.48 11.26 7.86 ;
         LAYER m3 ;
         RECT  0.0 101.32 72.46 101.7 ;
         LAYER m4 ;
         RECT  83.64 0.0 84.02 139.78 ;
         LAYER m4 ;
         RECT  143.48 0.0 143.86 139.78 ;
         LAYER m3 ;
         RECT  101.3 71.395 101.79 71.885 ;
         LAYER m3 ;
         RECT  7.48 90.44 52.74 90.82 ;
         LAYER m4 ;
         RECT  78.2 0.0 78.58 112.58 ;
         LAYER m4 ;
         RECT  31.96 0.0 32.34 139.78 ;
         LAYER m3 ;
         RECT  28.56 27.88 122.78 28.26 ;
         LAYER m3 ;
         RECT  75.17 95.84 75.47 96.14 ;
         LAYER m4 ;
         RECT  34.68 17.0 35.06 139.78 ;
         LAYER m3 ;
         RECT  0.0 27.88 26.22 28.26 ;
         LAYER m3 ;
         RECT  0.0 52.36 7.86 52.74 ;
         LAYER m3 ;
         RECT  126.445 133.04 126.935 133.53 ;
         LAYER m3 ;
         RECT  42.84 0.68 152.02 1.06 ;
         LAYER m3 ;
         RECT  23.12 7.48 152.02 7.86 ;
         LAYER m3 ;
         RECT  9.52 99.96 152.02 100.34 ;
         LAYER m4 ;
         RECT  49.64 0.0 50.02 139.78 ;
         LAYER m3 ;
         RECT  86.36 65.96 98.3 66.34 ;
         LAYER m3 ;
         RECT  86.36 93.16 152.02 93.54 ;
         LAYER m3 ;
         RECT  109.115 67.41 109.605 67.9 ;
         LAYER m3 ;
         RECT  141.44 132.6 152.02 132.98 ;
         LAYER m3 ;
         RECT  0.0 94.52 67.02 94.9 ;
         LAYER m3 ;
         RECT  24.745 129.8 25.235 130.29 ;
         LAYER m3 ;
         RECT  25.84 108.12 86.06 108.5 ;
         LAYER m3 ;
         RECT  55.76 90.44 67.02 90.82 ;
         LAYER m3 ;
         RECT  78.29 95.84 78.59 96.14 ;
         LAYER m4 ;
         RECT  30.6 0.0 30.98 139.78 ;
         LAYER m3 ;
         RECT  86.36 72.76 98.3 73.14 ;
         LAYER m3 ;
         RECT  34.285 75.31 34.775 75.8 ;
         LAYER m3 ;
         RECT  86.36 85.0 98.3 85.38 ;
         LAYER m3 ;
         RECT  0.0 123.08 23.5 123.46 ;
         LAYER m3 ;
         RECT  0.0 119.0 26.22 119.38 ;
         LAYER m4 ;
         RECT  110.84 0.0 111.22 139.78 ;
         LAYER m3 ;
         RECT  70.04 91.8 83.34 92.18 ;
         LAYER m3 ;
         RECT  0.0 138.04 137.06 138.42 ;
         LAYER m4 ;
         RECT  7.48 0.0 7.86 139.78 ;
         LAYER m3 ;
         RECT  77.29 108.12 77.78 108.61 ;
         LAYER m3 ;
         RECT  70.04 72.76 83.34 73.14 ;
         LAYER m3 ;
         RECT  0.0 38.76 26.22 39.14 ;
         LAYER m3 ;
         RECT  55.225 83.21 55.715 83.7 ;
         LAYER m3 ;
         RECT  0.0 22.44 152.02 22.82 ;
         LAYER m3 ;
         RECT  0.0 26.52 152.02 26.9 ;
         LAYER m3 ;
         RECT  126.445 118.9 126.935 119.39 ;
         LAYER m3 ;
         RECT  55.76 71.4 67.02 71.78 ;
         LAYER m3 ;
         RECT  0.0 86.36 67.02 86.74 ;
         LAYER m3 ;
         RECT  86.36 71.4 98.3 71.78 ;
         LAYER m3 ;
         RECT  98.045 91.11 98.535 91.6 ;
         LAYER m3 ;
         RECT  98.045 75.31 98.535 75.8 ;
         LAYER m3 ;
         RECT  51.97 89.295 52.46 89.785 ;
         LAYER m3 ;
         RECT  105.4 91.8 152.02 92.18 ;
         LAYER m3 ;
         RECT  86.36 61.88 152.02 62.26 ;
         LAYER m3 ;
         RECT  75.17 58.63 75.47 58.93 ;
         LAYER m3 ;
         RECT  149.485 80.09 149.975 80.58 ;
         LAYER m3 ;
         RECT  70.04 70.04 83.34 70.42 ;
         LAYER m3 ;
         RECT  74.795 34.21 75.285 34.7 ;
         LAYER m3 ;
         RECT  105.4 76.84 142.5 77.22 ;
         LAYER m3 ;
         RECT  138.72 136.68 152.02 137.06 ;
         LAYER m3 ;
         RECT  0.0 109.48 152.02 109.86 ;
         LAYER m4 ;
         RECT  117.64 0.0 118.02 139.78 ;
         LAYER m3 ;
         RECT  70.04 85.0 83.34 85.38 ;
         LAYER m3 ;
         RECT  27.245 49.52 27.735 50.01 ;
         LAYER m3 ;
         RECT  0.0 46.92 152.02 47.3 ;
         LAYER m4 ;
         RECT  52.36 0.0 52.74 139.78 ;
         LAYER m3 ;
         RECT  55.76 91.8 67.02 92.18 ;
         LAYER m3 ;
         RECT  70.04 76.84 83.34 77.22 ;
         LAYER m3 ;
         RECT  0.0 97.24 124.82 97.62 ;
         LAYER m3 ;
         RECT  86.36 74.12 98.3 74.5 ;
         LAYER m3 ;
         RECT  27.245 21.24 27.735 21.73 ;
         LAYER m3 ;
         RECT  70.04 83.64 83.34 84.02 ;
         LAYER m4 ;
         RECT  17.0 0.0 17.38 139.78 ;
         LAYER m4 ;
         RECT  131.24 0.0 131.62 139.78 ;
         LAYER m4 ;
         RECT  70.04 0.0 70.42 139.78 ;
         LAYER m4 ;
         RECT  125.8 0.0 126.18 139.78 ;
         LAYER m3 ;
         RECT  98.045 73.335 98.535 73.825 ;
         LAYER m3 ;
         RECT  70.04 87.72 83.34 88.1 ;
         LAYER m3 ;
         RECT  70.04 75.48 83.34 75.86 ;
         LAYER m3 ;
         RECT  55.225 87.16 55.715 87.65 ;
         LAYER m3 ;
         RECT  55.225 89.135 55.715 89.625 ;
         LAYER m3 ;
         RECT  55.225 65.435 55.715 65.925 ;
         LAYER m3 ;
         RECT  0.0 42.84 10.58 43.22 ;
         LAYER m3 ;
         RECT  0.0 49.64 74.5 50.02 ;
         LAYER m3 ;
         RECT  28.56 56.44 152.02 56.82 ;
         LAYER m3 ;
         RECT  142.8 138.04 152.02 138.42 ;
         LAYER m4 ;
         RECT  26.52 0.0 26.9 139.78 ;
         LAYER m3 ;
         RECT  6.355 62.99 6.845 63.48 ;
         LAYER m4 ;
         RECT  21.08 0.0 21.46 139.78 ;
         LAYER m4 ;
         RECT  127.16 0.0 127.54 139.78 ;
         LAYER m3 ;
         RECT  77.855 34.21 78.345 34.7 ;
         LAYER m3 ;
         RECT  98.045 65.435 98.535 65.925 ;
         LAYER m3 ;
         RECT  55.76 80.92 67.02 81.3 ;
         LAYER m4 ;
         RECT  144.84 0.0 145.22 139.78 ;
         LAYER m3 ;
         RECT  51.97 85.345 52.46 85.835 ;
         LAYER m4 ;
         RECT  25.16 0.0 25.54 139.78 ;
         LAYER m3 ;
         RECT  9.52 93.16 67.02 93.54 ;
         LAYER m3 ;
         RECT  145.805 46.49 146.295 46.98 ;
         LAYER m3 ;
         RECT  74.48 98.7 74.97 99.19 ;
         LAYER m3 ;
         RECT  105.4 74.12 144.54 74.5 ;
         LAYER m4 ;
         RECT  45.56 0.0 45.94 139.78 ;
         LAYER m3 ;
         RECT  81.315 58.535 81.805 59.025 ;
         LAYER m3 ;
         RECT  105.4 87.72 142.5 88.1 ;
         LAYER m3 ;
         RECT  55.76 72.76 67.02 73.14 ;
         LAYER m3 ;
         RECT  145.805 80.09 146.295 80.58 ;
         LAYER m3 ;
         RECT  0.0 29.24 129.58 29.62 ;
         LAYER m3 ;
         RECT  70.04 89.08 83.34 89.46 ;
         LAYER m4 ;
         RECT  148.92 0.0 149.3 139.78 ;
         LAYER m3 ;
         RECT  51.97 67.445 52.46 67.935 ;
         LAYER m3 ;
         RECT  70.04 68.68 83.34 69.06 ;
         LAYER m3 ;
         RECT  101.3 79.295 101.79 79.785 ;
         LAYER m3 ;
         RECT  2.04 11.56 9.9 11.94 ;
         LAYER m3 ;
         RECT  0.0 113.56 72.46 113.94 ;
         LAYER m3 ;
         RECT  2.675 107.79 3.165 108.28 ;
         LAYER m4 ;
         RECT  37.4 0.0 37.78 139.78 ;
         LAYER m3 ;
         RECT  0.0 31.96 26.22 32.34 ;
         LAYER m3 ;
         RECT  44.155 63.46 44.645 63.95 ;
         LAYER m3 ;
         RECT  2.04 3.4 14.66 3.78 ;
         LAYER m3 ;
         RECT  70.04 71.4 83.34 71.78 ;
         LAYER m3 ;
         RECT  15.64 4.76 152.02 5.14 ;
         LAYER m3 ;
         RECT  51.97 87.195 52.46 87.685 ;
         LAYER m4 ;
         RECT  120.36 0.0 120.74 139.78 ;
         LAYER m4 ;
         RECT  108.12 0.0 108.5 139.78 ;
         LAYER m3 ;
         RECT  98.045 87.16 98.535 87.65 ;
         LAYER m3 ;
         RECT  86.36 91.8 98.3 92.18 ;
         LAYER m4 ;
         RECT  121.72 0.0 122.1 139.78 ;
         LAYER m3 ;
         RECT  27.245 7.1 27.735 7.59 ;
         LAYER m3 ;
         RECT  116.28 67.32 152.02 67.7 ;
         LAYER m3 ;
         RECT  0.0 53.72 26.22 54.1 ;
         LAYER m4 ;
         RECT  14.28 0.0 14.66 139.78 ;
         LAYER m3 ;
         RECT  0.0 8.84 152.02 9.22 ;
         LAYER m3 ;
         RECT  72.55 55.58 73.04 56.07 ;
         LAYER m3 ;
         RECT  86.36 68.68 152.02 69.06 ;
         LAYER m3 ;
         RECT  77.755 29.46 78.245 29.95 ;
         LAYER m3 ;
         RECT  6.355 85.39 6.845 85.88 ;
         LAYER m3 ;
         RECT  55.76 70.04 67.02 70.42 ;
         LAYER m4 ;
         RECT  140.76 0.0 141.14 139.78 ;
         LAYER m4 ;
         RECT  109.48 0.0 109.86 139.78 ;
         LAYER m3 ;
         RECT  0.0 74.12 48.66 74.5 ;
         LAYER m4 ;
         RECT  82.28 0.0 82.66 139.78 ;
         LAYER m4 ;
         RECT  112.2 0.0 112.58 139.78 ;
         LAYER m3 ;
         RECT  109.115 79.26 109.605 79.75 ;
         LAYER m3 ;
         RECT  0.0 2.04 152.02 2.42 ;
         LAYER m4 ;
         RECT  67.32 0.0 67.7 139.78 ;
         LAYER m4 ;
         RECT  2.04 0.0 2.42 139.78 ;
         LAYER m4 ;
         RECT  99.96 0.0 100.34 139.78 ;
         LAYER m3 ;
         RECT  0.0 124.44 152.02 124.82 ;
         LAYER m3 ;
         RECT  101.3 83.245 101.79 83.735 ;
         LAYER m3 ;
         RECT  44.155 75.31 44.645 75.8 ;
         LAYER m4 ;
         RECT  97.24 0.0 97.62 139.78 ;
         LAYER m3 ;
         RECT  40.9 67.445 41.39 67.935 ;
         LAYER m3 ;
         RECT  55.76 75.48 67.02 75.86 ;
         LAYER m3 ;
         RECT  27.245 35.38 27.735 35.87 ;
         LAYER m4 ;
         RECT  0.68 0.0 1.06 139.78 ;
         LAYER m3 ;
         RECT  81.6 51.0 152.02 51.38 ;
         LAYER m3 ;
         RECT  133.28 44.2 152.02 44.58 ;
         LAYER m4 ;
         RECT  75.48 0.0 75.86 139.78 ;
         LAYER m3 ;
         RECT  128.52 125.8 152.02 126.18 ;
         LAYER m3 ;
         RECT  75.36 46.16 75.85 46.65 ;
         LAYER m4 ;
         RECT  12.92 0.0 13.3 139.78 ;
         LAYER m3 ;
         RECT  101.3 73.495 101.79 73.985 ;
         LAYER m3 ;
         RECT  65.96 53.72 152.02 54.1 ;
         LAYER m4 ;
         RECT  68.68 0.0 69.06 139.78 ;
         LAYER m4 ;
         RECT  63.24 0.0 63.62 139.78 ;
         LAYER m3 ;
         RECT  98.045 69.385 98.535 69.875 ;
         LAYER m4 ;
         RECT  41.48 1.36 41.86 139.78 ;
         LAYER m3 ;
         RECT  23.8 120.36 152.02 120.74 ;
         LAYER m4 ;
         RECT  71.4 0.0 71.78 139.78 ;
         LAYER m4 ;
         RECT  76.84 0.0 77.22 139.78 ;
         LAYER m3 ;
         RECT  0.435 7.1 0.925 7.59 ;
         LAYER m4 ;
         RECT  56.44 0.0 56.82 139.78 ;
         LAYER m4 ;
         RECT  57.8 0.0 58.18 139.78 ;
         LAYER m3 ;
         RECT  101.3 63.495 101.79 63.985 ;
         LAYER m3 ;
         RECT  70.04 93.16 83.34 93.54 ;
         LAYER m3 ;
         RECT  79.56 31.96 127.54 32.34 ;
         LAYER m3 ;
         RECT  86.36 78.2 102.38 78.58 ;
         LAYER m3 ;
         RECT  105.4 85.0 152.02 85.38 ;
         LAYER m3 ;
         RECT  0.0 55.08 142.5 55.46 ;
         LAYER m3 ;
         RECT  89.76 104.04 152.02 104.42 ;
         LAYER m3 ;
         RECT  98.045 77.285 98.535 77.775 ;
         LAYER m3 ;
         RECT  98.045 81.235 98.535 81.725 ;
         LAYER m3 ;
         RECT  2.675 62.99 3.165 63.48 ;
         LAYER m3 ;
         RECT  78.88 49.64 142.5 50.02 ;
         LAYER m3 ;
         RECT  81.315 95.745 81.805 96.235 ;
         LAYER m3 ;
         RECT  51.97 83.245 52.46 83.735 ;
         LAYER m3 ;
         RECT  36.425 19.965 36.915 20.455 ;
         LAYER m3 ;
         RECT  0.0 48.28 152.02 48.66 ;
         LAYER m3 ;
         RECT  126.445 104.76 126.935 105.25 ;
         LAYER m3 ;
         RECT  1.36 0.68 13.3 1.06 ;
         LAYER m3 ;
         RECT  70.04 60.52 83.34 60.9 ;
         LAYER m3 ;
         RECT  30.6 112.2 124.82 112.58 ;
         LAYER m3 ;
         RECT  78.79 98.7 79.28 99.19 ;
         LAYER m3 ;
         RECT  0.0 17.0 127.54 17.38 ;
         LAYER m3 ;
         RECT  55.76 85.0 67.02 85.38 ;
         LAYER m3 ;
         RECT  86.36 83.64 98.3 84.02 ;
         LAYER m3 ;
         RECT  128.52 97.24 144.54 97.62 ;
         LAYER m3 ;
         RECT  1.36 14.28 26.22 14.66 ;
         LAYER m3 ;
         RECT  55.225 91.11 55.715 91.6 ;
         LAYER m4 ;
         RECT  123.08 0.0 123.46 139.78 ;
         LAYER m4 ;
         RECT  27.88 0.0 28.26 139.78 ;
         LAYER m3 ;
         RECT  127.84 21.08 152.02 21.46 ;
         LAYER m3 ;
         RECT  51.97 81.395 52.46 81.885 ;
         LAYER m3 ;
         RECT  51.97 69.545 52.46 70.035 ;
         LAYER m3 ;
         RECT  6.355 74.19 6.845 74.68 ;
         LAYER m3 ;
         RECT  0.0 104.04 72.46 104.42 ;
         LAYER m3 ;
         RECT  149.485 57.69 149.975 58.18 ;
         LAYER m3 ;
         RECT  40.9 79.295 41.39 79.785 ;
         LAYER m3 ;
         RECT  55.76 74.12 67.02 74.5 ;
         LAYER m3 ;
         RECT  0.0 135.32 136.38 135.7 ;
         LAYER m4 ;
         RECT  85.0 0.0 85.38 139.78 ;
         LAYER m3 ;
         RECT  0.0 37.4 152.02 37.78 ;
         LAYER m4 ;
         RECT  3.4 0.0 3.78 139.78 ;
         LAYER m4 ;
         RECT  119.0 0.0 119.38 139.78 ;
         LAYER m3 ;
         RECT  70.04 80.92 83.34 81.3 ;
         LAYER m3 ;
         RECT  89.115 77.14 89.605 77.63 ;
         LAYER m3 ;
         RECT  105.4 89.08 152.02 89.46 ;
         LAYER m4 ;
         RECT  89.08 0.0 89.46 139.78 ;
         LAYER m4 ;
         RECT  4.76 0.0 5.14 139.78 ;
         LAYER m3 ;
         RECT  40.9 63.495 41.39 63.985 ;
         LAYER m3 ;
         RECT  74.895 29.46 75.385 29.95 ;
         LAYER m4 ;
         RECT  80.92 0.0 81.3 139.78 ;
         LAYER m4 ;
         RECT  93.16 0.0 93.54 139.78 ;
         LAYER m3 ;
         RECT  0.0 136.68 23.5 137.06 ;
         LAYER m4 ;
         RECT  79.56 0.0 79.94 139.78 ;
         LAYER m4 ;
         RECT  33.32 0.0 33.7 139.78 ;
         LAYER m3 ;
         RECT  130.56 17.0 152.02 17.38 ;
         LAYER m3 ;
         RECT  0.0 23.8 152.02 24.18 ;
         LAYER m4 ;
         RECT  132.6 0.0 132.98 139.78 ;
         LAYER m3 ;
         RECT  70.04 63.24 83.34 63.62 ;
         LAYER m3 ;
         RECT  0.0 87.72 48.66 88.1 ;
         LAYER m4 ;
         RECT  138.04 0.0 138.42 139.78 ;
         LAYER m3 ;
         RECT  0.0 114.92 85.38 115.3 ;
         LAYER m4 ;
         RECT  65.96 0.0 66.34 139.78 ;
         LAYER m3 ;
         RECT  128.945 24.48 129.435 24.97 ;
         LAYER m3 ;
         RECT  127.84 101.32 152.02 101.7 ;
         LAYER m3 ;
         RECT  71.955 95.745 72.445 96.235 ;
         LAYER m3 ;
         RECT  0.0 116.28 152.02 116.66 ;
         LAYER m3 ;
         RECT  101.3 75.345 101.79 75.835 ;
         LAYER m3 ;
         RECT  55.76 83.64 67.02 84.02 ;
         LAYER m3 ;
         RECT  55.225 75.31 55.715 75.8 ;
         LAYER m3 ;
         RECT  109.115 75.31 109.605 75.8 ;
         LAYER m3 ;
         RECT  70.04 86.36 83.34 86.74 ;
         LAYER m4 ;
         RECT  44.2 0.0 44.58 139.78 ;
         LAYER m3 ;
         RECT  0.0 83.64 48.66 84.02 ;
         LAYER m3 ;
         RECT  122.4 75.48 152.02 75.86 ;
         LAYER m3 ;
         RECT  70.04 64.6 83.34 64.98 ;
         LAYER m3 ;
         RECT  7.48 102.68 78.58 103.06 ;
         LAYER m4 ;
         RECT  124.44 0.0 124.82 139.78 ;
         LAYER m3 ;
         RECT  2.675 74.19 3.165 74.68 ;
         LAYER m3 ;
         RECT  98.045 67.41 98.535 67.9 ;
         LAYER m3 ;
         RECT  149.485 91.29 149.975 91.78 ;
         LAYER m3 ;
         RECT  6.355 107.79 6.845 108.28 ;
         LAYER m3 ;
         RECT  14.28 10.2 152.02 10.58 ;
         LAYER m3 ;
         RECT  9.52 105.4 152.02 105.78 ;
         LAYER m4 ;
         RECT  116.28 0.0 116.66 139.78 ;
         LAYER m3 ;
         RECT  64.155 77.14 64.645 77.63 ;
         LAYER m4 ;
         RECT  106.76 0.0 107.14 139.78 ;
         LAYER m3 ;
         RECT  9.52 89.08 48.66 89.46 ;
         LAYER m3 ;
         RECT  70.04 90.44 83.34 90.82 ;
         LAYER m3 ;
         RECT  31.28 125.8 124.82 126.18 ;
         LAYER m3 ;
         RECT  34.285 63.46 34.775 63.95 ;
         LAYER m3 ;
         RECT  75.42 41.97 75.91 42.46 ;
         LAYER m4 ;
         RECT  53.72 0.0 54.1 139.78 ;
         LAYER m3 ;
         RECT  77.23 41.97 77.72 42.46 ;
         LAYER m3 ;
         RECT  51.97 75.345 52.46 75.835 ;
         LAYER m3 ;
         RECT  81.6 52.36 144.54 52.74 ;
         LAYER m3 ;
         RECT  51.97 79.295 52.46 79.785 ;
         LAYER m3 ;
         RECT  0.0 67.32 37.78 67.7 ;
         LAYER m3 ;
         RECT  101.3 81.395 101.79 81.885 ;
         LAYER m4 ;
         RECT  150.28 0.0 150.66 139.78 ;
         LAYER m3 ;
         RECT  0.0 18.36 152.02 18.74 ;
         LAYER m4 ;
         RECT  46.92 0.0 47.3 139.78 ;
         LAYER m3 ;
         RECT  0.0 15.64 33.02 16.02 ;
         LAYER m4 ;
         RECT  6.12 0.0 6.5 139.78 ;
         LAYER m3 ;
         RECT  128.52 112.2 152.02 112.58 ;
         LAYER m3 ;
         RECT  98.045 83.21 98.535 83.7 ;
         LAYER m3 ;
         RECT  0.0 139.4 127.54 139.78 ;
         LAYER m4 ;
         RECT  19.72 0.0 20.1 139.78 ;
         LAYER m3 ;
         RECT  0.0 33.32 73.82 33.7 ;
         LAYER m3 ;
         RECT  70.04 74.12 83.34 74.5 ;
         LAYER m3 ;
         RECT  0.0 34.68 122.78 35.06 ;
         LAYER m3 ;
         RECT  130.56 45.56 152.02 45.94 ;
         LAYER m3 ;
         RECT  29.92 110.84 152.02 111.22 ;
         LAYER m3 ;
         RECT  51.97 65.595 52.46 66.085 ;
         LAYER m3 ;
         RECT  40.9 75.345 41.39 75.835 ;
         LAYER m3 ;
         RECT  105.4 78.2 152.02 78.58 ;
         LAYER m4 ;
         RECT  101.32 0.0 101.7 139.78 ;
         LAYER m3 ;
         RECT  51.97 71.395 52.46 71.885 ;
         LAYER m3 ;
         RECT  98.045 89.135 98.535 89.625 ;
         LAYER m3 ;
         RECT  101.3 91.145 101.79 91.635 ;
         LAYER m3 ;
         RECT  0.0 78.2 48.66 78.58 ;
         LAYER m3 ;
         RECT  51.68 78.2 67.02 78.58 ;
         LAYER m3 ;
         RECT  86.36 90.44 98.3 90.82 ;
         LAYER m3 ;
         RECT  55.76 87.72 67.02 88.1 ;
         LAYER m4 ;
         RECT  146.2 0.0 146.58 139.78 ;
         LAYER m3 ;
         RECT  0.0 41.48 152.02 41.86 ;
         LAYER m4 ;
         RECT  61.88 0.0 62.26 139.78 ;
         LAYER m3 ;
         RECT  139.4 128.52 152.02 128.9 ;
         LAYER m3 ;
         RECT  55.225 85.185 55.715 85.675 ;
         LAYER m3 ;
         RECT  78.88 33.32 152.02 33.7 ;
         LAYER m4 ;
         RECT  90.44 0.0 90.82 139.78 ;
         LAYER m4 ;
         RECT  128.52 0.0 128.9 139.78 ;
         LAYER m3 ;
         RECT  0.0 19.72 129.58 20.1 ;
         LAYER m3 ;
         RECT  0.0 98.6 152.02 98.98 ;
         LAYER m3 ;
         RECT  128.945 38.62 129.435 39.11 ;
         LAYER m3 ;
         RECT  55.225 81.235 55.715 81.725 ;
         LAYER m4 ;
         RECT  147.56 0.0 147.94 139.78 ;
         LAYER m3 ;
         RECT  0.0 91.8 48.66 92.18 ;
         LAYER m3 ;
         RECT  75.36 108.12 75.85 108.61 ;
         LAYER m3 ;
         RECT  112.37 79.295 112.86 79.785 ;
         LAYER m3 ;
         RECT  55.225 79.26 55.715 79.75 ;
         LAYER m3 ;
         RECT  122.4 63.24 144.54 63.62 ;
         LAYER m3 ;
         RECT  145.805 68.89 146.295 69.38 ;
         LAYER m4 ;
         RECT  18.36 0.0 18.74 139.78 ;
         LAYER m3 ;
         RECT  51.97 77.445 52.46 77.935 ;
         LAYER m3 ;
         RECT  31.28 133.96 152.02 134.34 ;
         LAYER m3 ;
         RECT  70.04 79.56 83.34 79.94 ;
         LAYER m3 ;
         RECT  86.36 80.92 98.3 81.3 ;
         LAYER m3 ;
         RECT  149.485 68.89 149.975 69.38 ;
         LAYER m4 ;
         RECT  15.64 4.76 16.02 139.78 ;
         LAYER m4 ;
         RECT  42.84 0.0 43.22 139.78 ;
         LAYER m3 ;
         RECT  0.0 72.76 52.74 73.14 ;
         LAYER m3 ;
         RECT  112.37 67.445 112.86 67.935 ;
         LAYER m4 ;
         RECT  94.52 0.0 94.9 139.78 ;
         LAYER m3 ;
         RECT  55.225 73.335 55.715 73.825 ;
         LAYER m3 ;
         RECT  101.3 77.445 101.79 77.935 ;
         LAYER m4 ;
         RECT  129.88 0.0 130.26 139.78 ;
         LAYER m3 ;
         RECT  42.16 15.64 152.02 16.02 ;
         LAYER m3 ;
         RECT  93.69 77.06 94.18 77.55 ;
         LAYER m3 ;
         RECT  101.3 89.295 101.79 89.785 ;
         LAYER m3 ;
         RECT  55.225 77.285 55.715 77.775 ;
         LAYER m3 ;
         RECT  0.0 106.76 152.02 107.14 ;
         LAYER m3 ;
         RECT  6.355 96.59 6.845 97.08 ;
         LAYER m3 ;
         RECT  86.36 79.56 98.3 79.94 ;
         LAYER m3 ;
         RECT  70.04 78.2 83.34 78.58 ;
         LAYER m3 ;
         RECT  0.0 70.04 48.66 70.42 ;
         LAYER m3 ;
         RECT  74.48 55.58 74.97 56.07 ;
         LAYER m4 ;
         RECT  95.88 0.0 96.26 139.78 ;
         LAYER m3 ;
         RECT  0.0 56.44 26.22 56.82 ;
         LAYER m4 ;
         RECT  22.44 0.0 22.82 139.78 ;
         LAYER m3 ;
         RECT  145.805 57.69 146.295 58.18 ;
         LAYER m4 ;
         RECT  60.52 0.0 60.9 139.78 ;
         LAYER m3 ;
         RECT  2.675 96.59 3.165 97.08 ;
         LAYER m4 ;
         RECT  10.2 0.0 10.58 139.78 ;
         LAYER m3 ;
         RECT  86.36 94.52 142.5 94.9 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER m3 ;
         RECT  103.425 75.345 103.915 75.835 ;
         LAYER m3 ;
         RECT  49.845 71.395 50.335 71.885 ;
         LAYER m3 ;
         RECT  57.12 78.88 96.94 79.26 ;
         LAYER m3 ;
         RECT  0.0 115.6 23.5 115.98 ;
         LAYER m3 ;
         RECT  0.0 73.44 50.7 73.82 ;
         LAYER m3 ;
         RECT  0.0 136.0 136.38 136.38 ;
         LAYER m4 ;
         RECT  74.8 0.0 75.18 112.58 ;
         LAYER m3 ;
         RECT  74.85 36.395 75.34 36.885 ;
         LAYER m4 ;
         RECT  122.4 0.0 122.78 139.78 ;
         LAYER m3 ;
         RECT  0.0 57.12 144.54 57.5 ;
         LAYER m3 ;
         RECT  103.425 81.385 103.915 81.875 ;
         LAYER m3 ;
         RECT  103.36 77.52 142.5 77.9 ;
         LAYER m3 ;
         RECT  140.76 122.4 152.02 122.78 ;
         LAYER m3 ;
         RECT  84.89 77.235 85.19 77.535 ;
         LAYER m3 ;
         RECT  0.0 68.0 39.82 68.38 ;
         LAYER m3 ;
         RECT  14.28 9.52 152.02 9.9 ;
         LAYER m3 ;
         RECT  68.57 91.85 68.87 92.15 ;
         LAYER m3 ;
         RECT  29.92 110.16 152.02 110.54 ;
         LAYER m3 ;
         RECT  49.845 89.285 50.335 89.775 ;
         LAYER m3 ;
         RECT  110.475 67.41 110.965 67.9 ;
         LAYER m4 ;
         RECT  34.0 17.0 34.38 139.78 ;
         LAYER m3 ;
         RECT  25.84 115.6 85.38 115.98 ;
         LAYER m3 ;
         RECT  0.0 19.04 152.02 19.42 ;
         LAYER m3 ;
         RECT  53.865 89.135 54.355 89.625 ;
         LAYER m3 ;
         RECT  80.92 55.76 152.02 56.14 ;
         LAYER m3 ;
         RECT  53.865 71.36 54.355 71.85 ;
         LAYER m3 ;
         RECT  84.89 64.2 85.19 64.5 ;
         LAYER m3 ;
         RECT  79.56 34.0 129.58 34.38 ;
         LAYER m3 ;
         RECT  145.805 74.49 146.295 74.98 ;
         LAYER m3 ;
         RECT  0.0 138.72 152.02 139.1 ;
         LAYER m4 ;
         RECT  100.64 0.0 101.02 139.78 ;
         LAYER m4 ;
         RECT  110.16 0.0 110.54 139.78 ;
         LAYER m3 ;
         RECT  49.845 79.295 50.335 79.785 ;
         LAYER m3 ;
         RECT  57.12 65.28 96.94 65.66 ;
         LAYER m3 ;
         RECT  127.84 115.6 152.02 115.98 ;
         LAYER m4 ;
         RECT  28.56 0.0 28.94 139.78 ;
         LAYER m4 ;
         RECT  88.4 0.0 88.78 139.78 ;
         LAYER m3 ;
         RECT  103.425 87.195 103.915 87.685 ;
         LAYER m4 ;
         RECT  115.6 0.0 115.98 139.78 ;
         LAYER m3 ;
         RECT  17.0 4.08 152.02 4.46 ;
         LAYER m3 ;
         RECT  80.24 114.24 152.02 114.62 ;
         LAYER m4 ;
         RECT  35.36 1.36 35.74 139.78 ;
         LAYER m3 ;
         RECT  57.12 82.96 96.94 83.34 ;
         LAYER m3 ;
         RECT  9.52 66.64 152.02 67.02 ;
         LAYER m4 ;
         RECT  4.08 0.0 4.46 139.78 ;
         LAYER m3 ;
         RECT  84.89 70.52 85.19 70.82 ;
         LAYER m3 ;
         RECT  10.2 58.48 70.42 58.86 ;
         LAYER m4 ;
         RECT  69.36 0.0 69.74 139.78 ;
         LAYER m4 ;
         RECT  59.84 0.0 60.22 139.78 ;
         LAYER m3 ;
         RECT  0.0 106.08 152.02 106.46 ;
         LAYER m3 ;
         RECT  84.89 76.05 85.19 76.35 ;
         LAYER m3 ;
         RECT  78.88 112.88 152.02 113.26 ;
         LAYER m3 ;
         RECT  84.89 69.335 85.19 69.635 ;
         LAYER m3 ;
         RECT  53.865 65.435 54.355 65.925 ;
         LAYER m3 ;
         RECT  77.825 31.54 78.315 32.03 ;
         LAYER m4 ;
         RECT  138.72 0.0 139.1 139.78 ;
         LAYER m3 ;
         RECT  77.25 32.55 77.74 33.04 ;
         LAYER m3 ;
         RECT  0.0 55.76 71.1 56.14 ;
         LAYER m4 ;
         RECT  61.2 0.0 61.58 139.78 ;
         LAYER m4 ;
         RECT  130.56 0.0 130.94 139.78 ;
         LAYER m3 ;
         RECT  66.64 31.28 152.02 31.66 ;
         LAYER m3 ;
         RECT  0.0 48.96 26.22 49.34 ;
         LAYER m3 ;
         RECT  84.89 65.385 85.19 65.685 ;
         LAYER m3 ;
         RECT  84.89 73.285 85.19 73.585 ;
         LAYER m4 ;
         RECT  5.44 0.0 5.82 139.78 ;
         LAYER m3 ;
         RECT  114.495 63.495 114.985 63.985 ;
         LAYER m4 ;
         RECT  81.6 0.0 81.98 139.78 ;
         LAYER m3 ;
         RECT  99.405 83.21 99.895 83.7 ;
         LAYER m3 ;
         RECT  0.0 35.36 26.22 35.74 ;
         LAYER m3 ;
         RECT  82.96 95.2 141.82 95.58 ;
         LAYER m3 ;
         RECT  84.89 91.85 85.19 92.15 ;
         LAYER m3 ;
         RECT  28.56 35.36 122.78 35.74 ;
         LAYER m3 ;
         RECT  27.245 42.45 27.735 42.94 ;
         LAYER m4 ;
         RECT  99.28 0.0 99.66 139.78 ;
         LAYER m3 ;
         RECT  114.24 78.88 152.02 79.26 ;
         LAYER m3 ;
         RECT  99.405 69.385 99.895 69.875 ;
         LAYER m4 ;
         RECT  10.88 0.0 11.26 139.78 ;
         LAYER m3 ;
         RECT  53.865 79.26 54.355 79.75 ;
         LAYER m3 ;
         RECT  103.425 65.585 103.915 66.075 ;
         LAYER m3 ;
         RECT  6.355 68.59 6.845 69.08 ;
         LAYER m3 ;
         RECT  9.52 70.72 50.7 71.1 ;
         LAYER m3 ;
         RECT  139.4 129.2 152.02 129.58 ;
         LAYER m4 ;
         RECT  111.52 0.0 111.9 139.78 ;
         LAYER m3 ;
         RECT  103.36 65.28 152.02 65.66 ;
         LAYER m3 ;
         RECT  0.0 14.96 26.9 15.34 ;
         LAYER m3 ;
         RECT  78.88 42.16 123.46 42.54 ;
         LAYER m3 ;
         RECT  0.0 43.52 10.58 43.9 ;
         LAYER m3 ;
         RECT  0.0 137.36 135.02 137.74 ;
         LAYER m3 ;
         RECT  68.57 60.25 68.87 60.55 ;
         LAYER m3 ;
         RECT  74.825 31.54 75.315 32.03 ;
         LAYER m3 ;
         RECT  0.0 95.2 70.42 95.58 ;
         LAYER m3 ;
         RECT  23.12 8.16 152.02 8.54 ;
         LAYER m3 ;
         RECT  0.0 87.04 50.7 87.42 ;
         LAYER m3 ;
         RECT  49.845 75.345 50.335 75.835 ;
         LAYER m3 ;
         RECT  114.495 67.445 114.985 67.935 ;
         LAYER m3 ;
         RECT  0.0 84.32 152.02 84.7 ;
         LAYER m4 ;
         RECT  29.92 0.0 30.3 139.78 ;
         LAYER m3 ;
         RECT  53.865 75.31 54.355 75.8 ;
         LAYER m3 ;
         RECT  99.405 77.285 99.895 77.775 ;
         LAYER m3 ;
         RECT  27.245 56.59 27.735 57.08 ;
         LAYER m4 ;
         RECT  42.16 0.0 42.54 139.78 ;
         LAYER m3 ;
         RECT  121.04 63.92 152.02 64.3 ;
         LAYER m3 ;
         RECT  21.08 17.68 152.02 18.06 ;
         LAYER m3 ;
         RECT  68.57 82.37 68.87 82.67 ;
         LAYER m3 ;
         RECT  9.52 77.52 50.7 77.9 ;
         LAYER m3 ;
         RECT  84.89 62.62 85.19 62.92 ;
         LAYER m3 ;
         RECT  0.0 108.8 73.82 109.18 ;
         LAYER m4 ;
         RECT  68.0 0.0 68.38 139.78 ;
         LAYER m4 ;
         RECT  25.84 0.0 26.22 139.78 ;
         LAYER m3 ;
         RECT  127.84 35.36 152.02 35.74 ;
         LAYER m3 ;
         RECT  99.405 73.335 99.895 73.825 ;
         LAYER m4 ;
         RECT  96.56 0.0 96.94 139.78 ;
         LAYER m3 ;
         RECT  84.89 68.15 85.19 68.45 ;
         LAYER m3 ;
         RECT  103.425 73.485 103.915 73.975 ;
         LAYER m3 ;
         RECT  25.84 129.2 132.98 129.58 ;
         LAYER m3 ;
         RECT  145.805 52.09 146.295 52.58 ;
         LAYER m4 ;
         RECT  129.2 0.0 129.58 139.78 ;
         LAYER m3 ;
         RECT  0.0 31.28 26.22 31.66 ;
         LAYER m3 ;
         RECT  67.32 39.44 152.02 39.82 ;
         LAYER m4 ;
         RECT  40.8 17.0 41.18 139.78 ;
         LAYER m4 ;
         RECT  57.12 0.0 57.5 139.78 ;
         LAYER m3 ;
         RECT  78.88 107.44 152.02 107.82 ;
         LAYER m3 ;
         RECT  0.0 116.96 152.02 117.34 ;
         LAYER m3 ;
         RECT  0.0 42.16 73.82 42.54 ;
         LAYER m3 ;
         RECT  68.57 64.2 68.87 64.5 ;
         LAYER m3 ;
         RECT  127.84 100.64 152.02 101.02 ;
         LAYER m3 ;
         RECT  49.845 63.495 50.335 63.985 ;
         LAYER m3 ;
         RECT  149.485 74.49 149.975 74.98 ;
         LAYER m3 ;
         RECT  2.675 90.99 3.165 91.48 ;
         LAYER m4 ;
         RECT  126.48 0.0 126.86 139.78 ;
         LAYER m3 ;
         RECT  57.12 87.04 96.94 87.42 ;
         LAYER m3 ;
         RECT  151.725 140.12 152.215 140.61 ;
         LAYER m3 ;
         RECT  53.865 73.335 54.355 73.825 ;
         LAYER m4 ;
         RECT  106.08 0.0 106.46 139.78 ;
         LAYER m3 ;
         RECT  68.57 61.435 68.87 61.735 ;
         LAYER m3 ;
         RECT  0.0 54.4 142.5 54.78 ;
         LAYER m4 ;
         RECT  78.88 0.0 79.26 112.58 ;
         LAYER m3 ;
         RECT  74.8 51.68 152.02 52.06 ;
         LAYER m4 ;
         RECT  123.76 0.0 124.14 139.78 ;
         LAYER m3 ;
         RECT  103.425 63.495 103.915 63.985 ;
         LAYER m4 ;
         RECT  133.28 0.0 133.66 139.78 ;
         LAYER m3 ;
         RECT  57.12 81.6 96.94 81.98 ;
         LAYER m4 ;
         RECT  107.44 0.0 107.82 139.78 ;
         LAYER m3 ;
         RECT  126.445 140.11 126.935 140.6 ;
         LAYER m3 ;
         RECT  149.485 96.89 149.975 97.38 ;
         LAYER m4 ;
         RECT  148.24 0.0 148.62 139.78 ;
         LAYER m3 ;
         RECT  65.96 77.52 88.1 77.9 ;
         LAYER m3 ;
         RECT  0.0 28.56 122.78 28.94 ;
         LAYER m3 ;
         RECT  0.0 16.32 33.02 16.7 ;
         LAYER m3 ;
         RECT  103.425 79.295 103.915 79.785 ;
         LAYER m4 ;
         RECT  85.68 0.0 86.06 139.78 ;
         LAYER m3 ;
         RECT  77.8 36.395 78.29 36.885 ;
         LAYER m3 ;
         RECT  6.355 90.99 6.845 91.48 ;
         LAYER m3 ;
         RECT  103.425 91.145 103.915 91.635 ;
         LAYER m3 ;
         RECT  19.72 12.24 152.02 12.62 ;
         LAYER m3 ;
         RECT  30.6 111.52 152.02 111.9 ;
         LAYER m4 ;
         RECT  19.04 0.0 19.42 139.78 ;
         LAYER m4 ;
         RECT  116.96 0.0 117.34 139.78 ;
         LAYER m4 ;
         RECT  114.24 0.0 114.62 139.78 ;
         LAYER m3 ;
         RECT  126.445 111.83 126.935 112.32 ;
         LAYER m3 ;
         RECT  84.89 60.25 85.19 60.55 ;
         LAYER m3 ;
         RECT  53.865 85.185 54.355 85.675 ;
         LAYER m3 ;
         RECT  68.0 24.48 127.54 24.86 ;
         LAYER m3 ;
         RECT  23.8 134.64 152.02 135.02 ;
         LAYER m3 ;
         RECT  49.845 85.335 50.335 85.825 ;
         LAYER m3 ;
         RECT  7.48 74.8 33.02 75.18 ;
         LAYER m3 ;
         RECT  0.0 127.84 152.02 128.22 ;
         LAYER m3 ;
         RECT  0.0 38.08 127.54 38.46 ;
         LAYER m4 ;
         RECT  46.24 0.0 46.62 139.78 ;
         LAYER m3 ;
         RECT  49.845 65.585 50.335 66.075 ;
         LAYER m3 ;
         RECT  99.405 63.46 99.895 63.95 ;
         LAYER m3 ;
         RECT  53.865 77.285 54.355 77.775 ;
         LAYER m4 ;
         RECT  31.28 0.0 31.66 139.78 ;
         LAYER m3 ;
         RECT  0.0 110.16 20.78 110.54 ;
         LAYER m4 ;
         RECT  108.8 0.0 109.18 139.78 ;
         LAYER m3 ;
         RECT  0.0 76.16 152.02 76.54 ;
         LAYER m4 ;
         RECT  27.2 0.0 27.58 139.78 ;
         LAYER m3 ;
         RECT  99.405 87.16 99.895 87.65 ;
         LAYER m3 ;
         RECT  145.805 63.29 146.295 63.78 ;
         LAYER m3 ;
         RECT  0.0 121.04 152.02 121.42 ;
         LAYER m3 ;
         RECT  2.675 68.59 3.165 69.08 ;
         LAYER m3 ;
         RECT  6.355 102.19 6.845 102.68 ;
         LAYER m3 ;
         RECT  42.265 12.895 42.755 13.385 ;
         LAYER m4 ;
         RECT  63.92 0.0 64.3 139.78 ;
         LAYER m3 ;
         RECT  84.89 90.27 85.19 90.57 ;
         LAYER m3 ;
         RECT  128.945 45.69 129.435 46.18 ;
         LAYER m3 ;
         RECT  0.0 91.12 50.7 91.5 ;
         LAYER m3 ;
         RECT  149.485 85.69 149.975 86.18 ;
         LAYER m3 ;
         RECT  53.865 81.235 54.355 81.725 ;
         LAYER m4 ;
         RECT  144.16 0.0 144.54 139.78 ;
         LAYER m3 ;
         RECT  42.16 16.32 152.02 16.7 ;
         LAYER m3 ;
         RECT  7.48 62.56 152.02 62.94 ;
         LAYER m3 ;
         RECT  38.775 67.445 39.265 67.935 ;
         LAYER m3 ;
         RECT  42.795 75.31 43.285 75.8 ;
         LAYER m3 ;
         RECT  2.675 57.39 3.165 57.88 ;
         LAYER m3 ;
         RECT  128.945 31.55 129.435 32.04 ;
         LAYER m3 ;
         RECT  103.36 82.96 142.5 83.34 ;
         LAYER m3 ;
         RECT  28.56 6.8 152.02 7.18 ;
         LAYER m3 ;
         RECT  7.48 85.68 50.7 86.06 ;
         LAYER m3 ;
         RECT  128.52 118.32 152.02 118.7 ;
         LAYER m3 ;
         RECT  53.865 67.41 54.355 67.9 ;
         LAYER m3 ;
         RECT  84.89 61.435 85.19 61.735 ;
         LAYER m3 ;
         RECT  84.89 89.085 85.19 89.385 ;
         LAYER m3 ;
         RECT  68.57 80.0 68.87 80.3 ;
         LAYER m3 ;
         RECT  53.865 63.46 54.355 63.95 ;
         LAYER m3 ;
         RECT  103.425 69.535 103.915 70.025 ;
         LAYER m3 ;
         RECT  95.815 77.065 96.305 77.555 ;
         LAYER m3 ;
         RECT  0.0 27.2 152.02 27.58 ;
         LAYER m3 ;
         RECT  57.12 91.12 96.94 91.5 ;
         LAYER m4 ;
         RECT  65.28 0.0 65.66 139.78 ;
         LAYER m4 ;
         RECT  131.92 0.0 132.3 139.78 ;
         LAYER m4 ;
         RECT  141.44 0.0 141.82 139.78 ;
         LAYER m3 ;
         RECT  49.845 87.195 50.335 87.685 ;
         LAYER m3 ;
         RECT  6.355 57.39 6.845 57.88 ;
         LAYER m3 ;
         RECT  9.52 99.28 73.14 99.66 ;
         LAYER m3 ;
         RECT  0.0 53.04 26.22 53.42 ;
         LAYER m4 ;
         RECT  70.72 0.0 71.1 139.78 ;
         LAYER m3 ;
         RECT  0.0 21.76 26.22 22.14 ;
         LAYER m3 ;
         RECT  103.36 72.08 142.5 72.46 ;
         LAYER m3 ;
         RECT  17.68 43.52 129.58 43.9 ;
         LAYER m3 ;
         RECT  38.775 63.495 39.265 63.985 ;
         LAYER m4 ;
         RECT  39.44 0.0 39.82 139.78 ;
         LAYER m4 ;
         RECT  6.8 0.0 7.18 139.78 ;
         LAYER m3 ;
         RECT  27.245 28.31 27.735 28.8 ;
         LAYER m3 ;
         RECT  99.405 71.36 99.895 71.85 ;
         LAYER m3 ;
         RECT  0.0 50.32 62.94 50.7 ;
         LAYER m3 ;
         RECT  84.89 66.57 85.19 66.87 ;
         LAYER m3 ;
         RECT  53.865 83.21 54.355 83.7 ;
         LAYER m4 ;
         RECT  76.16 0.0 76.54 139.78 ;
         LAYER m3 ;
         RECT  28.56 48.96 142.5 49.34 ;
         LAYER m4 ;
         RECT  95.2 0.0 95.58 139.78 ;
         LAYER m3 ;
         RECT  99.405 85.185 99.895 85.675 ;
         LAYER m3 ;
         RECT  27.245 14.17 27.735 14.66 ;
         LAYER m3 ;
         RECT  57.12 89.76 96.94 90.14 ;
         LAYER m4 ;
         RECT  137.36 0.0 137.74 139.78 ;
         LAYER m3 ;
         RECT  130.56 38.08 152.02 38.46 ;
         LAYER m3 ;
         RECT  84.89 94.22 85.19 94.52 ;
         LAYER m3 ;
         RECT  103.425 67.445 103.915 67.935 ;
         LAYER m4 ;
         RECT  55.76 0.0 56.14 139.78 ;
         LAYER m3 ;
         RECT  110.475 75.31 110.965 75.8 ;
         LAYER m3 ;
         RECT  57.12 74.8 96.94 75.18 ;
         LAYER m3 ;
         RECT  9.52 59.84 152.02 60.22 ;
         LAYER m3 ;
         RECT  57.12 70.72 96.94 71.1 ;
         LAYER m3 ;
         RECT  0.0 46.24 73.82 46.62 ;
         LAYER m3 ;
         RECT  0.0 29.92 73.82 30.3 ;
         LAYER m3 ;
         RECT  0.0 32.64 152.02 33.02 ;
         LAYER m3 ;
         RECT  127.84 42.16 152.02 42.54 ;
         LAYER m3 ;
         RECT  25.84 130.56 152.02 130.94 ;
         LAYER m3 ;
         RECT  68.57 93.035 68.87 93.335 ;
         LAYER m3 ;
         RECT  68.57 94.22 68.87 94.52 ;
         LAYER m3 ;
         RECT  84.89 87.9 85.19 88.2 ;
         LAYER m4 ;
         RECT  104.72 0.0 105.1 139.78 ;
         LAYER m4 ;
         RECT  82.96 0.0 83.34 139.78 ;
         LAYER m3 ;
         RECT  31.28 126.48 152.02 126.86 ;
         LAYER m3 ;
         RECT  68.57 62.62 68.87 62.92 ;
         LAYER m3 ;
         RECT  84.89 93.035 85.19 93.335 ;
         LAYER m4 ;
         RECT  72.08 0.0 72.46 139.78 ;
         LAYER m3 ;
         RECT  114.495 75.345 114.985 75.835 ;
         LAYER m4 ;
         RECT  47.6 0.0 47.98 139.78 ;
         LAYER m4 ;
         RECT  142.8 0.0 143.18 139.78 ;
         LAYER m4 ;
         RECT  136.0 0.0 136.38 139.78 ;
         LAYER m3 ;
         RECT  99.405 75.31 99.895 75.8 ;
         LAYER m3 ;
         RECT  0.0 78.88 39.82 79.26 ;
         LAYER m3 ;
         RECT  57.455 77.065 57.945 77.555 ;
         LAYER m4 ;
         RECT  38.08 0.0 38.46 139.78 ;
         LAYER m3 ;
         RECT  77.23 113.92 77.72 114.41 ;
         LAYER m3 ;
         RECT  145.805 96.89 146.295 97.38 ;
         LAYER m3 ;
         RECT  82.28 99.28 152.02 99.66 ;
         LAYER m4 ;
         RECT  43.52 0.0 43.9 139.78 ;
         LAYER m4 ;
         RECT  146.88 0.0 147.26 139.78 ;
         LAYER m3 ;
         RECT  84.89 81.185 85.19 81.485 ;
         LAYER m3 ;
         RECT  28.56 21.76 152.02 22.14 ;
         LAYER m3 ;
         RECT  32.925 63.46 33.415 63.95 ;
         LAYER m4 ;
         RECT  50.32 0.0 50.7 139.78 ;
         LAYER m3 ;
         RECT  0.0 118.32 124.82 118.7 ;
         LAYER m3 ;
         RECT  0.0 1.36 13.3 1.74 ;
         LAYER m3 ;
         RECT  49.845 81.385 50.335 81.875 ;
         LAYER m3 ;
         RECT  0.0 81.6 50.7 81.98 ;
         LAYER m3 ;
         RECT  82.96 58.48 144.54 58.86 ;
         LAYER m3 ;
         RECT  57.12 85.68 96.94 86.06 ;
         LAYER m3 ;
         RECT  53.865 91.11 54.355 91.6 ;
         LAYER m4 ;
         RECT  13.6 0.0 13.98 139.78 ;
         LAYER m3 ;
         RECT  120.345 75.31 120.835 75.8 ;
         LAYER m3 ;
         RECT  110.475 79.26 110.965 79.75 ;
         LAYER m3 ;
         RECT  128.945 17.41 129.435 17.9 ;
         LAYER m3 ;
         RECT  127.84 108.8 152.02 109.18 ;
         LAYER m3 ;
         RECT  84.89 74.47 85.19 74.77 ;
         LAYER m3 ;
         RECT  68.57 87.9 68.87 88.2 ;
         LAYER m3 ;
         RECT  38.775 79.295 39.265 79.785 ;
         LAYER m3 ;
         RECT  75.77 50.03 76.26 50.52 ;
         LAYER m3 ;
         RECT  57.12 72.08 96.94 72.46 ;
         LAYER m4 ;
         RECT  44.88 0.0 45.26 139.78 ;
         LAYER m3 ;
         RECT  128.52 119.68 152.02 120.06 ;
         LAYER m3 ;
         RECT  0.435 14.18 0.925 14.67 ;
         LAYER m3 ;
         RECT  0.0 122.4 131.62 122.78 ;
         LAYER m4 ;
         RECT  36.72 0.0 37.1 139.78 ;
         LAYER m3 ;
         RECT  128.52 133.28 150.66 133.66 ;
         LAYER m3 ;
         RECT  2.675 102.19 3.165 102.68 ;
         LAYER m4 ;
         RECT  62.56 0.0 62.94 139.78 ;
         LAYER m3 ;
         RECT  42.795 67.41 43.285 67.9 ;
         LAYER m3 ;
         RECT  42.84 0.0 152.02 0.38 ;
         LAYER m3 ;
         RECT  84.89 72.1 85.19 72.4 ;
         LAYER m3 ;
         RECT  76.88 50.03 77.37 50.52 ;
         LAYER m4 ;
         RECT  121.04 0.0 121.42 139.78 ;
         LAYER m3 ;
         RECT  49.845 91.145 50.335 91.635 ;
         LAYER m3 ;
         RECT  68.57 86.32 68.87 86.62 ;
         LAYER m3 ;
         RECT  103.36 81.6 152.02 81.98 ;
         LAYER m3 ;
         RECT  0.0 13.6 152.02 13.98 ;
         LAYER m3 ;
         RECT  25.84 1.36 152.02 1.74 ;
         LAYER m3 ;
         RECT  27.245 0.03 27.735 0.52 ;
         LAYER m4 ;
         RECT  92.48 0.0 92.86 139.78 ;
         LAYER m3 ;
         RECT  53.865 69.385 54.355 69.875 ;
         LAYER m3 ;
         RECT  103.425 83.245 103.915 83.735 ;
         LAYER m3 ;
         RECT  103.36 73.44 152.02 73.82 ;
         LAYER m3 ;
         RECT  0.0 112.88 73.82 113.26 ;
         LAYER m3 ;
         RECT  89.76 103.36 152.02 103.74 ;
         LAYER m4 ;
         RECT  103.36 0.0 103.74 139.78 ;
         LAYER m3 ;
         RECT  68.57 81.185 68.87 81.485 ;
         LAYER m3 ;
         RECT  0.0 44.88 124.82 45.26 ;
         LAYER m4 ;
         RECT  1.36 0.0 1.74 139.78 ;
         LAYER m3 ;
         RECT  114.24 68.0 152.02 68.38 ;
         LAYER m3 ;
         RECT  68.57 76.05 68.87 76.35 ;
         LAYER m3 ;
         RECT  126.445 125.97 126.935 126.46 ;
         LAYER m4 ;
         RECT  80.24 0.0 80.62 139.78 ;
         LAYER m3 ;
         RECT  0.0 97.92 152.02 98.3 ;
         LAYER m4 ;
         RECT  91.12 0.0 91.5 139.78 ;
         LAYER m3 ;
         RECT  103.425 77.435 103.915 77.925 ;
         LAYER m3 ;
         RECT  75.77 104.25 76.26 104.74 ;
         LAYER m3 ;
         RECT  68.57 89.085 68.87 89.385 ;
         LAYER m3 ;
         RECT  84.89 80.0 85.19 80.3 ;
         LAYER m4 ;
         RECT  32.64 0.0 33.02 139.78 ;
         LAYER m3 ;
         RECT  68.57 72.1 68.87 72.4 ;
         LAYER m3 ;
         RECT  49.845 73.485 50.335 73.975 ;
         LAYER m3 ;
         RECT  0.0 61.2 142.5 61.58 ;
         LAYER m3 ;
         RECT  38.775 75.345 39.265 75.835 ;
         LAYER m3 ;
         RECT  68.57 77.235 68.87 77.535 ;
         LAYER m3 ;
         RECT  103.36 70.72 152.02 71.1 ;
         LAYER m3 ;
         RECT  0.0 72.08 50.7 72.46 ;
         LAYER m3 ;
         RECT  0.0 130.56 23.5 130.94 ;
         LAYER m3 ;
         RECT  2.04 10.88 152.02 11.26 ;
         LAYER m3 ;
         RECT  84.89 86.32 85.19 86.62 ;
         LAYER m4 ;
         RECT  84.32 0.0 84.7 139.78 ;
         LAYER m4 ;
         RECT  8.16 0.0 8.54 139.78 ;
         LAYER m4 ;
         RECT  0.0 0.0 0.38 139.78 ;
         LAYER m3 ;
         RECT  0.0 89.76 50.7 90.14 ;
         LAYER m3 ;
         RECT  75.4 32.55 75.89 33.04 ;
         LAYER m4 ;
         RECT  16.32 4.76 16.7 139.78 ;
         LAYER m3 ;
         RECT  103.36 69.36 144.54 69.74 ;
         LAYER m3 ;
         RECT  121.04 74.8 152.02 75.18 ;
         LAYER m3 ;
         RECT  23.8 125.12 152.02 125.5 ;
         LAYER m3 ;
         RECT  120.345 63.46 120.835 63.95 ;
         LAYER m4 ;
         RECT  23.12 0.0 23.5 139.78 ;
         LAYER m3 ;
         RECT  53.865 87.16 54.355 87.65 ;
         LAYER m4 ;
         RECT  140.08 0.0 140.46 139.78 ;
         LAYER m3 ;
         RECT  46.92 14.96 152.02 15.34 ;
         LAYER m3 ;
         RECT  126.445 97.69 126.935 98.18 ;
         LAYER m3 ;
         RECT  84.89 82.37 85.19 82.67 ;
         LAYER m3 ;
         RECT  49.845 83.245 50.335 83.735 ;
         LAYER m4 ;
         RECT  9.52 0.0 9.9 139.78 ;
         LAYER m3 ;
         RECT  99.405 91.11 99.895 91.6 ;
         LAYER m4 ;
         RECT  97.92 0.0 98.3 139.78 ;
         LAYER m3 ;
         RECT  0.0 34.0 73.14 34.38 ;
         LAYER m3 ;
         RECT  24.745 122.73 25.235 123.22 ;
         LAYER m3 ;
         RECT  103.36 87.04 152.02 87.42 ;
         LAYER m3 ;
         RECT  0.0 102.0 72.46 102.38 ;
         LAYER m3 ;
         RECT  57.12 69.36 96.94 69.74 ;
         LAYER m3 ;
         RECT  42.795 79.26 43.285 79.75 ;
         LAYER m3 ;
         RECT  24.745 108.59 25.235 109.08 ;
         LAYER m3 ;
         RECT  68.57 68.15 68.87 68.45 ;
         LAYER m3 ;
         RECT  42.795 63.46 43.285 63.95 ;
         LAYER m3 ;
         RECT  2.675 79.79 3.165 80.28 ;
         LAYER m4 ;
         RECT  149.6 0.0 149.98 139.78 ;
         LAYER m3 ;
         RECT  68.57 74.47 68.87 74.77 ;
         LAYER m3 ;
         RECT  6.355 79.79 6.845 80.28 ;
         LAYER m3 ;
         RECT  9.52 88.4 142.5 88.78 ;
         LAYER m3 ;
         RECT  99.405 79.26 99.895 79.75 ;
         LAYER m3 ;
         RECT  30.6 119.68 124.82 120.06 ;
         LAYER m3 ;
         RECT  0.0 69.36 50.7 69.74 ;
         LAYER m3 ;
         RECT  84.89 83.95 85.19 84.25 ;
         LAYER m3 ;
         RECT  24.745 136.87 25.235 137.36 ;
         LAYER m4 ;
         RECT  102.0 0.0 102.38 139.78 ;
         LAYER m3 ;
         RECT  84.89 78.42 85.19 78.72 ;
         LAYER m3 ;
         RECT  49.845 69.535 50.335 70.025 ;
         LAYER m4 ;
         RECT  119.68 0.0 120.06 139.78 ;
         LAYER m4 ;
         RECT  77.52 0.0 77.9 139.78 ;
         LAYER m3 ;
         RECT  0.0 40.8 152.02 41.18 ;
         LAYER m3 ;
         RECT  0.0 12.24 9.9 12.62 ;
         LAYER m3 ;
         RECT  99.405 81.235 99.895 81.725 ;
         LAYER m3 ;
         RECT  149.485 52.09 149.975 52.58 ;
         LAYER m3 ;
         RECT  68.57 70.52 68.87 70.82 ;
         LAYER m3 ;
         RECT  7.48 96.56 152.02 96.94 ;
         LAYER m3 ;
         RECT  0.0 36.72 152.02 37.1 ;
         LAYER m3 ;
         RECT  77.23 40.36 77.72 40.85 ;
         LAYER m4 ;
         RECT  145.52 0.0 145.9 139.78 ;
         LAYER m3 ;
         RECT  103.36 85.68 152.02 86.06 ;
         LAYER m3 ;
         RECT  130.56 24.48 152.02 24.86 ;
         LAYER m3 ;
         RECT  9.52 104.72 124.82 105.1 ;
         LAYER m4 ;
         RECT  73.44 0.0 73.82 139.78 ;
         LAYER m3 ;
         RECT  57.12 68.0 96.94 68.38 ;
         LAYER m3 ;
         RECT  9.52 93.84 142.5 94.22 ;
         LAYER m4 ;
         RECT  134.64 0.0 135.02 139.78 ;
         LAYER m4 ;
         RECT  125.12 0.0 125.5 139.78 ;
         LAYER m3 ;
         RECT  0.0 8.16 11.26 8.54 ;
         LAYER m4 ;
         RECT  21.76 0.0 22.14 139.78 ;
         LAYER m4 ;
         RECT  89.76 0.0 90.14 139.78 ;
         LAYER m3 ;
         RECT  103.425 71.395 103.915 71.885 ;
         LAYER m3 ;
         RECT  81.6 50.32 152.02 50.7 ;
         LAYER m3 ;
         RECT  103.425 85.335 103.915 85.825 ;
         LAYER m3 ;
         RECT  44.2 20.4 122.1 20.78 ;
         LAYER m4 ;
         RECT  14.96 0.0 15.34 139.78 ;
         LAYER m3 ;
         RECT  68.57 83.95 68.87 84.25 ;
         LAYER m3 ;
         RECT  145.805 85.69 146.295 86.18 ;
         LAYER m3 ;
         RECT  0.0 5.44 152.02 5.82 ;
         LAYER m4 ;
         RECT  54.4 0.0 54.78 139.78 ;
         LAYER m3 ;
         RECT  0.0 39.44 26.22 39.82 ;
         LAYER m3 ;
         RECT  114.495 79.295 114.985 79.785 ;
         LAYER m3 ;
         RECT  99.405 89.135 99.895 89.625 ;
         LAYER m3 ;
         RECT  84.89 85.135 85.19 85.435 ;
         LAYER m3 ;
         RECT  110.475 63.46 110.965 63.95 ;
         LAYER m3 ;
         RECT  0.0 23.12 152.02 23.5 ;
         LAYER m3 ;
         RECT  68.57 85.135 68.87 85.435 ;
         LAYER m3 ;
         RECT  57.12 73.44 96.94 73.82 ;
         LAYER m4 ;
         RECT  2.72 0.0 3.1 139.78 ;
         LAYER m4 ;
         RECT  66.64 0.0 67.02 139.78 ;
         LAYER m3 ;
         RECT  61.665 77.14 62.155 77.63 ;
         LAYER m3 ;
         RECT  0.435 0.02 0.925 0.51 ;
         LAYER m4 ;
         RECT  112.88 0.0 113.26 139.78 ;
         LAYER m3 ;
         RECT  0.0 126.48 26.22 126.86 ;
         LAYER m3 ;
         RECT  75.42 40.36 75.91 40.85 ;
         LAYER m3 ;
         RECT  0.0 51.68 7.86 52.06 ;
         LAYER m4 ;
         RECT  93.84 0.0 94.22 139.78 ;
         LAYER m3 ;
         RECT  103.36 91.12 144.54 91.5 ;
         LAYER m3 ;
         RECT  31.28 133.28 124.82 133.66 ;
         LAYER m3 ;
         RECT  0.0 17.68 11.94 18.06 ;
         LAYER m3 ;
         RECT  149.485 63.29 149.975 63.78 ;
         LAYER m3 ;
         RECT  127.84 44.88 152.02 45.26 ;
         LAYER m3 ;
         RECT  103.36 89.76 152.02 90.14 ;
         LAYER m3 ;
         RECT  0.0 129.2 23.5 129.58 ;
         LAYER m3 ;
         RECT  0.0 65.28 50.7 65.66 ;
         LAYER m3 ;
         RECT  68.57 90.27 68.87 90.57 ;
         LAYER m3 ;
         RECT  68.57 66.57 68.87 66.87 ;
         LAYER m3 ;
         RECT  68.57 69.335 68.87 69.635 ;
         LAYER m3 ;
         RECT  68.57 78.42 68.87 78.72 ;
         LAYER m3 ;
         RECT  99.405 67.41 99.895 67.9 ;
         LAYER m4 ;
         RECT  12.24 0.0 12.62 139.78 ;
         LAYER m3 ;
         RECT  7.48 107.44 73.82 107.82 ;
         LAYER m4 ;
         RECT  48.96 0.0 49.34 139.78 ;
         LAYER m3 ;
         RECT  75.42 113.92 75.91 114.41 ;
         LAYER m3 ;
         RECT  0.0 63.92 33.02 64.3 ;
         LAYER m3 ;
         RECT  0.0 123.76 152.02 124.14 ;
         LAYER m3 ;
         RECT  49.845 77.435 50.335 77.925 ;
         LAYER m3 ;
         RECT  79.56 29.92 152.02 30.3 ;
         LAYER m3 ;
         RECT  0.0 100.64 86.74 101.02 ;
         LAYER m3 ;
         RECT  0.0 114.24 72.46 114.62 ;
         LAYER m3 ;
         RECT  68.57 73.285 68.87 73.585 ;
         LAYER m3 ;
         RECT  103.425 89.285 103.915 89.775 ;
         LAYER m3 ;
         RECT  32.925 75.31 33.415 75.8 ;
         LAYER m3 ;
         RECT  76.88 104.25 77.37 104.74 ;
         LAYER m3 ;
         RECT  0.0 47.6 152.02 47.98 ;
         LAYER m3 ;
         RECT  1.36 6.8 26.22 7.18 ;
         LAYER m3 ;
         RECT  91.605 77.14 92.095 77.63 ;
         LAYER m4 ;
         RECT  150.96 0.0 151.34 139.78 ;
         LAYER m3 ;
         RECT  0.0 133.28 26.22 133.66 ;
         LAYER m4 ;
         RECT  53.04 0.0 53.42 139.78 ;
         LAYER m3 ;
         RECT  0.0 0.0 33.7 0.38 ;
         LAYER m4 ;
         RECT  20.4 0.0 20.78 139.78 ;
         LAYER m4 ;
         RECT  24.48 0.0 24.86 139.78 ;
         LAYER m4 ;
         RECT  51.68 0.0 52.06 139.78 ;
         LAYER m4 ;
         RECT  58.48 0.0 58.86 139.78 ;
         LAYER m3 ;
         RECT  0.0 24.48 26.22 24.86 ;
         LAYER m3 ;
         RECT  78.88 46.24 144.54 46.62 ;
         LAYER m3 ;
         RECT  0.0 80.24 144.54 80.62 ;
         LAYER m3 ;
         RECT  0.0 103.36 72.46 103.74 ;
         LAYER m4 ;
         RECT  87.04 0.0 87.42 139.78 ;
         LAYER m3 ;
         RECT  9.52 82.96 50.7 83.34 ;
         LAYER m4 ;
         RECT  17.68 0.0 18.06 139.78 ;
         LAYER m3 ;
         RECT  81.6 53.04 152.02 53.42 ;
         LAYER m3 ;
         RECT  57.12 63.92 96.94 64.3 ;
         LAYER m3 ;
         RECT  128.52 104.72 152.02 105.1 ;
         LAYER m3 ;
         RECT  0.0 92.48 152.02 92.86 ;
         LAYER m3 ;
         RECT  2.04 2.72 152.02 3.1 ;
         LAYER m3 ;
         RECT  49.845 67.445 50.335 67.935 ;
         LAYER m3 ;
         RECT  0.0 20.4 35.06 20.78 ;
         LAYER m4 ;
         RECT  118.32 0.0 118.7 139.78 ;
         LAYER m3 ;
         RECT  68.57 65.385 68.87 65.685 ;
         LAYER m3 ;
         RECT  0.0 131.92 129.58 132.3 ;
         LAYER m4 ;
         RECT  127.84 0.0 128.22 139.78 ;
         LAYER m3 ;
         RECT  36.425 12.895 36.915 13.385 ;
         LAYER m3 ;
         RECT  141.44 131.92 152.02 132.3 ;
         LAYER m3 ;
         RECT  99.405 65.435 99.895 65.925 ;
         LAYER m3 ;
         RECT  0.0 25.84 152.02 26.22 ;
      END
   END gnd
   OBS
   LAYER  m1 ;
      RECT  76.595 61.98 76.67 63.685 ;
      RECT  76.67 61.395 76.88 61.775 ;
      RECT  74.51 61.065 74.69 61.98 ;
      POLYGON  76.16 62.07 76.16 62.48 76.335 62.48 76.415 62.4 76.415 62.07 76.16 62.07 ;
      RECT  74.15 61.98 74.33 63.685 ;
      RECT  74.51 61.98 74.69 63.685 ;
      RECT  73.76 61.98 73.97 63.685 ;
      RECT  73.55 61.775 73.76 61.98 ;
      RECT  73.55 61.98 73.76 63.685 ;
      RECT  76.67 61.98 76.88 63.685 ;
      POLYGON  76.16 63.06 76.16 63.47 76.415 63.47 76.415 63.14 76.335 63.06 76.16 63.06 ;
      RECT  73.76 61.395 73.97 61.775 ;
      RECT  76.67 61.065 76.88 61.395 ;
      RECT  74.87 61.065 75.05 61.98 ;
      RECT  76.51 62.565 76.595 62.975 ;
      RECT  75.59 61.98 75.77 63.685 ;
      RECT  75.95 63.06 76.16 63.47 ;
      RECT  73.76 61.065 73.97 61.395 ;
      RECT  75.95 62.07 76.16 62.48 ;
      RECT  75.95 61.395 76.16 61.775 ;
      RECT  73.55 61.395 73.76 61.775 ;
      RECT  75.23 61.065 75.41 61.98 ;
      RECT  75.23 61.98 75.41 63.685 ;
      RECT  76.67 61.775 76.88 61.98 ;
      RECT  73.76 61.775 73.97 61.98 ;
      RECT  73.55 61.065 73.76 61.395 ;
      RECT  75.59 61.065 75.77 61.98 ;
      RECT  74.15 61.065 74.33 61.98 ;
      POLYGON  76.595 61.065 76.595 61.395 76.16 61.395 76.16 61.775 76.595 61.775 76.595 61.98 76.67 61.98 76.67 61.065 76.595 61.065 ;
      RECT  74.87 61.98 75.05 63.685 ;
      RECT  76.595 65.14 76.67 63.435 ;
      RECT  76.67 65.725 76.88 65.345 ;
      RECT  74.51 66.055 74.69 65.14 ;
      POLYGON  76.16 65.05 76.16 64.64 76.335 64.64 76.415 64.72 76.415 65.05 76.16 65.05 ;
      RECT  74.15 65.14 74.33 63.435 ;
      RECT  74.51 65.14 74.69 63.435 ;
      RECT  73.76 65.14 73.97 63.435 ;
      RECT  73.55 65.345 73.76 65.14 ;
      RECT  73.55 65.14 73.76 63.435 ;
      RECT  76.67 65.14 76.88 63.435 ;
      POLYGON  76.16 64.06 76.16 63.65 76.415 63.65 76.415 63.98 76.335 64.06 76.16 64.06 ;
      RECT  73.76 65.725 73.97 65.345 ;
      RECT  76.67 66.055 76.88 65.725 ;
      RECT  74.87 66.055 75.05 65.14 ;
      RECT  76.51 64.555 76.595 64.145 ;
      RECT  75.59 65.14 75.77 63.435 ;
      RECT  75.95 64.06 76.16 63.65 ;
      RECT  73.76 66.055 73.97 65.725 ;
      RECT  75.95 65.05 76.16 64.64 ;
      RECT  75.95 65.725 76.16 65.345 ;
      RECT  73.55 65.725 73.76 65.345 ;
      RECT  75.23 66.055 75.41 65.14 ;
      RECT  75.23 65.14 75.41 63.435 ;
      RECT  76.67 65.345 76.88 65.14 ;
      RECT  73.76 65.345 73.97 65.14 ;
      RECT  73.55 66.055 73.76 65.725 ;
      RECT  75.59 66.055 75.77 65.14 ;
      RECT  74.15 66.055 74.33 65.14 ;
      POLYGON  76.595 66.055 76.595 65.725 76.16 65.725 76.16 65.345 76.595 65.345 76.595 65.14 76.67 65.14 76.67 66.055 76.595 66.055 ;
      RECT  74.87 65.14 75.05 63.435 ;
      RECT  76.595 65.93 76.67 67.635 ;
      RECT  76.67 65.345 76.88 65.725 ;
      RECT  74.51 65.015 74.69 65.93 ;
      POLYGON  76.16 66.02 76.16 66.43 76.335 66.43 76.415 66.35 76.415 66.02 76.16 66.02 ;
      RECT  74.15 65.93 74.33 67.635 ;
      RECT  74.51 65.93 74.69 67.635 ;
      RECT  73.76 65.93 73.97 67.635 ;
      RECT  73.55 65.725 73.76 65.93 ;
      RECT  73.55 65.93 73.76 67.635 ;
      RECT  76.67 65.93 76.88 67.635 ;
      POLYGON  76.16 67.01 76.16 67.42 76.415 67.42 76.415 67.09 76.335 67.01 76.16 67.01 ;
      RECT  73.76 65.345 73.97 65.725 ;
      RECT  76.67 65.015 76.88 65.345 ;
      RECT  74.87 65.015 75.05 65.93 ;
      RECT  76.51 66.515 76.595 66.925 ;
      RECT  75.59 65.93 75.77 67.635 ;
      RECT  75.95 67.01 76.16 67.42 ;
      RECT  73.76 65.015 73.97 65.345 ;
      RECT  75.95 66.02 76.16 66.43 ;
      RECT  75.95 65.345 76.16 65.725 ;
      RECT  73.55 65.345 73.76 65.725 ;
      RECT  75.23 65.015 75.41 65.93 ;
      RECT  75.23 65.93 75.41 67.635 ;
      RECT  76.67 65.725 76.88 65.93 ;
      RECT  73.76 65.725 73.97 65.93 ;
      RECT  73.55 65.015 73.76 65.345 ;
      RECT  75.59 65.015 75.77 65.93 ;
      RECT  74.15 65.015 74.33 65.93 ;
      POLYGON  76.595 65.015 76.595 65.345 76.16 65.345 76.16 65.725 76.595 65.725 76.595 65.93 76.67 65.93 76.67 65.015 76.595 65.015 ;
      RECT  74.87 65.93 75.05 67.635 ;
      RECT  76.595 69.09 76.67 67.385 ;
      RECT  76.67 69.675 76.88 69.295 ;
      RECT  74.51 70.005 74.69 69.09 ;
      POLYGON  76.16 69.0 76.16 68.59 76.335 68.59 76.415 68.67 76.415 69.0 76.16 69.0 ;
      RECT  74.15 69.09 74.33 67.385 ;
      RECT  74.51 69.09 74.69 67.385 ;
      RECT  73.76 69.09 73.97 67.385 ;
      RECT  73.55 69.295 73.76 69.09 ;
      RECT  73.55 69.09 73.76 67.385 ;
      RECT  76.67 69.09 76.88 67.385 ;
      POLYGON  76.16 68.01 76.16 67.6 76.415 67.6 76.415 67.93 76.335 68.01 76.16 68.01 ;
      RECT  73.76 69.675 73.97 69.295 ;
      RECT  76.67 70.005 76.88 69.675 ;
      RECT  74.87 70.005 75.05 69.09 ;
      RECT  76.51 68.505 76.595 68.095 ;
      RECT  75.59 69.09 75.77 67.385 ;
      RECT  75.95 68.01 76.16 67.6 ;
      RECT  73.76 70.005 73.97 69.675 ;
      RECT  75.95 69.0 76.16 68.59 ;
      RECT  75.95 69.675 76.16 69.295 ;
      RECT  73.55 69.675 73.76 69.295 ;
      RECT  75.23 70.005 75.41 69.09 ;
      RECT  75.23 69.09 75.41 67.385 ;
      RECT  76.67 69.295 76.88 69.09 ;
      RECT  73.76 69.295 73.97 69.09 ;
      RECT  73.55 70.005 73.76 69.675 ;
      RECT  75.59 70.005 75.77 69.09 ;
      RECT  74.15 70.005 74.33 69.09 ;
      POLYGON  76.595 70.005 76.595 69.675 76.16 69.675 76.16 69.295 76.595 69.295 76.595 69.09 76.67 69.09 76.67 70.005 76.595 70.005 ;
      RECT  74.87 69.09 75.05 67.385 ;
      RECT  76.595 69.88 76.67 71.585 ;
      RECT  76.67 69.295 76.88 69.675 ;
      RECT  74.51 68.965 74.69 69.88 ;
      POLYGON  76.16 69.97 76.16 70.38 76.335 70.38 76.415 70.3 76.415 69.97 76.16 69.97 ;
      RECT  74.15 69.88 74.33 71.585 ;
      RECT  74.51 69.88 74.69 71.585 ;
      RECT  73.76 69.88 73.97 71.585 ;
      RECT  73.55 69.675 73.76 69.88 ;
      RECT  73.55 69.88 73.76 71.585 ;
      RECT  76.67 69.88 76.88 71.585 ;
      POLYGON  76.16 70.96 76.16 71.37 76.415 71.37 76.415 71.04 76.335 70.96 76.16 70.96 ;
      RECT  73.76 69.295 73.97 69.675 ;
      RECT  76.67 68.965 76.88 69.295 ;
      RECT  74.87 68.965 75.05 69.88 ;
      RECT  76.51 70.465 76.595 70.875 ;
      RECT  75.59 69.88 75.77 71.585 ;
      RECT  75.95 70.96 76.16 71.37 ;
      RECT  73.76 68.965 73.97 69.295 ;
      RECT  75.95 69.97 76.16 70.38 ;
      RECT  75.95 69.295 76.16 69.675 ;
      RECT  73.55 69.295 73.76 69.675 ;
      RECT  75.23 68.965 75.41 69.88 ;
      RECT  75.23 69.88 75.41 71.585 ;
      RECT  76.67 69.675 76.88 69.88 ;
      RECT  73.76 69.675 73.97 69.88 ;
      RECT  73.55 68.965 73.76 69.295 ;
      RECT  75.59 68.965 75.77 69.88 ;
      RECT  74.15 68.965 74.33 69.88 ;
      POLYGON  76.595 68.965 76.595 69.295 76.16 69.295 76.16 69.675 76.595 69.675 76.595 69.88 76.67 69.88 76.67 68.965 76.595 68.965 ;
      RECT  74.87 69.88 75.05 71.585 ;
      RECT  76.595 73.04 76.67 71.335 ;
      RECT  76.67 73.625 76.88 73.245 ;
      RECT  74.51 73.955 74.69 73.04 ;
      POLYGON  76.16 72.95 76.16 72.54 76.335 72.54 76.415 72.62 76.415 72.95 76.16 72.95 ;
      RECT  74.15 73.04 74.33 71.335 ;
      RECT  74.51 73.04 74.69 71.335 ;
      RECT  73.76 73.04 73.97 71.335 ;
      RECT  73.55 73.245 73.76 73.04 ;
      RECT  73.55 73.04 73.76 71.335 ;
      RECT  76.67 73.04 76.88 71.335 ;
      POLYGON  76.16 71.96 76.16 71.55 76.415 71.55 76.415 71.88 76.335 71.96 76.16 71.96 ;
      RECT  73.76 73.625 73.97 73.245 ;
      RECT  76.67 73.955 76.88 73.625 ;
      RECT  74.87 73.955 75.05 73.04 ;
      RECT  76.51 72.455 76.595 72.045 ;
      RECT  75.59 73.04 75.77 71.335 ;
      RECT  75.95 71.96 76.16 71.55 ;
      RECT  73.76 73.955 73.97 73.625 ;
      RECT  75.95 72.95 76.16 72.54 ;
      RECT  75.95 73.625 76.16 73.245 ;
      RECT  73.55 73.625 73.76 73.245 ;
      RECT  75.23 73.955 75.41 73.04 ;
      RECT  75.23 73.04 75.41 71.335 ;
      RECT  76.67 73.245 76.88 73.04 ;
      RECT  73.76 73.245 73.97 73.04 ;
      RECT  73.55 73.955 73.76 73.625 ;
      RECT  75.59 73.955 75.77 73.04 ;
      RECT  74.15 73.955 74.33 73.04 ;
      POLYGON  76.595 73.955 76.595 73.625 76.16 73.625 76.16 73.245 76.595 73.245 76.595 73.04 76.67 73.04 76.67 73.955 76.595 73.955 ;
      RECT  74.87 73.04 75.05 71.335 ;
      RECT  76.595 73.83 76.67 75.535 ;
      RECT  76.67 73.245 76.88 73.625 ;
      RECT  74.51 72.915 74.69 73.83 ;
      POLYGON  76.16 73.92 76.16 74.33 76.335 74.33 76.415 74.25 76.415 73.92 76.16 73.92 ;
      RECT  74.15 73.83 74.33 75.535 ;
      RECT  74.51 73.83 74.69 75.535 ;
      RECT  73.76 73.83 73.97 75.535 ;
      RECT  73.55 73.625 73.76 73.83 ;
      RECT  73.55 73.83 73.76 75.535 ;
      RECT  76.67 73.83 76.88 75.535 ;
      POLYGON  76.16 74.91 76.16 75.32 76.415 75.32 76.415 74.99 76.335 74.91 76.16 74.91 ;
      RECT  73.76 73.245 73.97 73.625 ;
      RECT  76.67 72.915 76.88 73.245 ;
      RECT  74.87 72.915 75.05 73.83 ;
      RECT  76.51 74.415 76.595 74.825 ;
      RECT  75.59 73.83 75.77 75.535 ;
      RECT  75.95 74.91 76.16 75.32 ;
      RECT  73.76 72.915 73.97 73.245 ;
      RECT  75.95 73.92 76.16 74.33 ;
      RECT  75.95 73.245 76.16 73.625 ;
      RECT  73.55 73.245 73.76 73.625 ;
      RECT  75.23 72.915 75.41 73.83 ;
      RECT  75.23 73.83 75.41 75.535 ;
      RECT  76.67 73.625 76.88 73.83 ;
      RECT  73.76 73.625 73.97 73.83 ;
      RECT  73.55 72.915 73.76 73.245 ;
      RECT  75.59 72.915 75.77 73.83 ;
      RECT  74.15 72.915 74.33 73.83 ;
      POLYGON  76.595 72.915 76.595 73.245 76.16 73.245 76.16 73.625 76.595 73.625 76.595 73.83 76.67 73.83 76.67 72.915 76.595 72.915 ;
      RECT  74.87 73.83 75.05 75.535 ;
      RECT  76.595 76.99 76.67 75.285 ;
      RECT  76.67 77.575 76.88 77.195 ;
      RECT  74.51 77.905 74.69 76.99 ;
      POLYGON  76.16 76.9 76.16 76.49 76.335 76.49 76.415 76.57 76.415 76.9 76.16 76.9 ;
      RECT  74.15 76.99 74.33 75.285 ;
      RECT  74.51 76.99 74.69 75.285 ;
      RECT  73.76 76.99 73.97 75.285 ;
      RECT  73.55 77.195 73.76 76.99 ;
      RECT  73.55 76.99 73.76 75.285 ;
      RECT  76.67 76.99 76.88 75.285 ;
      POLYGON  76.16 75.91 76.16 75.5 76.415 75.5 76.415 75.83 76.335 75.91 76.16 75.91 ;
      RECT  73.76 77.575 73.97 77.195 ;
      RECT  76.67 77.905 76.88 77.575 ;
      RECT  74.87 77.905 75.05 76.99 ;
      RECT  76.51 76.405 76.595 75.995 ;
      RECT  75.59 76.99 75.77 75.285 ;
      RECT  75.95 75.91 76.16 75.5 ;
      RECT  73.76 77.905 73.97 77.575 ;
      RECT  75.95 76.9 76.16 76.49 ;
      RECT  75.95 77.575 76.16 77.195 ;
      RECT  73.55 77.575 73.76 77.195 ;
      RECT  75.23 77.905 75.41 76.99 ;
      RECT  75.23 76.99 75.41 75.285 ;
      RECT  76.67 77.195 76.88 76.99 ;
      RECT  73.76 77.195 73.97 76.99 ;
      RECT  73.55 77.905 73.76 77.575 ;
      RECT  75.59 77.905 75.77 76.99 ;
      RECT  74.15 77.905 74.33 76.99 ;
      POLYGON  76.595 77.905 76.595 77.575 76.16 77.575 76.16 77.195 76.595 77.195 76.595 76.99 76.67 76.99 76.67 77.905 76.595 77.905 ;
      RECT  74.87 76.99 75.05 75.285 ;
      RECT  76.595 77.78 76.67 79.485 ;
      RECT  76.67 77.195 76.88 77.575 ;
      RECT  74.51 76.865 74.69 77.78 ;
      POLYGON  76.16 77.87 76.16 78.28 76.335 78.28 76.415 78.2 76.415 77.87 76.16 77.87 ;
      RECT  74.15 77.78 74.33 79.485 ;
      RECT  74.51 77.78 74.69 79.485 ;
      RECT  73.76 77.78 73.97 79.485 ;
      RECT  73.55 77.575 73.76 77.78 ;
      RECT  73.55 77.78 73.76 79.485 ;
      RECT  76.67 77.78 76.88 79.485 ;
      POLYGON  76.16 78.86 76.16 79.27 76.415 79.27 76.415 78.94 76.335 78.86 76.16 78.86 ;
      RECT  73.76 77.195 73.97 77.575 ;
      RECT  76.67 76.865 76.88 77.195 ;
      RECT  74.87 76.865 75.05 77.78 ;
      RECT  76.51 78.365 76.595 78.775 ;
      RECT  75.59 77.78 75.77 79.485 ;
      RECT  75.95 78.86 76.16 79.27 ;
      RECT  73.76 76.865 73.97 77.195 ;
      RECT  75.95 77.87 76.16 78.28 ;
      RECT  75.95 77.195 76.16 77.575 ;
      RECT  73.55 77.195 73.76 77.575 ;
      RECT  75.23 76.865 75.41 77.78 ;
      RECT  75.23 77.78 75.41 79.485 ;
      RECT  76.67 77.575 76.88 77.78 ;
      RECT  73.76 77.575 73.97 77.78 ;
      RECT  73.55 76.865 73.76 77.195 ;
      RECT  75.59 76.865 75.77 77.78 ;
      RECT  74.15 76.865 74.33 77.78 ;
      POLYGON  76.595 76.865 76.595 77.195 76.16 77.195 76.16 77.575 76.595 77.575 76.595 77.78 76.67 77.78 76.67 76.865 76.595 76.865 ;
      RECT  74.87 77.78 75.05 79.485 ;
      RECT  76.595 80.94 76.67 79.235 ;
      RECT  76.67 81.525 76.88 81.145 ;
      RECT  74.51 81.855 74.69 80.94 ;
      POLYGON  76.16 80.85 76.16 80.44 76.335 80.44 76.415 80.52 76.415 80.85 76.16 80.85 ;
      RECT  74.15 80.94 74.33 79.235 ;
      RECT  74.51 80.94 74.69 79.235 ;
      RECT  73.76 80.94 73.97 79.235 ;
      RECT  73.55 81.145 73.76 80.94 ;
      RECT  73.55 80.94 73.76 79.235 ;
      RECT  76.67 80.94 76.88 79.235 ;
      POLYGON  76.16 79.86 76.16 79.45 76.415 79.45 76.415 79.78 76.335 79.86 76.16 79.86 ;
      RECT  73.76 81.525 73.97 81.145 ;
      RECT  76.67 81.855 76.88 81.525 ;
      RECT  74.87 81.855 75.05 80.94 ;
      RECT  76.51 80.355 76.595 79.945 ;
      RECT  75.59 80.94 75.77 79.235 ;
      RECT  75.95 79.86 76.16 79.45 ;
      RECT  73.76 81.855 73.97 81.525 ;
      RECT  75.95 80.85 76.16 80.44 ;
      RECT  75.95 81.525 76.16 81.145 ;
      RECT  73.55 81.525 73.76 81.145 ;
      RECT  75.23 81.855 75.41 80.94 ;
      RECT  75.23 80.94 75.41 79.235 ;
      RECT  76.67 81.145 76.88 80.94 ;
      RECT  73.76 81.145 73.97 80.94 ;
      RECT  73.55 81.855 73.76 81.525 ;
      RECT  75.59 81.855 75.77 80.94 ;
      RECT  74.15 81.855 74.33 80.94 ;
      POLYGON  76.595 81.855 76.595 81.525 76.16 81.525 76.16 81.145 76.595 81.145 76.595 80.94 76.67 80.94 76.67 81.855 76.595 81.855 ;
      RECT  74.87 80.94 75.05 79.235 ;
      RECT  76.595 81.73 76.67 83.435 ;
      RECT  76.67 81.145 76.88 81.525 ;
      RECT  74.51 80.815 74.69 81.73 ;
      POLYGON  76.16 81.82 76.16 82.23 76.335 82.23 76.415 82.15 76.415 81.82 76.16 81.82 ;
      RECT  74.15 81.73 74.33 83.435 ;
      RECT  74.51 81.73 74.69 83.435 ;
      RECT  73.76 81.73 73.97 83.435 ;
      RECT  73.55 81.525 73.76 81.73 ;
      RECT  73.55 81.73 73.76 83.435 ;
      RECT  76.67 81.73 76.88 83.435 ;
      POLYGON  76.16 82.81 76.16 83.22 76.415 83.22 76.415 82.89 76.335 82.81 76.16 82.81 ;
      RECT  73.76 81.145 73.97 81.525 ;
      RECT  76.67 80.815 76.88 81.145 ;
      RECT  74.87 80.815 75.05 81.73 ;
      RECT  76.51 82.315 76.595 82.725 ;
      RECT  75.59 81.73 75.77 83.435 ;
      RECT  75.95 82.81 76.16 83.22 ;
      RECT  73.76 80.815 73.97 81.145 ;
      RECT  75.95 81.82 76.16 82.23 ;
      RECT  75.95 81.145 76.16 81.525 ;
      RECT  73.55 81.145 73.76 81.525 ;
      RECT  75.23 80.815 75.41 81.73 ;
      RECT  75.23 81.73 75.41 83.435 ;
      RECT  76.67 81.525 76.88 81.73 ;
      RECT  73.76 81.525 73.97 81.73 ;
      RECT  73.55 80.815 73.76 81.145 ;
      RECT  75.59 80.815 75.77 81.73 ;
      RECT  74.15 80.815 74.33 81.73 ;
      POLYGON  76.595 80.815 76.595 81.145 76.16 81.145 76.16 81.525 76.595 81.525 76.595 81.73 76.67 81.73 76.67 80.815 76.595 80.815 ;
      RECT  74.87 81.73 75.05 83.435 ;
      RECT  76.595 84.89 76.67 83.185 ;
      RECT  76.67 85.475 76.88 85.095 ;
      RECT  74.51 85.805 74.69 84.89 ;
      POLYGON  76.16 84.8 76.16 84.39 76.335 84.39 76.415 84.47 76.415 84.8 76.16 84.8 ;
      RECT  74.15 84.89 74.33 83.185 ;
      RECT  74.51 84.89 74.69 83.185 ;
      RECT  73.76 84.89 73.97 83.185 ;
      RECT  73.55 85.095 73.76 84.89 ;
      RECT  73.55 84.89 73.76 83.185 ;
      RECT  76.67 84.89 76.88 83.185 ;
      POLYGON  76.16 83.81 76.16 83.4 76.415 83.4 76.415 83.73 76.335 83.81 76.16 83.81 ;
      RECT  73.76 85.475 73.97 85.095 ;
      RECT  76.67 85.805 76.88 85.475 ;
      RECT  74.87 85.805 75.05 84.89 ;
      RECT  76.51 84.305 76.595 83.895 ;
      RECT  75.59 84.89 75.77 83.185 ;
      RECT  75.95 83.81 76.16 83.4 ;
      RECT  73.76 85.805 73.97 85.475 ;
      RECT  75.95 84.8 76.16 84.39 ;
      RECT  75.95 85.475 76.16 85.095 ;
      RECT  73.55 85.475 73.76 85.095 ;
      RECT  75.23 85.805 75.41 84.89 ;
      RECT  75.23 84.89 75.41 83.185 ;
      RECT  76.67 85.095 76.88 84.89 ;
      RECT  73.76 85.095 73.97 84.89 ;
      RECT  73.55 85.805 73.76 85.475 ;
      RECT  75.59 85.805 75.77 84.89 ;
      RECT  74.15 85.805 74.33 84.89 ;
      POLYGON  76.595 85.805 76.595 85.475 76.16 85.475 76.16 85.095 76.595 85.095 76.595 84.89 76.67 84.89 76.67 85.805 76.595 85.805 ;
      RECT  74.87 84.89 75.05 83.185 ;
      RECT  76.595 85.68 76.67 87.385 ;
      RECT  76.67 85.095 76.88 85.475 ;
      RECT  74.51 84.765 74.69 85.68 ;
      POLYGON  76.16 85.77 76.16 86.18 76.335 86.18 76.415 86.1 76.415 85.77 76.16 85.77 ;
      RECT  74.15 85.68 74.33 87.385 ;
      RECT  74.51 85.68 74.69 87.385 ;
      RECT  73.76 85.68 73.97 87.385 ;
      RECT  73.55 85.475 73.76 85.68 ;
      RECT  73.55 85.68 73.76 87.385 ;
      RECT  76.67 85.68 76.88 87.385 ;
      POLYGON  76.16 86.76 76.16 87.17 76.415 87.17 76.415 86.84 76.335 86.76 76.16 86.76 ;
      RECT  73.76 85.095 73.97 85.475 ;
      RECT  76.67 84.765 76.88 85.095 ;
      RECT  74.87 84.765 75.05 85.68 ;
      RECT  76.51 86.265 76.595 86.675 ;
      RECT  75.59 85.68 75.77 87.385 ;
      RECT  75.95 86.76 76.16 87.17 ;
      RECT  73.76 84.765 73.97 85.095 ;
      RECT  75.95 85.77 76.16 86.18 ;
      RECT  75.95 85.095 76.16 85.475 ;
      RECT  73.55 85.095 73.76 85.475 ;
      RECT  75.23 84.765 75.41 85.68 ;
      RECT  75.23 85.68 75.41 87.385 ;
      RECT  76.67 85.475 76.88 85.68 ;
      RECT  73.76 85.475 73.97 85.68 ;
      RECT  73.55 84.765 73.76 85.095 ;
      RECT  75.59 84.765 75.77 85.68 ;
      RECT  74.15 84.765 74.33 85.68 ;
      POLYGON  76.595 84.765 76.595 85.095 76.16 85.095 76.16 85.475 76.595 85.475 76.595 85.68 76.67 85.68 76.67 84.765 76.595 84.765 ;
      RECT  74.87 85.68 75.05 87.385 ;
      RECT  76.595 88.84 76.67 87.135 ;
      RECT  76.67 89.425 76.88 89.045 ;
      RECT  74.51 89.755 74.69 88.84 ;
      POLYGON  76.16 88.75 76.16 88.34 76.335 88.34 76.415 88.42 76.415 88.75 76.16 88.75 ;
      RECT  74.15 88.84 74.33 87.135 ;
      RECT  74.51 88.84 74.69 87.135 ;
      RECT  73.76 88.84 73.97 87.135 ;
      RECT  73.55 89.045 73.76 88.84 ;
      RECT  73.55 88.84 73.76 87.135 ;
      RECT  76.67 88.84 76.88 87.135 ;
      POLYGON  76.16 87.76 76.16 87.35 76.415 87.35 76.415 87.68 76.335 87.76 76.16 87.76 ;
      RECT  73.76 89.425 73.97 89.045 ;
      RECT  76.67 89.755 76.88 89.425 ;
      RECT  74.87 89.755 75.05 88.84 ;
      RECT  76.51 88.255 76.595 87.845 ;
      RECT  75.59 88.84 75.77 87.135 ;
      RECT  75.95 87.76 76.16 87.35 ;
      RECT  73.76 89.755 73.97 89.425 ;
      RECT  75.95 88.75 76.16 88.34 ;
      RECT  75.95 89.425 76.16 89.045 ;
      RECT  73.55 89.425 73.76 89.045 ;
      RECT  75.23 89.755 75.41 88.84 ;
      RECT  75.23 88.84 75.41 87.135 ;
      RECT  76.67 89.045 76.88 88.84 ;
      RECT  73.76 89.045 73.97 88.84 ;
      RECT  73.55 89.755 73.76 89.425 ;
      RECT  75.59 89.755 75.77 88.84 ;
      RECT  74.15 89.755 74.33 88.84 ;
      POLYGON  76.595 89.755 76.595 89.425 76.16 89.425 76.16 89.045 76.595 89.045 76.595 88.84 76.67 88.84 76.67 89.755 76.595 89.755 ;
      RECT  74.87 88.84 75.05 87.135 ;
      RECT  76.595 89.63 76.67 91.335 ;
      RECT  76.67 89.045 76.88 89.425 ;
      RECT  74.51 88.715 74.69 89.63 ;
      POLYGON  76.16 89.72 76.16 90.13 76.335 90.13 76.415 90.05 76.415 89.72 76.16 89.72 ;
      RECT  74.15 89.63 74.33 91.335 ;
      RECT  74.51 89.63 74.69 91.335 ;
      RECT  73.76 89.63 73.97 91.335 ;
      RECT  73.55 89.425 73.76 89.63 ;
      RECT  73.55 89.63 73.76 91.335 ;
      RECT  76.67 89.63 76.88 91.335 ;
      POLYGON  76.16 90.71 76.16 91.12 76.415 91.12 76.415 90.79 76.335 90.71 76.16 90.71 ;
      RECT  73.76 89.045 73.97 89.425 ;
      RECT  76.67 88.715 76.88 89.045 ;
      RECT  74.87 88.715 75.05 89.63 ;
      RECT  76.51 90.215 76.595 90.625 ;
      RECT  75.59 89.63 75.77 91.335 ;
      RECT  75.95 90.71 76.16 91.12 ;
      RECT  73.76 88.715 73.97 89.045 ;
      RECT  75.95 89.72 76.16 90.13 ;
      RECT  75.95 89.045 76.16 89.425 ;
      RECT  73.55 89.045 73.76 89.425 ;
      RECT  75.23 88.715 75.41 89.63 ;
      RECT  75.23 89.63 75.41 91.335 ;
      RECT  76.67 89.425 76.88 89.63 ;
      RECT  73.76 89.425 73.97 89.63 ;
      RECT  73.55 88.715 73.76 89.045 ;
      RECT  75.59 88.715 75.77 89.63 ;
      RECT  74.15 88.715 74.33 89.63 ;
      POLYGON  76.595 88.715 76.595 89.045 76.16 89.045 76.16 89.425 76.595 89.425 76.595 89.63 76.67 89.63 76.67 88.715 76.595 88.715 ;
      RECT  74.87 89.63 75.05 91.335 ;
      RECT  76.595 92.79 76.67 91.085 ;
      RECT  76.67 93.375 76.88 92.995 ;
      RECT  74.51 93.705 74.69 92.79 ;
      POLYGON  76.16 92.7 76.16 92.29 76.335 92.29 76.415 92.37 76.415 92.7 76.16 92.7 ;
      RECT  74.15 92.79 74.33 91.085 ;
      RECT  74.51 92.79 74.69 91.085 ;
      RECT  73.76 92.79 73.97 91.085 ;
      RECT  73.55 92.995 73.76 92.79 ;
      RECT  73.55 92.79 73.76 91.085 ;
      RECT  76.67 92.79 76.88 91.085 ;
      POLYGON  76.16 91.71 76.16 91.3 76.415 91.3 76.415 91.63 76.335 91.71 76.16 91.71 ;
      RECT  73.76 93.375 73.97 92.995 ;
      RECT  76.67 93.705 76.88 93.375 ;
      RECT  74.87 93.705 75.05 92.79 ;
      RECT  76.51 92.205 76.595 91.795 ;
      RECT  75.59 92.79 75.77 91.085 ;
      RECT  75.95 91.71 76.16 91.3 ;
      RECT  73.76 93.705 73.97 93.375 ;
      RECT  75.95 92.7 76.16 92.29 ;
      RECT  75.95 93.375 76.16 92.995 ;
      RECT  73.55 93.375 73.76 92.995 ;
      RECT  75.23 93.705 75.41 92.79 ;
      RECT  75.23 92.79 75.41 91.085 ;
      RECT  76.67 92.995 76.88 92.79 ;
      RECT  73.76 92.995 73.97 92.79 ;
      RECT  73.55 93.705 73.76 93.375 ;
      RECT  75.59 93.705 75.77 92.79 ;
      RECT  74.15 93.705 74.33 92.79 ;
      POLYGON  76.595 93.705 76.595 93.375 76.16 93.375 76.16 92.995 76.595 92.995 76.595 92.79 76.67 92.79 76.67 93.705 76.595 93.705 ;
      RECT  74.87 92.79 75.05 91.085 ;
      RECT  77.165 61.98 77.09 63.685 ;
      RECT  77.09 61.395 76.88 61.775 ;
      RECT  79.25 61.065 79.07 61.98 ;
      POLYGON  77.6 62.07 77.6 62.48 77.425 62.48 77.345 62.4 77.345 62.07 77.6 62.07 ;
      RECT  79.61 61.98 79.43 63.685 ;
      RECT  79.25 61.98 79.07 63.685 ;
      RECT  80.0 61.98 79.79 63.685 ;
      RECT  80.21 61.775 80.0 61.98 ;
      RECT  80.21 61.98 80.0 63.685 ;
      RECT  77.09 61.98 76.88 63.685 ;
      POLYGON  77.6 63.06 77.6 63.47 77.345 63.47 77.345 63.14 77.425 63.06 77.6 63.06 ;
      RECT  80.0 61.395 79.79 61.775 ;
      RECT  77.09 61.065 76.88 61.395 ;
      RECT  78.89 61.065 78.71 61.98 ;
      RECT  77.25 62.565 77.165 62.975 ;
      RECT  78.17 61.98 77.99 63.685 ;
      RECT  77.81 63.06 77.6 63.47 ;
      RECT  80.0 61.065 79.79 61.395 ;
      RECT  77.81 62.07 77.6 62.48 ;
      RECT  77.81 61.395 77.6 61.775 ;
      RECT  80.21 61.395 80.0 61.775 ;
      RECT  78.53 61.065 78.35 61.98 ;
      RECT  78.53 61.98 78.35 63.685 ;
      RECT  77.09 61.775 76.88 61.98 ;
      RECT  80.0 61.775 79.79 61.98 ;
      RECT  80.21 61.065 80.0 61.395 ;
      RECT  78.17 61.065 77.99 61.98 ;
      RECT  79.61 61.065 79.43 61.98 ;
      POLYGON  77.165 61.065 77.165 61.395 77.6 61.395 77.6 61.775 77.165 61.775 77.165 61.98 77.09 61.98 77.09 61.065 77.165 61.065 ;
      RECT  78.89 61.98 78.71 63.685 ;
      RECT  77.165 65.14 77.09 63.435 ;
      RECT  77.09 65.725 76.88 65.345 ;
      RECT  79.25 66.055 79.07 65.14 ;
      POLYGON  77.6 65.05 77.6 64.64 77.425 64.64 77.345 64.72 77.345 65.05 77.6 65.05 ;
      RECT  79.61 65.14 79.43 63.435 ;
      RECT  79.25 65.14 79.07 63.435 ;
      RECT  80.0 65.14 79.79 63.435 ;
      RECT  80.21 65.345 80.0 65.14 ;
      RECT  80.21 65.14 80.0 63.435 ;
      RECT  77.09 65.14 76.88 63.435 ;
      POLYGON  77.6 64.06 77.6 63.65 77.345 63.65 77.345 63.98 77.425 64.06 77.6 64.06 ;
      RECT  80.0 65.725 79.79 65.345 ;
      RECT  77.09 66.055 76.88 65.725 ;
      RECT  78.89 66.055 78.71 65.14 ;
      RECT  77.25 64.555 77.165 64.145 ;
      RECT  78.17 65.14 77.99 63.435 ;
      RECT  77.81 64.06 77.6 63.65 ;
      RECT  80.0 66.055 79.79 65.725 ;
      RECT  77.81 65.05 77.6 64.64 ;
      RECT  77.81 65.725 77.6 65.345 ;
      RECT  80.21 65.725 80.0 65.345 ;
      RECT  78.53 66.055 78.35 65.14 ;
      RECT  78.53 65.14 78.35 63.435 ;
      RECT  77.09 65.345 76.88 65.14 ;
      RECT  80.0 65.345 79.79 65.14 ;
      RECT  80.21 66.055 80.0 65.725 ;
      RECT  78.17 66.055 77.99 65.14 ;
      RECT  79.61 66.055 79.43 65.14 ;
      POLYGON  77.165 66.055 77.165 65.725 77.6 65.725 77.6 65.345 77.165 65.345 77.165 65.14 77.09 65.14 77.09 66.055 77.165 66.055 ;
      RECT  78.89 65.14 78.71 63.435 ;
      RECT  77.165 65.93 77.09 67.635 ;
      RECT  77.09 65.345 76.88 65.725 ;
      RECT  79.25 65.015 79.07 65.93 ;
      POLYGON  77.6 66.02 77.6 66.43 77.425 66.43 77.345 66.35 77.345 66.02 77.6 66.02 ;
      RECT  79.61 65.93 79.43 67.635 ;
      RECT  79.25 65.93 79.07 67.635 ;
      RECT  80.0 65.93 79.79 67.635 ;
      RECT  80.21 65.725 80.0 65.93 ;
      RECT  80.21 65.93 80.0 67.635 ;
      RECT  77.09 65.93 76.88 67.635 ;
      POLYGON  77.6 67.01 77.6 67.42 77.345 67.42 77.345 67.09 77.425 67.01 77.6 67.01 ;
      RECT  80.0 65.345 79.79 65.725 ;
      RECT  77.09 65.015 76.88 65.345 ;
      RECT  78.89 65.015 78.71 65.93 ;
      RECT  77.25 66.515 77.165 66.925 ;
      RECT  78.17 65.93 77.99 67.635 ;
      RECT  77.81 67.01 77.6 67.42 ;
      RECT  80.0 65.015 79.79 65.345 ;
      RECT  77.81 66.02 77.6 66.43 ;
      RECT  77.81 65.345 77.6 65.725 ;
      RECT  80.21 65.345 80.0 65.725 ;
      RECT  78.53 65.015 78.35 65.93 ;
      RECT  78.53 65.93 78.35 67.635 ;
      RECT  77.09 65.725 76.88 65.93 ;
      RECT  80.0 65.725 79.79 65.93 ;
      RECT  80.21 65.015 80.0 65.345 ;
      RECT  78.17 65.015 77.99 65.93 ;
      RECT  79.61 65.015 79.43 65.93 ;
      POLYGON  77.165 65.015 77.165 65.345 77.6 65.345 77.6 65.725 77.165 65.725 77.165 65.93 77.09 65.93 77.09 65.015 77.165 65.015 ;
      RECT  78.89 65.93 78.71 67.635 ;
      RECT  77.165 69.09 77.09 67.385 ;
      RECT  77.09 69.675 76.88 69.295 ;
      RECT  79.25 70.005 79.07 69.09 ;
      POLYGON  77.6 69.0 77.6 68.59 77.425 68.59 77.345 68.67 77.345 69.0 77.6 69.0 ;
      RECT  79.61 69.09 79.43 67.385 ;
      RECT  79.25 69.09 79.07 67.385 ;
      RECT  80.0 69.09 79.79 67.385 ;
      RECT  80.21 69.295 80.0 69.09 ;
      RECT  80.21 69.09 80.0 67.385 ;
      RECT  77.09 69.09 76.88 67.385 ;
      POLYGON  77.6 68.01 77.6 67.6 77.345 67.6 77.345 67.93 77.425 68.01 77.6 68.01 ;
      RECT  80.0 69.675 79.79 69.295 ;
      RECT  77.09 70.005 76.88 69.675 ;
      RECT  78.89 70.005 78.71 69.09 ;
      RECT  77.25 68.505 77.165 68.095 ;
      RECT  78.17 69.09 77.99 67.385 ;
      RECT  77.81 68.01 77.6 67.6 ;
      RECT  80.0 70.005 79.79 69.675 ;
      RECT  77.81 69.0 77.6 68.59 ;
      RECT  77.81 69.675 77.6 69.295 ;
      RECT  80.21 69.675 80.0 69.295 ;
      RECT  78.53 70.005 78.35 69.09 ;
      RECT  78.53 69.09 78.35 67.385 ;
      RECT  77.09 69.295 76.88 69.09 ;
      RECT  80.0 69.295 79.79 69.09 ;
      RECT  80.21 70.005 80.0 69.675 ;
      RECT  78.17 70.005 77.99 69.09 ;
      RECT  79.61 70.005 79.43 69.09 ;
      POLYGON  77.165 70.005 77.165 69.675 77.6 69.675 77.6 69.295 77.165 69.295 77.165 69.09 77.09 69.09 77.09 70.005 77.165 70.005 ;
      RECT  78.89 69.09 78.71 67.385 ;
      RECT  77.165 69.88 77.09 71.585 ;
      RECT  77.09 69.295 76.88 69.675 ;
      RECT  79.25 68.965 79.07 69.88 ;
      POLYGON  77.6 69.97 77.6 70.38 77.425 70.38 77.345 70.3 77.345 69.97 77.6 69.97 ;
      RECT  79.61 69.88 79.43 71.585 ;
      RECT  79.25 69.88 79.07 71.585 ;
      RECT  80.0 69.88 79.79 71.585 ;
      RECT  80.21 69.675 80.0 69.88 ;
      RECT  80.21 69.88 80.0 71.585 ;
      RECT  77.09 69.88 76.88 71.585 ;
      POLYGON  77.6 70.96 77.6 71.37 77.345 71.37 77.345 71.04 77.425 70.96 77.6 70.96 ;
      RECT  80.0 69.295 79.79 69.675 ;
      RECT  77.09 68.965 76.88 69.295 ;
      RECT  78.89 68.965 78.71 69.88 ;
      RECT  77.25 70.465 77.165 70.875 ;
      RECT  78.17 69.88 77.99 71.585 ;
      RECT  77.81 70.96 77.6 71.37 ;
      RECT  80.0 68.965 79.79 69.295 ;
      RECT  77.81 69.97 77.6 70.38 ;
      RECT  77.81 69.295 77.6 69.675 ;
      RECT  80.21 69.295 80.0 69.675 ;
      RECT  78.53 68.965 78.35 69.88 ;
      RECT  78.53 69.88 78.35 71.585 ;
      RECT  77.09 69.675 76.88 69.88 ;
      RECT  80.0 69.675 79.79 69.88 ;
      RECT  80.21 68.965 80.0 69.295 ;
      RECT  78.17 68.965 77.99 69.88 ;
      RECT  79.61 68.965 79.43 69.88 ;
      POLYGON  77.165 68.965 77.165 69.295 77.6 69.295 77.6 69.675 77.165 69.675 77.165 69.88 77.09 69.88 77.09 68.965 77.165 68.965 ;
      RECT  78.89 69.88 78.71 71.585 ;
      RECT  77.165 73.04 77.09 71.335 ;
      RECT  77.09 73.625 76.88 73.245 ;
      RECT  79.25 73.955 79.07 73.04 ;
      POLYGON  77.6 72.95 77.6 72.54 77.425 72.54 77.345 72.62 77.345 72.95 77.6 72.95 ;
      RECT  79.61 73.04 79.43 71.335 ;
      RECT  79.25 73.04 79.07 71.335 ;
      RECT  80.0 73.04 79.79 71.335 ;
      RECT  80.21 73.245 80.0 73.04 ;
      RECT  80.21 73.04 80.0 71.335 ;
      RECT  77.09 73.04 76.88 71.335 ;
      POLYGON  77.6 71.96 77.6 71.55 77.345 71.55 77.345 71.88 77.425 71.96 77.6 71.96 ;
      RECT  80.0 73.625 79.79 73.245 ;
      RECT  77.09 73.955 76.88 73.625 ;
      RECT  78.89 73.955 78.71 73.04 ;
      RECT  77.25 72.455 77.165 72.045 ;
      RECT  78.17 73.04 77.99 71.335 ;
      RECT  77.81 71.96 77.6 71.55 ;
      RECT  80.0 73.955 79.79 73.625 ;
      RECT  77.81 72.95 77.6 72.54 ;
      RECT  77.81 73.625 77.6 73.245 ;
      RECT  80.21 73.625 80.0 73.245 ;
      RECT  78.53 73.955 78.35 73.04 ;
      RECT  78.53 73.04 78.35 71.335 ;
      RECT  77.09 73.245 76.88 73.04 ;
      RECT  80.0 73.245 79.79 73.04 ;
      RECT  80.21 73.955 80.0 73.625 ;
      RECT  78.17 73.955 77.99 73.04 ;
      RECT  79.61 73.955 79.43 73.04 ;
      POLYGON  77.165 73.955 77.165 73.625 77.6 73.625 77.6 73.245 77.165 73.245 77.165 73.04 77.09 73.04 77.09 73.955 77.165 73.955 ;
      RECT  78.89 73.04 78.71 71.335 ;
      RECT  77.165 73.83 77.09 75.535 ;
      RECT  77.09 73.245 76.88 73.625 ;
      RECT  79.25 72.915 79.07 73.83 ;
      POLYGON  77.6 73.92 77.6 74.33 77.425 74.33 77.345 74.25 77.345 73.92 77.6 73.92 ;
      RECT  79.61 73.83 79.43 75.535 ;
      RECT  79.25 73.83 79.07 75.535 ;
      RECT  80.0 73.83 79.79 75.535 ;
      RECT  80.21 73.625 80.0 73.83 ;
      RECT  80.21 73.83 80.0 75.535 ;
      RECT  77.09 73.83 76.88 75.535 ;
      POLYGON  77.6 74.91 77.6 75.32 77.345 75.32 77.345 74.99 77.425 74.91 77.6 74.91 ;
      RECT  80.0 73.245 79.79 73.625 ;
      RECT  77.09 72.915 76.88 73.245 ;
      RECT  78.89 72.915 78.71 73.83 ;
      RECT  77.25 74.415 77.165 74.825 ;
      RECT  78.17 73.83 77.99 75.535 ;
      RECT  77.81 74.91 77.6 75.32 ;
      RECT  80.0 72.915 79.79 73.245 ;
      RECT  77.81 73.92 77.6 74.33 ;
      RECT  77.81 73.245 77.6 73.625 ;
      RECT  80.21 73.245 80.0 73.625 ;
      RECT  78.53 72.915 78.35 73.83 ;
      RECT  78.53 73.83 78.35 75.535 ;
      RECT  77.09 73.625 76.88 73.83 ;
      RECT  80.0 73.625 79.79 73.83 ;
      RECT  80.21 72.915 80.0 73.245 ;
      RECT  78.17 72.915 77.99 73.83 ;
      RECT  79.61 72.915 79.43 73.83 ;
      POLYGON  77.165 72.915 77.165 73.245 77.6 73.245 77.6 73.625 77.165 73.625 77.165 73.83 77.09 73.83 77.09 72.915 77.165 72.915 ;
      RECT  78.89 73.83 78.71 75.535 ;
      RECT  77.165 76.99 77.09 75.285 ;
      RECT  77.09 77.575 76.88 77.195 ;
      RECT  79.25 77.905 79.07 76.99 ;
      POLYGON  77.6 76.9 77.6 76.49 77.425 76.49 77.345 76.57 77.345 76.9 77.6 76.9 ;
      RECT  79.61 76.99 79.43 75.285 ;
      RECT  79.25 76.99 79.07 75.285 ;
      RECT  80.0 76.99 79.79 75.285 ;
      RECT  80.21 77.195 80.0 76.99 ;
      RECT  80.21 76.99 80.0 75.285 ;
      RECT  77.09 76.99 76.88 75.285 ;
      POLYGON  77.6 75.91 77.6 75.5 77.345 75.5 77.345 75.83 77.425 75.91 77.6 75.91 ;
      RECT  80.0 77.575 79.79 77.195 ;
      RECT  77.09 77.905 76.88 77.575 ;
      RECT  78.89 77.905 78.71 76.99 ;
      RECT  77.25 76.405 77.165 75.995 ;
      RECT  78.17 76.99 77.99 75.285 ;
      RECT  77.81 75.91 77.6 75.5 ;
      RECT  80.0 77.905 79.79 77.575 ;
      RECT  77.81 76.9 77.6 76.49 ;
      RECT  77.81 77.575 77.6 77.195 ;
      RECT  80.21 77.575 80.0 77.195 ;
      RECT  78.53 77.905 78.35 76.99 ;
      RECT  78.53 76.99 78.35 75.285 ;
      RECT  77.09 77.195 76.88 76.99 ;
      RECT  80.0 77.195 79.79 76.99 ;
      RECT  80.21 77.905 80.0 77.575 ;
      RECT  78.17 77.905 77.99 76.99 ;
      RECT  79.61 77.905 79.43 76.99 ;
      POLYGON  77.165 77.905 77.165 77.575 77.6 77.575 77.6 77.195 77.165 77.195 77.165 76.99 77.09 76.99 77.09 77.905 77.165 77.905 ;
      RECT  78.89 76.99 78.71 75.285 ;
      RECT  77.165 77.78 77.09 79.485 ;
      RECT  77.09 77.195 76.88 77.575 ;
      RECT  79.25 76.865 79.07 77.78 ;
      POLYGON  77.6 77.87 77.6 78.28 77.425 78.28 77.345 78.2 77.345 77.87 77.6 77.87 ;
      RECT  79.61 77.78 79.43 79.485 ;
      RECT  79.25 77.78 79.07 79.485 ;
      RECT  80.0 77.78 79.79 79.485 ;
      RECT  80.21 77.575 80.0 77.78 ;
      RECT  80.21 77.78 80.0 79.485 ;
      RECT  77.09 77.78 76.88 79.485 ;
      POLYGON  77.6 78.86 77.6 79.27 77.345 79.27 77.345 78.94 77.425 78.86 77.6 78.86 ;
      RECT  80.0 77.195 79.79 77.575 ;
      RECT  77.09 76.865 76.88 77.195 ;
      RECT  78.89 76.865 78.71 77.78 ;
      RECT  77.25 78.365 77.165 78.775 ;
      RECT  78.17 77.78 77.99 79.485 ;
      RECT  77.81 78.86 77.6 79.27 ;
      RECT  80.0 76.865 79.79 77.195 ;
      RECT  77.81 77.87 77.6 78.28 ;
      RECT  77.81 77.195 77.6 77.575 ;
      RECT  80.21 77.195 80.0 77.575 ;
      RECT  78.53 76.865 78.35 77.78 ;
      RECT  78.53 77.78 78.35 79.485 ;
      RECT  77.09 77.575 76.88 77.78 ;
      RECT  80.0 77.575 79.79 77.78 ;
      RECT  80.21 76.865 80.0 77.195 ;
      RECT  78.17 76.865 77.99 77.78 ;
      RECT  79.61 76.865 79.43 77.78 ;
      POLYGON  77.165 76.865 77.165 77.195 77.6 77.195 77.6 77.575 77.165 77.575 77.165 77.78 77.09 77.78 77.09 76.865 77.165 76.865 ;
      RECT  78.89 77.78 78.71 79.485 ;
      RECT  77.165 80.94 77.09 79.235 ;
      RECT  77.09 81.525 76.88 81.145 ;
      RECT  79.25 81.855 79.07 80.94 ;
      POLYGON  77.6 80.85 77.6 80.44 77.425 80.44 77.345 80.52 77.345 80.85 77.6 80.85 ;
      RECT  79.61 80.94 79.43 79.235 ;
      RECT  79.25 80.94 79.07 79.235 ;
      RECT  80.0 80.94 79.79 79.235 ;
      RECT  80.21 81.145 80.0 80.94 ;
      RECT  80.21 80.94 80.0 79.235 ;
      RECT  77.09 80.94 76.88 79.235 ;
      POLYGON  77.6 79.86 77.6 79.45 77.345 79.45 77.345 79.78 77.425 79.86 77.6 79.86 ;
      RECT  80.0 81.525 79.79 81.145 ;
      RECT  77.09 81.855 76.88 81.525 ;
      RECT  78.89 81.855 78.71 80.94 ;
      RECT  77.25 80.355 77.165 79.945 ;
      RECT  78.17 80.94 77.99 79.235 ;
      RECT  77.81 79.86 77.6 79.45 ;
      RECT  80.0 81.855 79.79 81.525 ;
      RECT  77.81 80.85 77.6 80.44 ;
      RECT  77.81 81.525 77.6 81.145 ;
      RECT  80.21 81.525 80.0 81.145 ;
      RECT  78.53 81.855 78.35 80.94 ;
      RECT  78.53 80.94 78.35 79.235 ;
      RECT  77.09 81.145 76.88 80.94 ;
      RECT  80.0 81.145 79.79 80.94 ;
      RECT  80.21 81.855 80.0 81.525 ;
      RECT  78.17 81.855 77.99 80.94 ;
      RECT  79.61 81.855 79.43 80.94 ;
      POLYGON  77.165 81.855 77.165 81.525 77.6 81.525 77.6 81.145 77.165 81.145 77.165 80.94 77.09 80.94 77.09 81.855 77.165 81.855 ;
      RECT  78.89 80.94 78.71 79.235 ;
      RECT  77.165 81.73 77.09 83.435 ;
      RECT  77.09 81.145 76.88 81.525 ;
      RECT  79.25 80.815 79.07 81.73 ;
      POLYGON  77.6 81.82 77.6 82.23 77.425 82.23 77.345 82.15 77.345 81.82 77.6 81.82 ;
      RECT  79.61 81.73 79.43 83.435 ;
      RECT  79.25 81.73 79.07 83.435 ;
      RECT  80.0 81.73 79.79 83.435 ;
      RECT  80.21 81.525 80.0 81.73 ;
      RECT  80.21 81.73 80.0 83.435 ;
      RECT  77.09 81.73 76.88 83.435 ;
      POLYGON  77.6 82.81 77.6 83.22 77.345 83.22 77.345 82.89 77.425 82.81 77.6 82.81 ;
      RECT  80.0 81.145 79.79 81.525 ;
      RECT  77.09 80.815 76.88 81.145 ;
      RECT  78.89 80.815 78.71 81.73 ;
      RECT  77.25 82.315 77.165 82.725 ;
      RECT  78.17 81.73 77.99 83.435 ;
      RECT  77.81 82.81 77.6 83.22 ;
      RECT  80.0 80.815 79.79 81.145 ;
      RECT  77.81 81.82 77.6 82.23 ;
      RECT  77.81 81.145 77.6 81.525 ;
      RECT  80.21 81.145 80.0 81.525 ;
      RECT  78.53 80.815 78.35 81.73 ;
      RECT  78.53 81.73 78.35 83.435 ;
      RECT  77.09 81.525 76.88 81.73 ;
      RECT  80.0 81.525 79.79 81.73 ;
      RECT  80.21 80.815 80.0 81.145 ;
      RECT  78.17 80.815 77.99 81.73 ;
      RECT  79.61 80.815 79.43 81.73 ;
      POLYGON  77.165 80.815 77.165 81.145 77.6 81.145 77.6 81.525 77.165 81.525 77.165 81.73 77.09 81.73 77.09 80.815 77.165 80.815 ;
      RECT  78.89 81.73 78.71 83.435 ;
      RECT  77.165 84.89 77.09 83.185 ;
      RECT  77.09 85.475 76.88 85.095 ;
      RECT  79.25 85.805 79.07 84.89 ;
      POLYGON  77.6 84.8 77.6 84.39 77.425 84.39 77.345 84.47 77.345 84.8 77.6 84.8 ;
      RECT  79.61 84.89 79.43 83.185 ;
      RECT  79.25 84.89 79.07 83.185 ;
      RECT  80.0 84.89 79.79 83.185 ;
      RECT  80.21 85.095 80.0 84.89 ;
      RECT  80.21 84.89 80.0 83.185 ;
      RECT  77.09 84.89 76.88 83.185 ;
      POLYGON  77.6 83.81 77.6 83.4 77.345 83.4 77.345 83.73 77.425 83.81 77.6 83.81 ;
      RECT  80.0 85.475 79.79 85.095 ;
      RECT  77.09 85.805 76.88 85.475 ;
      RECT  78.89 85.805 78.71 84.89 ;
      RECT  77.25 84.305 77.165 83.895 ;
      RECT  78.17 84.89 77.99 83.185 ;
      RECT  77.81 83.81 77.6 83.4 ;
      RECT  80.0 85.805 79.79 85.475 ;
      RECT  77.81 84.8 77.6 84.39 ;
      RECT  77.81 85.475 77.6 85.095 ;
      RECT  80.21 85.475 80.0 85.095 ;
      RECT  78.53 85.805 78.35 84.89 ;
      RECT  78.53 84.89 78.35 83.185 ;
      RECT  77.09 85.095 76.88 84.89 ;
      RECT  80.0 85.095 79.79 84.89 ;
      RECT  80.21 85.805 80.0 85.475 ;
      RECT  78.17 85.805 77.99 84.89 ;
      RECT  79.61 85.805 79.43 84.89 ;
      POLYGON  77.165 85.805 77.165 85.475 77.6 85.475 77.6 85.095 77.165 85.095 77.165 84.89 77.09 84.89 77.09 85.805 77.165 85.805 ;
      RECT  78.89 84.89 78.71 83.185 ;
      RECT  77.165 85.68 77.09 87.385 ;
      RECT  77.09 85.095 76.88 85.475 ;
      RECT  79.25 84.765 79.07 85.68 ;
      POLYGON  77.6 85.77 77.6 86.18 77.425 86.18 77.345 86.1 77.345 85.77 77.6 85.77 ;
      RECT  79.61 85.68 79.43 87.385 ;
      RECT  79.25 85.68 79.07 87.385 ;
      RECT  80.0 85.68 79.79 87.385 ;
      RECT  80.21 85.475 80.0 85.68 ;
      RECT  80.21 85.68 80.0 87.385 ;
      RECT  77.09 85.68 76.88 87.385 ;
      POLYGON  77.6 86.76 77.6 87.17 77.345 87.17 77.345 86.84 77.425 86.76 77.6 86.76 ;
      RECT  80.0 85.095 79.79 85.475 ;
      RECT  77.09 84.765 76.88 85.095 ;
      RECT  78.89 84.765 78.71 85.68 ;
      RECT  77.25 86.265 77.165 86.675 ;
      RECT  78.17 85.68 77.99 87.385 ;
      RECT  77.81 86.76 77.6 87.17 ;
      RECT  80.0 84.765 79.79 85.095 ;
      RECT  77.81 85.77 77.6 86.18 ;
      RECT  77.81 85.095 77.6 85.475 ;
      RECT  80.21 85.095 80.0 85.475 ;
      RECT  78.53 84.765 78.35 85.68 ;
      RECT  78.53 85.68 78.35 87.385 ;
      RECT  77.09 85.475 76.88 85.68 ;
      RECT  80.0 85.475 79.79 85.68 ;
      RECT  80.21 84.765 80.0 85.095 ;
      RECT  78.17 84.765 77.99 85.68 ;
      RECT  79.61 84.765 79.43 85.68 ;
      POLYGON  77.165 84.765 77.165 85.095 77.6 85.095 77.6 85.475 77.165 85.475 77.165 85.68 77.09 85.68 77.09 84.765 77.165 84.765 ;
      RECT  78.89 85.68 78.71 87.385 ;
      RECT  77.165 88.84 77.09 87.135 ;
      RECT  77.09 89.425 76.88 89.045 ;
      RECT  79.25 89.755 79.07 88.84 ;
      POLYGON  77.6 88.75 77.6 88.34 77.425 88.34 77.345 88.42 77.345 88.75 77.6 88.75 ;
      RECT  79.61 88.84 79.43 87.135 ;
      RECT  79.25 88.84 79.07 87.135 ;
      RECT  80.0 88.84 79.79 87.135 ;
      RECT  80.21 89.045 80.0 88.84 ;
      RECT  80.21 88.84 80.0 87.135 ;
      RECT  77.09 88.84 76.88 87.135 ;
      POLYGON  77.6 87.76 77.6 87.35 77.345 87.35 77.345 87.68 77.425 87.76 77.6 87.76 ;
      RECT  80.0 89.425 79.79 89.045 ;
      RECT  77.09 89.755 76.88 89.425 ;
      RECT  78.89 89.755 78.71 88.84 ;
      RECT  77.25 88.255 77.165 87.845 ;
      RECT  78.17 88.84 77.99 87.135 ;
      RECT  77.81 87.76 77.6 87.35 ;
      RECT  80.0 89.755 79.79 89.425 ;
      RECT  77.81 88.75 77.6 88.34 ;
      RECT  77.81 89.425 77.6 89.045 ;
      RECT  80.21 89.425 80.0 89.045 ;
      RECT  78.53 89.755 78.35 88.84 ;
      RECT  78.53 88.84 78.35 87.135 ;
      RECT  77.09 89.045 76.88 88.84 ;
      RECT  80.0 89.045 79.79 88.84 ;
      RECT  80.21 89.755 80.0 89.425 ;
      RECT  78.17 89.755 77.99 88.84 ;
      RECT  79.61 89.755 79.43 88.84 ;
      POLYGON  77.165 89.755 77.165 89.425 77.6 89.425 77.6 89.045 77.165 89.045 77.165 88.84 77.09 88.84 77.09 89.755 77.165 89.755 ;
      RECT  78.89 88.84 78.71 87.135 ;
      RECT  77.165 89.63 77.09 91.335 ;
      RECT  77.09 89.045 76.88 89.425 ;
      RECT  79.25 88.715 79.07 89.63 ;
      POLYGON  77.6 89.72 77.6 90.13 77.425 90.13 77.345 90.05 77.345 89.72 77.6 89.72 ;
      RECT  79.61 89.63 79.43 91.335 ;
      RECT  79.25 89.63 79.07 91.335 ;
      RECT  80.0 89.63 79.79 91.335 ;
      RECT  80.21 89.425 80.0 89.63 ;
      RECT  80.21 89.63 80.0 91.335 ;
      RECT  77.09 89.63 76.88 91.335 ;
      POLYGON  77.6 90.71 77.6 91.12 77.345 91.12 77.345 90.79 77.425 90.71 77.6 90.71 ;
      RECT  80.0 89.045 79.79 89.425 ;
      RECT  77.09 88.715 76.88 89.045 ;
      RECT  78.89 88.715 78.71 89.63 ;
      RECT  77.25 90.215 77.165 90.625 ;
      RECT  78.17 89.63 77.99 91.335 ;
      RECT  77.81 90.71 77.6 91.12 ;
      RECT  80.0 88.715 79.79 89.045 ;
      RECT  77.81 89.72 77.6 90.13 ;
      RECT  77.81 89.045 77.6 89.425 ;
      RECT  80.21 89.045 80.0 89.425 ;
      RECT  78.53 88.715 78.35 89.63 ;
      RECT  78.53 89.63 78.35 91.335 ;
      RECT  77.09 89.425 76.88 89.63 ;
      RECT  80.0 89.425 79.79 89.63 ;
      RECT  80.21 88.715 80.0 89.045 ;
      RECT  78.17 88.715 77.99 89.63 ;
      RECT  79.61 88.715 79.43 89.63 ;
      POLYGON  77.165 88.715 77.165 89.045 77.6 89.045 77.6 89.425 77.165 89.425 77.165 89.63 77.09 89.63 77.09 88.715 77.165 88.715 ;
      RECT  78.89 89.63 78.71 91.335 ;
      RECT  77.165 92.79 77.09 91.085 ;
      RECT  77.09 93.375 76.88 92.995 ;
      RECT  79.25 93.705 79.07 92.79 ;
      POLYGON  77.6 92.7 77.6 92.29 77.425 92.29 77.345 92.37 77.345 92.7 77.6 92.7 ;
      RECT  79.61 92.79 79.43 91.085 ;
      RECT  79.25 92.79 79.07 91.085 ;
      RECT  80.0 92.79 79.79 91.085 ;
      RECT  80.21 92.995 80.0 92.79 ;
      RECT  80.21 92.79 80.0 91.085 ;
      RECT  77.09 92.79 76.88 91.085 ;
      POLYGON  77.6 91.71 77.6 91.3 77.345 91.3 77.345 91.63 77.425 91.71 77.6 91.71 ;
      RECT  80.0 93.375 79.79 92.995 ;
      RECT  77.09 93.705 76.88 93.375 ;
      RECT  78.89 93.705 78.71 92.79 ;
      RECT  77.25 92.205 77.165 91.795 ;
      RECT  78.17 92.79 77.99 91.085 ;
      RECT  77.81 91.71 77.6 91.3 ;
      RECT  80.0 93.705 79.79 93.375 ;
      RECT  77.81 92.7 77.6 92.29 ;
      RECT  77.81 93.375 77.6 92.995 ;
      RECT  80.21 93.375 80.0 92.995 ;
      RECT  78.53 93.705 78.35 92.79 ;
      RECT  78.53 92.79 78.35 91.085 ;
      RECT  77.09 92.995 76.88 92.79 ;
      RECT  80.0 92.995 79.79 92.79 ;
      RECT  80.21 93.705 80.0 93.375 ;
      RECT  78.17 93.705 77.99 92.79 ;
      RECT  79.61 93.705 79.43 92.79 ;
      POLYGON  77.165 93.705 77.165 93.375 77.6 93.375 77.6 92.995 77.165 92.995 77.165 92.79 77.09 92.79 77.09 93.705 77.165 93.705 ;
      RECT  78.89 92.79 78.71 91.085 ;
      RECT  74.15 61.585 74.33 93.185 ;
      RECT  74.51 61.585 74.69 93.185 ;
      RECT  75.23 61.585 75.41 93.185 ;
      RECT  75.59 61.585 75.77 93.185 ;
      RECT  79.43 61.585 79.61 93.185 ;
      RECT  79.07 61.585 79.25 93.185 ;
      RECT  78.35 61.585 78.53 93.185 ;
      RECT  77.99 61.585 78.17 93.185 ;
      RECT  74.87 85.68 75.05 87.385 ;
      RECT  74.87 61.98 75.05 63.685 ;
      RECT  74.87 87.135 75.05 88.84 ;
      RECT  74.87 71.335 75.05 73.04 ;
      RECT  78.71 65.93 78.89 67.635 ;
      RECT  78.71 91.085 78.89 92.79 ;
      RECT  78.71 67.385 78.89 69.09 ;
      RECT  78.71 87.135 78.89 88.84 ;
      RECT  74.87 65.93 75.05 67.635 ;
      RECT  78.71 77.78 78.89 79.485 ;
      RECT  74.87 69.88 75.05 71.585 ;
      RECT  74.87 77.78 75.05 79.485 ;
      RECT  74.87 79.235 75.05 80.94 ;
      RECT  74.87 83.185 75.05 84.89 ;
      RECT  74.87 89.63 75.05 91.335 ;
      RECT  74.87 67.385 75.05 69.09 ;
      RECT  78.71 73.83 78.89 75.535 ;
      RECT  78.71 63.435 78.89 65.14 ;
      RECT  74.87 91.085 75.05 92.79 ;
      RECT  78.71 81.73 78.89 83.435 ;
      RECT  78.71 71.335 78.89 73.04 ;
      RECT  78.71 61.98 78.89 63.685 ;
      RECT  74.87 63.435 75.05 65.14 ;
      RECT  74.87 81.73 75.05 83.435 ;
      RECT  78.71 85.68 78.89 87.385 ;
      RECT  78.71 75.285 78.89 76.99 ;
      RECT  74.87 75.285 75.05 76.99 ;
      RECT  78.71 69.88 78.89 71.585 ;
      RECT  78.71 83.185 78.89 84.89 ;
      RECT  74.87 73.83 75.05 75.535 ;
      RECT  78.71 89.63 78.89 91.335 ;
      RECT  78.71 79.235 78.89 80.94 ;
      RECT  72.65 58.425 72.47 60.005 ;
      RECT  73.01 58.425 72.83 60.005 ;
      RECT  72.56 58.425 72.43 59.135 ;
      RECT  72.29 58.425 72.11 60.005 ;
      RECT  72.69 58.425 72.56 59.135 ;
      RECT  73.01 57.635 72.83 58.425 ;
      RECT  73.37 57.635 73.19 58.425 ;
      RECT  71.93 57.635 71.75 58.425 ;
      RECT  72.65 57.635 72.47 58.425 ;
      RECT  72.29 57.635 72.11 58.425 ;
      RECT  73.37 58.425 73.19 60.005 ;
      RECT  71.93 58.425 71.75 60.005 ;
      RECT  70.925 61.19 70.85 59.485 ;
      RECT  70.85 61.775 70.64 61.395 ;
      RECT  73.01 62.105 72.83 61.19 ;
      POLYGON  71.36 61.1 71.36 60.69 71.185 60.69 71.105 60.77 71.105 61.1 71.36 61.1 ;
      RECT  73.37 61.19 73.19 59.485 ;
      RECT  73.01 61.19 72.83 59.485 ;
      RECT  73.76 61.19 73.55 59.485 ;
      RECT  73.97 61.395 73.76 61.19 ;
      RECT  73.97 61.19 73.76 59.485 ;
      RECT  70.85 61.19 70.64 59.485 ;
      POLYGON  71.36 60.11 71.36 59.7 71.105 59.7 71.105 60.03 71.185 60.11 71.36 60.11 ;
      RECT  73.76 61.775 73.55 61.395 ;
      RECT  70.85 62.105 70.64 61.775 ;
      RECT  72.65 62.105 72.47 61.19 ;
      RECT  71.01 60.605 70.925 60.195 ;
      RECT  71.93 61.19 71.75 59.485 ;
      RECT  71.57 60.11 71.36 59.7 ;
      RECT  73.76 62.105 73.55 61.775 ;
      RECT  71.57 61.1 71.36 60.69 ;
      RECT  71.57 61.775 71.36 61.395 ;
      RECT  73.97 61.775 73.76 61.395 ;
      RECT  72.29 62.105 72.11 61.19 ;
      RECT  72.29 61.19 72.11 59.485 ;
      RECT  70.85 61.395 70.64 61.19 ;
      RECT  73.76 61.395 73.55 61.19 ;
      RECT  73.97 62.105 73.76 61.775 ;
      RECT  71.93 62.105 71.75 61.19 ;
      RECT  73.37 62.105 73.19 61.19 ;
      POLYGON  70.925 62.105 70.925 61.775 71.36 61.775 71.36 61.395 70.925 61.395 70.925 61.19 70.85 61.19 70.85 62.105 70.925 62.105 ;
      RECT  72.65 61.19 72.47 59.485 ;
      RECT  70.925 61.98 70.85 63.685 ;
      RECT  70.85 61.395 70.64 61.775 ;
      RECT  73.01 61.065 72.83 61.98 ;
      POLYGON  71.36 62.07 71.36 62.48 71.185 62.48 71.105 62.4 71.105 62.07 71.36 62.07 ;
      RECT  73.37 61.98 73.19 63.685 ;
      RECT  73.01 61.98 72.83 63.685 ;
      RECT  73.76 61.98 73.55 63.685 ;
      RECT  73.97 61.775 73.76 61.98 ;
      RECT  73.97 61.98 73.76 63.685 ;
      RECT  70.85 61.98 70.64 63.685 ;
      POLYGON  71.36 63.06 71.36 63.47 71.105 63.47 71.105 63.14 71.185 63.06 71.36 63.06 ;
      RECT  73.76 61.395 73.55 61.775 ;
      RECT  70.85 61.065 70.64 61.395 ;
      RECT  72.65 61.065 72.47 61.98 ;
      RECT  71.01 62.565 70.925 62.975 ;
      RECT  71.93 61.98 71.75 63.685 ;
      RECT  71.57 63.06 71.36 63.47 ;
      RECT  73.76 61.065 73.55 61.395 ;
      RECT  71.57 62.07 71.36 62.48 ;
      RECT  71.57 61.395 71.36 61.775 ;
      RECT  73.97 61.395 73.76 61.775 ;
      RECT  72.29 61.065 72.11 61.98 ;
      RECT  72.29 61.98 72.11 63.685 ;
      RECT  70.85 61.775 70.64 61.98 ;
      RECT  73.76 61.775 73.55 61.98 ;
      RECT  73.97 61.065 73.76 61.395 ;
      RECT  71.93 61.065 71.75 61.98 ;
      RECT  73.37 61.065 73.19 61.98 ;
      POLYGON  70.925 61.065 70.925 61.395 71.36 61.395 71.36 61.775 70.925 61.775 70.925 61.98 70.85 61.98 70.85 61.065 70.925 61.065 ;
      RECT  72.65 61.98 72.47 63.685 ;
      RECT  70.925 65.14 70.85 63.435 ;
      RECT  70.85 65.725 70.64 65.345 ;
      RECT  73.01 66.055 72.83 65.14 ;
      POLYGON  71.36 65.05 71.36 64.64 71.185 64.64 71.105 64.72 71.105 65.05 71.36 65.05 ;
      RECT  73.37 65.14 73.19 63.435 ;
      RECT  73.01 65.14 72.83 63.435 ;
      RECT  73.76 65.14 73.55 63.435 ;
      RECT  73.97 65.345 73.76 65.14 ;
      RECT  73.97 65.14 73.76 63.435 ;
      RECT  70.85 65.14 70.64 63.435 ;
      POLYGON  71.36 64.06 71.36 63.65 71.105 63.65 71.105 63.98 71.185 64.06 71.36 64.06 ;
      RECT  73.76 65.725 73.55 65.345 ;
      RECT  70.85 66.055 70.64 65.725 ;
      RECT  72.65 66.055 72.47 65.14 ;
      RECT  71.01 64.555 70.925 64.145 ;
      RECT  71.93 65.14 71.75 63.435 ;
      RECT  71.57 64.06 71.36 63.65 ;
      RECT  73.76 66.055 73.55 65.725 ;
      RECT  71.57 65.05 71.36 64.64 ;
      RECT  71.57 65.725 71.36 65.345 ;
      RECT  73.97 65.725 73.76 65.345 ;
      RECT  72.29 66.055 72.11 65.14 ;
      RECT  72.29 65.14 72.11 63.435 ;
      RECT  70.85 65.345 70.64 65.14 ;
      RECT  73.76 65.345 73.55 65.14 ;
      RECT  73.97 66.055 73.76 65.725 ;
      RECT  71.93 66.055 71.75 65.14 ;
      RECT  73.37 66.055 73.19 65.14 ;
      POLYGON  70.925 66.055 70.925 65.725 71.36 65.725 71.36 65.345 70.925 65.345 70.925 65.14 70.85 65.14 70.85 66.055 70.925 66.055 ;
      RECT  72.65 65.14 72.47 63.435 ;
      RECT  70.925 65.93 70.85 67.635 ;
      RECT  70.85 65.345 70.64 65.725 ;
      RECT  73.01 65.015 72.83 65.93 ;
      POLYGON  71.36 66.02 71.36 66.43 71.185 66.43 71.105 66.35 71.105 66.02 71.36 66.02 ;
      RECT  73.37 65.93 73.19 67.635 ;
      RECT  73.01 65.93 72.83 67.635 ;
      RECT  73.76 65.93 73.55 67.635 ;
      RECT  73.97 65.725 73.76 65.93 ;
      RECT  73.97 65.93 73.76 67.635 ;
      RECT  70.85 65.93 70.64 67.635 ;
      POLYGON  71.36 67.01 71.36 67.42 71.105 67.42 71.105 67.09 71.185 67.01 71.36 67.01 ;
      RECT  73.76 65.345 73.55 65.725 ;
      RECT  70.85 65.015 70.64 65.345 ;
      RECT  72.65 65.015 72.47 65.93 ;
      RECT  71.01 66.515 70.925 66.925 ;
      RECT  71.93 65.93 71.75 67.635 ;
      RECT  71.57 67.01 71.36 67.42 ;
      RECT  73.76 65.015 73.55 65.345 ;
      RECT  71.57 66.02 71.36 66.43 ;
      RECT  71.57 65.345 71.36 65.725 ;
      RECT  73.97 65.345 73.76 65.725 ;
      RECT  72.29 65.015 72.11 65.93 ;
      RECT  72.29 65.93 72.11 67.635 ;
      RECT  70.85 65.725 70.64 65.93 ;
      RECT  73.76 65.725 73.55 65.93 ;
      RECT  73.97 65.015 73.76 65.345 ;
      RECT  71.93 65.015 71.75 65.93 ;
      RECT  73.37 65.015 73.19 65.93 ;
      POLYGON  70.925 65.015 70.925 65.345 71.36 65.345 71.36 65.725 70.925 65.725 70.925 65.93 70.85 65.93 70.85 65.015 70.925 65.015 ;
      RECT  72.65 65.93 72.47 67.635 ;
      RECT  70.925 69.09 70.85 67.385 ;
      RECT  70.85 69.675 70.64 69.295 ;
      RECT  73.01 70.005 72.83 69.09 ;
      POLYGON  71.36 69.0 71.36 68.59 71.185 68.59 71.105 68.67 71.105 69.0 71.36 69.0 ;
      RECT  73.37 69.09 73.19 67.385 ;
      RECT  73.01 69.09 72.83 67.385 ;
      RECT  73.76 69.09 73.55 67.385 ;
      RECT  73.97 69.295 73.76 69.09 ;
      RECT  73.97 69.09 73.76 67.385 ;
      RECT  70.85 69.09 70.64 67.385 ;
      POLYGON  71.36 68.01 71.36 67.6 71.105 67.6 71.105 67.93 71.185 68.01 71.36 68.01 ;
      RECT  73.76 69.675 73.55 69.295 ;
      RECT  70.85 70.005 70.64 69.675 ;
      RECT  72.65 70.005 72.47 69.09 ;
      RECT  71.01 68.505 70.925 68.095 ;
      RECT  71.93 69.09 71.75 67.385 ;
      RECT  71.57 68.01 71.36 67.6 ;
      RECT  73.76 70.005 73.55 69.675 ;
      RECT  71.57 69.0 71.36 68.59 ;
      RECT  71.57 69.675 71.36 69.295 ;
      RECT  73.97 69.675 73.76 69.295 ;
      RECT  72.29 70.005 72.11 69.09 ;
      RECT  72.29 69.09 72.11 67.385 ;
      RECT  70.85 69.295 70.64 69.09 ;
      RECT  73.76 69.295 73.55 69.09 ;
      RECT  73.97 70.005 73.76 69.675 ;
      RECT  71.93 70.005 71.75 69.09 ;
      RECT  73.37 70.005 73.19 69.09 ;
      POLYGON  70.925 70.005 70.925 69.675 71.36 69.675 71.36 69.295 70.925 69.295 70.925 69.09 70.85 69.09 70.85 70.005 70.925 70.005 ;
      RECT  72.65 69.09 72.47 67.385 ;
      RECT  70.925 69.88 70.85 71.585 ;
      RECT  70.85 69.295 70.64 69.675 ;
      RECT  73.01 68.965 72.83 69.88 ;
      POLYGON  71.36 69.97 71.36 70.38 71.185 70.38 71.105 70.3 71.105 69.97 71.36 69.97 ;
      RECT  73.37 69.88 73.19 71.585 ;
      RECT  73.01 69.88 72.83 71.585 ;
      RECT  73.76 69.88 73.55 71.585 ;
      RECT  73.97 69.675 73.76 69.88 ;
      RECT  73.97 69.88 73.76 71.585 ;
      RECT  70.85 69.88 70.64 71.585 ;
      POLYGON  71.36 70.96 71.36 71.37 71.105 71.37 71.105 71.04 71.185 70.96 71.36 70.96 ;
      RECT  73.76 69.295 73.55 69.675 ;
      RECT  70.85 68.965 70.64 69.295 ;
      RECT  72.65 68.965 72.47 69.88 ;
      RECT  71.01 70.465 70.925 70.875 ;
      RECT  71.93 69.88 71.75 71.585 ;
      RECT  71.57 70.96 71.36 71.37 ;
      RECT  73.76 68.965 73.55 69.295 ;
      RECT  71.57 69.97 71.36 70.38 ;
      RECT  71.57 69.295 71.36 69.675 ;
      RECT  73.97 69.295 73.76 69.675 ;
      RECT  72.29 68.965 72.11 69.88 ;
      RECT  72.29 69.88 72.11 71.585 ;
      RECT  70.85 69.675 70.64 69.88 ;
      RECT  73.76 69.675 73.55 69.88 ;
      RECT  73.97 68.965 73.76 69.295 ;
      RECT  71.93 68.965 71.75 69.88 ;
      RECT  73.37 68.965 73.19 69.88 ;
      POLYGON  70.925 68.965 70.925 69.295 71.36 69.295 71.36 69.675 70.925 69.675 70.925 69.88 70.85 69.88 70.85 68.965 70.925 68.965 ;
      RECT  72.65 69.88 72.47 71.585 ;
      RECT  70.925 73.04 70.85 71.335 ;
      RECT  70.85 73.625 70.64 73.245 ;
      RECT  73.01 73.955 72.83 73.04 ;
      POLYGON  71.36 72.95 71.36 72.54 71.185 72.54 71.105 72.62 71.105 72.95 71.36 72.95 ;
      RECT  73.37 73.04 73.19 71.335 ;
      RECT  73.01 73.04 72.83 71.335 ;
      RECT  73.76 73.04 73.55 71.335 ;
      RECT  73.97 73.245 73.76 73.04 ;
      RECT  73.97 73.04 73.76 71.335 ;
      RECT  70.85 73.04 70.64 71.335 ;
      POLYGON  71.36 71.96 71.36 71.55 71.105 71.55 71.105 71.88 71.185 71.96 71.36 71.96 ;
      RECT  73.76 73.625 73.55 73.245 ;
      RECT  70.85 73.955 70.64 73.625 ;
      RECT  72.65 73.955 72.47 73.04 ;
      RECT  71.01 72.455 70.925 72.045 ;
      RECT  71.93 73.04 71.75 71.335 ;
      RECT  71.57 71.96 71.36 71.55 ;
      RECT  73.76 73.955 73.55 73.625 ;
      RECT  71.57 72.95 71.36 72.54 ;
      RECT  71.57 73.625 71.36 73.245 ;
      RECT  73.97 73.625 73.76 73.245 ;
      RECT  72.29 73.955 72.11 73.04 ;
      RECT  72.29 73.04 72.11 71.335 ;
      RECT  70.85 73.245 70.64 73.04 ;
      RECT  73.76 73.245 73.55 73.04 ;
      RECT  73.97 73.955 73.76 73.625 ;
      RECT  71.93 73.955 71.75 73.04 ;
      RECT  73.37 73.955 73.19 73.04 ;
      POLYGON  70.925 73.955 70.925 73.625 71.36 73.625 71.36 73.245 70.925 73.245 70.925 73.04 70.85 73.04 70.85 73.955 70.925 73.955 ;
      RECT  72.65 73.04 72.47 71.335 ;
      RECT  70.925 73.83 70.85 75.535 ;
      RECT  70.85 73.245 70.64 73.625 ;
      RECT  73.01 72.915 72.83 73.83 ;
      POLYGON  71.36 73.92 71.36 74.33 71.185 74.33 71.105 74.25 71.105 73.92 71.36 73.92 ;
      RECT  73.37 73.83 73.19 75.535 ;
      RECT  73.01 73.83 72.83 75.535 ;
      RECT  73.76 73.83 73.55 75.535 ;
      RECT  73.97 73.625 73.76 73.83 ;
      RECT  73.97 73.83 73.76 75.535 ;
      RECT  70.85 73.83 70.64 75.535 ;
      POLYGON  71.36 74.91 71.36 75.32 71.105 75.32 71.105 74.99 71.185 74.91 71.36 74.91 ;
      RECT  73.76 73.245 73.55 73.625 ;
      RECT  70.85 72.915 70.64 73.245 ;
      RECT  72.65 72.915 72.47 73.83 ;
      RECT  71.01 74.415 70.925 74.825 ;
      RECT  71.93 73.83 71.75 75.535 ;
      RECT  71.57 74.91 71.36 75.32 ;
      RECT  73.76 72.915 73.55 73.245 ;
      RECT  71.57 73.92 71.36 74.33 ;
      RECT  71.57 73.245 71.36 73.625 ;
      RECT  73.97 73.245 73.76 73.625 ;
      RECT  72.29 72.915 72.11 73.83 ;
      RECT  72.29 73.83 72.11 75.535 ;
      RECT  70.85 73.625 70.64 73.83 ;
      RECT  73.76 73.625 73.55 73.83 ;
      RECT  73.97 72.915 73.76 73.245 ;
      RECT  71.93 72.915 71.75 73.83 ;
      RECT  73.37 72.915 73.19 73.83 ;
      POLYGON  70.925 72.915 70.925 73.245 71.36 73.245 71.36 73.625 70.925 73.625 70.925 73.83 70.85 73.83 70.85 72.915 70.925 72.915 ;
      RECT  72.65 73.83 72.47 75.535 ;
      RECT  70.925 76.99 70.85 75.285 ;
      RECT  70.85 77.575 70.64 77.195 ;
      RECT  73.01 77.905 72.83 76.99 ;
      POLYGON  71.36 76.9 71.36 76.49 71.185 76.49 71.105 76.57 71.105 76.9 71.36 76.9 ;
      RECT  73.37 76.99 73.19 75.285 ;
      RECT  73.01 76.99 72.83 75.285 ;
      RECT  73.76 76.99 73.55 75.285 ;
      RECT  73.97 77.195 73.76 76.99 ;
      RECT  73.97 76.99 73.76 75.285 ;
      RECT  70.85 76.99 70.64 75.285 ;
      POLYGON  71.36 75.91 71.36 75.5 71.105 75.5 71.105 75.83 71.185 75.91 71.36 75.91 ;
      RECT  73.76 77.575 73.55 77.195 ;
      RECT  70.85 77.905 70.64 77.575 ;
      RECT  72.65 77.905 72.47 76.99 ;
      RECT  71.01 76.405 70.925 75.995 ;
      RECT  71.93 76.99 71.75 75.285 ;
      RECT  71.57 75.91 71.36 75.5 ;
      RECT  73.76 77.905 73.55 77.575 ;
      RECT  71.57 76.9 71.36 76.49 ;
      RECT  71.57 77.575 71.36 77.195 ;
      RECT  73.97 77.575 73.76 77.195 ;
      RECT  72.29 77.905 72.11 76.99 ;
      RECT  72.29 76.99 72.11 75.285 ;
      RECT  70.85 77.195 70.64 76.99 ;
      RECT  73.76 77.195 73.55 76.99 ;
      RECT  73.97 77.905 73.76 77.575 ;
      RECT  71.93 77.905 71.75 76.99 ;
      RECT  73.37 77.905 73.19 76.99 ;
      POLYGON  70.925 77.905 70.925 77.575 71.36 77.575 71.36 77.195 70.925 77.195 70.925 76.99 70.85 76.99 70.85 77.905 70.925 77.905 ;
      RECT  72.65 76.99 72.47 75.285 ;
      RECT  70.925 77.78 70.85 79.485 ;
      RECT  70.85 77.195 70.64 77.575 ;
      RECT  73.01 76.865 72.83 77.78 ;
      POLYGON  71.36 77.87 71.36 78.28 71.185 78.28 71.105 78.2 71.105 77.87 71.36 77.87 ;
      RECT  73.37 77.78 73.19 79.485 ;
      RECT  73.01 77.78 72.83 79.485 ;
      RECT  73.76 77.78 73.55 79.485 ;
      RECT  73.97 77.575 73.76 77.78 ;
      RECT  73.97 77.78 73.76 79.485 ;
      RECT  70.85 77.78 70.64 79.485 ;
      POLYGON  71.36 78.86 71.36 79.27 71.105 79.27 71.105 78.94 71.185 78.86 71.36 78.86 ;
      RECT  73.76 77.195 73.55 77.575 ;
      RECT  70.85 76.865 70.64 77.195 ;
      RECT  72.65 76.865 72.47 77.78 ;
      RECT  71.01 78.365 70.925 78.775 ;
      RECT  71.93 77.78 71.75 79.485 ;
      RECT  71.57 78.86 71.36 79.27 ;
      RECT  73.76 76.865 73.55 77.195 ;
      RECT  71.57 77.87 71.36 78.28 ;
      RECT  71.57 77.195 71.36 77.575 ;
      RECT  73.97 77.195 73.76 77.575 ;
      RECT  72.29 76.865 72.11 77.78 ;
      RECT  72.29 77.78 72.11 79.485 ;
      RECT  70.85 77.575 70.64 77.78 ;
      RECT  73.76 77.575 73.55 77.78 ;
      RECT  73.97 76.865 73.76 77.195 ;
      RECT  71.93 76.865 71.75 77.78 ;
      RECT  73.37 76.865 73.19 77.78 ;
      POLYGON  70.925 76.865 70.925 77.195 71.36 77.195 71.36 77.575 70.925 77.575 70.925 77.78 70.85 77.78 70.85 76.865 70.925 76.865 ;
      RECT  72.65 77.78 72.47 79.485 ;
      RECT  70.925 80.94 70.85 79.235 ;
      RECT  70.85 81.525 70.64 81.145 ;
      RECT  73.01 81.855 72.83 80.94 ;
      POLYGON  71.36 80.85 71.36 80.44 71.185 80.44 71.105 80.52 71.105 80.85 71.36 80.85 ;
      RECT  73.37 80.94 73.19 79.235 ;
      RECT  73.01 80.94 72.83 79.235 ;
      RECT  73.76 80.94 73.55 79.235 ;
      RECT  73.97 81.145 73.76 80.94 ;
      RECT  73.97 80.94 73.76 79.235 ;
      RECT  70.85 80.94 70.64 79.235 ;
      POLYGON  71.36 79.86 71.36 79.45 71.105 79.45 71.105 79.78 71.185 79.86 71.36 79.86 ;
      RECT  73.76 81.525 73.55 81.145 ;
      RECT  70.85 81.855 70.64 81.525 ;
      RECT  72.65 81.855 72.47 80.94 ;
      RECT  71.01 80.355 70.925 79.945 ;
      RECT  71.93 80.94 71.75 79.235 ;
      RECT  71.57 79.86 71.36 79.45 ;
      RECT  73.76 81.855 73.55 81.525 ;
      RECT  71.57 80.85 71.36 80.44 ;
      RECT  71.57 81.525 71.36 81.145 ;
      RECT  73.97 81.525 73.76 81.145 ;
      RECT  72.29 81.855 72.11 80.94 ;
      RECT  72.29 80.94 72.11 79.235 ;
      RECT  70.85 81.145 70.64 80.94 ;
      RECT  73.76 81.145 73.55 80.94 ;
      RECT  73.97 81.855 73.76 81.525 ;
      RECT  71.93 81.855 71.75 80.94 ;
      RECT  73.37 81.855 73.19 80.94 ;
      POLYGON  70.925 81.855 70.925 81.525 71.36 81.525 71.36 81.145 70.925 81.145 70.925 80.94 70.85 80.94 70.85 81.855 70.925 81.855 ;
      RECT  72.65 80.94 72.47 79.235 ;
      RECT  70.925 81.73 70.85 83.435 ;
      RECT  70.85 81.145 70.64 81.525 ;
      RECT  73.01 80.815 72.83 81.73 ;
      POLYGON  71.36 81.82 71.36 82.23 71.185 82.23 71.105 82.15 71.105 81.82 71.36 81.82 ;
      RECT  73.37 81.73 73.19 83.435 ;
      RECT  73.01 81.73 72.83 83.435 ;
      RECT  73.76 81.73 73.55 83.435 ;
      RECT  73.97 81.525 73.76 81.73 ;
      RECT  73.97 81.73 73.76 83.435 ;
      RECT  70.85 81.73 70.64 83.435 ;
      POLYGON  71.36 82.81 71.36 83.22 71.105 83.22 71.105 82.89 71.185 82.81 71.36 82.81 ;
      RECT  73.76 81.145 73.55 81.525 ;
      RECT  70.85 80.815 70.64 81.145 ;
      RECT  72.65 80.815 72.47 81.73 ;
      RECT  71.01 82.315 70.925 82.725 ;
      RECT  71.93 81.73 71.75 83.435 ;
      RECT  71.57 82.81 71.36 83.22 ;
      RECT  73.76 80.815 73.55 81.145 ;
      RECT  71.57 81.82 71.36 82.23 ;
      RECT  71.57 81.145 71.36 81.525 ;
      RECT  73.97 81.145 73.76 81.525 ;
      RECT  72.29 80.815 72.11 81.73 ;
      RECT  72.29 81.73 72.11 83.435 ;
      RECT  70.85 81.525 70.64 81.73 ;
      RECT  73.76 81.525 73.55 81.73 ;
      RECT  73.97 80.815 73.76 81.145 ;
      RECT  71.93 80.815 71.75 81.73 ;
      RECT  73.37 80.815 73.19 81.73 ;
      POLYGON  70.925 80.815 70.925 81.145 71.36 81.145 71.36 81.525 70.925 81.525 70.925 81.73 70.85 81.73 70.85 80.815 70.925 80.815 ;
      RECT  72.65 81.73 72.47 83.435 ;
      RECT  70.925 84.89 70.85 83.185 ;
      RECT  70.85 85.475 70.64 85.095 ;
      RECT  73.01 85.805 72.83 84.89 ;
      POLYGON  71.36 84.8 71.36 84.39 71.185 84.39 71.105 84.47 71.105 84.8 71.36 84.8 ;
      RECT  73.37 84.89 73.19 83.185 ;
      RECT  73.01 84.89 72.83 83.185 ;
      RECT  73.76 84.89 73.55 83.185 ;
      RECT  73.97 85.095 73.76 84.89 ;
      RECT  73.97 84.89 73.76 83.185 ;
      RECT  70.85 84.89 70.64 83.185 ;
      POLYGON  71.36 83.81 71.36 83.4 71.105 83.4 71.105 83.73 71.185 83.81 71.36 83.81 ;
      RECT  73.76 85.475 73.55 85.095 ;
      RECT  70.85 85.805 70.64 85.475 ;
      RECT  72.65 85.805 72.47 84.89 ;
      RECT  71.01 84.305 70.925 83.895 ;
      RECT  71.93 84.89 71.75 83.185 ;
      RECT  71.57 83.81 71.36 83.4 ;
      RECT  73.76 85.805 73.55 85.475 ;
      RECT  71.57 84.8 71.36 84.39 ;
      RECT  71.57 85.475 71.36 85.095 ;
      RECT  73.97 85.475 73.76 85.095 ;
      RECT  72.29 85.805 72.11 84.89 ;
      RECT  72.29 84.89 72.11 83.185 ;
      RECT  70.85 85.095 70.64 84.89 ;
      RECT  73.76 85.095 73.55 84.89 ;
      RECT  73.97 85.805 73.76 85.475 ;
      RECT  71.93 85.805 71.75 84.89 ;
      RECT  73.37 85.805 73.19 84.89 ;
      POLYGON  70.925 85.805 70.925 85.475 71.36 85.475 71.36 85.095 70.925 85.095 70.925 84.89 70.85 84.89 70.85 85.805 70.925 85.805 ;
      RECT  72.65 84.89 72.47 83.185 ;
      RECT  70.925 85.68 70.85 87.385 ;
      RECT  70.85 85.095 70.64 85.475 ;
      RECT  73.01 84.765 72.83 85.68 ;
      POLYGON  71.36 85.77 71.36 86.18 71.185 86.18 71.105 86.1 71.105 85.77 71.36 85.77 ;
      RECT  73.37 85.68 73.19 87.385 ;
      RECT  73.01 85.68 72.83 87.385 ;
      RECT  73.76 85.68 73.55 87.385 ;
      RECT  73.97 85.475 73.76 85.68 ;
      RECT  73.97 85.68 73.76 87.385 ;
      RECT  70.85 85.68 70.64 87.385 ;
      POLYGON  71.36 86.76 71.36 87.17 71.105 87.17 71.105 86.84 71.185 86.76 71.36 86.76 ;
      RECT  73.76 85.095 73.55 85.475 ;
      RECT  70.85 84.765 70.64 85.095 ;
      RECT  72.65 84.765 72.47 85.68 ;
      RECT  71.01 86.265 70.925 86.675 ;
      RECT  71.93 85.68 71.75 87.385 ;
      RECT  71.57 86.76 71.36 87.17 ;
      RECT  73.76 84.765 73.55 85.095 ;
      RECT  71.57 85.77 71.36 86.18 ;
      RECT  71.57 85.095 71.36 85.475 ;
      RECT  73.97 85.095 73.76 85.475 ;
      RECT  72.29 84.765 72.11 85.68 ;
      RECT  72.29 85.68 72.11 87.385 ;
      RECT  70.85 85.475 70.64 85.68 ;
      RECT  73.76 85.475 73.55 85.68 ;
      RECT  73.97 84.765 73.76 85.095 ;
      RECT  71.93 84.765 71.75 85.68 ;
      RECT  73.37 84.765 73.19 85.68 ;
      POLYGON  70.925 84.765 70.925 85.095 71.36 85.095 71.36 85.475 70.925 85.475 70.925 85.68 70.85 85.68 70.85 84.765 70.925 84.765 ;
      RECT  72.65 85.68 72.47 87.385 ;
      RECT  70.925 88.84 70.85 87.135 ;
      RECT  70.85 89.425 70.64 89.045 ;
      RECT  73.01 89.755 72.83 88.84 ;
      POLYGON  71.36 88.75 71.36 88.34 71.185 88.34 71.105 88.42 71.105 88.75 71.36 88.75 ;
      RECT  73.37 88.84 73.19 87.135 ;
      RECT  73.01 88.84 72.83 87.135 ;
      RECT  73.76 88.84 73.55 87.135 ;
      RECT  73.97 89.045 73.76 88.84 ;
      RECT  73.97 88.84 73.76 87.135 ;
      RECT  70.85 88.84 70.64 87.135 ;
      POLYGON  71.36 87.76 71.36 87.35 71.105 87.35 71.105 87.68 71.185 87.76 71.36 87.76 ;
      RECT  73.76 89.425 73.55 89.045 ;
      RECT  70.85 89.755 70.64 89.425 ;
      RECT  72.65 89.755 72.47 88.84 ;
      RECT  71.01 88.255 70.925 87.845 ;
      RECT  71.93 88.84 71.75 87.135 ;
      RECT  71.57 87.76 71.36 87.35 ;
      RECT  73.76 89.755 73.55 89.425 ;
      RECT  71.57 88.75 71.36 88.34 ;
      RECT  71.57 89.425 71.36 89.045 ;
      RECT  73.97 89.425 73.76 89.045 ;
      RECT  72.29 89.755 72.11 88.84 ;
      RECT  72.29 88.84 72.11 87.135 ;
      RECT  70.85 89.045 70.64 88.84 ;
      RECT  73.76 89.045 73.55 88.84 ;
      RECT  73.97 89.755 73.76 89.425 ;
      RECT  71.93 89.755 71.75 88.84 ;
      RECT  73.37 89.755 73.19 88.84 ;
      POLYGON  70.925 89.755 70.925 89.425 71.36 89.425 71.36 89.045 70.925 89.045 70.925 88.84 70.85 88.84 70.85 89.755 70.925 89.755 ;
      RECT  72.65 88.84 72.47 87.135 ;
      RECT  70.925 89.63 70.85 91.335 ;
      RECT  70.85 89.045 70.64 89.425 ;
      RECT  73.01 88.715 72.83 89.63 ;
      POLYGON  71.36 89.72 71.36 90.13 71.185 90.13 71.105 90.05 71.105 89.72 71.36 89.72 ;
      RECT  73.37 89.63 73.19 91.335 ;
      RECT  73.01 89.63 72.83 91.335 ;
      RECT  73.76 89.63 73.55 91.335 ;
      RECT  73.97 89.425 73.76 89.63 ;
      RECT  73.97 89.63 73.76 91.335 ;
      RECT  70.85 89.63 70.64 91.335 ;
      POLYGON  71.36 90.71 71.36 91.12 71.105 91.12 71.105 90.79 71.185 90.71 71.36 90.71 ;
      RECT  73.76 89.045 73.55 89.425 ;
      RECT  70.85 88.715 70.64 89.045 ;
      RECT  72.65 88.715 72.47 89.63 ;
      RECT  71.01 90.215 70.925 90.625 ;
      RECT  71.93 89.63 71.75 91.335 ;
      RECT  71.57 90.71 71.36 91.12 ;
      RECT  73.76 88.715 73.55 89.045 ;
      RECT  71.57 89.72 71.36 90.13 ;
      RECT  71.57 89.045 71.36 89.425 ;
      RECT  73.97 89.045 73.76 89.425 ;
      RECT  72.29 88.715 72.11 89.63 ;
      RECT  72.29 89.63 72.11 91.335 ;
      RECT  70.85 89.425 70.64 89.63 ;
      RECT  73.76 89.425 73.55 89.63 ;
      RECT  73.97 88.715 73.76 89.045 ;
      RECT  71.93 88.715 71.75 89.63 ;
      RECT  73.37 88.715 73.19 89.63 ;
      POLYGON  70.925 88.715 70.925 89.045 71.36 89.045 71.36 89.425 70.925 89.425 70.925 89.63 70.85 89.63 70.85 88.715 70.925 88.715 ;
      RECT  72.65 89.63 72.47 91.335 ;
      RECT  70.925 92.79 70.85 91.085 ;
      RECT  70.85 93.375 70.64 92.995 ;
      RECT  73.01 93.705 72.83 92.79 ;
      POLYGON  71.36 92.7 71.36 92.29 71.185 92.29 71.105 92.37 71.105 92.7 71.36 92.7 ;
      RECT  73.37 92.79 73.19 91.085 ;
      RECT  73.01 92.79 72.83 91.085 ;
      RECT  73.76 92.79 73.55 91.085 ;
      RECT  73.97 92.995 73.76 92.79 ;
      RECT  73.97 92.79 73.76 91.085 ;
      RECT  70.85 92.79 70.64 91.085 ;
      POLYGON  71.36 91.71 71.36 91.3 71.105 91.3 71.105 91.63 71.185 91.71 71.36 91.71 ;
      RECT  73.76 93.375 73.55 92.995 ;
      RECT  70.85 93.705 70.64 93.375 ;
      RECT  72.65 93.705 72.47 92.79 ;
      RECT  71.01 92.205 70.925 91.795 ;
      RECT  71.93 92.79 71.75 91.085 ;
      RECT  71.57 91.71 71.36 91.3 ;
      RECT  73.76 93.705 73.55 93.375 ;
      RECT  71.57 92.7 71.36 92.29 ;
      RECT  71.57 93.375 71.36 92.995 ;
      RECT  73.97 93.375 73.76 92.995 ;
      RECT  72.29 93.705 72.11 92.79 ;
      RECT  72.29 92.79 72.11 91.085 ;
      RECT  70.85 92.995 70.64 92.79 ;
      RECT  73.76 92.995 73.55 92.79 ;
      RECT  73.97 93.705 73.76 93.375 ;
      RECT  71.93 93.705 71.75 92.79 ;
      RECT  73.37 93.705 73.19 92.79 ;
      POLYGON  70.925 93.705 70.925 93.375 71.36 93.375 71.36 92.995 70.925 92.995 70.925 92.79 70.85 92.79 70.85 93.705 70.925 93.705 ;
      RECT  72.65 92.79 72.47 91.085 ;
      RECT  70.925 93.58 70.85 95.285 ;
      RECT  70.85 92.995 70.64 93.375 ;
      RECT  73.01 92.665 72.83 93.58 ;
      POLYGON  71.36 93.67 71.36 94.08 71.185 94.08 71.105 94.0 71.105 93.67 71.36 93.67 ;
      RECT  73.37 93.58 73.19 95.285 ;
      RECT  73.01 93.58 72.83 95.285 ;
      RECT  73.76 93.58 73.55 95.285 ;
      RECT  73.97 93.375 73.76 93.58 ;
      RECT  73.97 93.58 73.76 95.285 ;
      RECT  70.85 93.58 70.64 95.285 ;
      POLYGON  71.36 94.66 71.36 95.07 71.105 95.07 71.105 94.74 71.185 94.66 71.36 94.66 ;
      RECT  73.76 92.995 73.55 93.375 ;
      RECT  70.85 92.665 70.64 92.995 ;
      RECT  72.65 92.665 72.47 93.58 ;
      RECT  71.01 94.165 70.925 94.575 ;
      RECT  71.93 93.58 71.75 95.285 ;
      RECT  71.57 94.66 71.36 95.07 ;
      RECT  73.76 92.665 73.55 92.995 ;
      RECT  71.57 93.67 71.36 94.08 ;
      RECT  71.57 92.995 71.36 93.375 ;
      RECT  73.97 92.995 73.76 93.375 ;
      RECT  72.29 92.665 72.11 93.58 ;
      RECT  72.29 93.58 72.11 95.285 ;
      RECT  70.85 93.375 70.64 93.58 ;
      RECT  73.76 93.375 73.55 93.58 ;
      RECT  73.97 92.665 73.76 92.995 ;
      RECT  71.93 92.665 71.75 93.58 ;
      RECT  73.37 92.665 73.19 93.58 ;
      POLYGON  70.925 92.665 70.925 92.995 71.36 92.995 71.36 93.375 70.925 93.375 70.925 93.58 70.85 93.58 70.85 92.665 70.925 92.665 ;
      RECT  72.65 93.58 72.47 95.285 ;
      RECT  72.65 96.345 72.47 94.765 ;
      RECT  73.01 96.345 72.83 94.765 ;
      RECT  72.56 96.345 72.43 95.635 ;
      RECT  72.29 96.345 72.11 94.765 ;
      RECT  72.69 96.345 72.56 95.635 ;
      RECT  73.01 97.135 72.83 96.345 ;
      RECT  73.37 97.135 73.19 96.345 ;
      RECT  71.93 97.135 71.75 96.345 ;
      RECT  72.65 97.135 72.47 96.345 ;
      RECT  72.29 97.135 72.11 96.345 ;
      RECT  73.37 96.345 73.19 94.765 ;
      RECT  71.93 96.345 71.75 94.765 ;
      RECT  72.47 91.085 72.65 92.79 ;
      RECT  72.47 93.58 72.65 95.285 ;
      RECT  72.47 71.335 72.65 73.04 ;
      RECT  72.47 75.285 72.65 76.99 ;
      RECT  72.47 85.68 72.65 87.385 ;
      RECT  72.47 67.385 72.65 69.09 ;
      RECT  72.47 73.83 72.65 75.535 ;
      RECT  72.47 81.73 72.65 83.435 ;
      RECT  72.47 63.435 72.65 65.14 ;
      RECT  72.47 65.93 72.65 67.635 ;
      RECT  72.47 83.185 72.65 84.89 ;
      RECT  72.47 87.135 72.65 88.84 ;
      RECT  72.47 69.88 72.65 71.585 ;
      RECT  72.47 61.98 72.65 63.685 ;
      RECT  72.47 77.78 72.65 79.485 ;
      RECT  72.47 79.235 72.65 80.94 ;
      RECT  72.47 89.63 72.65 91.335 ;
      RECT  72.47 59.485 72.65 61.19 ;
      RECT  81.11 58.425 81.29 60.005 ;
      RECT  80.75 58.425 80.93 60.005 ;
      RECT  81.2 58.425 81.33 59.135 ;
      RECT  81.47 58.425 81.65 60.005 ;
      RECT  81.07 58.425 81.2 59.135 ;
      RECT  80.75 57.635 80.93 58.425 ;
      RECT  80.39 57.635 80.57 58.425 ;
      RECT  81.83 57.635 82.01 58.425 ;
      RECT  81.11 57.635 81.29 58.425 ;
      RECT  81.47 57.635 81.65 58.425 ;
      RECT  80.39 58.425 80.57 60.005 ;
      RECT  81.83 58.425 82.01 60.005 ;
      RECT  82.835 61.19 82.91 59.485 ;
      RECT  82.91 61.775 83.12 61.395 ;
      RECT  80.75 62.105 80.93 61.19 ;
      POLYGON  82.4 61.1 82.4 60.69 82.575 60.69 82.655 60.77 82.655 61.1 82.4 61.1 ;
      RECT  80.39 61.19 80.57 59.485 ;
      RECT  80.75 61.19 80.93 59.485 ;
      RECT  80.0 61.19 80.21 59.485 ;
      RECT  79.79 61.395 80.0 61.19 ;
      RECT  79.79 61.19 80.0 59.485 ;
      RECT  82.91 61.19 83.12 59.485 ;
      POLYGON  82.4 60.11 82.4 59.7 82.655 59.7 82.655 60.03 82.575 60.11 82.4 60.11 ;
      RECT  80.0 61.775 80.21 61.395 ;
      RECT  82.91 62.105 83.12 61.775 ;
      RECT  81.11 62.105 81.29 61.19 ;
      RECT  82.75 60.605 82.835 60.195 ;
      RECT  81.83 61.19 82.01 59.485 ;
      RECT  82.19 60.11 82.4 59.7 ;
      RECT  80.0 62.105 80.21 61.775 ;
      RECT  82.19 61.1 82.4 60.69 ;
      RECT  82.19 61.775 82.4 61.395 ;
      RECT  79.79 61.775 80.0 61.395 ;
      RECT  81.47 62.105 81.65 61.19 ;
      RECT  81.47 61.19 81.65 59.485 ;
      RECT  82.91 61.395 83.12 61.19 ;
      RECT  80.0 61.395 80.21 61.19 ;
      RECT  79.79 62.105 80.0 61.775 ;
      RECT  81.83 62.105 82.01 61.19 ;
      RECT  80.39 62.105 80.57 61.19 ;
      POLYGON  82.835 62.105 82.835 61.775 82.4 61.775 82.4 61.395 82.835 61.395 82.835 61.19 82.91 61.19 82.91 62.105 82.835 62.105 ;
      RECT  81.11 61.19 81.29 59.485 ;
      RECT  82.835 61.98 82.91 63.685 ;
      RECT  82.91 61.395 83.12 61.775 ;
      RECT  80.75 61.065 80.93 61.98 ;
      POLYGON  82.4 62.07 82.4 62.48 82.575 62.48 82.655 62.4 82.655 62.07 82.4 62.07 ;
      RECT  80.39 61.98 80.57 63.685 ;
      RECT  80.75 61.98 80.93 63.685 ;
      RECT  80.0 61.98 80.21 63.685 ;
      RECT  79.79 61.775 80.0 61.98 ;
      RECT  79.79 61.98 80.0 63.685 ;
      RECT  82.91 61.98 83.12 63.685 ;
      POLYGON  82.4 63.06 82.4 63.47 82.655 63.47 82.655 63.14 82.575 63.06 82.4 63.06 ;
      RECT  80.0 61.395 80.21 61.775 ;
      RECT  82.91 61.065 83.12 61.395 ;
      RECT  81.11 61.065 81.29 61.98 ;
      RECT  82.75 62.565 82.835 62.975 ;
      RECT  81.83 61.98 82.01 63.685 ;
      RECT  82.19 63.06 82.4 63.47 ;
      RECT  80.0 61.065 80.21 61.395 ;
      RECT  82.19 62.07 82.4 62.48 ;
      RECT  82.19 61.395 82.4 61.775 ;
      RECT  79.79 61.395 80.0 61.775 ;
      RECT  81.47 61.065 81.65 61.98 ;
      RECT  81.47 61.98 81.65 63.685 ;
      RECT  82.91 61.775 83.12 61.98 ;
      RECT  80.0 61.775 80.21 61.98 ;
      RECT  79.79 61.065 80.0 61.395 ;
      RECT  81.83 61.065 82.01 61.98 ;
      RECT  80.39 61.065 80.57 61.98 ;
      POLYGON  82.835 61.065 82.835 61.395 82.4 61.395 82.4 61.775 82.835 61.775 82.835 61.98 82.91 61.98 82.91 61.065 82.835 61.065 ;
      RECT  81.11 61.98 81.29 63.685 ;
      RECT  82.835 65.14 82.91 63.435 ;
      RECT  82.91 65.725 83.12 65.345 ;
      RECT  80.75 66.055 80.93 65.14 ;
      POLYGON  82.4 65.05 82.4 64.64 82.575 64.64 82.655 64.72 82.655 65.05 82.4 65.05 ;
      RECT  80.39 65.14 80.57 63.435 ;
      RECT  80.75 65.14 80.93 63.435 ;
      RECT  80.0 65.14 80.21 63.435 ;
      RECT  79.79 65.345 80.0 65.14 ;
      RECT  79.79 65.14 80.0 63.435 ;
      RECT  82.91 65.14 83.12 63.435 ;
      POLYGON  82.4 64.06 82.4 63.65 82.655 63.65 82.655 63.98 82.575 64.06 82.4 64.06 ;
      RECT  80.0 65.725 80.21 65.345 ;
      RECT  82.91 66.055 83.12 65.725 ;
      RECT  81.11 66.055 81.29 65.14 ;
      RECT  82.75 64.555 82.835 64.145 ;
      RECT  81.83 65.14 82.01 63.435 ;
      RECT  82.19 64.06 82.4 63.65 ;
      RECT  80.0 66.055 80.21 65.725 ;
      RECT  82.19 65.05 82.4 64.64 ;
      RECT  82.19 65.725 82.4 65.345 ;
      RECT  79.79 65.725 80.0 65.345 ;
      RECT  81.47 66.055 81.65 65.14 ;
      RECT  81.47 65.14 81.65 63.435 ;
      RECT  82.91 65.345 83.12 65.14 ;
      RECT  80.0 65.345 80.21 65.14 ;
      RECT  79.79 66.055 80.0 65.725 ;
      RECT  81.83 66.055 82.01 65.14 ;
      RECT  80.39 66.055 80.57 65.14 ;
      POLYGON  82.835 66.055 82.835 65.725 82.4 65.725 82.4 65.345 82.835 65.345 82.835 65.14 82.91 65.14 82.91 66.055 82.835 66.055 ;
      RECT  81.11 65.14 81.29 63.435 ;
      RECT  82.835 65.93 82.91 67.635 ;
      RECT  82.91 65.345 83.12 65.725 ;
      RECT  80.75 65.015 80.93 65.93 ;
      POLYGON  82.4 66.02 82.4 66.43 82.575 66.43 82.655 66.35 82.655 66.02 82.4 66.02 ;
      RECT  80.39 65.93 80.57 67.635 ;
      RECT  80.75 65.93 80.93 67.635 ;
      RECT  80.0 65.93 80.21 67.635 ;
      RECT  79.79 65.725 80.0 65.93 ;
      RECT  79.79 65.93 80.0 67.635 ;
      RECT  82.91 65.93 83.12 67.635 ;
      POLYGON  82.4 67.01 82.4 67.42 82.655 67.42 82.655 67.09 82.575 67.01 82.4 67.01 ;
      RECT  80.0 65.345 80.21 65.725 ;
      RECT  82.91 65.015 83.12 65.345 ;
      RECT  81.11 65.015 81.29 65.93 ;
      RECT  82.75 66.515 82.835 66.925 ;
      RECT  81.83 65.93 82.01 67.635 ;
      RECT  82.19 67.01 82.4 67.42 ;
      RECT  80.0 65.015 80.21 65.345 ;
      RECT  82.19 66.02 82.4 66.43 ;
      RECT  82.19 65.345 82.4 65.725 ;
      RECT  79.79 65.345 80.0 65.725 ;
      RECT  81.47 65.015 81.65 65.93 ;
      RECT  81.47 65.93 81.65 67.635 ;
      RECT  82.91 65.725 83.12 65.93 ;
      RECT  80.0 65.725 80.21 65.93 ;
      RECT  79.79 65.015 80.0 65.345 ;
      RECT  81.83 65.015 82.01 65.93 ;
      RECT  80.39 65.015 80.57 65.93 ;
      POLYGON  82.835 65.015 82.835 65.345 82.4 65.345 82.4 65.725 82.835 65.725 82.835 65.93 82.91 65.93 82.91 65.015 82.835 65.015 ;
      RECT  81.11 65.93 81.29 67.635 ;
      RECT  82.835 69.09 82.91 67.385 ;
      RECT  82.91 69.675 83.12 69.295 ;
      RECT  80.75 70.005 80.93 69.09 ;
      POLYGON  82.4 69.0 82.4 68.59 82.575 68.59 82.655 68.67 82.655 69.0 82.4 69.0 ;
      RECT  80.39 69.09 80.57 67.385 ;
      RECT  80.75 69.09 80.93 67.385 ;
      RECT  80.0 69.09 80.21 67.385 ;
      RECT  79.79 69.295 80.0 69.09 ;
      RECT  79.79 69.09 80.0 67.385 ;
      RECT  82.91 69.09 83.12 67.385 ;
      POLYGON  82.4 68.01 82.4 67.6 82.655 67.6 82.655 67.93 82.575 68.01 82.4 68.01 ;
      RECT  80.0 69.675 80.21 69.295 ;
      RECT  82.91 70.005 83.12 69.675 ;
      RECT  81.11 70.005 81.29 69.09 ;
      RECT  82.75 68.505 82.835 68.095 ;
      RECT  81.83 69.09 82.01 67.385 ;
      RECT  82.19 68.01 82.4 67.6 ;
      RECT  80.0 70.005 80.21 69.675 ;
      RECT  82.19 69.0 82.4 68.59 ;
      RECT  82.19 69.675 82.4 69.295 ;
      RECT  79.79 69.675 80.0 69.295 ;
      RECT  81.47 70.005 81.65 69.09 ;
      RECT  81.47 69.09 81.65 67.385 ;
      RECT  82.91 69.295 83.12 69.09 ;
      RECT  80.0 69.295 80.21 69.09 ;
      RECT  79.79 70.005 80.0 69.675 ;
      RECT  81.83 70.005 82.01 69.09 ;
      RECT  80.39 70.005 80.57 69.09 ;
      POLYGON  82.835 70.005 82.835 69.675 82.4 69.675 82.4 69.295 82.835 69.295 82.835 69.09 82.91 69.09 82.91 70.005 82.835 70.005 ;
      RECT  81.11 69.09 81.29 67.385 ;
      RECT  82.835 69.88 82.91 71.585 ;
      RECT  82.91 69.295 83.12 69.675 ;
      RECT  80.75 68.965 80.93 69.88 ;
      POLYGON  82.4 69.97 82.4 70.38 82.575 70.38 82.655 70.3 82.655 69.97 82.4 69.97 ;
      RECT  80.39 69.88 80.57 71.585 ;
      RECT  80.75 69.88 80.93 71.585 ;
      RECT  80.0 69.88 80.21 71.585 ;
      RECT  79.79 69.675 80.0 69.88 ;
      RECT  79.79 69.88 80.0 71.585 ;
      RECT  82.91 69.88 83.12 71.585 ;
      POLYGON  82.4 70.96 82.4 71.37 82.655 71.37 82.655 71.04 82.575 70.96 82.4 70.96 ;
      RECT  80.0 69.295 80.21 69.675 ;
      RECT  82.91 68.965 83.12 69.295 ;
      RECT  81.11 68.965 81.29 69.88 ;
      RECT  82.75 70.465 82.835 70.875 ;
      RECT  81.83 69.88 82.01 71.585 ;
      RECT  82.19 70.96 82.4 71.37 ;
      RECT  80.0 68.965 80.21 69.295 ;
      RECT  82.19 69.97 82.4 70.38 ;
      RECT  82.19 69.295 82.4 69.675 ;
      RECT  79.79 69.295 80.0 69.675 ;
      RECT  81.47 68.965 81.65 69.88 ;
      RECT  81.47 69.88 81.65 71.585 ;
      RECT  82.91 69.675 83.12 69.88 ;
      RECT  80.0 69.675 80.21 69.88 ;
      RECT  79.79 68.965 80.0 69.295 ;
      RECT  81.83 68.965 82.01 69.88 ;
      RECT  80.39 68.965 80.57 69.88 ;
      POLYGON  82.835 68.965 82.835 69.295 82.4 69.295 82.4 69.675 82.835 69.675 82.835 69.88 82.91 69.88 82.91 68.965 82.835 68.965 ;
      RECT  81.11 69.88 81.29 71.585 ;
      RECT  82.835 73.04 82.91 71.335 ;
      RECT  82.91 73.625 83.12 73.245 ;
      RECT  80.75 73.955 80.93 73.04 ;
      POLYGON  82.4 72.95 82.4 72.54 82.575 72.54 82.655 72.62 82.655 72.95 82.4 72.95 ;
      RECT  80.39 73.04 80.57 71.335 ;
      RECT  80.75 73.04 80.93 71.335 ;
      RECT  80.0 73.04 80.21 71.335 ;
      RECT  79.79 73.245 80.0 73.04 ;
      RECT  79.79 73.04 80.0 71.335 ;
      RECT  82.91 73.04 83.12 71.335 ;
      POLYGON  82.4 71.96 82.4 71.55 82.655 71.55 82.655 71.88 82.575 71.96 82.4 71.96 ;
      RECT  80.0 73.625 80.21 73.245 ;
      RECT  82.91 73.955 83.12 73.625 ;
      RECT  81.11 73.955 81.29 73.04 ;
      RECT  82.75 72.455 82.835 72.045 ;
      RECT  81.83 73.04 82.01 71.335 ;
      RECT  82.19 71.96 82.4 71.55 ;
      RECT  80.0 73.955 80.21 73.625 ;
      RECT  82.19 72.95 82.4 72.54 ;
      RECT  82.19 73.625 82.4 73.245 ;
      RECT  79.79 73.625 80.0 73.245 ;
      RECT  81.47 73.955 81.65 73.04 ;
      RECT  81.47 73.04 81.65 71.335 ;
      RECT  82.91 73.245 83.12 73.04 ;
      RECT  80.0 73.245 80.21 73.04 ;
      RECT  79.79 73.955 80.0 73.625 ;
      RECT  81.83 73.955 82.01 73.04 ;
      RECT  80.39 73.955 80.57 73.04 ;
      POLYGON  82.835 73.955 82.835 73.625 82.4 73.625 82.4 73.245 82.835 73.245 82.835 73.04 82.91 73.04 82.91 73.955 82.835 73.955 ;
      RECT  81.11 73.04 81.29 71.335 ;
      RECT  82.835 73.83 82.91 75.535 ;
      RECT  82.91 73.245 83.12 73.625 ;
      RECT  80.75 72.915 80.93 73.83 ;
      POLYGON  82.4 73.92 82.4 74.33 82.575 74.33 82.655 74.25 82.655 73.92 82.4 73.92 ;
      RECT  80.39 73.83 80.57 75.535 ;
      RECT  80.75 73.83 80.93 75.535 ;
      RECT  80.0 73.83 80.21 75.535 ;
      RECT  79.79 73.625 80.0 73.83 ;
      RECT  79.79 73.83 80.0 75.535 ;
      RECT  82.91 73.83 83.12 75.535 ;
      POLYGON  82.4 74.91 82.4 75.32 82.655 75.32 82.655 74.99 82.575 74.91 82.4 74.91 ;
      RECT  80.0 73.245 80.21 73.625 ;
      RECT  82.91 72.915 83.12 73.245 ;
      RECT  81.11 72.915 81.29 73.83 ;
      RECT  82.75 74.415 82.835 74.825 ;
      RECT  81.83 73.83 82.01 75.535 ;
      RECT  82.19 74.91 82.4 75.32 ;
      RECT  80.0 72.915 80.21 73.245 ;
      RECT  82.19 73.92 82.4 74.33 ;
      RECT  82.19 73.245 82.4 73.625 ;
      RECT  79.79 73.245 80.0 73.625 ;
      RECT  81.47 72.915 81.65 73.83 ;
      RECT  81.47 73.83 81.65 75.535 ;
      RECT  82.91 73.625 83.12 73.83 ;
      RECT  80.0 73.625 80.21 73.83 ;
      RECT  79.79 72.915 80.0 73.245 ;
      RECT  81.83 72.915 82.01 73.83 ;
      RECT  80.39 72.915 80.57 73.83 ;
      POLYGON  82.835 72.915 82.835 73.245 82.4 73.245 82.4 73.625 82.835 73.625 82.835 73.83 82.91 73.83 82.91 72.915 82.835 72.915 ;
      RECT  81.11 73.83 81.29 75.535 ;
      RECT  82.835 76.99 82.91 75.285 ;
      RECT  82.91 77.575 83.12 77.195 ;
      RECT  80.75 77.905 80.93 76.99 ;
      POLYGON  82.4 76.9 82.4 76.49 82.575 76.49 82.655 76.57 82.655 76.9 82.4 76.9 ;
      RECT  80.39 76.99 80.57 75.285 ;
      RECT  80.75 76.99 80.93 75.285 ;
      RECT  80.0 76.99 80.21 75.285 ;
      RECT  79.79 77.195 80.0 76.99 ;
      RECT  79.79 76.99 80.0 75.285 ;
      RECT  82.91 76.99 83.12 75.285 ;
      POLYGON  82.4 75.91 82.4 75.5 82.655 75.5 82.655 75.83 82.575 75.91 82.4 75.91 ;
      RECT  80.0 77.575 80.21 77.195 ;
      RECT  82.91 77.905 83.12 77.575 ;
      RECT  81.11 77.905 81.29 76.99 ;
      RECT  82.75 76.405 82.835 75.995 ;
      RECT  81.83 76.99 82.01 75.285 ;
      RECT  82.19 75.91 82.4 75.5 ;
      RECT  80.0 77.905 80.21 77.575 ;
      RECT  82.19 76.9 82.4 76.49 ;
      RECT  82.19 77.575 82.4 77.195 ;
      RECT  79.79 77.575 80.0 77.195 ;
      RECT  81.47 77.905 81.65 76.99 ;
      RECT  81.47 76.99 81.65 75.285 ;
      RECT  82.91 77.195 83.12 76.99 ;
      RECT  80.0 77.195 80.21 76.99 ;
      RECT  79.79 77.905 80.0 77.575 ;
      RECT  81.83 77.905 82.01 76.99 ;
      RECT  80.39 77.905 80.57 76.99 ;
      POLYGON  82.835 77.905 82.835 77.575 82.4 77.575 82.4 77.195 82.835 77.195 82.835 76.99 82.91 76.99 82.91 77.905 82.835 77.905 ;
      RECT  81.11 76.99 81.29 75.285 ;
      RECT  82.835 77.78 82.91 79.485 ;
      RECT  82.91 77.195 83.12 77.575 ;
      RECT  80.75 76.865 80.93 77.78 ;
      POLYGON  82.4 77.87 82.4 78.28 82.575 78.28 82.655 78.2 82.655 77.87 82.4 77.87 ;
      RECT  80.39 77.78 80.57 79.485 ;
      RECT  80.75 77.78 80.93 79.485 ;
      RECT  80.0 77.78 80.21 79.485 ;
      RECT  79.79 77.575 80.0 77.78 ;
      RECT  79.79 77.78 80.0 79.485 ;
      RECT  82.91 77.78 83.12 79.485 ;
      POLYGON  82.4 78.86 82.4 79.27 82.655 79.27 82.655 78.94 82.575 78.86 82.4 78.86 ;
      RECT  80.0 77.195 80.21 77.575 ;
      RECT  82.91 76.865 83.12 77.195 ;
      RECT  81.11 76.865 81.29 77.78 ;
      RECT  82.75 78.365 82.835 78.775 ;
      RECT  81.83 77.78 82.01 79.485 ;
      RECT  82.19 78.86 82.4 79.27 ;
      RECT  80.0 76.865 80.21 77.195 ;
      RECT  82.19 77.87 82.4 78.28 ;
      RECT  82.19 77.195 82.4 77.575 ;
      RECT  79.79 77.195 80.0 77.575 ;
      RECT  81.47 76.865 81.65 77.78 ;
      RECT  81.47 77.78 81.65 79.485 ;
      RECT  82.91 77.575 83.12 77.78 ;
      RECT  80.0 77.575 80.21 77.78 ;
      RECT  79.79 76.865 80.0 77.195 ;
      RECT  81.83 76.865 82.01 77.78 ;
      RECT  80.39 76.865 80.57 77.78 ;
      POLYGON  82.835 76.865 82.835 77.195 82.4 77.195 82.4 77.575 82.835 77.575 82.835 77.78 82.91 77.78 82.91 76.865 82.835 76.865 ;
      RECT  81.11 77.78 81.29 79.485 ;
      RECT  82.835 80.94 82.91 79.235 ;
      RECT  82.91 81.525 83.12 81.145 ;
      RECT  80.75 81.855 80.93 80.94 ;
      POLYGON  82.4 80.85 82.4 80.44 82.575 80.44 82.655 80.52 82.655 80.85 82.4 80.85 ;
      RECT  80.39 80.94 80.57 79.235 ;
      RECT  80.75 80.94 80.93 79.235 ;
      RECT  80.0 80.94 80.21 79.235 ;
      RECT  79.79 81.145 80.0 80.94 ;
      RECT  79.79 80.94 80.0 79.235 ;
      RECT  82.91 80.94 83.12 79.235 ;
      POLYGON  82.4 79.86 82.4 79.45 82.655 79.45 82.655 79.78 82.575 79.86 82.4 79.86 ;
      RECT  80.0 81.525 80.21 81.145 ;
      RECT  82.91 81.855 83.12 81.525 ;
      RECT  81.11 81.855 81.29 80.94 ;
      RECT  82.75 80.355 82.835 79.945 ;
      RECT  81.83 80.94 82.01 79.235 ;
      RECT  82.19 79.86 82.4 79.45 ;
      RECT  80.0 81.855 80.21 81.525 ;
      RECT  82.19 80.85 82.4 80.44 ;
      RECT  82.19 81.525 82.4 81.145 ;
      RECT  79.79 81.525 80.0 81.145 ;
      RECT  81.47 81.855 81.65 80.94 ;
      RECT  81.47 80.94 81.65 79.235 ;
      RECT  82.91 81.145 83.12 80.94 ;
      RECT  80.0 81.145 80.21 80.94 ;
      RECT  79.79 81.855 80.0 81.525 ;
      RECT  81.83 81.855 82.01 80.94 ;
      RECT  80.39 81.855 80.57 80.94 ;
      POLYGON  82.835 81.855 82.835 81.525 82.4 81.525 82.4 81.145 82.835 81.145 82.835 80.94 82.91 80.94 82.91 81.855 82.835 81.855 ;
      RECT  81.11 80.94 81.29 79.235 ;
      RECT  82.835 81.73 82.91 83.435 ;
      RECT  82.91 81.145 83.12 81.525 ;
      RECT  80.75 80.815 80.93 81.73 ;
      POLYGON  82.4 81.82 82.4 82.23 82.575 82.23 82.655 82.15 82.655 81.82 82.4 81.82 ;
      RECT  80.39 81.73 80.57 83.435 ;
      RECT  80.75 81.73 80.93 83.435 ;
      RECT  80.0 81.73 80.21 83.435 ;
      RECT  79.79 81.525 80.0 81.73 ;
      RECT  79.79 81.73 80.0 83.435 ;
      RECT  82.91 81.73 83.12 83.435 ;
      POLYGON  82.4 82.81 82.4 83.22 82.655 83.22 82.655 82.89 82.575 82.81 82.4 82.81 ;
      RECT  80.0 81.145 80.21 81.525 ;
      RECT  82.91 80.815 83.12 81.145 ;
      RECT  81.11 80.815 81.29 81.73 ;
      RECT  82.75 82.315 82.835 82.725 ;
      RECT  81.83 81.73 82.01 83.435 ;
      RECT  82.19 82.81 82.4 83.22 ;
      RECT  80.0 80.815 80.21 81.145 ;
      RECT  82.19 81.82 82.4 82.23 ;
      RECT  82.19 81.145 82.4 81.525 ;
      RECT  79.79 81.145 80.0 81.525 ;
      RECT  81.47 80.815 81.65 81.73 ;
      RECT  81.47 81.73 81.65 83.435 ;
      RECT  82.91 81.525 83.12 81.73 ;
      RECT  80.0 81.525 80.21 81.73 ;
      RECT  79.79 80.815 80.0 81.145 ;
      RECT  81.83 80.815 82.01 81.73 ;
      RECT  80.39 80.815 80.57 81.73 ;
      POLYGON  82.835 80.815 82.835 81.145 82.4 81.145 82.4 81.525 82.835 81.525 82.835 81.73 82.91 81.73 82.91 80.815 82.835 80.815 ;
      RECT  81.11 81.73 81.29 83.435 ;
      RECT  82.835 84.89 82.91 83.185 ;
      RECT  82.91 85.475 83.12 85.095 ;
      RECT  80.75 85.805 80.93 84.89 ;
      POLYGON  82.4 84.8 82.4 84.39 82.575 84.39 82.655 84.47 82.655 84.8 82.4 84.8 ;
      RECT  80.39 84.89 80.57 83.185 ;
      RECT  80.75 84.89 80.93 83.185 ;
      RECT  80.0 84.89 80.21 83.185 ;
      RECT  79.79 85.095 80.0 84.89 ;
      RECT  79.79 84.89 80.0 83.185 ;
      RECT  82.91 84.89 83.12 83.185 ;
      POLYGON  82.4 83.81 82.4 83.4 82.655 83.4 82.655 83.73 82.575 83.81 82.4 83.81 ;
      RECT  80.0 85.475 80.21 85.095 ;
      RECT  82.91 85.805 83.12 85.475 ;
      RECT  81.11 85.805 81.29 84.89 ;
      RECT  82.75 84.305 82.835 83.895 ;
      RECT  81.83 84.89 82.01 83.185 ;
      RECT  82.19 83.81 82.4 83.4 ;
      RECT  80.0 85.805 80.21 85.475 ;
      RECT  82.19 84.8 82.4 84.39 ;
      RECT  82.19 85.475 82.4 85.095 ;
      RECT  79.79 85.475 80.0 85.095 ;
      RECT  81.47 85.805 81.65 84.89 ;
      RECT  81.47 84.89 81.65 83.185 ;
      RECT  82.91 85.095 83.12 84.89 ;
      RECT  80.0 85.095 80.21 84.89 ;
      RECT  79.79 85.805 80.0 85.475 ;
      RECT  81.83 85.805 82.01 84.89 ;
      RECT  80.39 85.805 80.57 84.89 ;
      POLYGON  82.835 85.805 82.835 85.475 82.4 85.475 82.4 85.095 82.835 85.095 82.835 84.89 82.91 84.89 82.91 85.805 82.835 85.805 ;
      RECT  81.11 84.89 81.29 83.185 ;
      RECT  82.835 85.68 82.91 87.385 ;
      RECT  82.91 85.095 83.12 85.475 ;
      RECT  80.75 84.765 80.93 85.68 ;
      POLYGON  82.4 85.77 82.4 86.18 82.575 86.18 82.655 86.1 82.655 85.77 82.4 85.77 ;
      RECT  80.39 85.68 80.57 87.385 ;
      RECT  80.75 85.68 80.93 87.385 ;
      RECT  80.0 85.68 80.21 87.385 ;
      RECT  79.79 85.475 80.0 85.68 ;
      RECT  79.79 85.68 80.0 87.385 ;
      RECT  82.91 85.68 83.12 87.385 ;
      POLYGON  82.4 86.76 82.4 87.17 82.655 87.17 82.655 86.84 82.575 86.76 82.4 86.76 ;
      RECT  80.0 85.095 80.21 85.475 ;
      RECT  82.91 84.765 83.12 85.095 ;
      RECT  81.11 84.765 81.29 85.68 ;
      RECT  82.75 86.265 82.835 86.675 ;
      RECT  81.83 85.68 82.01 87.385 ;
      RECT  82.19 86.76 82.4 87.17 ;
      RECT  80.0 84.765 80.21 85.095 ;
      RECT  82.19 85.77 82.4 86.18 ;
      RECT  82.19 85.095 82.4 85.475 ;
      RECT  79.79 85.095 80.0 85.475 ;
      RECT  81.47 84.765 81.65 85.68 ;
      RECT  81.47 85.68 81.65 87.385 ;
      RECT  82.91 85.475 83.12 85.68 ;
      RECT  80.0 85.475 80.21 85.68 ;
      RECT  79.79 84.765 80.0 85.095 ;
      RECT  81.83 84.765 82.01 85.68 ;
      RECT  80.39 84.765 80.57 85.68 ;
      POLYGON  82.835 84.765 82.835 85.095 82.4 85.095 82.4 85.475 82.835 85.475 82.835 85.68 82.91 85.68 82.91 84.765 82.835 84.765 ;
      RECT  81.11 85.68 81.29 87.385 ;
      RECT  82.835 88.84 82.91 87.135 ;
      RECT  82.91 89.425 83.12 89.045 ;
      RECT  80.75 89.755 80.93 88.84 ;
      POLYGON  82.4 88.75 82.4 88.34 82.575 88.34 82.655 88.42 82.655 88.75 82.4 88.75 ;
      RECT  80.39 88.84 80.57 87.135 ;
      RECT  80.75 88.84 80.93 87.135 ;
      RECT  80.0 88.84 80.21 87.135 ;
      RECT  79.79 89.045 80.0 88.84 ;
      RECT  79.79 88.84 80.0 87.135 ;
      RECT  82.91 88.84 83.12 87.135 ;
      POLYGON  82.4 87.76 82.4 87.35 82.655 87.35 82.655 87.68 82.575 87.76 82.4 87.76 ;
      RECT  80.0 89.425 80.21 89.045 ;
      RECT  82.91 89.755 83.12 89.425 ;
      RECT  81.11 89.755 81.29 88.84 ;
      RECT  82.75 88.255 82.835 87.845 ;
      RECT  81.83 88.84 82.01 87.135 ;
      RECT  82.19 87.76 82.4 87.35 ;
      RECT  80.0 89.755 80.21 89.425 ;
      RECT  82.19 88.75 82.4 88.34 ;
      RECT  82.19 89.425 82.4 89.045 ;
      RECT  79.79 89.425 80.0 89.045 ;
      RECT  81.47 89.755 81.65 88.84 ;
      RECT  81.47 88.84 81.65 87.135 ;
      RECT  82.91 89.045 83.12 88.84 ;
      RECT  80.0 89.045 80.21 88.84 ;
      RECT  79.79 89.755 80.0 89.425 ;
      RECT  81.83 89.755 82.01 88.84 ;
      RECT  80.39 89.755 80.57 88.84 ;
      POLYGON  82.835 89.755 82.835 89.425 82.4 89.425 82.4 89.045 82.835 89.045 82.835 88.84 82.91 88.84 82.91 89.755 82.835 89.755 ;
      RECT  81.11 88.84 81.29 87.135 ;
      RECT  82.835 89.63 82.91 91.335 ;
      RECT  82.91 89.045 83.12 89.425 ;
      RECT  80.75 88.715 80.93 89.63 ;
      POLYGON  82.4 89.72 82.4 90.13 82.575 90.13 82.655 90.05 82.655 89.72 82.4 89.72 ;
      RECT  80.39 89.63 80.57 91.335 ;
      RECT  80.75 89.63 80.93 91.335 ;
      RECT  80.0 89.63 80.21 91.335 ;
      RECT  79.79 89.425 80.0 89.63 ;
      RECT  79.79 89.63 80.0 91.335 ;
      RECT  82.91 89.63 83.12 91.335 ;
      POLYGON  82.4 90.71 82.4 91.12 82.655 91.12 82.655 90.79 82.575 90.71 82.4 90.71 ;
      RECT  80.0 89.045 80.21 89.425 ;
      RECT  82.91 88.715 83.12 89.045 ;
      RECT  81.11 88.715 81.29 89.63 ;
      RECT  82.75 90.215 82.835 90.625 ;
      RECT  81.83 89.63 82.01 91.335 ;
      RECT  82.19 90.71 82.4 91.12 ;
      RECT  80.0 88.715 80.21 89.045 ;
      RECT  82.19 89.72 82.4 90.13 ;
      RECT  82.19 89.045 82.4 89.425 ;
      RECT  79.79 89.045 80.0 89.425 ;
      RECT  81.47 88.715 81.65 89.63 ;
      RECT  81.47 89.63 81.65 91.335 ;
      RECT  82.91 89.425 83.12 89.63 ;
      RECT  80.0 89.425 80.21 89.63 ;
      RECT  79.79 88.715 80.0 89.045 ;
      RECT  81.83 88.715 82.01 89.63 ;
      RECT  80.39 88.715 80.57 89.63 ;
      POLYGON  82.835 88.715 82.835 89.045 82.4 89.045 82.4 89.425 82.835 89.425 82.835 89.63 82.91 89.63 82.91 88.715 82.835 88.715 ;
      RECT  81.11 89.63 81.29 91.335 ;
      RECT  82.835 92.79 82.91 91.085 ;
      RECT  82.91 93.375 83.12 92.995 ;
      RECT  80.75 93.705 80.93 92.79 ;
      POLYGON  82.4 92.7 82.4 92.29 82.575 92.29 82.655 92.37 82.655 92.7 82.4 92.7 ;
      RECT  80.39 92.79 80.57 91.085 ;
      RECT  80.75 92.79 80.93 91.085 ;
      RECT  80.0 92.79 80.21 91.085 ;
      RECT  79.79 92.995 80.0 92.79 ;
      RECT  79.79 92.79 80.0 91.085 ;
      RECT  82.91 92.79 83.12 91.085 ;
      POLYGON  82.4 91.71 82.4 91.3 82.655 91.3 82.655 91.63 82.575 91.71 82.4 91.71 ;
      RECT  80.0 93.375 80.21 92.995 ;
      RECT  82.91 93.705 83.12 93.375 ;
      RECT  81.11 93.705 81.29 92.79 ;
      RECT  82.75 92.205 82.835 91.795 ;
      RECT  81.83 92.79 82.01 91.085 ;
      RECT  82.19 91.71 82.4 91.3 ;
      RECT  80.0 93.705 80.21 93.375 ;
      RECT  82.19 92.7 82.4 92.29 ;
      RECT  82.19 93.375 82.4 92.995 ;
      RECT  79.79 93.375 80.0 92.995 ;
      RECT  81.47 93.705 81.65 92.79 ;
      RECT  81.47 92.79 81.65 91.085 ;
      RECT  82.91 92.995 83.12 92.79 ;
      RECT  80.0 92.995 80.21 92.79 ;
      RECT  79.79 93.705 80.0 93.375 ;
      RECT  81.83 93.705 82.01 92.79 ;
      RECT  80.39 93.705 80.57 92.79 ;
      POLYGON  82.835 93.705 82.835 93.375 82.4 93.375 82.4 92.995 82.835 92.995 82.835 92.79 82.91 92.79 82.91 93.705 82.835 93.705 ;
      RECT  81.11 92.79 81.29 91.085 ;
      RECT  82.835 93.58 82.91 95.285 ;
      RECT  82.91 92.995 83.12 93.375 ;
      RECT  80.75 92.665 80.93 93.58 ;
      POLYGON  82.4 93.67 82.4 94.08 82.575 94.08 82.655 94.0 82.655 93.67 82.4 93.67 ;
      RECT  80.39 93.58 80.57 95.285 ;
      RECT  80.75 93.58 80.93 95.285 ;
      RECT  80.0 93.58 80.21 95.285 ;
      RECT  79.79 93.375 80.0 93.58 ;
      RECT  79.79 93.58 80.0 95.285 ;
      RECT  82.91 93.58 83.12 95.285 ;
      POLYGON  82.4 94.66 82.4 95.07 82.655 95.07 82.655 94.74 82.575 94.66 82.4 94.66 ;
      RECT  80.0 92.995 80.21 93.375 ;
      RECT  82.91 92.665 83.12 92.995 ;
      RECT  81.11 92.665 81.29 93.58 ;
      RECT  82.75 94.165 82.835 94.575 ;
      RECT  81.83 93.58 82.01 95.285 ;
      RECT  82.19 94.66 82.4 95.07 ;
      RECT  80.0 92.665 80.21 92.995 ;
      RECT  82.19 93.67 82.4 94.08 ;
      RECT  82.19 92.995 82.4 93.375 ;
      RECT  79.79 92.995 80.0 93.375 ;
      RECT  81.47 92.665 81.65 93.58 ;
      RECT  81.47 93.58 81.65 95.285 ;
      RECT  82.91 93.375 83.12 93.58 ;
      RECT  80.0 93.375 80.21 93.58 ;
      RECT  79.79 92.665 80.0 92.995 ;
      RECT  81.83 92.665 82.01 93.58 ;
      RECT  80.39 92.665 80.57 93.58 ;
      POLYGON  82.835 92.665 82.835 92.995 82.4 92.995 82.4 93.375 82.835 93.375 82.835 93.58 82.91 93.58 82.91 92.665 82.835 92.665 ;
      RECT  81.11 93.58 81.29 95.285 ;
      RECT  81.11 96.345 81.29 94.765 ;
      RECT  80.75 96.345 80.93 94.765 ;
      RECT  81.2 96.345 81.33 95.635 ;
      RECT  81.47 96.345 81.65 94.765 ;
      RECT  81.07 96.345 81.2 95.635 ;
      RECT  80.75 97.135 80.93 96.345 ;
      RECT  80.39 97.135 80.57 96.345 ;
      RECT  81.83 97.135 82.01 96.345 ;
      RECT  81.11 97.135 81.29 96.345 ;
      RECT  81.47 97.135 81.65 96.345 ;
      RECT  80.39 96.345 80.57 94.765 ;
      RECT  81.83 96.345 82.01 94.765 ;
      RECT  81.11 61.98 81.29 63.685 ;
      RECT  81.11 91.085 81.29 92.79 ;
      RECT  81.11 65.93 81.29 67.635 ;
      RECT  81.11 81.73 81.29 83.435 ;
      RECT  81.11 87.135 81.29 88.84 ;
      RECT  81.11 73.83 81.29 75.535 ;
      RECT  81.11 75.285 81.29 76.99 ;
      RECT  81.11 83.185 81.29 84.89 ;
      RECT  81.11 93.58 81.29 95.285 ;
      RECT  81.11 79.235 81.29 80.94 ;
      RECT  81.11 59.485 81.29 61.19 ;
      RECT  81.11 67.385 81.29 69.09 ;
      RECT  81.11 77.78 81.29 79.485 ;
      RECT  81.11 63.435 81.29 65.14 ;
      RECT  81.11 69.88 81.29 71.585 ;
      RECT  81.11 85.68 81.29 87.385 ;
      RECT  81.11 71.335 81.29 73.04 ;
      RECT  81.11 89.63 81.29 91.335 ;
      RECT  76.595 61.19 76.67 59.485 ;
      RECT  76.67 61.775 76.88 61.395 ;
      RECT  74.51 62.105 74.69 61.19 ;
      POLYGON  76.16 61.1 76.16 60.69 76.335 60.69 76.415 60.77 76.415 61.1 76.16 61.1 ;
      RECT  74.15 61.19 74.33 59.485 ;
      RECT  74.51 61.19 74.69 59.485 ;
      RECT  73.76 61.19 73.97 59.485 ;
      RECT  73.55 61.395 73.76 61.19 ;
      RECT  73.55 61.19 73.76 59.485 ;
      RECT  76.67 61.19 76.88 59.485 ;
      POLYGON  76.16 60.11 76.16 59.7 76.415 59.7 76.415 60.03 76.335 60.11 76.16 60.11 ;
      RECT  73.76 61.775 73.97 61.395 ;
      RECT  76.67 62.105 76.88 61.775 ;
      RECT  74.87 62.105 75.05 61.19 ;
      RECT  76.51 60.605 76.595 60.195 ;
      RECT  75.59 61.19 75.77 59.485 ;
      RECT  75.95 60.11 76.16 59.7 ;
      RECT  73.76 62.105 73.97 61.775 ;
      RECT  75.95 61.1 76.16 60.69 ;
      RECT  75.95 61.775 76.16 61.395 ;
      RECT  73.55 61.775 73.76 61.395 ;
      RECT  75.23 62.105 75.41 61.19 ;
      RECT  75.23 61.19 75.41 59.485 ;
      RECT  76.67 61.395 76.88 61.19 ;
      RECT  73.76 61.395 73.97 61.19 ;
      RECT  73.55 62.105 73.76 61.775 ;
      RECT  75.59 62.105 75.77 61.19 ;
      RECT  74.15 62.105 74.33 61.19 ;
      POLYGON  76.595 62.105 76.595 61.775 76.16 61.775 76.16 61.395 76.595 61.395 76.595 61.19 76.67 61.19 76.67 62.105 76.595 62.105 ;
      RECT  74.87 61.19 75.05 59.485 ;
      RECT  77.165 61.19 77.09 59.485 ;
      RECT  77.09 61.775 76.88 61.395 ;
      RECT  79.25 62.105 79.07 61.19 ;
      POLYGON  77.6 61.1 77.6 60.69 77.425 60.69 77.345 60.77 77.345 61.1 77.6 61.1 ;
      RECT  79.61 61.19 79.43 59.485 ;
      RECT  79.25 61.19 79.07 59.485 ;
      RECT  80.0 61.19 79.79 59.485 ;
      RECT  80.21 61.395 80.0 61.19 ;
      RECT  80.21 61.19 80.0 59.485 ;
      RECT  77.09 61.19 76.88 59.485 ;
      POLYGON  77.6 60.11 77.6 59.7 77.345 59.7 77.345 60.03 77.425 60.11 77.6 60.11 ;
      RECT  80.0 61.775 79.79 61.395 ;
      RECT  77.09 62.105 76.88 61.775 ;
      RECT  78.89 62.105 78.71 61.19 ;
      RECT  77.25 60.605 77.165 60.195 ;
      RECT  78.17 61.19 77.99 59.485 ;
      RECT  77.81 60.11 77.6 59.7 ;
      RECT  80.0 62.105 79.79 61.775 ;
      RECT  77.81 61.1 77.6 60.69 ;
      RECT  77.81 61.775 77.6 61.395 ;
      RECT  80.21 61.775 80.0 61.395 ;
      RECT  78.53 62.105 78.35 61.19 ;
      RECT  78.53 61.19 78.35 59.485 ;
      RECT  77.09 61.395 76.88 61.19 ;
      RECT  80.0 61.395 79.79 61.19 ;
      RECT  80.21 62.105 80.0 61.775 ;
      RECT  78.17 62.105 77.99 61.19 ;
      RECT  79.61 62.105 79.43 61.19 ;
      POLYGON  77.165 62.105 77.165 61.775 77.6 61.775 77.6 61.395 77.165 61.395 77.165 61.19 77.09 61.19 77.09 62.105 77.165 62.105 ;
      RECT  78.89 61.19 78.71 59.485 ;
      RECT  74.15 61.585 74.33 59.61 ;
      RECT  74.51 61.585 74.69 59.61 ;
      RECT  75.23 61.585 75.41 59.61 ;
      RECT  75.59 61.585 75.77 59.61 ;
      RECT  79.43 61.585 79.61 59.61 ;
      RECT  79.07 61.585 79.25 59.61 ;
      RECT  78.35 61.585 78.53 59.61 ;
      RECT  77.99 61.585 78.17 59.61 ;
      RECT  78.71 61.19 78.89 59.485 ;
      RECT  74.87 61.19 75.05 59.485 ;
      RECT  76.595 93.58 76.67 95.285 ;
      RECT  76.67 92.995 76.88 93.375 ;
      RECT  74.51 92.665 74.69 93.58 ;
      POLYGON  76.16 93.67 76.16 94.08 76.335 94.08 76.415 94.0 76.415 93.67 76.16 93.67 ;
      RECT  74.15 93.58 74.33 95.285 ;
      RECT  74.51 93.58 74.69 95.285 ;
      RECT  73.76 93.58 73.97 95.285 ;
      RECT  73.55 93.375 73.76 93.58 ;
      RECT  73.55 93.58 73.76 95.285 ;
      RECT  76.67 93.58 76.88 95.285 ;
      POLYGON  76.16 94.66 76.16 95.07 76.415 95.07 76.415 94.74 76.335 94.66 76.16 94.66 ;
      RECT  73.76 92.995 73.97 93.375 ;
      RECT  76.67 92.665 76.88 92.995 ;
      RECT  74.87 92.665 75.05 93.58 ;
      RECT  76.51 94.165 76.595 94.575 ;
      RECT  75.59 93.58 75.77 95.285 ;
      RECT  75.95 94.66 76.16 95.07 ;
      RECT  73.76 92.665 73.97 92.995 ;
      RECT  75.95 93.67 76.16 94.08 ;
      RECT  75.95 92.995 76.16 93.375 ;
      RECT  73.55 92.995 73.76 93.375 ;
      RECT  75.23 92.665 75.41 93.58 ;
      RECT  75.23 93.58 75.41 95.285 ;
      RECT  76.67 93.375 76.88 93.58 ;
      RECT  73.76 93.375 73.97 93.58 ;
      RECT  73.55 92.665 73.76 92.995 ;
      RECT  75.59 92.665 75.77 93.58 ;
      RECT  74.15 92.665 74.33 93.58 ;
      POLYGON  76.595 92.665 76.595 92.995 76.16 92.995 76.16 93.375 76.595 93.375 76.595 93.58 76.67 93.58 76.67 92.665 76.595 92.665 ;
      RECT  74.87 93.58 75.05 95.285 ;
      RECT  77.165 93.58 77.09 95.285 ;
      RECT  77.09 92.995 76.88 93.375 ;
      RECT  79.25 92.665 79.07 93.58 ;
      POLYGON  77.6 93.67 77.6 94.08 77.425 94.08 77.345 94.0 77.345 93.67 77.6 93.67 ;
      RECT  79.61 93.58 79.43 95.285 ;
      RECT  79.25 93.58 79.07 95.285 ;
      RECT  80.0 93.58 79.79 95.285 ;
      RECT  80.21 93.375 80.0 93.58 ;
      RECT  80.21 93.58 80.0 95.285 ;
      RECT  77.09 93.58 76.88 95.285 ;
      POLYGON  77.6 94.66 77.6 95.07 77.345 95.07 77.345 94.74 77.425 94.66 77.6 94.66 ;
      RECT  80.0 92.995 79.79 93.375 ;
      RECT  77.09 92.665 76.88 92.995 ;
      RECT  78.89 92.665 78.71 93.58 ;
      RECT  77.25 94.165 77.165 94.575 ;
      RECT  78.17 93.58 77.99 95.285 ;
      RECT  77.81 94.66 77.6 95.07 ;
      RECT  80.0 92.665 79.79 92.995 ;
      RECT  77.81 93.67 77.6 94.08 ;
      RECT  77.81 92.995 77.6 93.375 ;
      RECT  80.21 92.995 80.0 93.375 ;
      RECT  78.53 92.665 78.35 93.58 ;
      RECT  78.53 93.58 78.35 95.285 ;
      RECT  77.09 93.375 76.88 93.58 ;
      RECT  80.0 93.375 79.79 93.58 ;
      RECT  80.21 92.665 80.0 92.995 ;
      RECT  78.17 92.665 77.99 93.58 ;
      RECT  79.61 92.665 79.43 93.58 ;
      POLYGON  77.165 92.665 77.165 92.995 77.6 92.995 77.6 93.375 77.165 93.375 77.165 93.58 77.09 93.58 77.09 92.665 77.165 92.665 ;
      RECT  78.89 93.58 78.71 95.285 ;
      RECT  74.15 93.185 74.33 95.16 ;
      RECT  74.51 93.185 74.69 95.16 ;
      RECT  75.23 93.185 75.41 95.16 ;
      RECT  75.59 93.185 75.77 95.16 ;
      RECT  79.43 93.185 79.61 95.16 ;
      RECT  79.07 93.185 79.25 95.16 ;
      RECT  78.35 93.185 78.53 95.16 ;
      RECT  77.99 93.185 78.17 95.16 ;
      RECT  78.71 93.58 78.89 95.285 ;
      RECT  74.87 93.58 75.05 95.285 ;
      RECT  74.87 58.425 75.05 60.005 ;
      RECT  74.51 58.425 74.69 60.005 ;
      RECT  74.96 58.425 75.09 59.135 ;
      RECT  75.23 58.425 75.41 60.005 ;
      RECT  74.83 58.425 74.96 59.135 ;
      RECT  74.51 57.635 74.69 58.425 ;
      RECT  74.15 57.635 74.33 58.425 ;
      RECT  75.59 57.635 75.77 58.425 ;
      RECT  74.87 57.635 75.05 58.425 ;
      RECT  75.23 57.635 75.41 58.425 ;
      RECT  74.15 58.425 74.33 60.005 ;
      RECT  75.59 58.425 75.77 60.005 ;
      RECT  78.89 58.425 78.71 60.005 ;
      RECT  79.25 58.425 79.07 60.005 ;
      RECT  78.8 58.425 78.67 59.135 ;
      RECT  78.53 58.425 78.35 60.005 ;
      RECT  78.93 58.425 78.8 59.135 ;
      RECT  79.25 57.635 79.07 58.425 ;
      RECT  79.61 57.635 79.43 58.425 ;
      RECT  78.17 57.635 77.99 58.425 ;
      RECT  78.89 57.635 78.71 58.425 ;
      RECT  78.53 57.635 78.35 58.425 ;
      RECT  79.61 58.425 79.43 60.005 ;
      RECT  78.17 58.425 77.99 60.005 ;
      RECT  74.15 57.635 74.33 59.61 ;
      RECT  74.51 57.635 74.69 59.61 ;
      RECT  75.23 57.635 75.41 59.61 ;
      RECT  75.59 57.635 75.77 59.61 ;
      RECT  79.43 57.635 79.61 59.61 ;
      RECT  79.07 57.635 79.25 59.61 ;
      RECT  78.35 57.635 78.53 59.61 ;
      RECT  77.99 57.635 78.17 59.61 ;
      RECT  74.87 96.345 75.05 94.765 ;
      RECT  74.51 96.345 74.69 94.765 ;
      RECT  74.96 96.345 75.09 95.635 ;
      RECT  75.23 96.345 75.41 94.765 ;
      RECT  74.83 96.345 74.96 95.635 ;
      RECT  74.51 97.135 74.69 96.345 ;
      RECT  74.15 97.135 74.33 96.345 ;
      RECT  75.59 97.135 75.77 96.345 ;
      RECT  74.87 97.135 75.05 96.345 ;
      RECT  75.23 97.135 75.41 96.345 ;
      RECT  74.15 96.345 74.33 94.765 ;
      RECT  75.59 96.345 75.77 94.765 ;
      RECT  78.89 96.345 78.71 94.765 ;
      RECT  79.25 96.345 79.07 94.765 ;
      RECT  78.8 96.345 78.67 95.635 ;
      RECT  78.53 96.345 78.35 94.765 ;
      RECT  78.93 96.345 78.8 95.635 ;
      RECT  79.25 97.135 79.07 96.345 ;
      RECT  79.61 97.135 79.43 96.345 ;
      RECT  78.17 97.135 77.99 96.345 ;
      RECT  78.89 97.135 78.71 96.345 ;
      RECT  78.53 97.135 78.35 96.345 ;
      RECT  79.61 96.345 79.43 94.765 ;
      RECT  78.17 96.345 77.99 94.765 ;
      RECT  74.15 97.135 74.33 95.16 ;
      RECT  74.51 97.135 74.69 95.16 ;
      RECT  75.23 97.135 75.41 95.16 ;
      RECT  75.59 97.135 75.77 95.16 ;
      RECT  79.43 97.135 79.61 95.16 ;
      RECT  79.07 97.135 79.25 95.16 ;
      RECT  78.35 97.135 78.53 95.16 ;
      RECT  77.99 97.135 78.17 95.16 ;
      RECT  74.15 57.635 74.33 97.135 ;
      RECT  74.51 57.635 74.69 97.135 ;
      RECT  75.23 57.635 75.41 97.135 ;
      RECT  75.59 57.635 75.77 97.135 ;
      RECT  79.43 57.635 79.61 97.135 ;
      RECT  79.07 57.635 79.25 97.135 ;
      RECT  78.35 57.635 78.53 97.135 ;
      RECT  77.99 57.635 78.17 97.135 ;
      RECT  73.19 57.635 73.37 97.135 ;
      RECT  72.83 57.635 73.01 97.135 ;
      RECT  81.47 57.635 81.65 97.135 ;
      RECT  81.83 57.635 82.01 97.135 ;
      RECT  72.47 91.085 72.65 92.79 ;
      RECT  81.11 79.235 81.29 80.94 ;
      RECT  81.11 93.58 81.29 95.285 ;
      RECT  81.11 71.335 81.29 73.04 ;
      RECT  72.47 61.98 72.65 63.685 ;
      RECT  81.11 69.88 81.29 71.585 ;
      RECT  72.47 63.435 72.65 65.14 ;
      RECT  72.47 83.185 72.65 84.89 ;
      RECT  81.11 63.435 81.29 65.14 ;
      RECT  72.47 73.83 72.65 75.535 ;
      RECT  81.11 75.285 81.29 76.99 ;
      RECT  72.47 69.88 72.65 71.585 ;
      RECT  81.11 59.485 81.29 61.19 ;
      RECT  72.47 59.485 72.65 61.19 ;
      RECT  81.11 85.68 81.29 87.385 ;
      RECT  81.11 61.98 81.29 63.685 ;
      RECT  81.11 77.78 81.29 79.485 ;
      RECT  72.47 77.78 72.65 79.485 ;
      RECT  81.11 91.085 81.29 92.79 ;
      RECT  72.47 67.385 72.65 69.09 ;
      RECT  72.47 81.73 72.65 83.435 ;
      RECT  72.47 71.335 72.65 73.04 ;
      RECT  81.11 87.135 81.29 88.84 ;
      RECT  81.11 67.385 81.29 69.09 ;
      RECT  81.11 81.73 81.29 83.435 ;
      RECT  72.47 65.93 72.65 67.635 ;
      RECT  81.11 89.63 81.29 91.335 ;
      RECT  81.11 65.93 81.29 67.635 ;
      RECT  72.47 93.58 72.65 95.285 ;
      RECT  81.11 83.185 81.29 84.89 ;
      RECT  72.47 79.235 72.65 80.94 ;
      RECT  72.47 89.63 72.65 91.335 ;
      RECT  81.11 73.83 81.29 75.535 ;
      RECT  72.47 85.68 72.65 87.385 ;
      RECT  72.47 87.135 72.65 88.84 ;
      RECT  72.47 75.285 72.65 76.99 ;
      RECT  73.43 52.605 73.29 56.375 ;
      RECT  71.11 52.605 70.97 56.375 ;
      RECT  74.09 52.605 74.23 56.375 ;
      RECT  76.41 52.605 76.55 56.375 ;
      RECT  79.67 52.605 79.53 56.375 ;
      RECT  77.35 52.605 77.21 56.375 ;
      RECT  73.29 52.605 73.43 56.375 ;
      RECT  70.97 52.605 71.11 56.375 ;
      RECT  74.09 52.605 74.23 56.375 ;
      RECT  76.41 52.605 76.55 56.375 ;
      RECT  79.53 52.605 79.67 56.375 ;
      RECT  77.21 52.605 77.35 56.375 ;
      RECT  74.74 45.715 74.91 51.345 ;
      RECT  75.12 40.065 75.26 45.485 ;
      RECT  75.55 40.42 75.78 40.79 ;
      RECT  75.55 42.025 75.78 42.405 ;
      RECT  75.9 50.09 76.13 50.46 ;
      RECT  74.28 40.065 74.51 41.335 ;
      RECT  75.12 45.485 75.46 45.775 ;
      RECT  74.74 40.065 74.91 45.485 ;
      RECT  74.68 45.485 74.97 45.715 ;
      RECT  75.45 46.235 75.76 46.575 ;
      RECT  75.12 45.775 75.26 51.345 ;
      RECT  74.23 50.885 74.52 51.185 ;
      RECT  78.4 45.715 78.23 51.345 ;
      RECT  78.02 40.065 77.88 45.485 ;
      RECT  77.59 40.42 77.36 40.79 ;
      RECT  77.59 42.025 77.36 42.405 ;
      RECT  77.24 50.09 77.01 50.46 ;
      RECT  78.86 40.065 78.63 41.335 ;
      RECT  78.02 45.485 77.68 45.775 ;
      RECT  78.4 40.065 78.23 45.485 ;
      RECT  78.46 45.485 78.17 45.715 ;
      RECT  77.69 46.235 77.38 46.575 ;
      RECT  78.02 45.775 77.88 51.345 ;
      RECT  78.91 50.885 78.62 51.185 ;
      RECT  74.28 40.065 74.51 41.335 ;
      RECT  74.74 45.715 74.91 51.345 ;
      RECT  75.12 45.775 75.26 51.345 ;
      RECT  78.63 40.065 78.86 41.335 ;
      RECT  78.23 45.715 78.4 51.345 ;
      RECT  77.88 45.775 78.02 51.345 ;
      RECT  74.825 36.555 75.365 36.725 ;
      RECT  74.925 29.59 75.355 29.82 ;
      RECT  75.27 38.255 75.555 38.545 ;
      RECT  74.255 29.22 76.26 29.39 ;
      RECT  75.4 38.545 75.55 38.805 ;
      RECT  75.035 28.77 75.335 29.05 ;
      RECT  74.255 29.39 74.545 29.53 ;
      RECT  74.39 38.545 74.54 38.805 ;
      RECT  74.825 36.525 75.255 36.555 ;
      RECT  74.825 34.34 75.255 34.57 ;
      RECT  75.43 32.695 75.86 32.9 ;
      RECT  74.825 36.725 75.255 36.755 ;
      RECT  74.385 38.255 74.67 38.545 ;
      RECT  74.855 31.67 75.285 31.9 ;
      RECT  75.495 32.67 75.86 32.695 ;
      RECT  78.315 36.555 77.775 36.725 ;
      RECT  78.215 29.59 77.785 29.82 ;
      RECT  77.87 38.255 77.585 38.545 ;
      RECT  78.885 29.22 76.88 29.39 ;
      RECT  77.74 38.545 77.59 38.805 ;
      RECT  78.105 28.77 77.805 29.05 ;
      RECT  78.885 29.39 78.595 29.53 ;
      RECT  78.75 38.545 78.6 38.805 ;
      RECT  78.315 36.525 77.885 36.555 ;
      RECT  78.315 34.34 77.885 34.57 ;
      RECT  77.71 32.695 77.28 32.9 ;
      RECT  78.315 36.725 77.885 36.755 ;
      RECT  78.755 38.255 78.47 38.545 ;
      RECT  78.285 31.67 77.855 31.9 ;
      RECT  77.645 32.67 77.28 32.695 ;
      RECT  75.035 28.77 75.335 29.05 ;
      RECT  77.805 28.77 78.105 29.05 ;
      RECT  74.39 38.545 74.54 38.805 ;
      RECT  75.4 38.545 75.55 38.805 ;
      RECT  78.6 38.545 78.75 38.805 ;
      RECT  77.59 38.545 77.74 38.805 ;
      RECT  73.76 29.22 80.0 29.36 ;
      RECT  73.29 56.375 73.43 52.605 ;
      RECT  70.97 56.375 71.11 52.605 ;
      RECT  74.28 41.335 74.51 40.065 ;
      RECT  78.63 41.335 78.86 40.065 ;
      RECT  75.035 29.05 75.335 28.77 ;
      RECT  77.805 29.05 78.105 28.77 ;
      RECT  73.76 29.36 80.0 29.22 ;
      RECT  74.09 102.165 74.23 98.395 ;
      RECT  76.41 102.165 76.55 98.395 ;
      RECT  79.67 102.165 79.53 98.395 ;
      RECT  77.35 102.165 77.21 98.395 ;
      RECT  80.33 102.165 80.47 98.395 ;
      RECT  82.65 102.165 82.79 98.395 ;
      RECT  74.09 102.165 74.23 98.395 ;
      RECT  76.41 102.165 76.55 98.395 ;
      RECT  79.53 102.165 79.67 98.395 ;
      RECT  77.21 102.165 77.35 98.395 ;
      RECT  80.33 102.165 80.47 98.395 ;
      RECT  82.65 102.165 82.79 98.395 ;
      RECT  74.74 109.055 74.91 103.425 ;
      RECT  75.12 114.705 75.26 109.285 ;
      RECT  75.55 114.35 75.78 113.98 ;
      RECT  75.55 112.745 75.78 112.365 ;
      RECT  75.9 104.68 76.13 104.31 ;
      RECT  74.28 114.705 74.51 113.435 ;
      RECT  75.12 109.285 75.46 108.995 ;
      RECT  74.74 114.705 74.91 109.285 ;
      RECT  74.68 109.285 74.97 109.055 ;
      RECT  75.45 108.535 75.76 108.195 ;
      RECT  75.12 108.995 75.26 103.425 ;
      RECT  74.23 103.885 74.52 103.585 ;
      RECT  78.4 109.055 78.23 103.425 ;
      RECT  78.02 114.705 77.88 109.285 ;
      RECT  77.59 114.35 77.36 113.98 ;
      RECT  77.59 112.745 77.36 112.365 ;
      RECT  77.24 104.68 77.01 104.31 ;
      RECT  78.86 114.705 78.63 113.435 ;
      RECT  78.02 109.285 77.68 108.995 ;
      RECT  78.4 114.705 78.23 109.285 ;
      RECT  78.46 109.285 78.17 109.055 ;
      RECT  77.69 108.535 77.38 108.195 ;
      RECT  78.02 108.995 77.88 103.425 ;
      RECT  78.91 103.885 78.62 103.585 ;
      RECT  74.28 114.705 74.51 113.435 ;
      RECT  74.74 109.055 74.91 103.425 ;
      RECT  75.12 108.995 75.26 103.425 ;
      RECT  78.63 114.705 78.86 113.435 ;
      RECT  78.23 109.055 78.4 103.425 ;
      RECT  77.88 108.995 78.02 103.425 ;
      RECT  80.33 98.395 80.47 102.165 ;
      RECT  82.65 98.395 82.79 102.165 ;
      RECT  74.28 113.435 74.51 114.705 ;
      RECT  78.63 113.435 78.86 114.705 ;
      RECT  34.46 61.73 34.6 63.705 ;
      RECT  33.1 61.73 33.24 63.705 ;
      RECT  34.46 65.68 34.6 63.705 ;
      RECT  33.1 65.68 33.24 63.705 ;
      RECT  41.02 61.57 41.27 63.74 ;
      RECT  38.9 61.58 39.14 63.74 ;
      RECT  44.33 61.73 44.47 63.705 ;
      RECT  42.97 61.73 43.11 63.705 ;
      RECT  41.02 61.57 41.27 63.74 ;
      RECT  44.33 61.73 44.47 63.705 ;
      RECT  38.9 61.58 39.14 63.74 ;
      RECT  42.97 61.73 43.11 63.705 ;
      RECT  41.02 65.84 41.27 63.67 ;
      RECT  38.9 65.83 39.14 63.67 ;
      RECT  44.33 65.68 44.47 63.705 ;
      RECT  42.97 65.68 43.11 63.705 ;
      RECT  41.02 65.84 41.27 63.67 ;
      RECT  44.33 65.68 44.47 63.705 ;
      RECT  38.9 65.83 39.14 63.67 ;
      RECT  42.97 65.68 43.11 63.705 ;
      RECT  41.02 65.52 41.27 67.69 ;
      RECT  38.9 65.53 39.14 67.69 ;
      RECT  44.33 65.68 44.47 67.655 ;
      RECT  42.97 65.68 43.11 67.655 ;
      RECT  41.02 65.52 41.27 67.69 ;
      RECT  44.33 65.68 44.47 67.655 ;
      RECT  38.9 65.53 39.14 67.69 ;
      RECT  42.97 65.68 43.11 67.655 ;
      RECT  41.02 69.79 41.27 67.62 ;
      RECT  38.9 69.78 39.14 67.62 ;
      RECT  44.33 69.63 44.47 67.655 ;
      RECT  42.97 69.63 43.11 67.655 ;
      RECT  41.02 69.79 41.27 67.62 ;
      RECT  44.33 69.63 44.47 67.655 ;
      RECT  38.9 69.78 39.14 67.62 ;
      RECT  42.97 69.63 43.11 67.655 ;
      RECT  30.92 62.555 31.18 62.875 ;
      RECT  31.32 64.535 31.58 64.855 ;
      RECT  34.46 73.58 34.6 75.555 ;
      RECT  33.1 73.58 33.24 75.555 ;
      RECT  34.46 77.53 34.6 75.555 ;
      RECT  33.1 77.53 33.24 75.555 ;
      RECT  41.02 73.42 41.27 75.59 ;
      RECT  38.9 73.43 39.14 75.59 ;
      RECT  44.33 73.58 44.47 75.555 ;
      RECT  42.97 73.58 43.11 75.555 ;
      RECT  41.02 73.42 41.27 75.59 ;
      RECT  44.33 73.58 44.47 75.555 ;
      RECT  38.9 73.43 39.14 75.59 ;
      RECT  42.97 73.58 43.11 75.555 ;
      RECT  41.02 77.69 41.27 75.52 ;
      RECT  38.9 77.68 39.14 75.52 ;
      RECT  44.33 77.53 44.47 75.555 ;
      RECT  42.97 77.53 43.11 75.555 ;
      RECT  41.02 77.69 41.27 75.52 ;
      RECT  44.33 77.53 44.47 75.555 ;
      RECT  38.9 77.68 39.14 75.52 ;
      RECT  42.97 77.53 43.11 75.555 ;
      RECT  41.02 77.37 41.27 79.54 ;
      RECT  38.9 77.38 39.14 79.54 ;
      RECT  44.33 77.53 44.47 79.505 ;
      RECT  42.97 77.53 43.11 79.505 ;
      RECT  41.02 77.37 41.27 79.54 ;
      RECT  44.33 77.53 44.47 79.505 ;
      RECT  38.9 77.38 39.14 79.54 ;
      RECT  42.97 77.53 43.11 79.505 ;
      RECT  41.02 81.64 41.27 79.47 ;
      RECT  38.9 81.63 39.14 79.47 ;
      RECT  44.33 81.48 44.47 79.505 ;
      RECT  42.97 81.48 43.11 79.505 ;
      RECT  41.02 81.64 41.27 79.47 ;
      RECT  44.33 81.48 44.47 79.505 ;
      RECT  38.9 81.63 39.14 79.47 ;
      RECT  42.97 81.48 43.11 79.505 ;
      RECT  30.92 74.405 31.18 74.725 ;
      RECT  31.32 76.385 31.58 76.705 ;
      RECT  52.09 61.57 52.34 63.74 ;
      RECT  49.97 61.58 50.21 63.74 ;
      RECT  55.4 61.73 55.54 63.705 ;
      RECT  54.04 61.73 54.18 63.705 ;
      RECT  52.09 61.57 52.34 63.74 ;
      RECT  55.4 61.73 55.54 63.705 ;
      RECT  49.97 61.58 50.21 63.74 ;
      RECT  54.04 61.73 54.18 63.705 ;
      RECT  52.09 65.84 52.34 63.67 ;
      RECT  49.97 65.83 50.21 63.67 ;
      RECT  55.4 65.68 55.54 63.705 ;
      RECT  54.04 65.68 54.18 63.705 ;
      RECT  52.09 65.84 52.34 63.67 ;
      RECT  55.4 65.68 55.54 63.705 ;
      RECT  49.97 65.83 50.21 63.67 ;
      RECT  54.04 65.68 54.18 63.705 ;
      RECT  52.09 65.52 52.34 67.69 ;
      RECT  49.97 65.53 50.21 67.69 ;
      RECT  55.4 65.68 55.54 67.655 ;
      RECT  54.04 65.68 54.18 67.655 ;
      RECT  52.09 65.52 52.34 67.69 ;
      RECT  55.4 65.68 55.54 67.655 ;
      RECT  49.97 65.53 50.21 67.69 ;
      RECT  54.04 65.68 54.18 67.655 ;
      RECT  52.09 69.79 52.34 67.62 ;
      RECT  49.97 69.78 50.21 67.62 ;
      RECT  55.4 69.63 55.54 67.655 ;
      RECT  54.04 69.63 54.18 67.655 ;
      RECT  52.09 69.79 52.34 67.62 ;
      RECT  55.4 69.63 55.54 67.655 ;
      RECT  49.97 69.78 50.21 67.62 ;
      RECT  54.04 69.63 54.18 67.655 ;
      RECT  52.09 69.47 52.34 71.64 ;
      RECT  49.97 69.48 50.21 71.64 ;
      RECT  55.4 69.63 55.54 71.605 ;
      RECT  54.04 69.63 54.18 71.605 ;
      RECT  52.09 69.47 52.34 71.64 ;
      RECT  55.4 69.63 55.54 71.605 ;
      RECT  49.97 69.48 50.21 71.64 ;
      RECT  54.04 69.63 54.18 71.605 ;
      RECT  52.09 73.74 52.34 71.57 ;
      RECT  49.97 73.73 50.21 71.57 ;
      RECT  55.4 73.58 55.54 71.605 ;
      RECT  54.04 73.58 54.18 71.605 ;
      RECT  52.09 73.74 52.34 71.57 ;
      RECT  55.4 73.58 55.54 71.605 ;
      RECT  49.97 73.73 50.21 71.57 ;
      RECT  54.04 73.58 54.18 71.605 ;
      RECT  52.09 73.42 52.34 75.59 ;
      RECT  49.97 73.43 50.21 75.59 ;
      RECT  55.4 73.58 55.54 75.555 ;
      RECT  54.04 73.58 54.18 75.555 ;
      RECT  52.09 73.42 52.34 75.59 ;
      RECT  55.4 73.58 55.54 75.555 ;
      RECT  49.97 73.43 50.21 75.59 ;
      RECT  54.04 73.58 54.18 75.555 ;
      RECT  52.09 77.69 52.34 75.52 ;
      RECT  49.97 77.68 50.21 75.52 ;
      RECT  55.4 77.53 55.54 75.555 ;
      RECT  54.04 77.53 54.18 75.555 ;
      RECT  52.09 77.69 52.34 75.52 ;
      RECT  55.4 77.53 55.54 75.555 ;
      RECT  49.97 77.68 50.21 75.52 ;
      RECT  54.04 77.53 54.18 75.555 ;
      RECT  52.09 77.37 52.34 79.54 ;
      RECT  49.97 77.38 50.21 79.54 ;
      RECT  55.4 77.53 55.54 79.505 ;
      RECT  54.04 77.53 54.18 79.505 ;
      RECT  52.09 77.37 52.34 79.54 ;
      RECT  55.4 77.53 55.54 79.505 ;
      RECT  49.97 77.38 50.21 79.54 ;
      RECT  54.04 77.53 54.18 79.505 ;
      RECT  52.09 81.64 52.34 79.47 ;
      RECT  49.97 81.63 50.21 79.47 ;
      RECT  55.4 81.48 55.54 79.505 ;
      RECT  54.04 81.48 54.18 79.505 ;
      RECT  52.09 81.64 52.34 79.47 ;
      RECT  55.4 81.48 55.54 79.505 ;
      RECT  49.97 81.63 50.21 79.47 ;
      RECT  54.04 81.48 54.18 79.505 ;
      RECT  52.09 81.32 52.34 83.49 ;
      RECT  49.97 81.33 50.21 83.49 ;
      RECT  55.4 81.48 55.54 83.455 ;
      RECT  54.04 81.48 54.18 83.455 ;
      RECT  52.09 81.32 52.34 83.49 ;
      RECT  55.4 81.48 55.54 83.455 ;
      RECT  49.97 81.33 50.21 83.49 ;
      RECT  54.04 81.48 54.18 83.455 ;
      RECT  52.09 85.59 52.34 83.42 ;
      RECT  49.97 85.58 50.21 83.42 ;
      RECT  55.4 85.43 55.54 83.455 ;
      RECT  54.04 85.43 54.18 83.455 ;
      RECT  52.09 85.59 52.34 83.42 ;
      RECT  55.4 85.43 55.54 83.455 ;
      RECT  49.97 85.58 50.21 83.42 ;
      RECT  54.04 85.43 54.18 83.455 ;
      RECT  52.09 85.27 52.34 87.44 ;
      RECT  49.97 85.28 50.21 87.44 ;
      RECT  55.4 85.43 55.54 87.405 ;
      RECT  54.04 85.43 54.18 87.405 ;
      RECT  52.09 85.27 52.34 87.44 ;
      RECT  55.4 85.43 55.54 87.405 ;
      RECT  49.97 85.28 50.21 87.44 ;
      RECT  54.04 85.43 54.18 87.405 ;
      RECT  52.09 89.54 52.34 87.37 ;
      RECT  49.97 89.53 50.21 87.37 ;
      RECT  55.4 89.38 55.54 87.405 ;
      RECT  54.04 89.38 54.18 87.405 ;
      RECT  52.09 89.54 52.34 87.37 ;
      RECT  55.4 89.38 55.54 87.405 ;
      RECT  49.97 89.53 50.21 87.37 ;
      RECT  54.04 89.38 54.18 87.405 ;
      RECT  52.09 89.22 52.34 91.39 ;
      RECT  49.97 89.23 50.21 91.39 ;
      RECT  55.4 89.38 55.54 91.355 ;
      RECT  54.04 89.38 54.18 91.355 ;
      RECT  52.09 89.22 52.34 91.39 ;
      RECT  55.4 89.38 55.54 91.355 ;
      RECT  49.97 89.23 50.21 91.39 ;
      RECT  54.04 89.38 54.18 91.355 ;
      RECT  52.09 93.49 52.34 91.32 ;
      RECT  49.97 93.48 50.21 91.32 ;
      RECT  55.4 93.33 55.54 91.355 ;
      RECT  54.04 93.33 54.18 91.355 ;
      RECT  52.09 93.49 52.34 91.32 ;
      RECT  55.4 93.33 55.54 91.355 ;
      RECT  49.97 93.48 50.21 91.32 ;
      RECT  54.04 93.33 54.18 91.355 ;
      RECT  28.84 61.73 28.98 81.48 ;
      RECT  29.24 61.73 29.38 81.48 ;
      RECT  29.64 61.73 29.78 81.48 ;
      RECT  30.04 61.73 30.18 81.48 ;
      RECT  59.7 61.425 59.95 63.595 ;
      RECT  57.58 61.435 57.82 63.595 ;
      RECT  64.33 61.585 64.47 63.56 ;
      RECT  61.84 61.585 61.98 63.56 ;
      RECT  59.7 61.425 59.95 63.595 ;
      RECT  64.33 61.585 64.47 63.56 ;
      RECT  57.58 61.435 57.82 63.595 ;
      RECT  61.84 61.585 61.98 63.56 ;
      RECT  59.7 65.695 59.95 63.525 ;
      RECT  57.58 65.685 57.82 63.525 ;
      RECT  64.33 65.535 64.47 63.56 ;
      RECT  61.84 65.535 61.98 63.56 ;
      RECT  59.7 65.695 59.95 63.525 ;
      RECT  64.33 65.535 64.47 63.56 ;
      RECT  57.58 65.685 57.82 63.525 ;
      RECT  61.84 65.535 61.98 63.56 ;
      RECT  59.7 65.375 59.95 67.545 ;
      RECT  57.58 65.385 57.82 67.545 ;
      RECT  64.33 65.535 64.47 67.51 ;
      RECT  61.84 65.535 61.98 67.51 ;
      RECT  59.7 65.375 59.95 67.545 ;
      RECT  64.33 65.535 64.47 67.51 ;
      RECT  57.58 65.385 57.82 67.545 ;
      RECT  61.84 65.535 61.98 67.51 ;
      RECT  59.7 69.645 59.95 67.475 ;
      RECT  57.58 69.635 57.82 67.475 ;
      RECT  64.33 69.485 64.47 67.51 ;
      RECT  61.84 69.485 61.98 67.51 ;
      RECT  59.7 69.645 59.95 67.475 ;
      RECT  64.33 69.485 64.47 67.51 ;
      RECT  57.58 69.635 57.82 67.475 ;
      RECT  61.84 69.485 61.98 67.51 ;
      RECT  59.7 69.325 59.95 71.495 ;
      RECT  57.58 69.335 57.82 71.495 ;
      RECT  64.33 69.485 64.47 71.46 ;
      RECT  61.84 69.485 61.98 71.46 ;
      RECT  59.7 69.325 59.95 71.495 ;
      RECT  64.33 69.485 64.47 71.46 ;
      RECT  57.58 69.335 57.82 71.495 ;
      RECT  61.84 69.485 61.98 71.46 ;
      RECT  59.7 73.595 59.95 71.425 ;
      RECT  57.58 73.585 57.82 71.425 ;
      RECT  64.33 73.435 64.47 71.46 ;
      RECT  61.84 73.435 61.98 71.46 ;
      RECT  59.7 73.595 59.95 71.425 ;
      RECT  64.33 73.435 64.47 71.46 ;
      RECT  57.58 73.585 57.82 71.425 ;
      RECT  61.84 73.435 61.98 71.46 ;
      RECT  59.7 73.275 59.95 75.445 ;
      RECT  57.58 73.285 57.82 75.445 ;
      RECT  64.33 73.435 64.47 75.41 ;
      RECT  61.84 73.435 61.98 75.41 ;
      RECT  59.7 73.275 59.95 75.445 ;
      RECT  64.33 73.435 64.47 75.41 ;
      RECT  57.58 73.285 57.82 75.445 ;
      RECT  61.84 73.435 61.98 75.41 ;
      RECT  59.7 77.545 59.95 75.375 ;
      RECT  57.58 77.535 57.82 75.375 ;
      RECT  64.33 77.385 64.47 75.41 ;
      RECT  61.84 77.385 61.98 75.41 ;
      RECT  59.7 77.545 59.95 75.375 ;
      RECT  64.33 77.385 64.47 75.41 ;
      RECT  57.58 77.535 57.82 75.375 ;
      RECT  61.84 77.385 61.98 75.41 ;
      RECT  59.7 77.225 59.95 79.395 ;
      RECT  57.58 77.235 57.82 79.395 ;
      RECT  64.33 77.385 64.47 79.36 ;
      RECT  61.84 77.385 61.98 79.36 ;
      RECT  59.7 77.225 59.95 79.395 ;
      RECT  64.33 77.385 64.47 79.36 ;
      RECT  57.58 77.235 57.82 79.395 ;
      RECT  61.84 77.385 61.98 79.36 ;
      RECT  59.7 81.495 59.95 79.325 ;
      RECT  57.58 81.485 57.82 79.325 ;
      RECT  64.33 81.335 64.47 79.36 ;
      RECT  61.84 81.335 61.98 79.36 ;
      RECT  59.7 81.495 59.95 79.325 ;
      RECT  64.33 81.335 64.47 79.36 ;
      RECT  57.58 81.485 57.82 79.325 ;
      RECT  61.84 81.335 61.98 79.36 ;
      RECT  59.7 81.175 59.95 83.345 ;
      RECT  57.58 81.185 57.82 83.345 ;
      RECT  64.33 81.335 64.47 83.31 ;
      RECT  61.84 81.335 61.98 83.31 ;
      RECT  59.7 81.175 59.95 83.345 ;
      RECT  64.33 81.335 64.47 83.31 ;
      RECT  57.58 81.185 57.82 83.345 ;
      RECT  61.84 81.335 61.98 83.31 ;
      RECT  59.7 85.445 59.95 83.275 ;
      RECT  57.58 85.435 57.82 83.275 ;
      RECT  64.33 85.285 64.47 83.31 ;
      RECT  61.84 85.285 61.98 83.31 ;
      RECT  59.7 85.445 59.95 83.275 ;
      RECT  64.33 85.285 64.47 83.31 ;
      RECT  57.58 85.435 57.82 83.275 ;
      RECT  61.84 85.285 61.98 83.31 ;
      RECT  59.7 85.125 59.95 87.295 ;
      RECT  57.58 85.135 57.82 87.295 ;
      RECT  64.33 85.285 64.47 87.26 ;
      RECT  61.84 85.285 61.98 87.26 ;
      RECT  59.7 85.125 59.95 87.295 ;
      RECT  64.33 85.285 64.47 87.26 ;
      RECT  57.58 85.135 57.82 87.295 ;
      RECT  61.84 85.285 61.98 87.26 ;
      RECT  59.7 89.395 59.95 87.225 ;
      RECT  57.58 89.385 57.82 87.225 ;
      RECT  64.33 89.235 64.47 87.26 ;
      RECT  61.84 89.235 61.98 87.26 ;
      RECT  59.7 89.395 59.95 87.225 ;
      RECT  64.33 89.235 64.47 87.26 ;
      RECT  57.58 89.385 57.82 87.225 ;
      RECT  61.84 89.235 61.98 87.26 ;
      RECT  59.7 89.075 59.95 91.245 ;
      RECT  57.58 89.085 57.82 91.245 ;
      RECT  64.33 89.235 64.47 91.21 ;
      RECT  61.84 89.235 61.98 91.21 ;
      RECT  59.7 89.075 59.95 91.245 ;
      RECT  64.33 89.235 64.47 91.21 ;
      RECT  57.58 89.085 57.82 91.245 ;
      RECT  61.84 89.235 61.98 91.21 ;
      RECT  59.7 93.345 59.95 91.175 ;
      RECT  57.58 93.335 57.82 91.175 ;
      RECT  64.33 93.185 64.47 91.21 ;
      RECT  61.84 93.185 61.98 91.21 ;
      RECT  59.7 93.345 59.95 91.175 ;
      RECT  64.33 93.185 64.47 91.21 ;
      RECT  57.58 93.335 57.82 91.175 ;
      RECT  61.84 93.185 61.98 91.21 ;
      RECT  64.33 61.585 64.47 93.185 ;
      RECT  59.755 61.425 59.895 93.185 ;
      RECT  61.84 61.585 61.98 93.185 ;
      RECT  57.63 61.435 57.77 93.185 ;
      RECT  28.84 61.73 28.98 81.48 ;
      RECT  29.24 61.73 29.38 81.48 ;
      RECT  29.64 61.73 29.78 81.48 ;
      RECT  30.04 61.73 30.18 81.48 ;
      RECT  119.3 61.73 119.16 63.705 ;
      RECT  120.66 61.73 120.52 63.705 ;
      RECT  119.3 65.68 119.16 63.705 ;
      RECT  120.66 65.68 120.52 63.705 ;
      RECT  112.74 61.57 112.49 63.74 ;
      RECT  114.86 61.58 114.62 63.74 ;
      RECT  109.43 61.73 109.29 63.705 ;
      RECT  110.79 61.73 110.65 63.705 ;
      RECT  112.74 61.57 112.49 63.74 ;
      RECT  109.43 61.73 109.29 63.705 ;
      RECT  114.86 61.58 114.62 63.74 ;
      RECT  110.79 61.73 110.65 63.705 ;
      RECT  112.74 65.84 112.49 63.67 ;
      RECT  114.86 65.83 114.62 63.67 ;
      RECT  109.43 65.68 109.29 63.705 ;
      RECT  110.79 65.68 110.65 63.705 ;
      RECT  112.74 65.84 112.49 63.67 ;
      RECT  109.43 65.68 109.29 63.705 ;
      RECT  114.86 65.83 114.62 63.67 ;
      RECT  110.79 65.68 110.65 63.705 ;
      RECT  112.74 65.52 112.49 67.69 ;
      RECT  114.86 65.53 114.62 67.69 ;
      RECT  109.43 65.68 109.29 67.655 ;
      RECT  110.79 65.68 110.65 67.655 ;
      RECT  112.74 65.52 112.49 67.69 ;
      RECT  109.43 65.68 109.29 67.655 ;
      RECT  114.86 65.53 114.62 67.69 ;
      RECT  110.79 65.68 110.65 67.655 ;
      RECT  112.74 69.79 112.49 67.62 ;
      RECT  114.86 69.78 114.62 67.62 ;
      RECT  109.43 69.63 109.29 67.655 ;
      RECT  110.79 69.63 110.65 67.655 ;
      RECT  112.74 69.79 112.49 67.62 ;
      RECT  109.43 69.63 109.29 67.655 ;
      RECT  114.86 69.78 114.62 67.62 ;
      RECT  110.79 69.63 110.65 67.655 ;
      RECT  122.84 62.555 122.58 62.875 ;
      RECT  122.44 64.535 122.18 64.855 ;
      RECT  119.3 73.58 119.16 75.555 ;
      RECT  120.66 73.58 120.52 75.555 ;
      RECT  119.3 77.53 119.16 75.555 ;
      RECT  120.66 77.53 120.52 75.555 ;
      RECT  112.74 73.42 112.49 75.59 ;
      RECT  114.86 73.43 114.62 75.59 ;
      RECT  109.43 73.58 109.29 75.555 ;
      RECT  110.79 73.58 110.65 75.555 ;
      RECT  112.74 73.42 112.49 75.59 ;
      RECT  109.43 73.58 109.29 75.555 ;
      RECT  114.86 73.43 114.62 75.59 ;
      RECT  110.79 73.58 110.65 75.555 ;
      RECT  112.74 77.69 112.49 75.52 ;
      RECT  114.86 77.68 114.62 75.52 ;
      RECT  109.43 77.53 109.29 75.555 ;
      RECT  110.79 77.53 110.65 75.555 ;
      RECT  112.74 77.69 112.49 75.52 ;
      RECT  109.43 77.53 109.29 75.555 ;
      RECT  114.86 77.68 114.62 75.52 ;
      RECT  110.79 77.53 110.65 75.555 ;
      RECT  112.74 77.37 112.49 79.54 ;
      RECT  114.86 77.38 114.62 79.54 ;
      RECT  109.43 77.53 109.29 79.505 ;
      RECT  110.79 77.53 110.65 79.505 ;
      RECT  112.74 77.37 112.49 79.54 ;
      RECT  109.43 77.53 109.29 79.505 ;
      RECT  114.86 77.38 114.62 79.54 ;
      RECT  110.79 77.53 110.65 79.505 ;
      RECT  112.74 81.64 112.49 79.47 ;
      RECT  114.86 81.63 114.62 79.47 ;
      RECT  109.43 81.48 109.29 79.505 ;
      RECT  110.79 81.48 110.65 79.505 ;
      RECT  112.74 81.64 112.49 79.47 ;
      RECT  109.43 81.48 109.29 79.505 ;
      RECT  114.86 81.63 114.62 79.47 ;
      RECT  110.79 81.48 110.65 79.505 ;
      RECT  122.84 74.405 122.58 74.725 ;
      RECT  122.44 76.385 122.18 76.705 ;
      RECT  101.67 61.57 101.42 63.74 ;
      RECT  103.79 61.58 103.55 63.74 ;
      RECT  98.36 61.73 98.22 63.705 ;
      RECT  99.72 61.73 99.58 63.705 ;
      RECT  101.67 61.57 101.42 63.74 ;
      RECT  98.36 61.73 98.22 63.705 ;
      RECT  103.79 61.58 103.55 63.74 ;
      RECT  99.72 61.73 99.58 63.705 ;
      RECT  101.67 65.84 101.42 63.67 ;
      RECT  103.79 65.83 103.55 63.67 ;
      RECT  98.36 65.68 98.22 63.705 ;
      RECT  99.72 65.68 99.58 63.705 ;
      RECT  101.67 65.84 101.42 63.67 ;
      RECT  98.36 65.68 98.22 63.705 ;
      RECT  103.79 65.83 103.55 63.67 ;
      RECT  99.72 65.68 99.58 63.705 ;
      RECT  101.67 65.52 101.42 67.69 ;
      RECT  103.79 65.53 103.55 67.69 ;
      RECT  98.36 65.68 98.22 67.655 ;
      RECT  99.72 65.68 99.58 67.655 ;
      RECT  101.67 65.52 101.42 67.69 ;
      RECT  98.36 65.68 98.22 67.655 ;
      RECT  103.79 65.53 103.55 67.69 ;
      RECT  99.72 65.68 99.58 67.655 ;
      RECT  101.67 69.79 101.42 67.62 ;
      RECT  103.79 69.78 103.55 67.62 ;
      RECT  98.36 69.63 98.22 67.655 ;
      RECT  99.72 69.63 99.58 67.655 ;
      RECT  101.67 69.79 101.42 67.62 ;
      RECT  98.36 69.63 98.22 67.655 ;
      RECT  103.79 69.78 103.55 67.62 ;
      RECT  99.72 69.63 99.58 67.655 ;
      RECT  101.67 69.47 101.42 71.64 ;
      RECT  103.79 69.48 103.55 71.64 ;
      RECT  98.36 69.63 98.22 71.605 ;
      RECT  99.72 69.63 99.58 71.605 ;
      RECT  101.67 69.47 101.42 71.64 ;
      RECT  98.36 69.63 98.22 71.605 ;
      RECT  103.79 69.48 103.55 71.64 ;
      RECT  99.72 69.63 99.58 71.605 ;
      RECT  101.67 73.74 101.42 71.57 ;
      RECT  103.79 73.73 103.55 71.57 ;
      RECT  98.36 73.58 98.22 71.605 ;
      RECT  99.72 73.58 99.58 71.605 ;
      RECT  101.67 73.74 101.42 71.57 ;
      RECT  98.36 73.58 98.22 71.605 ;
      RECT  103.79 73.73 103.55 71.57 ;
      RECT  99.72 73.58 99.58 71.605 ;
      RECT  101.67 73.42 101.42 75.59 ;
      RECT  103.79 73.43 103.55 75.59 ;
      RECT  98.36 73.58 98.22 75.555 ;
      RECT  99.72 73.58 99.58 75.555 ;
      RECT  101.67 73.42 101.42 75.59 ;
      RECT  98.36 73.58 98.22 75.555 ;
      RECT  103.79 73.43 103.55 75.59 ;
      RECT  99.72 73.58 99.58 75.555 ;
      RECT  101.67 77.69 101.42 75.52 ;
      RECT  103.79 77.68 103.55 75.52 ;
      RECT  98.36 77.53 98.22 75.555 ;
      RECT  99.72 77.53 99.58 75.555 ;
      RECT  101.67 77.69 101.42 75.52 ;
      RECT  98.36 77.53 98.22 75.555 ;
      RECT  103.79 77.68 103.55 75.52 ;
      RECT  99.72 77.53 99.58 75.555 ;
      RECT  101.67 77.37 101.42 79.54 ;
      RECT  103.79 77.38 103.55 79.54 ;
      RECT  98.36 77.53 98.22 79.505 ;
      RECT  99.72 77.53 99.58 79.505 ;
      RECT  101.67 77.37 101.42 79.54 ;
      RECT  98.36 77.53 98.22 79.505 ;
      RECT  103.79 77.38 103.55 79.54 ;
      RECT  99.72 77.53 99.58 79.505 ;
      RECT  101.67 81.64 101.42 79.47 ;
      RECT  103.79 81.63 103.55 79.47 ;
      RECT  98.36 81.48 98.22 79.505 ;
      RECT  99.72 81.48 99.58 79.505 ;
      RECT  101.67 81.64 101.42 79.47 ;
      RECT  98.36 81.48 98.22 79.505 ;
      RECT  103.79 81.63 103.55 79.47 ;
      RECT  99.72 81.48 99.58 79.505 ;
      RECT  101.67 81.32 101.42 83.49 ;
      RECT  103.79 81.33 103.55 83.49 ;
      RECT  98.36 81.48 98.22 83.455 ;
      RECT  99.72 81.48 99.58 83.455 ;
      RECT  101.67 81.32 101.42 83.49 ;
      RECT  98.36 81.48 98.22 83.455 ;
      RECT  103.79 81.33 103.55 83.49 ;
      RECT  99.72 81.48 99.58 83.455 ;
      RECT  101.67 85.59 101.42 83.42 ;
      RECT  103.79 85.58 103.55 83.42 ;
      RECT  98.36 85.43 98.22 83.455 ;
      RECT  99.72 85.43 99.58 83.455 ;
      RECT  101.67 85.59 101.42 83.42 ;
      RECT  98.36 85.43 98.22 83.455 ;
      RECT  103.79 85.58 103.55 83.42 ;
      RECT  99.72 85.43 99.58 83.455 ;
      RECT  101.67 85.27 101.42 87.44 ;
      RECT  103.79 85.28 103.55 87.44 ;
      RECT  98.36 85.43 98.22 87.405 ;
      RECT  99.72 85.43 99.58 87.405 ;
      RECT  101.67 85.27 101.42 87.44 ;
      RECT  98.36 85.43 98.22 87.405 ;
      RECT  103.79 85.28 103.55 87.44 ;
      RECT  99.72 85.43 99.58 87.405 ;
      RECT  101.67 89.54 101.42 87.37 ;
      RECT  103.79 89.53 103.55 87.37 ;
      RECT  98.36 89.38 98.22 87.405 ;
      RECT  99.72 89.38 99.58 87.405 ;
      RECT  101.67 89.54 101.42 87.37 ;
      RECT  98.36 89.38 98.22 87.405 ;
      RECT  103.79 89.53 103.55 87.37 ;
      RECT  99.72 89.38 99.58 87.405 ;
      RECT  101.67 89.22 101.42 91.39 ;
      RECT  103.79 89.23 103.55 91.39 ;
      RECT  98.36 89.38 98.22 91.355 ;
      RECT  99.72 89.38 99.58 91.355 ;
      RECT  101.67 89.22 101.42 91.39 ;
      RECT  98.36 89.38 98.22 91.355 ;
      RECT  103.79 89.23 103.55 91.39 ;
      RECT  99.72 89.38 99.58 91.355 ;
      RECT  101.67 93.49 101.42 91.32 ;
      RECT  103.79 93.48 103.55 91.32 ;
      RECT  98.36 93.33 98.22 91.355 ;
      RECT  99.72 93.33 99.58 91.355 ;
      RECT  101.67 93.49 101.42 91.32 ;
      RECT  98.36 93.33 98.22 91.355 ;
      RECT  103.79 93.48 103.55 91.32 ;
      RECT  99.72 93.33 99.58 91.355 ;
      RECT  124.92 61.73 124.78 81.48 ;
      RECT  124.52 61.73 124.38 81.48 ;
      RECT  124.12 61.73 123.98 81.48 ;
      RECT  123.72 61.73 123.58 81.48 ;
      RECT  94.06 61.425 93.81 63.595 ;
      RECT  96.18 61.435 95.94 63.595 ;
      RECT  89.43 61.585 89.29 63.56 ;
      RECT  91.92 61.585 91.78 63.56 ;
      RECT  94.06 61.425 93.81 63.595 ;
      RECT  89.43 61.585 89.29 63.56 ;
      RECT  96.18 61.435 95.94 63.595 ;
      RECT  91.92 61.585 91.78 63.56 ;
      RECT  94.06 65.695 93.81 63.525 ;
      RECT  96.18 65.685 95.94 63.525 ;
      RECT  89.43 65.535 89.29 63.56 ;
      RECT  91.92 65.535 91.78 63.56 ;
      RECT  94.06 65.695 93.81 63.525 ;
      RECT  89.43 65.535 89.29 63.56 ;
      RECT  96.18 65.685 95.94 63.525 ;
      RECT  91.92 65.535 91.78 63.56 ;
      RECT  94.06 65.375 93.81 67.545 ;
      RECT  96.18 65.385 95.94 67.545 ;
      RECT  89.43 65.535 89.29 67.51 ;
      RECT  91.92 65.535 91.78 67.51 ;
      RECT  94.06 65.375 93.81 67.545 ;
      RECT  89.43 65.535 89.29 67.51 ;
      RECT  96.18 65.385 95.94 67.545 ;
      RECT  91.92 65.535 91.78 67.51 ;
      RECT  94.06 69.645 93.81 67.475 ;
      RECT  96.18 69.635 95.94 67.475 ;
      RECT  89.43 69.485 89.29 67.51 ;
      RECT  91.92 69.485 91.78 67.51 ;
      RECT  94.06 69.645 93.81 67.475 ;
      RECT  89.43 69.485 89.29 67.51 ;
      RECT  96.18 69.635 95.94 67.475 ;
      RECT  91.92 69.485 91.78 67.51 ;
      RECT  94.06 69.325 93.81 71.495 ;
      RECT  96.18 69.335 95.94 71.495 ;
      RECT  89.43 69.485 89.29 71.46 ;
      RECT  91.92 69.485 91.78 71.46 ;
      RECT  94.06 69.325 93.81 71.495 ;
      RECT  89.43 69.485 89.29 71.46 ;
      RECT  96.18 69.335 95.94 71.495 ;
      RECT  91.92 69.485 91.78 71.46 ;
      RECT  94.06 73.595 93.81 71.425 ;
      RECT  96.18 73.585 95.94 71.425 ;
      RECT  89.43 73.435 89.29 71.46 ;
      RECT  91.92 73.435 91.78 71.46 ;
      RECT  94.06 73.595 93.81 71.425 ;
      RECT  89.43 73.435 89.29 71.46 ;
      RECT  96.18 73.585 95.94 71.425 ;
      RECT  91.92 73.435 91.78 71.46 ;
      RECT  94.06 73.275 93.81 75.445 ;
      RECT  96.18 73.285 95.94 75.445 ;
      RECT  89.43 73.435 89.29 75.41 ;
      RECT  91.92 73.435 91.78 75.41 ;
      RECT  94.06 73.275 93.81 75.445 ;
      RECT  89.43 73.435 89.29 75.41 ;
      RECT  96.18 73.285 95.94 75.445 ;
      RECT  91.92 73.435 91.78 75.41 ;
      RECT  94.06 77.545 93.81 75.375 ;
      RECT  96.18 77.535 95.94 75.375 ;
      RECT  89.43 77.385 89.29 75.41 ;
      RECT  91.92 77.385 91.78 75.41 ;
      RECT  94.06 77.545 93.81 75.375 ;
      RECT  89.43 77.385 89.29 75.41 ;
      RECT  96.18 77.535 95.94 75.375 ;
      RECT  91.92 77.385 91.78 75.41 ;
      RECT  94.06 77.225 93.81 79.395 ;
      RECT  96.18 77.235 95.94 79.395 ;
      RECT  89.43 77.385 89.29 79.36 ;
      RECT  91.92 77.385 91.78 79.36 ;
      RECT  94.06 77.225 93.81 79.395 ;
      RECT  89.43 77.385 89.29 79.36 ;
      RECT  96.18 77.235 95.94 79.395 ;
      RECT  91.92 77.385 91.78 79.36 ;
      RECT  94.06 81.495 93.81 79.325 ;
      RECT  96.18 81.485 95.94 79.325 ;
      RECT  89.43 81.335 89.29 79.36 ;
      RECT  91.92 81.335 91.78 79.36 ;
      RECT  94.06 81.495 93.81 79.325 ;
      RECT  89.43 81.335 89.29 79.36 ;
      RECT  96.18 81.485 95.94 79.325 ;
      RECT  91.92 81.335 91.78 79.36 ;
      RECT  94.06 81.175 93.81 83.345 ;
      RECT  96.18 81.185 95.94 83.345 ;
      RECT  89.43 81.335 89.29 83.31 ;
      RECT  91.92 81.335 91.78 83.31 ;
      RECT  94.06 81.175 93.81 83.345 ;
      RECT  89.43 81.335 89.29 83.31 ;
      RECT  96.18 81.185 95.94 83.345 ;
      RECT  91.92 81.335 91.78 83.31 ;
      RECT  94.06 85.445 93.81 83.275 ;
      RECT  96.18 85.435 95.94 83.275 ;
      RECT  89.43 85.285 89.29 83.31 ;
      RECT  91.92 85.285 91.78 83.31 ;
      RECT  94.06 85.445 93.81 83.275 ;
      RECT  89.43 85.285 89.29 83.31 ;
      RECT  96.18 85.435 95.94 83.275 ;
      RECT  91.92 85.285 91.78 83.31 ;
      RECT  94.06 85.125 93.81 87.295 ;
      RECT  96.18 85.135 95.94 87.295 ;
      RECT  89.43 85.285 89.29 87.26 ;
      RECT  91.92 85.285 91.78 87.26 ;
      RECT  94.06 85.125 93.81 87.295 ;
      RECT  89.43 85.285 89.29 87.26 ;
      RECT  96.18 85.135 95.94 87.295 ;
      RECT  91.92 85.285 91.78 87.26 ;
      RECT  94.06 89.395 93.81 87.225 ;
      RECT  96.18 89.385 95.94 87.225 ;
      RECT  89.43 89.235 89.29 87.26 ;
      RECT  91.92 89.235 91.78 87.26 ;
      RECT  94.06 89.395 93.81 87.225 ;
      RECT  89.43 89.235 89.29 87.26 ;
      RECT  96.18 89.385 95.94 87.225 ;
      RECT  91.92 89.235 91.78 87.26 ;
      RECT  94.06 89.075 93.81 91.245 ;
      RECT  96.18 89.085 95.94 91.245 ;
      RECT  89.43 89.235 89.29 91.21 ;
      RECT  91.92 89.235 91.78 91.21 ;
      RECT  94.06 89.075 93.81 91.245 ;
      RECT  89.43 89.235 89.29 91.21 ;
      RECT  96.18 89.085 95.94 91.245 ;
      RECT  91.92 89.235 91.78 91.21 ;
      RECT  94.06 93.345 93.81 91.175 ;
      RECT  96.18 93.335 95.94 91.175 ;
      RECT  89.43 93.185 89.29 91.21 ;
      RECT  91.92 93.185 91.78 91.21 ;
      RECT  94.06 93.345 93.81 91.175 ;
      RECT  89.43 93.185 89.29 91.21 ;
      RECT  96.18 93.335 95.94 91.175 ;
      RECT  91.92 93.185 91.78 91.21 ;
      RECT  89.43 61.585 89.29 93.185 ;
      RECT  94.005 61.425 93.865 93.185 ;
      RECT  91.92 61.585 91.78 93.185 ;
      RECT  96.13 61.435 95.99 93.185 ;
      RECT  124.92 61.73 124.78 81.48 ;
      RECT  124.52 61.73 124.38 81.48 ;
      RECT  124.12 61.73 123.98 81.48 ;
      RECT  123.72 61.73 123.58 81.48 ;
      RECT  74.28 40.065 74.51 41.335 ;
      RECT  78.63 40.065 78.86 41.335 ;
      RECT  74.28 113.435 74.51 114.705 ;
      RECT  78.63 113.435 78.86 114.705 ;
      RECT  75.035 28.77 75.335 29.05 ;
      RECT  77.805 28.77 78.105 29.05 ;
      RECT  28.84 61.73 28.98 81.48 ;
      RECT  29.24 61.73 29.38 81.48 ;
      RECT  29.64 61.73 29.78 81.48 ;
      RECT  30.04 61.73 30.18 81.48 ;
      RECT  124.78 61.73 124.92 81.48 ;
      RECT  124.38 61.73 124.52 81.48 ;
      RECT  123.98 61.73 124.12 81.48 ;
      RECT  123.58 61.73 123.72 81.48 ;
      RECT  1.185 3.38 1.475 3.41 ;
      RECT  0.86 1.61 1.03 2.58 ;
      RECT  5.16 1.38 5.45 1.61 ;
      RECT  3.855 1.38 4.145 1.61 ;
      RECT  2.575 2.455 2.745 3.735 ;
      RECT  0.8 4.18 1.09 4.41 ;
      RECT  0.8 2.58 1.09 2.81 ;
      RECT  2.525 4.01 2.795 4.055 ;
      RECT  2.525 2.41 2.795 2.455 ;
      RECT  5.16 4.18 5.45 4.41 ;
      RECT  5.16 2.58 5.45 2.81 ;
      RECT  2.105 4.18 2.395 4.41 ;
      RECT  0.86 2.81 1.03 4.18 ;
      RECT  0.8 1.38 1.09 1.61 ;
      RECT  1.185 3.58 1.475 3.61 ;
      RECT  5.22 2.81 5.39 4.18 ;
      RECT  6.09 3.32 6.42 3.58 ;
      RECT  3.915 1.61 4.085 4.18 ;
      RECT  1.185 3.41 2.335 3.58 ;
      RECT  1.365 2.965 1.695 3.225 ;
      RECT  6.11 4.18 6.4 4.41 ;
      RECT  5.7 2.565 6.03 2.825 ;
      RECT  2.165 3.58 2.335 4.18 ;
      RECT  2.525 3.735 2.795 3.78 ;
      RECT  2.525 2.135 2.795 2.18 ;
      RECT  3.855 4.18 4.145 4.41 ;
      RECT  2.515 3.78 2.805 4.01 ;
      RECT  2.515 2.18 2.805 2.41 ;
      RECT  2.105 1.38 2.395 1.61 ;
      RECT  6.17 3.58 6.34 4.18 ;
      RECT  5.22 1.61 5.39 2.58 ;
      RECT  6.17 1.61 6.34 3.32 ;
      RECT  6.11 1.38 6.4 1.61 ;
      RECT  2.165 1.61 2.335 3.41 ;
      RECT  1.185 11.31 1.475 11.28 ;
      RECT  0.86 13.08 1.03 12.11 ;
      RECT  5.16 13.31 5.45 13.08 ;
      RECT  3.855 13.31 4.145 13.08 ;
      RECT  2.575 12.235 2.745 10.955 ;
      RECT  0.8 10.51 1.09 10.28 ;
      RECT  0.8 12.11 1.09 11.88 ;
      RECT  2.525 10.68 2.795 10.635 ;
      RECT  2.525 12.28 2.795 12.235 ;
      RECT  5.16 10.51 5.45 10.28 ;
      RECT  5.16 12.11 5.45 11.88 ;
      RECT  2.105 10.51 2.395 10.28 ;
      RECT  0.86 11.88 1.03 10.51 ;
      RECT  0.8 13.31 1.09 13.08 ;
      RECT  1.185 11.11 1.475 11.08 ;
      RECT  5.22 11.88 5.39 10.51 ;
      RECT  6.09 11.37 6.42 11.11 ;
      RECT  3.915 13.08 4.085 10.51 ;
      RECT  1.185 11.28 2.335 11.11 ;
      RECT  1.365 11.725 1.695 11.465 ;
      RECT  6.11 10.51 6.4 10.28 ;
      RECT  5.7 12.125 6.03 11.865 ;
      RECT  2.165 11.11 2.335 10.51 ;
      RECT  2.525 10.955 2.795 10.91 ;
      RECT  2.525 12.555 2.795 12.51 ;
      RECT  3.855 10.51 4.145 10.28 ;
      RECT  2.515 10.91 2.805 10.68 ;
      RECT  2.515 12.51 2.805 12.28 ;
      RECT  2.105 13.31 2.395 13.08 ;
      RECT  6.17 11.11 6.34 10.51 ;
      RECT  5.22 13.08 5.39 12.11 ;
      RECT  6.17 13.08 6.34 11.37 ;
      RECT  6.11 13.31 6.4 13.08 ;
      RECT  2.165 13.08 2.335 11.28 ;
      RECT  151.465 137.25 151.175 137.22 ;
      RECT  151.79 139.02 151.62 138.05 ;
      RECT  147.49 139.25 147.2 139.02 ;
      RECT  148.795 139.25 148.505 139.02 ;
      RECT  150.075 138.175 149.905 136.895 ;
      RECT  151.85 136.45 151.56 136.22 ;
      RECT  151.85 138.05 151.56 137.82 ;
      RECT  150.125 136.62 149.855 136.575 ;
      RECT  150.125 138.22 149.855 138.175 ;
      RECT  147.49 136.45 147.2 136.22 ;
      RECT  147.49 138.05 147.2 137.82 ;
      RECT  150.545 136.45 150.255 136.22 ;
      RECT  151.79 137.82 151.62 136.45 ;
      RECT  151.85 139.25 151.56 139.02 ;
      RECT  151.465 137.05 151.175 137.02 ;
      RECT  147.43 137.82 147.26 136.45 ;
      RECT  146.56 137.31 146.23 137.05 ;
      RECT  148.735 139.02 148.565 136.45 ;
      RECT  151.465 137.22 150.315 137.05 ;
      RECT  151.285 137.665 150.955 137.405 ;
      RECT  146.54 136.45 146.25 136.22 ;
      RECT  146.95 138.065 146.62 137.805 ;
      RECT  150.485 137.05 150.315 136.45 ;
      RECT  150.125 136.895 149.855 136.85 ;
      RECT  150.125 138.495 149.855 138.45 ;
      RECT  148.795 136.45 148.505 136.22 ;
      RECT  150.135 136.85 149.845 136.62 ;
      RECT  150.135 138.45 149.845 138.22 ;
      RECT  150.545 139.25 150.255 139.02 ;
      RECT  146.48 137.05 146.31 136.45 ;
      RECT  147.43 139.02 147.26 138.05 ;
      RECT  146.48 139.02 146.31 137.31 ;
      RECT  146.54 139.25 146.25 139.02 ;
      RECT  150.485 139.02 150.315 137.22 ;
      RECT  22.575 111.94 22.865 111.97 ;
      RECT  22.25 110.17 22.42 111.14 ;
      RECT  26.55 109.94 26.84 110.17 ;
      RECT  25.245 109.94 25.535 110.17 ;
      RECT  23.965 111.015 24.135 112.295 ;
      RECT  22.19 112.74 22.48 112.97 ;
      RECT  22.19 111.14 22.48 111.37 ;
      RECT  23.915 112.57 24.185 112.615 ;
      RECT  23.915 110.97 24.185 111.015 ;
      RECT  26.55 112.74 26.84 112.97 ;
      RECT  26.55 111.14 26.84 111.37 ;
      RECT  23.495 112.74 23.785 112.97 ;
      RECT  22.25 111.37 22.42 112.74 ;
      RECT  22.19 109.94 22.48 110.17 ;
      RECT  22.575 112.14 22.865 112.17 ;
      RECT  26.61 111.37 26.78 112.74 ;
      RECT  27.48 111.88 27.81 112.14 ;
      RECT  25.305 110.17 25.475 112.74 ;
      RECT  22.575 111.97 23.725 112.14 ;
      RECT  22.755 111.525 23.085 111.785 ;
      RECT  27.5 112.74 27.79 112.97 ;
      RECT  27.09 111.125 27.42 111.385 ;
      RECT  23.555 112.14 23.725 112.74 ;
      RECT  23.915 112.295 24.185 112.34 ;
      RECT  23.915 110.695 24.185 110.74 ;
      RECT  25.245 112.74 25.535 112.97 ;
      RECT  23.905 112.34 24.195 112.57 ;
      RECT  23.905 110.74 24.195 110.97 ;
      RECT  23.495 109.94 23.785 110.17 ;
      RECT  27.56 112.14 27.73 112.74 ;
      RECT  26.61 110.17 26.78 111.14 ;
      RECT  27.56 110.17 27.73 111.88 ;
      RECT  27.5 109.94 27.79 110.17 ;
      RECT  23.555 110.17 23.725 111.97 ;
      RECT  22.575 119.87 22.865 119.84 ;
      RECT  22.25 121.64 22.42 120.67 ;
      RECT  26.55 121.87 26.84 121.64 ;
      RECT  25.245 121.87 25.535 121.64 ;
      RECT  23.965 120.795 24.135 119.515 ;
      RECT  22.19 119.07 22.48 118.84 ;
      RECT  22.19 120.67 22.48 120.44 ;
      RECT  23.915 119.24 24.185 119.195 ;
      RECT  23.915 120.84 24.185 120.795 ;
      RECT  26.55 119.07 26.84 118.84 ;
      RECT  26.55 120.67 26.84 120.44 ;
      RECT  23.495 119.07 23.785 118.84 ;
      RECT  22.25 120.44 22.42 119.07 ;
      RECT  22.19 121.87 22.48 121.64 ;
      RECT  22.575 119.67 22.865 119.64 ;
      RECT  26.61 120.44 26.78 119.07 ;
      RECT  27.48 119.93 27.81 119.67 ;
      RECT  25.305 121.64 25.475 119.07 ;
      RECT  22.575 119.84 23.725 119.67 ;
      RECT  22.755 120.285 23.085 120.025 ;
      RECT  27.5 119.07 27.79 118.84 ;
      RECT  27.09 120.685 27.42 120.425 ;
      RECT  23.555 119.67 23.725 119.07 ;
      RECT  23.915 119.515 24.185 119.47 ;
      RECT  23.915 121.115 24.185 121.07 ;
      RECT  25.245 119.07 25.535 118.84 ;
      RECT  23.905 119.47 24.195 119.24 ;
      RECT  23.905 121.07 24.195 120.84 ;
      RECT  23.495 121.87 23.785 121.64 ;
      RECT  27.56 119.67 27.73 119.07 ;
      RECT  26.61 121.64 26.78 120.67 ;
      RECT  27.56 121.64 27.73 119.93 ;
      RECT  27.5 121.87 27.79 121.64 ;
      RECT  23.555 121.64 23.725 119.84 ;
      RECT  22.575 126.08 22.865 126.11 ;
      RECT  22.25 124.31 22.42 125.28 ;
      RECT  26.55 124.08 26.84 124.31 ;
      RECT  25.245 124.08 25.535 124.31 ;
      RECT  23.965 125.155 24.135 126.435 ;
      RECT  22.19 126.88 22.48 127.11 ;
      RECT  22.19 125.28 22.48 125.51 ;
      RECT  23.915 126.71 24.185 126.755 ;
      RECT  23.915 125.11 24.185 125.155 ;
      RECT  26.55 126.88 26.84 127.11 ;
      RECT  26.55 125.28 26.84 125.51 ;
      RECT  23.495 126.88 23.785 127.11 ;
      RECT  22.25 125.51 22.42 126.88 ;
      RECT  22.19 124.08 22.48 124.31 ;
      RECT  22.575 126.28 22.865 126.31 ;
      RECT  26.61 125.51 26.78 126.88 ;
      RECT  27.48 126.02 27.81 126.28 ;
      RECT  25.305 124.31 25.475 126.88 ;
      RECT  22.575 126.11 23.725 126.28 ;
      RECT  22.755 125.665 23.085 125.925 ;
      RECT  27.5 126.88 27.79 127.11 ;
      RECT  27.09 125.265 27.42 125.525 ;
      RECT  23.555 126.28 23.725 126.88 ;
      RECT  23.915 126.435 24.185 126.48 ;
      RECT  23.915 124.835 24.185 124.88 ;
      RECT  25.245 126.88 25.535 127.11 ;
      RECT  23.905 126.48 24.195 126.71 ;
      RECT  23.905 124.88 24.195 125.11 ;
      RECT  23.495 124.08 23.785 124.31 ;
      RECT  27.56 126.28 27.73 126.88 ;
      RECT  26.61 124.31 26.78 125.28 ;
      RECT  27.56 124.31 27.73 126.02 ;
      RECT  27.5 124.08 27.79 124.31 ;
      RECT  23.555 124.31 23.725 126.11 ;
      RECT  22.575 134.01 22.865 133.98 ;
      RECT  22.25 135.78 22.42 134.81 ;
      RECT  26.55 136.01 26.84 135.78 ;
      RECT  25.245 136.01 25.535 135.78 ;
      RECT  23.965 134.935 24.135 133.655 ;
      RECT  22.19 133.21 22.48 132.98 ;
      RECT  22.19 134.81 22.48 134.58 ;
      RECT  23.915 133.38 24.185 133.335 ;
      RECT  23.915 134.98 24.185 134.935 ;
      RECT  26.55 133.21 26.84 132.98 ;
      RECT  26.55 134.81 26.84 134.58 ;
      RECT  23.495 133.21 23.785 132.98 ;
      RECT  22.25 134.58 22.42 133.21 ;
      RECT  22.19 136.01 22.48 135.78 ;
      RECT  22.575 133.81 22.865 133.78 ;
      RECT  26.61 134.58 26.78 133.21 ;
      RECT  27.48 134.07 27.81 133.81 ;
      RECT  25.305 135.78 25.475 133.21 ;
      RECT  22.575 133.98 23.725 133.81 ;
      RECT  22.755 134.425 23.085 134.165 ;
      RECT  27.5 133.21 27.79 132.98 ;
      RECT  27.09 134.825 27.42 134.565 ;
      RECT  23.555 133.81 23.725 133.21 ;
      RECT  23.915 133.655 24.185 133.61 ;
      RECT  23.915 135.255 24.185 135.21 ;
      RECT  25.245 133.21 25.535 132.98 ;
      RECT  23.905 133.61 24.195 133.38 ;
      RECT  23.905 135.21 24.195 134.98 ;
      RECT  23.495 136.01 23.785 135.78 ;
      RECT  27.56 133.81 27.73 133.21 ;
      RECT  26.61 135.78 26.78 134.81 ;
      RECT  27.56 135.78 27.73 134.07 ;
      RECT  27.5 136.01 27.79 135.78 ;
      RECT  23.555 135.78 23.725 133.98 ;
      RECT  131.605 42.83 131.315 42.8 ;
      RECT  131.93 44.6 131.76 43.63 ;
      RECT  127.63 44.83 127.34 44.6 ;
      RECT  128.935 44.83 128.645 44.6 ;
      RECT  130.215 43.755 130.045 42.475 ;
      RECT  131.99 42.03 131.7 41.8 ;
      RECT  131.99 43.63 131.7 43.4 ;
      RECT  130.265 42.2 129.995 42.155 ;
      RECT  130.265 43.8 129.995 43.755 ;
      RECT  127.63 42.03 127.34 41.8 ;
      RECT  127.63 43.63 127.34 43.4 ;
      RECT  130.685 42.03 130.395 41.8 ;
      RECT  131.93 43.4 131.76 42.03 ;
      RECT  131.99 44.83 131.7 44.6 ;
      RECT  131.605 42.63 131.315 42.6 ;
      RECT  127.57 43.4 127.4 42.03 ;
      RECT  126.7 42.89 126.37 42.63 ;
      RECT  128.875 44.6 128.705 42.03 ;
      RECT  131.605 42.8 130.455 42.63 ;
      RECT  131.425 43.245 131.095 42.985 ;
      RECT  126.68 42.03 126.39 41.8 ;
      RECT  127.09 43.645 126.76 43.385 ;
      RECT  130.625 42.63 130.455 42.03 ;
      RECT  130.265 42.475 129.995 42.43 ;
      RECT  130.265 44.075 129.995 44.03 ;
      RECT  128.935 42.03 128.645 41.8 ;
      RECT  130.275 42.43 129.985 42.2 ;
      RECT  130.275 44.03 129.985 43.8 ;
      RECT  130.685 44.83 130.395 44.6 ;
      RECT  126.62 42.63 126.45 42.03 ;
      RECT  127.57 44.6 127.4 43.63 ;
      RECT  126.62 44.6 126.45 42.89 ;
      RECT  126.68 44.83 126.39 44.6 ;
      RECT  130.625 44.6 130.455 42.8 ;
      RECT  131.605 34.9 131.315 34.93 ;
      RECT  131.93 33.13 131.76 34.1 ;
      RECT  127.63 32.9 127.34 33.13 ;
      RECT  128.935 32.9 128.645 33.13 ;
      RECT  130.215 33.975 130.045 35.255 ;
      RECT  131.99 35.7 131.7 35.93 ;
      RECT  131.99 34.1 131.7 34.33 ;
      RECT  130.265 35.53 129.995 35.575 ;
      RECT  130.265 33.93 129.995 33.975 ;
      RECT  127.63 35.7 127.34 35.93 ;
      RECT  127.63 34.1 127.34 34.33 ;
      RECT  130.685 35.7 130.395 35.93 ;
      RECT  131.93 34.33 131.76 35.7 ;
      RECT  131.99 32.9 131.7 33.13 ;
      RECT  131.605 35.1 131.315 35.13 ;
      RECT  127.57 34.33 127.4 35.7 ;
      RECT  126.7 34.84 126.37 35.1 ;
      RECT  128.875 33.13 128.705 35.7 ;
      RECT  131.605 34.93 130.455 35.1 ;
      RECT  131.425 34.485 131.095 34.745 ;
      RECT  126.68 35.7 126.39 35.93 ;
      RECT  127.09 34.085 126.76 34.345 ;
      RECT  130.625 35.1 130.455 35.7 ;
      RECT  130.265 35.255 129.995 35.3 ;
      RECT  130.265 33.655 129.995 33.7 ;
      RECT  128.935 35.7 128.645 35.93 ;
      RECT  130.275 35.3 129.985 35.53 ;
      RECT  130.275 33.7 129.985 33.93 ;
      RECT  130.685 32.9 130.395 33.13 ;
      RECT  126.62 35.1 126.45 35.7 ;
      RECT  127.57 33.13 127.4 34.1 ;
      RECT  126.62 33.13 126.45 34.84 ;
      RECT  126.68 32.9 126.39 33.13 ;
      RECT  130.625 33.13 130.455 34.93 ;
      RECT  131.605 28.69 131.315 28.66 ;
      RECT  131.93 30.46 131.76 29.49 ;
      RECT  127.63 30.69 127.34 30.46 ;
      RECT  128.935 30.69 128.645 30.46 ;
      RECT  130.215 29.615 130.045 28.335 ;
      RECT  131.99 27.89 131.7 27.66 ;
      RECT  131.99 29.49 131.7 29.26 ;
      RECT  130.265 28.06 129.995 28.015 ;
      RECT  130.265 29.66 129.995 29.615 ;
      RECT  127.63 27.89 127.34 27.66 ;
      RECT  127.63 29.49 127.34 29.26 ;
      RECT  130.685 27.89 130.395 27.66 ;
      RECT  131.93 29.26 131.76 27.89 ;
      RECT  131.99 30.69 131.7 30.46 ;
      RECT  131.605 28.49 131.315 28.46 ;
      RECT  127.57 29.26 127.4 27.89 ;
      RECT  126.7 28.75 126.37 28.49 ;
      RECT  128.875 30.46 128.705 27.89 ;
      RECT  131.605 28.66 130.455 28.49 ;
      RECT  131.425 29.105 131.095 28.845 ;
      RECT  126.68 27.89 126.39 27.66 ;
      RECT  127.09 29.505 126.76 29.245 ;
      RECT  130.625 28.49 130.455 27.89 ;
      RECT  130.265 28.335 129.995 28.29 ;
      RECT  130.265 29.935 129.995 29.89 ;
      RECT  128.935 27.89 128.645 27.66 ;
      RECT  130.275 28.29 129.985 28.06 ;
      RECT  130.275 29.89 129.985 29.66 ;
      RECT  130.685 30.69 130.395 30.46 ;
      RECT  126.62 28.49 126.45 27.89 ;
      RECT  127.57 30.46 127.4 29.49 ;
      RECT  126.62 30.46 126.45 28.75 ;
      RECT  126.68 30.69 126.39 30.46 ;
      RECT  130.625 30.46 130.455 28.66 ;
      RECT  131.605 20.76 131.315 20.79 ;
      RECT  131.93 18.99 131.76 19.96 ;
      RECT  127.63 18.76 127.34 18.99 ;
      RECT  128.935 18.76 128.645 18.99 ;
      RECT  130.215 19.835 130.045 21.115 ;
      RECT  131.99 21.56 131.7 21.79 ;
      RECT  131.99 19.96 131.7 20.19 ;
      RECT  130.265 21.39 129.995 21.435 ;
      RECT  130.265 19.79 129.995 19.835 ;
      RECT  127.63 21.56 127.34 21.79 ;
      RECT  127.63 19.96 127.34 20.19 ;
      RECT  130.685 21.56 130.395 21.79 ;
      RECT  131.93 20.19 131.76 21.56 ;
      RECT  131.99 18.76 131.7 18.99 ;
      RECT  131.605 20.96 131.315 20.99 ;
      RECT  127.57 20.19 127.4 21.56 ;
      RECT  126.7 20.7 126.37 20.96 ;
      RECT  128.875 18.99 128.705 21.56 ;
      RECT  131.605 20.79 130.455 20.96 ;
      RECT  131.425 20.345 131.095 20.605 ;
      RECT  126.68 21.56 126.39 21.79 ;
      RECT  127.09 19.945 126.76 20.205 ;
      RECT  130.625 20.96 130.455 21.56 ;
      RECT  130.265 21.115 129.995 21.16 ;
      RECT  130.265 19.515 129.995 19.56 ;
      RECT  128.935 21.56 128.645 21.79 ;
      RECT  130.275 21.16 129.985 21.39 ;
      RECT  130.275 19.56 129.985 19.79 ;
      RECT  130.685 18.76 130.395 18.99 ;
      RECT  126.62 20.96 126.45 21.56 ;
      RECT  127.57 18.99 127.4 19.96 ;
      RECT  126.62 18.99 126.45 20.7 ;
      RECT  126.68 18.76 126.39 18.99 ;
      RECT  130.625 18.99 130.455 20.79 ;
      RECT  34.255 16.245 34.545 16.275 ;
      RECT  33.93 14.475 34.1 15.445 ;
      RECT  38.23 14.245 38.52 14.475 ;
      RECT  36.925 14.245 37.215 14.475 ;
      RECT  35.645 15.32 35.815 16.6 ;
      RECT  33.87 17.045 34.16 17.275 ;
      RECT  33.87 15.445 34.16 15.675 ;
      RECT  35.595 16.875 35.865 16.92 ;
      RECT  35.595 15.275 35.865 15.32 ;
      RECT  38.23 17.045 38.52 17.275 ;
      RECT  38.23 15.445 38.52 15.675 ;
      RECT  35.175 17.045 35.465 17.275 ;
      RECT  33.93 15.675 34.1 17.045 ;
      RECT  33.87 14.245 34.16 14.475 ;
      RECT  34.255 16.445 34.545 16.475 ;
      RECT  38.29 15.675 38.46 17.045 ;
      RECT  39.16 16.185 39.49 16.445 ;
      RECT  36.985 14.475 37.155 17.045 ;
      RECT  34.255 16.275 35.405 16.445 ;
      RECT  34.435 15.83 34.765 16.09 ;
      RECT  39.18 17.045 39.47 17.275 ;
      RECT  38.77 15.43 39.1 15.69 ;
      RECT  35.235 16.445 35.405 17.045 ;
      RECT  35.595 16.6 35.865 16.645 ;
      RECT  35.595 15.0 35.865 15.045 ;
      RECT  36.925 17.045 37.215 17.275 ;
      RECT  35.585 16.645 35.875 16.875 ;
      RECT  35.585 15.045 35.875 15.275 ;
      RECT  35.175 14.245 35.465 14.475 ;
      RECT  39.24 16.445 39.41 17.045 ;
      RECT  38.29 14.475 38.46 15.445 ;
      RECT  39.24 14.475 39.41 16.185 ;
      RECT  39.18 14.245 39.47 14.475 ;
      RECT  35.235 14.475 35.405 16.275 ;
      RECT  40.095 16.245 40.385 16.275 ;
      RECT  39.77 14.475 39.94 15.445 ;
      RECT  44.07 14.245 44.36 14.475 ;
      RECT  42.765 14.245 43.055 14.475 ;
      RECT  41.485 15.32 41.655 16.6 ;
      RECT  39.71 17.045 40.0 17.275 ;
      RECT  39.71 15.445 40.0 15.675 ;
      RECT  41.435 16.875 41.705 16.92 ;
      RECT  41.435 15.275 41.705 15.32 ;
      RECT  44.07 17.045 44.36 17.275 ;
      RECT  44.07 15.445 44.36 15.675 ;
      RECT  41.015 17.045 41.305 17.275 ;
      RECT  39.77 15.675 39.94 17.045 ;
      RECT  39.71 14.245 40.0 14.475 ;
      RECT  40.095 16.445 40.385 16.475 ;
      RECT  44.13 15.675 44.3 17.045 ;
      RECT  45.0 16.185 45.33 16.445 ;
      RECT  42.825 14.475 42.995 17.045 ;
      RECT  40.095 16.275 41.245 16.445 ;
      RECT  40.275 15.83 40.605 16.09 ;
      RECT  45.02 17.045 45.31 17.275 ;
      RECT  44.61 15.43 44.94 15.69 ;
      RECT  41.075 16.445 41.245 17.045 ;
      RECT  41.435 16.6 41.705 16.645 ;
      RECT  41.435 15.0 41.705 15.045 ;
      RECT  42.765 17.045 43.055 17.275 ;
      RECT  41.425 16.645 41.715 16.875 ;
      RECT  41.425 15.045 41.715 15.275 ;
      RECT  41.015 14.245 41.305 14.475 ;
      RECT  45.08 16.445 45.25 17.045 ;
      RECT  44.13 14.475 44.3 15.445 ;
      RECT  45.08 14.475 45.25 16.185 ;
      RECT  45.02 14.245 45.31 14.475 ;
      RECT  41.075 14.475 41.245 16.275 ;
   LAYER  m2 ;
      RECT  76.16 63.2 76.67 63.44 ;
      RECT  76.16 63.13 76.36 63.2 ;
      RECT  74.69 62.58 75.23 62.96 ;
      RECT  73.76 61.31 74.69 61.86 ;
      RECT  73.55 63.2 73.76 63.44 ;
      RECT  76.67 63.2 76.88 63.44 ;
      RECT  73.76 63.2 76.16 63.44 ;
      RECT  75.95 62.34 76.16 62.41 ;
      RECT  76.67 62.58 76.88 62.96 ;
      RECT  75.95 63.13 76.16 63.2 ;
      RECT  76.16 62.34 76.36 62.41 ;
      RECT  73.76 62.1 76.16 62.34 ;
      RECT  76.67 62.1 76.88 62.34 ;
      RECT  74.69 61.31 75.23 61.86 ;
      RECT  73.55 62.58 74.69 62.96 ;
      RECT  73.55 61.31 73.76 61.86 ;
      POLYGON  76.53 62.58 76.53 62.65 76.16 62.65 76.16 62.89 76.53 62.89 76.53 62.96 76.67 62.96 76.67 62.58 76.53 62.58 ;
      RECT  76.16 62.1 76.67 62.34 ;
      RECT  75.23 61.31 76.88 61.86 ;
      POLYGON  75.23 62.58 75.23 62.96 75.78 62.96 75.78 62.89 76.16 62.89 76.16 62.65 75.78 62.65 75.78 62.58 75.23 62.58 ;
      RECT  73.55 62.1 73.76 62.34 ;
      RECT  76.16 63.92 76.67 63.68 ;
      RECT  76.16 63.99 76.36 63.92 ;
      RECT  74.69 64.54 75.23 64.16 ;
      RECT  73.76 65.81 74.69 65.26 ;
      RECT  73.55 63.92 73.76 63.68 ;
      RECT  76.67 63.92 76.88 63.68 ;
      RECT  73.76 63.92 76.16 63.68 ;
      RECT  75.95 64.78 76.16 64.71 ;
      RECT  76.67 64.54 76.88 64.16 ;
      RECT  75.95 63.99 76.16 63.92 ;
      RECT  76.16 64.78 76.36 64.71 ;
      RECT  73.76 65.02 76.16 64.78 ;
      RECT  76.67 65.02 76.88 64.78 ;
      RECT  74.69 65.81 75.23 65.26 ;
      RECT  73.55 64.54 74.69 64.16 ;
      RECT  73.55 65.81 73.76 65.26 ;
      POLYGON  76.53 64.54 76.53 64.47 76.16 64.47 76.16 64.23 76.53 64.23 76.53 64.16 76.67 64.16 76.67 64.54 76.53 64.54 ;
      RECT  76.16 65.02 76.67 64.78 ;
      RECT  75.23 65.81 76.88 65.26 ;
      POLYGON  75.23 64.54 75.23 64.16 75.78 64.16 75.78 64.23 76.16 64.23 76.16 64.47 75.78 64.47 75.78 64.54 75.23 64.54 ;
      RECT  73.55 65.02 73.76 64.78 ;
      RECT  76.16 67.15 76.67 67.39 ;
      RECT  76.16 67.08 76.36 67.15 ;
      RECT  74.69 66.53 75.23 66.91 ;
      RECT  73.76 65.26 74.69 65.81 ;
      RECT  73.55 67.15 73.76 67.39 ;
      RECT  76.67 67.15 76.88 67.39 ;
      RECT  73.76 67.15 76.16 67.39 ;
      RECT  75.95 66.29 76.16 66.36 ;
      RECT  76.67 66.53 76.88 66.91 ;
      RECT  75.95 67.08 76.16 67.15 ;
      RECT  76.16 66.29 76.36 66.36 ;
      RECT  73.76 66.05 76.16 66.29 ;
      RECT  76.67 66.05 76.88 66.29 ;
      RECT  74.69 65.26 75.23 65.81 ;
      RECT  73.55 66.53 74.69 66.91 ;
      RECT  73.55 65.26 73.76 65.81 ;
      POLYGON  76.53 66.53 76.53 66.6 76.16 66.6 76.16 66.84 76.53 66.84 76.53 66.91 76.67 66.91 76.67 66.53 76.53 66.53 ;
      RECT  76.16 66.05 76.67 66.29 ;
      RECT  75.23 65.26 76.88 65.81 ;
      POLYGON  75.23 66.53 75.23 66.91 75.78 66.91 75.78 66.84 76.16 66.84 76.16 66.6 75.78 66.6 75.78 66.53 75.23 66.53 ;
      RECT  73.55 66.05 73.76 66.29 ;
      RECT  76.16 67.87 76.67 67.63 ;
      RECT  76.16 67.94 76.36 67.87 ;
      RECT  74.69 68.49 75.23 68.11 ;
      RECT  73.76 69.76 74.69 69.21 ;
      RECT  73.55 67.87 73.76 67.63 ;
      RECT  76.67 67.87 76.88 67.63 ;
      RECT  73.76 67.87 76.16 67.63 ;
      RECT  75.95 68.73 76.16 68.66 ;
      RECT  76.67 68.49 76.88 68.11 ;
      RECT  75.95 67.94 76.16 67.87 ;
      RECT  76.16 68.73 76.36 68.66 ;
      RECT  73.76 68.97 76.16 68.73 ;
      RECT  76.67 68.97 76.88 68.73 ;
      RECT  74.69 69.76 75.23 69.21 ;
      RECT  73.55 68.49 74.69 68.11 ;
      RECT  73.55 69.76 73.76 69.21 ;
      POLYGON  76.53 68.49 76.53 68.42 76.16 68.42 76.16 68.18 76.53 68.18 76.53 68.11 76.67 68.11 76.67 68.49 76.53 68.49 ;
      RECT  76.16 68.97 76.67 68.73 ;
      RECT  75.23 69.76 76.88 69.21 ;
      POLYGON  75.23 68.49 75.23 68.11 75.78 68.11 75.78 68.18 76.16 68.18 76.16 68.42 75.78 68.42 75.78 68.49 75.23 68.49 ;
      RECT  73.55 68.97 73.76 68.73 ;
      RECT  76.16 71.1 76.67 71.34 ;
      RECT  76.16 71.03 76.36 71.1 ;
      RECT  74.69 70.48 75.23 70.86 ;
      RECT  73.76 69.21 74.69 69.76 ;
      RECT  73.55 71.1 73.76 71.34 ;
      RECT  76.67 71.1 76.88 71.34 ;
      RECT  73.76 71.1 76.16 71.34 ;
      RECT  75.95 70.24 76.16 70.31 ;
      RECT  76.67 70.48 76.88 70.86 ;
      RECT  75.95 71.03 76.16 71.1 ;
      RECT  76.16 70.24 76.36 70.31 ;
      RECT  73.76 70.0 76.16 70.24 ;
      RECT  76.67 70.0 76.88 70.24 ;
      RECT  74.69 69.21 75.23 69.76 ;
      RECT  73.55 70.48 74.69 70.86 ;
      RECT  73.55 69.21 73.76 69.76 ;
      POLYGON  76.53 70.48 76.53 70.55 76.16 70.55 76.16 70.79 76.53 70.79 76.53 70.86 76.67 70.86 76.67 70.48 76.53 70.48 ;
      RECT  76.16 70.0 76.67 70.24 ;
      RECT  75.23 69.21 76.88 69.76 ;
      POLYGON  75.23 70.48 75.23 70.86 75.78 70.86 75.78 70.79 76.16 70.79 76.16 70.55 75.78 70.55 75.78 70.48 75.23 70.48 ;
      RECT  73.55 70.0 73.76 70.24 ;
      RECT  76.16 71.82 76.67 71.58 ;
      RECT  76.16 71.89 76.36 71.82 ;
      RECT  74.69 72.44 75.23 72.06 ;
      RECT  73.76 73.71 74.69 73.16 ;
      RECT  73.55 71.82 73.76 71.58 ;
      RECT  76.67 71.82 76.88 71.58 ;
      RECT  73.76 71.82 76.16 71.58 ;
      RECT  75.95 72.68 76.16 72.61 ;
      RECT  76.67 72.44 76.88 72.06 ;
      RECT  75.95 71.89 76.16 71.82 ;
      RECT  76.16 72.68 76.36 72.61 ;
      RECT  73.76 72.92 76.16 72.68 ;
      RECT  76.67 72.92 76.88 72.68 ;
      RECT  74.69 73.71 75.23 73.16 ;
      RECT  73.55 72.44 74.69 72.06 ;
      RECT  73.55 73.71 73.76 73.16 ;
      POLYGON  76.53 72.44 76.53 72.37 76.16 72.37 76.16 72.13 76.53 72.13 76.53 72.06 76.67 72.06 76.67 72.44 76.53 72.44 ;
      RECT  76.16 72.92 76.67 72.68 ;
      RECT  75.23 73.71 76.88 73.16 ;
      POLYGON  75.23 72.44 75.23 72.06 75.78 72.06 75.78 72.13 76.16 72.13 76.16 72.37 75.78 72.37 75.78 72.44 75.23 72.44 ;
      RECT  73.55 72.92 73.76 72.68 ;
      RECT  76.16 75.05 76.67 75.29 ;
      RECT  76.16 74.98 76.36 75.05 ;
      RECT  74.69 74.43 75.23 74.81 ;
      RECT  73.76 73.16 74.69 73.71 ;
      RECT  73.55 75.05 73.76 75.29 ;
      RECT  76.67 75.05 76.88 75.29 ;
      RECT  73.76 75.05 76.16 75.29 ;
      RECT  75.95 74.19 76.16 74.26 ;
      RECT  76.67 74.43 76.88 74.81 ;
      RECT  75.95 74.98 76.16 75.05 ;
      RECT  76.16 74.19 76.36 74.26 ;
      RECT  73.76 73.95 76.16 74.19 ;
      RECT  76.67 73.95 76.88 74.19 ;
      RECT  74.69 73.16 75.23 73.71 ;
      RECT  73.55 74.43 74.69 74.81 ;
      RECT  73.55 73.16 73.76 73.71 ;
      POLYGON  76.53 74.43 76.53 74.5 76.16 74.5 76.16 74.74 76.53 74.74 76.53 74.81 76.67 74.81 76.67 74.43 76.53 74.43 ;
      RECT  76.16 73.95 76.67 74.19 ;
      RECT  75.23 73.16 76.88 73.71 ;
      POLYGON  75.23 74.43 75.23 74.81 75.78 74.81 75.78 74.74 76.16 74.74 76.16 74.5 75.78 74.5 75.78 74.43 75.23 74.43 ;
      RECT  73.55 73.95 73.76 74.19 ;
      RECT  76.16 75.77 76.67 75.53 ;
      RECT  76.16 75.84 76.36 75.77 ;
      RECT  74.69 76.39 75.23 76.01 ;
      RECT  73.76 77.66 74.69 77.11 ;
      RECT  73.55 75.77 73.76 75.53 ;
      RECT  76.67 75.77 76.88 75.53 ;
      RECT  73.76 75.77 76.16 75.53 ;
      RECT  75.95 76.63 76.16 76.56 ;
      RECT  76.67 76.39 76.88 76.01 ;
      RECT  75.95 75.84 76.16 75.77 ;
      RECT  76.16 76.63 76.36 76.56 ;
      RECT  73.76 76.87 76.16 76.63 ;
      RECT  76.67 76.87 76.88 76.63 ;
      RECT  74.69 77.66 75.23 77.11 ;
      RECT  73.55 76.39 74.69 76.01 ;
      RECT  73.55 77.66 73.76 77.11 ;
      POLYGON  76.53 76.39 76.53 76.32 76.16 76.32 76.16 76.08 76.53 76.08 76.53 76.01 76.67 76.01 76.67 76.39 76.53 76.39 ;
      RECT  76.16 76.87 76.67 76.63 ;
      RECT  75.23 77.66 76.88 77.11 ;
      POLYGON  75.23 76.39 75.23 76.01 75.78 76.01 75.78 76.08 76.16 76.08 76.16 76.32 75.78 76.32 75.78 76.39 75.23 76.39 ;
      RECT  73.55 76.87 73.76 76.63 ;
      RECT  76.16 79.0 76.67 79.24 ;
      RECT  76.16 78.93 76.36 79.0 ;
      RECT  74.69 78.38 75.23 78.76 ;
      RECT  73.76 77.11 74.69 77.66 ;
      RECT  73.55 79.0 73.76 79.24 ;
      RECT  76.67 79.0 76.88 79.24 ;
      RECT  73.76 79.0 76.16 79.24 ;
      RECT  75.95 78.14 76.16 78.21 ;
      RECT  76.67 78.38 76.88 78.76 ;
      RECT  75.95 78.93 76.16 79.0 ;
      RECT  76.16 78.14 76.36 78.21 ;
      RECT  73.76 77.9 76.16 78.14 ;
      RECT  76.67 77.9 76.88 78.14 ;
      RECT  74.69 77.11 75.23 77.66 ;
      RECT  73.55 78.38 74.69 78.76 ;
      RECT  73.55 77.11 73.76 77.66 ;
      POLYGON  76.53 78.38 76.53 78.45 76.16 78.45 76.16 78.69 76.53 78.69 76.53 78.76 76.67 78.76 76.67 78.38 76.53 78.38 ;
      RECT  76.16 77.9 76.67 78.14 ;
      RECT  75.23 77.11 76.88 77.66 ;
      POLYGON  75.23 78.38 75.23 78.76 75.78 78.76 75.78 78.69 76.16 78.69 76.16 78.45 75.78 78.45 75.78 78.38 75.23 78.38 ;
      RECT  73.55 77.9 73.76 78.14 ;
      RECT  76.16 79.72 76.67 79.48 ;
      RECT  76.16 79.79 76.36 79.72 ;
      RECT  74.69 80.34 75.23 79.96 ;
      RECT  73.76 81.61 74.69 81.06 ;
      RECT  73.55 79.72 73.76 79.48 ;
      RECT  76.67 79.72 76.88 79.48 ;
      RECT  73.76 79.72 76.16 79.48 ;
      RECT  75.95 80.58 76.16 80.51 ;
      RECT  76.67 80.34 76.88 79.96 ;
      RECT  75.95 79.79 76.16 79.72 ;
      RECT  76.16 80.58 76.36 80.51 ;
      RECT  73.76 80.82 76.16 80.58 ;
      RECT  76.67 80.82 76.88 80.58 ;
      RECT  74.69 81.61 75.23 81.06 ;
      RECT  73.55 80.34 74.69 79.96 ;
      RECT  73.55 81.61 73.76 81.06 ;
      POLYGON  76.53 80.34 76.53 80.27 76.16 80.27 76.16 80.03 76.53 80.03 76.53 79.96 76.67 79.96 76.67 80.34 76.53 80.34 ;
      RECT  76.16 80.82 76.67 80.58 ;
      RECT  75.23 81.61 76.88 81.06 ;
      POLYGON  75.23 80.34 75.23 79.96 75.78 79.96 75.78 80.03 76.16 80.03 76.16 80.27 75.78 80.27 75.78 80.34 75.23 80.34 ;
      RECT  73.55 80.82 73.76 80.58 ;
      RECT  76.16 82.95 76.67 83.19 ;
      RECT  76.16 82.88 76.36 82.95 ;
      RECT  74.69 82.33 75.23 82.71 ;
      RECT  73.76 81.06 74.69 81.61 ;
      RECT  73.55 82.95 73.76 83.19 ;
      RECT  76.67 82.95 76.88 83.19 ;
      RECT  73.76 82.95 76.16 83.19 ;
      RECT  75.95 82.09 76.16 82.16 ;
      RECT  76.67 82.33 76.88 82.71 ;
      RECT  75.95 82.88 76.16 82.95 ;
      RECT  76.16 82.09 76.36 82.16 ;
      RECT  73.76 81.85 76.16 82.09 ;
      RECT  76.67 81.85 76.88 82.09 ;
      RECT  74.69 81.06 75.23 81.61 ;
      RECT  73.55 82.33 74.69 82.71 ;
      RECT  73.55 81.06 73.76 81.61 ;
      POLYGON  76.53 82.33 76.53 82.4 76.16 82.4 76.16 82.64 76.53 82.64 76.53 82.71 76.67 82.71 76.67 82.33 76.53 82.33 ;
      RECT  76.16 81.85 76.67 82.09 ;
      RECT  75.23 81.06 76.88 81.61 ;
      POLYGON  75.23 82.33 75.23 82.71 75.78 82.71 75.78 82.64 76.16 82.64 76.16 82.4 75.78 82.4 75.78 82.33 75.23 82.33 ;
      RECT  73.55 81.85 73.76 82.09 ;
      RECT  76.16 83.67 76.67 83.43 ;
      RECT  76.16 83.74 76.36 83.67 ;
      RECT  74.69 84.29 75.23 83.91 ;
      RECT  73.76 85.56 74.69 85.01 ;
      RECT  73.55 83.67 73.76 83.43 ;
      RECT  76.67 83.67 76.88 83.43 ;
      RECT  73.76 83.67 76.16 83.43 ;
      RECT  75.95 84.53 76.16 84.46 ;
      RECT  76.67 84.29 76.88 83.91 ;
      RECT  75.95 83.74 76.16 83.67 ;
      RECT  76.16 84.53 76.36 84.46 ;
      RECT  73.76 84.77 76.16 84.53 ;
      RECT  76.67 84.77 76.88 84.53 ;
      RECT  74.69 85.56 75.23 85.01 ;
      RECT  73.55 84.29 74.69 83.91 ;
      RECT  73.55 85.56 73.76 85.01 ;
      POLYGON  76.53 84.29 76.53 84.22 76.16 84.22 76.16 83.98 76.53 83.98 76.53 83.91 76.67 83.91 76.67 84.29 76.53 84.29 ;
      RECT  76.16 84.77 76.67 84.53 ;
      RECT  75.23 85.56 76.88 85.01 ;
      POLYGON  75.23 84.29 75.23 83.91 75.78 83.91 75.78 83.98 76.16 83.98 76.16 84.22 75.78 84.22 75.78 84.29 75.23 84.29 ;
      RECT  73.55 84.77 73.76 84.53 ;
      RECT  76.16 86.9 76.67 87.14 ;
      RECT  76.16 86.83 76.36 86.9 ;
      RECT  74.69 86.28 75.23 86.66 ;
      RECT  73.76 85.01 74.69 85.56 ;
      RECT  73.55 86.9 73.76 87.14 ;
      RECT  76.67 86.9 76.88 87.14 ;
      RECT  73.76 86.9 76.16 87.14 ;
      RECT  75.95 86.04 76.16 86.11 ;
      RECT  76.67 86.28 76.88 86.66 ;
      RECT  75.95 86.83 76.16 86.9 ;
      RECT  76.16 86.04 76.36 86.11 ;
      RECT  73.76 85.8 76.16 86.04 ;
      RECT  76.67 85.8 76.88 86.04 ;
      RECT  74.69 85.01 75.23 85.56 ;
      RECT  73.55 86.28 74.69 86.66 ;
      RECT  73.55 85.01 73.76 85.56 ;
      POLYGON  76.53 86.28 76.53 86.35 76.16 86.35 76.16 86.59 76.53 86.59 76.53 86.66 76.67 86.66 76.67 86.28 76.53 86.28 ;
      RECT  76.16 85.8 76.67 86.04 ;
      RECT  75.23 85.01 76.88 85.56 ;
      POLYGON  75.23 86.28 75.23 86.66 75.78 86.66 75.78 86.59 76.16 86.59 76.16 86.35 75.78 86.35 75.78 86.28 75.23 86.28 ;
      RECT  73.55 85.8 73.76 86.04 ;
      RECT  76.16 87.62 76.67 87.38 ;
      RECT  76.16 87.69 76.36 87.62 ;
      RECT  74.69 88.24 75.23 87.86 ;
      RECT  73.76 89.51 74.69 88.96 ;
      RECT  73.55 87.62 73.76 87.38 ;
      RECT  76.67 87.62 76.88 87.38 ;
      RECT  73.76 87.62 76.16 87.38 ;
      RECT  75.95 88.48 76.16 88.41 ;
      RECT  76.67 88.24 76.88 87.86 ;
      RECT  75.95 87.69 76.16 87.62 ;
      RECT  76.16 88.48 76.36 88.41 ;
      RECT  73.76 88.72 76.16 88.48 ;
      RECT  76.67 88.72 76.88 88.48 ;
      RECT  74.69 89.51 75.23 88.96 ;
      RECT  73.55 88.24 74.69 87.86 ;
      RECT  73.55 89.51 73.76 88.96 ;
      POLYGON  76.53 88.24 76.53 88.17 76.16 88.17 76.16 87.93 76.53 87.93 76.53 87.86 76.67 87.86 76.67 88.24 76.53 88.24 ;
      RECT  76.16 88.72 76.67 88.48 ;
      RECT  75.23 89.51 76.88 88.96 ;
      POLYGON  75.23 88.24 75.23 87.86 75.78 87.86 75.78 87.93 76.16 87.93 76.16 88.17 75.78 88.17 75.78 88.24 75.23 88.24 ;
      RECT  73.55 88.72 73.76 88.48 ;
      RECT  76.16 90.85 76.67 91.09 ;
      RECT  76.16 90.78 76.36 90.85 ;
      RECT  74.69 90.23 75.23 90.61 ;
      RECT  73.76 88.96 74.69 89.51 ;
      RECT  73.55 90.85 73.76 91.09 ;
      RECT  76.67 90.85 76.88 91.09 ;
      RECT  73.76 90.85 76.16 91.09 ;
      RECT  75.95 89.99 76.16 90.06 ;
      RECT  76.67 90.23 76.88 90.61 ;
      RECT  75.95 90.78 76.16 90.85 ;
      RECT  76.16 89.99 76.36 90.06 ;
      RECT  73.76 89.75 76.16 89.99 ;
      RECT  76.67 89.75 76.88 89.99 ;
      RECT  74.69 88.96 75.23 89.51 ;
      RECT  73.55 90.23 74.69 90.61 ;
      RECT  73.55 88.96 73.76 89.51 ;
      POLYGON  76.53 90.23 76.53 90.3 76.16 90.3 76.16 90.54 76.53 90.54 76.53 90.61 76.67 90.61 76.67 90.23 76.53 90.23 ;
      RECT  76.16 89.75 76.67 89.99 ;
      RECT  75.23 88.96 76.88 89.51 ;
      POLYGON  75.23 90.23 75.23 90.61 75.78 90.61 75.78 90.54 76.16 90.54 76.16 90.3 75.78 90.3 75.78 90.23 75.23 90.23 ;
      RECT  73.55 89.75 73.76 89.99 ;
      RECT  76.16 91.57 76.67 91.33 ;
      RECT  76.16 91.64 76.36 91.57 ;
      RECT  74.69 92.19 75.23 91.81 ;
      RECT  73.76 93.46 74.69 92.91 ;
      RECT  73.55 91.57 73.76 91.33 ;
      RECT  76.67 91.57 76.88 91.33 ;
      RECT  73.76 91.57 76.16 91.33 ;
      RECT  75.95 92.43 76.16 92.36 ;
      RECT  76.67 92.19 76.88 91.81 ;
      RECT  75.95 91.64 76.16 91.57 ;
      RECT  76.16 92.43 76.36 92.36 ;
      RECT  73.76 92.67 76.16 92.43 ;
      RECT  76.67 92.67 76.88 92.43 ;
      RECT  74.69 93.46 75.23 92.91 ;
      RECT  73.55 92.19 74.69 91.81 ;
      RECT  73.55 93.46 73.76 92.91 ;
      POLYGON  76.53 92.19 76.53 92.12 76.16 92.12 76.16 91.88 76.53 91.88 76.53 91.81 76.67 91.81 76.67 92.19 76.53 92.19 ;
      RECT  76.16 92.67 76.67 92.43 ;
      RECT  75.23 93.46 76.88 92.91 ;
      POLYGON  75.23 92.19 75.23 91.81 75.78 91.81 75.78 91.88 76.16 91.88 76.16 92.12 75.78 92.12 75.78 92.19 75.23 92.19 ;
      RECT  73.55 92.67 73.76 92.43 ;
      RECT  77.6 63.2 77.09 63.44 ;
      RECT  77.6 63.13 77.4 63.2 ;
      RECT  79.07 62.58 78.53 62.96 ;
      RECT  80.0 61.31 79.07 61.86 ;
      RECT  80.21 63.2 80.0 63.44 ;
      RECT  77.09 63.2 76.88 63.44 ;
      RECT  80.0 63.2 77.6 63.44 ;
      RECT  77.81 62.34 77.6 62.41 ;
      RECT  77.09 62.58 76.88 62.96 ;
      RECT  77.81 63.13 77.6 63.2 ;
      RECT  77.6 62.34 77.4 62.41 ;
      RECT  80.0 62.1 77.6 62.34 ;
      RECT  77.09 62.1 76.88 62.34 ;
      RECT  79.07 61.31 78.53 61.86 ;
      RECT  80.21 62.58 79.07 62.96 ;
      RECT  80.21 61.31 80.0 61.86 ;
      POLYGON  77.23 62.58 77.23 62.65 77.6 62.65 77.6 62.89 77.23 62.89 77.23 62.96 77.09 62.96 77.09 62.58 77.23 62.58 ;
      RECT  77.6 62.1 77.09 62.34 ;
      RECT  78.53 61.31 76.88 61.86 ;
      POLYGON  78.53 62.58 78.53 62.96 77.98 62.96 77.98 62.89 77.6 62.89 77.6 62.65 77.98 62.65 77.98 62.58 78.53 62.58 ;
      RECT  80.21 62.1 80.0 62.34 ;
      RECT  77.6 63.92 77.09 63.68 ;
      RECT  77.6 63.99 77.4 63.92 ;
      RECT  79.07 64.54 78.53 64.16 ;
      RECT  80.0 65.81 79.07 65.26 ;
      RECT  80.21 63.92 80.0 63.68 ;
      RECT  77.09 63.92 76.88 63.68 ;
      RECT  80.0 63.92 77.6 63.68 ;
      RECT  77.81 64.78 77.6 64.71 ;
      RECT  77.09 64.54 76.88 64.16 ;
      RECT  77.81 63.99 77.6 63.92 ;
      RECT  77.6 64.78 77.4 64.71 ;
      RECT  80.0 65.02 77.6 64.78 ;
      RECT  77.09 65.02 76.88 64.78 ;
      RECT  79.07 65.81 78.53 65.26 ;
      RECT  80.21 64.54 79.07 64.16 ;
      RECT  80.21 65.81 80.0 65.26 ;
      POLYGON  77.23 64.54 77.23 64.47 77.6 64.47 77.6 64.23 77.23 64.23 77.23 64.16 77.09 64.16 77.09 64.54 77.23 64.54 ;
      RECT  77.6 65.02 77.09 64.78 ;
      RECT  78.53 65.81 76.88 65.26 ;
      POLYGON  78.53 64.54 78.53 64.16 77.98 64.16 77.98 64.23 77.6 64.23 77.6 64.47 77.98 64.47 77.98 64.54 78.53 64.54 ;
      RECT  80.21 65.02 80.0 64.78 ;
      RECT  77.6 67.15 77.09 67.39 ;
      RECT  77.6 67.08 77.4 67.15 ;
      RECT  79.07 66.53 78.53 66.91 ;
      RECT  80.0 65.26 79.07 65.81 ;
      RECT  80.21 67.15 80.0 67.39 ;
      RECT  77.09 67.15 76.88 67.39 ;
      RECT  80.0 67.15 77.6 67.39 ;
      RECT  77.81 66.29 77.6 66.36 ;
      RECT  77.09 66.53 76.88 66.91 ;
      RECT  77.81 67.08 77.6 67.15 ;
      RECT  77.6 66.29 77.4 66.36 ;
      RECT  80.0 66.05 77.6 66.29 ;
      RECT  77.09 66.05 76.88 66.29 ;
      RECT  79.07 65.26 78.53 65.81 ;
      RECT  80.21 66.53 79.07 66.91 ;
      RECT  80.21 65.26 80.0 65.81 ;
      POLYGON  77.23 66.53 77.23 66.6 77.6 66.6 77.6 66.84 77.23 66.84 77.23 66.91 77.09 66.91 77.09 66.53 77.23 66.53 ;
      RECT  77.6 66.05 77.09 66.29 ;
      RECT  78.53 65.26 76.88 65.81 ;
      POLYGON  78.53 66.53 78.53 66.91 77.98 66.91 77.98 66.84 77.6 66.84 77.6 66.6 77.98 66.6 77.98 66.53 78.53 66.53 ;
      RECT  80.21 66.05 80.0 66.29 ;
      RECT  77.6 67.87 77.09 67.63 ;
      RECT  77.6 67.94 77.4 67.87 ;
      RECT  79.07 68.49 78.53 68.11 ;
      RECT  80.0 69.76 79.07 69.21 ;
      RECT  80.21 67.87 80.0 67.63 ;
      RECT  77.09 67.87 76.88 67.63 ;
      RECT  80.0 67.87 77.6 67.63 ;
      RECT  77.81 68.73 77.6 68.66 ;
      RECT  77.09 68.49 76.88 68.11 ;
      RECT  77.81 67.94 77.6 67.87 ;
      RECT  77.6 68.73 77.4 68.66 ;
      RECT  80.0 68.97 77.6 68.73 ;
      RECT  77.09 68.97 76.88 68.73 ;
      RECT  79.07 69.76 78.53 69.21 ;
      RECT  80.21 68.49 79.07 68.11 ;
      RECT  80.21 69.76 80.0 69.21 ;
      POLYGON  77.23 68.49 77.23 68.42 77.6 68.42 77.6 68.18 77.23 68.18 77.23 68.11 77.09 68.11 77.09 68.49 77.23 68.49 ;
      RECT  77.6 68.97 77.09 68.73 ;
      RECT  78.53 69.76 76.88 69.21 ;
      POLYGON  78.53 68.49 78.53 68.11 77.98 68.11 77.98 68.18 77.6 68.18 77.6 68.42 77.98 68.42 77.98 68.49 78.53 68.49 ;
      RECT  80.21 68.97 80.0 68.73 ;
      RECT  77.6 71.1 77.09 71.34 ;
      RECT  77.6 71.03 77.4 71.1 ;
      RECT  79.07 70.48 78.53 70.86 ;
      RECT  80.0 69.21 79.07 69.76 ;
      RECT  80.21 71.1 80.0 71.34 ;
      RECT  77.09 71.1 76.88 71.34 ;
      RECT  80.0 71.1 77.6 71.34 ;
      RECT  77.81 70.24 77.6 70.31 ;
      RECT  77.09 70.48 76.88 70.86 ;
      RECT  77.81 71.03 77.6 71.1 ;
      RECT  77.6 70.24 77.4 70.31 ;
      RECT  80.0 70.0 77.6 70.24 ;
      RECT  77.09 70.0 76.88 70.24 ;
      RECT  79.07 69.21 78.53 69.76 ;
      RECT  80.21 70.48 79.07 70.86 ;
      RECT  80.21 69.21 80.0 69.76 ;
      POLYGON  77.23 70.48 77.23 70.55 77.6 70.55 77.6 70.79 77.23 70.79 77.23 70.86 77.09 70.86 77.09 70.48 77.23 70.48 ;
      RECT  77.6 70.0 77.09 70.24 ;
      RECT  78.53 69.21 76.88 69.76 ;
      POLYGON  78.53 70.48 78.53 70.86 77.98 70.86 77.98 70.79 77.6 70.79 77.6 70.55 77.98 70.55 77.98 70.48 78.53 70.48 ;
      RECT  80.21 70.0 80.0 70.24 ;
      RECT  77.6 71.82 77.09 71.58 ;
      RECT  77.6 71.89 77.4 71.82 ;
      RECT  79.07 72.44 78.53 72.06 ;
      RECT  80.0 73.71 79.07 73.16 ;
      RECT  80.21 71.82 80.0 71.58 ;
      RECT  77.09 71.82 76.88 71.58 ;
      RECT  80.0 71.82 77.6 71.58 ;
      RECT  77.81 72.68 77.6 72.61 ;
      RECT  77.09 72.44 76.88 72.06 ;
      RECT  77.81 71.89 77.6 71.82 ;
      RECT  77.6 72.68 77.4 72.61 ;
      RECT  80.0 72.92 77.6 72.68 ;
      RECT  77.09 72.92 76.88 72.68 ;
      RECT  79.07 73.71 78.53 73.16 ;
      RECT  80.21 72.44 79.07 72.06 ;
      RECT  80.21 73.71 80.0 73.16 ;
      POLYGON  77.23 72.44 77.23 72.37 77.6 72.37 77.6 72.13 77.23 72.13 77.23 72.06 77.09 72.06 77.09 72.44 77.23 72.44 ;
      RECT  77.6 72.92 77.09 72.68 ;
      RECT  78.53 73.71 76.88 73.16 ;
      POLYGON  78.53 72.44 78.53 72.06 77.98 72.06 77.98 72.13 77.6 72.13 77.6 72.37 77.98 72.37 77.98 72.44 78.53 72.44 ;
      RECT  80.21 72.92 80.0 72.68 ;
      RECT  77.6 75.05 77.09 75.29 ;
      RECT  77.6 74.98 77.4 75.05 ;
      RECT  79.07 74.43 78.53 74.81 ;
      RECT  80.0 73.16 79.07 73.71 ;
      RECT  80.21 75.05 80.0 75.29 ;
      RECT  77.09 75.05 76.88 75.29 ;
      RECT  80.0 75.05 77.6 75.29 ;
      RECT  77.81 74.19 77.6 74.26 ;
      RECT  77.09 74.43 76.88 74.81 ;
      RECT  77.81 74.98 77.6 75.05 ;
      RECT  77.6 74.19 77.4 74.26 ;
      RECT  80.0 73.95 77.6 74.19 ;
      RECT  77.09 73.95 76.88 74.19 ;
      RECT  79.07 73.16 78.53 73.71 ;
      RECT  80.21 74.43 79.07 74.81 ;
      RECT  80.21 73.16 80.0 73.71 ;
      POLYGON  77.23 74.43 77.23 74.5 77.6 74.5 77.6 74.74 77.23 74.74 77.23 74.81 77.09 74.81 77.09 74.43 77.23 74.43 ;
      RECT  77.6 73.95 77.09 74.19 ;
      RECT  78.53 73.16 76.88 73.71 ;
      POLYGON  78.53 74.43 78.53 74.81 77.98 74.81 77.98 74.74 77.6 74.74 77.6 74.5 77.98 74.5 77.98 74.43 78.53 74.43 ;
      RECT  80.21 73.95 80.0 74.19 ;
      RECT  77.6 75.77 77.09 75.53 ;
      RECT  77.6 75.84 77.4 75.77 ;
      RECT  79.07 76.39 78.53 76.01 ;
      RECT  80.0 77.66 79.07 77.11 ;
      RECT  80.21 75.77 80.0 75.53 ;
      RECT  77.09 75.77 76.88 75.53 ;
      RECT  80.0 75.77 77.6 75.53 ;
      RECT  77.81 76.63 77.6 76.56 ;
      RECT  77.09 76.39 76.88 76.01 ;
      RECT  77.81 75.84 77.6 75.77 ;
      RECT  77.6 76.63 77.4 76.56 ;
      RECT  80.0 76.87 77.6 76.63 ;
      RECT  77.09 76.87 76.88 76.63 ;
      RECT  79.07 77.66 78.53 77.11 ;
      RECT  80.21 76.39 79.07 76.01 ;
      RECT  80.21 77.66 80.0 77.11 ;
      POLYGON  77.23 76.39 77.23 76.32 77.6 76.32 77.6 76.08 77.23 76.08 77.23 76.01 77.09 76.01 77.09 76.39 77.23 76.39 ;
      RECT  77.6 76.87 77.09 76.63 ;
      RECT  78.53 77.66 76.88 77.11 ;
      POLYGON  78.53 76.39 78.53 76.01 77.98 76.01 77.98 76.08 77.6 76.08 77.6 76.32 77.98 76.32 77.98 76.39 78.53 76.39 ;
      RECT  80.21 76.87 80.0 76.63 ;
      RECT  77.6 79.0 77.09 79.24 ;
      RECT  77.6 78.93 77.4 79.0 ;
      RECT  79.07 78.38 78.53 78.76 ;
      RECT  80.0 77.11 79.07 77.66 ;
      RECT  80.21 79.0 80.0 79.24 ;
      RECT  77.09 79.0 76.88 79.24 ;
      RECT  80.0 79.0 77.6 79.24 ;
      RECT  77.81 78.14 77.6 78.21 ;
      RECT  77.09 78.38 76.88 78.76 ;
      RECT  77.81 78.93 77.6 79.0 ;
      RECT  77.6 78.14 77.4 78.21 ;
      RECT  80.0 77.9 77.6 78.14 ;
      RECT  77.09 77.9 76.88 78.14 ;
      RECT  79.07 77.11 78.53 77.66 ;
      RECT  80.21 78.38 79.07 78.76 ;
      RECT  80.21 77.11 80.0 77.66 ;
      POLYGON  77.23 78.38 77.23 78.45 77.6 78.45 77.6 78.69 77.23 78.69 77.23 78.76 77.09 78.76 77.09 78.38 77.23 78.38 ;
      RECT  77.6 77.9 77.09 78.14 ;
      RECT  78.53 77.11 76.88 77.66 ;
      POLYGON  78.53 78.38 78.53 78.76 77.98 78.76 77.98 78.69 77.6 78.69 77.6 78.45 77.98 78.45 77.98 78.38 78.53 78.38 ;
      RECT  80.21 77.9 80.0 78.14 ;
      RECT  77.6 79.72 77.09 79.48 ;
      RECT  77.6 79.79 77.4 79.72 ;
      RECT  79.07 80.34 78.53 79.96 ;
      RECT  80.0 81.61 79.07 81.06 ;
      RECT  80.21 79.72 80.0 79.48 ;
      RECT  77.09 79.72 76.88 79.48 ;
      RECT  80.0 79.72 77.6 79.48 ;
      RECT  77.81 80.58 77.6 80.51 ;
      RECT  77.09 80.34 76.88 79.96 ;
      RECT  77.81 79.79 77.6 79.72 ;
      RECT  77.6 80.58 77.4 80.51 ;
      RECT  80.0 80.82 77.6 80.58 ;
      RECT  77.09 80.82 76.88 80.58 ;
      RECT  79.07 81.61 78.53 81.06 ;
      RECT  80.21 80.34 79.07 79.96 ;
      RECT  80.21 81.61 80.0 81.06 ;
      POLYGON  77.23 80.34 77.23 80.27 77.6 80.27 77.6 80.03 77.23 80.03 77.23 79.96 77.09 79.96 77.09 80.34 77.23 80.34 ;
      RECT  77.6 80.82 77.09 80.58 ;
      RECT  78.53 81.61 76.88 81.06 ;
      POLYGON  78.53 80.34 78.53 79.96 77.98 79.96 77.98 80.03 77.6 80.03 77.6 80.27 77.98 80.27 77.98 80.34 78.53 80.34 ;
      RECT  80.21 80.82 80.0 80.58 ;
      RECT  77.6 82.95 77.09 83.19 ;
      RECT  77.6 82.88 77.4 82.95 ;
      RECT  79.07 82.33 78.53 82.71 ;
      RECT  80.0 81.06 79.07 81.61 ;
      RECT  80.21 82.95 80.0 83.19 ;
      RECT  77.09 82.95 76.88 83.19 ;
      RECT  80.0 82.95 77.6 83.19 ;
      RECT  77.81 82.09 77.6 82.16 ;
      RECT  77.09 82.33 76.88 82.71 ;
      RECT  77.81 82.88 77.6 82.95 ;
      RECT  77.6 82.09 77.4 82.16 ;
      RECT  80.0 81.85 77.6 82.09 ;
      RECT  77.09 81.85 76.88 82.09 ;
      RECT  79.07 81.06 78.53 81.61 ;
      RECT  80.21 82.33 79.07 82.71 ;
      RECT  80.21 81.06 80.0 81.61 ;
      POLYGON  77.23 82.33 77.23 82.4 77.6 82.4 77.6 82.64 77.23 82.64 77.23 82.71 77.09 82.71 77.09 82.33 77.23 82.33 ;
      RECT  77.6 81.85 77.09 82.09 ;
      RECT  78.53 81.06 76.88 81.61 ;
      POLYGON  78.53 82.33 78.53 82.71 77.98 82.71 77.98 82.64 77.6 82.64 77.6 82.4 77.98 82.4 77.98 82.33 78.53 82.33 ;
      RECT  80.21 81.85 80.0 82.09 ;
      RECT  77.6 83.67 77.09 83.43 ;
      RECT  77.6 83.74 77.4 83.67 ;
      RECT  79.07 84.29 78.53 83.91 ;
      RECT  80.0 85.56 79.07 85.01 ;
      RECT  80.21 83.67 80.0 83.43 ;
      RECT  77.09 83.67 76.88 83.43 ;
      RECT  80.0 83.67 77.6 83.43 ;
      RECT  77.81 84.53 77.6 84.46 ;
      RECT  77.09 84.29 76.88 83.91 ;
      RECT  77.81 83.74 77.6 83.67 ;
      RECT  77.6 84.53 77.4 84.46 ;
      RECT  80.0 84.77 77.6 84.53 ;
      RECT  77.09 84.77 76.88 84.53 ;
      RECT  79.07 85.56 78.53 85.01 ;
      RECT  80.21 84.29 79.07 83.91 ;
      RECT  80.21 85.56 80.0 85.01 ;
      POLYGON  77.23 84.29 77.23 84.22 77.6 84.22 77.6 83.98 77.23 83.98 77.23 83.91 77.09 83.91 77.09 84.29 77.23 84.29 ;
      RECT  77.6 84.77 77.09 84.53 ;
      RECT  78.53 85.56 76.88 85.01 ;
      POLYGON  78.53 84.29 78.53 83.91 77.98 83.91 77.98 83.98 77.6 83.98 77.6 84.22 77.98 84.22 77.98 84.29 78.53 84.29 ;
      RECT  80.21 84.77 80.0 84.53 ;
      RECT  77.6 86.9 77.09 87.14 ;
      RECT  77.6 86.83 77.4 86.9 ;
      RECT  79.07 86.28 78.53 86.66 ;
      RECT  80.0 85.01 79.07 85.56 ;
      RECT  80.21 86.9 80.0 87.14 ;
      RECT  77.09 86.9 76.88 87.14 ;
      RECT  80.0 86.9 77.6 87.14 ;
      RECT  77.81 86.04 77.6 86.11 ;
      RECT  77.09 86.28 76.88 86.66 ;
      RECT  77.81 86.83 77.6 86.9 ;
      RECT  77.6 86.04 77.4 86.11 ;
      RECT  80.0 85.8 77.6 86.04 ;
      RECT  77.09 85.8 76.88 86.04 ;
      RECT  79.07 85.01 78.53 85.56 ;
      RECT  80.21 86.28 79.07 86.66 ;
      RECT  80.21 85.01 80.0 85.56 ;
      POLYGON  77.23 86.28 77.23 86.35 77.6 86.35 77.6 86.59 77.23 86.59 77.23 86.66 77.09 86.66 77.09 86.28 77.23 86.28 ;
      RECT  77.6 85.8 77.09 86.04 ;
      RECT  78.53 85.01 76.88 85.56 ;
      POLYGON  78.53 86.28 78.53 86.66 77.98 86.66 77.98 86.59 77.6 86.59 77.6 86.35 77.98 86.35 77.98 86.28 78.53 86.28 ;
      RECT  80.21 85.8 80.0 86.04 ;
      RECT  77.6 87.62 77.09 87.38 ;
      RECT  77.6 87.69 77.4 87.62 ;
      RECT  79.07 88.24 78.53 87.86 ;
      RECT  80.0 89.51 79.07 88.96 ;
      RECT  80.21 87.62 80.0 87.38 ;
      RECT  77.09 87.62 76.88 87.38 ;
      RECT  80.0 87.62 77.6 87.38 ;
      RECT  77.81 88.48 77.6 88.41 ;
      RECT  77.09 88.24 76.88 87.86 ;
      RECT  77.81 87.69 77.6 87.62 ;
      RECT  77.6 88.48 77.4 88.41 ;
      RECT  80.0 88.72 77.6 88.48 ;
      RECT  77.09 88.72 76.88 88.48 ;
      RECT  79.07 89.51 78.53 88.96 ;
      RECT  80.21 88.24 79.07 87.86 ;
      RECT  80.21 89.51 80.0 88.96 ;
      POLYGON  77.23 88.24 77.23 88.17 77.6 88.17 77.6 87.93 77.23 87.93 77.23 87.86 77.09 87.86 77.09 88.24 77.23 88.24 ;
      RECT  77.6 88.72 77.09 88.48 ;
      RECT  78.53 89.51 76.88 88.96 ;
      POLYGON  78.53 88.24 78.53 87.86 77.98 87.86 77.98 87.93 77.6 87.93 77.6 88.17 77.98 88.17 77.98 88.24 78.53 88.24 ;
      RECT  80.21 88.72 80.0 88.48 ;
      RECT  77.6 90.85 77.09 91.09 ;
      RECT  77.6 90.78 77.4 90.85 ;
      RECT  79.07 90.23 78.53 90.61 ;
      RECT  80.0 88.96 79.07 89.51 ;
      RECT  80.21 90.85 80.0 91.09 ;
      RECT  77.09 90.85 76.88 91.09 ;
      RECT  80.0 90.85 77.6 91.09 ;
      RECT  77.81 89.99 77.6 90.06 ;
      RECT  77.09 90.23 76.88 90.61 ;
      RECT  77.81 90.78 77.6 90.85 ;
      RECT  77.6 89.99 77.4 90.06 ;
      RECT  80.0 89.75 77.6 89.99 ;
      RECT  77.09 89.75 76.88 89.99 ;
      RECT  79.07 88.96 78.53 89.51 ;
      RECT  80.21 90.23 79.07 90.61 ;
      RECT  80.21 88.96 80.0 89.51 ;
      POLYGON  77.23 90.23 77.23 90.3 77.6 90.3 77.6 90.54 77.23 90.54 77.23 90.61 77.09 90.61 77.09 90.23 77.23 90.23 ;
      RECT  77.6 89.75 77.09 89.99 ;
      RECT  78.53 88.96 76.88 89.51 ;
      POLYGON  78.53 90.23 78.53 90.61 77.98 90.61 77.98 90.54 77.6 90.54 77.6 90.3 77.98 90.3 77.98 90.23 78.53 90.23 ;
      RECT  80.21 89.75 80.0 89.99 ;
      RECT  77.6 91.57 77.09 91.33 ;
      RECT  77.6 91.64 77.4 91.57 ;
      RECT  79.07 92.19 78.53 91.81 ;
      RECT  80.0 93.46 79.07 92.91 ;
      RECT  80.21 91.57 80.0 91.33 ;
      RECT  77.09 91.57 76.88 91.33 ;
      RECT  80.0 91.57 77.6 91.33 ;
      RECT  77.81 92.43 77.6 92.36 ;
      RECT  77.09 92.19 76.88 91.81 ;
      RECT  77.81 91.64 77.6 91.57 ;
      RECT  77.6 92.43 77.4 92.36 ;
      RECT  80.0 92.67 77.6 92.43 ;
      RECT  77.09 92.67 76.88 92.43 ;
      RECT  79.07 93.46 78.53 92.91 ;
      RECT  80.21 92.19 79.07 91.81 ;
      RECT  80.21 93.46 80.0 92.91 ;
      POLYGON  77.23 92.19 77.23 92.12 77.6 92.12 77.6 91.88 77.23 91.88 77.23 91.81 77.09 91.81 77.09 92.19 77.23 92.19 ;
      RECT  77.6 92.67 77.09 92.43 ;
      RECT  78.53 93.46 76.88 92.91 ;
      POLYGON  78.53 92.19 78.53 91.81 77.98 91.81 77.98 91.88 77.6 91.88 77.6 92.12 77.98 92.12 77.98 92.19 78.53 92.19 ;
      RECT  80.21 92.67 80.0 92.43 ;
      RECT  73.76 63.2 80.0 63.44 ;
      RECT  73.76 62.1 80.0 62.34 ;
      RECT  73.76 63.68 80.0 63.92 ;
      RECT  73.76 64.78 80.0 65.02 ;
      RECT  73.76 67.15 80.0 67.39 ;
      RECT  73.76 66.05 80.0 66.29 ;
      RECT  73.76 67.63 80.0 67.87 ;
      RECT  73.76 68.73 80.0 68.97 ;
      RECT  73.76 71.1 80.0 71.34 ;
      RECT  73.76 70.0 80.0 70.24 ;
      RECT  73.76 71.58 80.0 71.82 ;
      RECT  73.76 72.68 80.0 72.92 ;
      RECT  73.76 75.05 80.0 75.29 ;
      RECT  73.76 73.95 80.0 74.19 ;
      RECT  73.76 75.53 80.0 75.77 ;
      RECT  73.76 76.63 80.0 76.87 ;
      RECT  73.76 79.0 80.0 79.24 ;
      RECT  73.76 77.9 80.0 78.14 ;
      RECT  73.76 79.48 80.0 79.72 ;
      RECT  73.76 80.58 80.0 80.82 ;
      RECT  73.76 82.95 80.0 83.19 ;
      RECT  73.76 81.85 80.0 82.09 ;
      RECT  73.76 83.43 80.0 83.67 ;
      RECT  73.76 84.53 80.0 84.77 ;
      RECT  73.76 86.9 80.0 87.14 ;
      RECT  73.76 85.8 80.0 86.04 ;
      RECT  73.76 87.38 80.0 87.62 ;
      RECT  73.76 88.48 80.0 88.72 ;
      RECT  73.76 90.85 80.0 91.09 ;
      RECT  73.76 89.75 80.0 89.99 ;
      RECT  73.76 91.33 80.0 91.57 ;
      RECT  73.76 92.43 80.0 92.67 ;
      RECT  78.53 74.43 79.07 74.81 ;
      RECT  74.69 85.01 75.23 85.56 ;
      RECT  74.69 66.53 75.23 66.91 ;
      RECT  78.53 61.31 79.07 61.86 ;
      RECT  78.53 87.86 79.07 88.24 ;
      RECT  74.69 90.23 75.23 90.61 ;
      RECT  74.69 61.31 75.23 61.86 ;
      RECT  74.69 74.43 75.23 74.81 ;
      RECT  74.69 78.38 75.23 78.76 ;
      RECT  78.53 85.01 79.07 85.56 ;
      RECT  74.69 65.26 75.23 65.81 ;
      RECT  74.69 70.48 75.23 70.86 ;
      RECT  78.53 90.23 79.07 90.61 ;
      RECT  74.69 82.33 75.23 82.71 ;
      RECT  78.53 76.01 79.07 76.39 ;
      RECT  78.53 65.26 79.07 65.81 ;
      RECT  74.69 87.86 75.23 88.24 ;
      RECT  78.53 64.16 79.07 64.54 ;
      RECT  74.69 86.28 75.23 86.66 ;
      RECT  74.69 91.81 75.23 92.19 ;
      RECT  78.53 66.53 79.07 66.91 ;
      RECT  78.53 72.06 79.07 72.44 ;
      RECT  74.69 76.01 75.23 76.39 ;
      RECT  78.53 79.96 79.07 80.34 ;
      RECT  78.53 82.33 79.07 82.71 ;
      RECT  78.53 70.48 79.07 70.86 ;
      RECT  74.69 69.21 75.23 69.76 ;
      RECT  78.53 78.38 79.07 78.76 ;
      RECT  74.69 77.11 75.23 77.66 ;
      RECT  78.53 86.28 79.07 86.66 ;
      RECT  74.69 73.16 75.23 73.71 ;
      RECT  78.53 88.96 79.07 89.51 ;
      RECT  74.69 64.16 75.23 64.54 ;
      RECT  78.53 62.58 79.07 62.96 ;
      RECT  78.53 91.81 79.07 92.19 ;
      RECT  78.53 73.16 79.07 73.71 ;
      RECT  78.53 68.11 79.07 68.49 ;
      RECT  74.69 81.06 75.23 81.61 ;
      RECT  74.69 72.06 75.23 72.44 ;
      RECT  78.53 81.06 79.07 81.61 ;
      RECT  78.53 83.91 79.07 84.29 ;
      RECT  74.69 62.58 75.23 62.96 ;
      RECT  78.53 77.11 79.07 77.66 ;
      RECT  78.53 92.91 79.07 93.46 ;
      RECT  74.69 79.96 75.23 80.34 ;
      RECT  74.69 92.91 75.23 93.46 ;
      RECT  78.53 69.21 79.07 69.76 ;
      RECT  74.69 88.96 75.23 89.51 ;
      RECT  74.69 83.91 75.23 84.29 ;
      RECT  74.69 68.11 75.23 68.49 ;
      RECT  73.76 58.505 70.64 59.055 ;
      RECT  71.36 59.97 70.85 59.73 ;
      RECT  71.36 60.04 71.16 59.97 ;
      RECT  72.83 60.59 72.29 60.21 ;
      RECT  73.76 61.86 72.83 61.31 ;
      RECT  73.97 59.97 73.76 59.73 ;
      RECT  70.85 59.97 70.64 59.73 ;
      RECT  73.76 59.97 71.36 59.73 ;
      RECT  71.57 60.83 71.36 60.76 ;
      RECT  70.85 60.59 70.64 60.21 ;
      RECT  71.57 60.04 71.36 59.97 ;
      RECT  71.36 60.83 71.16 60.76 ;
      RECT  73.76 61.07 71.36 60.83 ;
      RECT  70.85 61.07 70.64 60.83 ;
      RECT  72.83 61.86 72.29 61.31 ;
      RECT  73.97 60.59 72.83 60.21 ;
      RECT  73.97 61.86 73.76 61.31 ;
      POLYGON  70.99 60.59 70.99 60.52 71.36 60.52 71.36 60.28 70.99 60.28 70.99 60.21 70.85 60.21 70.85 60.59 70.99 60.59 ;
      RECT  71.36 61.07 70.85 60.83 ;
      RECT  72.29 61.86 70.64 61.31 ;
      POLYGON  72.29 60.59 72.29 60.21 71.74 60.21 71.74 60.28 71.36 60.28 71.36 60.52 71.74 60.52 71.74 60.59 72.29 60.59 ;
      RECT  73.97 61.07 73.76 60.83 ;
      RECT  71.36 63.2 70.85 63.44 ;
      RECT  71.36 63.13 71.16 63.2 ;
      RECT  72.83 62.58 72.29 62.96 ;
      RECT  73.76 61.31 72.83 61.86 ;
      RECT  73.97 63.2 73.76 63.44 ;
      RECT  70.85 63.2 70.64 63.44 ;
      RECT  73.76 63.2 71.36 63.44 ;
      RECT  71.57 62.34 71.36 62.41 ;
      RECT  70.85 62.58 70.64 62.96 ;
      RECT  71.57 63.13 71.36 63.2 ;
      RECT  71.36 62.34 71.16 62.41 ;
      RECT  73.76 62.1 71.36 62.34 ;
      RECT  70.85 62.1 70.64 62.34 ;
      RECT  72.83 61.31 72.29 61.86 ;
      RECT  73.97 62.58 72.83 62.96 ;
      RECT  73.97 61.31 73.76 61.86 ;
      POLYGON  70.99 62.58 70.99 62.65 71.36 62.65 71.36 62.89 70.99 62.89 70.99 62.96 70.85 62.96 70.85 62.58 70.99 62.58 ;
      RECT  71.36 62.1 70.85 62.34 ;
      RECT  72.29 61.31 70.64 61.86 ;
      POLYGON  72.29 62.58 72.29 62.96 71.74 62.96 71.74 62.89 71.36 62.89 71.36 62.65 71.74 62.65 71.74 62.58 72.29 62.58 ;
      RECT  73.97 62.1 73.76 62.34 ;
      RECT  71.36 63.92 70.85 63.68 ;
      RECT  71.36 63.99 71.16 63.92 ;
      RECT  72.83 64.54 72.29 64.16 ;
      RECT  73.76 65.81 72.83 65.26 ;
      RECT  73.97 63.92 73.76 63.68 ;
      RECT  70.85 63.92 70.64 63.68 ;
      RECT  73.76 63.92 71.36 63.68 ;
      RECT  71.57 64.78 71.36 64.71 ;
      RECT  70.85 64.54 70.64 64.16 ;
      RECT  71.57 63.99 71.36 63.92 ;
      RECT  71.36 64.78 71.16 64.71 ;
      RECT  73.76 65.02 71.36 64.78 ;
      RECT  70.85 65.02 70.64 64.78 ;
      RECT  72.83 65.81 72.29 65.26 ;
      RECT  73.97 64.54 72.83 64.16 ;
      RECT  73.97 65.81 73.76 65.26 ;
      POLYGON  70.99 64.54 70.99 64.47 71.36 64.47 71.36 64.23 70.99 64.23 70.99 64.16 70.85 64.16 70.85 64.54 70.99 64.54 ;
      RECT  71.36 65.02 70.85 64.78 ;
      RECT  72.29 65.81 70.64 65.26 ;
      POLYGON  72.29 64.54 72.29 64.16 71.74 64.16 71.74 64.23 71.36 64.23 71.36 64.47 71.74 64.47 71.74 64.54 72.29 64.54 ;
      RECT  73.97 65.02 73.76 64.78 ;
      RECT  71.36 67.15 70.85 67.39 ;
      RECT  71.36 67.08 71.16 67.15 ;
      RECT  72.83 66.53 72.29 66.91 ;
      RECT  73.76 65.26 72.83 65.81 ;
      RECT  73.97 67.15 73.76 67.39 ;
      RECT  70.85 67.15 70.64 67.39 ;
      RECT  73.76 67.15 71.36 67.39 ;
      RECT  71.57 66.29 71.36 66.36 ;
      RECT  70.85 66.53 70.64 66.91 ;
      RECT  71.57 67.08 71.36 67.15 ;
      RECT  71.36 66.29 71.16 66.36 ;
      RECT  73.76 66.05 71.36 66.29 ;
      RECT  70.85 66.05 70.64 66.29 ;
      RECT  72.83 65.26 72.29 65.81 ;
      RECT  73.97 66.53 72.83 66.91 ;
      RECT  73.97 65.26 73.76 65.81 ;
      POLYGON  70.99 66.53 70.99 66.6 71.36 66.6 71.36 66.84 70.99 66.84 70.99 66.91 70.85 66.91 70.85 66.53 70.99 66.53 ;
      RECT  71.36 66.05 70.85 66.29 ;
      RECT  72.29 65.26 70.64 65.81 ;
      POLYGON  72.29 66.53 72.29 66.91 71.74 66.91 71.74 66.84 71.36 66.84 71.36 66.6 71.74 66.6 71.74 66.53 72.29 66.53 ;
      RECT  73.97 66.05 73.76 66.29 ;
      RECT  71.36 67.87 70.85 67.63 ;
      RECT  71.36 67.94 71.16 67.87 ;
      RECT  72.83 68.49 72.29 68.11 ;
      RECT  73.76 69.76 72.83 69.21 ;
      RECT  73.97 67.87 73.76 67.63 ;
      RECT  70.85 67.87 70.64 67.63 ;
      RECT  73.76 67.87 71.36 67.63 ;
      RECT  71.57 68.73 71.36 68.66 ;
      RECT  70.85 68.49 70.64 68.11 ;
      RECT  71.57 67.94 71.36 67.87 ;
      RECT  71.36 68.73 71.16 68.66 ;
      RECT  73.76 68.97 71.36 68.73 ;
      RECT  70.85 68.97 70.64 68.73 ;
      RECT  72.83 69.76 72.29 69.21 ;
      RECT  73.97 68.49 72.83 68.11 ;
      RECT  73.97 69.76 73.76 69.21 ;
      POLYGON  70.99 68.49 70.99 68.42 71.36 68.42 71.36 68.18 70.99 68.18 70.99 68.11 70.85 68.11 70.85 68.49 70.99 68.49 ;
      RECT  71.36 68.97 70.85 68.73 ;
      RECT  72.29 69.76 70.64 69.21 ;
      POLYGON  72.29 68.49 72.29 68.11 71.74 68.11 71.74 68.18 71.36 68.18 71.36 68.42 71.74 68.42 71.74 68.49 72.29 68.49 ;
      RECT  73.97 68.97 73.76 68.73 ;
      RECT  71.36 71.1 70.85 71.34 ;
      RECT  71.36 71.03 71.16 71.1 ;
      RECT  72.83 70.48 72.29 70.86 ;
      RECT  73.76 69.21 72.83 69.76 ;
      RECT  73.97 71.1 73.76 71.34 ;
      RECT  70.85 71.1 70.64 71.34 ;
      RECT  73.76 71.1 71.36 71.34 ;
      RECT  71.57 70.24 71.36 70.31 ;
      RECT  70.85 70.48 70.64 70.86 ;
      RECT  71.57 71.03 71.36 71.1 ;
      RECT  71.36 70.24 71.16 70.31 ;
      RECT  73.76 70.0 71.36 70.24 ;
      RECT  70.85 70.0 70.64 70.24 ;
      RECT  72.83 69.21 72.29 69.76 ;
      RECT  73.97 70.48 72.83 70.86 ;
      RECT  73.97 69.21 73.76 69.76 ;
      POLYGON  70.99 70.48 70.99 70.55 71.36 70.55 71.36 70.79 70.99 70.79 70.99 70.86 70.85 70.86 70.85 70.48 70.99 70.48 ;
      RECT  71.36 70.0 70.85 70.24 ;
      RECT  72.29 69.21 70.64 69.76 ;
      POLYGON  72.29 70.48 72.29 70.86 71.74 70.86 71.74 70.79 71.36 70.79 71.36 70.55 71.74 70.55 71.74 70.48 72.29 70.48 ;
      RECT  73.97 70.0 73.76 70.24 ;
      RECT  71.36 71.82 70.85 71.58 ;
      RECT  71.36 71.89 71.16 71.82 ;
      RECT  72.83 72.44 72.29 72.06 ;
      RECT  73.76 73.71 72.83 73.16 ;
      RECT  73.97 71.82 73.76 71.58 ;
      RECT  70.85 71.82 70.64 71.58 ;
      RECT  73.76 71.82 71.36 71.58 ;
      RECT  71.57 72.68 71.36 72.61 ;
      RECT  70.85 72.44 70.64 72.06 ;
      RECT  71.57 71.89 71.36 71.82 ;
      RECT  71.36 72.68 71.16 72.61 ;
      RECT  73.76 72.92 71.36 72.68 ;
      RECT  70.85 72.92 70.64 72.68 ;
      RECT  72.83 73.71 72.29 73.16 ;
      RECT  73.97 72.44 72.83 72.06 ;
      RECT  73.97 73.71 73.76 73.16 ;
      POLYGON  70.99 72.44 70.99 72.37 71.36 72.37 71.36 72.13 70.99 72.13 70.99 72.06 70.85 72.06 70.85 72.44 70.99 72.44 ;
      RECT  71.36 72.92 70.85 72.68 ;
      RECT  72.29 73.71 70.64 73.16 ;
      POLYGON  72.29 72.44 72.29 72.06 71.74 72.06 71.74 72.13 71.36 72.13 71.36 72.37 71.74 72.37 71.74 72.44 72.29 72.44 ;
      RECT  73.97 72.92 73.76 72.68 ;
      RECT  71.36 75.05 70.85 75.29 ;
      RECT  71.36 74.98 71.16 75.05 ;
      RECT  72.83 74.43 72.29 74.81 ;
      RECT  73.76 73.16 72.83 73.71 ;
      RECT  73.97 75.05 73.76 75.29 ;
      RECT  70.85 75.05 70.64 75.29 ;
      RECT  73.76 75.05 71.36 75.29 ;
      RECT  71.57 74.19 71.36 74.26 ;
      RECT  70.85 74.43 70.64 74.81 ;
      RECT  71.57 74.98 71.36 75.05 ;
      RECT  71.36 74.19 71.16 74.26 ;
      RECT  73.76 73.95 71.36 74.19 ;
      RECT  70.85 73.95 70.64 74.19 ;
      RECT  72.83 73.16 72.29 73.71 ;
      RECT  73.97 74.43 72.83 74.81 ;
      RECT  73.97 73.16 73.76 73.71 ;
      POLYGON  70.99 74.43 70.99 74.5 71.36 74.5 71.36 74.74 70.99 74.74 70.99 74.81 70.85 74.81 70.85 74.43 70.99 74.43 ;
      RECT  71.36 73.95 70.85 74.19 ;
      RECT  72.29 73.16 70.64 73.71 ;
      POLYGON  72.29 74.43 72.29 74.81 71.74 74.81 71.74 74.74 71.36 74.74 71.36 74.5 71.74 74.5 71.74 74.43 72.29 74.43 ;
      RECT  73.97 73.95 73.76 74.19 ;
      RECT  71.36 75.77 70.85 75.53 ;
      RECT  71.36 75.84 71.16 75.77 ;
      RECT  72.83 76.39 72.29 76.01 ;
      RECT  73.76 77.66 72.83 77.11 ;
      RECT  73.97 75.77 73.76 75.53 ;
      RECT  70.85 75.77 70.64 75.53 ;
      RECT  73.76 75.77 71.36 75.53 ;
      RECT  71.57 76.63 71.36 76.56 ;
      RECT  70.85 76.39 70.64 76.01 ;
      RECT  71.57 75.84 71.36 75.77 ;
      RECT  71.36 76.63 71.16 76.56 ;
      RECT  73.76 76.87 71.36 76.63 ;
      RECT  70.85 76.87 70.64 76.63 ;
      RECT  72.83 77.66 72.29 77.11 ;
      RECT  73.97 76.39 72.83 76.01 ;
      RECT  73.97 77.66 73.76 77.11 ;
      POLYGON  70.99 76.39 70.99 76.32 71.36 76.32 71.36 76.08 70.99 76.08 70.99 76.01 70.85 76.01 70.85 76.39 70.99 76.39 ;
      RECT  71.36 76.87 70.85 76.63 ;
      RECT  72.29 77.66 70.64 77.11 ;
      POLYGON  72.29 76.39 72.29 76.01 71.74 76.01 71.74 76.08 71.36 76.08 71.36 76.32 71.74 76.32 71.74 76.39 72.29 76.39 ;
      RECT  73.97 76.87 73.76 76.63 ;
      RECT  71.36 79.0 70.85 79.24 ;
      RECT  71.36 78.93 71.16 79.0 ;
      RECT  72.83 78.38 72.29 78.76 ;
      RECT  73.76 77.11 72.83 77.66 ;
      RECT  73.97 79.0 73.76 79.24 ;
      RECT  70.85 79.0 70.64 79.24 ;
      RECT  73.76 79.0 71.36 79.24 ;
      RECT  71.57 78.14 71.36 78.21 ;
      RECT  70.85 78.38 70.64 78.76 ;
      RECT  71.57 78.93 71.36 79.0 ;
      RECT  71.36 78.14 71.16 78.21 ;
      RECT  73.76 77.9 71.36 78.14 ;
      RECT  70.85 77.9 70.64 78.14 ;
      RECT  72.83 77.11 72.29 77.66 ;
      RECT  73.97 78.38 72.83 78.76 ;
      RECT  73.97 77.11 73.76 77.66 ;
      POLYGON  70.99 78.38 70.99 78.45 71.36 78.45 71.36 78.69 70.99 78.69 70.99 78.76 70.85 78.76 70.85 78.38 70.99 78.38 ;
      RECT  71.36 77.9 70.85 78.14 ;
      RECT  72.29 77.11 70.64 77.66 ;
      POLYGON  72.29 78.38 72.29 78.76 71.74 78.76 71.74 78.69 71.36 78.69 71.36 78.45 71.74 78.45 71.74 78.38 72.29 78.38 ;
      RECT  73.97 77.9 73.76 78.14 ;
      RECT  71.36 79.72 70.85 79.48 ;
      RECT  71.36 79.79 71.16 79.72 ;
      RECT  72.83 80.34 72.29 79.96 ;
      RECT  73.76 81.61 72.83 81.06 ;
      RECT  73.97 79.72 73.76 79.48 ;
      RECT  70.85 79.72 70.64 79.48 ;
      RECT  73.76 79.72 71.36 79.48 ;
      RECT  71.57 80.58 71.36 80.51 ;
      RECT  70.85 80.34 70.64 79.96 ;
      RECT  71.57 79.79 71.36 79.72 ;
      RECT  71.36 80.58 71.16 80.51 ;
      RECT  73.76 80.82 71.36 80.58 ;
      RECT  70.85 80.82 70.64 80.58 ;
      RECT  72.83 81.61 72.29 81.06 ;
      RECT  73.97 80.34 72.83 79.96 ;
      RECT  73.97 81.61 73.76 81.06 ;
      POLYGON  70.99 80.34 70.99 80.27 71.36 80.27 71.36 80.03 70.99 80.03 70.99 79.96 70.85 79.96 70.85 80.34 70.99 80.34 ;
      RECT  71.36 80.82 70.85 80.58 ;
      RECT  72.29 81.61 70.64 81.06 ;
      POLYGON  72.29 80.34 72.29 79.96 71.74 79.96 71.74 80.03 71.36 80.03 71.36 80.27 71.74 80.27 71.74 80.34 72.29 80.34 ;
      RECT  73.97 80.82 73.76 80.58 ;
      RECT  71.36 82.95 70.85 83.19 ;
      RECT  71.36 82.88 71.16 82.95 ;
      RECT  72.83 82.33 72.29 82.71 ;
      RECT  73.76 81.06 72.83 81.61 ;
      RECT  73.97 82.95 73.76 83.19 ;
      RECT  70.85 82.95 70.64 83.19 ;
      RECT  73.76 82.95 71.36 83.19 ;
      RECT  71.57 82.09 71.36 82.16 ;
      RECT  70.85 82.33 70.64 82.71 ;
      RECT  71.57 82.88 71.36 82.95 ;
      RECT  71.36 82.09 71.16 82.16 ;
      RECT  73.76 81.85 71.36 82.09 ;
      RECT  70.85 81.85 70.64 82.09 ;
      RECT  72.83 81.06 72.29 81.61 ;
      RECT  73.97 82.33 72.83 82.71 ;
      RECT  73.97 81.06 73.76 81.61 ;
      POLYGON  70.99 82.33 70.99 82.4 71.36 82.4 71.36 82.64 70.99 82.64 70.99 82.71 70.85 82.71 70.85 82.33 70.99 82.33 ;
      RECT  71.36 81.85 70.85 82.09 ;
      RECT  72.29 81.06 70.64 81.61 ;
      POLYGON  72.29 82.33 72.29 82.71 71.74 82.71 71.74 82.64 71.36 82.64 71.36 82.4 71.74 82.4 71.74 82.33 72.29 82.33 ;
      RECT  73.97 81.85 73.76 82.09 ;
      RECT  71.36 83.67 70.85 83.43 ;
      RECT  71.36 83.74 71.16 83.67 ;
      RECT  72.83 84.29 72.29 83.91 ;
      RECT  73.76 85.56 72.83 85.01 ;
      RECT  73.97 83.67 73.76 83.43 ;
      RECT  70.85 83.67 70.64 83.43 ;
      RECT  73.76 83.67 71.36 83.43 ;
      RECT  71.57 84.53 71.36 84.46 ;
      RECT  70.85 84.29 70.64 83.91 ;
      RECT  71.57 83.74 71.36 83.67 ;
      RECT  71.36 84.53 71.16 84.46 ;
      RECT  73.76 84.77 71.36 84.53 ;
      RECT  70.85 84.77 70.64 84.53 ;
      RECT  72.83 85.56 72.29 85.01 ;
      RECT  73.97 84.29 72.83 83.91 ;
      RECT  73.97 85.56 73.76 85.01 ;
      POLYGON  70.99 84.29 70.99 84.22 71.36 84.22 71.36 83.98 70.99 83.98 70.99 83.91 70.85 83.91 70.85 84.29 70.99 84.29 ;
      RECT  71.36 84.77 70.85 84.53 ;
      RECT  72.29 85.56 70.64 85.01 ;
      POLYGON  72.29 84.29 72.29 83.91 71.74 83.91 71.74 83.98 71.36 83.98 71.36 84.22 71.74 84.22 71.74 84.29 72.29 84.29 ;
      RECT  73.97 84.77 73.76 84.53 ;
      RECT  71.36 86.9 70.85 87.14 ;
      RECT  71.36 86.83 71.16 86.9 ;
      RECT  72.83 86.28 72.29 86.66 ;
      RECT  73.76 85.01 72.83 85.56 ;
      RECT  73.97 86.9 73.76 87.14 ;
      RECT  70.85 86.9 70.64 87.14 ;
      RECT  73.76 86.9 71.36 87.14 ;
      RECT  71.57 86.04 71.36 86.11 ;
      RECT  70.85 86.28 70.64 86.66 ;
      RECT  71.57 86.83 71.36 86.9 ;
      RECT  71.36 86.04 71.16 86.11 ;
      RECT  73.76 85.8 71.36 86.04 ;
      RECT  70.85 85.8 70.64 86.04 ;
      RECT  72.83 85.01 72.29 85.56 ;
      RECT  73.97 86.28 72.83 86.66 ;
      RECT  73.97 85.01 73.76 85.56 ;
      POLYGON  70.99 86.28 70.99 86.35 71.36 86.35 71.36 86.59 70.99 86.59 70.99 86.66 70.85 86.66 70.85 86.28 70.99 86.28 ;
      RECT  71.36 85.8 70.85 86.04 ;
      RECT  72.29 85.01 70.64 85.56 ;
      POLYGON  72.29 86.28 72.29 86.66 71.74 86.66 71.74 86.59 71.36 86.59 71.36 86.35 71.74 86.35 71.74 86.28 72.29 86.28 ;
      RECT  73.97 85.8 73.76 86.04 ;
      RECT  71.36 87.62 70.85 87.38 ;
      RECT  71.36 87.69 71.16 87.62 ;
      RECT  72.83 88.24 72.29 87.86 ;
      RECT  73.76 89.51 72.83 88.96 ;
      RECT  73.97 87.62 73.76 87.38 ;
      RECT  70.85 87.62 70.64 87.38 ;
      RECT  73.76 87.62 71.36 87.38 ;
      RECT  71.57 88.48 71.36 88.41 ;
      RECT  70.85 88.24 70.64 87.86 ;
      RECT  71.57 87.69 71.36 87.62 ;
      RECT  71.36 88.48 71.16 88.41 ;
      RECT  73.76 88.72 71.36 88.48 ;
      RECT  70.85 88.72 70.64 88.48 ;
      RECT  72.83 89.51 72.29 88.96 ;
      RECT  73.97 88.24 72.83 87.86 ;
      RECT  73.97 89.51 73.76 88.96 ;
      POLYGON  70.99 88.24 70.99 88.17 71.36 88.17 71.36 87.93 70.99 87.93 70.99 87.86 70.85 87.86 70.85 88.24 70.99 88.24 ;
      RECT  71.36 88.72 70.85 88.48 ;
      RECT  72.29 89.51 70.64 88.96 ;
      POLYGON  72.29 88.24 72.29 87.86 71.74 87.86 71.74 87.93 71.36 87.93 71.36 88.17 71.74 88.17 71.74 88.24 72.29 88.24 ;
      RECT  73.97 88.72 73.76 88.48 ;
      RECT  71.36 90.85 70.85 91.09 ;
      RECT  71.36 90.78 71.16 90.85 ;
      RECT  72.83 90.23 72.29 90.61 ;
      RECT  73.76 88.96 72.83 89.51 ;
      RECT  73.97 90.85 73.76 91.09 ;
      RECT  70.85 90.85 70.64 91.09 ;
      RECT  73.76 90.85 71.36 91.09 ;
      RECT  71.57 89.99 71.36 90.06 ;
      RECT  70.85 90.23 70.64 90.61 ;
      RECT  71.57 90.78 71.36 90.85 ;
      RECT  71.36 89.99 71.16 90.06 ;
      RECT  73.76 89.75 71.36 89.99 ;
      RECT  70.85 89.75 70.64 89.99 ;
      RECT  72.83 88.96 72.29 89.51 ;
      RECT  73.97 90.23 72.83 90.61 ;
      RECT  73.97 88.96 73.76 89.51 ;
      POLYGON  70.99 90.23 70.99 90.3 71.36 90.3 71.36 90.54 70.99 90.54 70.99 90.61 70.85 90.61 70.85 90.23 70.99 90.23 ;
      RECT  71.36 89.75 70.85 89.99 ;
      RECT  72.29 88.96 70.64 89.51 ;
      POLYGON  72.29 90.23 72.29 90.61 71.74 90.61 71.74 90.54 71.36 90.54 71.36 90.3 71.74 90.3 71.74 90.23 72.29 90.23 ;
      RECT  73.97 89.75 73.76 89.99 ;
      RECT  71.36 91.57 70.85 91.33 ;
      RECT  71.36 91.64 71.16 91.57 ;
      RECT  72.83 92.19 72.29 91.81 ;
      RECT  73.76 93.46 72.83 92.91 ;
      RECT  73.97 91.57 73.76 91.33 ;
      RECT  70.85 91.57 70.64 91.33 ;
      RECT  73.76 91.57 71.36 91.33 ;
      RECT  71.57 92.43 71.36 92.36 ;
      RECT  70.85 92.19 70.64 91.81 ;
      RECT  71.57 91.64 71.36 91.57 ;
      RECT  71.36 92.43 71.16 92.36 ;
      RECT  73.76 92.67 71.36 92.43 ;
      RECT  70.85 92.67 70.64 92.43 ;
      RECT  72.83 93.46 72.29 92.91 ;
      RECT  73.97 92.19 72.83 91.81 ;
      RECT  73.97 93.46 73.76 92.91 ;
      POLYGON  70.99 92.19 70.99 92.12 71.36 92.12 71.36 91.88 70.99 91.88 70.99 91.81 70.85 91.81 70.85 92.19 70.99 92.19 ;
      RECT  71.36 92.67 70.85 92.43 ;
      RECT  72.29 93.46 70.64 92.91 ;
      POLYGON  72.29 92.19 72.29 91.81 71.74 91.81 71.74 91.88 71.36 91.88 71.36 92.12 71.74 92.12 71.74 92.19 72.29 92.19 ;
      RECT  73.97 92.67 73.76 92.43 ;
      RECT  71.36 94.8 70.85 95.04 ;
      RECT  71.36 94.73 71.16 94.8 ;
      RECT  72.83 94.18 72.29 94.56 ;
      RECT  73.76 92.91 72.83 93.46 ;
      RECT  73.97 94.8 73.76 95.04 ;
      RECT  70.85 94.8 70.64 95.04 ;
      RECT  73.76 94.8 71.36 95.04 ;
      RECT  71.57 93.94 71.36 94.01 ;
      RECT  70.85 94.18 70.64 94.56 ;
      RECT  71.57 94.73 71.36 94.8 ;
      RECT  71.36 93.94 71.16 94.01 ;
      RECT  73.76 93.7 71.36 93.94 ;
      RECT  70.85 93.7 70.64 93.94 ;
      RECT  72.83 92.91 72.29 93.46 ;
      RECT  73.97 94.18 72.83 94.56 ;
      RECT  73.97 92.91 73.76 93.46 ;
      POLYGON  70.99 94.18 70.99 94.25 71.36 94.25 71.36 94.49 70.99 94.49 70.99 94.56 70.85 94.56 70.85 94.18 70.99 94.18 ;
      RECT  71.36 93.7 70.85 93.94 ;
      RECT  72.29 92.91 70.64 93.46 ;
      POLYGON  72.29 94.18 72.29 94.56 71.74 94.56 71.74 94.49 71.36 94.49 71.36 94.25 71.74 94.25 71.74 94.18 72.29 94.18 ;
      RECT  73.97 93.7 73.76 93.94 ;
      RECT  73.76 96.265 70.64 95.715 ;
      RECT  70.64 59.73 73.76 59.97 ;
      RECT  70.64 60.83 73.76 61.07 ;
      RECT  70.64 63.2 73.76 63.44 ;
      RECT  70.64 62.1 73.76 62.34 ;
      RECT  70.64 63.68 73.76 63.92 ;
      RECT  70.64 64.78 73.76 65.02 ;
      RECT  70.64 67.15 73.76 67.39 ;
      RECT  70.64 66.05 73.76 66.29 ;
      RECT  70.64 67.63 73.76 67.87 ;
      RECT  70.64 68.73 73.76 68.97 ;
      RECT  70.64 71.1 73.76 71.34 ;
      RECT  70.64 70.0 73.76 70.24 ;
      RECT  70.64 71.58 73.76 71.82 ;
      RECT  70.64 72.68 73.76 72.92 ;
      RECT  70.64 75.05 73.76 75.29 ;
      RECT  70.64 73.95 73.76 74.19 ;
      RECT  70.64 75.53 73.76 75.77 ;
      RECT  70.64 76.63 73.76 76.87 ;
      RECT  70.64 79.0 73.76 79.24 ;
      RECT  70.64 77.9 73.76 78.14 ;
      RECT  70.64 79.48 73.76 79.72 ;
      RECT  70.64 80.58 73.76 80.82 ;
      RECT  70.64 82.95 73.76 83.19 ;
      RECT  70.64 81.85 73.76 82.09 ;
      RECT  70.64 83.43 73.76 83.67 ;
      RECT  70.64 84.53 73.76 84.77 ;
      RECT  70.64 86.9 73.76 87.14 ;
      RECT  70.64 85.8 73.76 86.04 ;
      RECT  70.64 87.38 73.76 87.62 ;
      RECT  70.64 88.48 73.76 88.72 ;
      RECT  70.64 90.85 73.76 91.09 ;
      RECT  70.64 89.75 73.76 89.99 ;
      RECT  70.64 91.33 73.76 91.57 ;
      RECT  70.64 92.43 73.76 92.67 ;
      RECT  70.64 94.8 73.76 95.04 ;
      RECT  70.64 93.7 73.76 93.94 ;
      RECT  72.29 87.86 72.83 88.24 ;
      RECT  72.29 69.21 72.83 69.76 ;
      RECT  72.29 65.26 72.83 65.81 ;
      RECT  72.29 90.23 72.83 90.61 ;
      RECT  72.29 70.48 72.83 70.86 ;
      RECT  72.29 78.38 72.83 78.76 ;
      RECT  72.29 73.16 72.83 73.71 ;
      RECT  72.29 82.33 72.83 82.71 ;
      RECT  72.29 83.91 72.83 84.29 ;
      RECT  72.29 64.16 72.83 64.54 ;
      RECT  72.29 81.06 72.83 81.61 ;
      RECT  72.29 92.91 72.83 93.46 ;
      RECT  72.29 72.06 72.83 72.44 ;
      RECT  72.29 60.21 72.83 60.59 ;
      RECT  72.29 74.43 72.83 74.81 ;
      RECT  72.29 61.31 72.83 61.86 ;
      RECT  72.29 76.01 72.83 76.39 ;
      RECT  72.29 79.96 72.83 80.34 ;
      RECT  72.29 91.81 72.83 92.19 ;
      RECT  72.29 85.01 72.83 85.56 ;
      RECT  72.29 86.28 72.83 86.66 ;
      RECT  72.29 62.58 72.83 62.96 ;
      RECT  72.29 94.18 72.83 94.56 ;
      RECT  72.29 66.53 72.83 66.91 ;
      RECT  72.29 77.11 72.83 77.66 ;
      RECT  72.29 68.11 72.83 68.49 ;
      RECT  72.29 88.96 72.83 89.51 ;
      RECT  80.0 58.505 83.12 59.055 ;
      RECT  82.4 59.97 82.91 59.73 ;
      RECT  82.4 60.04 82.6 59.97 ;
      RECT  80.93 60.59 81.47 60.21 ;
      RECT  80.0 61.86 80.93 61.31 ;
      RECT  79.79 59.97 80.0 59.73 ;
      RECT  82.91 59.97 83.12 59.73 ;
      RECT  80.0 59.97 82.4 59.73 ;
      RECT  82.19 60.83 82.4 60.76 ;
      RECT  82.91 60.59 83.12 60.21 ;
      RECT  82.19 60.04 82.4 59.97 ;
      RECT  82.4 60.83 82.6 60.76 ;
      RECT  80.0 61.07 82.4 60.83 ;
      RECT  82.91 61.07 83.12 60.83 ;
      RECT  80.93 61.86 81.47 61.31 ;
      RECT  79.79 60.59 80.93 60.21 ;
      RECT  79.79 61.86 80.0 61.31 ;
      POLYGON  82.77 60.59 82.77 60.52 82.4 60.52 82.4 60.28 82.77 60.28 82.77 60.21 82.91 60.21 82.91 60.59 82.77 60.59 ;
      RECT  82.4 61.07 82.91 60.83 ;
      RECT  81.47 61.86 83.12 61.31 ;
      POLYGON  81.47 60.59 81.47 60.21 82.02 60.21 82.02 60.28 82.4 60.28 82.4 60.52 82.02 60.52 82.02 60.59 81.47 60.59 ;
      RECT  79.79 61.07 80.0 60.83 ;
      RECT  82.4 63.2 82.91 63.44 ;
      RECT  82.4 63.13 82.6 63.2 ;
      RECT  80.93 62.58 81.47 62.96 ;
      RECT  80.0 61.31 80.93 61.86 ;
      RECT  79.79 63.2 80.0 63.44 ;
      RECT  82.91 63.2 83.12 63.44 ;
      RECT  80.0 63.2 82.4 63.44 ;
      RECT  82.19 62.34 82.4 62.41 ;
      RECT  82.91 62.58 83.12 62.96 ;
      RECT  82.19 63.13 82.4 63.2 ;
      RECT  82.4 62.34 82.6 62.41 ;
      RECT  80.0 62.1 82.4 62.34 ;
      RECT  82.91 62.1 83.12 62.34 ;
      RECT  80.93 61.31 81.47 61.86 ;
      RECT  79.79 62.58 80.93 62.96 ;
      RECT  79.79 61.31 80.0 61.86 ;
      POLYGON  82.77 62.58 82.77 62.65 82.4 62.65 82.4 62.89 82.77 62.89 82.77 62.96 82.91 62.96 82.91 62.58 82.77 62.58 ;
      RECT  82.4 62.1 82.91 62.34 ;
      RECT  81.47 61.31 83.12 61.86 ;
      POLYGON  81.47 62.58 81.47 62.96 82.02 62.96 82.02 62.89 82.4 62.89 82.4 62.65 82.02 62.65 82.02 62.58 81.47 62.58 ;
      RECT  79.79 62.1 80.0 62.34 ;
      RECT  82.4 63.92 82.91 63.68 ;
      RECT  82.4 63.99 82.6 63.92 ;
      RECT  80.93 64.54 81.47 64.16 ;
      RECT  80.0 65.81 80.93 65.26 ;
      RECT  79.79 63.92 80.0 63.68 ;
      RECT  82.91 63.92 83.12 63.68 ;
      RECT  80.0 63.92 82.4 63.68 ;
      RECT  82.19 64.78 82.4 64.71 ;
      RECT  82.91 64.54 83.12 64.16 ;
      RECT  82.19 63.99 82.4 63.92 ;
      RECT  82.4 64.78 82.6 64.71 ;
      RECT  80.0 65.02 82.4 64.78 ;
      RECT  82.91 65.02 83.12 64.78 ;
      RECT  80.93 65.81 81.47 65.26 ;
      RECT  79.79 64.54 80.93 64.16 ;
      RECT  79.79 65.81 80.0 65.26 ;
      POLYGON  82.77 64.54 82.77 64.47 82.4 64.47 82.4 64.23 82.77 64.23 82.77 64.16 82.91 64.16 82.91 64.54 82.77 64.54 ;
      RECT  82.4 65.02 82.91 64.78 ;
      RECT  81.47 65.81 83.12 65.26 ;
      POLYGON  81.47 64.54 81.47 64.16 82.02 64.16 82.02 64.23 82.4 64.23 82.4 64.47 82.02 64.47 82.02 64.54 81.47 64.54 ;
      RECT  79.79 65.02 80.0 64.78 ;
      RECT  82.4 67.15 82.91 67.39 ;
      RECT  82.4 67.08 82.6 67.15 ;
      RECT  80.93 66.53 81.47 66.91 ;
      RECT  80.0 65.26 80.93 65.81 ;
      RECT  79.79 67.15 80.0 67.39 ;
      RECT  82.91 67.15 83.12 67.39 ;
      RECT  80.0 67.15 82.4 67.39 ;
      RECT  82.19 66.29 82.4 66.36 ;
      RECT  82.91 66.53 83.12 66.91 ;
      RECT  82.19 67.08 82.4 67.15 ;
      RECT  82.4 66.29 82.6 66.36 ;
      RECT  80.0 66.05 82.4 66.29 ;
      RECT  82.91 66.05 83.12 66.29 ;
      RECT  80.93 65.26 81.47 65.81 ;
      RECT  79.79 66.53 80.93 66.91 ;
      RECT  79.79 65.26 80.0 65.81 ;
      POLYGON  82.77 66.53 82.77 66.6 82.4 66.6 82.4 66.84 82.77 66.84 82.77 66.91 82.91 66.91 82.91 66.53 82.77 66.53 ;
      RECT  82.4 66.05 82.91 66.29 ;
      RECT  81.47 65.26 83.12 65.81 ;
      POLYGON  81.47 66.53 81.47 66.91 82.02 66.91 82.02 66.84 82.4 66.84 82.4 66.6 82.02 66.6 82.02 66.53 81.47 66.53 ;
      RECT  79.79 66.05 80.0 66.29 ;
      RECT  82.4 67.87 82.91 67.63 ;
      RECT  82.4 67.94 82.6 67.87 ;
      RECT  80.93 68.49 81.47 68.11 ;
      RECT  80.0 69.76 80.93 69.21 ;
      RECT  79.79 67.87 80.0 67.63 ;
      RECT  82.91 67.87 83.12 67.63 ;
      RECT  80.0 67.87 82.4 67.63 ;
      RECT  82.19 68.73 82.4 68.66 ;
      RECT  82.91 68.49 83.12 68.11 ;
      RECT  82.19 67.94 82.4 67.87 ;
      RECT  82.4 68.73 82.6 68.66 ;
      RECT  80.0 68.97 82.4 68.73 ;
      RECT  82.91 68.97 83.12 68.73 ;
      RECT  80.93 69.76 81.47 69.21 ;
      RECT  79.79 68.49 80.93 68.11 ;
      RECT  79.79 69.76 80.0 69.21 ;
      POLYGON  82.77 68.49 82.77 68.42 82.4 68.42 82.4 68.18 82.77 68.18 82.77 68.11 82.91 68.11 82.91 68.49 82.77 68.49 ;
      RECT  82.4 68.97 82.91 68.73 ;
      RECT  81.47 69.76 83.12 69.21 ;
      POLYGON  81.47 68.49 81.47 68.11 82.02 68.11 82.02 68.18 82.4 68.18 82.4 68.42 82.02 68.42 82.02 68.49 81.47 68.49 ;
      RECT  79.79 68.97 80.0 68.73 ;
      RECT  82.4 71.1 82.91 71.34 ;
      RECT  82.4 71.03 82.6 71.1 ;
      RECT  80.93 70.48 81.47 70.86 ;
      RECT  80.0 69.21 80.93 69.76 ;
      RECT  79.79 71.1 80.0 71.34 ;
      RECT  82.91 71.1 83.12 71.34 ;
      RECT  80.0 71.1 82.4 71.34 ;
      RECT  82.19 70.24 82.4 70.31 ;
      RECT  82.91 70.48 83.12 70.86 ;
      RECT  82.19 71.03 82.4 71.1 ;
      RECT  82.4 70.24 82.6 70.31 ;
      RECT  80.0 70.0 82.4 70.24 ;
      RECT  82.91 70.0 83.12 70.24 ;
      RECT  80.93 69.21 81.47 69.76 ;
      RECT  79.79 70.48 80.93 70.86 ;
      RECT  79.79 69.21 80.0 69.76 ;
      POLYGON  82.77 70.48 82.77 70.55 82.4 70.55 82.4 70.79 82.77 70.79 82.77 70.86 82.91 70.86 82.91 70.48 82.77 70.48 ;
      RECT  82.4 70.0 82.91 70.24 ;
      RECT  81.47 69.21 83.12 69.76 ;
      POLYGON  81.47 70.48 81.47 70.86 82.02 70.86 82.02 70.79 82.4 70.79 82.4 70.55 82.02 70.55 82.02 70.48 81.47 70.48 ;
      RECT  79.79 70.0 80.0 70.24 ;
      RECT  82.4 71.82 82.91 71.58 ;
      RECT  82.4 71.89 82.6 71.82 ;
      RECT  80.93 72.44 81.47 72.06 ;
      RECT  80.0 73.71 80.93 73.16 ;
      RECT  79.79 71.82 80.0 71.58 ;
      RECT  82.91 71.82 83.12 71.58 ;
      RECT  80.0 71.82 82.4 71.58 ;
      RECT  82.19 72.68 82.4 72.61 ;
      RECT  82.91 72.44 83.12 72.06 ;
      RECT  82.19 71.89 82.4 71.82 ;
      RECT  82.4 72.68 82.6 72.61 ;
      RECT  80.0 72.92 82.4 72.68 ;
      RECT  82.91 72.92 83.12 72.68 ;
      RECT  80.93 73.71 81.47 73.16 ;
      RECT  79.79 72.44 80.93 72.06 ;
      RECT  79.79 73.71 80.0 73.16 ;
      POLYGON  82.77 72.44 82.77 72.37 82.4 72.37 82.4 72.13 82.77 72.13 82.77 72.06 82.91 72.06 82.91 72.44 82.77 72.44 ;
      RECT  82.4 72.92 82.91 72.68 ;
      RECT  81.47 73.71 83.12 73.16 ;
      POLYGON  81.47 72.44 81.47 72.06 82.02 72.06 82.02 72.13 82.4 72.13 82.4 72.37 82.02 72.37 82.02 72.44 81.47 72.44 ;
      RECT  79.79 72.92 80.0 72.68 ;
      RECT  82.4 75.05 82.91 75.29 ;
      RECT  82.4 74.98 82.6 75.05 ;
      RECT  80.93 74.43 81.47 74.81 ;
      RECT  80.0 73.16 80.93 73.71 ;
      RECT  79.79 75.05 80.0 75.29 ;
      RECT  82.91 75.05 83.12 75.29 ;
      RECT  80.0 75.05 82.4 75.29 ;
      RECT  82.19 74.19 82.4 74.26 ;
      RECT  82.91 74.43 83.12 74.81 ;
      RECT  82.19 74.98 82.4 75.05 ;
      RECT  82.4 74.19 82.6 74.26 ;
      RECT  80.0 73.95 82.4 74.19 ;
      RECT  82.91 73.95 83.12 74.19 ;
      RECT  80.93 73.16 81.47 73.71 ;
      RECT  79.79 74.43 80.93 74.81 ;
      RECT  79.79 73.16 80.0 73.71 ;
      POLYGON  82.77 74.43 82.77 74.5 82.4 74.5 82.4 74.74 82.77 74.74 82.77 74.81 82.91 74.81 82.91 74.43 82.77 74.43 ;
      RECT  82.4 73.95 82.91 74.19 ;
      RECT  81.47 73.16 83.12 73.71 ;
      POLYGON  81.47 74.43 81.47 74.81 82.02 74.81 82.02 74.74 82.4 74.74 82.4 74.5 82.02 74.5 82.02 74.43 81.47 74.43 ;
      RECT  79.79 73.95 80.0 74.19 ;
      RECT  82.4 75.77 82.91 75.53 ;
      RECT  82.4 75.84 82.6 75.77 ;
      RECT  80.93 76.39 81.47 76.01 ;
      RECT  80.0 77.66 80.93 77.11 ;
      RECT  79.79 75.77 80.0 75.53 ;
      RECT  82.91 75.77 83.12 75.53 ;
      RECT  80.0 75.77 82.4 75.53 ;
      RECT  82.19 76.63 82.4 76.56 ;
      RECT  82.91 76.39 83.12 76.01 ;
      RECT  82.19 75.84 82.4 75.77 ;
      RECT  82.4 76.63 82.6 76.56 ;
      RECT  80.0 76.87 82.4 76.63 ;
      RECT  82.91 76.87 83.12 76.63 ;
      RECT  80.93 77.66 81.47 77.11 ;
      RECT  79.79 76.39 80.93 76.01 ;
      RECT  79.79 77.66 80.0 77.11 ;
      POLYGON  82.77 76.39 82.77 76.32 82.4 76.32 82.4 76.08 82.77 76.08 82.77 76.01 82.91 76.01 82.91 76.39 82.77 76.39 ;
      RECT  82.4 76.87 82.91 76.63 ;
      RECT  81.47 77.66 83.12 77.11 ;
      POLYGON  81.47 76.39 81.47 76.01 82.02 76.01 82.02 76.08 82.4 76.08 82.4 76.32 82.02 76.32 82.02 76.39 81.47 76.39 ;
      RECT  79.79 76.87 80.0 76.63 ;
      RECT  82.4 79.0 82.91 79.24 ;
      RECT  82.4 78.93 82.6 79.0 ;
      RECT  80.93 78.38 81.47 78.76 ;
      RECT  80.0 77.11 80.93 77.66 ;
      RECT  79.79 79.0 80.0 79.24 ;
      RECT  82.91 79.0 83.12 79.24 ;
      RECT  80.0 79.0 82.4 79.24 ;
      RECT  82.19 78.14 82.4 78.21 ;
      RECT  82.91 78.38 83.12 78.76 ;
      RECT  82.19 78.93 82.4 79.0 ;
      RECT  82.4 78.14 82.6 78.21 ;
      RECT  80.0 77.9 82.4 78.14 ;
      RECT  82.91 77.9 83.12 78.14 ;
      RECT  80.93 77.11 81.47 77.66 ;
      RECT  79.79 78.38 80.93 78.76 ;
      RECT  79.79 77.11 80.0 77.66 ;
      POLYGON  82.77 78.38 82.77 78.45 82.4 78.45 82.4 78.69 82.77 78.69 82.77 78.76 82.91 78.76 82.91 78.38 82.77 78.38 ;
      RECT  82.4 77.9 82.91 78.14 ;
      RECT  81.47 77.11 83.12 77.66 ;
      POLYGON  81.47 78.38 81.47 78.76 82.02 78.76 82.02 78.69 82.4 78.69 82.4 78.45 82.02 78.45 82.02 78.38 81.47 78.38 ;
      RECT  79.79 77.9 80.0 78.14 ;
      RECT  82.4 79.72 82.91 79.48 ;
      RECT  82.4 79.79 82.6 79.72 ;
      RECT  80.93 80.34 81.47 79.96 ;
      RECT  80.0 81.61 80.93 81.06 ;
      RECT  79.79 79.72 80.0 79.48 ;
      RECT  82.91 79.72 83.12 79.48 ;
      RECT  80.0 79.72 82.4 79.48 ;
      RECT  82.19 80.58 82.4 80.51 ;
      RECT  82.91 80.34 83.12 79.96 ;
      RECT  82.19 79.79 82.4 79.72 ;
      RECT  82.4 80.58 82.6 80.51 ;
      RECT  80.0 80.82 82.4 80.58 ;
      RECT  82.91 80.82 83.12 80.58 ;
      RECT  80.93 81.61 81.47 81.06 ;
      RECT  79.79 80.34 80.93 79.96 ;
      RECT  79.79 81.61 80.0 81.06 ;
      POLYGON  82.77 80.34 82.77 80.27 82.4 80.27 82.4 80.03 82.77 80.03 82.77 79.96 82.91 79.96 82.91 80.34 82.77 80.34 ;
      RECT  82.4 80.82 82.91 80.58 ;
      RECT  81.47 81.61 83.12 81.06 ;
      POLYGON  81.47 80.34 81.47 79.96 82.02 79.96 82.02 80.03 82.4 80.03 82.4 80.27 82.02 80.27 82.02 80.34 81.47 80.34 ;
      RECT  79.79 80.82 80.0 80.58 ;
      RECT  82.4 82.95 82.91 83.19 ;
      RECT  82.4 82.88 82.6 82.95 ;
      RECT  80.93 82.33 81.47 82.71 ;
      RECT  80.0 81.06 80.93 81.61 ;
      RECT  79.79 82.95 80.0 83.19 ;
      RECT  82.91 82.95 83.12 83.19 ;
      RECT  80.0 82.95 82.4 83.19 ;
      RECT  82.19 82.09 82.4 82.16 ;
      RECT  82.91 82.33 83.12 82.71 ;
      RECT  82.19 82.88 82.4 82.95 ;
      RECT  82.4 82.09 82.6 82.16 ;
      RECT  80.0 81.85 82.4 82.09 ;
      RECT  82.91 81.85 83.12 82.09 ;
      RECT  80.93 81.06 81.47 81.61 ;
      RECT  79.79 82.33 80.93 82.71 ;
      RECT  79.79 81.06 80.0 81.61 ;
      POLYGON  82.77 82.33 82.77 82.4 82.4 82.4 82.4 82.64 82.77 82.64 82.77 82.71 82.91 82.71 82.91 82.33 82.77 82.33 ;
      RECT  82.4 81.85 82.91 82.09 ;
      RECT  81.47 81.06 83.12 81.61 ;
      POLYGON  81.47 82.33 81.47 82.71 82.02 82.71 82.02 82.64 82.4 82.64 82.4 82.4 82.02 82.4 82.02 82.33 81.47 82.33 ;
      RECT  79.79 81.85 80.0 82.09 ;
      RECT  82.4 83.67 82.91 83.43 ;
      RECT  82.4 83.74 82.6 83.67 ;
      RECT  80.93 84.29 81.47 83.91 ;
      RECT  80.0 85.56 80.93 85.01 ;
      RECT  79.79 83.67 80.0 83.43 ;
      RECT  82.91 83.67 83.12 83.43 ;
      RECT  80.0 83.67 82.4 83.43 ;
      RECT  82.19 84.53 82.4 84.46 ;
      RECT  82.91 84.29 83.12 83.91 ;
      RECT  82.19 83.74 82.4 83.67 ;
      RECT  82.4 84.53 82.6 84.46 ;
      RECT  80.0 84.77 82.4 84.53 ;
      RECT  82.91 84.77 83.12 84.53 ;
      RECT  80.93 85.56 81.47 85.01 ;
      RECT  79.79 84.29 80.93 83.91 ;
      RECT  79.79 85.56 80.0 85.01 ;
      POLYGON  82.77 84.29 82.77 84.22 82.4 84.22 82.4 83.98 82.77 83.98 82.77 83.91 82.91 83.91 82.91 84.29 82.77 84.29 ;
      RECT  82.4 84.77 82.91 84.53 ;
      RECT  81.47 85.56 83.12 85.01 ;
      POLYGON  81.47 84.29 81.47 83.91 82.02 83.91 82.02 83.98 82.4 83.98 82.4 84.22 82.02 84.22 82.02 84.29 81.47 84.29 ;
      RECT  79.79 84.77 80.0 84.53 ;
      RECT  82.4 86.9 82.91 87.14 ;
      RECT  82.4 86.83 82.6 86.9 ;
      RECT  80.93 86.28 81.47 86.66 ;
      RECT  80.0 85.01 80.93 85.56 ;
      RECT  79.79 86.9 80.0 87.14 ;
      RECT  82.91 86.9 83.12 87.14 ;
      RECT  80.0 86.9 82.4 87.14 ;
      RECT  82.19 86.04 82.4 86.11 ;
      RECT  82.91 86.28 83.12 86.66 ;
      RECT  82.19 86.83 82.4 86.9 ;
      RECT  82.4 86.04 82.6 86.11 ;
      RECT  80.0 85.8 82.4 86.04 ;
      RECT  82.91 85.8 83.12 86.04 ;
      RECT  80.93 85.01 81.47 85.56 ;
      RECT  79.79 86.28 80.93 86.66 ;
      RECT  79.79 85.01 80.0 85.56 ;
      POLYGON  82.77 86.28 82.77 86.35 82.4 86.35 82.4 86.59 82.77 86.59 82.77 86.66 82.91 86.66 82.91 86.28 82.77 86.28 ;
      RECT  82.4 85.8 82.91 86.04 ;
      RECT  81.47 85.01 83.12 85.56 ;
      POLYGON  81.47 86.28 81.47 86.66 82.02 86.66 82.02 86.59 82.4 86.59 82.4 86.35 82.02 86.35 82.02 86.28 81.47 86.28 ;
      RECT  79.79 85.8 80.0 86.04 ;
      RECT  82.4 87.62 82.91 87.38 ;
      RECT  82.4 87.69 82.6 87.62 ;
      RECT  80.93 88.24 81.47 87.86 ;
      RECT  80.0 89.51 80.93 88.96 ;
      RECT  79.79 87.62 80.0 87.38 ;
      RECT  82.91 87.62 83.12 87.38 ;
      RECT  80.0 87.62 82.4 87.38 ;
      RECT  82.19 88.48 82.4 88.41 ;
      RECT  82.91 88.24 83.12 87.86 ;
      RECT  82.19 87.69 82.4 87.62 ;
      RECT  82.4 88.48 82.6 88.41 ;
      RECT  80.0 88.72 82.4 88.48 ;
      RECT  82.91 88.72 83.12 88.48 ;
      RECT  80.93 89.51 81.47 88.96 ;
      RECT  79.79 88.24 80.93 87.86 ;
      RECT  79.79 89.51 80.0 88.96 ;
      POLYGON  82.77 88.24 82.77 88.17 82.4 88.17 82.4 87.93 82.77 87.93 82.77 87.86 82.91 87.86 82.91 88.24 82.77 88.24 ;
      RECT  82.4 88.72 82.91 88.48 ;
      RECT  81.47 89.51 83.12 88.96 ;
      POLYGON  81.47 88.24 81.47 87.86 82.02 87.86 82.02 87.93 82.4 87.93 82.4 88.17 82.02 88.17 82.02 88.24 81.47 88.24 ;
      RECT  79.79 88.72 80.0 88.48 ;
      RECT  82.4 90.85 82.91 91.09 ;
      RECT  82.4 90.78 82.6 90.85 ;
      RECT  80.93 90.23 81.47 90.61 ;
      RECT  80.0 88.96 80.93 89.51 ;
      RECT  79.79 90.85 80.0 91.09 ;
      RECT  82.91 90.85 83.12 91.09 ;
      RECT  80.0 90.85 82.4 91.09 ;
      RECT  82.19 89.99 82.4 90.06 ;
      RECT  82.91 90.23 83.12 90.61 ;
      RECT  82.19 90.78 82.4 90.85 ;
      RECT  82.4 89.99 82.6 90.06 ;
      RECT  80.0 89.75 82.4 89.99 ;
      RECT  82.91 89.75 83.12 89.99 ;
      RECT  80.93 88.96 81.47 89.51 ;
      RECT  79.79 90.23 80.93 90.61 ;
      RECT  79.79 88.96 80.0 89.51 ;
      POLYGON  82.77 90.23 82.77 90.3 82.4 90.3 82.4 90.54 82.77 90.54 82.77 90.61 82.91 90.61 82.91 90.23 82.77 90.23 ;
      RECT  82.4 89.75 82.91 89.99 ;
      RECT  81.47 88.96 83.12 89.51 ;
      POLYGON  81.47 90.23 81.47 90.61 82.02 90.61 82.02 90.54 82.4 90.54 82.4 90.3 82.02 90.3 82.02 90.23 81.47 90.23 ;
      RECT  79.79 89.75 80.0 89.99 ;
      RECT  82.4 91.57 82.91 91.33 ;
      RECT  82.4 91.64 82.6 91.57 ;
      RECT  80.93 92.19 81.47 91.81 ;
      RECT  80.0 93.46 80.93 92.91 ;
      RECT  79.79 91.57 80.0 91.33 ;
      RECT  82.91 91.57 83.12 91.33 ;
      RECT  80.0 91.57 82.4 91.33 ;
      RECT  82.19 92.43 82.4 92.36 ;
      RECT  82.91 92.19 83.12 91.81 ;
      RECT  82.19 91.64 82.4 91.57 ;
      RECT  82.4 92.43 82.6 92.36 ;
      RECT  80.0 92.67 82.4 92.43 ;
      RECT  82.91 92.67 83.12 92.43 ;
      RECT  80.93 93.46 81.47 92.91 ;
      RECT  79.79 92.19 80.93 91.81 ;
      RECT  79.79 93.46 80.0 92.91 ;
      POLYGON  82.77 92.19 82.77 92.12 82.4 92.12 82.4 91.88 82.77 91.88 82.77 91.81 82.91 91.81 82.91 92.19 82.77 92.19 ;
      RECT  82.4 92.67 82.91 92.43 ;
      RECT  81.47 93.46 83.12 92.91 ;
      POLYGON  81.47 92.19 81.47 91.81 82.02 91.81 82.02 91.88 82.4 91.88 82.4 92.12 82.02 92.12 82.02 92.19 81.47 92.19 ;
      RECT  79.79 92.67 80.0 92.43 ;
      RECT  82.4 94.8 82.91 95.04 ;
      RECT  82.4 94.73 82.6 94.8 ;
      RECT  80.93 94.18 81.47 94.56 ;
      RECT  80.0 92.91 80.93 93.46 ;
      RECT  79.79 94.8 80.0 95.04 ;
      RECT  82.91 94.8 83.12 95.04 ;
      RECT  80.0 94.8 82.4 95.04 ;
      RECT  82.19 93.94 82.4 94.01 ;
      RECT  82.91 94.18 83.12 94.56 ;
      RECT  82.19 94.73 82.4 94.8 ;
      RECT  82.4 93.94 82.6 94.01 ;
      RECT  80.0 93.7 82.4 93.94 ;
      RECT  82.91 93.7 83.12 93.94 ;
      RECT  80.93 92.91 81.47 93.46 ;
      RECT  79.79 94.18 80.93 94.56 ;
      RECT  79.79 92.91 80.0 93.46 ;
      POLYGON  82.77 94.18 82.77 94.25 82.4 94.25 82.4 94.49 82.77 94.49 82.77 94.56 82.91 94.56 82.91 94.18 82.77 94.18 ;
      RECT  82.4 93.7 82.91 93.94 ;
      RECT  81.47 92.91 83.12 93.46 ;
      POLYGON  81.47 94.18 81.47 94.56 82.02 94.56 82.02 94.49 82.4 94.49 82.4 94.25 82.02 94.25 82.02 94.18 81.47 94.18 ;
      RECT  79.79 93.7 80.0 93.94 ;
      RECT  80.0 96.265 83.12 95.715 ;
      RECT  80.0 59.73 83.12 59.97 ;
      RECT  80.0 60.83 83.12 61.07 ;
      RECT  80.0 63.2 83.12 63.44 ;
      RECT  80.0 62.1 83.12 62.34 ;
      RECT  80.0 63.68 83.12 63.92 ;
      RECT  80.0 64.78 83.12 65.02 ;
      RECT  80.0 67.15 83.12 67.39 ;
      RECT  80.0 66.05 83.12 66.29 ;
      RECT  80.0 67.63 83.12 67.87 ;
      RECT  80.0 68.73 83.12 68.97 ;
      RECT  80.0 71.1 83.12 71.34 ;
      RECT  80.0 70.0 83.12 70.24 ;
      RECT  80.0 71.58 83.12 71.82 ;
      RECT  80.0 72.68 83.12 72.92 ;
      RECT  80.0 75.05 83.12 75.29 ;
      RECT  80.0 73.95 83.12 74.19 ;
      RECT  80.0 75.53 83.12 75.77 ;
      RECT  80.0 76.63 83.12 76.87 ;
      RECT  80.0 79.0 83.12 79.24 ;
      RECT  80.0 77.9 83.12 78.14 ;
      RECT  80.0 79.48 83.12 79.72 ;
      RECT  80.0 80.58 83.12 80.82 ;
      RECT  80.0 82.95 83.12 83.19 ;
      RECT  80.0 81.85 83.12 82.09 ;
      RECT  80.0 83.43 83.12 83.67 ;
      RECT  80.0 84.53 83.12 84.77 ;
      RECT  80.0 86.9 83.12 87.14 ;
      RECT  80.0 85.8 83.12 86.04 ;
      RECT  80.0 87.38 83.12 87.62 ;
      RECT  80.0 88.48 83.12 88.72 ;
      RECT  80.0 90.85 83.12 91.09 ;
      RECT  80.0 89.75 83.12 89.99 ;
      RECT  80.0 91.33 83.12 91.57 ;
      RECT  80.0 92.43 83.12 92.67 ;
      RECT  80.0 94.8 83.12 95.04 ;
      RECT  80.0 93.7 83.12 93.94 ;
      RECT  80.93 81.06 81.47 81.61 ;
      RECT  80.93 62.58 81.47 62.96 ;
      RECT  80.93 86.28 81.47 86.66 ;
      RECT  80.93 70.48 81.47 70.86 ;
      RECT  80.93 74.43 81.47 74.81 ;
      RECT  80.93 61.31 81.47 61.86 ;
      RECT  80.93 90.23 81.47 90.61 ;
      RECT  80.93 66.53 81.47 66.91 ;
      RECT  80.93 92.91 81.47 93.46 ;
      RECT  80.93 78.38 81.47 78.76 ;
      RECT  80.93 83.91 81.47 84.29 ;
      RECT  80.93 91.81 81.47 92.19 ;
      RECT  80.93 82.33 81.47 82.71 ;
      RECT  80.93 87.86 81.47 88.24 ;
      RECT  80.93 72.06 81.47 72.44 ;
      RECT  80.93 94.18 81.47 94.56 ;
      RECT  80.93 65.26 81.47 65.81 ;
      RECT  80.93 73.16 81.47 73.71 ;
      RECT  80.93 69.21 81.47 69.76 ;
      RECT  80.93 60.21 81.47 60.59 ;
      RECT  80.93 77.11 81.47 77.66 ;
      RECT  80.93 68.11 81.47 68.49 ;
      RECT  80.93 76.01 81.47 76.39 ;
      RECT  80.93 88.96 81.47 89.51 ;
      RECT  80.93 85.01 81.47 85.56 ;
      RECT  80.93 79.96 81.47 80.34 ;
      RECT  80.93 64.16 81.47 64.54 ;
      RECT  76.16 59.97 76.67 59.73 ;
      RECT  76.16 60.04 76.36 59.97 ;
      RECT  74.69 60.59 75.23 60.21 ;
      RECT  73.76 61.86 74.69 61.31 ;
      RECT  73.55 59.97 73.76 59.73 ;
      RECT  76.67 59.97 76.88 59.73 ;
      RECT  73.76 59.97 76.16 59.73 ;
      RECT  75.95 60.83 76.16 60.76 ;
      RECT  76.67 60.59 76.88 60.21 ;
      RECT  75.95 60.04 76.16 59.97 ;
      RECT  76.16 60.83 76.36 60.76 ;
      RECT  73.76 61.07 76.16 60.83 ;
      RECT  76.67 61.07 76.88 60.83 ;
      RECT  74.69 61.86 75.23 61.31 ;
      RECT  73.55 60.59 74.69 60.21 ;
      RECT  73.55 61.86 73.76 61.31 ;
      POLYGON  76.53 60.59 76.53 60.52 76.16 60.52 76.16 60.28 76.53 60.28 76.53 60.21 76.67 60.21 76.67 60.59 76.53 60.59 ;
      RECT  76.16 61.07 76.67 60.83 ;
      RECT  75.23 61.86 76.88 61.31 ;
      POLYGON  75.23 60.59 75.23 60.21 75.78 60.21 75.78 60.28 76.16 60.28 76.16 60.52 75.78 60.52 75.78 60.59 75.23 60.59 ;
      RECT  73.55 61.07 73.76 60.83 ;
      RECT  77.6 59.97 77.09 59.73 ;
      RECT  77.6 60.04 77.4 59.97 ;
      RECT  79.07 60.59 78.53 60.21 ;
      RECT  80.0 61.86 79.07 61.31 ;
      RECT  80.21 59.97 80.0 59.73 ;
      RECT  77.09 59.97 76.88 59.73 ;
      RECT  80.0 59.97 77.6 59.73 ;
      RECT  77.81 60.83 77.6 60.76 ;
      RECT  77.09 60.59 76.88 60.21 ;
      RECT  77.81 60.04 77.6 59.97 ;
      RECT  77.6 60.83 77.4 60.76 ;
      RECT  80.0 61.07 77.6 60.83 ;
      RECT  77.09 61.07 76.88 60.83 ;
      RECT  79.07 61.86 78.53 61.31 ;
      RECT  80.21 60.59 79.07 60.21 ;
      RECT  80.21 61.86 80.0 61.31 ;
      POLYGON  77.23 60.59 77.23 60.52 77.6 60.52 77.6 60.28 77.23 60.28 77.23 60.21 77.09 60.21 77.09 60.59 77.23 60.59 ;
      RECT  77.6 61.07 77.09 60.83 ;
      RECT  78.53 61.86 76.88 61.31 ;
      POLYGON  78.53 60.59 78.53 60.21 77.98 60.21 77.98 60.28 77.6 60.28 77.6 60.52 77.98 60.52 77.98 60.59 78.53 60.59 ;
      RECT  80.21 61.07 80.0 60.83 ;
      RECT  73.76 59.97 80.0 59.73 ;
      RECT  73.76 61.07 80.0 60.83 ;
      RECT  74.69 61.86 75.23 61.31 ;
      RECT  74.69 60.59 75.23 60.21 ;
      RECT  78.53 60.59 79.07 60.21 ;
      RECT  78.53 61.86 79.07 61.31 ;
      RECT  76.16 94.8 76.67 95.04 ;
      RECT  76.16 94.73 76.36 94.8 ;
      RECT  74.69 94.18 75.23 94.56 ;
      RECT  73.76 92.91 74.69 93.46 ;
      RECT  73.55 94.8 73.76 95.04 ;
      RECT  76.67 94.8 76.88 95.04 ;
      RECT  73.76 94.8 76.16 95.04 ;
      RECT  75.95 93.94 76.16 94.01 ;
      RECT  76.67 94.18 76.88 94.56 ;
      RECT  75.95 94.73 76.16 94.8 ;
      RECT  76.16 93.94 76.36 94.01 ;
      RECT  73.76 93.7 76.16 93.94 ;
      RECT  76.67 93.7 76.88 93.94 ;
      RECT  74.69 92.91 75.23 93.46 ;
      RECT  73.55 94.18 74.69 94.56 ;
      RECT  73.55 92.91 73.76 93.46 ;
      POLYGON  76.53 94.18 76.53 94.25 76.16 94.25 76.16 94.49 76.53 94.49 76.53 94.56 76.67 94.56 76.67 94.18 76.53 94.18 ;
      RECT  76.16 93.7 76.67 93.94 ;
      RECT  75.23 92.91 76.88 93.46 ;
      POLYGON  75.23 94.18 75.23 94.56 75.78 94.56 75.78 94.49 76.16 94.49 76.16 94.25 75.78 94.25 75.78 94.18 75.23 94.18 ;
      RECT  73.55 93.7 73.76 93.94 ;
      RECT  77.6 94.8 77.09 95.04 ;
      RECT  77.6 94.73 77.4 94.8 ;
      RECT  79.07 94.18 78.53 94.56 ;
      RECT  80.0 92.91 79.07 93.46 ;
      RECT  80.21 94.8 80.0 95.04 ;
      RECT  77.09 94.8 76.88 95.04 ;
      RECT  80.0 94.8 77.6 95.04 ;
      RECT  77.81 93.94 77.6 94.01 ;
      RECT  77.09 94.18 76.88 94.56 ;
      RECT  77.81 94.73 77.6 94.8 ;
      RECT  77.6 93.94 77.4 94.01 ;
      RECT  80.0 93.7 77.6 93.94 ;
      RECT  77.09 93.7 76.88 93.94 ;
      RECT  79.07 92.91 78.53 93.46 ;
      RECT  80.21 94.18 79.07 94.56 ;
      RECT  80.21 92.91 80.0 93.46 ;
      POLYGON  77.23 94.18 77.23 94.25 77.6 94.25 77.6 94.49 77.23 94.49 77.23 94.56 77.09 94.56 77.09 94.18 77.23 94.18 ;
      RECT  77.6 93.7 77.09 93.94 ;
      RECT  78.53 92.91 76.88 93.46 ;
      POLYGON  78.53 94.18 78.53 94.56 77.98 94.56 77.98 94.49 77.6 94.49 77.6 94.25 77.98 94.25 77.98 94.18 78.53 94.18 ;
      RECT  80.21 93.7 80.0 93.94 ;
      RECT  73.76 94.8 80.0 95.04 ;
      RECT  73.76 93.7 80.0 93.94 ;
      RECT  74.69 92.91 75.23 93.46 ;
      RECT  74.69 94.18 75.23 94.56 ;
      RECT  78.53 94.18 79.07 94.56 ;
      RECT  78.53 92.91 79.07 93.46 ;
      RECT  73.76 58.505 76.88 59.055 ;
      RECT  80.0 58.505 76.88 59.055 ;
      RECT  73.76 96.265 76.88 95.715 ;
      RECT  80.0 96.265 76.88 95.715 ;
      RECT  69.92 59.97 70.43 59.73 ;
      RECT  69.92 60.04 70.12 59.97 ;
      RECT  68.45 60.59 68.99 60.21 ;
      RECT  67.52 61.86 68.45 61.31 ;
      RECT  67.31 59.97 67.52 59.73 ;
      RECT  70.43 59.97 70.64 59.73 ;
      RECT  67.52 59.97 69.92 59.73 ;
      RECT  69.71 60.83 69.92 60.76 ;
      RECT  70.43 60.59 70.64 60.21 ;
      RECT  69.71 60.04 69.92 59.97 ;
      RECT  69.92 60.83 70.12 60.76 ;
      RECT  67.52 61.07 69.92 60.83 ;
      RECT  70.43 61.07 70.64 60.83 ;
      RECT  68.45 61.86 68.99 61.31 ;
      RECT  67.31 60.59 68.45 60.21 ;
      RECT  67.31 61.86 67.52 61.31 ;
      POLYGON  70.29 60.59 70.29 60.52 69.92 60.52 69.92 60.28 70.29 60.28 70.29 60.21 70.43 60.21 70.43 60.59 70.29 60.59 ;
      RECT  69.92 61.07 70.43 60.83 ;
      RECT  68.99 61.86 70.64 61.31 ;
      POLYGON  68.99 60.59 68.99 60.21 69.54 60.21 69.54 60.28 69.92 60.28 69.92 60.52 69.54 60.52 69.54 60.59 68.99 60.59 ;
      RECT  67.31 61.07 67.52 60.83 ;
      RECT  69.92 63.2 70.43 63.44 ;
      RECT  69.92 63.13 70.12 63.2 ;
      RECT  68.45 62.58 68.99 62.96 ;
      RECT  67.52 61.31 68.45 61.86 ;
      RECT  67.31 63.2 67.52 63.44 ;
      RECT  70.43 63.2 70.64 63.44 ;
      RECT  67.52 63.2 69.92 63.44 ;
      RECT  69.71 62.34 69.92 62.41 ;
      RECT  70.43 62.58 70.64 62.96 ;
      RECT  69.71 63.13 69.92 63.2 ;
      RECT  69.92 62.34 70.12 62.41 ;
      RECT  67.52 62.1 69.92 62.34 ;
      RECT  70.43 62.1 70.64 62.34 ;
      RECT  68.45 61.31 68.99 61.86 ;
      RECT  67.31 62.58 68.45 62.96 ;
      RECT  67.31 61.31 67.52 61.86 ;
      POLYGON  70.29 62.58 70.29 62.65 69.92 62.65 69.92 62.89 70.29 62.89 70.29 62.96 70.43 62.96 70.43 62.58 70.29 62.58 ;
      RECT  69.92 62.1 70.43 62.34 ;
      RECT  68.99 61.31 70.64 61.86 ;
      POLYGON  68.99 62.58 68.99 62.96 69.54 62.96 69.54 62.89 69.92 62.89 69.92 62.65 69.54 62.65 69.54 62.58 68.99 62.58 ;
      RECT  67.31 62.1 67.52 62.34 ;
      RECT  69.92 63.92 70.43 63.68 ;
      RECT  69.92 63.99 70.12 63.92 ;
      RECT  68.45 64.54 68.99 64.16 ;
      RECT  67.52 65.81 68.45 65.26 ;
      RECT  67.31 63.92 67.52 63.68 ;
      RECT  70.43 63.92 70.64 63.68 ;
      RECT  67.52 63.92 69.92 63.68 ;
      RECT  69.71 64.78 69.92 64.71 ;
      RECT  70.43 64.54 70.64 64.16 ;
      RECT  69.71 63.99 69.92 63.92 ;
      RECT  69.92 64.78 70.12 64.71 ;
      RECT  67.52 65.02 69.92 64.78 ;
      RECT  70.43 65.02 70.64 64.78 ;
      RECT  68.45 65.81 68.99 65.26 ;
      RECT  67.31 64.54 68.45 64.16 ;
      RECT  67.31 65.81 67.52 65.26 ;
      POLYGON  70.29 64.54 70.29 64.47 69.92 64.47 69.92 64.23 70.29 64.23 70.29 64.16 70.43 64.16 70.43 64.54 70.29 64.54 ;
      RECT  69.92 65.02 70.43 64.78 ;
      RECT  68.99 65.81 70.64 65.26 ;
      POLYGON  68.99 64.54 68.99 64.16 69.54 64.16 69.54 64.23 69.92 64.23 69.92 64.47 69.54 64.47 69.54 64.54 68.99 64.54 ;
      RECT  67.31 65.02 67.52 64.78 ;
      RECT  69.92 67.15 70.43 67.39 ;
      RECT  69.92 67.08 70.12 67.15 ;
      RECT  68.45 66.53 68.99 66.91 ;
      RECT  67.52 65.26 68.45 65.81 ;
      RECT  67.31 67.15 67.52 67.39 ;
      RECT  70.43 67.15 70.64 67.39 ;
      RECT  67.52 67.15 69.92 67.39 ;
      RECT  69.71 66.29 69.92 66.36 ;
      RECT  70.43 66.53 70.64 66.91 ;
      RECT  69.71 67.08 69.92 67.15 ;
      RECT  69.92 66.29 70.12 66.36 ;
      RECT  67.52 66.05 69.92 66.29 ;
      RECT  70.43 66.05 70.64 66.29 ;
      RECT  68.45 65.26 68.99 65.81 ;
      RECT  67.31 66.53 68.45 66.91 ;
      RECT  67.31 65.26 67.52 65.81 ;
      POLYGON  70.29 66.53 70.29 66.6 69.92 66.6 69.92 66.84 70.29 66.84 70.29 66.91 70.43 66.91 70.43 66.53 70.29 66.53 ;
      RECT  69.92 66.05 70.43 66.29 ;
      RECT  68.99 65.26 70.64 65.81 ;
      POLYGON  68.99 66.53 68.99 66.91 69.54 66.91 69.54 66.84 69.92 66.84 69.92 66.6 69.54 66.6 69.54 66.53 68.99 66.53 ;
      RECT  67.31 66.05 67.52 66.29 ;
      RECT  69.92 67.87 70.43 67.63 ;
      RECT  69.92 67.94 70.12 67.87 ;
      RECT  68.45 68.49 68.99 68.11 ;
      RECT  67.52 69.76 68.45 69.21 ;
      RECT  67.31 67.87 67.52 67.63 ;
      RECT  70.43 67.87 70.64 67.63 ;
      RECT  67.52 67.87 69.92 67.63 ;
      RECT  69.71 68.73 69.92 68.66 ;
      RECT  70.43 68.49 70.64 68.11 ;
      RECT  69.71 67.94 69.92 67.87 ;
      RECT  69.92 68.73 70.12 68.66 ;
      RECT  67.52 68.97 69.92 68.73 ;
      RECT  70.43 68.97 70.64 68.73 ;
      RECT  68.45 69.76 68.99 69.21 ;
      RECT  67.31 68.49 68.45 68.11 ;
      RECT  67.31 69.76 67.52 69.21 ;
      POLYGON  70.29 68.49 70.29 68.42 69.92 68.42 69.92 68.18 70.29 68.18 70.29 68.11 70.43 68.11 70.43 68.49 70.29 68.49 ;
      RECT  69.92 68.97 70.43 68.73 ;
      RECT  68.99 69.76 70.64 69.21 ;
      POLYGON  68.99 68.49 68.99 68.11 69.54 68.11 69.54 68.18 69.92 68.18 69.92 68.42 69.54 68.42 69.54 68.49 68.99 68.49 ;
      RECT  67.31 68.97 67.52 68.73 ;
      RECT  69.92 71.1 70.43 71.34 ;
      RECT  69.92 71.03 70.12 71.1 ;
      RECT  68.45 70.48 68.99 70.86 ;
      RECT  67.52 69.21 68.45 69.76 ;
      RECT  67.31 71.1 67.52 71.34 ;
      RECT  70.43 71.1 70.64 71.34 ;
      RECT  67.52 71.1 69.92 71.34 ;
      RECT  69.71 70.24 69.92 70.31 ;
      RECT  70.43 70.48 70.64 70.86 ;
      RECT  69.71 71.03 69.92 71.1 ;
      RECT  69.92 70.24 70.12 70.31 ;
      RECT  67.52 70.0 69.92 70.24 ;
      RECT  70.43 70.0 70.64 70.24 ;
      RECT  68.45 69.21 68.99 69.76 ;
      RECT  67.31 70.48 68.45 70.86 ;
      RECT  67.31 69.21 67.52 69.76 ;
      POLYGON  70.29 70.48 70.29 70.55 69.92 70.55 69.92 70.79 70.29 70.79 70.29 70.86 70.43 70.86 70.43 70.48 70.29 70.48 ;
      RECT  69.92 70.0 70.43 70.24 ;
      RECT  68.99 69.21 70.64 69.76 ;
      POLYGON  68.99 70.48 68.99 70.86 69.54 70.86 69.54 70.79 69.92 70.79 69.92 70.55 69.54 70.55 69.54 70.48 68.99 70.48 ;
      RECT  67.31 70.0 67.52 70.24 ;
      RECT  69.92 71.82 70.43 71.58 ;
      RECT  69.92 71.89 70.12 71.82 ;
      RECT  68.45 72.44 68.99 72.06 ;
      RECT  67.52 73.71 68.45 73.16 ;
      RECT  67.31 71.82 67.52 71.58 ;
      RECT  70.43 71.82 70.64 71.58 ;
      RECT  67.52 71.82 69.92 71.58 ;
      RECT  69.71 72.68 69.92 72.61 ;
      RECT  70.43 72.44 70.64 72.06 ;
      RECT  69.71 71.89 69.92 71.82 ;
      RECT  69.92 72.68 70.12 72.61 ;
      RECT  67.52 72.92 69.92 72.68 ;
      RECT  70.43 72.92 70.64 72.68 ;
      RECT  68.45 73.71 68.99 73.16 ;
      RECT  67.31 72.44 68.45 72.06 ;
      RECT  67.31 73.71 67.52 73.16 ;
      POLYGON  70.29 72.44 70.29 72.37 69.92 72.37 69.92 72.13 70.29 72.13 70.29 72.06 70.43 72.06 70.43 72.44 70.29 72.44 ;
      RECT  69.92 72.92 70.43 72.68 ;
      RECT  68.99 73.71 70.64 73.16 ;
      POLYGON  68.99 72.44 68.99 72.06 69.54 72.06 69.54 72.13 69.92 72.13 69.92 72.37 69.54 72.37 69.54 72.44 68.99 72.44 ;
      RECT  67.31 72.92 67.52 72.68 ;
      RECT  69.92 75.05 70.43 75.29 ;
      RECT  69.92 74.98 70.12 75.05 ;
      RECT  68.45 74.43 68.99 74.81 ;
      RECT  67.52 73.16 68.45 73.71 ;
      RECT  67.31 75.05 67.52 75.29 ;
      RECT  70.43 75.05 70.64 75.29 ;
      RECT  67.52 75.05 69.92 75.29 ;
      RECT  69.71 74.19 69.92 74.26 ;
      RECT  70.43 74.43 70.64 74.81 ;
      RECT  69.71 74.98 69.92 75.05 ;
      RECT  69.92 74.19 70.12 74.26 ;
      RECT  67.52 73.95 69.92 74.19 ;
      RECT  70.43 73.95 70.64 74.19 ;
      RECT  68.45 73.16 68.99 73.71 ;
      RECT  67.31 74.43 68.45 74.81 ;
      RECT  67.31 73.16 67.52 73.71 ;
      POLYGON  70.29 74.43 70.29 74.5 69.92 74.5 69.92 74.74 70.29 74.74 70.29 74.81 70.43 74.81 70.43 74.43 70.29 74.43 ;
      RECT  69.92 73.95 70.43 74.19 ;
      RECT  68.99 73.16 70.64 73.71 ;
      POLYGON  68.99 74.43 68.99 74.81 69.54 74.81 69.54 74.74 69.92 74.74 69.92 74.5 69.54 74.5 69.54 74.43 68.99 74.43 ;
      RECT  67.31 73.95 67.52 74.19 ;
      RECT  69.92 75.77 70.43 75.53 ;
      RECT  69.92 75.84 70.12 75.77 ;
      RECT  68.45 76.39 68.99 76.01 ;
      RECT  67.52 77.66 68.45 77.11 ;
      RECT  67.31 75.77 67.52 75.53 ;
      RECT  70.43 75.77 70.64 75.53 ;
      RECT  67.52 75.77 69.92 75.53 ;
      RECT  69.71 76.63 69.92 76.56 ;
      RECT  70.43 76.39 70.64 76.01 ;
      RECT  69.71 75.84 69.92 75.77 ;
      RECT  69.92 76.63 70.12 76.56 ;
      RECT  67.52 76.87 69.92 76.63 ;
      RECT  70.43 76.87 70.64 76.63 ;
      RECT  68.45 77.66 68.99 77.11 ;
      RECT  67.31 76.39 68.45 76.01 ;
      RECT  67.31 77.66 67.52 77.11 ;
      POLYGON  70.29 76.39 70.29 76.32 69.92 76.32 69.92 76.08 70.29 76.08 70.29 76.01 70.43 76.01 70.43 76.39 70.29 76.39 ;
      RECT  69.92 76.87 70.43 76.63 ;
      RECT  68.99 77.66 70.64 77.11 ;
      POLYGON  68.99 76.39 68.99 76.01 69.54 76.01 69.54 76.08 69.92 76.08 69.92 76.32 69.54 76.32 69.54 76.39 68.99 76.39 ;
      RECT  67.31 76.87 67.52 76.63 ;
      RECT  69.92 79.0 70.43 79.24 ;
      RECT  69.92 78.93 70.12 79.0 ;
      RECT  68.45 78.38 68.99 78.76 ;
      RECT  67.52 77.11 68.45 77.66 ;
      RECT  67.31 79.0 67.52 79.24 ;
      RECT  70.43 79.0 70.64 79.24 ;
      RECT  67.52 79.0 69.92 79.24 ;
      RECT  69.71 78.14 69.92 78.21 ;
      RECT  70.43 78.38 70.64 78.76 ;
      RECT  69.71 78.93 69.92 79.0 ;
      RECT  69.92 78.14 70.12 78.21 ;
      RECT  67.52 77.9 69.92 78.14 ;
      RECT  70.43 77.9 70.64 78.14 ;
      RECT  68.45 77.11 68.99 77.66 ;
      RECT  67.31 78.38 68.45 78.76 ;
      RECT  67.31 77.11 67.52 77.66 ;
      POLYGON  70.29 78.38 70.29 78.45 69.92 78.45 69.92 78.69 70.29 78.69 70.29 78.76 70.43 78.76 70.43 78.38 70.29 78.38 ;
      RECT  69.92 77.9 70.43 78.14 ;
      RECT  68.99 77.11 70.64 77.66 ;
      POLYGON  68.99 78.38 68.99 78.76 69.54 78.76 69.54 78.69 69.92 78.69 69.92 78.45 69.54 78.45 69.54 78.38 68.99 78.38 ;
      RECT  67.31 77.9 67.52 78.14 ;
      RECT  69.92 79.72 70.43 79.48 ;
      RECT  69.92 79.79 70.12 79.72 ;
      RECT  68.45 80.34 68.99 79.96 ;
      RECT  67.52 81.61 68.45 81.06 ;
      RECT  67.31 79.72 67.52 79.48 ;
      RECT  70.43 79.72 70.64 79.48 ;
      RECT  67.52 79.72 69.92 79.48 ;
      RECT  69.71 80.58 69.92 80.51 ;
      RECT  70.43 80.34 70.64 79.96 ;
      RECT  69.71 79.79 69.92 79.72 ;
      RECT  69.92 80.58 70.12 80.51 ;
      RECT  67.52 80.82 69.92 80.58 ;
      RECT  70.43 80.82 70.64 80.58 ;
      RECT  68.45 81.61 68.99 81.06 ;
      RECT  67.31 80.34 68.45 79.96 ;
      RECT  67.31 81.61 67.52 81.06 ;
      POLYGON  70.29 80.34 70.29 80.27 69.92 80.27 69.92 80.03 70.29 80.03 70.29 79.96 70.43 79.96 70.43 80.34 70.29 80.34 ;
      RECT  69.92 80.82 70.43 80.58 ;
      RECT  68.99 81.61 70.64 81.06 ;
      POLYGON  68.99 80.34 68.99 79.96 69.54 79.96 69.54 80.03 69.92 80.03 69.92 80.27 69.54 80.27 69.54 80.34 68.99 80.34 ;
      RECT  67.31 80.82 67.52 80.58 ;
      RECT  69.92 82.95 70.43 83.19 ;
      RECT  69.92 82.88 70.12 82.95 ;
      RECT  68.45 82.33 68.99 82.71 ;
      RECT  67.52 81.06 68.45 81.61 ;
      RECT  67.31 82.95 67.52 83.19 ;
      RECT  70.43 82.95 70.64 83.19 ;
      RECT  67.52 82.95 69.92 83.19 ;
      RECT  69.71 82.09 69.92 82.16 ;
      RECT  70.43 82.33 70.64 82.71 ;
      RECT  69.71 82.88 69.92 82.95 ;
      RECT  69.92 82.09 70.12 82.16 ;
      RECT  67.52 81.85 69.92 82.09 ;
      RECT  70.43 81.85 70.64 82.09 ;
      RECT  68.45 81.06 68.99 81.61 ;
      RECT  67.31 82.33 68.45 82.71 ;
      RECT  67.31 81.06 67.52 81.61 ;
      POLYGON  70.29 82.33 70.29 82.4 69.92 82.4 69.92 82.64 70.29 82.64 70.29 82.71 70.43 82.71 70.43 82.33 70.29 82.33 ;
      RECT  69.92 81.85 70.43 82.09 ;
      RECT  68.99 81.06 70.64 81.61 ;
      POLYGON  68.99 82.33 68.99 82.71 69.54 82.71 69.54 82.64 69.92 82.64 69.92 82.4 69.54 82.4 69.54 82.33 68.99 82.33 ;
      RECT  67.31 81.85 67.52 82.09 ;
      RECT  69.92 83.67 70.43 83.43 ;
      RECT  69.92 83.74 70.12 83.67 ;
      RECT  68.45 84.29 68.99 83.91 ;
      RECT  67.52 85.56 68.45 85.01 ;
      RECT  67.31 83.67 67.52 83.43 ;
      RECT  70.43 83.67 70.64 83.43 ;
      RECT  67.52 83.67 69.92 83.43 ;
      RECT  69.71 84.53 69.92 84.46 ;
      RECT  70.43 84.29 70.64 83.91 ;
      RECT  69.71 83.74 69.92 83.67 ;
      RECT  69.92 84.53 70.12 84.46 ;
      RECT  67.52 84.77 69.92 84.53 ;
      RECT  70.43 84.77 70.64 84.53 ;
      RECT  68.45 85.56 68.99 85.01 ;
      RECT  67.31 84.29 68.45 83.91 ;
      RECT  67.31 85.56 67.52 85.01 ;
      POLYGON  70.29 84.29 70.29 84.22 69.92 84.22 69.92 83.98 70.29 83.98 70.29 83.91 70.43 83.91 70.43 84.29 70.29 84.29 ;
      RECT  69.92 84.77 70.43 84.53 ;
      RECT  68.99 85.56 70.64 85.01 ;
      POLYGON  68.99 84.29 68.99 83.91 69.54 83.91 69.54 83.98 69.92 83.98 69.92 84.22 69.54 84.22 69.54 84.29 68.99 84.29 ;
      RECT  67.31 84.77 67.52 84.53 ;
      RECT  69.92 86.9 70.43 87.14 ;
      RECT  69.92 86.83 70.12 86.9 ;
      RECT  68.45 86.28 68.99 86.66 ;
      RECT  67.52 85.01 68.45 85.56 ;
      RECT  67.31 86.9 67.52 87.14 ;
      RECT  70.43 86.9 70.64 87.14 ;
      RECT  67.52 86.9 69.92 87.14 ;
      RECT  69.71 86.04 69.92 86.11 ;
      RECT  70.43 86.28 70.64 86.66 ;
      RECT  69.71 86.83 69.92 86.9 ;
      RECT  69.92 86.04 70.12 86.11 ;
      RECT  67.52 85.8 69.92 86.04 ;
      RECT  70.43 85.8 70.64 86.04 ;
      RECT  68.45 85.01 68.99 85.56 ;
      RECT  67.31 86.28 68.45 86.66 ;
      RECT  67.31 85.01 67.52 85.56 ;
      POLYGON  70.29 86.28 70.29 86.35 69.92 86.35 69.92 86.59 70.29 86.59 70.29 86.66 70.43 86.66 70.43 86.28 70.29 86.28 ;
      RECT  69.92 85.8 70.43 86.04 ;
      RECT  68.99 85.01 70.64 85.56 ;
      POLYGON  68.99 86.28 68.99 86.66 69.54 86.66 69.54 86.59 69.92 86.59 69.92 86.35 69.54 86.35 69.54 86.28 68.99 86.28 ;
      RECT  67.31 85.8 67.52 86.04 ;
      RECT  69.92 87.62 70.43 87.38 ;
      RECT  69.92 87.69 70.12 87.62 ;
      RECT  68.45 88.24 68.99 87.86 ;
      RECT  67.52 89.51 68.45 88.96 ;
      RECT  67.31 87.62 67.52 87.38 ;
      RECT  70.43 87.62 70.64 87.38 ;
      RECT  67.52 87.62 69.92 87.38 ;
      RECT  69.71 88.48 69.92 88.41 ;
      RECT  70.43 88.24 70.64 87.86 ;
      RECT  69.71 87.69 69.92 87.62 ;
      RECT  69.92 88.48 70.12 88.41 ;
      RECT  67.52 88.72 69.92 88.48 ;
      RECT  70.43 88.72 70.64 88.48 ;
      RECT  68.45 89.51 68.99 88.96 ;
      RECT  67.31 88.24 68.45 87.86 ;
      RECT  67.31 89.51 67.52 88.96 ;
      POLYGON  70.29 88.24 70.29 88.17 69.92 88.17 69.92 87.93 70.29 87.93 70.29 87.86 70.43 87.86 70.43 88.24 70.29 88.24 ;
      RECT  69.92 88.72 70.43 88.48 ;
      RECT  68.99 89.51 70.64 88.96 ;
      POLYGON  68.99 88.24 68.99 87.86 69.54 87.86 69.54 87.93 69.92 87.93 69.92 88.17 69.54 88.17 69.54 88.24 68.99 88.24 ;
      RECT  67.31 88.72 67.52 88.48 ;
      RECT  69.92 90.85 70.43 91.09 ;
      RECT  69.92 90.78 70.12 90.85 ;
      RECT  68.45 90.23 68.99 90.61 ;
      RECT  67.52 88.96 68.45 89.51 ;
      RECT  67.31 90.85 67.52 91.09 ;
      RECT  70.43 90.85 70.64 91.09 ;
      RECT  67.52 90.85 69.92 91.09 ;
      RECT  69.71 89.99 69.92 90.06 ;
      RECT  70.43 90.23 70.64 90.61 ;
      RECT  69.71 90.78 69.92 90.85 ;
      RECT  69.92 89.99 70.12 90.06 ;
      RECT  67.52 89.75 69.92 89.99 ;
      RECT  70.43 89.75 70.64 89.99 ;
      RECT  68.45 88.96 68.99 89.51 ;
      RECT  67.31 90.23 68.45 90.61 ;
      RECT  67.31 88.96 67.52 89.51 ;
      POLYGON  70.29 90.23 70.29 90.3 69.92 90.3 69.92 90.54 70.29 90.54 70.29 90.61 70.43 90.61 70.43 90.23 70.29 90.23 ;
      RECT  69.92 89.75 70.43 89.99 ;
      RECT  68.99 88.96 70.64 89.51 ;
      POLYGON  68.99 90.23 68.99 90.61 69.54 90.61 69.54 90.54 69.92 90.54 69.92 90.3 69.54 90.3 69.54 90.23 68.99 90.23 ;
      RECT  67.31 89.75 67.52 89.99 ;
      RECT  69.92 91.57 70.43 91.33 ;
      RECT  69.92 91.64 70.12 91.57 ;
      RECT  68.45 92.19 68.99 91.81 ;
      RECT  67.52 93.46 68.45 92.91 ;
      RECT  67.31 91.57 67.52 91.33 ;
      RECT  70.43 91.57 70.64 91.33 ;
      RECT  67.52 91.57 69.92 91.33 ;
      RECT  69.71 92.43 69.92 92.36 ;
      RECT  70.43 92.19 70.64 91.81 ;
      RECT  69.71 91.64 69.92 91.57 ;
      RECT  69.92 92.43 70.12 92.36 ;
      RECT  67.52 92.67 69.92 92.43 ;
      RECT  70.43 92.67 70.64 92.43 ;
      RECT  68.45 93.46 68.99 92.91 ;
      RECT  67.31 92.19 68.45 91.81 ;
      RECT  67.31 93.46 67.52 92.91 ;
      POLYGON  70.29 92.19 70.29 92.12 69.92 92.12 69.92 91.88 70.29 91.88 70.29 91.81 70.43 91.81 70.43 92.19 70.29 92.19 ;
      RECT  69.92 92.67 70.43 92.43 ;
      RECT  68.99 93.46 70.64 92.91 ;
      POLYGON  68.99 92.19 68.99 91.81 69.54 91.81 69.54 91.88 69.92 91.88 69.92 92.12 69.54 92.12 69.54 92.19 68.99 92.19 ;
      RECT  67.31 92.67 67.52 92.43 ;
      RECT  69.92 94.8 70.43 95.04 ;
      RECT  69.92 94.73 70.12 94.8 ;
      RECT  68.45 94.18 68.99 94.56 ;
      RECT  67.52 92.91 68.45 93.46 ;
      RECT  67.31 94.8 67.52 95.04 ;
      RECT  70.43 94.8 70.64 95.04 ;
      RECT  67.52 94.8 69.92 95.04 ;
      RECT  69.71 93.94 69.92 94.01 ;
      RECT  70.43 94.18 70.64 94.56 ;
      RECT  69.71 94.73 69.92 94.8 ;
      RECT  69.92 93.94 70.12 94.01 ;
      RECT  67.52 93.7 69.92 93.94 ;
      RECT  70.43 93.7 70.64 93.94 ;
      RECT  68.45 92.91 68.99 93.46 ;
      RECT  67.31 94.18 68.45 94.56 ;
      RECT  67.31 92.91 67.52 93.46 ;
      POLYGON  70.29 94.18 70.29 94.25 69.92 94.25 69.92 94.49 70.29 94.49 70.29 94.56 70.43 94.56 70.43 94.18 70.29 94.18 ;
      RECT  69.92 93.7 70.43 93.94 ;
      RECT  68.99 92.91 70.64 93.46 ;
      POLYGON  68.99 94.18 68.99 94.56 69.54 94.56 69.54 94.49 69.92 94.49 69.92 94.25 69.54 94.25 69.54 94.18 68.99 94.18 ;
      RECT  67.31 93.7 67.52 93.94 ;
      RECT  67.52 59.73 70.64 59.97 ;
      RECT  67.52 60.83 70.64 61.07 ;
      RECT  67.52 63.2 70.64 63.44 ;
      RECT  67.52 62.1 70.64 62.34 ;
      RECT  67.52 63.68 70.64 63.92 ;
      RECT  67.52 64.78 70.64 65.02 ;
      RECT  67.52 67.15 70.64 67.39 ;
      RECT  67.52 66.05 70.64 66.29 ;
      RECT  67.52 67.63 70.64 67.87 ;
      RECT  67.52 68.73 70.64 68.97 ;
      RECT  67.52 71.1 70.64 71.34 ;
      RECT  67.52 70.0 70.64 70.24 ;
      RECT  67.52 71.58 70.64 71.82 ;
      RECT  67.52 72.68 70.64 72.92 ;
      RECT  67.52 75.05 70.64 75.29 ;
      RECT  67.52 73.95 70.64 74.19 ;
      RECT  67.52 75.53 70.64 75.77 ;
      RECT  67.52 76.63 70.64 76.87 ;
      RECT  67.52 79.0 70.64 79.24 ;
      RECT  67.52 77.9 70.64 78.14 ;
      RECT  67.52 79.48 70.64 79.72 ;
      RECT  67.52 80.58 70.64 80.82 ;
      RECT  67.52 82.95 70.64 83.19 ;
      RECT  67.52 81.85 70.64 82.09 ;
      RECT  67.52 83.43 70.64 83.67 ;
      RECT  67.52 84.53 70.64 84.77 ;
      RECT  67.52 86.9 70.64 87.14 ;
      RECT  67.52 85.8 70.64 86.04 ;
      RECT  67.52 87.38 70.64 87.62 ;
      RECT  67.52 88.48 70.64 88.72 ;
      RECT  67.52 90.85 70.64 91.09 ;
      RECT  67.52 89.75 70.64 89.99 ;
      RECT  67.52 91.33 70.64 91.57 ;
      RECT  67.52 92.43 70.64 92.67 ;
      RECT  67.52 94.8 70.64 95.04 ;
      RECT  67.52 93.7 70.64 93.94 ;
      RECT  83.84 59.97 83.33 59.73 ;
      RECT  83.84 60.04 83.64 59.97 ;
      RECT  85.31 60.59 84.77 60.21 ;
      RECT  86.24 61.86 85.31 61.31 ;
      RECT  86.45 59.97 86.24 59.73 ;
      RECT  83.33 59.97 83.12 59.73 ;
      RECT  86.24 59.97 83.84 59.73 ;
      RECT  84.05 60.83 83.84 60.76 ;
      RECT  83.33 60.59 83.12 60.21 ;
      RECT  84.05 60.04 83.84 59.97 ;
      RECT  83.84 60.83 83.64 60.76 ;
      RECT  86.24 61.07 83.84 60.83 ;
      RECT  83.33 61.07 83.12 60.83 ;
      RECT  85.31 61.86 84.77 61.31 ;
      RECT  86.45 60.59 85.31 60.21 ;
      RECT  86.45 61.86 86.24 61.31 ;
      POLYGON  83.47 60.59 83.47 60.52 83.84 60.52 83.84 60.28 83.47 60.28 83.47 60.21 83.33 60.21 83.33 60.59 83.47 60.59 ;
      RECT  83.84 61.07 83.33 60.83 ;
      RECT  84.77 61.86 83.12 61.31 ;
      POLYGON  84.77 60.59 84.77 60.21 84.22 60.21 84.22 60.28 83.84 60.28 83.84 60.52 84.22 60.52 84.22 60.59 84.77 60.59 ;
      RECT  86.45 61.07 86.24 60.83 ;
      RECT  83.84 63.2 83.33 63.44 ;
      RECT  83.84 63.13 83.64 63.2 ;
      RECT  85.31 62.58 84.77 62.96 ;
      RECT  86.24 61.31 85.31 61.86 ;
      RECT  86.45 63.2 86.24 63.44 ;
      RECT  83.33 63.2 83.12 63.44 ;
      RECT  86.24 63.2 83.84 63.44 ;
      RECT  84.05 62.34 83.84 62.41 ;
      RECT  83.33 62.58 83.12 62.96 ;
      RECT  84.05 63.13 83.84 63.2 ;
      RECT  83.84 62.34 83.64 62.41 ;
      RECT  86.24 62.1 83.84 62.34 ;
      RECT  83.33 62.1 83.12 62.34 ;
      RECT  85.31 61.31 84.77 61.86 ;
      RECT  86.45 62.58 85.31 62.96 ;
      RECT  86.45 61.31 86.24 61.86 ;
      POLYGON  83.47 62.58 83.47 62.65 83.84 62.65 83.84 62.89 83.47 62.89 83.47 62.96 83.33 62.96 83.33 62.58 83.47 62.58 ;
      RECT  83.84 62.1 83.33 62.34 ;
      RECT  84.77 61.31 83.12 61.86 ;
      POLYGON  84.77 62.58 84.77 62.96 84.22 62.96 84.22 62.89 83.84 62.89 83.84 62.65 84.22 62.65 84.22 62.58 84.77 62.58 ;
      RECT  86.45 62.1 86.24 62.34 ;
      RECT  83.84 63.92 83.33 63.68 ;
      RECT  83.84 63.99 83.64 63.92 ;
      RECT  85.31 64.54 84.77 64.16 ;
      RECT  86.24 65.81 85.31 65.26 ;
      RECT  86.45 63.92 86.24 63.68 ;
      RECT  83.33 63.92 83.12 63.68 ;
      RECT  86.24 63.92 83.84 63.68 ;
      RECT  84.05 64.78 83.84 64.71 ;
      RECT  83.33 64.54 83.12 64.16 ;
      RECT  84.05 63.99 83.84 63.92 ;
      RECT  83.84 64.78 83.64 64.71 ;
      RECT  86.24 65.02 83.84 64.78 ;
      RECT  83.33 65.02 83.12 64.78 ;
      RECT  85.31 65.81 84.77 65.26 ;
      RECT  86.45 64.54 85.31 64.16 ;
      RECT  86.45 65.81 86.24 65.26 ;
      POLYGON  83.47 64.54 83.47 64.47 83.84 64.47 83.84 64.23 83.47 64.23 83.47 64.16 83.33 64.16 83.33 64.54 83.47 64.54 ;
      RECT  83.84 65.02 83.33 64.78 ;
      RECT  84.77 65.81 83.12 65.26 ;
      POLYGON  84.77 64.54 84.77 64.16 84.22 64.16 84.22 64.23 83.84 64.23 83.84 64.47 84.22 64.47 84.22 64.54 84.77 64.54 ;
      RECT  86.45 65.02 86.24 64.78 ;
      RECT  83.84 67.15 83.33 67.39 ;
      RECT  83.84 67.08 83.64 67.15 ;
      RECT  85.31 66.53 84.77 66.91 ;
      RECT  86.24 65.26 85.31 65.81 ;
      RECT  86.45 67.15 86.24 67.39 ;
      RECT  83.33 67.15 83.12 67.39 ;
      RECT  86.24 67.15 83.84 67.39 ;
      RECT  84.05 66.29 83.84 66.36 ;
      RECT  83.33 66.53 83.12 66.91 ;
      RECT  84.05 67.08 83.84 67.15 ;
      RECT  83.84 66.29 83.64 66.36 ;
      RECT  86.24 66.05 83.84 66.29 ;
      RECT  83.33 66.05 83.12 66.29 ;
      RECT  85.31 65.26 84.77 65.81 ;
      RECT  86.45 66.53 85.31 66.91 ;
      RECT  86.45 65.26 86.24 65.81 ;
      POLYGON  83.47 66.53 83.47 66.6 83.84 66.6 83.84 66.84 83.47 66.84 83.47 66.91 83.33 66.91 83.33 66.53 83.47 66.53 ;
      RECT  83.84 66.05 83.33 66.29 ;
      RECT  84.77 65.26 83.12 65.81 ;
      POLYGON  84.77 66.53 84.77 66.91 84.22 66.91 84.22 66.84 83.84 66.84 83.84 66.6 84.22 66.6 84.22 66.53 84.77 66.53 ;
      RECT  86.45 66.05 86.24 66.29 ;
      RECT  83.84 67.87 83.33 67.63 ;
      RECT  83.84 67.94 83.64 67.87 ;
      RECT  85.31 68.49 84.77 68.11 ;
      RECT  86.24 69.76 85.31 69.21 ;
      RECT  86.45 67.87 86.24 67.63 ;
      RECT  83.33 67.87 83.12 67.63 ;
      RECT  86.24 67.87 83.84 67.63 ;
      RECT  84.05 68.73 83.84 68.66 ;
      RECT  83.33 68.49 83.12 68.11 ;
      RECT  84.05 67.94 83.84 67.87 ;
      RECT  83.84 68.73 83.64 68.66 ;
      RECT  86.24 68.97 83.84 68.73 ;
      RECT  83.33 68.97 83.12 68.73 ;
      RECT  85.31 69.76 84.77 69.21 ;
      RECT  86.45 68.49 85.31 68.11 ;
      RECT  86.45 69.76 86.24 69.21 ;
      POLYGON  83.47 68.49 83.47 68.42 83.84 68.42 83.84 68.18 83.47 68.18 83.47 68.11 83.33 68.11 83.33 68.49 83.47 68.49 ;
      RECT  83.84 68.97 83.33 68.73 ;
      RECT  84.77 69.76 83.12 69.21 ;
      POLYGON  84.77 68.49 84.77 68.11 84.22 68.11 84.22 68.18 83.84 68.18 83.84 68.42 84.22 68.42 84.22 68.49 84.77 68.49 ;
      RECT  86.45 68.97 86.24 68.73 ;
      RECT  83.84 71.1 83.33 71.34 ;
      RECT  83.84 71.03 83.64 71.1 ;
      RECT  85.31 70.48 84.77 70.86 ;
      RECT  86.24 69.21 85.31 69.76 ;
      RECT  86.45 71.1 86.24 71.34 ;
      RECT  83.33 71.1 83.12 71.34 ;
      RECT  86.24 71.1 83.84 71.34 ;
      RECT  84.05 70.24 83.84 70.31 ;
      RECT  83.33 70.48 83.12 70.86 ;
      RECT  84.05 71.03 83.84 71.1 ;
      RECT  83.84 70.24 83.64 70.31 ;
      RECT  86.24 70.0 83.84 70.24 ;
      RECT  83.33 70.0 83.12 70.24 ;
      RECT  85.31 69.21 84.77 69.76 ;
      RECT  86.45 70.48 85.31 70.86 ;
      RECT  86.45 69.21 86.24 69.76 ;
      POLYGON  83.47 70.48 83.47 70.55 83.84 70.55 83.84 70.79 83.47 70.79 83.47 70.86 83.33 70.86 83.33 70.48 83.47 70.48 ;
      RECT  83.84 70.0 83.33 70.24 ;
      RECT  84.77 69.21 83.12 69.76 ;
      POLYGON  84.77 70.48 84.77 70.86 84.22 70.86 84.22 70.79 83.84 70.79 83.84 70.55 84.22 70.55 84.22 70.48 84.77 70.48 ;
      RECT  86.45 70.0 86.24 70.24 ;
      RECT  83.84 71.82 83.33 71.58 ;
      RECT  83.84 71.89 83.64 71.82 ;
      RECT  85.31 72.44 84.77 72.06 ;
      RECT  86.24 73.71 85.31 73.16 ;
      RECT  86.45 71.82 86.24 71.58 ;
      RECT  83.33 71.82 83.12 71.58 ;
      RECT  86.24 71.82 83.84 71.58 ;
      RECT  84.05 72.68 83.84 72.61 ;
      RECT  83.33 72.44 83.12 72.06 ;
      RECT  84.05 71.89 83.84 71.82 ;
      RECT  83.84 72.68 83.64 72.61 ;
      RECT  86.24 72.92 83.84 72.68 ;
      RECT  83.33 72.92 83.12 72.68 ;
      RECT  85.31 73.71 84.77 73.16 ;
      RECT  86.45 72.44 85.31 72.06 ;
      RECT  86.45 73.71 86.24 73.16 ;
      POLYGON  83.47 72.44 83.47 72.37 83.84 72.37 83.84 72.13 83.47 72.13 83.47 72.06 83.33 72.06 83.33 72.44 83.47 72.44 ;
      RECT  83.84 72.92 83.33 72.68 ;
      RECT  84.77 73.71 83.12 73.16 ;
      POLYGON  84.77 72.44 84.77 72.06 84.22 72.06 84.22 72.13 83.84 72.13 83.84 72.37 84.22 72.37 84.22 72.44 84.77 72.44 ;
      RECT  86.45 72.92 86.24 72.68 ;
      RECT  83.84 75.05 83.33 75.29 ;
      RECT  83.84 74.98 83.64 75.05 ;
      RECT  85.31 74.43 84.77 74.81 ;
      RECT  86.24 73.16 85.31 73.71 ;
      RECT  86.45 75.05 86.24 75.29 ;
      RECT  83.33 75.05 83.12 75.29 ;
      RECT  86.24 75.05 83.84 75.29 ;
      RECT  84.05 74.19 83.84 74.26 ;
      RECT  83.33 74.43 83.12 74.81 ;
      RECT  84.05 74.98 83.84 75.05 ;
      RECT  83.84 74.19 83.64 74.26 ;
      RECT  86.24 73.95 83.84 74.19 ;
      RECT  83.33 73.95 83.12 74.19 ;
      RECT  85.31 73.16 84.77 73.71 ;
      RECT  86.45 74.43 85.31 74.81 ;
      RECT  86.45 73.16 86.24 73.71 ;
      POLYGON  83.47 74.43 83.47 74.5 83.84 74.5 83.84 74.74 83.47 74.74 83.47 74.81 83.33 74.81 83.33 74.43 83.47 74.43 ;
      RECT  83.84 73.95 83.33 74.19 ;
      RECT  84.77 73.16 83.12 73.71 ;
      POLYGON  84.77 74.43 84.77 74.81 84.22 74.81 84.22 74.74 83.84 74.74 83.84 74.5 84.22 74.5 84.22 74.43 84.77 74.43 ;
      RECT  86.45 73.95 86.24 74.19 ;
      RECT  83.84 75.77 83.33 75.53 ;
      RECT  83.84 75.84 83.64 75.77 ;
      RECT  85.31 76.39 84.77 76.01 ;
      RECT  86.24 77.66 85.31 77.11 ;
      RECT  86.45 75.77 86.24 75.53 ;
      RECT  83.33 75.77 83.12 75.53 ;
      RECT  86.24 75.77 83.84 75.53 ;
      RECT  84.05 76.63 83.84 76.56 ;
      RECT  83.33 76.39 83.12 76.01 ;
      RECT  84.05 75.84 83.84 75.77 ;
      RECT  83.84 76.63 83.64 76.56 ;
      RECT  86.24 76.87 83.84 76.63 ;
      RECT  83.33 76.87 83.12 76.63 ;
      RECT  85.31 77.66 84.77 77.11 ;
      RECT  86.45 76.39 85.31 76.01 ;
      RECT  86.45 77.66 86.24 77.11 ;
      POLYGON  83.47 76.39 83.47 76.32 83.84 76.32 83.84 76.08 83.47 76.08 83.47 76.01 83.33 76.01 83.33 76.39 83.47 76.39 ;
      RECT  83.84 76.87 83.33 76.63 ;
      RECT  84.77 77.66 83.12 77.11 ;
      POLYGON  84.77 76.39 84.77 76.01 84.22 76.01 84.22 76.08 83.84 76.08 83.84 76.32 84.22 76.32 84.22 76.39 84.77 76.39 ;
      RECT  86.45 76.87 86.24 76.63 ;
      RECT  83.84 79.0 83.33 79.24 ;
      RECT  83.84 78.93 83.64 79.0 ;
      RECT  85.31 78.38 84.77 78.76 ;
      RECT  86.24 77.11 85.31 77.66 ;
      RECT  86.45 79.0 86.24 79.24 ;
      RECT  83.33 79.0 83.12 79.24 ;
      RECT  86.24 79.0 83.84 79.24 ;
      RECT  84.05 78.14 83.84 78.21 ;
      RECT  83.33 78.38 83.12 78.76 ;
      RECT  84.05 78.93 83.84 79.0 ;
      RECT  83.84 78.14 83.64 78.21 ;
      RECT  86.24 77.9 83.84 78.14 ;
      RECT  83.33 77.9 83.12 78.14 ;
      RECT  85.31 77.11 84.77 77.66 ;
      RECT  86.45 78.38 85.31 78.76 ;
      RECT  86.45 77.11 86.24 77.66 ;
      POLYGON  83.47 78.38 83.47 78.45 83.84 78.45 83.84 78.69 83.47 78.69 83.47 78.76 83.33 78.76 83.33 78.38 83.47 78.38 ;
      RECT  83.84 77.9 83.33 78.14 ;
      RECT  84.77 77.11 83.12 77.66 ;
      POLYGON  84.77 78.38 84.77 78.76 84.22 78.76 84.22 78.69 83.84 78.69 83.84 78.45 84.22 78.45 84.22 78.38 84.77 78.38 ;
      RECT  86.45 77.9 86.24 78.14 ;
      RECT  83.84 79.72 83.33 79.48 ;
      RECT  83.84 79.79 83.64 79.72 ;
      RECT  85.31 80.34 84.77 79.96 ;
      RECT  86.24 81.61 85.31 81.06 ;
      RECT  86.45 79.72 86.24 79.48 ;
      RECT  83.33 79.72 83.12 79.48 ;
      RECT  86.24 79.72 83.84 79.48 ;
      RECT  84.05 80.58 83.84 80.51 ;
      RECT  83.33 80.34 83.12 79.96 ;
      RECT  84.05 79.79 83.84 79.72 ;
      RECT  83.84 80.58 83.64 80.51 ;
      RECT  86.24 80.82 83.84 80.58 ;
      RECT  83.33 80.82 83.12 80.58 ;
      RECT  85.31 81.61 84.77 81.06 ;
      RECT  86.45 80.34 85.31 79.96 ;
      RECT  86.45 81.61 86.24 81.06 ;
      POLYGON  83.47 80.34 83.47 80.27 83.84 80.27 83.84 80.03 83.47 80.03 83.47 79.96 83.33 79.96 83.33 80.34 83.47 80.34 ;
      RECT  83.84 80.82 83.33 80.58 ;
      RECT  84.77 81.61 83.12 81.06 ;
      POLYGON  84.77 80.34 84.77 79.96 84.22 79.96 84.22 80.03 83.84 80.03 83.84 80.27 84.22 80.27 84.22 80.34 84.77 80.34 ;
      RECT  86.45 80.82 86.24 80.58 ;
      RECT  83.84 82.95 83.33 83.19 ;
      RECT  83.84 82.88 83.64 82.95 ;
      RECT  85.31 82.33 84.77 82.71 ;
      RECT  86.24 81.06 85.31 81.61 ;
      RECT  86.45 82.95 86.24 83.19 ;
      RECT  83.33 82.95 83.12 83.19 ;
      RECT  86.24 82.95 83.84 83.19 ;
      RECT  84.05 82.09 83.84 82.16 ;
      RECT  83.33 82.33 83.12 82.71 ;
      RECT  84.05 82.88 83.84 82.95 ;
      RECT  83.84 82.09 83.64 82.16 ;
      RECT  86.24 81.85 83.84 82.09 ;
      RECT  83.33 81.85 83.12 82.09 ;
      RECT  85.31 81.06 84.77 81.61 ;
      RECT  86.45 82.33 85.31 82.71 ;
      RECT  86.45 81.06 86.24 81.61 ;
      POLYGON  83.47 82.33 83.47 82.4 83.84 82.4 83.84 82.64 83.47 82.64 83.47 82.71 83.33 82.71 83.33 82.33 83.47 82.33 ;
      RECT  83.84 81.85 83.33 82.09 ;
      RECT  84.77 81.06 83.12 81.61 ;
      POLYGON  84.77 82.33 84.77 82.71 84.22 82.71 84.22 82.64 83.84 82.64 83.84 82.4 84.22 82.4 84.22 82.33 84.77 82.33 ;
      RECT  86.45 81.85 86.24 82.09 ;
      RECT  83.84 83.67 83.33 83.43 ;
      RECT  83.84 83.74 83.64 83.67 ;
      RECT  85.31 84.29 84.77 83.91 ;
      RECT  86.24 85.56 85.31 85.01 ;
      RECT  86.45 83.67 86.24 83.43 ;
      RECT  83.33 83.67 83.12 83.43 ;
      RECT  86.24 83.67 83.84 83.43 ;
      RECT  84.05 84.53 83.84 84.46 ;
      RECT  83.33 84.29 83.12 83.91 ;
      RECT  84.05 83.74 83.84 83.67 ;
      RECT  83.84 84.53 83.64 84.46 ;
      RECT  86.24 84.77 83.84 84.53 ;
      RECT  83.33 84.77 83.12 84.53 ;
      RECT  85.31 85.56 84.77 85.01 ;
      RECT  86.45 84.29 85.31 83.91 ;
      RECT  86.45 85.56 86.24 85.01 ;
      POLYGON  83.47 84.29 83.47 84.22 83.84 84.22 83.84 83.98 83.47 83.98 83.47 83.91 83.33 83.91 83.33 84.29 83.47 84.29 ;
      RECT  83.84 84.77 83.33 84.53 ;
      RECT  84.77 85.56 83.12 85.01 ;
      POLYGON  84.77 84.29 84.77 83.91 84.22 83.91 84.22 83.98 83.84 83.98 83.84 84.22 84.22 84.22 84.22 84.29 84.77 84.29 ;
      RECT  86.45 84.77 86.24 84.53 ;
      RECT  83.84 86.9 83.33 87.14 ;
      RECT  83.84 86.83 83.64 86.9 ;
      RECT  85.31 86.28 84.77 86.66 ;
      RECT  86.24 85.01 85.31 85.56 ;
      RECT  86.45 86.9 86.24 87.14 ;
      RECT  83.33 86.9 83.12 87.14 ;
      RECT  86.24 86.9 83.84 87.14 ;
      RECT  84.05 86.04 83.84 86.11 ;
      RECT  83.33 86.28 83.12 86.66 ;
      RECT  84.05 86.83 83.84 86.9 ;
      RECT  83.84 86.04 83.64 86.11 ;
      RECT  86.24 85.8 83.84 86.04 ;
      RECT  83.33 85.8 83.12 86.04 ;
      RECT  85.31 85.01 84.77 85.56 ;
      RECT  86.45 86.28 85.31 86.66 ;
      RECT  86.45 85.01 86.24 85.56 ;
      POLYGON  83.47 86.28 83.47 86.35 83.84 86.35 83.84 86.59 83.47 86.59 83.47 86.66 83.33 86.66 83.33 86.28 83.47 86.28 ;
      RECT  83.84 85.8 83.33 86.04 ;
      RECT  84.77 85.01 83.12 85.56 ;
      POLYGON  84.77 86.28 84.77 86.66 84.22 86.66 84.22 86.59 83.84 86.59 83.84 86.35 84.22 86.35 84.22 86.28 84.77 86.28 ;
      RECT  86.45 85.8 86.24 86.04 ;
      RECT  83.84 87.62 83.33 87.38 ;
      RECT  83.84 87.69 83.64 87.62 ;
      RECT  85.31 88.24 84.77 87.86 ;
      RECT  86.24 89.51 85.31 88.96 ;
      RECT  86.45 87.62 86.24 87.38 ;
      RECT  83.33 87.62 83.12 87.38 ;
      RECT  86.24 87.62 83.84 87.38 ;
      RECT  84.05 88.48 83.84 88.41 ;
      RECT  83.33 88.24 83.12 87.86 ;
      RECT  84.05 87.69 83.84 87.62 ;
      RECT  83.84 88.48 83.64 88.41 ;
      RECT  86.24 88.72 83.84 88.48 ;
      RECT  83.33 88.72 83.12 88.48 ;
      RECT  85.31 89.51 84.77 88.96 ;
      RECT  86.45 88.24 85.31 87.86 ;
      RECT  86.45 89.51 86.24 88.96 ;
      POLYGON  83.47 88.24 83.47 88.17 83.84 88.17 83.84 87.93 83.47 87.93 83.47 87.86 83.33 87.86 83.33 88.24 83.47 88.24 ;
      RECT  83.84 88.72 83.33 88.48 ;
      RECT  84.77 89.51 83.12 88.96 ;
      POLYGON  84.77 88.24 84.77 87.86 84.22 87.86 84.22 87.93 83.84 87.93 83.84 88.17 84.22 88.17 84.22 88.24 84.77 88.24 ;
      RECT  86.45 88.72 86.24 88.48 ;
      RECT  83.84 90.85 83.33 91.09 ;
      RECT  83.84 90.78 83.64 90.85 ;
      RECT  85.31 90.23 84.77 90.61 ;
      RECT  86.24 88.96 85.31 89.51 ;
      RECT  86.45 90.85 86.24 91.09 ;
      RECT  83.33 90.85 83.12 91.09 ;
      RECT  86.24 90.85 83.84 91.09 ;
      RECT  84.05 89.99 83.84 90.06 ;
      RECT  83.33 90.23 83.12 90.61 ;
      RECT  84.05 90.78 83.84 90.85 ;
      RECT  83.84 89.99 83.64 90.06 ;
      RECT  86.24 89.75 83.84 89.99 ;
      RECT  83.33 89.75 83.12 89.99 ;
      RECT  85.31 88.96 84.77 89.51 ;
      RECT  86.45 90.23 85.31 90.61 ;
      RECT  86.45 88.96 86.24 89.51 ;
      POLYGON  83.47 90.23 83.47 90.3 83.84 90.3 83.84 90.54 83.47 90.54 83.47 90.61 83.33 90.61 83.33 90.23 83.47 90.23 ;
      RECT  83.84 89.75 83.33 89.99 ;
      RECT  84.77 88.96 83.12 89.51 ;
      POLYGON  84.77 90.23 84.77 90.61 84.22 90.61 84.22 90.54 83.84 90.54 83.84 90.3 84.22 90.3 84.22 90.23 84.77 90.23 ;
      RECT  86.45 89.75 86.24 89.99 ;
      RECT  83.84 91.57 83.33 91.33 ;
      RECT  83.84 91.64 83.64 91.57 ;
      RECT  85.31 92.19 84.77 91.81 ;
      RECT  86.24 93.46 85.31 92.91 ;
      RECT  86.45 91.57 86.24 91.33 ;
      RECT  83.33 91.57 83.12 91.33 ;
      RECT  86.24 91.57 83.84 91.33 ;
      RECT  84.05 92.43 83.84 92.36 ;
      RECT  83.33 92.19 83.12 91.81 ;
      RECT  84.05 91.64 83.84 91.57 ;
      RECT  83.84 92.43 83.64 92.36 ;
      RECT  86.24 92.67 83.84 92.43 ;
      RECT  83.33 92.67 83.12 92.43 ;
      RECT  85.31 93.46 84.77 92.91 ;
      RECT  86.45 92.19 85.31 91.81 ;
      RECT  86.45 93.46 86.24 92.91 ;
      POLYGON  83.47 92.19 83.47 92.12 83.84 92.12 83.84 91.88 83.47 91.88 83.47 91.81 83.33 91.81 83.33 92.19 83.47 92.19 ;
      RECT  83.84 92.67 83.33 92.43 ;
      RECT  84.77 93.46 83.12 92.91 ;
      POLYGON  84.77 92.19 84.77 91.81 84.22 91.81 84.22 91.88 83.84 91.88 83.84 92.12 84.22 92.12 84.22 92.19 84.77 92.19 ;
      RECT  86.45 92.67 86.24 92.43 ;
      RECT  83.84 94.8 83.33 95.04 ;
      RECT  83.84 94.73 83.64 94.8 ;
      RECT  85.31 94.18 84.77 94.56 ;
      RECT  86.24 92.91 85.31 93.46 ;
      RECT  86.45 94.8 86.24 95.04 ;
      RECT  83.33 94.8 83.12 95.04 ;
      RECT  86.24 94.8 83.84 95.04 ;
      RECT  84.05 93.94 83.84 94.01 ;
      RECT  83.33 94.18 83.12 94.56 ;
      RECT  84.05 94.73 83.84 94.8 ;
      RECT  83.84 93.94 83.64 94.01 ;
      RECT  86.24 93.7 83.84 93.94 ;
      RECT  83.33 93.7 83.12 93.94 ;
      RECT  85.31 92.91 84.77 93.46 ;
      RECT  86.45 94.18 85.31 94.56 ;
      RECT  86.45 92.91 86.24 93.46 ;
      POLYGON  83.47 94.18 83.47 94.25 83.84 94.25 83.84 94.49 83.47 94.49 83.47 94.56 83.33 94.56 83.33 94.18 83.47 94.18 ;
      RECT  83.84 93.7 83.33 93.94 ;
      RECT  84.77 92.91 83.12 93.46 ;
      POLYGON  84.77 94.18 84.77 94.56 84.22 94.56 84.22 94.49 83.84 94.49 83.84 94.25 84.22 94.25 84.22 94.18 84.77 94.18 ;
      RECT  86.45 93.7 86.24 93.94 ;
      RECT  83.12 59.73 86.24 59.97 ;
      RECT  83.12 60.83 86.24 61.07 ;
      RECT  83.12 63.2 86.24 63.44 ;
      RECT  83.12 62.1 86.24 62.34 ;
      RECT  83.12 63.68 86.24 63.92 ;
      RECT  83.12 64.78 86.24 65.02 ;
      RECT  83.12 67.15 86.24 67.39 ;
      RECT  83.12 66.05 86.24 66.29 ;
      RECT  83.12 67.63 86.24 67.87 ;
      RECT  83.12 68.73 86.24 68.97 ;
      RECT  83.12 71.1 86.24 71.34 ;
      RECT  83.12 70.0 86.24 70.24 ;
      RECT  83.12 71.58 86.24 71.82 ;
      RECT  83.12 72.68 86.24 72.92 ;
      RECT  83.12 75.05 86.24 75.29 ;
      RECT  83.12 73.95 86.24 74.19 ;
      RECT  83.12 75.53 86.24 75.77 ;
      RECT  83.12 76.63 86.24 76.87 ;
      RECT  83.12 79.0 86.24 79.24 ;
      RECT  83.12 77.9 86.24 78.14 ;
      RECT  83.12 79.48 86.24 79.72 ;
      RECT  83.12 80.58 86.24 80.82 ;
      RECT  83.12 82.95 86.24 83.19 ;
      RECT  83.12 81.85 86.24 82.09 ;
      RECT  83.12 83.43 86.24 83.67 ;
      RECT  83.12 84.53 86.24 84.77 ;
      RECT  83.12 86.9 86.24 87.14 ;
      RECT  83.12 85.8 86.24 86.04 ;
      RECT  83.12 87.38 86.24 87.62 ;
      RECT  83.12 88.48 86.24 88.72 ;
      RECT  83.12 90.85 86.24 91.09 ;
      RECT  83.12 89.75 86.24 89.99 ;
      RECT  83.12 91.33 86.24 91.57 ;
      RECT  83.12 92.43 86.24 92.67 ;
      RECT  83.12 94.8 86.24 95.04 ;
      RECT  83.12 93.7 86.24 93.94 ;
      RECT  67.52 63.2 86.24 63.44 ;
      RECT  67.52 62.1 86.24 62.34 ;
      RECT  67.52 63.68 86.24 63.92 ;
      RECT  67.52 64.78 86.24 65.02 ;
      RECT  67.52 67.15 86.24 67.39 ;
      RECT  67.52 66.05 86.24 66.29 ;
      RECT  67.52 67.63 86.24 67.87 ;
      RECT  67.52 68.73 86.24 68.97 ;
      RECT  67.52 71.1 86.24 71.34 ;
      RECT  67.52 70.0 86.24 70.24 ;
      RECT  67.52 71.58 86.24 71.82 ;
      RECT  67.52 72.68 86.24 72.92 ;
      RECT  67.52 75.05 86.24 75.29 ;
      RECT  67.52 73.95 86.24 74.19 ;
      RECT  67.52 75.53 86.24 75.77 ;
      RECT  67.52 76.63 86.24 76.87 ;
      RECT  67.52 79.0 86.24 79.24 ;
      RECT  67.52 77.9 86.24 78.14 ;
      RECT  67.52 79.48 86.24 79.72 ;
      RECT  67.52 80.58 86.24 80.82 ;
      RECT  67.52 82.95 86.24 83.19 ;
      RECT  67.52 81.85 86.24 82.09 ;
      RECT  67.52 83.43 86.24 83.67 ;
      RECT  67.52 84.53 86.24 84.77 ;
      RECT  67.52 86.9 86.24 87.14 ;
      RECT  67.52 85.8 86.24 86.04 ;
      RECT  67.52 87.38 86.24 87.62 ;
      RECT  67.52 88.48 86.24 88.72 ;
      RECT  67.52 90.85 86.24 91.09 ;
      RECT  67.52 89.75 86.24 89.99 ;
      RECT  67.52 91.33 86.24 91.57 ;
      RECT  67.52 92.43 86.24 92.67 ;
      RECT  67.52 59.73 86.24 59.97 ;
      RECT  67.52 93.7 86.24 93.94 ;
      RECT  72.29 83.91 72.83 84.29 ;
      RECT  72.29 81.06 72.83 81.61 ;
      RECT  80.93 69.21 81.47 69.76 ;
      RECT  80.93 66.53 81.47 66.91 ;
      RECT  72.29 61.31 72.83 61.86 ;
      RECT  72.29 62.58 72.83 62.96 ;
      RECT  72.29 76.01 72.83 76.39 ;
      RECT  72.29 87.86 72.83 88.24 ;
      RECT  80.93 91.81 81.47 92.19 ;
      RECT  72.29 94.18 72.83 94.56 ;
      RECT  72.29 77.11 72.83 77.66 ;
      RECT  80.93 62.58 81.47 62.96 ;
      RECT  80.93 86.28 81.47 86.66 ;
      RECT  80.93 94.18 81.47 94.56 ;
      RECT  72.29 78.38 72.83 78.76 ;
      RECT  72.29 69.21 72.83 69.76 ;
      RECT  72.29 64.16 72.83 64.54 ;
      RECT  80.93 60.21 81.47 60.59 ;
      RECT  80.93 74.43 81.47 74.81 ;
      RECT  72.29 73.16 72.83 73.71 ;
      RECT  72.29 88.96 72.83 89.51 ;
      RECT  72.29 65.26 72.83 65.81 ;
      RECT  72.29 70.48 72.83 70.86 ;
      RECT  80.93 73.16 81.47 73.71 ;
      RECT  80.93 87.86 81.47 88.24 ;
      RECT  72.29 90.23 72.83 90.61 ;
      RECT  80.93 81.06 81.47 81.61 ;
      RECT  80.93 70.48 81.47 70.86 ;
      RECT  80.93 72.06 81.47 72.44 ;
      RECT  80.93 88.96 81.47 89.51 ;
      RECT  80.93 64.16 81.47 64.54 ;
      RECT  80.93 79.96 81.47 80.34 ;
      RECT  72.29 74.43 72.83 74.81 ;
      RECT  72.29 85.01 72.83 85.56 ;
      RECT  72.29 82.33 72.83 82.71 ;
      RECT  80.93 68.11 81.47 68.49 ;
      RECT  72.29 79.96 72.83 80.34 ;
      RECT  80.93 92.91 81.47 93.46 ;
      RECT  80.93 78.38 81.47 78.76 ;
      RECT  72.29 92.91 72.83 93.46 ;
      RECT  72.29 91.81 72.83 92.19 ;
      RECT  80.93 83.91 81.47 84.29 ;
      RECT  72.29 86.28 72.83 86.66 ;
      RECT  80.93 61.31 81.47 61.86 ;
      RECT  72.29 72.06 72.83 72.44 ;
      RECT  72.29 60.21 72.83 60.59 ;
      RECT  80.93 85.01 81.47 85.56 ;
      RECT  72.29 68.11 72.83 68.49 ;
      RECT  72.29 66.53 72.83 66.91 ;
      RECT  80.93 65.26 81.47 65.81 ;
      RECT  80.93 77.11 81.47 77.66 ;
      RECT  80.93 90.23 81.47 90.61 ;
      RECT  80.93 82.33 81.47 82.71 ;
      RECT  80.93 76.01 81.47 76.39 ;
      RECT  73.76 52.66 70.64 52.8 ;
      RECT  73.76 52.66 76.88 52.8 ;
      RECT  80.0 52.66 76.88 52.8 ;
      RECT  73.76 102.11 76.88 101.97 ;
      RECT  80.0 102.11 76.88 101.97 ;
      RECT  80.0 102.11 83.12 101.97 ;
      RECT  56.7 61.585 56.84 93.185 ;
      RECT  56.7 61.585 56.84 93.185 ;
      RECT  97.06 61.585 96.92 93.185 ;
      RECT  97.06 61.585 96.92 93.185 ;
      RECT  64.42 28.75 64.56 60.785 ;
      RECT  88.1 93.985 88.24 115.125 ;
      RECT  65.66 28.75 65.8 60.785 ;
      RECT  87.48 93.985 87.62 115.125 ;
      RECT  65.04 28.75 65.18 60.785 ;
      RECT  66.28 28.75 66.42 60.785 ;
      RECT  86.86 93.985 87.0 115.125 ;
      RECT  6.09 3.32 6.42 3.58 ;
      RECT  1.365 2.965 1.695 3.225 ;
      RECT  5.7 2.565 6.03 2.825 ;
      RECT  2.525 3.735 2.795 4.055 ;
      RECT  1.365 2.965 1.695 3.225 ;
      RECT  11.05 2.72 11.19 2.86 ;
      RECT  8.52 4.63 8.66 4.77 ;
      RECT  2.525 3.735 2.795 4.055 ;
      RECT  6.09 11.37 6.42 11.11 ;
      RECT  1.365 11.725 1.695 11.465 ;
      RECT  5.7 12.125 6.03 11.865 ;
      RECT  2.525 10.955 2.795 10.635 ;
      RECT  1.365 11.725 1.695 11.465 ;
      RECT  11.05 11.97 11.19 11.83 ;
      RECT  8.52 10.06 8.66 9.92 ;
      RECT  2.525 10.955 2.795 10.635 ;
      RECT  1.365 2.965 1.695 3.225 ;
      RECT  1.365 11.465 1.695 11.725 ;
      RECT  11.05 2.72 11.19 2.86 ;
      RECT  8.52 4.63 8.66 4.77 ;
      RECT  11.05 11.83 11.19 11.97 ;
      RECT  8.52 9.92 8.66 10.06 ;
      RECT  2.525 0.275 2.665 14.415 ;
      RECT  9.56 57.635 9.42 60.245 ;
      RECT  1.765 57.635 1.625 105.045 ;
      RECT  1.365 2.965 1.695 3.225 ;
      RECT  1.365 11.465 1.695 11.725 ;
      RECT  16.115 3.55 16.255 3.69 ;
      RECT  9.42 57.635 9.56 60.245 ;
      RECT  19.17 53.36 27.91 53.5 ;
      RECT  20.25 32.02 27.91 32.16 ;
      RECT  20.94 39.28 27.91 39.42 ;
      RECT  22.27 24.95 27.91 25.09 ;
      RECT  25.0 3.74 27.91 3.88 ;
      RECT  146.56 137.31 146.23 137.05 ;
      RECT  151.285 137.665 150.955 137.405 ;
      RECT  146.95 138.065 146.62 137.805 ;
      RECT  150.125 136.895 149.855 136.575 ;
      RECT  151.285 137.665 150.955 137.405 ;
      RECT  141.6 137.91 141.46 137.77 ;
      RECT  144.13 136.0 143.99 135.86 ;
      RECT  150.125 136.895 149.855 136.575 ;
      RECT  151.285 137.665 150.955 137.405 ;
      RECT  141.6 137.91 141.46 137.77 ;
      RECT  144.13 136.0 143.99 135.86 ;
      RECT  150.125 140.355 149.985 133.285 ;
      RECT  143.09 97.135 143.23 94.525 ;
      RECT  150.885 97.135 151.025 49.725 ;
      RECT  151.285 137.665 150.955 137.405 ;
      RECT  136.955 137.08 136.815 136.94 ;
      RECT  143.23 97.135 143.09 94.525 ;
      RECT  133.9 101.41 126.27 101.27 ;
      RECT  132.13 108.8 126.27 108.66 ;
      RECT  130.8 115.68 126.27 115.54 ;
      RECT  129.14 136.97 126.27 136.83 ;
      RECT  27.48 111.88 27.81 112.14 ;
      RECT  22.755 111.525 23.085 111.785 ;
      RECT  27.09 111.125 27.42 111.385 ;
      RECT  23.915 112.295 24.185 112.615 ;
      RECT  27.48 119.93 27.81 119.67 ;
      RECT  22.755 120.285 23.085 120.025 ;
      RECT  27.09 120.685 27.42 120.425 ;
      RECT  23.915 119.515 24.185 119.195 ;
      RECT  27.48 126.02 27.81 126.28 ;
      RECT  22.755 125.665 23.085 125.925 ;
      RECT  27.09 125.265 27.42 125.525 ;
      RECT  23.915 126.435 24.185 126.755 ;
      RECT  27.48 134.07 27.81 133.81 ;
      RECT  22.755 134.425 23.085 134.165 ;
      RECT  27.09 134.825 27.42 134.565 ;
      RECT  23.915 133.655 24.185 133.335 ;
      RECT  22.755 111.525 23.085 111.785 ;
      RECT  22.755 120.025 23.085 120.285 ;
      RECT  22.755 125.665 23.085 125.925 ;
      RECT  22.755 134.165 23.085 134.425 ;
      RECT  27.48 111.88 27.81 112.14 ;
      RECT  27.48 119.67 27.81 119.93 ;
      RECT  27.48 126.02 27.81 126.28 ;
      RECT  27.48 133.81 27.81 134.07 ;
      RECT  126.7 42.89 126.37 42.63 ;
      RECT  131.425 43.245 131.095 42.985 ;
      RECT  127.09 43.645 126.76 43.385 ;
      RECT  130.265 42.475 129.995 42.155 ;
      RECT  126.7 34.84 126.37 35.1 ;
      RECT  131.425 34.485 131.095 34.745 ;
      RECT  127.09 34.085 126.76 34.345 ;
      RECT  130.265 35.255 129.995 35.575 ;
      RECT  126.7 28.75 126.37 28.49 ;
      RECT  131.425 29.105 131.095 28.845 ;
      RECT  127.09 29.505 126.76 29.245 ;
      RECT  130.265 28.335 129.995 28.015 ;
      RECT  126.7 20.7 126.37 20.96 ;
      RECT  131.425 20.345 131.095 20.605 ;
      RECT  127.09 19.945 126.76 20.205 ;
      RECT  130.265 21.115 129.995 21.435 ;
      RECT  131.425 43.245 131.095 42.985 ;
      RECT  131.425 34.745 131.095 34.485 ;
      RECT  131.425 29.105 131.095 28.845 ;
      RECT  131.425 20.605 131.095 20.345 ;
      RECT  126.7 42.89 126.37 42.63 ;
      RECT  126.7 35.1 126.37 34.84 ;
      RECT  126.7 28.75 126.37 28.49 ;
      RECT  126.7 20.96 126.37 20.7 ;
      RECT  39.16 16.185 39.49 16.445 ;
      RECT  34.435 15.83 34.765 16.09 ;
      RECT  38.77 15.43 39.1 15.69 ;
      RECT  35.595 16.6 35.865 16.92 ;
      RECT  45.0 16.185 45.33 16.445 ;
      RECT  40.275 15.83 40.605 16.09 ;
      RECT  44.61 15.43 44.94 15.69 ;
      RECT  41.435 16.6 41.705 16.92 ;
      RECT  34.435 15.83 34.765 16.09 ;
      RECT  40.275 15.83 40.605 16.09 ;
      RECT  39.16 16.185 39.49 16.445 ;
      RECT  45.0 16.185 45.33 16.445 ;
   LAYER  m3 ;
      RECT  71.955 95.745 72.445 96.235 ;
      RECT  71.955 58.535 72.445 59.025 ;
      RECT  81.315 95.745 81.805 96.235 ;
      RECT  81.315 58.535 81.805 59.025 ;
      RECT  75.075 58.535 75.565 59.025 ;
      RECT  78.195 58.535 78.685 59.025 ;
      RECT  75.075 96.235 75.565 95.745 ;
      RECT  78.195 96.235 78.685 95.745 ;
      RECT  68.475 74.375 68.965 74.865 ;
      RECT  68.475 73.19 68.965 73.68 ;
      RECT  68.475 81.09 68.965 81.58 ;
      RECT  68.475 85.04 68.965 85.53 ;
      RECT  68.475 70.425 68.965 70.915 ;
      RECT  68.475 88.99 68.965 89.48 ;
      RECT  68.475 75.955 68.965 76.445 ;
      RECT  68.475 78.325 68.965 78.815 ;
      RECT  68.475 61.34 68.965 61.83 ;
      RECT  68.475 91.755 68.965 92.245 ;
      RECT  68.475 79.905 68.965 80.395 ;
      RECT  68.475 94.125 68.965 94.615 ;
      RECT  68.475 87.805 68.965 88.295 ;
      RECT  68.475 66.475 68.965 66.965 ;
      RECT  68.475 62.525 68.965 63.015 ;
      RECT  68.475 65.29 68.965 65.78 ;
      RECT  68.475 90.175 68.965 90.665 ;
      RECT  68.475 82.275 68.965 82.765 ;
      RECT  68.475 83.855 68.965 84.345 ;
      RECT  68.475 86.225 68.965 86.715 ;
      RECT  68.475 64.105 68.965 64.595 ;
      RECT  68.475 72.005 68.965 72.495 ;
      RECT  68.475 68.055 68.965 68.545 ;
      RECT  68.475 92.94 68.965 93.43 ;
      RECT  68.475 69.24 68.965 69.73 ;
      RECT  68.475 77.14 68.965 77.63 ;
      RECT  68.475 60.155 68.965 60.645 ;
      RECT  84.795 94.125 85.285 94.615 ;
      RECT  84.795 73.19 85.285 73.68 ;
      RECT  84.795 86.225 85.285 86.715 ;
      RECT  84.795 69.24 85.285 69.73 ;
      RECT  84.795 75.955 85.285 76.445 ;
      RECT  84.795 62.525 85.285 63.015 ;
      RECT  84.795 64.105 85.285 64.595 ;
      RECT  84.795 87.805 85.285 88.295 ;
      RECT  84.795 60.155 85.285 60.645 ;
      RECT  84.795 72.005 85.285 72.495 ;
      RECT  84.795 88.99 85.285 89.48 ;
      RECT  84.795 78.325 85.285 78.815 ;
      RECT  84.795 66.475 85.285 66.965 ;
      RECT  84.795 83.855 85.285 84.345 ;
      RECT  84.795 90.175 85.285 90.665 ;
      RECT  84.795 81.09 85.285 81.58 ;
      RECT  84.795 70.425 85.285 70.915 ;
      RECT  84.795 82.275 85.285 82.765 ;
      RECT  84.795 68.055 85.285 68.545 ;
      RECT  84.795 65.29 85.285 65.78 ;
      RECT  84.795 74.375 85.285 74.865 ;
      RECT  84.795 92.94 85.285 93.43 ;
      RECT  84.795 91.755 85.285 92.245 ;
      RECT  84.795 61.34 85.285 61.83 ;
      RECT  84.795 79.905 85.285 80.395 ;
      RECT  84.795 85.04 85.285 85.53 ;
      RECT  84.795 77.14 85.285 77.63 ;
      RECT  81.315 58.535 81.805 59.025 ;
      RECT  75.17 58.63 75.47 58.93 ;
      RECT  71.955 58.535 72.445 59.025 ;
      RECT  71.955 95.745 72.445 96.235 ;
      RECT  78.29 58.63 78.59 58.93 ;
      RECT  78.29 95.84 78.59 96.14 ;
      RECT  75.17 95.84 75.47 96.14 ;
      RECT  81.315 95.745 81.805 96.235 ;
      RECT  68.57 65.385 68.87 65.685 ;
      RECT  84.89 66.57 85.19 66.87 ;
      RECT  68.57 68.15 68.87 68.45 ;
      RECT  68.57 64.2 68.87 64.5 ;
      RECT  84.89 86.32 85.19 86.62 ;
      RECT  68.57 85.135 68.87 85.435 ;
      RECT  84.89 64.2 85.19 64.5 ;
      RECT  84.89 91.85 85.19 92.15 ;
      RECT  68.57 78.42 68.87 78.72 ;
      RECT  84.89 89.085 85.19 89.385 ;
      RECT  84.89 77.235 85.19 77.535 ;
      RECT  68.57 90.27 68.87 90.57 ;
      RECT  84.89 73.285 85.19 73.585 ;
      RECT  68.57 70.52 68.87 70.82 ;
      RECT  84.89 61.435 85.19 61.735 ;
      RECT  68.57 69.335 68.87 69.635 ;
      RECT  84.89 65.385 85.19 65.685 ;
      RECT  84.89 90.27 85.19 90.57 ;
      RECT  84.89 68.15 85.19 68.45 ;
      RECT  68.57 77.235 68.87 77.535 ;
      RECT  84.89 94.22 85.19 94.52 ;
      RECT  68.57 89.085 68.87 89.385 ;
      RECT  68.57 82.37 68.87 82.67 ;
      RECT  68.57 81.185 68.87 81.485 ;
      RECT  84.89 82.37 85.19 82.67 ;
      RECT  84.89 72.1 85.19 72.4 ;
      RECT  84.89 69.335 85.19 69.635 ;
      RECT  68.57 60.25 68.87 60.55 ;
      RECT  84.89 74.47 85.19 74.77 ;
      RECT  84.89 62.62 85.19 62.92 ;
      RECT  84.89 78.42 85.19 78.72 ;
      RECT  84.89 60.25 85.19 60.55 ;
      RECT  84.89 83.95 85.19 84.25 ;
      RECT  84.89 87.9 85.19 88.2 ;
      RECT  68.57 94.22 68.87 94.52 ;
      RECT  84.89 76.05 85.19 76.35 ;
      RECT  68.57 86.32 68.87 86.62 ;
      RECT  68.57 83.95 68.87 84.25 ;
      RECT  68.57 87.9 68.87 88.2 ;
      RECT  68.57 66.57 68.87 66.87 ;
      RECT  68.57 76.05 68.87 76.35 ;
      RECT  84.89 93.035 85.19 93.335 ;
      RECT  68.57 73.285 68.87 73.585 ;
      RECT  68.57 61.435 68.87 61.735 ;
      RECT  68.57 74.47 68.87 74.77 ;
      RECT  84.89 81.185 85.19 81.485 ;
      RECT  84.89 85.135 85.19 85.435 ;
      RECT  68.57 93.035 68.87 93.335 ;
      RECT  68.57 62.62 68.87 62.92 ;
      RECT  68.57 72.1 68.87 72.4 ;
      RECT  68.57 80.0 68.87 80.3 ;
      RECT  84.89 80.0 85.19 80.3 ;
      RECT  68.57 91.85 68.87 92.15 ;
      RECT  84.89 70.52 85.19 70.82 ;
      RECT  73.04 55.58 72.55 56.07 ;
      RECT  74.48 55.58 74.97 56.07 ;
      RECT  79.28 55.58 78.79 56.07 ;
      RECT  70.64 52.58 80.0 52.88 ;
      RECT  72.55 55.58 73.04 56.07 ;
      RECT  78.79 55.58 79.28 56.07 ;
      RECT  74.48 55.58 74.97 56.07 ;
      RECT  73.76 50.885 80.0 51.185 ;
      RECT  77.29 46.16 77.78 46.65 ;
      RECT  77.23 41.97 77.72 42.46 ;
      RECT  75.36 46.16 75.85 46.65 ;
      RECT  75.42 41.97 75.91 42.46 ;
      RECT  76.88 50.03 77.37 50.52 ;
      RECT  75.42 40.36 75.91 40.85 ;
      RECT  77.23 40.36 77.72 40.85 ;
      RECT  75.77 50.03 76.26 50.52 ;
      RECT  74.795 34.21 75.285 34.7 ;
      RECT  77.755 29.46 78.245 29.95 ;
      RECT  74.895 29.46 75.385 29.95 ;
      RECT  77.855 34.21 78.345 34.7 ;
      RECT  74.85 36.395 75.34 36.885 ;
      RECT  75.4 32.55 75.89 33.04 ;
      RECT  77.825 31.54 78.315 32.03 ;
      RECT  77.8 36.395 78.29 36.885 ;
      RECT  74.825 31.54 75.315 32.03 ;
      RECT  77.25 32.55 77.74 33.04 ;
      RECT  73.76 51.185 80.0 50.885 ;
      RECT  70.64 52.88 80.0 52.58 ;
      RECT  74.895 29.95 75.385 29.46 ;
      RECT  72.55 56.07 73.04 55.58 ;
      RECT  77.855 34.7 78.345 34.21 ;
      RECT  75.42 42.46 75.91 41.97 ;
      RECT  77.29 46.65 77.78 46.16 ;
      RECT  74.48 56.07 74.97 55.58 ;
      RECT  75.36 46.65 75.85 46.16 ;
      RECT  74.795 34.7 75.285 34.21 ;
      RECT  78.79 56.07 79.28 55.58 ;
      RECT  77.755 29.95 78.245 29.46 ;
      RECT  77.23 42.46 77.72 41.97 ;
      RECT  74.85 36.885 75.34 36.395 ;
      RECT  77.8 36.885 78.29 36.395 ;
      RECT  75.42 40.85 75.91 40.36 ;
      RECT  77.25 33.04 77.74 32.55 ;
      RECT  75.4 33.04 75.89 32.55 ;
      RECT  75.77 50.52 76.26 50.03 ;
      RECT  77.825 32.03 78.315 31.54 ;
      RECT  77.23 40.85 77.72 40.36 ;
      RECT  74.825 32.03 75.315 31.54 ;
      RECT  76.88 50.52 77.37 50.03 ;
      RECT  74.48 99.19 74.97 98.7 ;
      RECT  79.28 99.19 78.79 98.7 ;
      RECT  80.72 99.19 81.21 98.7 ;
      RECT  73.76 102.19 83.12 101.89 ;
      RECT  80.72 99.19 81.21 98.7 ;
      RECT  78.79 99.19 79.28 98.7 ;
      RECT  74.48 99.19 74.97 98.7 ;
      RECT  73.76 103.885 80.0 103.585 ;
      RECT  77.29 108.61 77.78 108.12 ;
      RECT  77.23 112.8 77.72 112.31 ;
      RECT  75.36 108.61 75.85 108.12 ;
      RECT  75.42 112.8 75.91 112.31 ;
      RECT  76.88 104.74 77.37 104.25 ;
      RECT  75.42 114.41 75.91 113.92 ;
      RECT  77.23 114.41 77.72 113.92 ;
      RECT  75.77 104.74 76.26 104.25 ;
      RECT  73.76 103.585 80.0 103.885 ;
      RECT  73.76 101.89 83.12 102.19 ;
      RECT  77.29 108.12 77.78 108.61 ;
      RECT  74.48 98.7 74.97 99.19 ;
      RECT  77.23 112.31 77.72 112.8 ;
      RECT  75.36 108.12 75.85 108.61 ;
      RECT  78.79 98.7 79.28 99.19 ;
      RECT  80.72 98.7 81.21 99.19 ;
      RECT  75.42 112.31 75.91 112.8 ;
      RECT  75.77 104.25 76.26 104.74 ;
      RECT  76.88 104.25 77.37 104.74 ;
      RECT  75.42 113.92 75.91 114.41 ;
      RECT  77.23 113.92 77.72 114.41 ;
      RECT  40.9 63.495 41.39 63.985 ;
      RECT  34.285 63.46 34.775 63.95 ;
      RECT  44.155 63.46 44.645 63.95 ;
      RECT  44.155 67.41 44.645 67.9 ;
      RECT  40.9 67.445 41.39 67.935 ;
      RECT  42.795 67.41 43.285 67.9 ;
      RECT  38.775 67.445 39.265 67.935 ;
      RECT  32.925 63.46 33.415 63.95 ;
      RECT  42.795 63.46 43.285 63.95 ;
      RECT  38.775 63.495 39.265 63.985 ;
      RECT  40.9 75.345 41.39 75.835 ;
      RECT  34.285 75.31 34.775 75.8 ;
      RECT  44.155 75.31 44.645 75.8 ;
      RECT  44.155 79.26 44.645 79.75 ;
      RECT  40.9 79.295 41.39 79.785 ;
      RECT  42.795 79.26 43.285 79.75 ;
      RECT  38.775 79.295 39.265 79.785 ;
      RECT  32.925 75.31 33.415 75.8 ;
      RECT  42.795 75.31 43.285 75.8 ;
      RECT  38.775 75.345 39.265 75.835 ;
      RECT  51.97 69.545 52.46 70.035 ;
      RECT  44.155 63.46 44.645 63.95 ;
      RECT  51.97 71.395 52.46 71.885 ;
      RECT  55.225 65.435 55.715 65.925 ;
      RECT  55.225 81.235 55.715 81.725 ;
      RECT  55.225 87.16 55.715 87.65 ;
      RECT  55.225 75.31 55.715 75.8 ;
      RECT  44.155 67.41 44.645 67.9 ;
      RECT  34.285 75.31 34.775 75.8 ;
      RECT  55.225 77.285 55.715 77.775 ;
      RECT  55.225 73.335 55.715 73.825 ;
      RECT  44.155 75.31 44.645 75.8 ;
      RECT  51.97 67.445 52.46 67.935 ;
      RECT  51.97 79.295 52.46 79.785 ;
      RECT  51.97 89.295 52.46 89.785 ;
      RECT  55.225 83.21 55.715 83.7 ;
      RECT  55.225 69.385 55.715 69.875 ;
      RECT  51.97 81.395 52.46 81.885 ;
      RECT  51.97 75.345 52.46 75.835 ;
      RECT  55.225 63.46 55.715 63.95 ;
      RECT  55.225 91.11 55.715 91.6 ;
      RECT  51.97 63.495 52.46 63.985 ;
      RECT  40.9 63.495 41.39 63.985 ;
      RECT  40.9 67.445 41.39 67.935 ;
      RECT  40.9 79.295 41.39 79.785 ;
      RECT  51.97 83.245 52.46 83.735 ;
      RECT  51.97 73.495 52.46 73.985 ;
      RECT  55.225 85.185 55.715 85.675 ;
      RECT  55.225 71.36 55.715 71.85 ;
      RECT  44.155 79.26 44.645 79.75 ;
      RECT  34.285 63.46 34.775 63.95 ;
      RECT  51.97 87.195 52.46 87.685 ;
      RECT  51.97 85.345 52.46 85.835 ;
      RECT  55.225 79.26 55.715 79.75 ;
      RECT  55.225 89.135 55.715 89.625 ;
      RECT  51.97 91.145 52.46 91.635 ;
      RECT  40.9 75.345 41.39 75.835 ;
      RECT  51.97 77.445 52.46 77.935 ;
      RECT  51.97 65.595 52.46 66.085 ;
      RECT  55.225 67.41 55.715 67.9 ;
      RECT  49.845 73.485 50.335 73.975 ;
      RECT  49.845 89.285 50.335 89.775 ;
      RECT  38.775 75.345 39.265 75.835 ;
      RECT  49.845 81.385 50.335 81.875 ;
      RECT  53.865 73.335 54.355 73.825 ;
      RECT  49.845 69.535 50.335 70.025 ;
      RECT  42.795 75.31 43.285 75.8 ;
      RECT  53.865 71.36 54.355 71.85 ;
      RECT  53.865 77.285 54.355 77.775 ;
      RECT  53.865 89.135 54.355 89.625 ;
      RECT  38.775 79.295 39.265 79.785 ;
      RECT  42.795 63.46 43.285 63.95 ;
      RECT  49.845 67.445 50.335 67.935 ;
      RECT  49.845 79.295 50.335 79.785 ;
      RECT  53.865 81.235 54.355 81.725 ;
      RECT  53.865 85.185 54.355 85.675 ;
      RECT  53.865 91.11 54.355 91.6 ;
      RECT  42.795 67.41 43.285 67.9 ;
      RECT  53.865 79.26 54.355 79.75 ;
      RECT  49.845 85.335 50.335 85.825 ;
      RECT  32.925 63.46 33.415 63.95 ;
      RECT  49.845 87.195 50.335 87.685 ;
      RECT  42.795 79.26 43.285 79.75 ;
      RECT  53.865 75.31 54.355 75.8 ;
      RECT  49.845 77.435 50.335 77.925 ;
      RECT  53.865 69.385 54.355 69.875 ;
      RECT  53.865 83.21 54.355 83.7 ;
      RECT  38.775 67.445 39.265 67.935 ;
      RECT  38.775 63.495 39.265 63.985 ;
      RECT  49.845 71.395 50.335 71.885 ;
      RECT  49.845 75.345 50.335 75.835 ;
      RECT  49.845 63.495 50.335 63.985 ;
      RECT  53.865 65.435 54.355 65.925 ;
      RECT  49.845 83.245 50.335 83.735 ;
      RECT  53.865 87.16 54.355 87.65 ;
      RECT  49.845 91.145 50.335 91.635 ;
      RECT  49.845 65.585 50.335 66.075 ;
      RECT  53.865 63.46 54.355 63.95 ;
      RECT  53.865 67.41 54.355 67.9 ;
      RECT  32.925 75.31 33.415 75.8 ;
      RECT  55.225 71.36 55.715 71.85 ;
      RECT  40.9 63.495 41.39 63.985 ;
      RECT  40.9 75.345 41.39 75.835 ;
      RECT  51.97 91.145 52.46 91.635 ;
      RECT  51.97 77.445 52.46 77.935 ;
      RECT  40.9 67.445 41.39 67.935 ;
      RECT  51.97 87.195 52.46 87.685 ;
      RECT  51.97 89.295 52.46 89.785 ;
      RECT  55.225 83.21 55.715 83.7 ;
      RECT  51.97 81.395 52.46 81.885 ;
      RECT  51.97 67.445 52.46 67.935 ;
      RECT  55.225 79.26 55.715 79.75 ;
      RECT  44.155 67.41 44.645 67.9 ;
      RECT  51.97 75.345 52.46 75.835 ;
      RECT  55.225 63.46 55.715 63.95 ;
      RECT  51.97 79.295 52.46 79.785 ;
      RECT  51.97 83.245 52.46 83.735 ;
      RECT  55.225 81.235 55.715 81.725 ;
      RECT  51.97 73.495 52.46 73.985 ;
      RECT  55.225 87.16 55.715 87.65 ;
      RECT  51.97 65.595 52.46 66.085 ;
      RECT  44.155 75.31 44.645 75.8 ;
      RECT  64.155 77.14 64.645 77.63 ;
      RECT  55.225 67.41 55.715 67.9 ;
      RECT  51.97 85.345 52.46 85.835 ;
      RECT  34.285 63.46 34.775 63.95 ;
      RECT  55.225 65.435 55.715 65.925 ;
      RECT  51.97 63.495 52.46 63.985 ;
      RECT  55.225 89.135 55.715 89.625 ;
      RECT  55.225 75.31 55.715 75.8 ;
      RECT  44.155 79.26 44.645 79.75 ;
      RECT  34.285 75.31 34.775 75.8 ;
      RECT  59.58 77.06 60.07 77.55 ;
      RECT  55.225 69.385 55.715 69.875 ;
      RECT  44.155 63.46 44.645 63.95 ;
      RECT  55.225 77.285 55.715 77.775 ;
      RECT  55.225 85.185 55.715 85.675 ;
      RECT  51.97 69.545 52.46 70.035 ;
      RECT  40.9 79.295 41.39 79.785 ;
      RECT  55.225 91.11 55.715 91.6 ;
      RECT  51.97 71.395 52.46 71.885 ;
      RECT  55.225 73.335 55.715 73.825 ;
      RECT  49.845 91.145 50.335 91.635 ;
      RECT  49.845 87.195 50.335 87.685 ;
      RECT  53.865 81.235 54.355 81.725 ;
      RECT  53.865 91.11 54.355 91.6 ;
      RECT  49.845 89.285 50.335 89.775 ;
      RECT  49.845 63.495 50.335 63.985 ;
      RECT  49.845 67.445 50.335 67.935 ;
      RECT  49.845 79.295 50.335 79.785 ;
      RECT  49.845 69.535 50.335 70.025 ;
      RECT  53.865 67.41 54.355 67.9 ;
      RECT  57.455 77.065 57.945 77.555 ;
      RECT  53.865 79.26 54.355 79.75 ;
      RECT  42.795 67.41 43.285 67.9 ;
      RECT  49.845 75.345 50.335 75.835 ;
      RECT  49.845 83.245 50.335 83.735 ;
      RECT  49.845 71.395 50.335 71.885 ;
      RECT  42.795 79.26 43.285 79.75 ;
      RECT  38.775 63.495 39.265 63.985 ;
      RECT  53.865 85.185 54.355 85.675 ;
      RECT  53.865 83.21 54.355 83.7 ;
      RECT  49.845 85.335 50.335 85.825 ;
      RECT  49.845 73.485 50.335 73.975 ;
      RECT  53.865 65.435 54.355 65.925 ;
      RECT  42.795 75.31 43.285 75.8 ;
      RECT  49.845 65.585 50.335 66.075 ;
      RECT  53.865 71.36 54.355 71.85 ;
      RECT  32.925 63.46 33.415 63.95 ;
      RECT  42.795 63.46 43.285 63.95 ;
      RECT  49.845 81.385 50.335 81.875 ;
      RECT  53.865 77.285 54.355 77.775 ;
      RECT  53.865 73.335 54.355 73.825 ;
      RECT  61.665 77.14 62.155 77.63 ;
      RECT  38.775 67.445 39.265 67.935 ;
      RECT  53.865 87.16 54.355 87.65 ;
      RECT  38.775 79.295 39.265 79.785 ;
      RECT  53.865 69.385 54.355 69.875 ;
      RECT  38.775 75.345 39.265 75.835 ;
      RECT  49.845 77.435 50.335 77.925 ;
      RECT  53.865 75.31 54.355 75.8 ;
      RECT  53.865 89.135 54.355 89.625 ;
      RECT  32.925 75.31 33.415 75.8 ;
      RECT  53.865 63.46 54.355 63.95 ;
      RECT  112.86 63.495 112.37 63.985 ;
      RECT  119.475 63.46 118.985 63.95 ;
      RECT  109.605 63.46 109.115 63.95 ;
      RECT  109.605 67.41 109.115 67.9 ;
      RECT  112.86 67.445 112.37 67.935 ;
      RECT  110.965 67.41 110.475 67.9 ;
      RECT  114.985 67.445 114.495 67.935 ;
      RECT  120.835 63.46 120.345 63.95 ;
      RECT  110.965 63.46 110.475 63.95 ;
      RECT  114.985 63.495 114.495 63.985 ;
      RECT  112.86 75.345 112.37 75.835 ;
      RECT  119.475 75.31 118.985 75.8 ;
      RECT  109.605 75.31 109.115 75.8 ;
      RECT  109.605 79.26 109.115 79.75 ;
      RECT  112.86 79.295 112.37 79.785 ;
      RECT  110.965 79.26 110.475 79.75 ;
      RECT  114.985 79.295 114.495 79.785 ;
      RECT  120.835 75.31 120.345 75.8 ;
      RECT  110.965 75.31 110.475 75.8 ;
      RECT  114.985 75.345 114.495 75.835 ;
      RECT  101.79 69.545 101.3 70.035 ;
      RECT  109.605 63.46 109.115 63.95 ;
      RECT  101.79 71.395 101.3 71.885 ;
      RECT  98.535 65.435 98.045 65.925 ;
      RECT  98.535 81.235 98.045 81.725 ;
      RECT  98.535 87.16 98.045 87.65 ;
      RECT  98.535 75.31 98.045 75.8 ;
      RECT  109.605 67.41 109.115 67.9 ;
      RECT  119.475 75.31 118.985 75.8 ;
      RECT  98.535 77.285 98.045 77.775 ;
      RECT  98.535 73.335 98.045 73.825 ;
      RECT  109.605 75.31 109.115 75.8 ;
      RECT  101.79 67.445 101.3 67.935 ;
      RECT  101.79 79.295 101.3 79.785 ;
      RECT  101.79 89.295 101.3 89.785 ;
      RECT  98.535 83.21 98.045 83.7 ;
      RECT  98.535 69.385 98.045 69.875 ;
      RECT  101.79 81.395 101.3 81.885 ;
      RECT  101.79 75.345 101.3 75.835 ;
      RECT  98.535 63.46 98.045 63.95 ;
      RECT  98.535 91.11 98.045 91.6 ;
      RECT  101.79 63.495 101.3 63.985 ;
      RECT  112.86 63.495 112.37 63.985 ;
      RECT  112.86 67.445 112.37 67.935 ;
      RECT  112.86 79.295 112.37 79.785 ;
      RECT  101.79 83.245 101.3 83.735 ;
      RECT  101.79 73.495 101.3 73.985 ;
      RECT  98.535 85.185 98.045 85.675 ;
      RECT  98.535 71.36 98.045 71.85 ;
      RECT  109.605 79.26 109.115 79.75 ;
      RECT  119.475 63.46 118.985 63.95 ;
      RECT  101.79 87.195 101.3 87.685 ;
      RECT  101.79 85.345 101.3 85.835 ;
      RECT  98.535 79.26 98.045 79.75 ;
      RECT  98.535 89.135 98.045 89.625 ;
      RECT  101.79 91.145 101.3 91.635 ;
      RECT  112.86 75.345 112.37 75.835 ;
      RECT  101.79 77.445 101.3 77.935 ;
      RECT  101.79 65.595 101.3 66.085 ;
      RECT  98.535 67.41 98.045 67.9 ;
      RECT  103.915 73.485 103.425 73.975 ;
      RECT  103.915 89.285 103.425 89.775 ;
      RECT  114.985 75.345 114.495 75.835 ;
      RECT  103.915 81.385 103.425 81.875 ;
      RECT  99.895 73.335 99.405 73.825 ;
      RECT  103.915 69.535 103.425 70.025 ;
      RECT  110.965 75.31 110.475 75.8 ;
      RECT  99.895 71.36 99.405 71.85 ;
      RECT  99.895 77.285 99.405 77.775 ;
      RECT  99.895 89.135 99.405 89.625 ;
      RECT  114.985 79.295 114.495 79.785 ;
      RECT  110.965 63.46 110.475 63.95 ;
      RECT  103.915 67.445 103.425 67.935 ;
      RECT  103.915 79.295 103.425 79.785 ;
      RECT  99.895 81.235 99.405 81.725 ;
      RECT  99.895 85.185 99.405 85.675 ;
      RECT  99.895 91.11 99.405 91.6 ;
      RECT  110.965 67.41 110.475 67.9 ;
      RECT  99.895 79.26 99.405 79.75 ;
      RECT  103.915 85.335 103.425 85.825 ;
      RECT  120.835 63.46 120.345 63.95 ;
      RECT  103.915 87.195 103.425 87.685 ;
      RECT  110.965 79.26 110.475 79.75 ;
      RECT  99.895 75.31 99.405 75.8 ;
      RECT  103.915 77.435 103.425 77.925 ;
      RECT  99.895 69.385 99.405 69.875 ;
      RECT  99.895 83.21 99.405 83.7 ;
      RECT  114.985 67.445 114.495 67.935 ;
      RECT  114.985 63.495 114.495 63.985 ;
      RECT  103.915 71.395 103.425 71.885 ;
      RECT  103.915 75.345 103.425 75.835 ;
      RECT  103.915 63.495 103.425 63.985 ;
      RECT  99.895 65.435 99.405 65.925 ;
      RECT  103.915 83.245 103.425 83.735 ;
      RECT  99.895 87.16 99.405 87.65 ;
      RECT  103.915 91.145 103.425 91.635 ;
      RECT  103.915 65.585 103.425 66.075 ;
      RECT  99.895 63.46 99.405 63.95 ;
      RECT  99.895 67.41 99.405 67.9 ;
      RECT  120.835 75.31 120.345 75.8 ;
      RECT  98.535 71.36 98.045 71.85 ;
      RECT  112.86 63.495 112.37 63.985 ;
      RECT  112.86 75.345 112.37 75.835 ;
      RECT  101.79 91.145 101.3 91.635 ;
      RECT  101.79 77.445 101.3 77.935 ;
      RECT  112.86 67.445 112.37 67.935 ;
      RECT  101.79 87.195 101.3 87.685 ;
      RECT  101.79 89.295 101.3 89.785 ;
      RECT  98.535 83.21 98.045 83.7 ;
      RECT  101.79 81.395 101.3 81.885 ;
      RECT  101.79 67.445 101.3 67.935 ;
      RECT  98.535 79.26 98.045 79.75 ;
      RECT  109.605 67.41 109.115 67.9 ;
      RECT  101.79 75.345 101.3 75.835 ;
      RECT  98.535 63.46 98.045 63.95 ;
      RECT  101.79 79.295 101.3 79.785 ;
      RECT  101.79 83.245 101.3 83.735 ;
      RECT  98.535 81.235 98.045 81.725 ;
      RECT  101.79 73.495 101.3 73.985 ;
      RECT  98.535 87.16 98.045 87.65 ;
      RECT  101.79 65.595 101.3 66.085 ;
      RECT  109.605 75.31 109.115 75.8 ;
      RECT  89.605 77.14 89.115 77.63 ;
      RECT  98.535 67.41 98.045 67.9 ;
      RECT  101.79 85.345 101.3 85.835 ;
      RECT  119.475 63.46 118.985 63.95 ;
      RECT  98.535 65.435 98.045 65.925 ;
      RECT  101.79 63.495 101.3 63.985 ;
      RECT  98.535 89.135 98.045 89.625 ;
      RECT  98.535 75.31 98.045 75.8 ;
      RECT  109.605 79.26 109.115 79.75 ;
      RECT  119.475 75.31 118.985 75.8 ;
      RECT  94.18 77.06 93.69 77.55 ;
      RECT  98.535 69.385 98.045 69.875 ;
      RECT  109.605 63.46 109.115 63.95 ;
      RECT  98.535 77.285 98.045 77.775 ;
      RECT  98.535 85.185 98.045 85.675 ;
      RECT  101.79 69.545 101.3 70.035 ;
      RECT  112.86 79.295 112.37 79.785 ;
      RECT  98.535 91.11 98.045 91.6 ;
      RECT  101.79 71.395 101.3 71.885 ;
      RECT  98.535 73.335 98.045 73.825 ;
      RECT  103.915 91.145 103.425 91.635 ;
      RECT  103.915 87.195 103.425 87.685 ;
      RECT  99.895 81.235 99.405 81.725 ;
      RECT  99.895 91.11 99.405 91.6 ;
      RECT  103.915 89.285 103.425 89.775 ;
      RECT  103.915 63.495 103.425 63.985 ;
      RECT  103.915 67.445 103.425 67.935 ;
      RECT  103.915 79.295 103.425 79.785 ;
      RECT  103.915 69.535 103.425 70.025 ;
      RECT  99.895 67.41 99.405 67.9 ;
      RECT  96.305 77.065 95.815 77.555 ;
      RECT  99.895 79.26 99.405 79.75 ;
      RECT  110.965 67.41 110.475 67.9 ;
      RECT  103.915 75.345 103.425 75.835 ;
      RECT  103.915 83.245 103.425 83.735 ;
      RECT  103.915 71.395 103.425 71.885 ;
      RECT  110.965 79.26 110.475 79.75 ;
      RECT  114.985 63.495 114.495 63.985 ;
      RECT  99.895 85.185 99.405 85.675 ;
      RECT  99.895 83.21 99.405 83.7 ;
      RECT  103.915 85.335 103.425 85.825 ;
      RECT  103.915 73.485 103.425 73.975 ;
      RECT  99.895 65.435 99.405 65.925 ;
      RECT  110.965 75.31 110.475 75.8 ;
      RECT  103.915 65.585 103.425 66.075 ;
      RECT  99.895 71.36 99.405 71.85 ;
      RECT  120.835 63.46 120.345 63.95 ;
      RECT  110.965 63.46 110.475 63.95 ;
      RECT  103.915 81.385 103.425 81.875 ;
      RECT  99.895 77.285 99.405 77.775 ;
      RECT  99.895 73.335 99.405 73.825 ;
      RECT  92.095 77.14 91.605 77.63 ;
      RECT  114.985 67.445 114.495 67.935 ;
      RECT  99.895 87.16 99.405 87.65 ;
      RECT  114.985 79.295 114.495 79.785 ;
      RECT  99.895 69.385 99.405 69.875 ;
      RECT  114.985 75.345 114.495 75.835 ;
      RECT  103.915 77.435 103.425 77.925 ;
      RECT  99.895 75.31 99.405 75.8 ;
      RECT  99.895 89.135 99.405 89.625 ;
      RECT  120.835 75.31 120.345 75.8 ;
      RECT  99.895 63.46 99.405 63.95 ;
      RECT  77.29 108.12 77.78 108.61 ;
      RECT  75.17 58.63 75.47 58.93 ;
      RECT  101.3 79.295 101.79 79.785 ;
      RECT  98.045 83.21 98.535 83.7 ;
      RECT  51.97 65.595 52.46 66.085 ;
      RECT  98.045 65.435 98.535 65.925 ;
      RECT  75.42 41.97 75.91 42.46 ;
      RECT  55.225 65.435 55.715 65.925 ;
      RECT  112.37 67.445 112.86 67.935 ;
      RECT  109.115 63.46 109.605 63.95 ;
      RECT  44.155 63.46 44.645 63.95 ;
      RECT  101.3 71.395 101.79 71.885 ;
      RECT  75.36 46.16 75.85 46.65 ;
      RECT  55.225 67.41 55.715 67.9 ;
      RECT  98.045 85.185 98.535 85.675 ;
      RECT  101.3 69.545 101.79 70.035 ;
      RECT  98.045 67.41 98.535 67.9 ;
      RECT  109.115 79.26 109.605 79.75 ;
      RECT  55.225 91.11 55.715 91.6 ;
      RECT  51.97 81.395 52.46 81.885 ;
      RECT  101.3 73.495 101.79 73.985 ;
      RECT  44.155 67.41 44.645 67.9 ;
      RECT  109.115 75.31 109.605 75.8 ;
      RECT  51.97 79.295 52.46 79.785 ;
      RECT  55.225 69.385 55.715 69.875 ;
      RECT  98.045 75.31 98.535 75.8 ;
      RECT  55.225 89.135 55.715 89.625 ;
      RECT  51.97 69.545 52.46 70.035 ;
      RECT  51.97 89.295 52.46 89.785 ;
      RECT  89.115 77.14 89.605 77.63 ;
      RECT  101.3 87.195 101.79 87.685 ;
      RECT  55.225 63.46 55.715 63.95 ;
      RECT  98.045 71.36 98.535 71.85 ;
      RECT  44.155 75.31 44.645 75.8 ;
      RECT  78.29 95.84 78.59 96.14 ;
      RECT  80.72 98.7 81.21 99.19 ;
      RECT  77.855 34.21 78.345 34.7 ;
      RECT  98.045 91.11 98.535 91.6 ;
      RECT  51.97 91.145 52.46 91.635 ;
      RECT  101.3 63.495 101.79 63.985 ;
      RECT  34.285 75.31 34.775 75.8 ;
      RECT  51.97 63.495 52.46 63.985 ;
      RECT  112.37 75.345 112.86 75.835 ;
      RECT  44.155 79.26 44.645 79.75 ;
      RECT  55.225 75.31 55.715 75.8 ;
      RECT  77.23 41.97 77.72 42.46 ;
      RECT  64.155 77.14 64.645 77.63 ;
      RECT  51.97 77.445 52.46 77.935 ;
      RECT  74.48 98.7 74.97 99.19 ;
      RECT  78.79 98.7 79.28 99.19 ;
      RECT  74.895 29.46 75.385 29.95 ;
      RECT  93.69 77.06 94.18 77.55 ;
      RECT  101.3 89.295 101.79 89.785 ;
      RECT  55.225 73.335 55.715 73.825 ;
      RECT  98.045 89.135 98.535 89.625 ;
      RECT  51.97 71.395 52.46 71.885 ;
      RECT  55.225 87.16 55.715 87.65 ;
      RECT  71.955 95.745 72.445 96.235 ;
      RECT  98.045 77.285 98.535 77.775 ;
      RECT  40.9 75.345 41.39 75.835 ;
      RECT  101.3 83.245 101.79 83.735 ;
      RECT  51.97 75.345 52.46 75.835 ;
      RECT  101.3 75.345 101.79 75.835 ;
      RECT  112.37 63.495 112.86 63.985 ;
      RECT  51.97 67.445 52.46 67.935 ;
      RECT  78.29 58.63 78.59 58.93 ;
      RECT  55.225 79.26 55.715 79.75 ;
      RECT  40.9 63.495 41.39 63.985 ;
      RECT  72.55 55.58 73.04 56.07 ;
      RECT  59.58 77.06 60.07 77.55 ;
      RECT  78.79 55.58 79.28 56.07 ;
      RECT  75.36 108.12 75.85 108.61 ;
      RECT  77.23 112.31 77.72 112.8 ;
      RECT  40.9 67.445 41.39 67.935 ;
      RECT  55.225 85.185 55.715 85.675 ;
      RECT  101.3 81.395 101.79 81.885 ;
      RECT  118.985 63.46 119.475 63.95 ;
      RECT  81.315 58.535 81.805 59.025 ;
      RECT  51.97 83.245 52.46 83.735 ;
      RECT  51.97 87.195 52.46 87.685 ;
      RECT  77.29 46.16 77.78 46.65 ;
      RECT  51.97 85.345 52.46 85.835 ;
      RECT  98.045 63.46 98.535 63.95 ;
      RECT  101.3 65.595 101.79 66.085 ;
      RECT  118.985 75.31 119.475 75.8 ;
      RECT  101.3 91.145 101.79 91.635 ;
      RECT  40.9 79.295 41.39 79.785 ;
      RECT  55.225 81.235 55.715 81.725 ;
      RECT  55.225 83.21 55.715 83.7 ;
      RECT  55.225 77.285 55.715 77.775 ;
      RECT  98.045 81.235 98.535 81.725 ;
      RECT  71.955 58.535 72.445 59.025 ;
      RECT  74.795 34.21 75.285 34.7 ;
      RECT  98.045 87.16 98.535 87.65 ;
      RECT  112.37 79.295 112.86 79.785 ;
      RECT  98.045 79.26 98.535 79.75 ;
      RECT  109.115 67.41 109.605 67.9 ;
      RECT  98.045 69.385 98.535 69.875 ;
      RECT  101.3 85.345 101.79 85.835 ;
      RECT  75.42 112.31 75.91 112.8 ;
      RECT  98.045 73.335 98.535 73.825 ;
      RECT  75.17 95.84 75.47 96.14 ;
      RECT  34.285 63.46 34.775 63.95 ;
      RECT  74.48 55.58 74.97 56.07 ;
      RECT  101.3 77.445 101.79 77.935 ;
      RECT  101.3 67.445 101.79 67.935 ;
      RECT  55.225 71.36 55.715 71.85 ;
      RECT  51.97 73.495 52.46 73.985 ;
      RECT  81.315 95.745 81.805 96.235 ;
      RECT  77.755 29.46 78.245 29.95 ;
      RECT  68.57 65.385 68.87 65.685 ;
      RECT  49.845 71.395 50.335 71.885 ;
      RECT  84.89 66.57 85.19 66.87 ;
      RECT  53.865 83.21 54.355 83.7 ;
      RECT  103.425 81.385 103.915 81.875 ;
      RECT  68.57 68.15 68.87 68.45 ;
      RECT  68.57 64.2 68.87 64.5 ;
      RECT  84.89 86.32 85.19 86.62 ;
      RECT  68.57 85.135 68.87 85.435 ;
      RECT  84.89 64.2 85.19 64.5 ;
      RECT  99.405 91.11 99.895 91.6 ;
      RECT  84.89 91.85 85.19 92.15 ;
      RECT  53.865 69.385 54.355 69.875 ;
      RECT  68.57 78.42 68.87 78.72 ;
      RECT  84.89 89.085 85.19 89.385 ;
      RECT  84.89 77.235 85.19 77.535 ;
      RECT  103.425 65.585 103.915 66.075 ;
      RECT  68.57 90.27 68.87 90.57 ;
      RECT  53.865 89.135 54.355 89.625 ;
      RECT  53.865 75.31 54.355 75.8 ;
      RECT  99.405 71.36 99.895 71.85 ;
      RECT  84.89 73.285 85.19 73.585 ;
      RECT  42.795 79.26 43.285 79.75 ;
      RECT  103.425 63.495 103.915 63.985 ;
      RECT  68.57 70.52 68.87 70.82 ;
      RECT  84.89 61.435 85.19 61.735 ;
      RECT  68.57 69.335 68.87 69.635 ;
      RECT  84.89 65.385 85.19 65.685 ;
      RECT  84.89 90.27 85.19 90.57 ;
      RECT  103.425 87.195 103.915 87.685 ;
      RECT  99.405 87.16 99.895 87.65 ;
      RECT  84.89 68.15 85.19 68.45 ;
      RECT  53.865 87.16 54.355 87.65 ;
      RECT  49.845 81.385 50.335 81.875 ;
      RECT  68.57 77.235 68.87 77.535 ;
      RECT  77.825 31.54 78.315 32.03 ;
      RECT  120.345 75.31 120.835 75.8 ;
      RECT  84.89 94.22 85.19 94.52 ;
      RECT  120.345 63.46 120.835 63.95 ;
      RECT  68.57 89.085 68.87 89.385 ;
      RECT  75.42 40.36 75.91 40.85 ;
      RECT  68.57 82.37 68.87 82.67 ;
      RECT  99.405 73.335 99.895 73.825 ;
      RECT  49.845 69.535 50.335 70.025 ;
      RECT  103.425 79.295 103.915 79.785 ;
      RECT  77.23 113.92 77.72 114.41 ;
      RECT  42.795 67.41 43.285 67.9 ;
      RECT  53.865 85.185 54.355 85.675 ;
      RECT  38.775 63.495 39.265 63.985 ;
      RECT  114.495 75.345 114.985 75.835 ;
      RECT  68.57 81.185 68.87 81.485 ;
      RECT  103.425 83.245 103.915 83.735 ;
      RECT  84.89 82.37 85.19 82.67 ;
      RECT  84.89 72.1 85.19 72.4 ;
      RECT  53.865 73.335 54.355 73.825 ;
      RECT  38.775 67.445 39.265 67.935 ;
      RECT  84.89 69.335 85.19 69.635 ;
      RECT  114.495 63.495 114.985 63.985 ;
      RECT  49.845 73.485 50.335 73.975 ;
      RECT  68.57 60.25 68.87 60.55 ;
      RECT  49.845 63.495 50.335 63.985 ;
      RECT  53.865 71.36 54.355 71.85 ;
      RECT  84.89 74.47 85.19 74.77 ;
      RECT  49.845 65.585 50.335 66.075 ;
      RECT  32.925 63.46 33.415 63.95 ;
      RECT  103.425 71.395 103.915 71.885 ;
      RECT  49.845 87.195 50.335 87.685 ;
      RECT  84.89 78.42 85.19 78.72 ;
      RECT  84.89 62.62 85.19 62.92 ;
      RECT  84.89 60.25 85.19 60.55 ;
      RECT  84.89 83.95 85.19 84.25 ;
      RECT  84.89 87.9 85.19 88.2 ;
      RECT  68.57 94.22 68.87 94.52 ;
      RECT  84.89 76.05 85.19 76.35 ;
      RECT  53.865 79.26 54.355 79.75 ;
      RECT  68.57 86.32 68.87 86.62 ;
      RECT  99.405 67.41 99.895 67.9 ;
      RECT  75.77 50.03 76.26 50.52 ;
      RECT  53.865 81.235 54.355 81.725 ;
      RECT  103.425 73.485 103.915 73.975 ;
      RECT  68.57 83.95 68.87 84.25 ;
      RECT  110.475 67.41 110.965 67.9 ;
      RECT  95.815 77.065 96.305 77.555 ;
      RECT  74.85 36.395 75.34 36.885 ;
      RECT  103.425 89.285 103.915 89.775 ;
      RECT  49.845 75.345 50.335 75.835 ;
      RECT  53.865 65.435 54.355 65.925 ;
      RECT  103.425 75.345 103.915 75.835 ;
      RECT  99.405 69.385 99.895 69.875 ;
      RECT  91.605 77.14 92.095 77.63 ;
      RECT  68.57 87.9 68.87 88.2 ;
      RECT  49.845 91.145 50.335 91.635 ;
      RECT  38.775 75.345 39.265 75.835 ;
      RECT  76.88 50.03 77.37 50.52 ;
      RECT  99.405 77.285 99.895 77.775 ;
      RECT  68.57 66.57 68.87 66.87 ;
      RECT  99.405 83.21 99.895 83.7 ;
      RECT  49.845 85.335 50.335 85.825 ;
      RECT  99.405 65.435 99.895 65.925 ;
      RECT  77.8 36.395 78.29 36.885 ;
      RECT  110.475 75.31 110.965 75.8 ;
      RECT  68.57 76.05 68.87 76.35 ;
      RECT  99.405 81.235 99.895 81.725 ;
      RECT  114.495 79.295 114.985 79.785 ;
      RECT  38.775 79.295 39.265 79.785 ;
      RECT  49.845 79.295 50.335 79.785 ;
      RECT  42.795 63.46 43.285 63.95 ;
      RECT  75.77 104.25 76.26 104.74 ;
      RECT  75.42 113.92 75.91 114.41 ;
      RECT  53.865 91.11 54.355 91.6 ;
      RECT  84.89 93.035 85.19 93.335 ;
      RECT  53.865 67.41 54.355 67.9 ;
      RECT  61.665 77.14 62.155 77.63 ;
      RECT  99.405 75.31 99.895 75.8 ;
      RECT  74.825 31.54 75.315 32.03 ;
      RECT  68.57 73.285 68.87 73.585 ;
      RECT  68.57 61.435 68.87 61.735 ;
      RECT  114.495 67.445 114.985 67.935 ;
      RECT  103.425 67.445 103.915 67.935 ;
      RECT  42.795 75.31 43.285 75.8 ;
      RECT  76.88 104.25 77.37 104.74 ;
      RECT  49.845 67.445 50.335 67.935 ;
      RECT  49.845 89.285 50.335 89.775 ;
      RECT  110.475 79.26 110.965 79.75 ;
      RECT  49.845 83.245 50.335 83.735 ;
      RECT  103.425 77.435 103.915 77.925 ;
      RECT  110.475 63.46 110.965 63.95 ;
      RECT  103.425 91.145 103.915 91.635 ;
      RECT  49.845 77.435 50.335 77.925 ;
      RECT  103.425 85.335 103.915 85.825 ;
      RECT  68.57 74.47 68.87 74.77 ;
      RECT  99.405 79.26 99.895 79.75 ;
      RECT  77.25 32.55 77.74 33.04 ;
      RECT  99.405 89.135 99.895 89.625 ;
      RECT  57.455 77.065 57.945 77.555 ;
      RECT  84.89 81.185 85.19 81.485 ;
      RECT  84.89 85.135 85.19 85.435 ;
      RECT  68.57 93.035 68.87 93.335 ;
      RECT  103.425 69.535 103.915 70.025 ;
      RECT  53.865 63.46 54.355 63.95 ;
      RECT  68.57 62.62 68.87 62.92 ;
      RECT  68.57 72.1 68.87 72.4 ;
      RECT  53.865 77.285 54.355 77.775 ;
      RECT  77.23 40.36 77.72 40.85 ;
      RECT  99.405 85.185 99.895 85.675 ;
      RECT  68.57 80.0 68.87 80.3 ;
      RECT  84.89 80.0 85.19 80.3 ;
      RECT  68.57 91.85 68.87 92.15 ;
      RECT  75.4 32.55 75.89 33.04 ;
      RECT  99.405 63.46 99.895 63.95 ;
      RECT  32.925 75.31 33.415 75.8 ;
      RECT  84.89 70.52 85.19 70.82 ;
      RECT  0.435 7.1 0.925 7.59 ;
      RECT  0.435 0.02 0.925 0.51 ;
      RECT  0.435 14.18 0.925 14.67 ;
      RECT  6.845 62.99 6.355 63.48 ;
      RECT  3.165 62.99 2.675 63.48 ;
      RECT  6.845 62.99 6.355 63.48 ;
      RECT  3.165 74.19 2.675 74.68 ;
      RECT  3.165 62.99 2.675 63.48 ;
      RECT  3.165 74.19 2.675 74.68 ;
      RECT  3.165 85.39 2.675 85.88 ;
      RECT  3.165 107.79 2.675 108.28 ;
      RECT  6.845 74.19 6.355 74.68 ;
      RECT  6.845 74.19 6.355 74.68 ;
      RECT  6.845 85.39 6.355 85.88 ;
      RECT  6.845 96.59 6.355 97.08 ;
      RECT  3.165 96.59 2.675 97.08 ;
      RECT  6.845 107.79 6.355 108.28 ;
      RECT  6.845 68.59 6.355 69.08 ;
      RECT  3.165 102.19 2.675 102.68 ;
      RECT  6.845 79.79 6.355 80.28 ;
      RECT  6.845 90.99 6.355 91.48 ;
      RECT  3.165 90.99 2.675 91.48 ;
      RECT  6.845 102.19 6.355 102.68 ;
      RECT  3.165 79.79 2.675 80.28 ;
      RECT  6.845 57.39 6.355 57.88 ;
      RECT  3.165 68.59 2.675 69.08 ;
      RECT  3.165 57.39 2.675 57.88 ;
      RECT  27.245 49.52 27.735 50.01 ;
      RECT  6.355 74.19 6.845 74.68 ;
      RECT  2.675 62.99 3.165 63.48 ;
      RECT  27.245 35.38 27.735 35.87 ;
      RECT  27.245 7.1 27.735 7.59 ;
      RECT  2.675 96.59 3.165 97.08 ;
      RECT  6.355 85.39 6.845 85.88 ;
      RECT  6.355 62.99 6.845 63.48 ;
      RECT  2.675 107.79 3.165 108.28 ;
      RECT  6.355 107.79 6.845 108.28 ;
      RECT  0.435 7.1 0.925 7.59 ;
      RECT  27.245 21.24 27.735 21.73 ;
      RECT  2.675 74.19 3.165 74.68 ;
      RECT  6.355 96.59 6.845 97.08 ;
      RECT  2.675 85.39 3.165 85.88 ;
      RECT  27.245 42.45 27.735 42.94 ;
      RECT  6.355 79.79 6.845 80.28 ;
      RECT  27.245 0.03 27.735 0.52 ;
      RECT  6.355 68.59 6.845 69.08 ;
      RECT  6.355 102.19 6.845 102.68 ;
      RECT  2.675 68.59 3.165 69.08 ;
      RECT  6.355 57.39 6.845 57.88 ;
      RECT  2.675 57.39 3.165 57.88 ;
      RECT  0.435 0.02 0.925 0.51 ;
      RECT  6.355 90.99 6.845 91.48 ;
      RECT  27.245 56.59 27.735 57.08 ;
      RECT  27.245 28.31 27.735 28.8 ;
      RECT  2.675 102.19 3.165 102.68 ;
      RECT  2.675 90.99 3.165 91.48 ;
      RECT  2.675 79.79 3.165 80.28 ;
      RECT  0.435 14.18 0.925 14.67 ;
      RECT  27.245 14.17 27.735 14.66 ;
      RECT  152.215 133.53 151.725 133.04 ;
      RECT  152.215 140.61 151.725 140.12 ;
      RECT  145.805 91.78 146.295 91.29 ;
      RECT  149.485 91.78 149.975 91.29 ;
      RECT  145.805 91.78 146.295 91.29 ;
      RECT  149.485 80.58 149.975 80.09 ;
      RECT  149.485 91.78 149.975 91.29 ;
      RECT  149.485 80.58 149.975 80.09 ;
      RECT  149.485 69.38 149.975 68.89 ;
      RECT  149.485 46.98 149.975 46.49 ;
      RECT  145.805 80.58 146.295 80.09 ;
      RECT  145.805 80.58 146.295 80.09 ;
      RECT  145.805 69.38 146.295 68.89 ;
      RECT  145.805 58.18 146.295 57.69 ;
      RECT  149.485 58.18 149.975 57.69 ;
      RECT  145.805 46.98 146.295 46.49 ;
      RECT  145.805 86.18 146.295 85.69 ;
      RECT  149.485 52.58 149.975 52.09 ;
      RECT  145.805 74.98 146.295 74.49 ;
      RECT  145.805 63.78 146.295 63.29 ;
      RECT  149.485 63.78 149.975 63.29 ;
      RECT  145.805 52.58 146.295 52.09 ;
      RECT  149.485 74.98 149.975 74.49 ;
      RECT  145.805 97.38 146.295 96.89 ;
      RECT  149.485 86.18 149.975 85.69 ;
      RECT  149.485 97.38 149.975 96.89 ;
      RECT  146.295 69.38 145.805 68.89 ;
      RECT  146.295 58.18 145.805 57.69 ;
      RECT  126.935 133.53 126.445 133.04 ;
      RECT  149.975 46.98 149.485 46.49 ;
      RECT  149.975 58.18 149.485 57.69 ;
      RECT  126.935 119.39 126.445 118.9 ;
      RECT  146.295 91.78 145.805 91.29 ;
      RECT  146.295 46.98 145.805 46.49 ;
      RECT  146.295 80.58 145.805 80.09 ;
      RECT  149.975 91.78 149.485 91.29 ;
      RECT  149.975 80.58 149.485 80.09 ;
      RECT  126.935 105.25 126.445 104.76 ;
      RECT  152.215 133.53 151.725 133.04 ;
      RECT  149.975 69.38 149.485 68.89 ;
      RECT  146.295 86.18 145.805 85.69 ;
      RECT  126.935 98.18 126.445 97.69 ;
      RECT  126.935 126.46 126.445 125.97 ;
      RECT  146.295 74.98 145.805 74.49 ;
      RECT  146.295 63.78 145.805 63.29 ;
      RECT  149.975 74.98 149.485 74.49 ;
      RECT  146.295 97.38 145.805 96.89 ;
      RECT  152.215 140.61 151.725 140.12 ;
      RECT  149.975 86.18 149.485 85.69 ;
      RECT  149.975 97.38 149.485 96.89 ;
      RECT  146.295 52.58 145.805 52.09 ;
      RECT  149.975 52.58 149.485 52.09 ;
      RECT  126.935 112.32 126.445 111.83 ;
      RECT  149.975 63.78 149.485 63.29 ;
      RECT  126.935 140.6 126.445 140.11 ;
      RECT  22.07 110.225 27.91 110.525 ;
      RECT  24.745 115.66 25.235 116.15 ;
      RECT  24.745 129.8 25.235 130.29 ;
      RECT  24.745 136.87 25.235 137.36 ;
      RECT  24.745 122.73 25.235 123.22 ;
      RECT  24.745 108.59 25.235 109.08 ;
      RECT  132.11 44.545 126.27 44.245 ;
      RECT  129.435 39.11 128.945 38.62 ;
      RECT  129.435 24.97 128.945 24.48 ;
      RECT  129.435 17.9 128.945 17.41 ;
      RECT  129.435 32.04 128.945 31.55 ;
      RECT  129.435 46.18 128.945 45.69 ;
      RECT  33.75 14.53 45.43 14.83 ;
      RECT  42.265 19.965 42.755 20.455 ;
      RECT  36.425 19.965 36.915 20.455 ;
      RECT  42.265 12.895 42.755 13.385 ;
      RECT  36.425 12.895 36.915 13.385 ;
   LAYER  m4 ;
   END
   END    sram_1rw1r_2_16_sky130
END    LIBRARY
