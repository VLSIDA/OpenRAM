VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 1000 ;
END UNITS
SITE  MacroSite
   CLASS Core ;
   SIZE 2250.0 by 1200.0 ;
END  MacroSite
MACRO sram_2_16_1_scn3me_subm
   CLASS BLOCK ;
   SIZE 2250.0 BY 1200.0 ;
   SYMMETRY X Y R90 ;
   SITE MacroSite ;
   PIN DATA[0]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  180300.0 0.0 181200.0 1800.0 ;
      END
   END DATA[0]
   PIN DATA[1]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  190500.0 0.0 191400.0 1800.0 ;
      END
   END DATA[1]
   PIN ADDR[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  53100.0 75000.0 60300.0 76500.0 ;
      END
   END ADDR[0]
   PIN ADDR[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  53100.0 64800.0 60300.0 66300.0 ;
      END
   END ADDR[1]
   PIN ADDR[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  53100.0 54600.0 60300.0 56100.0 ;
      END
   END ADDR[2]
   PIN ADDR[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  53100.0 44400.0 60300.0 45900.0 ;
      END
   END ADDR[3]
   PIN CSb
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  14400.0 203100.0 16200.0 204900.0 ;
      END
   END CSb
   PIN WEb
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  24600.0 203100.0 26400.0 204900.0 ;
      END
   END WEb
   PIN OEb
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  4200.0 203100.0 6000.0 204900.0 ;
      END
   END OEb
   PIN clk
      DIRECTION INPUT ;
      PORT
         LAYER metal1 ;
         RECT  43050.0 202200.0 44250.0 205800.0 ;
      END
   END clk
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal1 ;
         RECT  198900.0 0.0 203400.0 444600.0 ;
         LAYER metal1 ;
         RECT  53100.0 0.0 57600.0 444600.0 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal2 ;
         RECT  148350.0 0.0 152850.0 444600.0 ;
      END
   END gnd
   OBS
   LAYER  metal1 ;
      RECT  54900.0 295650.0 55800.0 298350.0 ;
      RECT  97800.0 205200.0 98700.0 206100.0 ;
      RECT  97800.0 202950.0 98700.0 203850.0 ;
      RECT  96450.0 205200.0 98250.0 206100.0 ;
      RECT  97800.0 203400.0 98700.0 205650.0 ;
      RECT  98250.0 202950.0 100200.0 203850.0 ;
      RECT  155250.0 205200.0 156150.0 206100.0 ;
      RECT  155250.0 201450.0 156150.0 202350.0 ;
      RECT  136350.0 205200.0 155700.0 206100.0 ;
      RECT  155250.0 201900.0 156150.0 205650.0 ;
      RECT  155700.0 201450.0 175200.0 202350.0 ;
      RECT  97800.0 220500.0 98700.0 221400.0 ;
      RECT  97800.0 222750.0 98700.0 223650.0 ;
      RECT  96450.0 220500.0 98250.0 221400.0 ;
      RECT  97800.0 220950.0 98700.0 223200.0 ;
      RECT  98250.0 222750.0 100200.0 223650.0 ;
      RECT  155250.0 220500.0 156150.0 221400.0 ;
      RECT  155250.0 224250.0 156150.0 225150.0 ;
      RECT  136350.0 220500.0 155700.0 221400.0 ;
      RECT  155250.0 220950.0 156150.0 224700.0 ;
      RECT  155700.0 224250.0 175200.0 225150.0 ;
      RECT  97800.0 233400.0 98700.0 234300.0 ;
      RECT  97800.0 231150.0 98700.0 232050.0 ;
      RECT  96450.0 233400.0 98250.0 234300.0 ;
      RECT  97800.0 231600.0 98700.0 233850.0 ;
      RECT  98250.0 231150.0 100200.0 232050.0 ;
      RECT  155250.0 233400.0 156150.0 234300.0 ;
      RECT  155250.0 229650.0 156150.0 230550.0 ;
      RECT  136350.0 233400.0 155700.0 234300.0 ;
      RECT  155250.0 230100.0 156150.0 233850.0 ;
      RECT  155700.0 229650.0 175200.0 230550.0 ;
      RECT  97800.0 248700.0 98700.0 249600.0 ;
      RECT  97800.0 250950.0 98700.0 251850.0 ;
      RECT  96450.0 248700.0 98250.0 249600.0 ;
      RECT  97800.0 249150.0 98700.0 251400.0 ;
      RECT  98250.0 250950.0 100200.0 251850.0 ;
      RECT  155250.0 248700.0 156150.0 249600.0 ;
      RECT  155250.0 252450.0 156150.0 253350.0 ;
      RECT  136350.0 248700.0 155700.0 249600.0 ;
      RECT  155250.0 249150.0 156150.0 252900.0 ;
      RECT  155700.0 252450.0 175200.0 253350.0 ;
      RECT  97800.0 261600.0 98700.0 262500.0 ;
      RECT  97800.0 259350.0 98700.0 260250.0 ;
      RECT  96450.0 261600.0 98250.0 262500.0 ;
      RECT  97800.0 259800.0 98700.0 262050.0 ;
      RECT  98250.0 259350.0 100200.0 260250.0 ;
      RECT  155250.0 261600.0 156150.0 262500.0 ;
      RECT  155250.0 257850.0 156150.0 258750.0 ;
      RECT  136350.0 261600.0 155700.0 262500.0 ;
      RECT  155250.0 258300.0 156150.0 262050.0 ;
      RECT  155700.0 257850.0 175200.0 258750.0 ;
      RECT  97800.0 276900.0 98700.0 277800.0 ;
      RECT  97800.0 279150.0 98700.0 280050.0 ;
      RECT  96450.0 276900.0 98250.0 277800.0 ;
      RECT  97800.0 277350.0 98700.0 279600.0 ;
      RECT  98250.0 279150.0 100200.0 280050.0 ;
      RECT  155250.0 276900.0 156150.0 277800.0 ;
      RECT  155250.0 280650.0 156150.0 281550.0 ;
      RECT  136350.0 276900.0 155700.0 277800.0 ;
      RECT  155250.0 277350.0 156150.0 281100.0 ;
      RECT  155700.0 280650.0 175200.0 281550.0 ;
      RECT  97800.0 289800.0 98700.0 290700.0 ;
      RECT  97800.0 287550.0 98700.0 288450.0 ;
      RECT  96450.0 289800.0 98250.0 290700.0 ;
      RECT  97800.0 288000.0 98700.0 290250.0 ;
      RECT  98250.0 287550.0 100200.0 288450.0 ;
      RECT  155250.0 289800.0 156150.0 290700.0 ;
      RECT  155250.0 286050.0 156150.0 286950.0 ;
      RECT  136350.0 289800.0 155700.0 290700.0 ;
      RECT  155250.0 286500.0 156150.0 290250.0 ;
      RECT  155700.0 286050.0 175200.0 286950.0 ;
      RECT  97800.0 305100.0 98700.0 306000.0 ;
      RECT  97800.0 307350.0 98700.0 308250.0 ;
      RECT  96450.0 305100.0 98250.0 306000.0 ;
      RECT  97800.0 305550.0 98700.0 307800.0 ;
      RECT  98250.0 307350.0 100200.0 308250.0 ;
      RECT  155250.0 305100.0 156150.0 306000.0 ;
      RECT  155250.0 308850.0 156150.0 309750.0 ;
      RECT  136350.0 305100.0 155700.0 306000.0 ;
      RECT  155250.0 305550.0 156150.0 309300.0 ;
      RECT  155700.0 308850.0 175200.0 309750.0 ;
      RECT  97800.0 318000.0 98700.0 318900.0 ;
      RECT  97800.0 315750.0 98700.0 316650.0 ;
      RECT  96450.0 318000.0 98250.0 318900.0 ;
      RECT  97800.0 316200.0 98700.0 318450.0 ;
      RECT  98250.0 315750.0 100200.0 316650.0 ;
      RECT  155250.0 318000.0 156150.0 318900.0 ;
      RECT  155250.0 314250.0 156150.0 315150.0 ;
      RECT  136350.0 318000.0 155700.0 318900.0 ;
      RECT  155250.0 314700.0 156150.0 318450.0 ;
      RECT  155700.0 314250.0 175200.0 315150.0 ;
      RECT  97800.0 333300.0 98700.0 334200.0 ;
      RECT  97800.0 335550.0 98700.0 336450.0 ;
      RECT  96450.0 333300.0 98250.0 334200.0 ;
      RECT  97800.0 333750.0 98700.0 336000.0 ;
      RECT  98250.0 335550.0 100200.0 336450.0 ;
      RECT  155250.0 333300.0 156150.0 334200.0 ;
      RECT  155250.0 337050.0 156150.0 337950.0 ;
      RECT  136350.0 333300.0 155700.0 334200.0 ;
      RECT  155250.0 333750.0 156150.0 337500.0 ;
      RECT  155700.0 337050.0 175200.0 337950.0 ;
      RECT  97800.0 346200.0 98700.0 347100.0 ;
      RECT  97800.0 343950.0 98700.0 344850.0 ;
      RECT  96450.0 346200.0 98250.0 347100.0 ;
      RECT  97800.0 344400.0 98700.0 346650.0 ;
      RECT  98250.0 343950.0 100200.0 344850.0 ;
      RECT  155250.0 346200.0 156150.0 347100.0 ;
      RECT  155250.0 342450.0 156150.0 343350.0 ;
      RECT  136350.0 346200.0 155700.0 347100.0 ;
      RECT  155250.0 342900.0 156150.0 346650.0 ;
      RECT  155700.0 342450.0 175200.0 343350.0 ;
      RECT  97800.0 361500.0 98700.0 362400.0 ;
      RECT  97800.0 363750.0 98700.0 364650.0 ;
      RECT  96450.0 361500.0 98250.0 362400.0 ;
      RECT  97800.0 361950.0 98700.0 364200.0 ;
      RECT  98250.0 363750.0 100200.0 364650.0 ;
      RECT  155250.0 361500.0 156150.0 362400.0 ;
      RECT  155250.0 365250.0 156150.0 366150.0 ;
      RECT  136350.0 361500.0 155700.0 362400.0 ;
      RECT  155250.0 361950.0 156150.0 365700.0 ;
      RECT  155700.0 365250.0 175200.0 366150.0 ;
      RECT  97800.0 374400.0 98700.0 375300.0 ;
      RECT  97800.0 372150.0 98700.0 373050.0 ;
      RECT  96450.0 374400.0 98250.0 375300.0 ;
      RECT  97800.0 372600.0 98700.0 374850.0 ;
      RECT  98250.0 372150.0 100200.0 373050.0 ;
      RECT  155250.0 374400.0 156150.0 375300.0 ;
      RECT  155250.0 370650.0 156150.0 371550.0 ;
      RECT  136350.0 374400.0 155700.0 375300.0 ;
      RECT  155250.0 371100.0 156150.0 374850.0 ;
      RECT  155700.0 370650.0 175200.0 371550.0 ;
      RECT  97800.0 389700.0 98700.0 390600.0 ;
      RECT  97800.0 391950.0 98700.0 392850.0 ;
      RECT  96450.0 389700.0 98250.0 390600.0 ;
      RECT  97800.0 390150.0 98700.0 392400.0 ;
      RECT  98250.0 391950.0 100200.0 392850.0 ;
      RECT  155250.0 389700.0 156150.0 390600.0 ;
      RECT  155250.0 393450.0 156150.0 394350.0 ;
      RECT  136350.0 389700.0 155700.0 390600.0 ;
      RECT  155250.0 390150.0 156150.0 393900.0 ;
      RECT  155700.0 393450.0 175200.0 394350.0 ;
      RECT  97800.0 402600.0 98700.0 403500.0 ;
      RECT  97800.0 400350.0 98700.0 401250.0 ;
      RECT  96450.0 402600.0 98250.0 403500.0 ;
      RECT  97800.0 400800.0 98700.0 403050.0 ;
      RECT  98250.0 400350.0 100200.0 401250.0 ;
      RECT  155250.0 402600.0 156150.0 403500.0 ;
      RECT  155250.0 398850.0 156150.0 399750.0 ;
      RECT  136350.0 402600.0 155700.0 403500.0 ;
      RECT  155250.0 399300.0 156150.0 403050.0 ;
      RECT  155700.0 398850.0 175200.0 399750.0 ;
      RECT  97800.0 417900.0 98700.0 418800.0 ;
      RECT  97800.0 420150.0 98700.0 421050.0 ;
      RECT  96450.0 417900.0 98250.0 418800.0 ;
      RECT  97800.0 418350.0 98700.0 420600.0 ;
      RECT  98250.0 420150.0 100200.0 421050.0 ;
      RECT  155250.0 417900.0 156150.0 418800.0 ;
      RECT  155250.0 421650.0 156150.0 422550.0 ;
      RECT  136350.0 417900.0 155700.0 418800.0 ;
      RECT  155250.0 418350.0 156150.0 422100.0 ;
      RECT  155700.0 421650.0 175200.0 422550.0 ;
      RECT  106500.0 198750.0 175800.0 199650.0 ;
      RECT  106500.0 226950.0 175800.0 227850.0 ;
      RECT  106500.0 255150.0 175800.0 256050.0 ;
      RECT  106500.0 283350.0 175800.0 284250.0 ;
      RECT  106500.0 311550.0 175800.0 312450.0 ;
      RECT  106500.0 339750.0 175800.0 340650.0 ;
      RECT  106500.0 367950.0 175800.0 368850.0 ;
      RECT  106500.0 396150.0 175800.0 397050.0 ;
      RECT  106500.0 424350.0 175800.0 425250.0 ;
      RECT  53100.0 212850.0 203400.0 213750.0 ;
      RECT  53100.0 241050.0 203400.0 241950.0 ;
      RECT  53100.0 269250.0 203400.0 270150.0 ;
      RECT  53100.0 297450.0 203400.0 298350.0 ;
      RECT  53100.0 325650.0 203400.0 326550.0 ;
      RECT  53100.0 353850.0 203400.0 354750.0 ;
      RECT  53100.0 382050.0 203400.0 382950.0 ;
      RECT  53100.0 410250.0 203400.0 411150.0 ;
      RECT  130800.0 88650.0 135300.0 89550.0 ;
      RECT  127800.0 102750.0 138000.0 103650.0 ;
      RECT  130800.0 145050.0 140700.0 145950.0 ;
      RECT  127800.0 159150.0 143400.0 160050.0 ;
      RECT  130800.0 85950.0 132300.0 86850.0 ;
      RECT  130800.0 114150.0 132300.0 115050.0 ;
      RECT  130800.0 142350.0 132300.0 143250.0 ;
      RECT  130800.0 170550.0 132300.0 171450.0 ;
      RECT  53100.0 100050.0 130800.0 100950.0 ;
      RECT  53100.0 128250.0 130800.0 129150.0 ;
      RECT  53100.0 156450.0 130800.0 157350.0 ;
      RECT  53100.0 184650.0 130800.0 185550.0 ;
      RECT  119400.0 75450.0 135300.0 76350.0 ;
      RECT  119400.0 65250.0 138000.0 66150.0 ;
      RECT  119400.0 55050.0 140700.0 55950.0 ;
      RECT  119400.0 44850.0 143400.0 45750.0 ;
      RECT  119400.0 70350.0 149550.0 71250.0 ;
      RECT  119400.0 49950.0 149550.0 50850.0 ;
      RECT  115800.0 37650.0 116700.0 38550.0 ;
      RECT  115800.0 38100.0 116700.0 40200.0 ;
      RECT  53100.0 37650.0 116250.0 38550.0 ;
      RECT  164100.0 32400.0 175800.0 33300.0 ;
      RECT  158700.0 27900.0 175800.0 28800.0 ;
      RECT  161400.0 25500.0 175800.0 26400.0 ;
      RECT  164100.0 429600.0 175800.0 430500.0 ;
      RECT  166800.0 96900.0 175800.0 97800.0 ;
      RECT  169500.0 195000.0 175800.0 195900.0 ;
      RECT  61800.0 82650.0 62700.0 83550.0 ;
      RECT  61800.0 81000.0 62700.0 83100.0 ;
      RECT  62250.0 82650.0 156000.0 83550.0 ;
      RECT  103350.0 426450.0 156900.0 427350.0 ;
      RECT  175800.0 443700.0 198900.0 444600.0 ;
      RECT  175800.0 167700.0 198900.0 168600.0 ;
      RECT  175800.0 99000.0 198900.0 99900.0 ;
      RECT  175800.0 86400.0 198900.0 87300.0 ;
      RECT  175800.0 9600.0 198900.0 10500.0 ;
      RECT  152850.0 23400.0 175800.0 24300.0 ;
      RECT  152850.0 192900.0 175800.0 193800.0 ;
      RECT  152850.0 94800.0 175800.0 95700.0 ;
      RECT  175800.0 199200.0 186000.0 213300.0 ;
      RECT  175800.0 227400.0 186000.0 213300.0 ;
      RECT  175800.0 227400.0 186000.0 241500.0 ;
      RECT  175800.0 255600.0 186000.0 241500.0 ;
      RECT  175800.0 255600.0 186000.0 269700.0 ;
      RECT  175800.0 283800.0 186000.0 269700.0 ;
      RECT  175800.0 283800.0 186000.0 297900.0 ;
      RECT  175800.0 312000.0 186000.0 297900.0 ;
      RECT  175800.0 312000.0 186000.0 326100.0 ;
      RECT  175800.0 340200.0 186000.0 326100.0 ;
      RECT  175800.0 340200.0 186000.0 354300.0 ;
      RECT  175800.0 368400.0 186000.0 354300.0 ;
      RECT  175800.0 368400.0 186000.0 382500.0 ;
      RECT  175800.0 396600.0 186000.0 382500.0 ;
      RECT  175800.0 396600.0 186000.0 410700.0 ;
      RECT  175800.0 424800.0 186000.0 410700.0 ;
      RECT  186000.0 199200.0 196200.0 213300.0 ;
      RECT  186000.0 227400.0 196200.0 213300.0 ;
      RECT  186000.0 227400.0 196200.0 241500.0 ;
      RECT  186000.0 255600.0 196200.0 241500.0 ;
      RECT  186000.0 255600.0 196200.0 269700.0 ;
      RECT  186000.0 283800.0 196200.0 269700.0 ;
      RECT  186000.0 283800.0 196200.0 297900.0 ;
      RECT  186000.0 312000.0 196200.0 297900.0 ;
      RECT  186000.0 312000.0 196200.0 326100.0 ;
      RECT  186000.0 340200.0 196200.0 326100.0 ;
      RECT  186000.0 340200.0 196200.0 354300.0 ;
      RECT  186000.0 368400.0 196200.0 354300.0 ;
      RECT  186000.0 368400.0 196200.0 382500.0 ;
      RECT  186000.0 396600.0 196200.0 382500.0 ;
      RECT  186000.0 396600.0 196200.0 410700.0 ;
      RECT  186000.0 424800.0 196200.0 410700.0 ;
      RECT  175200.0 201300.0 196800.0 202500.0 ;
      RECT  175200.0 224100.0 196800.0 225300.0 ;
      RECT  175200.0 229500.0 196800.0 230700.0 ;
      RECT  175200.0 252300.0 196800.0 253500.0 ;
      RECT  175200.0 257700.0 196800.0 258900.0 ;
      RECT  175200.0 280500.0 196800.0 281700.0 ;
      RECT  175200.0 285900.0 196800.0 287100.0 ;
      RECT  175200.0 308700.0 196800.0 309900.0 ;
      RECT  175200.0 314100.0 196800.0 315300.0 ;
      RECT  175200.0 336900.0 196800.0 338100.0 ;
      RECT  175200.0 342300.0 196800.0 343500.0 ;
      RECT  175200.0 365100.0 196800.0 366300.0 ;
      RECT  175200.0 370500.0 196800.0 371700.0 ;
      RECT  175200.0 393300.0 196800.0 394500.0 ;
      RECT  175200.0 398700.0 196800.0 399900.0 ;
      RECT  175200.0 421500.0 196800.0 422700.0 ;
      RECT  175200.0 212700.0 196800.0 213600.0 ;
      RECT  175200.0 240900.0 196800.0 241800.0 ;
      RECT  175200.0 269100.0 196800.0 270000.0 ;
      RECT  175200.0 297300.0 196800.0 298200.0 ;
      RECT  175200.0 325500.0 196800.0 326400.0 ;
      RECT  175200.0 353700.0 196800.0 354600.0 ;
      RECT  175200.0 381900.0 196800.0 382800.0 ;
      RECT  175200.0 410100.0 196800.0 411000.0 ;
      RECT  181200.0 436200.0 182400.0 444600.0 ;
      RECT  178800.0 427200.0 180000.0 428400.0 ;
      RECT  181200.0 427200.0 182400.0 428400.0 ;
      RECT  181200.0 427200.0 182400.0 428400.0 ;
      RECT  178800.0 427200.0 180000.0 428400.0 ;
      RECT  178800.0 436200.0 180000.0 437400.0 ;
      RECT  181200.0 436200.0 182400.0 437400.0 ;
      RECT  181200.0 436200.0 182400.0 437400.0 ;
      RECT  178800.0 436200.0 180000.0 437400.0 ;
      RECT  181200.0 436200.0 182400.0 437400.0 ;
      RECT  183600.0 436200.0 184800.0 437400.0 ;
      RECT  183600.0 436200.0 184800.0 437400.0 ;
      RECT  181200.0 436200.0 182400.0 437400.0 ;
      RECT  180900.0 429450.0 179700.0 430650.0 ;
      RECT  181200.0 442800.0 182400.0 444000.0 ;
      RECT  178800.0 427200.0 180000.0 428400.0 ;
      RECT  181200.0 427200.0 182400.0 428400.0 ;
      RECT  178800.0 436200.0 180000.0 437400.0 ;
      RECT  183600.0 436200.0 184800.0 437400.0 ;
      RECT  178800.0 427200.0 180000.0 428400.0 ;
      RECT  181200.0 427200.0 182400.0 428400.0 ;
      RECT  178800.0 436200.0 180000.0 437400.0 ;
      RECT  183600.0 436200.0 184800.0 437400.0 ;
      RECT  175800.0 429600.0 186000.0 430500.0 ;
      RECT  175800.0 443700.0 186000.0 444600.0 ;
      RECT  191400.0 436200.0 192600.0 444600.0 ;
      RECT  189000.0 427200.0 190200.0 428400.0 ;
      RECT  191400.0 427200.0 192600.0 428400.0 ;
      RECT  191400.0 427200.0 192600.0 428400.0 ;
      RECT  189000.0 427200.0 190200.0 428400.0 ;
      RECT  189000.0 436200.0 190200.0 437400.0 ;
      RECT  191400.0 436200.0 192600.0 437400.0 ;
      RECT  191400.0 436200.0 192600.0 437400.0 ;
      RECT  189000.0 436200.0 190200.0 437400.0 ;
      RECT  191400.0 436200.0 192600.0 437400.0 ;
      RECT  193800.0 436200.0 195000.0 437400.0 ;
      RECT  193800.0 436200.0 195000.0 437400.0 ;
      RECT  191400.0 436200.0 192600.0 437400.0 ;
      RECT  191100.0 429450.0 189900.0 430650.0 ;
      RECT  191400.0 442800.0 192600.0 444000.0 ;
      RECT  189000.0 427200.0 190200.0 428400.0 ;
      RECT  191400.0 427200.0 192600.0 428400.0 ;
      RECT  189000.0 436200.0 190200.0 437400.0 ;
      RECT  193800.0 436200.0 195000.0 437400.0 ;
      RECT  189000.0 427200.0 190200.0 428400.0 ;
      RECT  191400.0 427200.0 192600.0 428400.0 ;
      RECT  189000.0 436200.0 190200.0 437400.0 ;
      RECT  193800.0 436200.0 195000.0 437400.0 ;
      RECT  186000.0 429600.0 196200.0 430500.0 ;
      RECT  186000.0 443700.0 196200.0 444600.0 ;
      RECT  175800.0 429600.0 196200.0 430500.0 ;
      RECT  175800.0 443700.0 196200.0 444600.0 ;
      RECT  175800.0 150300.0 186000.0 199200.0 ;
      RECT  186000.0 150300.0 196200.0 199200.0 ;
      RECT  175800.0 195000.0 196200.0 195900.0 ;
      RECT  175800.0 167700.0 196200.0 168600.0 ;
      RECT  175800.0 192900.0 196200.0 193800.0 ;
      RECT  175800.0 90000.0 186000.0 150300.0 ;
      RECT  186000.0 90000.0 196200.0 150300.0 ;
      RECT  175800.0 96900.0 196200.0 97800.0 ;
      RECT  175800.0 99000.0 196200.0 99900.0 ;
      RECT  175800.0 94800.0 196200.0 95700.0 ;
      RECT  175800.0 30000.0 186000.0 90000.0 ;
      RECT  196200.0 30000.0 186000.0 90000.0 ;
      RECT  175800.0 32400.0 196200.0 33300.0 ;
      RECT  175800.0 86400.0 196200.0 87300.0 ;
      RECT  175800.0 30000.0 186000.0 8100.0 ;
      RECT  186000.0 30000.0 196200.0 8100.0 ;
      RECT  175800.0 26400.0 196200.0 25500.0 ;
      RECT  175800.0 28800.0 196200.0 27900.0 ;
      RECT  175800.0 10500.0 196200.0 9600.0 ;
      RECT  175800.0 24300.0 196200.0 23400.0 ;
      RECT  88050.0 206550.0 88950.0 207450.0 ;
      RECT  88050.0 205200.0 88950.0 206100.0 ;
      RECT  84000.0 206550.0 88500.0 207450.0 ;
      RECT  88050.0 205650.0 88950.0 207000.0 ;
      RECT  88500.0 205200.0 93000.0 206100.0 ;
      RECT  88050.0 219150.0 88950.0 220050.0 ;
      RECT  88050.0 220500.0 88950.0 221400.0 ;
      RECT  84000.0 219150.0 88500.0 220050.0 ;
      RECT  88050.0 219600.0 88950.0 220950.0 ;
      RECT  88500.0 220500.0 93000.0 221400.0 ;
      RECT  88050.0 234750.0 88950.0 235650.0 ;
      RECT  88050.0 233400.0 88950.0 234300.0 ;
      RECT  84000.0 234750.0 88500.0 235650.0 ;
      RECT  88050.0 233850.0 88950.0 235200.0 ;
      RECT  88500.0 233400.0 93000.0 234300.0 ;
      RECT  88050.0 247350.0 88950.0 248250.0 ;
      RECT  88050.0 248700.0 88950.0 249600.0 ;
      RECT  84000.0 247350.0 88500.0 248250.0 ;
      RECT  88050.0 247800.0 88950.0 249150.0 ;
      RECT  88500.0 248700.0 93000.0 249600.0 ;
      RECT  88050.0 262950.0 88950.0 263850.0 ;
      RECT  88050.0 261600.0 88950.0 262500.0 ;
      RECT  84000.0 262950.0 88500.0 263850.0 ;
      RECT  88050.0 262050.0 88950.0 263400.0 ;
      RECT  88500.0 261600.0 93000.0 262500.0 ;
      RECT  88050.0 275550.0 88950.0 276450.0 ;
      RECT  88050.0 276900.0 88950.0 277800.0 ;
      RECT  84000.0 275550.0 88500.0 276450.0 ;
      RECT  88050.0 276000.0 88950.0 277350.0 ;
      RECT  88500.0 276900.0 93000.0 277800.0 ;
      RECT  88050.0 291150.0 88950.0 292050.0 ;
      RECT  88050.0 289800.0 88950.0 290700.0 ;
      RECT  84000.0 291150.0 88500.0 292050.0 ;
      RECT  88050.0 290250.0 88950.0 291600.0 ;
      RECT  88500.0 289800.0 93000.0 290700.0 ;
      RECT  88050.0 303750.0 88950.0 304650.0 ;
      RECT  88050.0 305100.0 88950.0 306000.0 ;
      RECT  84000.0 303750.0 88500.0 304650.0 ;
      RECT  88050.0 304200.0 88950.0 305550.0 ;
      RECT  88500.0 305100.0 93000.0 306000.0 ;
      RECT  88050.0 319350.0 88950.0 320250.0 ;
      RECT  88050.0 318000.0 88950.0 318900.0 ;
      RECT  84000.0 319350.0 88500.0 320250.0 ;
      RECT  88050.0 318450.0 88950.0 319800.0 ;
      RECT  88500.0 318000.0 93000.0 318900.0 ;
      RECT  88050.0 331950.0 88950.0 332850.0 ;
      RECT  88050.0 333300.0 88950.0 334200.0 ;
      RECT  84000.0 331950.0 88500.0 332850.0 ;
      RECT  88050.0 332400.0 88950.0 333750.0 ;
      RECT  88500.0 333300.0 93000.0 334200.0 ;
      RECT  88050.0 347550.0 88950.0 348450.0 ;
      RECT  88050.0 346200.0 88950.0 347100.0 ;
      RECT  84000.0 347550.0 88500.0 348450.0 ;
      RECT  88050.0 346650.0 88950.0 348000.0 ;
      RECT  88500.0 346200.0 93000.0 347100.0 ;
      RECT  88050.0 360150.0 88950.0 361050.0 ;
      RECT  88050.0 361500.0 88950.0 362400.0 ;
      RECT  84000.0 360150.0 88500.0 361050.0 ;
      RECT  88050.0 360600.0 88950.0 361950.0 ;
      RECT  88500.0 361500.0 93000.0 362400.0 ;
      RECT  88050.0 375750.0 88950.0 376650.0 ;
      RECT  88050.0 374400.0 88950.0 375300.0 ;
      RECT  84000.0 375750.0 88500.0 376650.0 ;
      RECT  88050.0 374850.0 88950.0 376200.0 ;
      RECT  88500.0 374400.0 93000.0 375300.0 ;
      RECT  88050.0 388350.0 88950.0 389250.0 ;
      RECT  88050.0 389700.0 88950.0 390600.0 ;
      RECT  84000.0 388350.0 88500.0 389250.0 ;
      RECT  88050.0 388800.0 88950.0 390150.0 ;
      RECT  88500.0 389700.0 93000.0 390600.0 ;
      RECT  88050.0 403950.0 88950.0 404850.0 ;
      RECT  88050.0 402600.0 88950.0 403500.0 ;
      RECT  84000.0 403950.0 88500.0 404850.0 ;
      RECT  88050.0 403050.0 88950.0 404400.0 ;
      RECT  88500.0 402600.0 93000.0 403500.0 ;
      RECT  88050.0 416550.0 88950.0 417450.0 ;
      RECT  88050.0 417900.0 88950.0 418800.0 ;
      RECT  84000.0 416550.0 88500.0 417450.0 ;
      RECT  88050.0 417000.0 88950.0 418350.0 ;
      RECT  88500.0 417900.0 93000.0 418800.0 ;
      RECT  59850.0 92400.0 76200.0 93300.0 ;
      RECT  61950.0 107700.0 76200.0 108600.0 ;
      RECT  64050.0 120600.0 76200.0 121500.0 ;
      RECT  66150.0 135900.0 76200.0 136800.0 ;
      RECT  68250.0 148800.0 76200.0 149700.0 ;
      RECT  70350.0 164100.0 76200.0 165000.0 ;
      RECT  72450.0 177000.0 76200.0 177900.0 ;
      RECT  74550.0 192300.0 76200.0 193200.0 ;
      RECT  59850.0 206550.0 78600.0 207450.0 ;
      RECT  68250.0 203850.0 81600.0 204750.0 ;
      RECT  59850.0 219150.0 78600.0 220050.0 ;
      RECT  70350.0 221850.0 81600.0 222750.0 ;
      RECT  59850.0 234750.0 78600.0 235650.0 ;
      RECT  72450.0 232050.0 81600.0 232950.0 ;
      RECT  59850.0 247350.0 78600.0 248250.0 ;
      RECT  74550.0 250050.0 81600.0 250950.0 ;
      RECT  61950.0 262950.0 78600.0 263850.0 ;
      RECT  68250.0 260250.0 81600.0 261150.0 ;
      RECT  61950.0 275550.0 78600.0 276450.0 ;
      RECT  70350.0 278250.0 81600.0 279150.0 ;
      RECT  61950.0 291150.0 78600.0 292050.0 ;
      RECT  72450.0 288450.0 81600.0 289350.0 ;
      RECT  61950.0 303750.0 78600.0 304650.0 ;
      RECT  74550.0 306450.0 81600.0 307350.0 ;
      RECT  64050.0 319350.0 78600.0 320250.0 ;
      RECT  68250.0 316650.0 81600.0 317550.0 ;
      RECT  64050.0 331950.0 78600.0 332850.0 ;
      RECT  70350.0 334650.0 81600.0 335550.0 ;
      RECT  64050.0 347550.0 78600.0 348450.0 ;
      RECT  72450.0 344850.0 81600.0 345750.0 ;
      RECT  64050.0 360150.0 78600.0 361050.0 ;
      RECT  74550.0 362850.0 81600.0 363750.0 ;
      RECT  66150.0 375750.0 78600.0 376650.0 ;
      RECT  68250.0 373050.0 81600.0 373950.0 ;
      RECT  66150.0 388350.0 78600.0 389250.0 ;
      RECT  70350.0 391050.0 81600.0 391950.0 ;
      RECT  66150.0 403950.0 78600.0 404850.0 ;
      RECT  72450.0 401250.0 81600.0 402150.0 ;
      RECT  66150.0 416550.0 78600.0 417450.0 ;
      RECT  74550.0 419250.0 81600.0 420150.0 ;
      RECT  114750.0 92400.0 113850.0 93300.0 ;
      RECT  114750.0 97350.0 113850.0 98250.0 ;
      RECT  118950.0 92400.0 114300.0 93300.0 ;
      RECT  114750.0 92850.0 113850.0 97800.0 ;
      RECT  114300.0 97350.0 111750.0 98250.0 ;
      RECT  130350.0 92400.0 122400.0 93300.0 ;
      RECT  114750.0 107700.0 113850.0 108600.0 ;
      RECT  114750.0 111450.0 113850.0 112350.0 ;
      RECT  118950.0 107700.0 114300.0 108600.0 ;
      RECT  114750.0 108150.0 113850.0 111900.0 ;
      RECT  114300.0 111450.0 108750.0 112350.0 ;
      RECT  127350.0 107700.0 122400.0 108600.0 ;
      RECT  130350.0 116250.0 105750.0 117150.0 ;
      RECT  127350.0 130350.0 102750.0 131250.0 ;
      RECT  111750.0 93750.0 97800.0 94650.0 ;
      RECT  108750.0 91050.0 94800.0 91950.0 ;
      RECT  105750.0 106350.0 97800.0 107250.0 ;
      RECT  108750.0 109050.0 94800.0 109950.0 ;
      RECT  111750.0 121950.0 97800.0 122850.0 ;
      RECT  102750.0 119250.0 94800.0 120150.0 ;
      RECT  105750.0 134550.0 97800.0 135450.0 ;
      RECT  102750.0 137250.0 94800.0 138150.0 ;
      RECT  88350.0 93750.0 87450.0 94650.0 ;
      RECT  88350.0 92400.0 87450.0 93300.0 ;
      RECT  92400.0 93750.0 87900.0 94650.0 ;
      RECT  88350.0 92850.0 87450.0 94200.0 ;
      RECT  87900.0 92400.0 83400.0 93300.0 ;
      RECT  88350.0 106350.0 87450.0 107250.0 ;
      RECT  88350.0 107700.0 87450.0 108600.0 ;
      RECT  92400.0 106350.0 87900.0 107250.0 ;
      RECT  88350.0 106800.0 87450.0 108150.0 ;
      RECT  87900.0 107700.0 83400.0 108600.0 ;
      RECT  88350.0 121950.0 87450.0 122850.0 ;
      RECT  88350.0 120600.0 87450.0 121500.0 ;
      RECT  92400.0 121950.0 87900.0 122850.0 ;
      RECT  88350.0 121050.0 87450.0 122400.0 ;
      RECT  87900.0 120600.0 83400.0 121500.0 ;
      RECT  88350.0 134550.0 87450.0 135450.0 ;
      RECT  88350.0 135900.0 87450.0 136800.0 ;
      RECT  92400.0 134550.0 87900.0 135450.0 ;
      RECT  88350.0 135000.0 87450.0 136350.0 ;
      RECT  87900.0 135900.0 83400.0 136800.0 ;
      RECT  118200.0 86400.0 117000.0 88350.0 ;
      RECT  118200.0 98550.0 117000.0 100500.0 ;
      RECT  123000.0 87750.0 121800.0 85950.0 ;
      RECT  123000.0 97350.0 121800.0 100950.0 ;
      RECT  120300.0 88950.0 119400.0 97350.0 ;
      RECT  123000.0 97350.0 121800.0 98550.0 ;
      RECT  120600.0 97350.0 119400.0 98550.0 ;
      RECT  120600.0 97350.0 119400.0 98550.0 ;
      RECT  123000.0 97350.0 121800.0 98550.0 ;
      RECT  123000.0 87750.0 121800.0 88950.0 ;
      RECT  120600.0 87750.0 119400.0 88950.0 ;
      RECT  120600.0 87750.0 119400.0 88950.0 ;
      RECT  123000.0 87750.0 121800.0 88950.0 ;
      RECT  118200.0 87750.0 117000.0 88950.0 ;
      RECT  118200.0 97950.0 117000.0 99150.0 ;
      RECT  122400.0 92250.0 121200.0 93450.0 ;
      RECT  122400.0 92250.0 121200.0 93450.0 ;
      RECT  119850.0 92400.0 118950.0 93300.0 ;
      RECT  124800.0 100050.0 115200.0 100950.0 ;
      RECT  124800.0 85950.0 115200.0 86850.0 ;
      RECT  118200.0 114600.0 117000.0 112650.0 ;
      RECT  118200.0 102450.0 117000.0 100500.0 ;
      RECT  123000.0 113250.0 121800.0 115050.0 ;
      RECT  123000.0 103650.0 121800.0 100050.0 ;
      RECT  120300.0 112050.0 119400.0 103650.0 ;
      RECT  123000.0 103650.0 121800.0 102450.0 ;
      RECT  120600.0 103650.0 119400.0 102450.0 ;
      RECT  120600.0 103650.0 119400.0 102450.0 ;
      RECT  123000.0 103650.0 121800.0 102450.0 ;
      RECT  123000.0 113250.0 121800.0 112050.0 ;
      RECT  120600.0 113250.0 119400.0 112050.0 ;
      RECT  120600.0 113250.0 119400.0 112050.0 ;
      RECT  123000.0 113250.0 121800.0 112050.0 ;
      RECT  118200.0 113250.0 117000.0 112050.0 ;
      RECT  118200.0 103050.0 117000.0 101850.0 ;
      RECT  122400.0 108750.0 121200.0 107550.0 ;
      RECT  122400.0 108750.0 121200.0 107550.0 ;
      RECT  119850.0 108600.0 118950.0 107700.0 ;
      RECT  124800.0 100950.0 115200.0 100050.0 ;
      RECT  124800.0 115050.0 115200.0 114150.0 ;
      RECT  79200.0 86400.0 78000.0 88350.0 ;
      RECT  79200.0 98550.0 78000.0 100500.0 ;
      RECT  84000.0 87750.0 82800.0 85950.0 ;
      RECT  84000.0 97350.0 82800.0 100950.0 ;
      RECT  81300.0 88950.0 80400.0 97350.0 ;
      RECT  84000.0 97350.0 82800.0 98550.0 ;
      RECT  81600.0 97350.0 80400.0 98550.0 ;
      RECT  81600.0 97350.0 80400.0 98550.0 ;
      RECT  84000.0 97350.0 82800.0 98550.0 ;
      RECT  84000.0 87750.0 82800.0 88950.0 ;
      RECT  81600.0 87750.0 80400.0 88950.0 ;
      RECT  81600.0 87750.0 80400.0 88950.0 ;
      RECT  84000.0 87750.0 82800.0 88950.0 ;
      RECT  79200.0 87750.0 78000.0 88950.0 ;
      RECT  79200.0 97950.0 78000.0 99150.0 ;
      RECT  83400.0 92250.0 82200.0 93450.0 ;
      RECT  83400.0 92250.0 82200.0 93450.0 ;
      RECT  80850.0 92400.0 79950.0 93300.0 ;
      RECT  85800.0 100050.0 76200.0 100950.0 ;
      RECT  85800.0 85950.0 76200.0 86850.0 ;
      RECT  79200.0 114600.0 78000.0 112650.0 ;
      RECT  79200.0 102450.0 78000.0 100500.0 ;
      RECT  84000.0 113250.0 82800.0 115050.0 ;
      RECT  84000.0 103650.0 82800.0 100050.0 ;
      RECT  81300.0 112050.0 80400.0 103650.0 ;
      RECT  84000.0 103650.0 82800.0 102450.0 ;
      RECT  81600.0 103650.0 80400.0 102450.0 ;
      RECT  81600.0 103650.0 80400.0 102450.0 ;
      RECT  84000.0 103650.0 82800.0 102450.0 ;
      RECT  84000.0 113250.0 82800.0 112050.0 ;
      RECT  81600.0 113250.0 80400.0 112050.0 ;
      RECT  81600.0 113250.0 80400.0 112050.0 ;
      RECT  84000.0 113250.0 82800.0 112050.0 ;
      RECT  79200.0 113250.0 78000.0 112050.0 ;
      RECT  79200.0 103050.0 78000.0 101850.0 ;
      RECT  83400.0 108750.0 82200.0 107550.0 ;
      RECT  83400.0 108750.0 82200.0 107550.0 ;
      RECT  80850.0 108600.0 79950.0 107700.0 ;
      RECT  85800.0 100950.0 76200.0 100050.0 ;
      RECT  85800.0 115050.0 76200.0 114150.0 ;
      RECT  79200.0 114600.0 78000.0 116550.0 ;
      RECT  79200.0 126750.0 78000.0 128700.0 ;
      RECT  84000.0 115950.0 82800.0 114150.0 ;
      RECT  84000.0 125550.0 82800.0 129150.0 ;
      RECT  81300.0 117150.0 80400.0 125550.0 ;
      RECT  84000.0 125550.0 82800.0 126750.0 ;
      RECT  81600.0 125550.0 80400.0 126750.0 ;
      RECT  81600.0 125550.0 80400.0 126750.0 ;
      RECT  84000.0 125550.0 82800.0 126750.0 ;
      RECT  84000.0 115950.0 82800.0 117150.0 ;
      RECT  81600.0 115950.0 80400.0 117150.0 ;
      RECT  81600.0 115950.0 80400.0 117150.0 ;
      RECT  84000.0 115950.0 82800.0 117150.0 ;
      RECT  79200.0 115950.0 78000.0 117150.0 ;
      RECT  79200.0 126150.0 78000.0 127350.0 ;
      RECT  83400.0 120450.0 82200.0 121650.0 ;
      RECT  83400.0 120450.0 82200.0 121650.0 ;
      RECT  80850.0 120600.0 79950.0 121500.0 ;
      RECT  85800.0 128250.0 76200.0 129150.0 ;
      RECT  85800.0 114150.0 76200.0 115050.0 ;
      RECT  79200.0 142800.0 78000.0 140850.0 ;
      RECT  79200.0 130650.0 78000.0 128700.0 ;
      RECT  84000.0 141450.0 82800.0 143250.0 ;
      RECT  84000.0 131850.0 82800.0 128250.0 ;
      RECT  81300.0 140250.0 80400.0 131850.0 ;
      RECT  84000.0 131850.0 82800.0 130650.0 ;
      RECT  81600.0 131850.0 80400.0 130650.0 ;
      RECT  81600.0 131850.0 80400.0 130650.0 ;
      RECT  84000.0 131850.0 82800.0 130650.0 ;
      RECT  84000.0 141450.0 82800.0 140250.0 ;
      RECT  81600.0 141450.0 80400.0 140250.0 ;
      RECT  81600.0 141450.0 80400.0 140250.0 ;
      RECT  84000.0 141450.0 82800.0 140250.0 ;
      RECT  79200.0 141450.0 78000.0 140250.0 ;
      RECT  79200.0 131250.0 78000.0 130050.0 ;
      RECT  83400.0 136950.0 82200.0 135750.0 ;
      RECT  83400.0 136950.0 82200.0 135750.0 ;
      RECT  80850.0 136800.0 79950.0 135900.0 ;
      RECT  85800.0 129150.0 76200.0 128250.0 ;
      RECT  85800.0 143250.0 76200.0 142350.0 ;
      RECT  91200.0 86400.0 90000.0 88350.0 ;
      RECT  91200.0 98550.0 90000.0 100500.0 ;
      RECT  98400.0 88350.0 97200.0 85950.0 ;
      RECT  98400.0 97350.0 97200.0 100950.0 ;
      RECT  93600.0 97350.0 92400.0 100950.0 ;
      RECT  98400.0 97350.0 97200.0 98550.0 ;
      RECT  96000.0 97350.0 94800.0 98550.0 ;
      RECT  96000.0 97350.0 94800.0 98550.0 ;
      RECT  98400.0 97350.0 97200.0 98550.0 ;
      RECT  96000.0 97350.0 94800.0 98550.0 ;
      RECT  93600.0 97350.0 92400.0 98550.0 ;
      RECT  93600.0 97350.0 92400.0 98550.0 ;
      RECT  96000.0 97350.0 94800.0 98550.0 ;
      RECT  98400.0 88350.0 97200.0 89550.0 ;
      RECT  96000.0 88350.0 94800.0 89550.0 ;
      RECT  96000.0 88350.0 94800.0 89550.0 ;
      RECT  98400.0 88350.0 97200.0 89550.0 ;
      RECT  96000.0 88350.0 94800.0 89550.0 ;
      RECT  93600.0 88350.0 92400.0 89550.0 ;
      RECT  93600.0 88350.0 92400.0 89550.0 ;
      RECT  96000.0 88350.0 94800.0 89550.0 ;
      RECT  91200.0 87750.0 90000.0 88950.0 ;
      RECT  91200.0 97950.0 90000.0 99150.0 ;
      RECT  93600.0 90900.0 94800.0 92100.0 ;
      RECT  96600.0 93600.0 97800.0 94800.0 ;
      RECT  96000.0 97350.0 94800.0 98550.0 ;
      RECT  93600.0 88350.0 92400.0 89550.0 ;
      RECT  92400.0 93600.0 93600.0 94800.0 ;
      RECT  97800.0 93600.0 96600.0 94800.0 ;
      RECT  94800.0 90900.0 93600.0 92100.0 ;
      RECT  93600.0 93600.0 92400.0 94800.0 ;
      RECT  100200.0 100050.0 85800.0 100950.0 ;
      RECT  100200.0 85950.0 85800.0 86850.0 ;
      RECT  91200.0 114600.0 90000.0 112650.0 ;
      RECT  91200.0 102450.0 90000.0 100500.0 ;
      RECT  98400.0 112650.0 97200.0 115050.0 ;
      RECT  98400.0 103650.0 97200.0 100050.0 ;
      RECT  93600.0 103650.0 92400.0 100050.0 ;
      RECT  98400.0 103650.0 97200.0 102450.0 ;
      RECT  96000.0 103650.0 94800.0 102450.0 ;
      RECT  96000.0 103650.0 94800.0 102450.0 ;
      RECT  98400.0 103650.0 97200.0 102450.0 ;
      RECT  96000.0 103650.0 94800.0 102450.0 ;
      RECT  93600.0 103650.0 92400.0 102450.0 ;
      RECT  93600.0 103650.0 92400.0 102450.0 ;
      RECT  96000.0 103650.0 94800.0 102450.0 ;
      RECT  98400.0 112650.0 97200.0 111450.0 ;
      RECT  96000.0 112650.0 94800.0 111450.0 ;
      RECT  96000.0 112650.0 94800.0 111450.0 ;
      RECT  98400.0 112650.0 97200.0 111450.0 ;
      RECT  96000.0 112650.0 94800.0 111450.0 ;
      RECT  93600.0 112650.0 92400.0 111450.0 ;
      RECT  93600.0 112650.0 92400.0 111450.0 ;
      RECT  96000.0 112650.0 94800.0 111450.0 ;
      RECT  91200.0 113250.0 90000.0 112050.0 ;
      RECT  91200.0 103050.0 90000.0 101850.0 ;
      RECT  93600.0 110100.0 94800.0 108900.0 ;
      RECT  96600.0 107400.0 97800.0 106200.0 ;
      RECT  96000.0 103650.0 94800.0 102450.0 ;
      RECT  93600.0 112650.0 92400.0 111450.0 ;
      RECT  92400.0 107400.0 93600.0 106200.0 ;
      RECT  97800.0 107400.0 96600.0 106200.0 ;
      RECT  94800.0 110100.0 93600.0 108900.0 ;
      RECT  93600.0 107400.0 92400.0 106200.0 ;
      RECT  100200.0 100950.0 85800.0 100050.0 ;
      RECT  100200.0 115050.0 85800.0 114150.0 ;
      RECT  91200.0 114600.0 90000.0 116550.0 ;
      RECT  91200.0 126750.0 90000.0 128700.0 ;
      RECT  98400.0 116550.0 97200.0 114150.0 ;
      RECT  98400.0 125550.0 97200.0 129150.0 ;
      RECT  93600.0 125550.0 92400.0 129150.0 ;
      RECT  98400.0 125550.0 97200.0 126750.0 ;
      RECT  96000.0 125550.0 94800.0 126750.0 ;
      RECT  96000.0 125550.0 94800.0 126750.0 ;
      RECT  98400.0 125550.0 97200.0 126750.0 ;
      RECT  96000.0 125550.0 94800.0 126750.0 ;
      RECT  93600.0 125550.0 92400.0 126750.0 ;
      RECT  93600.0 125550.0 92400.0 126750.0 ;
      RECT  96000.0 125550.0 94800.0 126750.0 ;
      RECT  98400.0 116550.0 97200.0 117750.0 ;
      RECT  96000.0 116550.0 94800.0 117750.0 ;
      RECT  96000.0 116550.0 94800.0 117750.0 ;
      RECT  98400.0 116550.0 97200.0 117750.0 ;
      RECT  96000.0 116550.0 94800.0 117750.0 ;
      RECT  93600.0 116550.0 92400.0 117750.0 ;
      RECT  93600.0 116550.0 92400.0 117750.0 ;
      RECT  96000.0 116550.0 94800.0 117750.0 ;
      RECT  91200.0 115950.0 90000.0 117150.0 ;
      RECT  91200.0 126150.0 90000.0 127350.0 ;
      RECT  93600.0 119100.0 94800.0 120300.0 ;
      RECT  96600.0 121800.0 97800.0 123000.0 ;
      RECT  96000.0 125550.0 94800.0 126750.0 ;
      RECT  93600.0 116550.0 92400.0 117750.0 ;
      RECT  92400.0 121800.0 93600.0 123000.0 ;
      RECT  97800.0 121800.0 96600.0 123000.0 ;
      RECT  94800.0 119100.0 93600.0 120300.0 ;
      RECT  93600.0 121800.0 92400.0 123000.0 ;
      RECT  100200.0 128250.0 85800.0 129150.0 ;
      RECT  100200.0 114150.0 85800.0 115050.0 ;
      RECT  91200.0 142800.0 90000.0 140850.0 ;
      RECT  91200.0 130650.0 90000.0 128700.0 ;
      RECT  98400.0 140850.0 97200.0 143250.0 ;
      RECT  98400.0 131850.0 97200.0 128250.0 ;
      RECT  93600.0 131850.0 92400.0 128250.0 ;
      RECT  98400.0 131850.0 97200.0 130650.0 ;
      RECT  96000.0 131850.0 94800.0 130650.0 ;
      RECT  96000.0 131850.0 94800.0 130650.0 ;
      RECT  98400.0 131850.0 97200.0 130650.0 ;
      RECT  96000.0 131850.0 94800.0 130650.0 ;
      RECT  93600.0 131850.0 92400.0 130650.0 ;
      RECT  93600.0 131850.0 92400.0 130650.0 ;
      RECT  96000.0 131850.0 94800.0 130650.0 ;
      RECT  98400.0 140850.0 97200.0 139650.0 ;
      RECT  96000.0 140850.0 94800.0 139650.0 ;
      RECT  96000.0 140850.0 94800.0 139650.0 ;
      RECT  98400.0 140850.0 97200.0 139650.0 ;
      RECT  96000.0 140850.0 94800.0 139650.0 ;
      RECT  93600.0 140850.0 92400.0 139650.0 ;
      RECT  93600.0 140850.0 92400.0 139650.0 ;
      RECT  96000.0 140850.0 94800.0 139650.0 ;
      RECT  91200.0 141450.0 90000.0 140250.0 ;
      RECT  91200.0 131250.0 90000.0 130050.0 ;
      RECT  93600.0 138300.0 94800.0 137100.0 ;
      RECT  96600.0 135600.0 97800.0 134400.0 ;
      RECT  96000.0 131850.0 94800.0 130650.0 ;
      RECT  93600.0 140850.0 92400.0 139650.0 ;
      RECT  92400.0 135600.0 93600.0 134400.0 ;
      RECT  97800.0 135600.0 96600.0 134400.0 ;
      RECT  94800.0 138300.0 93600.0 137100.0 ;
      RECT  93600.0 135600.0 92400.0 134400.0 ;
      RECT  100200.0 129150.0 85800.0 128250.0 ;
      RECT  100200.0 143250.0 85800.0 142350.0 ;
      RECT  111150.0 97200.0 112350.0 98400.0 ;
      RECT  129750.0 92250.0 130950.0 93450.0 ;
      RECT  108150.0 111300.0 109350.0 112500.0 ;
      RECT  126750.0 107550.0 127950.0 108750.0 ;
      RECT  129750.0 116100.0 130950.0 117300.0 ;
      RECT  105150.0 116100.0 106350.0 117300.0 ;
      RECT  126750.0 130200.0 127950.0 131400.0 ;
      RECT  102150.0 130200.0 103350.0 131400.0 ;
      RECT  111150.0 93600.0 112350.0 94800.0 ;
      RECT  108150.0 90900.0 109350.0 92100.0 ;
      RECT  105150.0 106200.0 106350.0 107400.0 ;
      RECT  108150.0 108900.0 109350.0 110100.0 ;
      RECT  111150.0 121800.0 112350.0 123000.0 ;
      RECT  102150.0 119100.0 103350.0 120300.0 ;
      RECT  105150.0 134400.0 106350.0 135600.0 ;
      RECT  102150.0 137100.0 103350.0 138300.0 ;
      RECT  79950.0 92400.0 76200.0 93300.0 ;
      RECT  79950.0 107700.0 76200.0 108600.0 ;
      RECT  79950.0 120600.0 76200.0 121500.0 ;
      RECT  79950.0 135900.0 76200.0 136800.0 ;
      RECT  130800.0 100050.0 76200.0 100950.0 ;
      RECT  130800.0 128250.0 76200.0 129150.0 ;
      RECT  130800.0 85950.0 76200.0 86850.0 ;
      RECT  130800.0 114150.0 76200.0 115050.0 ;
      RECT  130800.0 142350.0 76200.0 143250.0 ;
      RECT  114750.0 148800.0 113850.0 149700.0 ;
      RECT  114750.0 153750.0 113850.0 154650.0 ;
      RECT  118950.0 148800.0 114300.0 149700.0 ;
      RECT  114750.0 149250.0 113850.0 154200.0 ;
      RECT  114300.0 153750.0 111750.0 154650.0 ;
      RECT  130350.0 148800.0 122400.0 149700.0 ;
      RECT  114750.0 164100.0 113850.0 165000.0 ;
      RECT  114750.0 167850.0 113850.0 168750.0 ;
      RECT  118950.0 164100.0 114300.0 165000.0 ;
      RECT  114750.0 164550.0 113850.0 168300.0 ;
      RECT  114300.0 167850.0 108750.0 168750.0 ;
      RECT  127350.0 164100.0 122400.0 165000.0 ;
      RECT  130350.0 172650.0 105750.0 173550.0 ;
      RECT  127350.0 186750.0 102750.0 187650.0 ;
      RECT  111750.0 150150.0 97800.0 151050.0 ;
      RECT  108750.0 147450.0 94800.0 148350.0 ;
      RECT  105750.0 162750.0 97800.0 163650.0 ;
      RECT  108750.0 165450.0 94800.0 166350.0 ;
      RECT  111750.0 178350.0 97800.0 179250.0 ;
      RECT  102750.0 175650.0 94800.0 176550.0 ;
      RECT  105750.0 190950.0 97800.0 191850.0 ;
      RECT  102750.0 193650.0 94800.0 194550.0 ;
      RECT  88350.0 150150.0 87450.0 151050.0 ;
      RECT  88350.0 148800.0 87450.0 149700.0 ;
      RECT  92400.0 150150.0 87900.0 151050.0 ;
      RECT  88350.0 149250.0 87450.0 150600.0 ;
      RECT  87900.0 148800.0 83400.0 149700.0 ;
      RECT  88350.0 162750.0 87450.0 163650.0 ;
      RECT  88350.0 164100.0 87450.0 165000.0 ;
      RECT  92400.0 162750.0 87900.0 163650.0 ;
      RECT  88350.0 163200.0 87450.0 164550.0 ;
      RECT  87900.0 164100.0 83400.0 165000.0 ;
      RECT  88350.0 178350.0 87450.0 179250.0 ;
      RECT  88350.0 177000.0 87450.0 177900.0 ;
      RECT  92400.0 178350.0 87900.0 179250.0 ;
      RECT  88350.0 177450.0 87450.0 178800.0 ;
      RECT  87900.0 177000.0 83400.0 177900.0 ;
      RECT  88350.0 190950.0 87450.0 191850.0 ;
      RECT  88350.0 192300.0 87450.0 193200.0 ;
      RECT  92400.0 190950.0 87900.0 191850.0 ;
      RECT  88350.0 191400.0 87450.0 192750.0 ;
      RECT  87900.0 192300.0 83400.0 193200.0 ;
      RECT  118200.0 142800.0 117000.0 144750.0 ;
      RECT  118200.0 154950.0 117000.0 156900.0 ;
      RECT  123000.0 144150.0 121800.0 142350.0 ;
      RECT  123000.0 153750.0 121800.0 157350.0 ;
      RECT  120300.0 145350.0 119400.0 153750.0 ;
      RECT  123000.0 153750.0 121800.0 154950.0 ;
      RECT  120600.0 153750.0 119400.0 154950.0 ;
      RECT  120600.0 153750.0 119400.0 154950.0 ;
      RECT  123000.0 153750.0 121800.0 154950.0 ;
      RECT  123000.0 144150.0 121800.0 145350.0 ;
      RECT  120600.0 144150.0 119400.0 145350.0 ;
      RECT  120600.0 144150.0 119400.0 145350.0 ;
      RECT  123000.0 144150.0 121800.0 145350.0 ;
      RECT  118200.0 144150.0 117000.0 145350.0 ;
      RECT  118200.0 154350.0 117000.0 155550.0 ;
      RECT  122400.0 148650.0 121200.0 149850.0 ;
      RECT  122400.0 148650.0 121200.0 149850.0 ;
      RECT  119850.0 148800.0 118950.0 149700.0 ;
      RECT  124800.0 156450.0 115200.0 157350.0 ;
      RECT  124800.0 142350.0 115200.0 143250.0 ;
      RECT  118200.0 171000.0 117000.0 169050.0 ;
      RECT  118200.0 158850.0 117000.0 156900.0 ;
      RECT  123000.0 169650.0 121800.0 171450.0 ;
      RECT  123000.0 160050.0 121800.0 156450.0 ;
      RECT  120300.0 168450.0 119400.0 160050.0 ;
      RECT  123000.0 160050.0 121800.0 158850.0 ;
      RECT  120600.0 160050.0 119400.0 158850.0 ;
      RECT  120600.0 160050.0 119400.0 158850.0 ;
      RECT  123000.0 160050.0 121800.0 158850.0 ;
      RECT  123000.0 169650.0 121800.0 168450.0 ;
      RECT  120600.0 169650.0 119400.0 168450.0 ;
      RECT  120600.0 169650.0 119400.0 168450.0 ;
      RECT  123000.0 169650.0 121800.0 168450.0 ;
      RECT  118200.0 169650.0 117000.0 168450.0 ;
      RECT  118200.0 159450.0 117000.0 158250.0 ;
      RECT  122400.0 165150.0 121200.0 163950.0 ;
      RECT  122400.0 165150.0 121200.0 163950.0 ;
      RECT  119850.0 165000.0 118950.0 164100.0 ;
      RECT  124800.0 157350.0 115200.0 156450.0 ;
      RECT  124800.0 171450.0 115200.0 170550.0 ;
      RECT  79200.0 142800.0 78000.0 144750.0 ;
      RECT  79200.0 154950.0 78000.0 156900.0 ;
      RECT  84000.0 144150.0 82800.0 142350.0 ;
      RECT  84000.0 153750.0 82800.0 157350.0 ;
      RECT  81300.0 145350.0 80400.0 153750.0 ;
      RECT  84000.0 153750.0 82800.0 154950.0 ;
      RECT  81600.0 153750.0 80400.0 154950.0 ;
      RECT  81600.0 153750.0 80400.0 154950.0 ;
      RECT  84000.0 153750.0 82800.0 154950.0 ;
      RECT  84000.0 144150.0 82800.0 145350.0 ;
      RECT  81600.0 144150.0 80400.0 145350.0 ;
      RECT  81600.0 144150.0 80400.0 145350.0 ;
      RECT  84000.0 144150.0 82800.0 145350.0 ;
      RECT  79200.0 144150.0 78000.0 145350.0 ;
      RECT  79200.0 154350.0 78000.0 155550.0 ;
      RECT  83400.0 148650.0 82200.0 149850.0 ;
      RECT  83400.0 148650.0 82200.0 149850.0 ;
      RECT  80850.0 148800.0 79950.0 149700.0 ;
      RECT  85800.0 156450.0 76200.0 157350.0 ;
      RECT  85800.0 142350.0 76200.0 143250.0 ;
      RECT  79200.0 171000.0 78000.0 169050.0 ;
      RECT  79200.0 158850.0 78000.0 156900.0 ;
      RECT  84000.0 169650.0 82800.0 171450.0 ;
      RECT  84000.0 160050.0 82800.0 156450.0 ;
      RECT  81300.0 168450.0 80400.0 160050.0 ;
      RECT  84000.0 160050.0 82800.0 158850.0 ;
      RECT  81600.0 160050.0 80400.0 158850.0 ;
      RECT  81600.0 160050.0 80400.0 158850.0 ;
      RECT  84000.0 160050.0 82800.0 158850.0 ;
      RECT  84000.0 169650.0 82800.0 168450.0 ;
      RECT  81600.0 169650.0 80400.0 168450.0 ;
      RECT  81600.0 169650.0 80400.0 168450.0 ;
      RECT  84000.0 169650.0 82800.0 168450.0 ;
      RECT  79200.0 169650.0 78000.0 168450.0 ;
      RECT  79200.0 159450.0 78000.0 158250.0 ;
      RECT  83400.0 165150.0 82200.0 163950.0 ;
      RECT  83400.0 165150.0 82200.0 163950.0 ;
      RECT  80850.0 165000.0 79950.0 164100.0 ;
      RECT  85800.0 157350.0 76200.0 156450.0 ;
      RECT  85800.0 171450.0 76200.0 170550.0 ;
      RECT  79200.0 171000.0 78000.0 172950.0 ;
      RECT  79200.0 183150.0 78000.0 185100.0 ;
      RECT  84000.0 172350.0 82800.0 170550.0 ;
      RECT  84000.0 181950.0 82800.0 185550.0 ;
      RECT  81300.0 173550.0 80400.0 181950.0 ;
      RECT  84000.0 181950.0 82800.0 183150.0 ;
      RECT  81600.0 181950.0 80400.0 183150.0 ;
      RECT  81600.0 181950.0 80400.0 183150.0 ;
      RECT  84000.0 181950.0 82800.0 183150.0 ;
      RECT  84000.0 172350.0 82800.0 173550.0 ;
      RECT  81600.0 172350.0 80400.0 173550.0 ;
      RECT  81600.0 172350.0 80400.0 173550.0 ;
      RECT  84000.0 172350.0 82800.0 173550.0 ;
      RECT  79200.0 172350.0 78000.0 173550.0 ;
      RECT  79200.0 182550.0 78000.0 183750.0 ;
      RECT  83400.0 176850.0 82200.0 178050.0 ;
      RECT  83400.0 176850.0 82200.0 178050.0 ;
      RECT  80850.0 177000.0 79950.0 177900.0 ;
      RECT  85800.0 184650.0 76200.0 185550.0 ;
      RECT  85800.0 170550.0 76200.0 171450.0 ;
      RECT  79200.0 199200.0 78000.0 197250.0 ;
      RECT  79200.0 187050.0 78000.0 185100.0 ;
      RECT  84000.0 197850.0 82800.0 199650.0 ;
      RECT  84000.0 188250.0 82800.0 184650.0 ;
      RECT  81300.0 196650.0 80400.0 188250.0 ;
      RECT  84000.0 188250.0 82800.0 187050.0 ;
      RECT  81600.0 188250.0 80400.0 187050.0 ;
      RECT  81600.0 188250.0 80400.0 187050.0 ;
      RECT  84000.0 188250.0 82800.0 187050.0 ;
      RECT  84000.0 197850.0 82800.0 196650.0 ;
      RECT  81600.0 197850.0 80400.0 196650.0 ;
      RECT  81600.0 197850.0 80400.0 196650.0 ;
      RECT  84000.0 197850.0 82800.0 196650.0 ;
      RECT  79200.0 197850.0 78000.0 196650.0 ;
      RECT  79200.0 187650.0 78000.0 186450.0 ;
      RECT  83400.0 193350.0 82200.0 192150.0 ;
      RECT  83400.0 193350.0 82200.0 192150.0 ;
      RECT  80850.0 193200.0 79950.0 192300.0 ;
      RECT  85800.0 185550.0 76200.0 184650.0 ;
      RECT  85800.0 199650.0 76200.0 198750.0 ;
      RECT  91200.0 142800.0 90000.0 144750.0 ;
      RECT  91200.0 154950.0 90000.0 156900.0 ;
      RECT  98400.0 144750.0 97200.0 142350.0 ;
      RECT  98400.0 153750.0 97200.0 157350.0 ;
      RECT  93600.0 153750.0 92400.0 157350.0 ;
      RECT  98400.0 153750.0 97200.0 154950.0 ;
      RECT  96000.0 153750.0 94800.0 154950.0 ;
      RECT  96000.0 153750.0 94800.0 154950.0 ;
      RECT  98400.0 153750.0 97200.0 154950.0 ;
      RECT  96000.0 153750.0 94800.0 154950.0 ;
      RECT  93600.0 153750.0 92400.0 154950.0 ;
      RECT  93600.0 153750.0 92400.0 154950.0 ;
      RECT  96000.0 153750.0 94800.0 154950.0 ;
      RECT  98400.0 144750.0 97200.0 145950.0 ;
      RECT  96000.0 144750.0 94800.0 145950.0 ;
      RECT  96000.0 144750.0 94800.0 145950.0 ;
      RECT  98400.0 144750.0 97200.0 145950.0 ;
      RECT  96000.0 144750.0 94800.0 145950.0 ;
      RECT  93600.0 144750.0 92400.0 145950.0 ;
      RECT  93600.0 144750.0 92400.0 145950.0 ;
      RECT  96000.0 144750.0 94800.0 145950.0 ;
      RECT  91200.0 144150.0 90000.0 145350.0 ;
      RECT  91200.0 154350.0 90000.0 155550.0 ;
      RECT  93600.0 147300.0 94800.0 148500.0 ;
      RECT  96600.0 150000.0 97800.0 151200.0 ;
      RECT  96000.0 153750.0 94800.0 154950.0 ;
      RECT  93600.0 144750.0 92400.0 145950.0 ;
      RECT  92400.0 150000.0 93600.0 151200.0 ;
      RECT  97800.0 150000.0 96600.0 151200.0 ;
      RECT  94800.0 147300.0 93600.0 148500.0 ;
      RECT  93600.0 150000.0 92400.0 151200.0 ;
      RECT  100200.0 156450.0 85800.0 157350.0 ;
      RECT  100200.0 142350.0 85800.0 143250.0 ;
      RECT  91200.0 171000.0 90000.0 169050.0 ;
      RECT  91200.0 158850.0 90000.0 156900.0 ;
      RECT  98400.0 169050.0 97200.0 171450.0 ;
      RECT  98400.0 160050.0 97200.0 156450.0 ;
      RECT  93600.0 160050.0 92400.0 156450.0 ;
      RECT  98400.0 160050.0 97200.0 158850.0 ;
      RECT  96000.0 160050.0 94800.0 158850.0 ;
      RECT  96000.0 160050.0 94800.0 158850.0 ;
      RECT  98400.0 160050.0 97200.0 158850.0 ;
      RECT  96000.0 160050.0 94800.0 158850.0 ;
      RECT  93600.0 160050.0 92400.0 158850.0 ;
      RECT  93600.0 160050.0 92400.0 158850.0 ;
      RECT  96000.0 160050.0 94800.0 158850.0 ;
      RECT  98400.0 169050.0 97200.0 167850.0 ;
      RECT  96000.0 169050.0 94800.0 167850.0 ;
      RECT  96000.0 169050.0 94800.0 167850.0 ;
      RECT  98400.0 169050.0 97200.0 167850.0 ;
      RECT  96000.0 169050.0 94800.0 167850.0 ;
      RECT  93600.0 169050.0 92400.0 167850.0 ;
      RECT  93600.0 169050.0 92400.0 167850.0 ;
      RECT  96000.0 169050.0 94800.0 167850.0 ;
      RECT  91200.0 169650.0 90000.0 168450.0 ;
      RECT  91200.0 159450.0 90000.0 158250.0 ;
      RECT  93600.0 166500.0 94800.0 165300.0 ;
      RECT  96600.0 163800.0 97800.0 162600.0 ;
      RECT  96000.0 160050.0 94800.0 158850.0 ;
      RECT  93600.0 169050.0 92400.0 167850.0 ;
      RECT  92400.0 163800.0 93600.0 162600.0 ;
      RECT  97800.0 163800.0 96600.0 162600.0 ;
      RECT  94800.0 166500.0 93600.0 165300.0 ;
      RECT  93600.0 163800.0 92400.0 162600.0 ;
      RECT  100200.0 157350.0 85800.0 156450.0 ;
      RECT  100200.0 171450.0 85800.0 170550.0 ;
      RECT  91200.0 171000.0 90000.0 172950.0 ;
      RECT  91200.0 183150.0 90000.0 185100.0 ;
      RECT  98400.0 172950.0 97200.0 170550.0 ;
      RECT  98400.0 181950.0 97200.0 185550.0 ;
      RECT  93600.0 181950.0 92400.0 185550.0 ;
      RECT  98400.0 181950.0 97200.0 183150.0 ;
      RECT  96000.0 181950.0 94800.0 183150.0 ;
      RECT  96000.0 181950.0 94800.0 183150.0 ;
      RECT  98400.0 181950.0 97200.0 183150.0 ;
      RECT  96000.0 181950.0 94800.0 183150.0 ;
      RECT  93600.0 181950.0 92400.0 183150.0 ;
      RECT  93600.0 181950.0 92400.0 183150.0 ;
      RECT  96000.0 181950.0 94800.0 183150.0 ;
      RECT  98400.0 172950.0 97200.0 174150.0 ;
      RECT  96000.0 172950.0 94800.0 174150.0 ;
      RECT  96000.0 172950.0 94800.0 174150.0 ;
      RECT  98400.0 172950.0 97200.0 174150.0 ;
      RECT  96000.0 172950.0 94800.0 174150.0 ;
      RECT  93600.0 172950.0 92400.0 174150.0 ;
      RECT  93600.0 172950.0 92400.0 174150.0 ;
      RECT  96000.0 172950.0 94800.0 174150.0 ;
      RECT  91200.0 172350.0 90000.0 173550.0 ;
      RECT  91200.0 182550.0 90000.0 183750.0 ;
      RECT  93600.0 175500.0 94800.0 176700.0 ;
      RECT  96600.0 178200.0 97800.0 179400.0 ;
      RECT  96000.0 181950.0 94800.0 183150.0 ;
      RECT  93600.0 172950.0 92400.0 174150.0 ;
      RECT  92400.0 178200.0 93600.0 179400.0 ;
      RECT  97800.0 178200.0 96600.0 179400.0 ;
      RECT  94800.0 175500.0 93600.0 176700.0 ;
      RECT  93600.0 178200.0 92400.0 179400.0 ;
      RECT  100200.0 184650.0 85800.0 185550.0 ;
      RECT  100200.0 170550.0 85800.0 171450.0 ;
      RECT  91200.0 199200.0 90000.0 197250.0 ;
      RECT  91200.0 187050.0 90000.0 185100.0 ;
      RECT  98400.0 197250.0 97200.0 199650.0 ;
      RECT  98400.0 188250.0 97200.0 184650.0 ;
      RECT  93600.0 188250.0 92400.0 184650.0 ;
      RECT  98400.0 188250.0 97200.0 187050.0 ;
      RECT  96000.0 188250.0 94800.0 187050.0 ;
      RECT  96000.0 188250.0 94800.0 187050.0 ;
      RECT  98400.0 188250.0 97200.0 187050.0 ;
      RECT  96000.0 188250.0 94800.0 187050.0 ;
      RECT  93600.0 188250.0 92400.0 187050.0 ;
      RECT  93600.0 188250.0 92400.0 187050.0 ;
      RECT  96000.0 188250.0 94800.0 187050.0 ;
      RECT  98400.0 197250.0 97200.0 196050.0 ;
      RECT  96000.0 197250.0 94800.0 196050.0 ;
      RECT  96000.0 197250.0 94800.0 196050.0 ;
      RECT  98400.0 197250.0 97200.0 196050.0 ;
      RECT  96000.0 197250.0 94800.0 196050.0 ;
      RECT  93600.0 197250.0 92400.0 196050.0 ;
      RECT  93600.0 197250.0 92400.0 196050.0 ;
      RECT  96000.0 197250.0 94800.0 196050.0 ;
      RECT  91200.0 197850.0 90000.0 196650.0 ;
      RECT  91200.0 187650.0 90000.0 186450.0 ;
      RECT  93600.0 194700.0 94800.0 193500.0 ;
      RECT  96600.0 192000.0 97800.0 190800.0 ;
      RECT  96000.0 188250.0 94800.0 187050.0 ;
      RECT  93600.0 197250.0 92400.0 196050.0 ;
      RECT  92400.0 192000.0 93600.0 190800.0 ;
      RECT  97800.0 192000.0 96600.0 190800.0 ;
      RECT  94800.0 194700.0 93600.0 193500.0 ;
      RECT  93600.0 192000.0 92400.0 190800.0 ;
      RECT  100200.0 185550.0 85800.0 184650.0 ;
      RECT  100200.0 199650.0 85800.0 198750.0 ;
      RECT  111150.0 153600.0 112350.0 154800.0 ;
      RECT  129750.0 148650.0 130950.0 149850.0 ;
      RECT  108150.0 167700.0 109350.0 168900.0 ;
      RECT  126750.0 163950.0 127950.0 165150.0 ;
      RECT  129750.0 172500.0 130950.0 173700.0 ;
      RECT  105150.0 172500.0 106350.0 173700.0 ;
      RECT  126750.0 186600.0 127950.0 187800.0 ;
      RECT  102150.0 186600.0 103350.0 187800.0 ;
      RECT  111150.0 150000.0 112350.0 151200.0 ;
      RECT  108150.0 147300.0 109350.0 148500.0 ;
      RECT  105150.0 162600.0 106350.0 163800.0 ;
      RECT  108150.0 165300.0 109350.0 166500.0 ;
      RECT  111150.0 178200.0 112350.0 179400.0 ;
      RECT  102150.0 175500.0 103350.0 176700.0 ;
      RECT  105150.0 190800.0 106350.0 192000.0 ;
      RECT  102150.0 193500.0 103350.0 194700.0 ;
      RECT  79950.0 148800.0 76200.0 149700.0 ;
      RECT  79950.0 164100.0 76200.0 165000.0 ;
      RECT  79950.0 177000.0 76200.0 177900.0 ;
      RECT  79950.0 192300.0 76200.0 193200.0 ;
      RECT  130800.0 156450.0 76200.0 157350.0 ;
      RECT  130800.0 184650.0 76200.0 185550.0 ;
      RECT  130800.0 142350.0 76200.0 143250.0 ;
      RECT  130800.0 170550.0 76200.0 171450.0 ;
      RECT  130800.0 198750.0 76200.0 199650.0 ;
      RECT  85200.0 199200.0 86400.0 201150.0 ;
      RECT  85200.0 211350.0 86400.0 213300.0 ;
      RECT  78000.0 201150.0 79200.0 198750.0 ;
      RECT  78000.0 210150.0 79200.0 213750.0 ;
      RECT  82800.0 210150.0 84000.0 213750.0 ;
      RECT  78000.0 210150.0 79200.0 211350.0 ;
      RECT  80400.0 210150.0 81600.0 211350.0 ;
      RECT  80400.0 210150.0 81600.0 211350.0 ;
      RECT  78000.0 210150.0 79200.0 211350.0 ;
      RECT  80400.0 210150.0 81600.0 211350.0 ;
      RECT  82800.0 210150.0 84000.0 211350.0 ;
      RECT  82800.0 210150.0 84000.0 211350.0 ;
      RECT  80400.0 210150.0 81600.0 211350.0 ;
      RECT  78000.0 201150.0 79200.0 202350.0 ;
      RECT  80400.0 201150.0 81600.0 202350.0 ;
      RECT  80400.0 201150.0 81600.0 202350.0 ;
      RECT  78000.0 201150.0 79200.0 202350.0 ;
      RECT  80400.0 201150.0 81600.0 202350.0 ;
      RECT  82800.0 201150.0 84000.0 202350.0 ;
      RECT  82800.0 201150.0 84000.0 202350.0 ;
      RECT  80400.0 201150.0 81600.0 202350.0 ;
      RECT  85200.0 200550.0 86400.0 201750.0 ;
      RECT  85200.0 210750.0 86400.0 211950.0 ;
      RECT  82800.0 203700.0 81600.0 204900.0 ;
      RECT  79800.0 206400.0 78600.0 207600.0 ;
      RECT  80400.0 210150.0 81600.0 211350.0 ;
      RECT  82800.0 201150.0 84000.0 202350.0 ;
      RECT  84000.0 206400.0 82800.0 207600.0 ;
      RECT  78600.0 206400.0 79800.0 207600.0 ;
      RECT  81600.0 203700.0 82800.0 204900.0 ;
      RECT  82800.0 206400.0 84000.0 207600.0 ;
      RECT  76200.0 212850.0 90600.0 213750.0 ;
      RECT  76200.0 198750.0 90600.0 199650.0 ;
      RECT  85200.0 227400.0 86400.0 225450.0 ;
      RECT  85200.0 215250.0 86400.0 213300.0 ;
      RECT  78000.0 225450.0 79200.0 227850.0 ;
      RECT  78000.0 216450.0 79200.0 212850.0 ;
      RECT  82800.0 216450.0 84000.0 212850.0 ;
      RECT  78000.0 216450.0 79200.0 215250.0 ;
      RECT  80400.0 216450.0 81600.0 215250.0 ;
      RECT  80400.0 216450.0 81600.0 215250.0 ;
      RECT  78000.0 216450.0 79200.0 215250.0 ;
      RECT  80400.0 216450.0 81600.0 215250.0 ;
      RECT  82800.0 216450.0 84000.0 215250.0 ;
      RECT  82800.0 216450.0 84000.0 215250.0 ;
      RECT  80400.0 216450.0 81600.0 215250.0 ;
      RECT  78000.0 225450.0 79200.0 224250.0 ;
      RECT  80400.0 225450.0 81600.0 224250.0 ;
      RECT  80400.0 225450.0 81600.0 224250.0 ;
      RECT  78000.0 225450.0 79200.0 224250.0 ;
      RECT  80400.0 225450.0 81600.0 224250.0 ;
      RECT  82800.0 225450.0 84000.0 224250.0 ;
      RECT  82800.0 225450.0 84000.0 224250.0 ;
      RECT  80400.0 225450.0 81600.0 224250.0 ;
      RECT  85200.0 226050.0 86400.0 224850.0 ;
      RECT  85200.0 215850.0 86400.0 214650.0 ;
      RECT  82800.0 222900.0 81600.0 221700.0 ;
      RECT  79800.0 220200.0 78600.0 219000.0 ;
      RECT  80400.0 216450.0 81600.0 215250.0 ;
      RECT  82800.0 225450.0 84000.0 224250.0 ;
      RECT  84000.0 220200.0 82800.0 219000.0 ;
      RECT  78600.0 220200.0 79800.0 219000.0 ;
      RECT  81600.0 222900.0 82800.0 221700.0 ;
      RECT  82800.0 220200.0 84000.0 219000.0 ;
      RECT  76200.0 213750.0 90600.0 212850.0 ;
      RECT  76200.0 227850.0 90600.0 226950.0 ;
      RECT  85200.0 227400.0 86400.0 229350.0 ;
      RECT  85200.0 239550.0 86400.0 241500.0 ;
      RECT  78000.0 229350.0 79200.0 226950.0 ;
      RECT  78000.0 238350.0 79200.0 241950.0 ;
      RECT  82800.0 238350.0 84000.0 241950.0 ;
      RECT  78000.0 238350.0 79200.0 239550.0 ;
      RECT  80400.0 238350.0 81600.0 239550.0 ;
      RECT  80400.0 238350.0 81600.0 239550.0 ;
      RECT  78000.0 238350.0 79200.0 239550.0 ;
      RECT  80400.0 238350.0 81600.0 239550.0 ;
      RECT  82800.0 238350.0 84000.0 239550.0 ;
      RECT  82800.0 238350.0 84000.0 239550.0 ;
      RECT  80400.0 238350.0 81600.0 239550.0 ;
      RECT  78000.0 229350.0 79200.0 230550.0 ;
      RECT  80400.0 229350.0 81600.0 230550.0 ;
      RECT  80400.0 229350.0 81600.0 230550.0 ;
      RECT  78000.0 229350.0 79200.0 230550.0 ;
      RECT  80400.0 229350.0 81600.0 230550.0 ;
      RECT  82800.0 229350.0 84000.0 230550.0 ;
      RECT  82800.0 229350.0 84000.0 230550.0 ;
      RECT  80400.0 229350.0 81600.0 230550.0 ;
      RECT  85200.0 228750.0 86400.0 229950.0 ;
      RECT  85200.0 238950.0 86400.0 240150.0 ;
      RECT  82800.0 231900.0 81600.0 233100.0 ;
      RECT  79800.0 234600.0 78600.0 235800.0 ;
      RECT  80400.0 238350.0 81600.0 239550.0 ;
      RECT  82800.0 229350.0 84000.0 230550.0 ;
      RECT  84000.0 234600.0 82800.0 235800.0 ;
      RECT  78600.0 234600.0 79800.0 235800.0 ;
      RECT  81600.0 231900.0 82800.0 233100.0 ;
      RECT  82800.0 234600.0 84000.0 235800.0 ;
      RECT  76200.0 241050.0 90600.0 241950.0 ;
      RECT  76200.0 226950.0 90600.0 227850.0 ;
      RECT  85200.0 255600.0 86400.0 253650.0 ;
      RECT  85200.0 243450.0 86400.0 241500.0 ;
      RECT  78000.0 253650.0 79200.0 256050.0 ;
      RECT  78000.0 244650.0 79200.0 241050.0 ;
      RECT  82800.0 244650.0 84000.0 241050.0 ;
      RECT  78000.0 244650.0 79200.0 243450.0 ;
      RECT  80400.0 244650.0 81600.0 243450.0 ;
      RECT  80400.0 244650.0 81600.0 243450.0 ;
      RECT  78000.0 244650.0 79200.0 243450.0 ;
      RECT  80400.0 244650.0 81600.0 243450.0 ;
      RECT  82800.0 244650.0 84000.0 243450.0 ;
      RECT  82800.0 244650.0 84000.0 243450.0 ;
      RECT  80400.0 244650.0 81600.0 243450.0 ;
      RECT  78000.0 253650.0 79200.0 252450.0 ;
      RECT  80400.0 253650.0 81600.0 252450.0 ;
      RECT  80400.0 253650.0 81600.0 252450.0 ;
      RECT  78000.0 253650.0 79200.0 252450.0 ;
      RECT  80400.0 253650.0 81600.0 252450.0 ;
      RECT  82800.0 253650.0 84000.0 252450.0 ;
      RECT  82800.0 253650.0 84000.0 252450.0 ;
      RECT  80400.0 253650.0 81600.0 252450.0 ;
      RECT  85200.0 254250.0 86400.0 253050.0 ;
      RECT  85200.0 244050.0 86400.0 242850.0 ;
      RECT  82800.0 251100.0 81600.0 249900.0 ;
      RECT  79800.0 248400.0 78600.0 247200.0 ;
      RECT  80400.0 244650.0 81600.0 243450.0 ;
      RECT  82800.0 253650.0 84000.0 252450.0 ;
      RECT  84000.0 248400.0 82800.0 247200.0 ;
      RECT  78600.0 248400.0 79800.0 247200.0 ;
      RECT  81600.0 251100.0 82800.0 249900.0 ;
      RECT  82800.0 248400.0 84000.0 247200.0 ;
      RECT  76200.0 241950.0 90600.0 241050.0 ;
      RECT  76200.0 256050.0 90600.0 255150.0 ;
      RECT  85200.0 255600.0 86400.0 257550.0 ;
      RECT  85200.0 267750.0 86400.0 269700.0 ;
      RECT  78000.0 257550.0 79200.0 255150.0 ;
      RECT  78000.0 266550.0 79200.0 270150.0 ;
      RECT  82800.0 266550.0 84000.0 270150.0 ;
      RECT  78000.0 266550.0 79200.0 267750.0 ;
      RECT  80400.0 266550.0 81600.0 267750.0 ;
      RECT  80400.0 266550.0 81600.0 267750.0 ;
      RECT  78000.0 266550.0 79200.0 267750.0 ;
      RECT  80400.0 266550.0 81600.0 267750.0 ;
      RECT  82800.0 266550.0 84000.0 267750.0 ;
      RECT  82800.0 266550.0 84000.0 267750.0 ;
      RECT  80400.0 266550.0 81600.0 267750.0 ;
      RECT  78000.0 257550.0 79200.0 258750.0 ;
      RECT  80400.0 257550.0 81600.0 258750.0 ;
      RECT  80400.0 257550.0 81600.0 258750.0 ;
      RECT  78000.0 257550.0 79200.0 258750.0 ;
      RECT  80400.0 257550.0 81600.0 258750.0 ;
      RECT  82800.0 257550.0 84000.0 258750.0 ;
      RECT  82800.0 257550.0 84000.0 258750.0 ;
      RECT  80400.0 257550.0 81600.0 258750.0 ;
      RECT  85200.0 256950.0 86400.0 258150.0 ;
      RECT  85200.0 267150.0 86400.0 268350.0 ;
      RECT  82800.0 260100.0 81600.0 261300.0 ;
      RECT  79800.0 262800.0 78600.0 264000.0 ;
      RECT  80400.0 266550.0 81600.0 267750.0 ;
      RECT  82800.0 257550.0 84000.0 258750.0 ;
      RECT  84000.0 262800.0 82800.0 264000.0 ;
      RECT  78600.0 262800.0 79800.0 264000.0 ;
      RECT  81600.0 260100.0 82800.0 261300.0 ;
      RECT  82800.0 262800.0 84000.0 264000.0 ;
      RECT  76200.0 269250.0 90600.0 270150.0 ;
      RECT  76200.0 255150.0 90600.0 256050.0 ;
      RECT  85200.0 283800.0 86400.0 281850.0 ;
      RECT  85200.0 271650.0 86400.0 269700.0 ;
      RECT  78000.0 281850.0 79200.0 284250.0 ;
      RECT  78000.0 272850.0 79200.0 269250.0 ;
      RECT  82800.0 272850.0 84000.0 269250.0 ;
      RECT  78000.0 272850.0 79200.0 271650.0 ;
      RECT  80400.0 272850.0 81600.0 271650.0 ;
      RECT  80400.0 272850.0 81600.0 271650.0 ;
      RECT  78000.0 272850.0 79200.0 271650.0 ;
      RECT  80400.0 272850.0 81600.0 271650.0 ;
      RECT  82800.0 272850.0 84000.0 271650.0 ;
      RECT  82800.0 272850.0 84000.0 271650.0 ;
      RECT  80400.0 272850.0 81600.0 271650.0 ;
      RECT  78000.0 281850.0 79200.0 280650.0 ;
      RECT  80400.0 281850.0 81600.0 280650.0 ;
      RECT  80400.0 281850.0 81600.0 280650.0 ;
      RECT  78000.0 281850.0 79200.0 280650.0 ;
      RECT  80400.0 281850.0 81600.0 280650.0 ;
      RECT  82800.0 281850.0 84000.0 280650.0 ;
      RECT  82800.0 281850.0 84000.0 280650.0 ;
      RECT  80400.0 281850.0 81600.0 280650.0 ;
      RECT  85200.0 282450.0 86400.0 281250.0 ;
      RECT  85200.0 272250.0 86400.0 271050.0 ;
      RECT  82800.0 279300.0 81600.0 278100.0 ;
      RECT  79800.0 276600.0 78600.0 275400.0 ;
      RECT  80400.0 272850.0 81600.0 271650.0 ;
      RECT  82800.0 281850.0 84000.0 280650.0 ;
      RECT  84000.0 276600.0 82800.0 275400.0 ;
      RECT  78600.0 276600.0 79800.0 275400.0 ;
      RECT  81600.0 279300.0 82800.0 278100.0 ;
      RECT  82800.0 276600.0 84000.0 275400.0 ;
      RECT  76200.0 270150.0 90600.0 269250.0 ;
      RECT  76200.0 284250.0 90600.0 283350.0 ;
      RECT  85200.0 283800.0 86400.0 285750.0 ;
      RECT  85200.0 295950.0 86400.0 297900.0 ;
      RECT  78000.0 285750.0 79200.0 283350.0 ;
      RECT  78000.0 294750.0 79200.0 298350.0 ;
      RECT  82800.0 294750.0 84000.0 298350.0 ;
      RECT  78000.0 294750.0 79200.0 295950.0 ;
      RECT  80400.0 294750.0 81600.0 295950.0 ;
      RECT  80400.0 294750.0 81600.0 295950.0 ;
      RECT  78000.0 294750.0 79200.0 295950.0 ;
      RECT  80400.0 294750.0 81600.0 295950.0 ;
      RECT  82800.0 294750.0 84000.0 295950.0 ;
      RECT  82800.0 294750.0 84000.0 295950.0 ;
      RECT  80400.0 294750.0 81600.0 295950.0 ;
      RECT  78000.0 285750.0 79200.0 286950.0 ;
      RECT  80400.0 285750.0 81600.0 286950.0 ;
      RECT  80400.0 285750.0 81600.0 286950.0 ;
      RECT  78000.0 285750.0 79200.0 286950.0 ;
      RECT  80400.0 285750.0 81600.0 286950.0 ;
      RECT  82800.0 285750.0 84000.0 286950.0 ;
      RECT  82800.0 285750.0 84000.0 286950.0 ;
      RECT  80400.0 285750.0 81600.0 286950.0 ;
      RECT  85200.0 285150.0 86400.0 286350.0 ;
      RECT  85200.0 295350.0 86400.0 296550.0 ;
      RECT  82800.0 288300.0 81600.0 289500.0 ;
      RECT  79800.0 291000.0 78600.0 292200.0 ;
      RECT  80400.0 294750.0 81600.0 295950.0 ;
      RECT  82800.0 285750.0 84000.0 286950.0 ;
      RECT  84000.0 291000.0 82800.0 292200.0 ;
      RECT  78600.0 291000.0 79800.0 292200.0 ;
      RECT  81600.0 288300.0 82800.0 289500.0 ;
      RECT  82800.0 291000.0 84000.0 292200.0 ;
      RECT  76200.0 297450.0 90600.0 298350.0 ;
      RECT  76200.0 283350.0 90600.0 284250.0 ;
      RECT  85200.0 312000.0 86400.0 310050.0 ;
      RECT  85200.0 299850.0 86400.0 297900.0 ;
      RECT  78000.0 310050.0 79200.0 312450.0 ;
      RECT  78000.0 301050.0 79200.0 297450.0 ;
      RECT  82800.0 301050.0 84000.0 297450.0 ;
      RECT  78000.0 301050.0 79200.0 299850.0 ;
      RECT  80400.0 301050.0 81600.0 299850.0 ;
      RECT  80400.0 301050.0 81600.0 299850.0 ;
      RECT  78000.0 301050.0 79200.0 299850.0 ;
      RECT  80400.0 301050.0 81600.0 299850.0 ;
      RECT  82800.0 301050.0 84000.0 299850.0 ;
      RECT  82800.0 301050.0 84000.0 299850.0 ;
      RECT  80400.0 301050.0 81600.0 299850.0 ;
      RECT  78000.0 310050.0 79200.0 308850.0 ;
      RECT  80400.0 310050.0 81600.0 308850.0 ;
      RECT  80400.0 310050.0 81600.0 308850.0 ;
      RECT  78000.0 310050.0 79200.0 308850.0 ;
      RECT  80400.0 310050.0 81600.0 308850.0 ;
      RECT  82800.0 310050.0 84000.0 308850.0 ;
      RECT  82800.0 310050.0 84000.0 308850.0 ;
      RECT  80400.0 310050.0 81600.0 308850.0 ;
      RECT  85200.0 310650.0 86400.0 309450.0 ;
      RECT  85200.0 300450.0 86400.0 299250.0 ;
      RECT  82800.0 307500.0 81600.0 306300.0 ;
      RECT  79800.0 304800.0 78600.0 303600.0 ;
      RECT  80400.0 301050.0 81600.0 299850.0 ;
      RECT  82800.0 310050.0 84000.0 308850.0 ;
      RECT  84000.0 304800.0 82800.0 303600.0 ;
      RECT  78600.0 304800.0 79800.0 303600.0 ;
      RECT  81600.0 307500.0 82800.0 306300.0 ;
      RECT  82800.0 304800.0 84000.0 303600.0 ;
      RECT  76200.0 298350.0 90600.0 297450.0 ;
      RECT  76200.0 312450.0 90600.0 311550.0 ;
      RECT  85200.0 312000.0 86400.0 313950.0 ;
      RECT  85200.0 324150.0 86400.0 326100.0 ;
      RECT  78000.0 313950.0 79200.0 311550.0 ;
      RECT  78000.0 322950.0 79200.0 326550.0 ;
      RECT  82800.0 322950.0 84000.0 326550.0 ;
      RECT  78000.0 322950.0 79200.0 324150.0 ;
      RECT  80400.0 322950.0 81600.0 324150.0 ;
      RECT  80400.0 322950.0 81600.0 324150.0 ;
      RECT  78000.0 322950.0 79200.0 324150.0 ;
      RECT  80400.0 322950.0 81600.0 324150.0 ;
      RECT  82800.0 322950.0 84000.0 324150.0 ;
      RECT  82800.0 322950.0 84000.0 324150.0 ;
      RECT  80400.0 322950.0 81600.0 324150.0 ;
      RECT  78000.0 313950.0 79200.0 315150.0 ;
      RECT  80400.0 313950.0 81600.0 315150.0 ;
      RECT  80400.0 313950.0 81600.0 315150.0 ;
      RECT  78000.0 313950.0 79200.0 315150.0 ;
      RECT  80400.0 313950.0 81600.0 315150.0 ;
      RECT  82800.0 313950.0 84000.0 315150.0 ;
      RECT  82800.0 313950.0 84000.0 315150.0 ;
      RECT  80400.0 313950.0 81600.0 315150.0 ;
      RECT  85200.0 313350.0 86400.0 314550.0 ;
      RECT  85200.0 323550.0 86400.0 324750.0 ;
      RECT  82800.0 316500.0 81600.0 317700.0 ;
      RECT  79800.0 319200.0 78600.0 320400.0 ;
      RECT  80400.0 322950.0 81600.0 324150.0 ;
      RECT  82800.0 313950.0 84000.0 315150.0 ;
      RECT  84000.0 319200.0 82800.0 320400.0 ;
      RECT  78600.0 319200.0 79800.0 320400.0 ;
      RECT  81600.0 316500.0 82800.0 317700.0 ;
      RECT  82800.0 319200.0 84000.0 320400.0 ;
      RECT  76200.0 325650.0 90600.0 326550.0 ;
      RECT  76200.0 311550.0 90600.0 312450.0 ;
      RECT  85200.0 340200.0 86400.0 338250.0 ;
      RECT  85200.0 328050.0 86400.0 326100.0 ;
      RECT  78000.0 338250.0 79200.0 340650.0 ;
      RECT  78000.0 329250.0 79200.0 325650.0 ;
      RECT  82800.0 329250.0 84000.0 325650.0 ;
      RECT  78000.0 329250.0 79200.0 328050.0 ;
      RECT  80400.0 329250.0 81600.0 328050.0 ;
      RECT  80400.0 329250.0 81600.0 328050.0 ;
      RECT  78000.0 329250.0 79200.0 328050.0 ;
      RECT  80400.0 329250.0 81600.0 328050.0 ;
      RECT  82800.0 329250.0 84000.0 328050.0 ;
      RECT  82800.0 329250.0 84000.0 328050.0 ;
      RECT  80400.0 329250.0 81600.0 328050.0 ;
      RECT  78000.0 338250.0 79200.0 337050.0 ;
      RECT  80400.0 338250.0 81600.0 337050.0 ;
      RECT  80400.0 338250.0 81600.0 337050.0 ;
      RECT  78000.0 338250.0 79200.0 337050.0 ;
      RECT  80400.0 338250.0 81600.0 337050.0 ;
      RECT  82800.0 338250.0 84000.0 337050.0 ;
      RECT  82800.0 338250.0 84000.0 337050.0 ;
      RECT  80400.0 338250.0 81600.0 337050.0 ;
      RECT  85200.0 338850.0 86400.0 337650.0 ;
      RECT  85200.0 328650.0 86400.0 327450.0 ;
      RECT  82800.0 335700.0 81600.0 334500.0 ;
      RECT  79800.0 333000.0 78600.0 331800.0 ;
      RECT  80400.0 329250.0 81600.0 328050.0 ;
      RECT  82800.0 338250.0 84000.0 337050.0 ;
      RECT  84000.0 333000.0 82800.0 331800.0 ;
      RECT  78600.0 333000.0 79800.0 331800.0 ;
      RECT  81600.0 335700.0 82800.0 334500.0 ;
      RECT  82800.0 333000.0 84000.0 331800.0 ;
      RECT  76200.0 326550.0 90600.0 325650.0 ;
      RECT  76200.0 340650.0 90600.0 339750.0 ;
      RECT  85200.0 340200.0 86400.0 342150.0 ;
      RECT  85200.0 352350.0 86400.0 354300.0 ;
      RECT  78000.0 342150.0 79200.0 339750.0 ;
      RECT  78000.0 351150.0 79200.0 354750.0 ;
      RECT  82800.0 351150.0 84000.0 354750.0 ;
      RECT  78000.0 351150.0 79200.0 352350.0 ;
      RECT  80400.0 351150.0 81600.0 352350.0 ;
      RECT  80400.0 351150.0 81600.0 352350.0 ;
      RECT  78000.0 351150.0 79200.0 352350.0 ;
      RECT  80400.0 351150.0 81600.0 352350.0 ;
      RECT  82800.0 351150.0 84000.0 352350.0 ;
      RECT  82800.0 351150.0 84000.0 352350.0 ;
      RECT  80400.0 351150.0 81600.0 352350.0 ;
      RECT  78000.0 342150.0 79200.0 343350.0 ;
      RECT  80400.0 342150.0 81600.0 343350.0 ;
      RECT  80400.0 342150.0 81600.0 343350.0 ;
      RECT  78000.0 342150.0 79200.0 343350.0 ;
      RECT  80400.0 342150.0 81600.0 343350.0 ;
      RECT  82800.0 342150.0 84000.0 343350.0 ;
      RECT  82800.0 342150.0 84000.0 343350.0 ;
      RECT  80400.0 342150.0 81600.0 343350.0 ;
      RECT  85200.0 341550.0 86400.0 342750.0 ;
      RECT  85200.0 351750.0 86400.0 352950.0 ;
      RECT  82800.0 344700.0 81600.0 345900.0 ;
      RECT  79800.0 347400.0 78600.0 348600.0 ;
      RECT  80400.0 351150.0 81600.0 352350.0 ;
      RECT  82800.0 342150.0 84000.0 343350.0 ;
      RECT  84000.0 347400.0 82800.0 348600.0 ;
      RECT  78600.0 347400.0 79800.0 348600.0 ;
      RECT  81600.0 344700.0 82800.0 345900.0 ;
      RECT  82800.0 347400.0 84000.0 348600.0 ;
      RECT  76200.0 353850.0 90600.0 354750.0 ;
      RECT  76200.0 339750.0 90600.0 340650.0 ;
      RECT  85200.0 368400.0 86400.0 366450.0 ;
      RECT  85200.0 356250.0 86400.0 354300.0 ;
      RECT  78000.0 366450.0 79200.0 368850.0 ;
      RECT  78000.0 357450.0 79200.0 353850.0 ;
      RECT  82800.0 357450.0 84000.0 353850.0 ;
      RECT  78000.0 357450.0 79200.0 356250.0 ;
      RECT  80400.0 357450.0 81600.0 356250.0 ;
      RECT  80400.0 357450.0 81600.0 356250.0 ;
      RECT  78000.0 357450.0 79200.0 356250.0 ;
      RECT  80400.0 357450.0 81600.0 356250.0 ;
      RECT  82800.0 357450.0 84000.0 356250.0 ;
      RECT  82800.0 357450.0 84000.0 356250.0 ;
      RECT  80400.0 357450.0 81600.0 356250.0 ;
      RECT  78000.0 366450.0 79200.0 365250.0 ;
      RECT  80400.0 366450.0 81600.0 365250.0 ;
      RECT  80400.0 366450.0 81600.0 365250.0 ;
      RECT  78000.0 366450.0 79200.0 365250.0 ;
      RECT  80400.0 366450.0 81600.0 365250.0 ;
      RECT  82800.0 366450.0 84000.0 365250.0 ;
      RECT  82800.0 366450.0 84000.0 365250.0 ;
      RECT  80400.0 366450.0 81600.0 365250.0 ;
      RECT  85200.0 367050.0 86400.0 365850.0 ;
      RECT  85200.0 356850.0 86400.0 355650.0 ;
      RECT  82800.0 363900.0 81600.0 362700.0 ;
      RECT  79800.0 361200.0 78600.0 360000.0 ;
      RECT  80400.0 357450.0 81600.0 356250.0 ;
      RECT  82800.0 366450.0 84000.0 365250.0 ;
      RECT  84000.0 361200.0 82800.0 360000.0 ;
      RECT  78600.0 361200.0 79800.0 360000.0 ;
      RECT  81600.0 363900.0 82800.0 362700.0 ;
      RECT  82800.0 361200.0 84000.0 360000.0 ;
      RECT  76200.0 354750.0 90600.0 353850.0 ;
      RECT  76200.0 368850.0 90600.0 367950.0 ;
      RECT  85200.0 368400.0 86400.0 370350.0 ;
      RECT  85200.0 380550.0 86400.0 382500.0 ;
      RECT  78000.0 370350.0 79200.0 367950.0 ;
      RECT  78000.0 379350.0 79200.0 382950.0 ;
      RECT  82800.0 379350.0 84000.0 382950.0 ;
      RECT  78000.0 379350.0 79200.0 380550.0 ;
      RECT  80400.0 379350.0 81600.0 380550.0 ;
      RECT  80400.0 379350.0 81600.0 380550.0 ;
      RECT  78000.0 379350.0 79200.0 380550.0 ;
      RECT  80400.0 379350.0 81600.0 380550.0 ;
      RECT  82800.0 379350.0 84000.0 380550.0 ;
      RECT  82800.0 379350.0 84000.0 380550.0 ;
      RECT  80400.0 379350.0 81600.0 380550.0 ;
      RECT  78000.0 370350.0 79200.0 371550.0 ;
      RECT  80400.0 370350.0 81600.0 371550.0 ;
      RECT  80400.0 370350.0 81600.0 371550.0 ;
      RECT  78000.0 370350.0 79200.0 371550.0 ;
      RECT  80400.0 370350.0 81600.0 371550.0 ;
      RECT  82800.0 370350.0 84000.0 371550.0 ;
      RECT  82800.0 370350.0 84000.0 371550.0 ;
      RECT  80400.0 370350.0 81600.0 371550.0 ;
      RECT  85200.0 369750.0 86400.0 370950.0 ;
      RECT  85200.0 379950.0 86400.0 381150.0 ;
      RECT  82800.0 372900.0 81600.0 374100.0 ;
      RECT  79800.0 375600.0 78600.0 376800.0 ;
      RECT  80400.0 379350.0 81600.0 380550.0 ;
      RECT  82800.0 370350.0 84000.0 371550.0 ;
      RECT  84000.0 375600.0 82800.0 376800.0 ;
      RECT  78600.0 375600.0 79800.0 376800.0 ;
      RECT  81600.0 372900.0 82800.0 374100.0 ;
      RECT  82800.0 375600.0 84000.0 376800.0 ;
      RECT  76200.0 382050.0 90600.0 382950.0 ;
      RECT  76200.0 367950.0 90600.0 368850.0 ;
      RECT  85200.0 396600.0 86400.0 394650.0 ;
      RECT  85200.0 384450.0 86400.0 382500.0 ;
      RECT  78000.0 394650.0 79200.0 397050.0 ;
      RECT  78000.0 385650.0 79200.0 382050.0 ;
      RECT  82800.0 385650.0 84000.0 382050.0 ;
      RECT  78000.0 385650.0 79200.0 384450.0 ;
      RECT  80400.0 385650.0 81600.0 384450.0 ;
      RECT  80400.0 385650.0 81600.0 384450.0 ;
      RECT  78000.0 385650.0 79200.0 384450.0 ;
      RECT  80400.0 385650.0 81600.0 384450.0 ;
      RECT  82800.0 385650.0 84000.0 384450.0 ;
      RECT  82800.0 385650.0 84000.0 384450.0 ;
      RECT  80400.0 385650.0 81600.0 384450.0 ;
      RECT  78000.0 394650.0 79200.0 393450.0 ;
      RECT  80400.0 394650.0 81600.0 393450.0 ;
      RECT  80400.0 394650.0 81600.0 393450.0 ;
      RECT  78000.0 394650.0 79200.0 393450.0 ;
      RECT  80400.0 394650.0 81600.0 393450.0 ;
      RECT  82800.0 394650.0 84000.0 393450.0 ;
      RECT  82800.0 394650.0 84000.0 393450.0 ;
      RECT  80400.0 394650.0 81600.0 393450.0 ;
      RECT  85200.0 395250.0 86400.0 394050.0 ;
      RECT  85200.0 385050.0 86400.0 383850.0 ;
      RECT  82800.0 392100.0 81600.0 390900.0 ;
      RECT  79800.0 389400.0 78600.0 388200.0 ;
      RECT  80400.0 385650.0 81600.0 384450.0 ;
      RECT  82800.0 394650.0 84000.0 393450.0 ;
      RECT  84000.0 389400.0 82800.0 388200.0 ;
      RECT  78600.0 389400.0 79800.0 388200.0 ;
      RECT  81600.0 392100.0 82800.0 390900.0 ;
      RECT  82800.0 389400.0 84000.0 388200.0 ;
      RECT  76200.0 382950.0 90600.0 382050.0 ;
      RECT  76200.0 397050.0 90600.0 396150.0 ;
      RECT  85200.0 396600.0 86400.0 398550.0 ;
      RECT  85200.0 408750.0 86400.0 410700.0 ;
      RECT  78000.0 398550.0 79200.0 396150.0 ;
      RECT  78000.0 407550.0 79200.0 411150.0 ;
      RECT  82800.0 407550.0 84000.0 411150.0 ;
      RECT  78000.0 407550.0 79200.0 408750.0 ;
      RECT  80400.0 407550.0 81600.0 408750.0 ;
      RECT  80400.0 407550.0 81600.0 408750.0 ;
      RECT  78000.0 407550.0 79200.0 408750.0 ;
      RECT  80400.0 407550.0 81600.0 408750.0 ;
      RECT  82800.0 407550.0 84000.0 408750.0 ;
      RECT  82800.0 407550.0 84000.0 408750.0 ;
      RECT  80400.0 407550.0 81600.0 408750.0 ;
      RECT  78000.0 398550.0 79200.0 399750.0 ;
      RECT  80400.0 398550.0 81600.0 399750.0 ;
      RECT  80400.0 398550.0 81600.0 399750.0 ;
      RECT  78000.0 398550.0 79200.0 399750.0 ;
      RECT  80400.0 398550.0 81600.0 399750.0 ;
      RECT  82800.0 398550.0 84000.0 399750.0 ;
      RECT  82800.0 398550.0 84000.0 399750.0 ;
      RECT  80400.0 398550.0 81600.0 399750.0 ;
      RECT  85200.0 397950.0 86400.0 399150.0 ;
      RECT  85200.0 408150.0 86400.0 409350.0 ;
      RECT  82800.0 401100.0 81600.0 402300.0 ;
      RECT  79800.0 403800.0 78600.0 405000.0 ;
      RECT  80400.0 407550.0 81600.0 408750.0 ;
      RECT  82800.0 398550.0 84000.0 399750.0 ;
      RECT  84000.0 403800.0 82800.0 405000.0 ;
      RECT  78600.0 403800.0 79800.0 405000.0 ;
      RECT  81600.0 401100.0 82800.0 402300.0 ;
      RECT  82800.0 403800.0 84000.0 405000.0 ;
      RECT  76200.0 410250.0 90600.0 411150.0 ;
      RECT  76200.0 396150.0 90600.0 397050.0 ;
      RECT  85200.0 424800.0 86400.0 422850.0 ;
      RECT  85200.0 412650.0 86400.0 410700.0 ;
      RECT  78000.0 422850.0 79200.0 425250.0 ;
      RECT  78000.0 413850.0 79200.0 410250.0 ;
      RECT  82800.0 413850.0 84000.0 410250.0 ;
      RECT  78000.0 413850.0 79200.0 412650.0 ;
      RECT  80400.0 413850.0 81600.0 412650.0 ;
      RECT  80400.0 413850.0 81600.0 412650.0 ;
      RECT  78000.0 413850.0 79200.0 412650.0 ;
      RECT  80400.0 413850.0 81600.0 412650.0 ;
      RECT  82800.0 413850.0 84000.0 412650.0 ;
      RECT  82800.0 413850.0 84000.0 412650.0 ;
      RECT  80400.0 413850.0 81600.0 412650.0 ;
      RECT  78000.0 422850.0 79200.0 421650.0 ;
      RECT  80400.0 422850.0 81600.0 421650.0 ;
      RECT  80400.0 422850.0 81600.0 421650.0 ;
      RECT  78000.0 422850.0 79200.0 421650.0 ;
      RECT  80400.0 422850.0 81600.0 421650.0 ;
      RECT  82800.0 422850.0 84000.0 421650.0 ;
      RECT  82800.0 422850.0 84000.0 421650.0 ;
      RECT  80400.0 422850.0 81600.0 421650.0 ;
      RECT  85200.0 423450.0 86400.0 422250.0 ;
      RECT  85200.0 413250.0 86400.0 412050.0 ;
      RECT  82800.0 420300.0 81600.0 419100.0 ;
      RECT  79800.0 417600.0 78600.0 416400.0 ;
      RECT  80400.0 413850.0 81600.0 412650.0 ;
      RECT  82800.0 422850.0 84000.0 421650.0 ;
      RECT  84000.0 417600.0 82800.0 416400.0 ;
      RECT  78600.0 417600.0 79800.0 416400.0 ;
      RECT  81600.0 420300.0 82800.0 419100.0 ;
      RECT  82800.0 417600.0 84000.0 416400.0 ;
      RECT  76200.0 411150.0 90600.0 410250.0 ;
      RECT  76200.0 425250.0 90600.0 424350.0 ;
      RECT  97200.0 199200.0 98400.0 201150.0 ;
      RECT  97200.0 211350.0 98400.0 213300.0 ;
      RECT  92400.0 200550.0 93600.0 198750.0 ;
      RECT  92400.0 210150.0 93600.0 213750.0 ;
      RECT  95100.0 201750.0 96000.0 210150.0 ;
      RECT  92400.0 210150.0 93600.0 211350.0 ;
      RECT  94800.0 210150.0 96000.0 211350.0 ;
      RECT  94800.0 210150.0 96000.0 211350.0 ;
      RECT  92400.0 210150.0 93600.0 211350.0 ;
      RECT  92400.0 200550.0 93600.0 201750.0 ;
      RECT  94800.0 200550.0 96000.0 201750.0 ;
      RECT  94800.0 200550.0 96000.0 201750.0 ;
      RECT  92400.0 200550.0 93600.0 201750.0 ;
      RECT  97200.0 200550.0 98400.0 201750.0 ;
      RECT  97200.0 210750.0 98400.0 211950.0 ;
      RECT  93000.0 205050.0 94200.0 206250.0 ;
      RECT  93000.0 205050.0 94200.0 206250.0 ;
      RECT  95550.0 205200.0 96450.0 206100.0 ;
      RECT  90600.0 212850.0 100200.0 213750.0 ;
      RECT  90600.0 198750.0 100200.0 199650.0 ;
      RECT  97200.0 227400.0 98400.0 225450.0 ;
      RECT  97200.0 215250.0 98400.0 213300.0 ;
      RECT  92400.0 226050.0 93600.0 227850.0 ;
      RECT  92400.0 216450.0 93600.0 212850.0 ;
      RECT  95100.0 224850.0 96000.0 216450.0 ;
      RECT  92400.0 216450.0 93600.0 215250.0 ;
      RECT  94800.0 216450.0 96000.0 215250.0 ;
      RECT  94800.0 216450.0 96000.0 215250.0 ;
      RECT  92400.0 216450.0 93600.0 215250.0 ;
      RECT  92400.0 226050.0 93600.0 224850.0 ;
      RECT  94800.0 226050.0 96000.0 224850.0 ;
      RECT  94800.0 226050.0 96000.0 224850.0 ;
      RECT  92400.0 226050.0 93600.0 224850.0 ;
      RECT  97200.0 226050.0 98400.0 224850.0 ;
      RECT  97200.0 215850.0 98400.0 214650.0 ;
      RECT  93000.0 221550.0 94200.0 220350.0 ;
      RECT  93000.0 221550.0 94200.0 220350.0 ;
      RECT  95550.0 221400.0 96450.0 220500.0 ;
      RECT  90600.0 213750.0 100200.0 212850.0 ;
      RECT  90600.0 227850.0 100200.0 226950.0 ;
      RECT  97200.0 227400.0 98400.0 229350.0 ;
      RECT  97200.0 239550.0 98400.0 241500.0 ;
      RECT  92400.0 228750.0 93600.0 226950.0 ;
      RECT  92400.0 238350.0 93600.0 241950.0 ;
      RECT  95100.0 229950.0 96000.0 238350.0 ;
      RECT  92400.0 238350.0 93600.0 239550.0 ;
      RECT  94800.0 238350.0 96000.0 239550.0 ;
      RECT  94800.0 238350.0 96000.0 239550.0 ;
      RECT  92400.0 238350.0 93600.0 239550.0 ;
      RECT  92400.0 228750.0 93600.0 229950.0 ;
      RECT  94800.0 228750.0 96000.0 229950.0 ;
      RECT  94800.0 228750.0 96000.0 229950.0 ;
      RECT  92400.0 228750.0 93600.0 229950.0 ;
      RECT  97200.0 228750.0 98400.0 229950.0 ;
      RECT  97200.0 238950.0 98400.0 240150.0 ;
      RECT  93000.0 233250.0 94200.0 234450.0 ;
      RECT  93000.0 233250.0 94200.0 234450.0 ;
      RECT  95550.0 233400.0 96450.0 234300.0 ;
      RECT  90600.0 241050.0 100200.0 241950.0 ;
      RECT  90600.0 226950.0 100200.0 227850.0 ;
      RECT  97200.0 255600.0 98400.0 253650.0 ;
      RECT  97200.0 243450.0 98400.0 241500.0 ;
      RECT  92400.0 254250.0 93600.0 256050.0 ;
      RECT  92400.0 244650.0 93600.0 241050.0 ;
      RECT  95100.0 253050.0 96000.0 244650.0 ;
      RECT  92400.0 244650.0 93600.0 243450.0 ;
      RECT  94800.0 244650.0 96000.0 243450.0 ;
      RECT  94800.0 244650.0 96000.0 243450.0 ;
      RECT  92400.0 244650.0 93600.0 243450.0 ;
      RECT  92400.0 254250.0 93600.0 253050.0 ;
      RECT  94800.0 254250.0 96000.0 253050.0 ;
      RECT  94800.0 254250.0 96000.0 253050.0 ;
      RECT  92400.0 254250.0 93600.0 253050.0 ;
      RECT  97200.0 254250.0 98400.0 253050.0 ;
      RECT  97200.0 244050.0 98400.0 242850.0 ;
      RECT  93000.0 249750.0 94200.0 248550.0 ;
      RECT  93000.0 249750.0 94200.0 248550.0 ;
      RECT  95550.0 249600.0 96450.0 248700.0 ;
      RECT  90600.0 241950.0 100200.0 241050.0 ;
      RECT  90600.0 256050.0 100200.0 255150.0 ;
      RECT  97200.0 255600.0 98400.0 257550.0 ;
      RECT  97200.0 267750.0 98400.0 269700.0 ;
      RECT  92400.0 256950.0 93600.0 255150.0 ;
      RECT  92400.0 266550.0 93600.0 270150.0 ;
      RECT  95100.0 258150.0 96000.0 266550.0 ;
      RECT  92400.0 266550.0 93600.0 267750.0 ;
      RECT  94800.0 266550.0 96000.0 267750.0 ;
      RECT  94800.0 266550.0 96000.0 267750.0 ;
      RECT  92400.0 266550.0 93600.0 267750.0 ;
      RECT  92400.0 256950.0 93600.0 258150.0 ;
      RECT  94800.0 256950.0 96000.0 258150.0 ;
      RECT  94800.0 256950.0 96000.0 258150.0 ;
      RECT  92400.0 256950.0 93600.0 258150.0 ;
      RECT  97200.0 256950.0 98400.0 258150.0 ;
      RECT  97200.0 267150.0 98400.0 268350.0 ;
      RECT  93000.0 261450.0 94200.0 262650.0 ;
      RECT  93000.0 261450.0 94200.0 262650.0 ;
      RECT  95550.0 261600.0 96450.0 262500.0 ;
      RECT  90600.0 269250.0 100200.0 270150.0 ;
      RECT  90600.0 255150.0 100200.0 256050.0 ;
      RECT  97200.0 283800.0 98400.0 281850.0 ;
      RECT  97200.0 271650.0 98400.0 269700.0 ;
      RECT  92400.0 282450.0 93600.0 284250.0 ;
      RECT  92400.0 272850.0 93600.0 269250.0 ;
      RECT  95100.0 281250.0 96000.0 272850.0 ;
      RECT  92400.0 272850.0 93600.0 271650.0 ;
      RECT  94800.0 272850.0 96000.0 271650.0 ;
      RECT  94800.0 272850.0 96000.0 271650.0 ;
      RECT  92400.0 272850.0 93600.0 271650.0 ;
      RECT  92400.0 282450.0 93600.0 281250.0 ;
      RECT  94800.0 282450.0 96000.0 281250.0 ;
      RECT  94800.0 282450.0 96000.0 281250.0 ;
      RECT  92400.0 282450.0 93600.0 281250.0 ;
      RECT  97200.0 282450.0 98400.0 281250.0 ;
      RECT  97200.0 272250.0 98400.0 271050.0 ;
      RECT  93000.0 277950.0 94200.0 276750.0 ;
      RECT  93000.0 277950.0 94200.0 276750.0 ;
      RECT  95550.0 277800.0 96450.0 276900.0 ;
      RECT  90600.0 270150.0 100200.0 269250.0 ;
      RECT  90600.0 284250.0 100200.0 283350.0 ;
      RECT  97200.0 283800.0 98400.0 285750.0 ;
      RECT  97200.0 295950.0 98400.0 297900.0 ;
      RECT  92400.0 285150.0 93600.0 283350.0 ;
      RECT  92400.0 294750.0 93600.0 298350.0 ;
      RECT  95100.0 286350.0 96000.0 294750.0 ;
      RECT  92400.0 294750.0 93600.0 295950.0 ;
      RECT  94800.0 294750.0 96000.0 295950.0 ;
      RECT  94800.0 294750.0 96000.0 295950.0 ;
      RECT  92400.0 294750.0 93600.0 295950.0 ;
      RECT  92400.0 285150.0 93600.0 286350.0 ;
      RECT  94800.0 285150.0 96000.0 286350.0 ;
      RECT  94800.0 285150.0 96000.0 286350.0 ;
      RECT  92400.0 285150.0 93600.0 286350.0 ;
      RECT  97200.0 285150.0 98400.0 286350.0 ;
      RECT  97200.0 295350.0 98400.0 296550.0 ;
      RECT  93000.0 289650.0 94200.0 290850.0 ;
      RECT  93000.0 289650.0 94200.0 290850.0 ;
      RECT  95550.0 289800.0 96450.0 290700.0 ;
      RECT  90600.0 297450.0 100200.0 298350.0 ;
      RECT  90600.0 283350.0 100200.0 284250.0 ;
      RECT  97200.0 312000.0 98400.0 310050.0 ;
      RECT  97200.0 299850.0 98400.0 297900.0 ;
      RECT  92400.0 310650.0 93600.0 312450.0 ;
      RECT  92400.0 301050.0 93600.0 297450.0 ;
      RECT  95100.0 309450.0 96000.0 301050.0 ;
      RECT  92400.0 301050.0 93600.0 299850.0 ;
      RECT  94800.0 301050.0 96000.0 299850.0 ;
      RECT  94800.0 301050.0 96000.0 299850.0 ;
      RECT  92400.0 301050.0 93600.0 299850.0 ;
      RECT  92400.0 310650.0 93600.0 309450.0 ;
      RECT  94800.0 310650.0 96000.0 309450.0 ;
      RECT  94800.0 310650.0 96000.0 309450.0 ;
      RECT  92400.0 310650.0 93600.0 309450.0 ;
      RECT  97200.0 310650.0 98400.0 309450.0 ;
      RECT  97200.0 300450.0 98400.0 299250.0 ;
      RECT  93000.0 306150.0 94200.0 304950.0 ;
      RECT  93000.0 306150.0 94200.0 304950.0 ;
      RECT  95550.0 306000.0 96450.0 305100.0 ;
      RECT  90600.0 298350.0 100200.0 297450.0 ;
      RECT  90600.0 312450.0 100200.0 311550.0 ;
      RECT  97200.0 312000.0 98400.0 313950.0 ;
      RECT  97200.0 324150.0 98400.0 326100.0 ;
      RECT  92400.0 313350.0 93600.0 311550.0 ;
      RECT  92400.0 322950.0 93600.0 326550.0 ;
      RECT  95100.0 314550.0 96000.0 322950.0 ;
      RECT  92400.0 322950.0 93600.0 324150.0 ;
      RECT  94800.0 322950.0 96000.0 324150.0 ;
      RECT  94800.0 322950.0 96000.0 324150.0 ;
      RECT  92400.0 322950.0 93600.0 324150.0 ;
      RECT  92400.0 313350.0 93600.0 314550.0 ;
      RECT  94800.0 313350.0 96000.0 314550.0 ;
      RECT  94800.0 313350.0 96000.0 314550.0 ;
      RECT  92400.0 313350.0 93600.0 314550.0 ;
      RECT  97200.0 313350.0 98400.0 314550.0 ;
      RECT  97200.0 323550.0 98400.0 324750.0 ;
      RECT  93000.0 317850.0 94200.0 319050.0 ;
      RECT  93000.0 317850.0 94200.0 319050.0 ;
      RECT  95550.0 318000.0 96450.0 318900.0 ;
      RECT  90600.0 325650.0 100200.0 326550.0 ;
      RECT  90600.0 311550.0 100200.0 312450.0 ;
      RECT  97200.0 340200.0 98400.0 338250.0 ;
      RECT  97200.0 328050.0 98400.0 326100.0 ;
      RECT  92400.0 338850.0 93600.0 340650.0 ;
      RECT  92400.0 329250.0 93600.0 325650.0 ;
      RECT  95100.0 337650.0 96000.0 329250.0 ;
      RECT  92400.0 329250.0 93600.0 328050.0 ;
      RECT  94800.0 329250.0 96000.0 328050.0 ;
      RECT  94800.0 329250.0 96000.0 328050.0 ;
      RECT  92400.0 329250.0 93600.0 328050.0 ;
      RECT  92400.0 338850.0 93600.0 337650.0 ;
      RECT  94800.0 338850.0 96000.0 337650.0 ;
      RECT  94800.0 338850.0 96000.0 337650.0 ;
      RECT  92400.0 338850.0 93600.0 337650.0 ;
      RECT  97200.0 338850.0 98400.0 337650.0 ;
      RECT  97200.0 328650.0 98400.0 327450.0 ;
      RECT  93000.0 334350.0 94200.0 333150.0 ;
      RECT  93000.0 334350.0 94200.0 333150.0 ;
      RECT  95550.0 334200.0 96450.0 333300.0 ;
      RECT  90600.0 326550.0 100200.0 325650.0 ;
      RECT  90600.0 340650.0 100200.0 339750.0 ;
      RECT  97200.0 340200.0 98400.0 342150.0 ;
      RECT  97200.0 352350.0 98400.0 354300.0 ;
      RECT  92400.0 341550.0 93600.0 339750.0 ;
      RECT  92400.0 351150.0 93600.0 354750.0 ;
      RECT  95100.0 342750.0 96000.0 351150.0 ;
      RECT  92400.0 351150.0 93600.0 352350.0 ;
      RECT  94800.0 351150.0 96000.0 352350.0 ;
      RECT  94800.0 351150.0 96000.0 352350.0 ;
      RECT  92400.0 351150.0 93600.0 352350.0 ;
      RECT  92400.0 341550.0 93600.0 342750.0 ;
      RECT  94800.0 341550.0 96000.0 342750.0 ;
      RECT  94800.0 341550.0 96000.0 342750.0 ;
      RECT  92400.0 341550.0 93600.0 342750.0 ;
      RECT  97200.0 341550.0 98400.0 342750.0 ;
      RECT  97200.0 351750.0 98400.0 352950.0 ;
      RECT  93000.0 346050.0 94200.0 347250.0 ;
      RECT  93000.0 346050.0 94200.0 347250.0 ;
      RECT  95550.0 346200.0 96450.0 347100.0 ;
      RECT  90600.0 353850.0 100200.0 354750.0 ;
      RECT  90600.0 339750.0 100200.0 340650.0 ;
      RECT  97200.0 368400.0 98400.0 366450.0 ;
      RECT  97200.0 356250.0 98400.0 354300.0 ;
      RECT  92400.0 367050.0 93600.0 368850.0 ;
      RECT  92400.0 357450.0 93600.0 353850.0 ;
      RECT  95100.0 365850.0 96000.0 357450.0 ;
      RECT  92400.0 357450.0 93600.0 356250.0 ;
      RECT  94800.0 357450.0 96000.0 356250.0 ;
      RECT  94800.0 357450.0 96000.0 356250.0 ;
      RECT  92400.0 357450.0 93600.0 356250.0 ;
      RECT  92400.0 367050.0 93600.0 365850.0 ;
      RECT  94800.0 367050.0 96000.0 365850.0 ;
      RECT  94800.0 367050.0 96000.0 365850.0 ;
      RECT  92400.0 367050.0 93600.0 365850.0 ;
      RECT  97200.0 367050.0 98400.0 365850.0 ;
      RECT  97200.0 356850.0 98400.0 355650.0 ;
      RECT  93000.0 362550.0 94200.0 361350.0 ;
      RECT  93000.0 362550.0 94200.0 361350.0 ;
      RECT  95550.0 362400.0 96450.0 361500.0 ;
      RECT  90600.0 354750.0 100200.0 353850.0 ;
      RECT  90600.0 368850.0 100200.0 367950.0 ;
      RECT  97200.0 368400.0 98400.0 370350.0 ;
      RECT  97200.0 380550.0 98400.0 382500.0 ;
      RECT  92400.0 369750.0 93600.0 367950.0 ;
      RECT  92400.0 379350.0 93600.0 382950.0 ;
      RECT  95100.0 370950.0 96000.0 379350.0 ;
      RECT  92400.0 379350.0 93600.0 380550.0 ;
      RECT  94800.0 379350.0 96000.0 380550.0 ;
      RECT  94800.0 379350.0 96000.0 380550.0 ;
      RECT  92400.0 379350.0 93600.0 380550.0 ;
      RECT  92400.0 369750.0 93600.0 370950.0 ;
      RECT  94800.0 369750.0 96000.0 370950.0 ;
      RECT  94800.0 369750.0 96000.0 370950.0 ;
      RECT  92400.0 369750.0 93600.0 370950.0 ;
      RECT  97200.0 369750.0 98400.0 370950.0 ;
      RECT  97200.0 379950.0 98400.0 381150.0 ;
      RECT  93000.0 374250.0 94200.0 375450.0 ;
      RECT  93000.0 374250.0 94200.0 375450.0 ;
      RECT  95550.0 374400.0 96450.0 375300.0 ;
      RECT  90600.0 382050.0 100200.0 382950.0 ;
      RECT  90600.0 367950.0 100200.0 368850.0 ;
      RECT  97200.0 396600.0 98400.0 394650.0 ;
      RECT  97200.0 384450.0 98400.0 382500.0 ;
      RECT  92400.0 395250.0 93600.0 397050.0 ;
      RECT  92400.0 385650.0 93600.0 382050.0 ;
      RECT  95100.0 394050.0 96000.0 385650.0 ;
      RECT  92400.0 385650.0 93600.0 384450.0 ;
      RECT  94800.0 385650.0 96000.0 384450.0 ;
      RECT  94800.0 385650.0 96000.0 384450.0 ;
      RECT  92400.0 385650.0 93600.0 384450.0 ;
      RECT  92400.0 395250.0 93600.0 394050.0 ;
      RECT  94800.0 395250.0 96000.0 394050.0 ;
      RECT  94800.0 395250.0 96000.0 394050.0 ;
      RECT  92400.0 395250.0 93600.0 394050.0 ;
      RECT  97200.0 395250.0 98400.0 394050.0 ;
      RECT  97200.0 385050.0 98400.0 383850.0 ;
      RECT  93000.0 390750.0 94200.0 389550.0 ;
      RECT  93000.0 390750.0 94200.0 389550.0 ;
      RECT  95550.0 390600.0 96450.0 389700.0 ;
      RECT  90600.0 382950.0 100200.0 382050.0 ;
      RECT  90600.0 397050.0 100200.0 396150.0 ;
      RECT  97200.0 396600.0 98400.0 398550.0 ;
      RECT  97200.0 408750.0 98400.0 410700.0 ;
      RECT  92400.0 397950.0 93600.0 396150.0 ;
      RECT  92400.0 407550.0 93600.0 411150.0 ;
      RECT  95100.0 399150.0 96000.0 407550.0 ;
      RECT  92400.0 407550.0 93600.0 408750.0 ;
      RECT  94800.0 407550.0 96000.0 408750.0 ;
      RECT  94800.0 407550.0 96000.0 408750.0 ;
      RECT  92400.0 407550.0 93600.0 408750.0 ;
      RECT  92400.0 397950.0 93600.0 399150.0 ;
      RECT  94800.0 397950.0 96000.0 399150.0 ;
      RECT  94800.0 397950.0 96000.0 399150.0 ;
      RECT  92400.0 397950.0 93600.0 399150.0 ;
      RECT  97200.0 397950.0 98400.0 399150.0 ;
      RECT  97200.0 408150.0 98400.0 409350.0 ;
      RECT  93000.0 402450.0 94200.0 403650.0 ;
      RECT  93000.0 402450.0 94200.0 403650.0 ;
      RECT  95550.0 402600.0 96450.0 403500.0 ;
      RECT  90600.0 410250.0 100200.0 411150.0 ;
      RECT  90600.0 396150.0 100200.0 397050.0 ;
      RECT  97200.0 424800.0 98400.0 422850.0 ;
      RECT  97200.0 412650.0 98400.0 410700.0 ;
      RECT  92400.0 423450.0 93600.0 425250.0 ;
      RECT  92400.0 413850.0 93600.0 410250.0 ;
      RECT  95100.0 422250.0 96000.0 413850.0 ;
      RECT  92400.0 413850.0 93600.0 412650.0 ;
      RECT  94800.0 413850.0 96000.0 412650.0 ;
      RECT  94800.0 413850.0 96000.0 412650.0 ;
      RECT  92400.0 413850.0 93600.0 412650.0 ;
      RECT  92400.0 423450.0 93600.0 422250.0 ;
      RECT  94800.0 423450.0 96000.0 422250.0 ;
      RECT  94800.0 423450.0 96000.0 422250.0 ;
      RECT  92400.0 423450.0 93600.0 422250.0 ;
      RECT  97200.0 423450.0 98400.0 422250.0 ;
      RECT  97200.0 413250.0 98400.0 412050.0 ;
      RECT  93000.0 418950.0 94200.0 417750.0 ;
      RECT  93000.0 418950.0 94200.0 417750.0 ;
      RECT  95550.0 418800.0 96450.0 417900.0 ;
      RECT  90600.0 411150.0 100200.0 410250.0 ;
      RECT  90600.0 425250.0 100200.0 424350.0 ;
      RECT  60450.0 92250.0 59250.0 93450.0 ;
      RECT  62550.0 107550.0 61350.0 108750.0 ;
      RECT  64650.0 120450.0 63450.0 121650.0 ;
      RECT  66750.0 135750.0 65550.0 136950.0 ;
      RECT  68850.0 148650.0 67650.0 149850.0 ;
      RECT  70950.0 163950.0 69750.0 165150.0 ;
      RECT  73050.0 176850.0 71850.0 178050.0 ;
      RECT  75150.0 192150.0 73950.0 193350.0 ;
      RECT  60450.0 206400.0 59250.0 207600.0 ;
      RECT  68850.0 203700.0 67650.0 204900.0 ;
      RECT  60450.0 219000.0 59250.0 220200.0 ;
      RECT  70950.0 221700.0 69750.0 222900.0 ;
      RECT  60450.0 234600.0 59250.0 235800.0 ;
      RECT  73050.0 231900.0 71850.0 233100.0 ;
      RECT  60450.0 247200.0 59250.0 248400.0 ;
      RECT  75150.0 249900.0 73950.0 251100.0 ;
      RECT  62550.0 262800.0 61350.0 264000.0 ;
      RECT  68850.0 260100.0 67650.0 261300.0 ;
      RECT  62550.0 275400.0 61350.0 276600.0 ;
      RECT  70950.0 278100.0 69750.0 279300.0 ;
      RECT  62550.0 291000.0 61350.0 292200.0 ;
      RECT  73050.0 288300.0 71850.0 289500.0 ;
      RECT  62550.0 303600.0 61350.0 304800.0 ;
      RECT  75150.0 306300.0 73950.0 307500.0 ;
      RECT  64650.0 319200.0 63450.0 320400.0 ;
      RECT  68850.0 316500.0 67650.0 317700.0 ;
      RECT  64650.0 331800.0 63450.0 333000.0 ;
      RECT  70950.0 334500.0 69750.0 335700.0 ;
      RECT  64650.0 347400.0 63450.0 348600.0 ;
      RECT  73050.0 344700.0 71850.0 345900.0 ;
      RECT  64650.0 360000.0 63450.0 361200.0 ;
      RECT  75150.0 362700.0 73950.0 363900.0 ;
      RECT  66750.0 375600.0 65550.0 376800.0 ;
      RECT  68850.0 372900.0 67650.0 374100.0 ;
      RECT  66750.0 388200.0 65550.0 389400.0 ;
      RECT  70950.0 390900.0 69750.0 392100.0 ;
      RECT  66750.0 403800.0 65550.0 405000.0 ;
      RECT  73050.0 401100.0 71850.0 402300.0 ;
      RECT  66750.0 416400.0 65550.0 417600.0 ;
      RECT  75150.0 419100.0 73950.0 420300.0 ;
      RECT  95550.0 205200.0 96450.0 206100.0 ;
      RECT  95550.0 220500.0 96450.0 221400.0 ;
      RECT  95550.0 233400.0 96450.0 234300.0 ;
      RECT  95550.0 248700.0 96450.0 249600.0 ;
      RECT  95550.0 261600.0 96450.0 262500.0 ;
      RECT  95550.0 276900.0 96450.0 277800.0 ;
      RECT  95550.0 289800.0 96450.0 290700.0 ;
      RECT  95550.0 305100.0 96450.0 306000.0 ;
      RECT  95550.0 318000.0 96450.0 318900.0 ;
      RECT  95550.0 333300.0 96450.0 334200.0 ;
      RECT  95550.0 346200.0 96450.0 347100.0 ;
      RECT  95550.0 361500.0 96450.0 362400.0 ;
      RECT  95550.0 374400.0 96450.0 375300.0 ;
      RECT  95550.0 389700.0 96450.0 390600.0 ;
      RECT  95550.0 402600.0 96450.0 403500.0 ;
      RECT  95550.0 417900.0 96450.0 418800.0 ;
      RECT  59400.0 100050.0 130800.0 100950.0 ;
      RECT  59400.0 128250.0 130800.0 129150.0 ;
      RECT  59400.0 156450.0 130800.0 157350.0 ;
      RECT  59400.0 184650.0 130800.0 185550.0 ;
      RECT  59400.0 212850.0 130800.0 213750.0 ;
      RECT  59400.0 241050.0 130800.0 241950.0 ;
      RECT  59400.0 269250.0 130800.0 270150.0 ;
      RECT  59400.0 297450.0 130800.0 298350.0 ;
      RECT  59400.0 325650.0 130800.0 326550.0 ;
      RECT  59400.0 353850.0 130800.0 354750.0 ;
      RECT  59400.0 382050.0 130800.0 382950.0 ;
      RECT  59400.0 410250.0 130800.0 411150.0 ;
      RECT  59400.0 85950.0 130800.0 86850.0 ;
      RECT  59400.0 114150.0 130800.0 115050.0 ;
      RECT  59400.0 142350.0 130800.0 143250.0 ;
      RECT  59400.0 170550.0 130800.0 171450.0 ;
      RECT  59400.0 198750.0 130800.0 199650.0 ;
      RECT  59400.0 226950.0 130800.0 227850.0 ;
      RECT  59400.0 255150.0 130800.0 256050.0 ;
      RECT  59400.0 283350.0 130800.0 284250.0 ;
      RECT  59400.0 311550.0 130800.0 312450.0 ;
      RECT  59400.0 339750.0 130800.0 340650.0 ;
      RECT  59400.0 367950.0 130800.0 368850.0 ;
      RECT  59400.0 396150.0 130800.0 397050.0 ;
      RECT  59400.0 424350.0 130800.0 425250.0 ;
      RECT  103350.0 205200.0 108900.0 206100.0 ;
      RECT  111450.0 206550.0 112350.0 207450.0 ;
      RECT  111450.0 205200.0 112350.0 206100.0 ;
      RECT  111450.0 206100.0 112350.0 207000.0 ;
      RECT  111900.0 206550.0 118500.0 207450.0 ;
      RECT  118500.0 206550.0 119700.0 207450.0 ;
      RECT  127950.0 206550.0 128850.0 207450.0 ;
      RECT  127950.0 205200.0 128850.0 206100.0 ;
      RECT  123900.0 206550.0 128400.0 207450.0 ;
      RECT  127950.0 205650.0 128850.0 207000.0 ;
      RECT  128400.0 205200.0 132900.0 206100.0 ;
      RECT  103350.0 220500.0 108900.0 221400.0 ;
      RECT  111450.0 219150.0 112350.0 220050.0 ;
      RECT  111450.0 220500.0 112350.0 221400.0 ;
      RECT  111450.0 219600.0 112350.0 221400.0 ;
      RECT  111900.0 219150.0 118500.0 220050.0 ;
      RECT  118500.0 219150.0 119700.0 220050.0 ;
      RECT  127950.0 219150.0 128850.0 220050.0 ;
      RECT  127950.0 220500.0 128850.0 221400.0 ;
      RECT  123900.0 219150.0 128400.0 220050.0 ;
      RECT  127950.0 219600.0 128850.0 220950.0 ;
      RECT  128400.0 220500.0 132900.0 221400.0 ;
      RECT  103350.0 233400.0 108900.0 234300.0 ;
      RECT  111450.0 234750.0 112350.0 235650.0 ;
      RECT  111450.0 233400.0 112350.0 234300.0 ;
      RECT  111450.0 234300.0 112350.0 235200.0 ;
      RECT  111900.0 234750.0 118500.0 235650.0 ;
      RECT  118500.0 234750.0 119700.0 235650.0 ;
      RECT  127950.0 234750.0 128850.0 235650.0 ;
      RECT  127950.0 233400.0 128850.0 234300.0 ;
      RECT  123900.0 234750.0 128400.0 235650.0 ;
      RECT  127950.0 233850.0 128850.0 235200.0 ;
      RECT  128400.0 233400.0 132900.0 234300.0 ;
      RECT  103350.0 248700.0 108900.0 249600.0 ;
      RECT  111450.0 247350.0 112350.0 248250.0 ;
      RECT  111450.0 248700.0 112350.0 249600.0 ;
      RECT  111450.0 247800.0 112350.0 249600.0 ;
      RECT  111900.0 247350.0 118500.0 248250.0 ;
      RECT  118500.0 247350.0 119700.0 248250.0 ;
      RECT  127950.0 247350.0 128850.0 248250.0 ;
      RECT  127950.0 248700.0 128850.0 249600.0 ;
      RECT  123900.0 247350.0 128400.0 248250.0 ;
      RECT  127950.0 247800.0 128850.0 249150.0 ;
      RECT  128400.0 248700.0 132900.0 249600.0 ;
      RECT  103350.0 261600.0 108900.0 262500.0 ;
      RECT  111450.0 262950.0 112350.0 263850.0 ;
      RECT  111450.0 261600.0 112350.0 262500.0 ;
      RECT  111450.0 262500.0 112350.0 263400.0 ;
      RECT  111900.0 262950.0 118500.0 263850.0 ;
      RECT  118500.0 262950.0 119700.0 263850.0 ;
      RECT  127950.0 262950.0 128850.0 263850.0 ;
      RECT  127950.0 261600.0 128850.0 262500.0 ;
      RECT  123900.0 262950.0 128400.0 263850.0 ;
      RECT  127950.0 262050.0 128850.0 263400.0 ;
      RECT  128400.0 261600.0 132900.0 262500.0 ;
      RECT  103350.0 276900.0 108900.0 277800.0 ;
      RECT  111450.0 275550.0 112350.0 276450.0 ;
      RECT  111450.0 276900.0 112350.0 277800.0 ;
      RECT  111450.0 276000.0 112350.0 277800.0 ;
      RECT  111900.0 275550.0 118500.0 276450.0 ;
      RECT  118500.0 275550.0 119700.0 276450.0 ;
      RECT  127950.0 275550.0 128850.0 276450.0 ;
      RECT  127950.0 276900.0 128850.0 277800.0 ;
      RECT  123900.0 275550.0 128400.0 276450.0 ;
      RECT  127950.0 276000.0 128850.0 277350.0 ;
      RECT  128400.0 276900.0 132900.0 277800.0 ;
      RECT  103350.0 289800.0 108900.0 290700.0 ;
      RECT  111450.0 291150.0 112350.0 292050.0 ;
      RECT  111450.0 289800.0 112350.0 290700.0 ;
      RECT  111450.0 290700.0 112350.0 291600.0 ;
      RECT  111900.0 291150.0 118500.0 292050.0 ;
      RECT  118500.0 291150.0 119700.0 292050.0 ;
      RECT  127950.0 291150.0 128850.0 292050.0 ;
      RECT  127950.0 289800.0 128850.0 290700.0 ;
      RECT  123900.0 291150.0 128400.0 292050.0 ;
      RECT  127950.0 290250.0 128850.0 291600.0 ;
      RECT  128400.0 289800.0 132900.0 290700.0 ;
      RECT  103350.0 305100.0 108900.0 306000.0 ;
      RECT  111450.0 303750.0 112350.0 304650.0 ;
      RECT  111450.0 305100.0 112350.0 306000.0 ;
      RECT  111450.0 304200.0 112350.0 306000.0 ;
      RECT  111900.0 303750.0 118500.0 304650.0 ;
      RECT  118500.0 303750.0 119700.0 304650.0 ;
      RECT  127950.0 303750.0 128850.0 304650.0 ;
      RECT  127950.0 305100.0 128850.0 306000.0 ;
      RECT  123900.0 303750.0 128400.0 304650.0 ;
      RECT  127950.0 304200.0 128850.0 305550.0 ;
      RECT  128400.0 305100.0 132900.0 306000.0 ;
      RECT  103350.0 318000.0 108900.0 318900.0 ;
      RECT  111450.0 319350.0 112350.0 320250.0 ;
      RECT  111450.0 318000.0 112350.0 318900.0 ;
      RECT  111450.0 318900.0 112350.0 319800.0 ;
      RECT  111900.0 319350.0 118500.0 320250.0 ;
      RECT  118500.0 319350.0 119700.0 320250.0 ;
      RECT  127950.0 319350.0 128850.0 320250.0 ;
      RECT  127950.0 318000.0 128850.0 318900.0 ;
      RECT  123900.0 319350.0 128400.0 320250.0 ;
      RECT  127950.0 318450.0 128850.0 319800.0 ;
      RECT  128400.0 318000.0 132900.0 318900.0 ;
      RECT  103350.0 333300.0 108900.0 334200.0 ;
      RECT  111450.0 331950.0 112350.0 332850.0 ;
      RECT  111450.0 333300.0 112350.0 334200.0 ;
      RECT  111450.0 332400.0 112350.0 334200.0 ;
      RECT  111900.0 331950.0 118500.0 332850.0 ;
      RECT  118500.0 331950.0 119700.0 332850.0 ;
      RECT  127950.0 331950.0 128850.0 332850.0 ;
      RECT  127950.0 333300.0 128850.0 334200.0 ;
      RECT  123900.0 331950.0 128400.0 332850.0 ;
      RECT  127950.0 332400.0 128850.0 333750.0 ;
      RECT  128400.0 333300.0 132900.0 334200.0 ;
      RECT  103350.0 346200.0 108900.0 347100.0 ;
      RECT  111450.0 347550.0 112350.0 348450.0 ;
      RECT  111450.0 346200.0 112350.0 347100.0 ;
      RECT  111450.0 347100.0 112350.0 348000.0 ;
      RECT  111900.0 347550.0 118500.0 348450.0 ;
      RECT  118500.0 347550.0 119700.0 348450.0 ;
      RECT  127950.0 347550.0 128850.0 348450.0 ;
      RECT  127950.0 346200.0 128850.0 347100.0 ;
      RECT  123900.0 347550.0 128400.0 348450.0 ;
      RECT  127950.0 346650.0 128850.0 348000.0 ;
      RECT  128400.0 346200.0 132900.0 347100.0 ;
      RECT  103350.0 361500.0 108900.0 362400.0 ;
      RECT  111450.0 360150.0 112350.0 361050.0 ;
      RECT  111450.0 361500.0 112350.0 362400.0 ;
      RECT  111450.0 360600.0 112350.0 362400.0 ;
      RECT  111900.0 360150.0 118500.0 361050.0 ;
      RECT  118500.0 360150.0 119700.0 361050.0 ;
      RECT  127950.0 360150.0 128850.0 361050.0 ;
      RECT  127950.0 361500.0 128850.0 362400.0 ;
      RECT  123900.0 360150.0 128400.0 361050.0 ;
      RECT  127950.0 360600.0 128850.0 361950.0 ;
      RECT  128400.0 361500.0 132900.0 362400.0 ;
      RECT  103350.0 374400.0 108900.0 375300.0 ;
      RECT  111450.0 375750.0 112350.0 376650.0 ;
      RECT  111450.0 374400.0 112350.0 375300.0 ;
      RECT  111450.0 375300.0 112350.0 376200.0 ;
      RECT  111900.0 375750.0 118500.0 376650.0 ;
      RECT  118500.0 375750.0 119700.0 376650.0 ;
      RECT  127950.0 375750.0 128850.0 376650.0 ;
      RECT  127950.0 374400.0 128850.0 375300.0 ;
      RECT  123900.0 375750.0 128400.0 376650.0 ;
      RECT  127950.0 374850.0 128850.0 376200.0 ;
      RECT  128400.0 374400.0 132900.0 375300.0 ;
      RECT  103350.0 389700.0 108900.0 390600.0 ;
      RECT  111450.0 388350.0 112350.0 389250.0 ;
      RECT  111450.0 389700.0 112350.0 390600.0 ;
      RECT  111450.0 388800.0 112350.0 390600.0 ;
      RECT  111900.0 388350.0 118500.0 389250.0 ;
      RECT  118500.0 388350.0 119700.0 389250.0 ;
      RECT  127950.0 388350.0 128850.0 389250.0 ;
      RECT  127950.0 389700.0 128850.0 390600.0 ;
      RECT  123900.0 388350.0 128400.0 389250.0 ;
      RECT  127950.0 388800.0 128850.0 390150.0 ;
      RECT  128400.0 389700.0 132900.0 390600.0 ;
      RECT  103350.0 402600.0 108900.0 403500.0 ;
      RECT  111450.0 403950.0 112350.0 404850.0 ;
      RECT  111450.0 402600.0 112350.0 403500.0 ;
      RECT  111450.0 403500.0 112350.0 404400.0 ;
      RECT  111900.0 403950.0 118500.0 404850.0 ;
      RECT  118500.0 403950.0 119700.0 404850.0 ;
      RECT  127950.0 403950.0 128850.0 404850.0 ;
      RECT  127950.0 402600.0 128850.0 403500.0 ;
      RECT  123900.0 403950.0 128400.0 404850.0 ;
      RECT  127950.0 403050.0 128850.0 404400.0 ;
      RECT  128400.0 402600.0 132900.0 403500.0 ;
      RECT  103350.0 417900.0 108900.0 418800.0 ;
      RECT  111450.0 416550.0 112350.0 417450.0 ;
      RECT  111450.0 417900.0 112350.0 418800.0 ;
      RECT  111450.0 417000.0 112350.0 418800.0 ;
      RECT  111900.0 416550.0 118500.0 417450.0 ;
      RECT  118500.0 416550.0 119700.0 417450.0 ;
      RECT  127950.0 416550.0 128850.0 417450.0 ;
      RECT  127950.0 417900.0 128850.0 418800.0 ;
      RECT  123900.0 416550.0 128400.0 417450.0 ;
      RECT  127950.0 417000.0 128850.0 418350.0 ;
      RECT  128400.0 417900.0 132900.0 418800.0 ;
      RECT  113100.0 199200.0 114300.0 201150.0 ;
      RECT  113100.0 211350.0 114300.0 213300.0 ;
      RECT  108300.0 200550.0 109500.0 198750.0 ;
      RECT  108300.0 210150.0 109500.0 213750.0 ;
      RECT  111000.0 201750.0 111900.0 210150.0 ;
      RECT  108300.0 210150.0 109500.0 211350.0 ;
      RECT  110700.0 210150.0 111900.0 211350.0 ;
      RECT  110700.0 210150.0 111900.0 211350.0 ;
      RECT  108300.0 210150.0 109500.0 211350.0 ;
      RECT  108300.0 200550.0 109500.0 201750.0 ;
      RECT  110700.0 200550.0 111900.0 201750.0 ;
      RECT  110700.0 200550.0 111900.0 201750.0 ;
      RECT  108300.0 200550.0 109500.0 201750.0 ;
      RECT  113100.0 200550.0 114300.0 201750.0 ;
      RECT  113100.0 210750.0 114300.0 211950.0 ;
      RECT  108900.0 205050.0 110100.0 206250.0 ;
      RECT  108900.0 205050.0 110100.0 206250.0 ;
      RECT  111450.0 205200.0 112350.0 206100.0 ;
      RECT  106500.0 212850.0 116100.0 213750.0 ;
      RECT  106500.0 198750.0 116100.0 199650.0 ;
      RECT  125100.0 199200.0 126300.0 201150.0 ;
      RECT  125100.0 211350.0 126300.0 213300.0 ;
      RECT  117900.0 201150.0 119100.0 198750.0 ;
      RECT  117900.0 210150.0 119100.0 213750.0 ;
      RECT  122700.0 210150.0 123900.0 213750.0 ;
      RECT  117900.0 210150.0 119100.0 211350.0 ;
      RECT  120300.0 210150.0 121500.0 211350.0 ;
      RECT  120300.0 210150.0 121500.0 211350.0 ;
      RECT  117900.0 210150.0 119100.0 211350.0 ;
      RECT  120300.0 210150.0 121500.0 211350.0 ;
      RECT  122700.0 210150.0 123900.0 211350.0 ;
      RECT  122700.0 210150.0 123900.0 211350.0 ;
      RECT  120300.0 210150.0 121500.0 211350.0 ;
      RECT  117900.0 201150.0 119100.0 202350.0 ;
      RECT  120300.0 201150.0 121500.0 202350.0 ;
      RECT  120300.0 201150.0 121500.0 202350.0 ;
      RECT  117900.0 201150.0 119100.0 202350.0 ;
      RECT  120300.0 201150.0 121500.0 202350.0 ;
      RECT  122700.0 201150.0 123900.0 202350.0 ;
      RECT  122700.0 201150.0 123900.0 202350.0 ;
      RECT  120300.0 201150.0 121500.0 202350.0 ;
      RECT  125100.0 200550.0 126300.0 201750.0 ;
      RECT  125100.0 210750.0 126300.0 211950.0 ;
      RECT  122700.0 203700.0 121500.0 204900.0 ;
      RECT  119700.0 206400.0 118500.0 207600.0 ;
      RECT  120300.0 210150.0 121500.0 211350.0 ;
      RECT  122700.0 201150.0 123900.0 202350.0 ;
      RECT  123900.0 206400.0 122700.0 207600.0 ;
      RECT  118500.0 206400.0 119700.0 207600.0 ;
      RECT  121500.0 203700.0 122700.0 204900.0 ;
      RECT  122700.0 206400.0 123900.0 207600.0 ;
      RECT  116100.0 212850.0 130500.0 213750.0 ;
      RECT  116100.0 198750.0 130500.0 199650.0 ;
      RECT  137100.0 199200.0 138300.0 201150.0 ;
      RECT  137100.0 211350.0 138300.0 213300.0 ;
      RECT  132300.0 200550.0 133500.0 198750.0 ;
      RECT  132300.0 210150.0 133500.0 213750.0 ;
      RECT  135000.0 201750.0 135900.0 210150.0 ;
      RECT  132300.0 210150.0 133500.0 211350.0 ;
      RECT  134700.0 210150.0 135900.0 211350.0 ;
      RECT  134700.0 210150.0 135900.0 211350.0 ;
      RECT  132300.0 210150.0 133500.0 211350.0 ;
      RECT  132300.0 200550.0 133500.0 201750.0 ;
      RECT  134700.0 200550.0 135900.0 201750.0 ;
      RECT  134700.0 200550.0 135900.0 201750.0 ;
      RECT  132300.0 200550.0 133500.0 201750.0 ;
      RECT  137100.0 200550.0 138300.0 201750.0 ;
      RECT  137100.0 210750.0 138300.0 211950.0 ;
      RECT  132900.0 205050.0 134100.0 206250.0 ;
      RECT  132900.0 205050.0 134100.0 206250.0 ;
      RECT  135450.0 205200.0 136350.0 206100.0 ;
      RECT  130500.0 212850.0 140100.0 213750.0 ;
      RECT  130500.0 198750.0 140100.0 199650.0 ;
      RECT  102750.0 205050.0 103950.0 206250.0 ;
      RECT  104700.0 202800.0 105900.0 204000.0 ;
      RECT  121500.0 203700.0 120300.0 204900.0 ;
      RECT  113100.0 227400.0 114300.0 225450.0 ;
      RECT  113100.0 215250.0 114300.0 213300.0 ;
      RECT  108300.0 226050.0 109500.0 227850.0 ;
      RECT  108300.0 216450.0 109500.0 212850.0 ;
      RECT  111000.0 224850.0 111900.0 216450.0 ;
      RECT  108300.0 216450.0 109500.0 215250.0 ;
      RECT  110700.0 216450.0 111900.0 215250.0 ;
      RECT  110700.0 216450.0 111900.0 215250.0 ;
      RECT  108300.0 216450.0 109500.0 215250.0 ;
      RECT  108300.0 226050.0 109500.0 224850.0 ;
      RECT  110700.0 226050.0 111900.0 224850.0 ;
      RECT  110700.0 226050.0 111900.0 224850.0 ;
      RECT  108300.0 226050.0 109500.0 224850.0 ;
      RECT  113100.0 226050.0 114300.0 224850.0 ;
      RECT  113100.0 215850.0 114300.0 214650.0 ;
      RECT  108900.0 221550.0 110100.0 220350.0 ;
      RECT  108900.0 221550.0 110100.0 220350.0 ;
      RECT  111450.0 221400.0 112350.0 220500.0 ;
      RECT  106500.0 213750.0 116100.0 212850.0 ;
      RECT  106500.0 227850.0 116100.0 226950.0 ;
      RECT  125100.0 227400.0 126300.0 225450.0 ;
      RECT  125100.0 215250.0 126300.0 213300.0 ;
      RECT  117900.0 225450.0 119100.0 227850.0 ;
      RECT  117900.0 216450.0 119100.0 212850.0 ;
      RECT  122700.0 216450.0 123900.0 212850.0 ;
      RECT  117900.0 216450.0 119100.0 215250.0 ;
      RECT  120300.0 216450.0 121500.0 215250.0 ;
      RECT  120300.0 216450.0 121500.0 215250.0 ;
      RECT  117900.0 216450.0 119100.0 215250.0 ;
      RECT  120300.0 216450.0 121500.0 215250.0 ;
      RECT  122700.0 216450.0 123900.0 215250.0 ;
      RECT  122700.0 216450.0 123900.0 215250.0 ;
      RECT  120300.0 216450.0 121500.0 215250.0 ;
      RECT  117900.0 225450.0 119100.0 224250.0 ;
      RECT  120300.0 225450.0 121500.0 224250.0 ;
      RECT  120300.0 225450.0 121500.0 224250.0 ;
      RECT  117900.0 225450.0 119100.0 224250.0 ;
      RECT  120300.0 225450.0 121500.0 224250.0 ;
      RECT  122700.0 225450.0 123900.0 224250.0 ;
      RECT  122700.0 225450.0 123900.0 224250.0 ;
      RECT  120300.0 225450.0 121500.0 224250.0 ;
      RECT  125100.0 226050.0 126300.0 224850.0 ;
      RECT  125100.0 215850.0 126300.0 214650.0 ;
      RECT  122700.0 222900.0 121500.0 221700.0 ;
      RECT  119700.0 220200.0 118500.0 219000.0 ;
      RECT  120300.0 216450.0 121500.0 215250.0 ;
      RECT  122700.0 225450.0 123900.0 224250.0 ;
      RECT  123900.0 220200.0 122700.0 219000.0 ;
      RECT  118500.0 220200.0 119700.0 219000.0 ;
      RECT  121500.0 222900.0 122700.0 221700.0 ;
      RECT  122700.0 220200.0 123900.0 219000.0 ;
      RECT  116100.0 213750.0 130500.0 212850.0 ;
      RECT  116100.0 227850.0 130500.0 226950.0 ;
      RECT  137100.0 227400.0 138300.0 225450.0 ;
      RECT  137100.0 215250.0 138300.0 213300.0 ;
      RECT  132300.0 226050.0 133500.0 227850.0 ;
      RECT  132300.0 216450.0 133500.0 212850.0 ;
      RECT  135000.0 224850.0 135900.0 216450.0 ;
      RECT  132300.0 216450.0 133500.0 215250.0 ;
      RECT  134700.0 216450.0 135900.0 215250.0 ;
      RECT  134700.0 216450.0 135900.0 215250.0 ;
      RECT  132300.0 216450.0 133500.0 215250.0 ;
      RECT  132300.0 226050.0 133500.0 224850.0 ;
      RECT  134700.0 226050.0 135900.0 224850.0 ;
      RECT  134700.0 226050.0 135900.0 224850.0 ;
      RECT  132300.0 226050.0 133500.0 224850.0 ;
      RECT  137100.0 226050.0 138300.0 224850.0 ;
      RECT  137100.0 215850.0 138300.0 214650.0 ;
      RECT  132900.0 221550.0 134100.0 220350.0 ;
      RECT  132900.0 221550.0 134100.0 220350.0 ;
      RECT  135450.0 221400.0 136350.0 220500.0 ;
      RECT  130500.0 213750.0 140100.0 212850.0 ;
      RECT  130500.0 227850.0 140100.0 226950.0 ;
      RECT  102750.0 220350.0 103950.0 221550.0 ;
      RECT  104700.0 222600.0 105900.0 223800.0 ;
      RECT  121500.0 221700.0 120300.0 222900.0 ;
      RECT  113100.0 227400.0 114300.0 229350.0 ;
      RECT  113100.0 239550.0 114300.0 241500.0 ;
      RECT  108300.0 228750.0 109500.0 226950.0 ;
      RECT  108300.0 238350.0 109500.0 241950.0 ;
      RECT  111000.0 229950.0 111900.0 238350.0 ;
      RECT  108300.0 238350.0 109500.0 239550.0 ;
      RECT  110700.0 238350.0 111900.0 239550.0 ;
      RECT  110700.0 238350.0 111900.0 239550.0 ;
      RECT  108300.0 238350.0 109500.0 239550.0 ;
      RECT  108300.0 228750.0 109500.0 229950.0 ;
      RECT  110700.0 228750.0 111900.0 229950.0 ;
      RECT  110700.0 228750.0 111900.0 229950.0 ;
      RECT  108300.0 228750.0 109500.0 229950.0 ;
      RECT  113100.0 228750.0 114300.0 229950.0 ;
      RECT  113100.0 238950.0 114300.0 240150.0 ;
      RECT  108900.0 233250.0 110100.0 234450.0 ;
      RECT  108900.0 233250.0 110100.0 234450.0 ;
      RECT  111450.0 233400.0 112350.0 234300.0 ;
      RECT  106500.0 241050.0 116100.0 241950.0 ;
      RECT  106500.0 226950.0 116100.0 227850.0 ;
      RECT  125100.0 227400.0 126300.0 229350.0 ;
      RECT  125100.0 239550.0 126300.0 241500.0 ;
      RECT  117900.0 229350.0 119100.0 226950.0 ;
      RECT  117900.0 238350.0 119100.0 241950.0 ;
      RECT  122700.0 238350.0 123900.0 241950.0 ;
      RECT  117900.0 238350.0 119100.0 239550.0 ;
      RECT  120300.0 238350.0 121500.0 239550.0 ;
      RECT  120300.0 238350.0 121500.0 239550.0 ;
      RECT  117900.0 238350.0 119100.0 239550.0 ;
      RECT  120300.0 238350.0 121500.0 239550.0 ;
      RECT  122700.0 238350.0 123900.0 239550.0 ;
      RECT  122700.0 238350.0 123900.0 239550.0 ;
      RECT  120300.0 238350.0 121500.0 239550.0 ;
      RECT  117900.0 229350.0 119100.0 230550.0 ;
      RECT  120300.0 229350.0 121500.0 230550.0 ;
      RECT  120300.0 229350.0 121500.0 230550.0 ;
      RECT  117900.0 229350.0 119100.0 230550.0 ;
      RECT  120300.0 229350.0 121500.0 230550.0 ;
      RECT  122700.0 229350.0 123900.0 230550.0 ;
      RECT  122700.0 229350.0 123900.0 230550.0 ;
      RECT  120300.0 229350.0 121500.0 230550.0 ;
      RECT  125100.0 228750.0 126300.0 229950.0 ;
      RECT  125100.0 238950.0 126300.0 240150.0 ;
      RECT  122700.0 231900.0 121500.0 233100.0 ;
      RECT  119700.0 234600.0 118500.0 235800.0 ;
      RECT  120300.0 238350.0 121500.0 239550.0 ;
      RECT  122700.0 229350.0 123900.0 230550.0 ;
      RECT  123900.0 234600.0 122700.0 235800.0 ;
      RECT  118500.0 234600.0 119700.0 235800.0 ;
      RECT  121500.0 231900.0 122700.0 233100.0 ;
      RECT  122700.0 234600.0 123900.0 235800.0 ;
      RECT  116100.0 241050.0 130500.0 241950.0 ;
      RECT  116100.0 226950.0 130500.0 227850.0 ;
      RECT  137100.0 227400.0 138300.0 229350.0 ;
      RECT  137100.0 239550.0 138300.0 241500.0 ;
      RECT  132300.0 228750.0 133500.0 226950.0 ;
      RECT  132300.0 238350.0 133500.0 241950.0 ;
      RECT  135000.0 229950.0 135900.0 238350.0 ;
      RECT  132300.0 238350.0 133500.0 239550.0 ;
      RECT  134700.0 238350.0 135900.0 239550.0 ;
      RECT  134700.0 238350.0 135900.0 239550.0 ;
      RECT  132300.0 238350.0 133500.0 239550.0 ;
      RECT  132300.0 228750.0 133500.0 229950.0 ;
      RECT  134700.0 228750.0 135900.0 229950.0 ;
      RECT  134700.0 228750.0 135900.0 229950.0 ;
      RECT  132300.0 228750.0 133500.0 229950.0 ;
      RECT  137100.0 228750.0 138300.0 229950.0 ;
      RECT  137100.0 238950.0 138300.0 240150.0 ;
      RECT  132900.0 233250.0 134100.0 234450.0 ;
      RECT  132900.0 233250.0 134100.0 234450.0 ;
      RECT  135450.0 233400.0 136350.0 234300.0 ;
      RECT  130500.0 241050.0 140100.0 241950.0 ;
      RECT  130500.0 226950.0 140100.0 227850.0 ;
      RECT  102750.0 233250.0 103950.0 234450.0 ;
      RECT  104700.0 231000.0 105900.0 232200.0 ;
      RECT  121500.0 231900.0 120300.0 233100.0 ;
      RECT  113100.0 255600.0 114300.0 253650.0 ;
      RECT  113100.0 243450.0 114300.0 241500.0 ;
      RECT  108300.0 254250.0 109500.0 256050.0 ;
      RECT  108300.0 244650.0 109500.0 241050.0 ;
      RECT  111000.0 253050.0 111900.0 244650.0 ;
      RECT  108300.0 244650.0 109500.0 243450.0 ;
      RECT  110700.0 244650.0 111900.0 243450.0 ;
      RECT  110700.0 244650.0 111900.0 243450.0 ;
      RECT  108300.0 244650.0 109500.0 243450.0 ;
      RECT  108300.0 254250.0 109500.0 253050.0 ;
      RECT  110700.0 254250.0 111900.0 253050.0 ;
      RECT  110700.0 254250.0 111900.0 253050.0 ;
      RECT  108300.0 254250.0 109500.0 253050.0 ;
      RECT  113100.0 254250.0 114300.0 253050.0 ;
      RECT  113100.0 244050.0 114300.0 242850.0 ;
      RECT  108900.0 249750.0 110100.0 248550.0 ;
      RECT  108900.0 249750.0 110100.0 248550.0 ;
      RECT  111450.0 249600.0 112350.0 248700.0 ;
      RECT  106500.0 241950.0 116100.0 241050.0 ;
      RECT  106500.0 256050.0 116100.0 255150.0 ;
      RECT  125100.0 255600.0 126300.0 253650.0 ;
      RECT  125100.0 243450.0 126300.0 241500.0 ;
      RECT  117900.0 253650.0 119100.0 256050.0 ;
      RECT  117900.0 244650.0 119100.0 241050.0 ;
      RECT  122700.0 244650.0 123900.0 241050.0 ;
      RECT  117900.0 244650.0 119100.0 243450.0 ;
      RECT  120300.0 244650.0 121500.0 243450.0 ;
      RECT  120300.0 244650.0 121500.0 243450.0 ;
      RECT  117900.0 244650.0 119100.0 243450.0 ;
      RECT  120300.0 244650.0 121500.0 243450.0 ;
      RECT  122700.0 244650.0 123900.0 243450.0 ;
      RECT  122700.0 244650.0 123900.0 243450.0 ;
      RECT  120300.0 244650.0 121500.0 243450.0 ;
      RECT  117900.0 253650.0 119100.0 252450.0 ;
      RECT  120300.0 253650.0 121500.0 252450.0 ;
      RECT  120300.0 253650.0 121500.0 252450.0 ;
      RECT  117900.0 253650.0 119100.0 252450.0 ;
      RECT  120300.0 253650.0 121500.0 252450.0 ;
      RECT  122700.0 253650.0 123900.0 252450.0 ;
      RECT  122700.0 253650.0 123900.0 252450.0 ;
      RECT  120300.0 253650.0 121500.0 252450.0 ;
      RECT  125100.0 254250.0 126300.0 253050.0 ;
      RECT  125100.0 244050.0 126300.0 242850.0 ;
      RECT  122700.0 251100.0 121500.0 249900.0 ;
      RECT  119700.0 248400.0 118500.0 247200.0 ;
      RECT  120300.0 244650.0 121500.0 243450.0 ;
      RECT  122700.0 253650.0 123900.0 252450.0 ;
      RECT  123900.0 248400.0 122700.0 247200.0 ;
      RECT  118500.0 248400.0 119700.0 247200.0 ;
      RECT  121500.0 251100.0 122700.0 249900.0 ;
      RECT  122700.0 248400.0 123900.0 247200.0 ;
      RECT  116100.0 241950.0 130500.0 241050.0 ;
      RECT  116100.0 256050.0 130500.0 255150.0 ;
      RECT  137100.0 255600.0 138300.0 253650.0 ;
      RECT  137100.0 243450.0 138300.0 241500.0 ;
      RECT  132300.0 254250.0 133500.0 256050.0 ;
      RECT  132300.0 244650.0 133500.0 241050.0 ;
      RECT  135000.0 253050.0 135900.0 244650.0 ;
      RECT  132300.0 244650.0 133500.0 243450.0 ;
      RECT  134700.0 244650.0 135900.0 243450.0 ;
      RECT  134700.0 244650.0 135900.0 243450.0 ;
      RECT  132300.0 244650.0 133500.0 243450.0 ;
      RECT  132300.0 254250.0 133500.0 253050.0 ;
      RECT  134700.0 254250.0 135900.0 253050.0 ;
      RECT  134700.0 254250.0 135900.0 253050.0 ;
      RECT  132300.0 254250.0 133500.0 253050.0 ;
      RECT  137100.0 254250.0 138300.0 253050.0 ;
      RECT  137100.0 244050.0 138300.0 242850.0 ;
      RECT  132900.0 249750.0 134100.0 248550.0 ;
      RECT  132900.0 249750.0 134100.0 248550.0 ;
      RECT  135450.0 249600.0 136350.0 248700.0 ;
      RECT  130500.0 241950.0 140100.0 241050.0 ;
      RECT  130500.0 256050.0 140100.0 255150.0 ;
      RECT  102750.0 248550.0 103950.0 249750.0 ;
      RECT  104700.0 250800.0 105900.0 252000.0 ;
      RECT  121500.0 249900.0 120300.0 251100.0 ;
      RECT  113100.0 255600.0 114300.0 257550.0 ;
      RECT  113100.0 267750.0 114300.0 269700.0 ;
      RECT  108300.0 256950.0 109500.0 255150.0 ;
      RECT  108300.0 266550.0 109500.0 270150.0 ;
      RECT  111000.0 258150.0 111900.0 266550.0 ;
      RECT  108300.0 266550.0 109500.0 267750.0 ;
      RECT  110700.0 266550.0 111900.0 267750.0 ;
      RECT  110700.0 266550.0 111900.0 267750.0 ;
      RECT  108300.0 266550.0 109500.0 267750.0 ;
      RECT  108300.0 256950.0 109500.0 258150.0 ;
      RECT  110700.0 256950.0 111900.0 258150.0 ;
      RECT  110700.0 256950.0 111900.0 258150.0 ;
      RECT  108300.0 256950.0 109500.0 258150.0 ;
      RECT  113100.0 256950.0 114300.0 258150.0 ;
      RECT  113100.0 267150.0 114300.0 268350.0 ;
      RECT  108900.0 261450.0 110100.0 262650.0 ;
      RECT  108900.0 261450.0 110100.0 262650.0 ;
      RECT  111450.0 261600.0 112350.0 262500.0 ;
      RECT  106500.0 269250.0 116100.0 270150.0 ;
      RECT  106500.0 255150.0 116100.0 256050.0 ;
      RECT  125100.0 255600.0 126300.0 257550.0 ;
      RECT  125100.0 267750.0 126300.0 269700.0 ;
      RECT  117900.0 257550.0 119100.0 255150.0 ;
      RECT  117900.0 266550.0 119100.0 270150.0 ;
      RECT  122700.0 266550.0 123900.0 270150.0 ;
      RECT  117900.0 266550.0 119100.0 267750.0 ;
      RECT  120300.0 266550.0 121500.0 267750.0 ;
      RECT  120300.0 266550.0 121500.0 267750.0 ;
      RECT  117900.0 266550.0 119100.0 267750.0 ;
      RECT  120300.0 266550.0 121500.0 267750.0 ;
      RECT  122700.0 266550.0 123900.0 267750.0 ;
      RECT  122700.0 266550.0 123900.0 267750.0 ;
      RECT  120300.0 266550.0 121500.0 267750.0 ;
      RECT  117900.0 257550.0 119100.0 258750.0 ;
      RECT  120300.0 257550.0 121500.0 258750.0 ;
      RECT  120300.0 257550.0 121500.0 258750.0 ;
      RECT  117900.0 257550.0 119100.0 258750.0 ;
      RECT  120300.0 257550.0 121500.0 258750.0 ;
      RECT  122700.0 257550.0 123900.0 258750.0 ;
      RECT  122700.0 257550.0 123900.0 258750.0 ;
      RECT  120300.0 257550.0 121500.0 258750.0 ;
      RECT  125100.0 256950.0 126300.0 258150.0 ;
      RECT  125100.0 267150.0 126300.0 268350.0 ;
      RECT  122700.0 260100.0 121500.0 261300.0 ;
      RECT  119700.0 262800.0 118500.0 264000.0 ;
      RECT  120300.0 266550.0 121500.0 267750.0 ;
      RECT  122700.0 257550.0 123900.0 258750.0 ;
      RECT  123900.0 262800.0 122700.0 264000.0 ;
      RECT  118500.0 262800.0 119700.0 264000.0 ;
      RECT  121500.0 260100.0 122700.0 261300.0 ;
      RECT  122700.0 262800.0 123900.0 264000.0 ;
      RECT  116100.0 269250.0 130500.0 270150.0 ;
      RECT  116100.0 255150.0 130500.0 256050.0 ;
      RECT  137100.0 255600.0 138300.0 257550.0 ;
      RECT  137100.0 267750.0 138300.0 269700.0 ;
      RECT  132300.0 256950.0 133500.0 255150.0 ;
      RECT  132300.0 266550.0 133500.0 270150.0 ;
      RECT  135000.0 258150.0 135900.0 266550.0 ;
      RECT  132300.0 266550.0 133500.0 267750.0 ;
      RECT  134700.0 266550.0 135900.0 267750.0 ;
      RECT  134700.0 266550.0 135900.0 267750.0 ;
      RECT  132300.0 266550.0 133500.0 267750.0 ;
      RECT  132300.0 256950.0 133500.0 258150.0 ;
      RECT  134700.0 256950.0 135900.0 258150.0 ;
      RECT  134700.0 256950.0 135900.0 258150.0 ;
      RECT  132300.0 256950.0 133500.0 258150.0 ;
      RECT  137100.0 256950.0 138300.0 258150.0 ;
      RECT  137100.0 267150.0 138300.0 268350.0 ;
      RECT  132900.0 261450.0 134100.0 262650.0 ;
      RECT  132900.0 261450.0 134100.0 262650.0 ;
      RECT  135450.0 261600.0 136350.0 262500.0 ;
      RECT  130500.0 269250.0 140100.0 270150.0 ;
      RECT  130500.0 255150.0 140100.0 256050.0 ;
      RECT  102750.0 261450.0 103950.0 262650.0 ;
      RECT  104700.0 259200.0 105900.0 260400.0 ;
      RECT  121500.0 260100.0 120300.0 261300.0 ;
      RECT  113100.0 283800.0 114300.0 281850.0 ;
      RECT  113100.0 271650.0 114300.0 269700.0 ;
      RECT  108300.0 282450.0 109500.0 284250.0 ;
      RECT  108300.0 272850.0 109500.0 269250.0 ;
      RECT  111000.0 281250.0 111900.0 272850.0 ;
      RECT  108300.0 272850.0 109500.0 271650.0 ;
      RECT  110700.0 272850.0 111900.0 271650.0 ;
      RECT  110700.0 272850.0 111900.0 271650.0 ;
      RECT  108300.0 272850.0 109500.0 271650.0 ;
      RECT  108300.0 282450.0 109500.0 281250.0 ;
      RECT  110700.0 282450.0 111900.0 281250.0 ;
      RECT  110700.0 282450.0 111900.0 281250.0 ;
      RECT  108300.0 282450.0 109500.0 281250.0 ;
      RECT  113100.0 282450.0 114300.0 281250.0 ;
      RECT  113100.0 272250.0 114300.0 271050.0 ;
      RECT  108900.0 277950.0 110100.0 276750.0 ;
      RECT  108900.0 277950.0 110100.0 276750.0 ;
      RECT  111450.0 277800.0 112350.0 276900.0 ;
      RECT  106500.0 270150.0 116100.0 269250.0 ;
      RECT  106500.0 284250.0 116100.0 283350.0 ;
      RECT  125100.0 283800.0 126300.0 281850.0 ;
      RECT  125100.0 271650.0 126300.0 269700.0 ;
      RECT  117900.0 281850.0 119100.0 284250.0 ;
      RECT  117900.0 272850.0 119100.0 269250.0 ;
      RECT  122700.0 272850.0 123900.0 269250.0 ;
      RECT  117900.0 272850.0 119100.0 271650.0 ;
      RECT  120300.0 272850.0 121500.0 271650.0 ;
      RECT  120300.0 272850.0 121500.0 271650.0 ;
      RECT  117900.0 272850.0 119100.0 271650.0 ;
      RECT  120300.0 272850.0 121500.0 271650.0 ;
      RECT  122700.0 272850.0 123900.0 271650.0 ;
      RECT  122700.0 272850.0 123900.0 271650.0 ;
      RECT  120300.0 272850.0 121500.0 271650.0 ;
      RECT  117900.0 281850.0 119100.0 280650.0 ;
      RECT  120300.0 281850.0 121500.0 280650.0 ;
      RECT  120300.0 281850.0 121500.0 280650.0 ;
      RECT  117900.0 281850.0 119100.0 280650.0 ;
      RECT  120300.0 281850.0 121500.0 280650.0 ;
      RECT  122700.0 281850.0 123900.0 280650.0 ;
      RECT  122700.0 281850.0 123900.0 280650.0 ;
      RECT  120300.0 281850.0 121500.0 280650.0 ;
      RECT  125100.0 282450.0 126300.0 281250.0 ;
      RECT  125100.0 272250.0 126300.0 271050.0 ;
      RECT  122700.0 279300.0 121500.0 278100.0 ;
      RECT  119700.0 276600.0 118500.0 275400.0 ;
      RECT  120300.0 272850.0 121500.0 271650.0 ;
      RECT  122700.0 281850.0 123900.0 280650.0 ;
      RECT  123900.0 276600.0 122700.0 275400.0 ;
      RECT  118500.0 276600.0 119700.0 275400.0 ;
      RECT  121500.0 279300.0 122700.0 278100.0 ;
      RECT  122700.0 276600.0 123900.0 275400.0 ;
      RECT  116100.0 270150.0 130500.0 269250.0 ;
      RECT  116100.0 284250.0 130500.0 283350.0 ;
      RECT  137100.0 283800.0 138300.0 281850.0 ;
      RECT  137100.0 271650.0 138300.0 269700.0 ;
      RECT  132300.0 282450.0 133500.0 284250.0 ;
      RECT  132300.0 272850.0 133500.0 269250.0 ;
      RECT  135000.0 281250.0 135900.0 272850.0 ;
      RECT  132300.0 272850.0 133500.0 271650.0 ;
      RECT  134700.0 272850.0 135900.0 271650.0 ;
      RECT  134700.0 272850.0 135900.0 271650.0 ;
      RECT  132300.0 272850.0 133500.0 271650.0 ;
      RECT  132300.0 282450.0 133500.0 281250.0 ;
      RECT  134700.0 282450.0 135900.0 281250.0 ;
      RECT  134700.0 282450.0 135900.0 281250.0 ;
      RECT  132300.0 282450.0 133500.0 281250.0 ;
      RECT  137100.0 282450.0 138300.0 281250.0 ;
      RECT  137100.0 272250.0 138300.0 271050.0 ;
      RECT  132900.0 277950.0 134100.0 276750.0 ;
      RECT  132900.0 277950.0 134100.0 276750.0 ;
      RECT  135450.0 277800.0 136350.0 276900.0 ;
      RECT  130500.0 270150.0 140100.0 269250.0 ;
      RECT  130500.0 284250.0 140100.0 283350.0 ;
      RECT  102750.0 276750.0 103950.0 277950.0 ;
      RECT  104700.0 279000.0 105900.0 280200.0 ;
      RECT  121500.0 278100.0 120300.0 279300.0 ;
      RECT  113100.0 283800.0 114300.0 285750.0 ;
      RECT  113100.0 295950.0 114300.0 297900.0 ;
      RECT  108300.0 285150.0 109500.0 283350.0 ;
      RECT  108300.0 294750.0 109500.0 298350.0 ;
      RECT  111000.0 286350.0 111900.0 294750.0 ;
      RECT  108300.0 294750.0 109500.0 295950.0 ;
      RECT  110700.0 294750.0 111900.0 295950.0 ;
      RECT  110700.0 294750.0 111900.0 295950.0 ;
      RECT  108300.0 294750.0 109500.0 295950.0 ;
      RECT  108300.0 285150.0 109500.0 286350.0 ;
      RECT  110700.0 285150.0 111900.0 286350.0 ;
      RECT  110700.0 285150.0 111900.0 286350.0 ;
      RECT  108300.0 285150.0 109500.0 286350.0 ;
      RECT  113100.0 285150.0 114300.0 286350.0 ;
      RECT  113100.0 295350.0 114300.0 296550.0 ;
      RECT  108900.0 289650.0 110100.0 290850.0 ;
      RECT  108900.0 289650.0 110100.0 290850.0 ;
      RECT  111450.0 289800.0 112350.0 290700.0 ;
      RECT  106500.0 297450.0 116100.0 298350.0 ;
      RECT  106500.0 283350.0 116100.0 284250.0 ;
      RECT  125100.0 283800.0 126300.0 285750.0 ;
      RECT  125100.0 295950.0 126300.0 297900.0 ;
      RECT  117900.0 285750.0 119100.0 283350.0 ;
      RECT  117900.0 294750.0 119100.0 298350.0 ;
      RECT  122700.0 294750.0 123900.0 298350.0 ;
      RECT  117900.0 294750.0 119100.0 295950.0 ;
      RECT  120300.0 294750.0 121500.0 295950.0 ;
      RECT  120300.0 294750.0 121500.0 295950.0 ;
      RECT  117900.0 294750.0 119100.0 295950.0 ;
      RECT  120300.0 294750.0 121500.0 295950.0 ;
      RECT  122700.0 294750.0 123900.0 295950.0 ;
      RECT  122700.0 294750.0 123900.0 295950.0 ;
      RECT  120300.0 294750.0 121500.0 295950.0 ;
      RECT  117900.0 285750.0 119100.0 286950.0 ;
      RECT  120300.0 285750.0 121500.0 286950.0 ;
      RECT  120300.0 285750.0 121500.0 286950.0 ;
      RECT  117900.0 285750.0 119100.0 286950.0 ;
      RECT  120300.0 285750.0 121500.0 286950.0 ;
      RECT  122700.0 285750.0 123900.0 286950.0 ;
      RECT  122700.0 285750.0 123900.0 286950.0 ;
      RECT  120300.0 285750.0 121500.0 286950.0 ;
      RECT  125100.0 285150.0 126300.0 286350.0 ;
      RECT  125100.0 295350.0 126300.0 296550.0 ;
      RECT  122700.0 288300.0 121500.0 289500.0 ;
      RECT  119700.0 291000.0 118500.0 292200.0 ;
      RECT  120300.0 294750.0 121500.0 295950.0 ;
      RECT  122700.0 285750.0 123900.0 286950.0 ;
      RECT  123900.0 291000.0 122700.0 292200.0 ;
      RECT  118500.0 291000.0 119700.0 292200.0 ;
      RECT  121500.0 288300.0 122700.0 289500.0 ;
      RECT  122700.0 291000.0 123900.0 292200.0 ;
      RECT  116100.0 297450.0 130500.0 298350.0 ;
      RECT  116100.0 283350.0 130500.0 284250.0 ;
      RECT  137100.0 283800.0 138300.0 285750.0 ;
      RECT  137100.0 295950.0 138300.0 297900.0 ;
      RECT  132300.0 285150.0 133500.0 283350.0 ;
      RECT  132300.0 294750.0 133500.0 298350.0 ;
      RECT  135000.0 286350.0 135900.0 294750.0 ;
      RECT  132300.0 294750.0 133500.0 295950.0 ;
      RECT  134700.0 294750.0 135900.0 295950.0 ;
      RECT  134700.0 294750.0 135900.0 295950.0 ;
      RECT  132300.0 294750.0 133500.0 295950.0 ;
      RECT  132300.0 285150.0 133500.0 286350.0 ;
      RECT  134700.0 285150.0 135900.0 286350.0 ;
      RECT  134700.0 285150.0 135900.0 286350.0 ;
      RECT  132300.0 285150.0 133500.0 286350.0 ;
      RECT  137100.0 285150.0 138300.0 286350.0 ;
      RECT  137100.0 295350.0 138300.0 296550.0 ;
      RECT  132900.0 289650.0 134100.0 290850.0 ;
      RECT  132900.0 289650.0 134100.0 290850.0 ;
      RECT  135450.0 289800.0 136350.0 290700.0 ;
      RECT  130500.0 297450.0 140100.0 298350.0 ;
      RECT  130500.0 283350.0 140100.0 284250.0 ;
      RECT  102750.0 289650.0 103950.0 290850.0 ;
      RECT  104700.0 287400.0 105900.0 288600.0 ;
      RECT  121500.0 288300.0 120300.0 289500.0 ;
      RECT  113100.0 312000.0 114300.0 310050.0 ;
      RECT  113100.0 299850.0 114300.0 297900.0 ;
      RECT  108300.0 310650.0 109500.0 312450.0 ;
      RECT  108300.0 301050.0 109500.0 297450.0 ;
      RECT  111000.0 309450.0 111900.0 301050.0 ;
      RECT  108300.0 301050.0 109500.0 299850.0 ;
      RECT  110700.0 301050.0 111900.0 299850.0 ;
      RECT  110700.0 301050.0 111900.0 299850.0 ;
      RECT  108300.0 301050.0 109500.0 299850.0 ;
      RECT  108300.0 310650.0 109500.0 309450.0 ;
      RECT  110700.0 310650.0 111900.0 309450.0 ;
      RECT  110700.0 310650.0 111900.0 309450.0 ;
      RECT  108300.0 310650.0 109500.0 309450.0 ;
      RECT  113100.0 310650.0 114300.0 309450.0 ;
      RECT  113100.0 300450.0 114300.0 299250.0 ;
      RECT  108900.0 306150.0 110100.0 304950.0 ;
      RECT  108900.0 306150.0 110100.0 304950.0 ;
      RECT  111450.0 306000.0 112350.0 305100.0 ;
      RECT  106500.0 298350.0 116100.0 297450.0 ;
      RECT  106500.0 312450.0 116100.0 311550.0 ;
      RECT  125100.0 312000.0 126300.0 310050.0 ;
      RECT  125100.0 299850.0 126300.0 297900.0 ;
      RECT  117900.0 310050.0 119100.0 312450.0 ;
      RECT  117900.0 301050.0 119100.0 297450.0 ;
      RECT  122700.0 301050.0 123900.0 297450.0 ;
      RECT  117900.0 301050.0 119100.0 299850.0 ;
      RECT  120300.0 301050.0 121500.0 299850.0 ;
      RECT  120300.0 301050.0 121500.0 299850.0 ;
      RECT  117900.0 301050.0 119100.0 299850.0 ;
      RECT  120300.0 301050.0 121500.0 299850.0 ;
      RECT  122700.0 301050.0 123900.0 299850.0 ;
      RECT  122700.0 301050.0 123900.0 299850.0 ;
      RECT  120300.0 301050.0 121500.0 299850.0 ;
      RECT  117900.0 310050.0 119100.0 308850.0 ;
      RECT  120300.0 310050.0 121500.0 308850.0 ;
      RECT  120300.0 310050.0 121500.0 308850.0 ;
      RECT  117900.0 310050.0 119100.0 308850.0 ;
      RECT  120300.0 310050.0 121500.0 308850.0 ;
      RECT  122700.0 310050.0 123900.0 308850.0 ;
      RECT  122700.0 310050.0 123900.0 308850.0 ;
      RECT  120300.0 310050.0 121500.0 308850.0 ;
      RECT  125100.0 310650.0 126300.0 309450.0 ;
      RECT  125100.0 300450.0 126300.0 299250.0 ;
      RECT  122700.0 307500.0 121500.0 306300.0 ;
      RECT  119700.0 304800.0 118500.0 303600.0 ;
      RECT  120300.0 301050.0 121500.0 299850.0 ;
      RECT  122700.0 310050.0 123900.0 308850.0 ;
      RECT  123900.0 304800.0 122700.0 303600.0 ;
      RECT  118500.0 304800.0 119700.0 303600.0 ;
      RECT  121500.0 307500.0 122700.0 306300.0 ;
      RECT  122700.0 304800.0 123900.0 303600.0 ;
      RECT  116100.0 298350.0 130500.0 297450.0 ;
      RECT  116100.0 312450.0 130500.0 311550.0 ;
      RECT  137100.0 312000.0 138300.0 310050.0 ;
      RECT  137100.0 299850.0 138300.0 297900.0 ;
      RECT  132300.0 310650.0 133500.0 312450.0 ;
      RECT  132300.0 301050.0 133500.0 297450.0 ;
      RECT  135000.0 309450.0 135900.0 301050.0 ;
      RECT  132300.0 301050.0 133500.0 299850.0 ;
      RECT  134700.0 301050.0 135900.0 299850.0 ;
      RECT  134700.0 301050.0 135900.0 299850.0 ;
      RECT  132300.0 301050.0 133500.0 299850.0 ;
      RECT  132300.0 310650.0 133500.0 309450.0 ;
      RECT  134700.0 310650.0 135900.0 309450.0 ;
      RECT  134700.0 310650.0 135900.0 309450.0 ;
      RECT  132300.0 310650.0 133500.0 309450.0 ;
      RECT  137100.0 310650.0 138300.0 309450.0 ;
      RECT  137100.0 300450.0 138300.0 299250.0 ;
      RECT  132900.0 306150.0 134100.0 304950.0 ;
      RECT  132900.0 306150.0 134100.0 304950.0 ;
      RECT  135450.0 306000.0 136350.0 305100.0 ;
      RECT  130500.0 298350.0 140100.0 297450.0 ;
      RECT  130500.0 312450.0 140100.0 311550.0 ;
      RECT  102750.0 304950.0 103950.0 306150.0 ;
      RECT  104700.0 307200.0 105900.0 308400.0 ;
      RECT  121500.0 306300.0 120300.0 307500.0 ;
      RECT  113100.0 312000.0 114300.0 313950.0 ;
      RECT  113100.0 324150.0 114300.0 326100.0 ;
      RECT  108300.0 313350.0 109500.0 311550.0 ;
      RECT  108300.0 322950.0 109500.0 326550.0 ;
      RECT  111000.0 314550.0 111900.0 322950.0 ;
      RECT  108300.0 322950.0 109500.0 324150.0 ;
      RECT  110700.0 322950.0 111900.0 324150.0 ;
      RECT  110700.0 322950.0 111900.0 324150.0 ;
      RECT  108300.0 322950.0 109500.0 324150.0 ;
      RECT  108300.0 313350.0 109500.0 314550.0 ;
      RECT  110700.0 313350.0 111900.0 314550.0 ;
      RECT  110700.0 313350.0 111900.0 314550.0 ;
      RECT  108300.0 313350.0 109500.0 314550.0 ;
      RECT  113100.0 313350.0 114300.0 314550.0 ;
      RECT  113100.0 323550.0 114300.0 324750.0 ;
      RECT  108900.0 317850.0 110100.0 319050.0 ;
      RECT  108900.0 317850.0 110100.0 319050.0 ;
      RECT  111450.0 318000.0 112350.0 318900.0 ;
      RECT  106500.0 325650.0 116100.0 326550.0 ;
      RECT  106500.0 311550.0 116100.0 312450.0 ;
      RECT  125100.0 312000.0 126300.0 313950.0 ;
      RECT  125100.0 324150.0 126300.0 326100.0 ;
      RECT  117900.0 313950.0 119100.0 311550.0 ;
      RECT  117900.0 322950.0 119100.0 326550.0 ;
      RECT  122700.0 322950.0 123900.0 326550.0 ;
      RECT  117900.0 322950.0 119100.0 324150.0 ;
      RECT  120300.0 322950.0 121500.0 324150.0 ;
      RECT  120300.0 322950.0 121500.0 324150.0 ;
      RECT  117900.0 322950.0 119100.0 324150.0 ;
      RECT  120300.0 322950.0 121500.0 324150.0 ;
      RECT  122700.0 322950.0 123900.0 324150.0 ;
      RECT  122700.0 322950.0 123900.0 324150.0 ;
      RECT  120300.0 322950.0 121500.0 324150.0 ;
      RECT  117900.0 313950.0 119100.0 315150.0 ;
      RECT  120300.0 313950.0 121500.0 315150.0 ;
      RECT  120300.0 313950.0 121500.0 315150.0 ;
      RECT  117900.0 313950.0 119100.0 315150.0 ;
      RECT  120300.0 313950.0 121500.0 315150.0 ;
      RECT  122700.0 313950.0 123900.0 315150.0 ;
      RECT  122700.0 313950.0 123900.0 315150.0 ;
      RECT  120300.0 313950.0 121500.0 315150.0 ;
      RECT  125100.0 313350.0 126300.0 314550.0 ;
      RECT  125100.0 323550.0 126300.0 324750.0 ;
      RECT  122700.0 316500.0 121500.0 317700.0 ;
      RECT  119700.0 319200.0 118500.0 320400.0 ;
      RECT  120300.0 322950.0 121500.0 324150.0 ;
      RECT  122700.0 313950.0 123900.0 315150.0 ;
      RECT  123900.0 319200.0 122700.0 320400.0 ;
      RECT  118500.0 319200.0 119700.0 320400.0 ;
      RECT  121500.0 316500.0 122700.0 317700.0 ;
      RECT  122700.0 319200.0 123900.0 320400.0 ;
      RECT  116100.0 325650.0 130500.0 326550.0 ;
      RECT  116100.0 311550.0 130500.0 312450.0 ;
      RECT  137100.0 312000.0 138300.0 313950.0 ;
      RECT  137100.0 324150.0 138300.0 326100.0 ;
      RECT  132300.0 313350.0 133500.0 311550.0 ;
      RECT  132300.0 322950.0 133500.0 326550.0 ;
      RECT  135000.0 314550.0 135900.0 322950.0 ;
      RECT  132300.0 322950.0 133500.0 324150.0 ;
      RECT  134700.0 322950.0 135900.0 324150.0 ;
      RECT  134700.0 322950.0 135900.0 324150.0 ;
      RECT  132300.0 322950.0 133500.0 324150.0 ;
      RECT  132300.0 313350.0 133500.0 314550.0 ;
      RECT  134700.0 313350.0 135900.0 314550.0 ;
      RECT  134700.0 313350.0 135900.0 314550.0 ;
      RECT  132300.0 313350.0 133500.0 314550.0 ;
      RECT  137100.0 313350.0 138300.0 314550.0 ;
      RECT  137100.0 323550.0 138300.0 324750.0 ;
      RECT  132900.0 317850.0 134100.0 319050.0 ;
      RECT  132900.0 317850.0 134100.0 319050.0 ;
      RECT  135450.0 318000.0 136350.0 318900.0 ;
      RECT  130500.0 325650.0 140100.0 326550.0 ;
      RECT  130500.0 311550.0 140100.0 312450.0 ;
      RECT  102750.0 317850.0 103950.0 319050.0 ;
      RECT  104700.0 315600.0 105900.0 316800.0 ;
      RECT  121500.0 316500.0 120300.0 317700.0 ;
      RECT  113100.0 340200.0 114300.0 338250.0 ;
      RECT  113100.0 328050.0 114300.0 326100.0 ;
      RECT  108300.0 338850.0 109500.0 340650.0 ;
      RECT  108300.0 329250.0 109500.0 325650.0 ;
      RECT  111000.0 337650.0 111900.0 329250.0 ;
      RECT  108300.0 329250.0 109500.0 328050.0 ;
      RECT  110700.0 329250.0 111900.0 328050.0 ;
      RECT  110700.0 329250.0 111900.0 328050.0 ;
      RECT  108300.0 329250.0 109500.0 328050.0 ;
      RECT  108300.0 338850.0 109500.0 337650.0 ;
      RECT  110700.0 338850.0 111900.0 337650.0 ;
      RECT  110700.0 338850.0 111900.0 337650.0 ;
      RECT  108300.0 338850.0 109500.0 337650.0 ;
      RECT  113100.0 338850.0 114300.0 337650.0 ;
      RECT  113100.0 328650.0 114300.0 327450.0 ;
      RECT  108900.0 334350.0 110100.0 333150.0 ;
      RECT  108900.0 334350.0 110100.0 333150.0 ;
      RECT  111450.0 334200.0 112350.0 333300.0 ;
      RECT  106500.0 326550.0 116100.0 325650.0 ;
      RECT  106500.0 340650.0 116100.0 339750.0 ;
      RECT  125100.0 340200.0 126300.0 338250.0 ;
      RECT  125100.0 328050.0 126300.0 326100.0 ;
      RECT  117900.0 338250.0 119100.0 340650.0 ;
      RECT  117900.0 329250.0 119100.0 325650.0 ;
      RECT  122700.0 329250.0 123900.0 325650.0 ;
      RECT  117900.0 329250.0 119100.0 328050.0 ;
      RECT  120300.0 329250.0 121500.0 328050.0 ;
      RECT  120300.0 329250.0 121500.0 328050.0 ;
      RECT  117900.0 329250.0 119100.0 328050.0 ;
      RECT  120300.0 329250.0 121500.0 328050.0 ;
      RECT  122700.0 329250.0 123900.0 328050.0 ;
      RECT  122700.0 329250.0 123900.0 328050.0 ;
      RECT  120300.0 329250.0 121500.0 328050.0 ;
      RECT  117900.0 338250.0 119100.0 337050.0 ;
      RECT  120300.0 338250.0 121500.0 337050.0 ;
      RECT  120300.0 338250.0 121500.0 337050.0 ;
      RECT  117900.0 338250.0 119100.0 337050.0 ;
      RECT  120300.0 338250.0 121500.0 337050.0 ;
      RECT  122700.0 338250.0 123900.0 337050.0 ;
      RECT  122700.0 338250.0 123900.0 337050.0 ;
      RECT  120300.0 338250.0 121500.0 337050.0 ;
      RECT  125100.0 338850.0 126300.0 337650.0 ;
      RECT  125100.0 328650.0 126300.0 327450.0 ;
      RECT  122700.0 335700.0 121500.0 334500.0 ;
      RECT  119700.0 333000.0 118500.0 331800.0 ;
      RECT  120300.0 329250.0 121500.0 328050.0 ;
      RECT  122700.0 338250.0 123900.0 337050.0 ;
      RECT  123900.0 333000.0 122700.0 331800.0 ;
      RECT  118500.0 333000.0 119700.0 331800.0 ;
      RECT  121500.0 335700.0 122700.0 334500.0 ;
      RECT  122700.0 333000.0 123900.0 331800.0 ;
      RECT  116100.0 326550.0 130500.0 325650.0 ;
      RECT  116100.0 340650.0 130500.0 339750.0 ;
      RECT  137100.0 340200.0 138300.0 338250.0 ;
      RECT  137100.0 328050.0 138300.0 326100.0 ;
      RECT  132300.0 338850.0 133500.0 340650.0 ;
      RECT  132300.0 329250.0 133500.0 325650.0 ;
      RECT  135000.0 337650.0 135900.0 329250.0 ;
      RECT  132300.0 329250.0 133500.0 328050.0 ;
      RECT  134700.0 329250.0 135900.0 328050.0 ;
      RECT  134700.0 329250.0 135900.0 328050.0 ;
      RECT  132300.0 329250.0 133500.0 328050.0 ;
      RECT  132300.0 338850.0 133500.0 337650.0 ;
      RECT  134700.0 338850.0 135900.0 337650.0 ;
      RECT  134700.0 338850.0 135900.0 337650.0 ;
      RECT  132300.0 338850.0 133500.0 337650.0 ;
      RECT  137100.0 338850.0 138300.0 337650.0 ;
      RECT  137100.0 328650.0 138300.0 327450.0 ;
      RECT  132900.0 334350.0 134100.0 333150.0 ;
      RECT  132900.0 334350.0 134100.0 333150.0 ;
      RECT  135450.0 334200.0 136350.0 333300.0 ;
      RECT  130500.0 326550.0 140100.0 325650.0 ;
      RECT  130500.0 340650.0 140100.0 339750.0 ;
      RECT  102750.0 333150.0 103950.0 334350.0 ;
      RECT  104700.0 335400.0 105900.0 336600.0 ;
      RECT  121500.0 334500.0 120300.0 335700.0 ;
      RECT  113100.0 340200.0 114300.0 342150.0 ;
      RECT  113100.0 352350.0 114300.0 354300.0 ;
      RECT  108300.0 341550.0 109500.0 339750.0 ;
      RECT  108300.0 351150.0 109500.0 354750.0 ;
      RECT  111000.0 342750.0 111900.0 351150.0 ;
      RECT  108300.0 351150.0 109500.0 352350.0 ;
      RECT  110700.0 351150.0 111900.0 352350.0 ;
      RECT  110700.0 351150.0 111900.0 352350.0 ;
      RECT  108300.0 351150.0 109500.0 352350.0 ;
      RECT  108300.0 341550.0 109500.0 342750.0 ;
      RECT  110700.0 341550.0 111900.0 342750.0 ;
      RECT  110700.0 341550.0 111900.0 342750.0 ;
      RECT  108300.0 341550.0 109500.0 342750.0 ;
      RECT  113100.0 341550.0 114300.0 342750.0 ;
      RECT  113100.0 351750.0 114300.0 352950.0 ;
      RECT  108900.0 346050.0 110100.0 347250.0 ;
      RECT  108900.0 346050.0 110100.0 347250.0 ;
      RECT  111450.0 346200.0 112350.0 347100.0 ;
      RECT  106500.0 353850.0 116100.0 354750.0 ;
      RECT  106500.0 339750.0 116100.0 340650.0 ;
      RECT  125100.0 340200.0 126300.0 342150.0 ;
      RECT  125100.0 352350.0 126300.0 354300.0 ;
      RECT  117900.0 342150.0 119100.0 339750.0 ;
      RECT  117900.0 351150.0 119100.0 354750.0 ;
      RECT  122700.0 351150.0 123900.0 354750.0 ;
      RECT  117900.0 351150.0 119100.0 352350.0 ;
      RECT  120300.0 351150.0 121500.0 352350.0 ;
      RECT  120300.0 351150.0 121500.0 352350.0 ;
      RECT  117900.0 351150.0 119100.0 352350.0 ;
      RECT  120300.0 351150.0 121500.0 352350.0 ;
      RECT  122700.0 351150.0 123900.0 352350.0 ;
      RECT  122700.0 351150.0 123900.0 352350.0 ;
      RECT  120300.0 351150.0 121500.0 352350.0 ;
      RECT  117900.0 342150.0 119100.0 343350.0 ;
      RECT  120300.0 342150.0 121500.0 343350.0 ;
      RECT  120300.0 342150.0 121500.0 343350.0 ;
      RECT  117900.0 342150.0 119100.0 343350.0 ;
      RECT  120300.0 342150.0 121500.0 343350.0 ;
      RECT  122700.0 342150.0 123900.0 343350.0 ;
      RECT  122700.0 342150.0 123900.0 343350.0 ;
      RECT  120300.0 342150.0 121500.0 343350.0 ;
      RECT  125100.0 341550.0 126300.0 342750.0 ;
      RECT  125100.0 351750.0 126300.0 352950.0 ;
      RECT  122700.0 344700.0 121500.0 345900.0 ;
      RECT  119700.0 347400.0 118500.0 348600.0 ;
      RECT  120300.0 351150.0 121500.0 352350.0 ;
      RECT  122700.0 342150.0 123900.0 343350.0 ;
      RECT  123900.0 347400.0 122700.0 348600.0 ;
      RECT  118500.0 347400.0 119700.0 348600.0 ;
      RECT  121500.0 344700.0 122700.0 345900.0 ;
      RECT  122700.0 347400.0 123900.0 348600.0 ;
      RECT  116100.0 353850.0 130500.0 354750.0 ;
      RECT  116100.0 339750.0 130500.0 340650.0 ;
      RECT  137100.0 340200.0 138300.0 342150.0 ;
      RECT  137100.0 352350.0 138300.0 354300.0 ;
      RECT  132300.0 341550.0 133500.0 339750.0 ;
      RECT  132300.0 351150.0 133500.0 354750.0 ;
      RECT  135000.0 342750.0 135900.0 351150.0 ;
      RECT  132300.0 351150.0 133500.0 352350.0 ;
      RECT  134700.0 351150.0 135900.0 352350.0 ;
      RECT  134700.0 351150.0 135900.0 352350.0 ;
      RECT  132300.0 351150.0 133500.0 352350.0 ;
      RECT  132300.0 341550.0 133500.0 342750.0 ;
      RECT  134700.0 341550.0 135900.0 342750.0 ;
      RECT  134700.0 341550.0 135900.0 342750.0 ;
      RECT  132300.0 341550.0 133500.0 342750.0 ;
      RECT  137100.0 341550.0 138300.0 342750.0 ;
      RECT  137100.0 351750.0 138300.0 352950.0 ;
      RECT  132900.0 346050.0 134100.0 347250.0 ;
      RECT  132900.0 346050.0 134100.0 347250.0 ;
      RECT  135450.0 346200.0 136350.0 347100.0 ;
      RECT  130500.0 353850.0 140100.0 354750.0 ;
      RECT  130500.0 339750.0 140100.0 340650.0 ;
      RECT  102750.0 346050.0 103950.0 347250.0 ;
      RECT  104700.0 343800.0 105900.0 345000.0 ;
      RECT  121500.0 344700.0 120300.0 345900.0 ;
      RECT  113100.0 368400.0 114300.0 366450.0 ;
      RECT  113100.0 356250.0 114300.0 354300.0 ;
      RECT  108300.0 367050.0 109500.0 368850.0 ;
      RECT  108300.0 357450.0 109500.0 353850.0 ;
      RECT  111000.0 365850.0 111900.0 357450.0 ;
      RECT  108300.0 357450.0 109500.0 356250.0 ;
      RECT  110700.0 357450.0 111900.0 356250.0 ;
      RECT  110700.0 357450.0 111900.0 356250.0 ;
      RECT  108300.0 357450.0 109500.0 356250.0 ;
      RECT  108300.0 367050.0 109500.0 365850.0 ;
      RECT  110700.0 367050.0 111900.0 365850.0 ;
      RECT  110700.0 367050.0 111900.0 365850.0 ;
      RECT  108300.0 367050.0 109500.0 365850.0 ;
      RECT  113100.0 367050.0 114300.0 365850.0 ;
      RECT  113100.0 356850.0 114300.0 355650.0 ;
      RECT  108900.0 362550.0 110100.0 361350.0 ;
      RECT  108900.0 362550.0 110100.0 361350.0 ;
      RECT  111450.0 362400.0 112350.0 361500.0 ;
      RECT  106500.0 354750.0 116100.0 353850.0 ;
      RECT  106500.0 368850.0 116100.0 367950.0 ;
      RECT  125100.0 368400.0 126300.0 366450.0 ;
      RECT  125100.0 356250.0 126300.0 354300.0 ;
      RECT  117900.0 366450.0 119100.0 368850.0 ;
      RECT  117900.0 357450.0 119100.0 353850.0 ;
      RECT  122700.0 357450.0 123900.0 353850.0 ;
      RECT  117900.0 357450.0 119100.0 356250.0 ;
      RECT  120300.0 357450.0 121500.0 356250.0 ;
      RECT  120300.0 357450.0 121500.0 356250.0 ;
      RECT  117900.0 357450.0 119100.0 356250.0 ;
      RECT  120300.0 357450.0 121500.0 356250.0 ;
      RECT  122700.0 357450.0 123900.0 356250.0 ;
      RECT  122700.0 357450.0 123900.0 356250.0 ;
      RECT  120300.0 357450.0 121500.0 356250.0 ;
      RECT  117900.0 366450.0 119100.0 365250.0 ;
      RECT  120300.0 366450.0 121500.0 365250.0 ;
      RECT  120300.0 366450.0 121500.0 365250.0 ;
      RECT  117900.0 366450.0 119100.0 365250.0 ;
      RECT  120300.0 366450.0 121500.0 365250.0 ;
      RECT  122700.0 366450.0 123900.0 365250.0 ;
      RECT  122700.0 366450.0 123900.0 365250.0 ;
      RECT  120300.0 366450.0 121500.0 365250.0 ;
      RECT  125100.0 367050.0 126300.0 365850.0 ;
      RECT  125100.0 356850.0 126300.0 355650.0 ;
      RECT  122700.0 363900.0 121500.0 362700.0 ;
      RECT  119700.0 361200.0 118500.0 360000.0 ;
      RECT  120300.0 357450.0 121500.0 356250.0 ;
      RECT  122700.0 366450.0 123900.0 365250.0 ;
      RECT  123900.0 361200.0 122700.0 360000.0 ;
      RECT  118500.0 361200.0 119700.0 360000.0 ;
      RECT  121500.0 363900.0 122700.0 362700.0 ;
      RECT  122700.0 361200.0 123900.0 360000.0 ;
      RECT  116100.0 354750.0 130500.0 353850.0 ;
      RECT  116100.0 368850.0 130500.0 367950.0 ;
      RECT  137100.0 368400.0 138300.0 366450.0 ;
      RECT  137100.0 356250.0 138300.0 354300.0 ;
      RECT  132300.0 367050.0 133500.0 368850.0 ;
      RECT  132300.0 357450.0 133500.0 353850.0 ;
      RECT  135000.0 365850.0 135900.0 357450.0 ;
      RECT  132300.0 357450.0 133500.0 356250.0 ;
      RECT  134700.0 357450.0 135900.0 356250.0 ;
      RECT  134700.0 357450.0 135900.0 356250.0 ;
      RECT  132300.0 357450.0 133500.0 356250.0 ;
      RECT  132300.0 367050.0 133500.0 365850.0 ;
      RECT  134700.0 367050.0 135900.0 365850.0 ;
      RECT  134700.0 367050.0 135900.0 365850.0 ;
      RECT  132300.0 367050.0 133500.0 365850.0 ;
      RECT  137100.0 367050.0 138300.0 365850.0 ;
      RECT  137100.0 356850.0 138300.0 355650.0 ;
      RECT  132900.0 362550.0 134100.0 361350.0 ;
      RECT  132900.0 362550.0 134100.0 361350.0 ;
      RECT  135450.0 362400.0 136350.0 361500.0 ;
      RECT  130500.0 354750.0 140100.0 353850.0 ;
      RECT  130500.0 368850.0 140100.0 367950.0 ;
      RECT  102750.0 361350.0 103950.0 362550.0 ;
      RECT  104700.0 363600.0 105900.0 364800.0 ;
      RECT  121500.0 362700.0 120300.0 363900.0 ;
      RECT  113100.0 368400.0 114300.0 370350.0 ;
      RECT  113100.0 380550.0 114300.0 382500.0 ;
      RECT  108300.0 369750.0 109500.0 367950.0 ;
      RECT  108300.0 379350.0 109500.0 382950.0 ;
      RECT  111000.0 370950.0 111900.0 379350.0 ;
      RECT  108300.0 379350.0 109500.0 380550.0 ;
      RECT  110700.0 379350.0 111900.0 380550.0 ;
      RECT  110700.0 379350.0 111900.0 380550.0 ;
      RECT  108300.0 379350.0 109500.0 380550.0 ;
      RECT  108300.0 369750.0 109500.0 370950.0 ;
      RECT  110700.0 369750.0 111900.0 370950.0 ;
      RECT  110700.0 369750.0 111900.0 370950.0 ;
      RECT  108300.0 369750.0 109500.0 370950.0 ;
      RECT  113100.0 369750.0 114300.0 370950.0 ;
      RECT  113100.0 379950.0 114300.0 381150.0 ;
      RECT  108900.0 374250.0 110100.0 375450.0 ;
      RECT  108900.0 374250.0 110100.0 375450.0 ;
      RECT  111450.0 374400.0 112350.0 375300.0 ;
      RECT  106500.0 382050.0 116100.0 382950.0 ;
      RECT  106500.0 367950.0 116100.0 368850.0 ;
      RECT  125100.0 368400.0 126300.0 370350.0 ;
      RECT  125100.0 380550.0 126300.0 382500.0 ;
      RECT  117900.0 370350.0 119100.0 367950.0 ;
      RECT  117900.0 379350.0 119100.0 382950.0 ;
      RECT  122700.0 379350.0 123900.0 382950.0 ;
      RECT  117900.0 379350.0 119100.0 380550.0 ;
      RECT  120300.0 379350.0 121500.0 380550.0 ;
      RECT  120300.0 379350.0 121500.0 380550.0 ;
      RECT  117900.0 379350.0 119100.0 380550.0 ;
      RECT  120300.0 379350.0 121500.0 380550.0 ;
      RECT  122700.0 379350.0 123900.0 380550.0 ;
      RECT  122700.0 379350.0 123900.0 380550.0 ;
      RECT  120300.0 379350.0 121500.0 380550.0 ;
      RECT  117900.0 370350.0 119100.0 371550.0 ;
      RECT  120300.0 370350.0 121500.0 371550.0 ;
      RECT  120300.0 370350.0 121500.0 371550.0 ;
      RECT  117900.0 370350.0 119100.0 371550.0 ;
      RECT  120300.0 370350.0 121500.0 371550.0 ;
      RECT  122700.0 370350.0 123900.0 371550.0 ;
      RECT  122700.0 370350.0 123900.0 371550.0 ;
      RECT  120300.0 370350.0 121500.0 371550.0 ;
      RECT  125100.0 369750.0 126300.0 370950.0 ;
      RECT  125100.0 379950.0 126300.0 381150.0 ;
      RECT  122700.0 372900.0 121500.0 374100.0 ;
      RECT  119700.0 375600.0 118500.0 376800.0 ;
      RECT  120300.0 379350.0 121500.0 380550.0 ;
      RECT  122700.0 370350.0 123900.0 371550.0 ;
      RECT  123900.0 375600.0 122700.0 376800.0 ;
      RECT  118500.0 375600.0 119700.0 376800.0 ;
      RECT  121500.0 372900.0 122700.0 374100.0 ;
      RECT  122700.0 375600.0 123900.0 376800.0 ;
      RECT  116100.0 382050.0 130500.0 382950.0 ;
      RECT  116100.0 367950.0 130500.0 368850.0 ;
      RECT  137100.0 368400.0 138300.0 370350.0 ;
      RECT  137100.0 380550.0 138300.0 382500.0 ;
      RECT  132300.0 369750.0 133500.0 367950.0 ;
      RECT  132300.0 379350.0 133500.0 382950.0 ;
      RECT  135000.0 370950.0 135900.0 379350.0 ;
      RECT  132300.0 379350.0 133500.0 380550.0 ;
      RECT  134700.0 379350.0 135900.0 380550.0 ;
      RECT  134700.0 379350.0 135900.0 380550.0 ;
      RECT  132300.0 379350.0 133500.0 380550.0 ;
      RECT  132300.0 369750.0 133500.0 370950.0 ;
      RECT  134700.0 369750.0 135900.0 370950.0 ;
      RECT  134700.0 369750.0 135900.0 370950.0 ;
      RECT  132300.0 369750.0 133500.0 370950.0 ;
      RECT  137100.0 369750.0 138300.0 370950.0 ;
      RECT  137100.0 379950.0 138300.0 381150.0 ;
      RECT  132900.0 374250.0 134100.0 375450.0 ;
      RECT  132900.0 374250.0 134100.0 375450.0 ;
      RECT  135450.0 374400.0 136350.0 375300.0 ;
      RECT  130500.0 382050.0 140100.0 382950.0 ;
      RECT  130500.0 367950.0 140100.0 368850.0 ;
      RECT  102750.0 374250.0 103950.0 375450.0 ;
      RECT  104700.0 372000.0 105900.0 373200.0 ;
      RECT  121500.0 372900.0 120300.0 374100.0 ;
      RECT  113100.0 396600.0 114300.0 394650.0 ;
      RECT  113100.0 384450.0 114300.0 382500.0 ;
      RECT  108300.0 395250.0 109500.0 397050.0 ;
      RECT  108300.0 385650.0 109500.0 382050.0 ;
      RECT  111000.0 394050.0 111900.0 385650.0 ;
      RECT  108300.0 385650.0 109500.0 384450.0 ;
      RECT  110700.0 385650.0 111900.0 384450.0 ;
      RECT  110700.0 385650.0 111900.0 384450.0 ;
      RECT  108300.0 385650.0 109500.0 384450.0 ;
      RECT  108300.0 395250.0 109500.0 394050.0 ;
      RECT  110700.0 395250.0 111900.0 394050.0 ;
      RECT  110700.0 395250.0 111900.0 394050.0 ;
      RECT  108300.0 395250.0 109500.0 394050.0 ;
      RECT  113100.0 395250.0 114300.0 394050.0 ;
      RECT  113100.0 385050.0 114300.0 383850.0 ;
      RECT  108900.0 390750.0 110100.0 389550.0 ;
      RECT  108900.0 390750.0 110100.0 389550.0 ;
      RECT  111450.0 390600.0 112350.0 389700.0 ;
      RECT  106500.0 382950.0 116100.0 382050.0 ;
      RECT  106500.0 397050.0 116100.0 396150.0 ;
      RECT  125100.0 396600.0 126300.0 394650.0 ;
      RECT  125100.0 384450.0 126300.0 382500.0 ;
      RECT  117900.0 394650.0 119100.0 397050.0 ;
      RECT  117900.0 385650.0 119100.0 382050.0 ;
      RECT  122700.0 385650.0 123900.0 382050.0 ;
      RECT  117900.0 385650.0 119100.0 384450.0 ;
      RECT  120300.0 385650.0 121500.0 384450.0 ;
      RECT  120300.0 385650.0 121500.0 384450.0 ;
      RECT  117900.0 385650.0 119100.0 384450.0 ;
      RECT  120300.0 385650.0 121500.0 384450.0 ;
      RECT  122700.0 385650.0 123900.0 384450.0 ;
      RECT  122700.0 385650.0 123900.0 384450.0 ;
      RECT  120300.0 385650.0 121500.0 384450.0 ;
      RECT  117900.0 394650.0 119100.0 393450.0 ;
      RECT  120300.0 394650.0 121500.0 393450.0 ;
      RECT  120300.0 394650.0 121500.0 393450.0 ;
      RECT  117900.0 394650.0 119100.0 393450.0 ;
      RECT  120300.0 394650.0 121500.0 393450.0 ;
      RECT  122700.0 394650.0 123900.0 393450.0 ;
      RECT  122700.0 394650.0 123900.0 393450.0 ;
      RECT  120300.0 394650.0 121500.0 393450.0 ;
      RECT  125100.0 395250.0 126300.0 394050.0 ;
      RECT  125100.0 385050.0 126300.0 383850.0 ;
      RECT  122700.0 392100.0 121500.0 390900.0 ;
      RECT  119700.0 389400.0 118500.0 388200.0 ;
      RECT  120300.0 385650.0 121500.0 384450.0 ;
      RECT  122700.0 394650.0 123900.0 393450.0 ;
      RECT  123900.0 389400.0 122700.0 388200.0 ;
      RECT  118500.0 389400.0 119700.0 388200.0 ;
      RECT  121500.0 392100.0 122700.0 390900.0 ;
      RECT  122700.0 389400.0 123900.0 388200.0 ;
      RECT  116100.0 382950.0 130500.0 382050.0 ;
      RECT  116100.0 397050.0 130500.0 396150.0 ;
      RECT  137100.0 396600.0 138300.0 394650.0 ;
      RECT  137100.0 384450.0 138300.0 382500.0 ;
      RECT  132300.0 395250.0 133500.0 397050.0 ;
      RECT  132300.0 385650.0 133500.0 382050.0 ;
      RECT  135000.0 394050.0 135900.0 385650.0 ;
      RECT  132300.0 385650.0 133500.0 384450.0 ;
      RECT  134700.0 385650.0 135900.0 384450.0 ;
      RECT  134700.0 385650.0 135900.0 384450.0 ;
      RECT  132300.0 385650.0 133500.0 384450.0 ;
      RECT  132300.0 395250.0 133500.0 394050.0 ;
      RECT  134700.0 395250.0 135900.0 394050.0 ;
      RECT  134700.0 395250.0 135900.0 394050.0 ;
      RECT  132300.0 395250.0 133500.0 394050.0 ;
      RECT  137100.0 395250.0 138300.0 394050.0 ;
      RECT  137100.0 385050.0 138300.0 383850.0 ;
      RECT  132900.0 390750.0 134100.0 389550.0 ;
      RECT  132900.0 390750.0 134100.0 389550.0 ;
      RECT  135450.0 390600.0 136350.0 389700.0 ;
      RECT  130500.0 382950.0 140100.0 382050.0 ;
      RECT  130500.0 397050.0 140100.0 396150.0 ;
      RECT  102750.0 389550.0 103950.0 390750.0 ;
      RECT  104700.0 391800.0 105900.0 393000.0 ;
      RECT  121500.0 390900.0 120300.0 392100.0 ;
      RECT  113100.0 396600.0 114300.0 398550.0 ;
      RECT  113100.0 408750.0 114300.0 410700.0 ;
      RECT  108300.0 397950.0 109500.0 396150.0 ;
      RECT  108300.0 407550.0 109500.0 411150.0 ;
      RECT  111000.0 399150.0 111900.0 407550.0 ;
      RECT  108300.0 407550.0 109500.0 408750.0 ;
      RECT  110700.0 407550.0 111900.0 408750.0 ;
      RECT  110700.0 407550.0 111900.0 408750.0 ;
      RECT  108300.0 407550.0 109500.0 408750.0 ;
      RECT  108300.0 397950.0 109500.0 399150.0 ;
      RECT  110700.0 397950.0 111900.0 399150.0 ;
      RECT  110700.0 397950.0 111900.0 399150.0 ;
      RECT  108300.0 397950.0 109500.0 399150.0 ;
      RECT  113100.0 397950.0 114300.0 399150.0 ;
      RECT  113100.0 408150.0 114300.0 409350.0 ;
      RECT  108900.0 402450.0 110100.0 403650.0 ;
      RECT  108900.0 402450.0 110100.0 403650.0 ;
      RECT  111450.0 402600.0 112350.0 403500.0 ;
      RECT  106500.0 410250.0 116100.0 411150.0 ;
      RECT  106500.0 396150.0 116100.0 397050.0 ;
      RECT  125100.0 396600.0 126300.0 398550.0 ;
      RECT  125100.0 408750.0 126300.0 410700.0 ;
      RECT  117900.0 398550.0 119100.0 396150.0 ;
      RECT  117900.0 407550.0 119100.0 411150.0 ;
      RECT  122700.0 407550.0 123900.0 411150.0 ;
      RECT  117900.0 407550.0 119100.0 408750.0 ;
      RECT  120300.0 407550.0 121500.0 408750.0 ;
      RECT  120300.0 407550.0 121500.0 408750.0 ;
      RECT  117900.0 407550.0 119100.0 408750.0 ;
      RECT  120300.0 407550.0 121500.0 408750.0 ;
      RECT  122700.0 407550.0 123900.0 408750.0 ;
      RECT  122700.0 407550.0 123900.0 408750.0 ;
      RECT  120300.0 407550.0 121500.0 408750.0 ;
      RECT  117900.0 398550.0 119100.0 399750.0 ;
      RECT  120300.0 398550.0 121500.0 399750.0 ;
      RECT  120300.0 398550.0 121500.0 399750.0 ;
      RECT  117900.0 398550.0 119100.0 399750.0 ;
      RECT  120300.0 398550.0 121500.0 399750.0 ;
      RECT  122700.0 398550.0 123900.0 399750.0 ;
      RECT  122700.0 398550.0 123900.0 399750.0 ;
      RECT  120300.0 398550.0 121500.0 399750.0 ;
      RECT  125100.0 397950.0 126300.0 399150.0 ;
      RECT  125100.0 408150.0 126300.0 409350.0 ;
      RECT  122700.0 401100.0 121500.0 402300.0 ;
      RECT  119700.0 403800.0 118500.0 405000.0 ;
      RECT  120300.0 407550.0 121500.0 408750.0 ;
      RECT  122700.0 398550.0 123900.0 399750.0 ;
      RECT  123900.0 403800.0 122700.0 405000.0 ;
      RECT  118500.0 403800.0 119700.0 405000.0 ;
      RECT  121500.0 401100.0 122700.0 402300.0 ;
      RECT  122700.0 403800.0 123900.0 405000.0 ;
      RECT  116100.0 410250.0 130500.0 411150.0 ;
      RECT  116100.0 396150.0 130500.0 397050.0 ;
      RECT  137100.0 396600.0 138300.0 398550.0 ;
      RECT  137100.0 408750.0 138300.0 410700.0 ;
      RECT  132300.0 397950.0 133500.0 396150.0 ;
      RECT  132300.0 407550.0 133500.0 411150.0 ;
      RECT  135000.0 399150.0 135900.0 407550.0 ;
      RECT  132300.0 407550.0 133500.0 408750.0 ;
      RECT  134700.0 407550.0 135900.0 408750.0 ;
      RECT  134700.0 407550.0 135900.0 408750.0 ;
      RECT  132300.0 407550.0 133500.0 408750.0 ;
      RECT  132300.0 397950.0 133500.0 399150.0 ;
      RECT  134700.0 397950.0 135900.0 399150.0 ;
      RECT  134700.0 397950.0 135900.0 399150.0 ;
      RECT  132300.0 397950.0 133500.0 399150.0 ;
      RECT  137100.0 397950.0 138300.0 399150.0 ;
      RECT  137100.0 408150.0 138300.0 409350.0 ;
      RECT  132900.0 402450.0 134100.0 403650.0 ;
      RECT  132900.0 402450.0 134100.0 403650.0 ;
      RECT  135450.0 402600.0 136350.0 403500.0 ;
      RECT  130500.0 410250.0 140100.0 411150.0 ;
      RECT  130500.0 396150.0 140100.0 397050.0 ;
      RECT  102750.0 402450.0 103950.0 403650.0 ;
      RECT  104700.0 400200.0 105900.0 401400.0 ;
      RECT  121500.0 401100.0 120300.0 402300.0 ;
      RECT  113100.0 424800.0 114300.0 422850.0 ;
      RECT  113100.0 412650.0 114300.0 410700.0 ;
      RECT  108300.0 423450.0 109500.0 425250.0 ;
      RECT  108300.0 413850.0 109500.0 410250.0 ;
      RECT  111000.0 422250.0 111900.0 413850.0 ;
      RECT  108300.0 413850.0 109500.0 412650.0 ;
      RECT  110700.0 413850.0 111900.0 412650.0 ;
      RECT  110700.0 413850.0 111900.0 412650.0 ;
      RECT  108300.0 413850.0 109500.0 412650.0 ;
      RECT  108300.0 423450.0 109500.0 422250.0 ;
      RECT  110700.0 423450.0 111900.0 422250.0 ;
      RECT  110700.0 423450.0 111900.0 422250.0 ;
      RECT  108300.0 423450.0 109500.0 422250.0 ;
      RECT  113100.0 423450.0 114300.0 422250.0 ;
      RECT  113100.0 413250.0 114300.0 412050.0 ;
      RECT  108900.0 418950.0 110100.0 417750.0 ;
      RECT  108900.0 418950.0 110100.0 417750.0 ;
      RECT  111450.0 418800.0 112350.0 417900.0 ;
      RECT  106500.0 411150.0 116100.0 410250.0 ;
      RECT  106500.0 425250.0 116100.0 424350.0 ;
      RECT  125100.0 424800.0 126300.0 422850.0 ;
      RECT  125100.0 412650.0 126300.0 410700.0 ;
      RECT  117900.0 422850.0 119100.0 425250.0 ;
      RECT  117900.0 413850.0 119100.0 410250.0 ;
      RECT  122700.0 413850.0 123900.0 410250.0 ;
      RECT  117900.0 413850.0 119100.0 412650.0 ;
      RECT  120300.0 413850.0 121500.0 412650.0 ;
      RECT  120300.0 413850.0 121500.0 412650.0 ;
      RECT  117900.0 413850.0 119100.0 412650.0 ;
      RECT  120300.0 413850.0 121500.0 412650.0 ;
      RECT  122700.0 413850.0 123900.0 412650.0 ;
      RECT  122700.0 413850.0 123900.0 412650.0 ;
      RECT  120300.0 413850.0 121500.0 412650.0 ;
      RECT  117900.0 422850.0 119100.0 421650.0 ;
      RECT  120300.0 422850.0 121500.0 421650.0 ;
      RECT  120300.0 422850.0 121500.0 421650.0 ;
      RECT  117900.0 422850.0 119100.0 421650.0 ;
      RECT  120300.0 422850.0 121500.0 421650.0 ;
      RECT  122700.0 422850.0 123900.0 421650.0 ;
      RECT  122700.0 422850.0 123900.0 421650.0 ;
      RECT  120300.0 422850.0 121500.0 421650.0 ;
      RECT  125100.0 423450.0 126300.0 422250.0 ;
      RECT  125100.0 413250.0 126300.0 412050.0 ;
      RECT  122700.0 420300.0 121500.0 419100.0 ;
      RECT  119700.0 417600.0 118500.0 416400.0 ;
      RECT  120300.0 413850.0 121500.0 412650.0 ;
      RECT  122700.0 422850.0 123900.0 421650.0 ;
      RECT  123900.0 417600.0 122700.0 416400.0 ;
      RECT  118500.0 417600.0 119700.0 416400.0 ;
      RECT  121500.0 420300.0 122700.0 419100.0 ;
      RECT  122700.0 417600.0 123900.0 416400.0 ;
      RECT  116100.0 411150.0 130500.0 410250.0 ;
      RECT  116100.0 425250.0 130500.0 424350.0 ;
      RECT  137100.0 424800.0 138300.0 422850.0 ;
      RECT  137100.0 412650.0 138300.0 410700.0 ;
      RECT  132300.0 423450.0 133500.0 425250.0 ;
      RECT  132300.0 413850.0 133500.0 410250.0 ;
      RECT  135000.0 422250.0 135900.0 413850.0 ;
      RECT  132300.0 413850.0 133500.0 412650.0 ;
      RECT  134700.0 413850.0 135900.0 412650.0 ;
      RECT  134700.0 413850.0 135900.0 412650.0 ;
      RECT  132300.0 413850.0 133500.0 412650.0 ;
      RECT  132300.0 423450.0 133500.0 422250.0 ;
      RECT  134700.0 423450.0 135900.0 422250.0 ;
      RECT  134700.0 423450.0 135900.0 422250.0 ;
      RECT  132300.0 423450.0 133500.0 422250.0 ;
      RECT  137100.0 423450.0 138300.0 422250.0 ;
      RECT  137100.0 413250.0 138300.0 412050.0 ;
      RECT  132900.0 418950.0 134100.0 417750.0 ;
      RECT  132900.0 418950.0 134100.0 417750.0 ;
      RECT  135450.0 418800.0 136350.0 417900.0 ;
      RECT  130500.0 411150.0 140100.0 410250.0 ;
      RECT  130500.0 425250.0 140100.0 424350.0 ;
      RECT  102750.0 417750.0 103950.0 418950.0 ;
      RECT  104700.0 420000.0 105900.0 421200.0 ;
      RECT  121500.0 419100.0 120300.0 420300.0 ;
      RECT  100200.0 202950.0 105300.0 203850.0 ;
      RECT  100200.0 222750.0 105300.0 223650.0 ;
      RECT  100200.0 231150.0 105300.0 232050.0 ;
      RECT  100200.0 250950.0 105300.0 251850.0 ;
      RECT  100200.0 259350.0 105300.0 260250.0 ;
      RECT  100200.0 279150.0 105300.0 280050.0 ;
      RECT  100200.0 287550.0 105300.0 288450.0 ;
      RECT  100200.0 307350.0 105300.0 308250.0 ;
      RECT  100200.0 315750.0 105300.0 316650.0 ;
      RECT  100200.0 335550.0 105300.0 336450.0 ;
      RECT  100200.0 343950.0 105300.0 344850.0 ;
      RECT  100200.0 363750.0 105300.0 364650.0 ;
      RECT  100200.0 372150.0 105300.0 373050.0 ;
      RECT  100200.0 391950.0 105300.0 392850.0 ;
      RECT  100200.0 400350.0 105300.0 401250.0 ;
      RECT  100200.0 420150.0 105300.0 421050.0 ;
      RECT  135450.0 205200.0 136350.0 206100.0 ;
      RECT  135450.0 220500.0 136350.0 221400.0 ;
      RECT  135450.0 233400.0 136350.0 234300.0 ;
      RECT  135450.0 248700.0 136350.0 249600.0 ;
      RECT  135450.0 261600.0 136350.0 262500.0 ;
      RECT  135450.0 276900.0 136350.0 277800.0 ;
      RECT  135450.0 289800.0 136350.0 290700.0 ;
      RECT  135450.0 305100.0 136350.0 306000.0 ;
      RECT  135450.0 318000.0 136350.0 318900.0 ;
      RECT  135450.0 333300.0 136350.0 334200.0 ;
      RECT  135450.0 346200.0 136350.0 347100.0 ;
      RECT  135450.0 361500.0 136350.0 362400.0 ;
      RECT  135450.0 374400.0 136350.0 375300.0 ;
      RECT  135450.0 389700.0 136350.0 390600.0 ;
      RECT  135450.0 402600.0 136350.0 403500.0 ;
      RECT  135450.0 417900.0 136350.0 418800.0 ;
      RECT  100200.0 212850.0 106500.0 213750.0 ;
      RECT  100200.0 241050.0 106500.0 241950.0 ;
      RECT  100200.0 269250.0 106500.0 270150.0 ;
      RECT  100200.0 297450.0 106500.0 298350.0 ;
      RECT  100200.0 325650.0 106500.0 326550.0 ;
      RECT  100200.0 353850.0 106500.0 354750.0 ;
      RECT  100200.0 382050.0 106500.0 382950.0 ;
      RECT  100200.0 410250.0 106500.0 411150.0 ;
      RECT  100200.0 198750.0 106500.0 199650.0 ;
      RECT  100200.0 226950.0 106500.0 227850.0 ;
      RECT  100200.0 255150.0 106500.0 256050.0 ;
      RECT  100200.0 283350.0 106500.0 284250.0 ;
      RECT  100200.0 311550.0 106500.0 312450.0 ;
      RECT  100200.0 339750.0 106500.0 340650.0 ;
      RECT  100200.0 367950.0 106500.0 368850.0 ;
      RECT  100200.0 396150.0 106500.0 397050.0 ;
      RECT  100200.0 424350.0 106500.0 425250.0 ;
      RECT  59400.0 81000.0 119400.0 70800.0 ;
      RECT  59400.0 60600.0 119400.0 70800.0 ;
      RECT  59400.0 60600.0 119400.0 50400.0 ;
      RECT  59400.0 40200.0 119400.0 50400.0 ;
      RECT  61800.0 81000.0 62700.0 40200.0 ;
      RECT  115800.0 81000.0 116700.0 40200.0 ;
      RECT  148350.0 199800.0 149550.0 198600.0 ;
      RECT  148350.0 228000.0 149550.0 226800.0 ;
      RECT  148350.0 256200.0 149550.0 255000.0 ;
      RECT  148350.0 284400.0 149550.0 283200.0 ;
      RECT  148350.0 312600.0 149550.0 311400.0 ;
      RECT  148350.0 340800.0 149550.0 339600.0 ;
      RECT  148350.0 369000.0 149550.0 367800.0 ;
      RECT  148350.0 397200.0 149550.0 396000.0 ;
      RECT  148350.0 425400.0 149550.0 424200.0 ;
      RECT  130800.0 88650.0 129600.0 89850.0 ;
      RECT  135900.0 88500.0 134700.0 89700.0 ;
      RECT  127800.0 102750.0 126600.0 103950.0 ;
      RECT  138600.0 102600.0 137400.0 103800.0 ;
      RECT  130800.0 145050.0 129600.0 146250.0 ;
      RECT  141300.0 144900.0 140100.0 146100.0 ;
      RECT  127800.0 159150.0 126600.0 160350.0 ;
      RECT  144000.0 159000.0 142800.0 160200.0 ;
      RECT  132900.0 85800.0 131700.0 87000.0 ;
      RECT  132900.0 114000.0 131700.0 115200.0 ;
      RECT  132900.0 142200.0 131700.0 143400.0 ;
      RECT  132900.0 170400.0 131700.0 171600.0 ;
      RECT  120000.0 75300.0 118800.0 76500.0 ;
      RECT  135900.0 75300.0 134700.0 76500.0 ;
      RECT  120000.0 65100.0 118800.0 66300.0 ;
      RECT  138600.0 65100.0 137400.0 66300.0 ;
      RECT  120000.0 54900.0 118800.0 56100.0 ;
      RECT  141300.0 54900.0 140100.0 56100.0 ;
      RECT  120000.0 44700.0 118800.0 45900.0 ;
      RECT  144000.0 44700.0 142800.0 45900.0 ;
      RECT  120600.0 70200.0 119400.0 71400.0 ;
      RECT  149550.0 70350.0 148350.0 71550.0 ;
      RECT  120600.0 49800.0 119400.0 51000.0 ;
      RECT  149550.0 49950.0 148350.0 51150.0 ;
      RECT  164700.0 32250.0 163500.0 33450.0 ;
      RECT  159300.0 27750.0 158100.0 28950.0 ;
      RECT  162000.0 25350.0 160800.0 26550.0 ;
      RECT  164700.0 429450.0 163500.0 430650.0 ;
      RECT  167400.0 96750.0 166200.0 97950.0 ;
      RECT  170100.0 194850.0 168900.0 196050.0 ;
      RECT  156600.0 82500.0 155400.0 83700.0 ;
      RECT  103950.0 426300.0 102750.0 427500.0 ;
      RECT  156600.0 426300.0 155400.0 427500.0 ;
      RECT  152850.0 23400.0 151650.0 24600.0 ;
      RECT  152850.0 192900.0 151650.0 194100.0 ;
      RECT  152850.0 94800.0 151650.0 96000.0 ;
      RECT  198900.0 0.0 203400.0 444600.0 ;
      RECT  53100.0 0.0 57600.0 444600.0 ;
      RECT  44250.0 207150.0 43350.0 208050.0 ;
      RECT  43800.0 207150.0 43650.0 208050.0 ;
      RECT  44250.0 207600.0 43350.0 217200.0 ;
      RECT  44400.0 223950.0 43500.0 224850.0 ;
      RECT  43950.0 223950.0 43800.0 224850.0 ;
      RECT  44400.0 224400.0 43500.0 231600.0 ;
      RECT  44400.0 243600.0 43500.0 250800.0 ;
      RECT  35550.0 258600.0 30600.0 259500.0 ;
      RECT  44100.0 207150.0 43200.0 208050.0 ;
      RECT  44250.0 223950.0 43350.0 224850.0 ;
      RECT  28800.0 362100.0 27900.0 375450.0 ;
      RECT  44400.0 272850.0 43500.0 284850.0 ;
      RECT  33300.0 204600.0 30600.0 205500.0 ;
      RECT  29400.0 284850.0 28500.0 311700.0 ;
      RECT  26700.0 290250.0 25800.0 314700.0 ;
      RECT  41250.0 303750.0 40350.0 312300.0 ;
      RECT  43200.0 301050.0 42300.0 314700.0 ;
      RECT  45150.0 292950.0 44250.0 317100.0 ;
      RECT  41250.0 326850.0 40350.0 327750.0 ;
      RECT  41250.0 318300.0 40350.0 327300.0 ;
      RECT  43650.0 326850.0 40800.0 327750.0 ;
      RECT  44250.0 329250.0 43350.0 330150.0 ;
      RECT  43800.0 329250.0 43650.0 330150.0 ;
      RECT  44250.0 329700.0 43350.0 387300.0 ;
      RECT  13050.0 303750.0 12150.0 321900.0 ;
      RECT  15000.0 292950.0 14100.0 324300.0 ;
      RECT  16950.0 295650.0 16050.0 326700.0 ;
      RECT  13050.0 336450.0 12150.0 337350.0 ;
      RECT  13050.0 327900.0 12150.0 336900.0 ;
      RECT  15450.0 336450.0 12600.0 337350.0 ;
      RECT  15900.0 339300.0 15000.0 346500.0 ;
      RECT  15900.0 348900.0 15000.0 356100.0 ;
      RECT  28800.0 361650.0 27900.0 362550.0 ;
      RECT  28350.0 361650.0 27900.0 362550.0 ;
      RECT  28800.0 359700.0 27900.0 362100.0 ;
      RECT  28800.0 349500.0 27900.0 356700.0 ;
      RECT  29400.0 316800.0 28500.0 323100.0 ;
      RECT  30150.0 333000.0 29250.0 340200.0 ;
      RECT  15900.0 358500.0 15000.0 362700.0 ;
      RECT  28800.0 342900.0 27900.0 347100.0 ;
      RECT  50550.0 202200.0 49650.0 362100.0 ;
      RECT  50550.0 287550.0 49650.0 308700.0 ;
      RECT  36450.0 202200.0 35550.0 362100.0 ;
      RECT  36450.0 298350.0 35550.0 308700.0 ;
      RECT  22350.0 308700.0 21450.0 362100.0 ;
      RECT  22350.0 287550.0 21450.0 308700.0 ;
      RECT  8250.0 308700.0 7350.0 362100.0 ;
      RECT  8250.0 298350.0 7350.0 308700.0 ;
      RECT  8250.0 361650.0 7350.0 362550.0 ;
      RECT  8250.0 360000.0 7350.0 362100.0 ;
      RECT  7800.0 361650.0 3300.0 362550.0 ;
      RECT  0.0 202200.0 10200.0 262200.0 ;
      RECT  20400.0 202200.0 10200.0 262200.0 ;
      RECT  20400.0 202200.0 30600.0 262200.0 ;
      RECT  0.0 204600.0 30600.0 205500.0 ;
      RECT  7.1054273576e-12 258600.0 30600.0 259500.0 ;
      RECT  50100.0 211200.0 48150.0 212400.0 ;
      RECT  37950.0 211200.0 36000.0 212400.0 ;
      RECT  47550.0 206700.0 39150.0 207600.0 ;
      RECT  38550.0 204150.0 36600.0 205050.0 ;
      RECT  38550.0 208950.0 36600.0 209850.0 ;
      RECT  39150.0 204000.0 37950.0 205200.0 ;
      RECT  39150.0 208800.0 37950.0 210000.0 ;
      RECT  39150.0 206400.0 37950.0 207600.0 ;
      RECT  39150.0 206400.0 37950.0 207600.0 ;
      RECT  37050.0 204000.0 36150.0 210000.0 ;
      RECT  50100.0 204150.0 48150.0 205050.0 ;
      RECT  50100.0 208950.0 48150.0 209850.0 ;
      RECT  48750.0 204000.0 47550.0 205200.0 ;
      RECT  48750.0 208800.0 47550.0 210000.0 ;
      RECT  48750.0 206400.0 47550.0 207600.0 ;
      RECT  48750.0 206400.0 47550.0 207600.0 ;
      RECT  50550.0 204000.0 49650.0 210000.0 ;
      RECT  48750.0 211200.0 47550.0 212400.0 ;
      RECT  38550.0 211200.0 37350.0 212400.0 ;
      RECT  44250.0 204600.0 43050.0 205800.0 ;
      RECT  44250.0 204600.0 43050.0 205800.0 ;
      RECT  44100.0 207150.0 43200.0 208050.0 ;
      RECT  36450.0 202200.0 35550.0 214200.0 ;
      RECT  50550.0 202200.0 49650.0 214200.0 ;
      RECT  50100.0 225600.0 48150.0 226800.0 ;
      RECT  37950.0 225600.0 36000.0 226800.0 ;
      RECT  37350.0 216000.0 35550.0 222000.0 ;
      RECT  45450.0 223500.0 41250.0 224400.0 ;
      RECT  38850.0 216150.0 36900.0 217050.0 ;
      RECT  38850.0 220950.0 36900.0 221850.0 ;
      RECT  40800.0 218550.0 38850.0 219450.0 ;
      RECT  40800.0 223350.0 38850.0 224250.0 ;
      RECT  39450.0 216000.0 38250.0 217200.0 ;
      RECT  39450.0 220800.0 38250.0 222000.0 ;
      RECT  39450.0 218400.0 38250.0 219600.0 ;
      RECT  39450.0 223200.0 38250.0 224400.0 ;
      RECT  41250.0 218400.0 40350.0 224400.0 ;
      RECT  37350.0 216000.0 36450.0 222000.0 ;
      RECT  49800.0 216150.0 47850.0 217050.0 ;
      RECT  49800.0 220950.0 47850.0 221850.0 ;
      RECT  47850.0 218550.0 45900.0 219450.0 ;
      RECT  47850.0 223350.0 45900.0 224250.0 ;
      RECT  48450.0 216000.0 47250.0 217200.0 ;
      RECT  48450.0 220800.0 47250.0 222000.0 ;
      RECT  48450.0 218400.0 47250.0 219600.0 ;
      RECT  48450.0 223200.0 47250.0 224400.0 ;
      RECT  46350.0 218400.0 45450.0 224400.0 ;
      RECT  50250.0 216000.0 49350.0 222000.0 ;
      RECT  48750.0 225600.0 47550.0 226800.0 ;
      RECT  38550.0 225600.0 37350.0 226800.0 ;
      RECT  44400.0 216600.0 43200.0 217800.0 ;
      RECT  44400.0 216600.0 43200.0 217800.0 ;
      RECT  44250.0 223950.0 43350.0 224850.0 ;
      RECT  36450.0 214200.0 35550.0 228600.0 ;
      RECT  50550.0 214200.0 49650.0 228600.0 ;
      RECT  50100.0 244800.0 48150.0 246000.0 ;
      RECT  37950.0 244800.0 36000.0 246000.0 ;
      RECT  37800.0 230400.0 35550.0 241200.0 ;
      RECT  45300.0 242700.0 41700.0 243600.0 ;
      RECT  39300.0 230550.0 37350.0 231450.0 ;
      RECT  39300.0 235350.0 37350.0 236250.0 ;
      RECT  39300.0 240150.0 37350.0 241050.0 ;
      RECT  41250.0 232950.0 39300.0 233850.0 ;
      RECT  41250.0 237750.0 39300.0 238650.0 ;
      RECT  41250.0 242550.0 39300.0 243450.0 ;
      RECT  39900.0 230400.0 38700.0 231600.0 ;
      RECT  39900.0 235200.0 38700.0 236400.0 ;
      RECT  39900.0 240000.0 38700.0 241200.0 ;
      RECT  39900.0 232800.0 38700.0 234000.0 ;
      RECT  39900.0 237600.0 38700.0 238800.0 ;
      RECT  39900.0 242400.0 38700.0 243600.0 ;
      RECT  41700.0 232800.0 40800.0 243600.0 ;
      RECT  37800.0 230400.0 36900.0 241200.0 ;
      RECT  49650.0 230550.0 47700.0 231450.0 ;
      RECT  49650.0 235350.0 47700.0 236250.0 ;
      RECT  49650.0 240150.0 47700.0 241050.0 ;
      RECT  47700.0 232950.0 45750.0 233850.0 ;
      RECT  47700.0 237750.0 45750.0 238650.0 ;
      RECT  47700.0 242550.0 45750.0 243450.0 ;
      RECT  48300.0 230400.0 47100.0 231600.0 ;
      RECT  48300.0 235200.0 47100.0 236400.0 ;
      RECT  48300.0 240000.0 47100.0 241200.0 ;
      RECT  48300.0 232800.0 47100.0 234000.0 ;
      RECT  48300.0 237600.0 47100.0 238800.0 ;
      RECT  48300.0 242400.0 47100.0 243600.0 ;
      RECT  46200.0 232800.0 45300.0 243600.0 ;
      RECT  50100.0 230400.0 49200.0 241200.0 ;
      RECT  48750.0 244800.0 47550.0 246000.0 ;
      RECT  38550.0 244800.0 37350.0 246000.0 ;
      RECT  44550.0 231000.0 43350.0 232200.0 ;
      RECT  44550.0 231000.0 43350.0 232200.0 ;
      RECT  44400.0 243150.0 43500.0 244050.0 ;
      RECT  36450.0 228600.0 35550.0 247800.0 ;
      RECT  50550.0 228600.0 49650.0 247800.0 ;
      RECT  50100.0 276000.0 48150.0 277200.0 ;
      RECT  37950.0 276000.0 36000.0 277200.0 ;
      RECT  37800.0 249600.0 35550.0 274800.0 ;
      RECT  45300.0 271500.0 41700.0 272400.0 ;
      RECT  39300.0 249750.0 37350.0 250650.0 ;
      RECT  39300.0 254550.0 37350.0 255450.0 ;
      RECT  39300.0 259350.0 37350.0 260250.0 ;
      RECT  39300.0 264150.0 37350.0 265050.0 ;
      RECT  39300.0 268950.0 37350.0 269850.0 ;
      RECT  39300.0 273750.0 37350.0 274650.0 ;
      RECT  41250.0 252150.0 39300.0 253050.0 ;
      RECT  41250.0 256950.0 39300.0 257850.0 ;
      RECT  41250.0 261750.0 39300.0 262650.0 ;
      RECT  41250.0 266550.0 39300.0 267450.0 ;
      RECT  41250.0 271350.0 39300.0 272250.0 ;
      RECT  39900.0 249600.0 38700.0 250800.0 ;
      RECT  39900.0 254400.0 38700.0 255600.0 ;
      RECT  39900.0 259200.0 38700.0 260400.0 ;
      RECT  39900.0 264000.0 38700.0 265200.0 ;
      RECT  39900.0 268800.0 38700.0 270000.0 ;
      RECT  39900.0 273600.0 38700.0 274800.0 ;
      RECT  39900.0 252000.0 38700.0 253200.0 ;
      RECT  39900.0 256800.0 38700.0 258000.0 ;
      RECT  39900.0 261600.0 38700.0 262800.0 ;
      RECT  39900.0 266400.0 38700.0 267600.0 ;
      RECT  39900.0 271200.0 38700.0 272400.0 ;
      RECT  41700.0 252000.0 40800.0 272400.0 ;
      RECT  37800.0 249600.0 36900.0 274800.0 ;
      RECT  49650.0 249750.0 47700.0 250650.0 ;
      RECT  49650.0 254550.0 47700.0 255450.0 ;
      RECT  49650.0 259350.0 47700.0 260250.0 ;
      RECT  49650.0 264150.0 47700.0 265050.0 ;
      RECT  49650.0 268950.0 47700.0 269850.0 ;
      RECT  49650.0 273750.0 47700.0 274650.0 ;
      RECT  47700.0 252150.0 45750.0 253050.0 ;
      RECT  47700.0 256950.0 45750.0 257850.0 ;
      RECT  47700.0 261750.0 45750.0 262650.0 ;
      RECT  47700.0 266550.0 45750.0 267450.0 ;
      RECT  47700.0 271350.0 45750.0 272250.0 ;
      RECT  48300.0 249600.0 47100.0 250800.0 ;
      RECT  48300.0 254400.0 47100.0 255600.0 ;
      RECT  48300.0 259200.0 47100.0 260400.0 ;
      RECT  48300.0 264000.0 47100.0 265200.0 ;
      RECT  48300.0 268800.0 47100.0 270000.0 ;
      RECT  48300.0 273600.0 47100.0 274800.0 ;
      RECT  48300.0 252000.0 47100.0 253200.0 ;
      RECT  48300.0 256800.0 47100.0 258000.0 ;
      RECT  48300.0 261600.0 47100.0 262800.0 ;
      RECT  48300.0 266400.0 47100.0 267600.0 ;
      RECT  48300.0 271200.0 47100.0 272400.0 ;
      RECT  46200.0 252000.0 45300.0 272400.0 ;
      RECT  50100.0 249600.0 49200.0 274800.0 ;
      RECT  48750.0 276000.0 47550.0 277200.0 ;
      RECT  38550.0 276000.0 37350.0 277200.0 ;
      RECT  44550.0 250200.0 43350.0 251400.0 ;
      RECT  44550.0 250200.0 43350.0 251400.0 ;
      RECT  44400.0 271950.0 43500.0 272850.0 ;
      RECT  36450.0 247800.0 35550.0 279000.0 ;
      RECT  50550.0 247800.0 49650.0 279000.0 ;
      RECT  50100.0 320100.0 48600.0 321300.0 ;
      RECT  37500.0 320100.0 36000.0 321300.0 ;
      RECT  48000.0 310500.0 50550.0 311700.0 ;
      RECT  38700.0 310500.0 35550.0 311700.0 ;
      RECT  38700.0 315300.0 35550.0 316500.0 ;
      RECT  38700.0 310500.0 37500.0 311700.0 ;
      RECT  38700.0 312900.0 37500.0 314100.0 ;
      RECT  38700.0 312900.0 37500.0 314100.0 ;
      RECT  38700.0 310500.0 37500.0 311700.0 ;
      RECT  38700.0 312900.0 37500.0 314100.0 ;
      RECT  38700.0 315300.0 37500.0 316500.0 ;
      RECT  38700.0 315300.0 37500.0 316500.0 ;
      RECT  38700.0 312900.0 37500.0 314100.0 ;
      RECT  38700.0 315300.0 37500.0 316500.0 ;
      RECT  38700.0 317700.0 37500.0 318900.0 ;
      RECT  38700.0 317700.0 37500.0 318900.0 ;
      RECT  38700.0 315300.0 37500.0 316500.0 ;
      RECT  48000.0 310500.0 46800.0 311700.0 ;
      RECT  48000.0 312900.0 46800.0 314100.0 ;
      RECT  48000.0 312900.0 46800.0 314100.0 ;
      RECT  48000.0 310500.0 46800.0 311700.0 ;
      RECT  48000.0 312900.0 46800.0 314100.0 ;
      RECT  48000.0 315300.0 46800.0 316500.0 ;
      RECT  48000.0 315300.0 46800.0 316500.0 ;
      RECT  48000.0 312900.0 46800.0 314100.0 ;
      RECT  48000.0 315300.0 46800.0 316500.0 ;
      RECT  48000.0 317700.0 46800.0 318900.0 ;
      RECT  48000.0 317700.0 46800.0 318900.0 ;
      RECT  48000.0 315300.0 46800.0 316500.0 ;
      RECT  49200.0 320100.0 48000.0 321300.0 ;
      RECT  38100.0 320100.0 36900.0 321300.0 ;
      RECT  45300.0 317700.0 44100.0 316500.0 ;
      RECT  43350.0 315300.0 42150.0 314100.0 ;
      RECT  41400.0 312900.0 40200.0 311700.0 ;
      RECT  38700.0 312900.0 37500.0 314100.0 ;
      RECT  38700.0 317700.0 37500.0 318900.0 ;
      RECT  48000.0 317700.0 46800.0 318900.0 ;
      RECT  41400.0 317700.0 40200.0 318900.0 ;
      RECT  41400.0 311700.0 40200.0 312900.0 ;
      RECT  43350.0 314100.0 42150.0 315300.0 ;
      RECT  45300.0 316500.0 44100.0 317700.0 ;
      RECT  41400.0 317700.0 40200.0 318900.0 ;
      RECT  36450.0 308700.0 35550.0 324300.0 ;
      RECT  50550.0 308700.0 49650.0 324300.0 ;
      RECT  50100.0 330900.0 48150.0 332100.0 ;
      RECT  37950.0 330900.0 36000.0 332100.0 ;
      RECT  48750.0 326100.0 50550.0 327300.0 ;
      RECT  39150.0 326100.0 35550.0 327300.0 ;
      RECT  47550.0 328800.0 39150.0 329700.0 ;
      RECT  39150.0 326100.0 37950.0 327300.0 ;
      RECT  39150.0 328500.0 37950.0 329700.0 ;
      RECT  39150.0 328500.0 37950.0 329700.0 ;
      RECT  39150.0 326100.0 37950.0 327300.0 ;
      RECT  48750.0 326100.0 47550.0 327300.0 ;
      RECT  48750.0 328500.0 47550.0 329700.0 ;
      RECT  48750.0 328500.0 47550.0 329700.0 ;
      RECT  48750.0 326100.0 47550.0 327300.0 ;
      RECT  48750.0 330900.0 47550.0 332100.0 ;
      RECT  38550.0 330900.0 37350.0 332100.0 ;
      RECT  44250.0 326700.0 43050.0 327900.0 ;
      RECT  44250.0 326700.0 43050.0 327900.0 ;
      RECT  44100.0 329250.0 43200.0 330150.0 ;
      RECT  36450.0 324300.0 35550.0 333900.0 ;
      RECT  50550.0 324300.0 49650.0 333900.0 ;
      RECT  21900.0 317700.0 23850.0 318900.0 ;
      RECT  34050.0 317700.0 36000.0 318900.0 ;
      RECT  23250.0 310500.0 21450.0 311700.0 ;
      RECT  23250.0 315300.0 21450.0 316500.0 ;
      RECT  32250.0 310500.0 36450.0 311700.0 ;
      RECT  32250.0 310500.0 33450.0 311700.0 ;
      RECT  32250.0 312900.0 33450.0 314100.0 ;
      RECT  32250.0 312900.0 33450.0 314100.0 ;
      RECT  32250.0 310500.0 33450.0 311700.0 ;
      RECT  32250.0 312900.0 33450.0 314100.0 ;
      RECT  32250.0 315300.0 33450.0 316500.0 ;
      RECT  32250.0 315300.0 33450.0 316500.0 ;
      RECT  32250.0 312900.0 33450.0 314100.0 ;
      RECT  23250.0 310500.0 24450.0 311700.0 ;
      RECT  23250.0 312900.0 24450.0 314100.0 ;
      RECT  23250.0 312900.0 24450.0 314100.0 ;
      RECT  23250.0 310500.0 24450.0 311700.0 ;
      RECT  23250.0 312900.0 24450.0 314100.0 ;
      RECT  23250.0 315300.0 24450.0 316500.0 ;
      RECT  23250.0 315300.0 24450.0 316500.0 ;
      RECT  23250.0 312900.0 24450.0 314100.0 ;
      RECT  23250.0 317700.0 24450.0 318900.0 ;
      RECT  33450.0 317700.0 34650.0 318900.0 ;
      RECT  25650.0 315300.0 26850.0 314100.0 ;
      RECT  28350.0 312300.0 29550.0 311100.0 ;
      RECT  32250.0 315300.0 33450.0 316500.0 ;
      RECT  23250.0 314100.0 24450.0 312900.0 ;
      RECT  28350.0 317400.0 29550.0 316200.0 ;
      RECT  28350.0 311100.0 29550.0 312300.0 ;
      RECT  25650.0 314100.0 26850.0 315300.0 ;
      RECT  28350.0 316200.0 29550.0 317400.0 ;
      RECT  35550.0 308700.0 36450.0 323100.0 ;
      RECT  21450.0 308700.0 22350.0 323100.0 ;
      RECT  21900.0 334800.0 23850.0 336000.0 ;
      RECT  34050.0 334800.0 36000.0 336000.0 ;
      RECT  23850.0 327600.0 21450.0 328800.0 ;
      RECT  32850.0 327600.0 36450.0 328800.0 ;
      RECT  32850.0 332400.0 36450.0 333600.0 ;
      RECT  32850.0 327600.0 34050.0 328800.0 ;
      RECT  32850.0 330000.0 34050.0 331200.0 ;
      RECT  32850.0 330000.0 34050.0 331200.0 ;
      RECT  32850.0 327600.0 34050.0 328800.0 ;
      RECT  32850.0 330000.0 34050.0 331200.0 ;
      RECT  32850.0 332400.0 34050.0 333600.0 ;
      RECT  32850.0 332400.0 34050.0 333600.0 ;
      RECT  32850.0 330000.0 34050.0 331200.0 ;
      RECT  23850.0 327600.0 25050.0 328800.0 ;
      RECT  23850.0 330000.0 25050.0 331200.0 ;
      RECT  23850.0 330000.0 25050.0 331200.0 ;
      RECT  23850.0 327600.0 25050.0 328800.0 ;
      RECT  23850.0 330000.0 25050.0 331200.0 ;
      RECT  23850.0 332400.0 25050.0 333600.0 ;
      RECT  23850.0 332400.0 25050.0 333600.0 ;
      RECT  23850.0 330000.0 25050.0 331200.0 ;
      RECT  23250.0 334800.0 24450.0 336000.0 ;
      RECT  33450.0 334800.0 34650.0 336000.0 ;
      RECT  26400.0 332400.0 27600.0 331200.0 ;
      RECT  29100.0 329400.0 30300.0 328200.0 ;
      RECT  32850.0 330000.0 34050.0 331200.0 ;
      RECT  23850.0 332400.0 25050.0 333600.0 ;
      RECT  29100.0 333600.0 30300.0 332400.0 ;
      RECT  29100.0 328200.0 30300.0 329400.0 ;
      RECT  26400.0 331200.0 27600.0 332400.0 ;
      RECT  29100.0 332400.0 30300.0 333600.0 ;
      RECT  35550.0 325800.0 36450.0 340200.0 ;
      RECT  21450.0 325800.0 22350.0 340200.0 ;
      RECT  21900.0 345900.0 23850.0 344700.0 ;
      RECT  34050.0 345900.0 36000.0 344700.0 ;
      RECT  23250.0 350700.0 21450.0 349500.0 ;
      RECT  32850.0 350700.0 36450.0 349500.0 ;
      RECT  24450.0 348000.0 32850.0 347100.0 ;
      RECT  32850.0 350700.0 34050.0 349500.0 ;
      RECT  32850.0 348300.0 34050.0 347100.0 ;
      RECT  32850.0 348300.0 34050.0 347100.0 ;
      RECT  32850.0 350700.0 34050.0 349500.0 ;
      RECT  23250.0 350700.0 24450.0 349500.0 ;
      RECT  23250.0 348300.0 24450.0 347100.0 ;
      RECT  23250.0 348300.0 24450.0 347100.0 ;
      RECT  23250.0 350700.0 24450.0 349500.0 ;
      RECT  23250.0 345900.0 24450.0 344700.0 ;
      RECT  33450.0 345900.0 34650.0 344700.0 ;
      RECT  27750.0 350100.0 28950.0 348900.0 ;
      RECT  27750.0 350100.0 28950.0 348900.0 ;
      RECT  27900.0 347550.0 28800.0 346650.0 ;
      RECT  35550.0 352500.0 36450.0 342900.0 ;
      RECT  21450.0 352500.0 22350.0 342900.0 ;
      RECT  21900.0 355500.0 23850.0 354300.0 ;
      RECT  34050.0 355500.0 36000.0 354300.0 ;
      RECT  23250.0 360300.0 21450.0 359100.0 ;
      RECT  32850.0 360300.0 36450.0 359100.0 ;
      RECT  24450.0 357600.0 32850.0 356700.0 ;
      RECT  32850.0 360300.0 34050.0 359100.0 ;
      RECT  32850.0 357900.0 34050.0 356700.0 ;
      RECT  32850.0 357900.0 34050.0 356700.0 ;
      RECT  32850.0 360300.0 34050.0 359100.0 ;
      RECT  23250.0 360300.0 24450.0 359100.0 ;
      RECT  23250.0 357900.0 24450.0 356700.0 ;
      RECT  23250.0 357900.0 24450.0 356700.0 ;
      RECT  23250.0 360300.0 24450.0 359100.0 ;
      RECT  23250.0 355500.0 24450.0 354300.0 ;
      RECT  33450.0 355500.0 34650.0 354300.0 ;
      RECT  27750.0 359700.0 28950.0 358500.0 ;
      RECT  27750.0 359700.0 28950.0 358500.0 ;
      RECT  27900.0 357150.0 28800.0 356250.0 ;
      RECT  35550.0 362100.0 36450.0 352500.0 ;
      RECT  21450.0 362100.0 22350.0 352500.0 ;
      RECT  21900.0 329700.0 20400.0 330900.0 ;
      RECT  9300.0 329700.0 7800.0 330900.0 ;
      RECT  19800.0 320100.0 22350.0 321300.0 ;
      RECT  10500.0 320100.0 7350.0 321300.0 ;
      RECT  10500.0 324900.0 7350.0 326100.0 ;
      RECT  10500.0 320100.0 9300.0 321300.0 ;
      RECT  10500.0 322500.0 9300.0 323700.0 ;
      RECT  10500.0 322500.0 9300.0 323700.0 ;
      RECT  10500.0 320100.0 9300.0 321300.0 ;
      RECT  10500.0 322500.0 9300.0 323700.0 ;
      RECT  10500.0 324900.0 9300.0 326100.0 ;
      RECT  10500.0 324900.0 9300.0 326100.0 ;
      RECT  10500.0 322500.0 9300.0 323700.0 ;
      RECT  10500.0 324900.0 9300.0 326100.0 ;
      RECT  10500.0 327300.0 9300.0 328500.0 ;
      RECT  10500.0 327300.0 9300.0 328500.0 ;
      RECT  10500.0 324900.0 9300.0 326100.0 ;
      RECT  19800.0 320100.0 18600.0 321300.0 ;
      RECT  19800.0 322500.0 18600.0 323700.0 ;
      RECT  19800.0 322500.0 18600.0 323700.0 ;
      RECT  19800.0 320100.0 18600.0 321300.0 ;
      RECT  19800.0 322500.0 18600.0 323700.0 ;
      RECT  19800.0 324900.0 18600.0 326100.0 ;
      RECT  19800.0 324900.0 18600.0 326100.0 ;
      RECT  19800.0 322500.0 18600.0 323700.0 ;
      RECT  19800.0 324900.0 18600.0 326100.0 ;
      RECT  19800.0 327300.0 18600.0 328500.0 ;
      RECT  19800.0 327300.0 18600.0 328500.0 ;
      RECT  19800.0 324900.0 18600.0 326100.0 ;
      RECT  21000.0 329700.0 19800.0 330900.0 ;
      RECT  9900.0 329700.0 8700.0 330900.0 ;
      RECT  17100.0 327300.0 15900.0 326100.0 ;
      RECT  15150.0 324900.0 13950.0 323700.0 ;
      RECT  13200.0 322500.0 12000.0 321300.0 ;
      RECT  10500.0 322500.0 9300.0 323700.0 ;
      RECT  10500.0 327300.0 9300.0 328500.0 ;
      RECT  19800.0 327300.0 18600.0 328500.0 ;
      RECT  13200.0 327300.0 12000.0 328500.0 ;
      RECT  13200.0 321300.0 12000.0 322500.0 ;
      RECT  15150.0 323700.0 13950.0 324900.0 ;
      RECT  17100.0 326100.0 15900.0 327300.0 ;
      RECT  13200.0 327300.0 12000.0 328500.0 ;
      RECT  8250.0 318300.0 7350.0 333900.0 ;
      RECT  22350.0 318300.0 21450.0 333900.0 ;
      RECT  21900.0 340500.0 19950.0 341700.0 ;
      RECT  9750.0 340500.0 7800.0 341700.0 ;
      RECT  20550.0 335700.0 22350.0 336900.0 ;
      RECT  10950.0 335700.0 7350.0 336900.0 ;
      RECT  19350.0 338400.0 10950.0 339300.0 ;
      RECT  10950.0 335700.0 9750.0 336900.0 ;
      RECT  10950.0 338100.0 9750.0 339300.0 ;
      RECT  10950.0 338100.0 9750.0 339300.0 ;
      RECT  10950.0 335700.0 9750.0 336900.0 ;
      RECT  20550.0 335700.0 19350.0 336900.0 ;
      RECT  20550.0 338100.0 19350.0 339300.0 ;
      RECT  20550.0 338100.0 19350.0 339300.0 ;
      RECT  20550.0 335700.0 19350.0 336900.0 ;
      RECT  20550.0 340500.0 19350.0 341700.0 ;
      RECT  10350.0 340500.0 9150.0 341700.0 ;
      RECT  16050.0 336300.0 14850.0 337500.0 ;
      RECT  16050.0 336300.0 14850.0 337500.0 ;
      RECT  15900.0 338850.0 15000.0 339750.0 ;
      RECT  8250.0 333900.0 7350.0 343500.0 ;
      RECT  22350.0 333900.0 21450.0 343500.0 ;
      RECT  21900.0 350100.0 19950.0 351300.0 ;
      RECT  9750.0 350100.0 7800.0 351300.0 ;
      RECT  20550.0 345300.0 22350.0 346500.0 ;
      RECT  10950.0 345300.0 7350.0 346500.0 ;
      RECT  19350.0 348000.0 10950.0 348900.0 ;
      RECT  10950.0 345300.0 9750.0 346500.0 ;
      RECT  10950.0 347700.0 9750.0 348900.0 ;
      RECT  10950.0 347700.0 9750.0 348900.0 ;
      RECT  10950.0 345300.0 9750.0 346500.0 ;
      RECT  20550.0 345300.0 19350.0 346500.0 ;
      RECT  20550.0 347700.0 19350.0 348900.0 ;
      RECT  20550.0 347700.0 19350.0 348900.0 ;
      RECT  20550.0 345300.0 19350.0 346500.0 ;
      RECT  20550.0 350100.0 19350.0 351300.0 ;
      RECT  10350.0 350100.0 9150.0 351300.0 ;
      RECT  16050.0 345900.0 14850.0 347100.0 ;
      RECT  16050.0 345900.0 14850.0 347100.0 ;
      RECT  15900.0 348450.0 15000.0 349350.0 ;
      RECT  8250.0 343500.0 7350.0 353100.0 ;
      RECT  22350.0 343500.0 21450.0 353100.0 ;
      RECT  21900.0 359700.0 19950.0 360900.0 ;
      RECT  9750.0 359700.0 7800.0 360900.0 ;
      RECT  20550.0 354900.0 22350.0 356100.0 ;
      RECT  10950.0 354900.0 7350.0 356100.0 ;
      RECT  19350.0 357600.0 10950.0 358500.0 ;
      RECT  10950.0 354900.0 9750.0 356100.0 ;
      RECT  10950.0 357300.0 9750.0 358500.0 ;
      RECT  10950.0 357300.0 9750.0 358500.0 ;
      RECT  10950.0 354900.0 9750.0 356100.0 ;
      RECT  20550.0 354900.0 19350.0 356100.0 ;
      RECT  20550.0 357300.0 19350.0 358500.0 ;
      RECT  20550.0 357300.0 19350.0 358500.0 ;
      RECT  20550.0 354900.0 19350.0 356100.0 ;
      RECT  20550.0 359700.0 19350.0 360900.0 ;
      RECT  10350.0 359700.0 9150.0 360900.0 ;
      RECT  16050.0 355500.0 14850.0 356700.0 ;
      RECT  16050.0 355500.0 14850.0 356700.0 ;
      RECT  15900.0 358050.0 15000.0 358950.0 ;
      RECT  8250.0 353100.0 7350.0 362700.0 ;
      RECT  22350.0 353100.0 21450.0 362700.0 ;
      RECT  22350.0 398100.0 16500.0 399000.0 ;
      RECT  22350.0 420900.0 16500.0 421800.0 ;
      RECT  21900.0 426450.0 6300.0 427350.0 ;
      RECT  4200.0 409500.0 16500.0 410400.0 ;
      RECT  4200.0 381300.0 16500.0 382200.0 ;
      RECT  28800.0 397500.0 27900.0 410100.0 ;
      RECT  28800.0 392850.0 27900.0 393750.0 ;
      RECT  28800.0 393300.0 27900.0 397500.0 ;
      RECT  28350.0 392850.0 16500.0 393750.0 ;
      RECT  36000.0 398250.0 33600.0 399150.0 ;
      RECT  33450.0 383550.0 32550.0 384450.0 ;
      RECT  28800.0 383550.0 27900.0 384450.0 ;
      RECT  33450.0 384000.0 32550.0 395700.0 ;
      RECT  33000.0 383550.0 28350.0 384450.0 ;
      RECT  28800.0 378900.0 27900.0 384000.0 ;
      RECT  28350.0 383550.0 19650.0 384450.0 ;
      RECT  19650.0 376050.0 12900.0 376950.0 ;
      RECT  28950.0 377700.0 27750.0 378900.0 ;
      RECT  28800.0 410100.0 27900.0 413850.0 ;
      RECT  21900.0 374700.0 23850.0 373500.0 ;
      RECT  34050.0 374700.0 36000.0 373500.0 ;
      RECT  23250.0 379500.0 21450.0 378300.0 ;
      RECT  32850.0 379500.0 36450.0 378300.0 ;
      RECT  24450.0 376800.0 32850.0 375900.0 ;
      RECT  32850.0 379500.0 34050.0 378300.0 ;
      RECT  32850.0 377100.0 34050.0 375900.0 ;
      RECT  32850.0 377100.0 34050.0 375900.0 ;
      RECT  32850.0 379500.0 34050.0 378300.0 ;
      RECT  23250.0 379500.0 24450.0 378300.0 ;
      RECT  23250.0 377100.0 24450.0 375900.0 ;
      RECT  23250.0 377100.0 24450.0 375900.0 ;
      RECT  23250.0 379500.0 24450.0 378300.0 ;
      RECT  23250.0 374700.0 24450.0 373500.0 ;
      RECT  33450.0 374700.0 34650.0 373500.0 ;
      RECT  27750.0 378900.0 28950.0 377700.0 ;
      RECT  27750.0 378900.0 28950.0 377700.0 ;
      RECT  27900.0 376350.0 28800.0 375450.0 ;
      RECT  35550.0 381300.0 36450.0 371700.0 ;
      RECT  21450.0 381300.0 22350.0 371700.0 ;
      RECT  32400.0 395700.0 33600.0 396900.0 ;
      RECT  32400.0 398100.0 33600.0 399300.0 ;
      RECT  32400.0 398100.0 33600.0 399300.0 ;
      RECT  32400.0 395700.0 33600.0 396900.0 ;
      RECT  21450.0 430650.0 22350.0 431550.0 ;
      RECT  49650.0 430650.0 50550.0 431550.0 ;
      RECT  21450.0 429300.0 22350.0 431100.0 ;
      RECT  21900.0 430650.0 50100.0 431550.0 ;
      RECT  49650.0 429300.0 50550.0 431100.0 ;
      RECT  50100.0 416700.0 48150.0 417900.0 ;
      RECT  37950.0 416700.0 36000.0 417900.0 ;
      RECT  48750.0 411900.0 50550.0 413100.0 ;
      RECT  39150.0 411900.0 35550.0 413100.0 ;
      RECT  47550.0 414600.0 39150.0 415500.0 ;
      RECT  39150.0 411900.0 37950.0 413100.0 ;
      RECT  39150.0 414300.0 37950.0 415500.0 ;
      RECT  39150.0 414300.0 37950.0 415500.0 ;
      RECT  39150.0 411900.0 37950.0 413100.0 ;
      RECT  48750.0 411900.0 47550.0 413100.0 ;
      RECT  48750.0 414300.0 47550.0 415500.0 ;
      RECT  48750.0 414300.0 47550.0 415500.0 ;
      RECT  48750.0 411900.0 47550.0 413100.0 ;
      RECT  48750.0 416700.0 47550.0 417900.0 ;
      RECT  38550.0 416700.0 37350.0 417900.0 ;
      RECT  44250.0 412500.0 43050.0 413700.0 ;
      RECT  44250.0 412500.0 43050.0 413700.0 ;
      RECT  44100.0 415050.0 43200.0 415950.0 ;
      RECT  36450.0 410100.0 35550.0 419700.0 ;
      RECT  50550.0 410100.0 49650.0 419700.0 ;
      RECT  50100.0 426300.0 48150.0 427500.0 ;
      RECT  37950.0 426300.0 36000.0 427500.0 ;
      RECT  48750.0 421500.0 50550.0 422700.0 ;
      RECT  39150.0 421500.0 35550.0 422700.0 ;
      RECT  47550.0 424200.0 39150.0 425100.0 ;
      RECT  39150.0 421500.0 37950.0 422700.0 ;
      RECT  39150.0 423900.0 37950.0 425100.0 ;
      RECT  39150.0 423900.0 37950.0 425100.0 ;
      RECT  39150.0 421500.0 37950.0 422700.0 ;
      RECT  48750.0 421500.0 47550.0 422700.0 ;
      RECT  48750.0 423900.0 47550.0 425100.0 ;
      RECT  48750.0 423900.0 47550.0 425100.0 ;
      RECT  48750.0 421500.0 47550.0 422700.0 ;
      RECT  48750.0 426300.0 47550.0 427500.0 ;
      RECT  38550.0 426300.0 37350.0 427500.0 ;
      RECT  44250.0 422100.0 43050.0 423300.0 ;
      RECT  44250.0 422100.0 43050.0 423300.0 ;
      RECT  44100.0 424650.0 43200.0 425550.0 ;
      RECT  36450.0 419700.0 35550.0 429300.0 ;
      RECT  50550.0 419700.0 49650.0 429300.0 ;
      RECT  43050.0 422100.0 44250.0 423300.0 ;
      RECT  21900.0 422700.0 23850.0 421500.0 ;
      RECT  34050.0 422700.0 36000.0 421500.0 ;
      RECT  23250.0 427500.0 21450.0 426300.0 ;
      RECT  32850.0 427500.0 36450.0 426300.0 ;
      RECT  24450.0 424800.0 32850.0 423900.0 ;
      RECT  32850.0 427500.0 34050.0 426300.0 ;
      RECT  32850.0 425100.0 34050.0 423900.0 ;
      RECT  32850.0 425100.0 34050.0 423900.0 ;
      RECT  32850.0 427500.0 34050.0 426300.0 ;
      RECT  23250.0 427500.0 24450.0 426300.0 ;
      RECT  23250.0 425100.0 24450.0 423900.0 ;
      RECT  23250.0 425100.0 24450.0 423900.0 ;
      RECT  23250.0 427500.0 24450.0 426300.0 ;
      RECT  23250.0 422700.0 24450.0 421500.0 ;
      RECT  33450.0 422700.0 34650.0 421500.0 ;
      RECT  27750.0 426900.0 28950.0 425700.0 ;
      RECT  27750.0 426900.0 28950.0 425700.0 ;
      RECT  27900.0 424350.0 28800.0 423450.0 ;
      RECT  35550.0 429300.0 36450.0 419700.0 ;
      RECT  21450.0 429300.0 22350.0 419700.0 ;
      RECT  27750.0 425700.0 28950.0 426900.0 ;
      RECT  21900.0 413100.0 23850.0 411900.0 ;
      RECT  34050.0 413100.0 36000.0 411900.0 ;
      RECT  23250.0 417900.0 21450.0 416700.0 ;
      RECT  32850.0 417900.0 36450.0 416700.0 ;
      RECT  24450.0 415200.0 32850.0 414300.0 ;
      RECT  32850.0 417900.0 34050.0 416700.0 ;
      RECT  32850.0 415500.0 34050.0 414300.0 ;
      RECT  32850.0 415500.0 34050.0 414300.0 ;
      RECT  32850.0 417900.0 34050.0 416700.0 ;
      RECT  23250.0 417900.0 24450.0 416700.0 ;
      RECT  23250.0 415500.0 24450.0 414300.0 ;
      RECT  23250.0 415500.0 24450.0 414300.0 ;
      RECT  23250.0 417900.0 24450.0 416700.0 ;
      RECT  23250.0 413100.0 24450.0 411900.0 ;
      RECT  33450.0 413100.0 34650.0 411900.0 ;
      RECT  27750.0 417300.0 28950.0 416100.0 ;
      RECT  27750.0 417300.0 28950.0 416100.0 ;
      RECT  27900.0 414750.0 28800.0 413850.0 ;
      RECT  35550.0 419700.0 36450.0 410100.0 ;
      RECT  21450.0 419700.0 22350.0 410100.0 ;
      RECT  27750.0 416100.0 28950.0 417300.0 ;
      RECT  43050.0 414900.0 44250.0 416100.0 ;
      RECT  43050.0 424500.0 44250.0 425700.0 ;
      RECT  27750.0 423300.0 28950.0 424500.0 ;
      RECT  43050.0 412500.0 44250.0 413700.0 ;
      RECT  27900.0 410100.0 28800.0 413850.0 ;
      RECT  35550.0 410100.0 36450.0 429300.0 ;
      RECT  21450.0 410100.0 22350.0 429300.0 ;
      RECT  49650.0 410100.0 50550.0 429300.0 ;
      RECT  16500.0 396000.0 6300.0 381300.0 ;
      RECT  16500.0 396000.0 6300.0 410100.0 ;
      RECT  16500.0 424200.0 6300.0 410100.0 ;
      RECT  17100.0 398100.0 5700.0 399300.0 ;
      RECT  17100.0 420900.0 5700.0 422100.0 ;
      RECT  17100.0 409500.0 5700.0 410400.0 ;
      RECT  22350.0 398100.0 21150.0 399300.0 ;
      RECT  22350.0 420900.0 21150.0 422100.0 ;
      RECT  22350.0 410100.0 21150.0 411300.0 ;
      RECT  22350.0 370500.0 21150.0 371700.0 ;
      RECT  21300.0 426300.0 22500.0 427500.0 ;
      RECT  5700.0 426300.0 6900.0 427500.0 ;
      RECT  28950.0 396900.0 27750.0 398100.0 ;
      RECT  19050.0 383400.0 20250.0 384600.0 ;
      RECT  19050.0 375900.0 20250.0 377100.0 ;
      RECT  12300.0 375900.0 13500.0 377100.0 ;
      RECT  44250.0 362100.0 43350.0 412500.0 ;
      RECT  28800.0 362100.0 27900.0 375450.0 ;
      RECT  4200.0 362100.0 3300.0 424650.0 ;
      RECT  36450.0 362100.0 35550.0 410100.0 ;
      RECT  22350.0 362100.0 21450.0 381300.0 ;
      RECT  50550.0 362100.0 49650.0 410100.0 ;
      RECT  44550.0 285450.0 43350.0 284250.0 ;
      RECT  44550.0 244650.0 43350.0 243450.0 ;
      RECT  33900.0 205650.0 32700.0 204450.0 ;
      RECT  29550.0 285450.0 28350.0 284250.0 ;
      RECT  26850.0 290850.0 25650.0 289650.0 ;
      RECT  30300.0 328200.0 29100.0 327000.0 ;
      RECT  27600.0 331200.0 26400.0 330000.0 ;
      RECT  41400.0 304350.0 40200.0 303150.0 ;
      RECT  43350.0 301650.0 42150.0 300450.0 ;
      RECT  45300.0 293550.0 44100.0 292350.0 ;
      RECT  13200.0 304350.0 12000.0 303150.0 ;
      RECT  15150.0 293550.0 13950.0 292350.0 ;
      RECT  17100.0 296250.0 15900.0 295050.0 ;
      RECT  29550.0 322500.0 28350.0 323700.0 ;
      RECT  30300.0 339600.0 29100.0 340800.0 ;
      RECT  16050.0 362100.0 14850.0 363300.0 ;
      RECT  28950.0 342300.0 27750.0 343500.0 ;
      RECT  50700.0 288150.0 49500.0 286950.0 ;
      RECT  36600.0 298950.0 35400.0 297750.0 ;
      RECT  22500.0 288150.0 21300.0 286950.0 ;
      RECT  8400.0 298950.0 7200.0 297750.0 ;
      RECT  44250.0 202200.0 43050.0 205800.0 ;
      RECT  36450.0 202200.0 35550.0 203100.0 ;
      RECT  50550.0 202200.0 49650.0 203100.0 ;
      RECT  55950.0 297750.0 54750.0 298950.0 ;
   LAYER  metal2 ;
      RECT  169050.0 340200.0 169950.0 342900.0 ;
      RECT  166350.0 360000.0 167250.0 362700.0 ;
      RECT  160950.0 320400.0 161850.0 323100.0 ;
      RECT  158250.0 337500.0 159150.0 340200.0 ;
      RECT  163650.0 301050.0 164550.0 303750.0 ;
      RECT  155550.0 282150.0 156450.0 284850.0 ;
      RECT  50100.0 297900.0 55350.0 298800.0 ;
      RECT  150150.0 284850.0 151050.0 287550.0 ;
      RECT  155550.0 0.0 156450.0 444600.0 ;
      RECT  158250.0 0.0 159150.0 444600.0 ;
      RECT  160950.0 0.0 161850.0 444600.0 ;
      RECT  163650.0 0.0 164550.0 444600.0 ;
      RECT  166350.0 0.0 167250.0 444600.0 ;
      RECT  169050.0 0.0 169950.0 444600.0 ;
      RECT  134850.0 34800.0 135750.0 199200.0 ;
      RECT  137550.0 34800.0 138450.0 199200.0 ;
      RECT  140250.0 34800.0 141150.0 199200.0 ;
      RECT  142950.0 34800.0 143850.0 199200.0 ;
      RECT  180450.0 5850.0 181350.0 6750.0 ;
      RECT  177300.0 5850.0 180900.0 6750.0 ;
      RECT  180450.0 6300.0 181350.0 8100.0 ;
      RECT  190650.0 5850.0 191550.0 6750.0 ;
      RECT  187500.0 5850.0 191100.0 6750.0 ;
      RECT  190650.0 6300.0 191550.0 8100.0 ;
      RECT  102900.0 424800.0 103800.0 426900.0 ;
      RECT  175800.0 199200.0 186000.0 213300.0 ;
      RECT  175800.0 227400.0 186000.0 213300.0 ;
      RECT  175800.0 227400.0 186000.0 241500.0 ;
      RECT  175800.0 255600.0 186000.0 241500.0 ;
      RECT  175800.0 255600.0 186000.0 269700.0 ;
      RECT  175800.0 283800.0 186000.0 269700.0 ;
      RECT  175800.0 283800.0 186000.0 297900.0 ;
      RECT  175800.0 312000.0 186000.0 297900.0 ;
      RECT  175800.0 312000.0 186000.0 326100.0 ;
      RECT  175800.0 340200.0 186000.0 326100.0 ;
      RECT  175800.0 340200.0 186000.0 354300.0 ;
      RECT  175800.0 368400.0 186000.0 354300.0 ;
      RECT  175800.0 368400.0 186000.0 382500.0 ;
      RECT  175800.0 396600.0 186000.0 382500.0 ;
      RECT  175800.0 396600.0 186000.0 410700.0 ;
      RECT  175800.0 424800.0 186000.0 410700.0 ;
      RECT  186000.0 199200.0 196200.0 213300.0 ;
      RECT  186000.0 227400.0 196200.0 213300.0 ;
      RECT  186000.0 227400.0 196200.0 241500.0 ;
      RECT  186000.0 255600.0 196200.0 241500.0 ;
      RECT  186000.0 255600.0 196200.0 269700.0 ;
      RECT  186000.0 283800.0 196200.0 269700.0 ;
      RECT  186000.0 283800.0 196200.0 297900.0 ;
      RECT  186000.0 312000.0 196200.0 297900.0 ;
      RECT  186000.0 312000.0 196200.0 326100.0 ;
      RECT  186000.0 340200.0 196200.0 326100.0 ;
      RECT  186000.0 340200.0 196200.0 354300.0 ;
      RECT  186000.0 368400.0 196200.0 354300.0 ;
      RECT  186000.0 368400.0 196200.0 382500.0 ;
      RECT  186000.0 396600.0 196200.0 382500.0 ;
      RECT  186000.0 396600.0 196200.0 410700.0 ;
      RECT  186000.0 424800.0 196200.0 410700.0 ;
      RECT  178800.0 199200.0 180000.0 424800.0 ;
      RECT  181800.0 199200.0 183000.0 424800.0 ;
      RECT  189000.0 199200.0 190200.0 424800.0 ;
      RECT  192000.0 199200.0 193200.0 424800.0 ;
      RECT  185400.0 199200.0 186600.0 424800.0 ;
      RECT  178800.0 427200.0 180000.0 428400.0 ;
      RECT  181200.0 427200.0 182850.0 428400.0 ;
      RECT  178800.0 436200.0 180000.0 437400.0 ;
      RECT  181950.0 436200.0 184800.0 437400.0 ;
      RECT  178800.0 427200.0 180000.0 428400.0 ;
      RECT  181200.0 427200.0 182400.0 428400.0 ;
      RECT  178800.0 436200.0 180000.0 437400.0 ;
      RECT  183600.0 436200.0 184800.0 437400.0 ;
      RECT  178950.0 424800.0 179850.0 444600.0 ;
      RECT  181950.0 424800.0 182850.0 444600.0 ;
      RECT  189000.0 427200.0 190200.0 428400.0 ;
      RECT  191400.0 427200.0 193050.0 428400.0 ;
      RECT  189000.0 436200.0 190200.0 437400.0 ;
      RECT  192150.0 436200.0 195000.0 437400.0 ;
      RECT  189000.0 427200.0 190200.0 428400.0 ;
      RECT  191400.0 427200.0 192600.0 428400.0 ;
      RECT  189000.0 436200.0 190200.0 437400.0 ;
      RECT  193800.0 436200.0 195000.0 437400.0 ;
      RECT  189150.0 424800.0 190050.0 444600.0 ;
      RECT  192150.0 424800.0 193050.0 444600.0 ;
      RECT  178950.0 424800.0 179850.0 444600.0 ;
      RECT  181950.0 424800.0 182850.0 444600.0 ;
      RECT  189150.0 424800.0 190050.0 444600.0 ;
      RECT  192150.0 424800.0 193050.0 444600.0 ;
      RECT  175800.0 150300.0 186000.0 199200.0 ;
      RECT  186000.0 150300.0 196200.0 199200.0 ;
      RECT  178800.0 150300.0 180000.0 163500.0 ;
      RECT  181800.0 150300.0 183000.0 163500.0 ;
      RECT  189000.0 150300.0 190200.0 163500.0 ;
      RECT  192000.0 150300.0 193200.0 163500.0 ;
      RECT  175800.0 90000.0 186000.0 150300.0 ;
      RECT  186000.0 90000.0 196200.0 150300.0 ;
      RECT  180300.0 90000.0 181500.0 92700.0 ;
      RECT  190500.0 90000.0 191700.0 92700.0 ;
      RECT  178800.0 148200.0 180000.0 150300.0 ;
      RECT  181800.0 142800.0 183000.0 150300.0 ;
      RECT  189000.0 148200.0 190200.0 150300.0 ;
      RECT  192000.0 142800.0 193200.0 150300.0 ;
      RECT  175800.0 30000.0 186000.0 90000.0 ;
      RECT  196200.0 30000.0 186000.0 90000.0 ;
      RECT  180300.0 30000.0 181500.0 31200.0 ;
      RECT  190500.0 30000.0 191700.0 31200.0 ;
      RECT  180300.0 88800.0 181500.0 90000.0 ;
      RECT  177600.0 85500.0 178800.0 90000.0 ;
      RECT  190500.0 88800.0 191700.0 90000.0 ;
      RECT  193200.0 85500.0 194400.0 90000.0 ;
      RECT  185400.0 30000.0 186600.0 90000.0 ;
      RECT  175800.0 30000.0 186000.0 8100.0 ;
      RECT  186000.0 30000.0 196200.0 8100.0 ;
      RECT  180300.0 15000.0 181500.0 8100.0 ;
      RECT  190500.0 15000.0 191700.0 8100.0 ;
      RECT  180300.0 30000.0 181500.0 28500.0 ;
      RECT  190500.0 30000.0 191700.0 28500.0 ;
      RECT  59400.0 86400.0 60300.0 424800.0 ;
      RECT  61500.0 86400.0 62400.0 424800.0 ;
      RECT  63600.0 86400.0 64500.0 424800.0 ;
      RECT  65700.0 86400.0 66600.0 424800.0 ;
      RECT  67800.0 86400.0 68700.0 424800.0 ;
      RECT  69900.0 86400.0 70800.0 424800.0 ;
      RECT  72000.0 86400.0 72900.0 424800.0 ;
      RECT  74100.0 86400.0 75000.0 424800.0 ;
      RECT  106200.0 86400.0 105300.0 141000.0 ;
      RECT  103200.0 86400.0 102300.0 141000.0 ;
      RECT  112200.0 86400.0 111300.0 141000.0 ;
      RECT  109200.0 86400.0 108300.0 141000.0 ;
      RECT  95850.0 93750.0 94950.0 94650.0 ;
      RECT  93450.0 93750.0 92550.0 94650.0 ;
      RECT  95850.0 94200.0 94950.0 97350.0 ;
      RECT  95400.0 93750.0 93000.0 94650.0 ;
      RECT  93450.0 89550.0 92550.0 94200.0 ;
      RECT  96000.0 97350.0 94800.0 98550.0 ;
      RECT  93600.0 88350.0 92400.0 89550.0 ;
      RECT  92400.0 93600.0 93600.0 94800.0 ;
      RECT  95850.0 107250.0 94950.0 106350.0 ;
      RECT  93450.0 107250.0 92550.0 106350.0 ;
      RECT  95850.0 106800.0 94950.0 103650.0 ;
      RECT  95400.0 107250.0 93000.0 106350.0 ;
      RECT  93450.0 111450.0 92550.0 106800.0 ;
      RECT  96000.0 103650.0 94800.0 102450.0 ;
      RECT  93600.0 112650.0 92400.0 111450.0 ;
      RECT  92400.0 107400.0 93600.0 106200.0 ;
      RECT  95850.0 121950.0 94950.0 122850.0 ;
      RECT  93450.0 121950.0 92550.0 122850.0 ;
      RECT  95850.0 122400.0 94950.0 125550.0 ;
      RECT  95400.0 121950.0 93000.0 122850.0 ;
      RECT  93450.0 117750.0 92550.0 122400.0 ;
      RECT  96000.0 125550.0 94800.0 126750.0 ;
      RECT  93600.0 116550.0 92400.0 117750.0 ;
      RECT  92400.0 121800.0 93600.0 123000.0 ;
      RECT  95850.0 135450.0 94950.0 134550.0 ;
      RECT  93450.0 135450.0 92550.0 134550.0 ;
      RECT  95850.0 135000.0 94950.0 131850.0 ;
      RECT  95400.0 135450.0 93000.0 134550.0 ;
      RECT  93450.0 139650.0 92550.0 135000.0 ;
      RECT  96000.0 131850.0 94800.0 130650.0 ;
      RECT  93600.0 140850.0 92400.0 139650.0 ;
      RECT  92400.0 135600.0 93600.0 134400.0 ;
      RECT  111150.0 97200.0 112350.0 98400.0 ;
      RECT  129750.0 92250.0 130950.0 93450.0 ;
      RECT  108150.0 111300.0 109350.0 112500.0 ;
      RECT  126750.0 107550.0 127950.0 108750.0 ;
      RECT  129750.0 116100.0 130950.0 117300.0 ;
      RECT  105150.0 116100.0 106350.0 117300.0 ;
      RECT  126750.0 130200.0 127950.0 131400.0 ;
      RECT  102150.0 130200.0 103350.0 131400.0 ;
      RECT  111150.0 93600.0 112350.0 94800.0 ;
      RECT  108150.0 90900.0 109350.0 92100.0 ;
      RECT  105150.0 106200.0 106350.0 107400.0 ;
      RECT  108150.0 108900.0 109350.0 110100.0 ;
      RECT  111150.0 121800.0 112350.0 123000.0 ;
      RECT  102150.0 119100.0 103350.0 120300.0 ;
      RECT  105150.0 134400.0 106350.0 135600.0 ;
      RECT  102150.0 137100.0 103350.0 138300.0 ;
      RECT  130800.0 86400.0 129900.0 141000.0 ;
      RECT  127800.0 86400.0 126900.0 141000.0 ;
      RECT  106200.0 142800.0 105300.0 197400.0 ;
      RECT  103200.0 142800.0 102300.0 197400.0 ;
      RECT  112200.0 142800.0 111300.0 197400.0 ;
      RECT  109200.0 142800.0 108300.0 197400.0 ;
      RECT  95850.0 150150.0 94950.0 151050.0 ;
      RECT  93450.0 150150.0 92550.0 151050.0 ;
      RECT  95850.0 150600.0 94950.0 153750.0 ;
      RECT  95400.0 150150.0 93000.0 151050.0 ;
      RECT  93450.0 145950.0 92550.0 150600.0 ;
      RECT  96000.0 153750.0 94800.0 154950.0 ;
      RECT  93600.0 144750.0 92400.0 145950.0 ;
      RECT  92400.0 150000.0 93600.0 151200.0 ;
      RECT  95850.0 163650.0 94950.0 162750.0 ;
      RECT  93450.0 163650.0 92550.0 162750.0 ;
      RECT  95850.0 163200.0 94950.0 160050.0 ;
      RECT  95400.0 163650.0 93000.0 162750.0 ;
      RECT  93450.0 167850.0 92550.0 163200.0 ;
      RECT  96000.0 160050.0 94800.0 158850.0 ;
      RECT  93600.0 169050.0 92400.0 167850.0 ;
      RECT  92400.0 163800.0 93600.0 162600.0 ;
      RECT  95850.0 178350.0 94950.0 179250.0 ;
      RECT  93450.0 178350.0 92550.0 179250.0 ;
      RECT  95850.0 178800.0 94950.0 181950.0 ;
      RECT  95400.0 178350.0 93000.0 179250.0 ;
      RECT  93450.0 174150.0 92550.0 178800.0 ;
      RECT  96000.0 181950.0 94800.0 183150.0 ;
      RECT  93600.0 172950.0 92400.0 174150.0 ;
      RECT  92400.0 178200.0 93600.0 179400.0 ;
      RECT  95850.0 191850.0 94950.0 190950.0 ;
      RECT  93450.0 191850.0 92550.0 190950.0 ;
      RECT  95850.0 191400.0 94950.0 188250.0 ;
      RECT  95400.0 191850.0 93000.0 190950.0 ;
      RECT  93450.0 196050.0 92550.0 191400.0 ;
      RECT  96000.0 188250.0 94800.0 187050.0 ;
      RECT  93600.0 197250.0 92400.0 196050.0 ;
      RECT  92400.0 192000.0 93600.0 190800.0 ;
      RECT  111150.0 153600.0 112350.0 154800.0 ;
      RECT  129750.0 148650.0 130950.0 149850.0 ;
      RECT  108150.0 167700.0 109350.0 168900.0 ;
      RECT  126750.0 163950.0 127950.0 165150.0 ;
      RECT  129750.0 172500.0 130950.0 173700.0 ;
      RECT  105150.0 172500.0 106350.0 173700.0 ;
      RECT  126750.0 186600.0 127950.0 187800.0 ;
      RECT  102150.0 186600.0 103350.0 187800.0 ;
      RECT  111150.0 150000.0 112350.0 151200.0 ;
      RECT  108150.0 147300.0 109350.0 148500.0 ;
      RECT  105150.0 162600.0 106350.0 163800.0 ;
      RECT  108150.0 165300.0 109350.0 166500.0 ;
      RECT  111150.0 178200.0 112350.0 179400.0 ;
      RECT  102150.0 175500.0 103350.0 176700.0 ;
      RECT  105150.0 190800.0 106350.0 192000.0 ;
      RECT  102150.0 193500.0 103350.0 194700.0 ;
      RECT  130800.0 142800.0 129900.0 197400.0 ;
      RECT  127800.0 142800.0 126900.0 197400.0 ;
      RECT  80550.0 206550.0 81450.0 207450.0 ;
      RECT  82950.0 206550.0 83850.0 207450.0 ;
      RECT  80550.0 207000.0 81450.0 210150.0 ;
      RECT  81000.0 206550.0 83400.0 207450.0 ;
      RECT  82950.0 202350.0 83850.0 207000.0 ;
      RECT  80400.0 210150.0 81600.0 211350.0 ;
      RECT  82800.0 201150.0 84000.0 202350.0 ;
      RECT  84000.0 206400.0 82800.0 207600.0 ;
      RECT  80550.0 220050.0 81450.0 219150.0 ;
      RECT  82950.0 220050.0 83850.0 219150.0 ;
      RECT  80550.0 219600.0 81450.0 216450.0 ;
      RECT  81000.0 220050.0 83400.0 219150.0 ;
      RECT  82950.0 224250.0 83850.0 219600.0 ;
      RECT  80400.0 216450.0 81600.0 215250.0 ;
      RECT  82800.0 225450.0 84000.0 224250.0 ;
      RECT  84000.0 220200.0 82800.0 219000.0 ;
      RECT  80550.0 234750.0 81450.0 235650.0 ;
      RECT  82950.0 234750.0 83850.0 235650.0 ;
      RECT  80550.0 235200.0 81450.0 238350.0 ;
      RECT  81000.0 234750.0 83400.0 235650.0 ;
      RECT  82950.0 230550.0 83850.0 235200.0 ;
      RECT  80400.0 238350.0 81600.0 239550.0 ;
      RECT  82800.0 229350.0 84000.0 230550.0 ;
      RECT  84000.0 234600.0 82800.0 235800.0 ;
      RECT  80550.0 248250.0 81450.0 247350.0 ;
      RECT  82950.0 248250.0 83850.0 247350.0 ;
      RECT  80550.0 247800.0 81450.0 244650.0 ;
      RECT  81000.0 248250.0 83400.0 247350.0 ;
      RECT  82950.0 252450.0 83850.0 247800.0 ;
      RECT  80400.0 244650.0 81600.0 243450.0 ;
      RECT  82800.0 253650.0 84000.0 252450.0 ;
      RECT  84000.0 248400.0 82800.0 247200.0 ;
      RECT  80550.0 262950.0 81450.0 263850.0 ;
      RECT  82950.0 262950.0 83850.0 263850.0 ;
      RECT  80550.0 263400.0 81450.0 266550.0 ;
      RECT  81000.0 262950.0 83400.0 263850.0 ;
      RECT  82950.0 258750.0 83850.0 263400.0 ;
      RECT  80400.0 266550.0 81600.0 267750.0 ;
      RECT  82800.0 257550.0 84000.0 258750.0 ;
      RECT  84000.0 262800.0 82800.0 264000.0 ;
      RECT  80550.0 276450.0 81450.0 275550.0 ;
      RECT  82950.0 276450.0 83850.0 275550.0 ;
      RECT  80550.0 276000.0 81450.0 272850.0 ;
      RECT  81000.0 276450.0 83400.0 275550.0 ;
      RECT  82950.0 280650.0 83850.0 276000.0 ;
      RECT  80400.0 272850.0 81600.0 271650.0 ;
      RECT  82800.0 281850.0 84000.0 280650.0 ;
      RECT  84000.0 276600.0 82800.0 275400.0 ;
      RECT  80550.0 291150.0 81450.0 292050.0 ;
      RECT  82950.0 291150.0 83850.0 292050.0 ;
      RECT  80550.0 291600.0 81450.0 294750.0 ;
      RECT  81000.0 291150.0 83400.0 292050.0 ;
      RECT  82950.0 286950.0 83850.0 291600.0 ;
      RECT  80400.0 294750.0 81600.0 295950.0 ;
      RECT  82800.0 285750.0 84000.0 286950.0 ;
      RECT  84000.0 291000.0 82800.0 292200.0 ;
      RECT  80550.0 304650.0 81450.0 303750.0 ;
      RECT  82950.0 304650.0 83850.0 303750.0 ;
      RECT  80550.0 304200.0 81450.0 301050.0 ;
      RECT  81000.0 304650.0 83400.0 303750.0 ;
      RECT  82950.0 308850.0 83850.0 304200.0 ;
      RECT  80400.0 301050.0 81600.0 299850.0 ;
      RECT  82800.0 310050.0 84000.0 308850.0 ;
      RECT  84000.0 304800.0 82800.0 303600.0 ;
      RECT  80550.0 319350.0 81450.0 320250.0 ;
      RECT  82950.0 319350.0 83850.0 320250.0 ;
      RECT  80550.0 319800.0 81450.0 322950.0 ;
      RECT  81000.0 319350.0 83400.0 320250.0 ;
      RECT  82950.0 315150.0 83850.0 319800.0 ;
      RECT  80400.0 322950.0 81600.0 324150.0 ;
      RECT  82800.0 313950.0 84000.0 315150.0 ;
      RECT  84000.0 319200.0 82800.0 320400.0 ;
      RECT  80550.0 332850.0 81450.0 331950.0 ;
      RECT  82950.0 332850.0 83850.0 331950.0 ;
      RECT  80550.0 332400.0 81450.0 329250.0 ;
      RECT  81000.0 332850.0 83400.0 331950.0 ;
      RECT  82950.0 337050.0 83850.0 332400.0 ;
      RECT  80400.0 329250.0 81600.0 328050.0 ;
      RECT  82800.0 338250.0 84000.0 337050.0 ;
      RECT  84000.0 333000.0 82800.0 331800.0 ;
      RECT  80550.0 347550.0 81450.0 348450.0 ;
      RECT  82950.0 347550.0 83850.0 348450.0 ;
      RECT  80550.0 348000.0 81450.0 351150.0 ;
      RECT  81000.0 347550.0 83400.0 348450.0 ;
      RECT  82950.0 343350.0 83850.0 348000.0 ;
      RECT  80400.0 351150.0 81600.0 352350.0 ;
      RECT  82800.0 342150.0 84000.0 343350.0 ;
      RECT  84000.0 347400.0 82800.0 348600.0 ;
      RECT  80550.0 361050.0 81450.0 360150.0 ;
      RECT  82950.0 361050.0 83850.0 360150.0 ;
      RECT  80550.0 360600.0 81450.0 357450.0 ;
      RECT  81000.0 361050.0 83400.0 360150.0 ;
      RECT  82950.0 365250.0 83850.0 360600.0 ;
      RECT  80400.0 357450.0 81600.0 356250.0 ;
      RECT  82800.0 366450.0 84000.0 365250.0 ;
      RECT  84000.0 361200.0 82800.0 360000.0 ;
      RECT  80550.0 375750.0 81450.0 376650.0 ;
      RECT  82950.0 375750.0 83850.0 376650.0 ;
      RECT  80550.0 376200.0 81450.0 379350.0 ;
      RECT  81000.0 375750.0 83400.0 376650.0 ;
      RECT  82950.0 371550.0 83850.0 376200.0 ;
      RECT  80400.0 379350.0 81600.0 380550.0 ;
      RECT  82800.0 370350.0 84000.0 371550.0 ;
      RECT  84000.0 375600.0 82800.0 376800.0 ;
      RECT  80550.0 389250.0 81450.0 388350.0 ;
      RECT  82950.0 389250.0 83850.0 388350.0 ;
      RECT  80550.0 388800.0 81450.0 385650.0 ;
      RECT  81000.0 389250.0 83400.0 388350.0 ;
      RECT  82950.0 393450.0 83850.0 388800.0 ;
      RECT  80400.0 385650.0 81600.0 384450.0 ;
      RECT  82800.0 394650.0 84000.0 393450.0 ;
      RECT  84000.0 389400.0 82800.0 388200.0 ;
      RECT  80550.0 403950.0 81450.0 404850.0 ;
      RECT  82950.0 403950.0 83850.0 404850.0 ;
      RECT  80550.0 404400.0 81450.0 407550.0 ;
      RECT  81000.0 403950.0 83400.0 404850.0 ;
      RECT  82950.0 399750.0 83850.0 404400.0 ;
      RECT  80400.0 407550.0 81600.0 408750.0 ;
      RECT  82800.0 398550.0 84000.0 399750.0 ;
      RECT  84000.0 403800.0 82800.0 405000.0 ;
      RECT  80550.0 417450.0 81450.0 416550.0 ;
      RECT  82950.0 417450.0 83850.0 416550.0 ;
      RECT  80550.0 417000.0 81450.0 413850.0 ;
      RECT  81000.0 417450.0 83400.0 416550.0 ;
      RECT  82950.0 421650.0 83850.0 417000.0 ;
      RECT  80400.0 413850.0 81600.0 412650.0 ;
      RECT  82800.0 422850.0 84000.0 421650.0 ;
      RECT  84000.0 417600.0 82800.0 416400.0 ;
      RECT  60450.0 92250.0 59250.0 93450.0 ;
      RECT  62550.0 107550.0 61350.0 108750.0 ;
      RECT  64650.0 120450.0 63450.0 121650.0 ;
      RECT  66750.0 135750.0 65550.0 136950.0 ;
      RECT  68850.0 148650.0 67650.0 149850.0 ;
      RECT  70950.0 163950.0 69750.0 165150.0 ;
      RECT  73050.0 176850.0 71850.0 178050.0 ;
      RECT  75150.0 192150.0 73950.0 193350.0 ;
      RECT  60450.0 206400.0 59250.0 207600.0 ;
      RECT  68850.0 203700.0 67650.0 204900.0 ;
      RECT  60450.0 219000.0 59250.0 220200.0 ;
      RECT  70950.0 221700.0 69750.0 222900.0 ;
      RECT  60450.0 234600.0 59250.0 235800.0 ;
      RECT  73050.0 231900.0 71850.0 233100.0 ;
      RECT  60450.0 247200.0 59250.0 248400.0 ;
      RECT  75150.0 249900.0 73950.0 251100.0 ;
      RECT  62550.0 262800.0 61350.0 264000.0 ;
      RECT  68850.0 260100.0 67650.0 261300.0 ;
      RECT  62550.0 275400.0 61350.0 276600.0 ;
      RECT  70950.0 278100.0 69750.0 279300.0 ;
      RECT  62550.0 291000.0 61350.0 292200.0 ;
      RECT  73050.0 288300.0 71850.0 289500.0 ;
      RECT  62550.0 303600.0 61350.0 304800.0 ;
      RECT  75150.0 306300.0 73950.0 307500.0 ;
      RECT  64650.0 319200.0 63450.0 320400.0 ;
      RECT  68850.0 316500.0 67650.0 317700.0 ;
      RECT  64650.0 331800.0 63450.0 333000.0 ;
      RECT  70950.0 334500.0 69750.0 335700.0 ;
      RECT  64650.0 347400.0 63450.0 348600.0 ;
      RECT  73050.0 344700.0 71850.0 345900.0 ;
      RECT  64650.0 360000.0 63450.0 361200.0 ;
      RECT  75150.0 362700.0 73950.0 363900.0 ;
      RECT  66750.0 375600.0 65550.0 376800.0 ;
      RECT  68850.0 372900.0 67650.0 374100.0 ;
      RECT  66750.0 388200.0 65550.0 389400.0 ;
      RECT  70950.0 390900.0 69750.0 392100.0 ;
      RECT  66750.0 403800.0 65550.0 405000.0 ;
      RECT  73050.0 401100.0 71850.0 402300.0 ;
      RECT  66750.0 416400.0 65550.0 417600.0 ;
      RECT  75150.0 419100.0 73950.0 420300.0 ;
      RECT  129900.0 86400.0 130800.0 141000.0 ;
      RECT  126900.0 86400.0 127800.0 141000.0 ;
      RECT  129900.0 142800.0 130800.0 197400.0 ;
      RECT  126900.0 142800.0 127800.0 197400.0 ;
      RECT  104850.0 203850.0 105750.0 204750.0 ;
      RECT  104850.0 203400.0 105750.0 204300.0 ;
      RECT  105300.0 203850.0 121500.0 204750.0 ;
      RECT  104850.0 221850.0 105750.0 222750.0 ;
      RECT  104850.0 222300.0 105750.0 223200.0 ;
      RECT  105300.0 221850.0 121500.0 222750.0 ;
      RECT  104850.0 232050.0 105750.0 232950.0 ;
      RECT  104850.0 231600.0 105750.0 232500.0 ;
      RECT  105300.0 232050.0 121500.0 232950.0 ;
      RECT  104850.0 250050.0 105750.0 250950.0 ;
      RECT  104850.0 250500.0 105750.0 251400.0 ;
      RECT  105300.0 250050.0 121500.0 250950.0 ;
      RECT  104850.0 260250.0 105750.0 261150.0 ;
      RECT  104850.0 259800.0 105750.0 260700.0 ;
      RECT  105300.0 260250.0 121500.0 261150.0 ;
      RECT  104850.0 278250.0 105750.0 279150.0 ;
      RECT  104850.0 278700.0 105750.0 279600.0 ;
      RECT  105300.0 278250.0 121500.0 279150.0 ;
      RECT  104850.0 288450.0 105750.0 289350.0 ;
      RECT  104850.0 288000.0 105750.0 288900.0 ;
      RECT  105300.0 288450.0 121500.0 289350.0 ;
      RECT  104850.0 306450.0 105750.0 307350.0 ;
      RECT  104850.0 306900.0 105750.0 307800.0 ;
      RECT  105300.0 306450.0 121500.0 307350.0 ;
      RECT  104850.0 316650.0 105750.0 317550.0 ;
      RECT  104850.0 316200.0 105750.0 317100.0 ;
      RECT  105300.0 316650.0 121500.0 317550.0 ;
      RECT  104850.0 334650.0 105750.0 335550.0 ;
      RECT  104850.0 335100.0 105750.0 336000.0 ;
      RECT  105300.0 334650.0 121500.0 335550.0 ;
      RECT  104850.0 344850.0 105750.0 345750.0 ;
      RECT  104850.0 344400.0 105750.0 345300.0 ;
      RECT  105300.0 344850.0 121500.0 345750.0 ;
      RECT  104850.0 362850.0 105750.0 363750.0 ;
      RECT  104850.0 363300.0 105750.0 364200.0 ;
      RECT  105300.0 362850.0 121500.0 363750.0 ;
      RECT  104850.0 373050.0 105750.0 373950.0 ;
      RECT  104850.0 372600.0 105750.0 373500.0 ;
      RECT  105300.0 373050.0 121500.0 373950.0 ;
      RECT  104850.0 391050.0 105750.0 391950.0 ;
      RECT  104850.0 391500.0 105750.0 392400.0 ;
      RECT  105300.0 391050.0 121500.0 391950.0 ;
      RECT  104850.0 401250.0 105750.0 402150.0 ;
      RECT  104850.0 400800.0 105750.0 401700.0 ;
      RECT  105300.0 401250.0 121500.0 402150.0 ;
      RECT  104850.0 419250.0 105750.0 420150.0 ;
      RECT  104850.0 419700.0 105750.0 420600.0 ;
      RECT  105300.0 419250.0 121500.0 420150.0 ;
      RECT  120450.0 206550.0 121350.0 207450.0 ;
      RECT  122850.0 206550.0 123750.0 207450.0 ;
      RECT  120450.0 207000.0 121350.0 210150.0 ;
      RECT  120900.0 206550.0 123300.0 207450.0 ;
      RECT  122850.0 202350.0 123750.0 207000.0 ;
      RECT  120300.0 210150.0 121500.0 211350.0 ;
      RECT  122700.0 201150.0 123900.0 202350.0 ;
      RECT  123900.0 206400.0 122700.0 207600.0 ;
      RECT  102750.0 205050.0 103950.0 206250.0 ;
      RECT  104700.0 202800.0 105900.0 204000.0 ;
      RECT  121500.0 203700.0 120300.0 204900.0 ;
      RECT  120450.0 220050.0 121350.0 219150.0 ;
      RECT  122850.0 220050.0 123750.0 219150.0 ;
      RECT  120450.0 219600.0 121350.0 216450.0 ;
      RECT  120900.0 220050.0 123300.0 219150.0 ;
      RECT  122850.0 224250.0 123750.0 219600.0 ;
      RECT  120300.0 216450.0 121500.0 215250.0 ;
      RECT  122700.0 225450.0 123900.0 224250.0 ;
      RECT  123900.0 220200.0 122700.0 219000.0 ;
      RECT  102750.0 220350.0 103950.0 221550.0 ;
      RECT  104700.0 222600.0 105900.0 223800.0 ;
      RECT  121500.0 221700.0 120300.0 222900.0 ;
      RECT  120450.0 234750.0 121350.0 235650.0 ;
      RECT  122850.0 234750.0 123750.0 235650.0 ;
      RECT  120450.0 235200.0 121350.0 238350.0 ;
      RECT  120900.0 234750.0 123300.0 235650.0 ;
      RECT  122850.0 230550.0 123750.0 235200.0 ;
      RECT  120300.0 238350.0 121500.0 239550.0 ;
      RECT  122700.0 229350.0 123900.0 230550.0 ;
      RECT  123900.0 234600.0 122700.0 235800.0 ;
      RECT  102750.0 233250.0 103950.0 234450.0 ;
      RECT  104700.0 231000.0 105900.0 232200.0 ;
      RECT  121500.0 231900.0 120300.0 233100.0 ;
      RECT  120450.0 248250.0 121350.0 247350.0 ;
      RECT  122850.0 248250.0 123750.0 247350.0 ;
      RECT  120450.0 247800.0 121350.0 244650.0 ;
      RECT  120900.0 248250.0 123300.0 247350.0 ;
      RECT  122850.0 252450.0 123750.0 247800.0 ;
      RECT  120300.0 244650.0 121500.0 243450.0 ;
      RECT  122700.0 253650.0 123900.0 252450.0 ;
      RECT  123900.0 248400.0 122700.0 247200.0 ;
      RECT  102750.0 248550.0 103950.0 249750.0 ;
      RECT  104700.0 250800.0 105900.0 252000.0 ;
      RECT  121500.0 249900.0 120300.0 251100.0 ;
      RECT  120450.0 262950.0 121350.0 263850.0 ;
      RECT  122850.0 262950.0 123750.0 263850.0 ;
      RECT  120450.0 263400.0 121350.0 266550.0 ;
      RECT  120900.0 262950.0 123300.0 263850.0 ;
      RECT  122850.0 258750.0 123750.0 263400.0 ;
      RECT  120300.0 266550.0 121500.0 267750.0 ;
      RECT  122700.0 257550.0 123900.0 258750.0 ;
      RECT  123900.0 262800.0 122700.0 264000.0 ;
      RECT  102750.0 261450.0 103950.0 262650.0 ;
      RECT  104700.0 259200.0 105900.0 260400.0 ;
      RECT  121500.0 260100.0 120300.0 261300.0 ;
      RECT  120450.0 276450.0 121350.0 275550.0 ;
      RECT  122850.0 276450.0 123750.0 275550.0 ;
      RECT  120450.0 276000.0 121350.0 272850.0 ;
      RECT  120900.0 276450.0 123300.0 275550.0 ;
      RECT  122850.0 280650.0 123750.0 276000.0 ;
      RECT  120300.0 272850.0 121500.0 271650.0 ;
      RECT  122700.0 281850.0 123900.0 280650.0 ;
      RECT  123900.0 276600.0 122700.0 275400.0 ;
      RECT  102750.0 276750.0 103950.0 277950.0 ;
      RECT  104700.0 279000.0 105900.0 280200.0 ;
      RECT  121500.0 278100.0 120300.0 279300.0 ;
      RECT  120450.0 291150.0 121350.0 292050.0 ;
      RECT  122850.0 291150.0 123750.0 292050.0 ;
      RECT  120450.0 291600.0 121350.0 294750.0 ;
      RECT  120900.0 291150.0 123300.0 292050.0 ;
      RECT  122850.0 286950.0 123750.0 291600.0 ;
      RECT  120300.0 294750.0 121500.0 295950.0 ;
      RECT  122700.0 285750.0 123900.0 286950.0 ;
      RECT  123900.0 291000.0 122700.0 292200.0 ;
      RECT  102750.0 289650.0 103950.0 290850.0 ;
      RECT  104700.0 287400.0 105900.0 288600.0 ;
      RECT  121500.0 288300.0 120300.0 289500.0 ;
      RECT  120450.0 304650.0 121350.0 303750.0 ;
      RECT  122850.0 304650.0 123750.0 303750.0 ;
      RECT  120450.0 304200.0 121350.0 301050.0 ;
      RECT  120900.0 304650.0 123300.0 303750.0 ;
      RECT  122850.0 308850.0 123750.0 304200.0 ;
      RECT  120300.0 301050.0 121500.0 299850.0 ;
      RECT  122700.0 310050.0 123900.0 308850.0 ;
      RECT  123900.0 304800.0 122700.0 303600.0 ;
      RECT  102750.0 304950.0 103950.0 306150.0 ;
      RECT  104700.0 307200.0 105900.0 308400.0 ;
      RECT  121500.0 306300.0 120300.0 307500.0 ;
      RECT  120450.0 319350.0 121350.0 320250.0 ;
      RECT  122850.0 319350.0 123750.0 320250.0 ;
      RECT  120450.0 319800.0 121350.0 322950.0 ;
      RECT  120900.0 319350.0 123300.0 320250.0 ;
      RECT  122850.0 315150.0 123750.0 319800.0 ;
      RECT  120300.0 322950.0 121500.0 324150.0 ;
      RECT  122700.0 313950.0 123900.0 315150.0 ;
      RECT  123900.0 319200.0 122700.0 320400.0 ;
      RECT  102750.0 317850.0 103950.0 319050.0 ;
      RECT  104700.0 315600.0 105900.0 316800.0 ;
      RECT  121500.0 316500.0 120300.0 317700.0 ;
      RECT  120450.0 332850.0 121350.0 331950.0 ;
      RECT  122850.0 332850.0 123750.0 331950.0 ;
      RECT  120450.0 332400.0 121350.0 329250.0 ;
      RECT  120900.0 332850.0 123300.0 331950.0 ;
      RECT  122850.0 337050.0 123750.0 332400.0 ;
      RECT  120300.0 329250.0 121500.0 328050.0 ;
      RECT  122700.0 338250.0 123900.0 337050.0 ;
      RECT  123900.0 333000.0 122700.0 331800.0 ;
      RECT  102750.0 333150.0 103950.0 334350.0 ;
      RECT  104700.0 335400.0 105900.0 336600.0 ;
      RECT  121500.0 334500.0 120300.0 335700.0 ;
      RECT  120450.0 347550.0 121350.0 348450.0 ;
      RECT  122850.0 347550.0 123750.0 348450.0 ;
      RECT  120450.0 348000.0 121350.0 351150.0 ;
      RECT  120900.0 347550.0 123300.0 348450.0 ;
      RECT  122850.0 343350.0 123750.0 348000.0 ;
      RECT  120300.0 351150.0 121500.0 352350.0 ;
      RECT  122700.0 342150.0 123900.0 343350.0 ;
      RECT  123900.0 347400.0 122700.0 348600.0 ;
      RECT  102750.0 346050.0 103950.0 347250.0 ;
      RECT  104700.0 343800.0 105900.0 345000.0 ;
      RECT  121500.0 344700.0 120300.0 345900.0 ;
      RECT  120450.0 361050.0 121350.0 360150.0 ;
      RECT  122850.0 361050.0 123750.0 360150.0 ;
      RECT  120450.0 360600.0 121350.0 357450.0 ;
      RECT  120900.0 361050.0 123300.0 360150.0 ;
      RECT  122850.0 365250.0 123750.0 360600.0 ;
      RECT  120300.0 357450.0 121500.0 356250.0 ;
      RECT  122700.0 366450.0 123900.0 365250.0 ;
      RECT  123900.0 361200.0 122700.0 360000.0 ;
      RECT  102750.0 361350.0 103950.0 362550.0 ;
      RECT  104700.0 363600.0 105900.0 364800.0 ;
      RECT  121500.0 362700.0 120300.0 363900.0 ;
      RECT  120450.0 375750.0 121350.0 376650.0 ;
      RECT  122850.0 375750.0 123750.0 376650.0 ;
      RECT  120450.0 376200.0 121350.0 379350.0 ;
      RECT  120900.0 375750.0 123300.0 376650.0 ;
      RECT  122850.0 371550.0 123750.0 376200.0 ;
      RECT  120300.0 379350.0 121500.0 380550.0 ;
      RECT  122700.0 370350.0 123900.0 371550.0 ;
      RECT  123900.0 375600.0 122700.0 376800.0 ;
      RECT  102750.0 374250.0 103950.0 375450.0 ;
      RECT  104700.0 372000.0 105900.0 373200.0 ;
      RECT  121500.0 372900.0 120300.0 374100.0 ;
      RECT  120450.0 389250.0 121350.0 388350.0 ;
      RECT  122850.0 389250.0 123750.0 388350.0 ;
      RECT  120450.0 388800.0 121350.0 385650.0 ;
      RECT  120900.0 389250.0 123300.0 388350.0 ;
      RECT  122850.0 393450.0 123750.0 388800.0 ;
      RECT  120300.0 385650.0 121500.0 384450.0 ;
      RECT  122700.0 394650.0 123900.0 393450.0 ;
      RECT  123900.0 389400.0 122700.0 388200.0 ;
      RECT  102750.0 389550.0 103950.0 390750.0 ;
      RECT  104700.0 391800.0 105900.0 393000.0 ;
      RECT  121500.0 390900.0 120300.0 392100.0 ;
      RECT  120450.0 403950.0 121350.0 404850.0 ;
      RECT  122850.0 403950.0 123750.0 404850.0 ;
      RECT  120450.0 404400.0 121350.0 407550.0 ;
      RECT  120900.0 403950.0 123300.0 404850.0 ;
      RECT  122850.0 399750.0 123750.0 404400.0 ;
      RECT  120300.0 407550.0 121500.0 408750.0 ;
      RECT  122700.0 398550.0 123900.0 399750.0 ;
      RECT  123900.0 403800.0 122700.0 405000.0 ;
      RECT  102750.0 402450.0 103950.0 403650.0 ;
      RECT  104700.0 400200.0 105900.0 401400.0 ;
      RECT  121500.0 401100.0 120300.0 402300.0 ;
      RECT  120450.0 417450.0 121350.0 416550.0 ;
      RECT  122850.0 417450.0 123750.0 416550.0 ;
      RECT  120450.0 417000.0 121350.0 413850.0 ;
      RECT  120900.0 417450.0 123300.0 416550.0 ;
      RECT  122850.0 421650.0 123750.0 417000.0 ;
      RECT  120300.0 413850.0 121500.0 412650.0 ;
      RECT  122700.0 422850.0 123900.0 421650.0 ;
      RECT  123900.0 417600.0 122700.0 416400.0 ;
      RECT  102750.0 417750.0 103950.0 418950.0 ;
      RECT  104700.0 420000.0 105900.0 421200.0 ;
      RECT  121500.0 419100.0 120300.0 420300.0 ;
      RECT  102900.0 199200.0 103800.0 424800.0 ;
      RECT  59400.0 81000.0 119400.0 70800.0 ;
      RECT  59400.0 60600.0 119400.0 70800.0 ;
      RECT  59400.0 60600.0 119400.0 50400.0 ;
      RECT  59400.0 40200.0 119400.0 50400.0 ;
      RECT  59400.0 76500.0 60600.0 75300.0 ;
      RECT  59400.0 66300.0 60600.0 65100.0 ;
      RECT  59400.0 56100.0 60600.0 54900.0 ;
      RECT  59400.0 45900.0 60600.0 44700.0 ;
      RECT  118200.0 76500.0 119400.0 75300.0 ;
      RECT  114900.0 79200.0 119400.0 78000.0 ;
      RECT  118200.0 66300.0 119400.0 65100.0 ;
      RECT  114900.0 63600.0 119400.0 62400.0 ;
      RECT  118200.0 56100.0 119400.0 54900.0 ;
      RECT  114900.0 58800.0 119400.0 57600.0 ;
      RECT  118200.0 45900.0 119400.0 44700.0 ;
      RECT  114900.0 43200.0 119400.0 42000.0 ;
      RECT  59400.0 71400.0 119400.0 70200.0 ;
      RECT  59400.0 51000.0 119400.0 49800.0 ;
      RECT  176850.0 5850.0 178050.0 7050.0 ;
      RECT  187050.0 5850.0 188250.0 7050.0 ;
      RECT  180600.0 300.0 181800.0 1500.0 ;
      RECT  190800.0 300.0 192000.0 1500.0 ;
      RECT  148350.0 199800.0 149550.0 198600.0 ;
      RECT  148350.0 228000.0 149550.0 226800.0 ;
      RECT  148350.0 256200.0 149550.0 255000.0 ;
      RECT  148350.0 284400.0 149550.0 283200.0 ;
      RECT  148350.0 312600.0 149550.0 311400.0 ;
      RECT  148350.0 340800.0 149550.0 339600.0 ;
      RECT  148350.0 369000.0 149550.0 367800.0 ;
      RECT  148350.0 397200.0 149550.0 396000.0 ;
      RECT  148350.0 425400.0 149550.0 424200.0 ;
      RECT  130800.0 88650.0 129600.0 89850.0 ;
      RECT  135900.0 88500.0 134700.0 89700.0 ;
      RECT  127800.0 102750.0 126600.0 103950.0 ;
      RECT  138600.0 102600.0 137400.0 103800.0 ;
      RECT  130800.0 145050.0 129600.0 146250.0 ;
      RECT  141300.0 144900.0 140100.0 146100.0 ;
      RECT  127800.0 159150.0 126600.0 160350.0 ;
      RECT  144000.0 159000.0 142800.0 160200.0 ;
      RECT  132900.0 85800.0 131700.0 87000.0 ;
      RECT  132900.0 85800.0 131700.0 87000.0 ;
      RECT  147750.0 87000.0 148950.0 85800.0 ;
      RECT  132900.0 114000.0 131700.0 115200.0 ;
      RECT  132900.0 114000.0 131700.0 115200.0 ;
      RECT  147750.0 115200.0 148950.0 114000.0 ;
      RECT  132900.0 142200.0 131700.0 143400.0 ;
      RECT  132900.0 142200.0 131700.0 143400.0 ;
      RECT  147750.0 143400.0 148950.0 142200.0 ;
      RECT  132900.0 170400.0 131700.0 171600.0 ;
      RECT  132900.0 170400.0 131700.0 171600.0 ;
      RECT  147750.0 171600.0 148950.0 170400.0 ;
      RECT  120000.0 75300.0 118800.0 76500.0 ;
      RECT  135900.0 75300.0 134700.0 76500.0 ;
      RECT  120000.0 65100.0 118800.0 66300.0 ;
      RECT  138600.0 65100.0 137400.0 66300.0 ;
      RECT  120000.0 54900.0 118800.0 56100.0 ;
      RECT  141300.0 54900.0 140100.0 56100.0 ;
      RECT  120000.0 44700.0 118800.0 45900.0 ;
      RECT  144000.0 44700.0 142800.0 45900.0 ;
      RECT  120600.0 70200.0 119400.0 71400.0 ;
      RECT  149550.0 70350.0 148350.0 71550.0 ;
      RECT  120600.0 49800.0 119400.0 51000.0 ;
      RECT  149550.0 49950.0 148350.0 51150.0 ;
      RECT  164700.0 32250.0 163500.0 33450.0 ;
      RECT  159300.0 27750.0 158100.0 28950.0 ;
      RECT  162000.0 25350.0 160800.0 26550.0 ;
      RECT  164700.0 429450.0 163500.0 430650.0 ;
      RECT  167400.0 96750.0 166200.0 97950.0 ;
      RECT  170100.0 194850.0 168900.0 196050.0 ;
      RECT  156600.0 82500.0 155400.0 83700.0 ;
      RECT  103950.0 426300.0 102750.0 427500.0 ;
      RECT  156600.0 426300.0 155400.0 427500.0 ;
      RECT  152850.0 23400.0 151650.0 24600.0 ;
      RECT  152850.0 192900.0 151650.0 194100.0 ;
      RECT  152850.0 94800.0 151650.0 96000.0 ;
      RECT  180300.0 0.0 181200.0 1800.0 ;
      RECT  190500.0 0.0 191400.0 1800.0 ;
      RECT  169050.0 0.0 169950.0 444600.0 ;
      RECT  166350.0 0.0 167250.0 444600.0 ;
      RECT  158250.0 0.0 159150.0 444600.0 ;
      RECT  160950.0 0.0 161850.0 444600.0 ;
      RECT  163650.0 0.0 164550.0 444600.0 ;
      RECT  155550.0 0.0 156450.0 444600.0 ;
      RECT  148350.0 0.0 152850.0 444600.0 ;
      RECT  50100.0 289800.0 7.1054273576e-12 290700.0 ;
      RECT  50100.0 292500.0 7.1054273576e-12 293400.0 ;
      RECT  50100.0 295200.0 7.1054273576e-12 296100.0 ;
      RECT  50100.0 300600.0 7.1054273576e-12 301500.0 ;
      RECT  33750.0 205050.0 32850.0 284850.0 ;
      RECT  50100.0 287100.0 47400.0 288000.0 ;
      RECT  38700.0 297900.0 36000.0 298800.0 ;
      RECT  24600.0 287100.0 21900.0 288000.0 ;
      RECT  10500.0 297900.0 7800.0 298800.0 ;
      RECT  0.0 202200.0 10200.0 262200.0 ;
      RECT  20400.0 202200.0 10200.0 262200.0 ;
      RECT  20400.0 202200.0 30600.0 262200.0 ;
      RECT  4500.0 202200.0 5700.0 203400.0 ;
      RECT  14700.0 202200.0 15900.0 203400.0 ;
      RECT  24900.0 202200.0 26100.0 203400.0 ;
      RECT  4500.0 261000.0 5700.0 262200.0 ;
      RECT  1800.0 257700.0 3000.0 262200.0 ;
      RECT  14700.0 261000.0 15900.0 262200.0 ;
      RECT  17400.0 257700.0 18600.0 262200.0 ;
      RECT  24900.0 261000.0 26100.0 262200.0 ;
      RECT  22200.0 257700.0 23400.0 262200.0 ;
      RECT  9600.0 202200.0 10800.0 262200.0 ;
      RECT  30000.0 202200.0 31200.0 262200.0 ;
      RECT  46800.0 317850.0 38700.0 318750.0 ;
      RECT  41250.0 313050.0 40350.0 313950.0 ;
      RECT  41250.0 317850.0 40350.0 318750.0 ;
      RECT  40800.0 313050.0 38700.0 313950.0 ;
      RECT  41250.0 313500.0 40350.0 318300.0 ;
      RECT  46800.0 317850.0 40800.0 318750.0 ;
      RECT  38700.0 312900.0 37500.0 314100.0 ;
      RECT  38700.0 317700.0 37500.0 318900.0 ;
      RECT  48000.0 317700.0 46800.0 318900.0 ;
      RECT  41400.0 317700.0 40200.0 318900.0 ;
      RECT  28500.0 315450.0 29400.0 316350.0 ;
      RECT  28950.0 315450.0 32250.0 316350.0 ;
      RECT  28500.0 315900.0 29400.0 316800.0 ;
      RECT  23400.0 315450.0 24300.0 316350.0 ;
      RECT  23400.0 314100.0 24300.0 315900.0 ;
      RECT  23850.0 315450.0 28950.0 316350.0 ;
      RECT  32250.0 315300.0 33450.0 316500.0 ;
      RECT  23250.0 314100.0 24450.0 312900.0 ;
      RECT  28350.0 317400.0 29550.0 316200.0 ;
      RECT  29250.0 330150.0 30150.0 331050.0 ;
      RECT  29250.0 332550.0 30150.0 333450.0 ;
      RECT  29700.0 330150.0 32850.0 331050.0 ;
      RECT  29250.0 330600.0 30150.0 333000.0 ;
      RECT  25050.0 332550.0 29700.0 333450.0 ;
      RECT  32850.0 330000.0 34050.0 331200.0 ;
      RECT  23850.0 332400.0 25050.0 333600.0 ;
      RECT  29100.0 333600.0 30300.0 332400.0 ;
      RECT  18600.0 327450.0 10500.0 328350.0 ;
      RECT  13050.0 322650.0 12150.0 323550.0 ;
      RECT  13050.0 327450.0 12150.0 328350.0 ;
      RECT  12600.0 322650.0 10500.0 323550.0 ;
      RECT  13050.0 323100.0 12150.0 327900.0 ;
      RECT  18600.0 327450.0 12600.0 328350.0 ;
      RECT  10500.0 322500.0 9300.0 323700.0 ;
      RECT  10500.0 327300.0 9300.0 328500.0 ;
      RECT  19800.0 327300.0 18600.0 328500.0 ;
      RECT  13200.0 327300.0 12000.0 328500.0 ;
      RECT  3000.0 262800.0 1800.0 261600.0 ;
      RECT  3000.0 301650.0 1800.0 300450.0 ;
      RECT  5700.0 262800.0 4500.0 261600.0 ;
      RECT  5700.0 290850.0 4500.0 289650.0 ;
      RECT  18600.0 262800.0 17400.0 261600.0 ;
      RECT  18600.0 293550.0 17400.0 292350.0 ;
      RECT  23400.0 262800.0 22200.0 261600.0 ;
      RECT  23400.0 296250.0 22200.0 295050.0 ;
      RECT  10800.0 262800.0 9600.0 261600.0 ;
      RECT  10800.0 288150.0 9600.0 286950.0 ;
      RECT  31200.0 262800.0 30000.0 261600.0 ;
      RECT  31200.0 288150.0 30000.0 286950.0 ;
      RECT  22350.0 371700.0 21450.0 426900.0 ;
      RECT  22350.0 381300.0 21450.0 384000.0 ;
      RECT  22350.0 384000.0 21450.0 426900.0 ;
      RECT  6750.0 424200.0 5850.0 426900.0 ;
      RECT  20100.0 376500.0 19200.0 384000.0 ;
      RECT  13350.0 376500.0 12450.0 381300.0 ;
      RECT  43200.0 415500.0 44100.0 422700.0 ;
      RECT  35550.0 424650.0 36450.0 425550.0 ;
      RECT  35550.0 425850.0 36450.0 426750.0 ;
      RECT  36000.0 424650.0 43650.0 425550.0 ;
      RECT  35550.0 425100.0 36450.0 426300.0 ;
      RECT  28350.0 425850.0 36000.0 426750.0 ;
      RECT  27900.0 416700.0 28800.0 423900.0 ;
      RECT  43050.0 422100.0 44250.0 423300.0 ;
      RECT  27750.0 425700.0 28950.0 426900.0 ;
      RECT  27750.0 416100.0 28950.0 417300.0 ;
      RECT  43050.0 414900.0 44250.0 416100.0 ;
      RECT  43050.0 424500.0 44250.0 425700.0 ;
      RECT  27750.0 423300.0 28950.0 424500.0 ;
      RECT  16500.0 396000.0 6300.0 381300.0 ;
      RECT  16500.0 396000.0 6300.0 410100.0 ;
      RECT  16500.0 424200.0 6300.0 410100.0 ;
      RECT  13500.0 396000.0 12300.0 424200.0 ;
      RECT  10500.0 396000.0 9300.0 424200.0 ;
      RECT  6900.0 396000.0 5700.0 424200.0 ;
      RECT  22350.0 398100.0 21150.0 399300.0 ;
      RECT  22350.0 420900.0 21150.0 422100.0 ;
      RECT  22350.0 410100.0 21150.0 411300.0 ;
      RECT  22350.0 370500.0 21150.0 371700.0 ;
      RECT  21300.0 426300.0 22500.0 427500.0 ;
      RECT  5700.0 426300.0 6900.0 427500.0 ;
      RECT  19050.0 383400.0 20250.0 384600.0 ;
      RECT  19050.0 375900.0 20250.0 377100.0 ;
      RECT  12300.0 375900.0 13500.0 377100.0 ;
      RECT  44550.0 285450.0 43350.0 284250.0 ;
      RECT  44550.0 244650.0 43350.0 243450.0 ;
      RECT  44550.0 304350.0 43350.0 303150.0 ;
      RECT  44550.0 244650.0 43350.0 243450.0 ;
      RECT  33900.0 205650.0 32700.0 204450.0 ;
      RECT  29550.0 285450.0 28350.0 284250.0 ;
      RECT  26850.0 290850.0 25650.0 289650.0 ;
      RECT  30300.0 328200.0 29100.0 327000.0 ;
      RECT  30300.0 328200.0 29100.0 327000.0 ;
      RECT  30300.0 304350.0 29100.0 303150.0 ;
      RECT  27600.0 331200.0 26400.0 330000.0 ;
      RECT  27600.0 331200.0 26400.0 330000.0 ;
      RECT  27600.0 301650.0 26400.0 300450.0 ;
      RECT  41400.0 304350.0 40200.0 303150.0 ;
      RECT  43350.0 301650.0 42150.0 300450.0 ;
      RECT  45300.0 293550.0 44100.0 292350.0 ;
      RECT  13200.0 304350.0 12000.0 303150.0 ;
      RECT  15150.0 293550.0 13950.0 292350.0 ;
      RECT  17100.0 296250.0 15900.0 295050.0 ;
      RECT  29550.0 322500.0 28350.0 323700.0 ;
      RECT  30300.0 339600.0 29100.0 340800.0 ;
      RECT  16050.0 362100.0 14850.0 363300.0 ;
      RECT  28950.0 342300.0 27750.0 343500.0 ;
      RECT  50700.0 288150.0 49500.0 286950.0 ;
      RECT  36600.0 298950.0 35400.0 297750.0 ;
      RECT  22500.0 288150.0 21300.0 286950.0 ;
      RECT  8400.0 298950.0 7200.0 297750.0 ;
      RECT  50100.0 342450.0 28350.0 343350.0 ;
      RECT  50100.0 362250.0 15450.0 363150.0 ;
      RECT  50100.0 322650.0 28950.0 323550.0 ;
      RECT  50100.0 339750.0 29700.0 340650.0 ;
      RECT  50100.0 303300.0 7.1054273576e-12 304200.0 ;
      RECT  50100.0 284400.0 7.1054273576e-12 285300.0 ;
      RECT  50100.0 297900.0 7.1054273576e-12 298800.0 ;
      RECT  50100.0 287100.0 7.1054273576e-12 288000.0 ;
      RECT  170100.0 342300.0 168900.0 343500.0 ;
      RECT  49800.0 342450.0 48600.0 343650.0 ;
      RECT  167400.0 362100.0 166200.0 363300.0 ;
      RECT  49800.0 362250.0 48600.0 363450.0 ;
      RECT  162000.0 322500.0 160800.0 323700.0 ;
      RECT  49800.0 322650.0 48600.0 323850.0 ;
      RECT  159300.0 339600.0 158100.0 340800.0 ;
      RECT  49800.0 339750.0 48600.0 340950.0 ;
      RECT  164700.0 303150.0 163500.0 304350.0 ;
      RECT  49800.0 303300.0 48600.0 304500.0 ;
      RECT  156600.0 284250.0 155400.0 285450.0 ;
      RECT  49800.0 284400.0 48600.0 285600.0 ;
      RECT  55950.0 297750.0 54750.0 298950.0 ;
      RECT  151200.0 286950.0 150000.0 288150.0 ;
      RECT  49800.0 287100.0 48600.0 288300.0 ;
   LAYER  metal3 ;
      RECT  50100.0 342150.0 169500.0 343650.0 ;
      RECT  50100.0 361950.0 166800.0 363450.0 ;
      RECT  50100.0 322350.0 161400.0 323850.0 ;
      RECT  50100.0 339450.0 158700.0 340950.0 ;
      RECT  50100.0 303000.0 164100.0 304500.0 ;
      RECT  50100.0 284100.0 156000.0 285600.0 ;
      RECT  50100.0 286800.0 150600.0 288300.0 ;
      RECT  176550.0 6300.0 178050.0 151200.0 ;
      RECT  186750.0 6300.0 188250.0 151200.0 ;
      RECT  180300.0 0.0 181800.0 30000.0 ;
      RECT  190500.0 0.0 192000.0 30000.0 ;
      RECT  132300.0 85650.0 148350.0 87150.0 ;
      RECT  132300.0 113850.0 148350.0 115350.0 ;
      RECT  132300.0 142050.0 148350.0 143550.0 ;
      RECT  132300.0 170250.0 148350.0 171750.0 ;
      RECT  176400.0 151200.0 178200.0 153000.0 ;
      RECT  186600.0 151200.0 188400.0 153000.0 ;
      RECT  180000.0 30900.0 181800.0 32700.0 ;
      RECT  190200.0 30900.0 192000.0 32700.0 ;
      RECT  60300.0 76800.0 62100.0 75000.0 ;
      RECT  60300.0 66600.0 62100.0 64800.0 ;
      RECT  60300.0 56400.0 62100.0 54600.0 ;
      RECT  60300.0 46200.0 62100.0 44400.0 ;
      RECT  176550.0 5550.0 178350.0 7350.0 ;
      RECT  186750.0 5550.0 188550.0 7350.0 ;
      RECT  180300.0 0.0 182100.0 1800.0 ;
      RECT  190500.0 0.0 192300.0 1800.0 ;
      RECT  133200.0 85500.0 131400.0 87300.0 ;
      RECT  147450.0 87300.0 149250.0 85500.0 ;
      RECT  133200.0 113700.0 131400.0 115500.0 ;
      RECT  147450.0 115500.0 149250.0 113700.0 ;
      RECT  133200.0 141900.0 131400.0 143700.0 ;
      RECT  147450.0 143700.0 149250.0 141900.0 ;
      RECT  133200.0 170100.0 131400.0 171900.0 ;
      RECT  147450.0 171900.0 149250.0 170100.0 ;
      RECT  53100.0 75000.0 60300.0 76500.0 ;
      RECT  53100.0 64800.0 60300.0 66300.0 ;
      RECT  53100.0 54600.0 60300.0 56100.0 ;
      RECT  53100.0 44400.0 60300.0 45900.0 ;
      RECT  3150.0 262200.0 1650.0 301050.0 ;
      RECT  5850.0 262200.0 4350.0 290250.0 ;
      RECT  18750.0 262200.0 17250.0 292950.0 ;
      RECT  23550.0 262200.0 22050.0 295650.0 ;
      RECT  10950.0 262200.0 9450.0 287550.0 ;
      RECT  31350.0 262200.0 29850.0 287550.0 ;
      RECT  44700.0 244050.0 43200.0 303750.0 ;
      RECT  30450.0 303750.0 28950.0 327600.0 ;
      RECT  27750.0 301050.0 26250.0 330600.0 ;
      RECT  4200.0 203100.0 6000.0 204900.0 ;
      RECT  14400.0 203100.0 16200.0 204900.0 ;
      RECT  24600.0 203100.0 26400.0 204900.0 ;
      RECT  3300.0 263100.0 1500.0 261300.0 ;
      RECT  3300.0 301950.0 1500.0 300150.0 ;
      RECT  6000.0 263100.0 4200.0 261300.0 ;
      RECT  6000.0 291150.0 4200.0 289350.0 ;
      RECT  18900.0 263100.0 17100.0 261300.0 ;
      RECT  18900.0 293850.0 17100.0 292050.0 ;
      RECT  23700.0 263100.0 21900.0 261300.0 ;
      RECT  23700.0 296550.0 21900.0 294750.0 ;
      RECT  11100.0 263100.0 9300.0 261300.0 ;
      RECT  11100.0 288450.0 9300.0 286650.0 ;
      RECT  31500.0 263100.0 29700.0 261300.0 ;
      RECT  31500.0 288450.0 29700.0 286650.0 ;
      RECT  44850.0 244950.0 43050.0 243150.0 ;
      RECT  44850.0 304650.0 43050.0 302850.0 ;
      RECT  30600.0 328500.0 28800.0 326700.0 ;
      RECT  30600.0 304650.0 28800.0 302850.0 ;
      RECT  27900.0 331500.0 26100.0 329700.0 ;
      RECT  27900.0 301950.0 26100.0 300150.0 ;
      RECT  16200.0 203100.0 14400.0 204900.0 ;
      RECT  26400.0 203100.0 24600.0 204900.0 ;
      RECT  6000.0 203100.0 4200.0 204900.0 ;
      RECT  170400.0 342000.0 168600.0 343800.0 ;
      RECT  50100.0 342150.0 48300.0 343950.0 ;
      RECT  167700.0 361800.0 165900.0 363600.0 ;
      RECT  50100.0 361950.0 48300.0 363750.0 ;
      RECT  162300.0 322200.0 160500.0 324000.0 ;
      RECT  50100.0 322350.0 48300.0 324150.0 ;
      RECT  159600.0 339300.0 157800.0 341100.0 ;
      RECT  50100.0 339450.0 48300.0 341250.0 ;
      RECT  165000.0 302850.0 163200.0 304650.0 ;
      RECT  50100.0 303000.0 48300.0 304800.0 ;
      RECT  156900.0 283950.0 155100.0 285750.0 ;
      RECT  50100.0 284100.0 48300.0 285900.0 ;
      RECT  151500.0 286650.0 149700.0 288450.0 ;
      RECT  50100.0 286800.0 48300.0 288600.0 ;
   END
   END    sram_2_16_1_scn3me_subm
END    LIBRARY
