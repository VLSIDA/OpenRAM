MACRO sram_2_16_1_scn3me_subm
    CLASS RING ;
    ORIGIN 66.9 0.0 ;
    FOREIGN  sram 0.0 0.0 ;
    SIZE 222.3 BY 459.3 ;
    SYMMETRY X Y R90 ;
    PIN vdd 
        DIRECTION INOUT ; 
        USE POWER ; 
        SHAPE ABUTMENT ; 
        PORT             
        Layer metal1 ; 
        RECT  0.45 0.0 9.45 459.3 ;
        RECT  147.45 0.0 156.45 459.3 ;
        END             
    END vdd 
    PIN gnd 
        DIRECTION INOUT ; 
        USE GROUND ; 
        SHAPE ABUTMENT ; 
        PORT             
        Layer metal2 ; 
        RECT  95.55 0.0 104.55 459.3 ;
        END             
    END gnd 
    PIN DATA[0] 
        DIRECTION INOUT ; 
        PORT             
        Layer metal3 ; 
        RECT  128.7 0.0 130.2 30.15 ;
        RECT  128.7 0.0 130.5 1.8 ;
        END             
    END DATA[0] 
    PIN DATA[1] 
        DIRECTION INOUT ; 
        PORT             
        Layer metal3 ; 
        RECT  138.9 0.0 140.4 30.15 ;
        RECT  138.9 0.0 140.7 1.8 ;
        END             
    END DATA[1] 
    PIN ADDR[0] 
        DIRECTION INPUT ; 
        PORT             
        Layer metal3 ; 
        RECT  0.45 73.95 17.55 75.45 ;
        END             
    END ADDR[0] 
    PIN ADDR[1] 
        DIRECTION INPUT ; 
        PORT             
        Layer metal3 ; 
        RECT  0.45 63.75 17.55 65.25 ;
        END             
    END ADDR[1] 
    PIN ADDR[2] 
        DIRECTION INPUT ; 
        PORT             
        Layer metal3 ; 
        RECT  0.45 53.55 17.55 55.05 ;
        END             
    END ADDR[2] 
    PIN ADDR[3] 
        DIRECTION INPUT ; 
        PORT             
        Layer metal3 ; 
        RECT  0.45 43.35 17.55 44.85 ;
        END             
    END ADDR[3] 
    PIN CSb 
        DIRECTION INPUT ; 
        PORT             
        Layer metal3 ; 
        RECT  -62.1 86.4 -60.3 88.2 ;
        END             
    END CSb 
    PIN OEb 
        DIRECTION INPUT ; 
        PORT             
        Layer metal3 ; 
        RECT  -41.7 86.4 -39.9 88.2 ;
        END             
    END OEb 
    PIN WEb 
        DIRECTION INPUT ; 
        PORT             
        Layer metal3 ; 
        RECT  -51.9 86.4 -50.1 88.2 ;
        END             
    END WEb 
    PIN clk 
        DIRECTION INPUT ; 
        PORT             
        Layer metal3 ; 
        RECT  -27.15 85.5 106.35 87.0 ;
        RECT  -27.6 85.5 -25.8 87.3 ;
        END             
    END clk 
    OBS 
        Layer  metal1 ; 
        RECT  -10.2 293.55 0.45 294.45 ;
        RECT  147.45 0.0 156.45 459.3 ;
        RECT  0.45 0.0 9.45 459.3 ;
        RECT  51.45 206.4 52.35 209.7 ;
        RECT  88.95 202.35 89.85 203.25 ;
        RECT  89.4 202.35 124.8 203.25 ;
        RECT  88.95 202.8 89.85 208.2 ;
        RECT  51.45 219.9 52.35 223.2 ;
        RECT  88.95 226.35 89.85 227.25 ;
        RECT  89.4 226.35 124.8 227.25 ;
        RECT  88.95 221.4 89.85 226.8 ;
        RECT  51.45 235.8 52.35 239.1 ;
        RECT  88.95 231.75 89.85 232.65 ;
        RECT  89.4 231.75 124.8 232.65 ;
        RECT  88.95 232.2 89.85 237.6 ;
        RECT  51.45 249.3 52.35 252.6 ;
        RECT  88.95 255.75 89.85 256.65 ;
        RECT  89.4 255.75 124.8 256.65 ;
        RECT  88.95 250.8 89.85 256.2 ;
        RECT  51.45 265.2 52.35 268.5 ;
        RECT  88.95 261.15 89.85 262.05 ;
        RECT  89.4 261.15 124.8 262.05 ;
        RECT  88.95 261.6 89.85 267.0 ;
        RECT  51.45 278.7 52.35 282.0 ;
        RECT  88.95 285.15 89.85 286.05 ;
        RECT  89.4 285.15 124.8 286.05 ;
        RECT  88.95 280.2 89.85 285.6 ;
        RECT  51.45 294.6 52.35 297.9 ;
        RECT  88.95 290.55 89.85 291.45 ;
        RECT  89.4 290.55 124.8 291.45 ;
        RECT  88.95 291.0 89.85 296.4 ;
        RECT  51.45 308.1 52.35 311.4 ;
        RECT  88.95 314.55 89.85 315.45 ;
        RECT  89.4 314.55 124.8 315.45 ;
        RECT  88.95 309.6 89.85 315.0 ;
        RECT  51.45 324.0 52.35 327.3 ;
        RECT  88.95 319.95 89.85 320.85 ;
        RECT  89.4 319.95 124.8 320.85 ;
        RECT  88.95 320.4 89.85 325.8 ;
        RECT  51.45 337.5 52.35 340.8 ;
        RECT  88.95 343.95 89.85 344.85 ;
        RECT  89.4 343.95 124.8 344.85 ;
        RECT  88.95 339.0 89.85 344.4 ;
        RECT  51.45 353.4 52.35 356.7 ;
        RECT  88.95 349.35 89.85 350.25 ;
        RECT  89.4 349.35 124.8 350.25 ;
        RECT  88.95 349.8 89.85 355.2 ;
        RECT  51.45 366.9 52.35 370.2 ;
        RECT  88.95 373.35 89.85 374.25 ;
        RECT  89.4 373.35 124.8 374.25 ;
        RECT  88.95 368.4 89.85 373.8 ;
        RECT  51.45 382.8 52.35 386.1 ;
        RECT  88.95 378.75 89.85 379.65 ;
        RECT  89.4 378.75 124.8 379.65 ;
        RECT  88.95 379.2 89.85 384.6 ;
        RECT  51.45 396.3 52.35 399.6 ;
        RECT  88.95 402.75 89.85 403.65 ;
        RECT  89.4 402.75 124.8 403.65 ;
        RECT  88.95 397.8 89.85 403.2 ;
        RECT  51.45 412.2 52.35 415.5 ;
        RECT  88.95 408.15 89.85 409.05 ;
        RECT  89.4 408.15 124.8 409.05 ;
        RECT  88.95 408.6 89.85 414.0 ;
        RECT  51.45 425.7 52.35 429.0 ;
        RECT  88.95 432.15 89.85 433.05 ;
        RECT  89.4 432.15 124.8 433.05 ;
        RECT  88.95 427.2 89.85 432.6 ;
        RECT  88.95 214.35 124.35 215.25 ;
        RECT  88.95 243.75 124.35 244.65 ;
        RECT  88.95 273.15 124.35 274.05 ;
        RECT  88.95 302.55 124.35 303.45 ;
        RECT  88.95 331.95 124.35 332.85 ;
        RECT  88.95 361.35 124.35 362.25 ;
        RECT  88.95 390.75 124.35 391.65 ;
        RECT  88.95 420.15 124.35 421.05 ;
        RECT  74.85 88.8 91.95 89.7 ;
        RECT  74.85 104.7 89.25 105.6 ;
        RECT  74.85 147.6 86.55 148.5 ;
        RECT  74.85 163.5 83.85 164.4 ;
        RECT  114.45 33.3 129.45 34.2 ;
        RECT  109.05 28.65 129.75 29.55 ;
        RECT  111.75 26.25 129.75 27.15 ;
        RECT  114.45 446.4 124.35 447.3 ;
        RECT  117.15 97.95 124.35 98.85 ;
        RECT  119.85 196.05 124.35 196.95 ;
        RECT  54.15 456.6 55.05 457.5 ;
        RECT  54.15 435.3 55.05 457.05 ;
        RECT  54.6 456.6 107.25 457.5 ;
        RECT  124.35 213.75 147.45 214.65 ;
        RECT  124.35 243.15 147.45 244.05 ;
        RECT  124.35 272.55 147.45 273.45 ;
        RECT  124.35 301.95 147.45 302.85 ;
        RECT  124.35 331.35 147.45 332.25 ;
        RECT  124.35 360.75 147.45 361.65 ;
        RECT  124.35 390.15 147.45 391.05 ;
        RECT  124.35 419.55 147.45 420.45 ;
        RECT  124.35 458.4 147.45 459.3 ;
        RECT  124.35 168.75 147.45 169.65 ;
        RECT  124.35 100.05 147.45 100.95 ;
        RECT  124.35 87.3 147.45 88.2 ;
        RECT  129.75 10.35 147.45 11.25 ;
        RECT  139.35 10.35 147.45 11.25 ;
        RECT  0.45 214.35 29.85 215.25 ;
        RECT  0.45 243.75 29.85 244.65 ;
        RECT  0.45 273.15 29.85 274.05 ;
        RECT  0.45 302.55 29.85 303.45 ;
        RECT  0.45 331.95 29.85 332.85 ;
        RECT  0.45 361.35 29.85 362.25 ;
        RECT  0.45 390.75 29.85 391.65 ;
        RECT  0.45 420.15 29.85 421.05 ;
        RECT  0.45 126.15 29.85 127.05 ;
        RECT  0.45 184.95 29.85 185.85 ;
        RECT  0.0 36.3 0.9 37.2 ;
        RECT  72.15 36.3 73.05 37.2 ;
        RECT  0.0 36.3 0.9 36.75 ;
        RECT  0.45 36.3 72.6 37.2 ;
        RECT  72.15 36.75 73.05 39.0 ;
        RECT  95.55 437.1 144.75 438.0 ;
        RECT  102.15 8.1 144.75 9.0 ;
        RECT  29.85 140.85 95.55 141.75 ;
        RECT  29.85 199.65 95.55 200.55 ;
        RECT  75.75 69.15 95.55 70.05 ;
        RECT  75.75 69.15 95.55 70.05 ;
        RECT  75.75 48.75 95.55 49.65 ;
        RECT  75.75 48.75 95.55 49.65 ;
        RECT  123.75 213.6 135.15 214.8 ;
        RECT  124.95 211.5 126.15 213.6 ;
        RECT  127.95 211.5 129.15 212.7 ;
        RECT  130.95 211.5 132.15 212.7 ;
        RECT  133.95 211.5 135.15 213.6 ;
        RECT  127.65 210.6 128.85 211.5 ;
        RECT  124.95 204.9 126.15 210.6 ;
        RECT  127.65 209.4 130.05 210.6 ;
        RECT  127.65 206.1 128.85 209.4 ;
        RECT  131.25 207.9 132.45 211.5 ;
        RECT  130.65 206.7 132.45 207.9 ;
        RECT  131.25 206.1 132.45 206.7 ;
        RECT  127.35 204.9 128.55 206.1 ;
        RECT  131.55 204.9 132.75 206.1 ;
        RECT  133.95 204.9 135.15 210.6 ;
        RECT  129.45 203.4 130.65 203.7 ;
        RECT  123.75 202.2 135.15 203.4 ;
        RECT  125.85 200.1 128.55 201.3 ;
        RECT  130.05 200.1 132.75 201.3 ;
        RECT  123.75 214.8 135.15 216.0 ;
        RECT  124.95 216.0 126.15 218.1 ;
        RECT  127.95 216.9 129.15 218.1 ;
        RECT  130.95 216.9 132.15 218.1 ;
        RECT  133.95 216.0 135.15 218.1 ;
        RECT  127.65 218.1 128.85 219.0 ;
        RECT  124.95 219.0 126.15 224.7 ;
        RECT  127.65 219.0 130.05 220.2 ;
        RECT  127.65 220.2 128.85 223.5 ;
        RECT  131.25 218.1 132.45 221.7 ;
        RECT  130.65 221.7 132.45 222.9 ;
        RECT  131.25 222.9 132.45 223.5 ;
        RECT  127.35 223.5 128.55 224.7 ;
        RECT  131.55 223.5 132.75 224.7 ;
        RECT  133.95 219.0 135.15 224.7 ;
        RECT  129.45 225.9 130.65 226.2 ;
        RECT  123.75 226.2 135.15 227.4 ;
        RECT  125.85 228.3 128.55 229.5 ;
        RECT  130.05 228.3 132.75 229.5 ;
        RECT  123.75 243.0 135.15 244.2 ;
        RECT  124.95 240.9 126.15 243.0 ;
        RECT  127.95 240.9 129.15 242.1 ;
        RECT  130.95 240.9 132.15 242.1 ;
        RECT  133.95 240.9 135.15 243.0 ;
        RECT  127.65 240.0 128.85 240.9 ;
        RECT  124.95 234.3 126.15 240.0 ;
        RECT  127.65 238.8 130.05 240.0 ;
        RECT  127.65 235.5 128.85 238.8 ;
        RECT  131.25 237.3 132.45 240.9 ;
        RECT  130.65 236.1 132.45 237.3 ;
        RECT  131.25 235.5 132.45 236.1 ;
        RECT  127.35 234.3 128.55 235.5 ;
        RECT  131.55 234.3 132.75 235.5 ;
        RECT  133.95 234.3 135.15 240.0 ;
        RECT  129.45 232.8 130.65 233.1 ;
        RECT  123.75 231.6 135.15 232.8 ;
        RECT  125.85 229.5 128.55 230.7 ;
        RECT  130.05 229.5 132.75 230.7 ;
        RECT  123.75 244.2 135.15 245.4 ;
        RECT  124.95 245.4 126.15 247.5 ;
        RECT  127.95 246.3 129.15 247.5 ;
        RECT  130.95 246.3 132.15 247.5 ;
        RECT  133.95 245.4 135.15 247.5 ;
        RECT  127.65 247.5 128.85 248.4 ;
        RECT  124.95 248.4 126.15 254.1 ;
        RECT  127.65 248.4 130.05 249.6 ;
        RECT  127.65 249.6 128.85 252.9 ;
        RECT  131.25 247.5 132.45 251.1 ;
        RECT  130.65 251.1 132.45 252.3 ;
        RECT  131.25 252.3 132.45 252.9 ;
        RECT  127.35 252.9 128.55 254.1 ;
        RECT  131.55 252.9 132.75 254.1 ;
        RECT  133.95 248.4 135.15 254.1 ;
        RECT  129.45 255.3 130.65 255.6 ;
        RECT  123.75 255.6 135.15 256.8 ;
        RECT  125.85 257.7 128.55 258.9 ;
        RECT  130.05 257.7 132.75 258.9 ;
        RECT  123.75 272.4 135.15 273.6 ;
        RECT  124.95 270.3 126.15 272.4 ;
        RECT  127.95 270.3 129.15 271.5 ;
        RECT  130.95 270.3 132.15 271.5 ;
        RECT  133.95 270.3 135.15 272.4 ;
        RECT  127.65 269.4 128.85 270.3 ;
        RECT  124.95 263.7 126.15 269.4 ;
        RECT  127.65 268.2 130.05 269.4 ;
        RECT  127.65 264.9 128.85 268.2 ;
        RECT  131.25 266.7 132.45 270.3 ;
        RECT  130.65 265.5 132.45 266.7 ;
        RECT  131.25 264.9 132.45 265.5 ;
        RECT  127.35 263.7 128.55 264.9 ;
        RECT  131.55 263.7 132.75 264.9 ;
        RECT  133.95 263.7 135.15 269.4 ;
        RECT  129.45 262.2 130.65 262.5 ;
        RECT  123.75 261.0 135.15 262.2 ;
        RECT  125.85 258.9 128.55 260.1 ;
        RECT  130.05 258.9 132.75 260.1 ;
        RECT  123.75 273.6 135.15 274.8 ;
        RECT  124.95 274.8 126.15 276.9 ;
        RECT  127.95 275.7 129.15 276.9 ;
        RECT  130.95 275.7 132.15 276.9 ;
        RECT  133.95 274.8 135.15 276.9 ;
        RECT  127.65 276.9 128.85 277.8 ;
        RECT  124.95 277.8 126.15 283.5 ;
        RECT  127.65 277.8 130.05 279.0 ;
        RECT  127.65 279.0 128.85 282.3 ;
        RECT  131.25 276.9 132.45 280.5 ;
        RECT  130.65 280.5 132.45 281.7 ;
        RECT  131.25 281.7 132.45 282.3 ;
        RECT  127.35 282.3 128.55 283.5 ;
        RECT  131.55 282.3 132.75 283.5 ;
        RECT  133.95 277.8 135.15 283.5 ;
        RECT  129.45 284.7 130.65 285.0 ;
        RECT  123.75 285.0 135.15 286.2 ;
        RECT  125.85 287.1 128.55 288.3 ;
        RECT  130.05 287.1 132.75 288.3 ;
        RECT  123.75 301.8 135.15 303.0 ;
        RECT  124.95 299.7 126.15 301.8 ;
        RECT  127.95 299.7 129.15 300.9 ;
        RECT  130.95 299.7 132.15 300.9 ;
        RECT  133.95 299.7 135.15 301.8 ;
        RECT  127.65 298.8 128.85 299.7 ;
        RECT  124.95 293.1 126.15 298.8 ;
        RECT  127.65 297.6 130.05 298.8 ;
        RECT  127.65 294.3 128.85 297.6 ;
        RECT  131.25 296.1 132.45 299.7 ;
        RECT  130.65 294.9 132.45 296.1 ;
        RECT  131.25 294.3 132.45 294.9 ;
        RECT  127.35 293.1 128.55 294.3 ;
        RECT  131.55 293.1 132.75 294.3 ;
        RECT  133.95 293.1 135.15 298.8 ;
        RECT  129.45 291.6 130.65 291.9 ;
        RECT  123.75 290.4 135.15 291.6 ;
        RECT  125.85 288.3 128.55 289.5 ;
        RECT  130.05 288.3 132.75 289.5 ;
        RECT  123.75 303.0 135.15 304.2 ;
        RECT  124.95 304.2 126.15 306.3 ;
        RECT  127.95 305.1 129.15 306.3 ;
        RECT  130.95 305.1 132.15 306.3 ;
        RECT  133.95 304.2 135.15 306.3 ;
        RECT  127.65 306.3 128.85 307.2 ;
        RECT  124.95 307.2 126.15 312.9 ;
        RECT  127.65 307.2 130.05 308.4 ;
        RECT  127.65 308.4 128.85 311.7 ;
        RECT  131.25 306.3 132.45 309.9 ;
        RECT  130.65 309.9 132.45 311.1 ;
        RECT  131.25 311.1 132.45 311.7 ;
        RECT  127.35 311.7 128.55 312.9 ;
        RECT  131.55 311.7 132.75 312.9 ;
        RECT  133.95 307.2 135.15 312.9 ;
        RECT  129.45 314.1 130.65 314.4 ;
        RECT  123.75 314.4 135.15 315.6 ;
        RECT  125.85 316.5 128.55 317.7 ;
        RECT  130.05 316.5 132.75 317.7 ;
        RECT  123.75 331.2 135.15 332.4 ;
        RECT  124.95 329.1 126.15 331.2 ;
        RECT  127.95 329.1 129.15 330.3 ;
        RECT  130.95 329.1 132.15 330.3 ;
        RECT  133.95 329.1 135.15 331.2 ;
        RECT  127.65 328.2 128.85 329.1 ;
        RECT  124.95 322.5 126.15 328.2 ;
        RECT  127.65 327.0 130.05 328.2 ;
        RECT  127.65 323.7 128.85 327.0 ;
        RECT  131.25 325.5 132.45 329.1 ;
        RECT  130.65 324.3 132.45 325.5 ;
        RECT  131.25 323.7 132.45 324.3 ;
        RECT  127.35 322.5 128.55 323.7 ;
        RECT  131.55 322.5 132.75 323.7 ;
        RECT  133.95 322.5 135.15 328.2 ;
        RECT  129.45 321.0 130.65 321.3 ;
        RECT  123.75 319.8 135.15 321.0 ;
        RECT  125.85 317.7 128.55 318.9 ;
        RECT  130.05 317.7 132.75 318.9 ;
        RECT  123.75 332.4 135.15 333.6 ;
        RECT  124.95 333.6 126.15 335.7 ;
        RECT  127.95 334.5 129.15 335.7 ;
        RECT  130.95 334.5 132.15 335.7 ;
        RECT  133.95 333.6 135.15 335.7 ;
        RECT  127.65 335.7 128.85 336.6 ;
        RECT  124.95 336.6 126.15 342.3 ;
        RECT  127.65 336.6 130.05 337.8 ;
        RECT  127.65 337.8 128.85 341.1 ;
        RECT  131.25 335.7 132.45 339.3 ;
        RECT  130.65 339.3 132.45 340.5 ;
        RECT  131.25 340.5 132.45 341.1 ;
        RECT  127.35 341.1 128.55 342.3 ;
        RECT  131.55 341.1 132.75 342.3 ;
        RECT  133.95 336.6 135.15 342.3 ;
        RECT  129.45 343.5 130.65 343.8 ;
        RECT  123.75 343.8 135.15 345.0 ;
        RECT  125.85 345.9 128.55 347.1 ;
        RECT  130.05 345.9 132.75 347.1 ;
        RECT  123.75 360.6 135.15 361.8 ;
        RECT  124.95 358.5 126.15 360.6 ;
        RECT  127.95 358.5 129.15 359.7 ;
        RECT  130.95 358.5 132.15 359.7 ;
        RECT  133.95 358.5 135.15 360.6 ;
        RECT  127.65 357.6 128.85 358.5 ;
        RECT  124.95 351.9 126.15 357.6 ;
        RECT  127.65 356.4 130.05 357.6 ;
        RECT  127.65 353.1 128.85 356.4 ;
        RECT  131.25 354.9 132.45 358.5 ;
        RECT  130.65 353.7 132.45 354.9 ;
        RECT  131.25 353.1 132.45 353.7 ;
        RECT  127.35 351.9 128.55 353.1 ;
        RECT  131.55 351.9 132.75 353.1 ;
        RECT  133.95 351.9 135.15 357.6 ;
        RECT  129.45 350.4 130.65 350.7 ;
        RECT  123.75 349.2 135.15 350.4 ;
        RECT  125.85 347.1 128.55 348.3 ;
        RECT  130.05 347.1 132.75 348.3 ;
        RECT  123.75 361.8 135.15 363.0 ;
        RECT  124.95 363.0 126.15 365.1 ;
        RECT  127.95 363.9 129.15 365.1 ;
        RECT  130.95 363.9 132.15 365.1 ;
        RECT  133.95 363.0 135.15 365.1 ;
        RECT  127.65 365.1 128.85 366.0 ;
        RECT  124.95 366.0 126.15 371.7 ;
        RECT  127.65 366.0 130.05 367.2 ;
        RECT  127.65 367.2 128.85 370.5 ;
        RECT  131.25 365.1 132.45 368.7 ;
        RECT  130.65 368.7 132.45 369.9 ;
        RECT  131.25 369.9 132.45 370.5 ;
        RECT  127.35 370.5 128.55 371.7 ;
        RECT  131.55 370.5 132.75 371.7 ;
        RECT  133.95 366.0 135.15 371.7 ;
        RECT  129.45 372.9 130.65 373.2 ;
        RECT  123.75 373.2 135.15 374.4 ;
        RECT  125.85 375.3 128.55 376.5 ;
        RECT  130.05 375.3 132.75 376.5 ;
        RECT  123.75 390.0 135.15 391.2 ;
        RECT  124.95 387.9 126.15 390.0 ;
        RECT  127.95 387.9 129.15 389.1 ;
        RECT  130.95 387.9 132.15 389.1 ;
        RECT  133.95 387.9 135.15 390.0 ;
        RECT  127.65 387.0 128.85 387.9 ;
        RECT  124.95 381.3 126.15 387.0 ;
        RECT  127.65 385.8 130.05 387.0 ;
        RECT  127.65 382.5 128.85 385.8 ;
        RECT  131.25 384.3 132.45 387.9 ;
        RECT  130.65 383.1 132.45 384.3 ;
        RECT  131.25 382.5 132.45 383.1 ;
        RECT  127.35 381.3 128.55 382.5 ;
        RECT  131.55 381.3 132.75 382.5 ;
        RECT  133.95 381.3 135.15 387.0 ;
        RECT  129.45 379.8 130.65 380.1 ;
        RECT  123.75 378.6 135.15 379.8 ;
        RECT  125.85 376.5 128.55 377.7 ;
        RECT  130.05 376.5 132.75 377.7 ;
        RECT  123.75 391.2 135.15 392.4 ;
        RECT  124.95 392.4 126.15 394.5 ;
        RECT  127.95 393.3 129.15 394.5 ;
        RECT  130.95 393.3 132.15 394.5 ;
        RECT  133.95 392.4 135.15 394.5 ;
        RECT  127.65 394.5 128.85 395.4 ;
        RECT  124.95 395.4 126.15 401.1 ;
        RECT  127.65 395.4 130.05 396.6 ;
        RECT  127.65 396.6 128.85 399.9 ;
        RECT  131.25 394.5 132.45 398.1 ;
        RECT  130.65 398.1 132.45 399.3 ;
        RECT  131.25 399.3 132.45 399.9 ;
        RECT  127.35 399.9 128.55 401.1 ;
        RECT  131.55 399.9 132.75 401.1 ;
        RECT  133.95 395.4 135.15 401.1 ;
        RECT  129.45 402.3 130.65 402.6 ;
        RECT  123.75 402.6 135.15 403.8 ;
        RECT  125.85 404.7 128.55 405.9 ;
        RECT  130.05 404.7 132.75 405.9 ;
        RECT  123.75 419.4 135.15 420.6 ;
        RECT  124.95 417.3 126.15 419.4 ;
        RECT  127.95 417.3 129.15 418.5 ;
        RECT  130.95 417.3 132.15 418.5 ;
        RECT  133.95 417.3 135.15 419.4 ;
        RECT  127.65 416.4 128.85 417.3 ;
        RECT  124.95 410.7 126.15 416.4 ;
        RECT  127.65 415.2 130.05 416.4 ;
        RECT  127.65 411.9 128.85 415.2 ;
        RECT  131.25 413.7 132.45 417.3 ;
        RECT  130.65 412.5 132.45 413.7 ;
        RECT  131.25 411.9 132.45 412.5 ;
        RECT  127.35 410.7 128.55 411.9 ;
        RECT  131.55 410.7 132.75 411.9 ;
        RECT  133.95 410.7 135.15 416.4 ;
        RECT  129.45 409.2 130.65 409.5 ;
        RECT  123.75 408.0 135.15 409.2 ;
        RECT  125.85 405.9 128.55 407.1 ;
        RECT  130.05 405.9 132.75 407.1 ;
        RECT  123.75 420.6 135.15 421.8 ;
        RECT  124.95 421.8 126.15 423.9 ;
        RECT  127.95 422.7 129.15 423.9 ;
        RECT  130.95 422.7 132.15 423.9 ;
        RECT  133.95 421.8 135.15 423.9 ;
        RECT  127.65 423.9 128.85 424.8 ;
        RECT  124.95 424.8 126.15 430.5 ;
        RECT  127.65 424.8 130.05 426.0 ;
        RECT  127.65 426.0 128.85 429.3 ;
        RECT  131.25 423.9 132.45 427.5 ;
        RECT  130.65 427.5 132.45 428.7 ;
        RECT  131.25 428.7 132.45 429.3 ;
        RECT  127.35 429.3 128.55 430.5 ;
        RECT  131.55 429.3 132.75 430.5 ;
        RECT  133.95 424.8 135.15 430.5 ;
        RECT  129.45 431.7 130.65 432.0 ;
        RECT  123.75 432.0 135.15 433.2 ;
        RECT  125.85 434.1 128.55 435.3 ;
        RECT  130.05 434.1 132.75 435.3 ;
        RECT  133.95 213.6 145.35 214.8 ;
        RECT  135.15 211.5 136.35 213.6 ;
        RECT  138.15 211.5 139.35 212.7 ;
        RECT  141.15 211.5 142.35 212.7 ;
        RECT  144.15 211.5 145.35 213.6 ;
        RECT  137.85 210.6 139.05 211.5 ;
        RECT  135.15 204.9 136.35 210.6 ;
        RECT  137.85 209.4 140.25 210.6 ;
        RECT  137.85 206.1 139.05 209.4 ;
        RECT  141.45 207.9 142.65 211.5 ;
        RECT  140.85 206.7 142.65 207.9 ;
        RECT  141.45 206.1 142.65 206.7 ;
        RECT  137.55 204.9 138.75 206.1 ;
        RECT  141.75 204.9 142.95 206.1 ;
        RECT  144.15 204.9 145.35 210.6 ;
        RECT  139.65 203.4 140.85 203.7 ;
        RECT  133.95 202.2 145.35 203.4 ;
        RECT  136.05 200.1 138.75 201.3 ;
        RECT  140.25 200.1 142.95 201.3 ;
        RECT  133.95 214.8 145.35 216.0 ;
        RECT  135.15 216.0 136.35 218.1 ;
        RECT  138.15 216.9 139.35 218.1 ;
        RECT  141.15 216.9 142.35 218.1 ;
        RECT  144.15 216.0 145.35 218.1 ;
        RECT  137.85 218.1 139.05 219.0 ;
        RECT  135.15 219.0 136.35 224.7 ;
        RECT  137.85 219.0 140.25 220.2 ;
        RECT  137.85 220.2 139.05 223.5 ;
        RECT  141.45 218.1 142.65 221.7 ;
        RECT  140.85 221.7 142.65 222.9 ;
        RECT  141.45 222.9 142.65 223.5 ;
        RECT  137.55 223.5 138.75 224.7 ;
        RECT  141.75 223.5 142.95 224.7 ;
        RECT  144.15 219.0 145.35 224.7 ;
        RECT  139.65 225.9 140.85 226.2 ;
        RECT  133.95 226.2 145.35 227.4 ;
        RECT  136.05 228.3 138.75 229.5 ;
        RECT  140.25 228.3 142.95 229.5 ;
        RECT  133.95 243.0 145.35 244.2 ;
        RECT  135.15 240.9 136.35 243.0 ;
        RECT  138.15 240.9 139.35 242.1 ;
        RECT  141.15 240.9 142.35 242.1 ;
        RECT  144.15 240.9 145.35 243.0 ;
        RECT  137.85 240.0 139.05 240.9 ;
        RECT  135.15 234.3 136.35 240.0 ;
        RECT  137.85 238.8 140.25 240.0 ;
        RECT  137.85 235.5 139.05 238.8 ;
        RECT  141.45 237.3 142.65 240.9 ;
        RECT  140.85 236.1 142.65 237.3 ;
        RECT  141.45 235.5 142.65 236.1 ;
        RECT  137.55 234.3 138.75 235.5 ;
        RECT  141.75 234.3 142.95 235.5 ;
        RECT  144.15 234.3 145.35 240.0 ;
        RECT  139.65 232.8 140.85 233.1 ;
        RECT  133.95 231.6 145.35 232.8 ;
        RECT  136.05 229.5 138.75 230.7 ;
        RECT  140.25 229.5 142.95 230.7 ;
        RECT  133.95 244.2 145.35 245.4 ;
        RECT  135.15 245.4 136.35 247.5 ;
        RECT  138.15 246.3 139.35 247.5 ;
        RECT  141.15 246.3 142.35 247.5 ;
        RECT  144.15 245.4 145.35 247.5 ;
        RECT  137.85 247.5 139.05 248.4 ;
        RECT  135.15 248.4 136.35 254.1 ;
        RECT  137.85 248.4 140.25 249.6 ;
        RECT  137.85 249.6 139.05 252.9 ;
        RECT  141.45 247.5 142.65 251.1 ;
        RECT  140.85 251.1 142.65 252.3 ;
        RECT  141.45 252.3 142.65 252.9 ;
        RECT  137.55 252.9 138.75 254.1 ;
        RECT  141.75 252.9 142.95 254.1 ;
        RECT  144.15 248.4 145.35 254.1 ;
        RECT  139.65 255.3 140.85 255.6 ;
        RECT  133.95 255.6 145.35 256.8 ;
        RECT  136.05 257.7 138.75 258.9 ;
        RECT  140.25 257.7 142.95 258.9 ;
        RECT  133.95 272.4 145.35 273.6 ;
        RECT  135.15 270.3 136.35 272.4 ;
        RECT  138.15 270.3 139.35 271.5 ;
        RECT  141.15 270.3 142.35 271.5 ;
        RECT  144.15 270.3 145.35 272.4 ;
        RECT  137.85 269.4 139.05 270.3 ;
        RECT  135.15 263.7 136.35 269.4 ;
        RECT  137.85 268.2 140.25 269.4 ;
        RECT  137.85 264.9 139.05 268.2 ;
        RECT  141.45 266.7 142.65 270.3 ;
        RECT  140.85 265.5 142.65 266.7 ;
        RECT  141.45 264.9 142.65 265.5 ;
        RECT  137.55 263.7 138.75 264.9 ;
        RECT  141.75 263.7 142.95 264.9 ;
        RECT  144.15 263.7 145.35 269.4 ;
        RECT  139.65 262.2 140.85 262.5 ;
        RECT  133.95 261.0 145.35 262.2 ;
        RECT  136.05 258.9 138.75 260.1 ;
        RECT  140.25 258.9 142.95 260.1 ;
        RECT  133.95 273.6 145.35 274.8 ;
        RECT  135.15 274.8 136.35 276.9 ;
        RECT  138.15 275.7 139.35 276.9 ;
        RECT  141.15 275.7 142.35 276.9 ;
        RECT  144.15 274.8 145.35 276.9 ;
        RECT  137.85 276.9 139.05 277.8 ;
        RECT  135.15 277.8 136.35 283.5 ;
        RECT  137.85 277.8 140.25 279.0 ;
        RECT  137.85 279.0 139.05 282.3 ;
        RECT  141.45 276.9 142.65 280.5 ;
        RECT  140.85 280.5 142.65 281.7 ;
        RECT  141.45 281.7 142.65 282.3 ;
        RECT  137.55 282.3 138.75 283.5 ;
        RECT  141.75 282.3 142.95 283.5 ;
        RECT  144.15 277.8 145.35 283.5 ;
        RECT  139.65 284.7 140.85 285.0 ;
        RECT  133.95 285.0 145.35 286.2 ;
        RECT  136.05 287.1 138.75 288.3 ;
        RECT  140.25 287.1 142.95 288.3 ;
        RECT  133.95 301.8 145.35 303.0 ;
        RECT  135.15 299.7 136.35 301.8 ;
        RECT  138.15 299.7 139.35 300.9 ;
        RECT  141.15 299.7 142.35 300.9 ;
        RECT  144.15 299.7 145.35 301.8 ;
        RECT  137.85 298.8 139.05 299.7 ;
        RECT  135.15 293.1 136.35 298.8 ;
        RECT  137.85 297.6 140.25 298.8 ;
        RECT  137.85 294.3 139.05 297.6 ;
        RECT  141.45 296.1 142.65 299.7 ;
        RECT  140.85 294.9 142.65 296.1 ;
        RECT  141.45 294.3 142.65 294.9 ;
        RECT  137.55 293.1 138.75 294.3 ;
        RECT  141.75 293.1 142.95 294.3 ;
        RECT  144.15 293.1 145.35 298.8 ;
        RECT  139.65 291.6 140.85 291.9 ;
        RECT  133.95 290.4 145.35 291.6 ;
        RECT  136.05 288.3 138.75 289.5 ;
        RECT  140.25 288.3 142.95 289.5 ;
        RECT  133.95 303.0 145.35 304.2 ;
        RECT  135.15 304.2 136.35 306.3 ;
        RECT  138.15 305.1 139.35 306.3 ;
        RECT  141.15 305.1 142.35 306.3 ;
        RECT  144.15 304.2 145.35 306.3 ;
        RECT  137.85 306.3 139.05 307.2 ;
        RECT  135.15 307.2 136.35 312.9 ;
        RECT  137.85 307.2 140.25 308.4 ;
        RECT  137.85 308.4 139.05 311.7 ;
        RECT  141.45 306.3 142.65 309.9 ;
        RECT  140.85 309.9 142.65 311.1 ;
        RECT  141.45 311.1 142.65 311.7 ;
        RECT  137.55 311.7 138.75 312.9 ;
        RECT  141.75 311.7 142.95 312.9 ;
        RECT  144.15 307.2 145.35 312.9 ;
        RECT  139.65 314.1 140.85 314.4 ;
        RECT  133.95 314.4 145.35 315.6 ;
        RECT  136.05 316.5 138.75 317.7 ;
        RECT  140.25 316.5 142.95 317.7 ;
        RECT  133.95 331.2 145.35 332.4 ;
        RECT  135.15 329.1 136.35 331.2 ;
        RECT  138.15 329.1 139.35 330.3 ;
        RECT  141.15 329.1 142.35 330.3 ;
        RECT  144.15 329.1 145.35 331.2 ;
        RECT  137.85 328.2 139.05 329.1 ;
        RECT  135.15 322.5 136.35 328.2 ;
        RECT  137.85 327.0 140.25 328.2 ;
        RECT  137.85 323.7 139.05 327.0 ;
        RECT  141.45 325.5 142.65 329.1 ;
        RECT  140.85 324.3 142.65 325.5 ;
        RECT  141.45 323.7 142.65 324.3 ;
        RECT  137.55 322.5 138.75 323.7 ;
        RECT  141.75 322.5 142.95 323.7 ;
        RECT  144.15 322.5 145.35 328.2 ;
        RECT  139.65 321.0 140.85 321.3 ;
        RECT  133.95 319.8 145.35 321.0 ;
        RECT  136.05 317.7 138.75 318.9 ;
        RECT  140.25 317.7 142.95 318.9 ;
        RECT  133.95 332.4 145.35 333.6 ;
        RECT  135.15 333.6 136.35 335.7 ;
        RECT  138.15 334.5 139.35 335.7 ;
        RECT  141.15 334.5 142.35 335.7 ;
        RECT  144.15 333.6 145.35 335.7 ;
        RECT  137.85 335.7 139.05 336.6 ;
        RECT  135.15 336.6 136.35 342.3 ;
        RECT  137.85 336.6 140.25 337.8 ;
        RECT  137.85 337.8 139.05 341.1 ;
        RECT  141.45 335.7 142.65 339.3 ;
        RECT  140.85 339.3 142.65 340.5 ;
        RECT  141.45 340.5 142.65 341.1 ;
        RECT  137.55 341.1 138.75 342.3 ;
        RECT  141.75 341.1 142.95 342.3 ;
        RECT  144.15 336.6 145.35 342.3 ;
        RECT  139.65 343.5 140.85 343.8 ;
        RECT  133.95 343.8 145.35 345.0 ;
        RECT  136.05 345.9 138.75 347.1 ;
        RECT  140.25 345.9 142.95 347.1 ;
        RECT  133.95 360.6 145.35 361.8 ;
        RECT  135.15 358.5 136.35 360.6 ;
        RECT  138.15 358.5 139.35 359.7 ;
        RECT  141.15 358.5 142.35 359.7 ;
        RECT  144.15 358.5 145.35 360.6 ;
        RECT  137.85 357.6 139.05 358.5 ;
        RECT  135.15 351.9 136.35 357.6 ;
        RECT  137.85 356.4 140.25 357.6 ;
        RECT  137.85 353.1 139.05 356.4 ;
        RECT  141.45 354.9 142.65 358.5 ;
        RECT  140.85 353.7 142.65 354.9 ;
        RECT  141.45 353.1 142.65 353.7 ;
        RECT  137.55 351.9 138.75 353.1 ;
        RECT  141.75 351.9 142.95 353.1 ;
        RECT  144.15 351.9 145.35 357.6 ;
        RECT  139.65 350.4 140.85 350.7 ;
        RECT  133.95 349.2 145.35 350.4 ;
        RECT  136.05 347.1 138.75 348.3 ;
        RECT  140.25 347.1 142.95 348.3 ;
        RECT  133.95 361.8 145.35 363.0 ;
        RECT  135.15 363.0 136.35 365.1 ;
        RECT  138.15 363.9 139.35 365.1 ;
        RECT  141.15 363.9 142.35 365.1 ;
        RECT  144.15 363.0 145.35 365.1 ;
        RECT  137.85 365.1 139.05 366.0 ;
        RECT  135.15 366.0 136.35 371.7 ;
        RECT  137.85 366.0 140.25 367.2 ;
        RECT  137.85 367.2 139.05 370.5 ;
        RECT  141.45 365.1 142.65 368.7 ;
        RECT  140.85 368.7 142.65 369.9 ;
        RECT  141.45 369.9 142.65 370.5 ;
        RECT  137.55 370.5 138.75 371.7 ;
        RECT  141.75 370.5 142.95 371.7 ;
        RECT  144.15 366.0 145.35 371.7 ;
        RECT  139.65 372.9 140.85 373.2 ;
        RECT  133.95 373.2 145.35 374.4 ;
        RECT  136.05 375.3 138.75 376.5 ;
        RECT  140.25 375.3 142.95 376.5 ;
        RECT  133.95 390.0 145.35 391.2 ;
        RECT  135.15 387.9 136.35 390.0 ;
        RECT  138.15 387.9 139.35 389.1 ;
        RECT  141.15 387.9 142.35 389.1 ;
        RECT  144.15 387.9 145.35 390.0 ;
        RECT  137.85 387.0 139.05 387.9 ;
        RECT  135.15 381.3 136.35 387.0 ;
        RECT  137.85 385.8 140.25 387.0 ;
        RECT  137.85 382.5 139.05 385.8 ;
        RECT  141.45 384.3 142.65 387.9 ;
        RECT  140.85 383.1 142.65 384.3 ;
        RECT  141.45 382.5 142.65 383.1 ;
        RECT  137.55 381.3 138.75 382.5 ;
        RECT  141.75 381.3 142.95 382.5 ;
        RECT  144.15 381.3 145.35 387.0 ;
        RECT  139.65 379.8 140.85 380.1 ;
        RECT  133.95 378.6 145.35 379.8 ;
        RECT  136.05 376.5 138.75 377.7 ;
        RECT  140.25 376.5 142.95 377.7 ;
        RECT  133.95 391.2 145.35 392.4 ;
        RECT  135.15 392.4 136.35 394.5 ;
        RECT  138.15 393.3 139.35 394.5 ;
        RECT  141.15 393.3 142.35 394.5 ;
        RECT  144.15 392.4 145.35 394.5 ;
        RECT  137.85 394.5 139.05 395.4 ;
        RECT  135.15 395.4 136.35 401.1 ;
        RECT  137.85 395.4 140.25 396.6 ;
        RECT  137.85 396.6 139.05 399.9 ;
        RECT  141.45 394.5 142.65 398.1 ;
        RECT  140.85 398.1 142.65 399.3 ;
        RECT  141.45 399.3 142.65 399.9 ;
        RECT  137.55 399.9 138.75 401.1 ;
        RECT  141.75 399.9 142.95 401.1 ;
        RECT  144.15 395.4 145.35 401.1 ;
        RECT  139.65 402.3 140.85 402.6 ;
        RECT  133.95 402.6 145.35 403.8 ;
        RECT  136.05 404.7 138.75 405.9 ;
        RECT  140.25 404.7 142.95 405.9 ;
        RECT  133.95 419.4 145.35 420.6 ;
        RECT  135.15 417.3 136.35 419.4 ;
        RECT  138.15 417.3 139.35 418.5 ;
        RECT  141.15 417.3 142.35 418.5 ;
        RECT  144.15 417.3 145.35 419.4 ;
        RECT  137.85 416.4 139.05 417.3 ;
        RECT  135.15 410.7 136.35 416.4 ;
        RECT  137.85 415.2 140.25 416.4 ;
        RECT  137.85 411.9 139.05 415.2 ;
        RECT  141.45 413.7 142.65 417.3 ;
        RECT  140.85 412.5 142.65 413.7 ;
        RECT  141.45 411.9 142.65 412.5 ;
        RECT  137.55 410.7 138.75 411.9 ;
        RECT  141.75 410.7 142.95 411.9 ;
        RECT  144.15 410.7 145.35 416.4 ;
        RECT  139.65 409.2 140.85 409.5 ;
        RECT  133.95 408.0 145.35 409.2 ;
        RECT  136.05 405.9 138.75 407.1 ;
        RECT  140.25 405.9 142.95 407.1 ;
        RECT  133.95 420.6 145.35 421.8 ;
        RECT  135.15 421.8 136.35 423.9 ;
        RECT  138.15 422.7 139.35 423.9 ;
        RECT  141.15 422.7 142.35 423.9 ;
        RECT  144.15 421.8 145.35 423.9 ;
        RECT  137.85 423.9 139.05 424.8 ;
        RECT  135.15 424.8 136.35 430.5 ;
        RECT  137.85 424.8 140.25 426.0 ;
        RECT  137.85 426.0 139.05 429.3 ;
        RECT  141.45 423.9 142.65 427.5 ;
        RECT  140.85 427.5 142.65 428.7 ;
        RECT  141.45 428.7 142.65 429.3 ;
        RECT  137.55 429.3 138.75 430.5 ;
        RECT  141.75 429.3 142.95 430.5 ;
        RECT  144.15 424.8 145.35 430.5 ;
        RECT  139.65 431.7 140.85 432.0 ;
        RECT  133.95 432.0 145.35 433.2 ;
        RECT  136.05 434.1 138.75 435.3 ;
        RECT  140.25 434.1 142.95 435.3 ;
        RECT  124.35 458.4 144.75 459.3 ;
        RECT  124.35 446.4 144.75 447.3 ;
        RECT  124.35 446.4 134.55 447.3 ;
        RECT  124.35 458.4 134.55 459.3 ;
        RECT  129.75 450.9 130.65 459.3 ;
        RECT  127.35 442.5 128.55 443.7 ;
        RECT  129.75 442.5 130.95 443.7 ;
        RECT  127.35 450.9 128.55 452.1 ;
        RECT  129.75 450.9 130.95 452.1 ;
        RECT  129.75 450.9 130.95 452.1 ;
        RECT  132.15 450.9 133.35 452.1 ;
        RECT  128.25 446.4 129.45 447.6 ;
        RECT  129.75 456.3 130.95 457.5 ;
        RECT  127.35 450.9 128.55 452.1 ;
        RECT  132.15 450.9 133.35 452.1 ;
        RECT  127.35 442.5 128.55 443.7 ;
        RECT  129.75 442.5 130.95 443.7 ;
        RECT  134.55 446.4 144.75 447.3 ;
        RECT  134.55 458.4 144.75 459.3 ;
        RECT  139.95 450.9 140.85 459.3 ;
        RECT  137.55 442.5 138.75 443.7 ;
        RECT  139.95 442.5 141.15 443.7 ;
        RECT  137.55 450.9 138.75 452.1 ;
        RECT  139.95 450.9 141.15 452.1 ;
        RECT  139.95 450.9 141.15 452.1 ;
        RECT  142.35 450.9 143.55 452.1 ;
        RECT  138.45 446.4 139.65 447.6 ;
        RECT  139.95 456.3 141.15 457.5 ;
        RECT  137.55 450.9 138.75 452.1 ;
        RECT  142.35 450.9 143.55 452.1 ;
        RECT  137.55 442.5 138.75 443.7 ;
        RECT  139.95 442.5 141.15 443.7 ;
        RECT  124.35 168.75 144.75 169.65 ;
        RECT  124.35 193.95 144.75 194.85 ;
        RECT  124.35 196.05 144.75 196.95 ;
        RECT  123.75 195.9 135.15 197.1 ;
        RECT  123.75 193.8 135.15 195.0 ;
        RECT  129.15 190.2 130.35 192.9 ;
        RECT  131.55 190.2 132.75 193.8 ;
        RECT  133.95 192.6 135.15 193.8 ;
        RECT  129.15 186.3 130.05 190.2 ;
        RECT  126.45 171.9 127.65 186.3 ;
        RECT  128.85 183.6 130.05 186.3 ;
        RECT  131.25 182.7 132.45 186.3 ;
        RECT  131.25 181.5 133.35 182.7 ;
        RECT  128.85 174.6 130.05 180.0 ;
        RECT  131.25 174.6 132.45 181.5 ;
        RECT  128.85 173.7 129.75 174.6 ;
        RECT  128.85 172.8 130.65 173.7 ;
        RECT  126.45 170.7 128.25 171.9 ;
        RECT  129.75 171.0 130.65 172.8 ;
        RECT  129.75 169.8 130.95 171.0 ;
        RECT  123.75 168.6 135.15 169.8 ;
        RECT  127.05 167.4 128.25 167.7 ;
        RECT  126.15 166.5 128.25 167.4 ;
        RECT  133.05 166.5 134.55 167.7 ;
        RECT  126.15 164.4 127.05 166.5 ;
        RECT  128.25 164.4 129.45 165.6 ;
        RECT  126.15 158.1 127.35 164.4 ;
        RECT  125.25 157.2 127.35 158.1 ;
        RECT  128.55 157.2 129.75 164.4 ;
        RECT  130.95 157.2 132.15 165.6 ;
        RECT  133.65 164.4 134.55 166.5 ;
        RECT  133.35 157.2 134.55 164.4 ;
        RECT  125.25 154.5 126.45 157.2 ;
        RECT  133.95 195.9 145.35 197.1 ;
        RECT  133.95 193.8 145.35 195.0 ;
        RECT  139.35 190.2 140.55 192.9 ;
        RECT  141.75 190.2 142.95 193.8 ;
        RECT  144.15 192.6 145.35 193.8 ;
        RECT  139.35 186.3 140.25 190.2 ;
        RECT  136.65 171.9 137.85 186.3 ;
        RECT  139.05 183.6 140.25 186.3 ;
        RECT  141.45 182.7 142.65 186.3 ;
        RECT  141.45 181.5 143.55 182.7 ;
        RECT  139.05 174.6 140.25 180.0 ;
        RECT  141.45 174.6 142.65 181.5 ;
        RECT  139.05 173.7 139.95 174.6 ;
        RECT  139.05 172.8 140.85 173.7 ;
        RECT  136.65 170.7 138.45 171.9 ;
        RECT  139.95 171.0 140.85 172.8 ;
        RECT  139.95 169.8 141.15 171.0 ;
        RECT  133.95 168.6 145.35 169.8 ;
        RECT  137.25 167.4 138.45 167.7 ;
        RECT  136.35 166.5 138.45 167.4 ;
        RECT  143.25 166.5 144.75 167.7 ;
        RECT  136.35 164.4 137.25 166.5 ;
        RECT  138.45 164.4 139.65 165.6 ;
        RECT  136.35 158.1 137.55 164.4 ;
        RECT  135.45 157.2 137.55 158.1 ;
        RECT  138.75 157.2 139.95 164.4 ;
        RECT  141.15 157.2 142.35 165.6 ;
        RECT  143.85 164.4 144.75 166.5 ;
        RECT  143.55 157.2 144.75 164.4 ;
        RECT  135.45 154.5 136.65 157.2 ;
        RECT  124.35 97.95 144.75 98.85 ;
        RECT  124.35 100.05 144.75 100.95 ;
        RECT  124.35 95.85 144.75 96.75 ;
        RECT  125.85 147.9 127.05 149.1 ;
        RECT  125.85 147.3 126.75 147.9 ;
        RECT  125.55 143.7 126.75 147.3 ;
        RECT  127.95 143.7 129.15 147.3 ;
        RECT  130.35 143.7 131.55 148.5 ;
        RECT  132.75 144.9 134.25 146.1 ;
        RECT  128.25 141.3 129.15 143.7 ;
        RECT  125.55 128.1 126.75 140.7 ;
        RECT  128.25 140.1 132.45 141.3 ;
        RECT  127.65 137.7 132.45 138.9 ;
        RECT  127.95 133.8 129.15 137.7 ;
        RECT  130.35 133.2 131.55 135.0 ;
        RECT  133.35 133.2 134.25 144.9 ;
        RECT  130.35 132.0 134.25 133.2 ;
        RECT  127.95 127.2 129.15 130.2 ;
        RECT  130.35 128.1 131.55 132.0 ;
        RECT  124.35 126.0 135.15 127.2 ;
        RECT  125.85 121.8 127.05 124.8 ;
        RECT  128.25 122.7 129.45 126.0 ;
        RECT  130.65 121.8 131.85 124.8 ;
        RECT  125.85 120.9 131.85 121.8 ;
        RECT  125.85 115.2 127.05 120.9 ;
        RECT  130.65 120.6 131.85 120.9 ;
        RECT  130.65 119.4 132.45 120.6 ;
        RECT  128.25 115.2 129.45 117.3 ;
        RECT  130.65 116.4 131.85 117.3 ;
        RECT  130.65 115.2 134.55 116.4 ;
        RECT  131.25 113.1 133.65 114.3 ;
        RECT  125.25 111.9 126.45 113.1 ;
        RECT  125.55 109.8 126.45 111.9 ;
        RECT  125.25 105.9 126.45 109.8 ;
        RECT  127.65 107.7 128.85 109.8 ;
        RECT  130.05 107.7 131.25 111.0 ;
        RECT  125.25 105.0 128.85 105.9 ;
        RECT  125.25 101.1 126.45 104.1 ;
        RECT  127.65 102.0 128.85 105.0 ;
        RECT  130.05 101.1 131.25 104.1 ;
        RECT  132.45 102.0 133.65 113.1 ;
        RECT  124.35 99.9 135.15 101.1 ;
        RECT  124.35 97.8 135.15 99.0 ;
        RECT  124.35 95.7 135.15 96.9 ;
        RECT  127.95 93.6 130.35 94.8 ;
        RECT  136.05 147.9 137.25 149.1 ;
        RECT  136.05 147.3 136.95 147.9 ;
        RECT  135.75 143.7 136.95 147.3 ;
        RECT  138.15 143.7 139.35 147.3 ;
        RECT  140.55 143.7 141.75 148.5 ;
        RECT  142.95 144.9 144.45 146.1 ;
        RECT  138.45 141.3 139.35 143.7 ;
        RECT  135.75 128.1 136.95 140.7 ;
        RECT  138.45 140.1 142.65 141.3 ;
        RECT  137.85 137.7 142.65 138.9 ;
        RECT  138.15 133.8 139.35 137.7 ;
        RECT  140.55 133.2 141.75 135.0 ;
        RECT  143.55 133.2 144.45 144.9 ;
        RECT  140.55 132.0 144.45 133.2 ;
        RECT  138.15 127.2 139.35 130.2 ;
        RECT  140.55 128.1 141.75 132.0 ;
        RECT  134.55 126.0 145.35 127.2 ;
        RECT  136.05 121.8 137.25 124.8 ;
        RECT  138.45 122.7 139.65 126.0 ;
        RECT  140.85 121.8 142.05 124.8 ;
        RECT  136.05 120.9 142.05 121.8 ;
        RECT  136.05 115.2 137.25 120.9 ;
        RECT  140.85 120.6 142.05 120.9 ;
        RECT  140.85 119.4 142.65 120.6 ;
        RECT  138.45 115.2 139.65 117.3 ;
        RECT  140.85 116.4 142.05 117.3 ;
        RECT  140.85 115.2 144.75 116.4 ;
        RECT  141.45 113.1 143.85 114.3 ;
        RECT  135.45 111.9 136.65 113.1 ;
        RECT  135.75 109.8 136.65 111.9 ;
        RECT  135.45 105.9 136.65 109.8 ;
        RECT  137.85 107.7 139.05 109.8 ;
        RECT  140.25 107.7 141.45 111.0 ;
        RECT  135.45 105.0 139.05 105.9 ;
        RECT  135.45 101.1 136.65 104.1 ;
        RECT  137.85 102.0 139.05 105.0 ;
        RECT  140.25 101.1 141.45 104.1 ;
        RECT  142.65 102.0 143.85 113.1 ;
        RECT  134.55 99.9 145.35 101.1 ;
        RECT  134.55 97.8 145.35 99.0 ;
        RECT  134.55 95.7 145.35 96.9 ;
        RECT  138.15 93.6 140.55 94.8 ;
        RECT  124.35 32.85 144.75 33.75 ;
        RECT  124.35 87.3 144.75 88.2 ;
        RECT  123.75 87.3 135.15 88.2 ;
        RECT  123.75 84.0 124.95 87.3 ;
        RECT  126.15 85.5 132.75 86.4 ;
        RECT  126.15 85.2 129.15 85.5 ;
        RECT  131.55 85.2 132.75 85.5 ;
        RECT  123.75 82.8 127.95 84.0 ;
        RECT  131.55 82.8 135.15 84.0 ;
        RECT  123.75 79.2 124.95 82.8 ;
        RECT  129.15 81.9 130.35 82.8 ;
        RECT  129.15 81.6 131.55 81.9 ;
        RECT  126.15 80.7 132.75 81.6 ;
        RECT  126.15 80.4 127.95 80.7 ;
        RECT  131.55 80.4 132.75 80.7 ;
        RECT  123.75 78.0 127.95 79.2 ;
        RECT  123.75 64.2 124.95 78.0 ;
        RECT  129.45 77.4 130.65 79.8 ;
        RECT  134.25 79.2 135.15 82.8 ;
        RECT  131.55 78.0 135.15 79.2 ;
        RECT  133.95 76.8 135.15 78.0 ;
        RECT  126.15 74.4 127.35 75.6 ;
        RECT  128.25 75.3 130.65 76.5 ;
        RECT  126.15 73.5 132.75 74.4 ;
        RECT  126.15 73.2 127.95 73.5 ;
        RECT  131.55 73.2 132.75 73.5 ;
        RECT  126.15 71.1 132.75 72.0 ;
        RECT  126.15 70.8 127.95 71.1 ;
        RECT  130.35 70.8 132.75 71.1 ;
        RECT  126.15 68.7 132.75 69.6 ;
        RECT  126.15 68.4 127.95 68.7 ;
        RECT  130.35 68.4 132.75 68.7 ;
        RECT  129.15 66.6 130.35 67.5 ;
        RECT  126.15 65.7 132.75 66.6 ;
        RECT  126.15 65.4 129.15 65.7 ;
        RECT  131.55 65.4 132.75 65.7 ;
        RECT  123.75 63.0 127.95 64.2 ;
        RECT  123.75 58.5 124.95 63.0 ;
        RECT  128.85 62.1 130.05 64.5 ;
        RECT  134.25 64.2 135.15 76.8 ;
        RECT  131.55 63.0 135.15 64.2 ;
        RECT  126.15 60.9 127.35 62.1 ;
        RECT  126.15 60.0 132.75 60.9 ;
        RECT  126.15 59.7 127.95 60.0 ;
        RECT  131.55 59.7 132.75 60.0 ;
        RECT  134.25 58.5 135.15 63.0 ;
        RECT  123.75 57.3 127.95 58.5 ;
        RECT  123.75 53.7 124.95 57.3 ;
        RECT  129.45 56.4 130.65 57.6 ;
        RECT  131.55 57.3 135.15 58.5 ;
        RECT  126.15 56.1 131.55 56.4 ;
        RECT  126.15 55.5 132.75 56.1 ;
        RECT  126.15 54.9 127.95 55.5 ;
        RECT  130.35 55.2 132.75 55.5 ;
        RECT  131.55 54.9 132.75 55.2 ;
        RECT  123.75 52.5 127.95 53.7 ;
        RECT  123.75 37.5 124.95 52.5 ;
        RECT  129.45 51.9 130.65 54.3 ;
        RECT  134.25 53.7 135.15 57.3 ;
        RECT  131.55 52.5 135.15 53.7 ;
        RECT  133.95 51.3 135.15 52.5 ;
        RECT  126.15 48.0 127.35 49.2 ;
        RECT  128.25 48.9 130.65 50.1 ;
        RECT  126.15 47.1 132.75 48.0 ;
        RECT  126.15 46.8 127.95 47.1 ;
        RECT  131.55 46.8 132.75 47.1 ;
        RECT  126.15 44.7 132.75 45.6 ;
        RECT  126.15 44.4 127.95 44.7 ;
        RECT  130.35 44.4 132.75 44.7 ;
        RECT  126.15 42.3 132.75 43.2 ;
        RECT  126.15 42.0 127.95 42.3 ;
        RECT  130.35 42.0 132.75 42.3 ;
        RECT  129.15 40.2 130.35 41.1 ;
        RECT  126.15 39.3 132.75 40.2 ;
        RECT  126.15 39.0 129.15 39.3 ;
        RECT  131.55 39.0 132.75 39.3 ;
        RECT  134.25 37.8 135.15 51.3 ;
        RECT  126.15 37.5 127.95 37.8 ;
        RECT  123.75 36.6 127.95 37.5 ;
        RECT  131.55 36.9 135.15 37.8 ;
        RECT  131.55 36.6 132.75 36.9 ;
        RECT  126.75 35.1 127.95 36.6 ;
        RECT  128.85 34.2 130.05 35.1 ;
        RECT  123.75 33.3 135.15 34.2 ;
        RECT  133.95 87.3 145.35 88.2 ;
        RECT  144.15 84.0 145.35 87.3 ;
        RECT  136.35 85.5 142.95 86.4 ;
        RECT  139.95 85.2 142.95 85.5 ;
        RECT  136.35 85.2 137.55 85.5 ;
        RECT  141.15 82.8 145.35 84.0 ;
        RECT  133.95 82.8 137.55 84.0 ;
        RECT  144.15 79.2 145.35 82.8 ;
        RECT  138.75 81.9 139.95 82.8 ;
        RECT  137.55 81.6 139.95 81.9 ;
        RECT  136.35 80.7 142.95 81.6 ;
        RECT  141.15 80.4 142.95 80.7 ;
        RECT  136.35 80.4 137.55 80.7 ;
        RECT  141.15 78.0 145.35 79.2 ;
        RECT  144.15 64.2 145.35 78.0 ;
        RECT  138.45 77.4 139.65 79.8 ;
        RECT  133.95 79.2 134.85 82.8 ;
        RECT  133.95 78.0 137.55 79.2 ;
        RECT  133.95 76.8 135.15 78.0 ;
        RECT  141.75 74.4 142.95 75.6 ;
        RECT  138.45 75.3 140.85 76.5 ;
        RECT  136.35 73.5 142.95 74.4 ;
        RECT  141.15 73.2 142.95 73.5 ;
        RECT  136.35 73.2 137.55 73.5 ;
        RECT  136.35 71.1 142.95 72.0 ;
        RECT  141.15 70.8 142.95 71.1 ;
        RECT  136.35 70.8 138.75 71.1 ;
        RECT  136.35 68.7 142.95 69.6 ;
        RECT  141.15 68.4 142.95 68.7 ;
        RECT  136.35 68.4 138.75 68.7 ;
        RECT  138.75 66.6 139.95 67.5 ;
        RECT  136.35 65.7 142.95 66.6 ;
        RECT  139.95 65.4 142.95 65.7 ;
        RECT  136.35 65.4 137.55 65.7 ;
        RECT  141.15 63.0 145.35 64.2 ;
        RECT  144.15 58.5 145.35 63.0 ;
        RECT  139.05 62.1 140.25 64.5 ;
        RECT  133.95 64.2 134.85 76.8 ;
        RECT  133.95 63.0 137.55 64.2 ;
        RECT  141.75 60.9 142.95 62.1 ;
        RECT  136.35 60.0 142.95 60.9 ;
        RECT  141.15 59.7 142.95 60.0 ;
        RECT  136.35 59.7 137.55 60.0 ;
        RECT  133.95 58.5 134.85 63.0 ;
        RECT  141.15 57.3 145.35 58.5 ;
        RECT  144.15 53.7 145.35 57.3 ;
        RECT  138.45 56.4 139.65 57.6 ;
        RECT  133.95 57.3 137.55 58.5 ;
        RECT  137.55 56.1 142.95 56.4 ;
        RECT  136.35 55.5 142.95 56.1 ;
        RECT  141.15 54.9 142.95 55.5 ;
        RECT  136.35 55.2 138.75 55.5 ;
        RECT  136.35 54.9 137.55 55.2 ;
        RECT  141.15 52.5 145.35 53.7 ;
        RECT  144.15 37.5 145.35 52.5 ;
        RECT  138.45 51.9 139.65 54.3 ;
        RECT  133.95 53.7 134.85 57.3 ;
        RECT  133.95 52.5 137.55 53.7 ;
        RECT  133.95 51.3 135.15 52.5 ;
        RECT  141.75 48.0 142.95 49.2 ;
        RECT  138.45 48.9 140.85 50.1 ;
        RECT  136.35 47.1 142.95 48.0 ;
        RECT  141.15 46.8 142.95 47.1 ;
        RECT  136.35 46.8 137.55 47.1 ;
        RECT  136.35 44.7 142.95 45.6 ;
        RECT  141.15 44.4 142.95 44.7 ;
        RECT  136.35 44.4 138.75 44.7 ;
        RECT  136.35 42.3 142.95 43.2 ;
        RECT  141.15 42.0 142.95 42.3 ;
        RECT  136.35 42.0 138.75 42.3 ;
        RECT  138.75 40.2 139.95 41.1 ;
        RECT  136.35 39.3 142.95 40.2 ;
        RECT  139.95 39.0 142.95 39.3 ;
        RECT  136.35 39.0 137.55 39.3 ;
        RECT  133.95 37.8 134.85 51.3 ;
        RECT  141.15 37.5 142.95 37.8 ;
        RECT  141.15 36.6 145.35 37.5 ;
        RECT  133.95 36.9 137.55 37.8 ;
        RECT  136.35 36.6 137.55 36.9 ;
        RECT  141.15 35.1 142.35 36.6 ;
        RECT  139.05 34.2 140.25 35.1 ;
        RECT  133.95 33.3 145.35 34.2 ;
        RECT  124.35 26.25 144.75 27.15 ;
        RECT  124.35 28.65 144.75 29.55 ;
        RECT  124.35 10.35 144.75 11.25 ;
        RECT  124.35 50.4 135.15 51.6 ;
        RECT  125.25 46.8 126.75 49.2 ;
        RECT  127.95 46.8 129.15 50.4 ;
        RECT  130.35 46.8 131.55 49.2 ;
        RECT  132.75 46.8 133.95 49.2 ;
        RECT  125.25 43.5 126.15 46.8 ;
        RECT  127.05 44.7 128.25 45.9 ;
        RECT  125.25 42.3 130.35 43.5 ;
        RECT  133.05 42.3 133.95 46.8 ;
        RECT  125.25 40.2 126.15 42.3 ;
        RECT  131.85 41.1 133.95 42.3 ;
        RECT  133.05 40.2 133.95 41.1 ;
        RECT  125.25 39.0 126.75 40.2 ;
        RECT  127.95 37.8 129.15 40.2 ;
        RECT  130.35 39.0 131.55 40.2 ;
        RECT  132.75 39.0 133.95 40.2 ;
        RECT  124.35 36.6 135.15 37.8 ;
        RECT  124.35 34.5 135.15 35.7 ;
        RECT  124.35 32.1 135.15 33.3 ;
        RECT  133.95 50.4 144.75 51.6 ;
        RECT  142.35 46.8 143.85 49.2 ;
        RECT  139.95 46.8 141.15 50.4 ;
        RECT  137.55 46.8 138.75 49.2 ;
        RECT  135.15 46.8 136.35 49.2 ;
        RECT  142.95 43.5 143.85 46.8 ;
        RECT  140.85 44.7 142.05 45.9 ;
        RECT  138.75 42.3 143.85 43.5 ;
        RECT  135.15 42.3 136.05 46.8 ;
        RECT  142.95 40.2 143.85 42.3 ;
        RECT  135.15 41.1 137.25 42.3 ;
        RECT  135.15 40.2 136.05 41.1 ;
        RECT  142.35 39.0 143.85 40.2 ;
        RECT  139.95 37.8 141.15 40.2 ;
        RECT  137.55 39.0 138.75 40.2 ;
        RECT  135.15 39.0 136.35 40.2 ;
        RECT  133.95 36.6 144.75 37.8 ;
        RECT  133.95 34.5 144.75 35.7 ;
        RECT  133.95 32.1 144.75 33.3 ;
        RECT  41.85 206.4 42.75 207.3 ;
        RECT  41.85 222.3 42.75 223.2 ;
        RECT  41.85 235.8 42.75 236.7 ;
        RECT  41.85 251.7 42.75 252.6 ;
        RECT  41.85 265.2 42.75 266.1 ;
        RECT  41.85 281.1 42.75 282.0 ;
        RECT  41.85 294.6 42.75 295.5 ;
        RECT  41.85 310.5 42.75 311.4 ;
        RECT  41.85 324.0 42.75 324.9 ;
        RECT  41.85 339.9 42.75 340.8 ;
        RECT  41.85 353.4 42.75 354.3 ;
        RECT  41.85 369.3 42.75 370.2 ;
        RECT  41.85 382.8 42.75 383.7 ;
        RECT  41.85 398.7 42.75 399.6 ;
        RECT  41.85 412.2 42.75 413.1 ;
        RECT  41.85 428.1 42.75 429.0 ;
        RECT  13.05 88.8 29.85 89.7 ;
        RECT  15.15 104.7 29.85 105.6 ;
        RECT  17.25 118.2 29.85 119.1 ;
        RECT  19.35 134.1 29.85 135.0 ;
        RECT  21.45 147.6 29.85 148.5 ;
        RECT  23.55 163.5 29.85 164.4 ;
        RECT  25.65 177.0 29.85 177.9 ;
        RECT  27.75 192.9 29.85 193.8 ;
        RECT  13.05 208.8 29.85 209.7 ;
        RECT  21.45 205.5 29.85 206.4 ;
        RECT  13.05 219.9 29.85 220.8 ;
        RECT  23.55 223.2 29.85 224.1 ;
        RECT  13.05 238.2 29.85 239.1 ;
        RECT  25.65 234.9 29.85 235.8 ;
        RECT  13.05 249.3 29.85 250.2 ;
        RECT  27.75 252.6 29.85 253.5 ;
        RECT  15.15 267.6 29.85 268.5 ;
        RECT  21.45 264.3 29.85 265.2 ;
        RECT  15.15 278.7 29.85 279.6 ;
        RECT  23.55 282.0 29.85 282.9 ;
        RECT  15.15 297.0 29.85 297.9 ;
        RECT  25.65 293.7 29.85 294.6 ;
        RECT  15.15 308.1 29.85 309.0 ;
        RECT  27.75 311.4 29.85 312.3 ;
        RECT  17.25 326.4 29.85 327.3 ;
        RECT  21.45 323.1 29.85 324.0 ;
        RECT  17.25 337.5 29.85 338.4 ;
        RECT  23.55 340.8 29.85 341.7 ;
        RECT  17.25 355.8 29.85 356.7 ;
        RECT  25.65 352.5 29.85 353.4 ;
        RECT  17.25 366.9 29.85 367.8 ;
        RECT  27.75 370.2 29.85 371.1 ;
        RECT  19.35 385.2 29.85 386.1 ;
        RECT  21.45 381.9 29.85 382.8 ;
        RECT  19.35 396.3 29.85 397.2 ;
        RECT  23.55 399.6 29.85 400.5 ;
        RECT  19.35 414.6 29.85 415.5 ;
        RECT  25.65 411.3 29.85 412.2 ;
        RECT  19.35 425.7 29.85 426.6 ;
        RECT  27.75 429.0 29.85 429.9 ;
        RECT  38.55 88.8 39.45 89.7 ;
        RECT  38.55 104.7 39.45 105.6 ;
        RECT  38.55 118.2 39.45 119.1 ;
        RECT  38.55 134.1 39.45 135.0 ;
        RECT  64.35 88.8 65.25 94.95 ;
        RECT  58.95 94.05 65.25 94.95 ;
        RECT  73.95 88.8 79.05 89.7 ;
        RECT  63.15 96.75 74.85 97.65 ;
        RECT  61.05 82.05 74.85 82.95 ;
        RECT  64.35 99.45 65.25 105.6 ;
        RECT  56.85 99.45 65.25 100.35 ;
        RECT  73.95 104.7 76.95 105.6 ;
        RECT  63.15 96.75 74.85 97.65 ;
        RECT  61.05 111.45 74.85 112.35 ;
        RECT  51.45 91.2 59.85 92.1 ;
        RECT  51.45 87.9 57.75 88.8 ;
        RECT  51.45 102.3 55.65 103.2 ;
        RECT  51.45 105.6 57.75 106.5 ;
        RECT  51.45 120.6 59.85 121.5 ;
        RECT  51.45 117.3 53.55 118.2 ;
        RECT  51.45 131.7 55.65 132.6 ;
        RECT  51.45 131.7 79.05 132.6 ;
        RECT  51.45 135.0 53.55 135.9 ;
        RECT  51.45 135.0 76.95 135.9 ;
        RECT  51.45 82.05 61.95 82.95 ;
        RECT  51.45 96.75 64.05 97.65 ;
        RECT  51.45 111.45 61.95 112.35 ;
        RECT  51.45 126.15 64.05 127.05 ;
        RECT  51.45 140.85 61.95 141.75 ;
        RECT  61.05 138.6 61.95 140.85 ;
        RECT  65.25 82.05 74.85 82.95 ;
        RECT  65.25 67.35 74.85 68.25 ;
        RECT  67.05 68.25 68.25 70.65 ;
        RECT  67.05 80.25 68.25 82.05 ;
        RECT  71.85 81.15 73.05 82.05 ;
        RECT  71.85 68.25 73.05 69.45 ;
        RECT  69.45 70.5 70.65 79.95 ;
        RECT  72.75 75.3 74.85 76.2 ;
        RECT  65.25 75.3 69.45 76.2 ;
        RECT  71.85 78.75 73.05 79.95 ;
        RECT  69.45 78.75 70.65 79.95 ;
        RECT  71.85 69.45 73.05 70.65 ;
        RECT  69.45 69.45 70.65 70.65 ;
        RECT  67.05 69.45 68.25 70.65 ;
        RECT  67.05 79.95 68.25 81.15 ;
        RECT  71.55 75.15 72.75 76.35 ;
        RECT  65.25 111.45 74.85 112.35 ;
        RECT  65.25 126.15 74.85 127.05 ;
        RECT  67.05 123.75 68.25 126.15 ;
        RECT  67.05 112.35 68.25 114.15 ;
        RECT  71.85 112.35 73.05 113.25 ;
        RECT  71.85 124.95 73.05 126.15 ;
        RECT  69.45 114.45 70.65 123.9 ;
        RECT  72.75 118.2 74.85 119.1 ;
        RECT  65.25 118.2 69.45 119.1 ;
        RECT  71.85 116.85 73.05 118.05 ;
        RECT  69.45 116.85 70.65 118.05 ;
        RECT  71.85 117.75 73.05 118.95 ;
        RECT  69.45 117.75 70.65 118.95 ;
        RECT  67.05 122.55 68.25 123.75 ;
        RECT  67.05 112.05 68.25 113.25 ;
        RECT  71.55 116.85 72.75 118.05 ;
        RECT  29.85 82.05 39.45 82.95 ;
        RECT  29.85 67.35 39.45 68.25 ;
        RECT  31.65 68.25 32.85 70.65 ;
        RECT  31.65 80.25 32.85 82.05 ;
        RECT  36.45 81.15 37.65 82.05 ;
        RECT  36.45 68.25 37.65 69.45 ;
        RECT  34.05 70.5 35.25 79.95 ;
        RECT  37.35 75.3 39.45 76.2 ;
        RECT  29.85 75.3 34.05 76.2 ;
        RECT  36.45 78.75 37.65 79.95 ;
        RECT  34.05 78.75 35.25 79.95 ;
        RECT  36.45 69.45 37.65 70.65 ;
        RECT  34.05 69.45 35.25 70.65 ;
        RECT  31.65 69.45 32.85 70.65 ;
        RECT  31.65 79.95 32.85 81.15 ;
        RECT  36.15 75.15 37.35 76.35 ;
        RECT  29.85 111.45 39.45 112.35 ;
        RECT  29.85 126.15 39.45 127.05 ;
        RECT  31.65 123.75 32.85 126.15 ;
        RECT  31.65 112.35 32.85 114.15 ;
        RECT  36.45 112.35 37.65 113.25 ;
        RECT  36.45 124.95 37.65 126.15 ;
        RECT  34.05 114.45 35.25 123.9 ;
        RECT  37.35 118.2 39.45 119.1 ;
        RECT  29.85 118.2 34.05 119.1 ;
        RECT  36.45 116.85 37.65 118.05 ;
        RECT  34.05 116.85 35.25 118.05 ;
        RECT  36.45 117.75 37.65 118.95 ;
        RECT  34.05 117.75 35.25 118.95 ;
        RECT  31.65 122.55 32.85 123.75 ;
        RECT  31.65 112.05 32.85 113.25 ;
        RECT  36.15 116.85 37.35 118.05 ;
        RECT  29.85 111.45 39.45 112.35 ;
        RECT  29.85 96.75 39.45 97.65 ;
        RECT  31.65 97.65 32.85 100.05 ;
        RECT  31.65 109.65 32.85 111.45 ;
        RECT  36.45 110.55 37.65 111.45 ;
        RECT  36.45 97.65 37.65 98.85 ;
        RECT  34.05 99.9 35.25 109.35 ;
        RECT  37.35 104.7 39.45 105.6 ;
        RECT  29.85 104.7 34.05 105.6 ;
        RECT  36.45 108.15 37.65 109.35 ;
        RECT  34.05 108.15 35.25 109.35 ;
        RECT  36.45 98.85 37.65 100.05 ;
        RECT  34.05 98.85 35.25 100.05 ;
        RECT  31.65 98.85 32.85 100.05 ;
        RECT  31.65 109.35 32.85 110.55 ;
        RECT  36.15 104.55 37.35 105.75 ;
        RECT  29.85 140.85 39.45 141.75 ;
        RECT  29.85 155.55 39.45 156.45 ;
        RECT  31.65 153.15 32.85 155.55 ;
        RECT  31.65 141.75 32.85 143.55 ;
        RECT  36.45 141.75 37.65 142.65 ;
        RECT  36.45 154.35 37.65 155.55 ;
        RECT  34.05 143.85 35.25 153.3 ;
        RECT  37.35 147.6 39.45 148.5 ;
        RECT  29.85 147.6 34.05 148.5 ;
        RECT  36.45 146.25 37.65 147.45 ;
        RECT  34.05 146.25 35.25 147.45 ;
        RECT  36.45 147.15 37.65 148.35 ;
        RECT  34.05 147.15 35.25 148.35 ;
        RECT  31.65 151.95 32.85 153.15 ;
        RECT  31.65 141.45 32.85 142.65 ;
        RECT  36.15 146.25 37.35 147.45 ;
        RECT  39.45 82.05 51.45 82.95 ;
        RECT  39.45 67.35 51.45 68.25 ;
        RECT  41.55 67.8 42.45 70.65 ;
        RECT  41.55 80.1 42.45 82.5 ;
        RECT  48.6 67.8 49.5 70.65 ;
        RECT  43.8 67.8 44.7 70.65 ;
        RECT  48.6 79.65 49.5 82.5 ;
        RECT  43.35 72.9 44.25 73.8 ;
        RECT  46.35 72.9 47.25 73.8 ;
        RECT  43.35 73.35 44.25 80.85 ;
        RECT  43.8 72.9 46.8 73.8 ;
        RECT  46.35 70.65 47.25 73.35 ;
        RECT  49.35 72.9 51.45 73.8 ;
        RECT  46.35 76.2 51.45 77.1 ;
        RECT  39.45 75.3 43.8 76.2 ;
        RECT  48.45 78.45 49.65 79.65 ;
        RECT  46.05 78.45 47.25 79.65 ;
        RECT  46.05 78.45 47.25 79.65 ;
        RECT  43.65 78.45 44.85 79.65 ;
        RECT  48.45 69.45 49.65 70.65 ;
        RECT  46.05 69.45 47.25 70.65 ;
        RECT  46.05 69.45 47.25 70.65 ;
        RECT  43.65 69.45 44.85 70.65 ;
        RECT  41.25 69.45 42.45 70.65 ;
        RECT  41.25 79.65 42.45 80.85 ;
        RECT  48.15 72.9 49.35 74.1 ;
        RECT  45.15 76.2 46.35 77.4 ;
        RECT  39.45 111.45 51.45 112.35 ;
        RECT  39.45 126.15 51.45 127.05 ;
        RECT  41.55 123.75 42.45 126.6 ;
        RECT  41.55 111.9 42.45 114.3 ;
        RECT  48.6 123.75 49.5 126.6 ;
        RECT  43.8 123.75 44.7 126.6 ;
        RECT  48.6 111.9 49.5 114.75 ;
        RECT  43.35 120.6 44.25 121.5 ;
        RECT  46.35 120.6 47.25 121.5 ;
        RECT  43.35 113.55 44.25 121.05 ;
        RECT  43.8 120.6 46.8 121.5 ;
        RECT  46.35 121.05 47.25 123.75 ;
        RECT  49.35 120.6 51.45 121.5 ;
        RECT  46.35 117.3 51.45 118.2 ;
        RECT  39.45 118.2 43.8 119.1 ;
        RECT  48.45 118.35 49.65 119.55 ;
        RECT  46.05 118.35 47.25 119.55 ;
        RECT  46.05 118.35 47.25 119.55 ;
        RECT  43.65 118.35 44.85 119.55 ;
        RECT  48.45 117.75 49.65 118.95 ;
        RECT  46.05 117.75 47.25 118.95 ;
        RECT  46.05 117.75 47.25 118.95 ;
        RECT  43.65 117.75 44.85 118.95 ;
        RECT  41.25 122.55 42.45 123.75 ;
        RECT  41.25 112.35 42.45 113.55 ;
        RECT  48.15 119.1 49.35 120.3 ;
        RECT  45.15 115.8 46.35 117.0 ;
        RECT  39.45 111.45 51.45 112.35 ;
        RECT  39.45 96.75 51.45 97.65 ;
        RECT  41.55 97.2 42.45 100.05 ;
        RECT  41.55 109.5 42.45 111.9 ;
        RECT  48.6 97.2 49.5 100.05 ;
        RECT  43.8 97.2 44.7 100.05 ;
        RECT  48.6 109.05 49.5 111.9 ;
        RECT  43.35 102.3 44.25 103.2 ;
        RECT  46.35 102.3 47.25 103.2 ;
        RECT  43.35 102.75 44.25 110.25 ;
        RECT  43.8 102.3 46.8 103.2 ;
        RECT  46.35 100.05 47.25 102.75 ;
        RECT  49.35 102.3 51.45 103.2 ;
        RECT  46.35 105.6 51.45 106.5 ;
        RECT  39.45 104.7 43.8 105.6 ;
        RECT  48.45 107.85 49.65 109.05 ;
        RECT  46.05 107.85 47.25 109.05 ;
        RECT  46.05 107.85 47.25 109.05 ;
        RECT  43.65 107.85 44.85 109.05 ;
        RECT  48.45 98.85 49.65 100.05 ;
        RECT  46.05 98.85 47.25 100.05 ;
        RECT  46.05 98.85 47.25 100.05 ;
        RECT  43.65 98.85 44.85 100.05 ;
        RECT  41.25 98.85 42.45 100.05 ;
        RECT  41.25 109.05 42.45 110.25 ;
        RECT  48.15 102.3 49.35 103.5 ;
        RECT  45.15 105.6 46.35 106.8 ;
        RECT  39.45 140.85 51.45 141.75 ;
        RECT  39.45 155.55 51.45 156.45 ;
        RECT  41.55 153.15 42.45 156.0 ;
        RECT  41.55 141.3 42.45 143.7 ;
        RECT  48.6 153.15 49.5 156.0 ;
        RECT  43.8 153.15 44.7 156.0 ;
        RECT  48.6 141.3 49.5 144.15 ;
        RECT  43.35 150.0 44.25 150.9 ;
        RECT  46.35 150.0 47.25 150.9 ;
        RECT  43.35 142.95 44.25 150.45 ;
        RECT  43.8 150.0 46.8 150.9 ;
        RECT  46.35 150.45 47.25 153.15 ;
        RECT  49.35 150.0 51.45 150.9 ;
        RECT  46.35 146.7 51.45 147.6 ;
        RECT  39.45 147.6 43.8 148.5 ;
        RECT  48.45 147.75 49.65 148.95 ;
        RECT  46.05 147.75 47.25 148.95 ;
        RECT  46.05 147.75 47.25 148.95 ;
        RECT  43.65 147.75 44.85 148.95 ;
        RECT  48.45 147.15 49.65 148.35 ;
        RECT  46.05 147.15 47.25 148.35 ;
        RECT  46.05 147.15 47.25 148.35 ;
        RECT  43.65 147.15 44.85 148.35 ;
        RECT  41.25 151.95 42.45 153.15 ;
        RECT  41.25 141.75 42.45 142.95 ;
        RECT  48.15 148.5 49.35 149.7 ;
        RECT  45.15 145.2 46.35 146.4 ;
        RECT  58.65 92.85 59.85 94.05 ;
        RECT  77.85 87.6 79.05 88.8 ;
        RECT  56.55 98.25 57.75 99.45 ;
        RECT  75.75 103.5 76.95 104.7 ;
        RECT  58.65 90.0 59.85 91.2 ;
        RECT  56.55 86.7 57.75 87.9 ;
        RECT  54.45 101.1 55.65 102.3 ;
        RECT  56.55 104.4 57.75 105.6 ;
        RECT  58.65 119.4 59.85 120.6 ;
        RECT  52.35 116.1 53.55 117.3 ;
        RECT  54.45 130.5 55.65 131.7 ;
        RECT  77.85 130.5 79.05 131.7 ;
        RECT  52.35 133.8 53.55 135.0 ;
        RECT  75.75 133.8 76.95 135.0 ;
        RECT  60.75 80.85 61.95 82.05 ;
        RECT  62.85 95.55 64.05 96.75 ;
        RECT  60.75 110.25 61.95 111.45 ;
        RECT  62.85 124.95 64.05 126.15 ;
        RECT  60.75 137.4 61.95 138.6 ;
        RECT  38.55 147.6 39.45 148.5 ;
        RECT  38.55 163.5 39.45 164.4 ;
        RECT  38.55 177.0 39.45 177.9 ;
        RECT  38.55 192.9 39.45 193.8 ;
        RECT  64.35 147.6 65.25 153.75 ;
        RECT  58.95 152.85 65.25 153.75 ;
        RECT  73.95 147.6 79.05 148.5 ;
        RECT  63.15 155.55 74.85 156.45 ;
        RECT  61.05 140.85 74.85 141.75 ;
        RECT  64.35 158.25 65.25 164.4 ;
        RECT  56.85 158.25 65.25 159.15 ;
        RECT  73.95 163.5 76.95 164.4 ;
        RECT  63.15 155.55 74.85 156.45 ;
        RECT  61.05 170.25 74.85 171.15 ;
        RECT  51.45 150.0 59.85 150.9 ;
        RECT  51.45 146.7 57.75 147.6 ;
        RECT  51.45 161.1 55.65 162.0 ;
        RECT  51.45 164.4 57.75 165.3 ;
        RECT  51.45 179.4 59.85 180.3 ;
        RECT  51.45 176.1 53.55 177.0 ;
        RECT  51.45 190.5 55.65 191.4 ;
        RECT  51.45 190.5 79.05 191.4 ;
        RECT  51.45 193.8 53.55 194.7 ;
        RECT  51.45 193.8 76.95 194.7 ;
        RECT  51.45 140.85 61.95 141.75 ;
        RECT  51.45 155.55 64.05 156.45 ;
        RECT  51.45 170.25 61.95 171.15 ;
        RECT  51.45 184.95 64.05 185.85 ;
        RECT  51.45 199.65 61.95 200.55 ;
        RECT  61.05 197.4 61.95 199.65 ;
        RECT  65.25 140.85 74.85 141.75 ;
        RECT  65.25 126.15 74.85 127.05 ;
        RECT  67.05 127.05 68.25 129.45 ;
        RECT  67.05 139.05 68.25 140.85 ;
        RECT  71.85 139.95 73.05 140.85 ;
        RECT  71.85 127.05 73.05 128.25 ;
        RECT  69.45 129.3 70.65 138.75 ;
        RECT  72.75 134.1 74.85 135.0 ;
        RECT  65.25 134.1 69.45 135.0 ;
        RECT  71.85 137.55 73.05 138.75 ;
        RECT  69.45 137.55 70.65 138.75 ;
        RECT  71.85 128.25 73.05 129.45 ;
        RECT  69.45 128.25 70.65 129.45 ;
        RECT  67.05 128.25 68.25 129.45 ;
        RECT  67.05 138.75 68.25 139.95 ;
        RECT  71.55 133.95 72.75 135.15 ;
        RECT  65.25 170.25 74.85 171.15 ;
        RECT  65.25 184.95 74.85 185.85 ;
        RECT  67.05 182.55 68.25 184.95 ;
        RECT  67.05 171.15 68.25 172.95 ;
        RECT  71.85 171.15 73.05 172.05 ;
        RECT  71.85 183.75 73.05 184.95 ;
        RECT  69.45 173.25 70.65 182.7 ;
        RECT  72.75 177.0 74.85 177.9 ;
        RECT  65.25 177.0 69.45 177.9 ;
        RECT  71.85 175.65 73.05 176.85 ;
        RECT  69.45 175.65 70.65 176.85 ;
        RECT  71.85 176.55 73.05 177.75 ;
        RECT  69.45 176.55 70.65 177.75 ;
        RECT  67.05 181.35 68.25 182.55 ;
        RECT  67.05 170.85 68.25 172.05 ;
        RECT  71.55 175.65 72.75 176.85 ;
        RECT  29.85 140.85 39.45 141.75 ;
        RECT  29.85 126.15 39.45 127.05 ;
        RECT  31.65 127.05 32.85 129.45 ;
        RECT  31.65 139.05 32.85 140.85 ;
        RECT  36.45 139.95 37.65 140.85 ;
        RECT  36.45 127.05 37.65 128.25 ;
        RECT  34.05 129.3 35.25 138.75 ;
        RECT  37.35 134.1 39.45 135.0 ;
        RECT  29.85 134.1 34.05 135.0 ;
        RECT  36.45 137.55 37.65 138.75 ;
        RECT  34.05 137.55 35.25 138.75 ;
        RECT  36.45 128.25 37.65 129.45 ;
        RECT  34.05 128.25 35.25 129.45 ;
        RECT  31.65 128.25 32.85 129.45 ;
        RECT  31.65 138.75 32.85 139.95 ;
        RECT  36.15 133.95 37.35 135.15 ;
        RECT  29.85 170.25 39.45 171.15 ;
        RECT  29.85 184.95 39.45 185.85 ;
        RECT  31.65 182.55 32.85 184.95 ;
        RECT  31.65 171.15 32.85 172.95 ;
        RECT  36.45 171.15 37.65 172.05 ;
        RECT  36.45 183.75 37.65 184.95 ;
        RECT  34.05 173.25 35.25 182.7 ;
        RECT  37.35 177.0 39.45 177.9 ;
        RECT  29.85 177.0 34.05 177.9 ;
        RECT  36.45 175.65 37.65 176.85 ;
        RECT  34.05 175.65 35.25 176.85 ;
        RECT  36.45 176.55 37.65 177.75 ;
        RECT  34.05 176.55 35.25 177.75 ;
        RECT  31.65 181.35 32.85 182.55 ;
        RECT  31.65 170.85 32.85 172.05 ;
        RECT  36.15 175.65 37.35 176.85 ;
        RECT  29.85 170.25 39.45 171.15 ;
        RECT  29.85 155.55 39.45 156.45 ;
        RECT  31.65 156.45 32.85 158.85 ;
        RECT  31.65 168.45 32.85 170.25 ;
        RECT  36.45 169.35 37.65 170.25 ;
        RECT  36.45 156.45 37.65 157.65 ;
        RECT  34.05 158.7 35.25 168.15 ;
        RECT  37.35 163.5 39.45 164.4 ;
        RECT  29.85 163.5 34.05 164.4 ;
        RECT  36.45 166.95 37.65 168.15 ;
        RECT  34.05 166.95 35.25 168.15 ;
        RECT  36.45 157.65 37.65 158.85 ;
        RECT  34.05 157.65 35.25 158.85 ;
        RECT  31.65 157.65 32.85 158.85 ;
        RECT  31.65 168.15 32.85 169.35 ;
        RECT  36.15 163.35 37.35 164.55 ;
        RECT  29.85 199.65 39.45 200.55 ;
        RECT  29.85 214.35 39.45 215.25 ;
        RECT  31.65 211.95 32.85 214.35 ;
        RECT  31.65 200.55 32.85 202.35 ;
        RECT  36.45 200.55 37.65 201.45 ;
        RECT  36.45 213.15 37.65 214.35 ;
        RECT  34.05 202.65 35.25 212.1 ;
        RECT  37.35 206.4 39.45 207.3 ;
        RECT  29.85 206.4 34.05 207.3 ;
        RECT  36.45 205.05 37.65 206.25 ;
        RECT  34.05 205.05 35.25 206.25 ;
        RECT  36.45 205.95 37.65 207.15 ;
        RECT  34.05 205.95 35.25 207.15 ;
        RECT  31.65 210.75 32.85 211.95 ;
        RECT  31.65 200.25 32.85 201.45 ;
        RECT  36.15 205.05 37.35 206.25 ;
        RECT  39.45 140.85 51.45 141.75 ;
        RECT  39.45 126.15 51.45 127.05 ;
        RECT  41.55 126.6 42.45 129.45 ;
        RECT  41.55 138.9 42.45 141.3 ;
        RECT  48.6 126.6 49.5 129.45 ;
        RECT  43.8 126.6 44.7 129.45 ;
        RECT  48.6 138.45 49.5 141.3 ;
        RECT  43.35 131.7 44.25 132.6 ;
        RECT  46.35 131.7 47.25 132.6 ;
        RECT  43.35 132.15 44.25 139.65 ;
        RECT  43.8 131.7 46.8 132.6 ;
        RECT  46.35 129.45 47.25 132.15 ;
        RECT  49.35 131.7 51.45 132.6 ;
        RECT  46.35 135.0 51.45 135.9 ;
        RECT  39.45 134.1 43.8 135.0 ;
        RECT  48.45 137.25 49.65 138.45 ;
        RECT  46.05 137.25 47.25 138.45 ;
        RECT  46.05 137.25 47.25 138.45 ;
        RECT  43.65 137.25 44.85 138.45 ;
        RECT  48.45 128.25 49.65 129.45 ;
        RECT  46.05 128.25 47.25 129.45 ;
        RECT  46.05 128.25 47.25 129.45 ;
        RECT  43.65 128.25 44.85 129.45 ;
        RECT  41.25 128.25 42.45 129.45 ;
        RECT  41.25 138.45 42.45 139.65 ;
        RECT  48.15 131.7 49.35 132.9 ;
        RECT  45.15 135.0 46.35 136.2 ;
        RECT  39.45 170.25 51.45 171.15 ;
        RECT  39.45 184.95 51.45 185.85 ;
        RECT  41.55 182.55 42.45 185.4 ;
        RECT  41.55 170.7 42.45 173.1 ;
        RECT  48.6 182.55 49.5 185.4 ;
        RECT  43.8 182.55 44.7 185.4 ;
        RECT  48.6 170.7 49.5 173.55 ;
        RECT  43.35 179.4 44.25 180.3 ;
        RECT  46.35 179.4 47.25 180.3 ;
        RECT  43.35 172.35 44.25 179.85 ;
        RECT  43.8 179.4 46.8 180.3 ;
        RECT  46.35 179.85 47.25 182.55 ;
        RECT  49.35 179.4 51.45 180.3 ;
        RECT  46.35 176.1 51.45 177.0 ;
        RECT  39.45 177.0 43.8 177.9 ;
        RECT  48.45 177.15 49.65 178.35 ;
        RECT  46.05 177.15 47.25 178.35 ;
        RECT  46.05 177.15 47.25 178.35 ;
        RECT  43.65 177.15 44.85 178.35 ;
        RECT  48.45 176.55 49.65 177.75 ;
        RECT  46.05 176.55 47.25 177.75 ;
        RECT  46.05 176.55 47.25 177.75 ;
        RECT  43.65 176.55 44.85 177.75 ;
        RECT  41.25 181.35 42.45 182.55 ;
        RECT  41.25 171.15 42.45 172.35 ;
        RECT  48.15 177.9 49.35 179.1 ;
        RECT  45.15 174.6 46.35 175.8 ;
        RECT  39.45 170.25 51.45 171.15 ;
        RECT  39.45 155.55 51.45 156.45 ;
        RECT  41.55 156.0 42.45 158.85 ;
        RECT  41.55 168.3 42.45 170.7 ;
        RECT  48.6 156.0 49.5 158.85 ;
        RECT  43.8 156.0 44.7 158.85 ;
        RECT  48.6 167.85 49.5 170.7 ;
        RECT  43.35 161.1 44.25 162.0 ;
        RECT  46.35 161.1 47.25 162.0 ;
        RECT  43.35 161.55 44.25 169.05 ;
        RECT  43.8 161.1 46.8 162.0 ;
        RECT  46.35 158.85 47.25 161.55 ;
        RECT  49.35 161.1 51.45 162.0 ;
        RECT  46.35 164.4 51.45 165.3 ;
        RECT  39.45 163.5 43.8 164.4 ;
        RECT  48.45 166.65 49.65 167.85 ;
        RECT  46.05 166.65 47.25 167.85 ;
        RECT  46.05 166.65 47.25 167.85 ;
        RECT  43.65 166.65 44.85 167.85 ;
        RECT  48.45 157.65 49.65 158.85 ;
        RECT  46.05 157.65 47.25 158.85 ;
        RECT  46.05 157.65 47.25 158.85 ;
        RECT  43.65 157.65 44.85 158.85 ;
        RECT  41.25 157.65 42.45 158.85 ;
        RECT  41.25 167.85 42.45 169.05 ;
        RECT  48.15 161.1 49.35 162.3 ;
        RECT  45.15 164.4 46.35 165.6 ;
        RECT  39.45 199.65 51.45 200.55 ;
        RECT  39.45 214.35 51.45 215.25 ;
        RECT  41.55 211.95 42.45 214.8 ;
        RECT  41.55 200.1 42.45 202.5 ;
        RECT  48.6 211.95 49.5 214.8 ;
        RECT  43.8 211.95 44.7 214.8 ;
        RECT  48.6 200.1 49.5 202.95 ;
        RECT  43.35 208.8 44.25 209.7 ;
        RECT  46.35 208.8 47.25 209.7 ;
        RECT  43.35 201.75 44.25 209.25 ;
        RECT  43.8 208.8 46.8 209.7 ;
        RECT  46.35 209.25 47.25 211.95 ;
        RECT  49.35 208.8 51.45 209.7 ;
        RECT  46.35 205.5 51.45 206.4 ;
        RECT  39.45 206.4 43.8 207.3 ;
        RECT  48.45 206.55 49.65 207.75 ;
        RECT  46.05 206.55 47.25 207.75 ;
        RECT  46.05 206.55 47.25 207.75 ;
        RECT  43.65 206.55 44.85 207.75 ;
        RECT  48.45 205.95 49.65 207.15 ;
        RECT  46.05 205.95 47.25 207.15 ;
        RECT  46.05 205.95 47.25 207.15 ;
        RECT  43.65 205.95 44.85 207.15 ;
        RECT  41.25 210.75 42.45 211.95 ;
        RECT  41.25 200.55 42.45 201.75 ;
        RECT  48.15 207.3 49.35 208.5 ;
        RECT  45.15 204.0 46.35 205.2 ;
        RECT  58.65 151.65 59.85 152.85 ;
        RECT  77.85 146.4 79.05 147.6 ;
        RECT  56.55 157.05 57.75 158.25 ;
        RECT  75.75 162.3 76.95 163.5 ;
        RECT  58.65 148.8 59.85 150.0 ;
        RECT  56.55 145.5 57.75 146.7 ;
        RECT  54.45 159.9 55.65 161.1 ;
        RECT  56.55 163.2 57.75 164.4 ;
        RECT  58.65 178.2 59.85 179.4 ;
        RECT  52.35 174.9 53.55 176.1 ;
        RECT  54.45 189.3 55.65 190.5 ;
        RECT  77.85 189.3 79.05 190.5 ;
        RECT  52.35 192.6 53.55 193.8 ;
        RECT  75.75 192.6 76.95 193.8 ;
        RECT  60.75 139.65 61.95 140.85 ;
        RECT  62.85 154.35 64.05 155.55 ;
        RECT  60.75 169.05 61.95 170.25 ;
        RECT  62.85 183.75 64.05 184.95 ;
        RECT  60.75 196.2 61.95 197.4 ;
        RECT  29.85 199.65 41.85 200.55 ;
        RECT  29.85 214.35 41.85 215.25 ;
        RECT  38.85 211.95 39.75 214.8 ;
        RECT  38.85 200.1 39.75 202.5 ;
        RECT  31.8 211.95 32.7 214.8 ;
        RECT  36.6 211.95 37.5 214.8 ;
        RECT  31.8 200.1 32.7 202.95 ;
        RECT  37.05 208.8 37.95 209.7 ;
        RECT  34.05 208.8 34.95 209.7 ;
        RECT  37.05 201.75 37.95 209.25 ;
        RECT  34.5 208.8 37.5 209.7 ;
        RECT  34.05 209.25 34.95 211.95 ;
        RECT  29.85 208.8 31.95 209.7 ;
        RECT  29.85 205.5 34.95 206.4 ;
        RECT  37.5 206.4 41.85 207.3 ;
        RECT  31.65 202.95 32.85 204.15 ;
        RECT  34.05 202.95 35.25 204.15 ;
        RECT  34.05 202.95 35.25 204.15 ;
        RECT  36.45 202.95 37.65 204.15 ;
        RECT  31.65 211.95 32.85 213.15 ;
        RECT  34.05 211.95 35.25 213.15 ;
        RECT  34.05 211.95 35.25 213.15 ;
        RECT  36.45 211.95 37.65 213.15 ;
        RECT  38.85 211.95 40.05 213.15 ;
        RECT  38.85 201.75 40.05 202.95 ;
        RECT  31.95 208.5 33.15 209.7 ;
        RECT  34.95 205.2 36.15 206.4 ;
        RECT  29.85 229.05 41.85 229.95 ;
        RECT  29.85 214.35 41.85 215.25 ;
        RECT  38.85 214.8 39.75 217.65 ;
        RECT  38.85 227.1 39.75 229.5 ;
        RECT  31.8 214.8 32.7 217.65 ;
        RECT  36.6 214.8 37.5 217.65 ;
        RECT  31.8 226.65 32.7 229.5 ;
        RECT  37.05 219.9 37.95 220.8 ;
        RECT  34.05 219.9 34.95 220.8 ;
        RECT  37.05 220.35 37.95 227.85 ;
        RECT  34.5 219.9 37.5 220.8 ;
        RECT  34.05 217.65 34.95 220.35 ;
        RECT  29.85 219.9 31.95 220.8 ;
        RECT  29.85 223.2 34.95 224.1 ;
        RECT  37.5 222.3 41.85 223.2 ;
        RECT  31.65 221.85 32.85 223.05 ;
        RECT  34.05 221.85 35.25 223.05 ;
        RECT  34.05 221.85 35.25 223.05 ;
        RECT  36.45 221.85 37.65 223.05 ;
        RECT  31.65 222.45 32.85 223.65 ;
        RECT  34.05 222.45 35.25 223.65 ;
        RECT  34.05 222.45 35.25 223.65 ;
        RECT  36.45 222.45 37.65 223.65 ;
        RECT  38.85 217.65 40.05 218.85 ;
        RECT  38.85 227.85 40.05 229.05 ;
        RECT  31.95 221.1 33.15 222.3 ;
        RECT  34.95 224.4 36.15 225.6 ;
        RECT  29.85 229.05 41.85 229.95 ;
        RECT  29.85 243.75 41.85 244.65 ;
        RECT  38.85 241.35 39.75 244.2 ;
        RECT  38.85 229.5 39.75 231.9 ;
        RECT  31.8 241.35 32.7 244.2 ;
        RECT  36.6 241.35 37.5 244.2 ;
        RECT  31.8 229.5 32.7 232.35 ;
        RECT  37.05 238.2 37.95 239.1 ;
        RECT  34.05 238.2 34.95 239.1 ;
        RECT  37.05 231.15 37.95 238.65 ;
        RECT  34.5 238.2 37.5 239.1 ;
        RECT  34.05 238.65 34.95 241.35 ;
        RECT  29.85 238.2 31.95 239.1 ;
        RECT  29.85 234.9 34.95 235.8 ;
        RECT  37.5 235.8 41.85 236.7 ;
        RECT  31.65 232.35 32.85 233.55 ;
        RECT  34.05 232.35 35.25 233.55 ;
        RECT  34.05 232.35 35.25 233.55 ;
        RECT  36.45 232.35 37.65 233.55 ;
        RECT  31.65 241.35 32.85 242.55 ;
        RECT  34.05 241.35 35.25 242.55 ;
        RECT  34.05 241.35 35.25 242.55 ;
        RECT  36.45 241.35 37.65 242.55 ;
        RECT  38.85 241.35 40.05 242.55 ;
        RECT  38.85 231.15 40.05 232.35 ;
        RECT  31.95 237.9 33.15 239.1 ;
        RECT  34.95 234.6 36.15 235.8 ;
        RECT  29.85 258.45 41.85 259.35 ;
        RECT  29.85 243.75 41.85 244.65 ;
        RECT  38.85 244.2 39.75 247.05 ;
        RECT  38.85 256.5 39.75 258.9 ;
        RECT  31.8 244.2 32.7 247.05 ;
        RECT  36.6 244.2 37.5 247.05 ;
        RECT  31.8 256.05 32.7 258.9 ;
        RECT  37.05 249.3 37.95 250.2 ;
        RECT  34.05 249.3 34.95 250.2 ;
        RECT  37.05 249.75 37.95 257.25 ;
        RECT  34.5 249.3 37.5 250.2 ;
        RECT  34.05 247.05 34.95 249.75 ;
        RECT  29.85 249.3 31.95 250.2 ;
        RECT  29.85 252.6 34.95 253.5 ;
        RECT  37.5 251.7 41.85 252.6 ;
        RECT  31.65 251.25 32.85 252.45 ;
        RECT  34.05 251.25 35.25 252.45 ;
        RECT  34.05 251.25 35.25 252.45 ;
        RECT  36.45 251.25 37.65 252.45 ;
        RECT  31.65 251.85 32.85 253.05 ;
        RECT  34.05 251.85 35.25 253.05 ;
        RECT  34.05 251.85 35.25 253.05 ;
        RECT  36.45 251.85 37.65 253.05 ;
        RECT  38.85 247.05 40.05 248.25 ;
        RECT  38.85 257.25 40.05 258.45 ;
        RECT  31.95 250.5 33.15 251.7 ;
        RECT  34.95 253.8 36.15 255.0 ;
        RECT  29.85 258.45 41.85 259.35 ;
        RECT  29.85 273.15 41.85 274.05 ;
        RECT  38.85 270.75 39.75 273.6 ;
        RECT  38.85 258.9 39.75 261.3 ;
        RECT  31.8 270.75 32.7 273.6 ;
        RECT  36.6 270.75 37.5 273.6 ;
        RECT  31.8 258.9 32.7 261.75 ;
        RECT  37.05 267.6 37.95 268.5 ;
        RECT  34.05 267.6 34.95 268.5 ;
        RECT  37.05 260.55 37.95 268.05 ;
        RECT  34.5 267.6 37.5 268.5 ;
        RECT  34.05 268.05 34.95 270.75 ;
        RECT  29.85 267.6 31.95 268.5 ;
        RECT  29.85 264.3 34.95 265.2 ;
        RECT  37.5 265.2 41.85 266.1 ;
        RECT  31.65 261.75 32.85 262.95 ;
        RECT  34.05 261.75 35.25 262.95 ;
        RECT  34.05 261.75 35.25 262.95 ;
        RECT  36.45 261.75 37.65 262.95 ;
        RECT  31.65 270.75 32.85 271.95 ;
        RECT  34.05 270.75 35.25 271.95 ;
        RECT  34.05 270.75 35.25 271.95 ;
        RECT  36.45 270.75 37.65 271.95 ;
        RECT  38.85 270.75 40.05 271.95 ;
        RECT  38.85 260.55 40.05 261.75 ;
        RECT  31.95 267.3 33.15 268.5 ;
        RECT  34.95 264.0 36.15 265.2 ;
        RECT  29.85 287.85 41.85 288.75 ;
        RECT  29.85 273.15 41.85 274.05 ;
        RECT  38.85 273.6 39.75 276.45 ;
        RECT  38.85 285.9 39.75 288.3 ;
        RECT  31.8 273.6 32.7 276.45 ;
        RECT  36.6 273.6 37.5 276.45 ;
        RECT  31.8 285.45 32.7 288.3 ;
        RECT  37.05 278.7 37.95 279.6 ;
        RECT  34.05 278.7 34.95 279.6 ;
        RECT  37.05 279.15 37.95 286.65 ;
        RECT  34.5 278.7 37.5 279.6 ;
        RECT  34.05 276.45 34.95 279.15 ;
        RECT  29.85 278.7 31.95 279.6 ;
        RECT  29.85 282.0 34.95 282.9 ;
        RECT  37.5 281.1 41.85 282.0 ;
        RECT  31.65 280.65 32.85 281.85 ;
        RECT  34.05 280.65 35.25 281.85 ;
        RECT  34.05 280.65 35.25 281.85 ;
        RECT  36.45 280.65 37.65 281.85 ;
        RECT  31.65 281.25 32.85 282.45 ;
        RECT  34.05 281.25 35.25 282.45 ;
        RECT  34.05 281.25 35.25 282.45 ;
        RECT  36.45 281.25 37.65 282.45 ;
        RECT  38.85 276.45 40.05 277.65 ;
        RECT  38.85 286.65 40.05 287.85 ;
        RECT  31.95 279.9 33.15 281.1 ;
        RECT  34.95 283.2 36.15 284.4 ;
        RECT  29.85 287.85 41.85 288.75 ;
        RECT  29.85 302.55 41.85 303.45 ;
        RECT  38.85 300.15 39.75 303.0 ;
        RECT  38.85 288.3 39.75 290.7 ;
        RECT  31.8 300.15 32.7 303.0 ;
        RECT  36.6 300.15 37.5 303.0 ;
        RECT  31.8 288.3 32.7 291.15 ;
        RECT  37.05 297.0 37.95 297.9 ;
        RECT  34.05 297.0 34.95 297.9 ;
        RECT  37.05 289.95 37.95 297.45 ;
        RECT  34.5 297.0 37.5 297.9 ;
        RECT  34.05 297.45 34.95 300.15 ;
        RECT  29.85 297.0 31.95 297.9 ;
        RECT  29.85 293.7 34.95 294.6 ;
        RECT  37.5 294.6 41.85 295.5 ;
        RECT  31.65 291.15 32.85 292.35 ;
        RECT  34.05 291.15 35.25 292.35 ;
        RECT  34.05 291.15 35.25 292.35 ;
        RECT  36.45 291.15 37.65 292.35 ;
        RECT  31.65 300.15 32.85 301.35 ;
        RECT  34.05 300.15 35.25 301.35 ;
        RECT  34.05 300.15 35.25 301.35 ;
        RECT  36.45 300.15 37.65 301.35 ;
        RECT  38.85 300.15 40.05 301.35 ;
        RECT  38.85 289.95 40.05 291.15 ;
        RECT  31.95 296.7 33.15 297.9 ;
        RECT  34.95 293.4 36.15 294.6 ;
        RECT  29.85 317.25 41.85 318.15 ;
        RECT  29.85 302.55 41.85 303.45 ;
        RECT  38.85 303.0 39.75 305.85 ;
        RECT  38.85 315.3 39.75 317.7 ;
        RECT  31.8 303.0 32.7 305.85 ;
        RECT  36.6 303.0 37.5 305.85 ;
        RECT  31.8 314.85 32.7 317.7 ;
        RECT  37.05 308.1 37.95 309.0 ;
        RECT  34.05 308.1 34.95 309.0 ;
        RECT  37.05 308.55 37.95 316.05 ;
        RECT  34.5 308.1 37.5 309.0 ;
        RECT  34.05 305.85 34.95 308.55 ;
        RECT  29.85 308.1 31.95 309.0 ;
        RECT  29.85 311.4 34.95 312.3 ;
        RECT  37.5 310.5 41.85 311.4 ;
        RECT  31.65 310.05 32.85 311.25 ;
        RECT  34.05 310.05 35.25 311.25 ;
        RECT  34.05 310.05 35.25 311.25 ;
        RECT  36.45 310.05 37.65 311.25 ;
        RECT  31.65 310.65 32.85 311.85 ;
        RECT  34.05 310.65 35.25 311.85 ;
        RECT  34.05 310.65 35.25 311.85 ;
        RECT  36.45 310.65 37.65 311.85 ;
        RECT  38.85 305.85 40.05 307.05 ;
        RECT  38.85 316.05 40.05 317.25 ;
        RECT  31.95 309.3 33.15 310.5 ;
        RECT  34.95 312.6 36.15 313.8 ;
        RECT  29.85 317.25 41.85 318.15 ;
        RECT  29.85 331.95 41.85 332.85 ;
        RECT  38.85 329.55 39.75 332.4 ;
        RECT  38.85 317.7 39.75 320.1 ;
        RECT  31.8 329.55 32.7 332.4 ;
        RECT  36.6 329.55 37.5 332.4 ;
        RECT  31.8 317.7 32.7 320.55 ;
        RECT  37.05 326.4 37.95 327.3 ;
        RECT  34.05 326.4 34.95 327.3 ;
        RECT  37.05 319.35 37.95 326.85 ;
        RECT  34.5 326.4 37.5 327.3 ;
        RECT  34.05 326.85 34.95 329.55 ;
        RECT  29.85 326.4 31.95 327.3 ;
        RECT  29.85 323.1 34.95 324.0 ;
        RECT  37.5 324.0 41.85 324.9 ;
        RECT  31.65 320.55 32.85 321.75 ;
        RECT  34.05 320.55 35.25 321.75 ;
        RECT  34.05 320.55 35.25 321.75 ;
        RECT  36.45 320.55 37.65 321.75 ;
        RECT  31.65 329.55 32.85 330.75 ;
        RECT  34.05 329.55 35.25 330.75 ;
        RECT  34.05 329.55 35.25 330.75 ;
        RECT  36.45 329.55 37.65 330.75 ;
        RECT  38.85 329.55 40.05 330.75 ;
        RECT  38.85 319.35 40.05 320.55 ;
        RECT  31.95 326.1 33.15 327.3 ;
        RECT  34.95 322.8 36.15 324.0 ;
        RECT  29.85 346.65 41.85 347.55 ;
        RECT  29.85 331.95 41.85 332.85 ;
        RECT  38.85 332.4 39.75 335.25 ;
        RECT  38.85 344.7 39.75 347.1 ;
        RECT  31.8 332.4 32.7 335.25 ;
        RECT  36.6 332.4 37.5 335.25 ;
        RECT  31.8 344.25 32.7 347.1 ;
        RECT  37.05 337.5 37.95 338.4 ;
        RECT  34.05 337.5 34.95 338.4 ;
        RECT  37.05 337.95 37.95 345.45 ;
        RECT  34.5 337.5 37.5 338.4 ;
        RECT  34.05 335.25 34.95 337.95 ;
        RECT  29.85 337.5 31.95 338.4 ;
        RECT  29.85 340.8 34.95 341.7 ;
        RECT  37.5 339.9 41.85 340.8 ;
        RECT  31.65 339.45 32.85 340.65 ;
        RECT  34.05 339.45 35.25 340.65 ;
        RECT  34.05 339.45 35.25 340.65 ;
        RECT  36.45 339.45 37.65 340.65 ;
        RECT  31.65 340.05 32.85 341.25 ;
        RECT  34.05 340.05 35.25 341.25 ;
        RECT  34.05 340.05 35.25 341.25 ;
        RECT  36.45 340.05 37.65 341.25 ;
        RECT  38.85 335.25 40.05 336.45 ;
        RECT  38.85 345.45 40.05 346.65 ;
        RECT  31.95 338.7 33.15 339.9 ;
        RECT  34.95 342.0 36.15 343.2 ;
        RECT  29.85 346.65 41.85 347.55 ;
        RECT  29.85 361.35 41.85 362.25 ;
        RECT  38.85 358.95 39.75 361.8 ;
        RECT  38.85 347.1 39.75 349.5 ;
        RECT  31.8 358.95 32.7 361.8 ;
        RECT  36.6 358.95 37.5 361.8 ;
        RECT  31.8 347.1 32.7 349.95 ;
        RECT  37.05 355.8 37.95 356.7 ;
        RECT  34.05 355.8 34.95 356.7 ;
        RECT  37.05 348.75 37.95 356.25 ;
        RECT  34.5 355.8 37.5 356.7 ;
        RECT  34.05 356.25 34.95 358.95 ;
        RECT  29.85 355.8 31.95 356.7 ;
        RECT  29.85 352.5 34.95 353.4 ;
        RECT  37.5 353.4 41.85 354.3 ;
        RECT  31.65 349.95 32.85 351.15 ;
        RECT  34.05 349.95 35.25 351.15 ;
        RECT  34.05 349.95 35.25 351.15 ;
        RECT  36.45 349.95 37.65 351.15 ;
        RECT  31.65 358.95 32.85 360.15 ;
        RECT  34.05 358.95 35.25 360.15 ;
        RECT  34.05 358.95 35.25 360.15 ;
        RECT  36.45 358.95 37.65 360.15 ;
        RECT  38.85 358.95 40.05 360.15 ;
        RECT  38.85 348.75 40.05 349.95 ;
        RECT  31.95 355.5 33.15 356.7 ;
        RECT  34.95 352.2 36.15 353.4 ;
        RECT  29.85 376.05 41.85 376.95 ;
        RECT  29.85 361.35 41.85 362.25 ;
        RECT  38.85 361.8 39.75 364.65 ;
        RECT  38.85 374.1 39.75 376.5 ;
        RECT  31.8 361.8 32.7 364.65 ;
        RECT  36.6 361.8 37.5 364.65 ;
        RECT  31.8 373.65 32.7 376.5 ;
        RECT  37.05 366.9 37.95 367.8 ;
        RECT  34.05 366.9 34.95 367.8 ;
        RECT  37.05 367.35 37.95 374.85 ;
        RECT  34.5 366.9 37.5 367.8 ;
        RECT  34.05 364.65 34.95 367.35 ;
        RECT  29.85 366.9 31.95 367.8 ;
        RECT  29.85 370.2 34.95 371.1 ;
        RECT  37.5 369.3 41.85 370.2 ;
        RECT  31.65 368.85 32.85 370.05 ;
        RECT  34.05 368.85 35.25 370.05 ;
        RECT  34.05 368.85 35.25 370.05 ;
        RECT  36.45 368.85 37.65 370.05 ;
        RECT  31.65 369.45 32.85 370.65 ;
        RECT  34.05 369.45 35.25 370.65 ;
        RECT  34.05 369.45 35.25 370.65 ;
        RECT  36.45 369.45 37.65 370.65 ;
        RECT  38.85 364.65 40.05 365.85 ;
        RECT  38.85 374.85 40.05 376.05 ;
        RECT  31.95 368.1 33.15 369.3 ;
        RECT  34.95 371.4 36.15 372.6 ;
        RECT  29.85 376.05 41.85 376.95 ;
        RECT  29.85 390.75 41.85 391.65 ;
        RECT  38.85 388.35 39.75 391.2 ;
        RECT  38.85 376.5 39.75 378.9 ;
        RECT  31.8 388.35 32.7 391.2 ;
        RECT  36.6 388.35 37.5 391.2 ;
        RECT  31.8 376.5 32.7 379.35 ;
        RECT  37.05 385.2 37.95 386.1 ;
        RECT  34.05 385.2 34.95 386.1 ;
        RECT  37.05 378.15 37.95 385.65 ;
        RECT  34.5 385.2 37.5 386.1 ;
        RECT  34.05 385.65 34.95 388.35 ;
        RECT  29.85 385.2 31.95 386.1 ;
        RECT  29.85 381.9 34.95 382.8 ;
        RECT  37.5 382.8 41.85 383.7 ;
        RECT  31.65 379.35 32.85 380.55 ;
        RECT  34.05 379.35 35.25 380.55 ;
        RECT  34.05 379.35 35.25 380.55 ;
        RECT  36.45 379.35 37.65 380.55 ;
        RECT  31.65 388.35 32.85 389.55 ;
        RECT  34.05 388.35 35.25 389.55 ;
        RECT  34.05 388.35 35.25 389.55 ;
        RECT  36.45 388.35 37.65 389.55 ;
        RECT  38.85 388.35 40.05 389.55 ;
        RECT  38.85 378.15 40.05 379.35 ;
        RECT  31.95 384.9 33.15 386.1 ;
        RECT  34.95 381.6 36.15 382.8 ;
        RECT  29.85 405.45 41.85 406.35 ;
        RECT  29.85 390.75 41.85 391.65 ;
        RECT  38.85 391.2 39.75 394.05 ;
        RECT  38.85 403.5 39.75 405.9 ;
        RECT  31.8 391.2 32.7 394.05 ;
        RECT  36.6 391.2 37.5 394.05 ;
        RECT  31.8 403.05 32.7 405.9 ;
        RECT  37.05 396.3 37.95 397.2 ;
        RECT  34.05 396.3 34.95 397.2 ;
        RECT  37.05 396.75 37.95 404.25 ;
        RECT  34.5 396.3 37.5 397.2 ;
        RECT  34.05 394.05 34.95 396.75 ;
        RECT  29.85 396.3 31.95 397.2 ;
        RECT  29.85 399.6 34.95 400.5 ;
        RECT  37.5 398.7 41.85 399.6 ;
        RECT  31.65 398.25 32.85 399.45 ;
        RECT  34.05 398.25 35.25 399.45 ;
        RECT  34.05 398.25 35.25 399.45 ;
        RECT  36.45 398.25 37.65 399.45 ;
        RECT  31.65 398.85 32.85 400.05 ;
        RECT  34.05 398.85 35.25 400.05 ;
        RECT  34.05 398.85 35.25 400.05 ;
        RECT  36.45 398.85 37.65 400.05 ;
        RECT  38.85 394.05 40.05 395.25 ;
        RECT  38.85 404.25 40.05 405.45 ;
        RECT  31.95 397.5 33.15 398.7 ;
        RECT  34.95 400.8 36.15 402.0 ;
        RECT  29.85 405.45 41.85 406.35 ;
        RECT  29.85 420.15 41.85 421.05 ;
        RECT  38.85 417.75 39.75 420.6 ;
        RECT  38.85 405.9 39.75 408.3 ;
        RECT  31.8 417.75 32.7 420.6 ;
        RECT  36.6 417.75 37.5 420.6 ;
        RECT  31.8 405.9 32.7 408.75 ;
        RECT  37.05 414.6 37.95 415.5 ;
        RECT  34.05 414.6 34.95 415.5 ;
        RECT  37.05 407.55 37.95 415.05 ;
        RECT  34.5 414.6 37.5 415.5 ;
        RECT  34.05 415.05 34.95 417.75 ;
        RECT  29.85 414.6 31.95 415.5 ;
        RECT  29.85 411.3 34.95 412.2 ;
        RECT  37.5 412.2 41.85 413.1 ;
        RECT  31.65 408.75 32.85 409.95 ;
        RECT  34.05 408.75 35.25 409.95 ;
        RECT  34.05 408.75 35.25 409.95 ;
        RECT  36.45 408.75 37.65 409.95 ;
        RECT  31.65 417.75 32.85 418.95 ;
        RECT  34.05 417.75 35.25 418.95 ;
        RECT  34.05 417.75 35.25 418.95 ;
        RECT  36.45 417.75 37.65 418.95 ;
        RECT  38.85 417.75 40.05 418.95 ;
        RECT  38.85 407.55 40.05 408.75 ;
        RECT  31.95 414.3 33.15 415.5 ;
        RECT  34.95 411.0 36.15 412.2 ;
        RECT  29.85 434.85 41.85 435.75 ;
        RECT  29.85 420.15 41.85 421.05 ;
        RECT  38.85 420.6 39.75 423.45 ;
        RECT  38.85 432.9 39.75 435.3 ;
        RECT  31.8 420.6 32.7 423.45 ;
        RECT  36.6 420.6 37.5 423.45 ;
        RECT  31.8 432.45 32.7 435.3 ;
        RECT  37.05 425.7 37.95 426.6 ;
        RECT  34.05 425.7 34.95 426.6 ;
        RECT  37.05 426.15 37.95 433.65 ;
        RECT  34.5 425.7 37.5 426.6 ;
        RECT  34.05 423.45 34.95 426.15 ;
        RECT  29.85 425.7 31.95 426.6 ;
        RECT  29.85 429.0 34.95 429.9 ;
        RECT  37.5 428.1 41.85 429.0 ;
        RECT  31.65 427.65 32.85 428.85 ;
        RECT  34.05 427.65 35.25 428.85 ;
        RECT  34.05 427.65 35.25 428.85 ;
        RECT  36.45 427.65 37.65 428.85 ;
        RECT  31.65 428.25 32.85 429.45 ;
        RECT  34.05 428.25 35.25 429.45 ;
        RECT  34.05 428.25 35.25 429.45 ;
        RECT  36.45 428.25 37.65 429.45 ;
        RECT  38.85 423.45 40.05 424.65 ;
        RECT  38.85 433.65 40.05 434.85 ;
        RECT  31.95 426.9 33.15 428.1 ;
        RECT  34.95 430.2 36.15 431.4 ;
        RECT  41.85 199.65 51.45 200.55 ;
        RECT  41.85 214.35 51.45 215.25 ;
        RECT  48.45 211.95 49.65 214.35 ;
        RECT  48.45 200.55 49.65 202.35 ;
        RECT  43.65 200.55 44.85 201.45 ;
        RECT  43.65 213.15 44.85 214.35 ;
        RECT  46.05 202.65 47.25 212.1 ;
        RECT  41.85 206.4 43.95 207.3 ;
        RECT  47.25 206.4 51.45 207.3 ;
        RECT  43.65 202.65 44.85 203.85 ;
        RECT  46.05 202.65 47.25 203.85 ;
        RECT  43.65 211.95 44.85 213.15 ;
        RECT  46.05 211.95 47.25 213.15 ;
        RECT  48.45 211.95 49.65 213.15 ;
        RECT  48.45 201.45 49.65 202.65 ;
        RECT  43.95 206.25 45.15 207.45 ;
        RECT  41.85 229.05 51.45 229.95 ;
        RECT  41.85 214.35 51.45 215.25 ;
        RECT  48.45 215.25 49.65 217.65 ;
        RECT  48.45 227.25 49.65 229.05 ;
        RECT  43.65 228.15 44.85 229.05 ;
        RECT  43.65 215.25 44.85 216.45 ;
        RECT  46.05 217.5 47.25 226.95 ;
        RECT  41.85 222.3 43.95 223.2 ;
        RECT  47.25 222.3 51.45 223.2 ;
        RECT  43.65 223.35 44.85 224.55 ;
        RECT  46.05 223.35 47.25 224.55 ;
        RECT  43.65 222.45 44.85 223.65 ;
        RECT  46.05 222.45 47.25 223.65 ;
        RECT  48.45 217.65 49.65 218.85 ;
        RECT  48.45 228.15 49.65 229.35 ;
        RECT  43.95 223.35 45.15 224.55 ;
        RECT  41.85 229.05 51.45 229.95 ;
        RECT  41.85 243.75 51.45 244.65 ;
        RECT  48.45 241.35 49.65 243.75 ;
        RECT  48.45 229.95 49.65 231.75 ;
        RECT  43.65 229.95 44.85 230.85 ;
        RECT  43.65 242.55 44.85 243.75 ;
        RECT  46.05 232.05 47.25 241.5 ;
        RECT  41.85 235.8 43.95 236.7 ;
        RECT  47.25 235.8 51.45 236.7 ;
        RECT  43.65 232.05 44.85 233.25 ;
        RECT  46.05 232.05 47.25 233.25 ;
        RECT  43.65 241.35 44.85 242.55 ;
        RECT  46.05 241.35 47.25 242.55 ;
        RECT  48.45 241.35 49.65 242.55 ;
        RECT  48.45 230.85 49.65 232.05 ;
        RECT  43.95 235.65 45.15 236.85 ;
        RECT  41.85 258.45 51.45 259.35 ;
        RECT  41.85 243.75 51.45 244.65 ;
        RECT  48.45 244.65 49.65 247.05 ;
        RECT  48.45 256.65 49.65 258.45 ;
        RECT  43.65 257.55 44.85 258.45 ;
        RECT  43.65 244.65 44.85 245.85 ;
        RECT  46.05 246.9 47.25 256.35 ;
        RECT  41.85 251.7 43.95 252.6 ;
        RECT  47.25 251.7 51.45 252.6 ;
        RECT  43.65 252.75 44.85 253.95 ;
        RECT  46.05 252.75 47.25 253.95 ;
        RECT  43.65 251.85 44.85 253.05 ;
        RECT  46.05 251.85 47.25 253.05 ;
        RECT  48.45 247.05 49.65 248.25 ;
        RECT  48.45 257.55 49.65 258.75 ;
        RECT  43.95 252.75 45.15 253.95 ;
        RECT  41.85 258.45 51.45 259.35 ;
        RECT  41.85 273.15 51.45 274.05 ;
        RECT  48.45 270.75 49.65 273.15 ;
        RECT  48.45 259.35 49.65 261.15 ;
        RECT  43.65 259.35 44.85 260.25 ;
        RECT  43.65 271.95 44.85 273.15 ;
        RECT  46.05 261.45 47.25 270.9 ;
        RECT  41.85 265.2 43.95 266.1 ;
        RECT  47.25 265.2 51.45 266.1 ;
        RECT  43.65 261.45 44.85 262.65 ;
        RECT  46.05 261.45 47.25 262.65 ;
        RECT  43.65 270.75 44.85 271.95 ;
        RECT  46.05 270.75 47.25 271.95 ;
        RECT  48.45 270.75 49.65 271.95 ;
        RECT  48.45 260.25 49.65 261.45 ;
        RECT  43.95 265.05 45.15 266.25 ;
        RECT  41.85 287.85 51.45 288.75 ;
        RECT  41.85 273.15 51.45 274.05 ;
        RECT  48.45 274.05 49.65 276.45 ;
        RECT  48.45 286.05 49.65 287.85 ;
        RECT  43.65 286.95 44.85 287.85 ;
        RECT  43.65 274.05 44.85 275.25 ;
        RECT  46.05 276.3 47.25 285.75 ;
        RECT  41.85 281.1 43.95 282.0 ;
        RECT  47.25 281.1 51.45 282.0 ;
        RECT  43.65 282.15 44.85 283.35 ;
        RECT  46.05 282.15 47.25 283.35 ;
        RECT  43.65 281.25 44.85 282.45 ;
        RECT  46.05 281.25 47.25 282.45 ;
        RECT  48.45 276.45 49.65 277.65 ;
        RECT  48.45 286.95 49.65 288.15 ;
        RECT  43.95 282.15 45.15 283.35 ;
        RECT  41.85 287.85 51.45 288.75 ;
        RECT  41.85 302.55 51.45 303.45 ;
        RECT  48.45 300.15 49.65 302.55 ;
        RECT  48.45 288.75 49.65 290.55 ;
        RECT  43.65 288.75 44.85 289.65 ;
        RECT  43.65 301.35 44.85 302.55 ;
        RECT  46.05 290.85 47.25 300.3 ;
        RECT  41.85 294.6 43.95 295.5 ;
        RECT  47.25 294.6 51.45 295.5 ;
        RECT  43.65 290.85 44.85 292.05 ;
        RECT  46.05 290.85 47.25 292.05 ;
        RECT  43.65 300.15 44.85 301.35 ;
        RECT  46.05 300.15 47.25 301.35 ;
        RECT  48.45 300.15 49.65 301.35 ;
        RECT  48.45 289.65 49.65 290.85 ;
        RECT  43.95 294.45 45.15 295.65 ;
        RECT  41.85 317.25 51.45 318.15 ;
        RECT  41.85 302.55 51.45 303.45 ;
        RECT  48.45 303.45 49.65 305.85 ;
        RECT  48.45 315.45 49.65 317.25 ;
        RECT  43.65 316.35 44.85 317.25 ;
        RECT  43.65 303.45 44.85 304.65 ;
        RECT  46.05 305.7 47.25 315.15 ;
        RECT  41.85 310.5 43.95 311.4 ;
        RECT  47.25 310.5 51.45 311.4 ;
        RECT  43.65 311.55 44.85 312.75 ;
        RECT  46.05 311.55 47.25 312.75 ;
        RECT  43.65 310.65 44.85 311.85 ;
        RECT  46.05 310.65 47.25 311.85 ;
        RECT  48.45 305.85 49.65 307.05 ;
        RECT  48.45 316.35 49.65 317.55 ;
        RECT  43.95 311.55 45.15 312.75 ;
        RECT  41.85 317.25 51.45 318.15 ;
        RECT  41.85 331.95 51.45 332.85 ;
        RECT  48.45 329.55 49.65 331.95 ;
        RECT  48.45 318.15 49.65 319.95 ;
        RECT  43.65 318.15 44.85 319.05 ;
        RECT  43.65 330.75 44.85 331.95 ;
        RECT  46.05 320.25 47.25 329.7 ;
        RECT  41.85 324.0 43.95 324.9 ;
        RECT  47.25 324.0 51.45 324.9 ;
        RECT  43.65 320.25 44.85 321.45 ;
        RECT  46.05 320.25 47.25 321.45 ;
        RECT  43.65 329.55 44.85 330.75 ;
        RECT  46.05 329.55 47.25 330.75 ;
        RECT  48.45 329.55 49.65 330.75 ;
        RECT  48.45 319.05 49.65 320.25 ;
        RECT  43.95 323.85 45.15 325.05 ;
        RECT  41.85 346.65 51.45 347.55 ;
        RECT  41.85 331.95 51.45 332.85 ;
        RECT  48.45 332.85 49.65 335.25 ;
        RECT  48.45 344.85 49.65 346.65 ;
        RECT  43.65 345.75 44.85 346.65 ;
        RECT  43.65 332.85 44.85 334.05 ;
        RECT  46.05 335.1 47.25 344.55 ;
        RECT  41.85 339.9 43.95 340.8 ;
        RECT  47.25 339.9 51.45 340.8 ;
        RECT  43.65 340.95 44.85 342.15 ;
        RECT  46.05 340.95 47.25 342.15 ;
        RECT  43.65 340.05 44.85 341.25 ;
        RECT  46.05 340.05 47.25 341.25 ;
        RECT  48.45 335.25 49.65 336.45 ;
        RECT  48.45 345.75 49.65 346.95 ;
        RECT  43.95 340.95 45.15 342.15 ;
        RECT  41.85 346.65 51.45 347.55 ;
        RECT  41.85 361.35 51.45 362.25 ;
        RECT  48.45 358.95 49.65 361.35 ;
        RECT  48.45 347.55 49.65 349.35 ;
        RECT  43.65 347.55 44.85 348.45 ;
        RECT  43.65 360.15 44.85 361.35 ;
        RECT  46.05 349.65 47.25 359.1 ;
        RECT  41.85 353.4 43.95 354.3 ;
        RECT  47.25 353.4 51.45 354.3 ;
        RECT  43.65 349.65 44.85 350.85 ;
        RECT  46.05 349.65 47.25 350.85 ;
        RECT  43.65 358.95 44.85 360.15 ;
        RECT  46.05 358.95 47.25 360.15 ;
        RECT  48.45 358.95 49.65 360.15 ;
        RECT  48.45 348.45 49.65 349.65 ;
        RECT  43.95 353.25 45.15 354.45 ;
        RECT  41.85 376.05 51.45 376.95 ;
        RECT  41.85 361.35 51.45 362.25 ;
        RECT  48.45 362.25 49.65 364.65 ;
        RECT  48.45 374.25 49.65 376.05 ;
        RECT  43.65 375.15 44.85 376.05 ;
        RECT  43.65 362.25 44.85 363.45 ;
        RECT  46.05 364.5 47.25 373.95 ;
        RECT  41.85 369.3 43.95 370.2 ;
        RECT  47.25 369.3 51.45 370.2 ;
        RECT  43.65 370.35 44.85 371.55 ;
        RECT  46.05 370.35 47.25 371.55 ;
        RECT  43.65 369.45 44.85 370.65 ;
        RECT  46.05 369.45 47.25 370.65 ;
        RECT  48.45 364.65 49.65 365.85 ;
        RECT  48.45 375.15 49.65 376.35 ;
        RECT  43.95 370.35 45.15 371.55 ;
        RECT  41.85 376.05 51.45 376.95 ;
        RECT  41.85 390.75 51.45 391.65 ;
        RECT  48.45 388.35 49.65 390.75 ;
        RECT  48.45 376.95 49.65 378.75 ;
        RECT  43.65 376.95 44.85 377.85 ;
        RECT  43.65 389.55 44.85 390.75 ;
        RECT  46.05 379.05 47.25 388.5 ;
        RECT  41.85 382.8 43.95 383.7 ;
        RECT  47.25 382.8 51.45 383.7 ;
        RECT  43.65 379.05 44.85 380.25 ;
        RECT  46.05 379.05 47.25 380.25 ;
        RECT  43.65 388.35 44.85 389.55 ;
        RECT  46.05 388.35 47.25 389.55 ;
        RECT  48.45 388.35 49.65 389.55 ;
        RECT  48.45 377.85 49.65 379.05 ;
        RECT  43.95 382.65 45.15 383.85 ;
        RECT  41.85 405.45 51.45 406.35 ;
        RECT  41.85 390.75 51.45 391.65 ;
        RECT  48.45 391.65 49.65 394.05 ;
        RECT  48.45 403.65 49.65 405.45 ;
        RECT  43.65 404.55 44.85 405.45 ;
        RECT  43.65 391.65 44.85 392.85 ;
        RECT  46.05 393.9 47.25 403.35 ;
        RECT  41.85 398.7 43.95 399.6 ;
        RECT  47.25 398.7 51.45 399.6 ;
        RECT  43.65 399.75 44.85 400.95 ;
        RECT  46.05 399.75 47.25 400.95 ;
        RECT  43.65 398.85 44.85 400.05 ;
        RECT  46.05 398.85 47.25 400.05 ;
        RECT  48.45 394.05 49.65 395.25 ;
        RECT  48.45 404.55 49.65 405.75 ;
        RECT  43.95 399.75 45.15 400.95 ;
        RECT  41.85 405.45 51.45 406.35 ;
        RECT  41.85 420.15 51.45 421.05 ;
        RECT  48.45 417.75 49.65 420.15 ;
        RECT  48.45 406.35 49.65 408.15 ;
        RECT  43.65 406.35 44.85 407.25 ;
        RECT  43.65 418.95 44.85 420.15 ;
        RECT  46.05 408.45 47.25 417.9 ;
        RECT  41.85 412.2 43.95 413.1 ;
        RECT  47.25 412.2 51.45 413.1 ;
        RECT  43.65 408.45 44.85 409.65 ;
        RECT  46.05 408.45 47.25 409.65 ;
        RECT  43.65 417.75 44.85 418.95 ;
        RECT  46.05 417.75 47.25 418.95 ;
        RECT  48.45 417.75 49.65 418.95 ;
        RECT  48.45 407.25 49.65 408.45 ;
        RECT  43.95 412.05 45.15 413.25 ;
        RECT  41.85 434.85 51.45 435.75 ;
        RECT  41.85 420.15 51.45 421.05 ;
        RECT  48.45 421.05 49.65 423.45 ;
        RECT  48.45 433.05 49.65 434.85 ;
        RECT  43.65 433.95 44.85 434.85 ;
        RECT  43.65 421.05 44.85 422.25 ;
        RECT  46.05 423.3 47.25 432.75 ;
        RECT  41.85 428.1 43.95 429.0 ;
        RECT  47.25 428.1 51.45 429.0 ;
        RECT  43.65 429.15 44.85 430.35 ;
        RECT  46.05 429.15 47.25 430.35 ;
        RECT  43.65 428.25 44.85 429.45 ;
        RECT  46.05 428.25 47.25 429.45 ;
        RECT  48.45 423.45 49.65 424.65 ;
        RECT  48.45 433.95 49.65 435.15 ;
        RECT  43.95 429.15 45.15 430.35 ;
        RECT  13.05 88.8 14.25 90.0 ;
        RECT  15.15 104.7 16.35 105.9 ;
        RECT  17.25 118.2 18.45 119.4 ;
        RECT  19.35 134.1 20.55 135.3 ;
        RECT  21.45 147.6 22.65 148.8 ;
        RECT  23.55 163.5 24.75 164.7 ;
        RECT  25.65 177.0 26.85 178.2 ;
        RECT  27.75 192.9 28.95 194.1 ;
        RECT  13.05 208.8 14.25 210.0 ;
        RECT  21.45 205.5 22.65 206.7 ;
        RECT  13.05 219.9 14.25 221.1 ;
        RECT  23.55 223.2 24.75 224.4 ;
        RECT  13.05 238.2 14.25 239.4 ;
        RECT  25.65 234.9 26.85 236.1 ;
        RECT  13.05 249.3 14.25 250.5 ;
        RECT  27.75 252.6 28.95 253.8 ;
        RECT  15.15 267.6 16.35 268.8 ;
        RECT  21.45 264.3 22.65 265.5 ;
        RECT  15.15 278.7 16.35 279.9 ;
        RECT  23.55 282.0 24.75 283.2 ;
        RECT  15.15 297.0 16.35 298.2 ;
        RECT  25.65 293.7 26.85 294.9 ;
        RECT  15.15 308.1 16.35 309.3 ;
        RECT  27.75 311.4 28.95 312.6 ;
        RECT  17.25 326.4 18.45 327.6 ;
        RECT  21.45 323.1 22.65 324.3 ;
        RECT  17.25 337.5 18.45 338.7 ;
        RECT  23.55 340.8 24.75 342.0 ;
        RECT  17.25 355.8 18.45 357.0 ;
        RECT  25.65 352.5 26.85 353.7 ;
        RECT  17.25 366.9 18.45 368.1 ;
        RECT  27.75 370.2 28.95 371.4 ;
        RECT  19.35 385.2 20.55 386.4 ;
        RECT  21.45 381.9 22.65 383.1 ;
        RECT  19.35 396.3 20.55 397.5 ;
        RECT  23.55 399.6 24.75 400.8 ;
        RECT  19.35 414.6 20.55 415.8 ;
        RECT  25.65 411.3 26.85 412.5 ;
        RECT  19.35 425.7 20.55 426.9 ;
        RECT  27.75 429.0 28.95 430.2 ;
        RECT  54.15 201.9 55.05 440.7 ;
        RECT  54.15 206.4 58.65 207.3 ;
        RECT  66.45 205.5 67.35 207.3 ;
        RECT  79.35 206.4 80.25 207.3 ;
        RECT  88.95 206.4 89.85 207.3 ;
        RECT  54.15 222.3 58.65 223.2 ;
        RECT  66.45 222.3 67.35 224.1 ;
        RECT  79.35 222.3 80.25 223.2 ;
        RECT  88.05 222.3 88.95 223.2 ;
        RECT  54.15 235.8 58.65 236.7 ;
        RECT  66.45 234.9 67.35 236.7 ;
        RECT  79.35 235.8 80.25 236.7 ;
        RECT  88.95 235.8 89.85 236.7 ;
        RECT  54.15 251.7 58.65 252.6 ;
        RECT  66.45 251.7 67.35 253.5 ;
        RECT  79.35 251.7 80.25 252.6 ;
        RECT  88.05 251.7 88.95 252.6 ;
        RECT  54.15 265.2 58.65 266.1 ;
        RECT  66.45 264.3 67.35 266.1 ;
        RECT  79.35 265.2 80.25 266.1 ;
        RECT  88.95 265.2 89.85 266.1 ;
        RECT  54.15 281.1 58.65 282.0 ;
        RECT  66.45 281.1 67.35 282.9 ;
        RECT  79.35 281.1 80.25 282.0 ;
        RECT  88.05 281.1 88.95 282.0 ;
        RECT  54.15 294.6 58.65 295.5 ;
        RECT  66.45 293.7 67.35 295.5 ;
        RECT  79.35 294.6 80.25 295.5 ;
        RECT  88.95 294.6 89.85 295.5 ;
        RECT  54.15 310.5 58.65 311.4 ;
        RECT  66.45 310.5 67.35 312.3 ;
        RECT  79.35 310.5 80.25 311.4 ;
        RECT  88.05 310.5 88.95 311.4 ;
        RECT  54.15 324.0 58.65 324.9 ;
        RECT  66.45 323.1 67.35 324.9 ;
        RECT  79.35 324.0 80.25 324.9 ;
        RECT  88.95 324.0 89.85 324.9 ;
        RECT  54.15 339.9 58.65 340.8 ;
        RECT  66.45 339.9 67.35 341.7 ;
        RECT  79.35 339.9 80.25 340.8 ;
        RECT  88.05 339.9 88.95 340.8 ;
        RECT  54.15 353.4 58.65 354.3 ;
        RECT  66.45 352.5 67.35 354.3 ;
        RECT  79.35 353.4 80.25 354.3 ;
        RECT  88.95 353.4 89.85 354.3 ;
        RECT  54.15 369.3 58.65 370.2 ;
        RECT  66.45 369.3 67.35 371.1 ;
        RECT  79.35 369.3 80.25 370.2 ;
        RECT  88.05 369.3 88.95 370.2 ;
        RECT  54.15 382.8 58.65 383.7 ;
        RECT  66.45 381.9 67.35 383.7 ;
        RECT  79.35 382.8 80.25 383.7 ;
        RECT  88.95 382.8 89.85 383.7 ;
        RECT  54.15 398.7 58.65 399.6 ;
        RECT  66.45 398.7 67.35 400.5 ;
        RECT  79.35 398.7 80.25 399.6 ;
        RECT  88.05 398.7 88.95 399.6 ;
        RECT  54.15 412.2 58.65 413.1 ;
        RECT  66.45 411.3 67.35 413.1 ;
        RECT  79.35 412.2 80.25 413.1 ;
        RECT  88.95 412.2 89.85 413.1 ;
        RECT  54.15 428.1 58.65 429.0 ;
        RECT  66.45 428.1 67.35 429.9 ;
        RECT  79.35 428.1 80.25 429.0 ;
        RECT  88.05 428.1 88.95 429.0 ;
        RECT  51.15 214.35 52.35 215.55 ;
        RECT  57.45 214.35 58.65 215.55 ;
        RECT  57.75 199.65 67.35 200.55 ;
        RECT  57.75 214.35 67.35 215.25 ;
        RECT  64.35 211.95 65.55 214.35 ;
        RECT  64.35 200.55 65.55 202.35 ;
        RECT  59.55 200.55 60.75 201.45 ;
        RECT  59.55 213.15 60.75 214.35 ;
        RECT  61.95 202.65 63.15 212.1 ;
        RECT  57.75 206.4 59.85 207.3 ;
        RECT  63.15 206.4 67.35 207.3 ;
        RECT  59.55 202.65 60.75 203.85 ;
        RECT  61.95 202.65 63.15 203.85 ;
        RECT  59.55 211.95 60.75 213.15 ;
        RECT  61.95 211.95 63.15 213.15 ;
        RECT  64.35 211.95 65.55 213.15 ;
        RECT  64.35 201.45 65.55 202.65 ;
        RECT  59.85 206.25 61.05 207.45 ;
        RECT  67.35 199.65 79.35 200.55 ;
        RECT  67.35 214.35 79.35 215.25 ;
        RECT  76.35 211.95 77.25 214.8 ;
        RECT  76.35 200.1 77.25 202.5 ;
        RECT  69.3 211.95 70.2 214.8 ;
        RECT  74.1 211.95 75.0 214.8 ;
        RECT  69.3 200.1 70.2 202.95 ;
        RECT  74.55 208.8 75.45 209.7 ;
        RECT  71.55 208.8 72.45 209.7 ;
        RECT  74.55 201.75 75.45 209.25 ;
        RECT  72.0 208.8 75.0 209.7 ;
        RECT  71.55 209.25 72.45 211.95 ;
        RECT  67.35 208.8 69.45 209.7 ;
        RECT  67.35 205.5 72.45 206.4 ;
        RECT  75.0 206.4 79.35 207.3 ;
        RECT  69.15 202.95 70.35 204.15 ;
        RECT  71.55 202.95 72.75 204.15 ;
        RECT  71.55 202.95 72.75 204.15 ;
        RECT  73.95 202.95 75.15 204.15 ;
        RECT  69.15 211.95 70.35 213.15 ;
        RECT  71.55 211.95 72.75 213.15 ;
        RECT  71.55 211.95 72.75 213.15 ;
        RECT  73.95 211.95 75.15 213.15 ;
        RECT  76.35 211.95 77.55 213.15 ;
        RECT  76.35 201.75 77.55 202.95 ;
        RECT  69.45 208.5 70.65 209.7 ;
        RECT  72.45 205.2 73.65 206.4 ;
        RECT  79.35 199.65 88.95 200.55 ;
        RECT  79.35 214.35 88.95 215.25 ;
        RECT  85.95 211.95 87.15 214.35 ;
        RECT  85.95 200.55 87.15 202.35 ;
        RECT  81.15 200.55 82.35 201.45 ;
        RECT  81.15 213.15 82.35 214.35 ;
        RECT  83.55 202.65 84.75 212.1 ;
        RECT  79.35 206.4 81.45 207.3 ;
        RECT  84.75 206.4 88.95 207.3 ;
        RECT  81.15 202.65 82.35 203.85 ;
        RECT  83.55 202.65 84.75 203.85 ;
        RECT  81.15 211.95 82.35 213.15 ;
        RECT  83.55 211.95 84.75 213.15 ;
        RECT  85.95 211.95 87.15 213.15 ;
        RECT  85.95 201.45 87.15 202.65 ;
        RECT  81.45 206.25 82.65 207.45 ;
        RECT  67.35 208.8 68.55 210.0 ;
        RECT  51.45 208.8 52.65 210.0 ;
        RECT  51.15 229.05 52.35 230.25 ;
        RECT  57.45 229.05 58.65 230.25 ;
        RECT  57.75 229.05 67.35 229.95 ;
        RECT  57.75 214.35 67.35 215.25 ;
        RECT  64.35 215.25 65.55 217.65 ;
        RECT  64.35 227.25 65.55 229.05 ;
        RECT  59.55 228.15 60.75 229.05 ;
        RECT  59.55 215.25 60.75 216.45 ;
        RECT  61.95 217.5 63.15 226.95 ;
        RECT  57.75 222.3 59.85 223.2 ;
        RECT  63.15 222.3 67.35 223.2 ;
        RECT  59.55 223.35 60.75 224.55 ;
        RECT  61.95 223.35 63.15 224.55 ;
        RECT  59.55 222.45 60.75 223.65 ;
        RECT  61.95 222.45 63.15 223.65 ;
        RECT  64.35 217.65 65.55 218.85 ;
        RECT  64.35 228.15 65.55 229.35 ;
        RECT  59.85 223.35 61.05 224.55 ;
        RECT  67.35 229.05 79.35 229.95 ;
        RECT  67.35 214.35 79.35 215.25 ;
        RECT  76.35 214.8 77.25 217.65 ;
        RECT  76.35 227.1 77.25 229.5 ;
        RECT  69.3 214.8 70.2 217.65 ;
        RECT  74.1 214.8 75.0 217.65 ;
        RECT  69.3 226.65 70.2 229.5 ;
        RECT  74.55 219.9 75.45 220.8 ;
        RECT  71.55 219.9 72.45 220.8 ;
        RECT  74.55 220.35 75.45 227.85 ;
        RECT  72.0 219.9 75.0 220.8 ;
        RECT  71.55 217.65 72.45 220.35 ;
        RECT  67.35 219.9 69.45 220.8 ;
        RECT  67.35 223.2 72.45 224.1 ;
        RECT  75.0 222.3 79.35 223.2 ;
        RECT  69.15 221.85 70.35 223.05 ;
        RECT  71.55 221.85 72.75 223.05 ;
        RECT  71.55 221.85 72.75 223.05 ;
        RECT  73.95 221.85 75.15 223.05 ;
        RECT  69.15 222.45 70.35 223.65 ;
        RECT  71.55 222.45 72.75 223.65 ;
        RECT  71.55 222.45 72.75 223.65 ;
        RECT  73.95 222.45 75.15 223.65 ;
        RECT  76.35 217.65 77.55 218.85 ;
        RECT  76.35 227.85 77.55 229.05 ;
        RECT  69.45 221.1 70.65 222.3 ;
        RECT  72.45 224.4 73.65 225.6 ;
        RECT  79.35 229.05 88.95 229.95 ;
        RECT  79.35 214.35 88.95 215.25 ;
        RECT  85.95 215.25 87.15 217.65 ;
        RECT  85.95 227.25 87.15 229.05 ;
        RECT  81.15 228.15 82.35 229.05 ;
        RECT  81.15 215.25 82.35 216.45 ;
        RECT  83.55 217.5 84.75 226.95 ;
        RECT  79.35 222.3 81.45 223.2 ;
        RECT  84.75 222.3 88.95 223.2 ;
        RECT  81.15 223.35 82.35 224.55 ;
        RECT  83.55 223.35 84.75 224.55 ;
        RECT  81.15 222.45 82.35 223.65 ;
        RECT  83.55 222.45 84.75 223.65 ;
        RECT  85.95 217.65 87.15 218.85 ;
        RECT  85.95 228.15 87.15 229.35 ;
        RECT  81.45 223.35 82.65 224.55 ;
        RECT  67.35 219.6 68.55 220.8 ;
        RECT  51.45 219.6 52.65 220.8 ;
        RECT  51.15 243.75 52.35 244.95 ;
        RECT  57.45 243.75 58.65 244.95 ;
        RECT  57.75 229.05 67.35 229.95 ;
        RECT  57.75 243.75 67.35 244.65 ;
        RECT  64.35 241.35 65.55 243.75 ;
        RECT  64.35 229.95 65.55 231.75 ;
        RECT  59.55 229.95 60.75 230.85 ;
        RECT  59.55 242.55 60.75 243.75 ;
        RECT  61.95 232.05 63.15 241.5 ;
        RECT  57.75 235.8 59.85 236.7 ;
        RECT  63.15 235.8 67.35 236.7 ;
        RECT  59.55 232.05 60.75 233.25 ;
        RECT  61.95 232.05 63.15 233.25 ;
        RECT  59.55 241.35 60.75 242.55 ;
        RECT  61.95 241.35 63.15 242.55 ;
        RECT  64.35 241.35 65.55 242.55 ;
        RECT  64.35 230.85 65.55 232.05 ;
        RECT  59.85 235.65 61.05 236.85 ;
        RECT  67.35 229.05 79.35 229.95 ;
        RECT  67.35 243.75 79.35 244.65 ;
        RECT  76.35 241.35 77.25 244.2 ;
        RECT  76.35 229.5 77.25 231.9 ;
        RECT  69.3 241.35 70.2 244.2 ;
        RECT  74.1 241.35 75.0 244.2 ;
        RECT  69.3 229.5 70.2 232.35 ;
        RECT  74.55 238.2 75.45 239.1 ;
        RECT  71.55 238.2 72.45 239.1 ;
        RECT  74.55 231.15 75.45 238.65 ;
        RECT  72.0 238.2 75.0 239.1 ;
        RECT  71.55 238.65 72.45 241.35 ;
        RECT  67.35 238.2 69.45 239.1 ;
        RECT  67.35 234.9 72.45 235.8 ;
        RECT  75.0 235.8 79.35 236.7 ;
        RECT  69.15 232.35 70.35 233.55 ;
        RECT  71.55 232.35 72.75 233.55 ;
        RECT  71.55 232.35 72.75 233.55 ;
        RECT  73.95 232.35 75.15 233.55 ;
        RECT  69.15 241.35 70.35 242.55 ;
        RECT  71.55 241.35 72.75 242.55 ;
        RECT  71.55 241.35 72.75 242.55 ;
        RECT  73.95 241.35 75.15 242.55 ;
        RECT  76.35 241.35 77.55 242.55 ;
        RECT  76.35 231.15 77.55 232.35 ;
        RECT  69.45 237.9 70.65 239.1 ;
        RECT  72.45 234.6 73.65 235.8 ;
        RECT  79.35 229.05 88.95 229.95 ;
        RECT  79.35 243.75 88.95 244.65 ;
        RECT  85.95 241.35 87.15 243.75 ;
        RECT  85.95 229.95 87.15 231.75 ;
        RECT  81.15 229.95 82.35 230.85 ;
        RECT  81.15 242.55 82.35 243.75 ;
        RECT  83.55 232.05 84.75 241.5 ;
        RECT  79.35 235.8 81.45 236.7 ;
        RECT  84.75 235.8 88.95 236.7 ;
        RECT  81.15 232.05 82.35 233.25 ;
        RECT  83.55 232.05 84.75 233.25 ;
        RECT  81.15 241.35 82.35 242.55 ;
        RECT  83.55 241.35 84.75 242.55 ;
        RECT  85.95 241.35 87.15 242.55 ;
        RECT  85.95 230.85 87.15 232.05 ;
        RECT  81.45 235.65 82.65 236.85 ;
        RECT  67.35 238.2 68.55 239.4 ;
        RECT  51.45 238.2 52.65 239.4 ;
        RECT  51.15 258.45 52.35 259.65 ;
        RECT  57.45 258.45 58.65 259.65 ;
        RECT  57.75 258.45 67.35 259.35 ;
        RECT  57.75 243.75 67.35 244.65 ;
        RECT  64.35 244.65 65.55 247.05 ;
        RECT  64.35 256.65 65.55 258.45 ;
        RECT  59.55 257.55 60.75 258.45 ;
        RECT  59.55 244.65 60.75 245.85 ;
        RECT  61.95 246.9 63.15 256.35 ;
        RECT  57.75 251.7 59.85 252.6 ;
        RECT  63.15 251.7 67.35 252.6 ;
        RECT  59.55 252.75 60.75 253.95 ;
        RECT  61.95 252.75 63.15 253.95 ;
        RECT  59.55 251.85 60.75 253.05 ;
        RECT  61.95 251.85 63.15 253.05 ;
        RECT  64.35 247.05 65.55 248.25 ;
        RECT  64.35 257.55 65.55 258.75 ;
        RECT  59.85 252.75 61.05 253.95 ;
        RECT  67.35 258.45 79.35 259.35 ;
        RECT  67.35 243.75 79.35 244.65 ;
        RECT  76.35 244.2 77.25 247.05 ;
        RECT  76.35 256.5 77.25 258.9 ;
        RECT  69.3 244.2 70.2 247.05 ;
        RECT  74.1 244.2 75.0 247.05 ;
        RECT  69.3 256.05 70.2 258.9 ;
        RECT  74.55 249.3 75.45 250.2 ;
        RECT  71.55 249.3 72.45 250.2 ;
        RECT  74.55 249.75 75.45 257.25 ;
        RECT  72.0 249.3 75.0 250.2 ;
        RECT  71.55 247.05 72.45 249.75 ;
        RECT  67.35 249.3 69.45 250.2 ;
        RECT  67.35 252.6 72.45 253.5 ;
        RECT  75.0 251.7 79.35 252.6 ;
        RECT  69.15 251.25 70.35 252.45 ;
        RECT  71.55 251.25 72.75 252.45 ;
        RECT  71.55 251.25 72.75 252.45 ;
        RECT  73.95 251.25 75.15 252.45 ;
        RECT  69.15 251.85 70.35 253.05 ;
        RECT  71.55 251.85 72.75 253.05 ;
        RECT  71.55 251.85 72.75 253.05 ;
        RECT  73.95 251.85 75.15 253.05 ;
        RECT  76.35 247.05 77.55 248.25 ;
        RECT  76.35 257.25 77.55 258.45 ;
        RECT  69.45 250.5 70.65 251.7 ;
        RECT  72.45 253.8 73.65 255.0 ;
        RECT  79.35 258.45 88.95 259.35 ;
        RECT  79.35 243.75 88.95 244.65 ;
        RECT  85.95 244.65 87.15 247.05 ;
        RECT  85.95 256.65 87.15 258.45 ;
        RECT  81.15 257.55 82.35 258.45 ;
        RECT  81.15 244.65 82.35 245.85 ;
        RECT  83.55 246.9 84.75 256.35 ;
        RECT  79.35 251.7 81.45 252.6 ;
        RECT  84.75 251.7 88.95 252.6 ;
        RECT  81.15 252.75 82.35 253.95 ;
        RECT  83.55 252.75 84.75 253.95 ;
        RECT  81.15 251.85 82.35 253.05 ;
        RECT  83.55 251.85 84.75 253.05 ;
        RECT  85.95 247.05 87.15 248.25 ;
        RECT  85.95 257.55 87.15 258.75 ;
        RECT  81.45 252.75 82.65 253.95 ;
        RECT  67.35 249.0 68.55 250.2 ;
        RECT  51.45 249.0 52.65 250.2 ;
        RECT  51.15 273.15 52.35 274.35 ;
        RECT  57.45 273.15 58.65 274.35 ;
        RECT  57.75 258.45 67.35 259.35 ;
        RECT  57.75 273.15 67.35 274.05 ;
        RECT  64.35 270.75 65.55 273.15 ;
        RECT  64.35 259.35 65.55 261.15 ;
        RECT  59.55 259.35 60.75 260.25 ;
        RECT  59.55 271.95 60.75 273.15 ;
        RECT  61.95 261.45 63.15 270.9 ;
        RECT  57.75 265.2 59.85 266.1 ;
        RECT  63.15 265.2 67.35 266.1 ;
        RECT  59.55 261.45 60.75 262.65 ;
        RECT  61.95 261.45 63.15 262.65 ;
        RECT  59.55 270.75 60.75 271.95 ;
        RECT  61.95 270.75 63.15 271.95 ;
        RECT  64.35 270.75 65.55 271.95 ;
        RECT  64.35 260.25 65.55 261.45 ;
        RECT  59.85 265.05 61.05 266.25 ;
        RECT  67.35 258.45 79.35 259.35 ;
        RECT  67.35 273.15 79.35 274.05 ;
        RECT  76.35 270.75 77.25 273.6 ;
        RECT  76.35 258.9 77.25 261.3 ;
        RECT  69.3 270.75 70.2 273.6 ;
        RECT  74.1 270.75 75.0 273.6 ;
        RECT  69.3 258.9 70.2 261.75 ;
        RECT  74.55 267.6 75.45 268.5 ;
        RECT  71.55 267.6 72.45 268.5 ;
        RECT  74.55 260.55 75.45 268.05 ;
        RECT  72.0 267.6 75.0 268.5 ;
        RECT  71.55 268.05 72.45 270.75 ;
        RECT  67.35 267.6 69.45 268.5 ;
        RECT  67.35 264.3 72.45 265.2 ;
        RECT  75.0 265.2 79.35 266.1 ;
        RECT  69.15 261.75 70.35 262.95 ;
        RECT  71.55 261.75 72.75 262.95 ;
        RECT  71.55 261.75 72.75 262.95 ;
        RECT  73.95 261.75 75.15 262.95 ;
        RECT  69.15 270.75 70.35 271.95 ;
        RECT  71.55 270.75 72.75 271.95 ;
        RECT  71.55 270.75 72.75 271.95 ;
        RECT  73.95 270.75 75.15 271.95 ;
        RECT  76.35 270.75 77.55 271.95 ;
        RECT  76.35 260.55 77.55 261.75 ;
        RECT  69.45 267.3 70.65 268.5 ;
        RECT  72.45 264.0 73.65 265.2 ;
        RECT  79.35 258.45 88.95 259.35 ;
        RECT  79.35 273.15 88.95 274.05 ;
        RECT  85.95 270.75 87.15 273.15 ;
        RECT  85.95 259.35 87.15 261.15 ;
        RECT  81.15 259.35 82.35 260.25 ;
        RECT  81.15 271.95 82.35 273.15 ;
        RECT  83.55 261.45 84.75 270.9 ;
        RECT  79.35 265.2 81.45 266.1 ;
        RECT  84.75 265.2 88.95 266.1 ;
        RECT  81.15 261.45 82.35 262.65 ;
        RECT  83.55 261.45 84.75 262.65 ;
        RECT  81.15 270.75 82.35 271.95 ;
        RECT  83.55 270.75 84.75 271.95 ;
        RECT  85.95 270.75 87.15 271.95 ;
        RECT  85.95 260.25 87.15 261.45 ;
        RECT  81.45 265.05 82.65 266.25 ;
        RECT  67.35 267.6 68.55 268.8 ;
        RECT  51.45 267.6 52.65 268.8 ;
        RECT  51.15 287.85 52.35 289.05 ;
        RECT  57.45 287.85 58.65 289.05 ;
        RECT  57.75 287.85 67.35 288.75 ;
        RECT  57.75 273.15 67.35 274.05 ;
        RECT  64.35 274.05 65.55 276.45 ;
        RECT  64.35 286.05 65.55 287.85 ;
        RECT  59.55 286.95 60.75 287.85 ;
        RECT  59.55 274.05 60.75 275.25 ;
        RECT  61.95 276.3 63.15 285.75 ;
        RECT  57.75 281.1 59.85 282.0 ;
        RECT  63.15 281.1 67.35 282.0 ;
        RECT  59.55 282.15 60.75 283.35 ;
        RECT  61.95 282.15 63.15 283.35 ;
        RECT  59.55 281.25 60.75 282.45 ;
        RECT  61.95 281.25 63.15 282.45 ;
        RECT  64.35 276.45 65.55 277.65 ;
        RECT  64.35 286.95 65.55 288.15 ;
        RECT  59.85 282.15 61.05 283.35 ;
        RECT  67.35 287.85 79.35 288.75 ;
        RECT  67.35 273.15 79.35 274.05 ;
        RECT  76.35 273.6 77.25 276.45 ;
        RECT  76.35 285.9 77.25 288.3 ;
        RECT  69.3 273.6 70.2 276.45 ;
        RECT  74.1 273.6 75.0 276.45 ;
        RECT  69.3 285.45 70.2 288.3 ;
        RECT  74.55 278.7 75.45 279.6 ;
        RECT  71.55 278.7 72.45 279.6 ;
        RECT  74.55 279.15 75.45 286.65 ;
        RECT  72.0 278.7 75.0 279.6 ;
        RECT  71.55 276.45 72.45 279.15 ;
        RECT  67.35 278.7 69.45 279.6 ;
        RECT  67.35 282.0 72.45 282.9 ;
        RECT  75.0 281.1 79.35 282.0 ;
        RECT  69.15 280.65 70.35 281.85 ;
        RECT  71.55 280.65 72.75 281.85 ;
        RECT  71.55 280.65 72.75 281.85 ;
        RECT  73.95 280.65 75.15 281.85 ;
        RECT  69.15 281.25 70.35 282.45 ;
        RECT  71.55 281.25 72.75 282.45 ;
        RECT  71.55 281.25 72.75 282.45 ;
        RECT  73.95 281.25 75.15 282.45 ;
        RECT  76.35 276.45 77.55 277.65 ;
        RECT  76.35 286.65 77.55 287.85 ;
        RECT  69.45 279.9 70.65 281.1 ;
        RECT  72.45 283.2 73.65 284.4 ;
        RECT  79.35 287.85 88.95 288.75 ;
        RECT  79.35 273.15 88.95 274.05 ;
        RECT  85.95 274.05 87.15 276.45 ;
        RECT  85.95 286.05 87.15 287.85 ;
        RECT  81.15 286.95 82.35 287.85 ;
        RECT  81.15 274.05 82.35 275.25 ;
        RECT  83.55 276.3 84.75 285.75 ;
        RECT  79.35 281.1 81.45 282.0 ;
        RECT  84.75 281.1 88.95 282.0 ;
        RECT  81.15 282.15 82.35 283.35 ;
        RECT  83.55 282.15 84.75 283.35 ;
        RECT  81.15 281.25 82.35 282.45 ;
        RECT  83.55 281.25 84.75 282.45 ;
        RECT  85.95 276.45 87.15 277.65 ;
        RECT  85.95 286.95 87.15 288.15 ;
        RECT  81.45 282.15 82.65 283.35 ;
        RECT  67.35 278.4 68.55 279.6 ;
        RECT  51.45 278.4 52.65 279.6 ;
        RECT  51.15 302.55 52.35 303.75 ;
        RECT  57.45 302.55 58.65 303.75 ;
        RECT  57.75 287.85 67.35 288.75 ;
        RECT  57.75 302.55 67.35 303.45 ;
        RECT  64.35 300.15 65.55 302.55 ;
        RECT  64.35 288.75 65.55 290.55 ;
        RECT  59.55 288.75 60.75 289.65 ;
        RECT  59.55 301.35 60.75 302.55 ;
        RECT  61.95 290.85 63.15 300.3 ;
        RECT  57.75 294.6 59.85 295.5 ;
        RECT  63.15 294.6 67.35 295.5 ;
        RECT  59.55 290.85 60.75 292.05 ;
        RECT  61.95 290.85 63.15 292.05 ;
        RECT  59.55 300.15 60.75 301.35 ;
        RECT  61.95 300.15 63.15 301.35 ;
        RECT  64.35 300.15 65.55 301.35 ;
        RECT  64.35 289.65 65.55 290.85 ;
        RECT  59.85 294.45 61.05 295.65 ;
        RECT  67.35 287.85 79.35 288.75 ;
        RECT  67.35 302.55 79.35 303.45 ;
        RECT  76.35 300.15 77.25 303.0 ;
        RECT  76.35 288.3 77.25 290.7 ;
        RECT  69.3 300.15 70.2 303.0 ;
        RECT  74.1 300.15 75.0 303.0 ;
        RECT  69.3 288.3 70.2 291.15 ;
        RECT  74.55 297.0 75.45 297.9 ;
        RECT  71.55 297.0 72.45 297.9 ;
        RECT  74.55 289.95 75.45 297.45 ;
        RECT  72.0 297.0 75.0 297.9 ;
        RECT  71.55 297.45 72.45 300.15 ;
        RECT  67.35 297.0 69.45 297.9 ;
        RECT  67.35 293.7 72.45 294.6 ;
        RECT  75.0 294.6 79.35 295.5 ;
        RECT  69.15 291.15 70.35 292.35 ;
        RECT  71.55 291.15 72.75 292.35 ;
        RECT  71.55 291.15 72.75 292.35 ;
        RECT  73.95 291.15 75.15 292.35 ;
        RECT  69.15 300.15 70.35 301.35 ;
        RECT  71.55 300.15 72.75 301.35 ;
        RECT  71.55 300.15 72.75 301.35 ;
        RECT  73.95 300.15 75.15 301.35 ;
        RECT  76.35 300.15 77.55 301.35 ;
        RECT  76.35 289.95 77.55 291.15 ;
        RECT  69.45 296.7 70.65 297.9 ;
        RECT  72.45 293.4 73.65 294.6 ;
        RECT  79.35 287.85 88.95 288.75 ;
        RECT  79.35 302.55 88.95 303.45 ;
        RECT  85.95 300.15 87.15 302.55 ;
        RECT  85.95 288.75 87.15 290.55 ;
        RECT  81.15 288.75 82.35 289.65 ;
        RECT  81.15 301.35 82.35 302.55 ;
        RECT  83.55 290.85 84.75 300.3 ;
        RECT  79.35 294.6 81.45 295.5 ;
        RECT  84.75 294.6 88.95 295.5 ;
        RECT  81.15 290.85 82.35 292.05 ;
        RECT  83.55 290.85 84.75 292.05 ;
        RECT  81.15 300.15 82.35 301.35 ;
        RECT  83.55 300.15 84.75 301.35 ;
        RECT  85.95 300.15 87.15 301.35 ;
        RECT  85.95 289.65 87.15 290.85 ;
        RECT  81.45 294.45 82.65 295.65 ;
        RECT  67.35 297.0 68.55 298.2 ;
        RECT  51.45 297.0 52.65 298.2 ;
        RECT  51.15 317.25 52.35 318.45 ;
        RECT  57.45 317.25 58.65 318.45 ;
        RECT  57.75 317.25 67.35 318.15 ;
        RECT  57.75 302.55 67.35 303.45 ;
        RECT  64.35 303.45 65.55 305.85 ;
        RECT  64.35 315.45 65.55 317.25 ;
        RECT  59.55 316.35 60.75 317.25 ;
        RECT  59.55 303.45 60.75 304.65 ;
        RECT  61.95 305.7 63.15 315.15 ;
        RECT  57.75 310.5 59.85 311.4 ;
        RECT  63.15 310.5 67.35 311.4 ;
        RECT  59.55 311.55 60.75 312.75 ;
        RECT  61.95 311.55 63.15 312.75 ;
        RECT  59.55 310.65 60.75 311.85 ;
        RECT  61.95 310.65 63.15 311.85 ;
        RECT  64.35 305.85 65.55 307.05 ;
        RECT  64.35 316.35 65.55 317.55 ;
        RECT  59.85 311.55 61.05 312.75 ;
        RECT  67.35 317.25 79.35 318.15 ;
        RECT  67.35 302.55 79.35 303.45 ;
        RECT  76.35 303.0 77.25 305.85 ;
        RECT  76.35 315.3 77.25 317.7 ;
        RECT  69.3 303.0 70.2 305.85 ;
        RECT  74.1 303.0 75.0 305.85 ;
        RECT  69.3 314.85 70.2 317.7 ;
        RECT  74.55 308.1 75.45 309.0 ;
        RECT  71.55 308.1 72.45 309.0 ;
        RECT  74.55 308.55 75.45 316.05 ;
        RECT  72.0 308.1 75.0 309.0 ;
        RECT  71.55 305.85 72.45 308.55 ;
        RECT  67.35 308.1 69.45 309.0 ;
        RECT  67.35 311.4 72.45 312.3 ;
        RECT  75.0 310.5 79.35 311.4 ;
        RECT  69.15 310.05 70.35 311.25 ;
        RECT  71.55 310.05 72.75 311.25 ;
        RECT  71.55 310.05 72.75 311.25 ;
        RECT  73.95 310.05 75.15 311.25 ;
        RECT  69.15 310.65 70.35 311.85 ;
        RECT  71.55 310.65 72.75 311.85 ;
        RECT  71.55 310.65 72.75 311.85 ;
        RECT  73.95 310.65 75.15 311.85 ;
        RECT  76.35 305.85 77.55 307.05 ;
        RECT  76.35 316.05 77.55 317.25 ;
        RECT  69.45 309.3 70.65 310.5 ;
        RECT  72.45 312.6 73.65 313.8 ;
        RECT  79.35 317.25 88.95 318.15 ;
        RECT  79.35 302.55 88.95 303.45 ;
        RECT  85.95 303.45 87.15 305.85 ;
        RECT  85.95 315.45 87.15 317.25 ;
        RECT  81.15 316.35 82.35 317.25 ;
        RECT  81.15 303.45 82.35 304.65 ;
        RECT  83.55 305.7 84.75 315.15 ;
        RECT  79.35 310.5 81.45 311.4 ;
        RECT  84.75 310.5 88.95 311.4 ;
        RECT  81.15 311.55 82.35 312.75 ;
        RECT  83.55 311.55 84.75 312.75 ;
        RECT  81.15 310.65 82.35 311.85 ;
        RECT  83.55 310.65 84.75 311.85 ;
        RECT  85.95 305.85 87.15 307.05 ;
        RECT  85.95 316.35 87.15 317.55 ;
        RECT  81.45 311.55 82.65 312.75 ;
        RECT  67.35 307.8 68.55 309.0 ;
        RECT  51.45 307.8 52.65 309.0 ;
        RECT  51.15 331.95 52.35 333.15 ;
        RECT  57.45 331.95 58.65 333.15 ;
        RECT  57.75 317.25 67.35 318.15 ;
        RECT  57.75 331.95 67.35 332.85 ;
        RECT  64.35 329.55 65.55 331.95 ;
        RECT  64.35 318.15 65.55 319.95 ;
        RECT  59.55 318.15 60.75 319.05 ;
        RECT  59.55 330.75 60.75 331.95 ;
        RECT  61.95 320.25 63.15 329.7 ;
        RECT  57.75 324.0 59.85 324.9 ;
        RECT  63.15 324.0 67.35 324.9 ;
        RECT  59.55 320.25 60.75 321.45 ;
        RECT  61.95 320.25 63.15 321.45 ;
        RECT  59.55 329.55 60.75 330.75 ;
        RECT  61.95 329.55 63.15 330.75 ;
        RECT  64.35 329.55 65.55 330.75 ;
        RECT  64.35 319.05 65.55 320.25 ;
        RECT  59.85 323.85 61.05 325.05 ;
        RECT  67.35 317.25 79.35 318.15 ;
        RECT  67.35 331.95 79.35 332.85 ;
        RECT  76.35 329.55 77.25 332.4 ;
        RECT  76.35 317.7 77.25 320.1 ;
        RECT  69.3 329.55 70.2 332.4 ;
        RECT  74.1 329.55 75.0 332.4 ;
        RECT  69.3 317.7 70.2 320.55 ;
        RECT  74.55 326.4 75.45 327.3 ;
        RECT  71.55 326.4 72.45 327.3 ;
        RECT  74.55 319.35 75.45 326.85 ;
        RECT  72.0 326.4 75.0 327.3 ;
        RECT  71.55 326.85 72.45 329.55 ;
        RECT  67.35 326.4 69.45 327.3 ;
        RECT  67.35 323.1 72.45 324.0 ;
        RECT  75.0 324.0 79.35 324.9 ;
        RECT  69.15 320.55 70.35 321.75 ;
        RECT  71.55 320.55 72.75 321.75 ;
        RECT  71.55 320.55 72.75 321.75 ;
        RECT  73.95 320.55 75.15 321.75 ;
        RECT  69.15 329.55 70.35 330.75 ;
        RECT  71.55 329.55 72.75 330.75 ;
        RECT  71.55 329.55 72.75 330.75 ;
        RECT  73.95 329.55 75.15 330.75 ;
        RECT  76.35 329.55 77.55 330.75 ;
        RECT  76.35 319.35 77.55 320.55 ;
        RECT  69.45 326.1 70.65 327.3 ;
        RECT  72.45 322.8 73.65 324.0 ;
        RECT  79.35 317.25 88.95 318.15 ;
        RECT  79.35 331.95 88.95 332.85 ;
        RECT  85.95 329.55 87.15 331.95 ;
        RECT  85.95 318.15 87.15 319.95 ;
        RECT  81.15 318.15 82.35 319.05 ;
        RECT  81.15 330.75 82.35 331.95 ;
        RECT  83.55 320.25 84.75 329.7 ;
        RECT  79.35 324.0 81.45 324.9 ;
        RECT  84.75 324.0 88.95 324.9 ;
        RECT  81.15 320.25 82.35 321.45 ;
        RECT  83.55 320.25 84.75 321.45 ;
        RECT  81.15 329.55 82.35 330.75 ;
        RECT  83.55 329.55 84.75 330.75 ;
        RECT  85.95 329.55 87.15 330.75 ;
        RECT  85.95 319.05 87.15 320.25 ;
        RECT  81.45 323.85 82.65 325.05 ;
        RECT  67.35 326.4 68.55 327.6 ;
        RECT  51.45 326.4 52.65 327.6 ;
        RECT  51.15 346.65 52.35 347.85 ;
        RECT  57.45 346.65 58.65 347.85 ;
        RECT  57.75 346.65 67.35 347.55 ;
        RECT  57.75 331.95 67.35 332.85 ;
        RECT  64.35 332.85 65.55 335.25 ;
        RECT  64.35 344.85 65.55 346.65 ;
        RECT  59.55 345.75 60.75 346.65 ;
        RECT  59.55 332.85 60.75 334.05 ;
        RECT  61.95 335.1 63.15 344.55 ;
        RECT  57.75 339.9 59.85 340.8 ;
        RECT  63.15 339.9 67.35 340.8 ;
        RECT  59.55 340.95 60.75 342.15 ;
        RECT  61.95 340.95 63.15 342.15 ;
        RECT  59.55 340.05 60.75 341.25 ;
        RECT  61.95 340.05 63.15 341.25 ;
        RECT  64.35 335.25 65.55 336.45 ;
        RECT  64.35 345.75 65.55 346.95 ;
        RECT  59.85 340.95 61.05 342.15 ;
        RECT  67.35 346.65 79.35 347.55 ;
        RECT  67.35 331.95 79.35 332.85 ;
        RECT  76.35 332.4 77.25 335.25 ;
        RECT  76.35 344.7 77.25 347.1 ;
        RECT  69.3 332.4 70.2 335.25 ;
        RECT  74.1 332.4 75.0 335.25 ;
        RECT  69.3 344.25 70.2 347.1 ;
        RECT  74.55 337.5 75.45 338.4 ;
        RECT  71.55 337.5 72.45 338.4 ;
        RECT  74.55 337.95 75.45 345.45 ;
        RECT  72.0 337.5 75.0 338.4 ;
        RECT  71.55 335.25 72.45 337.95 ;
        RECT  67.35 337.5 69.45 338.4 ;
        RECT  67.35 340.8 72.45 341.7 ;
        RECT  75.0 339.9 79.35 340.8 ;
        RECT  69.15 339.45 70.35 340.65 ;
        RECT  71.55 339.45 72.75 340.65 ;
        RECT  71.55 339.45 72.75 340.65 ;
        RECT  73.95 339.45 75.15 340.65 ;
        RECT  69.15 340.05 70.35 341.25 ;
        RECT  71.55 340.05 72.75 341.25 ;
        RECT  71.55 340.05 72.75 341.25 ;
        RECT  73.95 340.05 75.15 341.25 ;
        RECT  76.35 335.25 77.55 336.45 ;
        RECT  76.35 345.45 77.55 346.65 ;
        RECT  69.45 338.7 70.65 339.9 ;
        RECT  72.45 342.0 73.65 343.2 ;
        RECT  79.35 346.65 88.95 347.55 ;
        RECT  79.35 331.95 88.95 332.85 ;
        RECT  85.95 332.85 87.15 335.25 ;
        RECT  85.95 344.85 87.15 346.65 ;
        RECT  81.15 345.75 82.35 346.65 ;
        RECT  81.15 332.85 82.35 334.05 ;
        RECT  83.55 335.1 84.75 344.55 ;
        RECT  79.35 339.9 81.45 340.8 ;
        RECT  84.75 339.9 88.95 340.8 ;
        RECT  81.15 340.95 82.35 342.15 ;
        RECT  83.55 340.95 84.75 342.15 ;
        RECT  81.15 340.05 82.35 341.25 ;
        RECT  83.55 340.05 84.75 341.25 ;
        RECT  85.95 335.25 87.15 336.45 ;
        RECT  85.95 345.75 87.15 346.95 ;
        RECT  81.45 340.95 82.65 342.15 ;
        RECT  67.35 337.2 68.55 338.4 ;
        RECT  51.45 337.2 52.65 338.4 ;
        RECT  51.15 361.35 52.35 362.55 ;
        RECT  57.45 361.35 58.65 362.55 ;
        RECT  57.75 346.65 67.35 347.55 ;
        RECT  57.75 361.35 67.35 362.25 ;
        RECT  64.35 358.95 65.55 361.35 ;
        RECT  64.35 347.55 65.55 349.35 ;
        RECT  59.55 347.55 60.75 348.45 ;
        RECT  59.55 360.15 60.75 361.35 ;
        RECT  61.95 349.65 63.15 359.1 ;
        RECT  57.75 353.4 59.85 354.3 ;
        RECT  63.15 353.4 67.35 354.3 ;
        RECT  59.55 349.65 60.75 350.85 ;
        RECT  61.95 349.65 63.15 350.85 ;
        RECT  59.55 358.95 60.75 360.15 ;
        RECT  61.95 358.95 63.15 360.15 ;
        RECT  64.35 358.95 65.55 360.15 ;
        RECT  64.35 348.45 65.55 349.65 ;
        RECT  59.85 353.25 61.05 354.45 ;
        RECT  67.35 346.65 79.35 347.55 ;
        RECT  67.35 361.35 79.35 362.25 ;
        RECT  76.35 358.95 77.25 361.8 ;
        RECT  76.35 347.1 77.25 349.5 ;
        RECT  69.3 358.95 70.2 361.8 ;
        RECT  74.1 358.95 75.0 361.8 ;
        RECT  69.3 347.1 70.2 349.95 ;
        RECT  74.55 355.8 75.45 356.7 ;
        RECT  71.55 355.8 72.45 356.7 ;
        RECT  74.55 348.75 75.45 356.25 ;
        RECT  72.0 355.8 75.0 356.7 ;
        RECT  71.55 356.25 72.45 358.95 ;
        RECT  67.35 355.8 69.45 356.7 ;
        RECT  67.35 352.5 72.45 353.4 ;
        RECT  75.0 353.4 79.35 354.3 ;
        RECT  69.15 349.95 70.35 351.15 ;
        RECT  71.55 349.95 72.75 351.15 ;
        RECT  71.55 349.95 72.75 351.15 ;
        RECT  73.95 349.95 75.15 351.15 ;
        RECT  69.15 358.95 70.35 360.15 ;
        RECT  71.55 358.95 72.75 360.15 ;
        RECT  71.55 358.95 72.75 360.15 ;
        RECT  73.95 358.95 75.15 360.15 ;
        RECT  76.35 358.95 77.55 360.15 ;
        RECT  76.35 348.75 77.55 349.95 ;
        RECT  69.45 355.5 70.65 356.7 ;
        RECT  72.45 352.2 73.65 353.4 ;
        RECT  79.35 346.65 88.95 347.55 ;
        RECT  79.35 361.35 88.95 362.25 ;
        RECT  85.95 358.95 87.15 361.35 ;
        RECT  85.95 347.55 87.15 349.35 ;
        RECT  81.15 347.55 82.35 348.45 ;
        RECT  81.15 360.15 82.35 361.35 ;
        RECT  83.55 349.65 84.75 359.1 ;
        RECT  79.35 353.4 81.45 354.3 ;
        RECT  84.75 353.4 88.95 354.3 ;
        RECT  81.15 349.65 82.35 350.85 ;
        RECT  83.55 349.65 84.75 350.85 ;
        RECT  81.15 358.95 82.35 360.15 ;
        RECT  83.55 358.95 84.75 360.15 ;
        RECT  85.95 358.95 87.15 360.15 ;
        RECT  85.95 348.45 87.15 349.65 ;
        RECT  81.45 353.25 82.65 354.45 ;
        RECT  67.35 355.8 68.55 357.0 ;
        RECT  51.45 355.8 52.65 357.0 ;
        RECT  51.15 376.05 52.35 377.25 ;
        RECT  57.45 376.05 58.65 377.25 ;
        RECT  57.75 376.05 67.35 376.95 ;
        RECT  57.75 361.35 67.35 362.25 ;
        RECT  64.35 362.25 65.55 364.65 ;
        RECT  64.35 374.25 65.55 376.05 ;
        RECT  59.55 375.15 60.75 376.05 ;
        RECT  59.55 362.25 60.75 363.45 ;
        RECT  61.95 364.5 63.15 373.95 ;
        RECT  57.75 369.3 59.85 370.2 ;
        RECT  63.15 369.3 67.35 370.2 ;
        RECT  59.55 370.35 60.75 371.55 ;
        RECT  61.95 370.35 63.15 371.55 ;
        RECT  59.55 369.45 60.75 370.65 ;
        RECT  61.95 369.45 63.15 370.65 ;
        RECT  64.35 364.65 65.55 365.85 ;
        RECT  64.35 375.15 65.55 376.35 ;
        RECT  59.85 370.35 61.05 371.55 ;
        RECT  67.35 376.05 79.35 376.95 ;
        RECT  67.35 361.35 79.35 362.25 ;
        RECT  76.35 361.8 77.25 364.65 ;
        RECT  76.35 374.1 77.25 376.5 ;
        RECT  69.3 361.8 70.2 364.65 ;
        RECT  74.1 361.8 75.0 364.65 ;
        RECT  69.3 373.65 70.2 376.5 ;
        RECT  74.55 366.9 75.45 367.8 ;
        RECT  71.55 366.9 72.45 367.8 ;
        RECT  74.55 367.35 75.45 374.85 ;
        RECT  72.0 366.9 75.0 367.8 ;
        RECT  71.55 364.65 72.45 367.35 ;
        RECT  67.35 366.9 69.45 367.8 ;
        RECT  67.35 370.2 72.45 371.1 ;
        RECT  75.0 369.3 79.35 370.2 ;
        RECT  69.15 368.85 70.35 370.05 ;
        RECT  71.55 368.85 72.75 370.05 ;
        RECT  71.55 368.85 72.75 370.05 ;
        RECT  73.95 368.85 75.15 370.05 ;
        RECT  69.15 369.45 70.35 370.65 ;
        RECT  71.55 369.45 72.75 370.65 ;
        RECT  71.55 369.45 72.75 370.65 ;
        RECT  73.95 369.45 75.15 370.65 ;
        RECT  76.35 364.65 77.55 365.85 ;
        RECT  76.35 374.85 77.55 376.05 ;
        RECT  69.45 368.1 70.65 369.3 ;
        RECT  72.45 371.4 73.65 372.6 ;
        RECT  79.35 376.05 88.95 376.95 ;
        RECT  79.35 361.35 88.95 362.25 ;
        RECT  85.95 362.25 87.15 364.65 ;
        RECT  85.95 374.25 87.15 376.05 ;
        RECT  81.15 375.15 82.35 376.05 ;
        RECT  81.15 362.25 82.35 363.45 ;
        RECT  83.55 364.5 84.75 373.95 ;
        RECT  79.35 369.3 81.45 370.2 ;
        RECT  84.75 369.3 88.95 370.2 ;
        RECT  81.15 370.35 82.35 371.55 ;
        RECT  83.55 370.35 84.75 371.55 ;
        RECT  81.15 369.45 82.35 370.65 ;
        RECT  83.55 369.45 84.75 370.65 ;
        RECT  85.95 364.65 87.15 365.85 ;
        RECT  85.95 375.15 87.15 376.35 ;
        RECT  81.45 370.35 82.65 371.55 ;
        RECT  67.35 366.6 68.55 367.8 ;
        RECT  51.45 366.6 52.65 367.8 ;
        RECT  51.15 390.75 52.35 391.95 ;
        RECT  57.45 390.75 58.65 391.95 ;
        RECT  57.75 376.05 67.35 376.95 ;
        RECT  57.75 390.75 67.35 391.65 ;
        RECT  64.35 388.35 65.55 390.75 ;
        RECT  64.35 376.95 65.55 378.75 ;
        RECT  59.55 376.95 60.75 377.85 ;
        RECT  59.55 389.55 60.75 390.75 ;
        RECT  61.95 379.05 63.15 388.5 ;
        RECT  57.75 382.8 59.85 383.7 ;
        RECT  63.15 382.8 67.35 383.7 ;
        RECT  59.55 379.05 60.75 380.25 ;
        RECT  61.95 379.05 63.15 380.25 ;
        RECT  59.55 388.35 60.75 389.55 ;
        RECT  61.95 388.35 63.15 389.55 ;
        RECT  64.35 388.35 65.55 389.55 ;
        RECT  64.35 377.85 65.55 379.05 ;
        RECT  59.85 382.65 61.05 383.85 ;
        RECT  67.35 376.05 79.35 376.95 ;
        RECT  67.35 390.75 79.35 391.65 ;
        RECT  76.35 388.35 77.25 391.2 ;
        RECT  76.35 376.5 77.25 378.9 ;
        RECT  69.3 388.35 70.2 391.2 ;
        RECT  74.1 388.35 75.0 391.2 ;
        RECT  69.3 376.5 70.2 379.35 ;
        RECT  74.55 385.2 75.45 386.1 ;
        RECT  71.55 385.2 72.45 386.1 ;
        RECT  74.55 378.15 75.45 385.65 ;
        RECT  72.0 385.2 75.0 386.1 ;
        RECT  71.55 385.65 72.45 388.35 ;
        RECT  67.35 385.2 69.45 386.1 ;
        RECT  67.35 381.9 72.45 382.8 ;
        RECT  75.0 382.8 79.35 383.7 ;
        RECT  69.15 379.35 70.35 380.55 ;
        RECT  71.55 379.35 72.75 380.55 ;
        RECT  71.55 379.35 72.75 380.55 ;
        RECT  73.95 379.35 75.15 380.55 ;
        RECT  69.15 388.35 70.35 389.55 ;
        RECT  71.55 388.35 72.75 389.55 ;
        RECT  71.55 388.35 72.75 389.55 ;
        RECT  73.95 388.35 75.15 389.55 ;
        RECT  76.35 388.35 77.55 389.55 ;
        RECT  76.35 378.15 77.55 379.35 ;
        RECT  69.45 384.9 70.65 386.1 ;
        RECT  72.45 381.6 73.65 382.8 ;
        RECT  79.35 376.05 88.95 376.95 ;
        RECT  79.35 390.75 88.95 391.65 ;
        RECT  85.95 388.35 87.15 390.75 ;
        RECT  85.95 376.95 87.15 378.75 ;
        RECT  81.15 376.95 82.35 377.85 ;
        RECT  81.15 389.55 82.35 390.75 ;
        RECT  83.55 379.05 84.75 388.5 ;
        RECT  79.35 382.8 81.45 383.7 ;
        RECT  84.75 382.8 88.95 383.7 ;
        RECT  81.15 379.05 82.35 380.25 ;
        RECT  83.55 379.05 84.75 380.25 ;
        RECT  81.15 388.35 82.35 389.55 ;
        RECT  83.55 388.35 84.75 389.55 ;
        RECT  85.95 388.35 87.15 389.55 ;
        RECT  85.95 377.85 87.15 379.05 ;
        RECT  81.45 382.65 82.65 383.85 ;
        RECT  67.35 385.2 68.55 386.4 ;
        RECT  51.45 385.2 52.65 386.4 ;
        RECT  51.15 405.45 52.35 406.65 ;
        RECT  57.45 405.45 58.65 406.65 ;
        RECT  57.75 405.45 67.35 406.35 ;
        RECT  57.75 390.75 67.35 391.65 ;
        RECT  64.35 391.65 65.55 394.05 ;
        RECT  64.35 403.65 65.55 405.45 ;
        RECT  59.55 404.55 60.75 405.45 ;
        RECT  59.55 391.65 60.75 392.85 ;
        RECT  61.95 393.9 63.15 403.35 ;
        RECT  57.75 398.7 59.85 399.6 ;
        RECT  63.15 398.7 67.35 399.6 ;
        RECT  59.55 399.75 60.75 400.95 ;
        RECT  61.95 399.75 63.15 400.95 ;
        RECT  59.55 398.85 60.75 400.05 ;
        RECT  61.95 398.85 63.15 400.05 ;
        RECT  64.35 394.05 65.55 395.25 ;
        RECT  64.35 404.55 65.55 405.75 ;
        RECT  59.85 399.75 61.05 400.95 ;
        RECT  67.35 405.45 79.35 406.35 ;
        RECT  67.35 390.75 79.35 391.65 ;
        RECT  76.35 391.2 77.25 394.05 ;
        RECT  76.35 403.5 77.25 405.9 ;
        RECT  69.3 391.2 70.2 394.05 ;
        RECT  74.1 391.2 75.0 394.05 ;
        RECT  69.3 403.05 70.2 405.9 ;
        RECT  74.55 396.3 75.45 397.2 ;
        RECT  71.55 396.3 72.45 397.2 ;
        RECT  74.55 396.75 75.45 404.25 ;
        RECT  72.0 396.3 75.0 397.2 ;
        RECT  71.55 394.05 72.45 396.75 ;
        RECT  67.35 396.3 69.45 397.2 ;
        RECT  67.35 399.6 72.45 400.5 ;
        RECT  75.0 398.7 79.35 399.6 ;
        RECT  69.15 398.25 70.35 399.45 ;
        RECT  71.55 398.25 72.75 399.45 ;
        RECT  71.55 398.25 72.75 399.45 ;
        RECT  73.95 398.25 75.15 399.45 ;
        RECT  69.15 398.85 70.35 400.05 ;
        RECT  71.55 398.85 72.75 400.05 ;
        RECT  71.55 398.85 72.75 400.05 ;
        RECT  73.95 398.85 75.15 400.05 ;
        RECT  76.35 394.05 77.55 395.25 ;
        RECT  76.35 404.25 77.55 405.45 ;
        RECT  69.45 397.5 70.65 398.7 ;
        RECT  72.45 400.8 73.65 402.0 ;
        RECT  79.35 405.45 88.95 406.35 ;
        RECT  79.35 390.75 88.95 391.65 ;
        RECT  85.95 391.65 87.15 394.05 ;
        RECT  85.95 403.65 87.15 405.45 ;
        RECT  81.15 404.55 82.35 405.45 ;
        RECT  81.15 391.65 82.35 392.85 ;
        RECT  83.55 393.9 84.75 403.35 ;
        RECT  79.35 398.7 81.45 399.6 ;
        RECT  84.75 398.7 88.95 399.6 ;
        RECT  81.15 399.75 82.35 400.95 ;
        RECT  83.55 399.75 84.75 400.95 ;
        RECT  81.15 398.85 82.35 400.05 ;
        RECT  83.55 398.85 84.75 400.05 ;
        RECT  85.95 394.05 87.15 395.25 ;
        RECT  85.95 404.55 87.15 405.75 ;
        RECT  81.45 399.75 82.65 400.95 ;
        RECT  67.35 396.0 68.55 397.2 ;
        RECT  51.45 396.0 52.65 397.2 ;
        RECT  51.15 420.15 52.35 421.35 ;
        RECT  57.45 420.15 58.65 421.35 ;
        RECT  57.75 405.45 67.35 406.35 ;
        RECT  57.75 420.15 67.35 421.05 ;
        RECT  64.35 417.75 65.55 420.15 ;
        RECT  64.35 406.35 65.55 408.15 ;
        RECT  59.55 406.35 60.75 407.25 ;
        RECT  59.55 418.95 60.75 420.15 ;
        RECT  61.95 408.45 63.15 417.9 ;
        RECT  57.75 412.2 59.85 413.1 ;
        RECT  63.15 412.2 67.35 413.1 ;
        RECT  59.55 408.45 60.75 409.65 ;
        RECT  61.95 408.45 63.15 409.65 ;
        RECT  59.55 417.75 60.75 418.95 ;
        RECT  61.95 417.75 63.15 418.95 ;
        RECT  64.35 417.75 65.55 418.95 ;
        RECT  64.35 407.25 65.55 408.45 ;
        RECT  59.85 412.05 61.05 413.25 ;
        RECT  67.35 405.45 79.35 406.35 ;
        RECT  67.35 420.15 79.35 421.05 ;
        RECT  76.35 417.75 77.25 420.6 ;
        RECT  76.35 405.9 77.25 408.3 ;
        RECT  69.3 417.75 70.2 420.6 ;
        RECT  74.1 417.75 75.0 420.6 ;
        RECT  69.3 405.9 70.2 408.75 ;
        RECT  74.55 414.6 75.45 415.5 ;
        RECT  71.55 414.6 72.45 415.5 ;
        RECT  74.55 407.55 75.45 415.05 ;
        RECT  72.0 414.6 75.0 415.5 ;
        RECT  71.55 415.05 72.45 417.75 ;
        RECT  67.35 414.6 69.45 415.5 ;
        RECT  67.35 411.3 72.45 412.2 ;
        RECT  75.0 412.2 79.35 413.1 ;
        RECT  69.15 408.75 70.35 409.95 ;
        RECT  71.55 408.75 72.75 409.95 ;
        RECT  71.55 408.75 72.75 409.95 ;
        RECT  73.95 408.75 75.15 409.95 ;
        RECT  69.15 417.75 70.35 418.95 ;
        RECT  71.55 417.75 72.75 418.95 ;
        RECT  71.55 417.75 72.75 418.95 ;
        RECT  73.95 417.75 75.15 418.95 ;
        RECT  76.35 417.75 77.55 418.95 ;
        RECT  76.35 407.55 77.55 408.75 ;
        RECT  69.45 414.3 70.65 415.5 ;
        RECT  72.45 411.0 73.65 412.2 ;
        RECT  79.35 405.45 88.95 406.35 ;
        RECT  79.35 420.15 88.95 421.05 ;
        RECT  85.95 417.75 87.15 420.15 ;
        RECT  85.95 406.35 87.15 408.15 ;
        RECT  81.15 406.35 82.35 407.25 ;
        RECT  81.15 418.95 82.35 420.15 ;
        RECT  83.55 408.45 84.75 417.9 ;
        RECT  79.35 412.2 81.45 413.1 ;
        RECT  84.75 412.2 88.95 413.1 ;
        RECT  81.15 408.45 82.35 409.65 ;
        RECT  83.55 408.45 84.75 409.65 ;
        RECT  81.15 417.75 82.35 418.95 ;
        RECT  83.55 417.75 84.75 418.95 ;
        RECT  85.95 417.75 87.15 418.95 ;
        RECT  85.95 407.25 87.15 408.45 ;
        RECT  81.45 412.05 82.65 413.25 ;
        RECT  67.35 414.6 68.55 415.8 ;
        RECT  51.45 414.6 52.65 415.8 ;
        RECT  51.15 434.85 52.35 436.05 ;
        RECT  57.45 434.85 58.65 436.05 ;
        RECT  57.75 434.85 67.35 435.75 ;
        RECT  57.75 420.15 67.35 421.05 ;
        RECT  64.35 421.05 65.55 423.45 ;
        RECT  64.35 433.05 65.55 434.85 ;
        RECT  59.55 433.95 60.75 434.85 ;
        RECT  59.55 421.05 60.75 422.25 ;
        RECT  61.95 423.3 63.15 432.75 ;
        RECT  57.75 428.1 59.85 429.0 ;
        RECT  63.15 428.1 67.35 429.0 ;
        RECT  59.55 429.15 60.75 430.35 ;
        RECT  61.95 429.15 63.15 430.35 ;
        RECT  59.55 428.25 60.75 429.45 ;
        RECT  61.95 428.25 63.15 429.45 ;
        RECT  64.35 423.45 65.55 424.65 ;
        RECT  64.35 433.95 65.55 435.15 ;
        RECT  59.85 429.15 61.05 430.35 ;
        RECT  67.35 434.85 79.35 435.75 ;
        RECT  67.35 420.15 79.35 421.05 ;
        RECT  76.35 420.6 77.25 423.45 ;
        RECT  76.35 432.9 77.25 435.3 ;
        RECT  69.3 420.6 70.2 423.45 ;
        RECT  74.1 420.6 75.0 423.45 ;
        RECT  69.3 432.45 70.2 435.3 ;
        RECT  74.55 425.7 75.45 426.6 ;
        RECT  71.55 425.7 72.45 426.6 ;
        RECT  74.55 426.15 75.45 433.65 ;
        RECT  72.0 425.7 75.0 426.6 ;
        RECT  71.55 423.45 72.45 426.15 ;
        RECT  67.35 425.7 69.45 426.6 ;
        RECT  67.35 429.0 72.45 429.9 ;
        RECT  75.0 428.1 79.35 429.0 ;
        RECT  69.15 427.65 70.35 428.85 ;
        RECT  71.55 427.65 72.75 428.85 ;
        RECT  71.55 427.65 72.75 428.85 ;
        RECT  73.95 427.65 75.15 428.85 ;
        RECT  69.15 428.25 70.35 429.45 ;
        RECT  71.55 428.25 72.75 429.45 ;
        RECT  71.55 428.25 72.75 429.45 ;
        RECT  73.95 428.25 75.15 429.45 ;
        RECT  76.35 423.45 77.55 424.65 ;
        RECT  76.35 433.65 77.55 434.85 ;
        RECT  69.45 426.9 70.65 428.1 ;
        RECT  72.45 430.2 73.65 431.4 ;
        RECT  79.35 434.85 88.95 435.75 ;
        RECT  79.35 420.15 88.95 421.05 ;
        RECT  85.95 421.05 87.15 423.45 ;
        RECT  85.95 433.05 87.15 434.85 ;
        RECT  81.15 433.95 82.35 434.85 ;
        RECT  81.15 421.05 82.35 422.25 ;
        RECT  83.55 423.3 84.75 432.75 ;
        RECT  79.35 428.1 81.45 429.0 ;
        RECT  84.75 428.1 88.95 429.0 ;
        RECT  81.15 429.15 82.35 430.35 ;
        RECT  83.55 429.15 84.75 430.35 ;
        RECT  81.15 428.25 82.35 429.45 ;
        RECT  83.55 428.25 84.75 429.45 ;
        RECT  85.95 423.45 87.15 424.65 ;
        RECT  85.95 433.95 87.15 435.15 ;
        RECT  81.45 429.15 82.65 430.35 ;
        RECT  67.35 425.4 68.55 426.6 ;
        RECT  51.45 425.4 52.65 426.6 ;
        RECT  17.7 39.0 18.6 79.8 ;
        RECT  72.15 39.0 73.05 79.8 ;
        RECT  72.15 69.0 73.05 80.4 ;
        RECT  68.85 79.2 72.15 80.4 ;
        RECT  70.35 71.4 71.25 78.0 ;
        RECT  70.05 75.0 70.35 78.0 ;
        RECT  70.05 71.4 70.35 72.6 ;
        RECT  67.65 76.2 68.85 80.4 ;
        RECT  67.65 69.0 68.85 72.6 ;
        RECT  64.05 79.2 67.65 80.4 ;
        RECT  66.75 73.8 67.65 75.0 ;
        RECT  66.45 72.6 66.75 75.0 ;
        RECT  65.55 71.4 66.45 78.0 ;
        RECT  65.25 76.2 65.55 78.0 ;
        RECT  65.25 71.4 65.55 72.6 ;
        RECT  62.85 76.2 64.05 80.4 ;
        RECT  49.05 79.2 62.85 80.4 ;
        RECT  62.25 73.5 64.65 74.7 ;
        RECT  64.05 69.0 67.65 69.9 ;
        RECT  62.85 69.0 64.05 72.6 ;
        RECT  61.65 69.0 62.85 70.2 ;
        RECT  59.25 76.8 60.45 78.0 ;
        RECT  60.15 73.5 61.35 75.9 ;
        RECT  58.35 71.4 59.25 78.0 ;
        RECT  58.05 76.2 58.35 78.0 ;
        RECT  58.05 71.4 58.35 72.6 ;
        RECT  55.95 71.4 56.85 78.0 ;
        RECT  55.65 76.2 55.95 78.0 ;
        RECT  55.65 71.4 55.95 73.8 ;
        RECT  53.55 71.4 54.45 78.0 ;
        RECT  53.25 76.2 53.55 78.0 ;
        RECT  53.25 71.4 53.55 73.8 ;
        RECT  51.45 73.8 52.35 75.0 ;
        RECT  50.55 71.4 51.45 78.0 ;
        RECT  50.25 75.0 50.55 78.0 ;
        RECT  50.25 71.4 50.55 72.6 ;
        RECT  47.85 76.2 49.05 80.4 ;
        RECT  43.35 79.2 47.85 80.4 ;
        RECT  46.95 74.1 49.35 75.3 ;
        RECT  49.05 69.0 61.65 69.9 ;
        RECT  47.85 69.0 49.05 72.6 ;
        RECT  45.75 76.8 46.95 78.0 ;
        RECT  44.85 71.4 45.75 78.0 ;
        RECT  44.55 76.2 44.85 78.0 ;
        RECT  44.55 71.4 44.85 72.6 ;
        RECT  43.35 69.0 47.85 69.9 ;
        RECT  42.15 76.2 43.35 80.4 ;
        RECT  38.55 79.2 42.15 80.4 ;
        RECT  41.25 73.5 42.45 74.7 ;
        RECT  42.15 69.0 43.35 72.6 ;
        RECT  40.95 72.6 41.25 78.0 ;
        RECT  40.35 71.4 40.95 78.0 ;
        RECT  39.75 76.2 40.35 78.0 ;
        RECT  40.05 71.4 40.35 73.8 ;
        RECT  39.75 71.4 40.05 72.6 ;
        RECT  37.35 76.2 38.55 80.4 ;
        RECT  22.35 79.2 37.35 80.4 ;
        RECT  36.75 73.5 39.15 74.7 ;
        RECT  38.55 69.0 42.15 69.9 ;
        RECT  37.35 69.0 38.55 72.6 ;
        RECT  36.15 69.0 37.35 70.2 ;
        RECT  32.85 76.8 34.05 78.0 ;
        RECT  33.75 73.5 34.95 75.9 ;
        RECT  31.95 71.4 32.85 78.0 ;
        RECT  31.65 76.2 31.95 78.0 ;
        RECT  31.65 71.4 31.95 72.6 ;
        RECT  29.55 71.4 30.45 78.0 ;
        RECT  29.25 76.2 29.55 78.0 ;
        RECT  29.25 71.4 29.55 73.8 ;
        RECT  27.15 71.4 28.05 78.0 ;
        RECT  26.85 76.2 27.15 78.0 ;
        RECT  26.85 71.4 27.15 73.8 ;
        RECT  25.05 73.8 25.95 75.0 ;
        RECT  24.15 71.4 25.05 78.0 ;
        RECT  23.85 75.0 24.15 78.0 ;
        RECT  23.85 71.4 24.15 72.6 ;
        RECT  22.65 69.0 36.15 69.9 ;
        RECT  22.35 76.2 22.65 78.0 ;
        RECT  21.45 76.2 22.35 80.4 ;
        RECT  21.75 69.0 22.65 72.6 ;
        RECT  21.45 71.4 21.75 72.6 ;
        RECT  19.95 76.2 21.45 77.4 ;
        RECT  19.05 74.1 19.95 75.3 ;
        RECT  18.15 69.0 19.05 80.4 ;
        RECT  72.15 58.8 73.05 70.2 ;
        RECT  68.85 58.8 72.15 60.0 ;
        RECT  70.35 61.2 71.25 67.8 ;
        RECT  70.05 61.2 70.35 64.2 ;
        RECT  70.05 66.6 70.35 67.8 ;
        RECT  67.65 58.8 68.85 63.0 ;
        RECT  67.65 66.6 68.85 70.2 ;
        RECT  64.05 58.8 67.65 60.0 ;
        RECT  66.75 64.2 67.65 65.4 ;
        RECT  66.45 64.2 66.75 66.6 ;
        RECT  65.55 61.2 66.45 67.8 ;
        RECT  65.25 61.2 65.55 63.0 ;
        RECT  65.25 66.6 65.55 67.8 ;
        RECT  62.85 58.8 64.05 63.0 ;
        RECT  49.05 58.8 62.85 60.0 ;
        RECT  62.25 64.5 64.65 65.7 ;
        RECT  64.05 69.3 67.65 70.2 ;
        RECT  62.85 66.6 64.05 70.2 ;
        RECT  61.65 69.0 62.85 70.2 ;
        RECT  59.25 61.2 60.45 62.4 ;
        RECT  60.15 63.3 61.35 65.7 ;
        RECT  58.35 61.2 59.25 67.8 ;
        RECT  58.05 61.2 58.35 63.0 ;
        RECT  58.05 66.6 58.35 67.8 ;
        RECT  55.95 61.2 56.85 67.8 ;
        RECT  55.65 61.2 55.95 63.0 ;
        RECT  55.65 65.4 55.95 67.8 ;
        RECT  53.55 61.2 54.45 67.8 ;
        RECT  53.25 61.2 53.55 63.0 ;
        RECT  53.25 65.4 53.55 67.8 ;
        RECT  51.45 64.2 52.35 65.4 ;
        RECT  50.55 61.2 51.45 67.8 ;
        RECT  50.25 61.2 50.55 64.2 ;
        RECT  50.25 66.6 50.55 67.8 ;
        RECT  47.85 58.8 49.05 63.0 ;
        RECT  43.35 58.8 47.85 60.0 ;
        RECT  46.95 63.9 49.35 65.1 ;
        RECT  49.05 69.3 61.65 70.2 ;
        RECT  47.85 66.6 49.05 70.2 ;
        RECT  45.75 61.2 46.95 62.4 ;
        RECT  44.85 61.2 45.75 67.8 ;
        RECT  44.55 61.2 44.85 63.0 ;
        RECT  44.55 66.6 44.85 67.8 ;
        RECT  43.35 69.3 47.85 70.2 ;
        RECT  42.15 58.8 43.35 63.0 ;
        RECT  38.55 58.8 42.15 60.0 ;
        RECT  41.25 64.5 42.45 65.7 ;
        RECT  42.15 66.6 43.35 70.2 ;
        RECT  40.95 61.2 41.25 66.6 ;
        RECT  40.35 61.2 40.95 67.8 ;
        RECT  39.75 61.2 40.35 63.0 ;
        RECT  40.05 65.4 40.35 67.8 ;
        RECT  39.75 66.6 40.05 67.8 ;
        RECT  37.35 58.8 38.55 63.0 ;
        RECT  22.35 58.8 37.35 60.0 ;
        RECT  36.75 64.5 39.15 65.7 ;
        RECT  38.55 69.3 42.15 70.2 ;
        RECT  37.35 66.6 38.55 70.2 ;
        RECT  36.15 69.0 37.35 70.2 ;
        RECT  32.85 61.2 34.05 62.4 ;
        RECT  33.75 63.3 34.95 65.7 ;
        RECT  31.95 61.2 32.85 67.8 ;
        RECT  31.65 61.2 31.95 63.0 ;
        RECT  31.65 66.6 31.95 67.8 ;
        RECT  29.55 61.2 30.45 67.8 ;
        RECT  29.25 61.2 29.55 63.0 ;
        RECT  29.25 65.4 29.55 67.8 ;
        RECT  27.15 61.2 28.05 67.8 ;
        RECT  26.85 61.2 27.15 63.0 ;
        RECT  26.85 65.4 27.15 67.8 ;
        RECT  25.05 64.2 25.95 65.4 ;
        RECT  24.15 61.2 25.05 67.8 ;
        RECT  23.85 61.2 24.15 64.2 ;
        RECT  23.85 66.6 24.15 67.8 ;
        RECT  22.65 69.3 36.15 70.2 ;
        RECT  22.35 61.2 22.65 63.0 ;
        RECT  21.45 58.8 22.35 63.0 ;
        RECT  21.75 66.6 22.65 70.2 ;
        RECT  21.45 66.6 21.75 67.8 ;
        RECT  19.95 61.8 21.45 63.0 ;
        RECT  19.05 63.9 19.95 65.1 ;
        RECT  18.15 58.8 19.05 70.2 ;
        RECT  72.15 48.6 73.05 60.0 ;
        RECT  68.85 58.8 72.15 60.0 ;
        RECT  70.35 51.0 71.25 57.6 ;
        RECT  70.05 54.6 70.35 57.6 ;
        RECT  70.05 51.0 70.35 52.2 ;
        RECT  67.65 55.8 68.85 60.0 ;
        RECT  67.65 48.6 68.85 52.2 ;
        RECT  64.05 58.8 67.65 60.0 ;
        RECT  66.75 53.4 67.65 54.6 ;
        RECT  66.45 52.2 66.75 54.6 ;
        RECT  65.55 51.0 66.45 57.6 ;
        RECT  65.25 55.8 65.55 57.6 ;
        RECT  65.25 51.0 65.55 52.2 ;
        RECT  62.85 55.8 64.05 60.0 ;
        RECT  49.05 58.8 62.85 60.0 ;
        RECT  62.25 53.1 64.65 54.3 ;
        RECT  64.05 48.6 67.65 49.5 ;
        RECT  62.85 48.6 64.05 52.2 ;
        RECT  61.65 48.6 62.85 49.8 ;
        RECT  59.25 56.4 60.45 57.6 ;
        RECT  60.15 53.1 61.35 55.5 ;
        RECT  58.35 51.0 59.25 57.6 ;
        RECT  58.05 55.8 58.35 57.6 ;
        RECT  58.05 51.0 58.35 52.2 ;
        RECT  55.95 51.0 56.85 57.6 ;
        RECT  55.65 55.8 55.95 57.6 ;
        RECT  55.65 51.0 55.95 53.4 ;
        RECT  53.55 51.0 54.45 57.6 ;
        RECT  53.25 55.8 53.55 57.6 ;
        RECT  53.25 51.0 53.55 53.4 ;
        RECT  51.45 53.4 52.35 54.6 ;
        RECT  50.55 51.0 51.45 57.6 ;
        RECT  50.25 54.6 50.55 57.6 ;
        RECT  50.25 51.0 50.55 52.2 ;
        RECT  47.85 55.8 49.05 60.0 ;
        RECT  43.35 58.8 47.85 60.0 ;
        RECT  46.95 53.7 49.35 54.9 ;
        RECT  49.05 48.6 61.65 49.5 ;
        RECT  47.85 48.6 49.05 52.2 ;
        RECT  45.75 56.4 46.95 57.6 ;
        RECT  44.85 51.0 45.75 57.6 ;
        RECT  44.55 55.8 44.85 57.6 ;
        RECT  44.55 51.0 44.85 52.2 ;
        RECT  43.35 48.6 47.85 49.5 ;
        RECT  42.15 55.8 43.35 60.0 ;
        RECT  38.55 58.8 42.15 60.0 ;
        RECT  41.25 53.1 42.45 54.3 ;
        RECT  42.15 48.6 43.35 52.2 ;
        RECT  40.95 52.2 41.25 57.6 ;
        RECT  40.35 51.0 40.95 57.6 ;
        RECT  39.75 55.8 40.35 57.6 ;
        RECT  40.05 51.0 40.35 53.4 ;
        RECT  39.75 51.0 40.05 52.2 ;
        RECT  37.35 55.8 38.55 60.0 ;
        RECT  22.35 58.8 37.35 60.0 ;
        RECT  36.75 53.1 39.15 54.3 ;
        RECT  38.55 48.6 42.15 49.5 ;
        RECT  37.35 48.6 38.55 52.2 ;
        RECT  36.15 48.6 37.35 49.8 ;
        RECT  32.85 56.4 34.05 57.6 ;
        RECT  33.75 53.1 34.95 55.5 ;
        RECT  31.95 51.0 32.85 57.6 ;
        RECT  31.65 55.8 31.95 57.6 ;
        RECT  31.65 51.0 31.95 52.2 ;
        RECT  29.55 51.0 30.45 57.6 ;
        RECT  29.25 55.8 29.55 57.6 ;
        RECT  29.25 51.0 29.55 53.4 ;
        RECT  27.15 51.0 28.05 57.6 ;
        RECT  26.85 55.8 27.15 57.6 ;
        RECT  26.85 51.0 27.15 53.4 ;
        RECT  25.05 53.4 25.95 54.6 ;
        RECT  24.15 51.0 25.05 57.6 ;
        RECT  23.85 54.6 24.15 57.6 ;
        RECT  23.85 51.0 24.15 52.2 ;
        RECT  22.65 48.6 36.15 49.5 ;
        RECT  22.35 55.8 22.65 57.6 ;
        RECT  21.45 55.8 22.35 60.0 ;
        RECT  21.75 48.6 22.65 52.2 ;
        RECT  21.45 51.0 21.75 52.2 ;
        RECT  19.95 55.8 21.45 57.0 ;
        RECT  19.05 53.7 19.95 54.9 ;
        RECT  18.15 48.6 19.05 60.0 ;
        RECT  72.15 38.4 73.05 49.8 ;
        RECT  68.85 38.4 72.15 39.6 ;
        RECT  70.35 40.8 71.25 47.4 ;
        RECT  70.05 40.8 70.35 43.8 ;
        RECT  70.05 46.2 70.35 47.4 ;
        RECT  67.65 38.4 68.85 42.6 ;
        RECT  67.65 46.2 68.85 49.8 ;
        RECT  64.05 38.4 67.65 39.6 ;
        RECT  66.75 43.8 67.65 45.0 ;
        RECT  66.45 43.8 66.75 46.2 ;
        RECT  65.55 40.8 66.45 47.4 ;
        RECT  65.25 40.8 65.55 42.6 ;
        RECT  65.25 46.2 65.55 47.4 ;
        RECT  62.85 38.4 64.05 42.6 ;
        RECT  49.05 38.4 62.85 39.6 ;
        RECT  62.25 44.1 64.65 45.3 ;
        RECT  64.05 48.9 67.65 49.8 ;
        RECT  62.85 46.2 64.05 49.8 ;
        RECT  61.65 48.6 62.85 49.8 ;
        RECT  59.25 40.8 60.45 42.0 ;
        RECT  60.15 42.9 61.35 45.3 ;
        RECT  58.35 40.8 59.25 47.4 ;
        RECT  58.05 40.8 58.35 42.6 ;
        RECT  58.05 46.2 58.35 47.4 ;
        RECT  55.95 40.8 56.85 47.4 ;
        RECT  55.65 40.8 55.95 42.6 ;
        RECT  55.65 45.0 55.95 47.4 ;
        RECT  53.55 40.8 54.45 47.4 ;
        RECT  53.25 40.8 53.55 42.6 ;
        RECT  53.25 45.0 53.55 47.4 ;
        RECT  51.45 43.8 52.35 45.0 ;
        RECT  50.55 40.8 51.45 47.4 ;
        RECT  50.25 40.8 50.55 43.8 ;
        RECT  50.25 46.2 50.55 47.4 ;
        RECT  47.85 38.4 49.05 42.6 ;
        RECT  43.35 38.4 47.85 39.6 ;
        RECT  46.95 43.5 49.35 44.7 ;
        RECT  49.05 48.9 61.65 49.8 ;
        RECT  47.85 46.2 49.05 49.8 ;
        RECT  45.75 40.8 46.95 42.0 ;
        RECT  44.85 40.8 45.75 47.4 ;
        RECT  44.55 40.8 44.85 42.6 ;
        RECT  44.55 46.2 44.85 47.4 ;
        RECT  43.35 48.9 47.85 49.8 ;
        RECT  42.15 38.4 43.35 42.6 ;
        RECT  38.55 38.4 42.15 39.6 ;
        RECT  41.25 44.1 42.45 45.3 ;
        RECT  42.15 46.2 43.35 49.8 ;
        RECT  40.95 40.8 41.25 46.2 ;
        RECT  40.35 40.8 40.95 47.4 ;
        RECT  39.75 40.8 40.35 42.6 ;
        RECT  40.05 45.0 40.35 47.4 ;
        RECT  39.75 46.2 40.05 47.4 ;
        RECT  37.35 38.4 38.55 42.6 ;
        RECT  22.35 38.4 37.35 39.6 ;
        RECT  36.75 44.1 39.15 45.3 ;
        RECT  38.55 48.9 42.15 49.8 ;
        RECT  37.35 46.2 38.55 49.8 ;
        RECT  36.15 48.6 37.35 49.8 ;
        RECT  32.85 40.8 34.05 42.0 ;
        RECT  33.75 42.9 34.95 45.3 ;
        RECT  31.95 40.8 32.85 47.4 ;
        RECT  31.65 40.8 31.95 42.6 ;
        RECT  31.65 46.2 31.95 47.4 ;
        RECT  29.55 40.8 30.45 47.4 ;
        RECT  29.25 40.8 29.55 42.6 ;
        RECT  29.25 45.0 29.55 47.4 ;
        RECT  27.15 40.8 28.05 47.4 ;
        RECT  26.85 40.8 27.15 42.6 ;
        RECT  26.85 45.0 27.15 47.4 ;
        RECT  25.05 43.8 25.95 45.0 ;
        RECT  24.15 40.8 25.05 47.4 ;
        RECT  23.85 40.8 24.15 43.8 ;
        RECT  23.85 46.2 24.15 47.4 ;
        RECT  22.65 48.9 36.15 49.8 ;
        RECT  22.35 40.8 22.65 42.6 ;
        RECT  21.45 38.4 22.35 42.6 ;
        RECT  21.75 46.2 22.65 49.8 ;
        RECT  21.45 46.2 21.75 47.4 ;
        RECT  19.95 41.4 21.45 42.6 ;
        RECT  19.05 43.5 19.95 44.7 ;
        RECT  18.15 38.4 19.05 49.8 ;
        RECT  91.05 88.8 92.25 90.0 ;
        RECT  88.35 104.7 89.55 105.9 ;
        RECT  85.65 147.6 86.85 148.8 ;
        RECT  82.95 163.5 84.15 164.7 ;
        RECT  114.45 33.3 115.65 34.5 ;
        RECT  109.05 28.65 110.25 29.85 ;
        RECT  111.75 26.25 112.95 27.45 ;
        RECT  114.45 446.4 115.65 447.6 ;
        RECT  117.15 97.95 118.35 99.15 ;
        RECT  119.85 196.05 121.05 197.25 ;
        RECT  16.95 76.5 18.15 77.7 ;
        RECT  106.35 456.6 107.55 457.8 ;
        RECT  95.55 437.1 97.95 438.3 ;
        RECT  134.25 437.1 135.45 438.3 ;
        RECT  144.45 437.1 145.65 438.3 ;
        RECT  123.15 437.1 124.35 438.3 ;
        RECT  102.15 8.1 104.55 9.3 ;
        RECT  133.95 8.1 135.15 9.3 ;
        RECT  133.95 8.1 135.15 9.3 ;
        RECT  88.2 229.05 89.4 230.25 ;
        RECT  88.2 258.45 89.4 259.65 ;
        RECT  88.2 287.85 89.4 289.05 ;
        RECT  88.2 317.25 89.4 318.45 ;
        RECT  88.2 346.65 89.4 347.85 ;
        RECT  88.2 376.05 89.4 377.25 ;
        RECT  88.2 405.45 89.4 406.65 ;
        RECT  88.2 434.85 89.4 436.05 ;
        RECT  95.55 140.55 97.95 141.75 ;
        RECT  95.55 199.35 97.95 200.55 ;
        RECT  75.45 69.15 76.65 70.35 ;
        RECT  95.55 69.15 97.95 70.35 ;
        RECT  75.45 69.15 76.65 70.35 ;
        RECT  95.55 69.15 97.95 70.35 ;
        RECT  75.45 48.75 76.65 49.95 ;
        RECT  95.55 48.75 97.95 49.95 ;
        RECT  75.45 48.75 76.65 49.95 ;
        RECT  95.55 48.75 97.95 49.95 ;
        RECT  -30.6 180.0 -28.95 180.9 ;
        RECT  -44.85 180.0 -43.2 180.9 ;
        RECT  -40.5 145.5 -39.6 151.8 ;
        RECT  -43.95 145.5 -43.05 154.5 ;
        RECT  -64.35 145.5 -63.45 157.2 ;
        RECT  -48.75 145.5 -47.85 159.9 ;
        RECT  -17.1 153.6 -16.2 164.4 ;
        RECT  -13.8 161.7 -12.9 164.4 ;
        RECT  -27.15 161.7 -26.25 164.4 ;
        RECT  -32.7 153.6 -31.8 164.4 ;
        RECT  -34.5 156.3 -33.6 164.4 ;
        RECT  -47.55 161.7 -46.65 164.4 ;
        RECT  -42.0 159.0 -41.1 164.4 ;
        RECT  -40.2 156.3 -39.3 164.4 ;
        RECT  -16.05 119.7 -15.15 121.5 ;
        RECT  -5.7 121.5 -4.8 151.35 ;
        RECT  -14.7 145.95 -13.8 146.85 ;
        RECT  -13.8 145.95 -12.9 146.85 ;
        RECT  -14.7 145.5 -13.8 146.4 ;
        RECT  -14.25 145.95 -13.35 146.85 ;
        RECT  -13.8 146.4 -12.9 164.4 ;
        RECT  -30.6 189.6 -29.7 215.1 ;
        RECT  -44.1 208.8 -43.2 212.4 ;
        RECT  -14.7 199.2 -13.8 217.8 ;
        RECT  -3.9 214.65 -3.0 265.8 ;
        RECT  -7.95 265.35 -3.0 266.25 ;
        RECT  -22.65 88.5 -21.75 223.5 ;
        RECT  -52.05 180.0 -51.15 220.5 ;
        RECT  -66.3 141.9 -21.75 142.8 ;
        RECT  -7.95 88.5 -7.05 233.4 ;
        RECT  -37.35 180.0 -36.45 231.3 ;
        RECT  -14.7 126.9 -13.8 128.7 ;
        RECT  -27.6 85.5 -26.7 126.9 ;
        RECT  -61.2 87.9 -27.15 88.8 ;
        RECT  -14.7 123.75 -13.8 124.65 ;
        RECT  -14.1 123.75 -13.2 124.65 ;
        RECT  -14.7 124.2 -13.8 126.9 ;
        RECT  -14.25 123.75 -13.65 124.65 ;
        RECT  -14.1 119.7 -13.2 124.2 ;
        RECT  -66.3 87.45 -35.7 88.35 ;
        RECT  -66.3 141.9 -35.7 142.8 ;
        RECT  -66.9 141.9 -55.5 142.8 ;
        RECT  -66.9 138.6 -65.7 141.9 ;
        RECT  -64.5 140.1 -57.9 141.0 ;
        RECT  -64.5 139.8 -61.5 140.1 ;
        RECT  -59.1 139.8 -57.9 140.1 ;
        RECT  -66.9 137.4 -62.7 138.6 ;
        RECT  -59.1 137.4 -55.5 138.6 ;
        RECT  -66.9 133.8 -65.7 137.4 ;
        RECT  -61.5 136.5 -60.3 137.4 ;
        RECT  -61.5 136.2 -59.1 136.5 ;
        RECT  -64.5 135.3 -57.9 136.2 ;
        RECT  -64.5 135.0 -62.7 135.3 ;
        RECT  -59.1 135.0 -57.9 135.3 ;
        RECT  -66.9 132.6 -62.7 133.8 ;
        RECT  -66.9 118.8 -65.7 132.6 ;
        RECT  -61.2 132.0 -60.0 134.4 ;
        RECT  -56.4 133.8 -55.5 137.4 ;
        RECT  -59.1 132.6 -55.5 133.8 ;
        RECT  -56.7 131.4 -55.5 132.6 ;
        RECT  -64.5 129.0 -63.3 130.2 ;
        RECT  -62.4 129.9 -60.0 131.1 ;
        RECT  -64.5 128.1 -57.9 129.0 ;
        RECT  -64.5 127.8 -62.7 128.1 ;
        RECT  -59.1 127.8 -57.9 128.1 ;
        RECT  -64.5 125.7 -57.9 126.6 ;
        RECT  -64.5 125.4 -62.7 125.7 ;
        RECT  -60.3 125.4 -57.9 125.7 ;
        RECT  -64.5 123.3 -57.9 124.2 ;
        RECT  -64.5 123.0 -62.7 123.3 ;
        RECT  -60.3 123.0 -57.9 123.3 ;
        RECT  -61.5 121.2 -60.3 122.1 ;
        RECT  -64.5 120.3 -57.9 121.2 ;
        RECT  -64.5 120.0 -61.5 120.3 ;
        RECT  -59.1 120.0 -57.9 120.3 ;
        RECT  -66.9 117.6 -62.7 118.8 ;
        RECT  -66.9 113.1 -65.7 117.6 ;
        RECT  -61.8 116.7 -60.6 119.1 ;
        RECT  -56.4 118.8 -55.5 131.4 ;
        RECT  -59.1 117.6 -55.5 118.8 ;
        RECT  -64.5 115.5 -63.3 116.7 ;
        RECT  -64.5 114.6 -57.9 115.5 ;
        RECT  -64.5 114.3 -62.7 114.6 ;
        RECT  -59.1 114.3 -57.9 114.6 ;
        RECT  -56.4 113.1 -55.5 117.6 ;
        RECT  -66.9 111.9 -62.7 113.1 ;
        RECT  -66.9 108.3 -65.7 111.9 ;
        RECT  -61.2 111.0 -60.0 112.2 ;
        RECT  -59.1 111.9 -55.5 113.1 ;
        RECT  -64.5 110.7 -59.1 111.0 ;
        RECT  -64.5 110.1 -57.9 110.7 ;
        RECT  -64.5 109.5 -62.7 110.1 ;
        RECT  -60.3 109.8 -57.9 110.1 ;
        RECT  -59.1 109.5 -57.9 109.8 ;
        RECT  -66.9 107.1 -62.7 108.3 ;
        RECT  -66.9 92.1 -65.7 107.1 ;
        RECT  -61.2 106.5 -60.0 108.9 ;
        RECT  -56.4 108.3 -55.5 111.9 ;
        RECT  -59.1 107.1 -55.5 108.3 ;
        RECT  -56.7 105.9 -55.5 107.1 ;
        RECT  -64.5 102.6 -63.3 103.8 ;
        RECT  -62.4 103.5 -60.0 104.7 ;
        RECT  -64.5 101.7 -57.9 102.6 ;
        RECT  -64.5 101.4 -62.7 101.7 ;
        RECT  -59.1 101.4 -57.9 101.7 ;
        RECT  -64.5 99.3 -57.9 100.2 ;
        RECT  -64.5 99.0 -62.7 99.3 ;
        RECT  -60.3 99.0 -57.9 99.3 ;
        RECT  -64.5 96.9 -57.9 97.8 ;
        RECT  -64.5 96.6 -62.7 96.9 ;
        RECT  -60.3 96.6 -57.9 96.9 ;
        RECT  -61.5 94.8 -60.3 95.7 ;
        RECT  -64.5 93.9 -57.9 94.8 ;
        RECT  -64.5 93.6 -61.5 93.9 ;
        RECT  -59.1 93.6 -57.9 93.9 ;
        RECT  -56.4 92.4 -55.5 105.9 ;
        RECT  -64.5 92.1 -62.7 92.4 ;
        RECT  -66.9 91.2 -62.7 92.1 ;
        RECT  -59.1 91.5 -55.5 92.4 ;
        RECT  -59.1 91.2 -57.9 91.5 ;
        RECT  -63.9 89.7 -62.7 91.2 ;
        RECT  -61.8 88.8 -60.6 89.7 ;
        RECT  -66.9 87.9 -55.5 88.8 ;
        RECT  -56.7 141.9 -45.3 142.8 ;
        RECT  -46.5 138.6 -45.3 141.9 ;
        RECT  -54.3 140.1 -47.7 141.0 ;
        RECT  -50.7 139.8 -47.7 140.1 ;
        RECT  -54.3 139.8 -53.1 140.1 ;
        RECT  -49.5 137.4 -45.3 138.6 ;
        RECT  -56.7 137.4 -53.1 138.6 ;
        RECT  -46.5 133.8 -45.3 137.4 ;
        RECT  -51.9 136.5 -50.7 137.4 ;
        RECT  -53.1 136.2 -50.7 136.5 ;
        RECT  -54.3 135.3 -47.7 136.2 ;
        RECT  -49.5 135.0 -47.7 135.3 ;
        RECT  -54.3 135.0 -53.1 135.3 ;
        RECT  -49.5 132.6 -45.3 133.8 ;
        RECT  -46.5 118.8 -45.3 132.6 ;
        RECT  -52.2 132.0 -51.0 134.4 ;
        RECT  -56.7 133.8 -55.8 137.4 ;
        RECT  -56.7 132.6 -53.1 133.8 ;
        RECT  -56.7 131.4 -55.5 132.6 ;
        RECT  -48.9 129.0 -47.7 130.2 ;
        RECT  -52.2 129.9 -49.8 131.1 ;
        RECT  -54.3 128.1 -47.7 129.0 ;
        RECT  -49.5 127.8 -47.7 128.1 ;
        RECT  -54.3 127.8 -53.1 128.1 ;
        RECT  -54.3 125.7 -47.7 126.6 ;
        RECT  -49.5 125.4 -47.7 125.7 ;
        RECT  -54.3 125.4 -51.9 125.7 ;
        RECT  -54.3 123.3 -47.7 124.2 ;
        RECT  -49.5 123.0 -47.7 123.3 ;
        RECT  -54.3 123.0 -51.9 123.3 ;
        RECT  -51.9 121.2 -50.7 122.1 ;
        RECT  -54.3 120.3 -47.7 121.2 ;
        RECT  -50.7 120.0 -47.7 120.3 ;
        RECT  -54.3 120.0 -53.1 120.3 ;
        RECT  -49.5 117.6 -45.3 118.8 ;
        RECT  -46.5 113.1 -45.3 117.6 ;
        RECT  -51.6 116.7 -50.4 119.1 ;
        RECT  -56.7 118.8 -55.8 131.4 ;
        RECT  -56.7 117.6 -53.1 118.8 ;
        RECT  -48.9 115.5 -47.7 116.7 ;
        RECT  -54.3 114.6 -47.7 115.5 ;
        RECT  -49.5 114.3 -47.7 114.6 ;
        RECT  -54.3 114.3 -53.1 114.6 ;
        RECT  -56.7 113.1 -55.8 117.6 ;
        RECT  -49.5 111.9 -45.3 113.1 ;
        RECT  -46.5 108.3 -45.3 111.9 ;
        RECT  -52.2 111.0 -51.0 112.2 ;
        RECT  -56.7 111.9 -53.1 113.1 ;
        RECT  -53.1 110.7 -47.7 111.0 ;
        RECT  -54.3 110.1 -47.7 110.7 ;
        RECT  -49.5 109.5 -47.7 110.1 ;
        RECT  -54.3 109.8 -51.9 110.1 ;
        RECT  -54.3 109.5 -53.1 109.8 ;
        RECT  -49.5 107.1 -45.3 108.3 ;
        RECT  -46.5 92.1 -45.3 107.1 ;
        RECT  -52.2 106.5 -51.0 108.9 ;
        RECT  -56.7 108.3 -55.8 111.9 ;
        RECT  -56.7 107.1 -53.1 108.3 ;
        RECT  -56.7 105.9 -55.5 107.1 ;
        RECT  -48.9 102.6 -47.7 103.8 ;
        RECT  -52.2 103.5 -49.8 104.7 ;
        RECT  -54.3 101.7 -47.7 102.6 ;
        RECT  -49.5 101.4 -47.7 101.7 ;
        RECT  -54.3 101.4 -53.1 101.7 ;
        RECT  -54.3 99.3 -47.7 100.2 ;
        RECT  -49.5 99.0 -47.7 99.3 ;
        RECT  -54.3 99.0 -51.9 99.3 ;
        RECT  -54.3 96.9 -47.7 97.8 ;
        RECT  -49.5 96.6 -47.7 96.9 ;
        RECT  -54.3 96.6 -51.9 96.9 ;
        RECT  -51.9 94.8 -50.7 95.7 ;
        RECT  -54.3 93.9 -47.7 94.8 ;
        RECT  -50.7 93.6 -47.7 93.9 ;
        RECT  -54.3 93.6 -53.1 93.9 ;
        RECT  -56.7 92.4 -55.8 105.9 ;
        RECT  -49.5 92.1 -47.7 92.4 ;
        RECT  -49.5 91.2 -45.3 92.1 ;
        RECT  -56.7 91.5 -53.1 92.4 ;
        RECT  -54.3 91.2 -53.1 91.5 ;
        RECT  -49.5 89.7 -48.3 91.2 ;
        RECT  -51.6 88.8 -50.4 89.7 ;
        RECT  -56.7 87.9 -45.3 88.8 ;
        RECT  -46.5 141.9 -35.1 142.8 ;
        RECT  -46.5 138.6 -45.3 141.9 ;
        RECT  -44.1 140.1 -37.5 141.0 ;
        RECT  -44.1 139.8 -41.1 140.1 ;
        RECT  -38.7 139.8 -37.5 140.1 ;
        RECT  -46.5 137.4 -42.3 138.6 ;
        RECT  -38.7 137.4 -35.1 138.6 ;
        RECT  -46.5 133.8 -45.3 137.4 ;
        RECT  -41.1 136.5 -39.9 137.4 ;
        RECT  -41.1 136.2 -38.7 136.5 ;
        RECT  -44.1 135.3 -37.5 136.2 ;
        RECT  -44.1 135.0 -42.3 135.3 ;
        RECT  -38.7 135.0 -37.5 135.3 ;
        RECT  -46.5 132.6 -42.3 133.8 ;
        RECT  -46.5 118.8 -45.3 132.6 ;
        RECT  -40.8 132.0 -39.6 134.4 ;
        RECT  -36.0 133.8 -35.1 137.4 ;
        RECT  -38.7 132.6 -35.1 133.8 ;
        RECT  -36.3 131.4 -35.1 132.6 ;
        RECT  -44.1 129.0 -42.9 130.2 ;
        RECT  -42.0 129.9 -39.6 131.1 ;
        RECT  -44.1 128.1 -37.5 129.0 ;
        RECT  -44.1 127.8 -42.3 128.1 ;
        RECT  -38.7 127.8 -37.5 128.1 ;
        RECT  -44.1 125.7 -37.5 126.6 ;
        RECT  -44.1 125.4 -42.3 125.7 ;
        RECT  -39.9 125.4 -37.5 125.7 ;
        RECT  -44.1 123.3 -37.5 124.2 ;
        RECT  -44.1 123.0 -42.3 123.3 ;
        RECT  -39.9 123.0 -37.5 123.3 ;
        RECT  -41.1 121.2 -39.9 122.1 ;
        RECT  -44.1 120.3 -37.5 121.2 ;
        RECT  -44.1 120.0 -41.1 120.3 ;
        RECT  -38.7 120.0 -37.5 120.3 ;
        RECT  -46.5 117.6 -42.3 118.8 ;
        RECT  -46.5 113.1 -45.3 117.6 ;
        RECT  -41.4 116.7 -40.2 119.1 ;
        RECT  -36.0 118.8 -35.1 131.4 ;
        RECT  -38.7 117.6 -35.1 118.8 ;
        RECT  -44.1 115.5 -42.9 116.7 ;
        RECT  -44.1 114.6 -37.5 115.5 ;
        RECT  -44.1 114.3 -42.3 114.6 ;
        RECT  -38.7 114.3 -37.5 114.6 ;
        RECT  -36.0 113.1 -35.1 117.6 ;
        RECT  -46.5 111.9 -42.3 113.1 ;
        RECT  -46.5 108.3 -45.3 111.9 ;
        RECT  -40.8 111.0 -39.6 112.2 ;
        RECT  -38.7 111.9 -35.1 113.1 ;
        RECT  -44.1 110.7 -38.7 111.0 ;
        RECT  -44.1 110.1 -37.5 110.7 ;
        RECT  -44.1 109.5 -42.3 110.1 ;
        RECT  -39.9 109.8 -37.5 110.1 ;
        RECT  -38.7 109.5 -37.5 109.8 ;
        RECT  -46.5 107.1 -42.3 108.3 ;
        RECT  -46.5 92.1 -45.3 107.1 ;
        RECT  -40.8 106.5 -39.6 108.9 ;
        RECT  -36.0 108.3 -35.1 111.9 ;
        RECT  -38.7 107.1 -35.1 108.3 ;
        RECT  -36.3 105.9 -35.1 107.1 ;
        RECT  -44.1 102.6 -42.9 103.8 ;
        RECT  -42.0 103.5 -39.6 104.7 ;
        RECT  -44.1 101.7 -37.5 102.6 ;
        RECT  -44.1 101.4 -42.3 101.7 ;
        RECT  -38.7 101.4 -37.5 101.7 ;
        RECT  -44.1 99.3 -37.5 100.2 ;
        RECT  -44.1 99.0 -42.3 99.3 ;
        RECT  -39.9 99.0 -37.5 99.3 ;
        RECT  -44.1 96.9 -37.5 97.8 ;
        RECT  -44.1 96.6 -42.3 96.9 ;
        RECT  -39.9 96.6 -37.5 96.9 ;
        RECT  -41.1 94.8 -39.9 95.7 ;
        RECT  -44.1 93.9 -37.5 94.8 ;
        RECT  -44.1 93.6 -41.1 93.9 ;
        RECT  -38.7 93.6 -37.5 93.9 ;
        RECT  -36.0 92.4 -35.1 105.9 ;
        RECT  -44.1 92.1 -42.3 92.4 ;
        RECT  -46.5 91.2 -42.3 92.1 ;
        RECT  -38.7 91.5 -35.1 92.4 ;
        RECT  -38.7 91.2 -37.5 91.5 ;
        RECT  -43.5 89.7 -42.3 91.2 ;
        RECT  -41.4 88.8 -40.2 89.7 ;
        RECT  -46.5 87.9 -35.1 88.8 ;
        RECT  -7.95 128.7 -7.05 145.5 ;
        RECT  -22.65 128.7 -21.75 145.5 ;
        RECT  -21.75 142.5 -19.35 143.7 ;
        RECT  -9.75 142.5 -7.95 143.7 ;
        RECT  -19.5 132.9 -10.05 134.1 ;
        RECT  -19.5 137.7 -10.05 138.9 ;
        RECT  -14.7 128.7 -13.8 130.8 ;
        RECT  -14.7 138.9 -13.8 145.5 ;
        RECT  -7.95 130.5 -7.05 131.4 ;
        RECT  -7.95 135.3 -7.05 136.2 ;
        RECT  -7.95 135.3 -7.05 136.2 ;
        RECT  -7.95 140.1 -7.05 141.0 ;
        RECT  -10.05 130.5 -7.95 131.4 ;
        RECT  -7.95 130.5 -7.5 131.4 ;
        RECT  -7.95 130.95 -7.05 135.75 ;
        RECT  -10.05 135.3 -7.5 136.2 ;
        RECT  -10.05 135.3 -7.95 136.2 ;
        RECT  -7.95 135.3 -7.5 136.2 ;
        RECT  -7.95 135.75 -7.05 140.55 ;
        RECT  -10.05 140.1 -7.5 141.0 ;
        RECT  -11.85 132.9 -10.95 133.8 ;
        RECT  -11.85 137.7 -10.95 138.6 ;
        RECT  -10.95 132.9 -10.05 133.8 ;
        RECT  -11.4 132.9 -10.95 133.8 ;
        RECT  -11.85 133.35 -10.95 138.15 ;
        RECT  -11.4 137.7 -10.05 138.6 ;
        RECT  -11.25 130.5 -10.05 131.7 ;
        RECT  -11.25 132.9 -10.05 134.1 ;
        RECT  -11.25 135.3 -10.05 136.5 ;
        RECT  -11.25 137.7 -10.05 138.9 ;
        RECT  -11.25 140.1 -10.05 141.3 ;
        RECT  -22.35 130.5 -21.45 131.4 ;
        RECT  -22.35 135.3 -21.45 136.2 ;
        RECT  -22.35 135.3 -21.45 136.2 ;
        RECT  -22.35 140.1 -21.45 141.0 ;
        RECT  -21.45 130.5 -19.35 131.4 ;
        RECT  -21.9 130.5 -21.45 131.4 ;
        RECT  -22.35 130.95 -21.45 135.75 ;
        RECT  -21.9 135.3 -19.35 136.2 ;
        RECT  -21.45 135.3 -19.35 136.2 ;
        RECT  -21.9 135.3 -21.45 136.2 ;
        RECT  -22.35 135.75 -21.45 140.55 ;
        RECT  -21.9 140.1 -19.35 141.0 ;
        RECT  -18.45 132.9 -17.55 133.8 ;
        RECT  -18.45 137.7 -17.55 138.6 ;
        RECT  -19.35 132.9 -18.45 133.8 ;
        RECT  -18.45 132.9 -18.0 133.8 ;
        RECT  -18.45 133.35 -17.55 138.15 ;
        RECT  -19.35 137.7 -18.0 138.6 ;
        RECT  -20.55 130.5 -19.35 131.7 ;
        RECT  -20.55 132.9 -19.35 134.1 ;
        RECT  -20.55 135.3 -19.35 136.5 ;
        RECT  -20.55 137.7 -19.35 138.9 ;
        RECT  -20.55 140.1 -19.35 141.3 ;
        RECT  -20.55 142.5 -19.35 143.7 ;
        RECT  -10.05 142.5 -8.85 143.7 ;
        RECT  -14.85 130.8 -13.65 132.0 ;
        RECT  -7.95 88.5 -7.05 119.7 ;
        RECT  -22.65 88.5 -21.75 119.7 ;
        RECT  -14.1 116.4 -13.2 119.7 ;
        RECT  -16.05 102.0 -15.15 119.7 ;
        RECT  -14.1 114.45 -13.2 115.35 ;
        RECT  -14.1 88.5 -13.2 114.9 ;
        RECT  -13.65 114.45 -8.85 115.35 ;
        RECT  -14.1 88.5 -13.2 100.5 ;
        RECT  -14.1 88.5 -13.2 95.7 ;
        RECT  -22.2 90.6 -19.65 91.5 ;
        RECT  -8.85 109.8 -7.5 110.7 ;
        RECT  -21.75 117.0 -19.65 117.9 ;
        RECT  -18.0 114.45 -17.1 115.35 ;
        RECT  -19.65 114.45 -17.55 115.35 ;
        RECT  -18.0 105.3 -17.1 114.9 ;
        RECT  -21.75 112.2 -19.65 113.1 ;
        RECT  -18.0 109.65 -17.1 110.55 ;
        RECT  -19.65 109.65 -17.55 110.55 ;
        RECT  -18.0 105.3 -17.1 110.1 ;
        RECT  -21.75 107.4 -19.65 108.3 ;
        RECT  -18.0 102.45 -17.1 103.35 ;
        RECT  -19.65 102.45 -17.55 103.35 ;
        RECT  -18.0 102.9 -17.1 105.3 ;
        RECT  -18.0 97.65 -17.1 98.55 ;
        RECT  -19.65 97.65 -17.55 98.55 ;
        RECT  -18.0 98.1 -17.1 105.3 ;
        RECT  -18.0 92.85 -17.1 93.75 ;
        RECT  -19.65 92.85 -17.55 93.75 ;
        RECT  -18.0 93.3 -17.1 105.3 ;
        RECT  -8.85 117.0 -7.05 117.9 ;
        RECT  -8.85 112.2 -7.05 113.1 ;
        RECT  -13.65 116.7 -12.45 117.9 ;
        RECT  -13.65 114.3 -12.45 115.5 ;
        RECT  -13.65 114.3 -12.45 115.5 ;
        RECT  -13.65 111.9 -12.45 113.1 ;
        RECT  -16.05 116.7 -14.85 117.9 ;
        RECT  -16.05 114.3 -14.85 115.5 ;
        RECT  -16.05 111.9 -14.85 113.1 ;
        RECT  -16.05 109.5 -14.85 110.7 ;
        RECT  -16.05 107.1 -14.85 108.3 ;
        RECT  -16.05 102.3 -14.85 103.5 ;
        RECT  -16.05 99.9 -14.85 101.1 ;
        RECT  -16.05 97.5 -14.85 98.7 ;
        RECT  -16.05 95.1 -14.85 96.3 ;
        RECT  -16.05 92.7 -14.85 93.9 ;
        RECT  -19.65 90.3 -18.45 91.5 ;
        RECT  -8.85 109.5 -7.65 110.7 ;
        RECT  -13.05 116.4 -11.85 117.6 ;
        RECT  -15.0 102.0 -13.8 103.2 ;
        RECT  -19.65 99.9 -18.45 101.1 ;
        RECT  -13.05 99.9 -11.85 101.1 ;
        RECT  -19.65 95.1 -18.45 96.3 ;
        RECT  -13.05 95.1 -11.85 96.3 ;
        RECT  -7.95 164.4 -7.05 176.4 ;
        RECT  -22.65 164.4 -21.75 176.4 ;
        RECT  -22.2 173.4 -19.35 174.3 ;
        RECT  -9.9 173.4 -7.5 174.3 ;
        RECT  -22.2 166.35 -19.35 167.25 ;
        RECT  -22.2 171.15 -19.35 172.05 ;
        RECT  -10.35 166.35 -7.5 167.25 ;
        RECT  -17.1 171.6 -16.2 172.5 ;
        RECT  -17.1 168.6 -16.2 169.5 ;
        RECT  -16.65 171.6 -9.15 172.5 ;
        RECT  -17.1 169.05 -16.2 172.05 ;
        RECT  -19.35 168.6 -16.65 169.5 ;
        RECT  -17.1 164.4 -16.2 166.5 ;
        RECT  -13.8 164.4 -12.9 169.5 ;
        RECT  -14.7 172.05 -13.8 176.4 ;
        RECT  -11.55 166.2 -10.35 167.4 ;
        RECT  -11.55 168.6 -10.35 169.8 ;
        RECT  -11.55 168.6 -10.35 169.8 ;
        RECT  -11.55 171.0 -10.35 172.2 ;
        RECT  -20.55 166.2 -19.35 167.4 ;
        RECT  -20.55 168.6 -19.35 169.8 ;
        RECT  -20.55 168.6 -19.35 169.8 ;
        RECT  -20.55 171.0 -19.35 172.2 ;
        RECT  -20.55 173.4 -19.35 174.6 ;
        RECT  -10.35 173.4 -9.15 174.6 ;
        RECT  -17.1 166.5 -15.9 167.7 ;
        RECT  -13.8 169.5 -12.6 170.7 ;
        RECT  -43.05 236.7 -41.85 237.9 ;
        RECT  -14.55 265.35 -13.65 266.25 ;
        RECT  -14.1 265.35 -7.95 266.25 ;
        RECT  -14.55 265.8 -13.65 267.6 ;
        RECT  -32.7 235.05 -31.8 237.15 ;
        RECT  -45.0 235.05 -44.1 237.15 ;
        RECT  -45.0 236.7 -44.1 237.6 ;
        RECT  -55.35 236.7 -44.55 237.6 ;
        RECT  -31.65 261.75 -13.2 262.65 ;
        RECT  -51.75 251.55 -49.2 252.45 ;
        RECT  -16.35 245.25 -15.45 246.15 ;
        RECT  -16.35 243.15 -15.45 245.7 ;
        RECT  -32.25 245.25 -15.9 246.15 ;
        RECT  -45.45 245.25 -32.25 246.15 ;
        RECT  -16.35 236.7 -15.45 237.6 ;
        RECT  -16.35 237.15 -15.45 240.75 ;
        RECT  -32.25 236.7 -15.9 237.6 ;
        RECT  -61.95 293.25 -7.95 294.15 ;
        RECT  -23.1 265.35 -22.2 266.25 ;
        RECT  -23.1 265.8 -22.2 267.6 ;
        RECT  -45.45 265.35 -22.65 266.25 ;
        RECT  -45.45 265.35 -22.65 266.25 ;
        RECT  -32.25 230.55 -7.95 231.45 ;
        RECT  -37.35 288.15 -7.95 289.05 ;
        RECT  -8.4 269.4 -7.5 288.6 ;
        RECT  -37.8 269.4 -36.9 288.6 ;
        RECT  -42.75 267.6 -36.9 268.5 ;
        RECT  -51.75 256.95 -42.75 257.85 ;
        RECT  -51.75 268.35 -45.45 269.25 ;
        RECT  -42.75 267.6 -36.9 268.5 ;
        RECT  -51.75 280.95 -42.75 281.85 ;
        RECT  -56.85 240.15 -45.45 241.05 ;
        RECT  -61.95 230.55 -22.65 231.45 ;
        RECT  -51.75 230.55 -22.65 231.45 ;
        RECT  -41.85 230.55 -32.25 231.45 ;
        RECT  -41.85 215.85 -32.25 216.75 ;
        RECT  -40.05 216.75 -38.85 220.5 ;
        RECT  -40.05 228.75 -38.85 230.55 ;
        RECT  -35.25 229.65 -34.05 230.55 ;
        RECT  -35.25 216.75 -34.05 217.8 ;
        RECT  -37.65 220.35 -36.45 228.45 ;
        RECT  -34.35 224.4 -32.25 225.3 ;
        RECT  -41.85 224.4 -37.65 225.3 ;
        RECT  -35.25 227.25 -34.05 228.45 ;
        RECT  -37.65 227.25 -36.45 228.45 ;
        RECT  -35.25 217.8 -34.05 220.5 ;
        RECT  -37.65 217.8 -36.45 220.5 ;
        RECT  -40.05 217.8 -38.85 220.5 ;
        RECT  -40.05 228.45 -38.85 229.65 ;
        RECT  -35.55 224.25 -34.35 225.45 ;
        RECT  -16.35 235.35 -15.15 236.55 ;
        RECT  -16.35 232.95 -15.15 234.15 ;
        RECT  -14.85 266.4 -13.65 267.6 ;
        RECT  -8.4 258.0 -7.5 267.6 ;
        RECT  -23.1 258.0 -22.2 267.6 ;
        RECT  -22.2 259.8 -18.45 261.0 ;
        RECT  -10.2 259.8 -8.4 261.0 ;
        RECT  -9.3 264.6 -8.4 265.8 ;
        RECT  -22.2 264.6 -21.15 265.8 ;
        RECT  -18.6 262.2 -10.5 263.4 ;
        RECT  -14.55 265.5 -13.65 267.6 ;
        RECT  -14.1 264.6 -12.9 265.8 ;
        RECT  -14.1 262.2 -12.9 263.4 ;
        RECT  -13.95 264.6 -11.25 265.8 ;
        RECT  -13.95 262.2 -11.25 263.4 ;
        RECT  -18.45 259.8 -15.75 261.0 ;
        RECT  -9.3 259.8 -8.1 261.0 ;
        RECT  -13.5 264.3 -12.3 265.5 ;
        RECT  -14.85 256.8 -13.65 258.0 ;
        RECT  -8.4 248.4 -7.5 258.0 ;
        RECT  -23.1 248.4 -22.2 258.0 ;
        RECT  -22.2 250.2 -18.45 251.4 ;
        RECT  -10.2 250.2 -8.4 251.4 ;
        RECT  -9.3 255.0 -8.4 256.2 ;
        RECT  -22.2 255.0 -21.15 256.2 ;
        RECT  -18.6 252.6 -10.5 253.8 ;
        RECT  -14.55 255.9 -13.65 258.0 ;
        RECT  -14.1 255.0 -12.9 256.2 ;
        RECT  -14.1 252.6 -12.9 253.8 ;
        RECT  -13.95 255.0 -11.25 256.2 ;
        RECT  -13.95 252.6 -11.25 253.8 ;
        RECT  -18.45 250.2 -15.75 251.4 ;
        RECT  -9.3 250.2 -8.1 251.4 ;
        RECT  -13.5 254.7 -12.3 255.9 ;
        RECT  -31.65 248.4 -30.45 249.6 ;
        RECT  -37.8 248.4 -36.9 258.0 ;
        RECT  -23.1 248.4 -22.2 258.0 ;
        RECT  -26.85 255.0 -23.1 256.2 ;
        RECT  -36.9 255.0 -35.1 256.2 ;
        RECT  -36.9 250.2 -36.0 251.4 ;
        RECT  -24.15 250.2 -23.1 251.4 ;
        RECT  -34.8 252.6 -26.7 253.8 ;
        RECT  -31.65 248.4 -30.75 250.5 ;
        RECT  -32.4 250.2 -31.2 251.4 ;
        RECT  -32.4 252.6 -31.2 253.8 ;
        RECT  -34.05 250.2 -31.35 251.4 ;
        RECT  -34.05 252.6 -31.35 253.8 ;
        RECT  -29.55 255.0 -26.85 256.2 ;
        RECT  -37.2 255.0 -36.0 256.2 ;
        RECT  -33.0 250.5 -31.8 251.7 ;
        RECT  -31.65 258.0 -30.45 259.2 ;
        RECT  -37.8 258.0 -36.9 267.6 ;
        RECT  -23.1 258.0 -22.2 267.6 ;
        RECT  -26.85 264.6 -23.1 265.8 ;
        RECT  -36.9 264.6 -35.1 265.8 ;
        RECT  -36.9 259.8 -36.0 261.0 ;
        RECT  -24.15 259.8 -23.1 261.0 ;
        RECT  -34.8 262.2 -26.7 263.4 ;
        RECT  -31.65 258.0 -30.75 260.1 ;
        RECT  -32.4 259.8 -31.2 261.0 ;
        RECT  -32.4 262.2 -31.2 263.4 ;
        RECT  -34.05 259.8 -31.35 261.0 ;
        RECT  -34.05 262.2 -31.35 263.4 ;
        RECT  -29.55 264.6 -26.85 265.8 ;
        RECT  -37.2 264.6 -36.0 265.8 ;
        RECT  -33.0 260.1 -31.8 261.3 ;
        RECT  -14.85 261.0 -13.65 262.2 ;
        RECT  -14.85 251.4 -13.65 252.6 ;
        RECT  -31.65 253.8 -30.45 255.0 ;
        RECT  -62.55 268.2 -51.75 269.4 ;
        RECT  -53.55 266.1 -52.35 268.2 ;
        RECT  -56.55 266.1 -55.35 267.3 ;
        RECT  -59.55 266.1 -58.35 267.3 ;
        RECT  -62.55 266.1 -61.35 268.2 ;
        RECT  -56.25 265.2 -55.05 266.1 ;
        RECT  -57.45 264.0 -52.35 265.2 ;
        RECT  -53.55 258.9 -52.35 264.0 ;
        RECT  -56.25 260.7 -55.05 264.0 ;
        RECT  -59.85 262.5 -58.65 266.1 ;
        RECT  -59.85 261.3 -58.05 262.5 ;
        RECT  -59.85 260.7 -58.65 261.3 ;
        RECT  -55.95 259.5 -54.75 260.7 ;
        RECT  -60.15 259.5 -58.95 260.7 ;
        RECT  -62.55 259.5 -61.35 265.2 ;
        RECT  -58.05 258.0 -56.85 258.3 ;
        RECT  -62.55 256.8 -51.75 258.0 ;
        RECT  -55.95 254.7 -53.25 255.9 ;
        RECT  -60.15 254.7 -57.45 255.9 ;
        RECT  -62.55 240.0 -51.15 241.2 ;
        RECT  -53.55 241.2 -52.35 243.3 ;
        RECT  -56.55 242.1 -55.35 243.3 ;
        RECT  -59.55 242.1 -58.35 243.3 ;
        RECT  -62.55 241.2 -61.35 243.3 ;
        RECT  -56.25 243.3 -55.05 244.2 ;
        RECT  -53.55 244.2 -52.35 249.9 ;
        RECT  -57.45 244.2 -55.05 245.4 ;
        RECT  -56.25 245.4 -55.05 248.7 ;
        RECT  -59.85 243.3 -58.65 246.9 ;
        RECT  -59.85 246.9 -58.05 248.1 ;
        RECT  -59.85 248.1 -58.65 248.7 ;
        RECT  -55.95 248.7 -54.75 249.9 ;
        RECT  -60.15 248.7 -58.95 249.9 ;
        RECT  -62.55 244.2 -61.35 249.9 ;
        RECT  -58.05 251.1 -56.85 251.4 ;
        RECT  -62.55 251.4 -51.15 252.6 ;
        RECT  -55.95 253.5 -53.25 254.7 ;
        RECT  -60.15 253.5 -57.45 254.7 ;
        RECT  -62.55 238.8 -51.15 240.0 ;
        RECT  -53.55 236.7 -52.35 238.8 ;
        RECT  -56.55 236.7 -55.35 237.9 ;
        RECT  -59.55 236.7 -58.35 237.9 ;
        RECT  -62.55 236.7 -61.35 238.8 ;
        RECT  -56.25 235.8 -55.05 236.7 ;
        RECT  -53.55 230.1 -52.35 235.8 ;
        RECT  -57.45 234.6 -55.05 235.8 ;
        RECT  -56.25 231.3 -55.05 234.6 ;
        RECT  -59.85 233.1 -58.65 236.7 ;
        RECT  -59.85 231.9 -58.05 233.1 ;
        RECT  -59.85 231.3 -58.65 231.9 ;
        RECT  -55.95 230.1 -54.75 231.3 ;
        RECT  -60.15 230.1 -58.95 231.3 ;
        RECT  -62.55 230.1 -61.35 235.8 ;
        RECT  -58.05 228.6 -56.85 228.9 ;
        RECT  -62.55 227.4 -51.15 228.6 ;
        RECT  -55.95 225.3 -53.25 226.5 ;
        RECT  -60.15 225.3 -57.45 226.5 ;
        RECT  -43.05 235.95 -41.85 237.15 ;
        RECT  -32.85 233.25 -31.65 234.45 ;
        RECT  -45.15 233.25 -43.95 234.45 ;
        RECT  -55.95 235.35 -54.75 236.55 ;
        RECT  -13.95 240.15 -12.75 241.35 ;
        RECT  -13.8 260.4 -12.6 261.6 ;
        RECT  -32.25 260.4 -31.05 261.6 ;
        RECT  -32.85 271.8 -31.65 273.0 ;
        RECT  -13.8 240.15 -12.6 241.35 ;
        RECT  -50.25 250.2 -49.05 251.4 ;
        RECT  -46.05 243.9 -44.85 245.1 ;
        RECT  -46.05 264.0 -44.85 265.2 ;
        RECT  -8.55 229.2 -7.35 230.4 ;
        RECT  -8.55 286.8 -7.35 288.0 ;
        RECT  -37.95 286.8 -36.75 288.0 ;
        RECT  -46.65 293.25 -45.45 294.45 ;
        RECT  -43.35 266.25 -42.15 267.45 ;
        RECT  -43.35 255.6 -42.15 256.8 ;
        RECT  -46.05 267.0 -44.85 268.2 ;
        RECT  -43.35 266.25 -42.15 267.45 ;
        RECT  -43.35 279.6 -42.15 280.8 ;
        RECT  -46.05 238.8 -44.85 240.0 ;
        RECT  -62.55 229.2 -61.35 230.4 ;
        RECT  -52.35 229.2 -51.15 230.4 ;
        RECT  -7.95 180.0 -7.05 189.6 ;
        RECT  -22.65 180.0 -21.75 189.6 ;
        RECT  -21.75 181.8 -19.35 183.0 ;
        RECT  -9.75 181.8 -7.95 183.0 ;
        RECT  -8.85 186.6 -7.95 187.8 ;
        RECT  -21.75 186.6 -20.55 187.8 ;
        RECT  -19.5 184.2 -10.05 185.4 ;
        RECT  -14.7 187.5 -13.8 189.6 ;
        RECT  -14.7 180.0 -13.8 184.2 ;
        RECT  -13.65 186.6 -12.45 187.8 ;
        RECT  -13.65 184.2 -12.45 185.4 ;
        RECT  -14.55 186.6 -13.35 187.8 ;
        RECT  -14.55 184.2 -13.35 185.4 ;
        RECT  -19.35 181.8 -18.15 183.0 ;
        RECT  -8.85 181.8 -7.65 183.0 ;
        RECT  -13.65 186.3 -12.45 187.5 ;
        RECT  -7.95 189.6 -7.05 199.2 ;
        RECT  -22.65 189.6 -21.75 199.2 ;
        RECT  -21.75 191.4 -19.35 192.6 ;
        RECT  -9.75 191.4 -7.95 192.6 ;
        RECT  -8.85 196.2 -7.95 197.4 ;
        RECT  -21.75 196.2 -20.55 197.4 ;
        RECT  -19.5 193.8 -10.05 195.0 ;
        RECT  -14.7 197.1 -13.8 199.2 ;
        RECT  -14.7 189.6 -13.8 193.8 ;
        RECT  -13.65 196.2 -12.45 197.4 ;
        RECT  -13.65 193.8 -12.45 195.0 ;
        RECT  -14.55 196.2 -13.35 197.4 ;
        RECT  -14.55 193.8 -13.35 195.0 ;
        RECT  -19.35 191.4 -18.15 192.6 ;
        RECT  -8.85 191.4 -7.65 192.6 ;
        RECT  -13.65 195.9 -12.45 197.1 ;
        RECT  -37.35 164.4 -36.45 180.0 ;
        RECT  -22.65 164.4 -21.75 180.0 ;
        RECT  -35.1 175.2 -24.0 176.1 ;
        RECT  -25.05 177.0 -22.2 177.9 ;
        RECT  -36.9 177.0 -33.3 177.9 ;
        RECT  -25.05 167.55 -22.2 168.45 ;
        RECT  -25.05 172.35 -22.2 173.25 ;
        RECT  -36.9 167.55 -34.05 168.45 ;
        RECT  -27.15 164.4 -26.25 168.6 ;
        RECT  -32.7 164.4 -31.8 166.5 ;
        RECT  -34.5 164.4 -33.6 166.5 ;
        RECT  -29.85 175.2 -28.95 180.0 ;
        RECT  -30.9 167.4 -28.2 168.6 ;
        RECT  -30.9 169.8 -28.2 171.0 ;
        RECT  -30.9 169.8 -28.2 171.0 ;
        RECT  -30.9 172.2 -28.2 173.4 ;
        RECT  -30.9 172.2 -28.2 173.4 ;
        RECT  -30.9 174.6 -28.2 175.8 ;
        RECT  -31.05 167.4 -29.85 168.6 ;
        RECT  -31.05 169.8 -29.85 171.0 ;
        RECT  -31.05 169.8 -29.85 171.0 ;
        RECT  -31.05 172.2 -29.85 173.4 ;
        RECT  -31.05 172.2 -29.85 173.4 ;
        RECT  -31.05 174.6 -29.85 175.8 ;
        RECT  -26.25 177.0 -25.05 178.2 ;
        RECT  -38.1 177.0 -35.4 178.2 ;
        RECT  -26.25 169.8 -25.05 171.0 ;
        RECT  -26.25 174.6 -25.05 175.8 ;
        RECT  -28.65 167.4 -27.45 168.6 ;
        RECT  -33.0 170.7 -31.8 171.9 ;
        RECT  -33.0 170.7 -31.8 171.9 ;
        RECT  -33.9 165.3 -32.7 166.5 ;
        RECT  -33.0 173.1 -31.8 174.3 ;
        RECT  -33.0 173.1 -31.8 174.3 ;
        RECT  -36.0 165.3 -34.8 166.5 ;
        RECT  -37.35 164.4 -36.45 180.0 ;
        RECT  -52.05 164.4 -51.15 180.0 ;
        RECT  -49.8 175.2 -38.7 176.1 ;
        RECT  -51.6 177.0 -48.75 177.9 ;
        RECT  -40.5 177.0 -36.9 177.9 ;
        RECT  -51.6 167.55 -48.75 168.45 ;
        RECT  -51.6 172.35 -48.75 173.25 ;
        RECT  -39.75 167.55 -36.9 168.45 ;
        RECT  -47.55 164.4 -46.65 168.6 ;
        RECT  -42.0 164.4 -41.1 166.5 ;
        RECT  -40.2 164.4 -39.3 166.5 ;
        RECT  -44.85 175.2 -43.95 180.0 ;
        RECT  -43.8 167.4 -41.1 168.6 ;
        RECT  -43.8 169.8 -41.1 171.0 ;
        RECT  -43.8 169.8 -41.1 171.0 ;
        RECT  -43.8 172.2 -41.1 173.4 ;
        RECT  -43.8 172.2 -41.1 173.4 ;
        RECT  -43.8 174.6 -41.1 175.8 ;
        RECT  -49.95 167.4 -48.75 168.6 ;
        RECT  -49.95 169.8 -48.75 171.0 ;
        RECT  -49.95 169.8 -48.75 171.0 ;
        RECT  -49.95 172.2 -48.75 173.4 ;
        RECT  -49.95 172.2 -48.75 173.4 ;
        RECT  -49.95 174.6 -48.75 175.8 ;
        RECT  -49.95 177.0 -48.75 178.2 ;
        RECT  -41.1 177.0 -38.4 178.2 ;
        RECT  -49.95 169.8 -48.75 171.0 ;
        RECT  -49.95 174.6 -48.75 175.8 ;
        RECT  -47.55 167.4 -46.35 168.6 ;
        RECT  -43.2 170.7 -42.0 171.9 ;
        RECT  -43.2 170.7 -42.0 171.9 ;
        RECT  -42.3 165.3 -41.1 166.5 ;
        RECT  -43.2 173.1 -42.0 174.3 ;
        RECT  -43.2 173.1 -42.0 174.3 ;
        RECT  -40.2 165.3 -39.0 166.5 ;
        RECT  -37.35 180.0 -36.45 189.6 ;
        RECT  -22.65 180.0 -21.75 189.6 ;
        RECT  -25.05 186.6 -22.65 187.8 ;
        RECT  -36.45 186.6 -34.65 187.8 ;
        RECT  -36.45 181.8 -35.55 183.0 ;
        RECT  -23.85 181.8 -22.65 183.0 ;
        RECT  -34.35 184.2 -24.9 185.4 ;
        RECT  -30.6 180.0 -29.7 182.1 ;
        RECT  -30.6 185.4 -29.7 189.6 ;
        RECT  -31.95 181.8 -30.75 183.0 ;
        RECT  -31.95 184.2 -30.75 185.4 ;
        RECT  -31.05 181.8 -29.85 183.0 ;
        RECT  -31.05 184.2 -29.85 185.4 ;
        RECT  -26.25 186.6 -25.05 187.8 ;
        RECT  -36.75 186.6 -35.55 187.8 ;
        RECT  -31.95 182.1 -30.75 183.3 ;
        RECT  -37.35 180.0 -36.45 189.6 ;
        RECT  -52.05 180.0 -51.15 189.6 ;
        RECT  -51.15 186.6 -48.75 187.8 ;
        RECT  -39.15 186.6 -37.35 187.8 ;
        RECT  -38.25 181.8 -37.35 183.0 ;
        RECT  -51.15 181.8 -49.95 183.0 ;
        RECT  -48.9 184.2 -39.45 185.4 ;
        RECT  -44.1 180.0 -43.2 182.1 ;
        RECT  -44.1 185.4 -43.2 189.6 ;
        RECT  -40.65 181.8 -39.45 183.0 ;
        RECT  -40.65 184.2 -39.45 185.4 ;
        RECT  -49.95 181.8 -48.75 183.0 ;
        RECT  -49.95 184.2 -48.75 185.4 ;
        RECT  -49.95 186.6 -48.75 187.8 ;
        RECT  -39.45 186.6 -38.25 187.8 ;
        RECT  -44.25 182.1 -43.05 183.3 ;
        RECT  -37.35 189.6 -36.45 199.2 ;
        RECT  -52.05 189.6 -51.15 199.2 ;
        RECT  -51.15 196.2 -48.75 197.4 ;
        RECT  -39.15 196.2 -37.35 197.4 ;
        RECT  -38.25 191.4 -37.35 192.6 ;
        RECT  -51.15 191.4 -49.95 192.6 ;
        RECT  -48.9 193.8 -39.45 195.0 ;
        RECT  -44.1 189.6 -43.2 191.7 ;
        RECT  -44.1 195.0 -43.2 199.2 ;
        RECT  -40.65 191.4 -39.45 192.6 ;
        RECT  -40.65 193.8 -39.45 195.0 ;
        RECT  -49.95 191.4 -48.75 192.6 ;
        RECT  -49.95 193.8 -48.75 195.0 ;
        RECT  -49.95 196.2 -48.75 197.4 ;
        RECT  -39.45 196.2 -38.25 197.4 ;
        RECT  -44.25 191.7 -43.05 192.9 ;
        RECT  -37.35 199.2 -36.45 208.8 ;
        RECT  -52.05 199.2 -51.15 208.8 ;
        RECT  -51.15 205.8 -48.75 207.0 ;
        RECT  -39.15 205.8 -37.35 207.0 ;
        RECT  -38.25 201.0 -37.35 202.2 ;
        RECT  -51.15 201.0 -49.95 202.2 ;
        RECT  -48.9 203.4 -39.45 204.6 ;
        RECT  -44.1 199.2 -43.2 201.3 ;
        RECT  -44.1 204.6 -43.2 208.8 ;
        RECT  -40.65 201.0 -39.45 202.2 ;
        RECT  -40.65 203.4 -39.45 204.6 ;
        RECT  -49.95 201.0 -48.75 202.2 ;
        RECT  -49.95 203.4 -48.75 204.6 ;
        RECT  -49.95 205.8 -48.75 207.0 ;
        RECT  -39.45 205.8 -38.25 207.0 ;
        RECT  -44.25 201.3 -43.05 202.5 ;
        RECT  -40.8 144.3 -39.6 145.5 ;
        RECT  -40.8 150.9 -39.6 152.1 ;
        RECT  -44.25 144.3 -43.05 145.5 ;
        RECT  -44.25 153.6 -43.05 154.8 ;
        RECT  -64.65 144.3 -63.45 145.5 ;
        RECT  -64.65 156.3 -63.45 157.5 ;
        RECT  -49.05 144.3 -47.85 145.5 ;
        RECT  -49.05 159.0 -47.85 160.2 ;
        RECT  -17.4 153.6 -16.2 154.8 ;
        RECT  -14.1 161.7 -12.9 162.9 ;
        RECT  -27.45 161.7 -26.25 162.9 ;
        RECT  -33.0 153.6 -31.8 154.8 ;
        RECT  -34.8 156.3 -33.6 157.5 ;
        RECT  -47.85 161.7 -46.65 162.9 ;
        RECT  -42.3 159.0 -41.1 160.2 ;
        RECT  -40.5 156.3 -39.3 157.5 ;
        RECT  -16.2 120.9 -15.0 122.1 ;
        RECT  -5.85 120.9 -4.65 122.1 ;
        RECT  -5.85 150.75 -4.65 151.95 ;
        RECT  -30.9 214.2 -29.7 215.4 ;
        RECT  -44.4 211.5 -43.2 212.7 ;
        RECT  -15.0 216.9 -13.8 218.1 ;
        RECT  -4.05 214.05 -2.85 215.25 ;
        RECT  -22.95 219.6 -21.75 220.8 ;
        RECT  -52.35 219.6 -51.15 220.8 ;
        RECT  -8.25 148.2 -7.05 149.4 ;
        RECT  -14.85 126.3 -13.65 127.5 ;
        RECT  -27.75 126.3 -26.55 127.5 ;
        RECT  -27.6 85.5 -26.4 86.7 ;
        RECT  -14.1 88.5 -12.9 89.7 ;
        RECT  -15.0 175.5 -13.8 176.7 ;
        RECT  -15.0 180.0 -13.8 181.2 ;
        RECT  0.45 219.6 2.85 220.8 ;
        Layer  via1 ; 
        RECT  125.25 209.7 125.85 210.3 ;
        RECT  134.25 209.7 134.85 210.3 ;
        RECT  126.15 200.4 126.75 201.0 ;
        RECT  130.35 200.4 130.95 201.0 ;
        RECT  125.25 219.3 125.85 219.9 ;
        RECT  134.25 219.3 134.85 219.9 ;
        RECT  126.15 228.6 126.75 229.2 ;
        RECT  130.35 228.6 130.95 229.2 ;
        RECT  125.25 239.1 125.85 239.7 ;
        RECT  134.25 239.1 134.85 239.7 ;
        RECT  126.15 229.8 126.75 230.4 ;
        RECT  130.35 229.8 130.95 230.4 ;
        RECT  125.25 248.7 125.85 249.3 ;
        RECT  134.25 248.7 134.85 249.3 ;
        RECT  126.15 258.0 126.75 258.6 ;
        RECT  130.35 258.0 130.95 258.6 ;
        RECT  125.25 268.5 125.85 269.1 ;
        RECT  134.25 268.5 134.85 269.1 ;
        RECT  126.15 259.2 126.75 259.8 ;
        RECT  130.35 259.2 130.95 259.8 ;
        RECT  125.25 278.1 125.85 278.7 ;
        RECT  134.25 278.1 134.85 278.7 ;
        RECT  126.15 287.4 126.75 288.0 ;
        RECT  130.35 287.4 130.95 288.0 ;
        RECT  125.25 297.9 125.85 298.5 ;
        RECT  134.25 297.9 134.85 298.5 ;
        RECT  126.15 288.6 126.75 289.2 ;
        RECT  130.35 288.6 130.95 289.2 ;
        RECT  125.25 307.5 125.85 308.1 ;
        RECT  134.25 307.5 134.85 308.1 ;
        RECT  126.15 316.8 126.75 317.4 ;
        RECT  130.35 316.8 130.95 317.4 ;
        RECT  125.25 327.3 125.85 327.9 ;
        RECT  134.25 327.3 134.85 327.9 ;
        RECT  126.15 318.0 126.75 318.6 ;
        RECT  130.35 318.0 130.95 318.6 ;
        RECT  125.25 336.9 125.85 337.5 ;
        RECT  134.25 336.9 134.85 337.5 ;
        RECT  126.15 346.2 126.75 346.8 ;
        RECT  130.35 346.2 130.95 346.8 ;
        RECT  125.25 356.7 125.85 357.3 ;
        RECT  134.25 356.7 134.85 357.3 ;
        RECT  126.15 347.4 126.75 348.0 ;
        RECT  130.35 347.4 130.95 348.0 ;
        RECT  125.25 366.3 125.85 366.9 ;
        RECT  134.25 366.3 134.85 366.9 ;
        RECT  126.15 375.6 126.75 376.2 ;
        RECT  130.35 375.6 130.95 376.2 ;
        RECT  125.25 386.1 125.85 386.7 ;
        RECT  134.25 386.1 134.85 386.7 ;
        RECT  126.15 376.8 126.75 377.4 ;
        RECT  130.35 376.8 130.95 377.4 ;
        RECT  125.25 395.7 125.85 396.3 ;
        RECT  134.25 395.7 134.85 396.3 ;
        RECT  126.15 405.0 126.75 405.6 ;
        RECT  130.35 405.0 130.95 405.6 ;
        RECT  125.25 415.5 125.85 416.1 ;
        RECT  134.25 415.5 134.85 416.1 ;
        RECT  126.15 406.2 126.75 406.8 ;
        RECT  130.35 406.2 130.95 406.8 ;
        RECT  125.25 425.1 125.85 425.7 ;
        RECT  134.25 425.1 134.85 425.7 ;
        RECT  126.15 434.4 126.75 435.0 ;
        RECT  130.35 434.4 130.95 435.0 ;
        RECT  135.45 209.7 136.05 210.3 ;
        RECT  144.45 209.7 145.05 210.3 ;
        RECT  136.35 200.4 136.95 201.0 ;
        RECT  140.55 200.4 141.15 201.0 ;
        RECT  135.45 219.3 136.05 219.9 ;
        RECT  144.45 219.3 145.05 219.9 ;
        RECT  136.35 228.6 136.95 229.2 ;
        RECT  140.55 228.6 141.15 229.2 ;
        RECT  135.45 239.1 136.05 239.7 ;
        RECT  144.45 239.1 145.05 239.7 ;
        RECT  136.35 229.8 136.95 230.4 ;
        RECT  140.55 229.8 141.15 230.4 ;
        RECT  135.45 248.7 136.05 249.3 ;
        RECT  144.45 248.7 145.05 249.3 ;
        RECT  136.35 258.0 136.95 258.6 ;
        RECT  140.55 258.0 141.15 258.6 ;
        RECT  135.45 268.5 136.05 269.1 ;
        RECT  144.45 268.5 145.05 269.1 ;
        RECT  136.35 259.2 136.95 259.8 ;
        RECT  140.55 259.2 141.15 259.8 ;
        RECT  135.45 278.1 136.05 278.7 ;
        RECT  144.45 278.1 145.05 278.7 ;
        RECT  136.35 287.4 136.95 288.0 ;
        RECT  140.55 287.4 141.15 288.0 ;
        RECT  135.45 297.9 136.05 298.5 ;
        RECT  144.45 297.9 145.05 298.5 ;
        RECT  136.35 288.6 136.95 289.2 ;
        RECT  140.55 288.6 141.15 289.2 ;
        RECT  135.45 307.5 136.05 308.1 ;
        RECT  144.45 307.5 145.05 308.1 ;
        RECT  136.35 316.8 136.95 317.4 ;
        RECT  140.55 316.8 141.15 317.4 ;
        RECT  135.45 327.3 136.05 327.9 ;
        RECT  144.45 327.3 145.05 327.9 ;
        RECT  136.35 318.0 136.95 318.6 ;
        RECT  140.55 318.0 141.15 318.6 ;
        RECT  135.45 336.9 136.05 337.5 ;
        RECT  144.45 336.9 145.05 337.5 ;
        RECT  136.35 346.2 136.95 346.8 ;
        RECT  140.55 346.2 141.15 346.8 ;
        RECT  135.45 356.7 136.05 357.3 ;
        RECT  144.45 356.7 145.05 357.3 ;
        RECT  136.35 347.4 136.95 348.0 ;
        RECT  140.55 347.4 141.15 348.0 ;
        RECT  135.45 366.3 136.05 366.9 ;
        RECT  144.45 366.3 145.05 366.9 ;
        RECT  136.35 375.6 136.95 376.2 ;
        RECT  140.55 375.6 141.15 376.2 ;
        RECT  135.45 386.1 136.05 386.7 ;
        RECT  144.45 386.1 145.05 386.7 ;
        RECT  136.35 376.8 136.95 377.4 ;
        RECT  140.55 376.8 141.15 377.4 ;
        RECT  135.45 395.7 136.05 396.3 ;
        RECT  144.45 395.7 145.05 396.3 ;
        RECT  136.35 405.0 136.95 405.6 ;
        RECT  140.55 405.0 141.15 405.6 ;
        RECT  135.45 415.5 136.05 416.1 ;
        RECT  144.45 415.5 145.05 416.1 ;
        RECT  136.35 406.2 136.95 406.8 ;
        RECT  140.55 406.2 141.15 406.8 ;
        RECT  135.45 425.1 136.05 425.7 ;
        RECT  144.45 425.1 145.05 425.7 ;
        RECT  136.35 434.4 136.95 435.0 ;
        RECT  140.55 434.4 141.15 435.0 ;
        RECT  127.65 451.2 128.25 451.8 ;
        RECT  132.45 451.2 133.05 451.8 ;
        RECT  127.65 442.8 128.25 443.4 ;
        RECT  130.05 442.8 130.65 443.4 ;
        RECT  137.85 451.2 138.45 451.8 ;
        RECT  142.65 451.2 143.25 451.8 ;
        RECT  137.85 442.8 138.45 443.4 ;
        RECT  140.25 442.8 140.85 443.4 ;
        RECT  134.25 194.1 134.85 194.7 ;
        RECT  128.55 164.7 129.15 165.3 ;
        RECT  131.25 164.7 131.85 165.3 ;
        RECT  125.55 154.8 126.15 155.4 ;
        RECT  144.45 194.1 145.05 194.7 ;
        RECT  138.75 164.7 139.35 165.3 ;
        RECT  141.45 164.7 142.05 165.3 ;
        RECT  135.75 154.8 136.35 155.4 ;
        RECT  126.15 148.2 126.75 148.8 ;
        RECT  130.65 147.6 131.25 148.2 ;
        RECT  127.95 138.0 128.55 138.6 ;
        RECT  127.05 126.3 127.65 126.9 ;
        RECT  133.65 115.5 134.25 116.1 ;
        RECT  130.35 110.1 130.95 110.7 ;
        RECT  127.05 100.2 127.65 100.8 ;
        RECT  134.25 96.0 134.85 96.6 ;
        RECT  128.25 93.9 128.85 94.5 ;
        RECT  136.35 148.2 136.95 148.8 ;
        RECT  140.85 147.6 141.45 148.2 ;
        RECT  138.15 138.0 138.75 138.6 ;
        RECT  137.25 126.3 137.85 126.9 ;
        RECT  143.85 115.5 144.45 116.1 ;
        RECT  140.55 110.1 141.15 110.7 ;
        RECT  137.25 100.2 137.85 100.8 ;
        RECT  144.45 96.0 145.05 96.6 ;
        RECT  138.45 93.9 139.05 94.5 ;
        RECT  128.25 85.5 128.85 86.1 ;
        RECT  130.65 81.0 131.25 81.6 ;
        RECT  129.75 77.7 130.35 78.3 ;
        RECT  134.25 77.1 134.85 77.7 ;
        RECT  129.75 75.6 130.35 76.2 ;
        RECT  126.45 74.7 127.05 75.3 ;
        RECT  130.65 71.1 131.25 71.7 ;
        RECT  130.65 68.7 131.25 69.3 ;
        RECT  128.25 65.7 128.85 66.3 ;
        RECT  129.15 62.4 129.75 63.0 ;
        RECT  126.45 61.2 127.05 61.8 ;
        RECT  130.65 55.5 131.25 56.1 ;
        RECT  129.75 52.2 130.35 52.8 ;
        RECT  134.25 51.6 134.85 52.2 ;
        RECT  129.75 49.2 130.35 49.8 ;
        RECT  126.45 48.3 127.05 48.9 ;
        RECT  130.65 44.7 131.25 45.3 ;
        RECT  130.65 42.3 131.25 42.9 ;
        RECT  128.25 39.3 128.85 39.9 ;
        RECT  140.25 85.5 140.85 86.1 ;
        RECT  137.85 81.0 138.45 81.6 ;
        RECT  138.75 77.7 139.35 78.3 ;
        RECT  134.25 77.1 134.85 77.7 ;
        RECT  138.75 75.6 139.35 76.2 ;
        RECT  142.05 74.7 142.65 75.3 ;
        RECT  137.85 71.1 138.45 71.7 ;
        RECT  137.85 68.7 138.45 69.3 ;
        RECT  140.25 65.7 140.85 66.3 ;
        RECT  139.35 62.4 139.95 63.0 ;
        RECT  142.05 61.2 142.65 61.8 ;
        RECT  137.85 55.5 138.45 56.1 ;
        RECT  138.75 52.2 139.35 52.8 ;
        RECT  134.25 51.6 134.85 52.2 ;
        RECT  138.75 49.2 139.35 49.8 ;
        RECT  142.05 48.3 142.65 48.9 ;
        RECT  137.85 44.7 138.45 45.3 ;
        RECT  137.85 42.3 138.45 42.9 ;
        RECT  140.25 39.3 140.85 39.9 ;
        RECT  127.35 45.0 127.95 45.6 ;
        RECT  132.15 41.4 132.75 42.0 ;
        RECT  134.25 36.9 134.85 37.5 ;
        RECT  141.15 45.0 141.75 45.6 ;
        RECT  136.35 41.4 136.95 42.0 ;
        RECT  134.25 36.9 134.85 37.5 ;
        RECT  58.95 93.15 59.55 93.75 ;
        RECT  78.15 87.9 78.75 88.5 ;
        RECT  56.85 98.55 57.45 99.15 ;
        RECT  76.05 103.8 76.65 104.4 ;
        RECT  58.95 90.3 59.55 90.9 ;
        RECT  56.85 87.0 57.45 87.6 ;
        RECT  54.75 101.4 55.35 102.0 ;
        RECT  56.85 104.7 57.45 105.3 ;
        RECT  58.95 119.7 59.55 120.3 ;
        RECT  52.65 116.4 53.25 117.0 ;
        RECT  54.75 130.8 55.35 131.4 ;
        RECT  78.15 130.8 78.75 131.4 ;
        RECT  52.65 134.1 53.25 134.7 ;
        RECT  76.05 134.1 76.65 134.7 ;
        RECT  61.05 81.15 61.65 81.75 ;
        RECT  63.15 95.85 63.75 96.45 ;
        RECT  61.05 110.55 61.65 111.15 ;
        RECT  63.15 125.25 63.75 125.85 ;
        RECT  61.05 137.7 61.65 138.3 ;
        RECT  58.95 151.95 59.55 152.55 ;
        RECT  78.15 146.7 78.75 147.3 ;
        RECT  56.85 157.35 57.45 157.95 ;
        RECT  76.05 162.6 76.65 163.2 ;
        RECT  58.95 149.1 59.55 149.7 ;
        RECT  56.85 145.8 57.45 146.4 ;
        RECT  54.75 160.2 55.35 160.8 ;
        RECT  56.85 163.5 57.45 164.1 ;
        RECT  58.95 178.5 59.55 179.1 ;
        RECT  52.65 175.2 53.25 175.8 ;
        RECT  54.75 189.6 55.35 190.2 ;
        RECT  78.15 189.6 78.75 190.2 ;
        RECT  52.65 192.9 53.25 193.5 ;
        RECT  76.05 192.9 76.65 193.5 ;
        RECT  61.05 139.95 61.65 140.55 ;
        RECT  63.15 154.65 63.75 155.25 ;
        RECT  61.05 169.35 61.65 169.95 ;
        RECT  63.15 184.05 63.75 184.65 ;
        RECT  61.05 196.5 61.65 197.1 ;
        RECT  13.35 89.1 13.95 89.7 ;
        RECT  15.45 105.0 16.05 105.6 ;
        RECT  17.55 118.5 18.15 119.1 ;
        RECT  19.65 134.4 20.25 135.0 ;
        RECT  21.75 147.9 22.35 148.5 ;
        RECT  23.85 163.8 24.45 164.4 ;
        RECT  25.95 177.3 26.55 177.9 ;
        RECT  28.05 193.2 28.65 193.8 ;
        RECT  13.35 209.1 13.95 209.7 ;
        RECT  21.75 205.8 22.35 206.4 ;
        RECT  13.35 220.2 13.95 220.8 ;
        RECT  23.85 223.5 24.45 224.1 ;
        RECT  13.35 238.5 13.95 239.1 ;
        RECT  25.95 235.2 26.55 235.8 ;
        RECT  13.35 249.6 13.95 250.2 ;
        RECT  28.05 252.9 28.65 253.5 ;
        RECT  15.45 267.9 16.05 268.5 ;
        RECT  21.75 264.6 22.35 265.2 ;
        RECT  15.45 279.0 16.05 279.6 ;
        RECT  23.85 282.3 24.45 282.9 ;
        RECT  15.45 297.3 16.05 297.9 ;
        RECT  25.95 294.0 26.55 294.6 ;
        RECT  15.45 308.4 16.05 309.0 ;
        RECT  28.05 311.7 28.65 312.3 ;
        RECT  17.55 326.7 18.15 327.3 ;
        RECT  21.75 323.4 22.35 324.0 ;
        RECT  17.55 337.8 18.15 338.4 ;
        RECT  23.85 341.1 24.45 341.7 ;
        RECT  17.55 356.1 18.15 356.7 ;
        RECT  25.95 352.8 26.55 353.4 ;
        RECT  17.55 367.2 18.15 367.8 ;
        RECT  28.05 370.5 28.65 371.1 ;
        RECT  19.65 385.5 20.25 386.1 ;
        RECT  21.75 382.2 22.35 382.8 ;
        RECT  19.65 396.6 20.25 397.2 ;
        RECT  23.85 399.9 24.45 400.5 ;
        RECT  19.65 414.9 20.25 415.5 ;
        RECT  25.95 411.6 26.55 412.2 ;
        RECT  19.65 426.0 20.25 426.6 ;
        RECT  28.05 429.3 28.65 429.9 ;
        RECT  51.45 214.65 52.05 215.25 ;
        RECT  57.75 214.65 58.35 215.25 ;
        RECT  67.65 209.1 68.25 209.7 ;
        RECT  51.75 209.1 52.35 209.7 ;
        RECT  51.45 229.35 52.05 229.95 ;
        RECT  57.75 229.35 58.35 229.95 ;
        RECT  67.65 219.9 68.25 220.5 ;
        RECT  51.75 219.9 52.35 220.5 ;
        RECT  51.45 244.05 52.05 244.65 ;
        RECT  57.75 244.05 58.35 244.65 ;
        RECT  67.65 238.5 68.25 239.1 ;
        RECT  51.75 238.5 52.35 239.1 ;
        RECT  51.45 258.75 52.05 259.35 ;
        RECT  57.75 258.75 58.35 259.35 ;
        RECT  67.65 249.3 68.25 249.9 ;
        RECT  51.75 249.3 52.35 249.9 ;
        RECT  51.45 273.45 52.05 274.05 ;
        RECT  57.75 273.45 58.35 274.05 ;
        RECT  67.65 267.9 68.25 268.5 ;
        RECT  51.75 267.9 52.35 268.5 ;
        RECT  51.45 288.15 52.05 288.75 ;
        RECT  57.75 288.15 58.35 288.75 ;
        RECT  67.65 278.7 68.25 279.3 ;
        RECT  51.75 278.7 52.35 279.3 ;
        RECT  51.45 302.85 52.05 303.45 ;
        RECT  57.75 302.85 58.35 303.45 ;
        RECT  67.65 297.3 68.25 297.9 ;
        RECT  51.75 297.3 52.35 297.9 ;
        RECT  51.45 317.55 52.05 318.15 ;
        RECT  57.75 317.55 58.35 318.15 ;
        RECT  67.65 308.1 68.25 308.7 ;
        RECT  51.75 308.1 52.35 308.7 ;
        RECT  51.45 332.25 52.05 332.85 ;
        RECT  57.75 332.25 58.35 332.85 ;
        RECT  67.65 326.7 68.25 327.3 ;
        RECT  51.75 326.7 52.35 327.3 ;
        RECT  51.45 346.95 52.05 347.55 ;
        RECT  57.75 346.95 58.35 347.55 ;
        RECT  67.65 337.5 68.25 338.1 ;
        RECT  51.75 337.5 52.35 338.1 ;
        RECT  51.45 361.65 52.05 362.25 ;
        RECT  57.75 361.65 58.35 362.25 ;
        RECT  67.65 356.1 68.25 356.7 ;
        RECT  51.75 356.1 52.35 356.7 ;
        RECT  51.45 376.35 52.05 376.95 ;
        RECT  57.75 376.35 58.35 376.95 ;
        RECT  67.65 366.9 68.25 367.5 ;
        RECT  51.75 366.9 52.35 367.5 ;
        RECT  51.45 391.05 52.05 391.65 ;
        RECT  57.75 391.05 58.35 391.65 ;
        RECT  67.65 385.5 68.25 386.1 ;
        RECT  51.75 385.5 52.35 386.1 ;
        RECT  51.45 405.75 52.05 406.35 ;
        RECT  57.75 405.75 58.35 406.35 ;
        RECT  67.65 396.3 68.25 396.9 ;
        RECT  51.75 396.3 52.35 396.9 ;
        RECT  51.45 420.45 52.05 421.05 ;
        RECT  57.75 420.45 58.35 421.05 ;
        RECT  67.65 414.9 68.25 415.5 ;
        RECT  51.75 414.9 52.35 415.5 ;
        RECT  51.45 435.15 52.05 435.75 ;
        RECT  57.75 435.15 58.35 435.75 ;
        RECT  67.65 425.7 68.25 426.3 ;
        RECT  51.75 425.7 52.35 426.3 ;
        RECT  70.35 75.3 70.95 75.9 ;
        RECT  65.85 72.9 66.45 73.5 ;
        RECT  62.55 73.8 63.15 74.4 ;
        RECT  61.95 69.3 62.55 69.9 ;
        RECT  60.45 73.8 61.05 74.4 ;
        RECT  59.55 77.1 60.15 77.7 ;
        RECT  55.95 72.9 56.55 73.5 ;
        RECT  53.55 72.9 54.15 73.5 ;
        RECT  50.55 75.3 51.15 75.9 ;
        RECT  47.25 74.4 47.85 75.0 ;
        RECT  46.05 77.1 46.65 77.7 ;
        RECT  40.35 72.9 40.95 73.5 ;
        RECT  37.05 73.8 37.65 74.4 ;
        RECT  36.45 69.3 37.05 69.9 ;
        RECT  34.05 73.8 34.65 74.4 ;
        RECT  33.15 77.1 33.75 77.7 ;
        RECT  29.55 72.9 30.15 73.5 ;
        RECT  27.15 72.9 27.75 73.5 ;
        RECT  24.15 75.3 24.75 75.9 ;
        RECT  70.35 63.3 70.95 63.9 ;
        RECT  65.85 65.7 66.45 66.3 ;
        RECT  62.55 64.8 63.15 65.4 ;
        RECT  61.95 69.3 62.55 69.9 ;
        RECT  60.45 64.8 61.05 65.4 ;
        RECT  59.55 61.5 60.15 62.1 ;
        RECT  55.95 65.7 56.55 66.3 ;
        RECT  53.55 65.7 54.15 66.3 ;
        RECT  50.55 63.3 51.15 63.9 ;
        RECT  47.25 64.2 47.85 64.8 ;
        RECT  46.05 61.5 46.65 62.1 ;
        RECT  40.35 65.7 40.95 66.3 ;
        RECT  37.05 64.8 37.65 65.4 ;
        RECT  36.45 69.3 37.05 69.9 ;
        RECT  34.05 64.8 34.65 65.4 ;
        RECT  33.15 61.5 33.75 62.1 ;
        RECT  29.55 65.7 30.15 66.3 ;
        RECT  27.15 65.7 27.75 66.3 ;
        RECT  24.15 63.3 24.75 63.9 ;
        RECT  70.35 54.9 70.95 55.5 ;
        RECT  65.85 52.5 66.45 53.1 ;
        RECT  62.55 53.4 63.15 54.0 ;
        RECT  61.95 48.9 62.55 49.5 ;
        RECT  60.45 53.4 61.05 54.0 ;
        RECT  59.55 56.7 60.15 57.3 ;
        RECT  55.95 52.5 56.55 53.1 ;
        RECT  53.55 52.5 54.15 53.1 ;
        RECT  50.55 54.9 51.15 55.5 ;
        RECT  47.25 54.0 47.85 54.6 ;
        RECT  46.05 56.7 46.65 57.3 ;
        RECT  40.35 52.5 40.95 53.1 ;
        RECT  37.05 53.4 37.65 54.0 ;
        RECT  36.45 48.9 37.05 49.5 ;
        RECT  34.05 53.4 34.65 54.0 ;
        RECT  33.15 56.7 33.75 57.3 ;
        RECT  29.55 52.5 30.15 53.1 ;
        RECT  27.15 52.5 27.75 53.1 ;
        RECT  24.15 54.9 24.75 55.5 ;
        RECT  70.35 42.9 70.95 43.5 ;
        RECT  65.85 45.3 66.45 45.9 ;
        RECT  62.55 44.4 63.15 45.0 ;
        RECT  61.95 48.9 62.55 49.5 ;
        RECT  60.45 44.4 61.05 45.0 ;
        RECT  59.55 41.1 60.15 41.7 ;
        RECT  55.95 45.3 56.55 45.9 ;
        RECT  53.55 45.3 54.15 45.9 ;
        RECT  50.55 42.9 51.15 43.5 ;
        RECT  47.25 43.8 47.85 44.4 ;
        RECT  46.05 41.1 46.65 41.7 ;
        RECT  40.35 45.3 40.95 45.9 ;
        RECT  37.05 44.4 37.65 45.0 ;
        RECT  36.45 48.9 37.05 49.5 ;
        RECT  34.05 44.4 34.65 45.0 ;
        RECT  33.15 41.1 33.75 41.7 ;
        RECT  29.55 45.3 30.15 45.9 ;
        RECT  27.15 45.3 27.75 45.9 ;
        RECT  24.15 42.9 24.75 43.5 ;
        RECT  91.35 89.1 91.95 89.7 ;
        RECT  88.65 105.0 89.25 105.6 ;
        RECT  85.95 147.9 86.55 148.5 ;
        RECT  83.25 163.8 83.85 164.4 ;
        RECT  114.75 33.6 115.35 34.2 ;
        RECT  109.35 28.95 109.95 29.55 ;
        RECT  112.05 26.55 112.65 27.15 ;
        RECT  114.75 446.7 115.35 447.3 ;
        RECT  117.45 98.25 118.05 98.85 ;
        RECT  120.15 196.35 120.75 196.95 ;
        RECT  17.25 76.8 17.85 77.4 ;
        RECT  106.65 456.9 107.25 457.5 ;
        RECT  95.85 437.4 96.45 438.0 ;
        RECT  97.05 437.4 97.65 438.0 ;
        RECT  134.55 437.4 135.15 438.0 ;
        RECT  144.75 437.4 145.35 438.0 ;
        RECT  123.45 437.4 124.05 438.0 ;
        RECT  102.45 8.4 103.05 9.0 ;
        RECT  103.65 8.4 104.25 9.0 ;
        RECT  134.25 8.4 134.85 9.0 ;
        RECT  134.25 8.4 134.85 9.0 ;
        RECT  88.5 229.35 89.1 229.95 ;
        RECT  88.5 258.75 89.1 259.35 ;
        RECT  88.5 288.15 89.1 288.75 ;
        RECT  88.5 317.55 89.1 318.15 ;
        RECT  88.5 346.95 89.1 347.55 ;
        RECT  88.5 376.35 89.1 376.95 ;
        RECT  88.5 405.75 89.1 406.35 ;
        RECT  88.5 435.15 89.1 435.75 ;
        RECT  95.85 140.85 96.45 141.45 ;
        RECT  97.05 140.85 97.65 141.45 ;
        RECT  95.85 199.65 96.45 200.25 ;
        RECT  97.05 199.65 97.65 200.25 ;
        RECT  75.75 69.45 76.35 70.05 ;
        RECT  95.85 69.45 96.45 70.05 ;
        RECT  97.05 69.45 97.65 70.05 ;
        RECT  75.75 69.45 76.35 70.05 ;
        RECT  95.85 69.45 96.45 70.05 ;
        RECT  97.05 69.45 97.65 70.05 ;
        RECT  75.75 49.05 76.35 49.65 ;
        RECT  95.85 49.05 96.45 49.65 ;
        RECT  97.05 49.05 97.65 49.65 ;
        RECT  75.75 49.05 76.35 49.65 ;
        RECT  95.85 49.05 96.45 49.65 ;
        RECT  97.05 49.05 97.65 49.65 ;
        RECT  -62.4 140.1 -61.8 140.7 ;
        RECT  -60.0 135.6 -59.4 136.2 ;
        RECT  -60.9 132.3 -60.3 132.9 ;
        RECT  -56.4 131.7 -55.8 132.3 ;
        RECT  -60.9 130.2 -60.3 130.8 ;
        RECT  -64.2 129.3 -63.6 129.9 ;
        RECT  -60.0 125.7 -59.4 126.3 ;
        RECT  -60.0 123.3 -59.4 123.9 ;
        RECT  -62.4 120.3 -61.8 120.9 ;
        RECT  -61.5 117.0 -60.9 117.6 ;
        RECT  -64.2 115.8 -63.6 116.4 ;
        RECT  -60.0 110.1 -59.4 110.7 ;
        RECT  -60.9 106.8 -60.3 107.4 ;
        RECT  -56.4 106.2 -55.8 106.8 ;
        RECT  -60.9 103.8 -60.3 104.4 ;
        RECT  -64.2 102.9 -63.6 103.5 ;
        RECT  -60.0 99.3 -59.4 99.9 ;
        RECT  -60.0 96.9 -59.4 97.5 ;
        RECT  -62.4 93.9 -61.8 94.5 ;
        RECT  -50.4 140.1 -49.8 140.7 ;
        RECT  -52.8 135.6 -52.2 136.2 ;
        RECT  -51.9 132.3 -51.3 132.9 ;
        RECT  -56.4 131.7 -55.8 132.3 ;
        RECT  -51.9 130.2 -51.3 130.8 ;
        RECT  -48.6 129.3 -48.0 129.9 ;
        RECT  -52.8 125.7 -52.2 126.3 ;
        RECT  -52.8 123.3 -52.2 123.9 ;
        RECT  -50.4 120.3 -49.8 120.9 ;
        RECT  -51.3 117.0 -50.7 117.6 ;
        RECT  -48.6 115.8 -48.0 116.4 ;
        RECT  -52.8 110.1 -52.2 110.7 ;
        RECT  -51.9 106.8 -51.3 107.4 ;
        RECT  -56.4 106.2 -55.8 106.8 ;
        RECT  -51.9 103.8 -51.3 104.4 ;
        RECT  -48.6 102.9 -48.0 103.5 ;
        RECT  -52.8 99.3 -52.2 99.9 ;
        RECT  -52.8 96.9 -52.2 97.5 ;
        RECT  -50.4 93.9 -49.8 94.5 ;
        RECT  -42.0 140.1 -41.4 140.7 ;
        RECT  -39.6 135.6 -39.0 136.2 ;
        RECT  -40.5 132.3 -39.9 132.9 ;
        RECT  -36.0 131.7 -35.4 132.3 ;
        RECT  -40.5 130.2 -39.9 130.8 ;
        RECT  -43.8 129.3 -43.2 129.9 ;
        RECT  -39.6 125.7 -39.0 126.3 ;
        RECT  -39.6 123.3 -39.0 123.9 ;
        RECT  -42.0 120.3 -41.4 120.9 ;
        RECT  -41.1 117.0 -40.5 117.6 ;
        RECT  -43.8 115.8 -43.2 116.4 ;
        RECT  -39.6 110.1 -39.0 110.7 ;
        RECT  -40.5 106.8 -39.9 107.4 ;
        RECT  -36.0 106.2 -35.4 106.8 ;
        RECT  -40.5 103.8 -39.9 104.4 ;
        RECT  -43.8 102.9 -43.2 103.5 ;
        RECT  -39.6 99.3 -39.0 99.9 ;
        RECT  -39.6 96.9 -39.0 97.5 ;
        RECT  -42.0 93.9 -41.4 94.5 ;
        RECT  -19.35 100.2 -18.75 100.8 ;
        RECT  -12.75 100.2 -12.15 100.8 ;
        RECT  -19.35 95.4 -18.75 96.0 ;
        RECT  -12.75 95.4 -12.15 96.0 ;
        RECT  -14.55 266.7 -13.95 267.3 ;
        RECT  -14.55 257.1 -13.95 257.7 ;
        RECT  -31.35 248.7 -30.75 249.3 ;
        RECT  -31.35 258.3 -30.75 258.9 ;
        RECT  -14.55 261.3 -13.95 261.9 ;
        RECT  -14.55 251.7 -13.95 252.3 ;
        RECT  -31.35 254.1 -30.75 254.7 ;
        RECT  -53.25 264.3 -52.65 264.9 ;
        RECT  -62.25 264.3 -61.65 264.9 ;
        RECT  -54.15 255.0 -53.55 255.6 ;
        RECT  -58.35 255.0 -57.75 255.6 ;
        RECT  -53.25 244.5 -52.65 245.1 ;
        RECT  -62.25 244.5 -61.65 245.1 ;
        RECT  -54.15 253.8 -53.55 254.4 ;
        RECT  -58.35 253.8 -57.75 254.4 ;
        RECT  -53.25 234.9 -52.65 235.5 ;
        RECT  -62.25 234.9 -61.65 235.5 ;
        RECT  -54.15 225.6 -53.55 226.2 ;
        RECT  -58.35 225.6 -57.75 226.2 ;
        RECT  -42.75 236.25 -42.15 236.85 ;
        RECT  -32.55 233.55 -31.95 234.15 ;
        RECT  -44.85 233.55 -44.25 234.15 ;
        RECT  -55.65 235.65 -55.05 236.25 ;
        RECT  -13.5 260.7 -12.9 261.3 ;
        RECT  -31.95 260.7 -31.35 261.3 ;
        RECT  -32.55 272.1 -31.95 272.7 ;
        RECT  -13.5 240.45 -12.9 241.05 ;
        RECT  -49.95 250.5 -49.35 251.1 ;
        RECT  -45.75 244.2 -45.15 244.8 ;
        RECT  -45.75 264.3 -45.15 264.9 ;
        RECT  -8.25 229.5 -7.65 230.1 ;
        RECT  -8.25 287.1 -7.65 287.7 ;
        RECT  -37.65 287.1 -37.05 287.7 ;
        RECT  -46.35 293.55 -45.75 294.15 ;
        RECT  -43.05 266.55 -42.45 267.15 ;
        RECT  -43.05 255.9 -42.45 256.5 ;
        RECT  -45.75 267.3 -45.15 267.9 ;
        RECT  -43.05 266.55 -42.45 267.15 ;
        RECT  -43.05 279.9 -42.45 280.5 ;
        RECT  -45.75 239.1 -45.15 239.7 ;
        RECT  -62.25 229.5 -61.65 230.1 ;
        RECT  -52.05 229.5 -51.45 230.1 ;
        RECT  -25.95 170.1 -25.35 170.7 ;
        RECT  -25.95 174.9 -25.35 175.5 ;
        RECT  -32.7 171.0 -32.1 171.6 ;
        RECT  -33.6 165.6 -33.0 166.2 ;
        RECT  -32.7 173.4 -32.1 174.0 ;
        RECT  -35.7 165.6 -35.1 166.2 ;
        RECT  -49.65 170.1 -49.05 170.7 ;
        RECT  -49.65 174.9 -49.05 175.5 ;
        RECT  -42.9 171.0 -42.3 171.6 ;
        RECT  -42.0 165.6 -41.4 166.2 ;
        RECT  -42.9 173.4 -42.3 174.0 ;
        RECT  -39.9 165.6 -39.3 166.2 ;
        RECT  -40.5 144.6 -39.9 145.2 ;
        RECT  -40.5 151.2 -39.9 151.8 ;
        RECT  -43.95 144.6 -43.35 145.2 ;
        RECT  -43.95 153.9 -43.35 154.5 ;
        RECT  -64.35 144.6 -63.75 145.2 ;
        RECT  -64.35 156.6 -63.75 157.2 ;
        RECT  -48.75 144.6 -48.15 145.2 ;
        RECT  -48.75 159.3 -48.15 159.9 ;
        RECT  -17.1 153.9 -16.5 154.5 ;
        RECT  -13.8 162.0 -13.2 162.6 ;
        RECT  -27.15 162.0 -26.55 162.6 ;
        RECT  -32.7 153.9 -32.1 154.5 ;
        RECT  -34.5 156.6 -33.9 157.2 ;
        RECT  -47.55 162.0 -46.95 162.6 ;
        RECT  -42.0 159.3 -41.4 159.9 ;
        RECT  -40.2 156.6 -39.6 157.2 ;
        RECT  -15.9 121.2 -15.3 121.8 ;
        RECT  -5.55 121.2 -4.95 121.8 ;
        RECT  -5.55 151.05 -4.95 151.65 ;
        RECT  -30.6 214.5 -30.0 215.1 ;
        RECT  -44.1 211.8 -43.5 212.4 ;
        RECT  -14.7 217.2 -14.1 217.8 ;
        RECT  -3.75 214.35 -3.15 214.95 ;
        RECT  -22.65 219.9 -22.05 220.5 ;
        RECT  -52.05 219.9 -51.45 220.5 ;
        RECT  -7.95 148.5 -7.35 149.1 ;
        RECT  -14.55 126.6 -13.95 127.2 ;
        RECT  -27.45 126.6 -26.85 127.2 ;
        RECT  -27.3 85.8 -26.7 86.4 ;
        RECT  -13.8 88.8 -13.2 89.4 ;
        RECT  -14.7 175.8 -14.1 176.4 ;
        RECT  -14.7 180.3 -14.1 180.9 ;
        RECT  0.75 219.9 1.35 220.5 ;
        RECT  1.95 219.9 2.55 220.5 ;
        Layer  metal2 ; 
        RECT  -7.5 219.6 0.45 220.5 ;
        RECT  95.55 0.0 104.55 459.3 ;
        RECT  119.85 0.0 120.75 459.3 ;
        RECT  117.15 0.0 118.05 459.3 ;
        RECT  114.45 0.0 115.35 459.3 ;
        RECT  111.75 0.0 112.65 459.3 ;
        RECT  109.05 0.0 109.95 459.3 ;
        RECT  106.35 0.0 107.25 459.3 ;
        RECT  91.05 39.0 91.95 196.5 ;
        RECT  88.35 39.0 89.25 196.5 ;
        RECT  85.65 39.0 86.55 196.5 ;
        RECT  82.95 39.0 83.85 196.5 ;
        RECT  127.5 435.3 128.4 439.8 ;
        RECT  130.5 435.3 131.4 439.8 ;
        RECT  137.7 435.3 138.6 439.8 ;
        RECT  140.7 435.3 141.6 439.8 ;
        RECT  129.0 6.0 129.9 6.9 ;
        RECT  124.95 6.0 129.45 6.9 ;
        RECT  129.0 6.45 129.9 12.45 ;
        RECT  139.2 6.0 140.1 6.9 ;
        RECT  135.15 6.0 139.65 6.9 ;
        RECT  139.2 6.45 140.1 12.45 ;
        RECT  114.45 200.1 115.35 448.2 ;
        RECT  134.1 435.3 135.0 438.0 ;
        RECT  144.3 435.3 145.2 438.0 ;
        RECT  123.45 200.1 124.35 438.0 ;
        RECT  88.95 229.05 95.55 229.95 ;
        RECT  88.95 258.45 95.55 259.35 ;
        RECT  88.95 287.85 95.55 288.75 ;
        RECT  88.95 317.25 95.55 318.15 ;
        RECT  88.95 346.65 95.55 347.55 ;
        RECT  88.95 376.05 95.55 376.95 ;
        RECT  88.95 405.45 95.55 406.35 ;
        RECT  88.95 434.85 95.55 435.75 ;
        RECT  123.75 204.3 126.15 214.8 ;
        RECT  127.35 201.3 128.55 214.8 ;
        RECT  130.35 201.3 131.55 214.8 ;
        RECT  125.85 200.1 128.55 201.3 ;
        RECT  130.05 200.1 131.55 201.3 ;
        RECT  133.95 200.1 135.15 214.8 ;
        RECT  123.75 214.8 126.15 225.3 ;
        RECT  127.35 214.8 128.55 228.3 ;
        RECT  130.35 214.8 131.55 228.3 ;
        RECT  125.85 228.3 128.55 229.5 ;
        RECT  130.05 228.3 131.55 229.5 ;
        RECT  133.95 214.8 135.15 229.5 ;
        RECT  123.75 233.7 126.15 244.2 ;
        RECT  127.35 230.7 128.55 244.2 ;
        RECT  130.35 230.7 131.55 244.2 ;
        RECT  125.85 229.5 128.55 230.7 ;
        RECT  130.05 229.5 131.55 230.7 ;
        RECT  133.95 229.5 135.15 244.2 ;
        RECT  123.75 244.2 126.15 254.7 ;
        RECT  127.35 244.2 128.55 257.7 ;
        RECT  130.35 244.2 131.55 257.7 ;
        RECT  125.85 257.7 128.55 258.9 ;
        RECT  130.05 257.7 131.55 258.9 ;
        RECT  133.95 244.2 135.15 258.9 ;
        RECT  123.75 263.1 126.15 273.6 ;
        RECT  127.35 260.1 128.55 273.6 ;
        RECT  130.35 260.1 131.55 273.6 ;
        RECT  125.85 258.9 128.55 260.1 ;
        RECT  130.05 258.9 131.55 260.1 ;
        RECT  133.95 258.9 135.15 273.6 ;
        RECT  123.75 273.6 126.15 284.1 ;
        RECT  127.35 273.6 128.55 287.1 ;
        RECT  130.35 273.6 131.55 287.1 ;
        RECT  125.85 287.1 128.55 288.3 ;
        RECT  130.05 287.1 131.55 288.3 ;
        RECT  133.95 273.6 135.15 288.3 ;
        RECT  123.75 292.5 126.15 303.0 ;
        RECT  127.35 289.5 128.55 303.0 ;
        RECT  130.35 289.5 131.55 303.0 ;
        RECT  125.85 288.3 128.55 289.5 ;
        RECT  130.05 288.3 131.55 289.5 ;
        RECT  133.95 288.3 135.15 303.0 ;
        RECT  123.75 303.0 126.15 313.5 ;
        RECT  127.35 303.0 128.55 316.5 ;
        RECT  130.35 303.0 131.55 316.5 ;
        RECT  125.85 316.5 128.55 317.7 ;
        RECT  130.05 316.5 131.55 317.7 ;
        RECT  133.95 303.0 135.15 317.7 ;
        RECT  123.75 321.9 126.15 332.4 ;
        RECT  127.35 318.9 128.55 332.4 ;
        RECT  130.35 318.9 131.55 332.4 ;
        RECT  125.85 317.7 128.55 318.9 ;
        RECT  130.05 317.7 131.55 318.9 ;
        RECT  133.95 317.7 135.15 332.4 ;
        RECT  123.75 332.4 126.15 342.9 ;
        RECT  127.35 332.4 128.55 345.9 ;
        RECT  130.35 332.4 131.55 345.9 ;
        RECT  125.85 345.9 128.55 347.1 ;
        RECT  130.05 345.9 131.55 347.1 ;
        RECT  133.95 332.4 135.15 347.1 ;
        RECT  123.75 351.3 126.15 361.8 ;
        RECT  127.35 348.3 128.55 361.8 ;
        RECT  130.35 348.3 131.55 361.8 ;
        RECT  125.85 347.1 128.55 348.3 ;
        RECT  130.05 347.1 131.55 348.3 ;
        RECT  133.95 347.1 135.15 361.8 ;
        RECT  123.75 361.8 126.15 372.3 ;
        RECT  127.35 361.8 128.55 375.3 ;
        RECT  130.35 361.8 131.55 375.3 ;
        RECT  125.85 375.3 128.55 376.5 ;
        RECT  130.05 375.3 131.55 376.5 ;
        RECT  133.95 361.8 135.15 376.5 ;
        RECT  123.75 380.7 126.15 391.2 ;
        RECT  127.35 377.7 128.55 391.2 ;
        RECT  130.35 377.7 131.55 391.2 ;
        RECT  125.85 376.5 128.55 377.7 ;
        RECT  130.05 376.5 131.55 377.7 ;
        RECT  133.95 376.5 135.15 391.2 ;
        RECT  123.75 391.2 126.15 401.7 ;
        RECT  127.35 391.2 128.55 404.7 ;
        RECT  130.35 391.2 131.55 404.7 ;
        RECT  125.85 404.7 128.55 405.9 ;
        RECT  130.05 404.7 131.55 405.9 ;
        RECT  133.95 391.2 135.15 405.9 ;
        RECT  123.75 410.1 126.15 420.6 ;
        RECT  127.35 407.1 128.55 420.6 ;
        RECT  130.35 407.1 131.55 420.6 ;
        RECT  125.85 405.9 128.55 407.1 ;
        RECT  130.05 405.9 131.55 407.1 ;
        RECT  133.95 405.9 135.15 420.6 ;
        RECT  123.75 420.6 126.15 431.1 ;
        RECT  127.35 420.6 128.55 434.1 ;
        RECT  130.35 420.6 131.55 434.1 ;
        RECT  125.85 434.1 128.55 435.3 ;
        RECT  130.05 434.1 131.55 435.3 ;
        RECT  133.95 420.6 135.15 435.3 ;
        RECT  133.95 204.3 136.35 214.8 ;
        RECT  137.55 201.3 138.75 214.8 ;
        RECT  140.55 201.3 141.75 214.8 ;
        RECT  136.05 200.1 138.75 201.3 ;
        RECT  140.25 200.1 141.75 201.3 ;
        RECT  144.15 200.1 145.35 214.8 ;
        RECT  133.95 214.8 136.35 225.3 ;
        RECT  137.55 214.8 138.75 228.3 ;
        RECT  140.55 214.8 141.75 228.3 ;
        RECT  136.05 228.3 138.75 229.5 ;
        RECT  140.25 228.3 141.75 229.5 ;
        RECT  144.15 214.8 145.35 229.5 ;
        RECT  133.95 233.7 136.35 244.2 ;
        RECT  137.55 230.7 138.75 244.2 ;
        RECT  140.55 230.7 141.75 244.2 ;
        RECT  136.05 229.5 138.75 230.7 ;
        RECT  140.25 229.5 141.75 230.7 ;
        RECT  144.15 229.5 145.35 244.2 ;
        RECT  133.95 244.2 136.35 254.7 ;
        RECT  137.55 244.2 138.75 257.7 ;
        RECT  140.55 244.2 141.75 257.7 ;
        RECT  136.05 257.7 138.75 258.9 ;
        RECT  140.25 257.7 141.75 258.9 ;
        RECT  144.15 244.2 145.35 258.9 ;
        RECT  133.95 263.1 136.35 273.6 ;
        RECT  137.55 260.1 138.75 273.6 ;
        RECT  140.55 260.1 141.75 273.6 ;
        RECT  136.05 258.9 138.75 260.1 ;
        RECT  140.25 258.9 141.75 260.1 ;
        RECT  144.15 258.9 145.35 273.6 ;
        RECT  133.95 273.6 136.35 284.1 ;
        RECT  137.55 273.6 138.75 287.1 ;
        RECT  140.55 273.6 141.75 287.1 ;
        RECT  136.05 287.1 138.75 288.3 ;
        RECT  140.25 287.1 141.75 288.3 ;
        RECT  144.15 273.6 145.35 288.3 ;
        RECT  133.95 292.5 136.35 303.0 ;
        RECT  137.55 289.5 138.75 303.0 ;
        RECT  140.55 289.5 141.75 303.0 ;
        RECT  136.05 288.3 138.75 289.5 ;
        RECT  140.25 288.3 141.75 289.5 ;
        RECT  144.15 288.3 145.35 303.0 ;
        RECT  133.95 303.0 136.35 313.5 ;
        RECT  137.55 303.0 138.75 316.5 ;
        RECT  140.55 303.0 141.75 316.5 ;
        RECT  136.05 316.5 138.75 317.7 ;
        RECT  140.25 316.5 141.75 317.7 ;
        RECT  144.15 303.0 145.35 317.7 ;
        RECT  133.95 321.9 136.35 332.4 ;
        RECT  137.55 318.9 138.75 332.4 ;
        RECT  140.55 318.9 141.75 332.4 ;
        RECT  136.05 317.7 138.75 318.9 ;
        RECT  140.25 317.7 141.75 318.9 ;
        RECT  144.15 317.7 145.35 332.4 ;
        RECT  133.95 332.4 136.35 342.9 ;
        RECT  137.55 332.4 138.75 345.9 ;
        RECT  140.55 332.4 141.75 345.9 ;
        RECT  136.05 345.9 138.75 347.1 ;
        RECT  140.25 345.9 141.75 347.1 ;
        RECT  144.15 332.4 145.35 347.1 ;
        RECT  133.95 351.3 136.35 361.8 ;
        RECT  137.55 348.3 138.75 361.8 ;
        RECT  140.55 348.3 141.75 361.8 ;
        RECT  136.05 347.1 138.75 348.3 ;
        RECT  140.25 347.1 141.75 348.3 ;
        RECT  144.15 347.1 145.35 361.8 ;
        RECT  133.95 361.8 136.35 372.3 ;
        RECT  137.55 361.8 138.75 375.3 ;
        RECT  140.55 361.8 141.75 375.3 ;
        RECT  136.05 375.3 138.75 376.5 ;
        RECT  140.25 375.3 141.75 376.5 ;
        RECT  144.15 361.8 145.35 376.5 ;
        RECT  133.95 380.7 136.35 391.2 ;
        RECT  137.55 377.7 138.75 391.2 ;
        RECT  140.55 377.7 141.75 391.2 ;
        RECT  136.05 376.5 138.75 377.7 ;
        RECT  140.25 376.5 141.75 377.7 ;
        RECT  144.15 376.5 145.35 391.2 ;
        RECT  133.95 391.2 136.35 401.7 ;
        RECT  137.55 391.2 138.75 404.7 ;
        RECT  140.55 391.2 141.75 404.7 ;
        RECT  136.05 404.7 138.75 405.9 ;
        RECT  140.25 404.7 141.75 405.9 ;
        RECT  144.15 391.2 145.35 405.9 ;
        RECT  133.95 410.1 136.35 420.6 ;
        RECT  137.55 407.1 138.75 420.6 ;
        RECT  140.55 407.1 141.75 420.6 ;
        RECT  136.05 405.9 138.75 407.1 ;
        RECT  140.25 405.9 141.75 407.1 ;
        RECT  144.15 405.9 145.35 420.6 ;
        RECT  133.95 420.6 136.35 431.1 ;
        RECT  137.55 420.6 138.75 434.1 ;
        RECT  140.55 420.6 141.75 434.1 ;
        RECT  136.05 434.1 138.75 435.3 ;
        RECT  140.25 434.1 141.75 435.3 ;
        RECT  144.15 420.6 145.35 435.3 ;
        RECT  127.5 439.8 128.4 459.3 ;
        RECT  130.5 439.8 131.4 459.3 ;
        RECT  127.8 450.9 127.95 452.1 ;
        RECT  130.5 450.9 132.15 452.1 ;
        RECT  127.8 442.5 127.95 443.7 ;
        RECT  129.75 442.5 130.5 443.7 ;
        RECT  127.35 450.9 128.55 452.1 ;
        RECT  132.15 450.9 133.35 452.1 ;
        RECT  127.35 442.5 128.55 443.7 ;
        RECT  129.75 442.5 130.95 443.7 ;
        RECT  137.7 439.8 138.6 459.3 ;
        RECT  140.7 439.8 141.6 459.3 ;
        RECT  138.0 450.9 138.15 452.1 ;
        RECT  140.7 450.9 142.35 452.1 ;
        RECT  138.0 442.5 138.15 443.7 ;
        RECT  139.95 442.5 140.7 443.7 ;
        RECT  137.55 450.9 138.75 452.1 ;
        RECT  142.35 450.9 143.55 452.1 ;
        RECT  137.55 442.5 138.75 443.7 ;
        RECT  139.95 442.5 141.15 443.7 ;
        RECT  127.35 165.6 128.55 200.1 ;
        RECT  130.35 165.6 131.55 200.1 ;
        RECT  133.95 192.6 135.15 200.1 ;
        RECT  127.35 164.4 129.45 165.6 ;
        RECT  130.35 164.4 132.15 165.6 ;
        RECT  125.25 151.2 126.45 155.7 ;
        RECT  127.35 151.2 128.55 164.4 ;
        RECT  130.35 151.2 131.55 164.4 ;
        RECT  137.55 165.6 138.75 200.1 ;
        RECT  140.55 165.6 141.75 200.1 ;
        RECT  144.15 192.6 145.35 200.1 ;
        RECT  137.55 164.4 139.65 165.6 ;
        RECT  140.55 164.4 142.35 165.6 ;
        RECT  135.45 151.2 136.65 155.7 ;
        RECT  137.55 151.2 138.75 164.4 ;
        RECT  140.55 151.2 141.75 164.4 ;
        RECT  127.35 149.1 128.55 151.2 ;
        RECT  125.85 147.9 128.55 149.1 ;
        RECT  130.35 143.7 131.55 151.2 ;
        RECT  133.95 138.9 135.15 149.4 ;
        RECT  127.65 137.7 135.15 138.9 ;
        RECT  126.75 99.9 127.95 127.2 ;
        RECT  133.95 116.4 135.15 137.7 ;
        RECT  133.35 115.2 135.15 116.4 ;
        RECT  133.95 112.2 135.15 115.2 ;
        RECT  130.05 111.0 135.15 112.2 ;
        RECT  130.05 109.8 131.25 111.0 ;
        RECT  127.95 93.6 130.35 94.8 ;
        RECT  128.85 90.9 130.05 93.6 ;
        RECT  133.95 90.9 135.15 111.0 ;
        RECT  137.55 149.1 138.75 151.2 ;
        RECT  136.05 147.9 138.75 149.1 ;
        RECT  140.55 143.7 141.75 151.2 ;
        RECT  144.15 138.9 145.35 149.4 ;
        RECT  137.85 137.7 145.35 138.9 ;
        RECT  136.95 99.9 138.15 127.2 ;
        RECT  144.15 116.4 145.35 137.7 ;
        RECT  143.55 115.2 145.35 116.4 ;
        RECT  144.15 112.2 145.35 115.2 ;
        RECT  140.25 111.0 145.35 112.2 ;
        RECT  140.25 109.8 141.45 111.0 ;
        RECT  138.15 93.6 140.55 94.8 ;
        RECT  139.05 90.9 140.25 93.6 ;
        RECT  144.15 90.9 145.35 111.0 ;
        RECT  126.15 86.4 127.35 90.9 ;
        RECT  128.85 89.7 130.05 90.9 ;
        RECT  128.85 88.5 131.55 89.7 ;
        RECT  126.15 85.2 129.15 86.4 ;
        RECT  126.15 75.6 127.05 85.2 ;
        RECT  130.35 80.7 131.55 88.5 ;
        RECT  129.45 77.4 132.45 78.6 ;
        RECT  126.15 74.4 127.35 75.6 ;
        RECT  129.45 75.3 130.65 76.5 ;
        RECT  129.75 73.8 130.65 75.3 ;
        RECT  128.25 72.9 130.65 73.8 ;
        RECT  128.25 66.6 129.15 72.9 ;
        RECT  131.55 72.0 132.45 77.4 ;
        RECT  130.35 70.8 132.45 72.0 ;
        RECT  130.35 68.4 132.45 69.6 ;
        RECT  127.95 65.4 129.15 66.6 ;
        RECT  125.85 60.9 127.35 62.1 ;
        RECT  125.85 49.2 126.75 60.9 ;
        RECT  128.85 58.8 130.05 63.3 ;
        RECT  127.65 57.9 130.05 58.8 ;
        RECT  127.65 51.0 128.55 57.9 ;
        RECT  131.55 56.4 132.45 68.4 ;
        RECT  130.35 55.2 132.45 56.4 ;
        RECT  129.45 51.9 132.45 53.1 ;
        RECT  127.65 50.1 129.15 51.0 ;
        RECT  125.85 48.0 127.35 49.2 ;
        RECT  128.25 48.9 130.65 50.1 ;
        RECT  128.25 40.2 129.15 48.9 ;
        RECT  131.55 45.6 132.45 51.9 ;
        RECT  130.35 44.4 132.45 45.6 ;
        RECT  130.35 42.0 132.45 43.2 ;
        RECT  127.95 39.0 129.15 40.2 ;
        RECT  131.55 33.3 132.45 42.0 ;
        RECT  128.85 32.1 132.45 33.3 ;
        RECT  128.85 30.9 130.05 32.1 ;
        RECT  133.95 30.9 135.15 90.9 ;
        RECT  141.75 86.4 142.95 90.9 ;
        RECT  139.05 89.7 140.25 90.9 ;
        RECT  137.55 88.5 140.25 89.7 ;
        RECT  139.95 85.2 142.95 86.4 ;
        RECT  142.05 75.6 142.95 85.2 ;
        RECT  137.55 80.7 138.75 88.5 ;
        RECT  136.65 77.4 139.65 78.6 ;
        RECT  141.75 74.4 142.95 75.6 ;
        RECT  138.45 75.3 139.65 76.5 ;
        RECT  138.45 73.8 139.35 75.3 ;
        RECT  138.45 72.9 140.85 73.8 ;
        RECT  139.95 66.6 140.85 72.9 ;
        RECT  136.65 72.0 137.55 77.4 ;
        RECT  136.65 70.8 138.75 72.0 ;
        RECT  136.65 68.4 138.75 69.6 ;
        RECT  139.95 65.4 141.15 66.6 ;
        RECT  141.75 60.9 143.25 62.1 ;
        RECT  142.35 49.2 143.25 60.9 ;
        RECT  139.05 58.8 140.25 63.3 ;
        RECT  139.05 57.9 141.45 58.8 ;
        RECT  140.55 51.0 141.45 57.9 ;
        RECT  136.65 56.4 137.55 68.4 ;
        RECT  136.65 55.2 138.75 56.4 ;
        RECT  136.65 51.9 139.65 53.1 ;
        RECT  139.95 50.1 141.45 51.0 ;
        RECT  141.75 48.0 143.25 49.2 ;
        RECT  138.45 48.9 140.85 50.1 ;
        RECT  139.95 40.2 140.85 48.9 ;
        RECT  136.65 45.6 137.55 51.9 ;
        RECT  136.65 44.4 138.75 45.6 ;
        RECT  136.65 42.0 138.75 43.2 ;
        RECT  139.95 39.0 141.15 40.2 ;
        RECT  136.65 33.3 137.55 42.0 ;
        RECT  136.65 32.1 140.25 33.3 ;
        RECT  139.05 30.9 140.25 32.1 ;
        RECT  133.95 30.9 135.15 90.9 ;
        RECT  128.85 45.9 130.05 52.8 ;
        RECT  127.05 44.7 130.05 45.9 ;
        RECT  128.85 41.1 133.05 42.3 ;
        RECT  128.85 33.6 130.05 41.1 ;
        RECT  128.85 32.4 130.35 33.6 ;
        RECT  128.85 30.9 130.05 32.4 ;
        RECT  133.95 30.9 135.15 52.8 ;
        RECT  139.05 45.9 140.25 52.8 ;
        RECT  139.05 44.7 142.05 45.9 ;
        RECT  136.05 41.1 140.25 42.3 ;
        RECT  139.05 33.6 140.25 41.1 ;
        RECT  138.75 32.4 140.25 33.6 ;
        RECT  139.05 30.9 140.25 32.4 ;
        RECT  133.95 30.9 135.15 52.8 ;
        RECT  27.75 82.5 28.65 435.3 ;
        RECT  25.65 82.5 26.55 435.3 ;
        RECT  23.55 82.5 24.45 435.3 ;
        RECT  21.45 82.5 22.35 435.3 ;
        RECT  19.35 82.5 20.25 435.3 ;
        RECT  17.25 82.5 18.15 435.3 ;
        RECT  15.15 82.5 16.05 435.3 ;
        RECT  13.05 82.5 13.95 435.3 ;
        RECT  78.15 82.5 79.05 138.6 ;
        RECT  76.05 82.5 76.95 138.6 ;
        RECT  63.15 82.5 64.05 138.6 ;
        RECT  61.05 82.5 61.95 138.6 ;
        RECT  58.95 82.5 59.85 138.6 ;
        RECT  56.85 82.5 57.75 138.6 ;
        RECT  54.75 82.5 55.65 138.6 ;
        RECT  52.65 82.5 53.55 138.6 ;
        RECT  58.65 92.85 59.85 94.05 ;
        RECT  77.85 87.6 79.05 88.8 ;
        RECT  56.55 98.25 57.75 99.45 ;
        RECT  75.75 103.5 76.95 104.7 ;
        RECT  58.65 90.0 59.85 91.2 ;
        RECT  56.55 86.7 57.75 87.9 ;
        RECT  54.45 101.1 55.65 102.3 ;
        RECT  56.55 104.4 57.75 105.6 ;
        RECT  58.65 119.4 59.85 120.6 ;
        RECT  52.35 116.1 53.55 117.3 ;
        RECT  54.45 130.5 55.65 131.7 ;
        RECT  77.85 130.5 79.05 131.7 ;
        RECT  52.35 133.8 53.55 135.0 ;
        RECT  75.75 133.8 76.95 135.0 ;
        RECT  60.75 80.85 61.95 82.05 ;
        RECT  62.85 95.55 64.05 96.75 ;
        RECT  60.75 110.25 61.95 111.45 ;
        RECT  62.85 124.95 64.05 126.15 ;
        RECT  60.75 137.4 61.95 138.6 ;
        RECT  78.15 141.3 79.05 197.4 ;
        RECT  76.05 141.3 76.95 197.4 ;
        RECT  63.15 141.3 64.05 197.4 ;
        RECT  61.05 141.3 61.95 197.4 ;
        RECT  58.95 141.3 59.85 197.4 ;
        RECT  56.85 141.3 57.75 197.4 ;
        RECT  54.75 141.3 55.65 197.4 ;
        RECT  52.65 141.3 53.55 197.4 ;
        RECT  58.65 151.65 59.85 152.85 ;
        RECT  77.85 146.4 79.05 147.6 ;
        RECT  56.55 157.05 57.75 158.25 ;
        RECT  75.75 162.3 76.95 163.5 ;
        RECT  58.65 148.8 59.85 150.0 ;
        RECT  56.55 145.5 57.75 146.7 ;
        RECT  54.45 159.9 55.65 161.1 ;
        RECT  56.55 163.2 57.75 164.4 ;
        RECT  58.65 178.2 59.85 179.4 ;
        RECT  52.35 174.9 53.55 176.1 ;
        RECT  54.45 189.3 55.65 190.5 ;
        RECT  77.85 189.3 79.05 190.5 ;
        RECT  52.35 192.6 53.55 193.8 ;
        RECT  75.75 192.6 76.95 193.8 ;
        RECT  60.75 139.65 61.95 140.85 ;
        RECT  62.85 154.35 64.05 155.55 ;
        RECT  60.75 169.05 61.95 170.25 ;
        RECT  62.85 183.75 64.05 184.95 ;
        RECT  60.75 196.2 61.95 197.4 ;
        RECT  13.05 88.8 14.25 90.0 ;
        RECT  15.15 104.7 16.35 105.9 ;
        RECT  17.25 118.2 18.45 119.4 ;
        RECT  19.35 134.1 20.55 135.3 ;
        RECT  21.45 147.6 22.65 148.8 ;
        RECT  23.55 163.5 24.75 164.7 ;
        RECT  25.65 177.0 26.85 178.2 ;
        RECT  27.75 192.9 28.95 194.1 ;
        RECT  13.05 208.8 14.25 210.0 ;
        RECT  21.45 205.5 22.65 206.7 ;
        RECT  13.05 219.9 14.25 221.1 ;
        RECT  23.55 223.2 24.75 224.4 ;
        RECT  13.05 238.2 14.25 239.4 ;
        RECT  25.65 234.9 26.85 236.1 ;
        RECT  13.05 249.3 14.25 250.5 ;
        RECT  27.75 252.6 28.95 253.8 ;
        RECT  15.15 267.6 16.35 268.8 ;
        RECT  21.45 264.3 22.65 265.5 ;
        RECT  15.15 278.7 16.35 279.9 ;
        RECT  23.55 282.0 24.75 283.2 ;
        RECT  15.15 297.0 16.35 298.2 ;
        RECT  25.65 293.7 26.85 294.9 ;
        RECT  15.15 308.1 16.35 309.3 ;
        RECT  27.75 311.4 28.95 312.6 ;
        RECT  17.25 326.4 18.45 327.6 ;
        RECT  21.45 323.1 22.65 324.3 ;
        RECT  17.25 337.5 18.45 338.7 ;
        RECT  23.55 340.8 24.75 342.0 ;
        RECT  17.25 355.8 18.45 357.0 ;
        RECT  25.65 352.5 26.85 353.7 ;
        RECT  17.25 366.9 18.45 368.1 ;
        RECT  27.75 370.2 28.95 371.4 ;
        RECT  19.35 385.2 20.55 386.4 ;
        RECT  21.45 381.9 22.65 383.1 ;
        RECT  19.35 396.3 20.55 397.5 ;
        RECT  23.55 399.6 24.75 400.8 ;
        RECT  19.35 414.6 20.55 415.8 ;
        RECT  25.65 411.3 26.85 412.5 ;
        RECT  19.35 425.7 20.55 426.9 ;
        RECT  27.75 429.0 28.95 430.2 ;
        RECT  51.45 214.35 57.75 215.25 ;
        RECT  51.45 208.8 67.35 209.7 ;
        RECT  51.45 229.05 57.75 229.95 ;
        RECT  51.45 219.9 67.35 220.8 ;
        RECT  51.45 243.75 57.75 244.65 ;
        RECT  51.45 238.2 67.35 239.1 ;
        RECT  51.45 258.45 57.75 259.35 ;
        RECT  51.45 249.3 67.35 250.2 ;
        RECT  51.45 273.15 57.75 274.05 ;
        RECT  51.45 267.6 67.35 268.5 ;
        RECT  51.45 287.85 57.75 288.75 ;
        RECT  51.45 278.7 67.35 279.6 ;
        RECT  51.45 302.55 57.75 303.45 ;
        RECT  51.45 297.0 67.35 297.9 ;
        RECT  51.45 317.25 57.75 318.15 ;
        RECT  51.45 308.1 67.35 309.0 ;
        RECT  51.45 331.95 57.75 332.85 ;
        RECT  51.45 326.4 67.35 327.3 ;
        RECT  51.45 346.65 57.75 347.55 ;
        RECT  51.45 337.5 67.35 338.4 ;
        RECT  51.45 361.35 57.75 362.25 ;
        RECT  51.45 355.8 67.35 356.7 ;
        RECT  51.45 376.05 57.75 376.95 ;
        RECT  51.45 366.9 67.35 367.8 ;
        RECT  51.45 390.75 57.75 391.65 ;
        RECT  51.45 385.2 67.35 386.1 ;
        RECT  51.45 405.45 57.75 406.35 ;
        RECT  51.45 396.3 67.35 397.2 ;
        RECT  51.45 420.15 57.75 421.05 ;
        RECT  51.45 414.6 67.35 415.5 ;
        RECT  51.45 434.85 57.75 435.75 ;
        RECT  51.45 425.7 67.35 426.6 ;
        RECT  51.15 214.35 52.35 215.55 ;
        RECT  57.45 214.35 58.65 215.55 ;
        RECT  67.35 208.8 68.55 210.0 ;
        RECT  51.45 208.8 52.65 210.0 ;
        RECT  51.15 229.05 52.35 230.25 ;
        RECT  57.45 229.05 58.65 230.25 ;
        RECT  67.35 219.6 68.55 220.8 ;
        RECT  51.45 219.6 52.65 220.8 ;
        RECT  51.15 243.75 52.35 244.95 ;
        RECT  57.45 243.75 58.65 244.95 ;
        RECT  67.35 238.2 68.55 239.4 ;
        RECT  51.45 238.2 52.65 239.4 ;
        RECT  51.15 258.45 52.35 259.65 ;
        RECT  57.45 258.45 58.65 259.65 ;
        RECT  67.35 249.0 68.55 250.2 ;
        RECT  51.45 249.0 52.65 250.2 ;
        RECT  51.15 273.15 52.35 274.35 ;
        RECT  57.45 273.15 58.65 274.35 ;
        RECT  67.35 267.6 68.55 268.8 ;
        RECT  51.45 267.6 52.65 268.8 ;
        RECT  51.15 287.85 52.35 289.05 ;
        RECT  57.45 287.85 58.65 289.05 ;
        RECT  67.35 278.4 68.55 279.6 ;
        RECT  51.45 278.4 52.65 279.6 ;
        RECT  51.15 302.55 52.35 303.75 ;
        RECT  57.45 302.55 58.65 303.75 ;
        RECT  67.35 297.0 68.55 298.2 ;
        RECT  51.45 297.0 52.65 298.2 ;
        RECT  51.15 317.25 52.35 318.45 ;
        RECT  57.45 317.25 58.65 318.45 ;
        RECT  67.35 307.8 68.55 309.0 ;
        RECT  51.45 307.8 52.65 309.0 ;
        RECT  51.15 331.95 52.35 333.15 ;
        RECT  57.45 331.95 58.65 333.15 ;
        RECT  67.35 326.4 68.55 327.6 ;
        RECT  51.45 326.4 52.65 327.6 ;
        RECT  51.15 346.65 52.35 347.85 ;
        RECT  57.45 346.65 58.65 347.85 ;
        RECT  67.35 337.2 68.55 338.4 ;
        RECT  51.45 337.2 52.65 338.4 ;
        RECT  51.15 361.35 52.35 362.55 ;
        RECT  57.45 361.35 58.65 362.55 ;
        RECT  67.35 355.8 68.55 357.0 ;
        RECT  51.45 355.8 52.65 357.0 ;
        RECT  51.15 376.05 52.35 377.25 ;
        RECT  57.45 376.05 58.65 377.25 ;
        RECT  67.35 366.6 68.55 367.8 ;
        RECT  51.45 366.6 52.65 367.8 ;
        RECT  51.15 390.75 52.35 391.95 ;
        RECT  57.45 390.75 58.65 391.95 ;
        RECT  67.35 385.2 68.55 386.4 ;
        RECT  51.45 385.2 52.65 386.4 ;
        RECT  51.15 405.45 52.35 406.65 ;
        RECT  57.45 405.45 58.65 406.65 ;
        RECT  67.35 396.0 68.55 397.2 ;
        RECT  51.45 396.0 52.65 397.2 ;
        RECT  51.15 420.15 52.35 421.35 ;
        RECT  57.45 420.15 58.65 421.35 ;
        RECT  67.35 414.6 68.55 415.8 ;
        RECT  51.45 414.6 52.65 415.8 ;
        RECT  51.15 434.85 52.35 436.05 ;
        RECT  57.45 434.85 58.65 436.05 ;
        RECT  67.35 425.4 68.55 426.6 ;
        RECT  51.45 425.4 52.65 426.6 ;
        RECT  71.25 76.8 75.75 78.0 ;
        RECT  74.55 74.1 75.75 75.3 ;
        RECT  73.35 72.6 74.55 75.3 ;
        RECT  70.05 75.0 71.25 78.0 ;
        RECT  60.45 77.1 70.05 78.0 ;
        RECT  65.55 72.6 73.35 73.8 ;
        RECT  62.25 71.7 63.45 74.7 ;
        RECT  59.25 76.8 60.45 78.0 ;
        RECT  60.15 73.5 61.35 74.7 ;
        RECT  58.65 73.5 60.15 74.4 ;
        RECT  57.75 73.5 58.65 75.9 ;
        RECT  51.45 75.0 57.75 75.9 ;
        RECT  56.85 71.7 62.25 72.6 ;
        RECT  55.65 71.7 56.85 73.8 ;
        RECT  53.25 71.7 54.45 73.8 ;
        RECT  50.25 75.0 51.45 76.2 ;
        RECT  45.75 76.8 46.95 78.3 ;
        RECT  34.05 77.4 45.75 78.3 ;
        RECT  43.65 74.1 48.15 75.3 ;
        RECT  42.75 74.1 43.65 76.5 ;
        RECT  35.85 75.6 42.75 76.5 ;
        RECT  41.25 71.7 53.25 72.6 ;
        RECT  40.05 71.7 41.25 73.8 ;
        RECT  36.75 71.7 37.95 74.7 ;
        RECT  34.95 75.0 35.85 76.5 ;
        RECT  32.85 76.8 34.05 78.3 ;
        RECT  33.75 73.5 34.95 75.9 ;
        RECT  25.05 75.0 33.75 75.9 ;
        RECT  30.45 71.7 36.75 72.6 ;
        RECT  29.25 71.7 30.45 73.8 ;
        RECT  26.85 71.7 28.05 73.8 ;
        RECT  23.85 75.0 25.05 76.2 ;
        RECT  18.15 71.7 26.85 72.6 ;
        RECT  16.95 71.7 18.15 75.3 ;
        RECT  15.75 74.1 16.95 75.3 ;
        RECT  15.75 69.0 75.75 70.2 ;
        RECT  71.25 61.2 75.75 62.4 ;
        RECT  74.55 63.9 75.75 65.1 ;
        RECT  73.35 63.9 74.55 66.6 ;
        RECT  70.05 61.2 71.25 64.2 ;
        RECT  60.45 61.2 70.05 62.1 ;
        RECT  65.55 65.4 73.35 66.6 ;
        RECT  62.25 64.5 63.45 67.5 ;
        RECT  59.25 61.2 60.45 62.4 ;
        RECT  60.15 64.5 61.35 65.7 ;
        RECT  58.65 64.8 60.15 65.7 ;
        RECT  57.75 63.3 58.65 65.7 ;
        RECT  51.45 63.3 57.75 64.2 ;
        RECT  56.85 66.6 62.25 67.5 ;
        RECT  55.65 65.4 56.85 67.5 ;
        RECT  53.25 65.4 54.45 67.5 ;
        RECT  50.25 63.0 51.45 64.2 ;
        RECT  45.75 60.9 46.95 62.4 ;
        RECT  34.05 60.9 45.75 61.8 ;
        RECT  43.65 63.9 48.15 65.1 ;
        RECT  42.75 62.7 43.65 65.1 ;
        RECT  35.85 62.7 42.75 63.6 ;
        RECT  41.25 66.6 53.25 67.5 ;
        RECT  40.05 65.4 41.25 67.5 ;
        RECT  36.75 64.5 37.95 67.5 ;
        RECT  34.95 62.7 35.85 64.2 ;
        RECT  32.85 60.9 34.05 62.4 ;
        RECT  33.75 63.3 34.95 65.7 ;
        RECT  25.05 63.3 33.75 64.2 ;
        RECT  30.45 66.6 36.75 67.5 ;
        RECT  29.25 65.4 30.45 67.5 ;
        RECT  26.85 65.4 28.05 67.5 ;
        RECT  23.85 63.0 25.05 64.2 ;
        RECT  18.15 66.6 26.85 67.5 ;
        RECT  16.95 63.9 18.15 67.5 ;
        RECT  15.75 63.9 16.95 65.1 ;
        RECT  15.75 69.0 75.75 70.2 ;
        RECT  71.25 56.4 75.75 57.6 ;
        RECT  74.55 53.7 75.75 54.9 ;
        RECT  73.35 52.2 74.55 54.9 ;
        RECT  70.05 54.6 71.25 57.6 ;
        RECT  60.45 56.7 70.05 57.6 ;
        RECT  65.55 52.2 73.35 53.4 ;
        RECT  62.25 51.3 63.45 54.3 ;
        RECT  59.25 56.4 60.45 57.6 ;
        RECT  60.15 53.1 61.35 54.3 ;
        RECT  58.65 53.1 60.15 54.0 ;
        RECT  57.75 53.1 58.65 55.5 ;
        RECT  51.45 54.6 57.75 55.5 ;
        RECT  56.85 51.3 62.25 52.2 ;
        RECT  55.65 51.3 56.85 53.4 ;
        RECT  53.25 51.3 54.45 53.4 ;
        RECT  50.25 54.6 51.45 55.8 ;
        RECT  45.75 56.4 46.95 57.9 ;
        RECT  34.05 57.0 45.75 57.9 ;
        RECT  43.65 53.7 48.15 54.9 ;
        RECT  42.75 53.7 43.65 56.1 ;
        RECT  35.85 55.2 42.75 56.1 ;
        RECT  41.25 51.3 53.25 52.2 ;
        RECT  40.05 51.3 41.25 53.4 ;
        RECT  36.75 51.3 37.95 54.3 ;
        RECT  34.95 54.6 35.85 56.1 ;
        RECT  32.85 56.4 34.05 57.9 ;
        RECT  33.75 53.1 34.95 55.5 ;
        RECT  25.05 54.6 33.75 55.5 ;
        RECT  30.45 51.3 36.75 52.2 ;
        RECT  29.25 51.3 30.45 53.4 ;
        RECT  26.85 51.3 28.05 53.4 ;
        RECT  23.85 54.6 25.05 55.8 ;
        RECT  18.15 51.3 26.85 52.2 ;
        RECT  16.95 51.3 18.15 54.9 ;
        RECT  15.75 53.7 16.95 54.9 ;
        RECT  15.75 48.6 75.75 49.8 ;
        RECT  71.25 40.8 75.75 42.0 ;
        RECT  74.55 43.5 75.75 44.7 ;
        RECT  73.35 43.5 74.55 46.2 ;
        RECT  70.05 40.8 71.25 43.8 ;
        RECT  60.45 40.8 70.05 41.7 ;
        RECT  65.55 45.0 73.35 46.2 ;
        RECT  62.25 44.1 63.45 47.1 ;
        RECT  59.25 40.8 60.45 42.0 ;
        RECT  60.15 44.1 61.35 45.3 ;
        RECT  58.65 44.4 60.15 45.3 ;
        RECT  57.75 42.9 58.65 45.3 ;
        RECT  51.45 42.9 57.75 43.8 ;
        RECT  56.85 46.2 62.25 47.1 ;
        RECT  55.65 45.0 56.85 47.1 ;
        RECT  53.25 45.0 54.45 47.1 ;
        RECT  50.25 42.6 51.45 43.8 ;
        RECT  45.75 40.5 46.95 42.0 ;
        RECT  34.05 40.5 45.75 41.4 ;
        RECT  43.65 43.5 48.15 44.7 ;
        RECT  42.75 42.3 43.65 44.7 ;
        RECT  35.85 42.3 42.75 43.2 ;
        RECT  41.25 46.2 53.25 47.1 ;
        RECT  40.05 45.0 41.25 47.1 ;
        RECT  36.75 44.1 37.95 47.1 ;
        RECT  34.95 42.3 35.85 43.8 ;
        RECT  32.85 40.5 34.05 42.0 ;
        RECT  33.75 42.9 34.95 45.3 ;
        RECT  25.05 42.9 33.75 43.8 ;
        RECT  30.45 46.2 36.75 47.1 ;
        RECT  29.25 45.0 30.45 47.1 ;
        RECT  26.85 45.0 28.05 47.1 ;
        RECT  23.85 42.6 25.05 43.8 ;
        RECT  18.15 46.2 26.85 47.1 ;
        RECT  16.95 43.5 18.15 47.1 ;
        RECT  15.75 43.5 16.95 44.7 ;
        RECT  15.75 48.6 75.75 49.8 ;
        RECT  124.5 6.0 125.7 7.2 ;
        RECT  134.7 6.0 135.9 7.2 ;
        RECT  129.0 0.3 130.2 1.5 ;
        RECT  139.2 0.3 140.4 1.5 ;
        RECT  91.05 88.8 92.25 90.0 ;
        RECT  91.35 73.5 92.55 74.7 ;
        RECT  72.45 73.5 73.65 74.7 ;
        RECT  88.35 104.7 89.55 105.9 ;
        RECT  88.65 64.8 89.85 66.0 ;
        RECT  72.45 64.8 73.65 66.0 ;
        RECT  85.65 147.6 86.85 148.8 ;
        RECT  85.95 53.1 87.15 54.3 ;
        RECT  72.45 53.1 73.65 54.3 ;
        RECT  82.95 163.5 84.15 164.7 ;
        RECT  83.25 44.4 84.45 45.6 ;
        RECT  72.45 44.4 73.65 45.6 ;
        RECT  114.45 33.3 115.65 34.5 ;
        RECT  109.05 28.65 110.25 29.85 ;
        RECT  111.75 26.25 112.95 27.45 ;
        RECT  114.45 446.4 115.65 447.6 ;
        RECT  117.15 97.95 118.35 99.15 ;
        RECT  119.85 196.05 121.05 197.25 ;
        RECT  16.95 76.5 18.15 77.7 ;
        RECT  16.65 76.8 17.85 78.0 ;
        RECT  106.65 83.1 107.85 84.3 ;
        RECT  106.35 456.6 107.55 457.8 ;
        RECT  95.55 437.1 97.95 438.3 ;
        RECT  134.25 437.1 135.45 438.3 ;
        RECT  144.45 437.1 145.65 438.3 ;
        RECT  123.15 437.1 124.35 438.3 ;
        RECT  102.15 8.1 104.55 9.3 ;
        RECT  133.95 8.1 135.15 9.3 ;
        RECT  133.95 8.1 135.15 9.3 ;
        RECT  88.2 229.05 89.4 230.25 ;
        RECT  88.2 258.45 89.4 259.65 ;
        RECT  88.2 287.85 89.4 289.05 ;
        RECT  88.2 317.25 89.4 318.45 ;
        RECT  88.2 346.65 89.4 347.85 ;
        RECT  88.2 376.05 89.4 377.25 ;
        RECT  88.2 405.45 89.4 406.65 ;
        RECT  88.2 434.85 89.4 436.05 ;
        RECT  95.55 140.55 97.95 141.75 ;
        RECT  95.55 199.35 97.95 200.55 ;
        RECT  75.45 69.15 76.65 70.35 ;
        RECT  95.55 69.15 97.95 70.35 ;
        RECT  75.45 69.15 76.65 70.35 ;
        RECT  95.55 69.15 97.95 70.35 ;
        RECT  75.45 48.75 76.65 49.95 ;
        RECT  95.55 48.75 97.95 49.95 ;
        RECT  75.45 48.75 76.65 49.95 ;
        RECT  95.55 48.75 97.95 49.95 ;
        RECT  -66.3 148.2 -7.5 149.1 ;
        RECT  -66.3 150.9 -7.5 151.8 ;
        RECT  -66.3 153.6 -7.5 154.5 ;
        RECT  -66.3 156.3 -7.5 157.2 ;
        RECT  -66.3 159.0 -7.5 159.9 ;
        RECT  -66.3 161.7 -7.5 162.6 ;
        RECT  -66.3 211.5 -7.5 212.4 ;
        RECT  -66.3 214.2 -7.5 215.1 ;
        RECT  -66.3 216.9 -7.5 217.8 ;
        RECT  -66.3 219.6 -7.5 220.5 ;
        RECT  -15.6 121.05 -5.25 121.95 ;
        RECT  -7.5 150.9 -5.25 151.8 ;
        RECT  -7.5 214.2 -3.45 215.1 ;
        RECT  -56.55 145.5 -55.65 149.1 ;
        RECT  -56.55 145.5 -55.65 149.1 ;
        RECT  -36.15 145.5 -35.25 149.1 ;
        RECT  -27.15 126.45 -14.25 127.35 ;
        RECT  -7.5 161.7 -3.0 162.6 ;
        RECT  -14.1 88.5 -3.0 89.4 ;
        RECT  -14.7 175.5 -3.0 176.4 ;
        RECT  -7.5 211.5 -3.0 212.4 ;
        RECT  -14.7 180.0 -3.0 180.9 ;
        RECT  -64.5 141.0 -63.3 145.5 ;
        RECT  -61.8 144.3 -60.6 145.5 ;
        RECT  -61.8 143.1 -59.1 144.3 ;
        RECT  -64.5 139.8 -61.5 141.0 ;
        RECT  -64.5 130.2 -63.6 139.8 ;
        RECT  -60.3 135.3 -59.1 143.1 ;
        RECT  -61.2 132.0 -58.2 133.2 ;
        RECT  -64.5 129.0 -63.3 130.2 ;
        RECT  -61.2 129.9 -60.0 131.1 ;
        RECT  -60.9 128.4 -60.0 129.9 ;
        RECT  -62.4 127.5 -60.0 128.4 ;
        RECT  -62.4 121.2 -61.5 127.5 ;
        RECT  -59.1 126.6 -58.2 132.0 ;
        RECT  -60.3 125.4 -58.2 126.6 ;
        RECT  -60.3 123.0 -58.2 124.2 ;
        RECT  -62.7 120.0 -61.5 121.2 ;
        RECT  -64.8 115.5 -63.3 116.7 ;
        RECT  -64.8 103.8 -63.9 115.5 ;
        RECT  -61.8 113.4 -60.6 117.9 ;
        RECT  -63.0 112.5 -60.6 113.4 ;
        RECT  -63.0 105.6 -62.1 112.5 ;
        RECT  -59.1 111.0 -58.2 123.0 ;
        RECT  -60.3 109.8 -58.2 111.0 ;
        RECT  -61.2 106.5 -58.2 107.7 ;
        RECT  -63.0 104.7 -61.5 105.6 ;
        RECT  -64.8 102.6 -63.3 103.8 ;
        RECT  -62.4 103.5 -60.0 104.7 ;
        RECT  -62.4 94.8 -61.5 103.5 ;
        RECT  -59.1 100.2 -58.2 106.5 ;
        RECT  -60.3 99.0 -58.2 100.2 ;
        RECT  -60.3 96.6 -58.2 97.8 ;
        RECT  -62.7 93.6 -61.5 94.8 ;
        RECT  -59.1 87.9 -58.2 96.6 ;
        RECT  -61.8 86.7 -58.2 87.9 ;
        RECT  -61.8 85.5 -60.6 86.7 ;
        RECT  -56.7 85.5 -55.5 145.5 ;
        RECT  -48.9 141.0 -47.7 145.5 ;
        RECT  -51.6 144.3 -50.4 145.5 ;
        RECT  -53.1 143.1 -50.4 144.3 ;
        RECT  -50.7 139.8 -47.7 141.0 ;
        RECT  -48.6 130.2 -47.7 139.8 ;
        RECT  -53.1 135.3 -51.9 143.1 ;
        RECT  -54.0 132.0 -51.0 133.2 ;
        RECT  -48.9 129.0 -47.7 130.2 ;
        RECT  -52.2 129.9 -51.0 131.1 ;
        RECT  -52.2 128.4 -51.3 129.9 ;
        RECT  -52.2 127.5 -49.8 128.4 ;
        RECT  -50.7 121.2 -49.8 127.5 ;
        RECT  -54.0 126.6 -53.1 132.0 ;
        RECT  -54.0 125.4 -51.9 126.6 ;
        RECT  -54.0 123.0 -51.9 124.2 ;
        RECT  -50.7 120.0 -49.5 121.2 ;
        RECT  -48.9 115.5 -47.4 116.7 ;
        RECT  -48.3 103.8 -47.4 115.5 ;
        RECT  -51.6 113.4 -50.4 117.9 ;
        RECT  -51.6 112.5 -49.2 113.4 ;
        RECT  -50.1 105.6 -49.2 112.5 ;
        RECT  -54.0 111.0 -53.1 123.0 ;
        RECT  -54.0 109.8 -51.9 111.0 ;
        RECT  -54.0 106.5 -51.0 107.7 ;
        RECT  -50.7 104.7 -49.2 105.6 ;
        RECT  -48.9 102.6 -47.4 103.8 ;
        RECT  -52.2 103.5 -49.8 104.7 ;
        RECT  -50.7 94.8 -49.8 103.5 ;
        RECT  -54.0 100.2 -53.1 106.5 ;
        RECT  -54.0 99.0 -51.9 100.2 ;
        RECT  -54.0 96.6 -51.9 97.8 ;
        RECT  -50.7 93.6 -49.5 94.8 ;
        RECT  -54.0 87.9 -53.1 96.6 ;
        RECT  -54.0 86.7 -50.4 87.9 ;
        RECT  -51.6 85.5 -50.4 86.7 ;
        RECT  -56.7 85.5 -55.5 145.5 ;
        RECT  -44.1 141.0 -42.9 145.5 ;
        RECT  -41.4 144.3 -40.2 145.5 ;
        RECT  -41.4 143.1 -38.7 144.3 ;
        RECT  -44.1 139.8 -41.1 141.0 ;
        RECT  -44.1 130.2 -43.2 139.8 ;
        RECT  -39.9 135.3 -38.7 143.1 ;
        RECT  -40.8 132.0 -37.8 133.2 ;
        RECT  -44.1 129.0 -42.9 130.2 ;
        RECT  -40.8 129.9 -39.6 131.1 ;
        RECT  -40.5 128.4 -39.6 129.9 ;
        RECT  -42.0 127.5 -39.6 128.4 ;
        RECT  -42.0 121.2 -41.1 127.5 ;
        RECT  -38.7 126.6 -37.8 132.0 ;
        RECT  -39.9 125.4 -37.8 126.6 ;
        RECT  -39.9 123.0 -37.8 124.2 ;
        RECT  -42.3 120.0 -41.1 121.2 ;
        RECT  -44.4 115.5 -42.9 116.7 ;
        RECT  -44.4 103.8 -43.5 115.5 ;
        RECT  -41.4 113.4 -40.2 117.9 ;
        RECT  -42.6 112.5 -40.2 113.4 ;
        RECT  -42.6 105.6 -41.7 112.5 ;
        RECT  -38.7 111.0 -37.8 123.0 ;
        RECT  -39.9 109.8 -37.8 111.0 ;
        RECT  -40.8 106.5 -37.8 107.7 ;
        RECT  -42.6 104.7 -41.1 105.6 ;
        RECT  -44.4 102.6 -42.9 103.8 ;
        RECT  -42.0 103.5 -39.6 104.7 ;
        RECT  -42.0 94.8 -41.1 103.5 ;
        RECT  -38.7 100.2 -37.8 106.5 ;
        RECT  -39.9 99.0 -37.8 100.2 ;
        RECT  -39.9 96.6 -37.8 97.8 ;
        RECT  -42.3 93.6 -41.1 94.8 ;
        RECT  -38.7 87.9 -37.8 96.6 ;
        RECT  -41.4 86.7 -37.8 87.9 ;
        RECT  -41.4 85.5 -40.2 86.7 ;
        RECT  -36.3 85.5 -35.1 145.5 ;
        RECT  -19.65 100.05 -13.65 100.95 ;
        RECT  -19.65 95.25 -13.65 96.15 ;
        RECT  -19.65 99.9 -18.45 101.1 ;
        RECT  -13.05 99.9 -11.85 101.1 ;
        RECT  -19.65 95.1 -18.45 96.3 ;
        RECT  -13.05 95.1 -11.85 96.3 ;
        RECT  -43.65 236.7 -41.85 238.5 ;
        RECT  -44.55 234.6 -32.25 235.5 ;
        RECT  -55.8 237.15 -54.9 254.7 ;
        RECT  -13.65 241.95 -12.75 262.2 ;
        RECT  -32.1 262.2 -31.2 271.8 ;
        RECT  -13.65 230.55 -12.75 231.45 ;
        RECT  -50.1 230.55 -49.2 231.45 ;
        RECT  -13.65 231.0 -12.75 241.95 ;
        RECT  -44.55 230.55 -13.2 231.45 ;
        RECT  -49.65 230.55 -44.55 231.45 ;
        RECT  -50.1 231.0 -49.2 252.0 ;
        RECT  -45.9 245.7 -45.0 293.25 ;
        RECT  -45.9 265.8 -45.0 293.25 ;
        RECT  -8.4 231.0 -7.5 288.6 ;
        RECT  -37.8 267.6 -36.9 288.6 ;
        RECT  -43.2 257.4 -42.3 268.05 ;
        RECT  -45.9 268.8 -45.0 293.25 ;
        RECT  -43.2 268.05 -42.3 281.4 ;
        RECT  -45.9 240.6 -45.0 293.25 ;
        RECT  -62.4 231.0 -61.5 284.1 ;
        RECT  -52.2 231.0 -51.3 284.1 ;
        RECT  -14.55 258.0 -13.65 262.2 ;
        RECT  -14.55 248.85 -13.65 252.6 ;
        RECT  -31.65 248.4 -30.75 248.85 ;
        RECT  -31.65 253.8 -30.75 258.0 ;
        RECT  -14.85 266.4 -13.65 267.6 ;
        RECT  -14.85 256.8 -13.65 258.0 ;
        RECT  -31.65 248.4 -30.45 249.6 ;
        RECT  -31.65 258.0 -30.45 259.2 ;
        RECT  -14.85 261.0 -13.65 262.2 ;
        RECT  -14.85 251.4 -13.65 252.6 ;
        RECT  -14.7 248.25 -13.5 249.45 ;
        RECT  -31.8 248.25 -30.6 249.45 ;
        RECT  -31.65 253.8 -30.45 255.0 ;
        RECT  -53.55 258.9 -51.75 269.4 ;
        RECT  -55.95 255.9 -54.75 269.4 ;
        RECT  -58.95 255.9 -57.75 269.4 ;
        RECT  -55.95 254.7 -53.25 255.9 ;
        RECT  -58.95 254.7 -57.45 255.9 ;
        RECT  -62.55 254.7 -61.35 269.4 ;
        RECT  -53.55 240.0 -51.15 250.5 ;
        RECT  -55.95 240.0 -54.75 253.5 ;
        RECT  -58.95 240.0 -57.75 253.5 ;
        RECT  -55.95 253.5 -53.25 254.7 ;
        RECT  -58.95 253.5 -57.45 254.7 ;
        RECT  -62.55 240.0 -61.35 254.7 ;
        RECT  -53.55 229.5 -51.15 240.0 ;
        RECT  -55.95 226.5 -54.75 240.0 ;
        RECT  -58.95 226.5 -57.75 240.0 ;
        RECT  -55.95 225.3 -53.25 226.5 ;
        RECT  -58.95 225.3 -57.45 226.5 ;
        RECT  -62.55 225.3 -61.35 240.0 ;
        RECT  -43.05 235.95 -41.85 237.15 ;
        RECT  -32.85 233.25 -31.65 234.45 ;
        RECT  -45.15 233.25 -43.95 234.45 ;
        RECT  -55.95 235.35 -54.75 236.55 ;
        RECT  -13.8 260.4 -12.6 261.6 ;
        RECT  -32.25 260.4 -31.05 261.6 ;
        RECT  -32.85 271.8 -31.65 273.0 ;
        RECT  -13.8 240.15 -12.6 241.35 ;
        RECT  -50.25 250.2 -49.05 251.4 ;
        RECT  -46.05 243.9 -44.85 245.1 ;
        RECT  -46.05 264.0 -44.85 265.2 ;
        RECT  -8.55 229.2 -7.35 230.4 ;
        RECT  -8.55 286.8 -7.35 288.0 ;
        RECT  -37.95 286.8 -36.75 288.0 ;
        RECT  -46.65 293.25 -45.45 294.45 ;
        RECT  -43.35 266.25 -42.15 267.45 ;
        RECT  -43.35 255.6 -42.15 256.8 ;
        RECT  -46.05 267.0 -44.85 268.2 ;
        RECT  -43.35 266.25 -42.15 267.45 ;
        RECT  -43.35 279.6 -42.15 280.8 ;
        RECT  -46.05 238.8 -44.85 240.0 ;
        RECT  -62.55 229.2 -61.35 230.4 ;
        RECT  -52.35 229.2 -51.15 230.4 ;
        RECT  -25.05 169.8 -23.85 175.8 ;
        RECT  -32.7 165.6 -31.8 171.9 ;
        RECT  -34.5 165.6 -33.6 174.3 ;
        RECT  -33.6 173.1 -31.8 174.3 ;
        RECT  -26.25 169.8 -25.05 171.0 ;
        RECT  -26.25 174.6 -25.05 175.8 ;
        RECT  -33.0 170.7 -31.8 171.9 ;
        RECT  -33.9 165.3 -32.7 166.5 ;
        RECT  -33.0 173.1 -31.8 174.3 ;
        RECT  -36.0 165.3 -34.8 166.5 ;
        RECT  -49.95 169.8 -48.75 175.8 ;
        RECT  -42.0 165.6 -41.1 171.9 ;
        RECT  -40.2 165.6 -39.3 174.3 ;
        RECT  -42.0 173.1 -40.2 174.3 ;
        RECT  -49.95 169.8 -48.75 171.0 ;
        RECT  -49.95 174.6 -48.75 175.8 ;
        RECT  -43.2 170.7 -42.0 171.9 ;
        RECT  -42.3 165.3 -41.1 166.5 ;
        RECT  -43.2 173.1 -42.0 174.3 ;
        RECT  -40.2 165.3 -39.0 166.5 ;
        RECT  -40.8 144.3 -39.6 145.5 ;
        RECT  -40.8 150.9 -39.6 152.1 ;
        RECT  -44.25 144.3 -43.05 145.5 ;
        RECT  -44.25 153.6 -43.05 154.8 ;
        RECT  -64.65 144.3 -63.45 145.5 ;
        RECT  -64.65 156.3 -63.45 157.5 ;
        RECT  -49.05 144.3 -47.85 145.5 ;
        RECT  -49.05 159.0 -47.85 160.2 ;
        RECT  -17.4 153.6 -16.2 154.8 ;
        RECT  -14.1 161.7 -12.9 162.9 ;
        RECT  -27.45 161.7 -26.25 162.9 ;
        RECT  -33.0 153.6 -31.8 154.8 ;
        RECT  -34.8 156.3 -33.6 157.5 ;
        RECT  -47.85 161.7 -46.65 162.9 ;
        RECT  -42.3 159.0 -41.1 160.2 ;
        RECT  -40.5 156.3 -39.3 157.5 ;
        RECT  -16.2 120.9 -15.0 122.1 ;
        RECT  -5.85 120.9 -4.65 122.1 ;
        RECT  -5.85 150.75 -4.65 151.95 ;
        RECT  -30.9 214.2 -29.7 215.4 ;
        RECT  -44.4 211.5 -43.2 212.7 ;
        RECT  -15.0 216.9 -13.8 218.1 ;
        RECT  -4.05 214.05 -2.85 215.25 ;
        RECT  -43.35 217.2 -42.15 218.4 ;
        RECT  -43.35 237.0 -42.15 238.2 ;
        RECT  -22.95 219.6 -21.75 220.8 ;
        RECT  -52.35 219.6 -51.15 220.8 ;
        RECT  -8.25 148.2 -7.05 149.4 ;
        RECT  -14.85 126.3 -13.65 127.5 ;
        RECT  -27.75 126.3 -26.55 127.5 ;
        RECT  -27.6 85.5 -26.4 86.7 ;
        RECT  -27.3 85.8 -26.1 87.0 ;
        RECT  -4.5 162.0 -3.3 163.2 ;
        RECT  -14.1 88.5 -12.9 89.7 ;
        RECT  -4.5 88.8 -3.3 90.0 ;
        RECT  -15.0 175.5 -13.8 176.7 ;
        RECT  -4.5 175.8 -3.3 177.0 ;
        RECT  -4.5 211.8 -3.3 213.0 ;
        RECT  -15.0 180.0 -13.8 181.2 ;
        RECT  -4.5 180.3 -3.3 181.5 ;
        RECT  105.75 85.8 106.95 87.0 ;
        RECT  113.85 162.0 115.05 163.2 ;
        RECT  111.15 88.8 112.35 90.0 ;
        RECT  108.45 175.8 109.65 177.0 ;
        RECT  116.55 211.8 117.75 213.0 ;
        RECT  119.25 180.3 120.45 181.5 ;
        RECT  0.45 219.6 2.85 220.8 ;
        RECT  95.85 230.7 98.55 231.9 ;
        RECT  -8.1 230.7 -6.9 231.9 ;
        Layer  via2 ; 
        RECT  125.55 152.7 126.15 153.3 ;
        RECT  135.75 152.7 136.35 153.3 ;
        RECT  129.15 32.4 129.75 33.0 ;
        RECT  139.35 32.4 139.95 33.0 ;
        RECT  129.15 32.7 129.75 33.3 ;
        RECT  139.35 32.7 139.95 33.3 ;
        RECT  17.25 74.4 17.85 75.0 ;
        RECT  17.25 64.2 17.85 64.8 ;
        RECT  17.25 54.0 17.85 54.6 ;
        RECT  17.25 43.8 17.85 44.4 ;
        RECT  124.8 6.3 125.4 6.9 ;
        RECT  135.0 6.3 135.6 6.9 ;
        RECT  129.3 0.6 129.9 1.2 ;
        RECT  139.5 0.6 140.1 1.2 ;
        RECT  91.65 73.8 92.25 74.4 ;
        RECT  72.75 73.8 73.35 74.4 ;
        RECT  88.95 65.1 89.55 65.7 ;
        RECT  72.75 65.1 73.35 65.7 ;
        RECT  86.25 53.4 86.85 54.0 ;
        RECT  72.75 53.4 73.35 54.0 ;
        RECT  83.55 44.7 84.15 45.3 ;
        RECT  72.75 44.7 73.35 45.3 ;
        RECT  16.95 77.1 17.55 77.7 ;
        RECT  106.95 83.4 107.55 84.0 ;
        RECT  -61.5 87.0 -60.9 87.6 ;
        RECT  -51.3 87.0 -50.7 87.6 ;
        RECT  -41.1 87.0 -40.5 87.6 ;
        RECT  -14.4 248.55 -13.8 249.15 ;
        RECT  -31.5 248.55 -30.9 249.15 ;
        RECT  -43.05 217.5 -42.45 218.1 ;
        RECT  -43.05 237.3 -42.45 237.9 ;
        RECT  -27.0 86.1 -26.4 86.7 ;
        RECT  -4.2 162.3 -3.6 162.9 ;
        RECT  -4.2 89.1 -3.6 89.7 ;
        RECT  -4.2 176.1 -3.6 176.7 ;
        RECT  -4.2 212.1 -3.6 212.7 ;
        RECT  -4.2 180.6 -3.6 181.2 ;
        RECT  106.05 86.1 106.65 86.7 ;
        RECT  114.15 162.3 114.75 162.9 ;
        RECT  111.45 89.1 112.05 89.7 ;
        RECT  108.75 176.1 109.35 176.7 ;
        RECT  116.85 212.1 117.45 212.7 ;
        RECT  119.55 180.6 120.15 181.2 ;
        RECT  96.15 231.0 96.75 231.6 ;
        RECT  97.65 231.0 98.25 231.6 ;
        RECT  -7.8 231.0 -7.2 231.6 ;
        Layer  metal3 ; 
        RECT  -27.15 85.5 106.35 87.0 ;
        RECT  -3.0 161.7 114.45 163.2 ;
        RECT  -3.0 88.5 111.75 90.0 ;
        RECT  -3.0 175.5 109.05 177.0 ;
        RECT  -3.0 211.5 117.15 213.0 ;
        RECT  -3.0 180.0 119.85 181.5 ;
        RECT  -6.6 230.4 95.55 231.9 ;
        RECT  124.2 153.75 125.7 155.25 ;
        RECT  124.2 6.45 125.7 154.5 ;
        RECT  124.95 153.75 126.6 155.25 ;
        RECT  134.4 153.75 135.9 155.25 ;
        RECT  134.4 6.45 135.9 154.5 ;
        RECT  135.15 153.75 136.8 155.25 ;
        RECT  128.7 0.0 130.2 30.15 ;
        RECT  138.9 0.0 140.4 30.15 ;
        RECT  73.95 73.2 91.95 74.7 ;
        RECT  73.95 64.5 89.25 66.0 ;
        RECT  73.95 52.8 86.55 54.3 ;
        RECT  73.95 44.1 83.85 45.6 ;
        RECT  0.45 73.95 17.55 75.45 ;
        RECT  0.45 63.75 17.55 65.25 ;
        RECT  0.45 53.55 17.55 55.05 ;
        RECT  0.45 43.35 17.55 44.85 ;
        RECT  17.4 82.8 18.9 84.3 ;
        RECT  17.4 76.5 18.9 83.55 ;
        RECT  18.15 82.8 106.65 84.3 ;
        RECT  124.95 152.1 126.75 153.9 ;
        RECT  135.15 152.1 136.95 153.9 ;
        RECT  128.55 31.8 130.35 33.6 ;
        RECT  138.75 31.8 140.55 33.6 ;
        RECT  128.55 32.1 130.35 33.9 ;
        RECT  138.75 32.1 140.55 33.9 ;
        RECT  16.65 73.8 18.45 75.6 ;
        RECT  16.65 63.6 18.45 65.4 ;
        RECT  16.65 53.4 18.45 55.2 ;
        RECT  16.65 43.2 18.45 45.0 ;
        RECT  124.2 5.7 126.0 7.5 ;
        RECT  134.4 5.7 136.2 7.5 ;
        RECT  128.7 0.0 130.5 1.8 ;
        RECT  138.9 0.0 140.7 1.8 ;
        RECT  91.05 73.2 92.85 75.0 ;
        RECT  72.15 73.2 73.95 75.0 ;
        RECT  88.35 64.5 90.15 66.3 ;
        RECT  72.15 64.5 73.95 66.3 ;
        RECT  85.65 52.8 87.45 54.6 ;
        RECT  72.15 52.8 73.95 54.6 ;
        RECT  82.95 44.1 84.75 45.9 ;
        RECT  72.15 44.1 73.95 45.9 ;
        RECT  16.35 76.5 18.15 78.3 ;
        RECT  106.35 82.8 108.15 84.6 ;
        RECT  -43.35 216.9 -41.85 237.15 ;
        RECT  -62.1 86.4 -60.3 88.2 ;
        RECT  -51.9 86.4 -50.1 88.2 ;
        RECT  -41.7 86.4 -39.9 88.2 ;
        RECT  -31.2 248.1 -14.1 249.6 ;
        RECT  -15.0 247.95 -13.2 249.75 ;
        RECT  -32.1 247.95 -30.3 249.75 ;
        RECT  -43.65 216.9 -41.85 218.7 ;
        RECT  -43.65 236.7 -41.85 238.5 ;
        RECT  -27.6 85.5 -25.8 87.3 ;
        RECT  -4.8 161.7 -3.0 163.5 ;
        RECT  -4.8 88.5 -3.0 90.3 ;
        RECT  -4.8 175.5 -3.0 177.3 ;
        RECT  -4.8 211.5 -3.0 213.3 ;
        RECT  -4.8 180.0 -3.0 181.8 ;
        RECT  105.45 85.5 107.25 87.3 ;
        RECT  113.55 161.7 115.35 163.5 ;
        RECT  110.85 88.5 112.65 90.3 ;
        RECT  108.15 175.5 109.95 177.3 ;
        RECT  116.25 211.5 118.05 213.3 ;
        RECT  118.95 180.0 120.75 181.8 ;
        RECT  95.55 230.4 98.85 232.2 ;
        RECT  -8.4 230.4 -6.6 232.2 ;
    END 
END    sram_2_16_1_scn3me_subm 
END    LIBRARY 
