MACRO sram_2_16_1_freepdk45
    CLASS RING ;
    ORIGIN 4.22 0.0 ;
    FOREIGN  sram 0.0 0.0 ;
    SIZE 16.475 BY 42.02 ;
    SYMMETRY X Y R90 ;
    PIN vdd
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  11.95 0.0 12.3 42.02 ;
        RECT  11.95 0.0 12.3 42.02 ;
        RECT  0.0 0.0 0.35 42.02 ;
        RECT  0.0 0.0 0.35 42.02 ;
        END
    END vdd
    PIN gnd
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal2 ;
        RECT  8.2525 0.0 8.6025 42.02 ;
        RECT  8.2525 0.0 8.6025 42.02 ;
        END
    END gnd
    PIN DATA[0]
        DIRECTION INOUT ;
        PORT
        LAYER metal2 ;
        RECT  10.6625 0.0 10.7325 0.14 ;
        RECT  10.6625 0.0 10.7325 0.14 ;
        RECT  10.6625 0.0 10.7325 0.135 ;
        END
    END DATA[0]
    PIN DATA[1]
        DIRECTION INOUT ;
        PORT
        LAYER metal2 ;
        RECT  11.3675 0.0 11.4375 0.14 ;
        RECT  11.3675 0.0 11.4375 0.14 ;
        RECT  11.3675 0.0 11.4375 0.135 ;
        END
    END DATA[1]
    PIN ADDR[0]
        DIRECTION INPUT ;
        PORT
        LAYER metal3 ;
        RECT  0.0 7.5325 0.48 7.6025 ;
        RECT  0.0 7.5325 0.48 7.6025 ;
        END
    END ADDR[0]
    PIN ADDR[1]
        DIRECTION INPUT ;
        PORT
        LAYER metal3 ;
        RECT  0.0 6.8275 0.48 6.8975 ;
        RECT  0.0 6.8275 0.48 6.8975 ;
        END
    END ADDR[1]
    PIN ADDR[2]
        DIRECTION INPUT ;
        PORT
        LAYER metal3 ;
        RECT  0.0 6.1225 0.48 6.1925 ;
        RECT  0.0 6.1225 0.48 6.1925 ;
        END
    END ADDR[2]
    PIN ADDR[3]
        DIRECTION INPUT ;
        PORT
        LAYER metal3 ;
        RECT  0.0 5.4175 0.48 5.4875 ;
        RECT  0.0 5.4175 0.48 5.4875 ;
        END
    END ADDR[3]
    PIN CSb
        DIRECTION INPUT ;
        PORT
        LAYER metal3 ;
        RECT  -2.9875 19.23 -2.9175 19.37 ;
        RECT  -2.9875 19.23 -2.9175 19.37 ;
        RECT  -2.9875 19.23 -2.9175 19.37 ;
        RECT  -2.9875 19.23 -2.9175 19.37 ;
        RECT  -2.9875 19.23 -2.9175 19.37 ;
        END
    END CSb
    PIN OEb
        DIRECTION INPUT ;
        PORT
        LAYER metal3 ;
        RECT  -3.6925 19.23 -3.6225 19.37 ;
        RECT  -3.6925 19.23 -3.6225 19.37 ;
        RECT  -3.6925 19.23 -3.6225 19.37 ;
        RECT  -3.6925 19.23 -3.6225 19.37 ;
        RECT  -3.6925 19.23 -3.6225 19.37 ;
        END
    END OEb
    PIN WEb
        DIRECTION INPUT ;
        PORT
        LAYER metal3 ;
        RECT  -2.2825 19.23 -2.2125 19.37 ;
        RECT  -2.2825 19.23 -2.2125 19.37 ;
        RECT  -2.2825 19.23 -2.2125 19.37 ;
        RECT  -2.2825 19.23 -2.2125 19.37 ;
        RECT  -2.2825 19.23 -2.2125 19.37 ;
        END
    END WEb
    PIN clk
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  -0.755 19.23 -0.69 19.295 ;
        RECT  -0.755 19.23 -0.69 19.295 ;
        RECT  -0.755 19.23 -0.69 19.265 ;
        END
    END clk
    OBS
        LAYER  metal1 ;
        RECT  0.1425 27.47 0.2075 27.675 ;
        RECT  -0.755 19.23 -0.69 19.295 ;
        RECT  11.95 0.0 12.3 42.02 ;
        RECT  0.0 0.0 0.35 42.02 ;
        RECT  4.435 19.64 4.5 19.705 ;
        RECT  4.435 20.0 4.5 20.065 ;
        RECT  4.1975 19.64 4.4675 19.705 ;
        RECT  4.435 19.6725 4.5 20.0325 ;
        RECT  4.4675 20.0 4.805 20.065 ;
        RECT  6.9325 19.64 6.9975 19.705 ;
        RECT  6.9325 19.1975 6.9975 19.2625 ;
        RECT  6.76 19.64 6.965 19.705 ;
        RECT  6.9325 19.23 6.9975 19.6725 ;
        RECT  6.965 19.1975 10.255 19.2625 ;
        RECT  4.435 21.165 4.5 21.23 ;
        RECT  4.435 20.805 4.5 20.87 ;
        RECT  4.1975 21.165 4.4675 21.23 ;
        RECT  4.435 20.8375 4.5 21.1975 ;
        RECT  4.4675 20.805 4.805 20.87 ;
        RECT  6.9325 21.165 6.9975 21.23 ;
        RECT  6.9325 21.6075 6.9975 21.6725 ;
        RECT  6.76 21.165 6.965 21.23 ;
        RECT  6.9325 21.1975 6.9975 21.64 ;
        RECT  6.965 21.6075 10.255 21.6725 ;
        RECT  4.435 22.33 4.5 22.395 ;
        RECT  4.435 22.69 4.5 22.755 ;
        RECT  4.1975 22.33 4.4675 22.395 ;
        RECT  4.435 22.3625 4.5 22.7225 ;
        RECT  4.4675 22.69 4.805 22.755 ;
        RECT  6.9325 22.33 6.9975 22.395 ;
        RECT  6.9325 21.8875 6.9975 21.9525 ;
        RECT  6.76 22.33 6.965 22.395 ;
        RECT  6.9325 21.92 6.9975 22.3625 ;
        RECT  6.965 21.8875 10.255 21.9525 ;
        RECT  4.435 23.855 4.5 23.92 ;
        RECT  4.435 23.495 4.5 23.56 ;
        RECT  4.1975 23.855 4.4675 23.92 ;
        RECT  4.435 23.5275 4.5 23.8875 ;
        RECT  4.4675 23.495 4.805 23.56 ;
        RECT  6.9325 23.855 6.9975 23.92 ;
        RECT  6.9325 24.2975 6.9975 24.3625 ;
        RECT  6.76 23.855 6.965 23.92 ;
        RECT  6.9325 23.8875 6.9975 24.33 ;
        RECT  6.965 24.2975 10.255 24.3625 ;
        RECT  4.435 25.02 4.5 25.085 ;
        RECT  4.435 25.38 4.5 25.445 ;
        RECT  4.1975 25.02 4.4675 25.085 ;
        RECT  4.435 25.0525 4.5 25.4125 ;
        RECT  4.4675 25.38 4.805 25.445 ;
        RECT  6.9325 25.02 6.9975 25.085 ;
        RECT  6.9325 24.5775 6.9975 24.6425 ;
        RECT  6.76 25.02 6.965 25.085 ;
        RECT  6.9325 24.61 6.9975 25.0525 ;
        RECT  6.965 24.5775 10.255 24.6425 ;
        RECT  4.435 26.545 4.5 26.61 ;
        RECT  4.435 26.185 4.5 26.25 ;
        RECT  4.1975 26.545 4.4675 26.61 ;
        RECT  4.435 26.2175 4.5 26.5775 ;
        RECT  4.4675 26.185 4.805 26.25 ;
        RECT  6.9325 26.545 6.9975 26.61 ;
        RECT  6.9325 26.9875 6.9975 27.0525 ;
        RECT  6.76 26.545 6.965 26.61 ;
        RECT  6.9325 26.5775 6.9975 27.02 ;
        RECT  6.965 26.9875 10.255 27.0525 ;
        RECT  4.435 27.71 4.5 27.775 ;
        RECT  4.435 28.07 4.5 28.135 ;
        RECT  4.1975 27.71 4.4675 27.775 ;
        RECT  4.435 27.7425 4.5 28.1025 ;
        RECT  4.4675 28.07 4.805 28.135 ;
        RECT  6.9325 27.71 6.9975 27.775 ;
        RECT  6.9325 27.2675 6.9975 27.3325 ;
        RECT  6.76 27.71 6.965 27.775 ;
        RECT  6.9325 27.3 6.9975 27.7425 ;
        RECT  6.965 27.2675 10.255 27.3325 ;
        RECT  4.435 29.235 4.5 29.3 ;
        RECT  4.435 28.875 4.5 28.94 ;
        RECT  4.1975 29.235 4.4675 29.3 ;
        RECT  4.435 28.9075 4.5 29.2675 ;
        RECT  4.4675 28.875 4.805 28.94 ;
        RECT  6.9325 29.235 6.9975 29.3 ;
        RECT  6.9325 29.6775 6.9975 29.7425 ;
        RECT  6.76 29.235 6.965 29.3 ;
        RECT  6.9325 29.2675 6.9975 29.71 ;
        RECT  6.965 29.6775 10.255 29.7425 ;
        RECT  4.435 30.4 4.5 30.465 ;
        RECT  4.435 30.76 4.5 30.825 ;
        RECT  4.1975 30.4 4.4675 30.465 ;
        RECT  4.435 30.4325 4.5 30.7925 ;
        RECT  4.4675 30.76 4.805 30.825 ;
        RECT  6.9325 30.4 6.9975 30.465 ;
        RECT  6.9325 29.9575 6.9975 30.0225 ;
        RECT  6.76 30.4 6.965 30.465 ;
        RECT  6.9325 29.99 6.9975 30.4325 ;
        RECT  6.965 29.9575 10.255 30.0225 ;
        RECT  4.435 31.925 4.5 31.99 ;
        RECT  4.435 31.565 4.5 31.63 ;
        RECT  4.1975 31.925 4.4675 31.99 ;
        RECT  4.435 31.5975 4.5 31.9575 ;
        RECT  4.4675 31.565 4.805 31.63 ;
        RECT  6.9325 31.925 6.9975 31.99 ;
        RECT  6.9325 32.3675 6.9975 32.4325 ;
        RECT  6.76 31.925 6.965 31.99 ;
        RECT  6.9325 31.9575 6.9975 32.4 ;
        RECT  6.965 32.3675 10.255 32.4325 ;
        RECT  4.435 33.09 4.5 33.155 ;
        RECT  4.435 33.45 4.5 33.515 ;
        RECT  4.1975 33.09 4.4675 33.155 ;
        RECT  4.435 33.1225 4.5 33.4825 ;
        RECT  4.4675 33.45 4.805 33.515 ;
        RECT  6.9325 33.09 6.9975 33.155 ;
        RECT  6.9325 32.6475 6.9975 32.7125 ;
        RECT  6.76 33.09 6.965 33.155 ;
        RECT  6.9325 32.68 6.9975 33.1225 ;
        RECT  6.965 32.6475 10.255 32.7125 ;
        RECT  4.435 34.615 4.5 34.68 ;
        RECT  4.435 34.255 4.5 34.32 ;
        RECT  4.1975 34.615 4.4675 34.68 ;
        RECT  4.435 34.2875 4.5 34.6475 ;
        RECT  4.4675 34.255 4.805 34.32 ;
        RECT  6.9325 34.615 6.9975 34.68 ;
        RECT  6.9325 35.0575 6.9975 35.1225 ;
        RECT  6.76 34.615 6.965 34.68 ;
        RECT  6.9325 34.6475 6.9975 35.09 ;
        RECT  6.965 35.0575 10.255 35.1225 ;
        RECT  4.435 35.78 4.5 35.845 ;
        RECT  4.435 36.14 4.5 36.205 ;
        RECT  4.1975 35.78 4.4675 35.845 ;
        RECT  4.435 35.8125 4.5 36.1725 ;
        RECT  4.4675 36.14 4.805 36.205 ;
        RECT  6.9325 35.78 6.9975 35.845 ;
        RECT  6.9325 35.3375 6.9975 35.4025 ;
        RECT  6.76 35.78 6.965 35.845 ;
        RECT  6.9325 35.37 6.9975 35.8125 ;
        RECT  6.965 35.3375 10.255 35.4025 ;
        RECT  4.435 37.305 4.5 37.37 ;
        RECT  4.435 36.945 4.5 37.01 ;
        RECT  4.1975 37.305 4.4675 37.37 ;
        RECT  4.435 36.9775 4.5 37.3375 ;
        RECT  4.4675 36.945 4.805 37.01 ;
        RECT  6.9325 37.305 6.9975 37.37 ;
        RECT  6.9325 37.7475 6.9975 37.8125 ;
        RECT  6.76 37.305 6.965 37.37 ;
        RECT  6.9325 37.3375 6.9975 37.78 ;
        RECT  6.965 37.7475 10.255 37.8125 ;
        RECT  4.435 38.47 4.5 38.535 ;
        RECT  4.435 38.83 4.5 38.895 ;
        RECT  4.1975 38.47 4.4675 38.535 ;
        RECT  4.435 38.5025 4.5 38.8625 ;
        RECT  4.4675 38.83 4.805 38.895 ;
        RECT  6.9325 38.47 6.9975 38.535 ;
        RECT  6.9325 38.0275 6.9975 38.0925 ;
        RECT  6.76 38.47 6.965 38.535 ;
        RECT  6.9325 38.06 6.9975 38.5025 ;
        RECT  6.965 38.0275 10.255 38.0925 ;
        RECT  4.435 39.995 4.5 40.06 ;
        RECT  4.435 39.635 4.5 39.7 ;
        RECT  4.1975 39.995 4.4675 40.06 ;
        RECT  4.435 39.6675 4.5 40.0275 ;
        RECT  4.4675 39.635 4.805 39.7 ;
        RECT  6.9325 39.995 6.9975 40.06 ;
        RECT  6.9325 40.4375 6.9975 40.5025 ;
        RECT  6.76 39.995 6.965 40.06 ;
        RECT  6.9325 40.0275 6.9975 40.47 ;
        RECT  6.965 40.4375 10.255 40.5025 ;
        RECT  4.89 19.0575 10.345 19.1225 ;
        RECT  4.89 21.7475 10.345 21.8125 ;
        RECT  4.89 24.4375 10.345 24.5025 ;
        RECT  4.89 27.1275 10.345 27.1925 ;
        RECT  4.89 29.8175 10.345 29.8825 ;
        RECT  4.89 32.5075 10.345 32.5725 ;
        RECT  4.89 35.1975 10.345 35.2625 ;
        RECT  4.89 37.8875 10.345 37.9525 ;
        RECT  4.89 40.5775 10.345 40.6425 ;
        RECT  0.0 20.4025 12.3 20.4675 ;
        RECT  0.0 23.0925 12.3 23.1575 ;
        RECT  0.0 25.7825 12.3 25.8475 ;
        RECT  0.0 28.4725 12.3 28.5375 ;
        RECT  0.0 31.1625 12.3 31.2275 ;
        RECT  0.0 33.8525 12.3 33.9175 ;
        RECT  0.0 36.5425 12.3 36.6075 ;
        RECT  0.0 39.2325 12.3 39.2975 ;
        RECT  6.92 8.5025 7.2975 8.5675 ;
        RECT  6.645 9.8475 7.5025 9.9125 ;
        RECT  6.92 13.8825 7.7075 13.9475 ;
        RECT  6.645 15.2275 7.9125 15.2925 ;
        RECT  6.92 8.2975 7.0575 8.3625 ;
        RECT  6.92 10.9875 7.0575 11.0525 ;
        RECT  6.92 13.6775 7.0575 13.7425 ;
        RECT  6.92 16.3675 7.0575 16.4325 ;
        RECT  0.0 9.6425 6.92 9.7075 ;
        RECT  0.0 12.3325 6.92 12.3975 ;
        RECT  0.0 15.0225 6.92 15.0875 ;
        RECT  0.0 17.7125 6.92 17.7775 ;
        RECT  6.92 7.535 7.2975 7.6 ;
        RECT  6.92 6.83 7.5025 6.895 ;
        RECT  6.92 6.125 7.7075 6.19 ;
        RECT  6.92 5.42 7.9125 5.485 ;
        RECT  6.92 7.8875 8.3875 7.9525 ;
        RECT  6.92 7.1825 8.3875 7.2475 ;
        RECT  6.92 6.4775 8.3875 6.5425 ;
        RECT  6.92 5.7725 8.3875 5.8375 ;
        RECT  6.92 5.0675 8.3875 5.1325 ;
        RECT  3.69 4.8625 3.755 4.9275 ;
        RECT  3.69 4.895 3.755 5.1 ;
        RECT  0.0 4.8625 3.7225 4.9275 ;
        RECT  6.65 4.8625 6.715 4.9275 ;
        RECT  6.65 4.895 6.715 5.1 ;
        RECT  0.0 4.8625 6.6825 4.9275 ;
        RECT  1.7 4.8625 1.765 4.9275 ;
        RECT  1.7 4.895 1.765 5.1 ;
        RECT  0.0 4.8625 1.7325 4.9275 ;
        RECT  4.66 4.8625 4.725 4.9275 ;
        RECT  4.66 4.895 4.725 5.1 ;
        RECT  0.0 4.8625 4.6925 4.9275 ;
        RECT  9.4575 3.795 10.345 3.86 ;
        RECT  9.0475 1.61 10.345 1.675 ;
        RECT  9.2525 3.1575 10.345 3.2225 ;
        RECT  9.4575 41.395 10.345 41.46 ;
        RECT  9.6625 10.2975 10.345 10.3625 ;
        RECT  9.8675 14.3225 10.345 14.3875 ;
        RECT  0.685 8.0925 0.75 8.1575 ;
        RECT  0.685 7.92 0.75 8.125 ;
        RECT  0.7175 8.0925 8.8725 8.1575 ;
        RECT  4.665 40.7825 8.8725 40.8475 ;
        RECT  10.345 41.955 11.95 42.02 ;
        RECT  10.345 18.895 11.95 18.96 ;
        RECT  10.345 10.4275 11.95 10.4925 ;
        RECT  10.345 6.8 11.95 6.865 ;
        RECT  10.345 9.76 11.95 9.825 ;
        RECT  10.345 4.81 11.95 4.875 ;
        RECT  10.345 7.77 11.95 7.835 ;
        RECT  10.345 1.74 11.95 1.805 ;
        RECT  8.6025 3.0275 10.345 3.0925 ;
        RECT  8.6025 14.4525 10.345 14.5175 ;
        RECT  8.6025 3.955 10.345 4.02 ;
        RECT  8.6025 11.23 10.345 11.295 ;
        RECT  11.95 0.0 12.3 42.02 ;
        RECT  0.0 0.0 0.35 42.02 ;
        RECT  10.255 24.5775 11.845 24.6425 ;
        RECT  10.255 19.1975 11.845 19.2625 ;
        RECT  10.255 21.8875 11.845 21.9525 ;
        RECT  10.255 40.4375 11.845 40.5025 ;
        RECT  10.255 29.9575 11.845 30.0225 ;
        RECT  10.255 27.2675 11.845 27.3325 ;
        RECT  10.255 37.7475 11.845 37.8125 ;
        RECT  10.255 35.0575 11.845 35.1225 ;
        RECT  10.255 24.2975 11.845 24.3625 ;
        RECT  10.255 26.9875 11.845 27.0525 ;
        RECT  10.255 21.6075 11.845 21.6725 ;
        RECT  10.255 38.0275 11.845 38.0925 ;
        RECT  10.255 32.6475 11.845 32.7125 ;
        RECT  10.255 32.3675 11.845 32.4325 ;
        RECT  10.255 20.4025 11.845 20.4675 ;
        RECT  10.255 23.0925 11.845 23.1575 ;
        RECT  10.255 25.7825 11.845 25.8475 ;
        RECT  10.255 28.4725 11.845 28.5375 ;
        RECT  10.255 31.1625 11.845 31.2275 ;
        RECT  10.255 33.8525 11.845 33.9175 ;
        RECT  10.255 36.5425 11.845 36.6075 ;
        RECT  10.255 39.2325 11.845 39.2975 ;
        RECT  10.255 19.0575 11.845 19.1225 ;
        RECT  10.255 21.7475 11.845 21.8125 ;
        RECT  10.255 24.4375 11.845 24.5025 ;
        RECT  10.255 27.1275 11.845 27.1925 ;
        RECT  10.255 29.8175 11.845 29.8825 ;
        RECT  10.255 32.5075 11.845 32.5725 ;
        RECT  10.255 35.1975 11.845 35.2625 ;
        RECT  10.255 37.8875 11.845 37.9525 ;
        RECT  10.255 40.5775 11.845 40.6425 ;
        RECT  10.255 35.3375 11.845 35.4025 ;
        RECT  10.255 29.6775 11.845 29.7425 ;
        RECT  11.015 20.2025 11.08 20.3375 ;
        RECT  10.83 20.2025 10.895 20.3375 ;
        RECT  10.315 20.2025 10.38 20.3375 ;
        RECT  10.5 20.2025 10.565 20.3375 ;
        RECT  10.83 19.7375 10.895 19.8725 ;
        RECT  11.015 19.7375 11.08 19.8725 ;
        RECT  10.5 19.7375 10.565 19.8725 ;
        RECT  10.315 19.7375 10.38 19.8725 ;
        RECT  10.935 19.3475 11.0 19.4825 ;
        RECT  10.75 19.3475 10.815 19.4825 ;
        RECT  10.58 19.3475 10.645 19.4825 ;
        RECT  10.395 19.3475 10.46 19.4825 ;
        RECT  11.0175 19.84 11.0825 19.975 ;
        RECT  11.0175 19.84 11.0825 19.975 ;
        RECT  11.0175 19.84 11.0825 19.975 ;
        RECT  11.0175 19.84 11.0825 19.975 ;
        RECT  11.0175 19.84 11.0825 19.975 ;
        RECT  11.0175 19.84 11.0825 19.975 ;
        RECT  10.625 20.4025 10.76 20.4675 ;
        RECT  10.2775 19.0575 10.4125 19.1225 ;
        RECT  10.9825 19.0575 11.1175 19.1225 ;
        RECT  10.6125 19.1975 10.7475 19.2625 ;
        RECT  11.0175 19.84 11.0825 19.975 ;
        RECT  11.0175 19.84 11.0825 19.975 ;
        RECT  11.0175 19.84 11.0825 19.975 ;
        RECT  11.0175 19.84 11.0825 19.975 ;
        RECT  10.5175 20.0875 10.6525 20.1525 ;
        RECT  10.5175 20.0875 10.6525 20.1525 ;
        RECT  10.7425 19.9375 10.8775 20.0025 ;
        RECT  10.7425 19.9375 10.8775 20.0025 ;
        RECT  11.0175 19.84 11.0825 19.975 ;
        RECT  11.0175 19.84 11.0825 19.975 ;
        RECT  11.0175 19.84 11.0825 19.975 ;
        RECT  11.0175 19.84 11.0825 19.975 ;
        RECT  10.5675 19.3475 10.6325 19.4825 ;
        RECT  10.3125 19.84 10.3775 19.975 ;
        RECT  10.3125 19.84 10.3775 19.975 ;
        RECT  10.3125 19.84 10.3775 19.975 ;
        RECT  10.3125 19.84 10.3775 19.975 ;
        RECT  10.3125 19.84 10.3775 19.975 ;
        RECT  10.3125 19.84 10.3775 19.975 ;
        RECT  11.0175 19.84 11.0825 19.975 ;
        RECT  11.0175 19.84 11.0825 19.975 ;
        RECT  11.0175 19.84 11.0825 19.975 ;
        RECT  11.0175 19.84 11.0825 19.975 ;
        RECT  10.7625 19.3475 10.8275 19.4825 ;
        RECT  10.63 19.0575 10.765 19.1225 ;
        RECT  10.63 19.0575 10.765 19.1225 ;
        RECT  10.9825 19.0575 11.1175 19.1225 ;
        RECT  10.625 20.4025 10.76 20.4675 ;
        RECT  10.9825 19.0575 11.1175 19.1225 ;
        RECT  10.9825 19.0575 11.1175 19.1225 ;
        RECT  11.0175 19.84 11.0825 19.975 ;
        RECT  11.0175 19.84 11.0825 19.975 ;
        RECT  11.0175 19.84 11.0825 19.975 ;
        RECT  11.0175 19.84 11.0825 19.975 ;
        RECT  11.0175 19.84 11.0825 19.975 ;
        RECT  11.0175 19.84 11.0825 19.975 ;
        RECT  10.2775 19.0575 10.4125 19.1225 ;
        RECT  10.6375 20.4025 10.7375 20.465 ;
        RECT  10.6375 20.405 10.7375 20.4675 ;
        RECT  10.965 19.2 11.0175 19.2625 ;
        RECT  10.6375 20.4025 10.7375 20.465 ;
        RECT  11.015 20.2025 11.085 20.4025 ;
        RECT  11.015 19.7375 11.085 19.8725 ;
        RECT  11.015 19.7375 11.085 19.8725 ;
        RECT  10.255 19.0575 11.14 19.1225 ;
        RECT  10.83 19.5725 11.005 19.6375 ;
        RECT  10.31 19.7375 10.38 19.8725 ;
        RECT  10.5 19.5725 10.565 20.3125 ;
        RECT  10.6375 20.405 10.7375 20.4675 ;
        RECT  10.26 19.2 10.3125 19.2625 ;
        RECT  11.015 19.7375 11.085 19.8725 ;
        RECT  10.255 20.4025 11.14 20.4675 ;
        RECT  10.83 19.5725 10.895 20.2025 ;
        RECT  11.015 19.7375 11.085 19.8725 ;
        RECT  11.015 19.7375 11.085 19.8725 ;
        RECT  10.395 19.3475 10.465 19.6375 ;
        RECT  10.31 19.7375 10.38 19.8725 ;
        RECT  10.255 19.1975 11.14 19.2625 ;
        RECT  11.015 19.7375 11.085 19.8725 ;
        RECT  11.015 20.2025 11.085 20.4025 ;
        RECT  10.31 20.2025 10.38 20.4025 ;
        RECT  10.935 19.3475 11.005 19.6375 ;
        RECT  10.395 19.5725 10.565 19.6375 ;
        RECT  10.255 19.1975 11.14 19.2625 ;
        RECT  10.255 19.0575 11.14 19.1225 ;
        RECT  10.255 20.4025 11.14 20.4675 ;
        RECT  11.015 20.5325 11.08 20.6675 ;
        RECT  10.83 20.5325 10.895 20.6675 ;
        RECT  10.315 20.5325 10.38 20.6675 ;
        RECT  10.5 20.5325 10.565 20.6675 ;
        RECT  10.83 20.9975 10.895 21.1325 ;
        RECT  11.015 20.9975 11.08 21.1325 ;
        RECT  10.5 20.9975 10.565 21.1325 ;
        RECT  10.315 20.9975 10.38 21.1325 ;
        RECT  10.935 21.3875 11.0 21.5225 ;
        RECT  10.75 21.3875 10.815 21.5225 ;
        RECT  10.58 21.3875 10.645 21.5225 ;
        RECT  10.395 21.3875 10.46 21.5225 ;
        RECT  11.0175 20.895 11.0825 21.03 ;
        RECT  11.0175 20.895 11.0825 21.03 ;
        RECT  11.0175 20.895 11.0825 21.03 ;
        RECT  11.0175 20.895 11.0825 21.03 ;
        RECT  11.0175 20.895 11.0825 21.03 ;
        RECT  11.0175 20.895 11.0825 21.03 ;
        RECT  10.625 20.4025 10.76 20.4675 ;
        RECT  10.2775 21.7475 10.4125 21.8125 ;
        RECT  10.9825 21.7475 11.1175 21.8125 ;
        RECT  10.6125 21.6075 10.7475 21.6725 ;
        RECT  11.0175 20.895 11.0825 21.03 ;
        RECT  11.0175 20.895 11.0825 21.03 ;
        RECT  11.0175 20.895 11.0825 21.03 ;
        RECT  11.0175 20.895 11.0825 21.03 ;
        RECT  10.5175 20.7175 10.6525 20.7825 ;
        RECT  10.5175 20.7175 10.6525 20.7825 ;
        RECT  10.7425 20.8675 10.8775 20.9325 ;
        RECT  10.7425 20.8675 10.8775 20.9325 ;
        RECT  11.0175 20.895 11.0825 21.03 ;
        RECT  11.0175 20.895 11.0825 21.03 ;
        RECT  11.0175 20.895 11.0825 21.03 ;
        RECT  11.0175 20.895 11.0825 21.03 ;
        RECT  10.5675 21.3875 10.6325 21.5225 ;
        RECT  10.3125 20.895 10.3775 21.03 ;
        RECT  10.3125 20.895 10.3775 21.03 ;
        RECT  10.3125 20.895 10.3775 21.03 ;
        RECT  10.3125 20.895 10.3775 21.03 ;
        RECT  10.3125 20.895 10.3775 21.03 ;
        RECT  10.3125 20.895 10.3775 21.03 ;
        RECT  11.0175 20.895 11.0825 21.03 ;
        RECT  11.0175 20.895 11.0825 21.03 ;
        RECT  11.0175 20.895 11.0825 21.03 ;
        RECT  11.0175 20.895 11.0825 21.03 ;
        RECT  10.7625 21.3875 10.8275 21.5225 ;
        RECT  10.63 21.7475 10.765 21.8125 ;
        RECT  10.63 21.7475 10.765 21.8125 ;
        RECT  10.9825 21.7475 11.1175 21.8125 ;
        RECT  10.625 20.4025 10.76 20.4675 ;
        RECT  10.9825 21.7475 11.1175 21.8125 ;
        RECT  10.9825 21.7475 11.1175 21.8125 ;
        RECT  11.0175 20.895 11.0825 21.03 ;
        RECT  11.0175 20.895 11.0825 21.03 ;
        RECT  11.0175 20.895 11.0825 21.03 ;
        RECT  11.0175 20.895 11.0825 21.03 ;
        RECT  11.0175 20.895 11.0825 21.03 ;
        RECT  11.0175 20.895 11.0825 21.03 ;
        RECT  10.2775 21.7475 10.4125 21.8125 ;
        RECT  10.6375 20.405 10.7375 20.4675 ;
        RECT  10.6375 20.4025 10.7375 20.465 ;
        RECT  10.965 21.6075 11.0175 21.67 ;
        RECT  10.6375 20.405 10.7375 20.4675 ;
        RECT  11.015 20.4675 11.085 20.6675 ;
        RECT  11.015 20.9975 11.085 21.1325 ;
        RECT  11.015 20.9975 11.085 21.1325 ;
        RECT  10.255 21.7475 11.14 21.8125 ;
        RECT  10.83 21.2325 11.005 21.2975 ;
        RECT  10.31 20.9975 10.38 21.1325 ;
        RECT  10.5 20.5575 10.565 21.2975 ;
        RECT  10.6375 20.4025 10.7375 20.465 ;
        RECT  10.26 21.6075 10.3125 21.67 ;
        RECT  11.015 20.9975 11.085 21.1325 ;
        RECT  10.255 20.4025 11.14 20.4675 ;
        RECT  10.83 20.6675 10.895 21.2975 ;
        RECT  11.015 20.9975 11.085 21.1325 ;
        RECT  11.015 20.9975 11.085 21.1325 ;
        RECT  10.395 21.2325 10.465 21.5225 ;
        RECT  10.31 20.9975 10.38 21.1325 ;
        RECT  10.255 21.6075 11.14 21.6725 ;
        RECT  11.015 20.9975 11.085 21.1325 ;
        RECT  11.015 20.4675 11.085 20.6675 ;
        RECT  10.31 20.4675 10.38 20.6675 ;
        RECT  10.935 21.2325 11.005 21.5225 ;
        RECT  10.395 21.2325 10.565 21.2975 ;
        RECT  10.255 21.6075 11.14 21.6725 ;
        RECT  10.255 21.7475 11.14 21.8125 ;
        RECT  10.255 20.4025 11.14 20.4675 ;
        RECT  11.015 22.8925 11.08 23.0275 ;
        RECT  10.83 22.8925 10.895 23.0275 ;
        RECT  10.315 22.8925 10.38 23.0275 ;
        RECT  10.5 22.8925 10.565 23.0275 ;
        RECT  10.83 22.4275 10.895 22.5625 ;
        RECT  11.015 22.4275 11.08 22.5625 ;
        RECT  10.5 22.4275 10.565 22.5625 ;
        RECT  10.315 22.4275 10.38 22.5625 ;
        RECT  10.935 22.0375 11.0 22.1725 ;
        RECT  10.75 22.0375 10.815 22.1725 ;
        RECT  10.58 22.0375 10.645 22.1725 ;
        RECT  10.395 22.0375 10.46 22.1725 ;
        RECT  11.0175 22.53 11.0825 22.665 ;
        RECT  11.0175 22.53 11.0825 22.665 ;
        RECT  11.0175 22.53 11.0825 22.665 ;
        RECT  11.0175 22.53 11.0825 22.665 ;
        RECT  11.0175 22.53 11.0825 22.665 ;
        RECT  11.0175 22.53 11.0825 22.665 ;
        RECT  10.625 23.0925 10.76 23.1575 ;
        RECT  10.2775 21.7475 10.4125 21.8125 ;
        RECT  10.9825 21.7475 11.1175 21.8125 ;
        RECT  10.6125 21.8875 10.7475 21.9525 ;
        RECT  11.0175 22.53 11.0825 22.665 ;
        RECT  11.0175 22.53 11.0825 22.665 ;
        RECT  11.0175 22.53 11.0825 22.665 ;
        RECT  11.0175 22.53 11.0825 22.665 ;
        RECT  10.5175 22.7775 10.6525 22.8425 ;
        RECT  10.5175 22.7775 10.6525 22.8425 ;
        RECT  10.7425 22.6275 10.8775 22.6925 ;
        RECT  10.7425 22.6275 10.8775 22.6925 ;
        RECT  11.0175 22.53 11.0825 22.665 ;
        RECT  11.0175 22.53 11.0825 22.665 ;
        RECT  11.0175 22.53 11.0825 22.665 ;
        RECT  11.0175 22.53 11.0825 22.665 ;
        RECT  10.5675 22.0375 10.6325 22.1725 ;
        RECT  10.3125 22.53 10.3775 22.665 ;
        RECT  10.3125 22.53 10.3775 22.665 ;
        RECT  10.3125 22.53 10.3775 22.665 ;
        RECT  10.3125 22.53 10.3775 22.665 ;
        RECT  10.3125 22.53 10.3775 22.665 ;
        RECT  10.3125 22.53 10.3775 22.665 ;
        RECT  11.0175 22.53 11.0825 22.665 ;
        RECT  11.0175 22.53 11.0825 22.665 ;
        RECT  11.0175 22.53 11.0825 22.665 ;
        RECT  11.0175 22.53 11.0825 22.665 ;
        RECT  10.7625 22.0375 10.8275 22.1725 ;
        RECT  10.63 21.7475 10.765 21.8125 ;
        RECT  10.63 21.7475 10.765 21.8125 ;
        RECT  10.9825 21.7475 11.1175 21.8125 ;
        RECT  10.625 23.0925 10.76 23.1575 ;
        RECT  10.9825 21.7475 11.1175 21.8125 ;
        RECT  10.9825 21.7475 11.1175 21.8125 ;
        RECT  11.0175 22.53 11.0825 22.665 ;
        RECT  11.0175 22.53 11.0825 22.665 ;
        RECT  11.0175 22.53 11.0825 22.665 ;
        RECT  11.0175 22.53 11.0825 22.665 ;
        RECT  11.0175 22.53 11.0825 22.665 ;
        RECT  11.0175 22.53 11.0825 22.665 ;
        RECT  10.2775 21.7475 10.4125 21.8125 ;
        RECT  10.6375 23.0925 10.7375 23.155 ;
        RECT  10.6375 23.095 10.7375 23.1575 ;
        RECT  10.965 21.89 11.0175 21.9525 ;
        RECT  10.6375 23.0925 10.7375 23.155 ;
        RECT  11.015 22.8925 11.085 23.0925 ;
        RECT  11.015 22.4275 11.085 22.5625 ;
        RECT  11.015 22.4275 11.085 22.5625 ;
        RECT  10.255 21.7475 11.14 21.8125 ;
        RECT  10.83 22.2625 11.005 22.3275 ;
        RECT  10.31 22.4275 10.38 22.5625 ;
        RECT  10.5 22.2625 10.565 23.0025 ;
        RECT  10.6375 23.095 10.7375 23.1575 ;
        RECT  10.26 21.89 10.3125 21.9525 ;
        RECT  11.015 22.4275 11.085 22.5625 ;
        RECT  10.255 23.0925 11.14 23.1575 ;
        RECT  10.83 22.2625 10.895 22.8925 ;
        RECT  11.015 22.4275 11.085 22.5625 ;
        RECT  11.015 22.4275 11.085 22.5625 ;
        RECT  10.395 22.0375 10.465 22.3275 ;
        RECT  10.31 22.4275 10.38 22.5625 ;
        RECT  10.255 21.8875 11.14 21.9525 ;
        RECT  11.015 22.4275 11.085 22.5625 ;
        RECT  11.015 22.8925 11.085 23.0925 ;
        RECT  10.31 22.8925 10.38 23.0925 ;
        RECT  10.935 22.0375 11.005 22.3275 ;
        RECT  10.395 22.2625 10.565 22.3275 ;
        RECT  10.255 21.8875 11.14 21.9525 ;
        RECT  10.255 21.7475 11.14 21.8125 ;
        RECT  10.255 23.0925 11.14 23.1575 ;
        RECT  11.015 23.2225 11.08 23.3575 ;
        RECT  10.83 23.2225 10.895 23.3575 ;
        RECT  10.315 23.2225 10.38 23.3575 ;
        RECT  10.5 23.2225 10.565 23.3575 ;
        RECT  10.83 23.6875 10.895 23.8225 ;
        RECT  11.015 23.6875 11.08 23.8225 ;
        RECT  10.5 23.6875 10.565 23.8225 ;
        RECT  10.315 23.6875 10.38 23.8225 ;
        RECT  10.935 24.0775 11.0 24.2125 ;
        RECT  10.75 24.0775 10.815 24.2125 ;
        RECT  10.58 24.0775 10.645 24.2125 ;
        RECT  10.395 24.0775 10.46 24.2125 ;
        RECT  11.0175 23.585 11.0825 23.72 ;
        RECT  11.0175 23.585 11.0825 23.72 ;
        RECT  11.0175 23.585 11.0825 23.72 ;
        RECT  11.0175 23.585 11.0825 23.72 ;
        RECT  11.0175 23.585 11.0825 23.72 ;
        RECT  11.0175 23.585 11.0825 23.72 ;
        RECT  10.625 23.0925 10.76 23.1575 ;
        RECT  10.2775 24.4375 10.4125 24.5025 ;
        RECT  10.9825 24.4375 11.1175 24.5025 ;
        RECT  10.6125 24.2975 10.7475 24.3625 ;
        RECT  11.0175 23.585 11.0825 23.72 ;
        RECT  11.0175 23.585 11.0825 23.72 ;
        RECT  11.0175 23.585 11.0825 23.72 ;
        RECT  11.0175 23.585 11.0825 23.72 ;
        RECT  10.5175 23.4075 10.6525 23.4725 ;
        RECT  10.5175 23.4075 10.6525 23.4725 ;
        RECT  10.7425 23.5575 10.8775 23.6225 ;
        RECT  10.7425 23.5575 10.8775 23.6225 ;
        RECT  11.0175 23.585 11.0825 23.72 ;
        RECT  11.0175 23.585 11.0825 23.72 ;
        RECT  11.0175 23.585 11.0825 23.72 ;
        RECT  11.0175 23.585 11.0825 23.72 ;
        RECT  10.5675 24.0775 10.6325 24.2125 ;
        RECT  10.3125 23.585 10.3775 23.72 ;
        RECT  10.3125 23.585 10.3775 23.72 ;
        RECT  10.3125 23.585 10.3775 23.72 ;
        RECT  10.3125 23.585 10.3775 23.72 ;
        RECT  10.3125 23.585 10.3775 23.72 ;
        RECT  10.3125 23.585 10.3775 23.72 ;
        RECT  11.0175 23.585 11.0825 23.72 ;
        RECT  11.0175 23.585 11.0825 23.72 ;
        RECT  11.0175 23.585 11.0825 23.72 ;
        RECT  11.0175 23.585 11.0825 23.72 ;
        RECT  10.7625 24.0775 10.8275 24.2125 ;
        RECT  10.63 24.4375 10.765 24.5025 ;
        RECT  10.63 24.4375 10.765 24.5025 ;
        RECT  10.9825 24.4375 11.1175 24.5025 ;
        RECT  10.625 23.0925 10.76 23.1575 ;
        RECT  10.9825 24.4375 11.1175 24.5025 ;
        RECT  10.9825 24.4375 11.1175 24.5025 ;
        RECT  11.0175 23.585 11.0825 23.72 ;
        RECT  11.0175 23.585 11.0825 23.72 ;
        RECT  11.0175 23.585 11.0825 23.72 ;
        RECT  11.0175 23.585 11.0825 23.72 ;
        RECT  11.0175 23.585 11.0825 23.72 ;
        RECT  11.0175 23.585 11.0825 23.72 ;
        RECT  10.2775 24.4375 10.4125 24.5025 ;
        RECT  10.6375 23.095 10.7375 23.1575 ;
        RECT  10.6375 23.0925 10.7375 23.155 ;
        RECT  10.965 24.2975 11.0175 24.36 ;
        RECT  10.6375 23.095 10.7375 23.1575 ;
        RECT  11.015 23.1575 11.085 23.3575 ;
        RECT  11.015 23.6875 11.085 23.8225 ;
        RECT  11.015 23.6875 11.085 23.8225 ;
        RECT  10.255 24.4375 11.14 24.5025 ;
        RECT  10.83 23.9225 11.005 23.9875 ;
        RECT  10.31 23.6875 10.38 23.8225 ;
        RECT  10.5 23.2475 10.565 23.9875 ;
        RECT  10.6375 23.0925 10.7375 23.155 ;
        RECT  10.26 24.2975 10.3125 24.36 ;
        RECT  11.015 23.6875 11.085 23.8225 ;
        RECT  10.255 23.0925 11.14 23.1575 ;
        RECT  10.83 23.3575 10.895 23.9875 ;
        RECT  11.015 23.6875 11.085 23.8225 ;
        RECT  11.015 23.6875 11.085 23.8225 ;
        RECT  10.395 23.9225 10.465 24.2125 ;
        RECT  10.31 23.6875 10.38 23.8225 ;
        RECT  10.255 24.2975 11.14 24.3625 ;
        RECT  11.015 23.6875 11.085 23.8225 ;
        RECT  11.015 23.1575 11.085 23.3575 ;
        RECT  10.31 23.1575 10.38 23.3575 ;
        RECT  10.935 23.9225 11.005 24.2125 ;
        RECT  10.395 23.9225 10.565 23.9875 ;
        RECT  10.255 24.2975 11.14 24.3625 ;
        RECT  10.255 24.4375 11.14 24.5025 ;
        RECT  10.255 23.0925 11.14 23.1575 ;
        RECT  11.015 25.5825 11.08 25.7175 ;
        RECT  10.83 25.5825 10.895 25.7175 ;
        RECT  10.315 25.5825 10.38 25.7175 ;
        RECT  10.5 25.5825 10.565 25.7175 ;
        RECT  10.83 25.1175 10.895 25.2525 ;
        RECT  11.015 25.1175 11.08 25.2525 ;
        RECT  10.5 25.1175 10.565 25.2525 ;
        RECT  10.315 25.1175 10.38 25.2525 ;
        RECT  10.935 24.7275 11.0 24.8625 ;
        RECT  10.75 24.7275 10.815 24.8625 ;
        RECT  10.58 24.7275 10.645 24.8625 ;
        RECT  10.395 24.7275 10.46 24.8625 ;
        RECT  11.0175 25.22 11.0825 25.355 ;
        RECT  11.0175 25.22 11.0825 25.355 ;
        RECT  11.0175 25.22 11.0825 25.355 ;
        RECT  11.0175 25.22 11.0825 25.355 ;
        RECT  11.0175 25.22 11.0825 25.355 ;
        RECT  11.0175 25.22 11.0825 25.355 ;
        RECT  10.625 25.7825 10.76 25.8475 ;
        RECT  10.2775 24.4375 10.4125 24.5025 ;
        RECT  10.9825 24.4375 11.1175 24.5025 ;
        RECT  10.6125 24.5775 10.7475 24.6425 ;
        RECT  11.0175 25.22 11.0825 25.355 ;
        RECT  11.0175 25.22 11.0825 25.355 ;
        RECT  11.0175 25.22 11.0825 25.355 ;
        RECT  11.0175 25.22 11.0825 25.355 ;
        RECT  10.5175 25.4675 10.6525 25.5325 ;
        RECT  10.5175 25.4675 10.6525 25.5325 ;
        RECT  10.7425 25.3175 10.8775 25.3825 ;
        RECT  10.7425 25.3175 10.8775 25.3825 ;
        RECT  11.0175 25.22 11.0825 25.355 ;
        RECT  11.0175 25.22 11.0825 25.355 ;
        RECT  11.0175 25.22 11.0825 25.355 ;
        RECT  11.0175 25.22 11.0825 25.355 ;
        RECT  10.5675 24.7275 10.6325 24.8625 ;
        RECT  10.3125 25.22 10.3775 25.355 ;
        RECT  10.3125 25.22 10.3775 25.355 ;
        RECT  10.3125 25.22 10.3775 25.355 ;
        RECT  10.3125 25.22 10.3775 25.355 ;
        RECT  10.3125 25.22 10.3775 25.355 ;
        RECT  10.3125 25.22 10.3775 25.355 ;
        RECT  11.0175 25.22 11.0825 25.355 ;
        RECT  11.0175 25.22 11.0825 25.355 ;
        RECT  11.0175 25.22 11.0825 25.355 ;
        RECT  11.0175 25.22 11.0825 25.355 ;
        RECT  10.7625 24.7275 10.8275 24.8625 ;
        RECT  10.63 24.4375 10.765 24.5025 ;
        RECT  10.63 24.4375 10.765 24.5025 ;
        RECT  10.9825 24.4375 11.1175 24.5025 ;
        RECT  10.625 25.7825 10.76 25.8475 ;
        RECT  10.9825 24.4375 11.1175 24.5025 ;
        RECT  10.9825 24.4375 11.1175 24.5025 ;
        RECT  11.0175 25.22 11.0825 25.355 ;
        RECT  11.0175 25.22 11.0825 25.355 ;
        RECT  11.0175 25.22 11.0825 25.355 ;
        RECT  11.0175 25.22 11.0825 25.355 ;
        RECT  11.0175 25.22 11.0825 25.355 ;
        RECT  11.0175 25.22 11.0825 25.355 ;
        RECT  10.2775 24.4375 10.4125 24.5025 ;
        RECT  10.6375 25.7825 10.7375 25.845 ;
        RECT  10.6375 25.785 10.7375 25.8475 ;
        RECT  10.965 24.58 11.0175 24.6425 ;
        RECT  10.6375 25.7825 10.7375 25.845 ;
        RECT  11.015 25.5825 11.085 25.7825 ;
        RECT  11.015 25.1175 11.085 25.2525 ;
        RECT  11.015 25.1175 11.085 25.2525 ;
        RECT  10.255 24.4375 11.14 24.5025 ;
        RECT  10.83 24.9525 11.005 25.0175 ;
        RECT  10.31 25.1175 10.38 25.2525 ;
        RECT  10.5 24.9525 10.565 25.6925 ;
        RECT  10.6375 25.785 10.7375 25.8475 ;
        RECT  10.26 24.58 10.3125 24.6425 ;
        RECT  11.015 25.1175 11.085 25.2525 ;
        RECT  10.255 25.7825 11.14 25.8475 ;
        RECT  10.83 24.9525 10.895 25.5825 ;
        RECT  11.015 25.1175 11.085 25.2525 ;
        RECT  11.015 25.1175 11.085 25.2525 ;
        RECT  10.395 24.7275 10.465 25.0175 ;
        RECT  10.31 25.1175 10.38 25.2525 ;
        RECT  10.255 24.5775 11.14 24.6425 ;
        RECT  11.015 25.1175 11.085 25.2525 ;
        RECT  11.015 25.5825 11.085 25.7825 ;
        RECT  10.31 25.5825 10.38 25.7825 ;
        RECT  10.935 24.7275 11.005 25.0175 ;
        RECT  10.395 24.9525 10.565 25.0175 ;
        RECT  10.255 24.5775 11.14 24.6425 ;
        RECT  10.255 24.4375 11.14 24.5025 ;
        RECT  10.255 25.7825 11.14 25.8475 ;
        RECT  11.015 25.9125 11.08 26.0475 ;
        RECT  10.83 25.9125 10.895 26.0475 ;
        RECT  10.315 25.9125 10.38 26.0475 ;
        RECT  10.5 25.9125 10.565 26.0475 ;
        RECT  10.83 26.3775 10.895 26.5125 ;
        RECT  11.015 26.3775 11.08 26.5125 ;
        RECT  10.5 26.3775 10.565 26.5125 ;
        RECT  10.315 26.3775 10.38 26.5125 ;
        RECT  10.935 26.7675 11.0 26.9025 ;
        RECT  10.75 26.7675 10.815 26.9025 ;
        RECT  10.58 26.7675 10.645 26.9025 ;
        RECT  10.395 26.7675 10.46 26.9025 ;
        RECT  11.0175 26.275 11.0825 26.41 ;
        RECT  11.0175 26.275 11.0825 26.41 ;
        RECT  11.0175 26.275 11.0825 26.41 ;
        RECT  11.0175 26.275 11.0825 26.41 ;
        RECT  11.0175 26.275 11.0825 26.41 ;
        RECT  11.0175 26.275 11.0825 26.41 ;
        RECT  10.625 25.7825 10.76 25.8475 ;
        RECT  10.2775 27.1275 10.4125 27.1925 ;
        RECT  10.9825 27.1275 11.1175 27.1925 ;
        RECT  10.6125 26.9875 10.7475 27.0525 ;
        RECT  11.0175 26.275 11.0825 26.41 ;
        RECT  11.0175 26.275 11.0825 26.41 ;
        RECT  11.0175 26.275 11.0825 26.41 ;
        RECT  11.0175 26.275 11.0825 26.41 ;
        RECT  10.5175 26.0975 10.6525 26.1625 ;
        RECT  10.5175 26.0975 10.6525 26.1625 ;
        RECT  10.7425 26.2475 10.8775 26.3125 ;
        RECT  10.7425 26.2475 10.8775 26.3125 ;
        RECT  11.0175 26.275 11.0825 26.41 ;
        RECT  11.0175 26.275 11.0825 26.41 ;
        RECT  11.0175 26.275 11.0825 26.41 ;
        RECT  11.0175 26.275 11.0825 26.41 ;
        RECT  10.5675 26.7675 10.6325 26.9025 ;
        RECT  10.3125 26.275 10.3775 26.41 ;
        RECT  10.3125 26.275 10.3775 26.41 ;
        RECT  10.3125 26.275 10.3775 26.41 ;
        RECT  10.3125 26.275 10.3775 26.41 ;
        RECT  10.3125 26.275 10.3775 26.41 ;
        RECT  10.3125 26.275 10.3775 26.41 ;
        RECT  11.0175 26.275 11.0825 26.41 ;
        RECT  11.0175 26.275 11.0825 26.41 ;
        RECT  11.0175 26.275 11.0825 26.41 ;
        RECT  11.0175 26.275 11.0825 26.41 ;
        RECT  10.7625 26.7675 10.8275 26.9025 ;
        RECT  10.63 27.1275 10.765 27.1925 ;
        RECT  10.63 27.1275 10.765 27.1925 ;
        RECT  10.9825 27.1275 11.1175 27.1925 ;
        RECT  10.625 25.7825 10.76 25.8475 ;
        RECT  10.9825 27.1275 11.1175 27.1925 ;
        RECT  10.9825 27.1275 11.1175 27.1925 ;
        RECT  11.0175 26.275 11.0825 26.41 ;
        RECT  11.0175 26.275 11.0825 26.41 ;
        RECT  11.0175 26.275 11.0825 26.41 ;
        RECT  11.0175 26.275 11.0825 26.41 ;
        RECT  11.0175 26.275 11.0825 26.41 ;
        RECT  11.0175 26.275 11.0825 26.41 ;
        RECT  10.2775 27.1275 10.4125 27.1925 ;
        RECT  10.6375 25.785 10.7375 25.8475 ;
        RECT  10.6375 25.7825 10.7375 25.845 ;
        RECT  10.965 26.9875 11.0175 27.05 ;
        RECT  10.6375 25.785 10.7375 25.8475 ;
        RECT  11.015 25.8475 11.085 26.0475 ;
        RECT  11.015 26.3775 11.085 26.5125 ;
        RECT  11.015 26.3775 11.085 26.5125 ;
        RECT  10.255 27.1275 11.14 27.1925 ;
        RECT  10.83 26.6125 11.005 26.6775 ;
        RECT  10.31 26.3775 10.38 26.5125 ;
        RECT  10.5 25.9375 10.565 26.6775 ;
        RECT  10.6375 25.7825 10.7375 25.845 ;
        RECT  10.26 26.9875 10.3125 27.05 ;
        RECT  11.015 26.3775 11.085 26.5125 ;
        RECT  10.255 25.7825 11.14 25.8475 ;
        RECT  10.83 26.0475 10.895 26.6775 ;
        RECT  11.015 26.3775 11.085 26.5125 ;
        RECT  11.015 26.3775 11.085 26.5125 ;
        RECT  10.395 26.6125 10.465 26.9025 ;
        RECT  10.31 26.3775 10.38 26.5125 ;
        RECT  10.255 26.9875 11.14 27.0525 ;
        RECT  11.015 26.3775 11.085 26.5125 ;
        RECT  11.015 25.8475 11.085 26.0475 ;
        RECT  10.31 25.8475 10.38 26.0475 ;
        RECT  10.935 26.6125 11.005 26.9025 ;
        RECT  10.395 26.6125 10.565 26.6775 ;
        RECT  10.255 26.9875 11.14 27.0525 ;
        RECT  10.255 27.1275 11.14 27.1925 ;
        RECT  10.255 25.7825 11.14 25.8475 ;
        RECT  11.015 28.2725 11.08 28.4075 ;
        RECT  10.83 28.2725 10.895 28.4075 ;
        RECT  10.315 28.2725 10.38 28.4075 ;
        RECT  10.5 28.2725 10.565 28.4075 ;
        RECT  10.83 27.8075 10.895 27.9425 ;
        RECT  11.015 27.8075 11.08 27.9425 ;
        RECT  10.5 27.8075 10.565 27.9425 ;
        RECT  10.315 27.8075 10.38 27.9425 ;
        RECT  10.935 27.4175 11.0 27.5525 ;
        RECT  10.75 27.4175 10.815 27.5525 ;
        RECT  10.58 27.4175 10.645 27.5525 ;
        RECT  10.395 27.4175 10.46 27.5525 ;
        RECT  11.0175 27.91 11.0825 28.045 ;
        RECT  11.0175 27.91 11.0825 28.045 ;
        RECT  11.0175 27.91 11.0825 28.045 ;
        RECT  11.0175 27.91 11.0825 28.045 ;
        RECT  11.0175 27.91 11.0825 28.045 ;
        RECT  11.0175 27.91 11.0825 28.045 ;
        RECT  10.625 28.4725 10.76 28.5375 ;
        RECT  10.2775 27.1275 10.4125 27.1925 ;
        RECT  10.9825 27.1275 11.1175 27.1925 ;
        RECT  10.6125 27.2675 10.7475 27.3325 ;
        RECT  11.0175 27.91 11.0825 28.045 ;
        RECT  11.0175 27.91 11.0825 28.045 ;
        RECT  11.0175 27.91 11.0825 28.045 ;
        RECT  11.0175 27.91 11.0825 28.045 ;
        RECT  10.5175 28.1575 10.6525 28.2225 ;
        RECT  10.5175 28.1575 10.6525 28.2225 ;
        RECT  10.7425 28.0075 10.8775 28.0725 ;
        RECT  10.7425 28.0075 10.8775 28.0725 ;
        RECT  11.0175 27.91 11.0825 28.045 ;
        RECT  11.0175 27.91 11.0825 28.045 ;
        RECT  11.0175 27.91 11.0825 28.045 ;
        RECT  11.0175 27.91 11.0825 28.045 ;
        RECT  10.5675 27.4175 10.6325 27.5525 ;
        RECT  10.3125 27.91 10.3775 28.045 ;
        RECT  10.3125 27.91 10.3775 28.045 ;
        RECT  10.3125 27.91 10.3775 28.045 ;
        RECT  10.3125 27.91 10.3775 28.045 ;
        RECT  10.3125 27.91 10.3775 28.045 ;
        RECT  10.3125 27.91 10.3775 28.045 ;
        RECT  11.0175 27.91 11.0825 28.045 ;
        RECT  11.0175 27.91 11.0825 28.045 ;
        RECT  11.0175 27.91 11.0825 28.045 ;
        RECT  11.0175 27.91 11.0825 28.045 ;
        RECT  10.7625 27.4175 10.8275 27.5525 ;
        RECT  10.63 27.1275 10.765 27.1925 ;
        RECT  10.63 27.1275 10.765 27.1925 ;
        RECT  10.9825 27.1275 11.1175 27.1925 ;
        RECT  10.625 28.4725 10.76 28.5375 ;
        RECT  10.9825 27.1275 11.1175 27.1925 ;
        RECT  10.9825 27.1275 11.1175 27.1925 ;
        RECT  11.0175 27.91 11.0825 28.045 ;
        RECT  11.0175 27.91 11.0825 28.045 ;
        RECT  11.0175 27.91 11.0825 28.045 ;
        RECT  11.0175 27.91 11.0825 28.045 ;
        RECT  11.0175 27.91 11.0825 28.045 ;
        RECT  11.0175 27.91 11.0825 28.045 ;
        RECT  10.2775 27.1275 10.4125 27.1925 ;
        RECT  10.6375 28.4725 10.7375 28.535 ;
        RECT  10.6375 28.475 10.7375 28.5375 ;
        RECT  10.965 27.27 11.0175 27.3325 ;
        RECT  10.6375 28.4725 10.7375 28.535 ;
        RECT  11.015 28.2725 11.085 28.4725 ;
        RECT  11.015 27.8075 11.085 27.9425 ;
        RECT  11.015 27.8075 11.085 27.9425 ;
        RECT  10.255 27.1275 11.14 27.1925 ;
        RECT  10.83 27.6425 11.005 27.7075 ;
        RECT  10.31 27.8075 10.38 27.9425 ;
        RECT  10.5 27.6425 10.565 28.3825 ;
        RECT  10.6375 28.475 10.7375 28.5375 ;
        RECT  10.26 27.27 10.3125 27.3325 ;
        RECT  11.015 27.8075 11.085 27.9425 ;
        RECT  10.255 28.4725 11.14 28.5375 ;
        RECT  10.83 27.6425 10.895 28.2725 ;
        RECT  11.015 27.8075 11.085 27.9425 ;
        RECT  11.015 27.8075 11.085 27.9425 ;
        RECT  10.395 27.4175 10.465 27.7075 ;
        RECT  10.31 27.8075 10.38 27.9425 ;
        RECT  10.255 27.2675 11.14 27.3325 ;
        RECT  11.015 27.8075 11.085 27.9425 ;
        RECT  11.015 28.2725 11.085 28.4725 ;
        RECT  10.31 28.2725 10.38 28.4725 ;
        RECT  10.935 27.4175 11.005 27.7075 ;
        RECT  10.395 27.6425 10.565 27.7075 ;
        RECT  10.255 27.2675 11.14 27.3325 ;
        RECT  10.255 27.1275 11.14 27.1925 ;
        RECT  10.255 28.4725 11.14 28.5375 ;
        RECT  11.015 28.6025 11.08 28.7375 ;
        RECT  10.83 28.6025 10.895 28.7375 ;
        RECT  10.315 28.6025 10.38 28.7375 ;
        RECT  10.5 28.6025 10.565 28.7375 ;
        RECT  10.83 29.0675 10.895 29.2025 ;
        RECT  11.015 29.0675 11.08 29.2025 ;
        RECT  10.5 29.0675 10.565 29.2025 ;
        RECT  10.315 29.0675 10.38 29.2025 ;
        RECT  10.935 29.4575 11.0 29.5925 ;
        RECT  10.75 29.4575 10.815 29.5925 ;
        RECT  10.58 29.4575 10.645 29.5925 ;
        RECT  10.395 29.4575 10.46 29.5925 ;
        RECT  11.0175 28.965 11.0825 29.1 ;
        RECT  11.0175 28.965 11.0825 29.1 ;
        RECT  11.0175 28.965 11.0825 29.1 ;
        RECT  11.0175 28.965 11.0825 29.1 ;
        RECT  11.0175 28.965 11.0825 29.1 ;
        RECT  11.0175 28.965 11.0825 29.1 ;
        RECT  10.625 28.4725 10.76 28.5375 ;
        RECT  10.2775 29.8175 10.4125 29.8825 ;
        RECT  10.9825 29.8175 11.1175 29.8825 ;
        RECT  10.6125 29.6775 10.7475 29.7425 ;
        RECT  11.0175 28.965 11.0825 29.1 ;
        RECT  11.0175 28.965 11.0825 29.1 ;
        RECT  11.0175 28.965 11.0825 29.1 ;
        RECT  11.0175 28.965 11.0825 29.1 ;
        RECT  10.5175 28.7875 10.6525 28.8525 ;
        RECT  10.5175 28.7875 10.6525 28.8525 ;
        RECT  10.7425 28.9375 10.8775 29.0025 ;
        RECT  10.7425 28.9375 10.8775 29.0025 ;
        RECT  11.0175 28.965 11.0825 29.1 ;
        RECT  11.0175 28.965 11.0825 29.1 ;
        RECT  11.0175 28.965 11.0825 29.1 ;
        RECT  11.0175 28.965 11.0825 29.1 ;
        RECT  10.5675 29.4575 10.6325 29.5925 ;
        RECT  10.3125 28.965 10.3775 29.1 ;
        RECT  10.3125 28.965 10.3775 29.1 ;
        RECT  10.3125 28.965 10.3775 29.1 ;
        RECT  10.3125 28.965 10.3775 29.1 ;
        RECT  10.3125 28.965 10.3775 29.1 ;
        RECT  10.3125 28.965 10.3775 29.1 ;
        RECT  11.0175 28.965 11.0825 29.1 ;
        RECT  11.0175 28.965 11.0825 29.1 ;
        RECT  11.0175 28.965 11.0825 29.1 ;
        RECT  11.0175 28.965 11.0825 29.1 ;
        RECT  10.7625 29.4575 10.8275 29.5925 ;
        RECT  10.63 29.8175 10.765 29.8825 ;
        RECT  10.63 29.8175 10.765 29.8825 ;
        RECT  10.9825 29.8175 11.1175 29.8825 ;
        RECT  10.625 28.4725 10.76 28.5375 ;
        RECT  10.9825 29.8175 11.1175 29.8825 ;
        RECT  10.9825 29.8175 11.1175 29.8825 ;
        RECT  11.0175 28.965 11.0825 29.1 ;
        RECT  11.0175 28.965 11.0825 29.1 ;
        RECT  11.0175 28.965 11.0825 29.1 ;
        RECT  11.0175 28.965 11.0825 29.1 ;
        RECT  11.0175 28.965 11.0825 29.1 ;
        RECT  11.0175 28.965 11.0825 29.1 ;
        RECT  10.2775 29.8175 10.4125 29.8825 ;
        RECT  10.6375 28.475 10.7375 28.5375 ;
        RECT  10.6375 28.4725 10.7375 28.535 ;
        RECT  10.965 29.6775 11.0175 29.74 ;
        RECT  10.6375 28.475 10.7375 28.5375 ;
        RECT  11.015 28.5375 11.085 28.7375 ;
        RECT  11.015 29.0675 11.085 29.2025 ;
        RECT  11.015 29.0675 11.085 29.2025 ;
        RECT  10.255 29.8175 11.14 29.8825 ;
        RECT  10.83 29.3025 11.005 29.3675 ;
        RECT  10.31 29.0675 10.38 29.2025 ;
        RECT  10.5 28.6275 10.565 29.3675 ;
        RECT  10.6375 28.4725 10.7375 28.535 ;
        RECT  10.26 29.6775 10.3125 29.74 ;
        RECT  11.015 29.0675 11.085 29.2025 ;
        RECT  10.255 28.4725 11.14 28.5375 ;
        RECT  10.83 28.7375 10.895 29.3675 ;
        RECT  11.015 29.0675 11.085 29.2025 ;
        RECT  11.015 29.0675 11.085 29.2025 ;
        RECT  10.395 29.3025 10.465 29.5925 ;
        RECT  10.31 29.0675 10.38 29.2025 ;
        RECT  10.255 29.6775 11.14 29.7425 ;
        RECT  11.015 29.0675 11.085 29.2025 ;
        RECT  11.015 28.5375 11.085 28.7375 ;
        RECT  10.31 28.5375 10.38 28.7375 ;
        RECT  10.935 29.3025 11.005 29.5925 ;
        RECT  10.395 29.3025 10.565 29.3675 ;
        RECT  10.255 29.6775 11.14 29.7425 ;
        RECT  10.255 29.8175 11.14 29.8825 ;
        RECT  10.255 28.4725 11.14 28.5375 ;
        RECT  11.015 30.9625 11.08 31.0975 ;
        RECT  10.83 30.9625 10.895 31.0975 ;
        RECT  10.315 30.9625 10.38 31.0975 ;
        RECT  10.5 30.9625 10.565 31.0975 ;
        RECT  10.83 30.4975 10.895 30.6325 ;
        RECT  11.015 30.4975 11.08 30.6325 ;
        RECT  10.5 30.4975 10.565 30.6325 ;
        RECT  10.315 30.4975 10.38 30.6325 ;
        RECT  10.935 30.1075 11.0 30.2425 ;
        RECT  10.75 30.1075 10.815 30.2425 ;
        RECT  10.58 30.1075 10.645 30.2425 ;
        RECT  10.395 30.1075 10.46 30.2425 ;
        RECT  11.0175 30.6 11.0825 30.735 ;
        RECT  11.0175 30.6 11.0825 30.735 ;
        RECT  11.0175 30.6 11.0825 30.735 ;
        RECT  11.0175 30.6 11.0825 30.735 ;
        RECT  11.0175 30.6 11.0825 30.735 ;
        RECT  11.0175 30.6 11.0825 30.735 ;
        RECT  10.625 31.1625 10.76 31.2275 ;
        RECT  10.2775 29.8175 10.4125 29.8825 ;
        RECT  10.9825 29.8175 11.1175 29.8825 ;
        RECT  10.6125 29.9575 10.7475 30.0225 ;
        RECT  11.0175 30.6 11.0825 30.735 ;
        RECT  11.0175 30.6 11.0825 30.735 ;
        RECT  11.0175 30.6 11.0825 30.735 ;
        RECT  11.0175 30.6 11.0825 30.735 ;
        RECT  10.5175 30.8475 10.6525 30.9125 ;
        RECT  10.5175 30.8475 10.6525 30.9125 ;
        RECT  10.7425 30.6975 10.8775 30.7625 ;
        RECT  10.7425 30.6975 10.8775 30.7625 ;
        RECT  11.0175 30.6 11.0825 30.735 ;
        RECT  11.0175 30.6 11.0825 30.735 ;
        RECT  11.0175 30.6 11.0825 30.735 ;
        RECT  11.0175 30.6 11.0825 30.735 ;
        RECT  10.5675 30.1075 10.6325 30.2425 ;
        RECT  10.3125 30.6 10.3775 30.735 ;
        RECT  10.3125 30.6 10.3775 30.735 ;
        RECT  10.3125 30.6 10.3775 30.735 ;
        RECT  10.3125 30.6 10.3775 30.735 ;
        RECT  10.3125 30.6 10.3775 30.735 ;
        RECT  10.3125 30.6 10.3775 30.735 ;
        RECT  11.0175 30.6 11.0825 30.735 ;
        RECT  11.0175 30.6 11.0825 30.735 ;
        RECT  11.0175 30.6 11.0825 30.735 ;
        RECT  11.0175 30.6 11.0825 30.735 ;
        RECT  10.7625 30.1075 10.8275 30.2425 ;
        RECT  10.63 29.8175 10.765 29.8825 ;
        RECT  10.63 29.8175 10.765 29.8825 ;
        RECT  10.9825 29.8175 11.1175 29.8825 ;
        RECT  10.625 31.1625 10.76 31.2275 ;
        RECT  10.9825 29.8175 11.1175 29.8825 ;
        RECT  10.9825 29.8175 11.1175 29.8825 ;
        RECT  11.0175 30.6 11.0825 30.735 ;
        RECT  11.0175 30.6 11.0825 30.735 ;
        RECT  11.0175 30.6 11.0825 30.735 ;
        RECT  11.0175 30.6 11.0825 30.735 ;
        RECT  11.0175 30.6 11.0825 30.735 ;
        RECT  11.0175 30.6 11.0825 30.735 ;
        RECT  10.2775 29.8175 10.4125 29.8825 ;
        RECT  10.6375 31.1625 10.7375 31.225 ;
        RECT  10.6375 31.165 10.7375 31.2275 ;
        RECT  10.965 29.96 11.0175 30.0225 ;
        RECT  10.6375 31.1625 10.7375 31.225 ;
        RECT  11.015 30.9625 11.085 31.1625 ;
        RECT  11.015 30.4975 11.085 30.6325 ;
        RECT  11.015 30.4975 11.085 30.6325 ;
        RECT  10.255 29.8175 11.14 29.8825 ;
        RECT  10.83 30.3325 11.005 30.3975 ;
        RECT  10.31 30.4975 10.38 30.6325 ;
        RECT  10.5 30.3325 10.565 31.0725 ;
        RECT  10.6375 31.165 10.7375 31.2275 ;
        RECT  10.26 29.96 10.3125 30.0225 ;
        RECT  11.015 30.4975 11.085 30.6325 ;
        RECT  10.255 31.1625 11.14 31.2275 ;
        RECT  10.83 30.3325 10.895 30.9625 ;
        RECT  11.015 30.4975 11.085 30.6325 ;
        RECT  11.015 30.4975 11.085 30.6325 ;
        RECT  10.395 30.1075 10.465 30.3975 ;
        RECT  10.31 30.4975 10.38 30.6325 ;
        RECT  10.255 29.9575 11.14 30.0225 ;
        RECT  11.015 30.4975 11.085 30.6325 ;
        RECT  11.015 30.9625 11.085 31.1625 ;
        RECT  10.31 30.9625 10.38 31.1625 ;
        RECT  10.935 30.1075 11.005 30.3975 ;
        RECT  10.395 30.3325 10.565 30.3975 ;
        RECT  10.255 29.9575 11.14 30.0225 ;
        RECT  10.255 29.8175 11.14 29.8825 ;
        RECT  10.255 31.1625 11.14 31.2275 ;
        RECT  11.015 31.2925 11.08 31.4275 ;
        RECT  10.83 31.2925 10.895 31.4275 ;
        RECT  10.315 31.2925 10.38 31.4275 ;
        RECT  10.5 31.2925 10.565 31.4275 ;
        RECT  10.83 31.7575 10.895 31.8925 ;
        RECT  11.015 31.7575 11.08 31.8925 ;
        RECT  10.5 31.7575 10.565 31.8925 ;
        RECT  10.315 31.7575 10.38 31.8925 ;
        RECT  10.935 32.1475 11.0 32.2825 ;
        RECT  10.75 32.1475 10.815 32.2825 ;
        RECT  10.58 32.1475 10.645 32.2825 ;
        RECT  10.395 32.1475 10.46 32.2825 ;
        RECT  11.0175 31.655 11.0825 31.79 ;
        RECT  11.0175 31.655 11.0825 31.79 ;
        RECT  11.0175 31.655 11.0825 31.79 ;
        RECT  11.0175 31.655 11.0825 31.79 ;
        RECT  11.0175 31.655 11.0825 31.79 ;
        RECT  11.0175 31.655 11.0825 31.79 ;
        RECT  10.625 31.1625 10.76 31.2275 ;
        RECT  10.2775 32.5075 10.4125 32.5725 ;
        RECT  10.9825 32.5075 11.1175 32.5725 ;
        RECT  10.6125 32.3675 10.7475 32.4325 ;
        RECT  11.0175 31.655 11.0825 31.79 ;
        RECT  11.0175 31.655 11.0825 31.79 ;
        RECT  11.0175 31.655 11.0825 31.79 ;
        RECT  11.0175 31.655 11.0825 31.79 ;
        RECT  10.5175 31.4775 10.6525 31.5425 ;
        RECT  10.5175 31.4775 10.6525 31.5425 ;
        RECT  10.7425 31.6275 10.8775 31.6925 ;
        RECT  10.7425 31.6275 10.8775 31.6925 ;
        RECT  11.0175 31.655 11.0825 31.79 ;
        RECT  11.0175 31.655 11.0825 31.79 ;
        RECT  11.0175 31.655 11.0825 31.79 ;
        RECT  11.0175 31.655 11.0825 31.79 ;
        RECT  10.5675 32.1475 10.6325 32.2825 ;
        RECT  10.3125 31.655 10.3775 31.79 ;
        RECT  10.3125 31.655 10.3775 31.79 ;
        RECT  10.3125 31.655 10.3775 31.79 ;
        RECT  10.3125 31.655 10.3775 31.79 ;
        RECT  10.3125 31.655 10.3775 31.79 ;
        RECT  10.3125 31.655 10.3775 31.79 ;
        RECT  11.0175 31.655 11.0825 31.79 ;
        RECT  11.0175 31.655 11.0825 31.79 ;
        RECT  11.0175 31.655 11.0825 31.79 ;
        RECT  11.0175 31.655 11.0825 31.79 ;
        RECT  10.7625 32.1475 10.8275 32.2825 ;
        RECT  10.63 32.5075 10.765 32.5725 ;
        RECT  10.63 32.5075 10.765 32.5725 ;
        RECT  10.9825 32.5075 11.1175 32.5725 ;
        RECT  10.625 31.1625 10.76 31.2275 ;
        RECT  10.9825 32.5075 11.1175 32.5725 ;
        RECT  10.9825 32.5075 11.1175 32.5725 ;
        RECT  11.0175 31.655 11.0825 31.79 ;
        RECT  11.0175 31.655 11.0825 31.79 ;
        RECT  11.0175 31.655 11.0825 31.79 ;
        RECT  11.0175 31.655 11.0825 31.79 ;
        RECT  11.0175 31.655 11.0825 31.79 ;
        RECT  11.0175 31.655 11.0825 31.79 ;
        RECT  10.2775 32.5075 10.4125 32.5725 ;
        RECT  10.6375 31.165 10.7375 31.2275 ;
        RECT  10.6375 31.1625 10.7375 31.225 ;
        RECT  10.965 32.3675 11.0175 32.43 ;
        RECT  10.6375 31.165 10.7375 31.2275 ;
        RECT  11.015 31.2275 11.085 31.4275 ;
        RECT  11.015 31.7575 11.085 31.8925 ;
        RECT  11.015 31.7575 11.085 31.8925 ;
        RECT  10.255 32.5075 11.14 32.5725 ;
        RECT  10.83 31.9925 11.005 32.0575 ;
        RECT  10.31 31.7575 10.38 31.8925 ;
        RECT  10.5 31.3175 10.565 32.0575 ;
        RECT  10.6375 31.1625 10.7375 31.225 ;
        RECT  10.26 32.3675 10.3125 32.43 ;
        RECT  11.015 31.7575 11.085 31.8925 ;
        RECT  10.255 31.1625 11.14 31.2275 ;
        RECT  10.83 31.4275 10.895 32.0575 ;
        RECT  11.015 31.7575 11.085 31.8925 ;
        RECT  11.015 31.7575 11.085 31.8925 ;
        RECT  10.395 31.9925 10.465 32.2825 ;
        RECT  10.31 31.7575 10.38 31.8925 ;
        RECT  10.255 32.3675 11.14 32.4325 ;
        RECT  11.015 31.7575 11.085 31.8925 ;
        RECT  11.015 31.2275 11.085 31.4275 ;
        RECT  10.31 31.2275 10.38 31.4275 ;
        RECT  10.935 31.9925 11.005 32.2825 ;
        RECT  10.395 31.9925 10.565 32.0575 ;
        RECT  10.255 32.3675 11.14 32.4325 ;
        RECT  10.255 32.5075 11.14 32.5725 ;
        RECT  10.255 31.1625 11.14 31.2275 ;
        RECT  11.015 33.6525 11.08 33.7875 ;
        RECT  10.83 33.6525 10.895 33.7875 ;
        RECT  10.315 33.6525 10.38 33.7875 ;
        RECT  10.5 33.6525 10.565 33.7875 ;
        RECT  10.83 33.1875 10.895 33.3225 ;
        RECT  11.015 33.1875 11.08 33.3225 ;
        RECT  10.5 33.1875 10.565 33.3225 ;
        RECT  10.315 33.1875 10.38 33.3225 ;
        RECT  10.935 32.7975 11.0 32.9325 ;
        RECT  10.75 32.7975 10.815 32.9325 ;
        RECT  10.58 32.7975 10.645 32.9325 ;
        RECT  10.395 32.7975 10.46 32.9325 ;
        RECT  11.0175 33.29 11.0825 33.425 ;
        RECT  11.0175 33.29 11.0825 33.425 ;
        RECT  11.0175 33.29 11.0825 33.425 ;
        RECT  11.0175 33.29 11.0825 33.425 ;
        RECT  11.0175 33.29 11.0825 33.425 ;
        RECT  11.0175 33.29 11.0825 33.425 ;
        RECT  10.625 33.8525 10.76 33.9175 ;
        RECT  10.2775 32.5075 10.4125 32.5725 ;
        RECT  10.9825 32.5075 11.1175 32.5725 ;
        RECT  10.6125 32.6475 10.7475 32.7125 ;
        RECT  11.0175 33.29 11.0825 33.425 ;
        RECT  11.0175 33.29 11.0825 33.425 ;
        RECT  11.0175 33.29 11.0825 33.425 ;
        RECT  11.0175 33.29 11.0825 33.425 ;
        RECT  10.5175 33.5375 10.6525 33.6025 ;
        RECT  10.5175 33.5375 10.6525 33.6025 ;
        RECT  10.7425 33.3875 10.8775 33.4525 ;
        RECT  10.7425 33.3875 10.8775 33.4525 ;
        RECT  11.0175 33.29 11.0825 33.425 ;
        RECT  11.0175 33.29 11.0825 33.425 ;
        RECT  11.0175 33.29 11.0825 33.425 ;
        RECT  11.0175 33.29 11.0825 33.425 ;
        RECT  10.5675 32.7975 10.6325 32.9325 ;
        RECT  10.3125 33.29 10.3775 33.425 ;
        RECT  10.3125 33.29 10.3775 33.425 ;
        RECT  10.3125 33.29 10.3775 33.425 ;
        RECT  10.3125 33.29 10.3775 33.425 ;
        RECT  10.3125 33.29 10.3775 33.425 ;
        RECT  10.3125 33.29 10.3775 33.425 ;
        RECT  11.0175 33.29 11.0825 33.425 ;
        RECT  11.0175 33.29 11.0825 33.425 ;
        RECT  11.0175 33.29 11.0825 33.425 ;
        RECT  11.0175 33.29 11.0825 33.425 ;
        RECT  10.7625 32.7975 10.8275 32.9325 ;
        RECT  10.63 32.5075 10.765 32.5725 ;
        RECT  10.63 32.5075 10.765 32.5725 ;
        RECT  10.9825 32.5075 11.1175 32.5725 ;
        RECT  10.625 33.8525 10.76 33.9175 ;
        RECT  10.9825 32.5075 11.1175 32.5725 ;
        RECT  10.9825 32.5075 11.1175 32.5725 ;
        RECT  11.0175 33.29 11.0825 33.425 ;
        RECT  11.0175 33.29 11.0825 33.425 ;
        RECT  11.0175 33.29 11.0825 33.425 ;
        RECT  11.0175 33.29 11.0825 33.425 ;
        RECT  11.0175 33.29 11.0825 33.425 ;
        RECT  11.0175 33.29 11.0825 33.425 ;
        RECT  10.2775 32.5075 10.4125 32.5725 ;
        RECT  10.6375 33.8525 10.7375 33.915 ;
        RECT  10.6375 33.855 10.7375 33.9175 ;
        RECT  10.965 32.65 11.0175 32.7125 ;
        RECT  10.6375 33.8525 10.7375 33.915 ;
        RECT  11.015 33.6525 11.085 33.8525 ;
        RECT  11.015 33.1875 11.085 33.3225 ;
        RECT  11.015 33.1875 11.085 33.3225 ;
        RECT  10.255 32.5075 11.14 32.5725 ;
        RECT  10.83 33.0225 11.005 33.0875 ;
        RECT  10.31 33.1875 10.38 33.3225 ;
        RECT  10.5 33.0225 10.565 33.7625 ;
        RECT  10.6375 33.855 10.7375 33.9175 ;
        RECT  10.26 32.65 10.3125 32.7125 ;
        RECT  11.015 33.1875 11.085 33.3225 ;
        RECT  10.255 33.8525 11.14 33.9175 ;
        RECT  10.83 33.0225 10.895 33.6525 ;
        RECT  11.015 33.1875 11.085 33.3225 ;
        RECT  11.015 33.1875 11.085 33.3225 ;
        RECT  10.395 32.7975 10.465 33.0875 ;
        RECT  10.31 33.1875 10.38 33.3225 ;
        RECT  10.255 32.6475 11.14 32.7125 ;
        RECT  11.015 33.1875 11.085 33.3225 ;
        RECT  11.015 33.6525 11.085 33.8525 ;
        RECT  10.31 33.6525 10.38 33.8525 ;
        RECT  10.935 32.7975 11.005 33.0875 ;
        RECT  10.395 33.0225 10.565 33.0875 ;
        RECT  10.255 32.6475 11.14 32.7125 ;
        RECT  10.255 32.5075 11.14 32.5725 ;
        RECT  10.255 33.8525 11.14 33.9175 ;
        RECT  11.015 33.9825 11.08 34.1175 ;
        RECT  10.83 33.9825 10.895 34.1175 ;
        RECT  10.315 33.9825 10.38 34.1175 ;
        RECT  10.5 33.9825 10.565 34.1175 ;
        RECT  10.83 34.4475 10.895 34.5825 ;
        RECT  11.015 34.4475 11.08 34.5825 ;
        RECT  10.5 34.4475 10.565 34.5825 ;
        RECT  10.315 34.4475 10.38 34.5825 ;
        RECT  10.935 34.8375 11.0 34.9725 ;
        RECT  10.75 34.8375 10.815 34.9725 ;
        RECT  10.58 34.8375 10.645 34.9725 ;
        RECT  10.395 34.8375 10.46 34.9725 ;
        RECT  11.0175 34.345 11.0825 34.48 ;
        RECT  11.0175 34.345 11.0825 34.48 ;
        RECT  11.0175 34.345 11.0825 34.48 ;
        RECT  11.0175 34.345 11.0825 34.48 ;
        RECT  11.0175 34.345 11.0825 34.48 ;
        RECT  11.0175 34.345 11.0825 34.48 ;
        RECT  10.625 33.8525 10.76 33.9175 ;
        RECT  10.2775 35.1975 10.4125 35.2625 ;
        RECT  10.9825 35.1975 11.1175 35.2625 ;
        RECT  10.6125 35.0575 10.7475 35.1225 ;
        RECT  11.0175 34.345 11.0825 34.48 ;
        RECT  11.0175 34.345 11.0825 34.48 ;
        RECT  11.0175 34.345 11.0825 34.48 ;
        RECT  11.0175 34.345 11.0825 34.48 ;
        RECT  10.5175 34.1675 10.6525 34.2325 ;
        RECT  10.5175 34.1675 10.6525 34.2325 ;
        RECT  10.7425 34.3175 10.8775 34.3825 ;
        RECT  10.7425 34.3175 10.8775 34.3825 ;
        RECT  11.0175 34.345 11.0825 34.48 ;
        RECT  11.0175 34.345 11.0825 34.48 ;
        RECT  11.0175 34.345 11.0825 34.48 ;
        RECT  11.0175 34.345 11.0825 34.48 ;
        RECT  10.5675 34.8375 10.6325 34.9725 ;
        RECT  10.3125 34.345 10.3775 34.48 ;
        RECT  10.3125 34.345 10.3775 34.48 ;
        RECT  10.3125 34.345 10.3775 34.48 ;
        RECT  10.3125 34.345 10.3775 34.48 ;
        RECT  10.3125 34.345 10.3775 34.48 ;
        RECT  10.3125 34.345 10.3775 34.48 ;
        RECT  11.0175 34.345 11.0825 34.48 ;
        RECT  11.0175 34.345 11.0825 34.48 ;
        RECT  11.0175 34.345 11.0825 34.48 ;
        RECT  11.0175 34.345 11.0825 34.48 ;
        RECT  10.7625 34.8375 10.8275 34.9725 ;
        RECT  10.63 35.1975 10.765 35.2625 ;
        RECT  10.63 35.1975 10.765 35.2625 ;
        RECT  10.9825 35.1975 11.1175 35.2625 ;
        RECT  10.625 33.8525 10.76 33.9175 ;
        RECT  10.9825 35.1975 11.1175 35.2625 ;
        RECT  10.9825 35.1975 11.1175 35.2625 ;
        RECT  11.0175 34.345 11.0825 34.48 ;
        RECT  11.0175 34.345 11.0825 34.48 ;
        RECT  11.0175 34.345 11.0825 34.48 ;
        RECT  11.0175 34.345 11.0825 34.48 ;
        RECT  11.0175 34.345 11.0825 34.48 ;
        RECT  11.0175 34.345 11.0825 34.48 ;
        RECT  10.2775 35.1975 10.4125 35.2625 ;
        RECT  10.6375 33.855 10.7375 33.9175 ;
        RECT  10.6375 33.8525 10.7375 33.915 ;
        RECT  10.965 35.0575 11.0175 35.12 ;
        RECT  10.6375 33.855 10.7375 33.9175 ;
        RECT  11.015 33.9175 11.085 34.1175 ;
        RECT  11.015 34.4475 11.085 34.5825 ;
        RECT  11.015 34.4475 11.085 34.5825 ;
        RECT  10.255 35.1975 11.14 35.2625 ;
        RECT  10.83 34.6825 11.005 34.7475 ;
        RECT  10.31 34.4475 10.38 34.5825 ;
        RECT  10.5 34.0075 10.565 34.7475 ;
        RECT  10.6375 33.8525 10.7375 33.915 ;
        RECT  10.26 35.0575 10.3125 35.12 ;
        RECT  11.015 34.4475 11.085 34.5825 ;
        RECT  10.255 33.8525 11.14 33.9175 ;
        RECT  10.83 34.1175 10.895 34.7475 ;
        RECT  11.015 34.4475 11.085 34.5825 ;
        RECT  11.015 34.4475 11.085 34.5825 ;
        RECT  10.395 34.6825 10.465 34.9725 ;
        RECT  10.31 34.4475 10.38 34.5825 ;
        RECT  10.255 35.0575 11.14 35.1225 ;
        RECT  11.015 34.4475 11.085 34.5825 ;
        RECT  11.015 33.9175 11.085 34.1175 ;
        RECT  10.31 33.9175 10.38 34.1175 ;
        RECT  10.935 34.6825 11.005 34.9725 ;
        RECT  10.395 34.6825 10.565 34.7475 ;
        RECT  10.255 35.0575 11.14 35.1225 ;
        RECT  10.255 35.1975 11.14 35.2625 ;
        RECT  10.255 33.8525 11.14 33.9175 ;
        RECT  11.015 36.3425 11.08 36.4775 ;
        RECT  10.83 36.3425 10.895 36.4775 ;
        RECT  10.315 36.3425 10.38 36.4775 ;
        RECT  10.5 36.3425 10.565 36.4775 ;
        RECT  10.83 35.8775 10.895 36.0125 ;
        RECT  11.015 35.8775 11.08 36.0125 ;
        RECT  10.5 35.8775 10.565 36.0125 ;
        RECT  10.315 35.8775 10.38 36.0125 ;
        RECT  10.935 35.4875 11.0 35.6225 ;
        RECT  10.75 35.4875 10.815 35.6225 ;
        RECT  10.58 35.4875 10.645 35.6225 ;
        RECT  10.395 35.4875 10.46 35.6225 ;
        RECT  11.0175 35.98 11.0825 36.115 ;
        RECT  11.0175 35.98 11.0825 36.115 ;
        RECT  11.0175 35.98 11.0825 36.115 ;
        RECT  11.0175 35.98 11.0825 36.115 ;
        RECT  11.0175 35.98 11.0825 36.115 ;
        RECT  11.0175 35.98 11.0825 36.115 ;
        RECT  10.625 36.5425 10.76 36.6075 ;
        RECT  10.2775 35.1975 10.4125 35.2625 ;
        RECT  10.9825 35.1975 11.1175 35.2625 ;
        RECT  10.6125 35.3375 10.7475 35.4025 ;
        RECT  11.0175 35.98 11.0825 36.115 ;
        RECT  11.0175 35.98 11.0825 36.115 ;
        RECT  11.0175 35.98 11.0825 36.115 ;
        RECT  11.0175 35.98 11.0825 36.115 ;
        RECT  10.5175 36.2275 10.6525 36.2925 ;
        RECT  10.5175 36.2275 10.6525 36.2925 ;
        RECT  10.7425 36.0775 10.8775 36.1425 ;
        RECT  10.7425 36.0775 10.8775 36.1425 ;
        RECT  11.0175 35.98 11.0825 36.115 ;
        RECT  11.0175 35.98 11.0825 36.115 ;
        RECT  11.0175 35.98 11.0825 36.115 ;
        RECT  11.0175 35.98 11.0825 36.115 ;
        RECT  10.5675 35.4875 10.6325 35.6225 ;
        RECT  10.3125 35.98 10.3775 36.115 ;
        RECT  10.3125 35.98 10.3775 36.115 ;
        RECT  10.3125 35.98 10.3775 36.115 ;
        RECT  10.3125 35.98 10.3775 36.115 ;
        RECT  10.3125 35.98 10.3775 36.115 ;
        RECT  10.3125 35.98 10.3775 36.115 ;
        RECT  11.0175 35.98 11.0825 36.115 ;
        RECT  11.0175 35.98 11.0825 36.115 ;
        RECT  11.0175 35.98 11.0825 36.115 ;
        RECT  11.0175 35.98 11.0825 36.115 ;
        RECT  10.7625 35.4875 10.8275 35.6225 ;
        RECT  10.63 35.1975 10.765 35.2625 ;
        RECT  10.63 35.1975 10.765 35.2625 ;
        RECT  10.9825 35.1975 11.1175 35.2625 ;
        RECT  10.625 36.5425 10.76 36.6075 ;
        RECT  10.9825 35.1975 11.1175 35.2625 ;
        RECT  10.9825 35.1975 11.1175 35.2625 ;
        RECT  11.0175 35.98 11.0825 36.115 ;
        RECT  11.0175 35.98 11.0825 36.115 ;
        RECT  11.0175 35.98 11.0825 36.115 ;
        RECT  11.0175 35.98 11.0825 36.115 ;
        RECT  11.0175 35.98 11.0825 36.115 ;
        RECT  11.0175 35.98 11.0825 36.115 ;
        RECT  10.2775 35.1975 10.4125 35.2625 ;
        RECT  10.6375 36.5425 10.7375 36.605 ;
        RECT  10.6375 36.545 10.7375 36.6075 ;
        RECT  10.965 35.34 11.0175 35.4025 ;
        RECT  10.6375 36.5425 10.7375 36.605 ;
        RECT  11.015 36.3425 11.085 36.5425 ;
        RECT  11.015 35.8775 11.085 36.0125 ;
        RECT  11.015 35.8775 11.085 36.0125 ;
        RECT  10.255 35.1975 11.14 35.2625 ;
        RECT  10.83 35.7125 11.005 35.7775 ;
        RECT  10.31 35.8775 10.38 36.0125 ;
        RECT  10.5 35.7125 10.565 36.4525 ;
        RECT  10.6375 36.545 10.7375 36.6075 ;
        RECT  10.26 35.34 10.3125 35.4025 ;
        RECT  11.015 35.8775 11.085 36.0125 ;
        RECT  10.255 36.5425 11.14 36.6075 ;
        RECT  10.83 35.7125 10.895 36.3425 ;
        RECT  11.015 35.8775 11.085 36.0125 ;
        RECT  11.015 35.8775 11.085 36.0125 ;
        RECT  10.395 35.4875 10.465 35.7775 ;
        RECT  10.31 35.8775 10.38 36.0125 ;
        RECT  10.255 35.3375 11.14 35.4025 ;
        RECT  11.015 35.8775 11.085 36.0125 ;
        RECT  11.015 36.3425 11.085 36.5425 ;
        RECT  10.31 36.3425 10.38 36.5425 ;
        RECT  10.935 35.4875 11.005 35.7775 ;
        RECT  10.395 35.7125 10.565 35.7775 ;
        RECT  10.255 35.3375 11.14 35.4025 ;
        RECT  10.255 35.1975 11.14 35.2625 ;
        RECT  10.255 36.5425 11.14 36.6075 ;
        RECT  11.015 36.6725 11.08 36.8075 ;
        RECT  10.83 36.6725 10.895 36.8075 ;
        RECT  10.315 36.6725 10.38 36.8075 ;
        RECT  10.5 36.6725 10.565 36.8075 ;
        RECT  10.83 37.1375 10.895 37.2725 ;
        RECT  11.015 37.1375 11.08 37.2725 ;
        RECT  10.5 37.1375 10.565 37.2725 ;
        RECT  10.315 37.1375 10.38 37.2725 ;
        RECT  10.935 37.5275 11.0 37.6625 ;
        RECT  10.75 37.5275 10.815 37.6625 ;
        RECT  10.58 37.5275 10.645 37.6625 ;
        RECT  10.395 37.5275 10.46 37.6625 ;
        RECT  11.0175 37.035 11.0825 37.17 ;
        RECT  11.0175 37.035 11.0825 37.17 ;
        RECT  11.0175 37.035 11.0825 37.17 ;
        RECT  11.0175 37.035 11.0825 37.17 ;
        RECT  11.0175 37.035 11.0825 37.17 ;
        RECT  11.0175 37.035 11.0825 37.17 ;
        RECT  10.625 36.5425 10.76 36.6075 ;
        RECT  10.2775 37.8875 10.4125 37.9525 ;
        RECT  10.9825 37.8875 11.1175 37.9525 ;
        RECT  10.6125 37.7475 10.7475 37.8125 ;
        RECT  11.0175 37.035 11.0825 37.17 ;
        RECT  11.0175 37.035 11.0825 37.17 ;
        RECT  11.0175 37.035 11.0825 37.17 ;
        RECT  11.0175 37.035 11.0825 37.17 ;
        RECT  10.5175 36.8575 10.6525 36.9225 ;
        RECT  10.5175 36.8575 10.6525 36.9225 ;
        RECT  10.7425 37.0075 10.8775 37.0725 ;
        RECT  10.7425 37.0075 10.8775 37.0725 ;
        RECT  11.0175 37.035 11.0825 37.17 ;
        RECT  11.0175 37.035 11.0825 37.17 ;
        RECT  11.0175 37.035 11.0825 37.17 ;
        RECT  11.0175 37.035 11.0825 37.17 ;
        RECT  10.5675 37.5275 10.6325 37.6625 ;
        RECT  10.3125 37.035 10.3775 37.17 ;
        RECT  10.3125 37.035 10.3775 37.17 ;
        RECT  10.3125 37.035 10.3775 37.17 ;
        RECT  10.3125 37.035 10.3775 37.17 ;
        RECT  10.3125 37.035 10.3775 37.17 ;
        RECT  10.3125 37.035 10.3775 37.17 ;
        RECT  11.0175 37.035 11.0825 37.17 ;
        RECT  11.0175 37.035 11.0825 37.17 ;
        RECT  11.0175 37.035 11.0825 37.17 ;
        RECT  11.0175 37.035 11.0825 37.17 ;
        RECT  10.7625 37.5275 10.8275 37.6625 ;
        RECT  10.63 37.8875 10.765 37.9525 ;
        RECT  10.63 37.8875 10.765 37.9525 ;
        RECT  10.9825 37.8875 11.1175 37.9525 ;
        RECT  10.625 36.5425 10.76 36.6075 ;
        RECT  10.9825 37.8875 11.1175 37.9525 ;
        RECT  10.9825 37.8875 11.1175 37.9525 ;
        RECT  11.0175 37.035 11.0825 37.17 ;
        RECT  11.0175 37.035 11.0825 37.17 ;
        RECT  11.0175 37.035 11.0825 37.17 ;
        RECT  11.0175 37.035 11.0825 37.17 ;
        RECT  11.0175 37.035 11.0825 37.17 ;
        RECT  11.0175 37.035 11.0825 37.17 ;
        RECT  10.2775 37.8875 10.4125 37.9525 ;
        RECT  10.6375 36.545 10.7375 36.6075 ;
        RECT  10.6375 36.5425 10.7375 36.605 ;
        RECT  10.965 37.7475 11.0175 37.81 ;
        RECT  10.6375 36.545 10.7375 36.6075 ;
        RECT  11.015 36.6075 11.085 36.8075 ;
        RECT  11.015 37.1375 11.085 37.2725 ;
        RECT  11.015 37.1375 11.085 37.2725 ;
        RECT  10.255 37.8875 11.14 37.9525 ;
        RECT  10.83 37.3725 11.005 37.4375 ;
        RECT  10.31 37.1375 10.38 37.2725 ;
        RECT  10.5 36.6975 10.565 37.4375 ;
        RECT  10.6375 36.5425 10.7375 36.605 ;
        RECT  10.26 37.7475 10.3125 37.81 ;
        RECT  11.015 37.1375 11.085 37.2725 ;
        RECT  10.255 36.5425 11.14 36.6075 ;
        RECT  10.83 36.8075 10.895 37.4375 ;
        RECT  11.015 37.1375 11.085 37.2725 ;
        RECT  11.015 37.1375 11.085 37.2725 ;
        RECT  10.395 37.3725 10.465 37.6625 ;
        RECT  10.31 37.1375 10.38 37.2725 ;
        RECT  10.255 37.7475 11.14 37.8125 ;
        RECT  11.015 37.1375 11.085 37.2725 ;
        RECT  11.015 36.6075 11.085 36.8075 ;
        RECT  10.31 36.6075 10.38 36.8075 ;
        RECT  10.935 37.3725 11.005 37.6625 ;
        RECT  10.395 37.3725 10.565 37.4375 ;
        RECT  10.255 37.7475 11.14 37.8125 ;
        RECT  10.255 37.8875 11.14 37.9525 ;
        RECT  10.255 36.5425 11.14 36.6075 ;
        RECT  11.015 39.0325 11.08 39.1675 ;
        RECT  10.83 39.0325 10.895 39.1675 ;
        RECT  10.315 39.0325 10.38 39.1675 ;
        RECT  10.5 39.0325 10.565 39.1675 ;
        RECT  10.83 38.5675 10.895 38.7025 ;
        RECT  11.015 38.5675 11.08 38.7025 ;
        RECT  10.5 38.5675 10.565 38.7025 ;
        RECT  10.315 38.5675 10.38 38.7025 ;
        RECT  10.935 38.1775 11.0 38.3125 ;
        RECT  10.75 38.1775 10.815 38.3125 ;
        RECT  10.58 38.1775 10.645 38.3125 ;
        RECT  10.395 38.1775 10.46 38.3125 ;
        RECT  11.0175 38.67 11.0825 38.805 ;
        RECT  11.0175 38.67 11.0825 38.805 ;
        RECT  11.0175 38.67 11.0825 38.805 ;
        RECT  11.0175 38.67 11.0825 38.805 ;
        RECT  11.0175 38.67 11.0825 38.805 ;
        RECT  11.0175 38.67 11.0825 38.805 ;
        RECT  10.625 39.2325 10.76 39.2975 ;
        RECT  10.2775 37.8875 10.4125 37.9525 ;
        RECT  10.9825 37.8875 11.1175 37.9525 ;
        RECT  10.6125 38.0275 10.7475 38.0925 ;
        RECT  11.0175 38.67 11.0825 38.805 ;
        RECT  11.0175 38.67 11.0825 38.805 ;
        RECT  11.0175 38.67 11.0825 38.805 ;
        RECT  11.0175 38.67 11.0825 38.805 ;
        RECT  10.5175 38.9175 10.6525 38.9825 ;
        RECT  10.5175 38.9175 10.6525 38.9825 ;
        RECT  10.7425 38.7675 10.8775 38.8325 ;
        RECT  10.7425 38.7675 10.8775 38.8325 ;
        RECT  11.0175 38.67 11.0825 38.805 ;
        RECT  11.0175 38.67 11.0825 38.805 ;
        RECT  11.0175 38.67 11.0825 38.805 ;
        RECT  11.0175 38.67 11.0825 38.805 ;
        RECT  10.5675 38.1775 10.6325 38.3125 ;
        RECT  10.3125 38.67 10.3775 38.805 ;
        RECT  10.3125 38.67 10.3775 38.805 ;
        RECT  10.3125 38.67 10.3775 38.805 ;
        RECT  10.3125 38.67 10.3775 38.805 ;
        RECT  10.3125 38.67 10.3775 38.805 ;
        RECT  10.3125 38.67 10.3775 38.805 ;
        RECT  11.0175 38.67 11.0825 38.805 ;
        RECT  11.0175 38.67 11.0825 38.805 ;
        RECT  11.0175 38.67 11.0825 38.805 ;
        RECT  11.0175 38.67 11.0825 38.805 ;
        RECT  10.7625 38.1775 10.8275 38.3125 ;
        RECT  10.63 37.8875 10.765 37.9525 ;
        RECT  10.63 37.8875 10.765 37.9525 ;
        RECT  10.9825 37.8875 11.1175 37.9525 ;
        RECT  10.625 39.2325 10.76 39.2975 ;
        RECT  10.9825 37.8875 11.1175 37.9525 ;
        RECT  10.9825 37.8875 11.1175 37.9525 ;
        RECT  11.0175 38.67 11.0825 38.805 ;
        RECT  11.0175 38.67 11.0825 38.805 ;
        RECT  11.0175 38.67 11.0825 38.805 ;
        RECT  11.0175 38.67 11.0825 38.805 ;
        RECT  11.0175 38.67 11.0825 38.805 ;
        RECT  11.0175 38.67 11.0825 38.805 ;
        RECT  10.2775 37.8875 10.4125 37.9525 ;
        RECT  10.6375 39.2325 10.7375 39.295 ;
        RECT  10.6375 39.235 10.7375 39.2975 ;
        RECT  10.965 38.03 11.0175 38.0925 ;
        RECT  10.6375 39.2325 10.7375 39.295 ;
        RECT  11.015 39.0325 11.085 39.2325 ;
        RECT  11.015 38.5675 11.085 38.7025 ;
        RECT  11.015 38.5675 11.085 38.7025 ;
        RECT  10.255 37.8875 11.14 37.9525 ;
        RECT  10.83 38.4025 11.005 38.4675 ;
        RECT  10.31 38.5675 10.38 38.7025 ;
        RECT  10.5 38.4025 10.565 39.1425 ;
        RECT  10.6375 39.235 10.7375 39.2975 ;
        RECT  10.26 38.03 10.3125 38.0925 ;
        RECT  11.015 38.5675 11.085 38.7025 ;
        RECT  10.255 39.2325 11.14 39.2975 ;
        RECT  10.83 38.4025 10.895 39.0325 ;
        RECT  11.015 38.5675 11.085 38.7025 ;
        RECT  11.015 38.5675 11.085 38.7025 ;
        RECT  10.395 38.1775 10.465 38.4675 ;
        RECT  10.31 38.5675 10.38 38.7025 ;
        RECT  10.255 38.0275 11.14 38.0925 ;
        RECT  11.015 38.5675 11.085 38.7025 ;
        RECT  11.015 39.0325 11.085 39.2325 ;
        RECT  10.31 39.0325 10.38 39.2325 ;
        RECT  10.935 38.1775 11.005 38.4675 ;
        RECT  10.395 38.4025 10.565 38.4675 ;
        RECT  10.255 38.0275 11.14 38.0925 ;
        RECT  10.255 37.8875 11.14 37.9525 ;
        RECT  10.255 39.2325 11.14 39.2975 ;
        RECT  11.015 39.3625 11.08 39.4975 ;
        RECT  10.83 39.3625 10.895 39.4975 ;
        RECT  10.315 39.3625 10.38 39.4975 ;
        RECT  10.5 39.3625 10.565 39.4975 ;
        RECT  10.83 39.8275 10.895 39.9625 ;
        RECT  11.015 39.8275 11.08 39.9625 ;
        RECT  10.5 39.8275 10.565 39.9625 ;
        RECT  10.315 39.8275 10.38 39.9625 ;
        RECT  10.935 40.2175 11.0 40.3525 ;
        RECT  10.75 40.2175 10.815 40.3525 ;
        RECT  10.58 40.2175 10.645 40.3525 ;
        RECT  10.395 40.2175 10.46 40.3525 ;
        RECT  11.0175 39.725 11.0825 39.86 ;
        RECT  11.0175 39.725 11.0825 39.86 ;
        RECT  11.0175 39.725 11.0825 39.86 ;
        RECT  11.0175 39.725 11.0825 39.86 ;
        RECT  11.0175 39.725 11.0825 39.86 ;
        RECT  11.0175 39.725 11.0825 39.86 ;
        RECT  10.625 39.2325 10.76 39.2975 ;
        RECT  10.2775 40.5775 10.4125 40.6425 ;
        RECT  10.9825 40.5775 11.1175 40.6425 ;
        RECT  10.6125 40.4375 10.7475 40.5025 ;
        RECT  11.0175 39.725 11.0825 39.86 ;
        RECT  11.0175 39.725 11.0825 39.86 ;
        RECT  11.0175 39.725 11.0825 39.86 ;
        RECT  11.0175 39.725 11.0825 39.86 ;
        RECT  10.5175 39.5475 10.6525 39.6125 ;
        RECT  10.5175 39.5475 10.6525 39.6125 ;
        RECT  10.7425 39.6975 10.8775 39.7625 ;
        RECT  10.7425 39.6975 10.8775 39.7625 ;
        RECT  11.0175 39.725 11.0825 39.86 ;
        RECT  11.0175 39.725 11.0825 39.86 ;
        RECT  11.0175 39.725 11.0825 39.86 ;
        RECT  11.0175 39.725 11.0825 39.86 ;
        RECT  10.5675 40.2175 10.6325 40.3525 ;
        RECT  10.3125 39.725 10.3775 39.86 ;
        RECT  10.3125 39.725 10.3775 39.86 ;
        RECT  10.3125 39.725 10.3775 39.86 ;
        RECT  10.3125 39.725 10.3775 39.86 ;
        RECT  10.3125 39.725 10.3775 39.86 ;
        RECT  10.3125 39.725 10.3775 39.86 ;
        RECT  11.0175 39.725 11.0825 39.86 ;
        RECT  11.0175 39.725 11.0825 39.86 ;
        RECT  11.0175 39.725 11.0825 39.86 ;
        RECT  11.0175 39.725 11.0825 39.86 ;
        RECT  10.7625 40.2175 10.8275 40.3525 ;
        RECT  10.63 40.5775 10.765 40.6425 ;
        RECT  10.63 40.5775 10.765 40.6425 ;
        RECT  10.9825 40.5775 11.1175 40.6425 ;
        RECT  10.625 39.2325 10.76 39.2975 ;
        RECT  10.9825 40.5775 11.1175 40.6425 ;
        RECT  10.9825 40.5775 11.1175 40.6425 ;
        RECT  11.0175 39.725 11.0825 39.86 ;
        RECT  11.0175 39.725 11.0825 39.86 ;
        RECT  11.0175 39.725 11.0825 39.86 ;
        RECT  11.0175 39.725 11.0825 39.86 ;
        RECT  11.0175 39.725 11.0825 39.86 ;
        RECT  11.0175 39.725 11.0825 39.86 ;
        RECT  10.2775 40.5775 10.4125 40.6425 ;
        RECT  10.6375 39.235 10.7375 39.2975 ;
        RECT  10.6375 39.2325 10.7375 39.295 ;
        RECT  10.965 40.4375 11.0175 40.5 ;
        RECT  10.6375 39.235 10.7375 39.2975 ;
        RECT  11.015 39.2975 11.085 39.4975 ;
        RECT  11.015 39.8275 11.085 39.9625 ;
        RECT  11.015 39.8275 11.085 39.9625 ;
        RECT  10.255 40.5775 11.14 40.6425 ;
        RECT  10.83 40.0625 11.005 40.1275 ;
        RECT  10.31 39.8275 10.38 39.9625 ;
        RECT  10.5 39.3875 10.565 40.1275 ;
        RECT  10.6375 39.2325 10.7375 39.295 ;
        RECT  10.26 40.4375 10.3125 40.5 ;
        RECT  11.015 39.8275 11.085 39.9625 ;
        RECT  10.255 39.2325 11.14 39.2975 ;
        RECT  10.83 39.4975 10.895 40.1275 ;
        RECT  11.015 39.8275 11.085 39.9625 ;
        RECT  11.015 39.8275 11.085 39.9625 ;
        RECT  10.395 40.0625 10.465 40.3525 ;
        RECT  10.31 39.8275 10.38 39.9625 ;
        RECT  10.255 40.4375 11.14 40.5025 ;
        RECT  11.015 39.8275 11.085 39.9625 ;
        RECT  11.015 39.2975 11.085 39.4975 ;
        RECT  10.31 39.2975 10.38 39.4975 ;
        RECT  10.935 40.0625 11.005 40.3525 ;
        RECT  10.395 40.0625 10.565 40.1275 ;
        RECT  10.255 40.4375 11.14 40.5025 ;
        RECT  10.255 40.5775 11.14 40.6425 ;
        RECT  10.255 39.2325 11.14 39.2975 ;
        RECT  11.72 20.2025 11.785 20.3375 ;
        RECT  11.535 20.2025 11.6 20.3375 ;
        RECT  11.02 20.2025 11.085 20.3375 ;
        RECT  11.205 20.2025 11.27 20.3375 ;
        RECT  11.535 19.7375 11.6 19.8725 ;
        RECT  11.72 19.7375 11.785 19.8725 ;
        RECT  11.205 19.7375 11.27 19.8725 ;
        RECT  11.02 19.7375 11.085 19.8725 ;
        RECT  11.64 19.3475 11.705 19.4825 ;
        RECT  11.455 19.3475 11.52 19.4825 ;
        RECT  11.285 19.3475 11.35 19.4825 ;
        RECT  11.1 19.3475 11.165 19.4825 ;
        RECT  11.7225 19.84 11.7875 19.975 ;
        RECT  11.7225 19.84 11.7875 19.975 ;
        RECT  11.7225 19.84 11.7875 19.975 ;
        RECT  11.7225 19.84 11.7875 19.975 ;
        RECT  11.7225 19.84 11.7875 19.975 ;
        RECT  11.7225 19.84 11.7875 19.975 ;
        RECT  11.33 20.4025 11.465 20.4675 ;
        RECT  10.9825 19.0575 11.1175 19.1225 ;
        RECT  11.6875 19.0575 11.8225 19.1225 ;
        RECT  11.3175 19.1975 11.4525 19.2625 ;
        RECT  11.7225 19.84 11.7875 19.975 ;
        RECT  11.7225 19.84 11.7875 19.975 ;
        RECT  11.7225 19.84 11.7875 19.975 ;
        RECT  11.7225 19.84 11.7875 19.975 ;
        RECT  11.2225 20.0875 11.3575 20.1525 ;
        RECT  11.2225 20.0875 11.3575 20.1525 ;
        RECT  11.4475 19.9375 11.5825 20.0025 ;
        RECT  11.4475 19.9375 11.5825 20.0025 ;
        RECT  11.7225 19.84 11.7875 19.975 ;
        RECT  11.7225 19.84 11.7875 19.975 ;
        RECT  11.7225 19.84 11.7875 19.975 ;
        RECT  11.7225 19.84 11.7875 19.975 ;
        RECT  11.2725 19.3475 11.3375 19.4825 ;
        RECT  11.0175 19.84 11.0825 19.975 ;
        RECT  11.0175 19.84 11.0825 19.975 ;
        RECT  11.0175 19.84 11.0825 19.975 ;
        RECT  11.0175 19.84 11.0825 19.975 ;
        RECT  11.0175 19.84 11.0825 19.975 ;
        RECT  11.0175 19.84 11.0825 19.975 ;
        RECT  11.7225 19.84 11.7875 19.975 ;
        RECT  11.7225 19.84 11.7875 19.975 ;
        RECT  11.7225 19.84 11.7875 19.975 ;
        RECT  11.7225 19.84 11.7875 19.975 ;
        RECT  11.4675 19.3475 11.5325 19.4825 ;
        RECT  11.335 19.0575 11.47 19.1225 ;
        RECT  11.335 19.0575 11.47 19.1225 ;
        RECT  11.6875 19.0575 11.8225 19.1225 ;
        RECT  11.33 20.4025 11.465 20.4675 ;
        RECT  11.6875 19.0575 11.8225 19.1225 ;
        RECT  11.6875 19.0575 11.8225 19.1225 ;
        RECT  11.7225 19.84 11.7875 19.975 ;
        RECT  11.7225 19.84 11.7875 19.975 ;
        RECT  11.7225 19.84 11.7875 19.975 ;
        RECT  11.7225 19.84 11.7875 19.975 ;
        RECT  11.7225 19.84 11.7875 19.975 ;
        RECT  11.7225 19.84 11.7875 19.975 ;
        RECT  10.9825 19.0575 11.1175 19.1225 ;
        RECT  11.3425 20.4025 11.4425 20.465 ;
        RECT  11.3425 20.405 11.4425 20.4675 ;
        RECT  11.67 19.2 11.7225 19.2625 ;
        RECT  11.3425 20.4025 11.4425 20.465 ;
        RECT  11.72 20.2025 11.79 20.4025 ;
        RECT  11.72 19.7375 11.79 19.8725 ;
        RECT  11.72 19.7375 11.79 19.8725 ;
        RECT  10.96 19.0575 11.845 19.1225 ;
        RECT  11.535 19.5725 11.71 19.6375 ;
        RECT  11.015 19.7375 11.085 19.8725 ;
        RECT  11.205 19.5725 11.27 20.3125 ;
        RECT  11.3425 20.405 11.4425 20.4675 ;
        RECT  10.965 19.2 11.0175 19.2625 ;
        RECT  11.72 19.7375 11.79 19.8725 ;
        RECT  10.96 20.4025 11.845 20.4675 ;
        RECT  11.535 19.5725 11.6 20.2025 ;
        RECT  11.72 19.7375 11.79 19.8725 ;
        RECT  11.72 19.7375 11.79 19.8725 ;
        RECT  11.1 19.3475 11.17 19.6375 ;
        RECT  11.015 19.7375 11.085 19.8725 ;
        RECT  10.96 19.1975 11.845 19.2625 ;
        RECT  11.72 19.7375 11.79 19.8725 ;
        RECT  11.72 20.2025 11.79 20.4025 ;
        RECT  11.015 20.2025 11.085 20.4025 ;
        RECT  11.64 19.3475 11.71 19.6375 ;
        RECT  11.1 19.5725 11.27 19.6375 ;
        RECT  10.96 19.1975 11.845 19.2625 ;
        RECT  10.96 19.0575 11.845 19.1225 ;
        RECT  10.96 20.4025 11.845 20.4675 ;
        RECT  11.72 20.5325 11.785 20.6675 ;
        RECT  11.535 20.5325 11.6 20.6675 ;
        RECT  11.02 20.5325 11.085 20.6675 ;
        RECT  11.205 20.5325 11.27 20.6675 ;
        RECT  11.535 20.9975 11.6 21.1325 ;
        RECT  11.72 20.9975 11.785 21.1325 ;
        RECT  11.205 20.9975 11.27 21.1325 ;
        RECT  11.02 20.9975 11.085 21.1325 ;
        RECT  11.64 21.3875 11.705 21.5225 ;
        RECT  11.455 21.3875 11.52 21.5225 ;
        RECT  11.285 21.3875 11.35 21.5225 ;
        RECT  11.1 21.3875 11.165 21.5225 ;
        RECT  11.7225 20.895 11.7875 21.03 ;
        RECT  11.7225 20.895 11.7875 21.03 ;
        RECT  11.7225 20.895 11.7875 21.03 ;
        RECT  11.7225 20.895 11.7875 21.03 ;
        RECT  11.7225 20.895 11.7875 21.03 ;
        RECT  11.7225 20.895 11.7875 21.03 ;
        RECT  11.33 20.4025 11.465 20.4675 ;
        RECT  10.9825 21.7475 11.1175 21.8125 ;
        RECT  11.6875 21.7475 11.8225 21.8125 ;
        RECT  11.3175 21.6075 11.4525 21.6725 ;
        RECT  11.7225 20.895 11.7875 21.03 ;
        RECT  11.7225 20.895 11.7875 21.03 ;
        RECT  11.7225 20.895 11.7875 21.03 ;
        RECT  11.7225 20.895 11.7875 21.03 ;
        RECT  11.2225 20.7175 11.3575 20.7825 ;
        RECT  11.2225 20.7175 11.3575 20.7825 ;
        RECT  11.4475 20.8675 11.5825 20.9325 ;
        RECT  11.4475 20.8675 11.5825 20.9325 ;
        RECT  11.7225 20.895 11.7875 21.03 ;
        RECT  11.7225 20.895 11.7875 21.03 ;
        RECT  11.7225 20.895 11.7875 21.03 ;
        RECT  11.7225 20.895 11.7875 21.03 ;
        RECT  11.2725 21.3875 11.3375 21.5225 ;
        RECT  11.0175 20.895 11.0825 21.03 ;
        RECT  11.0175 20.895 11.0825 21.03 ;
        RECT  11.0175 20.895 11.0825 21.03 ;
        RECT  11.0175 20.895 11.0825 21.03 ;
        RECT  11.0175 20.895 11.0825 21.03 ;
        RECT  11.0175 20.895 11.0825 21.03 ;
        RECT  11.7225 20.895 11.7875 21.03 ;
        RECT  11.7225 20.895 11.7875 21.03 ;
        RECT  11.7225 20.895 11.7875 21.03 ;
        RECT  11.7225 20.895 11.7875 21.03 ;
        RECT  11.4675 21.3875 11.5325 21.5225 ;
        RECT  11.335 21.7475 11.47 21.8125 ;
        RECT  11.335 21.7475 11.47 21.8125 ;
        RECT  11.6875 21.7475 11.8225 21.8125 ;
        RECT  11.33 20.4025 11.465 20.4675 ;
        RECT  11.6875 21.7475 11.8225 21.8125 ;
        RECT  11.6875 21.7475 11.8225 21.8125 ;
        RECT  11.7225 20.895 11.7875 21.03 ;
        RECT  11.7225 20.895 11.7875 21.03 ;
        RECT  11.7225 20.895 11.7875 21.03 ;
        RECT  11.7225 20.895 11.7875 21.03 ;
        RECT  11.7225 20.895 11.7875 21.03 ;
        RECT  11.7225 20.895 11.7875 21.03 ;
        RECT  10.9825 21.7475 11.1175 21.8125 ;
        RECT  11.3425 20.405 11.4425 20.4675 ;
        RECT  11.3425 20.4025 11.4425 20.465 ;
        RECT  11.67 21.6075 11.7225 21.67 ;
        RECT  11.3425 20.405 11.4425 20.4675 ;
        RECT  11.72 20.4675 11.79 20.6675 ;
        RECT  11.72 20.9975 11.79 21.1325 ;
        RECT  11.72 20.9975 11.79 21.1325 ;
        RECT  10.96 21.7475 11.845 21.8125 ;
        RECT  11.535 21.2325 11.71 21.2975 ;
        RECT  11.015 20.9975 11.085 21.1325 ;
        RECT  11.205 20.5575 11.27 21.2975 ;
        RECT  11.3425 20.4025 11.4425 20.465 ;
        RECT  10.965 21.6075 11.0175 21.67 ;
        RECT  11.72 20.9975 11.79 21.1325 ;
        RECT  10.96 20.4025 11.845 20.4675 ;
        RECT  11.535 20.6675 11.6 21.2975 ;
        RECT  11.72 20.9975 11.79 21.1325 ;
        RECT  11.72 20.9975 11.79 21.1325 ;
        RECT  11.1 21.2325 11.17 21.5225 ;
        RECT  11.015 20.9975 11.085 21.1325 ;
        RECT  10.96 21.6075 11.845 21.6725 ;
        RECT  11.72 20.9975 11.79 21.1325 ;
        RECT  11.72 20.4675 11.79 20.6675 ;
        RECT  11.015 20.4675 11.085 20.6675 ;
        RECT  11.64 21.2325 11.71 21.5225 ;
        RECT  11.1 21.2325 11.27 21.2975 ;
        RECT  10.96 21.6075 11.845 21.6725 ;
        RECT  10.96 21.7475 11.845 21.8125 ;
        RECT  10.96 20.4025 11.845 20.4675 ;
        RECT  11.72 22.8925 11.785 23.0275 ;
        RECT  11.535 22.8925 11.6 23.0275 ;
        RECT  11.02 22.8925 11.085 23.0275 ;
        RECT  11.205 22.8925 11.27 23.0275 ;
        RECT  11.535 22.4275 11.6 22.5625 ;
        RECT  11.72 22.4275 11.785 22.5625 ;
        RECT  11.205 22.4275 11.27 22.5625 ;
        RECT  11.02 22.4275 11.085 22.5625 ;
        RECT  11.64 22.0375 11.705 22.1725 ;
        RECT  11.455 22.0375 11.52 22.1725 ;
        RECT  11.285 22.0375 11.35 22.1725 ;
        RECT  11.1 22.0375 11.165 22.1725 ;
        RECT  11.7225 22.53 11.7875 22.665 ;
        RECT  11.7225 22.53 11.7875 22.665 ;
        RECT  11.7225 22.53 11.7875 22.665 ;
        RECT  11.7225 22.53 11.7875 22.665 ;
        RECT  11.7225 22.53 11.7875 22.665 ;
        RECT  11.7225 22.53 11.7875 22.665 ;
        RECT  11.33 23.0925 11.465 23.1575 ;
        RECT  10.9825 21.7475 11.1175 21.8125 ;
        RECT  11.6875 21.7475 11.8225 21.8125 ;
        RECT  11.3175 21.8875 11.4525 21.9525 ;
        RECT  11.7225 22.53 11.7875 22.665 ;
        RECT  11.7225 22.53 11.7875 22.665 ;
        RECT  11.7225 22.53 11.7875 22.665 ;
        RECT  11.7225 22.53 11.7875 22.665 ;
        RECT  11.2225 22.7775 11.3575 22.8425 ;
        RECT  11.2225 22.7775 11.3575 22.8425 ;
        RECT  11.4475 22.6275 11.5825 22.6925 ;
        RECT  11.4475 22.6275 11.5825 22.6925 ;
        RECT  11.7225 22.53 11.7875 22.665 ;
        RECT  11.7225 22.53 11.7875 22.665 ;
        RECT  11.7225 22.53 11.7875 22.665 ;
        RECT  11.7225 22.53 11.7875 22.665 ;
        RECT  11.2725 22.0375 11.3375 22.1725 ;
        RECT  11.0175 22.53 11.0825 22.665 ;
        RECT  11.0175 22.53 11.0825 22.665 ;
        RECT  11.0175 22.53 11.0825 22.665 ;
        RECT  11.0175 22.53 11.0825 22.665 ;
        RECT  11.0175 22.53 11.0825 22.665 ;
        RECT  11.0175 22.53 11.0825 22.665 ;
        RECT  11.7225 22.53 11.7875 22.665 ;
        RECT  11.7225 22.53 11.7875 22.665 ;
        RECT  11.7225 22.53 11.7875 22.665 ;
        RECT  11.7225 22.53 11.7875 22.665 ;
        RECT  11.4675 22.0375 11.5325 22.1725 ;
        RECT  11.335 21.7475 11.47 21.8125 ;
        RECT  11.335 21.7475 11.47 21.8125 ;
        RECT  11.6875 21.7475 11.8225 21.8125 ;
        RECT  11.33 23.0925 11.465 23.1575 ;
        RECT  11.6875 21.7475 11.8225 21.8125 ;
        RECT  11.6875 21.7475 11.8225 21.8125 ;
        RECT  11.7225 22.53 11.7875 22.665 ;
        RECT  11.7225 22.53 11.7875 22.665 ;
        RECT  11.7225 22.53 11.7875 22.665 ;
        RECT  11.7225 22.53 11.7875 22.665 ;
        RECT  11.7225 22.53 11.7875 22.665 ;
        RECT  11.7225 22.53 11.7875 22.665 ;
        RECT  10.9825 21.7475 11.1175 21.8125 ;
        RECT  11.3425 23.0925 11.4425 23.155 ;
        RECT  11.3425 23.095 11.4425 23.1575 ;
        RECT  11.67 21.89 11.7225 21.9525 ;
        RECT  11.3425 23.0925 11.4425 23.155 ;
        RECT  11.72 22.8925 11.79 23.0925 ;
        RECT  11.72 22.4275 11.79 22.5625 ;
        RECT  11.72 22.4275 11.79 22.5625 ;
        RECT  10.96 21.7475 11.845 21.8125 ;
        RECT  11.535 22.2625 11.71 22.3275 ;
        RECT  11.015 22.4275 11.085 22.5625 ;
        RECT  11.205 22.2625 11.27 23.0025 ;
        RECT  11.3425 23.095 11.4425 23.1575 ;
        RECT  10.965 21.89 11.0175 21.9525 ;
        RECT  11.72 22.4275 11.79 22.5625 ;
        RECT  10.96 23.0925 11.845 23.1575 ;
        RECT  11.535 22.2625 11.6 22.8925 ;
        RECT  11.72 22.4275 11.79 22.5625 ;
        RECT  11.72 22.4275 11.79 22.5625 ;
        RECT  11.1 22.0375 11.17 22.3275 ;
        RECT  11.015 22.4275 11.085 22.5625 ;
        RECT  10.96 21.8875 11.845 21.9525 ;
        RECT  11.72 22.4275 11.79 22.5625 ;
        RECT  11.72 22.8925 11.79 23.0925 ;
        RECT  11.015 22.8925 11.085 23.0925 ;
        RECT  11.64 22.0375 11.71 22.3275 ;
        RECT  11.1 22.2625 11.27 22.3275 ;
        RECT  10.96 21.8875 11.845 21.9525 ;
        RECT  10.96 21.7475 11.845 21.8125 ;
        RECT  10.96 23.0925 11.845 23.1575 ;
        RECT  11.72 23.2225 11.785 23.3575 ;
        RECT  11.535 23.2225 11.6 23.3575 ;
        RECT  11.02 23.2225 11.085 23.3575 ;
        RECT  11.205 23.2225 11.27 23.3575 ;
        RECT  11.535 23.6875 11.6 23.8225 ;
        RECT  11.72 23.6875 11.785 23.8225 ;
        RECT  11.205 23.6875 11.27 23.8225 ;
        RECT  11.02 23.6875 11.085 23.8225 ;
        RECT  11.64 24.0775 11.705 24.2125 ;
        RECT  11.455 24.0775 11.52 24.2125 ;
        RECT  11.285 24.0775 11.35 24.2125 ;
        RECT  11.1 24.0775 11.165 24.2125 ;
        RECT  11.7225 23.585 11.7875 23.72 ;
        RECT  11.7225 23.585 11.7875 23.72 ;
        RECT  11.7225 23.585 11.7875 23.72 ;
        RECT  11.7225 23.585 11.7875 23.72 ;
        RECT  11.7225 23.585 11.7875 23.72 ;
        RECT  11.7225 23.585 11.7875 23.72 ;
        RECT  11.33 23.0925 11.465 23.1575 ;
        RECT  10.9825 24.4375 11.1175 24.5025 ;
        RECT  11.6875 24.4375 11.8225 24.5025 ;
        RECT  11.3175 24.2975 11.4525 24.3625 ;
        RECT  11.7225 23.585 11.7875 23.72 ;
        RECT  11.7225 23.585 11.7875 23.72 ;
        RECT  11.7225 23.585 11.7875 23.72 ;
        RECT  11.7225 23.585 11.7875 23.72 ;
        RECT  11.2225 23.4075 11.3575 23.4725 ;
        RECT  11.2225 23.4075 11.3575 23.4725 ;
        RECT  11.4475 23.5575 11.5825 23.6225 ;
        RECT  11.4475 23.5575 11.5825 23.6225 ;
        RECT  11.7225 23.585 11.7875 23.72 ;
        RECT  11.7225 23.585 11.7875 23.72 ;
        RECT  11.7225 23.585 11.7875 23.72 ;
        RECT  11.7225 23.585 11.7875 23.72 ;
        RECT  11.2725 24.0775 11.3375 24.2125 ;
        RECT  11.0175 23.585 11.0825 23.72 ;
        RECT  11.0175 23.585 11.0825 23.72 ;
        RECT  11.0175 23.585 11.0825 23.72 ;
        RECT  11.0175 23.585 11.0825 23.72 ;
        RECT  11.0175 23.585 11.0825 23.72 ;
        RECT  11.0175 23.585 11.0825 23.72 ;
        RECT  11.7225 23.585 11.7875 23.72 ;
        RECT  11.7225 23.585 11.7875 23.72 ;
        RECT  11.7225 23.585 11.7875 23.72 ;
        RECT  11.7225 23.585 11.7875 23.72 ;
        RECT  11.4675 24.0775 11.5325 24.2125 ;
        RECT  11.335 24.4375 11.47 24.5025 ;
        RECT  11.335 24.4375 11.47 24.5025 ;
        RECT  11.6875 24.4375 11.8225 24.5025 ;
        RECT  11.33 23.0925 11.465 23.1575 ;
        RECT  11.6875 24.4375 11.8225 24.5025 ;
        RECT  11.6875 24.4375 11.8225 24.5025 ;
        RECT  11.7225 23.585 11.7875 23.72 ;
        RECT  11.7225 23.585 11.7875 23.72 ;
        RECT  11.7225 23.585 11.7875 23.72 ;
        RECT  11.7225 23.585 11.7875 23.72 ;
        RECT  11.7225 23.585 11.7875 23.72 ;
        RECT  11.7225 23.585 11.7875 23.72 ;
        RECT  10.9825 24.4375 11.1175 24.5025 ;
        RECT  11.3425 23.095 11.4425 23.1575 ;
        RECT  11.3425 23.0925 11.4425 23.155 ;
        RECT  11.67 24.2975 11.7225 24.36 ;
        RECT  11.3425 23.095 11.4425 23.1575 ;
        RECT  11.72 23.1575 11.79 23.3575 ;
        RECT  11.72 23.6875 11.79 23.8225 ;
        RECT  11.72 23.6875 11.79 23.8225 ;
        RECT  10.96 24.4375 11.845 24.5025 ;
        RECT  11.535 23.9225 11.71 23.9875 ;
        RECT  11.015 23.6875 11.085 23.8225 ;
        RECT  11.205 23.2475 11.27 23.9875 ;
        RECT  11.3425 23.0925 11.4425 23.155 ;
        RECT  10.965 24.2975 11.0175 24.36 ;
        RECT  11.72 23.6875 11.79 23.8225 ;
        RECT  10.96 23.0925 11.845 23.1575 ;
        RECT  11.535 23.3575 11.6 23.9875 ;
        RECT  11.72 23.6875 11.79 23.8225 ;
        RECT  11.72 23.6875 11.79 23.8225 ;
        RECT  11.1 23.9225 11.17 24.2125 ;
        RECT  11.015 23.6875 11.085 23.8225 ;
        RECT  10.96 24.2975 11.845 24.3625 ;
        RECT  11.72 23.6875 11.79 23.8225 ;
        RECT  11.72 23.1575 11.79 23.3575 ;
        RECT  11.015 23.1575 11.085 23.3575 ;
        RECT  11.64 23.9225 11.71 24.2125 ;
        RECT  11.1 23.9225 11.27 23.9875 ;
        RECT  10.96 24.2975 11.845 24.3625 ;
        RECT  10.96 24.4375 11.845 24.5025 ;
        RECT  10.96 23.0925 11.845 23.1575 ;
        RECT  11.72 25.5825 11.785 25.7175 ;
        RECT  11.535 25.5825 11.6 25.7175 ;
        RECT  11.02 25.5825 11.085 25.7175 ;
        RECT  11.205 25.5825 11.27 25.7175 ;
        RECT  11.535 25.1175 11.6 25.2525 ;
        RECT  11.72 25.1175 11.785 25.2525 ;
        RECT  11.205 25.1175 11.27 25.2525 ;
        RECT  11.02 25.1175 11.085 25.2525 ;
        RECT  11.64 24.7275 11.705 24.8625 ;
        RECT  11.455 24.7275 11.52 24.8625 ;
        RECT  11.285 24.7275 11.35 24.8625 ;
        RECT  11.1 24.7275 11.165 24.8625 ;
        RECT  11.7225 25.22 11.7875 25.355 ;
        RECT  11.7225 25.22 11.7875 25.355 ;
        RECT  11.7225 25.22 11.7875 25.355 ;
        RECT  11.7225 25.22 11.7875 25.355 ;
        RECT  11.7225 25.22 11.7875 25.355 ;
        RECT  11.7225 25.22 11.7875 25.355 ;
        RECT  11.33 25.7825 11.465 25.8475 ;
        RECT  10.9825 24.4375 11.1175 24.5025 ;
        RECT  11.6875 24.4375 11.8225 24.5025 ;
        RECT  11.3175 24.5775 11.4525 24.6425 ;
        RECT  11.7225 25.22 11.7875 25.355 ;
        RECT  11.7225 25.22 11.7875 25.355 ;
        RECT  11.7225 25.22 11.7875 25.355 ;
        RECT  11.7225 25.22 11.7875 25.355 ;
        RECT  11.2225 25.4675 11.3575 25.5325 ;
        RECT  11.2225 25.4675 11.3575 25.5325 ;
        RECT  11.4475 25.3175 11.5825 25.3825 ;
        RECT  11.4475 25.3175 11.5825 25.3825 ;
        RECT  11.7225 25.22 11.7875 25.355 ;
        RECT  11.7225 25.22 11.7875 25.355 ;
        RECT  11.7225 25.22 11.7875 25.355 ;
        RECT  11.7225 25.22 11.7875 25.355 ;
        RECT  11.2725 24.7275 11.3375 24.8625 ;
        RECT  11.0175 25.22 11.0825 25.355 ;
        RECT  11.0175 25.22 11.0825 25.355 ;
        RECT  11.0175 25.22 11.0825 25.355 ;
        RECT  11.0175 25.22 11.0825 25.355 ;
        RECT  11.0175 25.22 11.0825 25.355 ;
        RECT  11.0175 25.22 11.0825 25.355 ;
        RECT  11.7225 25.22 11.7875 25.355 ;
        RECT  11.7225 25.22 11.7875 25.355 ;
        RECT  11.7225 25.22 11.7875 25.355 ;
        RECT  11.7225 25.22 11.7875 25.355 ;
        RECT  11.4675 24.7275 11.5325 24.8625 ;
        RECT  11.335 24.4375 11.47 24.5025 ;
        RECT  11.335 24.4375 11.47 24.5025 ;
        RECT  11.6875 24.4375 11.8225 24.5025 ;
        RECT  11.33 25.7825 11.465 25.8475 ;
        RECT  11.6875 24.4375 11.8225 24.5025 ;
        RECT  11.6875 24.4375 11.8225 24.5025 ;
        RECT  11.7225 25.22 11.7875 25.355 ;
        RECT  11.7225 25.22 11.7875 25.355 ;
        RECT  11.7225 25.22 11.7875 25.355 ;
        RECT  11.7225 25.22 11.7875 25.355 ;
        RECT  11.7225 25.22 11.7875 25.355 ;
        RECT  11.7225 25.22 11.7875 25.355 ;
        RECT  10.9825 24.4375 11.1175 24.5025 ;
        RECT  11.3425 25.7825 11.4425 25.845 ;
        RECT  11.3425 25.785 11.4425 25.8475 ;
        RECT  11.67 24.58 11.7225 24.6425 ;
        RECT  11.3425 25.7825 11.4425 25.845 ;
        RECT  11.72 25.5825 11.79 25.7825 ;
        RECT  11.72 25.1175 11.79 25.2525 ;
        RECT  11.72 25.1175 11.79 25.2525 ;
        RECT  10.96 24.4375 11.845 24.5025 ;
        RECT  11.535 24.9525 11.71 25.0175 ;
        RECT  11.015 25.1175 11.085 25.2525 ;
        RECT  11.205 24.9525 11.27 25.6925 ;
        RECT  11.3425 25.785 11.4425 25.8475 ;
        RECT  10.965 24.58 11.0175 24.6425 ;
        RECT  11.72 25.1175 11.79 25.2525 ;
        RECT  10.96 25.7825 11.845 25.8475 ;
        RECT  11.535 24.9525 11.6 25.5825 ;
        RECT  11.72 25.1175 11.79 25.2525 ;
        RECT  11.72 25.1175 11.79 25.2525 ;
        RECT  11.1 24.7275 11.17 25.0175 ;
        RECT  11.015 25.1175 11.085 25.2525 ;
        RECT  10.96 24.5775 11.845 24.6425 ;
        RECT  11.72 25.1175 11.79 25.2525 ;
        RECT  11.72 25.5825 11.79 25.7825 ;
        RECT  11.015 25.5825 11.085 25.7825 ;
        RECT  11.64 24.7275 11.71 25.0175 ;
        RECT  11.1 24.9525 11.27 25.0175 ;
        RECT  10.96 24.5775 11.845 24.6425 ;
        RECT  10.96 24.4375 11.845 24.5025 ;
        RECT  10.96 25.7825 11.845 25.8475 ;
        RECT  11.72 25.9125 11.785 26.0475 ;
        RECT  11.535 25.9125 11.6 26.0475 ;
        RECT  11.02 25.9125 11.085 26.0475 ;
        RECT  11.205 25.9125 11.27 26.0475 ;
        RECT  11.535 26.3775 11.6 26.5125 ;
        RECT  11.72 26.3775 11.785 26.5125 ;
        RECT  11.205 26.3775 11.27 26.5125 ;
        RECT  11.02 26.3775 11.085 26.5125 ;
        RECT  11.64 26.7675 11.705 26.9025 ;
        RECT  11.455 26.7675 11.52 26.9025 ;
        RECT  11.285 26.7675 11.35 26.9025 ;
        RECT  11.1 26.7675 11.165 26.9025 ;
        RECT  11.7225 26.275 11.7875 26.41 ;
        RECT  11.7225 26.275 11.7875 26.41 ;
        RECT  11.7225 26.275 11.7875 26.41 ;
        RECT  11.7225 26.275 11.7875 26.41 ;
        RECT  11.7225 26.275 11.7875 26.41 ;
        RECT  11.7225 26.275 11.7875 26.41 ;
        RECT  11.33 25.7825 11.465 25.8475 ;
        RECT  10.9825 27.1275 11.1175 27.1925 ;
        RECT  11.6875 27.1275 11.8225 27.1925 ;
        RECT  11.3175 26.9875 11.4525 27.0525 ;
        RECT  11.7225 26.275 11.7875 26.41 ;
        RECT  11.7225 26.275 11.7875 26.41 ;
        RECT  11.7225 26.275 11.7875 26.41 ;
        RECT  11.7225 26.275 11.7875 26.41 ;
        RECT  11.2225 26.0975 11.3575 26.1625 ;
        RECT  11.2225 26.0975 11.3575 26.1625 ;
        RECT  11.4475 26.2475 11.5825 26.3125 ;
        RECT  11.4475 26.2475 11.5825 26.3125 ;
        RECT  11.7225 26.275 11.7875 26.41 ;
        RECT  11.7225 26.275 11.7875 26.41 ;
        RECT  11.7225 26.275 11.7875 26.41 ;
        RECT  11.7225 26.275 11.7875 26.41 ;
        RECT  11.2725 26.7675 11.3375 26.9025 ;
        RECT  11.0175 26.275 11.0825 26.41 ;
        RECT  11.0175 26.275 11.0825 26.41 ;
        RECT  11.0175 26.275 11.0825 26.41 ;
        RECT  11.0175 26.275 11.0825 26.41 ;
        RECT  11.0175 26.275 11.0825 26.41 ;
        RECT  11.0175 26.275 11.0825 26.41 ;
        RECT  11.7225 26.275 11.7875 26.41 ;
        RECT  11.7225 26.275 11.7875 26.41 ;
        RECT  11.7225 26.275 11.7875 26.41 ;
        RECT  11.7225 26.275 11.7875 26.41 ;
        RECT  11.4675 26.7675 11.5325 26.9025 ;
        RECT  11.335 27.1275 11.47 27.1925 ;
        RECT  11.335 27.1275 11.47 27.1925 ;
        RECT  11.6875 27.1275 11.8225 27.1925 ;
        RECT  11.33 25.7825 11.465 25.8475 ;
        RECT  11.6875 27.1275 11.8225 27.1925 ;
        RECT  11.6875 27.1275 11.8225 27.1925 ;
        RECT  11.7225 26.275 11.7875 26.41 ;
        RECT  11.7225 26.275 11.7875 26.41 ;
        RECT  11.7225 26.275 11.7875 26.41 ;
        RECT  11.7225 26.275 11.7875 26.41 ;
        RECT  11.7225 26.275 11.7875 26.41 ;
        RECT  11.7225 26.275 11.7875 26.41 ;
        RECT  10.9825 27.1275 11.1175 27.1925 ;
        RECT  11.3425 25.785 11.4425 25.8475 ;
        RECT  11.3425 25.7825 11.4425 25.845 ;
        RECT  11.67 26.9875 11.7225 27.05 ;
        RECT  11.3425 25.785 11.4425 25.8475 ;
        RECT  11.72 25.8475 11.79 26.0475 ;
        RECT  11.72 26.3775 11.79 26.5125 ;
        RECT  11.72 26.3775 11.79 26.5125 ;
        RECT  10.96 27.1275 11.845 27.1925 ;
        RECT  11.535 26.6125 11.71 26.6775 ;
        RECT  11.015 26.3775 11.085 26.5125 ;
        RECT  11.205 25.9375 11.27 26.6775 ;
        RECT  11.3425 25.7825 11.4425 25.845 ;
        RECT  10.965 26.9875 11.0175 27.05 ;
        RECT  11.72 26.3775 11.79 26.5125 ;
        RECT  10.96 25.7825 11.845 25.8475 ;
        RECT  11.535 26.0475 11.6 26.6775 ;
        RECT  11.72 26.3775 11.79 26.5125 ;
        RECT  11.72 26.3775 11.79 26.5125 ;
        RECT  11.1 26.6125 11.17 26.9025 ;
        RECT  11.015 26.3775 11.085 26.5125 ;
        RECT  10.96 26.9875 11.845 27.0525 ;
        RECT  11.72 26.3775 11.79 26.5125 ;
        RECT  11.72 25.8475 11.79 26.0475 ;
        RECT  11.015 25.8475 11.085 26.0475 ;
        RECT  11.64 26.6125 11.71 26.9025 ;
        RECT  11.1 26.6125 11.27 26.6775 ;
        RECT  10.96 26.9875 11.845 27.0525 ;
        RECT  10.96 27.1275 11.845 27.1925 ;
        RECT  10.96 25.7825 11.845 25.8475 ;
        RECT  11.72 28.2725 11.785 28.4075 ;
        RECT  11.535 28.2725 11.6 28.4075 ;
        RECT  11.02 28.2725 11.085 28.4075 ;
        RECT  11.205 28.2725 11.27 28.4075 ;
        RECT  11.535 27.8075 11.6 27.9425 ;
        RECT  11.72 27.8075 11.785 27.9425 ;
        RECT  11.205 27.8075 11.27 27.9425 ;
        RECT  11.02 27.8075 11.085 27.9425 ;
        RECT  11.64 27.4175 11.705 27.5525 ;
        RECT  11.455 27.4175 11.52 27.5525 ;
        RECT  11.285 27.4175 11.35 27.5525 ;
        RECT  11.1 27.4175 11.165 27.5525 ;
        RECT  11.7225 27.91 11.7875 28.045 ;
        RECT  11.7225 27.91 11.7875 28.045 ;
        RECT  11.7225 27.91 11.7875 28.045 ;
        RECT  11.7225 27.91 11.7875 28.045 ;
        RECT  11.7225 27.91 11.7875 28.045 ;
        RECT  11.7225 27.91 11.7875 28.045 ;
        RECT  11.33 28.4725 11.465 28.5375 ;
        RECT  10.9825 27.1275 11.1175 27.1925 ;
        RECT  11.6875 27.1275 11.8225 27.1925 ;
        RECT  11.3175 27.2675 11.4525 27.3325 ;
        RECT  11.7225 27.91 11.7875 28.045 ;
        RECT  11.7225 27.91 11.7875 28.045 ;
        RECT  11.7225 27.91 11.7875 28.045 ;
        RECT  11.7225 27.91 11.7875 28.045 ;
        RECT  11.2225 28.1575 11.3575 28.2225 ;
        RECT  11.2225 28.1575 11.3575 28.2225 ;
        RECT  11.4475 28.0075 11.5825 28.0725 ;
        RECT  11.4475 28.0075 11.5825 28.0725 ;
        RECT  11.7225 27.91 11.7875 28.045 ;
        RECT  11.7225 27.91 11.7875 28.045 ;
        RECT  11.7225 27.91 11.7875 28.045 ;
        RECT  11.7225 27.91 11.7875 28.045 ;
        RECT  11.2725 27.4175 11.3375 27.5525 ;
        RECT  11.0175 27.91 11.0825 28.045 ;
        RECT  11.0175 27.91 11.0825 28.045 ;
        RECT  11.0175 27.91 11.0825 28.045 ;
        RECT  11.0175 27.91 11.0825 28.045 ;
        RECT  11.0175 27.91 11.0825 28.045 ;
        RECT  11.0175 27.91 11.0825 28.045 ;
        RECT  11.7225 27.91 11.7875 28.045 ;
        RECT  11.7225 27.91 11.7875 28.045 ;
        RECT  11.7225 27.91 11.7875 28.045 ;
        RECT  11.7225 27.91 11.7875 28.045 ;
        RECT  11.4675 27.4175 11.5325 27.5525 ;
        RECT  11.335 27.1275 11.47 27.1925 ;
        RECT  11.335 27.1275 11.47 27.1925 ;
        RECT  11.6875 27.1275 11.8225 27.1925 ;
        RECT  11.33 28.4725 11.465 28.5375 ;
        RECT  11.6875 27.1275 11.8225 27.1925 ;
        RECT  11.6875 27.1275 11.8225 27.1925 ;
        RECT  11.7225 27.91 11.7875 28.045 ;
        RECT  11.7225 27.91 11.7875 28.045 ;
        RECT  11.7225 27.91 11.7875 28.045 ;
        RECT  11.7225 27.91 11.7875 28.045 ;
        RECT  11.7225 27.91 11.7875 28.045 ;
        RECT  11.7225 27.91 11.7875 28.045 ;
        RECT  10.9825 27.1275 11.1175 27.1925 ;
        RECT  11.3425 28.4725 11.4425 28.535 ;
        RECT  11.3425 28.475 11.4425 28.5375 ;
        RECT  11.67 27.27 11.7225 27.3325 ;
        RECT  11.3425 28.4725 11.4425 28.535 ;
        RECT  11.72 28.2725 11.79 28.4725 ;
        RECT  11.72 27.8075 11.79 27.9425 ;
        RECT  11.72 27.8075 11.79 27.9425 ;
        RECT  10.96 27.1275 11.845 27.1925 ;
        RECT  11.535 27.6425 11.71 27.7075 ;
        RECT  11.015 27.8075 11.085 27.9425 ;
        RECT  11.205 27.6425 11.27 28.3825 ;
        RECT  11.3425 28.475 11.4425 28.5375 ;
        RECT  10.965 27.27 11.0175 27.3325 ;
        RECT  11.72 27.8075 11.79 27.9425 ;
        RECT  10.96 28.4725 11.845 28.5375 ;
        RECT  11.535 27.6425 11.6 28.2725 ;
        RECT  11.72 27.8075 11.79 27.9425 ;
        RECT  11.72 27.8075 11.79 27.9425 ;
        RECT  11.1 27.4175 11.17 27.7075 ;
        RECT  11.015 27.8075 11.085 27.9425 ;
        RECT  10.96 27.2675 11.845 27.3325 ;
        RECT  11.72 27.8075 11.79 27.9425 ;
        RECT  11.72 28.2725 11.79 28.4725 ;
        RECT  11.015 28.2725 11.085 28.4725 ;
        RECT  11.64 27.4175 11.71 27.7075 ;
        RECT  11.1 27.6425 11.27 27.7075 ;
        RECT  10.96 27.2675 11.845 27.3325 ;
        RECT  10.96 27.1275 11.845 27.1925 ;
        RECT  10.96 28.4725 11.845 28.5375 ;
        RECT  11.72 28.6025 11.785 28.7375 ;
        RECT  11.535 28.6025 11.6 28.7375 ;
        RECT  11.02 28.6025 11.085 28.7375 ;
        RECT  11.205 28.6025 11.27 28.7375 ;
        RECT  11.535 29.0675 11.6 29.2025 ;
        RECT  11.72 29.0675 11.785 29.2025 ;
        RECT  11.205 29.0675 11.27 29.2025 ;
        RECT  11.02 29.0675 11.085 29.2025 ;
        RECT  11.64 29.4575 11.705 29.5925 ;
        RECT  11.455 29.4575 11.52 29.5925 ;
        RECT  11.285 29.4575 11.35 29.5925 ;
        RECT  11.1 29.4575 11.165 29.5925 ;
        RECT  11.7225 28.965 11.7875 29.1 ;
        RECT  11.7225 28.965 11.7875 29.1 ;
        RECT  11.7225 28.965 11.7875 29.1 ;
        RECT  11.7225 28.965 11.7875 29.1 ;
        RECT  11.7225 28.965 11.7875 29.1 ;
        RECT  11.7225 28.965 11.7875 29.1 ;
        RECT  11.33 28.4725 11.465 28.5375 ;
        RECT  10.9825 29.8175 11.1175 29.8825 ;
        RECT  11.6875 29.8175 11.8225 29.8825 ;
        RECT  11.3175 29.6775 11.4525 29.7425 ;
        RECT  11.7225 28.965 11.7875 29.1 ;
        RECT  11.7225 28.965 11.7875 29.1 ;
        RECT  11.7225 28.965 11.7875 29.1 ;
        RECT  11.7225 28.965 11.7875 29.1 ;
        RECT  11.2225 28.7875 11.3575 28.8525 ;
        RECT  11.2225 28.7875 11.3575 28.8525 ;
        RECT  11.4475 28.9375 11.5825 29.0025 ;
        RECT  11.4475 28.9375 11.5825 29.0025 ;
        RECT  11.7225 28.965 11.7875 29.1 ;
        RECT  11.7225 28.965 11.7875 29.1 ;
        RECT  11.7225 28.965 11.7875 29.1 ;
        RECT  11.7225 28.965 11.7875 29.1 ;
        RECT  11.2725 29.4575 11.3375 29.5925 ;
        RECT  11.0175 28.965 11.0825 29.1 ;
        RECT  11.0175 28.965 11.0825 29.1 ;
        RECT  11.0175 28.965 11.0825 29.1 ;
        RECT  11.0175 28.965 11.0825 29.1 ;
        RECT  11.0175 28.965 11.0825 29.1 ;
        RECT  11.0175 28.965 11.0825 29.1 ;
        RECT  11.7225 28.965 11.7875 29.1 ;
        RECT  11.7225 28.965 11.7875 29.1 ;
        RECT  11.7225 28.965 11.7875 29.1 ;
        RECT  11.7225 28.965 11.7875 29.1 ;
        RECT  11.4675 29.4575 11.5325 29.5925 ;
        RECT  11.335 29.8175 11.47 29.8825 ;
        RECT  11.335 29.8175 11.47 29.8825 ;
        RECT  11.6875 29.8175 11.8225 29.8825 ;
        RECT  11.33 28.4725 11.465 28.5375 ;
        RECT  11.6875 29.8175 11.8225 29.8825 ;
        RECT  11.6875 29.8175 11.8225 29.8825 ;
        RECT  11.7225 28.965 11.7875 29.1 ;
        RECT  11.7225 28.965 11.7875 29.1 ;
        RECT  11.7225 28.965 11.7875 29.1 ;
        RECT  11.7225 28.965 11.7875 29.1 ;
        RECT  11.7225 28.965 11.7875 29.1 ;
        RECT  11.7225 28.965 11.7875 29.1 ;
        RECT  10.9825 29.8175 11.1175 29.8825 ;
        RECT  11.3425 28.475 11.4425 28.5375 ;
        RECT  11.3425 28.4725 11.4425 28.535 ;
        RECT  11.67 29.6775 11.7225 29.74 ;
        RECT  11.3425 28.475 11.4425 28.5375 ;
        RECT  11.72 28.5375 11.79 28.7375 ;
        RECT  11.72 29.0675 11.79 29.2025 ;
        RECT  11.72 29.0675 11.79 29.2025 ;
        RECT  10.96 29.8175 11.845 29.8825 ;
        RECT  11.535 29.3025 11.71 29.3675 ;
        RECT  11.015 29.0675 11.085 29.2025 ;
        RECT  11.205 28.6275 11.27 29.3675 ;
        RECT  11.3425 28.4725 11.4425 28.535 ;
        RECT  10.965 29.6775 11.0175 29.74 ;
        RECT  11.72 29.0675 11.79 29.2025 ;
        RECT  10.96 28.4725 11.845 28.5375 ;
        RECT  11.535 28.7375 11.6 29.3675 ;
        RECT  11.72 29.0675 11.79 29.2025 ;
        RECT  11.72 29.0675 11.79 29.2025 ;
        RECT  11.1 29.3025 11.17 29.5925 ;
        RECT  11.015 29.0675 11.085 29.2025 ;
        RECT  10.96 29.6775 11.845 29.7425 ;
        RECT  11.72 29.0675 11.79 29.2025 ;
        RECT  11.72 28.5375 11.79 28.7375 ;
        RECT  11.015 28.5375 11.085 28.7375 ;
        RECT  11.64 29.3025 11.71 29.5925 ;
        RECT  11.1 29.3025 11.27 29.3675 ;
        RECT  10.96 29.6775 11.845 29.7425 ;
        RECT  10.96 29.8175 11.845 29.8825 ;
        RECT  10.96 28.4725 11.845 28.5375 ;
        RECT  11.72 30.9625 11.785 31.0975 ;
        RECT  11.535 30.9625 11.6 31.0975 ;
        RECT  11.02 30.9625 11.085 31.0975 ;
        RECT  11.205 30.9625 11.27 31.0975 ;
        RECT  11.535 30.4975 11.6 30.6325 ;
        RECT  11.72 30.4975 11.785 30.6325 ;
        RECT  11.205 30.4975 11.27 30.6325 ;
        RECT  11.02 30.4975 11.085 30.6325 ;
        RECT  11.64 30.1075 11.705 30.2425 ;
        RECT  11.455 30.1075 11.52 30.2425 ;
        RECT  11.285 30.1075 11.35 30.2425 ;
        RECT  11.1 30.1075 11.165 30.2425 ;
        RECT  11.7225 30.6 11.7875 30.735 ;
        RECT  11.7225 30.6 11.7875 30.735 ;
        RECT  11.7225 30.6 11.7875 30.735 ;
        RECT  11.7225 30.6 11.7875 30.735 ;
        RECT  11.7225 30.6 11.7875 30.735 ;
        RECT  11.7225 30.6 11.7875 30.735 ;
        RECT  11.33 31.1625 11.465 31.2275 ;
        RECT  10.9825 29.8175 11.1175 29.8825 ;
        RECT  11.6875 29.8175 11.8225 29.8825 ;
        RECT  11.3175 29.9575 11.4525 30.0225 ;
        RECT  11.7225 30.6 11.7875 30.735 ;
        RECT  11.7225 30.6 11.7875 30.735 ;
        RECT  11.7225 30.6 11.7875 30.735 ;
        RECT  11.7225 30.6 11.7875 30.735 ;
        RECT  11.2225 30.8475 11.3575 30.9125 ;
        RECT  11.2225 30.8475 11.3575 30.9125 ;
        RECT  11.4475 30.6975 11.5825 30.7625 ;
        RECT  11.4475 30.6975 11.5825 30.7625 ;
        RECT  11.7225 30.6 11.7875 30.735 ;
        RECT  11.7225 30.6 11.7875 30.735 ;
        RECT  11.7225 30.6 11.7875 30.735 ;
        RECT  11.7225 30.6 11.7875 30.735 ;
        RECT  11.2725 30.1075 11.3375 30.2425 ;
        RECT  11.0175 30.6 11.0825 30.735 ;
        RECT  11.0175 30.6 11.0825 30.735 ;
        RECT  11.0175 30.6 11.0825 30.735 ;
        RECT  11.0175 30.6 11.0825 30.735 ;
        RECT  11.0175 30.6 11.0825 30.735 ;
        RECT  11.0175 30.6 11.0825 30.735 ;
        RECT  11.7225 30.6 11.7875 30.735 ;
        RECT  11.7225 30.6 11.7875 30.735 ;
        RECT  11.7225 30.6 11.7875 30.735 ;
        RECT  11.7225 30.6 11.7875 30.735 ;
        RECT  11.4675 30.1075 11.5325 30.2425 ;
        RECT  11.335 29.8175 11.47 29.8825 ;
        RECT  11.335 29.8175 11.47 29.8825 ;
        RECT  11.6875 29.8175 11.8225 29.8825 ;
        RECT  11.33 31.1625 11.465 31.2275 ;
        RECT  11.6875 29.8175 11.8225 29.8825 ;
        RECT  11.6875 29.8175 11.8225 29.8825 ;
        RECT  11.7225 30.6 11.7875 30.735 ;
        RECT  11.7225 30.6 11.7875 30.735 ;
        RECT  11.7225 30.6 11.7875 30.735 ;
        RECT  11.7225 30.6 11.7875 30.735 ;
        RECT  11.7225 30.6 11.7875 30.735 ;
        RECT  11.7225 30.6 11.7875 30.735 ;
        RECT  10.9825 29.8175 11.1175 29.8825 ;
        RECT  11.3425 31.1625 11.4425 31.225 ;
        RECT  11.3425 31.165 11.4425 31.2275 ;
        RECT  11.67 29.96 11.7225 30.0225 ;
        RECT  11.3425 31.1625 11.4425 31.225 ;
        RECT  11.72 30.9625 11.79 31.1625 ;
        RECT  11.72 30.4975 11.79 30.6325 ;
        RECT  11.72 30.4975 11.79 30.6325 ;
        RECT  10.96 29.8175 11.845 29.8825 ;
        RECT  11.535 30.3325 11.71 30.3975 ;
        RECT  11.015 30.4975 11.085 30.6325 ;
        RECT  11.205 30.3325 11.27 31.0725 ;
        RECT  11.3425 31.165 11.4425 31.2275 ;
        RECT  10.965 29.96 11.0175 30.0225 ;
        RECT  11.72 30.4975 11.79 30.6325 ;
        RECT  10.96 31.1625 11.845 31.2275 ;
        RECT  11.535 30.3325 11.6 30.9625 ;
        RECT  11.72 30.4975 11.79 30.6325 ;
        RECT  11.72 30.4975 11.79 30.6325 ;
        RECT  11.1 30.1075 11.17 30.3975 ;
        RECT  11.015 30.4975 11.085 30.6325 ;
        RECT  10.96 29.9575 11.845 30.0225 ;
        RECT  11.72 30.4975 11.79 30.6325 ;
        RECT  11.72 30.9625 11.79 31.1625 ;
        RECT  11.015 30.9625 11.085 31.1625 ;
        RECT  11.64 30.1075 11.71 30.3975 ;
        RECT  11.1 30.3325 11.27 30.3975 ;
        RECT  10.96 29.9575 11.845 30.0225 ;
        RECT  10.96 29.8175 11.845 29.8825 ;
        RECT  10.96 31.1625 11.845 31.2275 ;
        RECT  11.72 31.2925 11.785 31.4275 ;
        RECT  11.535 31.2925 11.6 31.4275 ;
        RECT  11.02 31.2925 11.085 31.4275 ;
        RECT  11.205 31.2925 11.27 31.4275 ;
        RECT  11.535 31.7575 11.6 31.8925 ;
        RECT  11.72 31.7575 11.785 31.8925 ;
        RECT  11.205 31.7575 11.27 31.8925 ;
        RECT  11.02 31.7575 11.085 31.8925 ;
        RECT  11.64 32.1475 11.705 32.2825 ;
        RECT  11.455 32.1475 11.52 32.2825 ;
        RECT  11.285 32.1475 11.35 32.2825 ;
        RECT  11.1 32.1475 11.165 32.2825 ;
        RECT  11.7225 31.655 11.7875 31.79 ;
        RECT  11.7225 31.655 11.7875 31.79 ;
        RECT  11.7225 31.655 11.7875 31.79 ;
        RECT  11.7225 31.655 11.7875 31.79 ;
        RECT  11.7225 31.655 11.7875 31.79 ;
        RECT  11.7225 31.655 11.7875 31.79 ;
        RECT  11.33 31.1625 11.465 31.2275 ;
        RECT  10.9825 32.5075 11.1175 32.5725 ;
        RECT  11.6875 32.5075 11.8225 32.5725 ;
        RECT  11.3175 32.3675 11.4525 32.4325 ;
        RECT  11.7225 31.655 11.7875 31.79 ;
        RECT  11.7225 31.655 11.7875 31.79 ;
        RECT  11.7225 31.655 11.7875 31.79 ;
        RECT  11.7225 31.655 11.7875 31.79 ;
        RECT  11.2225 31.4775 11.3575 31.5425 ;
        RECT  11.2225 31.4775 11.3575 31.5425 ;
        RECT  11.4475 31.6275 11.5825 31.6925 ;
        RECT  11.4475 31.6275 11.5825 31.6925 ;
        RECT  11.7225 31.655 11.7875 31.79 ;
        RECT  11.7225 31.655 11.7875 31.79 ;
        RECT  11.7225 31.655 11.7875 31.79 ;
        RECT  11.7225 31.655 11.7875 31.79 ;
        RECT  11.2725 32.1475 11.3375 32.2825 ;
        RECT  11.0175 31.655 11.0825 31.79 ;
        RECT  11.0175 31.655 11.0825 31.79 ;
        RECT  11.0175 31.655 11.0825 31.79 ;
        RECT  11.0175 31.655 11.0825 31.79 ;
        RECT  11.0175 31.655 11.0825 31.79 ;
        RECT  11.0175 31.655 11.0825 31.79 ;
        RECT  11.7225 31.655 11.7875 31.79 ;
        RECT  11.7225 31.655 11.7875 31.79 ;
        RECT  11.7225 31.655 11.7875 31.79 ;
        RECT  11.7225 31.655 11.7875 31.79 ;
        RECT  11.4675 32.1475 11.5325 32.2825 ;
        RECT  11.335 32.5075 11.47 32.5725 ;
        RECT  11.335 32.5075 11.47 32.5725 ;
        RECT  11.6875 32.5075 11.8225 32.5725 ;
        RECT  11.33 31.1625 11.465 31.2275 ;
        RECT  11.6875 32.5075 11.8225 32.5725 ;
        RECT  11.6875 32.5075 11.8225 32.5725 ;
        RECT  11.7225 31.655 11.7875 31.79 ;
        RECT  11.7225 31.655 11.7875 31.79 ;
        RECT  11.7225 31.655 11.7875 31.79 ;
        RECT  11.7225 31.655 11.7875 31.79 ;
        RECT  11.7225 31.655 11.7875 31.79 ;
        RECT  11.7225 31.655 11.7875 31.79 ;
        RECT  10.9825 32.5075 11.1175 32.5725 ;
        RECT  11.3425 31.165 11.4425 31.2275 ;
        RECT  11.3425 31.1625 11.4425 31.225 ;
        RECT  11.67 32.3675 11.7225 32.43 ;
        RECT  11.3425 31.165 11.4425 31.2275 ;
        RECT  11.72 31.2275 11.79 31.4275 ;
        RECT  11.72 31.7575 11.79 31.8925 ;
        RECT  11.72 31.7575 11.79 31.8925 ;
        RECT  10.96 32.5075 11.845 32.5725 ;
        RECT  11.535 31.9925 11.71 32.0575 ;
        RECT  11.015 31.7575 11.085 31.8925 ;
        RECT  11.205 31.3175 11.27 32.0575 ;
        RECT  11.3425 31.1625 11.4425 31.225 ;
        RECT  10.965 32.3675 11.0175 32.43 ;
        RECT  11.72 31.7575 11.79 31.8925 ;
        RECT  10.96 31.1625 11.845 31.2275 ;
        RECT  11.535 31.4275 11.6 32.0575 ;
        RECT  11.72 31.7575 11.79 31.8925 ;
        RECT  11.72 31.7575 11.79 31.8925 ;
        RECT  11.1 31.9925 11.17 32.2825 ;
        RECT  11.015 31.7575 11.085 31.8925 ;
        RECT  10.96 32.3675 11.845 32.4325 ;
        RECT  11.72 31.7575 11.79 31.8925 ;
        RECT  11.72 31.2275 11.79 31.4275 ;
        RECT  11.015 31.2275 11.085 31.4275 ;
        RECT  11.64 31.9925 11.71 32.2825 ;
        RECT  11.1 31.9925 11.27 32.0575 ;
        RECT  10.96 32.3675 11.845 32.4325 ;
        RECT  10.96 32.5075 11.845 32.5725 ;
        RECT  10.96 31.1625 11.845 31.2275 ;
        RECT  11.72 33.6525 11.785 33.7875 ;
        RECT  11.535 33.6525 11.6 33.7875 ;
        RECT  11.02 33.6525 11.085 33.7875 ;
        RECT  11.205 33.6525 11.27 33.7875 ;
        RECT  11.535 33.1875 11.6 33.3225 ;
        RECT  11.72 33.1875 11.785 33.3225 ;
        RECT  11.205 33.1875 11.27 33.3225 ;
        RECT  11.02 33.1875 11.085 33.3225 ;
        RECT  11.64 32.7975 11.705 32.9325 ;
        RECT  11.455 32.7975 11.52 32.9325 ;
        RECT  11.285 32.7975 11.35 32.9325 ;
        RECT  11.1 32.7975 11.165 32.9325 ;
        RECT  11.7225 33.29 11.7875 33.425 ;
        RECT  11.7225 33.29 11.7875 33.425 ;
        RECT  11.7225 33.29 11.7875 33.425 ;
        RECT  11.7225 33.29 11.7875 33.425 ;
        RECT  11.7225 33.29 11.7875 33.425 ;
        RECT  11.7225 33.29 11.7875 33.425 ;
        RECT  11.33 33.8525 11.465 33.9175 ;
        RECT  10.9825 32.5075 11.1175 32.5725 ;
        RECT  11.6875 32.5075 11.8225 32.5725 ;
        RECT  11.3175 32.6475 11.4525 32.7125 ;
        RECT  11.7225 33.29 11.7875 33.425 ;
        RECT  11.7225 33.29 11.7875 33.425 ;
        RECT  11.7225 33.29 11.7875 33.425 ;
        RECT  11.7225 33.29 11.7875 33.425 ;
        RECT  11.2225 33.5375 11.3575 33.6025 ;
        RECT  11.2225 33.5375 11.3575 33.6025 ;
        RECT  11.4475 33.3875 11.5825 33.4525 ;
        RECT  11.4475 33.3875 11.5825 33.4525 ;
        RECT  11.7225 33.29 11.7875 33.425 ;
        RECT  11.7225 33.29 11.7875 33.425 ;
        RECT  11.7225 33.29 11.7875 33.425 ;
        RECT  11.7225 33.29 11.7875 33.425 ;
        RECT  11.2725 32.7975 11.3375 32.9325 ;
        RECT  11.0175 33.29 11.0825 33.425 ;
        RECT  11.0175 33.29 11.0825 33.425 ;
        RECT  11.0175 33.29 11.0825 33.425 ;
        RECT  11.0175 33.29 11.0825 33.425 ;
        RECT  11.0175 33.29 11.0825 33.425 ;
        RECT  11.0175 33.29 11.0825 33.425 ;
        RECT  11.7225 33.29 11.7875 33.425 ;
        RECT  11.7225 33.29 11.7875 33.425 ;
        RECT  11.7225 33.29 11.7875 33.425 ;
        RECT  11.7225 33.29 11.7875 33.425 ;
        RECT  11.4675 32.7975 11.5325 32.9325 ;
        RECT  11.335 32.5075 11.47 32.5725 ;
        RECT  11.335 32.5075 11.47 32.5725 ;
        RECT  11.6875 32.5075 11.8225 32.5725 ;
        RECT  11.33 33.8525 11.465 33.9175 ;
        RECT  11.6875 32.5075 11.8225 32.5725 ;
        RECT  11.6875 32.5075 11.8225 32.5725 ;
        RECT  11.7225 33.29 11.7875 33.425 ;
        RECT  11.7225 33.29 11.7875 33.425 ;
        RECT  11.7225 33.29 11.7875 33.425 ;
        RECT  11.7225 33.29 11.7875 33.425 ;
        RECT  11.7225 33.29 11.7875 33.425 ;
        RECT  11.7225 33.29 11.7875 33.425 ;
        RECT  10.9825 32.5075 11.1175 32.5725 ;
        RECT  11.3425 33.8525 11.4425 33.915 ;
        RECT  11.3425 33.855 11.4425 33.9175 ;
        RECT  11.67 32.65 11.7225 32.7125 ;
        RECT  11.3425 33.8525 11.4425 33.915 ;
        RECT  11.72 33.6525 11.79 33.8525 ;
        RECT  11.72 33.1875 11.79 33.3225 ;
        RECT  11.72 33.1875 11.79 33.3225 ;
        RECT  10.96 32.5075 11.845 32.5725 ;
        RECT  11.535 33.0225 11.71 33.0875 ;
        RECT  11.015 33.1875 11.085 33.3225 ;
        RECT  11.205 33.0225 11.27 33.7625 ;
        RECT  11.3425 33.855 11.4425 33.9175 ;
        RECT  10.965 32.65 11.0175 32.7125 ;
        RECT  11.72 33.1875 11.79 33.3225 ;
        RECT  10.96 33.8525 11.845 33.9175 ;
        RECT  11.535 33.0225 11.6 33.6525 ;
        RECT  11.72 33.1875 11.79 33.3225 ;
        RECT  11.72 33.1875 11.79 33.3225 ;
        RECT  11.1 32.7975 11.17 33.0875 ;
        RECT  11.015 33.1875 11.085 33.3225 ;
        RECT  10.96 32.6475 11.845 32.7125 ;
        RECT  11.72 33.1875 11.79 33.3225 ;
        RECT  11.72 33.6525 11.79 33.8525 ;
        RECT  11.015 33.6525 11.085 33.8525 ;
        RECT  11.64 32.7975 11.71 33.0875 ;
        RECT  11.1 33.0225 11.27 33.0875 ;
        RECT  10.96 32.6475 11.845 32.7125 ;
        RECT  10.96 32.5075 11.845 32.5725 ;
        RECT  10.96 33.8525 11.845 33.9175 ;
        RECT  11.72 33.9825 11.785 34.1175 ;
        RECT  11.535 33.9825 11.6 34.1175 ;
        RECT  11.02 33.9825 11.085 34.1175 ;
        RECT  11.205 33.9825 11.27 34.1175 ;
        RECT  11.535 34.4475 11.6 34.5825 ;
        RECT  11.72 34.4475 11.785 34.5825 ;
        RECT  11.205 34.4475 11.27 34.5825 ;
        RECT  11.02 34.4475 11.085 34.5825 ;
        RECT  11.64 34.8375 11.705 34.9725 ;
        RECT  11.455 34.8375 11.52 34.9725 ;
        RECT  11.285 34.8375 11.35 34.9725 ;
        RECT  11.1 34.8375 11.165 34.9725 ;
        RECT  11.7225 34.345 11.7875 34.48 ;
        RECT  11.7225 34.345 11.7875 34.48 ;
        RECT  11.7225 34.345 11.7875 34.48 ;
        RECT  11.7225 34.345 11.7875 34.48 ;
        RECT  11.7225 34.345 11.7875 34.48 ;
        RECT  11.7225 34.345 11.7875 34.48 ;
        RECT  11.33 33.8525 11.465 33.9175 ;
        RECT  10.9825 35.1975 11.1175 35.2625 ;
        RECT  11.6875 35.1975 11.8225 35.2625 ;
        RECT  11.3175 35.0575 11.4525 35.1225 ;
        RECT  11.7225 34.345 11.7875 34.48 ;
        RECT  11.7225 34.345 11.7875 34.48 ;
        RECT  11.7225 34.345 11.7875 34.48 ;
        RECT  11.7225 34.345 11.7875 34.48 ;
        RECT  11.2225 34.1675 11.3575 34.2325 ;
        RECT  11.2225 34.1675 11.3575 34.2325 ;
        RECT  11.4475 34.3175 11.5825 34.3825 ;
        RECT  11.4475 34.3175 11.5825 34.3825 ;
        RECT  11.7225 34.345 11.7875 34.48 ;
        RECT  11.7225 34.345 11.7875 34.48 ;
        RECT  11.7225 34.345 11.7875 34.48 ;
        RECT  11.7225 34.345 11.7875 34.48 ;
        RECT  11.2725 34.8375 11.3375 34.9725 ;
        RECT  11.0175 34.345 11.0825 34.48 ;
        RECT  11.0175 34.345 11.0825 34.48 ;
        RECT  11.0175 34.345 11.0825 34.48 ;
        RECT  11.0175 34.345 11.0825 34.48 ;
        RECT  11.0175 34.345 11.0825 34.48 ;
        RECT  11.0175 34.345 11.0825 34.48 ;
        RECT  11.7225 34.345 11.7875 34.48 ;
        RECT  11.7225 34.345 11.7875 34.48 ;
        RECT  11.7225 34.345 11.7875 34.48 ;
        RECT  11.7225 34.345 11.7875 34.48 ;
        RECT  11.4675 34.8375 11.5325 34.9725 ;
        RECT  11.335 35.1975 11.47 35.2625 ;
        RECT  11.335 35.1975 11.47 35.2625 ;
        RECT  11.6875 35.1975 11.8225 35.2625 ;
        RECT  11.33 33.8525 11.465 33.9175 ;
        RECT  11.6875 35.1975 11.8225 35.2625 ;
        RECT  11.6875 35.1975 11.8225 35.2625 ;
        RECT  11.7225 34.345 11.7875 34.48 ;
        RECT  11.7225 34.345 11.7875 34.48 ;
        RECT  11.7225 34.345 11.7875 34.48 ;
        RECT  11.7225 34.345 11.7875 34.48 ;
        RECT  11.7225 34.345 11.7875 34.48 ;
        RECT  11.7225 34.345 11.7875 34.48 ;
        RECT  10.9825 35.1975 11.1175 35.2625 ;
        RECT  11.3425 33.855 11.4425 33.9175 ;
        RECT  11.3425 33.8525 11.4425 33.915 ;
        RECT  11.67 35.0575 11.7225 35.12 ;
        RECT  11.3425 33.855 11.4425 33.9175 ;
        RECT  11.72 33.9175 11.79 34.1175 ;
        RECT  11.72 34.4475 11.79 34.5825 ;
        RECT  11.72 34.4475 11.79 34.5825 ;
        RECT  10.96 35.1975 11.845 35.2625 ;
        RECT  11.535 34.6825 11.71 34.7475 ;
        RECT  11.015 34.4475 11.085 34.5825 ;
        RECT  11.205 34.0075 11.27 34.7475 ;
        RECT  11.3425 33.8525 11.4425 33.915 ;
        RECT  10.965 35.0575 11.0175 35.12 ;
        RECT  11.72 34.4475 11.79 34.5825 ;
        RECT  10.96 33.8525 11.845 33.9175 ;
        RECT  11.535 34.1175 11.6 34.7475 ;
        RECT  11.72 34.4475 11.79 34.5825 ;
        RECT  11.72 34.4475 11.79 34.5825 ;
        RECT  11.1 34.6825 11.17 34.9725 ;
        RECT  11.015 34.4475 11.085 34.5825 ;
        RECT  10.96 35.0575 11.845 35.1225 ;
        RECT  11.72 34.4475 11.79 34.5825 ;
        RECT  11.72 33.9175 11.79 34.1175 ;
        RECT  11.015 33.9175 11.085 34.1175 ;
        RECT  11.64 34.6825 11.71 34.9725 ;
        RECT  11.1 34.6825 11.27 34.7475 ;
        RECT  10.96 35.0575 11.845 35.1225 ;
        RECT  10.96 35.1975 11.845 35.2625 ;
        RECT  10.96 33.8525 11.845 33.9175 ;
        RECT  11.72 36.3425 11.785 36.4775 ;
        RECT  11.535 36.3425 11.6 36.4775 ;
        RECT  11.02 36.3425 11.085 36.4775 ;
        RECT  11.205 36.3425 11.27 36.4775 ;
        RECT  11.535 35.8775 11.6 36.0125 ;
        RECT  11.72 35.8775 11.785 36.0125 ;
        RECT  11.205 35.8775 11.27 36.0125 ;
        RECT  11.02 35.8775 11.085 36.0125 ;
        RECT  11.64 35.4875 11.705 35.6225 ;
        RECT  11.455 35.4875 11.52 35.6225 ;
        RECT  11.285 35.4875 11.35 35.6225 ;
        RECT  11.1 35.4875 11.165 35.6225 ;
        RECT  11.7225 35.98 11.7875 36.115 ;
        RECT  11.7225 35.98 11.7875 36.115 ;
        RECT  11.7225 35.98 11.7875 36.115 ;
        RECT  11.7225 35.98 11.7875 36.115 ;
        RECT  11.7225 35.98 11.7875 36.115 ;
        RECT  11.7225 35.98 11.7875 36.115 ;
        RECT  11.33 36.5425 11.465 36.6075 ;
        RECT  10.9825 35.1975 11.1175 35.2625 ;
        RECT  11.6875 35.1975 11.8225 35.2625 ;
        RECT  11.3175 35.3375 11.4525 35.4025 ;
        RECT  11.7225 35.98 11.7875 36.115 ;
        RECT  11.7225 35.98 11.7875 36.115 ;
        RECT  11.7225 35.98 11.7875 36.115 ;
        RECT  11.7225 35.98 11.7875 36.115 ;
        RECT  11.2225 36.2275 11.3575 36.2925 ;
        RECT  11.2225 36.2275 11.3575 36.2925 ;
        RECT  11.4475 36.0775 11.5825 36.1425 ;
        RECT  11.4475 36.0775 11.5825 36.1425 ;
        RECT  11.7225 35.98 11.7875 36.115 ;
        RECT  11.7225 35.98 11.7875 36.115 ;
        RECT  11.7225 35.98 11.7875 36.115 ;
        RECT  11.7225 35.98 11.7875 36.115 ;
        RECT  11.2725 35.4875 11.3375 35.6225 ;
        RECT  11.0175 35.98 11.0825 36.115 ;
        RECT  11.0175 35.98 11.0825 36.115 ;
        RECT  11.0175 35.98 11.0825 36.115 ;
        RECT  11.0175 35.98 11.0825 36.115 ;
        RECT  11.0175 35.98 11.0825 36.115 ;
        RECT  11.0175 35.98 11.0825 36.115 ;
        RECT  11.7225 35.98 11.7875 36.115 ;
        RECT  11.7225 35.98 11.7875 36.115 ;
        RECT  11.7225 35.98 11.7875 36.115 ;
        RECT  11.7225 35.98 11.7875 36.115 ;
        RECT  11.4675 35.4875 11.5325 35.6225 ;
        RECT  11.335 35.1975 11.47 35.2625 ;
        RECT  11.335 35.1975 11.47 35.2625 ;
        RECT  11.6875 35.1975 11.8225 35.2625 ;
        RECT  11.33 36.5425 11.465 36.6075 ;
        RECT  11.6875 35.1975 11.8225 35.2625 ;
        RECT  11.6875 35.1975 11.8225 35.2625 ;
        RECT  11.7225 35.98 11.7875 36.115 ;
        RECT  11.7225 35.98 11.7875 36.115 ;
        RECT  11.7225 35.98 11.7875 36.115 ;
        RECT  11.7225 35.98 11.7875 36.115 ;
        RECT  11.7225 35.98 11.7875 36.115 ;
        RECT  11.7225 35.98 11.7875 36.115 ;
        RECT  10.9825 35.1975 11.1175 35.2625 ;
        RECT  11.3425 36.5425 11.4425 36.605 ;
        RECT  11.3425 36.545 11.4425 36.6075 ;
        RECT  11.67 35.34 11.7225 35.4025 ;
        RECT  11.3425 36.5425 11.4425 36.605 ;
        RECT  11.72 36.3425 11.79 36.5425 ;
        RECT  11.72 35.8775 11.79 36.0125 ;
        RECT  11.72 35.8775 11.79 36.0125 ;
        RECT  10.96 35.1975 11.845 35.2625 ;
        RECT  11.535 35.7125 11.71 35.7775 ;
        RECT  11.015 35.8775 11.085 36.0125 ;
        RECT  11.205 35.7125 11.27 36.4525 ;
        RECT  11.3425 36.545 11.4425 36.6075 ;
        RECT  10.965 35.34 11.0175 35.4025 ;
        RECT  11.72 35.8775 11.79 36.0125 ;
        RECT  10.96 36.5425 11.845 36.6075 ;
        RECT  11.535 35.7125 11.6 36.3425 ;
        RECT  11.72 35.8775 11.79 36.0125 ;
        RECT  11.72 35.8775 11.79 36.0125 ;
        RECT  11.1 35.4875 11.17 35.7775 ;
        RECT  11.015 35.8775 11.085 36.0125 ;
        RECT  10.96 35.3375 11.845 35.4025 ;
        RECT  11.72 35.8775 11.79 36.0125 ;
        RECT  11.72 36.3425 11.79 36.5425 ;
        RECT  11.015 36.3425 11.085 36.5425 ;
        RECT  11.64 35.4875 11.71 35.7775 ;
        RECT  11.1 35.7125 11.27 35.7775 ;
        RECT  10.96 35.3375 11.845 35.4025 ;
        RECT  10.96 35.1975 11.845 35.2625 ;
        RECT  10.96 36.5425 11.845 36.6075 ;
        RECT  11.72 36.6725 11.785 36.8075 ;
        RECT  11.535 36.6725 11.6 36.8075 ;
        RECT  11.02 36.6725 11.085 36.8075 ;
        RECT  11.205 36.6725 11.27 36.8075 ;
        RECT  11.535 37.1375 11.6 37.2725 ;
        RECT  11.72 37.1375 11.785 37.2725 ;
        RECT  11.205 37.1375 11.27 37.2725 ;
        RECT  11.02 37.1375 11.085 37.2725 ;
        RECT  11.64 37.5275 11.705 37.6625 ;
        RECT  11.455 37.5275 11.52 37.6625 ;
        RECT  11.285 37.5275 11.35 37.6625 ;
        RECT  11.1 37.5275 11.165 37.6625 ;
        RECT  11.7225 37.035 11.7875 37.17 ;
        RECT  11.7225 37.035 11.7875 37.17 ;
        RECT  11.7225 37.035 11.7875 37.17 ;
        RECT  11.7225 37.035 11.7875 37.17 ;
        RECT  11.7225 37.035 11.7875 37.17 ;
        RECT  11.7225 37.035 11.7875 37.17 ;
        RECT  11.33 36.5425 11.465 36.6075 ;
        RECT  10.9825 37.8875 11.1175 37.9525 ;
        RECT  11.6875 37.8875 11.8225 37.9525 ;
        RECT  11.3175 37.7475 11.4525 37.8125 ;
        RECT  11.7225 37.035 11.7875 37.17 ;
        RECT  11.7225 37.035 11.7875 37.17 ;
        RECT  11.7225 37.035 11.7875 37.17 ;
        RECT  11.7225 37.035 11.7875 37.17 ;
        RECT  11.2225 36.8575 11.3575 36.9225 ;
        RECT  11.2225 36.8575 11.3575 36.9225 ;
        RECT  11.4475 37.0075 11.5825 37.0725 ;
        RECT  11.4475 37.0075 11.5825 37.0725 ;
        RECT  11.7225 37.035 11.7875 37.17 ;
        RECT  11.7225 37.035 11.7875 37.17 ;
        RECT  11.7225 37.035 11.7875 37.17 ;
        RECT  11.7225 37.035 11.7875 37.17 ;
        RECT  11.2725 37.5275 11.3375 37.6625 ;
        RECT  11.0175 37.035 11.0825 37.17 ;
        RECT  11.0175 37.035 11.0825 37.17 ;
        RECT  11.0175 37.035 11.0825 37.17 ;
        RECT  11.0175 37.035 11.0825 37.17 ;
        RECT  11.0175 37.035 11.0825 37.17 ;
        RECT  11.0175 37.035 11.0825 37.17 ;
        RECT  11.7225 37.035 11.7875 37.17 ;
        RECT  11.7225 37.035 11.7875 37.17 ;
        RECT  11.7225 37.035 11.7875 37.17 ;
        RECT  11.7225 37.035 11.7875 37.17 ;
        RECT  11.4675 37.5275 11.5325 37.6625 ;
        RECT  11.335 37.8875 11.47 37.9525 ;
        RECT  11.335 37.8875 11.47 37.9525 ;
        RECT  11.6875 37.8875 11.8225 37.9525 ;
        RECT  11.33 36.5425 11.465 36.6075 ;
        RECT  11.6875 37.8875 11.8225 37.9525 ;
        RECT  11.6875 37.8875 11.8225 37.9525 ;
        RECT  11.7225 37.035 11.7875 37.17 ;
        RECT  11.7225 37.035 11.7875 37.17 ;
        RECT  11.7225 37.035 11.7875 37.17 ;
        RECT  11.7225 37.035 11.7875 37.17 ;
        RECT  11.7225 37.035 11.7875 37.17 ;
        RECT  11.7225 37.035 11.7875 37.17 ;
        RECT  10.9825 37.8875 11.1175 37.9525 ;
        RECT  11.3425 36.545 11.4425 36.6075 ;
        RECT  11.3425 36.5425 11.4425 36.605 ;
        RECT  11.67 37.7475 11.7225 37.81 ;
        RECT  11.3425 36.545 11.4425 36.6075 ;
        RECT  11.72 36.6075 11.79 36.8075 ;
        RECT  11.72 37.1375 11.79 37.2725 ;
        RECT  11.72 37.1375 11.79 37.2725 ;
        RECT  10.96 37.8875 11.845 37.9525 ;
        RECT  11.535 37.3725 11.71 37.4375 ;
        RECT  11.015 37.1375 11.085 37.2725 ;
        RECT  11.205 36.6975 11.27 37.4375 ;
        RECT  11.3425 36.5425 11.4425 36.605 ;
        RECT  10.965 37.7475 11.0175 37.81 ;
        RECT  11.72 37.1375 11.79 37.2725 ;
        RECT  10.96 36.5425 11.845 36.6075 ;
        RECT  11.535 36.8075 11.6 37.4375 ;
        RECT  11.72 37.1375 11.79 37.2725 ;
        RECT  11.72 37.1375 11.79 37.2725 ;
        RECT  11.1 37.3725 11.17 37.6625 ;
        RECT  11.015 37.1375 11.085 37.2725 ;
        RECT  10.96 37.7475 11.845 37.8125 ;
        RECT  11.72 37.1375 11.79 37.2725 ;
        RECT  11.72 36.6075 11.79 36.8075 ;
        RECT  11.015 36.6075 11.085 36.8075 ;
        RECT  11.64 37.3725 11.71 37.6625 ;
        RECT  11.1 37.3725 11.27 37.4375 ;
        RECT  10.96 37.7475 11.845 37.8125 ;
        RECT  10.96 37.8875 11.845 37.9525 ;
        RECT  10.96 36.5425 11.845 36.6075 ;
        RECT  11.72 39.0325 11.785 39.1675 ;
        RECT  11.535 39.0325 11.6 39.1675 ;
        RECT  11.02 39.0325 11.085 39.1675 ;
        RECT  11.205 39.0325 11.27 39.1675 ;
        RECT  11.535 38.5675 11.6 38.7025 ;
        RECT  11.72 38.5675 11.785 38.7025 ;
        RECT  11.205 38.5675 11.27 38.7025 ;
        RECT  11.02 38.5675 11.085 38.7025 ;
        RECT  11.64 38.1775 11.705 38.3125 ;
        RECT  11.455 38.1775 11.52 38.3125 ;
        RECT  11.285 38.1775 11.35 38.3125 ;
        RECT  11.1 38.1775 11.165 38.3125 ;
        RECT  11.7225 38.67 11.7875 38.805 ;
        RECT  11.7225 38.67 11.7875 38.805 ;
        RECT  11.7225 38.67 11.7875 38.805 ;
        RECT  11.7225 38.67 11.7875 38.805 ;
        RECT  11.7225 38.67 11.7875 38.805 ;
        RECT  11.7225 38.67 11.7875 38.805 ;
        RECT  11.33 39.2325 11.465 39.2975 ;
        RECT  10.9825 37.8875 11.1175 37.9525 ;
        RECT  11.6875 37.8875 11.8225 37.9525 ;
        RECT  11.3175 38.0275 11.4525 38.0925 ;
        RECT  11.7225 38.67 11.7875 38.805 ;
        RECT  11.7225 38.67 11.7875 38.805 ;
        RECT  11.7225 38.67 11.7875 38.805 ;
        RECT  11.7225 38.67 11.7875 38.805 ;
        RECT  11.2225 38.9175 11.3575 38.9825 ;
        RECT  11.2225 38.9175 11.3575 38.9825 ;
        RECT  11.4475 38.7675 11.5825 38.8325 ;
        RECT  11.4475 38.7675 11.5825 38.8325 ;
        RECT  11.7225 38.67 11.7875 38.805 ;
        RECT  11.7225 38.67 11.7875 38.805 ;
        RECT  11.7225 38.67 11.7875 38.805 ;
        RECT  11.7225 38.67 11.7875 38.805 ;
        RECT  11.2725 38.1775 11.3375 38.3125 ;
        RECT  11.0175 38.67 11.0825 38.805 ;
        RECT  11.0175 38.67 11.0825 38.805 ;
        RECT  11.0175 38.67 11.0825 38.805 ;
        RECT  11.0175 38.67 11.0825 38.805 ;
        RECT  11.0175 38.67 11.0825 38.805 ;
        RECT  11.0175 38.67 11.0825 38.805 ;
        RECT  11.7225 38.67 11.7875 38.805 ;
        RECT  11.7225 38.67 11.7875 38.805 ;
        RECT  11.7225 38.67 11.7875 38.805 ;
        RECT  11.7225 38.67 11.7875 38.805 ;
        RECT  11.4675 38.1775 11.5325 38.3125 ;
        RECT  11.335 37.8875 11.47 37.9525 ;
        RECT  11.335 37.8875 11.47 37.9525 ;
        RECT  11.6875 37.8875 11.8225 37.9525 ;
        RECT  11.33 39.2325 11.465 39.2975 ;
        RECT  11.6875 37.8875 11.8225 37.9525 ;
        RECT  11.6875 37.8875 11.8225 37.9525 ;
        RECT  11.7225 38.67 11.7875 38.805 ;
        RECT  11.7225 38.67 11.7875 38.805 ;
        RECT  11.7225 38.67 11.7875 38.805 ;
        RECT  11.7225 38.67 11.7875 38.805 ;
        RECT  11.7225 38.67 11.7875 38.805 ;
        RECT  11.7225 38.67 11.7875 38.805 ;
        RECT  10.9825 37.8875 11.1175 37.9525 ;
        RECT  11.3425 39.2325 11.4425 39.295 ;
        RECT  11.3425 39.235 11.4425 39.2975 ;
        RECT  11.67 38.03 11.7225 38.0925 ;
        RECT  11.3425 39.2325 11.4425 39.295 ;
        RECT  11.72 39.0325 11.79 39.2325 ;
        RECT  11.72 38.5675 11.79 38.7025 ;
        RECT  11.72 38.5675 11.79 38.7025 ;
        RECT  10.96 37.8875 11.845 37.9525 ;
        RECT  11.535 38.4025 11.71 38.4675 ;
        RECT  11.015 38.5675 11.085 38.7025 ;
        RECT  11.205 38.4025 11.27 39.1425 ;
        RECT  11.3425 39.235 11.4425 39.2975 ;
        RECT  10.965 38.03 11.0175 38.0925 ;
        RECT  11.72 38.5675 11.79 38.7025 ;
        RECT  10.96 39.2325 11.845 39.2975 ;
        RECT  11.535 38.4025 11.6 39.0325 ;
        RECT  11.72 38.5675 11.79 38.7025 ;
        RECT  11.72 38.5675 11.79 38.7025 ;
        RECT  11.1 38.1775 11.17 38.4675 ;
        RECT  11.015 38.5675 11.085 38.7025 ;
        RECT  10.96 38.0275 11.845 38.0925 ;
        RECT  11.72 38.5675 11.79 38.7025 ;
        RECT  11.72 39.0325 11.79 39.2325 ;
        RECT  11.015 39.0325 11.085 39.2325 ;
        RECT  11.64 38.1775 11.71 38.4675 ;
        RECT  11.1 38.4025 11.27 38.4675 ;
        RECT  10.96 38.0275 11.845 38.0925 ;
        RECT  10.96 37.8875 11.845 37.9525 ;
        RECT  10.96 39.2325 11.845 39.2975 ;
        RECT  11.72 39.3625 11.785 39.4975 ;
        RECT  11.535 39.3625 11.6 39.4975 ;
        RECT  11.02 39.3625 11.085 39.4975 ;
        RECT  11.205 39.3625 11.27 39.4975 ;
        RECT  11.535 39.8275 11.6 39.9625 ;
        RECT  11.72 39.8275 11.785 39.9625 ;
        RECT  11.205 39.8275 11.27 39.9625 ;
        RECT  11.02 39.8275 11.085 39.9625 ;
        RECT  11.64 40.2175 11.705 40.3525 ;
        RECT  11.455 40.2175 11.52 40.3525 ;
        RECT  11.285 40.2175 11.35 40.3525 ;
        RECT  11.1 40.2175 11.165 40.3525 ;
        RECT  11.7225 39.725 11.7875 39.86 ;
        RECT  11.7225 39.725 11.7875 39.86 ;
        RECT  11.7225 39.725 11.7875 39.86 ;
        RECT  11.7225 39.725 11.7875 39.86 ;
        RECT  11.7225 39.725 11.7875 39.86 ;
        RECT  11.7225 39.725 11.7875 39.86 ;
        RECT  11.33 39.2325 11.465 39.2975 ;
        RECT  10.9825 40.5775 11.1175 40.6425 ;
        RECT  11.6875 40.5775 11.8225 40.6425 ;
        RECT  11.3175 40.4375 11.4525 40.5025 ;
        RECT  11.7225 39.725 11.7875 39.86 ;
        RECT  11.7225 39.725 11.7875 39.86 ;
        RECT  11.7225 39.725 11.7875 39.86 ;
        RECT  11.7225 39.725 11.7875 39.86 ;
        RECT  11.2225 39.5475 11.3575 39.6125 ;
        RECT  11.2225 39.5475 11.3575 39.6125 ;
        RECT  11.4475 39.6975 11.5825 39.7625 ;
        RECT  11.4475 39.6975 11.5825 39.7625 ;
        RECT  11.7225 39.725 11.7875 39.86 ;
        RECT  11.7225 39.725 11.7875 39.86 ;
        RECT  11.7225 39.725 11.7875 39.86 ;
        RECT  11.7225 39.725 11.7875 39.86 ;
        RECT  11.2725 40.2175 11.3375 40.3525 ;
        RECT  11.0175 39.725 11.0825 39.86 ;
        RECT  11.0175 39.725 11.0825 39.86 ;
        RECT  11.0175 39.725 11.0825 39.86 ;
        RECT  11.0175 39.725 11.0825 39.86 ;
        RECT  11.0175 39.725 11.0825 39.86 ;
        RECT  11.0175 39.725 11.0825 39.86 ;
        RECT  11.7225 39.725 11.7875 39.86 ;
        RECT  11.7225 39.725 11.7875 39.86 ;
        RECT  11.7225 39.725 11.7875 39.86 ;
        RECT  11.7225 39.725 11.7875 39.86 ;
        RECT  11.4675 40.2175 11.5325 40.3525 ;
        RECT  11.335 40.5775 11.47 40.6425 ;
        RECT  11.335 40.5775 11.47 40.6425 ;
        RECT  11.6875 40.5775 11.8225 40.6425 ;
        RECT  11.33 39.2325 11.465 39.2975 ;
        RECT  11.6875 40.5775 11.8225 40.6425 ;
        RECT  11.6875 40.5775 11.8225 40.6425 ;
        RECT  11.7225 39.725 11.7875 39.86 ;
        RECT  11.7225 39.725 11.7875 39.86 ;
        RECT  11.7225 39.725 11.7875 39.86 ;
        RECT  11.7225 39.725 11.7875 39.86 ;
        RECT  11.7225 39.725 11.7875 39.86 ;
        RECT  11.7225 39.725 11.7875 39.86 ;
        RECT  10.9825 40.5775 11.1175 40.6425 ;
        RECT  11.3425 39.235 11.4425 39.2975 ;
        RECT  11.3425 39.2325 11.4425 39.295 ;
        RECT  11.67 40.4375 11.7225 40.5 ;
        RECT  11.3425 39.235 11.4425 39.2975 ;
        RECT  11.72 39.2975 11.79 39.4975 ;
        RECT  11.72 39.8275 11.79 39.9625 ;
        RECT  11.72 39.8275 11.79 39.9625 ;
        RECT  10.96 40.5775 11.845 40.6425 ;
        RECT  11.535 40.0625 11.71 40.1275 ;
        RECT  11.015 39.8275 11.085 39.9625 ;
        RECT  11.205 39.3875 11.27 40.1275 ;
        RECT  11.3425 39.2325 11.4425 39.295 ;
        RECT  10.965 40.4375 11.0175 40.5 ;
        RECT  11.72 39.8275 11.79 39.9625 ;
        RECT  10.96 39.2325 11.845 39.2975 ;
        RECT  11.535 39.4975 11.6 40.1275 ;
        RECT  11.72 39.8275 11.79 39.9625 ;
        RECT  11.72 39.8275 11.79 39.9625 ;
        RECT  11.1 40.0625 11.17 40.3525 ;
        RECT  11.015 39.8275 11.085 39.9625 ;
        RECT  10.96 40.4375 11.845 40.5025 ;
        RECT  11.72 39.8275 11.79 39.9625 ;
        RECT  11.72 39.2975 11.79 39.4975 ;
        RECT  11.015 39.2975 11.085 39.4975 ;
        RECT  11.64 40.0625 11.71 40.3525 ;
        RECT  11.1 40.0625 11.27 40.1275 ;
        RECT  10.96 40.4375 11.845 40.5025 ;
        RECT  10.96 40.5775 11.845 40.6425 ;
        RECT  10.96 39.2325 11.845 39.2975 ;
        RECT  10.345 41.395 11.755 41.46 ;
        RECT  10.345 41.955 11.755 42.02 ;
        RECT  10.73 41.6075 10.795 42.02 ;
        RECT  10.345 41.955 11.05 42.02 ;
        RECT  10.345 41.395 11.05 41.46 ;
        RECT  10.54 41.1575 10.605 41.2925 ;
        RECT  10.73 41.1575 10.795 41.2925 ;
        RECT  10.54 41.1575 10.605 41.2925 ;
        RECT  10.73 41.1575 10.795 41.2925 ;
        RECT  10.54 41.6075 10.605 41.7425 ;
        RECT  10.73 41.6075 10.795 41.7425 ;
        RECT  10.54 41.6075 10.605 41.7425 ;
        RECT  10.73 41.6075 10.795 41.7425 ;
        RECT  10.73 41.6075 10.795 41.7425 ;
        RECT  10.92 41.6075 10.985 41.7425 ;
        RECT  10.73 41.6075 10.795 41.7425 ;
        RECT  10.92 41.6075 10.985 41.7425 ;
        RECT  10.575 41.395 10.71 41.46 ;
        RECT  10.73 41.8525 10.795 41.9875 ;
        RECT  10.54 41.6075 10.605 41.7425 ;
        RECT  10.92 41.6075 10.985 41.7425 ;
        RECT  10.54 41.1575 10.605 41.2925 ;
        RECT  10.73 41.1575 10.795 41.2925 ;
        RECT  11.435 41.6075 11.5 42.02 ;
        RECT  11.05 41.955 11.755 42.02 ;
        RECT  11.05 41.395 11.755 41.46 ;
        RECT  11.245 41.1575 11.31 41.2925 ;
        RECT  11.435 41.1575 11.5 41.2925 ;
        RECT  11.245 41.1575 11.31 41.2925 ;
        RECT  11.435 41.1575 11.5 41.2925 ;
        RECT  11.245 41.6075 11.31 41.7425 ;
        RECT  11.435 41.6075 11.5 41.7425 ;
        RECT  11.245 41.6075 11.31 41.7425 ;
        RECT  11.435 41.6075 11.5 41.7425 ;
        RECT  11.435 41.6075 11.5 41.7425 ;
        RECT  11.625 41.6075 11.69 41.7425 ;
        RECT  11.435 41.6075 11.5 41.7425 ;
        RECT  11.625 41.6075 11.69 41.7425 ;
        RECT  11.28 41.395 11.415 41.46 ;
        RECT  11.435 41.8525 11.5 41.9875 ;
        RECT  11.245 41.6075 11.31 41.7425 ;
        RECT  11.625 41.6075 11.69 41.7425 ;
        RECT  11.245 41.1575 11.31 41.2925 ;
        RECT  11.435 41.1575 11.5 41.2925 ;
        RECT  10.345 14.3225 11.755 14.3875 ;
        RECT  10.345 18.895 11.755 18.96 ;
        RECT  10.345 14.4525 11.755 14.5175 ;
        RECT  10.31 14.3225 11.085 14.3875 ;
        RECT  10.8525 15.3925 10.9175 16.255 ;
        RECT  10.4775 15.3875 10.5425 16.255 ;
        RECT  10.4775 15.4925 10.7675 15.5575 ;
        RECT  10.6275 15.6925 10.9175 15.7575 ;
        RECT  10.31 18.895 11.085 18.96 ;
        RECT  10.4775 16.4175 10.5425 17.515 ;
        RECT  10.8525 16.415 10.9175 16.61 ;
        RECT  10.31 14.4525 11.085 14.5175 ;
        RECT  10.6275 14.8475 10.6975 15.175 ;
        RECT  10.6675 16.545 10.9175 16.61 ;
        RECT  10.6675 16.545 10.7325 16.74 ;
        RECT  10.4775 17.515 10.975 17.58 ;
        RECT  10.665 17.515 10.73 17.7125 ;
        RECT  10.6575 18.6925 10.975 18.7625 ;
        RECT  10.9375 14.4525 11.0025 14.6825 ;
        RECT  10.7625 14.5175 10.8275 14.67 ;
        RECT  10.4075 18.895 10.475 18.96 ;
        RECT  10.91 17.515 10.975 18.7625 ;
        RECT  10.4075 18.5575 10.765 18.6225 ;
        RECT  10.4075 18.6225 10.475 18.96 ;
        RECT  11.0025 14.5175 11.0175 14.5875 ;
        RECT  10.575 14.3225 10.64 14.3875 ;
        RECT  10.615 14.4525 10.675 14.5175 ;
        RECT  10.7225 15.4575 10.7875 15.5925 ;
        RECT  10.6075 15.6575 10.6725 15.7925 ;
        RECT  10.665 16.345 10.73 16.48 ;
        RECT  10.665 18.4875 10.73 18.6225 ;
        RECT  10.63 18.5575 10.765 18.6225 ;
        RECT  10.4725 17.645 10.5375 17.78 ;
        RECT  10.9375 14.6825 11.0025 14.8175 ;
        RECT  10.855 17.235 10.92 17.37 ;
        RECT  10.3125 14.4525 10.3775 14.5875 ;
        RECT  11.0175 14.4525 11.0825 14.5875 ;
        RECT  10.635 14.3225 10.77 14.3875 ;
        RECT  10.66 18.6925 10.725 18.8275 ;
        RECT  10.6675 16.675 10.7325 17.37 ;
        RECT  10.8525 16.675 10.9175 17.37 ;
        RECT  10.4775 17.645 10.5425 18.34 ;
        RECT  10.6625 17.645 10.7275 18.34 ;
        RECT  10.6675 15.8625 10.7325 16.4175 ;
        RECT  10.8525 15.8625 10.9175 16.4175 ;
        RECT  10.4775 15.8625 10.5425 16.4175 ;
        RECT  10.6625 15.8625 10.7275 16.4175 ;
        RECT  10.5775 14.66 10.6425 14.935 ;
        RECT  10.7625 14.66 10.8275 14.935 ;
        RECT  10.4775 15.1175 10.5425 15.3925 ;
        RECT  10.6625 15.1175 10.7275 15.3925 ;
        RECT  10.6675 15.1175 10.7325 15.3925 ;
        RECT  10.8525 15.1175 10.9175 15.3925 ;
        RECT  10.31 14.3225 11.085 14.3875 ;
        RECT  10.31 18.895 11.085 18.96 ;
        RECT  10.31 14.4525 11.085 14.5175 ;
        RECT  11.015 14.3225 11.79 14.3875 ;
        RECT  11.5575 15.3925 11.6225 16.255 ;
        RECT  11.1825 15.3875 11.2475 16.255 ;
        RECT  11.1825 15.4925 11.4725 15.5575 ;
        RECT  11.3325 15.6925 11.6225 15.7575 ;
        RECT  11.015 18.895 11.79 18.96 ;
        RECT  11.1825 16.4175 11.2475 17.515 ;
        RECT  11.5575 16.415 11.6225 16.61 ;
        RECT  11.015 14.4525 11.79 14.5175 ;
        RECT  11.3325 14.8475 11.4025 15.175 ;
        RECT  11.3725 16.545 11.6225 16.61 ;
        RECT  11.3725 16.545 11.4375 16.74 ;
        RECT  11.1825 17.515 11.68 17.58 ;
        RECT  11.37 17.515 11.435 17.7125 ;
        RECT  11.3625 18.6925 11.68 18.7625 ;
        RECT  11.6425 14.4525 11.7075 14.6825 ;
        RECT  11.4675 14.5175 11.5325 14.67 ;
        RECT  11.1125 18.895 11.18 18.96 ;
        RECT  11.615 17.515 11.68 18.7625 ;
        RECT  11.1125 18.5575 11.47 18.6225 ;
        RECT  11.1125 18.6225 11.18 18.96 ;
        RECT  11.7075 14.5175 11.7225 14.5875 ;
        RECT  11.28 14.3225 11.345 14.3875 ;
        RECT  11.32 14.4525 11.38 14.5175 ;
        RECT  11.4275 15.4575 11.4925 15.5925 ;
        RECT  11.3125 15.6575 11.3775 15.7925 ;
        RECT  11.37 16.345 11.435 16.48 ;
        RECT  11.37 18.4875 11.435 18.6225 ;
        RECT  11.335 18.5575 11.47 18.6225 ;
        RECT  11.1775 17.645 11.2425 17.78 ;
        RECT  11.6425 14.6825 11.7075 14.8175 ;
        RECT  11.56 17.235 11.625 17.37 ;
        RECT  11.0175 14.4525 11.0825 14.5875 ;
        RECT  11.7225 14.4525 11.7875 14.5875 ;
        RECT  11.34 14.3225 11.475 14.3875 ;
        RECT  11.365 18.6925 11.43 18.8275 ;
        RECT  11.3725 16.675 11.4375 17.37 ;
        RECT  11.5575 16.675 11.6225 17.37 ;
        RECT  11.1825 17.645 11.2475 18.34 ;
        RECT  11.3675 17.645 11.4325 18.34 ;
        RECT  11.3725 15.8625 11.4375 16.4175 ;
        RECT  11.5575 15.8625 11.6225 16.4175 ;
        RECT  11.1825 15.8625 11.2475 16.4175 ;
        RECT  11.3675 15.8625 11.4325 16.4175 ;
        RECT  11.2825 14.66 11.3475 14.935 ;
        RECT  11.4675 14.66 11.5325 14.935 ;
        RECT  11.1825 15.1175 11.2475 15.3925 ;
        RECT  11.3675 15.1175 11.4325 15.3925 ;
        RECT  11.3725 15.1175 11.4375 15.3925 ;
        RECT  11.5575 15.1175 11.6225 15.3925 ;
        RECT  11.015 14.3225 11.79 14.3875 ;
        RECT  11.015 18.895 11.79 18.96 ;
        RECT  11.015 14.4525 11.79 14.5175 ;
        RECT  10.345 10.2975 11.755 10.3625 ;
        RECT  10.345 10.4275 11.755 10.4925 ;
        RECT  10.345 11.23 11.755 11.295 ;
        RECT  10.765 13.6925 10.83 13.8275 ;
        RECT  10.39 13.6925 10.455 13.8275 ;
        RECT  10.39 11.765 10.455 11.9 ;
        RECT  10.765 11.765 10.83 11.9 ;
        RECT  10.765 12.8975 10.83 13.3125 ;
        RECT  10.39 12.8975 10.455 13.3125 ;
        RECT  10.39 12.28 10.455 12.695 ;
        RECT  10.765 12.28 10.83 12.695 ;
        RECT  10.575 10.71 10.64 11.125 ;
        RECT  10.39 10.71 10.455 11.125 ;
        RECT  10.73 10.71 10.795 11.125 ;
        RECT  10.915 10.71 10.98 11.125 ;
        RECT  10.575 11.4 10.64 11.535 ;
        RECT  10.39 11.4 10.455 11.535 ;
        RECT  10.73 11.4 10.795 11.535 ;
        RECT  10.915 11.4 10.98 11.535 ;
        RECT  10.5525 10.165 10.6875 10.23 ;
        RECT  10.6275 12.12 10.6925 12.255 ;
        RECT  11.0175 11.765 11.0825 11.9 ;
        RECT  10.93 11.765 10.995 11.9 ;
        RECT  10.3125 12.7275 10.3775 12.8625 ;
        RECT  11.0175 11.195 11.0825 11.33 ;
        RECT  10.3125 11.195 10.3775 11.33 ;
        RECT  10.7325 11.4 10.7975 11.535 ;
        RECT  11.0175 13.6925 11.0825 13.8275 ;
        RECT  10.9325 13.6925 10.9975 13.8275 ;
        RECT  10.7325 10.99 10.7975 11.125 ;
        RECT  10.5925 10.99 10.6575 11.125 ;
        RECT  10.615 10.5775 10.75 10.6425 ;
        RECT  10.4475 10.1675 10.5825 10.2325 ;
        RECT  10.7875 10.2975 10.9225 10.3625 ;
        RECT  11.0175 11.4 11.0825 11.535 ;
        RECT  10.3125 11.4 10.3775 11.535 ;
        RECT  10.45 10.4275 10.585 10.4925 ;
        RECT  10.5925 13.37 10.6575 13.505 ;
        RECT  10.7625 11.765 10.8275 11.9 ;
        RECT  10.4525 12.68 10.5175 12.815 ;
        RECT  10.5925 11.4 10.6575 11.535 ;
        RECT  10.53 13.37 10.595 13.505 ;
        RECT  10.3125 11.765 10.3775 11.9 ;
        RECT  10.7625 12.28 10.8275 12.415 ;
        RECT  10.4975 13.9025 10.5625 14.0375 ;
        RECT  10.3125 13.6925 10.3775 13.8275 ;
        RECT  10.9975 13.6925 11.0175 13.8275 ;
        RECT  10.995 11.765 11.0175 11.9 ;
        RECT  10.665 11.2325 10.7225 11.2925 ;
        RECT  10.64 10.2975 10.7125 10.3625 ;
        RECT  10.6425 10.4275 10.7125 10.4925 ;
        RECT  10.3725 13.6925 10.385 13.8275 ;
        RECT  10.3775 12.7275 10.52 12.8625 ;
        RECT  10.31 11.23 11.085 11.295 ;
        RECT  10.6475 10.4925 10.7125 10.6425 ;
        RECT  10.975 11.4 11.0175 11.535 ;
        RECT  10.915 10.4925 10.98 10.71 ;
        RECT  10.39 10.4925 10.455 10.71 ;
        RECT  10.31 10.4275 11.085 10.4925 ;
        RECT  10.31 10.2975 11.085 10.3625 ;
        RECT  10.3725 11.4 10.385 11.535 ;
        RECT  10.44 12.68 10.455 12.815 ;
        RECT  10.3725 11.765 10.385 11.9 ;
        RECT  10.39 12.695 10.455 12.8975 ;
        RECT  10.765 13.8275 10.83 13.9025 ;
        RECT  10.6275 11.6075 10.79 11.6725 ;
        RECT  10.38 13.6925 10.39 13.8275 ;
        RECT  10.38 11.765 10.39 11.9 ;
        RECT  10.725 11.4825 10.79 11.6075 ;
        RECT  10.6275 11.6075 10.6925 12.205 ;
        RECT  10.765 13.3125 10.83 13.6925 ;
        RECT  10.495 13.9025 10.83 13.9675 ;
        RECT  10.38 11.4 10.39 11.535 ;
        RECT  10.31 10.2975 11.085 10.3625 ;
        RECT  10.31 10.4275 11.085 10.4925 ;
        RECT  10.31 11.23 11.085 11.295 ;
        RECT  11.47 13.6925 11.535 13.8275 ;
        RECT  11.095 13.6925 11.16 13.8275 ;
        RECT  11.095 11.765 11.16 11.9 ;
        RECT  11.47 11.765 11.535 11.9 ;
        RECT  11.47 12.8975 11.535 13.3125 ;
        RECT  11.095 12.8975 11.16 13.3125 ;
        RECT  11.095 12.28 11.16 12.695 ;
        RECT  11.47 12.28 11.535 12.695 ;
        RECT  11.28 10.71 11.345 11.125 ;
        RECT  11.095 10.71 11.16 11.125 ;
        RECT  11.435 10.71 11.5 11.125 ;
        RECT  11.62 10.71 11.685 11.125 ;
        RECT  11.28 11.4 11.345 11.535 ;
        RECT  11.095 11.4 11.16 11.535 ;
        RECT  11.435 11.4 11.5 11.535 ;
        RECT  11.62 11.4 11.685 11.535 ;
        RECT  11.2575 10.165 11.3925 10.23 ;
        RECT  11.3325 12.12 11.3975 12.255 ;
        RECT  11.7225 11.765 11.7875 11.9 ;
        RECT  11.635 11.765 11.7 11.9 ;
        RECT  11.0175 12.7275 11.0825 12.8625 ;
        RECT  11.7225 11.195 11.7875 11.33 ;
        RECT  11.0175 11.195 11.0825 11.33 ;
        RECT  11.4375 11.4 11.5025 11.535 ;
        RECT  11.7225 13.6925 11.7875 13.8275 ;
        RECT  11.6375 13.6925 11.7025 13.8275 ;
        RECT  11.4375 10.99 11.5025 11.125 ;
        RECT  11.2975 10.99 11.3625 11.125 ;
        RECT  11.32 10.5775 11.455 10.6425 ;
        RECT  11.1525 10.1675 11.2875 10.2325 ;
        RECT  11.4925 10.2975 11.6275 10.3625 ;
        RECT  11.7225 11.4 11.7875 11.535 ;
        RECT  11.0175 11.4 11.0825 11.535 ;
        RECT  11.155 10.4275 11.29 10.4925 ;
        RECT  11.2975 13.37 11.3625 13.505 ;
        RECT  11.4675 11.765 11.5325 11.9 ;
        RECT  11.1575 12.68 11.2225 12.815 ;
        RECT  11.2975 11.4 11.3625 11.535 ;
        RECT  11.235 13.37 11.3 13.505 ;
        RECT  11.0175 11.765 11.0825 11.9 ;
        RECT  11.4675 12.28 11.5325 12.415 ;
        RECT  11.2025 13.9025 11.2675 14.0375 ;
        RECT  11.0175 13.6925 11.0825 13.8275 ;
        RECT  11.7025 13.6925 11.7225 13.8275 ;
        RECT  11.7 11.765 11.7225 11.9 ;
        RECT  11.37 11.2325 11.4275 11.2925 ;
        RECT  11.345 10.2975 11.4175 10.3625 ;
        RECT  11.3475 10.4275 11.4175 10.4925 ;
        RECT  11.0775 13.6925 11.09 13.8275 ;
        RECT  11.0825 12.7275 11.225 12.8625 ;
        RECT  11.015 11.23 11.79 11.295 ;
        RECT  11.3525 10.4925 11.4175 10.6425 ;
        RECT  11.68 11.4 11.7225 11.535 ;
        RECT  11.62 10.4925 11.685 10.71 ;
        RECT  11.095 10.4925 11.16 10.71 ;
        RECT  11.015 10.4275 11.79 10.4925 ;
        RECT  11.015 10.2975 11.79 10.3625 ;
        RECT  11.0775 11.4 11.09 11.535 ;
        RECT  11.145 12.68 11.16 12.815 ;
        RECT  11.0775 11.765 11.09 11.9 ;
        RECT  11.095 12.695 11.16 12.8975 ;
        RECT  11.47 13.8275 11.535 13.9025 ;
        RECT  11.3325 11.6075 11.495 11.6725 ;
        RECT  11.085 13.6925 11.095 13.8275 ;
        RECT  11.085 11.765 11.095 11.9 ;
        RECT  11.43 11.4825 11.495 11.6075 ;
        RECT  11.3325 11.6075 11.3975 12.205 ;
        RECT  11.47 13.3125 11.535 13.6925 ;
        RECT  11.2 13.9025 11.535 13.9675 ;
        RECT  11.085 11.4 11.095 11.535 ;
        RECT  11.015 10.2975 11.79 10.3625 ;
        RECT  11.015 10.4275 11.79 10.4925 ;
        RECT  11.015 11.23 11.79 11.295 ;
        RECT  10.345 3.795 11.755 3.86 ;
        RECT  10.345 6.8 11.755 6.865 ;
        RECT  10.345 9.76 11.755 9.825 ;
        RECT  10.345 4.81 11.755 4.875 ;
        RECT  10.345 7.77 11.755 7.835 ;
        RECT  10.345 3.955 11.755 4.02 ;
        RECT  10.885 6.28 10.95 6.415 ;
        RECT  10.7 6.28 10.765 6.415 ;
        RECT  10.885 5.045 10.95 5.18 ;
        RECT  10.7 5.045 10.765 5.18 ;
        RECT  10.695 6.28 10.76 6.415 ;
        RECT  10.51 6.28 10.575 6.415 ;
        RECT  10.695 9.24 10.76 9.375 ;
        RECT  10.51 9.24 10.575 9.375 ;
        RECT  10.695 5.045 10.76 5.18 ;
        RECT  10.51 5.045 10.575 5.18 ;
        RECT  10.885 9.24 10.95 9.375 ;
        RECT  10.7 9.24 10.765 9.375 ;
        RECT  10.695 4.51 10.76 4.645 ;
        RECT  10.51 4.51 10.575 4.645 ;
        RECT  10.835 7.47 10.9 7.605 ;
        RECT  10.65 7.47 10.715 7.605 ;
        RECT  10.885 8.005 10.95 8.14 ;
        RECT  10.7 8.005 10.765 8.14 ;
        RECT  10.695 8.005 10.76 8.14 ;
        RECT  10.51 8.005 10.575 8.14 ;
        RECT  10.885 8.43 10.95 8.565 ;
        RECT  10.7 8.43 10.765 8.565 ;
        RECT  10.885 5.47 10.95 5.605 ;
        RECT  10.7 5.47 10.765 5.605 ;
        RECT  10.885 8.815 10.95 8.95 ;
        RECT  10.7 8.815 10.765 8.95 ;
        RECT  10.695 8.815 10.76 8.95 ;
        RECT  10.51 8.815 10.575 8.95 ;
        RECT  10.695 5.47 10.76 5.605 ;
        RECT  10.51 5.47 10.575 5.605 ;
        RECT  10.695 8.43 10.76 8.565 ;
        RECT  10.51 8.43 10.575 8.565 ;
        RECT  10.695 5.855 10.76 5.99 ;
        RECT  10.51 5.855 10.575 5.99 ;
        RECT  10.885 5.855 10.95 5.99 ;
        RECT  10.7 5.855 10.765 5.99 ;
        RECT  10.695 4.085 10.76 4.22 ;
        RECT  10.51 4.085 10.575 4.22 ;
        RECT  10.77 7.06 10.835 7.195 ;
        RECT  10.585 7.06 10.65 7.195 ;
        RECT  10.5725 3.795 10.7075 3.86 ;
        RECT  10.51 9.2925 10.575 9.4275 ;
        RECT  10.4 7.4775 10.465 7.6125 ;
        RECT  10.51 6.5775 10.575 6.7125 ;
        RECT  10.9325 7.0525 10.9975 7.1875 ;
        RECT  10.51 9.6575 10.575 9.7925 ;
        RECT  11.0175 4.115 11.0825 4.25 ;
        RECT  10.875 8.1975 10.94 8.3325 ;
        RECT  10.8775 6.59 10.9425 6.725 ;
        RECT  10.8775 5.1925 10.9425 5.3275 ;
        RECT  10.3125 3.975 10.3775 4.11 ;
        RECT  10.8875 4.0925 10.9525 4.2275 ;
        RECT  10.8875 5.7025 11.0225 5.7675 ;
        RECT  10.9275 4.6175 10.9925 4.7525 ;
        RECT  10.8875 8.6625 11.0225 8.7275 ;
        RECT  10.835 9.55 10.9 9.685 ;
        RECT  10.755 6.08 10.82 6.215 ;
        RECT  10.745 9.04 10.81 9.175 ;
        RECT  10.5125 7.35 10.6475 7.415 ;
        RECT  11.0175 7.0525 11.0825 7.1875 ;
        RECT  10.4025 4.345 10.5375 4.41 ;
        RECT  10.5125 5.8575 10.5775 5.9925 ;
        RECT  10.8775 9.55 10.9425 9.685 ;
        RECT  10.7 9.04 10.765 9.175 ;
        RECT  11.0175 8.6275 11.0825 8.7625 ;
        RECT  11.0175 3.925 11.0825 4.06 ;
        RECT  10.8775 6.59 10.9425 6.725 ;
        RECT  11.0175 5.6675 11.0825 5.8025 ;
        RECT  10.5125 5.4675 10.5775 5.6025 ;
        RECT  10.7 5.4675 10.765 5.6025 ;
        RECT  10.7 6.08 10.765 6.215 ;
        RECT  10.51 8.4275 10.575 8.5625 ;
        RECT  10.7 8.4275 10.765 8.5625 ;
        RECT  10.31 3.795 11.085 3.86 ;
        RECT  10.38 6.865 10.445 9.76 ;
        RECT  10.885 9.375 10.95 9.685 ;
        RECT  10.51 8.95 10.575 9.24 ;
        RECT  10.51 8.14 10.575 8.43 ;
        RECT  10.65 9.7625 10.7225 9.825 ;
        RECT  10.695 9.375 10.765 9.76 ;
        RECT  10.695 8.14 10.765 8.43 ;
        RECT  10.695 8.66 10.765 8.8175 ;
        RECT  10.885 8.95 10.95 9.24 ;
        RECT  10.885 8.14 10.95 8.43 ;
        RECT  10.695 8.66 11.08 8.73 ;
        RECT  10.31 9.76 11.085 9.825 ;
        RECT  10.31 7.77 11.085 7.835 ;
        RECT  10.38 4.875 10.445 6.8 ;
        RECT  10.885 6.415 10.95 6.725 ;
        RECT  10.51 5.99 10.575 6.28 ;
        RECT  10.585 7.155 10.65 7.605 ;
        RECT  10.695 6.415 10.765 6.8 ;
        RECT  10.695 5.7 10.765 5.8575 ;
        RECT  10.51 6.7125 10.575 6.8 ;
        RECT  10.885 5.99 10.95 6.28 ;
        RECT  10.77 6.93 11.015 6.995 ;
        RECT  10.9325 6.93 11.015 7.0525 ;
        RECT  10.9525 7.0525 11.02 7.1875 ;
        RECT  10.31 6.8 11.085 6.865 ;
        RECT  10.51 5.18 10.575 5.47 ;
        RECT  10.695 4.6425 10.76 4.81 ;
        RECT  10.76 4.15 11.0175 4.22 ;
        RECT  10.51 4.085 10.575 4.51 ;
        RECT  10.695 5.18 10.765 5.47 ;
        RECT  10.4025 4.34 10.575 4.415 ;
        RECT  10.885 5.18 10.95 5.47 ;
        RECT  10.8875 4.02 10.9525 4.0925 ;
        RECT  10.695 5.7 11.08 5.77 ;
        RECT  10.9275 4.73 10.9925 4.845 ;
        RECT  10.31 3.955 11.085 4.02 ;
        RECT  10.31 4.81 11.085 4.875 ;
        RECT  10.45 3.8 10.515 3.8575 ;
        RECT  11.0175 4.04 11.0825 4.1625 ;
        RECT  10.835 7.6025 10.9 7.77 ;
        RECT  10.77 6.995 10.8375 7.0975 ;
        RECT  10.31 3.795 11.085 3.86 ;
        RECT  10.31 6.8 11.085 6.865 ;
        RECT  10.31 9.76 11.085 9.825 ;
        RECT  10.31 4.81 11.085 4.875 ;
        RECT  10.31 7.77 11.085 7.835 ;
        RECT  10.31 3.955 11.085 4.02 ;
        RECT  11.15 6.28 11.215 6.415 ;
        RECT  11.335 6.28 11.4 6.415 ;
        RECT  11.15 5.045 11.215 5.18 ;
        RECT  11.335 5.045 11.4 5.18 ;
        RECT  11.34 6.28 11.405 6.415 ;
        RECT  11.525 6.28 11.59 6.415 ;
        RECT  11.34 9.24 11.405 9.375 ;
        RECT  11.525 9.24 11.59 9.375 ;
        RECT  11.34 5.045 11.405 5.18 ;
        RECT  11.525 5.045 11.59 5.18 ;
        RECT  11.15 9.24 11.215 9.375 ;
        RECT  11.335 9.24 11.4 9.375 ;
        RECT  11.34 4.51 11.405 4.645 ;
        RECT  11.525 4.51 11.59 4.645 ;
        RECT  11.2 7.47 11.265 7.605 ;
        RECT  11.385 7.47 11.45 7.605 ;
        RECT  11.15 8.005 11.215 8.14 ;
        RECT  11.335 8.005 11.4 8.14 ;
        RECT  11.34 8.005 11.405 8.14 ;
        RECT  11.525 8.005 11.59 8.14 ;
        RECT  11.15 8.43 11.215 8.565 ;
        RECT  11.335 8.43 11.4 8.565 ;
        RECT  11.15 5.47 11.215 5.605 ;
        RECT  11.335 5.47 11.4 5.605 ;
        RECT  11.15 8.815 11.215 8.95 ;
        RECT  11.335 8.815 11.4 8.95 ;
        RECT  11.34 8.815 11.405 8.95 ;
        RECT  11.525 8.815 11.59 8.95 ;
        RECT  11.34 5.47 11.405 5.605 ;
        RECT  11.525 5.47 11.59 5.605 ;
        RECT  11.34 8.43 11.405 8.565 ;
        RECT  11.525 8.43 11.59 8.565 ;
        RECT  11.34 5.855 11.405 5.99 ;
        RECT  11.525 5.855 11.59 5.99 ;
        RECT  11.15 5.855 11.215 5.99 ;
        RECT  11.335 5.855 11.4 5.99 ;
        RECT  11.34 4.085 11.405 4.22 ;
        RECT  11.525 4.085 11.59 4.22 ;
        RECT  11.265 7.06 11.33 7.195 ;
        RECT  11.45 7.06 11.515 7.195 ;
        RECT  11.3925 3.795 11.5275 3.86 ;
        RECT  11.525 9.2925 11.59 9.4275 ;
        RECT  11.635 7.4775 11.7 7.6125 ;
        RECT  11.525 6.5775 11.59 6.7125 ;
        RECT  11.1025 7.0525 11.1675 7.1875 ;
        RECT  11.525 9.6575 11.59 9.7925 ;
        RECT  11.0175 4.115 11.0825 4.25 ;
        RECT  11.16 8.1975 11.225 8.3325 ;
        RECT  11.1575 6.59 11.2225 6.725 ;
        RECT  11.1575 5.1925 11.2225 5.3275 ;
        RECT  11.7225 3.975 11.7875 4.11 ;
        RECT  11.1475 4.0925 11.2125 4.2275 ;
        RECT  11.0775 5.7025 11.2125 5.7675 ;
        RECT  11.1075 4.6175 11.1725 4.7525 ;
        RECT  11.0775 8.6625 11.2125 8.7275 ;
        RECT  11.2 9.55 11.265 9.685 ;
        RECT  11.28 6.08 11.345 6.215 ;
        RECT  11.29 9.04 11.355 9.175 ;
        RECT  11.4525 7.35 11.5875 7.415 ;
        RECT  11.0175 7.0525 11.0825 7.1875 ;
        RECT  11.5625 4.345 11.6975 4.41 ;
        RECT  11.5225 5.8575 11.5875 5.9925 ;
        RECT  11.1575 9.55 11.2225 9.685 ;
        RECT  11.335 9.04 11.4 9.175 ;
        RECT  11.0175 8.6275 11.0825 8.7625 ;
        RECT  11.0175 3.925 11.0825 4.06 ;
        RECT  11.1575 6.59 11.2225 6.725 ;
        RECT  11.0175 5.6675 11.0825 5.8025 ;
        RECT  11.5225 5.4675 11.5875 5.6025 ;
        RECT  11.335 5.4675 11.4 5.6025 ;
        RECT  11.335 6.08 11.4 6.215 ;
        RECT  11.525 8.4275 11.59 8.5625 ;
        RECT  11.335 8.4275 11.4 8.5625 ;
        RECT  11.015 3.795 11.79 3.86 ;
        RECT  11.655 6.865 11.72 9.76 ;
        RECT  11.15 9.375 11.215 9.685 ;
        RECT  11.525 8.95 11.59 9.24 ;
        RECT  11.525 8.14 11.59 8.43 ;
        RECT  11.3775 9.7625 11.45 9.825 ;
        RECT  11.335 9.375 11.405 9.76 ;
        RECT  11.335 8.14 11.405 8.43 ;
        RECT  11.335 8.66 11.405 8.8175 ;
        RECT  11.15 8.95 11.215 9.24 ;
        RECT  11.15 8.14 11.215 8.43 ;
        RECT  11.02 8.66 11.405 8.73 ;
        RECT  11.015 9.76 11.79 9.825 ;
        RECT  11.015 7.77 11.79 7.835 ;
        RECT  11.655 4.875 11.72 6.8 ;
        RECT  11.15 6.415 11.215 6.725 ;
        RECT  11.525 5.99 11.59 6.28 ;
        RECT  11.45 7.155 11.515 7.605 ;
        RECT  11.335 6.415 11.405 6.8 ;
        RECT  11.335 5.7 11.405 5.8575 ;
        RECT  11.525 6.7125 11.59 6.8 ;
        RECT  11.15 5.99 11.215 6.28 ;
        RECT  11.085 6.93 11.33 6.995 ;
        RECT  11.085 6.93 11.1675 7.0525 ;
        RECT  11.08 7.0525 11.1475 7.1875 ;
        RECT  11.015 6.8 11.79 6.865 ;
        RECT  11.525 5.18 11.59 5.47 ;
        RECT  11.34 4.6425 11.405 4.81 ;
        RECT  11.0825 4.15 11.34 4.22 ;
        RECT  11.525 4.085 11.59 4.51 ;
        RECT  11.335 5.18 11.405 5.47 ;
        RECT  11.525 4.34 11.6975 4.415 ;
        RECT  11.15 5.18 11.215 5.47 ;
        RECT  11.1475 4.02 11.2125 4.0925 ;
        RECT  11.02 5.7 11.405 5.77 ;
        RECT  11.1075 4.73 11.1725 4.845 ;
        RECT  11.015 3.955 11.79 4.02 ;
        RECT  11.015 4.81 11.79 4.875 ;
        RECT  11.585 3.8 11.65 3.8575 ;
        RECT  11.0175 4.04 11.0825 4.1625 ;
        RECT  11.2 7.6025 11.265 7.77 ;
        RECT  11.2625 6.995 11.33 7.0975 ;
        RECT  11.015 3.795 11.79 3.86 ;
        RECT  11.015 6.8 11.79 6.865 ;
        RECT  11.015 9.76 11.79 9.825 ;
        RECT  11.015 4.81 11.79 4.875 ;
        RECT  11.015 7.77 11.79 7.835 ;
        RECT  11.015 3.955 11.79 4.02 ;
        RECT  10.345 3.1575 11.755 3.2225 ;
        RECT  10.345 1.74 11.755 1.805 ;
        RECT  10.345 3.0275 11.755 3.0925 ;
        RECT  10.345 1.61 11.755 1.675 ;
        RECT  10.4875 5.375 10.5525 5.44 ;
        RECT  10.8275 5.2825 10.8925 5.375 ;
        RECT  10.345 5.375 11.085 5.44 ;
        RECT  10.345 5.505 11.085 5.57 ;
        RECT  10.72 6.1475 11.0175 6.2825 ;
        RECT  10.8275 4.1525 10.8925 4.24 ;
        RECT  10.345 4.0875 11.085 4.1525 ;
        RECT  10.345 3.9575 11.085 4.0225 ;
        RECT  10.7625 4.5075 10.8975 4.5725 ;
        RECT  10.4525 4.3525 10.5175 4.8675 ;
        RECT  10.515 5.765 10.58 6.285 ;
        RECT  10.6225 5.505 10.685 5.57 ;
        RECT  10.67 3.9575 10.7275 4.0225 ;
        RECT  10.6975 5.68 10.7625 5.815 ;
        RECT  10.49 5.9575 10.555 6.0925 ;
        RECT  10.785 5.375 10.92 5.44 ;
        RECT  10.7625 5.975 10.8975 6.04 ;
        RECT  11.0175 6.1475 11.0825 6.2825 ;
        RECT  10.7625 6.015 10.8975 6.08 ;
        RECT  10.5075 3.9575 10.6425 4.0225 ;
        RECT  10.4025 5.505 10.5375 5.57 ;
        RECT  11.0175 4.0875 11.0825 4.2225 ;
        RECT  10.785 4.0875 10.92 4.1525 ;
        RECT  10.63 5.375 10.765 5.44 ;
        RECT  10.865 6.1575 10.93 6.2925 ;
        RECT  10.8425 4.5075 10.9775 4.5725 ;
        RECT  10.4525 4.8675 10.5175 5.2825 ;
        RECT  10.8275 4.8675 10.8925 5.2825 ;
        RECT  10.4525 4.24 10.5175 4.375 ;
        RECT  10.8275 4.24 10.8925 4.375 ;
        RECT  10.515 6.15 10.58 6.285 ;
        RECT  10.7 6.15 10.765 6.285 ;
        RECT  10.515 5.635 10.58 5.77 ;
        RECT  10.7 5.635 10.765 5.77 ;
        RECT  10.345 3.9575 11.085 4.0225 ;
        RECT  10.345 5.375 11.085 5.44 ;
        RECT  10.345 4.0875 11.085 4.1525 ;
        RECT  10.345 5.505 11.085 5.57 ;
        RECT  10.4525 4.24 10.5175 4.375 ;
        RECT  11.1925 5.375 11.2575 5.44 ;
        RECT  11.5325 5.2825 11.5975 5.375 ;
        RECT  11.05 5.375 11.79 5.44 ;
        RECT  11.05 5.505 11.79 5.57 ;
        RECT  11.425 6.1475 11.7225 6.2825 ;
        RECT  11.5325 4.1525 11.5975 4.24 ;
        RECT  11.05 4.0875 11.79 4.1525 ;
        RECT  11.05 3.9575 11.79 4.0225 ;
        RECT  11.4675 4.5075 11.6025 4.5725 ;
        RECT  11.1575 4.3525 11.2225 4.8675 ;
        RECT  11.22 5.765 11.285 6.285 ;
        RECT  11.3275 5.505 11.39 5.57 ;
        RECT  11.375 3.9575 11.4325 4.0225 ;
        RECT  11.4025 5.68 11.4675 5.815 ;
        RECT  11.195 5.9575 11.26 6.0925 ;
        RECT  11.49 5.375 11.625 5.44 ;
        RECT  11.4675 5.975 11.6025 6.04 ;
        RECT  11.7225 6.1475 11.7875 6.2825 ;
        RECT  11.4675 6.015 11.6025 6.08 ;
        RECT  11.2125 3.9575 11.3475 4.0225 ;
        RECT  11.1075 5.505 11.2425 5.57 ;
        RECT  11.7225 4.0875 11.7875 4.2225 ;
        RECT  11.49 4.0875 11.625 4.1525 ;
        RECT  11.335 5.375 11.47 5.44 ;
        RECT  11.57 6.1575 11.635 6.2925 ;
        RECT  11.5475 4.5075 11.6825 4.5725 ;
        RECT  11.1575 4.8675 11.2225 5.2825 ;
        RECT  11.5325 4.8675 11.5975 5.2825 ;
        RECT  11.1575 4.24 11.2225 4.375 ;
        RECT  11.5325 4.24 11.5975 4.375 ;
        RECT  11.22 6.15 11.285 6.285 ;
        RECT  11.405 6.15 11.47 6.285 ;
        RECT  11.22 5.635 11.285 5.77 ;
        RECT  11.405 5.635 11.47 5.77 ;
        RECT  11.05 3.9575 11.79 4.0225 ;
        RECT  11.05 5.375 11.79 5.44 ;
        RECT  11.05 4.0875 11.79 4.1525 ;
        RECT  11.05 5.505 11.79 5.57 ;
        RECT  11.1575 4.24 11.2225 4.375 ;
        RECT  3.875 19.64 3.94 19.7525 ;
        RECT  3.875 21.1175 3.94 21.23 ;
        RECT  3.875 22.33 3.94 22.4425 ;
        RECT  3.875 23.8075 3.94 23.92 ;
        RECT  3.875 25.02 3.94 25.1325 ;
        RECT  3.875 26.4975 3.94 26.61 ;
        RECT  3.875 27.71 3.94 27.8225 ;
        RECT  3.875 29.1875 3.94 29.3 ;
        RECT  3.875 30.4 3.94 30.5125 ;
        RECT  3.875 31.8775 3.94 31.99 ;
        RECT  3.875 33.09 3.94 33.2025 ;
        RECT  3.875 34.5675 3.94 34.68 ;
        RECT  3.875 35.78 3.94 35.8925 ;
        RECT  3.875 37.2575 3.94 37.37 ;
        RECT  3.875 38.47 3.94 38.5825 ;
        RECT  3.875 39.9475 3.94 40.06 ;
        RECT  1.725 8.88 3.125 8.945 ;
        RECT  1.9 10.405 3.125 10.47 ;
        RECT  2.075 11.57 3.125 11.635 ;
        RECT  2.25 13.095 3.125 13.16 ;
        RECT  2.425 14.26 3.125 14.325 ;
        RECT  2.6 15.785 3.125 15.85 ;
        RECT  2.775 16.95 3.125 17.015 ;
        RECT  2.95 18.475 3.125 18.54 ;
        RECT  1.725 20.0 3.125 20.065 ;
        RECT  2.425 19.47 3.125 19.535 ;
        RECT  1.725 20.805 3.125 20.87 ;
        RECT  2.6 21.335 3.125 21.4 ;
        RECT  1.725 22.69 3.125 22.755 ;
        RECT  2.775 22.16 3.125 22.225 ;
        RECT  1.725 23.495 3.125 23.56 ;
        RECT  2.95 24.025 3.125 24.09 ;
        RECT  1.9 25.38 3.125 25.445 ;
        RECT  2.425 24.85 3.125 24.915 ;
        RECT  1.9 26.185 3.125 26.25 ;
        RECT  2.6 26.715 3.125 26.78 ;
        RECT  1.9 28.07 3.125 28.135 ;
        RECT  2.775 27.54 3.125 27.605 ;
        RECT  1.9 28.875 3.125 28.94 ;
        RECT  2.95 29.405 3.125 29.47 ;
        RECT  2.075 30.76 3.125 30.825 ;
        RECT  2.425 30.23 3.125 30.295 ;
        RECT  2.075 31.565 3.125 31.63 ;
        RECT  2.6 32.095 3.125 32.16 ;
        RECT  2.075 33.45 3.125 33.515 ;
        RECT  2.775 32.92 3.125 32.985 ;
        RECT  2.075 34.255 3.125 34.32 ;
        RECT  2.95 34.785 3.125 34.85 ;
        RECT  2.25 36.14 3.125 36.205 ;
        RECT  2.425 35.61 3.125 35.675 ;
        RECT  2.25 36.945 3.125 37.01 ;
        RECT  2.6 37.475 3.125 37.54 ;
        RECT  2.25 38.83 3.125 38.895 ;
        RECT  2.775 38.3 3.125 38.365 ;
        RECT  2.25 39.635 3.125 39.7 ;
        RECT  2.95 40.165 3.125 40.23 ;
        RECT  4.1975 29.3 4.435 29.365 ;
        RECT  4.1975 26.61 4.435 26.675 ;
        RECT  4.1975 33.09 4.435 33.155 ;
        RECT  4.1975 21.23 4.435 21.295 ;
        RECT  4.1975 23.92 4.435 23.985 ;
        RECT  4.1975 35.78 4.435 35.845 ;
        RECT  4.1975 30.4 4.435 30.465 ;
        RECT  4.1975 38.47 4.435 38.535 ;
        RECT  4.1975 27.71 4.435 27.775 ;
        RECT  4.1975 19.64 4.435 19.705 ;
        RECT  4.1975 25.02 4.435 25.085 ;
        RECT  4.1975 22.33 4.435 22.395 ;
        RECT  4.1975 37.37 4.435 37.435 ;
        RECT  4.1975 31.99 4.435 32.055 ;
        RECT  4.1975 40.06 4.435 40.125 ;
        RECT  4.1975 34.68 4.435 34.745 ;
        RECT  1.725 9.6425 6.92 9.7075 ;
        RECT  1.725 12.3325 6.92 12.3975 ;
        RECT  1.725 15.0225 6.92 15.0875 ;
        RECT  1.725 17.7125 6.92 17.7775 ;
        RECT  1.725 20.4025 6.92 20.4675 ;
        RECT  1.725 23.0925 6.92 23.1575 ;
        RECT  1.725 25.7825 6.92 25.8475 ;
        RECT  1.725 28.4725 6.92 28.5375 ;
        RECT  1.725 31.1625 6.92 31.2275 ;
        RECT  1.725 33.8525 6.92 33.9175 ;
        RECT  1.725 36.5425 6.92 36.6075 ;
        RECT  1.725 39.2325 6.92 39.2975 ;
        RECT  1.725 8.2975 6.92 8.3625 ;
        RECT  1.725 10.9875 6.92 11.0525 ;
        RECT  1.725 13.6775 6.92 13.7425 ;
        RECT  1.725 16.3675 6.92 16.4325 ;
        RECT  1.725 19.0575 6.92 19.1225 ;
        RECT  1.725 21.7475 6.92 21.8125 ;
        RECT  1.725 24.4375 6.92 24.5025 ;
        RECT  1.725 27.1275 6.92 27.1925 ;
        RECT  1.725 29.8175 6.92 29.8825 ;
        RECT  1.725 32.5075 6.92 32.5725 ;
        RECT  1.725 35.1975 6.92 35.2625 ;
        RECT  1.725 37.8875 6.92 37.9525 ;
        RECT  1.725 40.5775 6.92 40.6425 ;
        RECT  3.62 8.88 3.685 8.9925 ;
        RECT  3.62 10.3575 3.685 10.47 ;
        RECT  3.62 11.57 3.685 11.6825 ;
        RECT  3.62 13.0475 3.685 13.16 ;
        RECT  5.465 9.48 5.81 9.545 ;
        RECT  5.745 8.88 5.81 9.48 ;
        RECT  6.37 8.88 6.92 8.945 ;
        RECT  5.19 10.825 5.81 10.89 ;
        RECT  5.745 10.405 5.81 10.825 ;
        RECT  6.37 10.405 6.645 10.47 ;
        RECT  4.915 11.15 6.92 11.215 ;
        RECT  4.64 12.495 6.645 12.56 ;
        RECT  4.435 9.24 5.535 9.305 ;
        RECT  4.435 8.71 5.26 8.775 ;
        RECT  4.435 10.045 4.985 10.11 ;
        RECT  4.435 10.575 5.26 10.64 ;
        RECT  4.435 11.93 5.535 11.995 ;
        RECT  4.435 11.4 4.71 11.465 ;
        RECT  4.435 12.735 4.985 12.8 ;
        RECT  4.435 13.265 4.71 13.33 ;
        RECT  3.125 13.095 3.3625 13.16 ;
        RECT  3.125 11.57 3.3625 11.635 ;
        RECT  3.125 8.88 3.3625 8.945 ;
        RECT  3.125 10.405 3.3625 10.47 ;
        RECT  3.055 9.6425 6.92 9.7075 ;
        RECT  3.055 12.3325 6.92 12.3975 ;
        RECT  3.055 8.2975 6.92 8.3625 ;
        RECT  3.055 10.9875 6.92 11.0525 ;
        RECT  3.055 13.6775 6.92 13.7425 ;
        RECT  5.8775 7.0175 5.9425 7.3825 ;
        RECT  5.8775 8.1625 5.9425 8.2975 ;
        RECT  6.2375 8.2275 6.3025 8.2975 ;
        RECT  6.2375 7.0175 6.3025 7.1075 ;
        RECT  6.0475 7.2475 6.1125 8.195 ;
        RECT  6.335 7.715 6.37 7.78 ;
        RECT  5.81 7.715 6.0475 7.78 ;
        RECT  5.81 6.9525 6.37 7.0175 ;
        RECT  5.81 8.2975 6.37 8.3625 ;
        RECT  6.2375 8.0925 6.3025 8.2275 ;
        RECT  6.0475 8.0925 6.1125 8.2275 ;
        RECT  6.2375 7.9575 6.3025 8.0925 ;
        RECT  6.0475 7.9575 6.1125 8.0925 ;
        RECT  6.2375 7.1075 6.3025 7.3825 ;
        RECT  6.0475 7.1075 6.1125 7.3825 ;
        RECT  6.2375 7.1075 6.3025 7.3825 ;
        RECT  6.0475 7.1075 6.1125 7.3825 ;
        RECT  5.8775 7.1075 5.9425 7.3825 ;
        RECT  5.8775 8.0925 5.9425 8.2275 ;
        RECT  6.2 7.715 6.335 7.78 ;
        RECT  5.8775 11.9675 5.9425 12.3325 ;
        RECT  5.8775 11.0525 5.9425 11.1875 ;
        RECT  6.2375 11.0525 6.3025 11.1225 ;
        RECT  6.2375 12.2425 6.3025 12.3325 ;
        RECT  6.0475 11.155 6.1125 12.1025 ;
        RECT  6.335 11.57 6.37 11.635 ;
        RECT  5.81 11.57 6.0475 11.635 ;
        RECT  5.81 12.3325 6.37 12.3975 ;
        RECT  5.81 10.9875 6.37 11.0525 ;
        RECT  6.2375 11.3225 6.3025 11.4575 ;
        RECT  6.0475 11.3225 6.1125 11.4575 ;
        RECT  6.2375 11.1875 6.3025 11.3225 ;
        RECT  6.0475 11.1875 6.1125 11.3225 ;
        RECT  6.2375 11.5875 6.3025 11.8625 ;
        RECT  6.0475 11.5875 6.1125 11.8625 ;
        RECT  6.2375 11.5875 6.3025 11.8625 ;
        RECT  6.0475 11.5875 6.1125 11.8625 ;
        RECT  5.8775 11.6925 5.9425 11.9675 ;
        RECT  5.8775 10.9875 5.9425 11.1225 ;
        RECT  6.2 11.495 6.335 11.56 ;
        RECT  3.1925 7.0175 3.2575 7.3825 ;
        RECT  3.1925 8.1625 3.2575 8.2975 ;
        RECT  3.5525 8.2275 3.6175 8.2975 ;
        RECT  3.5525 7.0175 3.6175 7.1075 ;
        RECT  3.3625 7.2475 3.4275 8.195 ;
        RECT  3.65 7.715 3.685 7.78 ;
        RECT  3.125 7.715 3.3625 7.78 ;
        RECT  3.125 6.9525 3.685 7.0175 ;
        RECT  3.125 8.2975 3.685 8.3625 ;
        RECT  3.5525 8.0925 3.6175 8.2275 ;
        RECT  3.3625 8.0925 3.4275 8.2275 ;
        RECT  3.5525 7.9575 3.6175 8.0925 ;
        RECT  3.3625 7.9575 3.4275 8.0925 ;
        RECT  3.5525 7.1075 3.6175 7.3825 ;
        RECT  3.3625 7.1075 3.4275 7.3825 ;
        RECT  3.5525 7.1075 3.6175 7.3825 ;
        RECT  3.3625 7.1075 3.4275 7.3825 ;
        RECT  3.1925 7.1075 3.2575 7.3825 ;
        RECT  3.1925 8.0925 3.2575 8.2275 ;
        RECT  3.515 7.715 3.65 7.78 ;
        RECT  3.1925 11.9675 3.2575 12.3325 ;
        RECT  3.1925 11.0525 3.2575 11.1875 ;
        RECT  3.5525 11.0525 3.6175 11.1225 ;
        RECT  3.5525 12.2425 3.6175 12.3325 ;
        RECT  3.3625 11.155 3.4275 12.1025 ;
        RECT  3.65 11.57 3.685 11.635 ;
        RECT  3.125 11.57 3.3625 11.635 ;
        RECT  3.125 12.3325 3.685 12.3975 ;
        RECT  3.125 10.9875 3.685 11.0525 ;
        RECT  3.5525 11.3225 3.6175 11.4575 ;
        RECT  3.3625 11.3225 3.4275 11.4575 ;
        RECT  3.5525 11.1875 3.6175 11.3225 ;
        RECT  3.3625 11.1875 3.4275 11.3225 ;
        RECT  3.5525 11.5875 3.6175 11.8625 ;
        RECT  3.3625 11.5875 3.4275 11.8625 ;
        RECT  3.5525 11.5875 3.6175 11.8625 ;
        RECT  3.3625 11.5875 3.4275 11.8625 ;
        RECT  3.1925 11.6925 3.2575 11.9675 ;
        RECT  3.1925 10.9875 3.2575 11.1225 ;
        RECT  3.515 11.495 3.65 11.56 ;
        RECT  3.1925 9.7075 3.2575 10.0725 ;
        RECT  3.1925 10.8525 3.2575 10.9875 ;
        RECT  3.5525 10.9175 3.6175 10.9875 ;
        RECT  3.5525 9.7075 3.6175 9.7975 ;
        RECT  3.3625 9.9375 3.4275 10.885 ;
        RECT  3.65 10.405 3.685 10.47 ;
        RECT  3.125 10.405 3.3625 10.47 ;
        RECT  3.125 9.6425 3.685 9.7075 ;
        RECT  3.125 10.9875 3.685 11.0525 ;
        RECT  3.5525 10.7825 3.6175 10.9175 ;
        RECT  3.3625 10.7825 3.4275 10.9175 ;
        RECT  3.5525 10.6475 3.6175 10.7825 ;
        RECT  3.3625 10.6475 3.4275 10.7825 ;
        RECT  3.5525 9.7975 3.6175 10.0725 ;
        RECT  3.3625 9.7975 3.4275 10.0725 ;
        RECT  3.5525 9.7975 3.6175 10.0725 ;
        RECT  3.3625 9.7975 3.4275 10.0725 ;
        RECT  3.1925 9.7975 3.2575 10.0725 ;
        RECT  3.1925 10.7825 3.2575 10.9175 ;
        RECT  3.515 10.405 3.65 10.47 ;
        RECT  3.1925 14.6575 3.2575 15.0225 ;
        RECT  3.1925 13.7425 3.2575 13.8775 ;
        RECT  3.5525 13.7425 3.6175 13.8125 ;
        RECT  3.5525 14.9325 3.6175 15.0225 ;
        RECT  3.3625 13.845 3.4275 14.7925 ;
        RECT  3.65 14.26 3.685 14.325 ;
        RECT  3.125 14.26 3.3625 14.325 ;
        RECT  3.125 15.0225 3.685 15.0875 ;
        RECT  3.125 13.6775 3.685 13.7425 ;
        RECT  3.5525 14.0125 3.6175 14.1475 ;
        RECT  3.3625 14.0125 3.4275 14.1475 ;
        RECT  3.5525 13.8775 3.6175 14.0125 ;
        RECT  3.3625 13.8775 3.4275 14.0125 ;
        RECT  3.5525 14.2775 3.6175 14.5525 ;
        RECT  3.3625 14.2775 3.4275 14.5525 ;
        RECT  3.5525 14.2775 3.6175 14.5525 ;
        RECT  3.3625 14.2775 3.4275 14.5525 ;
        RECT  3.1925 14.3825 3.2575 14.6575 ;
        RECT  3.1925 13.6775 3.2575 13.8125 ;
        RECT  3.515 14.185 3.65 14.25 ;
        RECT  3.7525 6.985 3.8175 7.2675 ;
        RECT  3.7525 8.15 3.8175 8.33 ;
        RECT  4.3025 6.985 4.3675 7.2675 ;
        RECT  3.9225 6.985 3.9875 7.2675 ;
        RECT  4.3025 8.0475 4.3675 8.33 ;
        RECT  3.89 7.37 3.955 7.435 ;
        RECT  4.1125 7.37 4.1775 7.435 ;
        RECT  3.89 7.4025 3.955 8.1825 ;
        RECT  3.9225 7.37 4.145 7.435 ;
        RECT  4.1125 7.2675 4.1775 7.4025 ;
        RECT  4.4 7.355 4.435 7.42 ;
        RECT  3.685 7.6675 3.9225 7.7325 ;
        RECT  4.16 7.885 4.435 7.95 ;
        RECT  3.685 6.9525 4.435 7.0175 ;
        RECT  3.685 8.2975 4.435 8.3625 ;
        RECT  4.3025 8.0475 4.3675 8.1825 ;
        RECT  4.1125 8.0475 4.1775 8.1825 ;
        RECT  4.3025 7.9125 4.3675 8.0475 ;
        RECT  4.1125 7.9125 4.1775 8.0475 ;
        RECT  4.1125 8.0475 4.1775 8.1825 ;
        RECT  3.9225 8.0475 3.9875 8.1825 ;
        RECT  4.1125 7.9125 4.1775 8.0475 ;
        RECT  3.9225 7.9125 3.9875 8.0475 ;
        RECT  4.3025 7.1325 4.3675 7.2675 ;
        RECT  4.1125 7.1325 4.1775 7.2675 ;
        RECT  4.3025 7.1325 4.3675 7.2675 ;
        RECT  4.1125 7.1325 4.1775 7.2675 ;
        RECT  4.1125 7.1325 4.1775 7.2675 ;
        RECT  3.9225 7.1325 3.9875 7.2675 ;
        RECT  4.1125 7.1325 4.1775 7.2675 ;
        RECT  3.9225 7.1325 3.9875 7.2675 ;
        RECT  3.7525 7.1325 3.8175 7.2675 ;
        RECT  3.7525 8.0475 3.8175 8.1825 ;
        RECT  4.265 7.355 4.4 7.42 ;
        RECT  4.025 7.885 4.16 7.95 ;
        RECT  3.7525 12.0825 3.8175 12.365 ;
        RECT  3.7525 11.02 3.8175 11.2 ;
        RECT  4.3025 12.0825 4.3675 12.365 ;
        RECT  3.9225 12.0825 3.9875 12.365 ;
        RECT  4.3025 11.02 4.3675 11.3025 ;
        RECT  3.89 11.915 3.955 11.98 ;
        RECT  4.1125 11.915 4.1775 11.98 ;
        RECT  3.89 11.1675 3.955 11.9475 ;
        RECT  3.9225 11.915 4.145 11.98 ;
        RECT  4.1125 11.9475 4.1775 12.0825 ;
        RECT  4.4 11.93 4.435 11.995 ;
        RECT  3.685 11.6175 3.9225 11.6825 ;
        RECT  4.16 11.4 4.435 11.465 ;
        RECT  3.685 12.3325 4.435 12.3975 ;
        RECT  3.685 10.9875 4.435 11.0525 ;
        RECT  4.3025 11.4575 4.3675 11.5925 ;
        RECT  4.1125 11.4575 4.1775 11.5925 ;
        RECT  4.3025 11.3225 4.3675 11.4575 ;
        RECT  4.1125 11.3225 4.1775 11.4575 ;
        RECT  4.1125 11.4575 4.1775 11.5925 ;
        RECT  3.9225 11.4575 3.9875 11.5925 ;
        RECT  4.1125 11.3225 4.1775 11.4575 ;
        RECT  3.9225 11.3225 3.9875 11.4575 ;
        RECT  4.3025 11.7925 4.3675 11.9275 ;
        RECT  4.1125 11.7925 4.1775 11.9275 ;
        RECT  4.3025 11.7925 4.3675 11.9275 ;
        RECT  4.1125 11.7925 4.1775 11.9275 ;
        RECT  4.1125 11.7925 4.1775 11.9275 ;
        RECT  3.9225 11.7925 3.9875 11.9275 ;
        RECT  4.1125 11.7925 4.1775 11.9275 ;
        RECT  3.9225 11.7925 3.9875 11.9275 ;
        RECT  3.7525 11.9475 3.8175 12.0825 ;
        RECT  3.7525 11.0325 3.8175 11.1675 ;
        RECT  4.265 11.855 4.4 11.92 ;
        RECT  4.025 11.325 4.16 11.39 ;
        RECT  3.7525 9.675 3.8175 9.9575 ;
        RECT  3.7525 10.84 3.8175 11.02 ;
        RECT  4.3025 9.675 4.3675 9.9575 ;
        RECT  3.9225 9.675 3.9875 9.9575 ;
        RECT  4.3025 10.7375 4.3675 11.02 ;
        RECT  3.89 10.06 3.955 10.125 ;
        RECT  4.1125 10.06 4.1775 10.125 ;
        RECT  3.89 10.0925 3.955 10.8725 ;
        RECT  3.9225 10.06 4.145 10.125 ;
        RECT  4.1125 9.9575 4.1775 10.0925 ;
        RECT  4.4 10.045 4.435 10.11 ;
        RECT  3.685 10.3575 3.9225 10.4225 ;
        RECT  4.16 10.575 4.435 10.64 ;
        RECT  3.685 9.6425 4.435 9.7075 ;
        RECT  3.685 10.9875 4.435 11.0525 ;
        RECT  4.3025 10.7375 4.3675 10.8725 ;
        RECT  4.1125 10.7375 4.1775 10.8725 ;
        RECT  4.3025 10.6025 4.3675 10.7375 ;
        RECT  4.1125 10.6025 4.1775 10.7375 ;
        RECT  4.1125 10.7375 4.1775 10.8725 ;
        RECT  3.9225 10.7375 3.9875 10.8725 ;
        RECT  4.1125 10.6025 4.1775 10.7375 ;
        RECT  3.9225 10.6025 3.9875 10.7375 ;
        RECT  4.3025 9.8225 4.3675 9.9575 ;
        RECT  4.1125 9.8225 4.1775 9.9575 ;
        RECT  4.3025 9.8225 4.3675 9.9575 ;
        RECT  4.1125 9.8225 4.1775 9.9575 ;
        RECT  4.1125 9.8225 4.1775 9.9575 ;
        RECT  3.9225 9.8225 3.9875 9.9575 ;
        RECT  4.1125 9.8225 4.1775 9.9575 ;
        RECT  3.9225 9.8225 3.9875 9.9575 ;
        RECT  3.7525 9.8225 3.8175 9.9575 ;
        RECT  3.7525 10.7375 3.8175 10.8725 ;
        RECT  4.265 10.045 4.4 10.11 ;
        RECT  4.025 10.575 4.16 10.64 ;
        RECT  3.7525 14.7725 3.8175 15.055 ;
        RECT  3.7525 13.71 3.8175 13.89 ;
        RECT  4.3025 14.7725 4.3675 15.055 ;
        RECT  3.9225 14.7725 3.9875 15.055 ;
        RECT  4.3025 13.71 4.3675 13.9925 ;
        RECT  3.89 14.605 3.955 14.67 ;
        RECT  4.1125 14.605 4.1775 14.67 ;
        RECT  3.89 13.8575 3.955 14.6375 ;
        RECT  3.9225 14.605 4.145 14.67 ;
        RECT  4.1125 14.6375 4.1775 14.7725 ;
        RECT  4.4 14.62 4.435 14.685 ;
        RECT  3.685 14.3075 3.9225 14.3725 ;
        RECT  4.16 14.09 4.435 14.155 ;
        RECT  3.685 15.0225 4.435 15.0875 ;
        RECT  3.685 13.6775 4.435 13.7425 ;
        RECT  4.3025 14.1475 4.3675 14.2825 ;
        RECT  4.1125 14.1475 4.1775 14.2825 ;
        RECT  4.3025 14.0125 4.3675 14.1475 ;
        RECT  4.1125 14.0125 4.1775 14.1475 ;
        RECT  4.1125 14.1475 4.1775 14.2825 ;
        RECT  3.9225 14.1475 3.9875 14.2825 ;
        RECT  4.1125 14.0125 4.1775 14.1475 ;
        RECT  3.9225 14.0125 3.9875 14.1475 ;
        RECT  4.3025 14.4825 4.3675 14.6175 ;
        RECT  4.1125 14.4825 4.1775 14.6175 ;
        RECT  4.3025 14.4825 4.3675 14.6175 ;
        RECT  4.1125 14.4825 4.1775 14.6175 ;
        RECT  4.1125 14.4825 4.1775 14.6175 ;
        RECT  3.9225 14.4825 3.9875 14.6175 ;
        RECT  4.1125 14.4825 4.1775 14.6175 ;
        RECT  3.9225 14.4825 3.9875 14.6175 ;
        RECT  3.7525 14.6375 3.8175 14.7725 ;
        RECT  3.7525 13.7225 3.8175 13.8575 ;
        RECT  4.265 14.545 4.4 14.61 ;
        RECT  4.025 14.015 4.16 14.08 ;
        RECT  5.435 9.41 5.57 9.475 ;
        RECT  6.82 8.81 6.955 8.875 ;
        RECT  5.16 10.755 5.295 10.82 ;
        RECT  6.545 10.335 6.68 10.4 ;
        RECT  6.82 11.08 6.955 11.145 ;
        RECT  4.885 11.08 5.02 11.145 ;
        RECT  6.545 12.425 6.68 12.49 ;
        RECT  4.61 12.425 4.745 12.49 ;
        RECT  5.435 9.17 5.57 9.235 ;
        RECT  5.16 8.64 5.295 8.705 ;
        RECT  4.885 9.975 5.02 10.04 ;
        RECT  5.16 10.505 5.295 10.57 ;
        RECT  5.435 11.86 5.57 11.925 ;
        RECT  4.61 11.33 4.745 11.395 ;
        RECT  4.885 12.665 5.02 12.73 ;
        RECT  4.61 13.195 4.745 13.26 ;
        RECT  3.62 14.26 3.685 14.3725 ;
        RECT  3.62 15.7375 3.685 15.85 ;
        RECT  3.62 16.95 3.685 17.0625 ;
        RECT  3.62 18.4275 3.685 18.54 ;
        RECT  5.465 14.86 5.81 14.925 ;
        RECT  5.745 14.26 5.81 14.86 ;
        RECT  6.37 14.26 6.92 14.325 ;
        RECT  5.19 16.205 5.81 16.27 ;
        RECT  5.745 15.785 5.81 16.205 ;
        RECT  6.37 15.785 6.645 15.85 ;
        RECT  4.915 16.53 6.92 16.595 ;
        RECT  4.64 17.875 6.645 17.94 ;
        RECT  4.435 14.62 5.535 14.685 ;
        RECT  4.435 14.09 5.26 14.155 ;
        RECT  4.435 15.425 4.985 15.49 ;
        RECT  4.435 15.955 5.26 16.02 ;
        RECT  4.435 17.31 5.535 17.375 ;
        RECT  4.435 16.78 4.71 16.845 ;
        RECT  4.435 18.115 4.985 18.18 ;
        RECT  4.435 18.645 4.71 18.71 ;
        RECT  3.125 18.475 3.3625 18.54 ;
        RECT  3.125 16.95 3.3625 17.015 ;
        RECT  3.125 14.26 3.3625 14.325 ;
        RECT  3.125 15.785 3.3625 15.85 ;
        RECT  3.055 15.0225 6.92 15.0875 ;
        RECT  3.055 17.7125 6.92 17.7775 ;
        RECT  3.055 13.6775 6.92 13.7425 ;
        RECT  3.055 16.3675 6.92 16.4325 ;
        RECT  3.055 19.0575 6.92 19.1225 ;
        RECT  5.8775 12.3975 5.9425 12.7625 ;
        RECT  5.8775 13.5425 5.9425 13.6775 ;
        RECT  6.2375 13.6075 6.3025 13.6775 ;
        RECT  6.2375 12.3975 6.3025 12.4875 ;
        RECT  6.0475 12.6275 6.1125 13.575 ;
        RECT  6.335 13.095 6.37 13.16 ;
        RECT  5.81 13.095 6.0475 13.16 ;
        RECT  5.81 12.3325 6.37 12.3975 ;
        RECT  5.81 13.6775 6.37 13.7425 ;
        RECT  6.2375 13.4725 6.3025 13.6075 ;
        RECT  6.0475 13.4725 6.1125 13.6075 ;
        RECT  6.2375 13.3375 6.3025 13.4725 ;
        RECT  6.0475 13.3375 6.1125 13.4725 ;
        RECT  6.2375 12.4875 6.3025 12.7625 ;
        RECT  6.0475 12.4875 6.1125 12.7625 ;
        RECT  6.2375 12.4875 6.3025 12.7625 ;
        RECT  6.0475 12.4875 6.1125 12.7625 ;
        RECT  5.8775 12.4875 5.9425 12.7625 ;
        RECT  5.8775 13.4725 5.9425 13.6075 ;
        RECT  6.2 13.095 6.335 13.16 ;
        RECT  5.8775 17.3475 5.9425 17.7125 ;
        RECT  5.8775 16.4325 5.9425 16.5675 ;
        RECT  6.2375 16.4325 6.3025 16.5025 ;
        RECT  6.2375 17.6225 6.3025 17.7125 ;
        RECT  6.0475 16.535 6.1125 17.4825 ;
        RECT  6.335 16.95 6.37 17.015 ;
        RECT  5.81 16.95 6.0475 17.015 ;
        RECT  5.81 17.7125 6.37 17.7775 ;
        RECT  5.81 16.3675 6.37 16.4325 ;
        RECT  6.2375 16.7025 6.3025 16.8375 ;
        RECT  6.0475 16.7025 6.1125 16.8375 ;
        RECT  6.2375 16.5675 6.3025 16.7025 ;
        RECT  6.0475 16.5675 6.1125 16.7025 ;
        RECT  6.2375 16.9675 6.3025 17.2425 ;
        RECT  6.0475 16.9675 6.1125 17.2425 ;
        RECT  6.2375 16.9675 6.3025 17.2425 ;
        RECT  6.0475 16.9675 6.1125 17.2425 ;
        RECT  5.8775 17.0725 5.9425 17.3475 ;
        RECT  5.8775 16.3675 5.9425 16.5025 ;
        RECT  6.2 16.875 6.335 16.94 ;
        RECT  3.1925 12.3975 3.2575 12.7625 ;
        RECT  3.1925 13.5425 3.2575 13.6775 ;
        RECT  3.5525 13.6075 3.6175 13.6775 ;
        RECT  3.5525 12.3975 3.6175 12.4875 ;
        RECT  3.3625 12.6275 3.4275 13.575 ;
        RECT  3.65 13.095 3.685 13.16 ;
        RECT  3.125 13.095 3.3625 13.16 ;
        RECT  3.125 12.3325 3.685 12.3975 ;
        RECT  3.125 13.6775 3.685 13.7425 ;
        RECT  3.5525 13.4725 3.6175 13.6075 ;
        RECT  3.3625 13.4725 3.4275 13.6075 ;
        RECT  3.5525 13.3375 3.6175 13.4725 ;
        RECT  3.3625 13.3375 3.4275 13.4725 ;
        RECT  3.5525 12.4875 3.6175 12.7625 ;
        RECT  3.3625 12.4875 3.4275 12.7625 ;
        RECT  3.5525 12.4875 3.6175 12.7625 ;
        RECT  3.3625 12.4875 3.4275 12.7625 ;
        RECT  3.1925 12.4875 3.2575 12.7625 ;
        RECT  3.1925 13.4725 3.2575 13.6075 ;
        RECT  3.515 13.095 3.65 13.16 ;
        RECT  3.1925 17.3475 3.2575 17.7125 ;
        RECT  3.1925 16.4325 3.2575 16.5675 ;
        RECT  3.5525 16.4325 3.6175 16.5025 ;
        RECT  3.5525 17.6225 3.6175 17.7125 ;
        RECT  3.3625 16.535 3.4275 17.4825 ;
        RECT  3.65 16.95 3.685 17.015 ;
        RECT  3.125 16.95 3.3625 17.015 ;
        RECT  3.125 17.7125 3.685 17.7775 ;
        RECT  3.125 16.3675 3.685 16.4325 ;
        RECT  3.5525 16.7025 3.6175 16.8375 ;
        RECT  3.3625 16.7025 3.4275 16.8375 ;
        RECT  3.5525 16.5675 3.6175 16.7025 ;
        RECT  3.3625 16.5675 3.4275 16.7025 ;
        RECT  3.5525 16.9675 3.6175 17.2425 ;
        RECT  3.3625 16.9675 3.4275 17.2425 ;
        RECT  3.5525 16.9675 3.6175 17.2425 ;
        RECT  3.3625 16.9675 3.4275 17.2425 ;
        RECT  3.1925 17.0725 3.2575 17.3475 ;
        RECT  3.1925 16.3675 3.2575 16.5025 ;
        RECT  3.515 16.875 3.65 16.94 ;
        RECT  3.1925 15.0875 3.2575 15.4525 ;
        RECT  3.1925 16.2325 3.2575 16.3675 ;
        RECT  3.5525 16.2975 3.6175 16.3675 ;
        RECT  3.5525 15.0875 3.6175 15.1775 ;
        RECT  3.3625 15.3175 3.4275 16.265 ;
        RECT  3.65 15.785 3.685 15.85 ;
        RECT  3.125 15.785 3.3625 15.85 ;
        RECT  3.125 15.0225 3.685 15.0875 ;
        RECT  3.125 16.3675 3.685 16.4325 ;
        RECT  3.5525 16.1625 3.6175 16.2975 ;
        RECT  3.3625 16.1625 3.4275 16.2975 ;
        RECT  3.5525 16.0275 3.6175 16.1625 ;
        RECT  3.3625 16.0275 3.4275 16.1625 ;
        RECT  3.5525 15.1775 3.6175 15.4525 ;
        RECT  3.3625 15.1775 3.4275 15.4525 ;
        RECT  3.5525 15.1775 3.6175 15.4525 ;
        RECT  3.3625 15.1775 3.4275 15.4525 ;
        RECT  3.1925 15.1775 3.2575 15.4525 ;
        RECT  3.1925 16.1625 3.2575 16.2975 ;
        RECT  3.515 15.785 3.65 15.85 ;
        RECT  3.1925 20.0375 3.2575 20.4025 ;
        RECT  3.1925 19.1225 3.2575 19.2575 ;
        RECT  3.5525 19.1225 3.6175 19.1925 ;
        RECT  3.5525 20.3125 3.6175 20.4025 ;
        RECT  3.3625 19.225 3.4275 20.1725 ;
        RECT  3.65 19.64 3.685 19.705 ;
        RECT  3.125 19.64 3.3625 19.705 ;
        RECT  3.125 20.4025 3.685 20.4675 ;
        RECT  3.125 19.0575 3.685 19.1225 ;
        RECT  3.5525 19.3925 3.6175 19.5275 ;
        RECT  3.3625 19.3925 3.4275 19.5275 ;
        RECT  3.5525 19.2575 3.6175 19.3925 ;
        RECT  3.3625 19.2575 3.4275 19.3925 ;
        RECT  3.5525 19.6575 3.6175 19.9325 ;
        RECT  3.3625 19.6575 3.4275 19.9325 ;
        RECT  3.5525 19.6575 3.6175 19.9325 ;
        RECT  3.3625 19.6575 3.4275 19.9325 ;
        RECT  3.1925 19.7625 3.2575 20.0375 ;
        RECT  3.1925 19.0575 3.2575 19.1925 ;
        RECT  3.515 19.565 3.65 19.63 ;
        RECT  3.7525 12.365 3.8175 12.6475 ;
        RECT  3.7525 13.53 3.8175 13.71 ;
        RECT  4.3025 12.365 4.3675 12.6475 ;
        RECT  3.9225 12.365 3.9875 12.6475 ;
        RECT  4.3025 13.4275 4.3675 13.71 ;
        RECT  3.89 12.75 3.955 12.815 ;
        RECT  4.1125 12.75 4.1775 12.815 ;
        RECT  3.89 12.7825 3.955 13.5625 ;
        RECT  3.9225 12.75 4.145 12.815 ;
        RECT  4.1125 12.6475 4.1775 12.7825 ;
        RECT  4.4 12.735 4.435 12.8 ;
        RECT  3.685 13.0475 3.9225 13.1125 ;
        RECT  4.16 13.265 4.435 13.33 ;
        RECT  3.685 12.3325 4.435 12.3975 ;
        RECT  3.685 13.6775 4.435 13.7425 ;
        RECT  4.3025 13.4275 4.3675 13.5625 ;
        RECT  4.1125 13.4275 4.1775 13.5625 ;
        RECT  4.3025 13.2925 4.3675 13.4275 ;
        RECT  4.1125 13.2925 4.1775 13.4275 ;
        RECT  4.1125 13.4275 4.1775 13.5625 ;
        RECT  3.9225 13.4275 3.9875 13.5625 ;
        RECT  4.1125 13.2925 4.1775 13.4275 ;
        RECT  3.9225 13.2925 3.9875 13.4275 ;
        RECT  4.3025 12.5125 4.3675 12.6475 ;
        RECT  4.1125 12.5125 4.1775 12.6475 ;
        RECT  4.3025 12.5125 4.3675 12.6475 ;
        RECT  4.1125 12.5125 4.1775 12.6475 ;
        RECT  4.1125 12.5125 4.1775 12.6475 ;
        RECT  3.9225 12.5125 3.9875 12.6475 ;
        RECT  4.1125 12.5125 4.1775 12.6475 ;
        RECT  3.9225 12.5125 3.9875 12.6475 ;
        RECT  3.7525 12.5125 3.8175 12.6475 ;
        RECT  3.7525 13.4275 3.8175 13.5625 ;
        RECT  4.265 12.735 4.4 12.8 ;
        RECT  4.025 13.265 4.16 13.33 ;
        RECT  3.7525 17.4625 3.8175 17.745 ;
        RECT  3.7525 16.4 3.8175 16.58 ;
        RECT  4.3025 17.4625 4.3675 17.745 ;
        RECT  3.9225 17.4625 3.9875 17.745 ;
        RECT  4.3025 16.4 4.3675 16.6825 ;
        RECT  3.89 17.295 3.955 17.36 ;
        RECT  4.1125 17.295 4.1775 17.36 ;
        RECT  3.89 16.5475 3.955 17.3275 ;
        RECT  3.9225 17.295 4.145 17.36 ;
        RECT  4.1125 17.3275 4.1775 17.4625 ;
        RECT  4.4 17.31 4.435 17.375 ;
        RECT  3.685 16.9975 3.9225 17.0625 ;
        RECT  4.16 16.78 4.435 16.845 ;
        RECT  3.685 17.7125 4.435 17.7775 ;
        RECT  3.685 16.3675 4.435 16.4325 ;
        RECT  4.3025 16.8375 4.3675 16.9725 ;
        RECT  4.1125 16.8375 4.1775 16.9725 ;
        RECT  4.3025 16.7025 4.3675 16.8375 ;
        RECT  4.1125 16.7025 4.1775 16.8375 ;
        RECT  4.1125 16.8375 4.1775 16.9725 ;
        RECT  3.9225 16.8375 3.9875 16.9725 ;
        RECT  4.1125 16.7025 4.1775 16.8375 ;
        RECT  3.9225 16.7025 3.9875 16.8375 ;
        RECT  4.3025 17.1725 4.3675 17.3075 ;
        RECT  4.1125 17.1725 4.1775 17.3075 ;
        RECT  4.3025 17.1725 4.3675 17.3075 ;
        RECT  4.1125 17.1725 4.1775 17.3075 ;
        RECT  4.1125 17.1725 4.1775 17.3075 ;
        RECT  3.9225 17.1725 3.9875 17.3075 ;
        RECT  4.1125 17.1725 4.1775 17.3075 ;
        RECT  3.9225 17.1725 3.9875 17.3075 ;
        RECT  3.7525 17.3275 3.8175 17.4625 ;
        RECT  3.7525 16.4125 3.8175 16.5475 ;
        RECT  4.265 17.235 4.4 17.3 ;
        RECT  4.025 16.705 4.16 16.77 ;
        RECT  3.7525 15.055 3.8175 15.3375 ;
        RECT  3.7525 16.22 3.8175 16.4 ;
        RECT  4.3025 15.055 4.3675 15.3375 ;
        RECT  3.9225 15.055 3.9875 15.3375 ;
        RECT  4.3025 16.1175 4.3675 16.4 ;
        RECT  3.89 15.44 3.955 15.505 ;
        RECT  4.1125 15.44 4.1775 15.505 ;
        RECT  3.89 15.4725 3.955 16.2525 ;
        RECT  3.9225 15.44 4.145 15.505 ;
        RECT  4.1125 15.3375 4.1775 15.4725 ;
        RECT  4.4 15.425 4.435 15.49 ;
        RECT  3.685 15.7375 3.9225 15.8025 ;
        RECT  4.16 15.955 4.435 16.02 ;
        RECT  3.685 15.0225 4.435 15.0875 ;
        RECT  3.685 16.3675 4.435 16.4325 ;
        RECT  4.3025 16.1175 4.3675 16.2525 ;
        RECT  4.1125 16.1175 4.1775 16.2525 ;
        RECT  4.3025 15.9825 4.3675 16.1175 ;
        RECT  4.1125 15.9825 4.1775 16.1175 ;
        RECT  4.1125 16.1175 4.1775 16.2525 ;
        RECT  3.9225 16.1175 3.9875 16.2525 ;
        RECT  4.1125 15.9825 4.1775 16.1175 ;
        RECT  3.9225 15.9825 3.9875 16.1175 ;
        RECT  4.3025 15.2025 4.3675 15.3375 ;
        RECT  4.1125 15.2025 4.1775 15.3375 ;
        RECT  4.3025 15.2025 4.3675 15.3375 ;
        RECT  4.1125 15.2025 4.1775 15.3375 ;
        RECT  4.1125 15.2025 4.1775 15.3375 ;
        RECT  3.9225 15.2025 3.9875 15.3375 ;
        RECT  4.1125 15.2025 4.1775 15.3375 ;
        RECT  3.9225 15.2025 3.9875 15.3375 ;
        RECT  3.7525 15.2025 3.8175 15.3375 ;
        RECT  3.7525 16.1175 3.8175 16.2525 ;
        RECT  4.265 15.425 4.4 15.49 ;
        RECT  4.025 15.955 4.16 16.02 ;
        RECT  3.7525 20.1525 3.8175 20.435 ;
        RECT  3.7525 19.09 3.8175 19.27 ;
        RECT  4.3025 20.1525 4.3675 20.435 ;
        RECT  3.9225 20.1525 3.9875 20.435 ;
        RECT  4.3025 19.09 4.3675 19.3725 ;
        RECT  3.89 19.985 3.955 20.05 ;
        RECT  4.1125 19.985 4.1775 20.05 ;
        RECT  3.89 19.2375 3.955 20.0175 ;
        RECT  3.9225 19.985 4.145 20.05 ;
        RECT  4.1125 20.0175 4.1775 20.1525 ;
        RECT  4.4 20.0 4.435 20.065 ;
        RECT  3.685 19.6875 3.9225 19.7525 ;
        RECT  4.16 19.47 4.435 19.535 ;
        RECT  3.685 20.4025 4.435 20.4675 ;
        RECT  3.685 19.0575 4.435 19.1225 ;
        RECT  4.3025 19.5275 4.3675 19.6625 ;
        RECT  4.1125 19.5275 4.1775 19.6625 ;
        RECT  4.3025 19.3925 4.3675 19.5275 ;
        RECT  4.1125 19.3925 4.1775 19.5275 ;
        RECT  4.1125 19.5275 4.1775 19.6625 ;
        RECT  3.9225 19.5275 3.9875 19.6625 ;
        RECT  4.1125 19.3925 4.1775 19.5275 ;
        RECT  3.9225 19.3925 3.9875 19.5275 ;
        RECT  4.3025 19.8625 4.3675 19.9975 ;
        RECT  4.1125 19.8625 4.1775 19.9975 ;
        RECT  4.3025 19.8625 4.3675 19.9975 ;
        RECT  4.1125 19.8625 4.1775 19.9975 ;
        RECT  4.1125 19.8625 4.1775 19.9975 ;
        RECT  3.9225 19.8625 3.9875 19.9975 ;
        RECT  4.1125 19.8625 4.1775 19.9975 ;
        RECT  3.9225 19.8625 3.9875 19.9975 ;
        RECT  3.7525 20.0175 3.8175 20.1525 ;
        RECT  3.7525 19.1025 3.8175 19.2375 ;
        RECT  4.265 19.925 4.4 19.99 ;
        RECT  4.025 19.395 4.16 19.46 ;
        RECT  5.435 14.79 5.57 14.855 ;
        RECT  6.82 14.19 6.955 14.255 ;
        RECT  5.16 16.135 5.295 16.2 ;
        RECT  6.545 15.715 6.68 15.78 ;
        RECT  6.82 16.46 6.955 16.525 ;
        RECT  4.885 16.46 5.02 16.525 ;
        RECT  6.545 17.805 6.68 17.87 ;
        RECT  4.61 17.805 4.745 17.87 ;
        RECT  5.435 14.55 5.57 14.615 ;
        RECT  5.16 14.02 5.295 14.085 ;
        RECT  4.885 15.355 5.02 15.42 ;
        RECT  5.16 15.885 5.295 15.95 ;
        RECT  5.435 17.24 5.57 17.305 ;
        RECT  4.61 16.71 4.745 16.775 ;
        RECT  4.885 18.045 5.02 18.11 ;
        RECT  4.61 18.575 4.745 18.64 ;
        RECT  3.7425 20.1525 3.8075 20.435 ;
        RECT  3.7425 19.09 3.8075 19.27 ;
        RECT  3.1925 20.1525 3.2575 20.435 ;
        RECT  3.5725 20.1525 3.6375 20.435 ;
        RECT  3.1925 19.09 3.2575 19.3725 ;
        RECT  3.605 19.985 3.67 20.05 ;
        RECT  3.3825 19.985 3.4475 20.05 ;
        RECT  3.605 19.2375 3.67 20.0175 ;
        RECT  3.415 19.985 3.6375 20.05 ;
        RECT  3.3825 20.0175 3.4475 20.1525 ;
        RECT  3.125 20.0 3.16 20.065 ;
        RECT  3.6375 19.6875 3.875 19.7525 ;
        RECT  3.125 19.47 3.4 19.535 ;
        RECT  3.125 20.4025 3.875 20.4675 ;
        RECT  3.125 19.0575 3.875 19.1225 ;
        RECT  3.1925 19.2375 3.2575 19.3725 ;
        RECT  3.3825 19.2375 3.4475 19.3725 ;
        RECT  3.1925 19.3725 3.2575 19.5075 ;
        RECT  3.3825 19.3725 3.4475 19.5075 ;
        RECT  3.3825 19.2375 3.4475 19.3725 ;
        RECT  3.5725 19.2375 3.6375 19.3725 ;
        RECT  3.3825 19.3725 3.4475 19.5075 ;
        RECT  3.5725 19.3725 3.6375 19.5075 ;
        RECT  3.1925 20.1525 3.2575 20.2875 ;
        RECT  3.3825 20.1525 3.4475 20.2875 ;
        RECT  3.1925 20.1525 3.2575 20.2875 ;
        RECT  3.3825 20.1525 3.4475 20.2875 ;
        RECT  3.3825 20.1525 3.4475 20.2875 ;
        RECT  3.5725 20.1525 3.6375 20.2875 ;
        RECT  3.3825 20.1525 3.4475 20.2875 ;
        RECT  3.5725 20.1525 3.6375 20.2875 ;
        RECT  3.7425 20.1525 3.8075 20.2875 ;
        RECT  3.7425 19.2375 3.8075 19.3725 ;
        RECT  3.16 20.0 3.295 20.065 ;
        RECT  3.4 19.47 3.535 19.535 ;
        RECT  3.7425 20.435 3.8075 20.7175 ;
        RECT  3.7425 21.6 3.8075 21.78 ;
        RECT  3.1925 20.435 3.2575 20.7175 ;
        RECT  3.5725 20.435 3.6375 20.7175 ;
        RECT  3.1925 21.4975 3.2575 21.78 ;
        RECT  3.605 20.82 3.67 20.885 ;
        RECT  3.3825 20.82 3.4475 20.885 ;
        RECT  3.605 20.8525 3.67 21.6325 ;
        RECT  3.415 20.82 3.6375 20.885 ;
        RECT  3.3825 20.7175 3.4475 20.8525 ;
        RECT  3.125 20.805 3.16 20.87 ;
        RECT  3.6375 21.1175 3.875 21.1825 ;
        RECT  3.125 21.335 3.4 21.4 ;
        RECT  3.125 20.4025 3.875 20.4675 ;
        RECT  3.125 21.7475 3.875 21.8125 ;
        RECT  3.1925 21.2075 3.2575 21.3425 ;
        RECT  3.3825 21.2075 3.4475 21.3425 ;
        RECT  3.1925 21.3425 3.2575 21.4775 ;
        RECT  3.3825 21.3425 3.4475 21.4775 ;
        RECT  3.3825 21.2075 3.4475 21.3425 ;
        RECT  3.5725 21.2075 3.6375 21.3425 ;
        RECT  3.3825 21.3425 3.4475 21.4775 ;
        RECT  3.5725 21.3425 3.6375 21.4775 ;
        RECT  3.1925 20.8725 3.2575 21.0075 ;
        RECT  3.3825 20.8725 3.4475 21.0075 ;
        RECT  3.1925 20.8725 3.2575 21.0075 ;
        RECT  3.3825 20.8725 3.4475 21.0075 ;
        RECT  3.3825 20.8725 3.4475 21.0075 ;
        RECT  3.5725 20.8725 3.6375 21.0075 ;
        RECT  3.3825 20.8725 3.4475 21.0075 ;
        RECT  3.5725 20.8725 3.6375 21.0075 ;
        RECT  3.7425 20.7175 3.8075 20.8525 ;
        RECT  3.7425 21.6325 3.8075 21.7675 ;
        RECT  3.16 20.88 3.295 20.945 ;
        RECT  3.4 21.41 3.535 21.475 ;
        RECT  3.7425 22.8425 3.8075 23.125 ;
        RECT  3.7425 21.78 3.8075 21.96 ;
        RECT  3.1925 22.8425 3.2575 23.125 ;
        RECT  3.5725 22.8425 3.6375 23.125 ;
        RECT  3.1925 21.78 3.2575 22.0625 ;
        RECT  3.605 22.675 3.67 22.74 ;
        RECT  3.3825 22.675 3.4475 22.74 ;
        RECT  3.605 21.9275 3.67 22.7075 ;
        RECT  3.415 22.675 3.6375 22.74 ;
        RECT  3.3825 22.7075 3.4475 22.8425 ;
        RECT  3.125 22.69 3.16 22.755 ;
        RECT  3.6375 22.3775 3.875 22.4425 ;
        RECT  3.125 22.16 3.4 22.225 ;
        RECT  3.125 23.0925 3.875 23.1575 ;
        RECT  3.125 21.7475 3.875 21.8125 ;
        RECT  3.1925 21.9275 3.2575 22.0625 ;
        RECT  3.3825 21.9275 3.4475 22.0625 ;
        RECT  3.1925 22.0625 3.2575 22.1975 ;
        RECT  3.3825 22.0625 3.4475 22.1975 ;
        RECT  3.3825 21.9275 3.4475 22.0625 ;
        RECT  3.5725 21.9275 3.6375 22.0625 ;
        RECT  3.3825 22.0625 3.4475 22.1975 ;
        RECT  3.5725 22.0625 3.6375 22.1975 ;
        RECT  3.1925 22.8425 3.2575 22.9775 ;
        RECT  3.3825 22.8425 3.4475 22.9775 ;
        RECT  3.1925 22.8425 3.2575 22.9775 ;
        RECT  3.3825 22.8425 3.4475 22.9775 ;
        RECT  3.3825 22.8425 3.4475 22.9775 ;
        RECT  3.5725 22.8425 3.6375 22.9775 ;
        RECT  3.3825 22.8425 3.4475 22.9775 ;
        RECT  3.5725 22.8425 3.6375 22.9775 ;
        RECT  3.7425 22.8425 3.8075 22.9775 ;
        RECT  3.7425 21.9275 3.8075 22.0625 ;
        RECT  3.16 22.69 3.295 22.755 ;
        RECT  3.4 22.16 3.535 22.225 ;
        RECT  3.7425 23.125 3.8075 23.4075 ;
        RECT  3.7425 24.29 3.8075 24.47 ;
        RECT  3.1925 23.125 3.2575 23.4075 ;
        RECT  3.5725 23.125 3.6375 23.4075 ;
        RECT  3.1925 24.1875 3.2575 24.47 ;
        RECT  3.605 23.51 3.67 23.575 ;
        RECT  3.3825 23.51 3.4475 23.575 ;
        RECT  3.605 23.5425 3.67 24.3225 ;
        RECT  3.415 23.51 3.6375 23.575 ;
        RECT  3.3825 23.4075 3.4475 23.5425 ;
        RECT  3.125 23.495 3.16 23.56 ;
        RECT  3.6375 23.8075 3.875 23.8725 ;
        RECT  3.125 24.025 3.4 24.09 ;
        RECT  3.125 23.0925 3.875 23.1575 ;
        RECT  3.125 24.4375 3.875 24.5025 ;
        RECT  3.1925 23.8975 3.2575 24.0325 ;
        RECT  3.3825 23.8975 3.4475 24.0325 ;
        RECT  3.1925 24.0325 3.2575 24.1675 ;
        RECT  3.3825 24.0325 3.4475 24.1675 ;
        RECT  3.3825 23.8975 3.4475 24.0325 ;
        RECT  3.5725 23.8975 3.6375 24.0325 ;
        RECT  3.3825 24.0325 3.4475 24.1675 ;
        RECT  3.5725 24.0325 3.6375 24.1675 ;
        RECT  3.1925 23.5625 3.2575 23.6975 ;
        RECT  3.3825 23.5625 3.4475 23.6975 ;
        RECT  3.1925 23.5625 3.2575 23.6975 ;
        RECT  3.3825 23.5625 3.4475 23.6975 ;
        RECT  3.3825 23.5625 3.4475 23.6975 ;
        RECT  3.5725 23.5625 3.6375 23.6975 ;
        RECT  3.3825 23.5625 3.4475 23.6975 ;
        RECT  3.5725 23.5625 3.6375 23.6975 ;
        RECT  3.7425 23.4075 3.8075 23.5425 ;
        RECT  3.7425 24.3225 3.8075 24.4575 ;
        RECT  3.16 23.57 3.295 23.635 ;
        RECT  3.4 24.1 3.535 24.165 ;
        RECT  3.7425 25.5325 3.8075 25.815 ;
        RECT  3.7425 24.47 3.8075 24.65 ;
        RECT  3.1925 25.5325 3.2575 25.815 ;
        RECT  3.5725 25.5325 3.6375 25.815 ;
        RECT  3.1925 24.47 3.2575 24.7525 ;
        RECT  3.605 25.365 3.67 25.43 ;
        RECT  3.3825 25.365 3.4475 25.43 ;
        RECT  3.605 24.6175 3.67 25.3975 ;
        RECT  3.415 25.365 3.6375 25.43 ;
        RECT  3.3825 25.3975 3.4475 25.5325 ;
        RECT  3.125 25.38 3.16 25.445 ;
        RECT  3.6375 25.0675 3.875 25.1325 ;
        RECT  3.125 24.85 3.4 24.915 ;
        RECT  3.125 25.7825 3.875 25.8475 ;
        RECT  3.125 24.4375 3.875 24.5025 ;
        RECT  3.1925 24.6175 3.2575 24.7525 ;
        RECT  3.3825 24.6175 3.4475 24.7525 ;
        RECT  3.1925 24.7525 3.2575 24.8875 ;
        RECT  3.3825 24.7525 3.4475 24.8875 ;
        RECT  3.3825 24.6175 3.4475 24.7525 ;
        RECT  3.5725 24.6175 3.6375 24.7525 ;
        RECT  3.3825 24.7525 3.4475 24.8875 ;
        RECT  3.5725 24.7525 3.6375 24.8875 ;
        RECT  3.1925 25.5325 3.2575 25.6675 ;
        RECT  3.3825 25.5325 3.4475 25.6675 ;
        RECT  3.1925 25.5325 3.2575 25.6675 ;
        RECT  3.3825 25.5325 3.4475 25.6675 ;
        RECT  3.3825 25.5325 3.4475 25.6675 ;
        RECT  3.5725 25.5325 3.6375 25.6675 ;
        RECT  3.3825 25.5325 3.4475 25.6675 ;
        RECT  3.5725 25.5325 3.6375 25.6675 ;
        RECT  3.7425 25.5325 3.8075 25.6675 ;
        RECT  3.7425 24.6175 3.8075 24.7525 ;
        RECT  3.16 25.38 3.295 25.445 ;
        RECT  3.4 24.85 3.535 24.915 ;
        RECT  3.7425 25.815 3.8075 26.0975 ;
        RECT  3.7425 26.98 3.8075 27.16 ;
        RECT  3.1925 25.815 3.2575 26.0975 ;
        RECT  3.5725 25.815 3.6375 26.0975 ;
        RECT  3.1925 26.8775 3.2575 27.16 ;
        RECT  3.605 26.2 3.67 26.265 ;
        RECT  3.3825 26.2 3.4475 26.265 ;
        RECT  3.605 26.2325 3.67 27.0125 ;
        RECT  3.415 26.2 3.6375 26.265 ;
        RECT  3.3825 26.0975 3.4475 26.2325 ;
        RECT  3.125 26.185 3.16 26.25 ;
        RECT  3.6375 26.4975 3.875 26.5625 ;
        RECT  3.125 26.715 3.4 26.78 ;
        RECT  3.125 25.7825 3.875 25.8475 ;
        RECT  3.125 27.1275 3.875 27.1925 ;
        RECT  3.1925 26.5875 3.2575 26.7225 ;
        RECT  3.3825 26.5875 3.4475 26.7225 ;
        RECT  3.1925 26.7225 3.2575 26.8575 ;
        RECT  3.3825 26.7225 3.4475 26.8575 ;
        RECT  3.3825 26.5875 3.4475 26.7225 ;
        RECT  3.5725 26.5875 3.6375 26.7225 ;
        RECT  3.3825 26.7225 3.4475 26.8575 ;
        RECT  3.5725 26.7225 3.6375 26.8575 ;
        RECT  3.1925 26.2525 3.2575 26.3875 ;
        RECT  3.3825 26.2525 3.4475 26.3875 ;
        RECT  3.1925 26.2525 3.2575 26.3875 ;
        RECT  3.3825 26.2525 3.4475 26.3875 ;
        RECT  3.3825 26.2525 3.4475 26.3875 ;
        RECT  3.5725 26.2525 3.6375 26.3875 ;
        RECT  3.3825 26.2525 3.4475 26.3875 ;
        RECT  3.5725 26.2525 3.6375 26.3875 ;
        RECT  3.7425 26.0975 3.8075 26.2325 ;
        RECT  3.7425 27.0125 3.8075 27.1475 ;
        RECT  3.16 26.26 3.295 26.325 ;
        RECT  3.4 26.79 3.535 26.855 ;
        RECT  3.7425 28.2225 3.8075 28.505 ;
        RECT  3.7425 27.16 3.8075 27.34 ;
        RECT  3.1925 28.2225 3.2575 28.505 ;
        RECT  3.5725 28.2225 3.6375 28.505 ;
        RECT  3.1925 27.16 3.2575 27.4425 ;
        RECT  3.605 28.055 3.67 28.12 ;
        RECT  3.3825 28.055 3.4475 28.12 ;
        RECT  3.605 27.3075 3.67 28.0875 ;
        RECT  3.415 28.055 3.6375 28.12 ;
        RECT  3.3825 28.0875 3.4475 28.2225 ;
        RECT  3.125 28.07 3.16 28.135 ;
        RECT  3.6375 27.7575 3.875 27.8225 ;
        RECT  3.125 27.54 3.4 27.605 ;
        RECT  3.125 28.4725 3.875 28.5375 ;
        RECT  3.125 27.1275 3.875 27.1925 ;
        RECT  3.1925 27.3075 3.2575 27.4425 ;
        RECT  3.3825 27.3075 3.4475 27.4425 ;
        RECT  3.1925 27.4425 3.2575 27.5775 ;
        RECT  3.3825 27.4425 3.4475 27.5775 ;
        RECT  3.3825 27.3075 3.4475 27.4425 ;
        RECT  3.5725 27.3075 3.6375 27.4425 ;
        RECT  3.3825 27.4425 3.4475 27.5775 ;
        RECT  3.5725 27.4425 3.6375 27.5775 ;
        RECT  3.1925 28.2225 3.2575 28.3575 ;
        RECT  3.3825 28.2225 3.4475 28.3575 ;
        RECT  3.1925 28.2225 3.2575 28.3575 ;
        RECT  3.3825 28.2225 3.4475 28.3575 ;
        RECT  3.3825 28.2225 3.4475 28.3575 ;
        RECT  3.5725 28.2225 3.6375 28.3575 ;
        RECT  3.3825 28.2225 3.4475 28.3575 ;
        RECT  3.5725 28.2225 3.6375 28.3575 ;
        RECT  3.7425 28.2225 3.8075 28.3575 ;
        RECT  3.7425 27.3075 3.8075 27.4425 ;
        RECT  3.16 28.07 3.295 28.135 ;
        RECT  3.4 27.54 3.535 27.605 ;
        RECT  3.7425 28.505 3.8075 28.7875 ;
        RECT  3.7425 29.67 3.8075 29.85 ;
        RECT  3.1925 28.505 3.2575 28.7875 ;
        RECT  3.5725 28.505 3.6375 28.7875 ;
        RECT  3.1925 29.5675 3.2575 29.85 ;
        RECT  3.605 28.89 3.67 28.955 ;
        RECT  3.3825 28.89 3.4475 28.955 ;
        RECT  3.605 28.9225 3.67 29.7025 ;
        RECT  3.415 28.89 3.6375 28.955 ;
        RECT  3.3825 28.7875 3.4475 28.9225 ;
        RECT  3.125 28.875 3.16 28.94 ;
        RECT  3.6375 29.1875 3.875 29.2525 ;
        RECT  3.125 29.405 3.4 29.47 ;
        RECT  3.125 28.4725 3.875 28.5375 ;
        RECT  3.125 29.8175 3.875 29.8825 ;
        RECT  3.1925 29.2775 3.2575 29.4125 ;
        RECT  3.3825 29.2775 3.4475 29.4125 ;
        RECT  3.1925 29.4125 3.2575 29.5475 ;
        RECT  3.3825 29.4125 3.4475 29.5475 ;
        RECT  3.3825 29.2775 3.4475 29.4125 ;
        RECT  3.5725 29.2775 3.6375 29.4125 ;
        RECT  3.3825 29.4125 3.4475 29.5475 ;
        RECT  3.5725 29.4125 3.6375 29.5475 ;
        RECT  3.1925 28.9425 3.2575 29.0775 ;
        RECT  3.3825 28.9425 3.4475 29.0775 ;
        RECT  3.1925 28.9425 3.2575 29.0775 ;
        RECT  3.3825 28.9425 3.4475 29.0775 ;
        RECT  3.3825 28.9425 3.4475 29.0775 ;
        RECT  3.5725 28.9425 3.6375 29.0775 ;
        RECT  3.3825 28.9425 3.4475 29.0775 ;
        RECT  3.5725 28.9425 3.6375 29.0775 ;
        RECT  3.7425 28.7875 3.8075 28.9225 ;
        RECT  3.7425 29.7025 3.8075 29.8375 ;
        RECT  3.16 28.95 3.295 29.015 ;
        RECT  3.4 29.48 3.535 29.545 ;
        RECT  3.7425 30.9125 3.8075 31.195 ;
        RECT  3.7425 29.85 3.8075 30.03 ;
        RECT  3.1925 30.9125 3.2575 31.195 ;
        RECT  3.5725 30.9125 3.6375 31.195 ;
        RECT  3.1925 29.85 3.2575 30.1325 ;
        RECT  3.605 30.745 3.67 30.81 ;
        RECT  3.3825 30.745 3.4475 30.81 ;
        RECT  3.605 29.9975 3.67 30.7775 ;
        RECT  3.415 30.745 3.6375 30.81 ;
        RECT  3.3825 30.7775 3.4475 30.9125 ;
        RECT  3.125 30.76 3.16 30.825 ;
        RECT  3.6375 30.4475 3.875 30.5125 ;
        RECT  3.125 30.23 3.4 30.295 ;
        RECT  3.125 31.1625 3.875 31.2275 ;
        RECT  3.125 29.8175 3.875 29.8825 ;
        RECT  3.1925 29.9975 3.2575 30.1325 ;
        RECT  3.3825 29.9975 3.4475 30.1325 ;
        RECT  3.1925 30.1325 3.2575 30.2675 ;
        RECT  3.3825 30.1325 3.4475 30.2675 ;
        RECT  3.3825 29.9975 3.4475 30.1325 ;
        RECT  3.5725 29.9975 3.6375 30.1325 ;
        RECT  3.3825 30.1325 3.4475 30.2675 ;
        RECT  3.5725 30.1325 3.6375 30.2675 ;
        RECT  3.1925 30.9125 3.2575 31.0475 ;
        RECT  3.3825 30.9125 3.4475 31.0475 ;
        RECT  3.1925 30.9125 3.2575 31.0475 ;
        RECT  3.3825 30.9125 3.4475 31.0475 ;
        RECT  3.3825 30.9125 3.4475 31.0475 ;
        RECT  3.5725 30.9125 3.6375 31.0475 ;
        RECT  3.3825 30.9125 3.4475 31.0475 ;
        RECT  3.5725 30.9125 3.6375 31.0475 ;
        RECT  3.7425 30.9125 3.8075 31.0475 ;
        RECT  3.7425 29.9975 3.8075 30.1325 ;
        RECT  3.16 30.76 3.295 30.825 ;
        RECT  3.4 30.23 3.535 30.295 ;
        RECT  3.7425 31.195 3.8075 31.4775 ;
        RECT  3.7425 32.36 3.8075 32.54 ;
        RECT  3.1925 31.195 3.2575 31.4775 ;
        RECT  3.5725 31.195 3.6375 31.4775 ;
        RECT  3.1925 32.2575 3.2575 32.54 ;
        RECT  3.605 31.58 3.67 31.645 ;
        RECT  3.3825 31.58 3.4475 31.645 ;
        RECT  3.605 31.6125 3.67 32.3925 ;
        RECT  3.415 31.58 3.6375 31.645 ;
        RECT  3.3825 31.4775 3.4475 31.6125 ;
        RECT  3.125 31.565 3.16 31.63 ;
        RECT  3.6375 31.8775 3.875 31.9425 ;
        RECT  3.125 32.095 3.4 32.16 ;
        RECT  3.125 31.1625 3.875 31.2275 ;
        RECT  3.125 32.5075 3.875 32.5725 ;
        RECT  3.1925 31.9675 3.2575 32.1025 ;
        RECT  3.3825 31.9675 3.4475 32.1025 ;
        RECT  3.1925 32.1025 3.2575 32.2375 ;
        RECT  3.3825 32.1025 3.4475 32.2375 ;
        RECT  3.3825 31.9675 3.4475 32.1025 ;
        RECT  3.5725 31.9675 3.6375 32.1025 ;
        RECT  3.3825 32.1025 3.4475 32.2375 ;
        RECT  3.5725 32.1025 3.6375 32.2375 ;
        RECT  3.1925 31.6325 3.2575 31.7675 ;
        RECT  3.3825 31.6325 3.4475 31.7675 ;
        RECT  3.1925 31.6325 3.2575 31.7675 ;
        RECT  3.3825 31.6325 3.4475 31.7675 ;
        RECT  3.3825 31.6325 3.4475 31.7675 ;
        RECT  3.5725 31.6325 3.6375 31.7675 ;
        RECT  3.3825 31.6325 3.4475 31.7675 ;
        RECT  3.5725 31.6325 3.6375 31.7675 ;
        RECT  3.7425 31.4775 3.8075 31.6125 ;
        RECT  3.7425 32.3925 3.8075 32.5275 ;
        RECT  3.16 31.64 3.295 31.705 ;
        RECT  3.4 32.17 3.535 32.235 ;
        RECT  3.7425 33.6025 3.8075 33.885 ;
        RECT  3.7425 32.54 3.8075 32.72 ;
        RECT  3.1925 33.6025 3.2575 33.885 ;
        RECT  3.5725 33.6025 3.6375 33.885 ;
        RECT  3.1925 32.54 3.2575 32.8225 ;
        RECT  3.605 33.435 3.67 33.5 ;
        RECT  3.3825 33.435 3.4475 33.5 ;
        RECT  3.605 32.6875 3.67 33.4675 ;
        RECT  3.415 33.435 3.6375 33.5 ;
        RECT  3.3825 33.4675 3.4475 33.6025 ;
        RECT  3.125 33.45 3.16 33.515 ;
        RECT  3.6375 33.1375 3.875 33.2025 ;
        RECT  3.125 32.92 3.4 32.985 ;
        RECT  3.125 33.8525 3.875 33.9175 ;
        RECT  3.125 32.5075 3.875 32.5725 ;
        RECT  3.1925 32.6875 3.2575 32.8225 ;
        RECT  3.3825 32.6875 3.4475 32.8225 ;
        RECT  3.1925 32.8225 3.2575 32.9575 ;
        RECT  3.3825 32.8225 3.4475 32.9575 ;
        RECT  3.3825 32.6875 3.4475 32.8225 ;
        RECT  3.5725 32.6875 3.6375 32.8225 ;
        RECT  3.3825 32.8225 3.4475 32.9575 ;
        RECT  3.5725 32.8225 3.6375 32.9575 ;
        RECT  3.1925 33.6025 3.2575 33.7375 ;
        RECT  3.3825 33.6025 3.4475 33.7375 ;
        RECT  3.1925 33.6025 3.2575 33.7375 ;
        RECT  3.3825 33.6025 3.4475 33.7375 ;
        RECT  3.3825 33.6025 3.4475 33.7375 ;
        RECT  3.5725 33.6025 3.6375 33.7375 ;
        RECT  3.3825 33.6025 3.4475 33.7375 ;
        RECT  3.5725 33.6025 3.6375 33.7375 ;
        RECT  3.7425 33.6025 3.8075 33.7375 ;
        RECT  3.7425 32.6875 3.8075 32.8225 ;
        RECT  3.16 33.45 3.295 33.515 ;
        RECT  3.4 32.92 3.535 32.985 ;
        RECT  3.7425 33.885 3.8075 34.1675 ;
        RECT  3.7425 35.05 3.8075 35.23 ;
        RECT  3.1925 33.885 3.2575 34.1675 ;
        RECT  3.5725 33.885 3.6375 34.1675 ;
        RECT  3.1925 34.9475 3.2575 35.23 ;
        RECT  3.605 34.27 3.67 34.335 ;
        RECT  3.3825 34.27 3.4475 34.335 ;
        RECT  3.605 34.3025 3.67 35.0825 ;
        RECT  3.415 34.27 3.6375 34.335 ;
        RECT  3.3825 34.1675 3.4475 34.3025 ;
        RECT  3.125 34.255 3.16 34.32 ;
        RECT  3.6375 34.5675 3.875 34.6325 ;
        RECT  3.125 34.785 3.4 34.85 ;
        RECT  3.125 33.8525 3.875 33.9175 ;
        RECT  3.125 35.1975 3.875 35.2625 ;
        RECT  3.1925 34.6575 3.2575 34.7925 ;
        RECT  3.3825 34.6575 3.4475 34.7925 ;
        RECT  3.1925 34.7925 3.2575 34.9275 ;
        RECT  3.3825 34.7925 3.4475 34.9275 ;
        RECT  3.3825 34.6575 3.4475 34.7925 ;
        RECT  3.5725 34.6575 3.6375 34.7925 ;
        RECT  3.3825 34.7925 3.4475 34.9275 ;
        RECT  3.5725 34.7925 3.6375 34.9275 ;
        RECT  3.1925 34.3225 3.2575 34.4575 ;
        RECT  3.3825 34.3225 3.4475 34.4575 ;
        RECT  3.1925 34.3225 3.2575 34.4575 ;
        RECT  3.3825 34.3225 3.4475 34.4575 ;
        RECT  3.3825 34.3225 3.4475 34.4575 ;
        RECT  3.5725 34.3225 3.6375 34.4575 ;
        RECT  3.3825 34.3225 3.4475 34.4575 ;
        RECT  3.5725 34.3225 3.6375 34.4575 ;
        RECT  3.7425 34.1675 3.8075 34.3025 ;
        RECT  3.7425 35.0825 3.8075 35.2175 ;
        RECT  3.16 34.33 3.295 34.395 ;
        RECT  3.4 34.86 3.535 34.925 ;
        RECT  3.7425 36.2925 3.8075 36.575 ;
        RECT  3.7425 35.23 3.8075 35.41 ;
        RECT  3.1925 36.2925 3.2575 36.575 ;
        RECT  3.5725 36.2925 3.6375 36.575 ;
        RECT  3.1925 35.23 3.2575 35.5125 ;
        RECT  3.605 36.125 3.67 36.19 ;
        RECT  3.3825 36.125 3.4475 36.19 ;
        RECT  3.605 35.3775 3.67 36.1575 ;
        RECT  3.415 36.125 3.6375 36.19 ;
        RECT  3.3825 36.1575 3.4475 36.2925 ;
        RECT  3.125 36.14 3.16 36.205 ;
        RECT  3.6375 35.8275 3.875 35.8925 ;
        RECT  3.125 35.61 3.4 35.675 ;
        RECT  3.125 36.5425 3.875 36.6075 ;
        RECT  3.125 35.1975 3.875 35.2625 ;
        RECT  3.1925 35.3775 3.2575 35.5125 ;
        RECT  3.3825 35.3775 3.4475 35.5125 ;
        RECT  3.1925 35.5125 3.2575 35.6475 ;
        RECT  3.3825 35.5125 3.4475 35.6475 ;
        RECT  3.3825 35.3775 3.4475 35.5125 ;
        RECT  3.5725 35.3775 3.6375 35.5125 ;
        RECT  3.3825 35.5125 3.4475 35.6475 ;
        RECT  3.5725 35.5125 3.6375 35.6475 ;
        RECT  3.1925 36.2925 3.2575 36.4275 ;
        RECT  3.3825 36.2925 3.4475 36.4275 ;
        RECT  3.1925 36.2925 3.2575 36.4275 ;
        RECT  3.3825 36.2925 3.4475 36.4275 ;
        RECT  3.3825 36.2925 3.4475 36.4275 ;
        RECT  3.5725 36.2925 3.6375 36.4275 ;
        RECT  3.3825 36.2925 3.4475 36.4275 ;
        RECT  3.5725 36.2925 3.6375 36.4275 ;
        RECT  3.7425 36.2925 3.8075 36.4275 ;
        RECT  3.7425 35.3775 3.8075 35.5125 ;
        RECT  3.16 36.14 3.295 36.205 ;
        RECT  3.4 35.61 3.535 35.675 ;
        RECT  3.7425 36.575 3.8075 36.8575 ;
        RECT  3.7425 37.74 3.8075 37.92 ;
        RECT  3.1925 36.575 3.2575 36.8575 ;
        RECT  3.5725 36.575 3.6375 36.8575 ;
        RECT  3.1925 37.6375 3.2575 37.92 ;
        RECT  3.605 36.96 3.67 37.025 ;
        RECT  3.3825 36.96 3.4475 37.025 ;
        RECT  3.605 36.9925 3.67 37.7725 ;
        RECT  3.415 36.96 3.6375 37.025 ;
        RECT  3.3825 36.8575 3.4475 36.9925 ;
        RECT  3.125 36.945 3.16 37.01 ;
        RECT  3.6375 37.2575 3.875 37.3225 ;
        RECT  3.125 37.475 3.4 37.54 ;
        RECT  3.125 36.5425 3.875 36.6075 ;
        RECT  3.125 37.8875 3.875 37.9525 ;
        RECT  3.1925 37.3475 3.2575 37.4825 ;
        RECT  3.3825 37.3475 3.4475 37.4825 ;
        RECT  3.1925 37.4825 3.2575 37.6175 ;
        RECT  3.3825 37.4825 3.4475 37.6175 ;
        RECT  3.3825 37.3475 3.4475 37.4825 ;
        RECT  3.5725 37.3475 3.6375 37.4825 ;
        RECT  3.3825 37.4825 3.4475 37.6175 ;
        RECT  3.5725 37.4825 3.6375 37.6175 ;
        RECT  3.1925 37.0125 3.2575 37.1475 ;
        RECT  3.3825 37.0125 3.4475 37.1475 ;
        RECT  3.1925 37.0125 3.2575 37.1475 ;
        RECT  3.3825 37.0125 3.4475 37.1475 ;
        RECT  3.3825 37.0125 3.4475 37.1475 ;
        RECT  3.5725 37.0125 3.6375 37.1475 ;
        RECT  3.3825 37.0125 3.4475 37.1475 ;
        RECT  3.5725 37.0125 3.6375 37.1475 ;
        RECT  3.7425 36.8575 3.8075 36.9925 ;
        RECT  3.7425 37.7725 3.8075 37.9075 ;
        RECT  3.16 37.02 3.295 37.085 ;
        RECT  3.4 37.55 3.535 37.615 ;
        RECT  3.7425 38.9825 3.8075 39.265 ;
        RECT  3.7425 37.92 3.8075 38.1 ;
        RECT  3.1925 38.9825 3.2575 39.265 ;
        RECT  3.5725 38.9825 3.6375 39.265 ;
        RECT  3.1925 37.92 3.2575 38.2025 ;
        RECT  3.605 38.815 3.67 38.88 ;
        RECT  3.3825 38.815 3.4475 38.88 ;
        RECT  3.605 38.0675 3.67 38.8475 ;
        RECT  3.415 38.815 3.6375 38.88 ;
        RECT  3.3825 38.8475 3.4475 38.9825 ;
        RECT  3.125 38.83 3.16 38.895 ;
        RECT  3.6375 38.5175 3.875 38.5825 ;
        RECT  3.125 38.3 3.4 38.365 ;
        RECT  3.125 39.2325 3.875 39.2975 ;
        RECT  3.125 37.8875 3.875 37.9525 ;
        RECT  3.1925 38.0675 3.2575 38.2025 ;
        RECT  3.3825 38.0675 3.4475 38.2025 ;
        RECT  3.1925 38.2025 3.2575 38.3375 ;
        RECT  3.3825 38.2025 3.4475 38.3375 ;
        RECT  3.3825 38.0675 3.4475 38.2025 ;
        RECT  3.5725 38.0675 3.6375 38.2025 ;
        RECT  3.3825 38.2025 3.4475 38.3375 ;
        RECT  3.5725 38.2025 3.6375 38.3375 ;
        RECT  3.1925 38.9825 3.2575 39.1175 ;
        RECT  3.3825 38.9825 3.4475 39.1175 ;
        RECT  3.1925 38.9825 3.2575 39.1175 ;
        RECT  3.3825 38.9825 3.4475 39.1175 ;
        RECT  3.3825 38.9825 3.4475 39.1175 ;
        RECT  3.5725 38.9825 3.6375 39.1175 ;
        RECT  3.3825 38.9825 3.4475 39.1175 ;
        RECT  3.5725 38.9825 3.6375 39.1175 ;
        RECT  3.7425 38.9825 3.8075 39.1175 ;
        RECT  3.7425 38.0675 3.8075 38.2025 ;
        RECT  3.16 38.83 3.295 38.895 ;
        RECT  3.4 38.3 3.535 38.365 ;
        RECT  3.7425 39.265 3.8075 39.5475 ;
        RECT  3.7425 40.43 3.8075 40.61 ;
        RECT  3.1925 39.265 3.2575 39.5475 ;
        RECT  3.5725 39.265 3.6375 39.5475 ;
        RECT  3.1925 40.3275 3.2575 40.61 ;
        RECT  3.605 39.65 3.67 39.715 ;
        RECT  3.3825 39.65 3.4475 39.715 ;
        RECT  3.605 39.6825 3.67 40.4625 ;
        RECT  3.415 39.65 3.6375 39.715 ;
        RECT  3.3825 39.5475 3.4475 39.6825 ;
        RECT  3.125 39.635 3.16 39.7 ;
        RECT  3.6375 39.9475 3.875 40.0125 ;
        RECT  3.125 40.165 3.4 40.23 ;
        RECT  3.125 39.2325 3.875 39.2975 ;
        RECT  3.125 40.5775 3.875 40.6425 ;
        RECT  3.1925 40.0375 3.2575 40.1725 ;
        RECT  3.3825 40.0375 3.4475 40.1725 ;
        RECT  3.1925 40.1725 3.2575 40.3075 ;
        RECT  3.3825 40.1725 3.4475 40.3075 ;
        RECT  3.3825 40.0375 3.4475 40.1725 ;
        RECT  3.5725 40.0375 3.6375 40.1725 ;
        RECT  3.3825 40.1725 3.4475 40.3075 ;
        RECT  3.5725 40.1725 3.6375 40.3075 ;
        RECT  3.1925 39.7025 3.2575 39.8375 ;
        RECT  3.3825 39.7025 3.4475 39.8375 ;
        RECT  3.1925 39.7025 3.2575 39.8375 ;
        RECT  3.3825 39.7025 3.4475 39.8375 ;
        RECT  3.3825 39.7025 3.4475 39.8375 ;
        RECT  3.5725 39.7025 3.6375 39.8375 ;
        RECT  3.3825 39.7025 3.4475 39.8375 ;
        RECT  3.5725 39.7025 3.6375 39.8375 ;
        RECT  3.7425 39.5475 3.8075 39.6825 ;
        RECT  3.7425 40.4625 3.8075 40.5975 ;
        RECT  3.16 39.71 3.295 39.775 ;
        RECT  3.4 40.24 3.535 40.305 ;
        RECT  4.3025 20.0375 4.3675 20.4025 ;
        RECT  4.3025 19.1225 4.3675 19.2575 ;
        RECT  3.9425 19.1225 4.0075 19.1925 ;
        RECT  3.9425 20.3125 4.0075 20.4025 ;
        RECT  4.1325 19.225 4.1975 20.1725 ;
        RECT  3.875 19.64 3.91 19.705 ;
        RECT  4.1975 19.64 4.435 19.705 ;
        RECT  3.875 20.4025 4.435 20.4675 ;
        RECT  3.875 19.0575 4.435 19.1225 ;
        RECT  3.9425 19.1925 4.0075 19.3275 ;
        RECT  4.1325 19.1925 4.1975 19.3275 ;
        RECT  3.9425 19.3275 4.0075 19.4625 ;
        RECT  4.1325 19.3275 4.1975 19.4625 ;
        RECT  3.9425 20.0375 4.0075 20.3125 ;
        RECT  4.1325 20.0375 4.1975 20.3125 ;
        RECT  3.9425 20.0375 4.0075 20.3125 ;
        RECT  4.1325 20.0375 4.1975 20.3125 ;
        RECT  4.3025 20.0375 4.3675 20.3125 ;
        RECT  4.3025 19.1925 4.3675 19.3275 ;
        RECT  3.91 19.64 4.045 19.705 ;
        RECT  4.3025 20.4675 4.3675 20.8325 ;
        RECT  4.3025 21.6125 4.3675 21.7475 ;
        RECT  3.9425 21.6775 4.0075 21.7475 ;
        RECT  3.9425 20.4675 4.0075 20.5575 ;
        RECT  4.1325 20.6975 4.1975 21.645 ;
        RECT  3.875 21.165 3.91 21.23 ;
        RECT  4.1975 21.165 4.435 21.23 ;
        RECT  3.875 20.4025 4.435 20.4675 ;
        RECT  3.875 21.7475 4.435 21.8125 ;
        RECT  3.9425 21.3425 4.0075 21.4775 ;
        RECT  4.1325 21.3425 4.1975 21.4775 ;
        RECT  3.9425 21.4775 4.0075 21.6125 ;
        RECT  4.1325 21.4775 4.1975 21.6125 ;
        RECT  3.9425 20.9375 4.0075 21.2125 ;
        RECT  4.1325 20.9375 4.1975 21.2125 ;
        RECT  3.9425 20.9375 4.0075 21.2125 ;
        RECT  4.1325 20.9375 4.1975 21.2125 ;
        RECT  4.3025 20.8325 4.3675 21.1075 ;
        RECT  4.3025 21.6775 4.3675 21.8125 ;
        RECT  3.91 21.24 4.045 21.305 ;
        RECT  4.3025 22.7275 4.3675 23.0925 ;
        RECT  4.3025 21.8125 4.3675 21.9475 ;
        RECT  3.9425 21.8125 4.0075 21.8825 ;
        RECT  3.9425 23.0025 4.0075 23.0925 ;
        RECT  4.1325 21.915 4.1975 22.8625 ;
        RECT  3.875 22.33 3.91 22.395 ;
        RECT  4.1975 22.33 4.435 22.395 ;
        RECT  3.875 23.0925 4.435 23.1575 ;
        RECT  3.875 21.7475 4.435 21.8125 ;
        RECT  3.9425 21.8825 4.0075 22.0175 ;
        RECT  4.1325 21.8825 4.1975 22.0175 ;
        RECT  3.9425 22.0175 4.0075 22.1525 ;
        RECT  4.1325 22.0175 4.1975 22.1525 ;
        RECT  3.9425 22.7275 4.0075 23.0025 ;
        RECT  4.1325 22.7275 4.1975 23.0025 ;
        RECT  3.9425 22.7275 4.0075 23.0025 ;
        RECT  4.1325 22.7275 4.1975 23.0025 ;
        RECT  4.3025 22.7275 4.3675 23.0025 ;
        RECT  4.3025 21.8825 4.3675 22.0175 ;
        RECT  3.91 22.33 4.045 22.395 ;
        RECT  4.3025 23.1575 4.3675 23.5225 ;
        RECT  4.3025 24.3025 4.3675 24.4375 ;
        RECT  3.9425 24.3675 4.0075 24.4375 ;
        RECT  3.9425 23.1575 4.0075 23.2475 ;
        RECT  4.1325 23.3875 4.1975 24.335 ;
        RECT  3.875 23.855 3.91 23.92 ;
        RECT  4.1975 23.855 4.435 23.92 ;
        RECT  3.875 23.0925 4.435 23.1575 ;
        RECT  3.875 24.4375 4.435 24.5025 ;
        RECT  3.9425 24.0325 4.0075 24.1675 ;
        RECT  4.1325 24.0325 4.1975 24.1675 ;
        RECT  3.9425 24.1675 4.0075 24.3025 ;
        RECT  4.1325 24.1675 4.1975 24.3025 ;
        RECT  3.9425 23.6275 4.0075 23.9025 ;
        RECT  4.1325 23.6275 4.1975 23.9025 ;
        RECT  3.9425 23.6275 4.0075 23.9025 ;
        RECT  4.1325 23.6275 4.1975 23.9025 ;
        RECT  4.3025 23.5225 4.3675 23.7975 ;
        RECT  4.3025 24.3675 4.3675 24.5025 ;
        RECT  3.91 23.93 4.045 23.995 ;
        RECT  4.3025 25.4175 4.3675 25.7825 ;
        RECT  4.3025 24.5025 4.3675 24.6375 ;
        RECT  3.9425 24.5025 4.0075 24.5725 ;
        RECT  3.9425 25.6925 4.0075 25.7825 ;
        RECT  4.1325 24.605 4.1975 25.5525 ;
        RECT  3.875 25.02 3.91 25.085 ;
        RECT  4.1975 25.02 4.435 25.085 ;
        RECT  3.875 25.7825 4.435 25.8475 ;
        RECT  3.875 24.4375 4.435 24.5025 ;
        RECT  3.9425 24.5725 4.0075 24.7075 ;
        RECT  4.1325 24.5725 4.1975 24.7075 ;
        RECT  3.9425 24.7075 4.0075 24.8425 ;
        RECT  4.1325 24.7075 4.1975 24.8425 ;
        RECT  3.9425 25.4175 4.0075 25.6925 ;
        RECT  4.1325 25.4175 4.1975 25.6925 ;
        RECT  3.9425 25.4175 4.0075 25.6925 ;
        RECT  4.1325 25.4175 4.1975 25.6925 ;
        RECT  4.3025 25.4175 4.3675 25.6925 ;
        RECT  4.3025 24.5725 4.3675 24.7075 ;
        RECT  3.91 25.02 4.045 25.085 ;
        RECT  4.3025 25.8475 4.3675 26.2125 ;
        RECT  4.3025 26.9925 4.3675 27.1275 ;
        RECT  3.9425 27.0575 4.0075 27.1275 ;
        RECT  3.9425 25.8475 4.0075 25.9375 ;
        RECT  4.1325 26.0775 4.1975 27.025 ;
        RECT  3.875 26.545 3.91 26.61 ;
        RECT  4.1975 26.545 4.435 26.61 ;
        RECT  3.875 25.7825 4.435 25.8475 ;
        RECT  3.875 27.1275 4.435 27.1925 ;
        RECT  3.9425 26.7225 4.0075 26.8575 ;
        RECT  4.1325 26.7225 4.1975 26.8575 ;
        RECT  3.9425 26.8575 4.0075 26.9925 ;
        RECT  4.1325 26.8575 4.1975 26.9925 ;
        RECT  3.9425 26.3175 4.0075 26.5925 ;
        RECT  4.1325 26.3175 4.1975 26.5925 ;
        RECT  3.9425 26.3175 4.0075 26.5925 ;
        RECT  4.1325 26.3175 4.1975 26.5925 ;
        RECT  4.3025 26.2125 4.3675 26.4875 ;
        RECT  4.3025 27.0575 4.3675 27.1925 ;
        RECT  3.91 26.62 4.045 26.685 ;
        RECT  4.3025 28.1075 4.3675 28.4725 ;
        RECT  4.3025 27.1925 4.3675 27.3275 ;
        RECT  3.9425 27.1925 4.0075 27.2625 ;
        RECT  3.9425 28.3825 4.0075 28.4725 ;
        RECT  4.1325 27.295 4.1975 28.2425 ;
        RECT  3.875 27.71 3.91 27.775 ;
        RECT  4.1975 27.71 4.435 27.775 ;
        RECT  3.875 28.4725 4.435 28.5375 ;
        RECT  3.875 27.1275 4.435 27.1925 ;
        RECT  3.9425 27.2625 4.0075 27.3975 ;
        RECT  4.1325 27.2625 4.1975 27.3975 ;
        RECT  3.9425 27.3975 4.0075 27.5325 ;
        RECT  4.1325 27.3975 4.1975 27.5325 ;
        RECT  3.9425 28.1075 4.0075 28.3825 ;
        RECT  4.1325 28.1075 4.1975 28.3825 ;
        RECT  3.9425 28.1075 4.0075 28.3825 ;
        RECT  4.1325 28.1075 4.1975 28.3825 ;
        RECT  4.3025 28.1075 4.3675 28.3825 ;
        RECT  4.3025 27.2625 4.3675 27.3975 ;
        RECT  3.91 27.71 4.045 27.775 ;
        RECT  4.3025 28.5375 4.3675 28.9025 ;
        RECT  4.3025 29.6825 4.3675 29.8175 ;
        RECT  3.9425 29.7475 4.0075 29.8175 ;
        RECT  3.9425 28.5375 4.0075 28.6275 ;
        RECT  4.1325 28.7675 4.1975 29.715 ;
        RECT  3.875 29.235 3.91 29.3 ;
        RECT  4.1975 29.235 4.435 29.3 ;
        RECT  3.875 28.4725 4.435 28.5375 ;
        RECT  3.875 29.8175 4.435 29.8825 ;
        RECT  3.9425 29.4125 4.0075 29.5475 ;
        RECT  4.1325 29.4125 4.1975 29.5475 ;
        RECT  3.9425 29.5475 4.0075 29.6825 ;
        RECT  4.1325 29.5475 4.1975 29.6825 ;
        RECT  3.9425 29.0075 4.0075 29.2825 ;
        RECT  4.1325 29.0075 4.1975 29.2825 ;
        RECT  3.9425 29.0075 4.0075 29.2825 ;
        RECT  4.1325 29.0075 4.1975 29.2825 ;
        RECT  4.3025 28.9025 4.3675 29.1775 ;
        RECT  4.3025 29.7475 4.3675 29.8825 ;
        RECT  3.91 29.31 4.045 29.375 ;
        RECT  4.3025 30.7975 4.3675 31.1625 ;
        RECT  4.3025 29.8825 4.3675 30.0175 ;
        RECT  3.9425 29.8825 4.0075 29.9525 ;
        RECT  3.9425 31.0725 4.0075 31.1625 ;
        RECT  4.1325 29.985 4.1975 30.9325 ;
        RECT  3.875 30.4 3.91 30.465 ;
        RECT  4.1975 30.4 4.435 30.465 ;
        RECT  3.875 31.1625 4.435 31.2275 ;
        RECT  3.875 29.8175 4.435 29.8825 ;
        RECT  3.9425 29.9525 4.0075 30.0875 ;
        RECT  4.1325 29.9525 4.1975 30.0875 ;
        RECT  3.9425 30.0875 4.0075 30.2225 ;
        RECT  4.1325 30.0875 4.1975 30.2225 ;
        RECT  3.9425 30.7975 4.0075 31.0725 ;
        RECT  4.1325 30.7975 4.1975 31.0725 ;
        RECT  3.9425 30.7975 4.0075 31.0725 ;
        RECT  4.1325 30.7975 4.1975 31.0725 ;
        RECT  4.3025 30.7975 4.3675 31.0725 ;
        RECT  4.3025 29.9525 4.3675 30.0875 ;
        RECT  3.91 30.4 4.045 30.465 ;
        RECT  4.3025 31.2275 4.3675 31.5925 ;
        RECT  4.3025 32.3725 4.3675 32.5075 ;
        RECT  3.9425 32.4375 4.0075 32.5075 ;
        RECT  3.9425 31.2275 4.0075 31.3175 ;
        RECT  4.1325 31.4575 4.1975 32.405 ;
        RECT  3.875 31.925 3.91 31.99 ;
        RECT  4.1975 31.925 4.435 31.99 ;
        RECT  3.875 31.1625 4.435 31.2275 ;
        RECT  3.875 32.5075 4.435 32.5725 ;
        RECT  3.9425 32.1025 4.0075 32.2375 ;
        RECT  4.1325 32.1025 4.1975 32.2375 ;
        RECT  3.9425 32.2375 4.0075 32.3725 ;
        RECT  4.1325 32.2375 4.1975 32.3725 ;
        RECT  3.9425 31.6975 4.0075 31.9725 ;
        RECT  4.1325 31.6975 4.1975 31.9725 ;
        RECT  3.9425 31.6975 4.0075 31.9725 ;
        RECT  4.1325 31.6975 4.1975 31.9725 ;
        RECT  4.3025 31.5925 4.3675 31.8675 ;
        RECT  4.3025 32.4375 4.3675 32.5725 ;
        RECT  3.91 32.0 4.045 32.065 ;
        RECT  4.3025 33.4875 4.3675 33.8525 ;
        RECT  4.3025 32.5725 4.3675 32.7075 ;
        RECT  3.9425 32.5725 4.0075 32.6425 ;
        RECT  3.9425 33.7625 4.0075 33.8525 ;
        RECT  4.1325 32.675 4.1975 33.6225 ;
        RECT  3.875 33.09 3.91 33.155 ;
        RECT  4.1975 33.09 4.435 33.155 ;
        RECT  3.875 33.8525 4.435 33.9175 ;
        RECT  3.875 32.5075 4.435 32.5725 ;
        RECT  3.9425 32.6425 4.0075 32.7775 ;
        RECT  4.1325 32.6425 4.1975 32.7775 ;
        RECT  3.9425 32.7775 4.0075 32.9125 ;
        RECT  4.1325 32.7775 4.1975 32.9125 ;
        RECT  3.9425 33.4875 4.0075 33.7625 ;
        RECT  4.1325 33.4875 4.1975 33.7625 ;
        RECT  3.9425 33.4875 4.0075 33.7625 ;
        RECT  4.1325 33.4875 4.1975 33.7625 ;
        RECT  4.3025 33.4875 4.3675 33.7625 ;
        RECT  4.3025 32.6425 4.3675 32.7775 ;
        RECT  3.91 33.09 4.045 33.155 ;
        RECT  4.3025 33.9175 4.3675 34.2825 ;
        RECT  4.3025 35.0625 4.3675 35.1975 ;
        RECT  3.9425 35.1275 4.0075 35.1975 ;
        RECT  3.9425 33.9175 4.0075 34.0075 ;
        RECT  4.1325 34.1475 4.1975 35.095 ;
        RECT  3.875 34.615 3.91 34.68 ;
        RECT  4.1975 34.615 4.435 34.68 ;
        RECT  3.875 33.8525 4.435 33.9175 ;
        RECT  3.875 35.1975 4.435 35.2625 ;
        RECT  3.9425 34.7925 4.0075 34.9275 ;
        RECT  4.1325 34.7925 4.1975 34.9275 ;
        RECT  3.9425 34.9275 4.0075 35.0625 ;
        RECT  4.1325 34.9275 4.1975 35.0625 ;
        RECT  3.9425 34.3875 4.0075 34.6625 ;
        RECT  4.1325 34.3875 4.1975 34.6625 ;
        RECT  3.9425 34.3875 4.0075 34.6625 ;
        RECT  4.1325 34.3875 4.1975 34.6625 ;
        RECT  4.3025 34.2825 4.3675 34.5575 ;
        RECT  4.3025 35.1275 4.3675 35.2625 ;
        RECT  3.91 34.69 4.045 34.755 ;
        RECT  4.3025 36.1775 4.3675 36.5425 ;
        RECT  4.3025 35.2625 4.3675 35.3975 ;
        RECT  3.9425 35.2625 4.0075 35.3325 ;
        RECT  3.9425 36.4525 4.0075 36.5425 ;
        RECT  4.1325 35.365 4.1975 36.3125 ;
        RECT  3.875 35.78 3.91 35.845 ;
        RECT  4.1975 35.78 4.435 35.845 ;
        RECT  3.875 36.5425 4.435 36.6075 ;
        RECT  3.875 35.1975 4.435 35.2625 ;
        RECT  3.9425 35.3325 4.0075 35.4675 ;
        RECT  4.1325 35.3325 4.1975 35.4675 ;
        RECT  3.9425 35.4675 4.0075 35.6025 ;
        RECT  4.1325 35.4675 4.1975 35.6025 ;
        RECT  3.9425 36.1775 4.0075 36.4525 ;
        RECT  4.1325 36.1775 4.1975 36.4525 ;
        RECT  3.9425 36.1775 4.0075 36.4525 ;
        RECT  4.1325 36.1775 4.1975 36.4525 ;
        RECT  4.3025 36.1775 4.3675 36.4525 ;
        RECT  4.3025 35.3325 4.3675 35.4675 ;
        RECT  3.91 35.78 4.045 35.845 ;
        RECT  4.3025 36.6075 4.3675 36.9725 ;
        RECT  4.3025 37.7525 4.3675 37.8875 ;
        RECT  3.9425 37.8175 4.0075 37.8875 ;
        RECT  3.9425 36.6075 4.0075 36.6975 ;
        RECT  4.1325 36.8375 4.1975 37.785 ;
        RECT  3.875 37.305 3.91 37.37 ;
        RECT  4.1975 37.305 4.435 37.37 ;
        RECT  3.875 36.5425 4.435 36.6075 ;
        RECT  3.875 37.8875 4.435 37.9525 ;
        RECT  3.9425 37.4825 4.0075 37.6175 ;
        RECT  4.1325 37.4825 4.1975 37.6175 ;
        RECT  3.9425 37.6175 4.0075 37.7525 ;
        RECT  4.1325 37.6175 4.1975 37.7525 ;
        RECT  3.9425 37.0775 4.0075 37.3525 ;
        RECT  4.1325 37.0775 4.1975 37.3525 ;
        RECT  3.9425 37.0775 4.0075 37.3525 ;
        RECT  4.1325 37.0775 4.1975 37.3525 ;
        RECT  4.3025 36.9725 4.3675 37.2475 ;
        RECT  4.3025 37.8175 4.3675 37.9525 ;
        RECT  3.91 37.38 4.045 37.445 ;
        RECT  4.3025 38.8675 4.3675 39.2325 ;
        RECT  4.3025 37.9525 4.3675 38.0875 ;
        RECT  3.9425 37.9525 4.0075 38.0225 ;
        RECT  3.9425 39.1425 4.0075 39.2325 ;
        RECT  4.1325 38.055 4.1975 39.0025 ;
        RECT  3.875 38.47 3.91 38.535 ;
        RECT  4.1975 38.47 4.435 38.535 ;
        RECT  3.875 39.2325 4.435 39.2975 ;
        RECT  3.875 37.8875 4.435 37.9525 ;
        RECT  3.9425 38.0225 4.0075 38.1575 ;
        RECT  4.1325 38.0225 4.1975 38.1575 ;
        RECT  3.9425 38.1575 4.0075 38.2925 ;
        RECT  4.1325 38.1575 4.1975 38.2925 ;
        RECT  3.9425 38.8675 4.0075 39.1425 ;
        RECT  4.1325 38.8675 4.1975 39.1425 ;
        RECT  3.9425 38.8675 4.0075 39.1425 ;
        RECT  4.1325 38.8675 4.1975 39.1425 ;
        RECT  4.3025 38.8675 4.3675 39.1425 ;
        RECT  4.3025 38.0225 4.3675 38.1575 ;
        RECT  3.91 38.47 4.045 38.535 ;
        RECT  4.3025 39.2975 4.3675 39.6625 ;
        RECT  4.3025 40.4425 4.3675 40.5775 ;
        RECT  3.9425 40.5075 4.0075 40.5775 ;
        RECT  3.9425 39.2975 4.0075 39.3875 ;
        RECT  4.1325 39.5275 4.1975 40.475 ;
        RECT  3.875 39.995 3.91 40.06 ;
        RECT  4.1975 39.995 4.435 40.06 ;
        RECT  3.875 39.2325 4.435 39.2975 ;
        RECT  3.875 40.5775 4.435 40.6425 ;
        RECT  3.9425 40.1725 4.0075 40.3075 ;
        RECT  4.1325 40.1725 4.1975 40.3075 ;
        RECT  3.9425 40.3075 4.0075 40.4425 ;
        RECT  4.1325 40.3075 4.1975 40.4425 ;
        RECT  3.9425 39.7675 4.0075 40.0425 ;
        RECT  4.1325 39.7675 4.1975 40.0425 ;
        RECT  3.9425 39.7675 4.0075 40.0425 ;
        RECT  4.1325 39.7675 4.1975 40.0425 ;
        RECT  4.3025 39.6625 4.3675 39.9375 ;
        RECT  4.3025 40.5075 4.3675 40.6425 ;
        RECT  3.91 40.07 4.045 40.135 ;
        RECT  1.695 8.88 1.83 8.945 ;
        RECT  1.87 10.405 2.005 10.47 ;
        RECT  2.045 11.57 2.18 11.635 ;
        RECT  2.22 13.095 2.355 13.16 ;
        RECT  2.395 14.26 2.53 14.325 ;
        RECT  2.57 15.785 2.705 15.85 ;
        RECT  2.745 16.95 2.88 17.015 ;
        RECT  2.92 18.475 3.055 18.54 ;
        RECT  1.695 20.0 1.83 20.065 ;
        RECT  2.395 19.47 2.53 19.535 ;
        RECT  1.695 20.805 1.83 20.87 ;
        RECT  2.57 21.335 2.705 21.4 ;
        RECT  1.695 22.69 1.83 22.755 ;
        RECT  2.745 22.16 2.88 22.225 ;
        RECT  1.695 23.495 1.83 23.56 ;
        RECT  2.92 24.025 3.055 24.09 ;
        RECT  1.87 25.38 2.005 25.445 ;
        RECT  2.395 24.85 2.53 24.915 ;
        RECT  1.87 26.185 2.005 26.25 ;
        RECT  2.57 26.715 2.705 26.78 ;
        RECT  1.87 28.07 2.005 28.135 ;
        RECT  2.745 27.54 2.88 27.605 ;
        RECT  1.87 28.875 2.005 28.94 ;
        RECT  2.92 29.405 3.055 29.47 ;
        RECT  2.045 30.76 2.18 30.825 ;
        RECT  2.395 30.23 2.53 30.295 ;
        RECT  2.045 31.565 2.18 31.63 ;
        RECT  2.57 32.095 2.705 32.16 ;
        RECT  2.045 33.45 2.18 33.515 ;
        RECT  2.745 32.92 2.88 32.985 ;
        RECT  2.045 34.255 2.18 34.32 ;
        RECT  2.92 34.785 3.055 34.85 ;
        RECT  2.22 36.14 2.355 36.205 ;
        RECT  2.395 35.61 2.53 35.675 ;
        RECT  2.22 36.945 2.355 37.01 ;
        RECT  2.57 37.475 2.705 37.54 ;
        RECT  2.22 38.83 2.355 38.895 ;
        RECT  2.745 38.3 2.88 38.365 ;
        RECT  2.22 39.635 2.355 39.7 ;
        RECT  2.92 40.165 3.055 40.23 ;
        RECT  4.665 19.64 4.89 19.705 ;
        RECT  5.4175 19.64 5.4825 19.705 ;
        RECT  5.4175 19.47 5.4825 19.535 ;
        RECT  5.2125 19.64 5.45 19.705 ;
        RECT  5.4175 19.5025 5.4825 19.6725 ;
        RECT  5.45 19.47 5.725 19.535 ;
        RECT  6.1675 19.6875 6.2325 19.7525 ;
        RECT  6.1675 19.64 6.2325 19.705 ;
        RECT  5.9625 19.6875 6.2 19.7525 ;
        RECT  6.1675 19.6725 6.2325 19.72 ;
        RECT  6.2 19.64 6.235 19.705 ;
        RECT  4.665 21.165 4.89 21.23 ;
        RECT  5.4175 21.165 5.4825 21.23 ;
        RECT  5.4175 21.335 5.4825 21.4 ;
        RECT  5.2125 21.165 5.45 21.23 ;
        RECT  5.4175 21.1975 5.4825 21.3675 ;
        RECT  5.45 21.335 5.725 21.4 ;
        RECT  6.1675 21.1175 6.2325 21.1825 ;
        RECT  6.1675 21.165 6.2325 21.23 ;
        RECT  5.9625 21.1175 6.2 21.1825 ;
        RECT  6.1675 21.15 6.2325 21.1975 ;
        RECT  6.2 21.165 6.235 21.23 ;
        RECT  4.665 22.33 4.89 22.395 ;
        RECT  5.4175 22.33 5.4825 22.395 ;
        RECT  5.4175 22.16 5.4825 22.225 ;
        RECT  5.2125 22.33 5.45 22.395 ;
        RECT  5.4175 22.1925 5.4825 22.3625 ;
        RECT  5.45 22.16 5.725 22.225 ;
        RECT  6.1675 22.3775 6.2325 22.4425 ;
        RECT  6.1675 22.33 6.2325 22.395 ;
        RECT  5.9625 22.3775 6.2 22.4425 ;
        RECT  6.1675 22.3625 6.2325 22.41 ;
        RECT  6.2 22.33 6.235 22.395 ;
        RECT  4.665 23.855 4.89 23.92 ;
        RECT  5.4175 23.855 5.4825 23.92 ;
        RECT  5.4175 24.025 5.4825 24.09 ;
        RECT  5.2125 23.855 5.45 23.92 ;
        RECT  5.4175 23.8875 5.4825 24.0575 ;
        RECT  5.45 24.025 5.725 24.09 ;
        RECT  6.1675 23.8075 6.2325 23.8725 ;
        RECT  6.1675 23.855 6.2325 23.92 ;
        RECT  5.9625 23.8075 6.2 23.8725 ;
        RECT  6.1675 23.84 6.2325 23.8875 ;
        RECT  6.2 23.855 6.235 23.92 ;
        RECT  4.665 25.02 4.89 25.085 ;
        RECT  5.4175 25.02 5.4825 25.085 ;
        RECT  5.4175 24.85 5.4825 24.915 ;
        RECT  5.2125 25.02 5.45 25.085 ;
        RECT  5.4175 24.8825 5.4825 25.0525 ;
        RECT  5.45 24.85 5.725 24.915 ;
        RECT  6.1675 25.0675 6.2325 25.1325 ;
        RECT  6.1675 25.02 6.2325 25.085 ;
        RECT  5.9625 25.0675 6.2 25.1325 ;
        RECT  6.1675 25.0525 6.2325 25.1 ;
        RECT  6.2 25.02 6.235 25.085 ;
        RECT  4.665 26.545 4.89 26.61 ;
        RECT  5.4175 26.545 5.4825 26.61 ;
        RECT  5.4175 26.715 5.4825 26.78 ;
        RECT  5.2125 26.545 5.45 26.61 ;
        RECT  5.4175 26.5775 5.4825 26.7475 ;
        RECT  5.45 26.715 5.725 26.78 ;
        RECT  6.1675 26.4975 6.2325 26.5625 ;
        RECT  6.1675 26.545 6.2325 26.61 ;
        RECT  5.9625 26.4975 6.2 26.5625 ;
        RECT  6.1675 26.53 6.2325 26.5775 ;
        RECT  6.2 26.545 6.235 26.61 ;
        RECT  4.665 27.71 4.89 27.775 ;
        RECT  5.4175 27.71 5.4825 27.775 ;
        RECT  5.4175 27.54 5.4825 27.605 ;
        RECT  5.2125 27.71 5.45 27.775 ;
        RECT  5.4175 27.5725 5.4825 27.7425 ;
        RECT  5.45 27.54 5.725 27.605 ;
        RECT  6.1675 27.7575 6.2325 27.8225 ;
        RECT  6.1675 27.71 6.2325 27.775 ;
        RECT  5.9625 27.7575 6.2 27.8225 ;
        RECT  6.1675 27.7425 6.2325 27.79 ;
        RECT  6.2 27.71 6.235 27.775 ;
        RECT  4.665 29.235 4.89 29.3 ;
        RECT  5.4175 29.235 5.4825 29.3 ;
        RECT  5.4175 29.405 5.4825 29.47 ;
        RECT  5.2125 29.235 5.45 29.3 ;
        RECT  5.4175 29.2675 5.4825 29.4375 ;
        RECT  5.45 29.405 5.725 29.47 ;
        RECT  6.1675 29.1875 6.2325 29.2525 ;
        RECT  6.1675 29.235 6.2325 29.3 ;
        RECT  5.9625 29.1875 6.2 29.2525 ;
        RECT  6.1675 29.22 6.2325 29.2675 ;
        RECT  6.2 29.235 6.235 29.3 ;
        RECT  4.665 30.4 4.89 30.465 ;
        RECT  5.4175 30.4 5.4825 30.465 ;
        RECT  5.4175 30.23 5.4825 30.295 ;
        RECT  5.2125 30.4 5.45 30.465 ;
        RECT  5.4175 30.2625 5.4825 30.4325 ;
        RECT  5.45 30.23 5.725 30.295 ;
        RECT  6.1675 30.4475 6.2325 30.5125 ;
        RECT  6.1675 30.4 6.2325 30.465 ;
        RECT  5.9625 30.4475 6.2 30.5125 ;
        RECT  6.1675 30.4325 6.2325 30.48 ;
        RECT  6.2 30.4 6.235 30.465 ;
        RECT  4.665 31.925 4.89 31.99 ;
        RECT  5.4175 31.925 5.4825 31.99 ;
        RECT  5.4175 32.095 5.4825 32.16 ;
        RECT  5.2125 31.925 5.45 31.99 ;
        RECT  5.4175 31.9575 5.4825 32.1275 ;
        RECT  5.45 32.095 5.725 32.16 ;
        RECT  6.1675 31.8775 6.2325 31.9425 ;
        RECT  6.1675 31.925 6.2325 31.99 ;
        RECT  5.9625 31.8775 6.2 31.9425 ;
        RECT  6.1675 31.91 6.2325 31.9575 ;
        RECT  6.2 31.925 6.235 31.99 ;
        RECT  4.665 33.09 4.89 33.155 ;
        RECT  5.4175 33.09 5.4825 33.155 ;
        RECT  5.4175 32.92 5.4825 32.985 ;
        RECT  5.2125 33.09 5.45 33.155 ;
        RECT  5.4175 32.9525 5.4825 33.1225 ;
        RECT  5.45 32.92 5.725 32.985 ;
        RECT  6.1675 33.1375 6.2325 33.2025 ;
        RECT  6.1675 33.09 6.2325 33.155 ;
        RECT  5.9625 33.1375 6.2 33.2025 ;
        RECT  6.1675 33.1225 6.2325 33.17 ;
        RECT  6.2 33.09 6.235 33.155 ;
        RECT  4.665 34.615 4.89 34.68 ;
        RECT  5.4175 34.615 5.4825 34.68 ;
        RECT  5.4175 34.785 5.4825 34.85 ;
        RECT  5.2125 34.615 5.45 34.68 ;
        RECT  5.4175 34.6475 5.4825 34.8175 ;
        RECT  5.45 34.785 5.725 34.85 ;
        RECT  6.1675 34.5675 6.2325 34.6325 ;
        RECT  6.1675 34.615 6.2325 34.68 ;
        RECT  5.9625 34.5675 6.2 34.6325 ;
        RECT  6.1675 34.6 6.2325 34.6475 ;
        RECT  6.2 34.615 6.235 34.68 ;
        RECT  4.665 35.78 4.89 35.845 ;
        RECT  5.4175 35.78 5.4825 35.845 ;
        RECT  5.4175 35.61 5.4825 35.675 ;
        RECT  5.2125 35.78 5.45 35.845 ;
        RECT  5.4175 35.6425 5.4825 35.8125 ;
        RECT  5.45 35.61 5.725 35.675 ;
        RECT  6.1675 35.8275 6.2325 35.8925 ;
        RECT  6.1675 35.78 6.2325 35.845 ;
        RECT  5.9625 35.8275 6.2 35.8925 ;
        RECT  6.1675 35.8125 6.2325 35.86 ;
        RECT  6.2 35.78 6.235 35.845 ;
        RECT  4.665 37.305 4.89 37.37 ;
        RECT  5.4175 37.305 5.4825 37.37 ;
        RECT  5.4175 37.475 5.4825 37.54 ;
        RECT  5.2125 37.305 5.45 37.37 ;
        RECT  5.4175 37.3375 5.4825 37.5075 ;
        RECT  5.45 37.475 5.725 37.54 ;
        RECT  6.1675 37.2575 6.2325 37.3225 ;
        RECT  6.1675 37.305 6.2325 37.37 ;
        RECT  5.9625 37.2575 6.2 37.3225 ;
        RECT  6.1675 37.29 6.2325 37.3375 ;
        RECT  6.2 37.305 6.235 37.37 ;
        RECT  4.665 38.47 4.89 38.535 ;
        RECT  5.4175 38.47 5.4825 38.535 ;
        RECT  5.4175 38.3 5.4825 38.365 ;
        RECT  5.2125 38.47 5.45 38.535 ;
        RECT  5.4175 38.3325 5.4825 38.5025 ;
        RECT  5.45 38.3 5.725 38.365 ;
        RECT  6.1675 38.5175 6.2325 38.5825 ;
        RECT  6.1675 38.47 6.2325 38.535 ;
        RECT  5.9625 38.5175 6.2 38.5825 ;
        RECT  6.1675 38.5025 6.2325 38.55 ;
        RECT  6.2 38.47 6.235 38.535 ;
        RECT  4.665 39.995 4.89 40.06 ;
        RECT  5.4175 39.995 5.4825 40.06 ;
        RECT  5.4175 40.165 5.4825 40.23 ;
        RECT  5.2125 39.995 5.45 40.06 ;
        RECT  5.4175 40.0275 5.4825 40.1975 ;
        RECT  5.45 40.165 5.725 40.23 ;
        RECT  6.1675 39.9475 6.2325 40.0125 ;
        RECT  6.1675 39.995 6.2325 40.06 ;
        RECT  5.9625 39.9475 6.2 40.0125 ;
        RECT  6.1675 39.98 6.2325 40.0275 ;
        RECT  6.2 39.995 6.235 40.06 ;
        RECT  6.695 25.02 6.76 25.085 ;
        RECT  4.435 23.495 4.805 23.56 ;
        RECT  6.695 19.64 6.76 19.705 ;
        RECT  4.435 28.875 4.805 28.94 ;
        RECT  6.695 22.33 6.76 22.395 ;
        RECT  4.435 20.805 4.805 20.87 ;
        RECT  4.435 26.185 4.805 26.25 ;
        RECT  4.435 30.76 4.805 30.825 ;
        RECT  6.695 39.995 6.76 40.06 ;
        RECT  4.435 33.45 4.805 33.515 ;
        RECT  6.695 30.4 6.76 30.465 ;
        RECT  4.435 38.83 4.805 38.895 ;
        RECT  4.435 36.14 4.805 36.205 ;
        RECT  6.695 27.71 6.76 27.775 ;
        RECT  6.695 37.305 6.76 37.37 ;
        RECT  6.695 34.615 6.76 34.68 ;
        RECT  6.695 23.855 6.76 23.92 ;
        RECT  4.435 22.69 4.805 22.755 ;
        RECT  6.695 26.545 6.76 26.61 ;
        RECT  6.695 21.165 6.76 21.23 ;
        RECT  4.435 20.0 4.805 20.065 ;
        RECT  4.435 25.38 4.805 25.445 ;
        RECT  4.435 28.07 4.805 28.135 ;
        RECT  4.435 31.565 4.805 31.63 ;
        RECT  4.435 34.255 4.805 34.32 ;
        RECT  6.695 38.47 6.76 38.535 ;
        RECT  4.435 39.635 4.805 39.7 ;
        RECT  6.695 33.09 6.76 33.155 ;
        RECT  6.695 31.925 6.76 31.99 ;
        RECT  4.435 20.4025 4.89 20.4675 ;
        RECT  4.435 23.0925 4.89 23.1575 ;
        RECT  4.435 25.7825 4.89 25.8475 ;
        RECT  4.435 28.4725 4.89 28.5375 ;
        RECT  4.435 31.1625 4.89 31.2275 ;
        RECT  4.435 33.8525 4.89 33.9175 ;
        RECT  4.435 36.5425 4.89 36.6075 ;
        RECT  4.435 39.2325 4.89 39.2975 ;
        RECT  4.435 19.0575 4.89 19.1225 ;
        RECT  4.435 21.7475 4.89 21.8125 ;
        RECT  4.435 24.4375 4.89 24.5025 ;
        RECT  4.435 27.1275 4.89 27.1925 ;
        RECT  4.435 29.8175 4.89 29.8825 ;
        RECT  4.435 32.5075 4.89 32.5725 ;
        RECT  4.435 35.1975 4.89 35.2625 ;
        RECT  4.435 37.8875 4.89 37.9525 ;
        RECT  4.435 40.5775 4.89 40.6425 ;
        RECT  4.435 36.945 4.805 37.01 ;
        RECT  6.695 35.78 6.76 35.845 ;
        RECT  6.695 29.235 6.76 29.3 ;
        RECT  5.3175 20.0375 5.3825 20.4025 ;
        RECT  5.3175 19.1225 5.3825 19.2575 ;
        RECT  4.9575 19.1225 5.0225 19.1925 ;
        RECT  4.9575 20.3125 5.0225 20.4025 ;
        RECT  5.1475 19.225 5.2125 20.1725 ;
        RECT  4.89 19.64 4.925 19.705 ;
        RECT  5.2125 19.64 5.45 19.705 ;
        RECT  4.89 20.4025 5.45 20.4675 ;
        RECT  4.89 19.0575 5.45 19.1225 ;
        RECT  4.9575 19.1925 5.0225 19.3275 ;
        RECT  5.1475 19.1925 5.2125 19.3275 ;
        RECT  4.9575 19.3275 5.0225 19.4625 ;
        RECT  5.1475 19.3275 5.2125 19.4625 ;
        RECT  4.9575 20.0375 5.0225 20.3125 ;
        RECT  5.1475 20.0375 5.2125 20.3125 ;
        RECT  4.9575 20.0375 5.0225 20.3125 ;
        RECT  5.1475 20.0375 5.2125 20.3125 ;
        RECT  5.3175 20.0375 5.3825 20.3125 ;
        RECT  5.3175 19.1925 5.3825 19.3275 ;
        RECT  4.925 19.64 5.06 19.705 ;
        RECT  6.0675 20.1525 6.1325 20.435 ;
        RECT  6.0675 19.09 6.1325 19.27 ;
        RECT  5.5175 20.1525 5.5825 20.435 ;
        RECT  5.8975 20.1525 5.9625 20.435 ;
        RECT  5.5175 19.09 5.5825 19.3725 ;
        RECT  5.93 19.985 5.995 20.05 ;
        RECT  5.7075 19.985 5.7725 20.05 ;
        RECT  5.93 19.2375 5.995 20.0175 ;
        RECT  5.74 19.985 5.9625 20.05 ;
        RECT  5.7075 20.0175 5.7725 20.1525 ;
        RECT  5.45 20.0 5.485 20.065 ;
        RECT  5.9625 19.6875 6.2 19.7525 ;
        RECT  5.45 19.47 5.725 19.535 ;
        RECT  5.45 20.4025 6.2 20.4675 ;
        RECT  5.45 19.0575 6.2 19.1225 ;
        RECT  5.5175 19.2375 5.5825 19.3725 ;
        RECT  5.7075 19.2375 5.7725 19.3725 ;
        RECT  5.5175 19.3725 5.5825 19.5075 ;
        RECT  5.7075 19.3725 5.7725 19.5075 ;
        RECT  5.7075 19.2375 5.7725 19.3725 ;
        RECT  5.8975 19.2375 5.9625 19.3725 ;
        RECT  5.7075 19.3725 5.7725 19.5075 ;
        RECT  5.8975 19.3725 5.9625 19.5075 ;
        RECT  5.5175 20.1525 5.5825 20.2875 ;
        RECT  5.7075 20.1525 5.7725 20.2875 ;
        RECT  5.5175 20.1525 5.5825 20.2875 ;
        RECT  5.7075 20.1525 5.7725 20.2875 ;
        RECT  5.7075 20.1525 5.7725 20.2875 ;
        RECT  5.8975 20.1525 5.9625 20.2875 ;
        RECT  5.7075 20.1525 5.7725 20.2875 ;
        RECT  5.8975 20.1525 5.9625 20.2875 ;
        RECT  6.0675 20.1525 6.1325 20.2875 ;
        RECT  6.0675 19.2375 6.1325 19.3725 ;
        RECT  5.485 20.0 5.62 20.065 ;
        RECT  5.725 19.47 5.86 19.535 ;
        RECT  6.6275 20.0375 6.6925 20.4025 ;
        RECT  6.6275 19.1225 6.6925 19.2575 ;
        RECT  6.2675 19.1225 6.3325 19.1925 ;
        RECT  6.2675 20.3125 6.3325 20.4025 ;
        RECT  6.4575 19.225 6.5225 20.1725 ;
        RECT  6.2 19.64 6.235 19.705 ;
        RECT  6.5225 19.64 6.76 19.705 ;
        RECT  6.2 20.4025 6.76 20.4675 ;
        RECT  6.2 19.0575 6.76 19.1225 ;
        RECT  6.2675 19.1925 6.3325 19.3275 ;
        RECT  6.4575 19.1925 6.5225 19.3275 ;
        RECT  6.2675 19.3275 6.3325 19.4625 ;
        RECT  6.4575 19.3275 6.5225 19.4625 ;
        RECT  6.2675 20.0375 6.3325 20.3125 ;
        RECT  6.4575 20.0375 6.5225 20.3125 ;
        RECT  6.2675 20.0375 6.3325 20.3125 ;
        RECT  6.4575 20.0375 6.5225 20.3125 ;
        RECT  6.6275 20.0375 6.6925 20.3125 ;
        RECT  6.6275 19.1925 6.6925 19.3275 ;
        RECT  6.235 19.64 6.37 19.705 ;
        RECT  4.6325 19.605 4.6975 19.74 ;
        RECT  4.7725 19.965 4.8375 20.1 ;
        RECT  5.45 20.0 5.585 20.065 ;
        RECT  5.3175 20.4675 5.3825 20.8325 ;
        RECT  5.3175 21.6125 5.3825 21.7475 ;
        RECT  4.9575 21.6775 5.0225 21.7475 ;
        RECT  4.9575 20.4675 5.0225 20.5575 ;
        RECT  5.1475 20.6975 5.2125 21.645 ;
        RECT  4.89 21.165 4.925 21.23 ;
        RECT  5.2125 21.165 5.45 21.23 ;
        RECT  4.89 20.4025 5.45 20.4675 ;
        RECT  4.89 21.7475 5.45 21.8125 ;
        RECT  4.9575 21.3425 5.0225 21.4775 ;
        RECT  5.1475 21.3425 5.2125 21.4775 ;
        RECT  4.9575 21.4775 5.0225 21.6125 ;
        RECT  5.1475 21.4775 5.2125 21.6125 ;
        RECT  4.9575 20.9375 5.0225 21.2125 ;
        RECT  5.1475 20.9375 5.2125 21.2125 ;
        RECT  4.9575 20.9375 5.0225 21.2125 ;
        RECT  5.1475 20.9375 5.2125 21.2125 ;
        RECT  5.3175 20.8325 5.3825 21.1075 ;
        RECT  5.3175 21.6775 5.3825 21.8125 ;
        RECT  4.925 21.24 5.06 21.305 ;
        RECT  6.0675 20.435 6.1325 20.7175 ;
        RECT  6.0675 21.6 6.1325 21.78 ;
        RECT  5.5175 20.435 5.5825 20.7175 ;
        RECT  5.8975 20.435 5.9625 20.7175 ;
        RECT  5.5175 21.4975 5.5825 21.78 ;
        RECT  5.93 20.82 5.995 20.885 ;
        RECT  5.7075 20.82 5.7725 20.885 ;
        RECT  5.93 20.8525 5.995 21.6325 ;
        RECT  5.74 20.82 5.9625 20.885 ;
        RECT  5.7075 20.7175 5.7725 20.8525 ;
        RECT  5.45 20.805 5.485 20.87 ;
        RECT  5.9625 21.1175 6.2 21.1825 ;
        RECT  5.45 21.335 5.725 21.4 ;
        RECT  5.45 20.4025 6.2 20.4675 ;
        RECT  5.45 21.7475 6.2 21.8125 ;
        RECT  5.5175 21.2075 5.5825 21.3425 ;
        RECT  5.7075 21.2075 5.7725 21.3425 ;
        RECT  5.5175 21.3425 5.5825 21.4775 ;
        RECT  5.7075 21.3425 5.7725 21.4775 ;
        RECT  5.7075 21.2075 5.7725 21.3425 ;
        RECT  5.8975 21.2075 5.9625 21.3425 ;
        RECT  5.7075 21.3425 5.7725 21.4775 ;
        RECT  5.8975 21.3425 5.9625 21.4775 ;
        RECT  5.5175 20.8725 5.5825 21.0075 ;
        RECT  5.7075 20.8725 5.7725 21.0075 ;
        RECT  5.5175 20.8725 5.5825 21.0075 ;
        RECT  5.7075 20.8725 5.7725 21.0075 ;
        RECT  5.7075 20.8725 5.7725 21.0075 ;
        RECT  5.8975 20.8725 5.9625 21.0075 ;
        RECT  5.7075 20.8725 5.7725 21.0075 ;
        RECT  5.8975 20.8725 5.9625 21.0075 ;
        RECT  6.0675 20.7175 6.1325 20.8525 ;
        RECT  6.0675 21.6325 6.1325 21.7675 ;
        RECT  5.485 20.88 5.62 20.945 ;
        RECT  5.725 21.41 5.86 21.475 ;
        RECT  6.6275 20.4675 6.6925 20.8325 ;
        RECT  6.6275 21.6125 6.6925 21.7475 ;
        RECT  6.2675 21.6775 6.3325 21.7475 ;
        RECT  6.2675 20.4675 6.3325 20.5575 ;
        RECT  6.4575 20.6975 6.5225 21.645 ;
        RECT  6.2 21.165 6.235 21.23 ;
        RECT  6.5225 21.165 6.76 21.23 ;
        RECT  6.2 20.4025 6.76 20.4675 ;
        RECT  6.2 21.7475 6.76 21.8125 ;
        RECT  6.2675 21.3425 6.3325 21.4775 ;
        RECT  6.4575 21.3425 6.5225 21.4775 ;
        RECT  6.2675 21.4775 6.3325 21.6125 ;
        RECT  6.4575 21.4775 6.5225 21.6125 ;
        RECT  6.2675 20.9375 6.3325 21.2125 ;
        RECT  6.4575 20.9375 6.5225 21.2125 ;
        RECT  6.2675 20.9375 6.3325 21.2125 ;
        RECT  6.4575 20.9375 6.5225 21.2125 ;
        RECT  6.6275 20.8325 6.6925 21.1075 ;
        RECT  6.6275 21.6775 6.6925 21.8125 ;
        RECT  6.235 21.24 6.37 21.305 ;
        RECT  4.6325 21.13 4.6975 21.265 ;
        RECT  4.7725 20.77 4.8375 20.905 ;
        RECT  5.45 20.805 5.585 20.87 ;
        RECT  5.3175 22.7275 5.3825 23.0925 ;
        RECT  5.3175 21.8125 5.3825 21.9475 ;
        RECT  4.9575 21.8125 5.0225 21.8825 ;
        RECT  4.9575 23.0025 5.0225 23.0925 ;
        RECT  5.1475 21.915 5.2125 22.8625 ;
        RECT  4.89 22.33 4.925 22.395 ;
        RECT  5.2125 22.33 5.45 22.395 ;
        RECT  4.89 23.0925 5.45 23.1575 ;
        RECT  4.89 21.7475 5.45 21.8125 ;
        RECT  4.9575 21.8825 5.0225 22.0175 ;
        RECT  5.1475 21.8825 5.2125 22.0175 ;
        RECT  4.9575 22.0175 5.0225 22.1525 ;
        RECT  5.1475 22.0175 5.2125 22.1525 ;
        RECT  4.9575 22.7275 5.0225 23.0025 ;
        RECT  5.1475 22.7275 5.2125 23.0025 ;
        RECT  4.9575 22.7275 5.0225 23.0025 ;
        RECT  5.1475 22.7275 5.2125 23.0025 ;
        RECT  5.3175 22.7275 5.3825 23.0025 ;
        RECT  5.3175 21.8825 5.3825 22.0175 ;
        RECT  4.925 22.33 5.06 22.395 ;
        RECT  6.0675 22.8425 6.1325 23.125 ;
        RECT  6.0675 21.78 6.1325 21.96 ;
        RECT  5.5175 22.8425 5.5825 23.125 ;
        RECT  5.8975 22.8425 5.9625 23.125 ;
        RECT  5.5175 21.78 5.5825 22.0625 ;
        RECT  5.93 22.675 5.995 22.74 ;
        RECT  5.7075 22.675 5.7725 22.74 ;
        RECT  5.93 21.9275 5.995 22.7075 ;
        RECT  5.74 22.675 5.9625 22.74 ;
        RECT  5.7075 22.7075 5.7725 22.8425 ;
        RECT  5.45 22.69 5.485 22.755 ;
        RECT  5.9625 22.3775 6.2 22.4425 ;
        RECT  5.45 22.16 5.725 22.225 ;
        RECT  5.45 23.0925 6.2 23.1575 ;
        RECT  5.45 21.7475 6.2 21.8125 ;
        RECT  5.5175 21.9275 5.5825 22.0625 ;
        RECT  5.7075 21.9275 5.7725 22.0625 ;
        RECT  5.5175 22.0625 5.5825 22.1975 ;
        RECT  5.7075 22.0625 5.7725 22.1975 ;
        RECT  5.7075 21.9275 5.7725 22.0625 ;
        RECT  5.8975 21.9275 5.9625 22.0625 ;
        RECT  5.7075 22.0625 5.7725 22.1975 ;
        RECT  5.8975 22.0625 5.9625 22.1975 ;
        RECT  5.5175 22.8425 5.5825 22.9775 ;
        RECT  5.7075 22.8425 5.7725 22.9775 ;
        RECT  5.5175 22.8425 5.5825 22.9775 ;
        RECT  5.7075 22.8425 5.7725 22.9775 ;
        RECT  5.7075 22.8425 5.7725 22.9775 ;
        RECT  5.8975 22.8425 5.9625 22.9775 ;
        RECT  5.7075 22.8425 5.7725 22.9775 ;
        RECT  5.8975 22.8425 5.9625 22.9775 ;
        RECT  6.0675 22.8425 6.1325 22.9775 ;
        RECT  6.0675 21.9275 6.1325 22.0625 ;
        RECT  5.485 22.69 5.62 22.755 ;
        RECT  5.725 22.16 5.86 22.225 ;
        RECT  6.6275 22.7275 6.6925 23.0925 ;
        RECT  6.6275 21.8125 6.6925 21.9475 ;
        RECT  6.2675 21.8125 6.3325 21.8825 ;
        RECT  6.2675 23.0025 6.3325 23.0925 ;
        RECT  6.4575 21.915 6.5225 22.8625 ;
        RECT  6.2 22.33 6.235 22.395 ;
        RECT  6.5225 22.33 6.76 22.395 ;
        RECT  6.2 23.0925 6.76 23.1575 ;
        RECT  6.2 21.7475 6.76 21.8125 ;
        RECT  6.2675 21.8825 6.3325 22.0175 ;
        RECT  6.4575 21.8825 6.5225 22.0175 ;
        RECT  6.2675 22.0175 6.3325 22.1525 ;
        RECT  6.4575 22.0175 6.5225 22.1525 ;
        RECT  6.2675 22.7275 6.3325 23.0025 ;
        RECT  6.4575 22.7275 6.5225 23.0025 ;
        RECT  6.2675 22.7275 6.3325 23.0025 ;
        RECT  6.4575 22.7275 6.5225 23.0025 ;
        RECT  6.6275 22.7275 6.6925 23.0025 ;
        RECT  6.6275 21.8825 6.6925 22.0175 ;
        RECT  6.235 22.33 6.37 22.395 ;
        RECT  4.6325 22.295 4.6975 22.43 ;
        RECT  4.7725 22.655 4.8375 22.79 ;
        RECT  5.45 22.69 5.585 22.755 ;
        RECT  5.3175 23.1575 5.3825 23.5225 ;
        RECT  5.3175 24.3025 5.3825 24.4375 ;
        RECT  4.9575 24.3675 5.0225 24.4375 ;
        RECT  4.9575 23.1575 5.0225 23.2475 ;
        RECT  5.1475 23.3875 5.2125 24.335 ;
        RECT  4.89 23.855 4.925 23.92 ;
        RECT  5.2125 23.855 5.45 23.92 ;
        RECT  4.89 23.0925 5.45 23.1575 ;
        RECT  4.89 24.4375 5.45 24.5025 ;
        RECT  4.9575 24.0325 5.0225 24.1675 ;
        RECT  5.1475 24.0325 5.2125 24.1675 ;
        RECT  4.9575 24.1675 5.0225 24.3025 ;
        RECT  5.1475 24.1675 5.2125 24.3025 ;
        RECT  4.9575 23.6275 5.0225 23.9025 ;
        RECT  5.1475 23.6275 5.2125 23.9025 ;
        RECT  4.9575 23.6275 5.0225 23.9025 ;
        RECT  5.1475 23.6275 5.2125 23.9025 ;
        RECT  5.3175 23.5225 5.3825 23.7975 ;
        RECT  5.3175 24.3675 5.3825 24.5025 ;
        RECT  4.925 23.93 5.06 23.995 ;
        RECT  6.0675 23.125 6.1325 23.4075 ;
        RECT  6.0675 24.29 6.1325 24.47 ;
        RECT  5.5175 23.125 5.5825 23.4075 ;
        RECT  5.8975 23.125 5.9625 23.4075 ;
        RECT  5.5175 24.1875 5.5825 24.47 ;
        RECT  5.93 23.51 5.995 23.575 ;
        RECT  5.7075 23.51 5.7725 23.575 ;
        RECT  5.93 23.5425 5.995 24.3225 ;
        RECT  5.74 23.51 5.9625 23.575 ;
        RECT  5.7075 23.4075 5.7725 23.5425 ;
        RECT  5.45 23.495 5.485 23.56 ;
        RECT  5.9625 23.8075 6.2 23.8725 ;
        RECT  5.45 24.025 5.725 24.09 ;
        RECT  5.45 23.0925 6.2 23.1575 ;
        RECT  5.45 24.4375 6.2 24.5025 ;
        RECT  5.5175 23.8975 5.5825 24.0325 ;
        RECT  5.7075 23.8975 5.7725 24.0325 ;
        RECT  5.5175 24.0325 5.5825 24.1675 ;
        RECT  5.7075 24.0325 5.7725 24.1675 ;
        RECT  5.7075 23.8975 5.7725 24.0325 ;
        RECT  5.8975 23.8975 5.9625 24.0325 ;
        RECT  5.7075 24.0325 5.7725 24.1675 ;
        RECT  5.8975 24.0325 5.9625 24.1675 ;
        RECT  5.5175 23.5625 5.5825 23.6975 ;
        RECT  5.7075 23.5625 5.7725 23.6975 ;
        RECT  5.5175 23.5625 5.5825 23.6975 ;
        RECT  5.7075 23.5625 5.7725 23.6975 ;
        RECT  5.7075 23.5625 5.7725 23.6975 ;
        RECT  5.8975 23.5625 5.9625 23.6975 ;
        RECT  5.7075 23.5625 5.7725 23.6975 ;
        RECT  5.8975 23.5625 5.9625 23.6975 ;
        RECT  6.0675 23.4075 6.1325 23.5425 ;
        RECT  6.0675 24.3225 6.1325 24.4575 ;
        RECT  5.485 23.57 5.62 23.635 ;
        RECT  5.725 24.1 5.86 24.165 ;
        RECT  6.6275 23.1575 6.6925 23.5225 ;
        RECT  6.6275 24.3025 6.6925 24.4375 ;
        RECT  6.2675 24.3675 6.3325 24.4375 ;
        RECT  6.2675 23.1575 6.3325 23.2475 ;
        RECT  6.4575 23.3875 6.5225 24.335 ;
        RECT  6.2 23.855 6.235 23.92 ;
        RECT  6.5225 23.855 6.76 23.92 ;
        RECT  6.2 23.0925 6.76 23.1575 ;
        RECT  6.2 24.4375 6.76 24.5025 ;
        RECT  6.2675 24.0325 6.3325 24.1675 ;
        RECT  6.4575 24.0325 6.5225 24.1675 ;
        RECT  6.2675 24.1675 6.3325 24.3025 ;
        RECT  6.4575 24.1675 6.5225 24.3025 ;
        RECT  6.2675 23.6275 6.3325 23.9025 ;
        RECT  6.4575 23.6275 6.5225 23.9025 ;
        RECT  6.2675 23.6275 6.3325 23.9025 ;
        RECT  6.4575 23.6275 6.5225 23.9025 ;
        RECT  6.6275 23.5225 6.6925 23.7975 ;
        RECT  6.6275 24.3675 6.6925 24.5025 ;
        RECT  6.235 23.93 6.37 23.995 ;
        RECT  4.6325 23.82 4.6975 23.955 ;
        RECT  4.7725 23.46 4.8375 23.595 ;
        RECT  5.45 23.495 5.585 23.56 ;
        RECT  5.3175 25.4175 5.3825 25.7825 ;
        RECT  5.3175 24.5025 5.3825 24.6375 ;
        RECT  4.9575 24.5025 5.0225 24.5725 ;
        RECT  4.9575 25.6925 5.0225 25.7825 ;
        RECT  5.1475 24.605 5.2125 25.5525 ;
        RECT  4.89 25.02 4.925 25.085 ;
        RECT  5.2125 25.02 5.45 25.085 ;
        RECT  4.89 25.7825 5.45 25.8475 ;
        RECT  4.89 24.4375 5.45 24.5025 ;
        RECT  4.9575 24.5725 5.0225 24.7075 ;
        RECT  5.1475 24.5725 5.2125 24.7075 ;
        RECT  4.9575 24.7075 5.0225 24.8425 ;
        RECT  5.1475 24.7075 5.2125 24.8425 ;
        RECT  4.9575 25.4175 5.0225 25.6925 ;
        RECT  5.1475 25.4175 5.2125 25.6925 ;
        RECT  4.9575 25.4175 5.0225 25.6925 ;
        RECT  5.1475 25.4175 5.2125 25.6925 ;
        RECT  5.3175 25.4175 5.3825 25.6925 ;
        RECT  5.3175 24.5725 5.3825 24.7075 ;
        RECT  4.925 25.02 5.06 25.085 ;
        RECT  6.0675 25.5325 6.1325 25.815 ;
        RECT  6.0675 24.47 6.1325 24.65 ;
        RECT  5.5175 25.5325 5.5825 25.815 ;
        RECT  5.8975 25.5325 5.9625 25.815 ;
        RECT  5.5175 24.47 5.5825 24.7525 ;
        RECT  5.93 25.365 5.995 25.43 ;
        RECT  5.7075 25.365 5.7725 25.43 ;
        RECT  5.93 24.6175 5.995 25.3975 ;
        RECT  5.74 25.365 5.9625 25.43 ;
        RECT  5.7075 25.3975 5.7725 25.5325 ;
        RECT  5.45 25.38 5.485 25.445 ;
        RECT  5.9625 25.0675 6.2 25.1325 ;
        RECT  5.45 24.85 5.725 24.915 ;
        RECT  5.45 25.7825 6.2 25.8475 ;
        RECT  5.45 24.4375 6.2 24.5025 ;
        RECT  5.5175 24.6175 5.5825 24.7525 ;
        RECT  5.7075 24.6175 5.7725 24.7525 ;
        RECT  5.5175 24.7525 5.5825 24.8875 ;
        RECT  5.7075 24.7525 5.7725 24.8875 ;
        RECT  5.7075 24.6175 5.7725 24.7525 ;
        RECT  5.8975 24.6175 5.9625 24.7525 ;
        RECT  5.7075 24.7525 5.7725 24.8875 ;
        RECT  5.8975 24.7525 5.9625 24.8875 ;
        RECT  5.5175 25.5325 5.5825 25.6675 ;
        RECT  5.7075 25.5325 5.7725 25.6675 ;
        RECT  5.5175 25.5325 5.5825 25.6675 ;
        RECT  5.7075 25.5325 5.7725 25.6675 ;
        RECT  5.7075 25.5325 5.7725 25.6675 ;
        RECT  5.8975 25.5325 5.9625 25.6675 ;
        RECT  5.7075 25.5325 5.7725 25.6675 ;
        RECT  5.8975 25.5325 5.9625 25.6675 ;
        RECT  6.0675 25.5325 6.1325 25.6675 ;
        RECT  6.0675 24.6175 6.1325 24.7525 ;
        RECT  5.485 25.38 5.62 25.445 ;
        RECT  5.725 24.85 5.86 24.915 ;
        RECT  6.6275 25.4175 6.6925 25.7825 ;
        RECT  6.6275 24.5025 6.6925 24.6375 ;
        RECT  6.2675 24.5025 6.3325 24.5725 ;
        RECT  6.2675 25.6925 6.3325 25.7825 ;
        RECT  6.4575 24.605 6.5225 25.5525 ;
        RECT  6.2 25.02 6.235 25.085 ;
        RECT  6.5225 25.02 6.76 25.085 ;
        RECT  6.2 25.7825 6.76 25.8475 ;
        RECT  6.2 24.4375 6.76 24.5025 ;
        RECT  6.2675 24.5725 6.3325 24.7075 ;
        RECT  6.4575 24.5725 6.5225 24.7075 ;
        RECT  6.2675 24.7075 6.3325 24.8425 ;
        RECT  6.4575 24.7075 6.5225 24.8425 ;
        RECT  6.2675 25.4175 6.3325 25.6925 ;
        RECT  6.4575 25.4175 6.5225 25.6925 ;
        RECT  6.2675 25.4175 6.3325 25.6925 ;
        RECT  6.4575 25.4175 6.5225 25.6925 ;
        RECT  6.6275 25.4175 6.6925 25.6925 ;
        RECT  6.6275 24.5725 6.6925 24.7075 ;
        RECT  6.235 25.02 6.37 25.085 ;
        RECT  4.6325 24.985 4.6975 25.12 ;
        RECT  4.7725 25.345 4.8375 25.48 ;
        RECT  5.45 25.38 5.585 25.445 ;
        RECT  5.3175 25.8475 5.3825 26.2125 ;
        RECT  5.3175 26.9925 5.3825 27.1275 ;
        RECT  4.9575 27.0575 5.0225 27.1275 ;
        RECT  4.9575 25.8475 5.0225 25.9375 ;
        RECT  5.1475 26.0775 5.2125 27.025 ;
        RECT  4.89 26.545 4.925 26.61 ;
        RECT  5.2125 26.545 5.45 26.61 ;
        RECT  4.89 25.7825 5.45 25.8475 ;
        RECT  4.89 27.1275 5.45 27.1925 ;
        RECT  4.9575 26.7225 5.0225 26.8575 ;
        RECT  5.1475 26.7225 5.2125 26.8575 ;
        RECT  4.9575 26.8575 5.0225 26.9925 ;
        RECT  5.1475 26.8575 5.2125 26.9925 ;
        RECT  4.9575 26.3175 5.0225 26.5925 ;
        RECT  5.1475 26.3175 5.2125 26.5925 ;
        RECT  4.9575 26.3175 5.0225 26.5925 ;
        RECT  5.1475 26.3175 5.2125 26.5925 ;
        RECT  5.3175 26.2125 5.3825 26.4875 ;
        RECT  5.3175 27.0575 5.3825 27.1925 ;
        RECT  4.925 26.62 5.06 26.685 ;
        RECT  6.0675 25.815 6.1325 26.0975 ;
        RECT  6.0675 26.98 6.1325 27.16 ;
        RECT  5.5175 25.815 5.5825 26.0975 ;
        RECT  5.8975 25.815 5.9625 26.0975 ;
        RECT  5.5175 26.8775 5.5825 27.16 ;
        RECT  5.93 26.2 5.995 26.265 ;
        RECT  5.7075 26.2 5.7725 26.265 ;
        RECT  5.93 26.2325 5.995 27.0125 ;
        RECT  5.74 26.2 5.9625 26.265 ;
        RECT  5.7075 26.0975 5.7725 26.2325 ;
        RECT  5.45 26.185 5.485 26.25 ;
        RECT  5.9625 26.4975 6.2 26.5625 ;
        RECT  5.45 26.715 5.725 26.78 ;
        RECT  5.45 25.7825 6.2 25.8475 ;
        RECT  5.45 27.1275 6.2 27.1925 ;
        RECT  5.5175 26.5875 5.5825 26.7225 ;
        RECT  5.7075 26.5875 5.7725 26.7225 ;
        RECT  5.5175 26.7225 5.5825 26.8575 ;
        RECT  5.7075 26.7225 5.7725 26.8575 ;
        RECT  5.7075 26.5875 5.7725 26.7225 ;
        RECT  5.8975 26.5875 5.9625 26.7225 ;
        RECT  5.7075 26.7225 5.7725 26.8575 ;
        RECT  5.8975 26.7225 5.9625 26.8575 ;
        RECT  5.5175 26.2525 5.5825 26.3875 ;
        RECT  5.7075 26.2525 5.7725 26.3875 ;
        RECT  5.5175 26.2525 5.5825 26.3875 ;
        RECT  5.7075 26.2525 5.7725 26.3875 ;
        RECT  5.7075 26.2525 5.7725 26.3875 ;
        RECT  5.8975 26.2525 5.9625 26.3875 ;
        RECT  5.7075 26.2525 5.7725 26.3875 ;
        RECT  5.8975 26.2525 5.9625 26.3875 ;
        RECT  6.0675 26.0975 6.1325 26.2325 ;
        RECT  6.0675 27.0125 6.1325 27.1475 ;
        RECT  5.485 26.26 5.62 26.325 ;
        RECT  5.725 26.79 5.86 26.855 ;
        RECT  6.6275 25.8475 6.6925 26.2125 ;
        RECT  6.6275 26.9925 6.6925 27.1275 ;
        RECT  6.2675 27.0575 6.3325 27.1275 ;
        RECT  6.2675 25.8475 6.3325 25.9375 ;
        RECT  6.4575 26.0775 6.5225 27.025 ;
        RECT  6.2 26.545 6.235 26.61 ;
        RECT  6.5225 26.545 6.76 26.61 ;
        RECT  6.2 25.7825 6.76 25.8475 ;
        RECT  6.2 27.1275 6.76 27.1925 ;
        RECT  6.2675 26.7225 6.3325 26.8575 ;
        RECT  6.4575 26.7225 6.5225 26.8575 ;
        RECT  6.2675 26.8575 6.3325 26.9925 ;
        RECT  6.4575 26.8575 6.5225 26.9925 ;
        RECT  6.2675 26.3175 6.3325 26.5925 ;
        RECT  6.4575 26.3175 6.5225 26.5925 ;
        RECT  6.2675 26.3175 6.3325 26.5925 ;
        RECT  6.4575 26.3175 6.5225 26.5925 ;
        RECT  6.6275 26.2125 6.6925 26.4875 ;
        RECT  6.6275 27.0575 6.6925 27.1925 ;
        RECT  6.235 26.62 6.37 26.685 ;
        RECT  4.6325 26.51 4.6975 26.645 ;
        RECT  4.7725 26.15 4.8375 26.285 ;
        RECT  5.45 26.185 5.585 26.25 ;
        RECT  5.3175 28.1075 5.3825 28.4725 ;
        RECT  5.3175 27.1925 5.3825 27.3275 ;
        RECT  4.9575 27.1925 5.0225 27.2625 ;
        RECT  4.9575 28.3825 5.0225 28.4725 ;
        RECT  5.1475 27.295 5.2125 28.2425 ;
        RECT  4.89 27.71 4.925 27.775 ;
        RECT  5.2125 27.71 5.45 27.775 ;
        RECT  4.89 28.4725 5.45 28.5375 ;
        RECT  4.89 27.1275 5.45 27.1925 ;
        RECT  4.9575 27.2625 5.0225 27.3975 ;
        RECT  5.1475 27.2625 5.2125 27.3975 ;
        RECT  4.9575 27.3975 5.0225 27.5325 ;
        RECT  5.1475 27.3975 5.2125 27.5325 ;
        RECT  4.9575 28.1075 5.0225 28.3825 ;
        RECT  5.1475 28.1075 5.2125 28.3825 ;
        RECT  4.9575 28.1075 5.0225 28.3825 ;
        RECT  5.1475 28.1075 5.2125 28.3825 ;
        RECT  5.3175 28.1075 5.3825 28.3825 ;
        RECT  5.3175 27.2625 5.3825 27.3975 ;
        RECT  4.925 27.71 5.06 27.775 ;
        RECT  6.0675 28.2225 6.1325 28.505 ;
        RECT  6.0675 27.16 6.1325 27.34 ;
        RECT  5.5175 28.2225 5.5825 28.505 ;
        RECT  5.8975 28.2225 5.9625 28.505 ;
        RECT  5.5175 27.16 5.5825 27.4425 ;
        RECT  5.93 28.055 5.995 28.12 ;
        RECT  5.7075 28.055 5.7725 28.12 ;
        RECT  5.93 27.3075 5.995 28.0875 ;
        RECT  5.74 28.055 5.9625 28.12 ;
        RECT  5.7075 28.0875 5.7725 28.2225 ;
        RECT  5.45 28.07 5.485 28.135 ;
        RECT  5.9625 27.7575 6.2 27.8225 ;
        RECT  5.45 27.54 5.725 27.605 ;
        RECT  5.45 28.4725 6.2 28.5375 ;
        RECT  5.45 27.1275 6.2 27.1925 ;
        RECT  5.5175 27.3075 5.5825 27.4425 ;
        RECT  5.7075 27.3075 5.7725 27.4425 ;
        RECT  5.5175 27.4425 5.5825 27.5775 ;
        RECT  5.7075 27.4425 5.7725 27.5775 ;
        RECT  5.7075 27.3075 5.7725 27.4425 ;
        RECT  5.8975 27.3075 5.9625 27.4425 ;
        RECT  5.7075 27.4425 5.7725 27.5775 ;
        RECT  5.8975 27.4425 5.9625 27.5775 ;
        RECT  5.5175 28.2225 5.5825 28.3575 ;
        RECT  5.7075 28.2225 5.7725 28.3575 ;
        RECT  5.5175 28.2225 5.5825 28.3575 ;
        RECT  5.7075 28.2225 5.7725 28.3575 ;
        RECT  5.7075 28.2225 5.7725 28.3575 ;
        RECT  5.8975 28.2225 5.9625 28.3575 ;
        RECT  5.7075 28.2225 5.7725 28.3575 ;
        RECT  5.8975 28.2225 5.9625 28.3575 ;
        RECT  6.0675 28.2225 6.1325 28.3575 ;
        RECT  6.0675 27.3075 6.1325 27.4425 ;
        RECT  5.485 28.07 5.62 28.135 ;
        RECT  5.725 27.54 5.86 27.605 ;
        RECT  6.6275 28.1075 6.6925 28.4725 ;
        RECT  6.6275 27.1925 6.6925 27.3275 ;
        RECT  6.2675 27.1925 6.3325 27.2625 ;
        RECT  6.2675 28.3825 6.3325 28.4725 ;
        RECT  6.4575 27.295 6.5225 28.2425 ;
        RECT  6.2 27.71 6.235 27.775 ;
        RECT  6.5225 27.71 6.76 27.775 ;
        RECT  6.2 28.4725 6.76 28.5375 ;
        RECT  6.2 27.1275 6.76 27.1925 ;
        RECT  6.2675 27.2625 6.3325 27.3975 ;
        RECT  6.4575 27.2625 6.5225 27.3975 ;
        RECT  6.2675 27.3975 6.3325 27.5325 ;
        RECT  6.4575 27.3975 6.5225 27.5325 ;
        RECT  6.2675 28.1075 6.3325 28.3825 ;
        RECT  6.4575 28.1075 6.5225 28.3825 ;
        RECT  6.2675 28.1075 6.3325 28.3825 ;
        RECT  6.4575 28.1075 6.5225 28.3825 ;
        RECT  6.6275 28.1075 6.6925 28.3825 ;
        RECT  6.6275 27.2625 6.6925 27.3975 ;
        RECT  6.235 27.71 6.37 27.775 ;
        RECT  4.6325 27.675 4.6975 27.81 ;
        RECT  4.7725 28.035 4.8375 28.17 ;
        RECT  5.45 28.07 5.585 28.135 ;
        RECT  5.3175 28.5375 5.3825 28.9025 ;
        RECT  5.3175 29.6825 5.3825 29.8175 ;
        RECT  4.9575 29.7475 5.0225 29.8175 ;
        RECT  4.9575 28.5375 5.0225 28.6275 ;
        RECT  5.1475 28.7675 5.2125 29.715 ;
        RECT  4.89 29.235 4.925 29.3 ;
        RECT  5.2125 29.235 5.45 29.3 ;
        RECT  4.89 28.4725 5.45 28.5375 ;
        RECT  4.89 29.8175 5.45 29.8825 ;
        RECT  4.9575 29.4125 5.0225 29.5475 ;
        RECT  5.1475 29.4125 5.2125 29.5475 ;
        RECT  4.9575 29.5475 5.0225 29.6825 ;
        RECT  5.1475 29.5475 5.2125 29.6825 ;
        RECT  4.9575 29.0075 5.0225 29.2825 ;
        RECT  5.1475 29.0075 5.2125 29.2825 ;
        RECT  4.9575 29.0075 5.0225 29.2825 ;
        RECT  5.1475 29.0075 5.2125 29.2825 ;
        RECT  5.3175 28.9025 5.3825 29.1775 ;
        RECT  5.3175 29.7475 5.3825 29.8825 ;
        RECT  4.925 29.31 5.06 29.375 ;
        RECT  6.0675 28.505 6.1325 28.7875 ;
        RECT  6.0675 29.67 6.1325 29.85 ;
        RECT  5.5175 28.505 5.5825 28.7875 ;
        RECT  5.8975 28.505 5.9625 28.7875 ;
        RECT  5.5175 29.5675 5.5825 29.85 ;
        RECT  5.93 28.89 5.995 28.955 ;
        RECT  5.7075 28.89 5.7725 28.955 ;
        RECT  5.93 28.9225 5.995 29.7025 ;
        RECT  5.74 28.89 5.9625 28.955 ;
        RECT  5.7075 28.7875 5.7725 28.9225 ;
        RECT  5.45 28.875 5.485 28.94 ;
        RECT  5.9625 29.1875 6.2 29.2525 ;
        RECT  5.45 29.405 5.725 29.47 ;
        RECT  5.45 28.4725 6.2 28.5375 ;
        RECT  5.45 29.8175 6.2 29.8825 ;
        RECT  5.5175 29.2775 5.5825 29.4125 ;
        RECT  5.7075 29.2775 5.7725 29.4125 ;
        RECT  5.5175 29.4125 5.5825 29.5475 ;
        RECT  5.7075 29.4125 5.7725 29.5475 ;
        RECT  5.7075 29.2775 5.7725 29.4125 ;
        RECT  5.8975 29.2775 5.9625 29.4125 ;
        RECT  5.7075 29.4125 5.7725 29.5475 ;
        RECT  5.8975 29.4125 5.9625 29.5475 ;
        RECT  5.5175 28.9425 5.5825 29.0775 ;
        RECT  5.7075 28.9425 5.7725 29.0775 ;
        RECT  5.5175 28.9425 5.5825 29.0775 ;
        RECT  5.7075 28.9425 5.7725 29.0775 ;
        RECT  5.7075 28.9425 5.7725 29.0775 ;
        RECT  5.8975 28.9425 5.9625 29.0775 ;
        RECT  5.7075 28.9425 5.7725 29.0775 ;
        RECT  5.8975 28.9425 5.9625 29.0775 ;
        RECT  6.0675 28.7875 6.1325 28.9225 ;
        RECT  6.0675 29.7025 6.1325 29.8375 ;
        RECT  5.485 28.95 5.62 29.015 ;
        RECT  5.725 29.48 5.86 29.545 ;
        RECT  6.6275 28.5375 6.6925 28.9025 ;
        RECT  6.6275 29.6825 6.6925 29.8175 ;
        RECT  6.2675 29.7475 6.3325 29.8175 ;
        RECT  6.2675 28.5375 6.3325 28.6275 ;
        RECT  6.4575 28.7675 6.5225 29.715 ;
        RECT  6.2 29.235 6.235 29.3 ;
        RECT  6.5225 29.235 6.76 29.3 ;
        RECT  6.2 28.4725 6.76 28.5375 ;
        RECT  6.2 29.8175 6.76 29.8825 ;
        RECT  6.2675 29.4125 6.3325 29.5475 ;
        RECT  6.4575 29.4125 6.5225 29.5475 ;
        RECT  6.2675 29.5475 6.3325 29.6825 ;
        RECT  6.4575 29.5475 6.5225 29.6825 ;
        RECT  6.2675 29.0075 6.3325 29.2825 ;
        RECT  6.4575 29.0075 6.5225 29.2825 ;
        RECT  6.2675 29.0075 6.3325 29.2825 ;
        RECT  6.4575 29.0075 6.5225 29.2825 ;
        RECT  6.6275 28.9025 6.6925 29.1775 ;
        RECT  6.6275 29.7475 6.6925 29.8825 ;
        RECT  6.235 29.31 6.37 29.375 ;
        RECT  4.6325 29.2 4.6975 29.335 ;
        RECT  4.7725 28.84 4.8375 28.975 ;
        RECT  5.45 28.875 5.585 28.94 ;
        RECT  5.3175 30.7975 5.3825 31.1625 ;
        RECT  5.3175 29.8825 5.3825 30.0175 ;
        RECT  4.9575 29.8825 5.0225 29.9525 ;
        RECT  4.9575 31.0725 5.0225 31.1625 ;
        RECT  5.1475 29.985 5.2125 30.9325 ;
        RECT  4.89 30.4 4.925 30.465 ;
        RECT  5.2125 30.4 5.45 30.465 ;
        RECT  4.89 31.1625 5.45 31.2275 ;
        RECT  4.89 29.8175 5.45 29.8825 ;
        RECT  4.9575 29.9525 5.0225 30.0875 ;
        RECT  5.1475 29.9525 5.2125 30.0875 ;
        RECT  4.9575 30.0875 5.0225 30.2225 ;
        RECT  5.1475 30.0875 5.2125 30.2225 ;
        RECT  4.9575 30.7975 5.0225 31.0725 ;
        RECT  5.1475 30.7975 5.2125 31.0725 ;
        RECT  4.9575 30.7975 5.0225 31.0725 ;
        RECT  5.1475 30.7975 5.2125 31.0725 ;
        RECT  5.3175 30.7975 5.3825 31.0725 ;
        RECT  5.3175 29.9525 5.3825 30.0875 ;
        RECT  4.925 30.4 5.06 30.465 ;
        RECT  6.0675 30.9125 6.1325 31.195 ;
        RECT  6.0675 29.85 6.1325 30.03 ;
        RECT  5.5175 30.9125 5.5825 31.195 ;
        RECT  5.8975 30.9125 5.9625 31.195 ;
        RECT  5.5175 29.85 5.5825 30.1325 ;
        RECT  5.93 30.745 5.995 30.81 ;
        RECT  5.7075 30.745 5.7725 30.81 ;
        RECT  5.93 29.9975 5.995 30.7775 ;
        RECT  5.74 30.745 5.9625 30.81 ;
        RECT  5.7075 30.7775 5.7725 30.9125 ;
        RECT  5.45 30.76 5.485 30.825 ;
        RECT  5.9625 30.4475 6.2 30.5125 ;
        RECT  5.45 30.23 5.725 30.295 ;
        RECT  5.45 31.1625 6.2 31.2275 ;
        RECT  5.45 29.8175 6.2 29.8825 ;
        RECT  5.5175 29.9975 5.5825 30.1325 ;
        RECT  5.7075 29.9975 5.7725 30.1325 ;
        RECT  5.5175 30.1325 5.5825 30.2675 ;
        RECT  5.7075 30.1325 5.7725 30.2675 ;
        RECT  5.7075 29.9975 5.7725 30.1325 ;
        RECT  5.8975 29.9975 5.9625 30.1325 ;
        RECT  5.7075 30.1325 5.7725 30.2675 ;
        RECT  5.8975 30.1325 5.9625 30.2675 ;
        RECT  5.5175 30.9125 5.5825 31.0475 ;
        RECT  5.7075 30.9125 5.7725 31.0475 ;
        RECT  5.5175 30.9125 5.5825 31.0475 ;
        RECT  5.7075 30.9125 5.7725 31.0475 ;
        RECT  5.7075 30.9125 5.7725 31.0475 ;
        RECT  5.8975 30.9125 5.9625 31.0475 ;
        RECT  5.7075 30.9125 5.7725 31.0475 ;
        RECT  5.8975 30.9125 5.9625 31.0475 ;
        RECT  6.0675 30.9125 6.1325 31.0475 ;
        RECT  6.0675 29.9975 6.1325 30.1325 ;
        RECT  5.485 30.76 5.62 30.825 ;
        RECT  5.725 30.23 5.86 30.295 ;
        RECT  6.6275 30.7975 6.6925 31.1625 ;
        RECT  6.6275 29.8825 6.6925 30.0175 ;
        RECT  6.2675 29.8825 6.3325 29.9525 ;
        RECT  6.2675 31.0725 6.3325 31.1625 ;
        RECT  6.4575 29.985 6.5225 30.9325 ;
        RECT  6.2 30.4 6.235 30.465 ;
        RECT  6.5225 30.4 6.76 30.465 ;
        RECT  6.2 31.1625 6.76 31.2275 ;
        RECT  6.2 29.8175 6.76 29.8825 ;
        RECT  6.2675 29.9525 6.3325 30.0875 ;
        RECT  6.4575 29.9525 6.5225 30.0875 ;
        RECT  6.2675 30.0875 6.3325 30.2225 ;
        RECT  6.4575 30.0875 6.5225 30.2225 ;
        RECT  6.2675 30.7975 6.3325 31.0725 ;
        RECT  6.4575 30.7975 6.5225 31.0725 ;
        RECT  6.2675 30.7975 6.3325 31.0725 ;
        RECT  6.4575 30.7975 6.5225 31.0725 ;
        RECT  6.6275 30.7975 6.6925 31.0725 ;
        RECT  6.6275 29.9525 6.6925 30.0875 ;
        RECT  6.235 30.4 6.37 30.465 ;
        RECT  4.6325 30.365 4.6975 30.5 ;
        RECT  4.7725 30.725 4.8375 30.86 ;
        RECT  5.45 30.76 5.585 30.825 ;
        RECT  5.3175 31.2275 5.3825 31.5925 ;
        RECT  5.3175 32.3725 5.3825 32.5075 ;
        RECT  4.9575 32.4375 5.0225 32.5075 ;
        RECT  4.9575 31.2275 5.0225 31.3175 ;
        RECT  5.1475 31.4575 5.2125 32.405 ;
        RECT  4.89 31.925 4.925 31.99 ;
        RECT  5.2125 31.925 5.45 31.99 ;
        RECT  4.89 31.1625 5.45 31.2275 ;
        RECT  4.89 32.5075 5.45 32.5725 ;
        RECT  4.9575 32.1025 5.0225 32.2375 ;
        RECT  5.1475 32.1025 5.2125 32.2375 ;
        RECT  4.9575 32.2375 5.0225 32.3725 ;
        RECT  5.1475 32.2375 5.2125 32.3725 ;
        RECT  4.9575 31.6975 5.0225 31.9725 ;
        RECT  5.1475 31.6975 5.2125 31.9725 ;
        RECT  4.9575 31.6975 5.0225 31.9725 ;
        RECT  5.1475 31.6975 5.2125 31.9725 ;
        RECT  5.3175 31.5925 5.3825 31.8675 ;
        RECT  5.3175 32.4375 5.3825 32.5725 ;
        RECT  4.925 32.0 5.06 32.065 ;
        RECT  6.0675 31.195 6.1325 31.4775 ;
        RECT  6.0675 32.36 6.1325 32.54 ;
        RECT  5.5175 31.195 5.5825 31.4775 ;
        RECT  5.8975 31.195 5.9625 31.4775 ;
        RECT  5.5175 32.2575 5.5825 32.54 ;
        RECT  5.93 31.58 5.995 31.645 ;
        RECT  5.7075 31.58 5.7725 31.645 ;
        RECT  5.93 31.6125 5.995 32.3925 ;
        RECT  5.74 31.58 5.9625 31.645 ;
        RECT  5.7075 31.4775 5.7725 31.6125 ;
        RECT  5.45 31.565 5.485 31.63 ;
        RECT  5.9625 31.8775 6.2 31.9425 ;
        RECT  5.45 32.095 5.725 32.16 ;
        RECT  5.45 31.1625 6.2 31.2275 ;
        RECT  5.45 32.5075 6.2 32.5725 ;
        RECT  5.5175 31.9675 5.5825 32.1025 ;
        RECT  5.7075 31.9675 5.7725 32.1025 ;
        RECT  5.5175 32.1025 5.5825 32.2375 ;
        RECT  5.7075 32.1025 5.7725 32.2375 ;
        RECT  5.7075 31.9675 5.7725 32.1025 ;
        RECT  5.8975 31.9675 5.9625 32.1025 ;
        RECT  5.7075 32.1025 5.7725 32.2375 ;
        RECT  5.8975 32.1025 5.9625 32.2375 ;
        RECT  5.5175 31.6325 5.5825 31.7675 ;
        RECT  5.7075 31.6325 5.7725 31.7675 ;
        RECT  5.5175 31.6325 5.5825 31.7675 ;
        RECT  5.7075 31.6325 5.7725 31.7675 ;
        RECT  5.7075 31.6325 5.7725 31.7675 ;
        RECT  5.8975 31.6325 5.9625 31.7675 ;
        RECT  5.7075 31.6325 5.7725 31.7675 ;
        RECT  5.8975 31.6325 5.9625 31.7675 ;
        RECT  6.0675 31.4775 6.1325 31.6125 ;
        RECT  6.0675 32.3925 6.1325 32.5275 ;
        RECT  5.485 31.64 5.62 31.705 ;
        RECT  5.725 32.17 5.86 32.235 ;
        RECT  6.6275 31.2275 6.6925 31.5925 ;
        RECT  6.6275 32.3725 6.6925 32.5075 ;
        RECT  6.2675 32.4375 6.3325 32.5075 ;
        RECT  6.2675 31.2275 6.3325 31.3175 ;
        RECT  6.4575 31.4575 6.5225 32.405 ;
        RECT  6.2 31.925 6.235 31.99 ;
        RECT  6.5225 31.925 6.76 31.99 ;
        RECT  6.2 31.1625 6.76 31.2275 ;
        RECT  6.2 32.5075 6.76 32.5725 ;
        RECT  6.2675 32.1025 6.3325 32.2375 ;
        RECT  6.4575 32.1025 6.5225 32.2375 ;
        RECT  6.2675 32.2375 6.3325 32.3725 ;
        RECT  6.4575 32.2375 6.5225 32.3725 ;
        RECT  6.2675 31.6975 6.3325 31.9725 ;
        RECT  6.4575 31.6975 6.5225 31.9725 ;
        RECT  6.2675 31.6975 6.3325 31.9725 ;
        RECT  6.4575 31.6975 6.5225 31.9725 ;
        RECT  6.6275 31.5925 6.6925 31.8675 ;
        RECT  6.6275 32.4375 6.6925 32.5725 ;
        RECT  6.235 32.0 6.37 32.065 ;
        RECT  4.6325 31.89 4.6975 32.025 ;
        RECT  4.7725 31.53 4.8375 31.665 ;
        RECT  5.45 31.565 5.585 31.63 ;
        RECT  5.3175 33.4875 5.3825 33.8525 ;
        RECT  5.3175 32.5725 5.3825 32.7075 ;
        RECT  4.9575 32.5725 5.0225 32.6425 ;
        RECT  4.9575 33.7625 5.0225 33.8525 ;
        RECT  5.1475 32.675 5.2125 33.6225 ;
        RECT  4.89 33.09 4.925 33.155 ;
        RECT  5.2125 33.09 5.45 33.155 ;
        RECT  4.89 33.8525 5.45 33.9175 ;
        RECT  4.89 32.5075 5.45 32.5725 ;
        RECT  4.9575 32.6425 5.0225 32.7775 ;
        RECT  5.1475 32.6425 5.2125 32.7775 ;
        RECT  4.9575 32.7775 5.0225 32.9125 ;
        RECT  5.1475 32.7775 5.2125 32.9125 ;
        RECT  4.9575 33.4875 5.0225 33.7625 ;
        RECT  5.1475 33.4875 5.2125 33.7625 ;
        RECT  4.9575 33.4875 5.0225 33.7625 ;
        RECT  5.1475 33.4875 5.2125 33.7625 ;
        RECT  5.3175 33.4875 5.3825 33.7625 ;
        RECT  5.3175 32.6425 5.3825 32.7775 ;
        RECT  4.925 33.09 5.06 33.155 ;
        RECT  6.0675 33.6025 6.1325 33.885 ;
        RECT  6.0675 32.54 6.1325 32.72 ;
        RECT  5.5175 33.6025 5.5825 33.885 ;
        RECT  5.8975 33.6025 5.9625 33.885 ;
        RECT  5.5175 32.54 5.5825 32.8225 ;
        RECT  5.93 33.435 5.995 33.5 ;
        RECT  5.7075 33.435 5.7725 33.5 ;
        RECT  5.93 32.6875 5.995 33.4675 ;
        RECT  5.74 33.435 5.9625 33.5 ;
        RECT  5.7075 33.4675 5.7725 33.6025 ;
        RECT  5.45 33.45 5.485 33.515 ;
        RECT  5.9625 33.1375 6.2 33.2025 ;
        RECT  5.45 32.92 5.725 32.985 ;
        RECT  5.45 33.8525 6.2 33.9175 ;
        RECT  5.45 32.5075 6.2 32.5725 ;
        RECT  5.5175 32.6875 5.5825 32.8225 ;
        RECT  5.7075 32.6875 5.7725 32.8225 ;
        RECT  5.5175 32.8225 5.5825 32.9575 ;
        RECT  5.7075 32.8225 5.7725 32.9575 ;
        RECT  5.7075 32.6875 5.7725 32.8225 ;
        RECT  5.8975 32.6875 5.9625 32.8225 ;
        RECT  5.7075 32.8225 5.7725 32.9575 ;
        RECT  5.8975 32.8225 5.9625 32.9575 ;
        RECT  5.5175 33.6025 5.5825 33.7375 ;
        RECT  5.7075 33.6025 5.7725 33.7375 ;
        RECT  5.5175 33.6025 5.5825 33.7375 ;
        RECT  5.7075 33.6025 5.7725 33.7375 ;
        RECT  5.7075 33.6025 5.7725 33.7375 ;
        RECT  5.8975 33.6025 5.9625 33.7375 ;
        RECT  5.7075 33.6025 5.7725 33.7375 ;
        RECT  5.8975 33.6025 5.9625 33.7375 ;
        RECT  6.0675 33.6025 6.1325 33.7375 ;
        RECT  6.0675 32.6875 6.1325 32.8225 ;
        RECT  5.485 33.45 5.62 33.515 ;
        RECT  5.725 32.92 5.86 32.985 ;
        RECT  6.6275 33.4875 6.6925 33.8525 ;
        RECT  6.6275 32.5725 6.6925 32.7075 ;
        RECT  6.2675 32.5725 6.3325 32.6425 ;
        RECT  6.2675 33.7625 6.3325 33.8525 ;
        RECT  6.4575 32.675 6.5225 33.6225 ;
        RECT  6.2 33.09 6.235 33.155 ;
        RECT  6.5225 33.09 6.76 33.155 ;
        RECT  6.2 33.8525 6.76 33.9175 ;
        RECT  6.2 32.5075 6.76 32.5725 ;
        RECT  6.2675 32.6425 6.3325 32.7775 ;
        RECT  6.4575 32.6425 6.5225 32.7775 ;
        RECT  6.2675 32.7775 6.3325 32.9125 ;
        RECT  6.4575 32.7775 6.5225 32.9125 ;
        RECT  6.2675 33.4875 6.3325 33.7625 ;
        RECT  6.4575 33.4875 6.5225 33.7625 ;
        RECT  6.2675 33.4875 6.3325 33.7625 ;
        RECT  6.4575 33.4875 6.5225 33.7625 ;
        RECT  6.6275 33.4875 6.6925 33.7625 ;
        RECT  6.6275 32.6425 6.6925 32.7775 ;
        RECT  6.235 33.09 6.37 33.155 ;
        RECT  4.6325 33.055 4.6975 33.19 ;
        RECT  4.7725 33.415 4.8375 33.55 ;
        RECT  5.45 33.45 5.585 33.515 ;
        RECT  5.3175 33.9175 5.3825 34.2825 ;
        RECT  5.3175 35.0625 5.3825 35.1975 ;
        RECT  4.9575 35.1275 5.0225 35.1975 ;
        RECT  4.9575 33.9175 5.0225 34.0075 ;
        RECT  5.1475 34.1475 5.2125 35.095 ;
        RECT  4.89 34.615 4.925 34.68 ;
        RECT  5.2125 34.615 5.45 34.68 ;
        RECT  4.89 33.8525 5.45 33.9175 ;
        RECT  4.89 35.1975 5.45 35.2625 ;
        RECT  4.9575 34.7925 5.0225 34.9275 ;
        RECT  5.1475 34.7925 5.2125 34.9275 ;
        RECT  4.9575 34.9275 5.0225 35.0625 ;
        RECT  5.1475 34.9275 5.2125 35.0625 ;
        RECT  4.9575 34.3875 5.0225 34.6625 ;
        RECT  5.1475 34.3875 5.2125 34.6625 ;
        RECT  4.9575 34.3875 5.0225 34.6625 ;
        RECT  5.1475 34.3875 5.2125 34.6625 ;
        RECT  5.3175 34.2825 5.3825 34.5575 ;
        RECT  5.3175 35.1275 5.3825 35.2625 ;
        RECT  4.925 34.69 5.06 34.755 ;
        RECT  6.0675 33.885 6.1325 34.1675 ;
        RECT  6.0675 35.05 6.1325 35.23 ;
        RECT  5.5175 33.885 5.5825 34.1675 ;
        RECT  5.8975 33.885 5.9625 34.1675 ;
        RECT  5.5175 34.9475 5.5825 35.23 ;
        RECT  5.93 34.27 5.995 34.335 ;
        RECT  5.7075 34.27 5.7725 34.335 ;
        RECT  5.93 34.3025 5.995 35.0825 ;
        RECT  5.74 34.27 5.9625 34.335 ;
        RECT  5.7075 34.1675 5.7725 34.3025 ;
        RECT  5.45 34.255 5.485 34.32 ;
        RECT  5.9625 34.5675 6.2 34.6325 ;
        RECT  5.45 34.785 5.725 34.85 ;
        RECT  5.45 33.8525 6.2 33.9175 ;
        RECT  5.45 35.1975 6.2 35.2625 ;
        RECT  5.5175 34.6575 5.5825 34.7925 ;
        RECT  5.7075 34.6575 5.7725 34.7925 ;
        RECT  5.5175 34.7925 5.5825 34.9275 ;
        RECT  5.7075 34.7925 5.7725 34.9275 ;
        RECT  5.7075 34.6575 5.7725 34.7925 ;
        RECT  5.8975 34.6575 5.9625 34.7925 ;
        RECT  5.7075 34.7925 5.7725 34.9275 ;
        RECT  5.8975 34.7925 5.9625 34.9275 ;
        RECT  5.5175 34.3225 5.5825 34.4575 ;
        RECT  5.7075 34.3225 5.7725 34.4575 ;
        RECT  5.5175 34.3225 5.5825 34.4575 ;
        RECT  5.7075 34.3225 5.7725 34.4575 ;
        RECT  5.7075 34.3225 5.7725 34.4575 ;
        RECT  5.8975 34.3225 5.9625 34.4575 ;
        RECT  5.7075 34.3225 5.7725 34.4575 ;
        RECT  5.8975 34.3225 5.9625 34.4575 ;
        RECT  6.0675 34.1675 6.1325 34.3025 ;
        RECT  6.0675 35.0825 6.1325 35.2175 ;
        RECT  5.485 34.33 5.62 34.395 ;
        RECT  5.725 34.86 5.86 34.925 ;
        RECT  6.6275 33.9175 6.6925 34.2825 ;
        RECT  6.6275 35.0625 6.6925 35.1975 ;
        RECT  6.2675 35.1275 6.3325 35.1975 ;
        RECT  6.2675 33.9175 6.3325 34.0075 ;
        RECT  6.4575 34.1475 6.5225 35.095 ;
        RECT  6.2 34.615 6.235 34.68 ;
        RECT  6.5225 34.615 6.76 34.68 ;
        RECT  6.2 33.8525 6.76 33.9175 ;
        RECT  6.2 35.1975 6.76 35.2625 ;
        RECT  6.2675 34.7925 6.3325 34.9275 ;
        RECT  6.4575 34.7925 6.5225 34.9275 ;
        RECT  6.2675 34.9275 6.3325 35.0625 ;
        RECT  6.4575 34.9275 6.5225 35.0625 ;
        RECT  6.2675 34.3875 6.3325 34.6625 ;
        RECT  6.4575 34.3875 6.5225 34.6625 ;
        RECT  6.2675 34.3875 6.3325 34.6625 ;
        RECT  6.4575 34.3875 6.5225 34.6625 ;
        RECT  6.6275 34.2825 6.6925 34.5575 ;
        RECT  6.6275 35.1275 6.6925 35.2625 ;
        RECT  6.235 34.69 6.37 34.755 ;
        RECT  4.6325 34.58 4.6975 34.715 ;
        RECT  4.7725 34.22 4.8375 34.355 ;
        RECT  5.45 34.255 5.585 34.32 ;
        RECT  5.3175 36.1775 5.3825 36.5425 ;
        RECT  5.3175 35.2625 5.3825 35.3975 ;
        RECT  4.9575 35.2625 5.0225 35.3325 ;
        RECT  4.9575 36.4525 5.0225 36.5425 ;
        RECT  5.1475 35.365 5.2125 36.3125 ;
        RECT  4.89 35.78 4.925 35.845 ;
        RECT  5.2125 35.78 5.45 35.845 ;
        RECT  4.89 36.5425 5.45 36.6075 ;
        RECT  4.89 35.1975 5.45 35.2625 ;
        RECT  4.9575 35.3325 5.0225 35.4675 ;
        RECT  5.1475 35.3325 5.2125 35.4675 ;
        RECT  4.9575 35.4675 5.0225 35.6025 ;
        RECT  5.1475 35.4675 5.2125 35.6025 ;
        RECT  4.9575 36.1775 5.0225 36.4525 ;
        RECT  5.1475 36.1775 5.2125 36.4525 ;
        RECT  4.9575 36.1775 5.0225 36.4525 ;
        RECT  5.1475 36.1775 5.2125 36.4525 ;
        RECT  5.3175 36.1775 5.3825 36.4525 ;
        RECT  5.3175 35.3325 5.3825 35.4675 ;
        RECT  4.925 35.78 5.06 35.845 ;
        RECT  6.0675 36.2925 6.1325 36.575 ;
        RECT  6.0675 35.23 6.1325 35.41 ;
        RECT  5.5175 36.2925 5.5825 36.575 ;
        RECT  5.8975 36.2925 5.9625 36.575 ;
        RECT  5.5175 35.23 5.5825 35.5125 ;
        RECT  5.93 36.125 5.995 36.19 ;
        RECT  5.7075 36.125 5.7725 36.19 ;
        RECT  5.93 35.3775 5.995 36.1575 ;
        RECT  5.74 36.125 5.9625 36.19 ;
        RECT  5.7075 36.1575 5.7725 36.2925 ;
        RECT  5.45 36.14 5.485 36.205 ;
        RECT  5.9625 35.8275 6.2 35.8925 ;
        RECT  5.45 35.61 5.725 35.675 ;
        RECT  5.45 36.5425 6.2 36.6075 ;
        RECT  5.45 35.1975 6.2 35.2625 ;
        RECT  5.5175 35.3775 5.5825 35.5125 ;
        RECT  5.7075 35.3775 5.7725 35.5125 ;
        RECT  5.5175 35.5125 5.5825 35.6475 ;
        RECT  5.7075 35.5125 5.7725 35.6475 ;
        RECT  5.7075 35.3775 5.7725 35.5125 ;
        RECT  5.8975 35.3775 5.9625 35.5125 ;
        RECT  5.7075 35.5125 5.7725 35.6475 ;
        RECT  5.8975 35.5125 5.9625 35.6475 ;
        RECT  5.5175 36.2925 5.5825 36.4275 ;
        RECT  5.7075 36.2925 5.7725 36.4275 ;
        RECT  5.5175 36.2925 5.5825 36.4275 ;
        RECT  5.7075 36.2925 5.7725 36.4275 ;
        RECT  5.7075 36.2925 5.7725 36.4275 ;
        RECT  5.8975 36.2925 5.9625 36.4275 ;
        RECT  5.7075 36.2925 5.7725 36.4275 ;
        RECT  5.8975 36.2925 5.9625 36.4275 ;
        RECT  6.0675 36.2925 6.1325 36.4275 ;
        RECT  6.0675 35.3775 6.1325 35.5125 ;
        RECT  5.485 36.14 5.62 36.205 ;
        RECT  5.725 35.61 5.86 35.675 ;
        RECT  6.6275 36.1775 6.6925 36.5425 ;
        RECT  6.6275 35.2625 6.6925 35.3975 ;
        RECT  6.2675 35.2625 6.3325 35.3325 ;
        RECT  6.2675 36.4525 6.3325 36.5425 ;
        RECT  6.4575 35.365 6.5225 36.3125 ;
        RECT  6.2 35.78 6.235 35.845 ;
        RECT  6.5225 35.78 6.76 35.845 ;
        RECT  6.2 36.5425 6.76 36.6075 ;
        RECT  6.2 35.1975 6.76 35.2625 ;
        RECT  6.2675 35.3325 6.3325 35.4675 ;
        RECT  6.4575 35.3325 6.5225 35.4675 ;
        RECT  6.2675 35.4675 6.3325 35.6025 ;
        RECT  6.4575 35.4675 6.5225 35.6025 ;
        RECT  6.2675 36.1775 6.3325 36.4525 ;
        RECT  6.4575 36.1775 6.5225 36.4525 ;
        RECT  6.2675 36.1775 6.3325 36.4525 ;
        RECT  6.4575 36.1775 6.5225 36.4525 ;
        RECT  6.6275 36.1775 6.6925 36.4525 ;
        RECT  6.6275 35.3325 6.6925 35.4675 ;
        RECT  6.235 35.78 6.37 35.845 ;
        RECT  4.6325 35.745 4.6975 35.88 ;
        RECT  4.7725 36.105 4.8375 36.24 ;
        RECT  5.45 36.14 5.585 36.205 ;
        RECT  5.3175 36.6075 5.3825 36.9725 ;
        RECT  5.3175 37.7525 5.3825 37.8875 ;
        RECT  4.9575 37.8175 5.0225 37.8875 ;
        RECT  4.9575 36.6075 5.0225 36.6975 ;
        RECT  5.1475 36.8375 5.2125 37.785 ;
        RECT  4.89 37.305 4.925 37.37 ;
        RECT  5.2125 37.305 5.45 37.37 ;
        RECT  4.89 36.5425 5.45 36.6075 ;
        RECT  4.89 37.8875 5.45 37.9525 ;
        RECT  4.9575 37.4825 5.0225 37.6175 ;
        RECT  5.1475 37.4825 5.2125 37.6175 ;
        RECT  4.9575 37.6175 5.0225 37.7525 ;
        RECT  5.1475 37.6175 5.2125 37.7525 ;
        RECT  4.9575 37.0775 5.0225 37.3525 ;
        RECT  5.1475 37.0775 5.2125 37.3525 ;
        RECT  4.9575 37.0775 5.0225 37.3525 ;
        RECT  5.1475 37.0775 5.2125 37.3525 ;
        RECT  5.3175 36.9725 5.3825 37.2475 ;
        RECT  5.3175 37.8175 5.3825 37.9525 ;
        RECT  4.925 37.38 5.06 37.445 ;
        RECT  6.0675 36.575 6.1325 36.8575 ;
        RECT  6.0675 37.74 6.1325 37.92 ;
        RECT  5.5175 36.575 5.5825 36.8575 ;
        RECT  5.8975 36.575 5.9625 36.8575 ;
        RECT  5.5175 37.6375 5.5825 37.92 ;
        RECT  5.93 36.96 5.995 37.025 ;
        RECT  5.7075 36.96 5.7725 37.025 ;
        RECT  5.93 36.9925 5.995 37.7725 ;
        RECT  5.74 36.96 5.9625 37.025 ;
        RECT  5.7075 36.8575 5.7725 36.9925 ;
        RECT  5.45 36.945 5.485 37.01 ;
        RECT  5.9625 37.2575 6.2 37.3225 ;
        RECT  5.45 37.475 5.725 37.54 ;
        RECT  5.45 36.5425 6.2 36.6075 ;
        RECT  5.45 37.8875 6.2 37.9525 ;
        RECT  5.5175 37.3475 5.5825 37.4825 ;
        RECT  5.7075 37.3475 5.7725 37.4825 ;
        RECT  5.5175 37.4825 5.5825 37.6175 ;
        RECT  5.7075 37.4825 5.7725 37.6175 ;
        RECT  5.7075 37.3475 5.7725 37.4825 ;
        RECT  5.8975 37.3475 5.9625 37.4825 ;
        RECT  5.7075 37.4825 5.7725 37.6175 ;
        RECT  5.8975 37.4825 5.9625 37.6175 ;
        RECT  5.5175 37.0125 5.5825 37.1475 ;
        RECT  5.7075 37.0125 5.7725 37.1475 ;
        RECT  5.5175 37.0125 5.5825 37.1475 ;
        RECT  5.7075 37.0125 5.7725 37.1475 ;
        RECT  5.7075 37.0125 5.7725 37.1475 ;
        RECT  5.8975 37.0125 5.9625 37.1475 ;
        RECT  5.7075 37.0125 5.7725 37.1475 ;
        RECT  5.8975 37.0125 5.9625 37.1475 ;
        RECT  6.0675 36.8575 6.1325 36.9925 ;
        RECT  6.0675 37.7725 6.1325 37.9075 ;
        RECT  5.485 37.02 5.62 37.085 ;
        RECT  5.725 37.55 5.86 37.615 ;
        RECT  6.6275 36.6075 6.6925 36.9725 ;
        RECT  6.6275 37.7525 6.6925 37.8875 ;
        RECT  6.2675 37.8175 6.3325 37.8875 ;
        RECT  6.2675 36.6075 6.3325 36.6975 ;
        RECT  6.4575 36.8375 6.5225 37.785 ;
        RECT  6.2 37.305 6.235 37.37 ;
        RECT  6.5225 37.305 6.76 37.37 ;
        RECT  6.2 36.5425 6.76 36.6075 ;
        RECT  6.2 37.8875 6.76 37.9525 ;
        RECT  6.2675 37.4825 6.3325 37.6175 ;
        RECT  6.4575 37.4825 6.5225 37.6175 ;
        RECT  6.2675 37.6175 6.3325 37.7525 ;
        RECT  6.4575 37.6175 6.5225 37.7525 ;
        RECT  6.2675 37.0775 6.3325 37.3525 ;
        RECT  6.4575 37.0775 6.5225 37.3525 ;
        RECT  6.2675 37.0775 6.3325 37.3525 ;
        RECT  6.4575 37.0775 6.5225 37.3525 ;
        RECT  6.6275 36.9725 6.6925 37.2475 ;
        RECT  6.6275 37.8175 6.6925 37.9525 ;
        RECT  6.235 37.38 6.37 37.445 ;
        RECT  4.6325 37.27 4.6975 37.405 ;
        RECT  4.7725 36.91 4.8375 37.045 ;
        RECT  5.45 36.945 5.585 37.01 ;
        RECT  5.3175 38.8675 5.3825 39.2325 ;
        RECT  5.3175 37.9525 5.3825 38.0875 ;
        RECT  4.9575 37.9525 5.0225 38.0225 ;
        RECT  4.9575 39.1425 5.0225 39.2325 ;
        RECT  5.1475 38.055 5.2125 39.0025 ;
        RECT  4.89 38.47 4.925 38.535 ;
        RECT  5.2125 38.47 5.45 38.535 ;
        RECT  4.89 39.2325 5.45 39.2975 ;
        RECT  4.89 37.8875 5.45 37.9525 ;
        RECT  4.9575 38.0225 5.0225 38.1575 ;
        RECT  5.1475 38.0225 5.2125 38.1575 ;
        RECT  4.9575 38.1575 5.0225 38.2925 ;
        RECT  5.1475 38.1575 5.2125 38.2925 ;
        RECT  4.9575 38.8675 5.0225 39.1425 ;
        RECT  5.1475 38.8675 5.2125 39.1425 ;
        RECT  4.9575 38.8675 5.0225 39.1425 ;
        RECT  5.1475 38.8675 5.2125 39.1425 ;
        RECT  5.3175 38.8675 5.3825 39.1425 ;
        RECT  5.3175 38.0225 5.3825 38.1575 ;
        RECT  4.925 38.47 5.06 38.535 ;
        RECT  6.0675 38.9825 6.1325 39.265 ;
        RECT  6.0675 37.92 6.1325 38.1 ;
        RECT  5.5175 38.9825 5.5825 39.265 ;
        RECT  5.8975 38.9825 5.9625 39.265 ;
        RECT  5.5175 37.92 5.5825 38.2025 ;
        RECT  5.93 38.815 5.995 38.88 ;
        RECT  5.7075 38.815 5.7725 38.88 ;
        RECT  5.93 38.0675 5.995 38.8475 ;
        RECT  5.74 38.815 5.9625 38.88 ;
        RECT  5.7075 38.8475 5.7725 38.9825 ;
        RECT  5.45 38.83 5.485 38.895 ;
        RECT  5.9625 38.5175 6.2 38.5825 ;
        RECT  5.45 38.3 5.725 38.365 ;
        RECT  5.45 39.2325 6.2 39.2975 ;
        RECT  5.45 37.8875 6.2 37.9525 ;
        RECT  5.5175 38.0675 5.5825 38.2025 ;
        RECT  5.7075 38.0675 5.7725 38.2025 ;
        RECT  5.5175 38.2025 5.5825 38.3375 ;
        RECT  5.7075 38.2025 5.7725 38.3375 ;
        RECT  5.7075 38.0675 5.7725 38.2025 ;
        RECT  5.8975 38.0675 5.9625 38.2025 ;
        RECT  5.7075 38.2025 5.7725 38.3375 ;
        RECT  5.8975 38.2025 5.9625 38.3375 ;
        RECT  5.5175 38.9825 5.5825 39.1175 ;
        RECT  5.7075 38.9825 5.7725 39.1175 ;
        RECT  5.5175 38.9825 5.5825 39.1175 ;
        RECT  5.7075 38.9825 5.7725 39.1175 ;
        RECT  5.7075 38.9825 5.7725 39.1175 ;
        RECT  5.8975 38.9825 5.9625 39.1175 ;
        RECT  5.7075 38.9825 5.7725 39.1175 ;
        RECT  5.8975 38.9825 5.9625 39.1175 ;
        RECT  6.0675 38.9825 6.1325 39.1175 ;
        RECT  6.0675 38.0675 6.1325 38.2025 ;
        RECT  5.485 38.83 5.62 38.895 ;
        RECT  5.725 38.3 5.86 38.365 ;
        RECT  6.6275 38.8675 6.6925 39.2325 ;
        RECT  6.6275 37.9525 6.6925 38.0875 ;
        RECT  6.2675 37.9525 6.3325 38.0225 ;
        RECT  6.2675 39.1425 6.3325 39.2325 ;
        RECT  6.4575 38.055 6.5225 39.0025 ;
        RECT  6.2 38.47 6.235 38.535 ;
        RECT  6.5225 38.47 6.76 38.535 ;
        RECT  6.2 39.2325 6.76 39.2975 ;
        RECT  6.2 37.8875 6.76 37.9525 ;
        RECT  6.2675 38.0225 6.3325 38.1575 ;
        RECT  6.4575 38.0225 6.5225 38.1575 ;
        RECT  6.2675 38.1575 6.3325 38.2925 ;
        RECT  6.4575 38.1575 6.5225 38.2925 ;
        RECT  6.2675 38.8675 6.3325 39.1425 ;
        RECT  6.4575 38.8675 6.5225 39.1425 ;
        RECT  6.2675 38.8675 6.3325 39.1425 ;
        RECT  6.4575 38.8675 6.5225 39.1425 ;
        RECT  6.6275 38.8675 6.6925 39.1425 ;
        RECT  6.6275 38.0225 6.6925 38.1575 ;
        RECT  6.235 38.47 6.37 38.535 ;
        RECT  4.6325 38.435 4.6975 38.57 ;
        RECT  4.7725 38.795 4.8375 38.93 ;
        RECT  5.45 38.83 5.585 38.895 ;
        RECT  5.3175 39.2975 5.3825 39.6625 ;
        RECT  5.3175 40.4425 5.3825 40.5775 ;
        RECT  4.9575 40.5075 5.0225 40.5775 ;
        RECT  4.9575 39.2975 5.0225 39.3875 ;
        RECT  5.1475 39.5275 5.2125 40.475 ;
        RECT  4.89 39.995 4.925 40.06 ;
        RECT  5.2125 39.995 5.45 40.06 ;
        RECT  4.89 39.2325 5.45 39.2975 ;
        RECT  4.89 40.5775 5.45 40.6425 ;
        RECT  4.9575 40.1725 5.0225 40.3075 ;
        RECT  5.1475 40.1725 5.2125 40.3075 ;
        RECT  4.9575 40.3075 5.0225 40.4425 ;
        RECT  5.1475 40.3075 5.2125 40.4425 ;
        RECT  4.9575 39.7675 5.0225 40.0425 ;
        RECT  5.1475 39.7675 5.2125 40.0425 ;
        RECT  4.9575 39.7675 5.0225 40.0425 ;
        RECT  5.1475 39.7675 5.2125 40.0425 ;
        RECT  5.3175 39.6625 5.3825 39.9375 ;
        RECT  5.3175 40.5075 5.3825 40.6425 ;
        RECT  4.925 40.07 5.06 40.135 ;
        RECT  6.0675 39.265 6.1325 39.5475 ;
        RECT  6.0675 40.43 6.1325 40.61 ;
        RECT  5.5175 39.265 5.5825 39.5475 ;
        RECT  5.8975 39.265 5.9625 39.5475 ;
        RECT  5.5175 40.3275 5.5825 40.61 ;
        RECT  5.93 39.65 5.995 39.715 ;
        RECT  5.7075 39.65 5.7725 39.715 ;
        RECT  5.93 39.6825 5.995 40.4625 ;
        RECT  5.74 39.65 5.9625 39.715 ;
        RECT  5.7075 39.5475 5.7725 39.6825 ;
        RECT  5.45 39.635 5.485 39.7 ;
        RECT  5.9625 39.9475 6.2 40.0125 ;
        RECT  5.45 40.165 5.725 40.23 ;
        RECT  5.45 39.2325 6.2 39.2975 ;
        RECT  5.45 40.5775 6.2 40.6425 ;
        RECT  5.5175 40.0375 5.5825 40.1725 ;
        RECT  5.7075 40.0375 5.7725 40.1725 ;
        RECT  5.5175 40.1725 5.5825 40.3075 ;
        RECT  5.7075 40.1725 5.7725 40.3075 ;
        RECT  5.7075 40.0375 5.7725 40.1725 ;
        RECT  5.8975 40.0375 5.9625 40.1725 ;
        RECT  5.7075 40.1725 5.7725 40.3075 ;
        RECT  5.8975 40.1725 5.9625 40.3075 ;
        RECT  5.5175 39.7025 5.5825 39.8375 ;
        RECT  5.7075 39.7025 5.7725 39.8375 ;
        RECT  5.5175 39.7025 5.5825 39.8375 ;
        RECT  5.7075 39.7025 5.7725 39.8375 ;
        RECT  5.7075 39.7025 5.7725 39.8375 ;
        RECT  5.8975 39.7025 5.9625 39.8375 ;
        RECT  5.7075 39.7025 5.7725 39.8375 ;
        RECT  5.8975 39.7025 5.9625 39.8375 ;
        RECT  6.0675 39.5475 6.1325 39.6825 ;
        RECT  6.0675 40.4625 6.1325 40.5975 ;
        RECT  5.485 39.71 5.62 39.775 ;
        RECT  5.725 40.24 5.86 40.305 ;
        RECT  6.6275 39.2975 6.6925 39.6625 ;
        RECT  6.6275 40.4425 6.6925 40.5775 ;
        RECT  6.2675 40.5075 6.3325 40.5775 ;
        RECT  6.2675 39.2975 6.3325 39.3875 ;
        RECT  6.4575 39.5275 6.5225 40.475 ;
        RECT  6.2 39.995 6.235 40.06 ;
        RECT  6.5225 39.995 6.76 40.06 ;
        RECT  6.2 39.2325 6.76 39.2975 ;
        RECT  6.2 40.5775 6.76 40.6425 ;
        RECT  6.2675 40.1725 6.3325 40.3075 ;
        RECT  6.4575 40.1725 6.5225 40.3075 ;
        RECT  6.2675 40.3075 6.3325 40.4425 ;
        RECT  6.4575 40.3075 6.5225 40.4425 ;
        RECT  6.2675 39.7675 6.3325 40.0425 ;
        RECT  6.4575 39.7675 6.5225 40.0425 ;
        RECT  6.2675 39.7675 6.3325 40.0425 ;
        RECT  6.4575 39.7675 6.5225 40.0425 ;
        RECT  6.6275 39.6625 6.6925 39.9375 ;
        RECT  6.6275 40.5075 6.6925 40.6425 ;
        RECT  6.235 40.07 6.37 40.135 ;
        RECT  4.6325 39.96 4.6975 40.095 ;
        RECT  4.7725 39.6 4.8375 39.735 ;
        RECT  5.45 39.635 5.585 39.7 ;
        RECT  0.685 5.1 0.75 7.92 ;
        RECT  0.845 5.1 0.91 7.92 ;
        RECT  3.69 5.1 3.755 7.92 ;
        RECT  6.65 5.1 6.715 7.92 ;
        RECT  1.7 5.1 1.765 7.92 ;
        RECT  4.66 5.1 4.725 7.92 ;
        RECT  3.17 7.315 3.305 7.38 ;
        RECT  3.17 7.5 3.305 7.565 ;
        RECT  1.935 7.315 2.07 7.38 ;
        RECT  1.935 7.5 2.07 7.565 ;
        RECT  3.17 7.505 3.305 7.57 ;
        RECT  3.17 7.69 3.305 7.755 ;
        RECT  6.13 7.505 6.265 7.57 ;
        RECT  6.13 7.69 6.265 7.755 ;
        RECT  1.935 7.505 2.07 7.57 ;
        RECT  1.935 7.69 2.07 7.755 ;
        RECT  6.13 7.315 6.265 7.38 ;
        RECT  6.13 7.5 6.265 7.565 ;
        RECT  1.4 7.505 1.535 7.57 ;
        RECT  1.4 7.69 1.535 7.755 ;
        RECT  4.36 7.365 4.495 7.43 ;
        RECT  4.36 7.55 4.495 7.615 ;
        RECT  4.895 7.315 5.03 7.38 ;
        RECT  4.895 7.5 5.03 7.565 ;
        RECT  4.895 7.505 5.03 7.57 ;
        RECT  4.895 7.69 5.03 7.755 ;
        RECT  5.32 7.315 5.455 7.38 ;
        RECT  5.32 7.5 5.455 7.565 ;
        RECT  2.36 7.315 2.495 7.38 ;
        RECT  2.36 7.5 2.495 7.565 ;
        RECT  5.705 7.315 5.84 7.38 ;
        RECT  5.705 7.5 5.84 7.565 ;
        RECT  5.705 7.505 5.84 7.57 ;
        RECT  5.705 7.69 5.84 7.755 ;
        RECT  2.36 7.505 2.495 7.57 ;
        RECT  2.36 7.69 2.495 7.755 ;
        RECT  5.32 7.505 5.455 7.57 ;
        RECT  5.32 7.69 5.455 7.755 ;
        RECT  2.745 7.505 2.88 7.57 ;
        RECT  2.745 7.69 2.88 7.755 ;
        RECT  2.745 7.315 2.88 7.38 ;
        RECT  2.745 7.5 2.88 7.565 ;
        RECT  0.975 7.505 1.11 7.57 ;
        RECT  0.975 7.69 1.11 7.755 ;
        RECT  3.95 7.43 4.085 7.495 ;
        RECT  3.95 7.615 4.085 7.68 ;
        RECT  0.685 7.5575 0.75 7.6925 ;
        RECT  6.1825 7.69 6.3175 7.755 ;
        RECT  4.3675 7.8 4.5025 7.865 ;
        RECT  3.4675 7.69 3.6025 7.755 ;
        RECT  3.9425 7.2675 4.0775 7.3325 ;
        RECT  6.5475 7.69 6.6825 7.755 ;
        RECT  1.005 7.1825 1.14 7.2475 ;
        RECT  5.0875 7.325 5.2225 7.39 ;
        RECT  3.48 7.3225 3.615 7.3875 ;
        RECT  2.0825 7.3225 2.2175 7.3875 ;
        RECT  0.865 7.8875 1.0 7.9525 ;
        RECT  0.9825 7.3125 1.1175 7.3775 ;
        RECT  2.5925 7.2425 2.6575 7.3775 ;
        RECT  1.5075 7.2725 1.6425 7.3375 ;
        RECT  5.5525 7.2425 5.6175 7.3775 ;
        RECT  6.44 7.365 6.575 7.43 ;
        RECT  2.97 7.445 3.105 7.51 ;
        RECT  5.93 7.455 6.065 7.52 ;
        RECT  4.24 7.6175 4.305 7.7525 ;
        RECT  3.9425 7.1825 4.0775 7.2475 ;
        RECT  1.235 7.7275 1.3 7.8625 ;
        RECT  2.7475 7.6875 2.8825 7.7525 ;
        RECT  6.44 7.3225 6.575 7.3875 ;
        RECT  5.93 7.5 6.065 7.565 ;
        RECT  5.5175 7.1825 5.6525 7.2475 ;
        RECT  0.815 7.1825 0.95 7.2475 ;
        RECT  3.48 7.3225 3.615 7.3875 ;
        RECT  2.5575 7.1825 2.6925 7.2475 ;
        RECT  2.3575 7.6875 2.4925 7.7525 ;
        RECT  2.3575 7.5 2.4925 7.565 ;
        RECT  2.97 7.5 3.105 7.565 ;
        RECT  5.3175 7.69 5.4525 7.755 ;
        RECT  5.3175 7.5 5.4525 7.565 ;
        RECT  0.685 7.18 0.75 7.955 ;
        RECT  3.755 7.82 6.65 7.885 ;
        RECT  6.265 7.315 6.575 7.38 ;
        RECT  5.84 7.69 6.13 7.755 ;
        RECT  5.03 7.69 5.32 7.755 ;
        RECT  6.6525 7.5425 6.715 7.615 ;
        RECT  6.265 7.5 6.65 7.57 ;
        RECT  5.03 7.5 5.32 7.57 ;
        RECT  5.55 7.5 5.7075 7.57 ;
        RECT  5.84 7.315 6.13 7.38 ;
        RECT  5.03 7.315 5.32 7.38 ;
        RECT  5.55 7.185 5.62 7.57 ;
        RECT  6.65 7.18 6.715 7.955 ;
        RECT  4.66 7.18 4.725 7.955 ;
        RECT  1.765 7.82 3.69 7.885 ;
        RECT  3.305 7.315 3.615 7.38 ;
        RECT  2.88 7.69 3.17 7.755 ;
        RECT  4.045 7.615 4.495 7.68 ;
        RECT  3.305 7.5 3.69 7.57 ;
        RECT  2.59 7.5 2.7475 7.57 ;
        RECT  3.6025 7.69 3.69 7.755 ;
        RECT  2.88 7.315 3.17 7.38 ;
        RECT  3.82 7.25 3.885 7.495 ;
        RECT  3.82 7.25 3.9425 7.3325 ;
        RECT  3.9425 7.245 4.0775 7.3125 ;
        RECT  3.69 7.18 3.755 7.955 ;
        RECT  2.07 7.69 2.36 7.755 ;
        RECT  1.5325 7.505 1.7 7.57 ;
        RECT  1.04 7.2475 1.11 7.505 ;
        RECT  0.975 7.69 1.4 7.755 ;
        RECT  2.07 7.5 2.36 7.57 ;
        RECT  1.23 7.69 1.305 7.8625 ;
        RECT  2.07 7.315 2.36 7.38 ;
        RECT  0.91 7.3125 0.9825 7.3775 ;
        RECT  2.59 7.185 2.66 7.57 ;
        RECT  1.62 7.2725 1.735 7.3375 ;
        RECT  0.845 7.18 0.91 7.955 ;
        RECT  1.7 7.18 1.765 7.955 ;
        RECT  0.69 7.75 0.7475 7.815 ;
        RECT  0.93 7.1825 1.0525 7.2475 ;
        RECT  4.4925 7.365 4.66 7.43 ;
        RECT  3.885 7.4275 3.9875 7.495 ;
        RECT  0.685 7.18 0.75 7.955 ;
        RECT  3.69 7.18 3.755 7.955 ;
        RECT  6.65 7.18 6.715 7.955 ;
        RECT  1.7 7.18 1.765 7.955 ;
        RECT  4.66 7.18 4.725 7.955 ;
        RECT  0.845 7.18 0.91 7.955 ;
        RECT  3.17 7.05 3.305 7.115 ;
        RECT  3.17 6.865 3.305 6.93 ;
        RECT  1.935 7.05 2.07 7.115 ;
        RECT  1.935 6.865 2.07 6.93 ;
        RECT  3.17 6.86 3.305 6.925 ;
        RECT  3.17 6.675 3.305 6.74 ;
        RECT  6.13 6.86 6.265 6.925 ;
        RECT  6.13 6.675 6.265 6.74 ;
        RECT  1.935 6.86 2.07 6.925 ;
        RECT  1.935 6.675 2.07 6.74 ;
        RECT  6.13 7.05 6.265 7.115 ;
        RECT  6.13 6.865 6.265 6.93 ;
        RECT  1.4 6.86 1.535 6.925 ;
        RECT  1.4 6.675 1.535 6.74 ;
        RECT  4.36 7.0 4.495 7.065 ;
        RECT  4.36 6.815 4.495 6.88 ;
        RECT  4.895 7.05 5.03 7.115 ;
        RECT  4.895 6.865 5.03 6.93 ;
        RECT  4.895 6.86 5.03 6.925 ;
        RECT  4.895 6.675 5.03 6.74 ;
        RECT  5.32 7.05 5.455 7.115 ;
        RECT  5.32 6.865 5.455 6.93 ;
        RECT  2.36 7.05 2.495 7.115 ;
        RECT  2.36 6.865 2.495 6.93 ;
        RECT  5.705 7.05 5.84 7.115 ;
        RECT  5.705 6.865 5.84 6.93 ;
        RECT  5.705 6.86 5.84 6.925 ;
        RECT  5.705 6.675 5.84 6.74 ;
        RECT  2.36 6.86 2.495 6.925 ;
        RECT  2.36 6.675 2.495 6.74 ;
        RECT  5.32 6.86 5.455 6.925 ;
        RECT  5.32 6.675 5.455 6.74 ;
        RECT  2.745 6.86 2.88 6.925 ;
        RECT  2.745 6.675 2.88 6.74 ;
        RECT  2.745 7.05 2.88 7.115 ;
        RECT  2.745 6.865 2.88 6.93 ;
        RECT  0.975 6.86 1.11 6.925 ;
        RECT  0.975 6.675 1.11 6.74 ;
        RECT  3.95 6.935 4.085 7.0 ;
        RECT  3.95 6.75 4.085 6.815 ;
        RECT  0.685 6.7375 0.75 6.8725 ;
        RECT  6.1825 6.675 6.3175 6.74 ;
        RECT  4.3675 6.565 4.5025 6.63 ;
        RECT  3.4675 6.675 3.6025 6.74 ;
        RECT  3.9425 7.0975 4.0775 7.1625 ;
        RECT  6.5475 6.675 6.6825 6.74 ;
        RECT  1.005 7.1825 1.14 7.2475 ;
        RECT  5.0875 7.04 5.2225 7.105 ;
        RECT  3.48 7.0425 3.615 7.1075 ;
        RECT  2.0825 7.0425 2.2175 7.1075 ;
        RECT  0.865 6.4775 1.0 6.5425 ;
        RECT  0.9825 7.0525 1.1175 7.1175 ;
        RECT  2.5925 7.0525 2.6575 7.1875 ;
        RECT  1.5075 7.0925 1.6425 7.1575 ;
        RECT  5.5525 7.0525 5.6175 7.1875 ;
        RECT  6.44 7.0 6.575 7.065 ;
        RECT  2.97 6.92 3.105 6.985 ;
        RECT  5.93 6.91 6.065 6.975 ;
        RECT  4.24 6.6775 4.305 6.8125 ;
        RECT  3.9425 7.1825 4.0775 7.2475 ;
        RECT  1.235 6.5675 1.3 6.7025 ;
        RECT  2.7475 6.6775 2.8825 6.7425 ;
        RECT  6.44 7.0425 6.575 7.1075 ;
        RECT  5.93 6.865 6.065 6.93 ;
        RECT  5.5175 7.1825 5.6525 7.2475 ;
        RECT  0.815 7.1825 0.95 7.2475 ;
        RECT  3.48 7.0425 3.615 7.1075 ;
        RECT  2.5575 7.1825 2.6925 7.2475 ;
        RECT  2.3575 6.6775 2.4925 6.7425 ;
        RECT  2.3575 6.865 2.4925 6.93 ;
        RECT  2.97 6.865 3.105 6.93 ;
        RECT  5.3175 6.675 5.4525 6.74 ;
        RECT  5.3175 6.865 5.4525 6.93 ;
        RECT  0.685 6.475 0.75 7.25 ;
        RECT  3.755 6.545 6.65 6.61 ;
        RECT  6.265 7.05 6.575 7.115 ;
        RECT  5.84 6.675 6.13 6.74 ;
        RECT  5.03 6.675 5.32 6.74 ;
        RECT  6.6525 6.815 6.715 6.8875 ;
        RECT  6.265 6.86 6.65 6.93 ;
        RECT  5.03 6.86 5.32 6.93 ;
        RECT  5.55 6.86 5.7075 6.93 ;
        RECT  5.84 7.05 6.13 7.115 ;
        RECT  5.03 7.05 5.32 7.115 ;
        RECT  5.55 6.86 5.62 7.245 ;
        RECT  6.65 6.475 6.715 7.25 ;
        RECT  4.66 6.475 4.725 7.25 ;
        RECT  1.765 6.545 3.69 6.61 ;
        RECT  3.305 7.05 3.615 7.115 ;
        RECT  2.88 6.675 3.17 6.74 ;
        RECT  4.045 6.75 4.495 6.815 ;
        RECT  3.305 6.86 3.69 6.93 ;
        RECT  2.59 6.86 2.7475 6.93 ;
        RECT  3.6025 6.675 3.69 6.74 ;
        RECT  2.88 7.05 3.17 7.115 ;
        RECT  3.82 6.935 3.885 7.18 ;
        RECT  3.82 7.0975 3.9425 7.18 ;
        RECT  3.9425 7.1175 4.0775 7.185 ;
        RECT  3.69 6.475 3.755 7.25 ;
        RECT  2.07 6.675 2.36 6.74 ;
        RECT  1.5325 6.86 1.7 6.925 ;
        RECT  1.04 6.925 1.11 7.1825 ;
        RECT  0.975 6.675 1.4 6.74 ;
        RECT  2.07 6.86 2.36 6.93 ;
        RECT  1.23 6.5675 1.305 6.74 ;
        RECT  2.07 7.05 2.36 7.115 ;
        RECT  0.91 7.0525 0.9825 7.1175 ;
        RECT  2.59 6.86 2.66 7.245 ;
        RECT  1.62 7.0925 1.735 7.1575 ;
        RECT  0.845 6.475 0.91 7.25 ;
        RECT  1.7 6.475 1.765 7.25 ;
        RECT  0.69 6.615 0.7475 6.68 ;
        RECT  0.93 7.1825 1.0525 7.2475 ;
        RECT  4.4925 7.0 4.66 7.065 ;
        RECT  3.885 6.935 3.9875 7.0025 ;
        RECT  0.685 6.475 0.75 7.25 ;
        RECT  3.69 6.475 3.755 7.25 ;
        RECT  6.65 6.475 6.715 7.25 ;
        RECT  1.7 6.475 1.765 7.25 ;
        RECT  4.66 6.475 4.725 7.25 ;
        RECT  0.845 6.475 0.91 7.25 ;
        RECT  3.17 5.905 3.305 5.97 ;
        RECT  3.17 6.09 3.305 6.155 ;
        RECT  1.935 5.905 2.07 5.97 ;
        RECT  1.935 6.09 2.07 6.155 ;
        RECT  3.17 6.095 3.305 6.16 ;
        RECT  3.17 6.28 3.305 6.345 ;
        RECT  6.13 6.095 6.265 6.16 ;
        RECT  6.13 6.28 6.265 6.345 ;
        RECT  1.935 6.095 2.07 6.16 ;
        RECT  1.935 6.28 2.07 6.345 ;
        RECT  6.13 5.905 6.265 5.97 ;
        RECT  6.13 6.09 6.265 6.155 ;
        RECT  1.4 6.095 1.535 6.16 ;
        RECT  1.4 6.28 1.535 6.345 ;
        RECT  4.36 5.955 4.495 6.02 ;
        RECT  4.36 6.14 4.495 6.205 ;
        RECT  4.895 5.905 5.03 5.97 ;
        RECT  4.895 6.09 5.03 6.155 ;
        RECT  4.895 6.095 5.03 6.16 ;
        RECT  4.895 6.28 5.03 6.345 ;
        RECT  5.32 5.905 5.455 5.97 ;
        RECT  5.32 6.09 5.455 6.155 ;
        RECT  2.36 5.905 2.495 5.97 ;
        RECT  2.36 6.09 2.495 6.155 ;
        RECT  5.705 5.905 5.84 5.97 ;
        RECT  5.705 6.09 5.84 6.155 ;
        RECT  5.705 6.095 5.84 6.16 ;
        RECT  5.705 6.28 5.84 6.345 ;
        RECT  2.36 6.095 2.495 6.16 ;
        RECT  2.36 6.28 2.495 6.345 ;
        RECT  5.32 6.095 5.455 6.16 ;
        RECT  5.32 6.28 5.455 6.345 ;
        RECT  2.745 6.095 2.88 6.16 ;
        RECT  2.745 6.28 2.88 6.345 ;
        RECT  2.745 5.905 2.88 5.97 ;
        RECT  2.745 6.09 2.88 6.155 ;
        RECT  0.975 6.095 1.11 6.16 ;
        RECT  0.975 6.28 1.11 6.345 ;
        RECT  3.95 6.02 4.085 6.085 ;
        RECT  3.95 6.205 4.085 6.27 ;
        RECT  0.685 6.1475 0.75 6.2825 ;
        RECT  6.1825 6.28 6.3175 6.345 ;
        RECT  4.3675 6.39 4.5025 6.455 ;
        RECT  3.4675 6.28 3.6025 6.345 ;
        RECT  3.9425 5.8575 4.0775 5.9225 ;
        RECT  6.5475 6.28 6.6825 6.345 ;
        RECT  1.005 5.7725 1.14 5.8375 ;
        RECT  5.0875 5.915 5.2225 5.98 ;
        RECT  3.48 5.9125 3.615 5.9775 ;
        RECT  2.0825 5.9125 2.2175 5.9775 ;
        RECT  0.865 6.4775 1.0 6.5425 ;
        RECT  0.9825 5.9025 1.1175 5.9675 ;
        RECT  2.5925 5.8325 2.6575 5.9675 ;
        RECT  1.5075 5.8625 1.6425 5.9275 ;
        RECT  5.5525 5.8325 5.6175 5.9675 ;
        RECT  6.44 5.955 6.575 6.02 ;
        RECT  2.97 6.035 3.105 6.1 ;
        RECT  5.93 6.045 6.065 6.11 ;
        RECT  4.24 6.2075 4.305 6.3425 ;
        RECT  3.9425 5.7725 4.0775 5.8375 ;
        RECT  1.235 6.3175 1.3 6.4525 ;
        RECT  2.7475 6.2775 2.8825 6.3425 ;
        RECT  6.44 5.9125 6.575 5.9775 ;
        RECT  5.93 6.09 6.065 6.155 ;
        RECT  5.5175 5.7725 5.6525 5.8375 ;
        RECT  0.815 5.7725 0.95 5.8375 ;
        RECT  3.48 5.9125 3.615 5.9775 ;
        RECT  2.5575 5.7725 2.6925 5.8375 ;
        RECT  2.3575 6.2775 2.4925 6.3425 ;
        RECT  2.3575 6.09 2.4925 6.155 ;
        RECT  2.97 6.09 3.105 6.155 ;
        RECT  5.3175 6.28 5.4525 6.345 ;
        RECT  5.3175 6.09 5.4525 6.155 ;
        RECT  0.685 5.77 0.75 6.545 ;
        RECT  3.755 6.41 6.65 6.475 ;
        RECT  6.265 5.905 6.575 5.97 ;
        RECT  5.84 6.28 6.13 6.345 ;
        RECT  5.03 6.28 5.32 6.345 ;
        RECT  6.6525 6.1325 6.715 6.205 ;
        RECT  6.265 6.09 6.65 6.16 ;
        RECT  5.03 6.09 5.32 6.16 ;
        RECT  5.55 6.09 5.7075 6.16 ;
        RECT  5.84 5.905 6.13 5.97 ;
        RECT  5.03 5.905 5.32 5.97 ;
        RECT  5.55 5.775 5.62 6.16 ;
        RECT  6.65 5.77 6.715 6.545 ;
        RECT  4.66 5.77 4.725 6.545 ;
        RECT  1.765 6.41 3.69 6.475 ;
        RECT  3.305 5.905 3.615 5.97 ;
        RECT  2.88 6.28 3.17 6.345 ;
        RECT  4.045 6.205 4.495 6.27 ;
        RECT  3.305 6.09 3.69 6.16 ;
        RECT  2.59 6.09 2.7475 6.16 ;
        RECT  3.6025 6.28 3.69 6.345 ;
        RECT  2.88 5.905 3.17 5.97 ;
        RECT  3.82 5.84 3.885 6.085 ;
        RECT  3.82 5.84 3.9425 5.9225 ;
        RECT  3.9425 5.835 4.0775 5.9025 ;
        RECT  3.69 5.77 3.755 6.545 ;
        RECT  2.07 6.28 2.36 6.345 ;
        RECT  1.5325 6.095 1.7 6.16 ;
        RECT  1.04 5.8375 1.11 6.095 ;
        RECT  0.975 6.28 1.4 6.345 ;
        RECT  2.07 6.09 2.36 6.16 ;
        RECT  1.23 6.28 1.305 6.4525 ;
        RECT  2.07 5.905 2.36 5.97 ;
        RECT  0.91 5.9025 0.9825 5.9675 ;
        RECT  2.59 5.775 2.66 6.16 ;
        RECT  1.62 5.8625 1.735 5.9275 ;
        RECT  0.845 5.77 0.91 6.545 ;
        RECT  1.7 5.77 1.765 6.545 ;
        RECT  0.69 6.34 0.7475 6.405 ;
        RECT  0.93 5.7725 1.0525 5.8375 ;
        RECT  4.4925 5.955 4.66 6.02 ;
        RECT  3.885 6.0175 3.9875 6.085 ;
        RECT  0.685 5.77 0.75 6.545 ;
        RECT  3.69 5.77 3.755 6.545 ;
        RECT  6.65 5.77 6.715 6.545 ;
        RECT  1.7 5.77 1.765 6.545 ;
        RECT  4.66 5.77 4.725 6.545 ;
        RECT  0.845 5.77 0.91 6.545 ;
        RECT  3.17 5.64 3.305 5.705 ;
        RECT  3.17 5.455 3.305 5.52 ;
        RECT  1.935 5.64 2.07 5.705 ;
        RECT  1.935 5.455 2.07 5.52 ;
        RECT  3.17 5.45 3.305 5.515 ;
        RECT  3.17 5.265 3.305 5.33 ;
        RECT  6.13 5.45 6.265 5.515 ;
        RECT  6.13 5.265 6.265 5.33 ;
        RECT  1.935 5.45 2.07 5.515 ;
        RECT  1.935 5.265 2.07 5.33 ;
        RECT  6.13 5.64 6.265 5.705 ;
        RECT  6.13 5.455 6.265 5.52 ;
        RECT  1.4 5.45 1.535 5.515 ;
        RECT  1.4 5.265 1.535 5.33 ;
        RECT  4.36 5.59 4.495 5.655 ;
        RECT  4.36 5.405 4.495 5.47 ;
        RECT  4.895 5.64 5.03 5.705 ;
        RECT  4.895 5.455 5.03 5.52 ;
        RECT  4.895 5.45 5.03 5.515 ;
        RECT  4.895 5.265 5.03 5.33 ;
        RECT  5.32 5.64 5.455 5.705 ;
        RECT  5.32 5.455 5.455 5.52 ;
        RECT  2.36 5.64 2.495 5.705 ;
        RECT  2.36 5.455 2.495 5.52 ;
        RECT  5.705 5.64 5.84 5.705 ;
        RECT  5.705 5.455 5.84 5.52 ;
        RECT  5.705 5.45 5.84 5.515 ;
        RECT  5.705 5.265 5.84 5.33 ;
        RECT  2.36 5.45 2.495 5.515 ;
        RECT  2.36 5.265 2.495 5.33 ;
        RECT  5.32 5.45 5.455 5.515 ;
        RECT  5.32 5.265 5.455 5.33 ;
        RECT  2.745 5.45 2.88 5.515 ;
        RECT  2.745 5.265 2.88 5.33 ;
        RECT  2.745 5.64 2.88 5.705 ;
        RECT  2.745 5.455 2.88 5.52 ;
        RECT  0.975 5.45 1.11 5.515 ;
        RECT  0.975 5.265 1.11 5.33 ;
        RECT  3.95 5.525 4.085 5.59 ;
        RECT  3.95 5.34 4.085 5.405 ;
        RECT  0.685 5.3275 0.75 5.4625 ;
        RECT  6.1825 5.265 6.3175 5.33 ;
        RECT  4.3675 5.155 4.5025 5.22 ;
        RECT  3.4675 5.265 3.6025 5.33 ;
        RECT  3.9425 5.6875 4.0775 5.7525 ;
        RECT  6.5475 5.265 6.6825 5.33 ;
        RECT  1.005 5.7725 1.14 5.8375 ;
        RECT  5.0875 5.63 5.2225 5.695 ;
        RECT  3.48 5.6325 3.615 5.6975 ;
        RECT  2.0825 5.6325 2.2175 5.6975 ;
        RECT  0.865 5.0675 1.0 5.1325 ;
        RECT  0.9825 5.6425 1.1175 5.7075 ;
        RECT  2.5925 5.6425 2.6575 5.7775 ;
        RECT  1.5075 5.6825 1.6425 5.7475 ;
        RECT  5.5525 5.6425 5.6175 5.7775 ;
        RECT  6.44 5.59 6.575 5.655 ;
        RECT  2.97 5.51 3.105 5.575 ;
        RECT  5.93 5.5 6.065 5.565 ;
        RECT  4.24 5.2675 4.305 5.4025 ;
        RECT  3.9425 5.7725 4.0775 5.8375 ;
        RECT  1.235 5.1575 1.3 5.2925 ;
        RECT  2.7475 5.2675 2.8825 5.3325 ;
        RECT  6.44 5.6325 6.575 5.6975 ;
        RECT  5.93 5.455 6.065 5.52 ;
        RECT  5.5175 5.7725 5.6525 5.8375 ;
        RECT  0.815 5.7725 0.95 5.8375 ;
        RECT  3.48 5.6325 3.615 5.6975 ;
        RECT  2.5575 5.7725 2.6925 5.8375 ;
        RECT  2.3575 5.2675 2.4925 5.3325 ;
        RECT  2.3575 5.455 2.4925 5.52 ;
        RECT  2.97 5.455 3.105 5.52 ;
        RECT  5.3175 5.265 5.4525 5.33 ;
        RECT  5.3175 5.455 5.4525 5.52 ;
        RECT  0.685 5.065 0.75 5.84 ;
        RECT  3.755 5.135 6.65 5.2 ;
        RECT  6.265 5.64 6.575 5.705 ;
        RECT  5.84 5.265 6.13 5.33 ;
        RECT  5.03 5.265 5.32 5.33 ;
        RECT  6.6525 5.405 6.715 5.4775 ;
        RECT  6.265 5.45 6.65 5.52 ;
        RECT  5.03 5.45 5.32 5.52 ;
        RECT  5.55 5.45 5.7075 5.52 ;
        RECT  5.84 5.64 6.13 5.705 ;
        RECT  5.03 5.64 5.32 5.705 ;
        RECT  5.55 5.45 5.62 5.835 ;
        RECT  6.65 5.065 6.715 5.84 ;
        RECT  4.66 5.065 4.725 5.84 ;
        RECT  1.765 5.135 3.69 5.2 ;
        RECT  3.305 5.64 3.615 5.705 ;
        RECT  2.88 5.265 3.17 5.33 ;
        RECT  4.045 5.34 4.495 5.405 ;
        RECT  3.305 5.45 3.69 5.52 ;
        RECT  2.59 5.45 2.7475 5.52 ;
        RECT  3.6025 5.265 3.69 5.33 ;
        RECT  2.88 5.64 3.17 5.705 ;
        RECT  3.82 5.525 3.885 5.77 ;
        RECT  3.82 5.6875 3.9425 5.77 ;
        RECT  3.9425 5.7075 4.0775 5.775 ;
        RECT  3.69 5.065 3.755 5.84 ;
        RECT  2.07 5.265 2.36 5.33 ;
        RECT  1.5325 5.45 1.7 5.515 ;
        RECT  1.04 5.515 1.11 5.7725 ;
        RECT  0.975 5.265 1.4 5.33 ;
        RECT  2.07 5.45 2.36 5.52 ;
        RECT  1.23 5.1575 1.305 5.33 ;
        RECT  2.07 5.64 2.36 5.705 ;
        RECT  0.91 5.6425 0.9825 5.7075 ;
        RECT  2.59 5.45 2.66 5.835 ;
        RECT  1.62 5.6825 1.735 5.7475 ;
        RECT  0.845 5.065 0.91 5.84 ;
        RECT  1.7 5.065 1.765 5.84 ;
        RECT  0.69 5.205 0.7475 5.27 ;
        RECT  0.93 5.7725 1.0525 5.8375 ;
        RECT  4.4925 5.59 4.66 5.655 ;
        RECT  3.885 5.525 3.9875 5.5925 ;
        RECT  0.685 5.065 0.75 5.84 ;
        RECT  3.69 5.065 3.755 5.84 ;
        RECT  6.65 5.065 6.715 5.84 ;
        RECT  1.7 5.065 1.765 5.84 ;
        RECT  4.66 5.065 4.725 5.84 ;
        RECT  0.845 5.065 0.91 5.84 ;
        RECT  8.2525 19.0575 8.3875 19.1225 ;
        RECT  8.2525 21.7475 8.3875 21.8125 ;
        RECT  8.2525 24.4375 8.3875 24.5025 ;
        RECT  8.2525 27.1275 8.3875 27.1925 ;
        RECT  8.2525 29.8175 8.3875 29.8825 ;
        RECT  8.2525 32.5075 8.3875 32.5725 ;
        RECT  8.2525 35.1975 8.3875 35.2625 ;
        RECT  8.2525 37.8875 8.3875 37.9525 ;
        RECT  8.2525 40.5775 8.3875 40.6425 ;
        RECT  6.785 8.5025 6.92 8.5675 ;
        RECT  7.1625 8.5025 7.2975 8.5675 ;
        RECT  6.51 9.8475 6.645 9.9125 ;
        RECT  7.3675 9.8475 7.5025 9.9125 ;
        RECT  6.785 13.8825 6.92 13.9475 ;
        RECT  7.5725 13.8825 7.7075 13.9475 ;
        RECT  6.51 15.2275 6.645 15.2925 ;
        RECT  7.7775 15.2275 7.9125 15.2925 ;
        RECT  6.99 8.2975 7.125 8.3625 ;
        RECT  6.99 10.9875 7.125 11.0525 ;
        RECT  6.99 13.6775 7.125 13.7425 ;
        RECT  6.99 16.3675 7.125 16.4325 ;
        RECT  6.92 7.535 7.055 7.6 ;
        RECT  7.1625 7.535 7.2975 7.6 ;
        RECT  6.92 6.83 7.055 6.895 ;
        RECT  7.3675 6.83 7.5025 6.895 ;
        RECT  6.92 6.125 7.055 6.19 ;
        RECT  7.5725 6.125 7.7075 6.19 ;
        RECT  6.92 5.42 7.055 5.485 ;
        RECT  7.7775 5.42 7.9125 5.485 ;
        RECT  6.92 7.8875 7.055 7.9525 ;
        RECT  8.2525 7.8875 8.3875 7.9525 ;
        RECT  6.92 7.1825 7.055 7.2475 ;
        RECT  8.2525 7.1825 8.3875 7.2475 ;
        RECT  6.92 6.4775 7.055 6.5425 ;
        RECT  8.2525 6.4775 8.3875 6.5425 ;
        RECT  6.92 5.7725 7.055 5.8375 ;
        RECT  8.2525 5.7725 8.3875 5.8375 ;
        RECT  6.92 5.0675 7.055 5.1325 ;
        RECT  8.2525 5.0675 8.3875 5.1325 ;
        RECT  9.39 3.795 9.525 3.86 ;
        RECT  8.98 1.61 9.115 1.675 ;
        RECT  9.185 3.1575 9.32 3.2225 ;
        RECT  9.39 41.395 9.525 41.46 ;
        RECT  9.595 10.2975 9.73 10.3625 ;
        RECT  9.8 14.3225 9.935 14.3875 ;
        RECT  8.81 8.09 8.875 8.225 ;
        RECT  4.5975 40.7825 4.7325 40.8475 ;
        RECT  8.81 40.78 8.875 40.915 ;
        RECT  8.4675 3.0275 8.6025 3.0925 ;
        RECT  8.4675 14.4525 8.6025 14.5175 ;
        RECT  8.4675 3.955 8.6025 4.02 ;
        RECT  8.4675 11.23 8.6025 11.295 ;
        RECT  -1.895 22.44 -1.5175 22.505 ;
        RECT  -1.895 25.4 -1.5175 25.465 ;
        RECT  -1.895 20.45 -1.5175 20.515 ;
        RECT  -1.895 23.41 -1.5175 23.475 ;
        RECT  -0.755 19.5525 -0.69 19.98 ;
        RECT  -0.755 20.6825 -0.69 21.11 ;
        RECT  -0.755 26.41 -0.69 26.65 ;
        RECT  -1.895 19.435 -1.69 19.5 ;
        RECT  -2.445 26.65 -2.38 28.46 ;
        RECT  -2.305 27.06 -2.24 28.46 ;
        RECT  -1.055 28.085 -0.99 28.46 ;
        RECT  -0.92 27.88 -0.855 28.46 ;
        RECT  -0.785 27.265 -0.72 28.46 ;
        RECT  -0.8575 29.5775 -0.69 29.6425 ;
        RECT  -0.755 30.17 -0.69 31.935 ;
        RECT  -3.745 28.085 -3.68 29.02 ;
        RECT  -3.61 27.47 -3.545 29.02 ;
        RECT  -3.475 27.265 -3.41 29.02 ;
        RECT  -3.5475 30.1375 -3.38 30.2025 ;
        RECT  -2.28 31.9025 -2.215 31.9675 ;
        RECT  -2.28 31.9025 -2.2475 31.9675 ;
        RECT  -2.28 31.73 -2.215 31.935 ;
        RECT  -0.1725 19.23 -0.1075 31.73 ;
        RECT  -0.1725 26.855 -0.1075 28.46 ;
        RECT  -1.5175 19.23 -1.4525 31.73 ;
        RECT  -1.5175 27.675 -1.4525 28.46 ;
        RECT  -2.8625 28.46 -2.7975 31.73 ;
        RECT  -2.8625 26.855 -2.7975 28.46 ;
        RECT  -4.2075 28.46 -4.1425 31.73 ;
        RECT  -4.2075 27.675 -4.1425 28.46 ;
        RECT  -0.1725 31.73 -0.1075 31.935 ;
        RECT  -1.5175 31.73 -1.4525 31.935 ;
        RECT  -2.8625 31.73 -2.7975 31.935 ;
        RECT  -4.2075 31.6975 -4.1425 31.7625 ;
        RECT  -4.22 31.6975 -4.155 31.7625 ;
        RECT  -4.2075 31.525 -4.1425 31.73 ;
        RECT  -4.1875 31.6975 -4.175 31.7625 ;
        RECT  -4.22 31.73 -4.155 31.935 ;
        RECT  -0.755 19.23 -0.69 19.295 ;
        RECT  -1.5175 19.23 -1.4525 19.295 ;
        RECT  -0.1725 19.23 -0.1075 19.295 ;
        RECT  -4.01 19.435 -1.895 19.5 ;
        RECT  -4.01 19.595 -1.895 19.66 ;
        RECT  -4.01 22.44 -1.895 22.505 ;
        RECT  -4.01 25.4 -1.895 25.465 ;
        RECT  -4.01 20.45 -1.895 20.515 ;
        RECT  -4.01 23.41 -1.895 23.475 ;
        RECT  -3.47 21.92 -3.405 22.055 ;
        RECT  -3.655 21.92 -3.59 22.055 ;
        RECT  -3.47 20.685 -3.405 20.82 ;
        RECT  -3.655 20.685 -3.59 20.82 ;
        RECT  -3.66 21.92 -3.595 22.055 ;
        RECT  -3.845 21.92 -3.78 22.055 ;
        RECT  -3.66 24.88 -3.595 25.015 ;
        RECT  -3.845 24.88 -3.78 25.015 ;
        RECT  -3.66 20.685 -3.595 20.82 ;
        RECT  -3.845 20.685 -3.78 20.82 ;
        RECT  -3.47 24.88 -3.405 25.015 ;
        RECT  -3.655 24.88 -3.59 25.015 ;
        RECT  -3.66 20.15 -3.595 20.285 ;
        RECT  -3.845 20.15 -3.78 20.285 ;
        RECT  -3.52 23.11 -3.455 23.245 ;
        RECT  -3.705 23.11 -3.64 23.245 ;
        RECT  -3.47 23.645 -3.405 23.78 ;
        RECT  -3.655 23.645 -3.59 23.78 ;
        RECT  -3.66 23.645 -3.595 23.78 ;
        RECT  -3.845 23.645 -3.78 23.78 ;
        RECT  -3.47 24.07 -3.405 24.205 ;
        RECT  -3.655 24.07 -3.59 24.205 ;
        RECT  -3.47 21.11 -3.405 21.245 ;
        RECT  -3.655 21.11 -3.59 21.245 ;
        RECT  -3.47 24.455 -3.405 24.59 ;
        RECT  -3.655 24.455 -3.59 24.59 ;
        RECT  -3.66 24.455 -3.595 24.59 ;
        RECT  -3.845 24.455 -3.78 24.59 ;
        RECT  -3.66 21.11 -3.595 21.245 ;
        RECT  -3.845 21.11 -3.78 21.245 ;
        RECT  -3.66 24.07 -3.595 24.205 ;
        RECT  -3.845 24.07 -3.78 24.205 ;
        RECT  -3.66 21.495 -3.595 21.63 ;
        RECT  -3.845 21.495 -3.78 21.63 ;
        RECT  -3.47 21.495 -3.405 21.63 ;
        RECT  -3.655 21.495 -3.59 21.63 ;
        RECT  -3.66 19.725 -3.595 19.86 ;
        RECT  -3.845 19.725 -3.78 19.86 ;
        RECT  -3.585 22.7 -3.52 22.835 ;
        RECT  -3.77 22.7 -3.705 22.835 ;
        RECT  -3.7825 19.435 -3.6475 19.5 ;
        RECT  -3.845 24.9325 -3.78 25.0675 ;
        RECT  -3.955 23.1175 -3.89 23.2525 ;
        RECT  -3.845 22.2175 -3.78 22.3525 ;
        RECT  -3.4225 22.6925 -3.3575 22.8275 ;
        RECT  -3.845 25.2975 -3.78 25.4325 ;
        RECT  -3.3375 19.755 -3.2725 19.89 ;
        RECT  -3.48 23.8375 -3.415 23.9725 ;
        RECT  -3.4775 22.23 -3.4125 22.365 ;
        RECT  -3.4775 20.8325 -3.4125 20.9675 ;
        RECT  -4.0425 19.615 -3.9775 19.75 ;
        RECT  -3.4675 19.7325 -3.4025 19.8675 ;
        RECT  -3.4675 21.3425 -3.3325 21.4075 ;
        RECT  -3.4275 20.2575 -3.3625 20.3925 ;
        RECT  -3.4675 24.3025 -3.3325 24.3675 ;
        RECT  -3.52 25.19 -3.455 25.325 ;
        RECT  -3.6 21.72 -3.535 21.855 ;
        RECT  -3.61 24.68 -3.545 24.815 ;
        RECT  -3.8425 22.99 -3.7075 23.055 ;
        RECT  -3.3375 22.6925 -3.2725 22.8275 ;
        RECT  -3.9525 19.985 -3.8175 20.05 ;
        RECT  -3.8425 21.4975 -3.7775 21.6325 ;
        RECT  -3.4775 25.19 -3.4125 25.325 ;
        RECT  -3.655 24.68 -3.59 24.815 ;
        RECT  -3.3375 24.2675 -3.2725 24.4025 ;
        RECT  -3.3375 19.565 -3.2725 19.7 ;
        RECT  -3.4775 22.23 -3.4125 22.365 ;
        RECT  -3.3375 21.3075 -3.2725 21.4425 ;
        RECT  -3.8425 21.1075 -3.7775 21.2425 ;
        RECT  -3.655 21.1075 -3.59 21.2425 ;
        RECT  -3.655 21.72 -3.59 21.855 ;
        RECT  -3.845 24.0675 -3.78 24.2025 ;
        RECT  -3.655 24.0675 -3.59 24.2025 ;
        RECT  -4.045 19.435 -3.27 19.5 ;
        RECT  -3.975 22.505 -3.91 25.4 ;
        RECT  -3.47 25.015 -3.405 25.325 ;
        RECT  -3.845 24.59 -3.78 24.88 ;
        RECT  -3.845 23.78 -3.78 24.07 ;
        RECT  -3.705 25.4025 -3.6325 25.465 ;
        RECT  -3.66 25.015 -3.59 25.4 ;
        RECT  -3.66 23.78 -3.59 24.07 ;
        RECT  -3.66 24.3 -3.59 24.4575 ;
        RECT  -3.47 24.59 -3.405 24.88 ;
        RECT  -3.47 23.78 -3.405 24.07 ;
        RECT  -3.66 24.3 -3.275 24.37 ;
        RECT  -4.045 25.4 -3.27 25.465 ;
        RECT  -4.045 23.41 -3.27 23.475 ;
        RECT  -3.975 20.515 -3.91 22.44 ;
        RECT  -3.47 22.055 -3.405 22.365 ;
        RECT  -3.845 21.63 -3.78 21.92 ;
        RECT  -3.77 22.795 -3.705 23.245 ;
        RECT  -3.66 22.055 -3.59 22.44 ;
        RECT  -3.66 21.34 -3.59 21.4975 ;
        RECT  -3.845 22.3525 -3.78 22.44 ;
        RECT  -3.47 21.63 -3.405 21.92 ;
        RECT  -3.585 22.57 -3.34 22.635 ;
        RECT  -3.4225 22.57 -3.34 22.6925 ;
        RECT  -3.4025 22.6925 -3.335 22.8275 ;
        RECT  -4.045 22.44 -3.27 22.505 ;
        RECT  -3.845 20.82 -3.78 21.11 ;
        RECT  -3.66 20.2825 -3.595 20.45 ;
        RECT  -3.595 19.79 -3.3375 19.86 ;
        RECT  -3.845 19.725 -3.78 20.15 ;
        RECT  -3.66 20.82 -3.59 21.11 ;
        RECT  -3.9525 19.98 -3.78 20.055 ;
        RECT  -3.47 20.82 -3.405 21.11 ;
        RECT  -3.4675 19.66 -3.4025 19.7325 ;
        RECT  -3.66 21.34 -3.275 21.41 ;
        RECT  -3.4275 20.37 -3.3625 20.485 ;
        RECT  -4.045 19.595 -3.27 19.66 ;
        RECT  -4.045 20.45 -3.27 20.515 ;
        RECT  -3.905 19.44 -3.84 19.4975 ;
        RECT  -3.3375 19.68 -3.2725 19.8025 ;
        RECT  -3.52 23.2425 -3.455 23.41 ;
        RECT  -3.585 22.635 -3.5175 22.7375 ;
        RECT  -4.045 19.435 -3.27 19.5 ;
        RECT  -4.045 22.44 -3.27 22.505 ;
        RECT  -4.045 25.4 -3.27 25.465 ;
        RECT  -4.045 20.45 -3.27 20.515 ;
        RECT  -4.045 23.41 -3.27 23.475 ;
        RECT  -4.045 19.595 -3.27 19.66 ;
        RECT  -3.205 21.92 -3.14 22.055 ;
        RECT  -3.02 21.92 -2.955 22.055 ;
        RECT  -3.205 20.685 -3.14 20.82 ;
        RECT  -3.02 20.685 -2.955 20.82 ;
        RECT  -3.015 21.92 -2.95 22.055 ;
        RECT  -2.83 21.92 -2.765 22.055 ;
        RECT  -3.015 24.88 -2.95 25.015 ;
        RECT  -2.83 24.88 -2.765 25.015 ;
        RECT  -3.015 20.685 -2.95 20.82 ;
        RECT  -2.83 20.685 -2.765 20.82 ;
        RECT  -3.205 24.88 -3.14 25.015 ;
        RECT  -3.02 24.88 -2.955 25.015 ;
        RECT  -3.015 20.15 -2.95 20.285 ;
        RECT  -2.83 20.15 -2.765 20.285 ;
        RECT  -3.155 23.11 -3.09 23.245 ;
        RECT  -2.97 23.11 -2.905 23.245 ;
        RECT  -3.205 23.645 -3.14 23.78 ;
        RECT  -3.02 23.645 -2.955 23.78 ;
        RECT  -3.015 23.645 -2.95 23.78 ;
        RECT  -2.83 23.645 -2.765 23.78 ;
        RECT  -3.205 24.07 -3.14 24.205 ;
        RECT  -3.02 24.07 -2.955 24.205 ;
        RECT  -3.205 21.11 -3.14 21.245 ;
        RECT  -3.02 21.11 -2.955 21.245 ;
        RECT  -3.205 24.455 -3.14 24.59 ;
        RECT  -3.02 24.455 -2.955 24.59 ;
        RECT  -3.015 24.455 -2.95 24.59 ;
        RECT  -2.83 24.455 -2.765 24.59 ;
        RECT  -3.015 21.11 -2.95 21.245 ;
        RECT  -2.83 21.11 -2.765 21.245 ;
        RECT  -3.015 24.07 -2.95 24.205 ;
        RECT  -2.83 24.07 -2.765 24.205 ;
        RECT  -3.015 21.495 -2.95 21.63 ;
        RECT  -2.83 21.495 -2.765 21.63 ;
        RECT  -3.205 21.495 -3.14 21.63 ;
        RECT  -3.02 21.495 -2.955 21.63 ;
        RECT  -3.015 19.725 -2.95 19.86 ;
        RECT  -2.83 19.725 -2.765 19.86 ;
        RECT  -3.09 22.7 -3.025 22.835 ;
        RECT  -2.905 22.7 -2.84 22.835 ;
        RECT  -2.9625 19.435 -2.8275 19.5 ;
        RECT  -2.83 24.9325 -2.765 25.0675 ;
        RECT  -2.72 23.1175 -2.655 23.2525 ;
        RECT  -2.83 22.2175 -2.765 22.3525 ;
        RECT  -3.2525 22.6925 -3.1875 22.8275 ;
        RECT  -2.83 25.2975 -2.765 25.4325 ;
        RECT  -3.3375 19.755 -3.2725 19.89 ;
        RECT  -3.195 23.8375 -3.13 23.9725 ;
        RECT  -3.1975 22.23 -3.1325 22.365 ;
        RECT  -3.1975 20.8325 -3.1325 20.9675 ;
        RECT  -2.6325 19.615 -2.5675 19.75 ;
        RECT  -3.2075 19.7325 -3.1425 19.8675 ;
        RECT  -3.2775 21.3425 -3.1425 21.4075 ;
        RECT  -3.2475 20.2575 -3.1825 20.3925 ;
        RECT  -3.2775 24.3025 -3.1425 24.3675 ;
        RECT  -3.155 25.19 -3.09 25.325 ;
        RECT  -3.075 21.72 -3.01 21.855 ;
        RECT  -3.065 24.68 -3.0 24.815 ;
        RECT  -2.9025 22.99 -2.7675 23.055 ;
        RECT  -3.3375 22.6925 -3.2725 22.8275 ;
        RECT  -2.7925 19.985 -2.6575 20.05 ;
        RECT  -2.8325 21.4975 -2.7675 21.6325 ;
        RECT  -3.1975 25.19 -3.1325 25.325 ;
        RECT  -3.02 24.68 -2.955 24.815 ;
        RECT  -3.3375 24.2675 -3.2725 24.4025 ;
        RECT  -3.3375 19.565 -3.2725 19.7 ;
        RECT  -3.1975 22.23 -3.1325 22.365 ;
        RECT  -3.3375 21.3075 -3.2725 21.4425 ;
        RECT  -2.8325 21.1075 -2.7675 21.2425 ;
        RECT  -3.02 21.1075 -2.955 21.2425 ;
        RECT  -3.02 21.72 -2.955 21.855 ;
        RECT  -2.83 24.0675 -2.765 24.2025 ;
        RECT  -3.02 24.0675 -2.955 24.2025 ;
        RECT  -3.34 19.435 -2.565 19.5 ;
        RECT  -2.7 22.505 -2.635 25.4 ;
        RECT  -3.205 25.015 -3.14 25.325 ;
        RECT  -2.83 24.59 -2.765 24.88 ;
        RECT  -2.83 23.78 -2.765 24.07 ;
        RECT  -2.9775 25.4025 -2.905 25.465 ;
        RECT  -3.02 25.015 -2.95 25.4 ;
        RECT  -3.02 23.78 -2.95 24.07 ;
        RECT  -3.02 24.3 -2.95 24.4575 ;
        RECT  -3.205 24.59 -3.14 24.88 ;
        RECT  -3.205 23.78 -3.14 24.07 ;
        RECT  -3.335 24.3 -2.95 24.37 ;
        RECT  -3.34 25.4 -2.565 25.465 ;
        RECT  -3.34 23.41 -2.565 23.475 ;
        RECT  -2.7 20.515 -2.635 22.44 ;
        RECT  -3.205 22.055 -3.14 22.365 ;
        RECT  -2.83 21.63 -2.765 21.92 ;
        RECT  -2.905 22.795 -2.84 23.245 ;
        RECT  -3.02 22.055 -2.95 22.44 ;
        RECT  -3.02 21.34 -2.95 21.4975 ;
        RECT  -2.83 22.3525 -2.765 22.44 ;
        RECT  -3.205 21.63 -3.14 21.92 ;
        RECT  -3.27 22.57 -3.025 22.635 ;
        RECT  -3.27 22.57 -3.1875 22.6925 ;
        RECT  -3.275 22.6925 -3.2075 22.8275 ;
        RECT  -3.34 22.44 -2.565 22.505 ;
        RECT  -2.83 20.82 -2.765 21.11 ;
        RECT  -3.015 20.2825 -2.95 20.45 ;
        RECT  -3.2725 19.79 -3.015 19.86 ;
        RECT  -2.83 19.725 -2.765 20.15 ;
        RECT  -3.02 20.82 -2.95 21.11 ;
        RECT  -2.83 19.98 -2.6575 20.055 ;
        RECT  -3.205 20.82 -3.14 21.11 ;
        RECT  -3.2075 19.66 -3.1425 19.7325 ;
        RECT  -3.335 21.34 -2.95 21.41 ;
        RECT  -3.2475 20.37 -3.1825 20.485 ;
        RECT  -3.34 19.595 -2.565 19.66 ;
        RECT  -3.34 20.45 -2.565 20.515 ;
        RECT  -2.77 19.44 -2.705 19.4975 ;
        RECT  -3.3375 19.68 -3.2725 19.8025 ;
        RECT  -3.155 23.2425 -3.09 23.41 ;
        RECT  -3.0925 22.635 -3.025 22.7375 ;
        RECT  -3.34 19.435 -2.565 19.5 ;
        RECT  -3.34 22.44 -2.565 22.505 ;
        RECT  -3.34 25.4 -2.565 25.465 ;
        RECT  -3.34 20.45 -2.565 20.515 ;
        RECT  -3.34 23.41 -2.565 23.475 ;
        RECT  -3.34 19.595 -2.565 19.66 ;
        RECT  -2.06 21.92 -1.995 22.055 ;
        RECT  -2.245 21.92 -2.18 22.055 ;
        RECT  -2.06 20.685 -1.995 20.82 ;
        RECT  -2.245 20.685 -2.18 20.82 ;
        RECT  -2.25 21.92 -2.185 22.055 ;
        RECT  -2.435 21.92 -2.37 22.055 ;
        RECT  -2.25 24.88 -2.185 25.015 ;
        RECT  -2.435 24.88 -2.37 25.015 ;
        RECT  -2.25 20.685 -2.185 20.82 ;
        RECT  -2.435 20.685 -2.37 20.82 ;
        RECT  -2.06 24.88 -1.995 25.015 ;
        RECT  -2.245 24.88 -2.18 25.015 ;
        RECT  -2.25 20.15 -2.185 20.285 ;
        RECT  -2.435 20.15 -2.37 20.285 ;
        RECT  -2.11 23.11 -2.045 23.245 ;
        RECT  -2.295 23.11 -2.23 23.245 ;
        RECT  -2.06 23.645 -1.995 23.78 ;
        RECT  -2.245 23.645 -2.18 23.78 ;
        RECT  -2.25 23.645 -2.185 23.78 ;
        RECT  -2.435 23.645 -2.37 23.78 ;
        RECT  -2.06 24.07 -1.995 24.205 ;
        RECT  -2.245 24.07 -2.18 24.205 ;
        RECT  -2.06 21.11 -1.995 21.245 ;
        RECT  -2.245 21.11 -2.18 21.245 ;
        RECT  -2.06 24.455 -1.995 24.59 ;
        RECT  -2.245 24.455 -2.18 24.59 ;
        RECT  -2.25 24.455 -2.185 24.59 ;
        RECT  -2.435 24.455 -2.37 24.59 ;
        RECT  -2.25 21.11 -2.185 21.245 ;
        RECT  -2.435 21.11 -2.37 21.245 ;
        RECT  -2.25 24.07 -2.185 24.205 ;
        RECT  -2.435 24.07 -2.37 24.205 ;
        RECT  -2.25 21.495 -2.185 21.63 ;
        RECT  -2.435 21.495 -2.37 21.63 ;
        RECT  -2.06 21.495 -1.995 21.63 ;
        RECT  -2.245 21.495 -2.18 21.63 ;
        RECT  -2.25 19.725 -2.185 19.86 ;
        RECT  -2.435 19.725 -2.37 19.86 ;
        RECT  -2.175 22.7 -2.11 22.835 ;
        RECT  -2.36 22.7 -2.295 22.835 ;
        RECT  -2.3725 19.435 -2.2375 19.5 ;
        RECT  -2.435 24.9325 -2.37 25.0675 ;
        RECT  -2.545 23.1175 -2.48 23.2525 ;
        RECT  -2.435 22.2175 -2.37 22.3525 ;
        RECT  -2.0125 22.6925 -1.9475 22.8275 ;
        RECT  -2.435 25.2975 -2.37 25.4325 ;
        RECT  -1.9275 19.755 -1.8625 19.89 ;
        RECT  -2.07 23.8375 -2.005 23.9725 ;
        RECT  -2.0675 22.23 -2.0025 22.365 ;
        RECT  -2.0675 20.8325 -2.0025 20.9675 ;
        RECT  -2.6325 19.615 -2.5675 19.75 ;
        RECT  -2.0575 19.7325 -1.9925 19.8675 ;
        RECT  -2.0575 21.3425 -1.9225 21.4075 ;
        RECT  -2.0175 20.2575 -1.9525 20.3925 ;
        RECT  -2.0575 24.3025 -1.9225 24.3675 ;
        RECT  -2.11 25.19 -2.045 25.325 ;
        RECT  -2.19 21.72 -2.125 21.855 ;
        RECT  -2.2 24.68 -2.135 24.815 ;
        RECT  -2.4325 22.99 -2.2975 23.055 ;
        RECT  -1.9275 22.6925 -1.8625 22.8275 ;
        RECT  -2.5425 19.985 -2.4075 20.05 ;
        RECT  -2.4325 21.4975 -2.3675 21.6325 ;
        RECT  -2.0675 25.19 -2.0025 25.325 ;
        RECT  -2.245 24.68 -2.18 24.815 ;
        RECT  -1.9275 24.2675 -1.8625 24.4025 ;
        RECT  -1.9275 19.565 -1.8625 19.7 ;
        RECT  -2.0675 22.23 -2.0025 22.365 ;
        RECT  -1.9275 21.3075 -1.8625 21.4425 ;
        RECT  -2.4325 21.1075 -2.3675 21.2425 ;
        RECT  -2.245 21.1075 -2.18 21.2425 ;
        RECT  -2.245 21.72 -2.18 21.855 ;
        RECT  -2.435 24.0675 -2.37 24.2025 ;
        RECT  -2.245 24.0675 -2.18 24.2025 ;
        RECT  -2.635 19.435 -1.86 19.5 ;
        RECT  -2.565 22.505 -2.5 25.4 ;
        RECT  -2.06 25.015 -1.995 25.325 ;
        RECT  -2.435 24.59 -2.37 24.88 ;
        RECT  -2.435 23.78 -2.37 24.07 ;
        RECT  -2.295 25.4025 -2.2225 25.465 ;
        RECT  -2.25 25.015 -2.18 25.4 ;
        RECT  -2.25 23.78 -2.18 24.07 ;
        RECT  -2.25 24.3 -2.18 24.4575 ;
        RECT  -2.06 24.59 -1.995 24.88 ;
        RECT  -2.06 23.78 -1.995 24.07 ;
        RECT  -2.25 24.3 -1.865 24.37 ;
        RECT  -2.635 25.4 -1.86 25.465 ;
        RECT  -2.635 23.41 -1.86 23.475 ;
        RECT  -2.565 20.515 -2.5 22.44 ;
        RECT  -2.06 22.055 -1.995 22.365 ;
        RECT  -2.435 21.63 -2.37 21.92 ;
        RECT  -2.36 22.795 -2.295 23.245 ;
        RECT  -2.25 22.055 -2.18 22.44 ;
        RECT  -2.25 21.34 -2.18 21.4975 ;
        RECT  -2.435 22.3525 -2.37 22.44 ;
        RECT  -2.06 21.63 -1.995 21.92 ;
        RECT  -2.175 22.57 -1.93 22.635 ;
        RECT  -2.0125 22.57 -1.93 22.6925 ;
        RECT  -1.9925 22.6925 -1.925 22.8275 ;
        RECT  -2.635 22.44 -1.86 22.505 ;
        RECT  -2.435 20.82 -2.37 21.11 ;
        RECT  -2.25 20.2825 -2.185 20.45 ;
        RECT  -2.185 19.79 -1.9275 19.86 ;
        RECT  -2.435 19.725 -2.37 20.15 ;
        RECT  -2.25 20.82 -2.18 21.11 ;
        RECT  -2.5425 19.98 -2.37 20.055 ;
        RECT  -2.06 20.82 -1.995 21.11 ;
        RECT  -2.0575 19.66 -1.9925 19.7325 ;
        RECT  -2.25 21.34 -1.865 21.41 ;
        RECT  -2.0175 20.37 -1.9525 20.485 ;
        RECT  -2.635 19.595 -1.86 19.66 ;
        RECT  -2.635 20.45 -1.86 20.515 ;
        RECT  -2.495 19.44 -2.43 19.4975 ;
        RECT  -1.9275 19.68 -1.8625 19.8025 ;
        RECT  -2.11 23.2425 -2.045 23.41 ;
        RECT  -2.175 22.635 -2.1075 22.7375 ;
        RECT  -2.635 19.435 -1.86 19.5 ;
        RECT  -2.635 22.44 -1.86 22.505 ;
        RECT  -2.635 25.4 -1.86 25.465 ;
        RECT  -2.635 20.45 -1.86 20.515 ;
        RECT  -2.635 23.41 -1.86 23.475 ;
        RECT  -2.635 19.595 -1.86 19.66 ;
        RECT  -1.4525 19.8475 -1.0875 19.9125 ;
        RECT  -0.3075 19.8475 -0.1725 19.9125 ;
        RECT  -1.2225 19.4875 -0.275 19.5525 ;
        RECT  -0.755 19.23 -0.69 19.265 ;
        RECT  -0.755 19.5525 -0.69 19.98 ;
        RECT  -1.5175 19.23 -1.4525 19.98 ;
        RECT  -0.1725 19.23 -0.1075 19.98 ;
        RECT  -0.3775 19.2975 -0.2425 19.3625 ;
        RECT  -0.3775 19.4875 -0.2425 19.5525 ;
        RECT  -0.3775 19.6775 -0.2425 19.7425 ;
        RECT  -0.175 19.2975 -0.11 19.3625 ;
        RECT  -0.175 19.6775 -0.11 19.7425 ;
        RECT  -0.3775 19.2975 -0.1775 19.3625 ;
        RECT  -0.1775 19.2975 -0.1425 19.3625 ;
        RECT  -0.175 19.33 -0.11 19.71 ;
        RECT  -0.3775 19.6775 -0.1425 19.7425 ;
        RECT  -0.175 19.2975 -0.11 19.7425 ;
        RECT  -0.5125 19.2975 -0.3775 19.3625 ;
        RECT  -0.5125 19.4875 -0.3775 19.5525 ;
        RECT  -0.5125 19.6775 -0.3775 19.7425 ;
        RECT  -1.3625 19.2975 -1.0875 19.3625 ;
        RECT  -1.3625 19.4875 -1.0875 19.5525 ;
        RECT  -1.3625 19.6775 -1.0875 19.7425 ;
        RECT  -1.495 19.2975 -1.43 19.3625 ;
        RECT  -1.495 19.6775 -1.43 19.7425 ;
        RECT  -1.4275 19.2975 -1.1575 19.3625 ;
        RECT  -1.4625 19.2975 -1.4275 19.3625 ;
        RECT  -1.495 19.33 -1.43 19.71 ;
        RECT  -1.4625 19.6775 -1.1575 19.7425 ;
        RECT  -1.495 19.2975 -1.43 19.7425 ;
        RECT  -1.3625 19.2975 -1.0875 19.3625 ;
        RECT  -1.3625 19.4875 -1.0875 19.5525 ;
        RECT  -1.3625 19.6775 -1.0875 19.7425 ;
        RECT  -1.3625 19.8475 -1.0875 19.9125 ;
        RECT  -0.3775 19.8475 -0.2425 19.9125 ;
        RECT  -0.755 19.265 -0.69 19.4 ;
        RECT  -1.4525 20.9775 -1.0875 21.0425 ;
        RECT  -0.3075 20.9775 -0.1725 21.0425 ;
        RECT  -1.2225 20.2375 -0.275 20.3025 ;
        RECT  -1.2225 20.6175 -0.275 20.6825 ;
        RECT  -0.755 19.98 -0.69 20.015 ;
        RECT  -0.755 20.6825 -0.69 21.11 ;
        RECT  -1.5175 19.98 -1.4525 21.11 ;
        RECT  -0.1725 19.98 -0.1075 21.11 ;
        RECT  -0.3775 20.0475 -0.2425 20.1125 ;
        RECT  -0.3775 20.2375 -0.2425 20.3025 ;
        RECT  -0.3775 20.4275 -0.2425 20.4925 ;
        RECT  -0.3775 20.6175 -0.2425 20.6825 ;
        RECT  -0.3775 20.8075 -0.2425 20.8725 ;
        RECT  -0.175 20.0475 -0.11 20.1125 ;
        RECT  -0.175 20.4275 -0.11 20.4925 ;
        RECT  -0.175 20.4275 -0.11 20.4925 ;
        RECT  -0.175 20.8075 -0.11 20.8725 ;
        RECT  -0.3775 20.0475 -0.1775 20.1125 ;
        RECT  -0.1775 20.0475 -0.1425 20.1125 ;
        RECT  -0.175 20.08 -0.11 20.46 ;
        RECT  -0.3775 20.4275 -0.1425 20.4925 ;
        RECT  -0.3775 20.4275 -0.1775 20.4925 ;
        RECT  -0.1775 20.4275 -0.1425 20.4925 ;
        RECT  -0.175 20.46 -0.11 20.84 ;
        RECT  -0.3775 20.8075 -0.1425 20.8725 ;
        RECT  -0.5075 20.2375 -0.4425 20.3025 ;
        RECT  -0.5075 20.6175 -0.4425 20.6825 ;
        RECT  -0.4425 20.2375 -0.3775 20.3025 ;
        RECT  -0.475 20.2375 -0.4425 20.3025 ;
        RECT  -0.5075 20.27 -0.4425 20.65 ;
        RECT  -0.475 20.6175 -0.3775 20.6825 ;
        RECT  -0.175 20.0475 -0.11 20.8725 ;
        RECT  -0.5075 20.2375 -0.4425 20.6825 ;
        RECT  -0.5125 20.0475 -0.3775 20.1125 ;
        RECT  -0.5125 20.2375 -0.3775 20.3025 ;
        RECT  -0.5125 20.4275 -0.3775 20.4925 ;
        RECT  -0.5125 20.6175 -0.3775 20.6825 ;
        RECT  -0.5125 20.8075 -0.3775 20.8725 ;
        RECT  -1.3625 20.0475 -1.0875 20.1125 ;
        RECT  -1.3625 20.2375 -1.0875 20.3025 ;
        RECT  -1.3625 20.4275 -1.0875 20.4925 ;
        RECT  -1.3625 20.6175 -1.0875 20.6825 ;
        RECT  -1.3625 20.8075 -1.0875 20.8725 ;
        RECT  -1.495 20.0475 -1.43 20.1125 ;
        RECT  -1.495 20.4275 -1.43 20.4925 ;
        RECT  -1.495 20.4275 -1.43 20.4925 ;
        RECT  -1.495 20.8075 -1.43 20.8725 ;
        RECT  -1.4275 20.0475 -1.1575 20.1125 ;
        RECT  -1.4625 20.0475 -1.4275 20.1125 ;
        RECT  -1.495 20.08 -1.43 20.46 ;
        RECT  -1.4625 20.4275 -1.1575 20.4925 ;
        RECT  -1.4275 20.4275 -1.1575 20.4925 ;
        RECT  -1.4625 20.4275 -1.4275 20.4925 ;
        RECT  -1.495 20.46 -1.43 20.84 ;
        RECT  -1.4625 20.8075 -1.1575 20.8725 ;
        RECT  -1.0225 20.2375 -0.9575 20.3025 ;
        RECT  -1.0225 20.6175 -0.9575 20.6825 ;
        RECT  -1.1575 20.2375 -1.0225 20.3025 ;
        RECT  -1.0225 20.2375 -0.99 20.3025 ;
        RECT  -1.0225 20.27 -0.9575 20.65 ;
        RECT  -1.1575 20.6175 -0.99 20.6825 ;
        RECT  -1.495 20.0475 -1.43 20.8725 ;
        RECT  -1.0225 20.2375 -0.9575 20.6825 ;
        RECT  -1.3625 20.0475 -1.0875 20.1125 ;
        RECT  -1.3625 20.2375 -1.0875 20.3025 ;
        RECT  -1.3625 20.4275 -1.0875 20.4925 ;
        RECT  -1.3625 20.6175 -1.0875 20.6825 ;
        RECT  -1.3625 20.8075 -1.0875 20.8725 ;
        RECT  -1.3625 20.9775 -1.0875 21.0425 ;
        RECT  -0.3775 20.9775 -0.2425 21.0425 ;
        RECT  -0.755 20.015 -0.69 20.15 ;
        RECT  -1.4525 22.8675 -1.0875 22.9325 ;
        RECT  -0.3075 22.8675 -0.1725 22.9325 ;
        RECT  -1.2225 21.3675 -0.275 21.4325 ;
        RECT  -1.2225 21.7475 -0.275 21.8125 ;
        RECT  -1.2225 22.1275 -0.275 22.1925 ;
        RECT  -1.2225 22.5075 -0.275 22.5725 ;
        RECT  -0.755 21.11 -0.69 21.145 ;
        RECT  -0.755 22.5725 -0.69 23.0 ;
        RECT  -1.5175 21.11 -1.4525 23.0 ;
        RECT  -0.1725 21.11 -0.1075 23.0 ;
        RECT  -0.3775 21.1775 -0.2425 21.2425 ;
        RECT  -0.3775 21.3675 -0.2425 21.4325 ;
        RECT  -0.3775 21.5575 -0.2425 21.6225 ;
        RECT  -0.3775 21.7475 -0.2425 21.8125 ;
        RECT  -0.3775 21.9375 -0.2425 22.0025 ;
        RECT  -0.3775 22.1275 -0.2425 22.1925 ;
        RECT  -0.3775 22.3175 -0.2425 22.3825 ;
        RECT  -0.3775 22.5075 -0.2425 22.5725 ;
        RECT  -0.3775 22.6975 -0.2425 22.7625 ;
        RECT  -0.175 21.1775 -0.11 21.2425 ;
        RECT  -0.175 21.5575 -0.11 21.6225 ;
        RECT  -0.175 21.5575 -0.11 21.6225 ;
        RECT  -0.175 21.9375 -0.11 22.0025 ;
        RECT  -0.175 21.9375 -0.11 22.0025 ;
        RECT  -0.175 22.3175 -0.11 22.3825 ;
        RECT  -0.175 22.3175 -0.11 22.3825 ;
        RECT  -0.175 22.6975 -0.11 22.7625 ;
        RECT  -0.3775 21.1775 -0.1775 21.2425 ;
        RECT  -0.1775 21.1775 -0.1425 21.2425 ;
        RECT  -0.175 21.21 -0.11 21.59 ;
        RECT  -0.3775 21.5575 -0.1425 21.6225 ;
        RECT  -0.3775 21.5575 -0.1775 21.6225 ;
        RECT  -0.1775 21.5575 -0.1425 21.6225 ;
        RECT  -0.175 21.59 -0.11 21.97 ;
        RECT  -0.3775 21.9375 -0.1425 22.0025 ;
        RECT  -0.3775 21.9375 -0.1775 22.0025 ;
        RECT  -0.1775 21.9375 -0.1425 22.0025 ;
        RECT  -0.175 21.97 -0.11 22.35 ;
        RECT  -0.3775 22.3175 -0.1425 22.3825 ;
        RECT  -0.3775 22.3175 -0.1775 22.3825 ;
        RECT  -0.1775 22.3175 -0.1425 22.3825 ;
        RECT  -0.175 22.35 -0.11 22.73 ;
        RECT  -0.3775 22.6975 -0.1425 22.7625 ;
        RECT  -0.5075 21.3675 -0.4425 21.4325 ;
        RECT  -0.5075 21.7475 -0.4425 21.8125 ;
        RECT  -0.5075 21.7475 -0.4425 21.8125 ;
        RECT  -0.5075 22.1275 -0.4425 22.1925 ;
        RECT  -0.5075 22.1275 -0.4425 22.1925 ;
        RECT  -0.5075 22.5075 -0.4425 22.5725 ;
        RECT  -0.4425 21.3675 -0.3775 21.4325 ;
        RECT  -0.475 21.3675 -0.4425 21.4325 ;
        RECT  -0.5075 21.4 -0.4425 21.78 ;
        RECT  -0.475 21.7475 -0.3775 21.8125 ;
        RECT  -0.4425 21.7475 -0.3775 21.8125 ;
        RECT  -0.475 21.7475 -0.4425 21.8125 ;
        RECT  -0.5075 21.78 -0.4425 22.16 ;
        RECT  -0.475 22.1275 -0.3775 22.1925 ;
        RECT  -0.4425 22.1275 -0.3775 22.1925 ;
        RECT  -0.475 22.1275 -0.4425 22.1925 ;
        RECT  -0.5075 22.16 -0.4425 22.54 ;
        RECT  -0.475 22.5075 -0.3775 22.5725 ;
        RECT  -0.175 21.1775 -0.11 22.7625 ;
        RECT  -0.5075 21.3675 -0.4425 22.5725 ;
        RECT  -0.5125 21.1775 -0.3775 21.2425 ;
        RECT  -0.5125 21.3675 -0.3775 21.4325 ;
        RECT  -0.5125 21.5575 -0.3775 21.6225 ;
        RECT  -0.5125 21.7475 -0.3775 21.8125 ;
        RECT  -0.5125 21.9375 -0.3775 22.0025 ;
        RECT  -0.5125 22.1275 -0.3775 22.1925 ;
        RECT  -0.5125 22.3175 -0.3775 22.3825 ;
        RECT  -0.5125 22.5075 -0.3775 22.5725 ;
        RECT  -0.5125 22.6975 -0.3775 22.7625 ;
        RECT  -1.3625 21.1775 -1.0875 21.2425 ;
        RECT  -1.3625 21.3675 -1.0875 21.4325 ;
        RECT  -1.3625 21.5575 -1.0875 21.6225 ;
        RECT  -1.3625 21.7475 -1.0875 21.8125 ;
        RECT  -1.3625 21.9375 -1.0875 22.0025 ;
        RECT  -1.3625 22.1275 -1.0875 22.1925 ;
        RECT  -1.3625 22.3175 -1.0875 22.3825 ;
        RECT  -1.3625 22.5075 -1.0875 22.5725 ;
        RECT  -1.3625 22.6975 -1.0875 22.7625 ;
        RECT  -1.495 21.1775 -1.43 21.2425 ;
        RECT  -1.495 21.5575 -1.43 21.6225 ;
        RECT  -1.495 21.5575 -1.43 21.6225 ;
        RECT  -1.495 21.9375 -1.43 22.0025 ;
        RECT  -1.495 21.9375 -1.43 22.0025 ;
        RECT  -1.495 22.3175 -1.43 22.3825 ;
        RECT  -1.495 22.3175 -1.43 22.3825 ;
        RECT  -1.495 22.6975 -1.43 22.7625 ;
        RECT  -1.4275 21.1775 -1.1575 21.2425 ;
        RECT  -1.4625 21.1775 -1.4275 21.2425 ;
        RECT  -1.495 21.21 -1.43 21.59 ;
        RECT  -1.4625 21.5575 -1.1575 21.6225 ;
        RECT  -1.4275 21.5575 -1.1575 21.6225 ;
        RECT  -1.4625 21.5575 -1.4275 21.6225 ;
        RECT  -1.495 21.59 -1.43 21.97 ;
        RECT  -1.4625 21.9375 -1.1575 22.0025 ;
        RECT  -1.4275 21.9375 -1.1575 22.0025 ;
        RECT  -1.4625 21.9375 -1.4275 22.0025 ;
        RECT  -1.495 21.97 -1.43 22.35 ;
        RECT  -1.4625 22.3175 -1.1575 22.3825 ;
        RECT  -1.4275 22.3175 -1.1575 22.3825 ;
        RECT  -1.4625 22.3175 -1.4275 22.3825 ;
        RECT  -1.495 22.35 -1.43 22.73 ;
        RECT  -1.4625 22.6975 -1.1575 22.7625 ;
        RECT  -1.0225 21.3675 -0.9575 21.4325 ;
        RECT  -1.0225 21.7475 -0.9575 21.8125 ;
        RECT  -1.0225 21.7475 -0.9575 21.8125 ;
        RECT  -1.0225 22.1275 -0.9575 22.1925 ;
        RECT  -1.0225 22.1275 -0.9575 22.1925 ;
        RECT  -1.0225 22.5075 -0.9575 22.5725 ;
        RECT  -1.1575 21.3675 -1.0225 21.4325 ;
        RECT  -1.0225 21.3675 -0.99 21.4325 ;
        RECT  -1.0225 21.4 -0.9575 21.78 ;
        RECT  -1.1575 21.7475 -0.99 21.8125 ;
        RECT  -1.1575 21.7475 -1.0225 21.8125 ;
        RECT  -1.0225 21.7475 -0.99 21.8125 ;
        RECT  -1.0225 21.78 -0.9575 22.16 ;
        RECT  -1.1575 22.1275 -0.99 22.1925 ;
        RECT  -1.1575 22.1275 -1.0225 22.1925 ;
        RECT  -1.0225 22.1275 -0.99 22.1925 ;
        RECT  -1.0225 22.16 -0.9575 22.54 ;
        RECT  -1.1575 22.5075 -0.99 22.5725 ;
        RECT  -1.495 21.1775 -1.43 22.7625 ;
        RECT  -1.0225 21.3675 -0.9575 22.5725 ;
        RECT  -1.3625 21.1775 -1.0875 21.2425 ;
        RECT  -1.3625 21.3675 -1.0875 21.4325 ;
        RECT  -1.3625 21.5575 -1.0875 21.6225 ;
        RECT  -1.3625 21.7475 -1.0875 21.8125 ;
        RECT  -1.3625 21.9375 -1.0875 22.0025 ;
        RECT  -1.3625 22.1275 -1.0875 22.1925 ;
        RECT  -1.3625 22.3175 -1.0875 22.3825 ;
        RECT  -1.3625 22.5075 -1.0875 22.5725 ;
        RECT  -1.3625 22.6975 -1.0875 22.7625 ;
        RECT  -1.3625 22.8675 -1.0875 22.9325 ;
        RECT  -0.3775 22.8675 -0.2425 22.9325 ;
        RECT  -0.755 21.145 -0.69 21.28 ;
        RECT  -1.4525 26.2775 -1.0875 26.3425 ;
        RECT  -0.3075 26.2775 -0.1725 26.3425 ;
        RECT  -1.2225 23.2575 -0.275 23.3225 ;
        RECT  -1.2225 23.6375 -0.275 23.7025 ;
        RECT  -1.2225 24.0175 -0.275 24.0825 ;
        RECT  -1.2225 24.3975 -0.275 24.4625 ;
        RECT  -1.2225 24.7775 -0.275 24.8425 ;
        RECT  -1.2225 25.1575 -0.275 25.2225 ;
        RECT  -1.2225 25.5375 -0.275 25.6025 ;
        RECT  -1.2225 25.9175 -0.275 25.9825 ;
        RECT  -0.755 23.0 -0.69 23.035 ;
        RECT  -0.755 25.9825 -0.69 26.41 ;
        RECT  -1.5175 23.0 -1.4525 26.41 ;
        RECT  -0.1725 23.0 -0.1075 26.41 ;
        RECT  -0.3775 23.0675 -0.2425 23.1325 ;
        RECT  -0.3775 23.2575 -0.2425 23.3225 ;
        RECT  -0.3775 23.4475 -0.2425 23.5125 ;
        RECT  -0.3775 23.6375 -0.2425 23.7025 ;
        RECT  -0.3775 23.8275 -0.2425 23.8925 ;
        RECT  -0.3775 24.0175 -0.2425 24.0825 ;
        RECT  -0.3775 24.2075 -0.2425 24.2725 ;
        RECT  -0.3775 24.3975 -0.2425 24.4625 ;
        RECT  -0.3775 24.5875 -0.2425 24.6525 ;
        RECT  -0.3775 24.7775 -0.2425 24.8425 ;
        RECT  -0.3775 24.9675 -0.2425 25.0325 ;
        RECT  -0.3775 25.1575 -0.2425 25.2225 ;
        RECT  -0.3775 25.3475 -0.2425 25.4125 ;
        RECT  -0.3775 25.5375 -0.2425 25.6025 ;
        RECT  -0.3775 25.7275 -0.2425 25.7925 ;
        RECT  -0.3775 25.9175 -0.2425 25.9825 ;
        RECT  -0.3775 26.1075 -0.2425 26.1725 ;
        RECT  -0.175 23.0675 -0.11 23.1325 ;
        RECT  -0.175 23.4475 -0.11 23.5125 ;
        RECT  -0.175 23.4475 -0.11 23.5125 ;
        RECT  -0.175 23.8275 -0.11 23.8925 ;
        RECT  -0.175 23.8275 -0.11 23.8925 ;
        RECT  -0.175 24.2075 -0.11 24.2725 ;
        RECT  -0.175 24.2075 -0.11 24.2725 ;
        RECT  -0.175 24.5875 -0.11 24.6525 ;
        RECT  -0.175 24.5875 -0.11 24.6525 ;
        RECT  -0.175 24.9675 -0.11 25.0325 ;
        RECT  -0.175 24.9675 -0.11 25.0325 ;
        RECT  -0.175 25.3475 -0.11 25.4125 ;
        RECT  -0.175 25.3475 -0.11 25.4125 ;
        RECT  -0.175 25.7275 -0.11 25.7925 ;
        RECT  -0.175 25.7275 -0.11 25.7925 ;
        RECT  -0.175 26.1075 -0.11 26.1725 ;
        RECT  -0.3775 23.0675 -0.1775 23.1325 ;
        RECT  -0.1775 23.0675 -0.1425 23.1325 ;
        RECT  -0.175 23.1 -0.11 23.48 ;
        RECT  -0.3775 23.4475 -0.1425 23.5125 ;
        RECT  -0.3775 23.4475 -0.1775 23.5125 ;
        RECT  -0.1775 23.4475 -0.1425 23.5125 ;
        RECT  -0.175 23.48 -0.11 23.86 ;
        RECT  -0.3775 23.8275 -0.1425 23.8925 ;
        RECT  -0.3775 23.8275 -0.1775 23.8925 ;
        RECT  -0.1775 23.8275 -0.1425 23.8925 ;
        RECT  -0.175 23.86 -0.11 24.24 ;
        RECT  -0.3775 24.2075 -0.1425 24.2725 ;
        RECT  -0.3775 24.2075 -0.1775 24.2725 ;
        RECT  -0.1775 24.2075 -0.1425 24.2725 ;
        RECT  -0.175 24.24 -0.11 24.62 ;
        RECT  -0.3775 24.5875 -0.1425 24.6525 ;
        RECT  -0.3775 24.5875 -0.1775 24.6525 ;
        RECT  -0.1775 24.5875 -0.1425 24.6525 ;
        RECT  -0.175 24.62 -0.11 25.0 ;
        RECT  -0.3775 24.9675 -0.1425 25.0325 ;
        RECT  -0.3775 24.9675 -0.1775 25.0325 ;
        RECT  -0.1775 24.9675 -0.1425 25.0325 ;
        RECT  -0.175 25.0 -0.11 25.38 ;
        RECT  -0.3775 25.3475 -0.1425 25.4125 ;
        RECT  -0.3775 25.3475 -0.1775 25.4125 ;
        RECT  -0.1775 25.3475 -0.1425 25.4125 ;
        RECT  -0.175 25.38 -0.11 25.76 ;
        RECT  -0.3775 25.7275 -0.1425 25.7925 ;
        RECT  -0.3775 25.7275 -0.1775 25.7925 ;
        RECT  -0.1775 25.7275 -0.1425 25.7925 ;
        RECT  -0.175 25.76 -0.11 26.14 ;
        RECT  -0.3775 26.1075 -0.1425 26.1725 ;
        RECT  -0.5075 23.2575 -0.4425 23.3225 ;
        RECT  -0.5075 23.6375 -0.4425 23.7025 ;
        RECT  -0.5075 23.6375 -0.4425 23.7025 ;
        RECT  -0.5075 24.0175 -0.4425 24.0825 ;
        RECT  -0.5075 24.0175 -0.4425 24.0825 ;
        RECT  -0.5075 24.3975 -0.4425 24.4625 ;
        RECT  -0.5075 24.3975 -0.4425 24.4625 ;
        RECT  -0.5075 24.7775 -0.4425 24.8425 ;
        RECT  -0.5075 24.7775 -0.4425 24.8425 ;
        RECT  -0.5075 25.1575 -0.4425 25.2225 ;
        RECT  -0.5075 25.1575 -0.4425 25.2225 ;
        RECT  -0.5075 25.5375 -0.4425 25.6025 ;
        RECT  -0.5075 25.5375 -0.4425 25.6025 ;
        RECT  -0.5075 25.9175 -0.4425 25.9825 ;
        RECT  -0.4425 23.2575 -0.3775 23.3225 ;
        RECT  -0.475 23.2575 -0.4425 23.3225 ;
        RECT  -0.5075 23.29 -0.4425 23.67 ;
        RECT  -0.475 23.6375 -0.3775 23.7025 ;
        RECT  -0.4425 23.6375 -0.3775 23.7025 ;
        RECT  -0.475 23.6375 -0.4425 23.7025 ;
        RECT  -0.5075 23.67 -0.4425 24.05 ;
        RECT  -0.475 24.0175 -0.3775 24.0825 ;
        RECT  -0.4425 24.0175 -0.3775 24.0825 ;
        RECT  -0.475 24.0175 -0.4425 24.0825 ;
        RECT  -0.5075 24.05 -0.4425 24.43 ;
        RECT  -0.475 24.3975 -0.3775 24.4625 ;
        RECT  -0.4425 24.3975 -0.3775 24.4625 ;
        RECT  -0.475 24.3975 -0.4425 24.4625 ;
        RECT  -0.5075 24.43 -0.4425 24.81 ;
        RECT  -0.475 24.7775 -0.3775 24.8425 ;
        RECT  -0.4425 24.7775 -0.3775 24.8425 ;
        RECT  -0.475 24.7775 -0.4425 24.8425 ;
        RECT  -0.5075 24.81 -0.4425 25.19 ;
        RECT  -0.475 25.1575 -0.3775 25.2225 ;
        RECT  -0.4425 25.1575 -0.3775 25.2225 ;
        RECT  -0.475 25.1575 -0.4425 25.2225 ;
        RECT  -0.5075 25.19 -0.4425 25.57 ;
        RECT  -0.475 25.5375 -0.3775 25.6025 ;
        RECT  -0.4425 25.5375 -0.3775 25.6025 ;
        RECT  -0.475 25.5375 -0.4425 25.6025 ;
        RECT  -0.5075 25.57 -0.4425 25.95 ;
        RECT  -0.475 25.9175 -0.3775 25.9825 ;
        RECT  -0.175 23.0675 -0.11 26.1725 ;
        RECT  -0.5075 23.2575 -0.4425 25.9825 ;
        RECT  -0.5125 23.0675 -0.3775 23.1325 ;
        RECT  -0.5125 23.2575 -0.3775 23.3225 ;
        RECT  -0.5125 23.4475 -0.3775 23.5125 ;
        RECT  -0.5125 23.6375 -0.3775 23.7025 ;
        RECT  -0.5125 23.8275 -0.3775 23.8925 ;
        RECT  -0.5125 24.0175 -0.3775 24.0825 ;
        RECT  -0.5125 24.2075 -0.3775 24.2725 ;
        RECT  -0.5125 24.3975 -0.3775 24.4625 ;
        RECT  -0.5125 24.5875 -0.3775 24.6525 ;
        RECT  -0.5125 24.7775 -0.3775 24.8425 ;
        RECT  -0.5125 24.9675 -0.3775 25.0325 ;
        RECT  -0.5125 25.1575 -0.3775 25.2225 ;
        RECT  -0.5125 25.3475 -0.3775 25.4125 ;
        RECT  -0.5125 25.5375 -0.3775 25.6025 ;
        RECT  -0.5125 25.7275 -0.3775 25.7925 ;
        RECT  -0.5125 25.9175 -0.3775 25.9825 ;
        RECT  -0.5125 26.1075 -0.3775 26.1725 ;
        RECT  -1.3625 23.0675 -1.0875 23.1325 ;
        RECT  -1.3625 23.2575 -1.0875 23.3225 ;
        RECT  -1.3625 23.4475 -1.0875 23.5125 ;
        RECT  -1.3625 23.6375 -1.0875 23.7025 ;
        RECT  -1.3625 23.8275 -1.0875 23.8925 ;
        RECT  -1.3625 24.0175 -1.0875 24.0825 ;
        RECT  -1.3625 24.2075 -1.0875 24.2725 ;
        RECT  -1.3625 24.3975 -1.0875 24.4625 ;
        RECT  -1.3625 24.5875 -1.0875 24.6525 ;
        RECT  -1.3625 24.7775 -1.0875 24.8425 ;
        RECT  -1.3625 24.9675 -1.0875 25.0325 ;
        RECT  -1.3625 25.1575 -1.0875 25.2225 ;
        RECT  -1.3625 25.3475 -1.0875 25.4125 ;
        RECT  -1.3625 25.5375 -1.0875 25.6025 ;
        RECT  -1.3625 25.7275 -1.0875 25.7925 ;
        RECT  -1.3625 25.9175 -1.0875 25.9825 ;
        RECT  -1.3625 26.1075 -1.0875 26.1725 ;
        RECT  -1.495 23.0675 -1.43 23.1325 ;
        RECT  -1.495 23.4475 -1.43 23.5125 ;
        RECT  -1.495 23.4475 -1.43 23.5125 ;
        RECT  -1.495 23.8275 -1.43 23.8925 ;
        RECT  -1.495 23.8275 -1.43 23.8925 ;
        RECT  -1.495 24.2075 -1.43 24.2725 ;
        RECT  -1.495 24.2075 -1.43 24.2725 ;
        RECT  -1.495 24.5875 -1.43 24.6525 ;
        RECT  -1.495 24.5875 -1.43 24.6525 ;
        RECT  -1.495 24.9675 -1.43 25.0325 ;
        RECT  -1.495 24.9675 -1.43 25.0325 ;
        RECT  -1.495 25.3475 -1.43 25.4125 ;
        RECT  -1.495 25.3475 -1.43 25.4125 ;
        RECT  -1.495 25.7275 -1.43 25.7925 ;
        RECT  -1.495 25.7275 -1.43 25.7925 ;
        RECT  -1.495 26.1075 -1.43 26.1725 ;
        RECT  -1.4275 23.0675 -1.1575 23.1325 ;
        RECT  -1.4625 23.0675 -1.4275 23.1325 ;
        RECT  -1.495 23.1 -1.43 23.48 ;
        RECT  -1.4625 23.4475 -1.1575 23.5125 ;
        RECT  -1.4275 23.4475 -1.1575 23.5125 ;
        RECT  -1.4625 23.4475 -1.4275 23.5125 ;
        RECT  -1.495 23.48 -1.43 23.86 ;
        RECT  -1.4625 23.8275 -1.1575 23.8925 ;
        RECT  -1.4275 23.8275 -1.1575 23.8925 ;
        RECT  -1.4625 23.8275 -1.4275 23.8925 ;
        RECT  -1.495 23.86 -1.43 24.24 ;
        RECT  -1.4625 24.2075 -1.1575 24.2725 ;
        RECT  -1.4275 24.2075 -1.1575 24.2725 ;
        RECT  -1.4625 24.2075 -1.4275 24.2725 ;
        RECT  -1.495 24.24 -1.43 24.62 ;
        RECT  -1.4625 24.5875 -1.1575 24.6525 ;
        RECT  -1.4275 24.5875 -1.1575 24.6525 ;
        RECT  -1.4625 24.5875 -1.4275 24.6525 ;
        RECT  -1.495 24.62 -1.43 25.0 ;
        RECT  -1.4625 24.9675 -1.1575 25.0325 ;
        RECT  -1.4275 24.9675 -1.1575 25.0325 ;
        RECT  -1.4625 24.9675 -1.4275 25.0325 ;
        RECT  -1.495 25.0 -1.43 25.38 ;
        RECT  -1.4625 25.3475 -1.1575 25.4125 ;
        RECT  -1.4275 25.3475 -1.1575 25.4125 ;
        RECT  -1.4625 25.3475 -1.4275 25.4125 ;
        RECT  -1.495 25.38 -1.43 25.76 ;
        RECT  -1.4625 25.7275 -1.1575 25.7925 ;
        RECT  -1.4275 25.7275 -1.1575 25.7925 ;
        RECT  -1.4625 25.7275 -1.4275 25.7925 ;
        RECT  -1.495 25.76 -1.43 26.14 ;
        RECT  -1.4625 26.1075 -1.1575 26.1725 ;
        RECT  -1.0225 23.2575 -0.9575 23.3225 ;
        RECT  -1.0225 23.6375 -0.9575 23.7025 ;
        RECT  -1.0225 23.6375 -0.9575 23.7025 ;
        RECT  -1.0225 24.0175 -0.9575 24.0825 ;
        RECT  -1.0225 24.0175 -0.9575 24.0825 ;
        RECT  -1.0225 24.3975 -0.9575 24.4625 ;
        RECT  -1.0225 24.3975 -0.9575 24.4625 ;
        RECT  -1.0225 24.7775 -0.9575 24.8425 ;
        RECT  -1.0225 24.7775 -0.9575 24.8425 ;
        RECT  -1.0225 25.1575 -0.9575 25.2225 ;
        RECT  -1.0225 25.1575 -0.9575 25.2225 ;
        RECT  -1.0225 25.5375 -0.9575 25.6025 ;
        RECT  -1.0225 25.5375 -0.9575 25.6025 ;
        RECT  -1.0225 25.9175 -0.9575 25.9825 ;
        RECT  -1.1575 23.2575 -1.0225 23.3225 ;
        RECT  -1.0225 23.2575 -0.99 23.3225 ;
        RECT  -1.0225 23.29 -0.9575 23.67 ;
        RECT  -1.1575 23.6375 -0.99 23.7025 ;
        RECT  -1.1575 23.6375 -1.0225 23.7025 ;
        RECT  -1.0225 23.6375 -0.99 23.7025 ;
        RECT  -1.0225 23.67 -0.9575 24.05 ;
        RECT  -1.1575 24.0175 -0.99 24.0825 ;
        RECT  -1.1575 24.0175 -1.0225 24.0825 ;
        RECT  -1.0225 24.0175 -0.99 24.0825 ;
        RECT  -1.0225 24.05 -0.9575 24.43 ;
        RECT  -1.1575 24.3975 -0.99 24.4625 ;
        RECT  -1.1575 24.3975 -1.0225 24.4625 ;
        RECT  -1.0225 24.3975 -0.99 24.4625 ;
        RECT  -1.0225 24.43 -0.9575 24.81 ;
        RECT  -1.1575 24.7775 -0.99 24.8425 ;
        RECT  -1.1575 24.7775 -1.0225 24.8425 ;
        RECT  -1.0225 24.7775 -0.99 24.8425 ;
        RECT  -1.0225 24.81 -0.9575 25.19 ;
        RECT  -1.1575 25.1575 -0.99 25.2225 ;
        RECT  -1.1575 25.1575 -1.0225 25.2225 ;
        RECT  -1.0225 25.1575 -0.99 25.2225 ;
        RECT  -1.0225 25.19 -0.9575 25.57 ;
        RECT  -1.1575 25.5375 -0.99 25.6025 ;
        RECT  -1.1575 25.5375 -1.0225 25.6025 ;
        RECT  -1.0225 25.5375 -0.99 25.6025 ;
        RECT  -1.0225 25.57 -0.9575 25.95 ;
        RECT  -1.1575 25.9175 -0.99 25.9825 ;
        RECT  -1.495 23.0675 -1.43 26.1725 ;
        RECT  -1.0225 23.2575 -0.9575 25.9825 ;
        RECT  -1.3625 23.0675 -1.0875 23.1325 ;
        RECT  -1.3625 23.2575 -1.0875 23.3225 ;
        RECT  -1.3625 23.4475 -1.0875 23.5125 ;
        RECT  -1.3625 23.6375 -1.0875 23.7025 ;
        RECT  -1.3625 23.8275 -1.0875 23.8925 ;
        RECT  -1.3625 24.0175 -1.0875 24.0825 ;
        RECT  -1.3625 24.2075 -1.0875 24.2725 ;
        RECT  -1.3625 24.3975 -1.0875 24.4625 ;
        RECT  -1.3625 24.5875 -1.0875 24.6525 ;
        RECT  -1.3625 24.7775 -1.0875 24.8425 ;
        RECT  -1.3625 24.9675 -1.0875 25.0325 ;
        RECT  -1.3625 25.1575 -1.0875 25.2225 ;
        RECT  -1.3625 25.3475 -1.0875 25.4125 ;
        RECT  -1.3625 25.5375 -1.0875 25.6025 ;
        RECT  -1.3625 25.7275 -1.0875 25.7925 ;
        RECT  -1.3625 25.9175 -1.0875 25.9825 ;
        RECT  -1.3625 26.1075 -1.0875 26.1725 ;
        RECT  -1.3625 26.2775 -1.0875 26.3425 ;
        RECT  -0.3775 26.2775 -0.2425 26.3425 ;
        RECT  -0.755 23.035 -0.69 23.17 ;
        RECT  -1.355 29.295 -0.27 29.36 ;
        RECT  -1.485 29.4325 -1.2025 29.4975 ;
        RECT  -0.41 29.4325 -0.14 29.4975 ;
        RECT  -1.485 28.6925 -1.2025 28.7575 ;
        RECT  -1.485 29.0725 -1.2025 29.1375 ;
        RECT  -0.4225 28.6925 -0.14 28.7575 ;
        RECT  -1.055 28.46 -0.99 28.795 ;
        RECT  -0.785 28.46 -0.72 29.175 ;
        RECT  -0.92 28.46 -0.855 28.985 ;
        RECT  -1.5175 28.46 -1.4525 29.61 ;
        RECT  -0.1725 28.46 -0.1075 29.61 ;
        RECT  -0.8575 29.295 -0.7925 29.61 ;
        RECT  -0.4675 28.6925 -0.3325 28.7575 ;
        RECT  -0.4675 28.8825 -0.3325 28.9475 ;
        RECT  -0.6025 28.6925 -0.4675 28.7575 ;
        RECT  -0.6025 28.8825 -0.4675 28.9475 ;
        RECT  -0.4675 28.8825 -0.3325 28.9475 ;
        RECT  -0.4675 29.0725 -0.3325 29.1375 ;
        RECT  -0.6025 28.8825 -0.4675 28.9475 ;
        RECT  -0.6025 29.0725 -0.4675 29.1375 ;
        RECT  -0.4675 29.0725 -0.3325 29.1375 ;
        RECT  -0.4675 29.2625 -0.3325 29.3275 ;
        RECT  -0.6025 29.0725 -0.4675 29.1375 ;
        RECT  -0.6025 29.2625 -0.4675 29.3275 ;
        RECT  -1.3375 28.6925 -1.2025 28.7575 ;
        RECT  -1.3375 28.8825 -1.2025 28.9475 ;
        RECT  -1.3375 28.6925 -1.2025 28.7575 ;
        RECT  -1.3375 28.8825 -1.2025 28.9475 ;
        RECT  -1.3375 28.8825 -1.2025 28.9475 ;
        RECT  -1.3375 29.0725 -1.2025 29.1375 ;
        RECT  -1.3375 28.8825 -1.2025 28.9475 ;
        RECT  -1.3375 29.0725 -1.2025 29.1375 ;
        RECT  -1.3375 29.0725 -1.2025 29.1375 ;
        RECT  -1.3375 29.2625 -1.2025 29.3275 ;
        RECT  -1.3375 29.0725 -1.2025 29.1375 ;
        RECT  -1.3375 29.2625 -1.2025 29.3275 ;
        RECT  -1.3375 29.4325 -1.2025 29.4975 ;
        RECT  -0.4675 29.4325 -0.3325 29.4975 ;
        RECT  -1.3375 28.8825 -1.2025 28.9475 ;
        RECT  -1.3375 29.2625 -1.2025 29.3275 ;
        RECT  -1.125 28.775 -0.99 28.84 ;
        RECT  -0.99 28.965 -0.855 29.03 ;
        RECT  -0.855 29.155 -0.72 29.22 ;
        RECT  -1.4525 30.0375 -1.0875 30.1025 ;
        RECT  -0.3075 30.0375 -0.1725 30.1025 ;
        RECT  -0.2425 29.6775 -0.1725 29.7425 ;
        RECT  -1.4525 29.6775 -1.3625 29.7425 ;
        RECT  -1.2225 29.8675 -0.275 29.9325 ;
        RECT  -0.755 29.61 -0.69 29.645 ;
        RECT  -0.755 29.9325 -0.69 30.17 ;
        RECT  -1.5175 29.61 -1.4525 30.17 ;
        RECT  -0.1725 29.61 -0.1075 30.17 ;
        RECT  -0.3775 29.6775 -0.2425 29.7425 ;
        RECT  -0.3775 29.8675 -0.2425 29.9325 ;
        RECT  -0.5125 29.6775 -0.3775 29.7425 ;
        RECT  -0.5125 29.8675 -0.3775 29.9325 ;
        RECT  -1.3625 29.6775 -1.0875 29.7425 ;
        RECT  -1.3625 29.8675 -1.0875 29.9325 ;
        RECT  -1.3625 29.6775 -1.0875 29.7425 ;
        RECT  -1.3625 29.8675 -1.0875 29.9325 ;
        RECT  -1.3625 30.0375 -1.0875 30.1025 ;
        RECT  -0.3775 30.0375 -0.2425 30.1025 ;
        RECT  -0.755 29.645 -0.69 29.78 ;
        RECT  -2.445 28.7175 -2.38 28.7825 ;
        RECT  -2.445 28.75 -2.38 29.41 ;
        RECT  -2.7275 28.7175 -2.4125 28.7825 ;
        RECT  -2.445 29.14 -2.38 29.41 ;
        RECT  -1.8825 29.2775 -1.485 29.3425 ;
        RECT  -2.83 29.0775 -2.7275 29.1425 ;
        RECT  -1.8825 28.5275 -1.5175 28.5925 ;
        RECT  -2.165 28.7175 -2.1 28.7825 ;
        RECT  -2.1325 28.7175 -1.8825 28.7825 ;
        RECT  -2.165 28.75 -2.1 28.85 ;
        RECT  -2.165 28.9175 -2.1 28.9825 ;
        RECT  -2.1325 28.9175 -1.8825 28.9825 ;
        RECT  -2.165 28.85 -2.1 28.95 ;
        RECT  -2.8625 28.5275 -2.7275 28.5925 ;
        RECT  -2.8625 28.9075 -2.7275 28.9725 ;
        RECT  -2.445 28.46 -2.38 28.63 ;
        RECT  -2.445 29.14 -2.38 29.41 ;
        RECT  -2.305 28.46 -2.24 29.02 ;
        RECT  -1.5175 28.46 -1.4525 29.41 ;
        RECT  -2.8625 28.46 -2.7975 29.41 ;
        RECT  -2.5275 28.5275 -2.3925 28.5925 ;
        RECT  -2.5275 28.7175 -2.3925 28.7825 ;
        RECT  -2.6625 28.5275 -2.5275 28.5925 ;
        RECT  -2.6625 28.7175 -2.5275 28.7825 ;
        RECT  -2.5275 28.7175 -2.3925 28.7825 ;
        RECT  -2.5275 28.9075 -2.3925 28.9725 ;
        RECT  -2.6625 28.7175 -2.5275 28.7825 ;
        RECT  -2.6625 28.9075 -2.5275 28.9725 ;
        RECT  -2.2625 28.5275 -1.9875 28.5925 ;
        RECT  -2.2625 28.7175 -1.9875 28.7825 ;
        RECT  -2.2625 28.5275 -1.9875 28.5925 ;
        RECT  -2.2625 28.7175 -1.9875 28.7825 ;
        RECT  -2.2625 28.9175 -1.9875 28.9825 ;
        RECT  -2.2625 29.1075 -1.9875 29.1725 ;
        RECT  -2.2625 28.9175 -1.9875 28.9825 ;
        RECT  -2.2625 29.1075 -1.9875 29.1725 ;
        RECT  -2.1575 29.2775 -1.8825 29.3425 ;
        RECT  -2.8625 29.0775 -2.7275 29.1425 ;
        RECT  -2.52 28.495 -2.455 28.63 ;
        RECT  -2.38 28.885 -2.315 29.02 ;
        RECT  -2.0175 29.1075 -1.8825 29.1725 ;
        RECT  -2.515 29.0725 -2.45 29.2075 ;
        RECT  -1.7675 30.2525 -1.485 30.3175 ;
        RECT  -2.83 30.2525 -2.65 30.3175 ;
        RECT  -1.7675 29.7025 -1.485 29.7675 ;
        RECT  -1.7675 30.0825 -1.485 30.1475 ;
        RECT  -2.83 29.7025 -2.5475 29.7675 ;
        RECT  -1.935 30.115 -1.87 30.18 ;
        RECT  -1.935 29.8925 -1.87 29.9575 ;
        RECT  -2.6825 30.115 -1.9025 30.18 ;
        RECT  -1.935 29.925 -1.87 30.1475 ;
        RECT  -1.9025 29.8925 -1.7675 29.9575 ;
        RECT  -1.92 29.635 -1.855 29.67 ;
        RECT  -2.2325 30.1475 -2.1675 30.385 ;
        RECT  -2.45 29.635 -2.385 29.91 ;
        RECT  -1.5175 29.635 -1.4525 30.385 ;
        RECT  -2.8625 29.635 -2.7975 30.385 ;
        RECT  -2.3925 29.7025 -2.2575 29.7675 ;
        RECT  -2.3925 29.8925 -2.2575 29.9575 ;
        RECT  -2.5275 29.7025 -2.3925 29.7675 ;
        RECT  -2.5275 29.8925 -2.3925 29.9575 ;
        RECT  -2.3925 29.8925 -2.2575 29.9575 ;
        RECT  -2.3925 30.0825 -2.2575 30.1475 ;
        RECT  -2.5275 29.8925 -2.3925 29.9575 ;
        RECT  -2.5275 30.0825 -2.3925 30.1475 ;
        RECT  -2.0575 29.7025 -1.9225 29.7675 ;
        RECT  -2.0575 29.8925 -1.9225 29.9575 ;
        RECT  -2.0575 29.7025 -1.9225 29.7675 ;
        RECT  -2.0575 29.8925 -1.9225 29.9575 ;
        RECT  -2.0575 29.8925 -1.9225 29.9575 ;
        RECT  -2.0575 30.0825 -1.9225 30.1475 ;
        RECT  -2.0575 29.8925 -1.9225 29.9575 ;
        RECT  -2.0575 30.0825 -1.9225 30.1475 ;
        RECT  -1.9025 30.2525 -1.7675 30.3175 ;
        RECT  -2.8175 30.2525 -2.6825 30.3175 ;
        RECT  -1.995 29.67 -1.93 29.805 ;
        RECT  -2.525 29.91 -2.46 30.045 ;
        RECT  -1.8825 30.6775 -1.5175 30.7425 ;
        RECT  -2.7975 30.6775 -2.6625 30.7425 ;
        RECT  -2.7975 31.0375 -2.7275 31.1025 ;
        RECT  -1.6075 31.0375 -1.5175 31.1025 ;
        RECT  -2.695 30.8475 -1.7475 30.9125 ;
        RECT  -2.28 31.135 -2.215 31.17 ;
        RECT  -2.28 30.61 -2.215 30.8475 ;
        RECT  -1.5175 30.61 -1.4525 31.17 ;
        RECT  -2.8625 30.61 -2.7975 31.17 ;
        RECT  -2.7275 31.0375 -2.5925 31.1025 ;
        RECT  -2.7275 30.8475 -2.5925 30.9125 ;
        RECT  -2.5925 31.0375 -2.4575 31.1025 ;
        RECT  -2.5925 30.8475 -2.4575 30.9125 ;
        RECT  -1.8825 31.0375 -1.6075 31.1025 ;
        RECT  -1.8825 30.8475 -1.6075 30.9125 ;
        RECT  -1.8825 31.0375 -1.6075 31.1025 ;
        RECT  -1.8825 30.8475 -1.6075 30.9125 ;
        RECT  -1.8825 30.6775 -1.6075 30.7425 ;
        RECT  -2.7275 30.6775 -2.5925 30.7425 ;
        RECT  -2.28 31.0 -2.215 31.135 ;
        RECT  -1.8825 31.2375 -1.5175 31.3025 ;
        RECT  -2.7975 31.2375 -2.6625 31.3025 ;
        RECT  -2.7975 31.5975 -2.7275 31.6625 ;
        RECT  -1.6075 31.5975 -1.5175 31.6625 ;
        RECT  -2.695 31.4075 -1.7475 31.4725 ;
        RECT  -2.28 31.695 -2.215 31.73 ;
        RECT  -2.28 31.17 -2.215 31.4075 ;
        RECT  -1.5175 31.17 -1.4525 31.73 ;
        RECT  -2.8625 31.17 -2.7975 31.73 ;
        RECT  -2.7275 31.5975 -2.5925 31.6625 ;
        RECT  -2.7275 31.4075 -2.5925 31.4725 ;
        RECT  -2.5925 31.5975 -2.4575 31.6625 ;
        RECT  -2.5925 31.4075 -2.4575 31.4725 ;
        RECT  -1.8825 31.5975 -1.6075 31.6625 ;
        RECT  -1.8825 31.4075 -1.6075 31.4725 ;
        RECT  -1.8825 31.5975 -1.6075 31.6625 ;
        RECT  -1.8825 31.4075 -1.6075 31.4725 ;
        RECT  -1.8825 31.2375 -1.6075 31.3025 ;
        RECT  -2.7275 31.2375 -2.5925 31.3025 ;
        RECT  -2.28 31.56 -2.215 31.695 ;
        RECT  -4.045 29.855 -2.96 29.92 ;
        RECT  -4.175 29.9925 -3.8925 30.0575 ;
        RECT  -3.1 29.9925 -2.83 30.0575 ;
        RECT  -4.175 29.2525 -3.8925 29.3175 ;
        RECT  -4.175 29.6325 -3.8925 29.6975 ;
        RECT  -3.1125 29.2525 -2.83 29.3175 ;
        RECT  -3.745 29.02 -3.68 29.355 ;
        RECT  -3.475 29.02 -3.41 29.735 ;
        RECT  -3.61 29.02 -3.545 29.545 ;
        RECT  -4.2075 29.02 -4.1425 30.17 ;
        RECT  -2.8625 29.02 -2.7975 30.17 ;
        RECT  -3.5475 29.855 -3.4825 30.17 ;
        RECT  -3.1575 29.2525 -3.0225 29.3175 ;
        RECT  -3.1575 29.4425 -3.0225 29.5075 ;
        RECT  -3.2925 29.2525 -3.1575 29.3175 ;
        RECT  -3.2925 29.4425 -3.1575 29.5075 ;
        RECT  -3.1575 29.4425 -3.0225 29.5075 ;
        RECT  -3.1575 29.6325 -3.0225 29.6975 ;
        RECT  -3.2925 29.4425 -3.1575 29.5075 ;
        RECT  -3.2925 29.6325 -3.1575 29.6975 ;
        RECT  -3.1575 29.6325 -3.0225 29.6975 ;
        RECT  -3.1575 29.8225 -3.0225 29.8875 ;
        RECT  -3.2925 29.6325 -3.1575 29.6975 ;
        RECT  -3.2925 29.8225 -3.1575 29.8875 ;
        RECT  -4.0275 29.2525 -3.8925 29.3175 ;
        RECT  -4.0275 29.4425 -3.8925 29.5075 ;
        RECT  -4.0275 29.2525 -3.8925 29.3175 ;
        RECT  -4.0275 29.4425 -3.8925 29.5075 ;
        RECT  -4.0275 29.4425 -3.8925 29.5075 ;
        RECT  -4.0275 29.6325 -3.8925 29.6975 ;
        RECT  -4.0275 29.4425 -3.8925 29.5075 ;
        RECT  -4.0275 29.6325 -3.8925 29.6975 ;
        RECT  -4.0275 29.6325 -3.8925 29.6975 ;
        RECT  -4.0275 29.8225 -3.8925 29.8875 ;
        RECT  -4.0275 29.6325 -3.8925 29.6975 ;
        RECT  -4.0275 29.8225 -3.8925 29.8875 ;
        RECT  -4.0275 29.9925 -3.8925 30.0575 ;
        RECT  -3.1575 29.9925 -3.0225 30.0575 ;
        RECT  -4.0275 29.4425 -3.8925 29.5075 ;
        RECT  -4.0275 29.8225 -3.8925 29.8875 ;
        RECT  -3.815 29.335 -3.68 29.4 ;
        RECT  -3.68 29.525 -3.545 29.59 ;
        RECT  -3.545 29.715 -3.41 29.78 ;
        RECT  -4.1425 30.5975 -3.7775 30.6625 ;
        RECT  -2.9975 30.5975 -2.8625 30.6625 ;
        RECT  -2.9325 30.2375 -2.8625 30.3025 ;
        RECT  -4.1425 30.2375 -4.0525 30.3025 ;
        RECT  -3.9125 30.4275 -2.965 30.4925 ;
        RECT  -3.445 30.17 -3.38 30.205 ;
        RECT  -3.445 30.4925 -3.38 30.73 ;
        RECT  -4.2075 30.17 -4.1425 30.73 ;
        RECT  -2.8625 30.17 -2.7975 30.73 ;
        RECT  -3.0675 30.2375 -2.9325 30.3025 ;
        RECT  -3.0675 30.4275 -2.9325 30.4925 ;
        RECT  -3.2025 30.2375 -3.0675 30.3025 ;
        RECT  -3.2025 30.4275 -3.0675 30.4925 ;
        RECT  -4.0525 30.2375 -3.7775 30.3025 ;
        RECT  -4.0525 30.4275 -3.7775 30.4925 ;
        RECT  -4.0525 30.2375 -3.7775 30.3025 ;
        RECT  -4.0525 30.4275 -3.7775 30.4925 ;
        RECT  -4.0525 30.5975 -3.7775 30.6625 ;
        RECT  -3.0675 30.5975 -2.9325 30.6625 ;
        RECT  -3.445 30.205 -3.38 30.34 ;
        RECT  -4.1425 31.1575 -3.7775 31.2225 ;
        RECT  -2.9975 31.1575 -2.8625 31.2225 ;
        RECT  -2.9325 30.7975 -2.8625 30.8625 ;
        RECT  -4.1425 30.7975 -4.0525 30.8625 ;
        RECT  -3.9125 30.9875 -2.965 31.0525 ;
        RECT  -3.445 30.73 -3.38 30.765 ;
        RECT  -3.445 31.0525 -3.38 31.29 ;
        RECT  -4.2075 30.73 -4.1425 31.29 ;
        RECT  -2.8625 30.73 -2.7975 31.29 ;
        RECT  -3.0675 30.7975 -2.9325 30.8625 ;
        RECT  -3.0675 30.9875 -2.9325 31.0525 ;
        RECT  -3.2025 30.7975 -3.0675 30.8625 ;
        RECT  -3.2025 30.9875 -3.0675 31.0525 ;
        RECT  -4.0525 30.7975 -3.7775 30.8625 ;
        RECT  -4.0525 30.9875 -3.7775 31.0525 ;
        RECT  -4.0525 30.7975 -3.7775 30.8625 ;
        RECT  -4.0525 30.9875 -3.7775 31.0525 ;
        RECT  -4.0525 31.1575 -3.7775 31.2225 ;
        RECT  -3.0675 31.1575 -2.9325 31.2225 ;
        RECT  -3.445 30.765 -3.38 30.9 ;
        RECT  -4.1425 31.7175 -3.7775 31.7825 ;
        RECT  -2.9975 31.7175 -2.8625 31.7825 ;
        RECT  -2.9325 31.3575 -2.8625 31.4225 ;
        RECT  -4.1425 31.3575 -4.0525 31.4225 ;
        RECT  -3.9125 31.5475 -2.965 31.6125 ;
        RECT  -3.445 31.29 -3.38 31.325 ;
        RECT  -3.445 31.6125 -3.38 31.85 ;
        RECT  -4.2075 31.29 -4.1425 31.85 ;
        RECT  -2.8625 31.29 -2.7975 31.85 ;
        RECT  -3.0675 31.3575 -2.9325 31.4225 ;
        RECT  -3.0675 31.5475 -2.9325 31.6125 ;
        RECT  -3.2025 31.3575 -3.0675 31.4225 ;
        RECT  -3.2025 31.5475 -3.0675 31.6125 ;
        RECT  -4.0525 31.3575 -3.7775 31.4225 ;
        RECT  -4.0525 31.5475 -3.7775 31.6125 ;
        RECT  -4.0525 31.3575 -3.7775 31.4225 ;
        RECT  -4.0525 31.5475 -3.7775 31.6125 ;
        RECT  -4.0525 31.7175 -3.7775 31.7825 ;
        RECT  -3.0675 31.7175 -2.9325 31.7825 ;
        RECT  -3.445 31.325 -3.38 31.46 ;
        RECT  -3.845 25.67 -3.78 25.805 ;
        RECT  -3.69 25.67 -3.625 25.805 ;
        RECT  -2.83 25.67 -2.765 25.805 ;
        RECT  -2.435 25.67 -2.37 25.805 ;
        RECT  -3.24 34.5075 -2.795 34.5725 ;
        RECT  -3.24 36.9175 -2.795 36.9825 ;
        RECT  -3.24 37.3625 -2.83 37.4275 ;
        RECT  -4.155 35.7125 -3.24 35.7775 ;
        RECT  -4.155 33.0225 -3.24 33.0875 ;
        RECT  -2.28 33.95 -2.215 34.735 ;
        RECT  -2.28 34.2275 -2.215 34.2925 ;
        RECT  -2.28 33.95 -2.215 34.26 ;
        RECT  -3.15 34.2275 -2.2475 34.2925 ;
        RECT  -2.08 34.0125 -1.485 34.0775 ;
        RECT  -2.09 33.2275 -2.025 33.2925 ;
        RECT  -2.28 33.2275 -2.215 33.2925 ;
        RECT  -2.09 33.26 -2.025 33.8475 ;
        RECT  -2.2475 33.2275 -2.0575 33.2925 ;
        RECT  -2.28 33.055 -2.215 33.26 ;
        RECT  -3.0025 33.2275 -2.2475 33.2925 ;
        RECT  -3.425 32.63 -3.0025 32.695 ;
        RECT  -0.755 31.935 -0.69 34.8 ;
        RECT  -4.22 31.935 -4.155 37.1225 ;
        RECT  -1.5175 31.935 -1.4525 34.735 ;
        RECT  -2.865 31.935 -2.795 33.055 ;
        RECT  -0.1725 31.935 -0.1075 34.735 ;
        RECT  -2.28 31.935 -2.215 32.495 ;
        RECT  -1.8825 33.4825 -1.5175 33.5475 ;
        RECT  -2.7975 33.4825 -2.6625 33.5475 ;
        RECT  -2.7975 33.1225 -2.7275 33.1875 ;
        RECT  -1.6075 33.1225 -1.5175 33.1875 ;
        RECT  -2.695 33.3125 -1.7475 33.3775 ;
        RECT  -2.28 33.055 -2.215 33.09 ;
        RECT  -2.28 33.3775 -2.215 33.615 ;
        RECT  -1.5175 33.055 -1.4525 33.615 ;
        RECT  -2.8625 33.055 -2.7975 33.615 ;
        RECT  -2.5275 33.1225 -2.3925 33.1875 ;
        RECT  -2.5275 33.3125 -2.3925 33.3775 ;
        RECT  -2.6625 33.1225 -2.5275 33.1875 ;
        RECT  -2.6625 33.3125 -2.5275 33.3775 ;
        RECT  -2.2625 33.1225 -1.9875 33.1875 ;
        RECT  -2.2625 33.3125 -1.9875 33.3775 ;
        RECT  -2.2625 33.1225 -1.9875 33.1875 ;
        RECT  -2.2625 33.3125 -1.9875 33.3775 ;
        RECT  -2.1575 33.4825 -1.8825 33.5475 ;
        RECT  -2.8625 33.4825 -2.7275 33.5475 ;
        RECT  -2.355 33.09 -2.29 33.225 ;
        RECT  -2.125 33.6225 -1.99 33.6875 ;
        RECT  -2.125 33.4325 -1.99 33.4975 ;
        RECT  -2.125 33.6225 -1.99 33.6875 ;
        RECT  -2.125 33.4325 -1.99 33.4975 ;
        RECT  -2.8625 33.4525 -2.7975 33.5175 ;
        RECT  -0.1725 33.4525 -0.1075 33.5175 ;
        RECT  -2.8625 33.485 -2.7975 33.615 ;
        RECT  -2.83 33.4525 -0.14 33.5175 ;
        RECT  -0.1725 33.485 -0.1075 33.615 ;
        RECT  -2.28 34.4975 -2.215 34.735 ;
        RECT  -1.5175 33.615 -1.4525 34.735 ;
        RECT  -2.8625 33.615 -2.7975 34.735 ;
        RECT  -0.1725 33.615 -0.1075 34.735 ;
        RECT  -0.755 34.67 -0.69 34.735 ;
        RECT  -0.7575 34.6 -0.6925 34.735 ;
        RECT  -1.4525 34.2425 -1.0875 34.3075 ;
        RECT  -0.3075 34.2425 -0.1725 34.3075 ;
        RECT  -0.2425 34.6025 -0.1725 34.6675 ;
        RECT  -1.4525 34.6025 -1.3625 34.6675 ;
        RECT  -1.2225 34.4125 -0.275 34.4775 ;
        RECT  -0.755 34.7 -0.69 34.735 ;
        RECT  -0.755 34.3475 -0.69 34.4125 ;
        RECT  -1.5175 34.175 -1.4525 34.735 ;
        RECT  -0.1725 34.175 -0.1075 34.735 ;
        RECT  -0.5775 34.6025 -0.4425 34.6675 ;
        RECT  -0.5775 34.4125 -0.4425 34.4775 ;
        RECT  -0.4425 34.6025 -0.3075 34.6675 ;
        RECT  -0.4425 34.4125 -0.3075 34.4775 ;
        RECT  -0.9825 34.6025 -0.7075 34.6675 ;
        RECT  -0.9825 34.4125 -0.7075 34.4775 ;
        RECT  -0.9825 34.6025 -0.7075 34.6675 ;
        RECT  -0.9825 34.4125 -0.7075 34.4775 ;
        RECT  -1.0875 34.2425 -0.8125 34.3075 ;
        RECT  -0.2425 34.2425 -0.1075 34.3075 ;
        RECT  -0.68 34.565 -0.615 34.7 ;
        RECT  -0.7575 34.04 -0.6925 34.175 ;
        RECT  -1.4525 33.6825 -1.0875 33.7475 ;
        RECT  -0.3075 33.6825 -0.1725 33.7475 ;
        RECT  -0.2425 34.0425 -0.1725 34.1075 ;
        RECT  -1.4525 34.0425 -1.3625 34.1075 ;
        RECT  -1.2225 33.8525 -0.275 33.9175 ;
        RECT  -0.755 34.14 -0.69 34.175 ;
        RECT  -0.755 33.7875 -0.69 33.8525 ;
        RECT  -1.5175 33.615 -1.4525 34.175 ;
        RECT  -0.1725 33.615 -0.1075 34.175 ;
        RECT  -0.5775 34.0425 -0.4425 34.1075 ;
        RECT  -0.5775 33.8525 -0.4425 33.9175 ;
        RECT  -0.4425 34.0425 -0.3075 34.1075 ;
        RECT  -0.4425 33.8525 -0.3075 33.9175 ;
        RECT  -0.9825 34.0425 -0.7075 34.1075 ;
        RECT  -0.9825 33.8525 -0.7075 33.9175 ;
        RECT  -0.9825 34.0425 -0.7075 34.1075 ;
        RECT  -0.9825 33.8525 -0.7075 33.9175 ;
        RECT  -1.0875 33.6825 -0.8125 33.7475 ;
        RECT  -0.2425 33.6825 -0.1075 33.7475 ;
        RECT  -0.68 34.005 -0.615 34.14 ;
        RECT  -2.2775 33.615 -2.2125 33.75 ;
        RECT  -1.8825 34.0425 -1.5175 34.1075 ;
        RECT  -2.7975 34.0425 -2.6625 34.1075 ;
        RECT  -2.7975 33.6825 -2.7275 33.7475 ;
        RECT  -1.6075 33.6825 -1.5175 33.7475 ;
        RECT  -2.695 33.8725 -1.7475 33.9375 ;
        RECT  -2.28 33.615 -2.215 33.65 ;
        RECT  -2.28 33.9375 -2.215 34.0025 ;
        RECT  -1.5175 33.615 -1.4525 34.175 ;
        RECT  -2.8625 33.615 -2.7975 34.175 ;
        RECT  -2.5275 33.6825 -2.3925 33.7475 ;
        RECT  -2.5275 33.8725 -2.3925 33.9375 ;
        RECT  -2.6625 33.6825 -2.5275 33.7475 ;
        RECT  -2.6625 33.8725 -2.5275 33.9375 ;
        RECT  -2.2625 33.6825 -1.9875 33.7475 ;
        RECT  -2.2625 33.8725 -1.9875 33.9375 ;
        RECT  -2.2625 33.6825 -1.9875 33.7475 ;
        RECT  -2.2625 33.8725 -1.9875 33.9375 ;
        RECT  -2.1575 34.0425 -1.8825 34.1075 ;
        RECT  -2.8625 34.0425 -2.7275 34.1075 ;
        RECT  -2.355 33.65 -2.29 33.785 ;
        RECT  -2.2775 34.175 -2.2125 34.31 ;
        RECT  -1.8825 34.6025 -1.5175 34.6675 ;
        RECT  -2.7975 34.6025 -2.6625 34.6675 ;
        RECT  -2.7975 34.2425 -2.7275 34.3075 ;
        RECT  -1.6075 34.2425 -1.5175 34.3075 ;
        RECT  -2.695 34.4325 -1.7475 34.4975 ;
        RECT  -2.28 34.175 -2.215 34.21 ;
        RECT  -2.28 34.4975 -2.215 34.5625 ;
        RECT  -1.5175 34.175 -1.4525 34.735 ;
        RECT  -2.8625 34.175 -2.7975 34.735 ;
        RECT  -2.5275 34.2425 -2.3925 34.3075 ;
        RECT  -2.5275 34.4325 -2.3925 34.4975 ;
        RECT  -2.6625 34.2425 -2.5275 34.3075 ;
        RECT  -2.6625 34.4325 -2.5275 34.4975 ;
        RECT  -2.2625 34.2425 -1.9875 34.3075 ;
        RECT  -2.2625 34.4325 -1.9875 34.4975 ;
        RECT  -2.2625 34.2425 -1.9875 34.3075 ;
        RECT  -2.2625 34.4325 -1.9875 34.4975 ;
        RECT  -2.1575 34.6025 -1.8825 34.6675 ;
        RECT  -2.8625 34.6025 -2.7275 34.6675 ;
        RECT  -2.355 34.21 -2.29 34.345 ;
        RECT  -0.7575 34.2775 -0.6925 34.4125 ;
        RECT  -0.7575 33.7175 -0.6925 33.8525 ;
        RECT  -2.2775 33.9375 -2.2125 34.0725 ;
        RECT  -3.895 34.6575 -3.83 34.7925 ;
        RECT  -3.71 34.6575 -3.645 34.7925 ;
        RECT  -3.54 34.6625 -3.475 34.7975 ;
        RECT  -3.355 34.6625 -3.29 34.7975 ;
        RECT  -3.975 35.0475 -3.91 35.1825 ;
        RECT  -3.79 35.0475 -3.725 35.1825 ;
        RECT  -3.46 35.0475 -3.395 35.1825 ;
        RECT  -3.275 35.0475 -3.21 35.1825 ;
        RECT  -3.975 35.5125 -3.91 35.6475 ;
        RECT  -3.79 35.5125 -3.725 35.6475 ;
        RECT  -3.46 35.5125 -3.395 35.6475 ;
        RECT  -3.275 35.5125 -3.21 35.6475 ;
        RECT  -3.2725 34.6625 -3.2075 34.7975 ;
        RECT  -3.9775 35.1375 -3.9125 35.2725 ;
        RECT  -3.2725 35.1375 -3.2075 35.2725 ;
        RECT  -3.725 34.6575 -3.66 34.7925 ;
        RECT  -3.525 34.6625 -3.46 34.7975 ;
        RECT  -3.7725 35.2525 -3.6375 35.3175 ;
        RECT  -3.5475 35.4025 -3.4125 35.4675 ;
        RECT  -3.65 34.5075 -3.515 34.5725 ;
        RECT  -3.6575 35.7125 -3.5225 35.7775 ;
        RECT  -3.655 34.3675 -3.52 34.4325 ;
        RECT  -4.0125 34.3675 -3.8775 34.4325 ;
        RECT  -3.2925 34.6625 -3.24 34.7975 ;
        RECT  -3.3075 34.3675 -3.1725 34.4325 ;
        RECT  -3.6225 35.7125 -3.5575 35.7775 ;
        RECT  -3.275 34.5075 -3.205 34.5725 ;
        RECT  -3.83 34.8825 -3.725 34.9475 ;
        RECT  -3.79 34.9475 -3.725 35.0475 ;
        RECT  -3.895 34.7925 -3.83 34.9475 ;
        RECT  -3.46 34.8825 -3.355 34.9475 ;
        RECT  -3.46 34.9475 -3.395 35.0475 ;
        RECT  -3.355 34.7975 -3.29 34.9475 ;
        RECT  -3.975 35.6475 -3.91 35.7125 ;
        RECT  -3.275 35.6475 -3.21 35.7125 ;
        RECT  -3.79 35.0475 -3.725 35.5375 ;
        RECT  -3.46 35.0475 -3.395 35.5375 ;
        RECT  -4.035 34.5075 -3.15 34.5725 ;
        RECT  -4.035 35.7125 -3.15 35.7775 ;
        RECT  -4.035 34.3675 -3.15 34.4325 ;
        RECT  -4.035 34.5075 -3.15 34.5725 ;
        RECT  -4.035 35.7125 -3.15 35.7775 ;
        RECT  -4.035 34.2275 -3.15 34.2925 ;
        RECT  -4.035 31.8175 -3.15 31.8825 ;
        RECT  -4.035 33.0225 -3.15 33.0875 ;
        RECT  -4.035 34.3675 -3.15 34.4325 ;
        RECT  -4.035 31.6775 -3.15 31.7425 ;
        RECT  -3.975 33.1525 -3.91 33.2875 ;
        RECT  -3.79 33.1525 -3.725 33.2875 ;
        RECT  -3.275 33.1525 -3.21 33.2875 ;
        RECT  -3.46 33.1525 -3.395 33.2875 ;
        RECT  -3.79 33.6175 -3.725 33.7525 ;
        RECT  -3.975 33.6175 -3.91 33.7525 ;
        RECT  -3.46 33.6175 -3.395 33.7525 ;
        RECT  -3.275 33.6175 -3.21 33.7525 ;
        RECT  -3.895 34.0075 -3.83 34.1425 ;
        RECT  -3.71 34.0075 -3.645 34.1425 ;
        RECT  -3.54 34.0075 -3.475 34.1425 ;
        RECT  -3.355 34.0075 -3.29 34.1425 ;
        RECT  -3.9775 33.515 -3.9125 33.65 ;
        RECT  -3.9775 33.515 -3.9125 33.65 ;
        RECT  -3.9775 33.515 -3.9125 33.65 ;
        RECT  -3.9775 33.515 -3.9125 33.65 ;
        RECT  -3.9775 33.515 -3.9125 33.65 ;
        RECT  -3.9775 33.515 -3.9125 33.65 ;
        RECT  -3.655 33.0225 -3.52 33.0875 ;
        RECT  -3.3075 34.3675 -3.1725 34.4325 ;
        RECT  -4.0125 34.3675 -3.8775 34.4325 ;
        RECT  -3.6425 34.2275 -3.5075 34.2925 ;
        RECT  -3.9775 33.515 -3.9125 33.65 ;
        RECT  -3.9775 33.515 -3.9125 33.65 ;
        RECT  -3.9775 33.515 -3.9125 33.65 ;
        RECT  -3.9775 33.515 -3.9125 33.65 ;
        RECT  -3.5475 33.3375 -3.4125 33.4025 ;
        RECT  -3.5475 33.3375 -3.4125 33.4025 ;
        RECT  -3.7725 33.4875 -3.6375 33.5525 ;
        RECT  -3.7725 33.4875 -3.6375 33.5525 ;
        RECT  -3.9775 33.515 -3.9125 33.65 ;
        RECT  -3.9775 33.515 -3.9125 33.65 ;
        RECT  -3.9775 33.515 -3.9125 33.65 ;
        RECT  -3.9775 33.515 -3.9125 33.65 ;
        RECT  -3.5275 34.0075 -3.4625 34.1425 ;
        RECT  -3.2725 33.515 -3.2075 33.65 ;
        RECT  -3.2725 33.515 -3.2075 33.65 ;
        RECT  -3.2725 33.515 -3.2075 33.65 ;
        RECT  -3.2725 33.515 -3.2075 33.65 ;
        RECT  -3.2725 33.515 -3.2075 33.65 ;
        RECT  -3.2725 33.515 -3.2075 33.65 ;
        RECT  -3.9775 33.515 -3.9125 33.65 ;
        RECT  -3.9775 33.515 -3.9125 33.65 ;
        RECT  -3.9775 33.515 -3.9125 33.65 ;
        RECT  -3.9775 33.515 -3.9125 33.65 ;
        RECT  -3.7225 34.0075 -3.6575 34.1425 ;
        RECT  -3.66 34.3675 -3.525 34.4325 ;
        RECT  -3.66 34.3675 -3.525 34.4325 ;
        RECT  -4.0125 34.3675 -3.8775 34.4325 ;
        RECT  -3.655 33.0225 -3.52 33.0875 ;
        RECT  -4.0125 34.3675 -3.8775 34.4325 ;
        RECT  -4.0125 34.3675 -3.8775 34.4325 ;
        RECT  -3.9775 33.515 -3.9125 33.65 ;
        RECT  -3.9775 33.515 -3.9125 33.65 ;
        RECT  -3.9775 33.515 -3.9125 33.65 ;
        RECT  -3.9775 33.515 -3.9125 33.65 ;
        RECT  -3.9775 33.515 -3.9125 33.65 ;
        RECT  -3.9775 33.515 -3.9125 33.65 ;
        RECT  -3.3075 34.3675 -3.1725 34.4325 ;
        RECT  -3.6325 33.025 -3.5325 33.0875 ;
        RECT  -3.6325 33.0225 -3.5325 33.085 ;
        RECT  -3.9125 34.2275 -3.86 34.29 ;
        RECT  -3.6325 33.025 -3.5325 33.0875 ;
        RECT  -3.98 33.0875 -3.91 33.2875 ;
        RECT  -3.98 33.6175 -3.91 33.7525 ;
        RECT  -3.98 33.6175 -3.91 33.7525 ;
        RECT  -4.035 34.3675 -3.15 34.4325 ;
        RECT  -3.9 33.8525 -3.725 33.9175 ;
        RECT  -3.275 33.6175 -3.205 33.7525 ;
        RECT  -3.46 33.1775 -3.395 33.9175 ;
        RECT  -3.6325 33.0225 -3.5325 33.085 ;
        RECT  -3.2075 34.2275 -3.155 34.29 ;
        RECT  -3.98 33.6175 -3.91 33.7525 ;
        RECT  -4.035 33.0225 -3.15 33.0875 ;
        RECT  -3.79 33.2875 -3.725 33.9175 ;
        RECT  -3.98 33.6175 -3.91 33.7525 ;
        RECT  -3.98 33.6175 -3.91 33.7525 ;
        RECT  -3.36 33.8525 -3.29 34.1425 ;
        RECT  -3.275 33.6175 -3.205 33.7525 ;
        RECT  -4.035 34.2275 -3.15 34.2925 ;
        RECT  -3.98 33.6175 -3.91 33.7525 ;
        RECT  -3.98 33.0875 -3.91 33.2875 ;
        RECT  -3.275 33.0875 -3.205 33.2875 ;
        RECT  -3.9 33.8525 -3.83 34.1425 ;
        RECT  -3.46 33.8525 -3.29 33.9175 ;
        RECT  -4.035 34.2275 -3.15 34.2925 ;
        RECT  -4.035 34.3675 -3.15 34.4325 ;
        RECT  -4.035 33.0225 -3.15 33.0875 ;
        RECT  -3.975 32.8225 -3.91 32.9575 ;
        RECT  -3.79 32.8225 -3.725 32.9575 ;
        RECT  -3.275 32.8225 -3.21 32.9575 ;
        RECT  -3.46 32.8225 -3.395 32.9575 ;
        RECT  -3.79 32.3575 -3.725 32.4925 ;
        RECT  -3.975 32.3575 -3.91 32.4925 ;
        RECT  -3.46 32.3575 -3.395 32.4925 ;
        RECT  -3.275 32.3575 -3.21 32.4925 ;
        RECT  -3.895 31.9675 -3.83 32.1025 ;
        RECT  -3.71 31.9675 -3.645 32.1025 ;
        RECT  -3.54 31.9675 -3.475 32.1025 ;
        RECT  -3.355 31.9675 -3.29 32.1025 ;
        RECT  -3.9775 32.46 -3.9125 32.595 ;
        RECT  -3.9775 32.46 -3.9125 32.595 ;
        RECT  -3.9775 32.46 -3.9125 32.595 ;
        RECT  -3.9775 32.46 -3.9125 32.595 ;
        RECT  -3.9775 32.46 -3.9125 32.595 ;
        RECT  -3.9775 32.46 -3.9125 32.595 ;
        RECT  -3.655 33.0225 -3.52 33.0875 ;
        RECT  -3.3075 31.6775 -3.1725 31.7425 ;
        RECT  -4.0125 31.6775 -3.8775 31.7425 ;
        RECT  -3.6425 31.8175 -3.5075 31.8825 ;
        RECT  -3.9775 32.46 -3.9125 32.595 ;
        RECT  -3.9775 32.46 -3.9125 32.595 ;
        RECT  -3.9775 32.46 -3.9125 32.595 ;
        RECT  -3.9775 32.46 -3.9125 32.595 ;
        RECT  -3.5475 32.7075 -3.4125 32.7725 ;
        RECT  -3.5475 32.7075 -3.4125 32.7725 ;
        RECT  -3.7725 32.5575 -3.6375 32.6225 ;
        RECT  -3.7725 32.5575 -3.6375 32.6225 ;
        RECT  -3.9775 32.46 -3.9125 32.595 ;
        RECT  -3.9775 32.46 -3.9125 32.595 ;
        RECT  -3.9775 32.46 -3.9125 32.595 ;
        RECT  -3.9775 32.46 -3.9125 32.595 ;
        RECT  -3.5275 31.9675 -3.4625 32.1025 ;
        RECT  -3.2725 32.46 -3.2075 32.595 ;
        RECT  -3.2725 32.46 -3.2075 32.595 ;
        RECT  -3.2725 32.46 -3.2075 32.595 ;
        RECT  -3.2725 32.46 -3.2075 32.595 ;
        RECT  -3.2725 32.46 -3.2075 32.595 ;
        RECT  -3.2725 32.46 -3.2075 32.595 ;
        RECT  -3.9775 32.46 -3.9125 32.595 ;
        RECT  -3.9775 32.46 -3.9125 32.595 ;
        RECT  -3.9775 32.46 -3.9125 32.595 ;
        RECT  -3.9775 32.46 -3.9125 32.595 ;
        RECT  -3.7225 31.9675 -3.6575 32.1025 ;
        RECT  -3.66 31.6775 -3.525 31.7425 ;
        RECT  -3.66 31.6775 -3.525 31.7425 ;
        RECT  -4.0125 31.6775 -3.8775 31.7425 ;
        RECT  -3.655 33.0225 -3.52 33.0875 ;
        RECT  -4.0125 31.6775 -3.8775 31.7425 ;
        RECT  -4.0125 31.6775 -3.8775 31.7425 ;
        RECT  -3.9775 32.46 -3.9125 32.595 ;
        RECT  -3.9775 32.46 -3.9125 32.595 ;
        RECT  -3.9775 32.46 -3.9125 32.595 ;
        RECT  -3.9775 32.46 -3.9125 32.595 ;
        RECT  -3.9775 32.46 -3.9125 32.595 ;
        RECT  -3.9775 32.46 -3.9125 32.595 ;
        RECT  -3.3075 31.6775 -3.1725 31.7425 ;
        RECT  -3.6325 33.0225 -3.5325 33.085 ;
        RECT  -3.6325 33.025 -3.5325 33.0875 ;
        RECT  -3.9125 31.82 -3.86 31.8825 ;
        RECT  -3.6325 33.0225 -3.5325 33.085 ;
        RECT  -3.98 32.8225 -3.91 33.0225 ;
        RECT  -3.98 32.3575 -3.91 32.4925 ;
        RECT  -3.98 32.3575 -3.91 32.4925 ;
        RECT  -4.035 31.6775 -3.15 31.7425 ;
        RECT  -3.9 32.1925 -3.725 32.2575 ;
        RECT  -3.275 32.3575 -3.205 32.4925 ;
        RECT  -3.46 32.1925 -3.395 32.9325 ;
        RECT  -3.6325 33.025 -3.5325 33.0875 ;
        RECT  -3.2075 31.82 -3.155 31.8825 ;
        RECT  -3.98 32.3575 -3.91 32.4925 ;
        RECT  -4.035 33.0225 -3.15 33.0875 ;
        RECT  -3.79 32.1925 -3.725 32.8225 ;
        RECT  -3.98 32.3575 -3.91 32.4925 ;
        RECT  -3.98 32.3575 -3.91 32.4925 ;
        RECT  -3.36 31.9675 -3.29 32.2575 ;
        RECT  -3.275 32.3575 -3.205 32.4925 ;
        RECT  -4.035 31.8175 -3.15 31.8825 ;
        RECT  -3.98 32.3575 -3.91 32.4925 ;
        RECT  -3.98 32.8225 -3.91 33.0225 ;
        RECT  -3.275 32.8225 -3.205 33.0225 ;
        RECT  -3.9 31.9675 -3.83 32.2575 ;
        RECT  -3.46 32.1925 -3.29 32.2575 ;
        RECT  -4.035 31.8175 -3.15 31.8825 ;
        RECT  -4.035 31.6775 -3.15 31.7425 ;
        RECT  -4.035 33.0225 -3.15 33.0875 ;
        RECT  -2.8625 34.3725 -2.7975 34.5075 ;
        RECT  -2.8625 36.7825 -2.7975 36.9175 ;
        RECT  -2.8625 34.6 -2.7975 34.735 ;
        RECT  -2.8625 32.225 -2.7975 32.36 ;
        RECT  -2.8975 37.2925 -2.7625 37.3575 ;
        RECT  -3.3075 37.2925 -3.1725 37.3575 ;
        RECT  -2.28 33.7475 -2.215 33.8825 ;
        RECT  -3.07 33.1575 -2.935 33.2225 ;
        RECT  -3.07 32.56 -2.935 32.625 ;
        RECT  -3.4925 32.56 -3.3575 32.625 ;
        RECT  -0.755 26.5825 -0.69 26.7175 ;
        RECT  -0.755 23.0 -0.69 23.135 ;
        RECT  -1.7225 19.4 -1.6575 19.535 ;
        RECT  -2.445 26.5825 -2.38 26.7175 ;
        RECT  -2.305 26.9925 -2.24 27.1275 ;
        RECT  -1.92 29.635 -1.855 29.77 ;
        RECT  -2.45 29.635 -2.385 29.77 ;
        RECT  -1.055 28.0175 -0.99 28.1525 ;
        RECT  -0.92 27.8125 -0.855 27.9475 ;
        RECT  -0.785 27.1975 -0.72 27.3325 ;
        RECT  -3.745 28.0175 -3.68 28.1525 ;
        RECT  -3.61 27.4025 -3.545 27.5375 ;
        RECT  -3.475 27.1975 -3.41 27.3325 ;
        RECT  -2.445 29.41 -2.38 29.545 ;
        RECT  -2.2325 30.385 -2.1675 30.52 ;
        RECT  -3.445 31.85 -3.38 31.985 ;
        RECT  -2.28 30.61 -2.215 30.745 ;
        RECT  -0.1725 26.7875 -0.1075 26.9225 ;
        RECT  -1.5175 27.6075 -1.4525 27.7425 ;
        RECT  -2.8625 26.7875 -2.7975 26.9225 ;
        RECT  -4.2075 27.6075 -4.1425 27.7425 ;
        RECT  0.1075 27.6425 0.2425 27.7075 ;
        LAYER  via1 ;
        RECT  11.0175 19.875 11.0825 19.94 ;
        RECT  11.0175 19.875 11.0825 19.94 ;
        RECT  11.0175 19.875 11.0825 19.94 ;
        RECT  11.0175 19.875 11.0825 19.94 ;
        RECT  11.0175 19.875 11.0825 19.94 ;
        RECT  11.0175 19.875 11.0825 19.94 ;
        RECT  10.3125 19.0575 10.3775 19.1225 ;
        RECT  11.0175 19.0575 11.0825 19.1225 ;
        RECT  11.0175 19.875 11.0825 19.94 ;
        RECT  11.0175 19.875 11.0825 19.94 ;
        RECT  11.0175 19.875 11.0825 19.94 ;
        RECT  11.0175 19.875 11.0825 19.94 ;
        RECT  11.0175 19.875 11.0825 19.94 ;
        RECT  11.0175 19.875 11.0825 19.94 ;
        RECT  11.0175 19.875 11.0825 19.94 ;
        RECT  11.0175 19.875 11.0825 19.94 ;
        RECT  10.5675 19.3825 10.6325 19.4475 ;
        RECT  10.3125 19.875 10.3775 19.94 ;
        RECT  10.3125 19.875 10.3775 19.94 ;
        RECT  10.3125 19.875 10.3775 19.94 ;
        RECT  10.3125 19.875 10.3775 19.94 ;
        RECT  10.3125 19.875 10.3775 19.94 ;
        RECT  10.3125 19.875 10.3775 19.94 ;
        RECT  11.0175 19.875 11.0825 19.94 ;
        RECT  11.0175 19.875 11.0825 19.94 ;
        RECT  11.0175 19.875 11.0825 19.94 ;
        RECT  11.0175 19.875 11.0825 19.94 ;
        RECT  10.7625 19.3825 10.8275 19.4475 ;
        RECT  11.0175 19.0575 11.0825 19.1225 ;
        RECT  11.0175 19.0575 11.0825 19.1225 ;
        RECT  11.0175 19.0575 11.0825 19.1225 ;
        RECT  11.0175 19.875 11.0825 19.94 ;
        RECT  11.0175 19.875 11.0825 19.94 ;
        RECT  11.0175 19.875 11.0825 19.94 ;
        RECT  11.0175 19.875 11.0825 19.94 ;
        RECT  11.0175 19.875 11.0825 19.94 ;
        RECT  11.0175 19.875 11.0825 19.94 ;
        RECT  10.3125 19.0575 10.3775 19.1225 ;
        RECT  11.0175 20.93 11.0825 20.995 ;
        RECT  11.0175 20.93 11.0825 20.995 ;
        RECT  11.0175 20.93 11.0825 20.995 ;
        RECT  11.0175 20.93 11.0825 20.995 ;
        RECT  11.0175 20.93 11.0825 20.995 ;
        RECT  11.0175 20.93 11.0825 20.995 ;
        RECT  10.3125 21.7475 10.3775 21.8125 ;
        RECT  11.0175 21.7475 11.0825 21.8125 ;
        RECT  11.0175 20.93 11.0825 20.995 ;
        RECT  11.0175 20.93 11.0825 20.995 ;
        RECT  11.0175 20.93 11.0825 20.995 ;
        RECT  11.0175 20.93 11.0825 20.995 ;
        RECT  11.0175 20.93 11.0825 20.995 ;
        RECT  11.0175 20.93 11.0825 20.995 ;
        RECT  11.0175 20.93 11.0825 20.995 ;
        RECT  11.0175 20.93 11.0825 20.995 ;
        RECT  10.5675 21.4225 10.6325 21.4875 ;
        RECT  10.3125 20.93 10.3775 20.995 ;
        RECT  10.3125 20.93 10.3775 20.995 ;
        RECT  10.3125 20.93 10.3775 20.995 ;
        RECT  10.3125 20.93 10.3775 20.995 ;
        RECT  10.3125 20.93 10.3775 20.995 ;
        RECT  10.3125 20.93 10.3775 20.995 ;
        RECT  11.0175 20.93 11.0825 20.995 ;
        RECT  11.0175 20.93 11.0825 20.995 ;
        RECT  11.0175 20.93 11.0825 20.995 ;
        RECT  11.0175 20.93 11.0825 20.995 ;
        RECT  10.7625 21.4225 10.8275 21.4875 ;
        RECT  11.0175 21.7475 11.0825 21.8125 ;
        RECT  11.0175 21.7475 11.0825 21.8125 ;
        RECT  11.0175 21.7475 11.0825 21.8125 ;
        RECT  11.0175 20.93 11.0825 20.995 ;
        RECT  11.0175 20.93 11.0825 20.995 ;
        RECT  11.0175 20.93 11.0825 20.995 ;
        RECT  11.0175 20.93 11.0825 20.995 ;
        RECT  11.0175 20.93 11.0825 20.995 ;
        RECT  11.0175 20.93 11.0825 20.995 ;
        RECT  10.3125 21.7475 10.3775 21.8125 ;
        RECT  11.0175 22.565 11.0825 22.63 ;
        RECT  11.0175 22.565 11.0825 22.63 ;
        RECT  11.0175 22.565 11.0825 22.63 ;
        RECT  11.0175 22.565 11.0825 22.63 ;
        RECT  11.0175 22.565 11.0825 22.63 ;
        RECT  11.0175 22.565 11.0825 22.63 ;
        RECT  10.3125 21.7475 10.3775 21.8125 ;
        RECT  11.0175 21.7475 11.0825 21.8125 ;
        RECT  11.0175 22.565 11.0825 22.63 ;
        RECT  11.0175 22.565 11.0825 22.63 ;
        RECT  11.0175 22.565 11.0825 22.63 ;
        RECT  11.0175 22.565 11.0825 22.63 ;
        RECT  11.0175 22.565 11.0825 22.63 ;
        RECT  11.0175 22.565 11.0825 22.63 ;
        RECT  11.0175 22.565 11.0825 22.63 ;
        RECT  11.0175 22.565 11.0825 22.63 ;
        RECT  10.5675 22.0725 10.6325 22.1375 ;
        RECT  10.3125 22.565 10.3775 22.63 ;
        RECT  10.3125 22.565 10.3775 22.63 ;
        RECT  10.3125 22.565 10.3775 22.63 ;
        RECT  10.3125 22.565 10.3775 22.63 ;
        RECT  10.3125 22.565 10.3775 22.63 ;
        RECT  10.3125 22.565 10.3775 22.63 ;
        RECT  11.0175 22.565 11.0825 22.63 ;
        RECT  11.0175 22.565 11.0825 22.63 ;
        RECT  11.0175 22.565 11.0825 22.63 ;
        RECT  11.0175 22.565 11.0825 22.63 ;
        RECT  10.7625 22.0725 10.8275 22.1375 ;
        RECT  11.0175 21.7475 11.0825 21.8125 ;
        RECT  11.0175 21.7475 11.0825 21.8125 ;
        RECT  11.0175 21.7475 11.0825 21.8125 ;
        RECT  11.0175 22.565 11.0825 22.63 ;
        RECT  11.0175 22.565 11.0825 22.63 ;
        RECT  11.0175 22.565 11.0825 22.63 ;
        RECT  11.0175 22.565 11.0825 22.63 ;
        RECT  11.0175 22.565 11.0825 22.63 ;
        RECT  11.0175 22.565 11.0825 22.63 ;
        RECT  10.3125 21.7475 10.3775 21.8125 ;
        RECT  11.0175 23.62 11.0825 23.685 ;
        RECT  11.0175 23.62 11.0825 23.685 ;
        RECT  11.0175 23.62 11.0825 23.685 ;
        RECT  11.0175 23.62 11.0825 23.685 ;
        RECT  11.0175 23.62 11.0825 23.685 ;
        RECT  11.0175 23.62 11.0825 23.685 ;
        RECT  10.3125 24.4375 10.3775 24.5025 ;
        RECT  11.0175 24.4375 11.0825 24.5025 ;
        RECT  11.0175 23.62 11.0825 23.685 ;
        RECT  11.0175 23.62 11.0825 23.685 ;
        RECT  11.0175 23.62 11.0825 23.685 ;
        RECT  11.0175 23.62 11.0825 23.685 ;
        RECT  11.0175 23.62 11.0825 23.685 ;
        RECT  11.0175 23.62 11.0825 23.685 ;
        RECT  11.0175 23.62 11.0825 23.685 ;
        RECT  11.0175 23.62 11.0825 23.685 ;
        RECT  10.5675 24.1125 10.6325 24.1775 ;
        RECT  10.3125 23.62 10.3775 23.685 ;
        RECT  10.3125 23.62 10.3775 23.685 ;
        RECT  10.3125 23.62 10.3775 23.685 ;
        RECT  10.3125 23.62 10.3775 23.685 ;
        RECT  10.3125 23.62 10.3775 23.685 ;
        RECT  10.3125 23.62 10.3775 23.685 ;
        RECT  11.0175 23.62 11.0825 23.685 ;
        RECT  11.0175 23.62 11.0825 23.685 ;
        RECT  11.0175 23.62 11.0825 23.685 ;
        RECT  11.0175 23.62 11.0825 23.685 ;
        RECT  10.7625 24.1125 10.8275 24.1775 ;
        RECT  11.0175 24.4375 11.0825 24.5025 ;
        RECT  11.0175 24.4375 11.0825 24.5025 ;
        RECT  11.0175 24.4375 11.0825 24.5025 ;
        RECT  11.0175 23.62 11.0825 23.685 ;
        RECT  11.0175 23.62 11.0825 23.685 ;
        RECT  11.0175 23.62 11.0825 23.685 ;
        RECT  11.0175 23.62 11.0825 23.685 ;
        RECT  11.0175 23.62 11.0825 23.685 ;
        RECT  11.0175 23.62 11.0825 23.685 ;
        RECT  10.3125 24.4375 10.3775 24.5025 ;
        RECT  11.0175 25.255 11.0825 25.32 ;
        RECT  11.0175 25.255 11.0825 25.32 ;
        RECT  11.0175 25.255 11.0825 25.32 ;
        RECT  11.0175 25.255 11.0825 25.32 ;
        RECT  11.0175 25.255 11.0825 25.32 ;
        RECT  11.0175 25.255 11.0825 25.32 ;
        RECT  10.3125 24.4375 10.3775 24.5025 ;
        RECT  11.0175 24.4375 11.0825 24.5025 ;
        RECT  11.0175 25.255 11.0825 25.32 ;
        RECT  11.0175 25.255 11.0825 25.32 ;
        RECT  11.0175 25.255 11.0825 25.32 ;
        RECT  11.0175 25.255 11.0825 25.32 ;
        RECT  11.0175 25.255 11.0825 25.32 ;
        RECT  11.0175 25.255 11.0825 25.32 ;
        RECT  11.0175 25.255 11.0825 25.32 ;
        RECT  11.0175 25.255 11.0825 25.32 ;
        RECT  10.5675 24.7625 10.6325 24.8275 ;
        RECT  10.3125 25.255 10.3775 25.32 ;
        RECT  10.3125 25.255 10.3775 25.32 ;
        RECT  10.3125 25.255 10.3775 25.32 ;
        RECT  10.3125 25.255 10.3775 25.32 ;
        RECT  10.3125 25.255 10.3775 25.32 ;
        RECT  10.3125 25.255 10.3775 25.32 ;
        RECT  11.0175 25.255 11.0825 25.32 ;
        RECT  11.0175 25.255 11.0825 25.32 ;
        RECT  11.0175 25.255 11.0825 25.32 ;
        RECT  11.0175 25.255 11.0825 25.32 ;
        RECT  10.7625 24.7625 10.8275 24.8275 ;
        RECT  11.0175 24.4375 11.0825 24.5025 ;
        RECT  11.0175 24.4375 11.0825 24.5025 ;
        RECT  11.0175 24.4375 11.0825 24.5025 ;
        RECT  11.0175 25.255 11.0825 25.32 ;
        RECT  11.0175 25.255 11.0825 25.32 ;
        RECT  11.0175 25.255 11.0825 25.32 ;
        RECT  11.0175 25.255 11.0825 25.32 ;
        RECT  11.0175 25.255 11.0825 25.32 ;
        RECT  11.0175 25.255 11.0825 25.32 ;
        RECT  10.3125 24.4375 10.3775 24.5025 ;
        RECT  11.0175 26.31 11.0825 26.375 ;
        RECT  11.0175 26.31 11.0825 26.375 ;
        RECT  11.0175 26.31 11.0825 26.375 ;
        RECT  11.0175 26.31 11.0825 26.375 ;
        RECT  11.0175 26.31 11.0825 26.375 ;
        RECT  11.0175 26.31 11.0825 26.375 ;
        RECT  10.3125 27.1275 10.3775 27.1925 ;
        RECT  11.0175 27.1275 11.0825 27.1925 ;
        RECT  11.0175 26.31 11.0825 26.375 ;
        RECT  11.0175 26.31 11.0825 26.375 ;
        RECT  11.0175 26.31 11.0825 26.375 ;
        RECT  11.0175 26.31 11.0825 26.375 ;
        RECT  11.0175 26.31 11.0825 26.375 ;
        RECT  11.0175 26.31 11.0825 26.375 ;
        RECT  11.0175 26.31 11.0825 26.375 ;
        RECT  11.0175 26.31 11.0825 26.375 ;
        RECT  10.5675 26.8025 10.6325 26.8675 ;
        RECT  10.3125 26.31 10.3775 26.375 ;
        RECT  10.3125 26.31 10.3775 26.375 ;
        RECT  10.3125 26.31 10.3775 26.375 ;
        RECT  10.3125 26.31 10.3775 26.375 ;
        RECT  10.3125 26.31 10.3775 26.375 ;
        RECT  10.3125 26.31 10.3775 26.375 ;
        RECT  11.0175 26.31 11.0825 26.375 ;
        RECT  11.0175 26.31 11.0825 26.375 ;
        RECT  11.0175 26.31 11.0825 26.375 ;
        RECT  11.0175 26.31 11.0825 26.375 ;
        RECT  10.7625 26.8025 10.8275 26.8675 ;
        RECT  11.0175 27.1275 11.0825 27.1925 ;
        RECT  11.0175 27.1275 11.0825 27.1925 ;
        RECT  11.0175 27.1275 11.0825 27.1925 ;
        RECT  11.0175 26.31 11.0825 26.375 ;
        RECT  11.0175 26.31 11.0825 26.375 ;
        RECT  11.0175 26.31 11.0825 26.375 ;
        RECT  11.0175 26.31 11.0825 26.375 ;
        RECT  11.0175 26.31 11.0825 26.375 ;
        RECT  11.0175 26.31 11.0825 26.375 ;
        RECT  10.3125 27.1275 10.3775 27.1925 ;
        RECT  11.0175 27.945 11.0825 28.01 ;
        RECT  11.0175 27.945 11.0825 28.01 ;
        RECT  11.0175 27.945 11.0825 28.01 ;
        RECT  11.0175 27.945 11.0825 28.01 ;
        RECT  11.0175 27.945 11.0825 28.01 ;
        RECT  11.0175 27.945 11.0825 28.01 ;
        RECT  10.3125 27.1275 10.3775 27.1925 ;
        RECT  11.0175 27.1275 11.0825 27.1925 ;
        RECT  11.0175 27.945 11.0825 28.01 ;
        RECT  11.0175 27.945 11.0825 28.01 ;
        RECT  11.0175 27.945 11.0825 28.01 ;
        RECT  11.0175 27.945 11.0825 28.01 ;
        RECT  11.0175 27.945 11.0825 28.01 ;
        RECT  11.0175 27.945 11.0825 28.01 ;
        RECT  11.0175 27.945 11.0825 28.01 ;
        RECT  11.0175 27.945 11.0825 28.01 ;
        RECT  10.5675 27.4525 10.6325 27.5175 ;
        RECT  10.3125 27.945 10.3775 28.01 ;
        RECT  10.3125 27.945 10.3775 28.01 ;
        RECT  10.3125 27.945 10.3775 28.01 ;
        RECT  10.3125 27.945 10.3775 28.01 ;
        RECT  10.3125 27.945 10.3775 28.01 ;
        RECT  10.3125 27.945 10.3775 28.01 ;
        RECT  11.0175 27.945 11.0825 28.01 ;
        RECT  11.0175 27.945 11.0825 28.01 ;
        RECT  11.0175 27.945 11.0825 28.01 ;
        RECT  11.0175 27.945 11.0825 28.01 ;
        RECT  10.7625 27.4525 10.8275 27.5175 ;
        RECT  11.0175 27.1275 11.0825 27.1925 ;
        RECT  11.0175 27.1275 11.0825 27.1925 ;
        RECT  11.0175 27.1275 11.0825 27.1925 ;
        RECT  11.0175 27.945 11.0825 28.01 ;
        RECT  11.0175 27.945 11.0825 28.01 ;
        RECT  11.0175 27.945 11.0825 28.01 ;
        RECT  11.0175 27.945 11.0825 28.01 ;
        RECT  11.0175 27.945 11.0825 28.01 ;
        RECT  11.0175 27.945 11.0825 28.01 ;
        RECT  10.3125 27.1275 10.3775 27.1925 ;
        RECT  11.0175 29.0 11.0825 29.065 ;
        RECT  11.0175 29.0 11.0825 29.065 ;
        RECT  11.0175 29.0 11.0825 29.065 ;
        RECT  11.0175 29.0 11.0825 29.065 ;
        RECT  11.0175 29.0 11.0825 29.065 ;
        RECT  11.0175 29.0 11.0825 29.065 ;
        RECT  10.3125 29.8175 10.3775 29.8825 ;
        RECT  11.0175 29.8175 11.0825 29.8825 ;
        RECT  11.0175 29.0 11.0825 29.065 ;
        RECT  11.0175 29.0 11.0825 29.065 ;
        RECT  11.0175 29.0 11.0825 29.065 ;
        RECT  11.0175 29.0 11.0825 29.065 ;
        RECT  11.0175 29.0 11.0825 29.065 ;
        RECT  11.0175 29.0 11.0825 29.065 ;
        RECT  11.0175 29.0 11.0825 29.065 ;
        RECT  11.0175 29.0 11.0825 29.065 ;
        RECT  10.5675 29.4925 10.6325 29.5575 ;
        RECT  10.3125 29.0 10.3775 29.065 ;
        RECT  10.3125 29.0 10.3775 29.065 ;
        RECT  10.3125 29.0 10.3775 29.065 ;
        RECT  10.3125 29.0 10.3775 29.065 ;
        RECT  10.3125 29.0 10.3775 29.065 ;
        RECT  10.3125 29.0 10.3775 29.065 ;
        RECT  11.0175 29.0 11.0825 29.065 ;
        RECT  11.0175 29.0 11.0825 29.065 ;
        RECT  11.0175 29.0 11.0825 29.065 ;
        RECT  11.0175 29.0 11.0825 29.065 ;
        RECT  10.7625 29.4925 10.8275 29.5575 ;
        RECT  11.0175 29.8175 11.0825 29.8825 ;
        RECT  11.0175 29.8175 11.0825 29.8825 ;
        RECT  11.0175 29.8175 11.0825 29.8825 ;
        RECT  11.0175 29.0 11.0825 29.065 ;
        RECT  11.0175 29.0 11.0825 29.065 ;
        RECT  11.0175 29.0 11.0825 29.065 ;
        RECT  11.0175 29.0 11.0825 29.065 ;
        RECT  11.0175 29.0 11.0825 29.065 ;
        RECT  11.0175 29.0 11.0825 29.065 ;
        RECT  10.3125 29.8175 10.3775 29.8825 ;
        RECT  11.0175 30.635 11.0825 30.7 ;
        RECT  11.0175 30.635 11.0825 30.7 ;
        RECT  11.0175 30.635 11.0825 30.7 ;
        RECT  11.0175 30.635 11.0825 30.7 ;
        RECT  11.0175 30.635 11.0825 30.7 ;
        RECT  11.0175 30.635 11.0825 30.7 ;
        RECT  10.3125 29.8175 10.3775 29.8825 ;
        RECT  11.0175 29.8175 11.0825 29.8825 ;
        RECT  11.0175 30.635 11.0825 30.7 ;
        RECT  11.0175 30.635 11.0825 30.7 ;
        RECT  11.0175 30.635 11.0825 30.7 ;
        RECT  11.0175 30.635 11.0825 30.7 ;
        RECT  11.0175 30.635 11.0825 30.7 ;
        RECT  11.0175 30.635 11.0825 30.7 ;
        RECT  11.0175 30.635 11.0825 30.7 ;
        RECT  11.0175 30.635 11.0825 30.7 ;
        RECT  10.5675 30.1425 10.6325 30.2075 ;
        RECT  10.3125 30.635 10.3775 30.7 ;
        RECT  10.3125 30.635 10.3775 30.7 ;
        RECT  10.3125 30.635 10.3775 30.7 ;
        RECT  10.3125 30.635 10.3775 30.7 ;
        RECT  10.3125 30.635 10.3775 30.7 ;
        RECT  10.3125 30.635 10.3775 30.7 ;
        RECT  11.0175 30.635 11.0825 30.7 ;
        RECT  11.0175 30.635 11.0825 30.7 ;
        RECT  11.0175 30.635 11.0825 30.7 ;
        RECT  11.0175 30.635 11.0825 30.7 ;
        RECT  10.7625 30.1425 10.8275 30.2075 ;
        RECT  11.0175 29.8175 11.0825 29.8825 ;
        RECT  11.0175 29.8175 11.0825 29.8825 ;
        RECT  11.0175 29.8175 11.0825 29.8825 ;
        RECT  11.0175 30.635 11.0825 30.7 ;
        RECT  11.0175 30.635 11.0825 30.7 ;
        RECT  11.0175 30.635 11.0825 30.7 ;
        RECT  11.0175 30.635 11.0825 30.7 ;
        RECT  11.0175 30.635 11.0825 30.7 ;
        RECT  11.0175 30.635 11.0825 30.7 ;
        RECT  10.3125 29.8175 10.3775 29.8825 ;
        RECT  11.0175 31.69 11.0825 31.755 ;
        RECT  11.0175 31.69 11.0825 31.755 ;
        RECT  11.0175 31.69 11.0825 31.755 ;
        RECT  11.0175 31.69 11.0825 31.755 ;
        RECT  11.0175 31.69 11.0825 31.755 ;
        RECT  11.0175 31.69 11.0825 31.755 ;
        RECT  10.3125 32.5075 10.3775 32.5725 ;
        RECT  11.0175 32.5075 11.0825 32.5725 ;
        RECT  11.0175 31.69 11.0825 31.755 ;
        RECT  11.0175 31.69 11.0825 31.755 ;
        RECT  11.0175 31.69 11.0825 31.755 ;
        RECT  11.0175 31.69 11.0825 31.755 ;
        RECT  11.0175 31.69 11.0825 31.755 ;
        RECT  11.0175 31.69 11.0825 31.755 ;
        RECT  11.0175 31.69 11.0825 31.755 ;
        RECT  11.0175 31.69 11.0825 31.755 ;
        RECT  10.5675 32.1825 10.6325 32.2475 ;
        RECT  10.3125 31.69 10.3775 31.755 ;
        RECT  10.3125 31.69 10.3775 31.755 ;
        RECT  10.3125 31.69 10.3775 31.755 ;
        RECT  10.3125 31.69 10.3775 31.755 ;
        RECT  10.3125 31.69 10.3775 31.755 ;
        RECT  10.3125 31.69 10.3775 31.755 ;
        RECT  11.0175 31.69 11.0825 31.755 ;
        RECT  11.0175 31.69 11.0825 31.755 ;
        RECT  11.0175 31.69 11.0825 31.755 ;
        RECT  11.0175 31.69 11.0825 31.755 ;
        RECT  10.7625 32.1825 10.8275 32.2475 ;
        RECT  11.0175 32.5075 11.0825 32.5725 ;
        RECT  11.0175 32.5075 11.0825 32.5725 ;
        RECT  11.0175 32.5075 11.0825 32.5725 ;
        RECT  11.0175 31.69 11.0825 31.755 ;
        RECT  11.0175 31.69 11.0825 31.755 ;
        RECT  11.0175 31.69 11.0825 31.755 ;
        RECT  11.0175 31.69 11.0825 31.755 ;
        RECT  11.0175 31.69 11.0825 31.755 ;
        RECT  11.0175 31.69 11.0825 31.755 ;
        RECT  10.3125 32.5075 10.3775 32.5725 ;
        RECT  11.0175 33.325 11.0825 33.39 ;
        RECT  11.0175 33.325 11.0825 33.39 ;
        RECT  11.0175 33.325 11.0825 33.39 ;
        RECT  11.0175 33.325 11.0825 33.39 ;
        RECT  11.0175 33.325 11.0825 33.39 ;
        RECT  11.0175 33.325 11.0825 33.39 ;
        RECT  10.3125 32.5075 10.3775 32.5725 ;
        RECT  11.0175 32.5075 11.0825 32.5725 ;
        RECT  11.0175 33.325 11.0825 33.39 ;
        RECT  11.0175 33.325 11.0825 33.39 ;
        RECT  11.0175 33.325 11.0825 33.39 ;
        RECT  11.0175 33.325 11.0825 33.39 ;
        RECT  11.0175 33.325 11.0825 33.39 ;
        RECT  11.0175 33.325 11.0825 33.39 ;
        RECT  11.0175 33.325 11.0825 33.39 ;
        RECT  11.0175 33.325 11.0825 33.39 ;
        RECT  10.5675 32.8325 10.6325 32.8975 ;
        RECT  10.3125 33.325 10.3775 33.39 ;
        RECT  10.3125 33.325 10.3775 33.39 ;
        RECT  10.3125 33.325 10.3775 33.39 ;
        RECT  10.3125 33.325 10.3775 33.39 ;
        RECT  10.3125 33.325 10.3775 33.39 ;
        RECT  10.3125 33.325 10.3775 33.39 ;
        RECT  11.0175 33.325 11.0825 33.39 ;
        RECT  11.0175 33.325 11.0825 33.39 ;
        RECT  11.0175 33.325 11.0825 33.39 ;
        RECT  11.0175 33.325 11.0825 33.39 ;
        RECT  10.7625 32.8325 10.8275 32.8975 ;
        RECT  11.0175 32.5075 11.0825 32.5725 ;
        RECT  11.0175 32.5075 11.0825 32.5725 ;
        RECT  11.0175 32.5075 11.0825 32.5725 ;
        RECT  11.0175 33.325 11.0825 33.39 ;
        RECT  11.0175 33.325 11.0825 33.39 ;
        RECT  11.0175 33.325 11.0825 33.39 ;
        RECT  11.0175 33.325 11.0825 33.39 ;
        RECT  11.0175 33.325 11.0825 33.39 ;
        RECT  11.0175 33.325 11.0825 33.39 ;
        RECT  10.3125 32.5075 10.3775 32.5725 ;
        RECT  11.0175 34.38 11.0825 34.445 ;
        RECT  11.0175 34.38 11.0825 34.445 ;
        RECT  11.0175 34.38 11.0825 34.445 ;
        RECT  11.0175 34.38 11.0825 34.445 ;
        RECT  11.0175 34.38 11.0825 34.445 ;
        RECT  11.0175 34.38 11.0825 34.445 ;
        RECT  10.3125 35.1975 10.3775 35.2625 ;
        RECT  11.0175 35.1975 11.0825 35.2625 ;
        RECT  11.0175 34.38 11.0825 34.445 ;
        RECT  11.0175 34.38 11.0825 34.445 ;
        RECT  11.0175 34.38 11.0825 34.445 ;
        RECT  11.0175 34.38 11.0825 34.445 ;
        RECT  11.0175 34.38 11.0825 34.445 ;
        RECT  11.0175 34.38 11.0825 34.445 ;
        RECT  11.0175 34.38 11.0825 34.445 ;
        RECT  11.0175 34.38 11.0825 34.445 ;
        RECT  10.5675 34.8725 10.6325 34.9375 ;
        RECT  10.3125 34.38 10.3775 34.445 ;
        RECT  10.3125 34.38 10.3775 34.445 ;
        RECT  10.3125 34.38 10.3775 34.445 ;
        RECT  10.3125 34.38 10.3775 34.445 ;
        RECT  10.3125 34.38 10.3775 34.445 ;
        RECT  10.3125 34.38 10.3775 34.445 ;
        RECT  11.0175 34.38 11.0825 34.445 ;
        RECT  11.0175 34.38 11.0825 34.445 ;
        RECT  11.0175 34.38 11.0825 34.445 ;
        RECT  11.0175 34.38 11.0825 34.445 ;
        RECT  10.7625 34.8725 10.8275 34.9375 ;
        RECT  11.0175 35.1975 11.0825 35.2625 ;
        RECT  11.0175 35.1975 11.0825 35.2625 ;
        RECT  11.0175 35.1975 11.0825 35.2625 ;
        RECT  11.0175 34.38 11.0825 34.445 ;
        RECT  11.0175 34.38 11.0825 34.445 ;
        RECT  11.0175 34.38 11.0825 34.445 ;
        RECT  11.0175 34.38 11.0825 34.445 ;
        RECT  11.0175 34.38 11.0825 34.445 ;
        RECT  11.0175 34.38 11.0825 34.445 ;
        RECT  10.3125 35.1975 10.3775 35.2625 ;
        RECT  11.0175 36.015 11.0825 36.08 ;
        RECT  11.0175 36.015 11.0825 36.08 ;
        RECT  11.0175 36.015 11.0825 36.08 ;
        RECT  11.0175 36.015 11.0825 36.08 ;
        RECT  11.0175 36.015 11.0825 36.08 ;
        RECT  11.0175 36.015 11.0825 36.08 ;
        RECT  10.3125 35.1975 10.3775 35.2625 ;
        RECT  11.0175 35.1975 11.0825 35.2625 ;
        RECT  11.0175 36.015 11.0825 36.08 ;
        RECT  11.0175 36.015 11.0825 36.08 ;
        RECT  11.0175 36.015 11.0825 36.08 ;
        RECT  11.0175 36.015 11.0825 36.08 ;
        RECT  11.0175 36.015 11.0825 36.08 ;
        RECT  11.0175 36.015 11.0825 36.08 ;
        RECT  11.0175 36.015 11.0825 36.08 ;
        RECT  11.0175 36.015 11.0825 36.08 ;
        RECT  10.5675 35.5225 10.6325 35.5875 ;
        RECT  10.3125 36.015 10.3775 36.08 ;
        RECT  10.3125 36.015 10.3775 36.08 ;
        RECT  10.3125 36.015 10.3775 36.08 ;
        RECT  10.3125 36.015 10.3775 36.08 ;
        RECT  10.3125 36.015 10.3775 36.08 ;
        RECT  10.3125 36.015 10.3775 36.08 ;
        RECT  11.0175 36.015 11.0825 36.08 ;
        RECT  11.0175 36.015 11.0825 36.08 ;
        RECT  11.0175 36.015 11.0825 36.08 ;
        RECT  11.0175 36.015 11.0825 36.08 ;
        RECT  10.7625 35.5225 10.8275 35.5875 ;
        RECT  11.0175 35.1975 11.0825 35.2625 ;
        RECT  11.0175 35.1975 11.0825 35.2625 ;
        RECT  11.0175 35.1975 11.0825 35.2625 ;
        RECT  11.0175 36.015 11.0825 36.08 ;
        RECT  11.0175 36.015 11.0825 36.08 ;
        RECT  11.0175 36.015 11.0825 36.08 ;
        RECT  11.0175 36.015 11.0825 36.08 ;
        RECT  11.0175 36.015 11.0825 36.08 ;
        RECT  11.0175 36.015 11.0825 36.08 ;
        RECT  10.3125 35.1975 10.3775 35.2625 ;
        RECT  11.0175 37.07 11.0825 37.135 ;
        RECT  11.0175 37.07 11.0825 37.135 ;
        RECT  11.0175 37.07 11.0825 37.135 ;
        RECT  11.0175 37.07 11.0825 37.135 ;
        RECT  11.0175 37.07 11.0825 37.135 ;
        RECT  11.0175 37.07 11.0825 37.135 ;
        RECT  10.3125 37.8875 10.3775 37.9525 ;
        RECT  11.0175 37.8875 11.0825 37.9525 ;
        RECT  11.0175 37.07 11.0825 37.135 ;
        RECT  11.0175 37.07 11.0825 37.135 ;
        RECT  11.0175 37.07 11.0825 37.135 ;
        RECT  11.0175 37.07 11.0825 37.135 ;
        RECT  11.0175 37.07 11.0825 37.135 ;
        RECT  11.0175 37.07 11.0825 37.135 ;
        RECT  11.0175 37.07 11.0825 37.135 ;
        RECT  11.0175 37.07 11.0825 37.135 ;
        RECT  10.5675 37.5625 10.6325 37.6275 ;
        RECT  10.3125 37.07 10.3775 37.135 ;
        RECT  10.3125 37.07 10.3775 37.135 ;
        RECT  10.3125 37.07 10.3775 37.135 ;
        RECT  10.3125 37.07 10.3775 37.135 ;
        RECT  10.3125 37.07 10.3775 37.135 ;
        RECT  10.3125 37.07 10.3775 37.135 ;
        RECT  11.0175 37.07 11.0825 37.135 ;
        RECT  11.0175 37.07 11.0825 37.135 ;
        RECT  11.0175 37.07 11.0825 37.135 ;
        RECT  11.0175 37.07 11.0825 37.135 ;
        RECT  10.7625 37.5625 10.8275 37.6275 ;
        RECT  11.0175 37.8875 11.0825 37.9525 ;
        RECT  11.0175 37.8875 11.0825 37.9525 ;
        RECT  11.0175 37.8875 11.0825 37.9525 ;
        RECT  11.0175 37.07 11.0825 37.135 ;
        RECT  11.0175 37.07 11.0825 37.135 ;
        RECT  11.0175 37.07 11.0825 37.135 ;
        RECT  11.0175 37.07 11.0825 37.135 ;
        RECT  11.0175 37.07 11.0825 37.135 ;
        RECT  11.0175 37.07 11.0825 37.135 ;
        RECT  10.3125 37.8875 10.3775 37.9525 ;
        RECT  11.0175 38.705 11.0825 38.77 ;
        RECT  11.0175 38.705 11.0825 38.77 ;
        RECT  11.0175 38.705 11.0825 38.77 ;
        RECT  11.0175 38.705 11.0825 38.77 ;
        RECT  11.0175 38.705 11.0825 38.77 ;
        RECT  11.0175 38.705 11.0825 38.77 ;
        RECT  10.3125 37.8875 10.3775 37.9525 ;
        RECT  11.0175 37.8875 11.0825 37.9525 ;
        RECT  11.0175 38.705 11.0825 38.77 ;
        RECT  11.0175 38.705 11.0825 38.77 ;
        RECT  11.0175 38.705 11.0825 38.77 ;
        RECT  11.0175 38.705 11.0825 38.77 ;
        RECT  11.0175 38.705 11.0825 38.77 ;
        RECT  11.0175 38.705 11.0825 38.77 ;
        RECT  11.0175 38.705 11.0825 38.77 ;
        RECT  11.0175 38.705 11.0825 38.77 ;
        RECT  10.5675 38.2125 10.6325 38.2775 ;
        RECT  10.3125 38.705 10.3775 38.77 ;
        RECT  10.3125 38.705 10.3775 38.77 ;
        RECT  10.3125 38.705 10.3775 38.77 ;
        RECT  10.3125 38.705 10.3775 38.77 ;
        RECT  10.3125 38.705 10.3775 38.77 ;
        RECT  10.3125 38.705 10.3775 38.77 ;
        RECT  11.0175 38.705 11.0825 38.77 ;
        RECT  11.0175 38.705 11.0825 38.77 ;
        RECT  11.0175 38.705 11.0825 38.77 ;
        RECT  11.0175 38.705 11.0825 38.77 ;
        RECT  10.7625 38.2125 10.8275 38.2775 ;
        RECT  11.0175 37.8875 11.0825 37.9525 ;
        RECT  11.0175 37.8875 11.0825 37.9525 ;
        RECT  11.0175 37.8875 11.0825 37.9525 ;
        RECT  11.0175 38.705 11.0825 38.77 ;
        RECT  11.0175 38.705 11.0825 38.77 ;
        RECT  11.0175 38.705 11.0825 38.77 ;
        RECT  11.0175 38.705 11.0825 38.77 ;
        RECT  11.0175 38.705 11.0825 38.77 ;
        RECT  11.0175 38.705 11.0825 38.77 ;
        RECT  10.3125 37.8875 10.3775 37.9525 ;
        RECT  11.0175 39.76 11.0825 39.825 ;
        RECT  11.0175 39.76 11.0825 39.825 ;
        RECT  11.0175 39.76 11.0825 39.825 ;
        RECT  11.0175 39.76 11.0825 39.825 ;
        RECT  11.0175 39.76 11.0825 39.825 ;
        RECT  11.0175 39.76 11.0825 39.825 ;
        RECT  10.3125 40.5775 10.3775 40.6425 ;
        RECT  11.0175 40.5775 11.0825 40.6425 ;
        RECT  11.0175 39.76 11.0825 39.825 ;
        RECT  11.0175 39.76 11.0825 39.825 ;
        RECT  11.0175 39.76 11.0825 39.825 ;
        RECT  11.0175 39.76 11.0825 39.825 ;
        RECT  11.0175 39.76 11.0825 39.825 ;
        RECT  11.0175 39.76 11.0825 39.825 ;
        RECT  11.0175 39.76 11.0825 39.825 ;
        RECT  11.0175 39.76 11.0825 39.825 ;
        RECT  10.5675 40.2525 10.6325 40.3175 ;
        RECT  10.3125 39.76 10.3775 39.825 ;
        RECT  10.3125 39.76 10.3775 39.825 ;
        RECT  10.3125 39.76 10.3775 39.825 ;
        RECT  10.3125 39.76 10.3775 39.825 ;
        RECT  10.3125 39.76 10.3775 39.825 ;
        RECT  10.3125 39.76 10.3775 39.825 ;
        RECT  11.0175 39.76 11.0825 39.825 ;
        RECT  11.0175 39.76 11.0825 39.825 ;
        RECT  11.0175 39.76 11.0825 39.825 ;
        RECT  11.0175 39.76 11.0825 39.825 ;
        RECT  10.7625 40.2525 10.8275 40.3175 ;
        RECT  11.0175 40.5775 11.0825 40.6425 ;
        RECT  11.0175 40.5775 11.0825 40.6425 ;
        RECT  11.0175 40.5775 11.0825 40.6425 ;
        RECT  11.0175 39.76 11.0825 39.825 ;
        RECT  11.0175 39.76 11.0825 39.825 ;
        RECT  11.0175 39.76 11.0825 39.825 ;
        RECT  11.0175 39.76 11.0825 39.825 ;
        RECT  11.0175 39.76 11.0825 39.825 ;
        RECT  11.0175 39.76 11.0825 39.825 ;
        RECT  10.3125 40.5775 10.3775 40.6425 ;
        RECT  11.7225 19.875 11.7875 19.94 ;
        RECT  11.7225 19.875 11.7875 19.94 ;
        RECT  11.7225 19.875 11.7875 19.94 ;
        RECT  11.7225 19.875 11.7875 19.94 ;
        RECT  11.7225 19.875 11.7875 19.94 ;
        RECT  11.7225 19.875 11.7875 19.94 ;
        RECT  11.0175 19.0575 11.0825 19.1225 ;
        RECT  11.7225 19.0575 11.7875 19.1225 ;
        RECT  11.7225 19.875 11.7875 19.94 ;
        RECT  11.7225 19.875 11.7875 19.94 ;
        RECT  11.7225 19.875 11.7875 19.94 ;
        RECT  11.7225 19.875 11.7875 19.94 ;
        RECT  11.7225 19.875 11.7875 19.94 ;
        RECT  11.7225 19.875 11.7875 19.94 ;
        RECT  11.7225 19.875 11.7875 19.94 ;
        RECT  11.7225 19.875 11.7875 19.94 ;
        RECT  11.2725 19.3825 11.3375 19.4475 ;
        RECT  11.0175 19.875 11.0825 19.94 ;
        RECT  11.0175 19.875 11.0825 19.94 ;
        RECT  11.0175 19.875 11.0825 19.94 ;
        RECT  11.0175 19.875 11.0825 19.94 ;
        RECT  11.0175 19.875 11.0825 19.94 ;
        RECT  11.0175 19.875 11.0825 19.94 ;
        RECT  11.7225 19.875 11.7875 19.94 ;
        RECT  11.7225 19.875 11.7875 19.94 ;
        RECT  11.7225 19.875 11.7875 19.94 ;
        RECT  11.7225 19.875 11.7875 19.94 ;
        RECT  11.4675 19.3825 11.5325 19.4475 ;
        RECT  11.7225 19.0575 11.7875 19.1225 ;
        RECT  11.7225 19.0575 11.7875 19.1225 ;
        RECT  11.7225 19.0575 11.7875 19.1225 ;
        RECT  11.7225 19.875 11.7875 19.94 ;
        RECT  11.7225 19.875 11.7875 19.94 ;
        RECT  11.7225 19.875 11.7875 19.94 ;
        RECT  11.7225 19.875 11.7875 19.94 ;
        RECT  11.7225 19.875 11.7875 19.94 ;
        RECT  11.7225 19.875 11.7875 19.94 ;
        RECT  11.0175 19.0575 11.0825 19.1225 ;
        RECT  11.7225 20.93 11.7875 20.995 ;
        RECT  11.7225 20.93 11.7875 20.995 ;
        RECT  11.7225 20.93 11.7875 20.995 ;
        RECT  11.7225 20.93 11.7875 20.995 ;
        RECT  11.7225 20.93 11.7875 20.995 ;
        RECT  11.7225 20.93 11.7875 20.995 ;
        RECT  11.0175 21.7475 11.0825 21.8125 ;
        RECT  11.7225 21.7475 11.7875 21.8125 ;
        RECT  11.7225 20.93 11.7875 20.995 ;
        RECT  11.7225 20.93 11.7875 20.995 ;
        RECT  11.7225 20.93 11.7875 20.995 ;
        RECT  11.7225 20.93 11.7875 20.995 ;
        RECT  11.7225 20.93 11.7875 20.995 ;
        RECT  11.7225 20.93 11.7875 20.995 ;
        RECT  11.7225 20.93 11.7875 20.995 ;
        RECT  11.7225 20.93 11.7875 20.995 ;
        RECT  11.2725 21.4225 11.3375 21.4875 ;
        RECT  11.0175 20.93 11.0825 20.995 ;
        RECT  11.0175 20.93 11.0825 20.995 ;
        RECT  11.0175 20.93 11.0825 20.995 ;
        RECT  11.0175 20.93 11.0825 20.995 ;
        RECT  11.0175 20.93 11.0825 20.995 ;
        RECT  11.0175 20.93 11.0825 20.995 ;
        RECT  11.7225 20.93 11.7875 20.995 ;
        RECT  11.7225 20.93 11.7875 20.995 ;
        RECT  11.7225 20.93 11.7875 20.995 ;
        RECT  11.7225 20.93 11.7875 20.995 ;
        RECT  11.4675 21.4225 11.5325 21.4875 ;
        RECT  11.7225 21.7475 11.7875 21.8125 ;
        RECT  11.7225 21.7475 11.7875 21.8125 ;
        RECT  11.7225 21.7475 11.7875 21.8125 ;
        RECT  11.7225 20.93 11.7875 20.995 ;
        RECT  11.7225 20.93 11.7875 20.995 ;
        RECT  11.7225 20.93 11.7875 20.995 ;
        RECT  11.7225 20.93 11.7875 20.995 ;
        RECT  11.7225 20.93 11.7875 20.995 ;
        RECT  11.7225 20.93 11.7875 20.995 ;
        RECT  11.0175 21.7475 11.0825 21.8125 ;
        RECT  11.7225 22.565 11.7875 22.63 ;
        RECT  11.7225 22.565 11.7875 22.63 ;
        RECT  11.7225 22.565 11.7875 22.63 ;
        RECT  11.7225 22.565 11.7875 22.63 ;
        RECT  11.7225 22.565 11.7875 22.63 ;
        RECT  11.7225 22.565 11.7875 22.63 ;
        RECT  11.0175 21.7475 11.0825 21.8125 ;
        RECT  11.7225 21.7475 11.7875 21.8125 ;
        RECT  11.7225 22.565 11.7875 22.63 ;
        RECT  11.7225 22.565 11.7875 22.63 ;
        RECT  11.7225 22.565 11.7875 22.63 ;
        RECT  11.7225 22.565 11.7875 22.63 ;
        RECT  11.7225 22.565 11.7875 22.63 ;
        RECT  11.7225 22.565 11.7875 22.63 ;
        RECT  11.7225 22.565 11.7875 22.63 ;
        RECT  11.7225 22.565 11.7875 22.63 ;
        RECT  11.2725 22.0725 11.3375 22.1375 ;
        RECT  11.0175 22.565 11.0825 22.63 ;
        RECT  11.0175 22.565 11.0825 22.63 ;
        RECT  11.0175 22.565 11.0825 22.63 ;
        RECT  11.0175 22.565 11.0825 22.63 ;
        RECT  11.0175 22.565 11.0825 22.63 ;
        RECT  11.0175 22.565 11.0825 22.63 ;
        RECT  11.7225 22.565 11.7875 22.63 ;
        RECT  11.7225 22.565 11.7875 22.63 ;
        RECT  11.7225 22.565 11.7875 22.63 ;
        RECT  11.7225 22.565 11.7875 22.63 ;
        RECT  11.4675 22.0725 11.5325 22.1375 ;
        RECT  11.7225 21.7475 11.7875 21.8125 ;
        RECT  11.7225 21.7475 11.7875 21.8125 ;
        RECT  11.7225 21.7475 11.7875 21.8125 ;
        RECT  11.7225 22.565 11.7875 22.63 ;
        RECT  11.7225 22.565 11.7875 22.63 ;
        RECT  11.7225 22.565 11.7875 22.63 ;
        RECT  11.7225 22.565 11.7875 22.63 ;
        RECT  11.7225 22.565 11.7875 22.63 ;
        RECT  11.7225 22.565 11.7875 22.63 ;
        RECT  11.0175 21.7475 11.0825 21.8125 ;
        RECT  11.7225 23.62 11.7875 23.685 ;
        RECT  11.7225 23.62 11.7875 23.685 ;
        RECT  11.7225 23.62 11.7875 23.685 ;
        RECT  11.7225 23.62 11.7875 23.685 ;
        RECT  11.7225 23.62 11.7875 23.685 ;
        RECT  11.7225 23.62 11.7875 23.685 ;
        RECT  11.0175 24.4375 11.0825 24.5025 ;
        RECT  11.7225 24.4375 11.7875 24.5025 ;
        RECT  11.7225 23.62 11.7875 23.685 ;
        RECT  11.7225 23.62 11.7875 23.685 ;
        RECT  11.7225 23.62 11.7875 23.685 ;
        RECT  11.7225 23.62 11.7875 23.685 ;
        RECT  11.7225 23.62 11.7875 23.685 ;
        RECT  11.7225 23.62 11.7875 23.685 ;
        RECT  11.7225 23.62 11.7875 23.685 ;
        RECT  11.7225 23.62 11.7875 23.685 ;
        RECT  11.2725 24.1125 11.3375 24.1775 ;
        RECT  11.0175 23.62 11.0825 23.685 ;
        RECT  11.0175 23.62 11.0825 23.685 ;
        RECT  11.0175 23.62 11.0825 23.685 ;
        RECT  11.0175 23.62 11.0825 23.685 ;
        RECT  11.0175 23.62 11.0825 23.685 ;
        RECT  11.0175 23.62 11.0825 23.685 ;
        RECT  11.7225 23.62 11.7875 23.685 ;
        RECT  11.7225 23.62 11.7875 23.685 ;
        RECT  11.7225 23.62 11.7875 23.685 ;
        RECT  11.7225 23.62 11.7875 23.685 ;
        RECT  11.4675 24.1125 11.5325 24.1775 ;
        RECT  11.7225 24.4375 11.7875 24.5025 ;
        RECT  11.7225 24.4375 11.7875 24.5025 ;
        RECT  11.7225 24.4375 11.7875 24.5025 ;
        RECT  11.7225 23.62 11.7875 23.685 ;
        RECT  11.7225 23.62 11.7875 23.685 ;
        RECT  11.7225 23.62 11.7875 23.685 ;
        RECT  11.7225 23.62 11.7875 23.685 ;
        RECT  11.7225 23.62 11.7875 23.685 ;
        RECT  11.7225 23.62 11.7875 23.685 ;
        RECT  11.0175 24.4375 11.0825 24.5025 ;
        RECT  11.7225 25.255 11.7875 25.32 ;
        RECT  11.7225 25.255 11.7875 25.32 ;
        RECT  11.7225 25.255 11.7875 25.32 ;
        RECT  11.7225 25.255 11.7875 25.32 ;
        RECT  11.7225 25.255 11.7875 25.32 ;
        RECT  11.7225 25.255 11.7875 25.32 ;
        RECT  11.0175 24.4375 11.0825 24.5025 ;
        RECT  11.7225 24.4375 11.7875 24.5025 ;
        RECT  11.7225 25.255 11.7875 25.32 ;
        RECT  11.7225 25.255 11.7875 25.32 ;
        RECT  11.7225 25.255 11.7875 25.32 ;
        RECT  11.7225 25.255 11.7875 25.32 ;
        RECT  11.7225 25.255 11.7875 25.32 ;
        RECT  11.7225 25.255 11.7875 25.32 ;
        RECT  11.7225 25.255 11.7875 25.32 ;
        RECT  11.7225 25.255 11.7875 25.32 ;
        RECT  11.2725 24.7625 11.3375 24.8275 ;
        RECT  11.0175 25.255 11.0825 25.32 ;
        RECT  11.0175 25.255 11.0825 25.32 ;
        RECT  11.0175 25.255 11.0825 25.32 ;
        RECT  11.0175 25.255 11.0825 25.32 ;
        RECT  11.0175 25.255 11.0825 25.32 ;
        RECT  11.0175 25.255 11.0825 25.32 ;
        RECT  11.7225 25.255 11.7875 25.32 ;
        RECT  11.7225 25.255 11.7875 25.32 ;
        RECT  11.7225 25.255 11.7875 25.32 ;
        RECT  11.7225 25.255 11.7875 25.32 ;
        RECT  11.4675 24.7625 11.5325 24.8275 ;
        RECT  11.7225 24.4375 11.7875 24.5025 ;
        RECT  11.7225 24.4375 11.7875 24.5025 ;
        RECT  11.7225 24.4375 11.7875 24.5025 ;
        RECT  11.7225 25.255 11.7875 25.32 ;
        RECT  11.7225 25.255 11.7875 25.32 ;
        RECT  11.7225 25.255 11.7875 25.32 ;
        RECT  11.7225 25.255 11.7875 25.32 ;
        RECT  11.7225 25.255 11.7875 25.32 ;
        RECT  11.7225 25.255 11.7875 25.32 ;
        RECT  11.0175 24.4375 11.0825 24.5025 ;
        RECT  11.7225 26.31 11.7875 26.375 ;
        RECT  11.7225 26.31 11.7875 26.375 ;
        RECT  11.7225 26.31 11.7875 26.375 ;
        RECT  11.7225 26.31 11.7875 26.375 ;
        RECT  11.7225 26.31 11.7875 26.375 ;
        RECT  11.7225 26.31 11.7875 26.375 ;
        RECT  11.0175 27.1275 11.0825 27.1925 ;
        RECT  11.7225 27.1275 11.7875 27.1925 ;
        RECT  11.7225 26.31 11.7875 26.375 ;
        RECT  11.7225 26.31 11.7875 26.375 ;
        RECT  11.7225 26.31 11.7875 26.375 ;
        RECT  11.7225 26.31 11.7875 26.375 ;
        RECT  11.7225 26.31 11.7875 26.375 ;
        RECT  11.7225 26.31 11.7875 26.375 ;
        RECT  11.7225 26.31 11.7875 26.375 ;
        RECT  11.7225 26.31 11.7875 26.375 ;
        RECT  11.2725 26.8025 11.3375 26.8675 ;
        RECT  11.0175 26.31 11.0825 26.375 ;
        RECT  11.0175 26.31 11.0825 26.375 ;
        RECT  11.0175 26.31 11.0825 26.375 ;
        RECT  11.0175 26.31 11.0825 26.375 ;
        RECT  11.0175 26.31 11.0825 26.375 ;
        RECT  11.0175 26.31 11.0825 26.375 ;
        RECT  11.7225 26.31 11.7875 26.375 ;
        RECT  11.7225 26.31 11.7875 26.375 ;
        RECT  11.7225 26.31 11.7875 26.375 ;
        RECT  11.7225 26.31 11.7875 26.375 ;
        RECT  11.4675 26.8025 11.5325 26.8675 ;
        RECT  11.7225 27.1275 11.7875 27.1925 ;
        RECT  11.7225 27.1275 11.7875 27.1925 ;
        RECT  11.7225 27.1275 11.7875 27.1925 ;
        RECT  11.7225 26.31 11.7875 26.375 ;
        RECT  11.7225 26.31 11.7875 26.375 ;
        RECT  11.7225 26.31 11.7875 26.375 ;
        RECT  11.7225 26.31 11.7875 26.375 ;
        RECT  11.7225 26.31 11.7875 26.375 ;
        RECT  11.7225 26.31 11.7875 26.375 ;
        RECT  11.0175 27.1275 11.0825 27.1925 ;
        RECT  11.7225 27.945 11.7875 28.01 ;
        RECT  11.7225 27.945 11.7875 28.01 ;
        RECT  11.7225 27.945 11.7875 28.01 ;
        RECT  11.7225 27.945 11.7875 28.01 ;
        RECT  11.7225 27.945 11.7875 28.01 ;
        RECT  11.7225 27.945 11.7875 28.01 ;
        RECT  11.0175 27.1275 11.0825 27.1925 ;
        RECT  11.7225 27.1275 11.7875 27.1925 ;
        RECT  11.7225 27.945 11.7875 28.01 ;
        RECT  11.7225 27.945 11.7875 28.01 ;
        RECT  11.7225 27.945 11.7875 28.01 ;
        RECT  11.7225 27.945 11.7875 28.01 ;
        RECT  11.7225 27.945 11.7875 28.01 ;
        RECT  11.7225 27.945 11.7875 28.01 ;
        RECT  11.7225 27.945 11.7875 28.01 ;
        RECT  11.7225 27.945 11.7875 28.01 ;
        RECT  11.2725 27.4525 11.3375 27.5175 ;
        RECT  11.0175 27.945 11.0825 28.01 ;
        RECT  11.0175 27.945 11.0825 28.01 ;
        RECT  11.0175 27.945 11.0825 28.01 ;
        RECT  11.0175 27.945 11.0825 28.01 ;
        RECT  11.0175 27.945 11.0825 28.01 ;
        RECT  11.0175 27.945 11.0825 28.01 ;
        RECT  11.7225 27.945 11.7875 28.01 ;
        RECT  11.7225 27.945 11.7875 28.01 ;
        RECT  11.7225 27.945 11.7875 28.01 ;
        RECT  11.7225 27.945 11.7875 28.01 ;
        RECT  11.4675 27.4525 11.5325 27.5175 ;
        RECT  11.7225 27.1275 11.7875 27.1925 ;
        RECT  11.7225 27.1275 11.7875 27.1925 ;
        RECT  11.7225 27.1275 11.7875 27.1925 ;
        RECT  11.7225 27.945 11.7875 28.01 ;
        RECT  11.7225 27.945 11.7875 28.01 ;
        RECT  11.7225 27.945 11.7875 28.01 ;
        RECT  11.7225 27.945 11.7875 28.01 ;
        RECT  11.7225 27.945 11.7875 28.01 ;
        RECT  11.7225 27.945 11.7875 28.01 ;
        RECT  11.0175 27.1275 11.0825 27.1925 ;
        RECT  11.7225 29.0 11.7875 29.065 ;
        RECT  11.7225 29.0 11.7875 29.065 ;
        RECT  11.7225 29.0 11.7875 29.065 ;
        RECT  11.7225 29.0 11.7875 29.065 ;
        RECT  11.7225 29.0 11.7875 29.065 ;
        RECT  11.7225 29.0 11.7875 29.065 ;
        RECT  11.0175 29.8175 11.0825 29.8825 ;
        RECT  11.7225 29.8175 11.7875 29.8825 ;
        RECT  11.7225 29.0 11.7875 29.065 ;
        RECT  11.7225 29.0 11.7875 29.065 ;
        RECT  11.7225 29.0 11.7875 29.065 ;
        RECT  11.7225 29.0 11.7875 29.065 ;
        RECT  11.7225 29.0 11.7875 29.065 ;
        RECT  11.7225 29.0 11.7875 29.065 ;
        RECT  11.7225 29.0 11.7875 29.065 ;
        RECT  11.7225 29.0 11.7875 29.065 ;
        RECT  11.2725 29.4925 11.3375 29.5575 ;
        RECT  11.0175 29.0 11.0825 29.065 ;
        RECT  11.0175 29.0 11.0825 29.065 ;
        RECT  11.0175 29.0 11.0825 29.065 ;
        RECT  11.0175 29.0 11.0825 29.065 ;
        RECT  11.0175 29.0 11.0825 29.065 ;
        RECT  11.0175 29.0 11.0825 29.065 ;
        RECT  11.7225 29.0 11.7875 29.065 ;
        RECT  11.7225 29.0 11.7875 29.065 ;
        RECT  11.7225 29.0 11.7875 29.065 ;
        RECT  11.7225 29.0 11.7875 29.065 ;
        RECT  11.4675 29.4925 11.5325 29.5575 ;
        RECT  11.7225 29.8175 11.7875 29.8825 ;
        RECT  11.7225 29.8175 11.7875 29.8825 ;
        RECT  11.7225 29.8175 11.7875 29.8825 ;
        RECT  11.7225 29.0 11.7875 29.065 ;
        RECT  11.7225 29.0 11.7875 29.065 ;
        RECT  11.7225 29.0 11.7875 29.065 ;
        RECT  11.7225 29.0 11.7875 29.065 ;
        RECT  11.7225 29.0 11.7875 29.065 ;
        RECT  11.7225 29.0 11.7875 29.065 ;
        RECT  11.0175 29.8175 11.0825 29.8825 ;
        RECT  11.7225 30.635 11.7875 30.7 ;
        RECT  11.7225 30.635 11.7875 30.7 ;
        RECT  11.7225 30.635 11.7875 30.7 ;
        RECT  11.7225 30.635 11.7875 30.7 ;
        RECT  11.7225 30.635 11.7875 30.7 ;
        RECT  11.7225 30.635 11.7875 30.7 ;
        RECT  11.0175 29.8175 11.0825 29.8825 ;
        RECT  11.7225 29.8175 11.7875 29.8825 ;
        RECT  11.7225 30.635 11.7875 30.7 ;
        RECT  11.7225 30.635 11.7875 30.7 ;
        RECT  11.7225 30.635 11.7875 30.7 ;
        RECT  11.7225 30.635 11.7875 30.7 ;
        RECT  11.7225 30.635 11.7875 30.7 ;
        RECT  11.7225 30.635 11.7875 30.7 ;
        RECT  11.7225 30.635 11.7875 30.7 ;
        RECT  11.7225 30.635 11.7875 30.7 ;
        RECT  11.2725 30.1425 11.3375 30.2075 ;
        RECT  11.0175 30.635 11.0825 30.7 ;
        RECT  11.0175 30.635 11.0825 30.7 ;
        RECT  11.0175 30.635 11.0825 30.7 ;
        RECT  11.0175 30.635 11.0825 30.7 ;
        RECT  11.0175 30.635 11.0825 30.7 ;
        RECT  11.0175 30.635 11.0825 30.7 ;
        RECT  11.7225 30.635 11.7875 30.7 ;
        RECT  11.7225 30.635 11.7875 30.7 ;
        RECT  11.7225 30.635 11.7875 30.7 ;
        RECT  11.7225 30.635 11.7875 30.7 ;
        RECT  11.4675 30.1425 11.5325 30.2075 ;
        RECT  11.7225 29.8175 11.7875 29.8825 ;
        RECT  11.7225 29.8175 11.7875 29.8825 ;
        RECT  11.7225 29.8175 11.7875 29.8825 ;
        RECT  11.7225 30.635 11.7875 30.7 ;
        RECT  11.7225 30.635 11.7875 30.7 ;
        RECT  11.7225 30.635 11.7875 30.7 ;
        RECT  11.7225 30.635 11.7875 30.7 ;
        RECT  11.7225 30.635 11.7875 30.7 ;
        RECT  11.7225 30.635 11.7875 30.7 ;
        RECT  11.0175 29.8175 11.0825 29.8825 ;
        RECT  11.7225 31.69 11.7875 31.755 ;
        RECT  11.7225 31.69 11.7875 31.755 ;
        RECT  11.7225 31.69 11.7875 31.755 ;
        RECT  11.7225 31.69 11.7875 31.755 ;
        RECT  11.7225 31.69 11.7875 31.755 ;
        RECT  11.7225 31.69 11.7875 31.755 ;
        RECT  11.0175 32.5075 11.0825 32.5725 ;
        RECT  11.7225 32.5075 11.7875 32.5725 ;
        RECT  11.7225 31.69 11.7875 31.755 ;
        RECT  11.7225 31.69 11.7875 31.755 ;
        RECT  11.7225 31.69 11.7875 31.755 ;
        RECT  11.7225 31.69 11.7875 31.755 ;
        RECT  11.7225 31.69 11.7875 31.755 ;
        RECT  11.7225 31.69 11.7875 31.755 ;
        RECT  11.7225 31.69 11.7875 31.755 ;
        RECT  11.7225 31.69 11.7875 31.755 ;
        RECT  11.2725 32.1825 11.3375 32.2475 ;
        RECT  11.0175 31.69 11.0825 31.755 ;
        RECT  11.0175 31.69 11.0825 31.755 ;
        RECT  11.0175 31.69 11.0825 31.755 ;
        RECT  11.0175 31.69 11.0825 31.755 ;
        RECT  11.0175 31.69 11.0825 31.755 ;
        RECT  11.0175 31.69 11.0825 31.755 ;
        RECT  11.7225 31.69 11.7875 31.755 ;
        RECT  11.7225 31.69 11.7875 31.755 ;
        RECT  11.7225 31.69 11.7875 31.755 ;
        RECT  11.7225 31.69 11.7875 31.755 ;
        RECT  11.4675 32.1825 11.5325 32.2475 ;
        RECT  11.7225 32.5075 11.7875 32.5725 ;
        RECT  11.7225 32.5075 11.7875 32.5725 ;
        RECT  11.7225 32.5075 11.7875 32.5725 ;
        RECT  11.7225 31.69 11.7875 31.755 ;
        RECT  11.7225 31.69 11.7875 31.755 ;
        RECT  11.7225 31.69 11.7875 31.755 ;
        RECT  11.7225 31.69 11.7875 31.755 ;
        RECT  11.7225 31.69 11.7875 31.755 ;
        RECT  11.7225 31.69 11.7875 31.755 ;
        RECT  11.0175 32.5075 11.0825 32.5725 ;
        RECT  11.7225 33.325 11.7875 33.39 ;
        RECT  11.7225 33.325 11.7875 33.39 ;
        RECT  11.7225 33.325 11.7875 33.39 ;
        RECT  11.7225 33.325 11.7875 33.39 ;
        RECT  11.7225 33.325 11.7875 33.39 ;
        RECT  11.7225 33.325 11.7875 33.39 ;
        RECT  11.0175 32.5075 11.0825 32.5725 ;
        RECT  11.7225 32.5075 11.7875 32.5725 ;
        RECT  11.7225 33.325 11.7875 33.39 ;
        RECT  11.7225 33.325 11.7875 33.39 ;
        RECT  11.7225 33.325 11.7875 33.39 ;
        RECT  11.7225 33.325 11.7875 33.39 ;
        RECT  11.7225 33.325 11.7875 33.39 ;
        RECT  11.7225 33.325 11.7875 33.39 ;
        RECT  11.7225 33.325 11.7875 33.39 ;
        RECT  11.7225 33.325 11.7875 33.39 ;
        RECT  11.2725 32.8325 11.3375 32.8975 ;
        RECT  11.0175 33.325 11.0825 33.39 ;
        RECT  11.0175 33.325 11.0825 33.39 ;
        RECT  11.0175 33.325 11.0825 33.39 ;
        RECT  11.0175 33.325 11.0825 33.39 ;
        RECT  11.0175 33.325 11.0825 33.39 ;
        RECT  11.0175 33.325 11.0825 33.39 ;
        RECT  11.7225 33.325 11.7875 33.39 ;
        RECT  11.7225 33.325 11.7875 33.39 ;
        RECT  11.7225 33.325 11.7875 33.39 ;
        RECT  11.7225 33.325 11.7875 33.39 ;
        RECT  11.4675 32.8325 11.5325 32.8975 ;
        RECT  11.7225 32.5075 11.7875 32.5725 ;
        RECT  11.7225 32.5075 11.7875 32.5725 ;
        RECT  11.7225 32.5075 11.7875 32.5725 ;
        RECT  11.7225 33.325 11.7875 33.39 ;
        RECT  11.7225 33.325 11.7875 33.39 ;
        RECT  11.7225 33.325 11.7875 33.39 ;
        RECT  11.7225 33.325 11.7875 33.39 ;
        RECT  11.7225 33.325 11.7875 33.39 ;
        RECT  11.7225 33.325 11.7875 33.39 ;
        RECT  11.0175 32.5075 11.0825 32.5725 ;
        RECT  11.7225 34.38 11.7875 34.445 ;
        RECT  11.7225 34.38 11.7875 34.445 ;
        RECT  11.7225 34.38 11.7875 34.445 ;
        RECT  11.7225 34.38 11.7875 34.445 ;
        RECT  11.7225 34.38 11.7875 34.445 ;
        RECT  11.7225 34.38 11.7875 34.445 ;
        RECT  11.0175 35.1975 11.0825 35.2625 ;
        RECT  11.7225 35.1975 11.7875 35.2625 ;
        RECT  11.7225 34.38 11.7875 34.445 ;
        RECT  11.7225 34.38 11.7875 34.445 ;
        RECT  11.7225 34.38 11.7875 34.445 ;
        RECT  11.7225 34.38 11.7875 34.445 ;
        RECT  11.7225 34.38 11.7875 34.445 ;
        RECT  11.7225 34.38 11.7875 34.445 ;
        RECT  11.7225 34.38 11.7875 34.445 ;
        RECT  11.7225 34.38 11.7875 34.445 ;
        RECT  11.2725 34.8725 11.3375 34.9375 ;
        RECT  11.0175 34.38 11.0825 34.445 ;
        RECT  11.0175 34.38 11.0825 34.445 ;
        RECT  11.0175 34.38 11.0825 34.445 ;
        RECT  11.0175 34.38 11.0825 34.445 ;
        RECT  11.0175 34.38 11.0825 34.445 ;
        RECT  11.0175 34.38 11.0825 34.445 ;
        RECT  11.7225 34.38 11.7875 34.445 ;
        RECT  11.7225 34.38 11.7875 34.445 ;
        RECT  11.7225 34.38 11.7875 34.445 ;
        RECT  11.7225 34.38 11.7875 34.445 ;
        RECT  11.4675 34.8725 11.5325 34.9375 ;
        RECT  11.7225 35.1975 11.7875 35.2625 ;
        RECT  11.7225 35.1975 11.7875 35.2625 ;
        RECT  11.7225 35.1975 11.7875 35.2625 ;
        RECT  11.7225 34.38 11.7875 34.445 ;
        RECT  11.7225 34.38 11.7875 34.445 ;
        RECT  11.7225 34.38 11.7875 34.445 ;
        RECT  11.7225 34.38 11.7875 34.445 ;
        RECT  11.7225 34.38 11.7875 34.445 ;
        RECT  11.7225 34.38 11.7875 34.445 ;
        RECT  11.0175 35.1975 11.0825 35.2625 ;
        RECT  11.7225 36.015 11.7875 36.08 ;
        RECT  11.7225 36.015 11.7875 36.08 ;
        RECT  11.7225 36.015 11.7875 36.08 ;
        RECT  11.7225 36.015 11.7875 36.08 ;
        RECT  11.7225 36.015 11.7875 36.08 ;
        RECT  11.7225 36.015 11.7875 36.08 ;
        RECT  11.0175 35.1975 11.0825 35.2625 ;
        RECT  11.7225 35.1975 11.7875 35.2625 ;
        RECT  11.7225 36.015 11.7875 36.08 ;
        RECT  11.7225 36.015 11.7875 36.08 ;
        RECT  11.7225 36.015 11.7875 36.08 ;
        RECT  11.7225 36.015 11.7875 36.08 ;
        RECT  11.7225 36.015 11.7875 36.08 ;
        RECT  11.7225 36.015 11.7875 36.08 ;
        RECT  11.7225 36.015 11.7875 36.08 ;
        RECT  11.7225 36.015 11.7875 36.08 ;
        RECT  11.2725 35.5225 11.3375 35.5875 ;
        RECT  11.0175 36.015 11.0825 36.08 ;
        RECT  11.0175 36.015 11.0825 36.08 ;
        RECT  11.0175 36.015 11.0825 36.08 ;
        RECT  11.0175 36.015 11.0825 36.08 ;
        RECT  11.0175 36.015 11.0825 36.08 ;
        RECT  11.0175 36.015 11.0825 36.08 ;
        RECT  11.7225 36.015 11.7875 36.08 ;
        RECT  11.7225 36.015 11.7875 36.08 ;
        RECT  11.7225 36.015 11.7875 36.08 ;
        RECT  11.7225 36.015 11.7875 36.08 ;
        RECT  11.4675 35.5225 11.5325 35.5875 ;
        RECT  11.7225 35.1975 11.7875 35.2625 ;
        RECT  11.7225 35.1975 11.7875 35.2625 ;
        RECT  11.7225 35.1975 11.7875 35.2625 ;
        RECT  11.7225 36.015 11.7875 36.08 ;
        RECT  11.7225 36.015 11.7875 36.08 ;
        RECT  11.7225 36.015 11.7875 36.08 ;
        RECT  11.7225 36.015 11.7875 36.08 ;
        RECT  11.7225 36.015 11.7875 36.08 ;
        RECT  11.7225 36.015 11.7875 36.08 ;
        RECT  11.0175 35.1975 11.0825 35.2625 ;
        RECT  11.7225 37.07 11.7875 37.135 ;
        RECT  11.7225 37.07 11.7875 37.135 ;
        RECT  11.7225 37.07 11.7875 37.135 ;
        RECT  11.7225 37.07 11.7875 37.135 ;
        RECT  11.7225 37.07 11.7875 37.135 ;
        RECT  11.7225 37.07 11.7875 37.135 ;
        RECT  11.0175 37.8875 11.0825 37.9525 ;
        RECT  11.7225 37.8875 11.7875 37.9525 ;
        RECT  11.7225 37.07 11.7875 37.135 ;
        RECT  11.7225 37.07 11.7875 37.135 ;
        RECT  11.7225 37.07 11.7875 37.135 ;
        RECT  11.7225 37.07 11.7875 37.135 ;
        RECT  11.7225 37.07 11.7875 37.135 ;
        RECT  11.7225 37.07 11.7875 37.135 ;
        RECT  11.7225 37.07 11.7875 37.135 ;
        RECT  11.7225 37.07 11.7875 37.135 ;
        RECT  11.2725 37.5625 11.3375 37.6275 ;
        RECT  11.0175 37.07 11.0825 37.135 ;
        RECT  11.0175 37.07 11.0825 37.135 ;
        RECT  11.0175 37.07 11.0825 37.135 ;
        RECT  11.0175 37.07 11.0825 37.135 ;
        RECT  11.0175 37.07 11.0825 37.135 ;
        RECT  11.0175 37.07 11.0825 37.135 ;
        RECT  11.7225 37.07 11.7875 37.135 ;
        RECT  11.7225 37.07 11.7875 37.135 ;
        RECT  11.7225 37.07 11.7875 37.135 ;
        RECT  11.7225 37.07 11.7875 37.135 ;
        RECT  11.4675 37.5625 11.5325 37.6275 ;
        RECT  11.7225 37.8875 11.7875 37.9525 ;
        RECT  11.7225 37.8875 11.7875 37.9525 ;
        RECT  11.7225 37.8875 11.7875 37.9525 ;
        RECT  11.7225 37.07 11.7875 37.135 ;
        RECT  11.7225 37.07 11.7875 37.135 ;
        RECT  11.7225 37.07 11.7875 37.135 ;
        RECT  11.7225 37.07 11.7875 37.135 ;
        RECT  11.7225 37.07 11.7875 37.135 ;
        RECT  11.7225 37.07 11.7875 37.135 ;
        RECT  11.0175 37.8875 11.0825 37.9525 ;
        RECT  11.7225 38.705 11.7875 38.77 ;
        RECT  11.7225 38.705 11.7875 38.77 ;
        RECT  11.7225 38.705 11.7875 38.77 ;
        RECT  11.7225 38.705 11.7875 38.77 ;
        RECT  11.7225 38.705 11.7875 38.77 ;
        RECT  11.7225 38.705 11.7875 38.77 ;
        RECT  11.0175 37.8875 11.0825 37.9525 ;
        RECT  11.7225 37.8875 11.7875 37.9525 ;
        RECT  11.7225 38.705 11.7875 38.77 ;
        RECT  11.7225 38.705 11.7875 38.77 ;
        RECT  11.7225 38.705 11.7875 38.77 ;
        RECT  11.7225 38.705 11.7875 38.77 ;
        RECT  11.7225 38.705 11.7875 38.77 ;
        RECT  11.7225 38.705 11.7875 38.77 ;
        RECT  11.7225 38.705 11.7875 38.77 ;
        RECT  11.7225 38.705 11.7875 38.77 ;
        RECT  11.2725 38.2125 11.3375 38.2775 ;
        RECT  11.0175 38.705 11.0825 38.77 ;
        RECT  11.0175 38.705 11.0825 38.77 ;
        RECT  11.0175 38.705 11.0825 38.77 ;
        RECT  11.0175 38.705 11.0825 38.77 ;
        RECT  11.0175 38.705 11.0825 38.77 ;
        RECT  11.0175 38.705 11.0825 38.77 ;
        RECT  11.7225 38.705 11.7875 38.77 ;
        RECT  11.7225 38.705 11.7875 38.77 ;
        RECT  11.7225 38.705 11.7875 38.77 ;
        RECT  11.7225 38.705 11.7875 38.77 ;
        RECT  11.4675 38.2125 11.5325 38.2775 ;
        RECT  11.7225 37.8875 11.7875 37.9525 ;
        RECT  11.7225 37.8875 11.7875 37.9525 ;
        RECT  11.7225 37.8875 11.7875 37.9525 ;
        RECT  11.7225 38.705 11.7875 38.77 ;
        RECT  11.7225 38.705 11.7875 38.77 ;
        RECT  11.7225 38.705 11.7875 38.77 ;
        RECT  11.7225 38.705 11.7875 38.77 ;
        RECT  11.7225 38.705 11.7875 38.77 ;
        RECT  11.7225 38.705 11.7875 38.77 ;
        RECT  11.0175 37.8875 11.0825 37.9525 ;
        RECT  11.7225 39.76 11.7875 39.825 ;
        RECT  11.7225 39.76 11.7875 39.825 ;
        RECT  11.7225 39.76 11.7875 39.825 ;
        RECT  11.7225 39.76 11.7875 39.825 ;
        RECT  11.7225 39.76 11.7875 39.825 ;
        RECT  11.7225 39.76 11.7875 39.825 ;
        RECT  11.0175 40.5775 11.0825 40.6425 ;
        RECT  11.7225 40.5775 11.7875 40.6425 ;
        RECT  11.7225 39.76 11.7875 39.825 ;
        RECT  11.7225 39.76 11.7875 39.825 ;
        RECT  11.7225 39.76 11.7875 39.825 ;
        RECT  11.7225 39.76 11.7875 39.825 ;
        RECT  11.7225 39.76 11.7875 39.825 ;
        RECT  11.7225 39.76 11.7875 39.825 ;
        RECT  11.7225 39.76 11.7875 39.825 ;
        RECT  11.7225 39.76 11.7875 39.825 ;
        RECT  11.2725 40.2525 11.3375 40.3175 ;
        RECT  11.0175 39.76 11.0825 39.825 ;
        RECT  11.0175 39.76 11.0825 39.825 ;
        RECT  11.0175 39.76 11.0825 39.825 ;
        RECT  11.0175 39.76 11.0825 39.825 ;
        RECT  11.0175 39.76 11.0825 39.825 ;
        RECT  11.0175 39.76 11.0825 39.825 ;
        RECT  11.7225 39.76 11.7875 39.825 ;
        RECT  11.7225 39.76 11.7875 39.825 ;
        RECT  11.7225 39.76 11.7875 39.825 ;
        RECT  11.7225 39.76 11.7875 39.825 ;
        RECT  11.4675 40.2525 11.5325 40.3175 ;
        RECT  11.7225 40.5775 11.7875 40.6425 ;
        RECT  11.7225 40.5775 11.7875 40.6425 ;
        RECT  11.7225 40.5775 11.7875 40.6425 ;
        RECT  11.7225 39.76 11.7875 39.825 ;
        RECT  11.7225 39.76 11.7875 39.825 ;
        RECT  11.7225 39.76 11.7875 39.825 ;
        RECT  11.7225 39.76 11.7875 39.825 ;
        RECT  11.7225 39.76 11.7875 39.825 ;
        RECT  11.7225 39.76 11.7875 39.825 ;
        RECT  11.0175 40.5775 11.0825 40.6425 ;
        RECT  10.54 41.6425 10.605 41.7075 ;
        RECT  10.92 41.6425 10.985 41.7075 ;
        RECT  10.54 41.1925 10.605 41.2575 ;
        RECT  10.73 41.1925 10.795 41.2575 ;
        RECT  11.245 41.6425 11.31 41.7075 ;
        RECT  11.625 41.6425 11.69 41.7075 ;
        RECT  11.245 41.1925 11.31 41.2575 ;
        RECT  11.435 41.1925 11.5 41.2575 ;
        RECT  10.665 16.38 10.73 16.445 ;
        RECT  10.665 18.5225 10.73 18.5875 ;
        RECT  10.4725 17.68 10.5375 17.745 ;
        RECT  10.855 17.27 10.92 17.335 ;
        RECT  10.3125 14.4875 10.3775 14.5525 ;
        RECT  11.0175 14.4875 11.0825 14.5525 ;
        RECT  10.66 18.7275 10.725 18.7925 ;
        RECT  11.37 16.38 11.435 16.445 ;
        RECT  11.37 18.5225 11.435 18.5875 ;
        RECT  11.1775 17.68 11.2425 17.745 ;
        RECT  11.56 17.27 11.625 17.335 ;
        RECT  11.0175 14.4875 11.0825 14.5525 ;
        RECT  11.7225 14.4875 11.7875 14.5525 ;
        RECT  11.365 18.7275 11.43 18.7925 ;
        RECT  10.5875 10.165 10.6525 10.23 ;
        RECT  11.0175 11.8 11.0825 11.865 ;
        RECT  11.0175 11.23 11.0825 11.295 ;
        RECT  10.3125 11.23 10.3775 11.295 ;
        RECT  10.7325 11.435 10.7975 11.5 ;
        RECT  11.0175 13.7275 11.0825 13.7925 ;
        RECT  10.7325 11.025 10.7975 11.09 ;
        RECT  10.5925 11.025 10.6575 11.09 ;
        RECT  11.0175 11.435 11.0825 11.5 ;
        RECT  10.3125 11.435 10.3775 11.5 ;
        RECT  10.485 10.4275 10.55 10.4925 ;
        RECT  10.5925 13.405 10.6575 13.47 ;
        RECT  10.7625 11.8 10.8275 11.865 ;
        RECT  10.4525 12.715 10.5175 12.78 ;
        RECT  10.5925 11.435 10.6575 11.5 ;
        RECT  10.3125 11.8 10.3775 11.865 ;
        RECT  10.7625 12.315 10.8275 12.38 ;
        RECT  10.4975 13.9375 10.5625 14.0025 ;
        RECT  10.3125 13.7275 10.3775 13.7925 ;
        RECT  11.2925 10.165 11.3575 10.23 ;
        RECT  11.7225 11.8 11.7875 11.865 ;
        RECT  11.7225 11.23 11.7875 11.295 ;
        RECT  11.0175 11.23 11.0825 11.295 ;
        RECT  11.4375 11.435 11.5025 11.5 ;
        RECT  11.7225 13.7275 11.7875 13.7925 ;
        RECT  11.4375 11.025 11.5025 11.09 ;
        RECT  11.2975 11.025 11.3625 11.09 ;
        RECT  11.7225 11.435 11.7875 11.5 ;
        RECT  11.0175 11.435 11.0825 11.5 ;
        RECT  11.19 10.4275 11.255 10.4925 ;
        RECT  11.2975 13.405 11.3625 13.47 ;
        RECT  11.4675 11.8 11.5325 11.865 ;
        RECT  11.1575 12.715 11.2225 12.78 ;
        RECT  11.2975 11.435 11.3625 11.5 ;
        RECT  11.0175 11.8 11.0825 11.865 ;
        RECT  11.4675 12.315 11.5325 12.38 ;
        RECT  11.2025 13.9375 11.2675 14.0025 ;
        RECT  11.0175 13.7275 11.0825 13.7925 ;
        RECT  10.51 9.3275 10.575 9.3925 ;
        RECT  11.0175 4.15 11.0825 4.215 ;
        RECT  10.875 8.2325 10.94 8.2975 ;
        RECT  10.8775 6.625 10.9425 6.69 ;
        RECT  10.8775 5.2275 10.9425 5.2925 ;
        RECT  10.3125 4.01 10.3775 4.075 ;
        RECT  11.0175 7.0875 11.0825 7.1525 ;
        RECT  10.5125 5.8925 10.5775 5.9575 ;
        RECT  10.8775 9.585 10.9425 9.65 ;
        RECT  10.7 9.075 10.765 9.14 ;
        RECT  11.0175 8.6625 11.0825 8.7275 ;
        RECT  11.0175 3.96 11.0825 4.025 ;
        RECT  11.0175 5.7025 11.0825 5.7675 ;
        RECT  10.5125 5.5025 10.5775 5.5675 ;
        RECT  10.7 5.5025 10.765 5.5675 ;
        RECT  10.7 6.115 10.765 6.18 ;
        RECT  10.51 8.4625 10.575 8.5275 ;
        RECT  10.7 8.4625 10.765 8.5275 ;
        RECT  11.525 9.3275 11.59 9.3925 ;
        RECT  11.0175 4.15 11.0825 4.215 ;
        RECT  11.16 8.2325 11.225 8.2975 ;
        RECT  11.1575 6.625 11.2225 6.69 ;
        RECT  11.1575 5.2275 11.2225 5.2925 ;
        RECT  11.7225 4.01 11.7875 4.075 ;
        RECT  11.0175 7.0875 11.0825 7.1525 ;
        RECT  11.5225 5.8925 11.5875 5.9575 ;
        RECT  11.1575 9.585 11.2225 9.65 ;
        RECT  11.335 9.075 11.4 9.14 ;
        RECT  11.0175 8.6625 11.0825 8.7275 ;
        RECT  11.0175 3.96 11.0825 4.025 ;
        RECT  11.0175 5.7025 11.0825 5.7675 ;
        RECT  11.5225 5.5025 11.5875 5.5675 ;
        RECT  11.335 5.5025 11.4 5.5675 ;
        RECT  11.335 6.115 11.4 6.18 ;
        RECT  11.525 8.4625 11.59 8.5275 ;
        RECT  11.335 8.4625 11.4 8.5275 ;
        RECT  10.7975 4.5075 10.8625 4.5725 ;
        RECT  10.6975 5.715 10.7625 5.78 ;
        RECT  10.49 5.9925 10.555 6.0575 ;
        RECT  11.0175 6.1825 11.0825 6.2475 ;
        RECT  10.7975 6.015 10.8625 6.08 ;
        RECT  11.0175 4.1225 11.0825 4.1875 ;
        RECT  10.665 5.375 10.73 5.44 ;
        RECT  10.4525 4.275 10.5175 4.34 ;
        RECT  11.5025 4.5075 11.5675 4.5725 ;
        RECT  11.4025 5.715 11.4675 5.78 ;
        RECT  11.195 5.9925 11.26 6.0575 ;
        RECT  11.7225 6.1825 11.7875 6.2475 ;
        RECT  11.5025 6.015 11.5675 6.08 ;
        RECT  11.7225 4.1225 11.7875 4.1875 ;
        RECT  11.37 5.375 11.435 5.44 ;
        RECT  11.1575 4.275 11.2225 4.34 ;
        RECT  5.47 9.41 5.535 9.475 ;
        RECT  6.855 8.81 6.92 8.875 ;
        RECT  5.195 10.755 5.26 10.82 ;
        RECT  6.58 10.335 6.645 10.4 ;
        RECT  6.855 11.08 6.92 11.145 ;
        RECT  4.92 11.08 4.985 11.145 ;
        RECT  6.58 12.425 6.645 12.49 ;
        RECT  4.645 12.425 4.71 12.49 ;
        RECT  5.47 9.17 5.535 9.235 ;
        RECT  5.195 8.64 5.26 8.705 ;
        RECT  4.92 9.975 4.985 10.04 ;
        RECT  5.195 10.505 5.26 10.57 ;
        RECT  5.47 11.86 5.535 11.925 ;
        RECT  4.645 11.33 4.71 11.395 ;
        RECT  4.92 12.665 4.985 12.73 ;
        RECT  4.645 13.195 4.71 13.26 ;
        RECT  5.47 14.79 5.535 14.855 ;
        RECT  6.855 14.19 6.92 14.255 ;
        RECT  5.195 16.135 5.26 16.2 ;
        RECT  6.58 15.715 6.645 15.78 ;
        RECT  6.855 16.46 6.92 16.525 ;
        RECT  4.92 16.46 4.985 16.525 ;
        RECT  6.58 17.805 6.645 17.87 ;
        RECT  4.645 17.805 4.71 17.87 ;
        RECT  5.47 14.55 5.535 14.615 ;
        RECT  5.195 14.02 5.26 14.085 ;
        RECT  4.92 15.355 4.985 15.42 ;
        RECT  5.195 15.885 5.26 15.95 ;
        RECT  5.47 17.24 5.535 17.305 ;
        RECT  4.645 16.71 4.71 16.775 ;
        RECT  4.92 18.045 4.985 18.11 ;
        RECT  4.645 18.575 4.71 18.64 ;
        RECT  1.73 8.88 1.795 8.945 ;
        RECT  1.905 10.405 1.97 10.47 ;
        RECT  2.08 11.57 2.145 11.635 ;
        RECT  2.255 13.095 2.32 13.16 ;
        RECT  2.43 14.26 2.495 14.325 ;
        RECT  2.605 15.785 2.67 15.85 ;
        RECT  2.78 16.95 2.845 17.015 ;
        RECT  2.955 18.475 3.02 18.54 ;
        RECT  1.73 20.0 1.795 20.065 ;
        RECT  2.43 19.47 2.495 19.535 ;
        RECT  1.73 20.805 1.795 20.87 ;
        RECT  2.605 21.335 2.67 21.4 ;
        RECT  1.73 22.69 1.795 22.755 ;
        RECT  2.78 22.16 2.845 22.225 ;
        RECT  1.73 23.495 1.795 23.56 ;
        RECT  2.955 24.025 3.02 24.09 ;
        RECT  1.905 25.38 1.97 25.445 ;
        RECT  2.43 24.85 2.495 24.915 ;
        RECT  1.905 26.185 1.97 26.25 ;
        RECT  2.605 26.715 2.67 26.78 ;
        RECT  1.905 28.07 1.97 28.135 ;
        RECT  2.78 27.54 2.845 27.605 ;
        RECT  1.905 28.875 1.97 28.94 ;
        RECT  2.955 29.405 3.02 29.47 ;
        RECT  2.08 30.76 2.145 30.825 ;
        RECT  2.43 30.23 2.495 30.295 ;
        RECT  2.08 31.565 2.145 31.63 ;
        RECT  2.605 32.095 2.67 32.16 ;
        RECT  2.08 33.45 2.145 33.515 ;
        RECT  2.78 32.92 2.845 32.985 ;
        RECT  2.08 34.255 2.145 34.32 ;
        RECT  2.955 34.785 3.02 34.85 ;
        RECT  2.255 36.14 2.32 36.205 ;
        RECT  2.43 35.61 2.495 35.675 ;
        RECT  2.255 36.945 2.32 37.01 ;
        RECT  2.605 37.475 2.67 37.54 ;
        RECT  2.255 38.83 2.32 38.895 ;
        RECT  2.78 38.3 2.845 38.365 ;
        RECT  2.255 39.635 2.32 39.7 ;
        RECT  2.955 40.165 3.02 40.23 ;
        RECT  4.6325 19.64 4.6975 19.705 ;
        RECT  4.7725 20.0 4.8375 20.065 ;
        RECT  5.485 20.0 5.55 20.065 ;
        RECT  4.6325 21.165 4.6975 21.23 ;
        RECT  4.7725 20.805 4.8375 20.87 ;
        RECT  5.485 20.805 5.55 20.87 ;
        RECT  4.6325 22.33 4.6975 22.395 ;
        RECT  4.7725 22.69 4.8375 22.755 ;
        RECT  5.485 22.69 5.55 22.755 ;
        RECT  4.6325 23.855 4.6975 23.92 ;
        RECT  4.7725 23.495 4.8375 23.56 ;
        RECT  5.485 23.495 5.55 23.56 ;
        RECT  4.6325 25.02 4.6975 25.085 ;
        RECT  4.7725 25.38 4.8375 25.445 ;
        RECT  5.485 25.38 5.55 25.445 ;
        RECT  4.6325 26.545 4.6975 26.61 ;
        RECT  4.7725 26.185 4.8375 26.25 ;
        RECT  5.485 26.185 5.55 26.25 ;
        RECT  4.6325 27.71 4.6975 27.775 ;
        RECT  4.7725 28.07 4.8375 28.135 ;
        RECT  5.485 28.07 5.55 28.135 ;
        RECT  4.6325 29.235 4.6975 29.3 ;
        RECT  4.7725 28.875 4.8375 28.94 ;
        RECT  5.485 28.875 5.55 28.94 ;
        RECT  4.6325 30.4 4.6975 30.465 ;
        RECT  4.7725 30.76 4.8375 30.825 ;
        RECT  5.485 30.76 5.55 30.825 ;
        RECT  4.6325 31.925 4.6975 31.99 ;
        RECT  4.7725 31.565 4.8375 31.63 ;
        RECT  5.485 31.565 5.55 31.63 ;
        RECT  4.6325 33.09 4.6975 33.155 ;
        RECT  4.7725 33.45 4.8375 33.515 ;
        RECT  5.485 33.45 5.55 33.515 ;
        RECT  4.6325 34.615 4.6975 34.68 ;
        RECT  4.7725 34.255 4.8375 34.32 ;
        RECT  5.485 34.255 5.55 34.32 ;
        RECT  4.6325 35.78 4.6975 35.845 ;
        RECT  4.7725 36.14 4.8375 36.205 ;
        RECT  5.485 36.14 5.55 36.205 ;
        RECT  4.6325 37.305 4.6975 37.37 ;
        RECT  4.7725 36.945 4.8375 37.01 ;
        RECT  5.485 36.945 5.55 37.01 ;
        RECT  4.6325 38.47 4.6975 38.535 ;
        RECT  4.7725 38.83 4.8375 38.895 ;
        RECT  5.485 38.83 5.55 38.895 ;
        RECT  4.6325 39.995 4.6975 40.06 ;
        RECT  4.7725 39.635 4.8375 39.7 ;
        RECT  5.485 39.635 5.55 39.7 ;
        RECT  6.2175 7.69 6.2825 7.755 ;
        RECT  1.04 7.1825 1.105 7.2475 ;
        RECT  5.1225 7.325 5.1875 7.39 ;
        RECT  3.515 7.3225 3.58 7.3875 ;
        RECT  2.1175 7.3225 2.1825 7.3875 ;
        RECT  0.9 7.8875 0.965 7.9525 ;
        RECT  3.9775 7.1825 4.0425 7.2475 ;
        RECT  2.7825 7.6875 2.8475 7.7525 ;
        RECT  6.475 7.3225 6.54 7.3875 ;
        RECT  5.965 7.5 6.03 7.565 ;
        RECT  5.5525 7.1825 5.6175 7.2475 ;
        RECT  0.85 7.1825 0.915 7.2475 ;
        RECT  2.5925 7.1825 2.6575 7.2475 ;
        RECT  2.3925 7.6875 2.4575 7.7525 ;
        RECT  2.3925 7.5 2.4575 7.565 ;
        RECT  3.005 7.5 3.07 7.565 ;
        RECT  5.3525 7.69 5.4175 7.755 ;
        RECT  5.3525 7.5 5.4175 7.565 ;
        RECT  6.2175 6.675 6.2825 6.74 ;
        RECT  1.04 7.1825 1.105 7.2475 ;
        RECT  5.1225 7.04 5.1875 7.105 ;
        RECT  3.515 7.0425 3.58 7.1075 ;
        RECT  2.1175 7.0425 2.1825 7.1075 ;
        RECT  0.9 6.4775 0.965 6.5425 ;
        RECT  3.9775 7.1825 4.0425 7.2475 ;
        RECT  2.7825 6.6775 2.8475 6.7425 ;
        RECT  6.475 7.0425 6.54 7.1075 ;
        RECT  5.965 6.865 6.03 6.93 ;
        RECT  5.5525 7.1825 5.6175 7.2475 ;
        RECT  0.85 7.1825 0.915 7.2475 ;
        RECT  2.5925 7.1825 2.6575 7.2475 ;
        RECT  2.3925 6.6775 2.4575 6.7425 ;
        RECT  2.3925 6.865 2.4575 6.93 ;
        RECT  3.005 6.865 3.07 6.93 ;
        RECT  5.3525 6.675 5.4175 6.74 ;
        RECT  5.3525 6.865 5.4175 6.93 ;
        RECT  6.2175 6.28 6.2825 6.345 ;
        RECT  1.04 5.7725 1.105 5.8375 ;
        RECT  5.1225 5.915 5.1875 5.98 ;
        RECT  3.515 5.9125 3.58 5.9775 ;
        RECT  2.1175 5.9125 2.1825 5.9775 ;
        RECT  0.9 6.4775 0.965 6.5425 ;
        RECT  3.9775 5.7725 4.0425 5.8375 ;
        RECT  2.7825 6.2775 2.8475 6.3425 ;
        RECT  6.475 5.9125 6.54 5.9775 ;
        RECT  5.965 6.09 6.03 6.155 ;
        RECT  5.5525 5.7725 5.6175 5.8375 ;
        RECT  0.85 5.7725 0.915 5.8375 ;
        RECT  2.5925 5.7725 2.6575 5.8375 ;
        RECT  2.3925 6.2775 2.4575 6.3425 ;
        RECT  2.3925 6.09 2.4575 6.155 ;
        RECT  3.005 6.09 3.07 6.155 ;
        RECT  5.3525 6.28 5.4175 6.345 ;
        RECT  5.3525 6.09 5.4175 6.155 ;
        RECT  6.2175 5.265 6.2825 5.33 ;
        RECT  1.04 5.7725 1.105 5.8375 ;
        RECT  5.1225 5.63 5.1875 5.695 ;
        RECT  3.515 5.6325 3.58 5.6975 ;
        RECT  2.1175 5.6325 2.1825 5.6975 ;
        RECT  0.9 5.0675 0.965 5.1325 ;
        RECT  3.9775 5.7725 4.0425 5.8375 ;
        RECT  2.7825 5.2675 2.8475 5.3325 ;
        RECT  6.475 5.6325 6.54 5.6975 ;
        RECT  5.965 5.455 6.03 5.52 ;
        RECT  5.5525 5.7725 5.6175 5.8375 ;
        RECT  0.85 5.7725 0.915 5.8375 ;
        RECT  2.5925 5.7725 2.6575 5.8375 ;
        RECT  2.3925 5.2675 2.4575 5.3325 ;
        RECT  2.3925 5.455 2.4575 5.52 ;
        RECT  3.005 5.455 3.07 5.52 ;
        RECT  5.3525 5.265 5.4175 5.33 ;
        RECT  5.3525 5.455 5.4175 5.52 ;
        RECT  8.2875 19.0575 8.3525 19.1225 ;
        RECT  8.2875 21.7475 8.3525 21.8125 ;
        RECT  8.2875 24.4375 8.3525 24.5025 ;
        RECT  8.2875 27.1275 8.3525 27.1925 ;
        RECT  8.2875 29.8175 8.3525 29.8825 ;
        RECT  8.2875 32.5075 8.3525 32.5725 ;
        RECT  8.2875 35.1975 8.3525 35.2625 ;
        RECT  8.2875 37.8875 8.3525 37.9525 ;
        RECT  8.2875 40.5775 8.3525 40.6425 ;
        RECT  6.82 8.5025 6.885 8.5675 ;
        RECT  7.1975 8.5025 7.2625 8.5675 ;
        RECT  6.545 9.8475 6.61 9.9125 ;
        RECT  7.4025 9.8475 7.4675 9.9125 ;
        RECT  6.82 13.8825 6.885 13.9475 ;
        RECT  7.6075 13.8825 7.6725 13.9475 ;
        RECT  6.545 15.2275 6.61 15.2925 ;
        RECT  7.8125 15.2275 7.8775 15.2925 ;
        RECT  7.025 8.2975 7.09 8.3625 ;
        RECT  7.025 10.9875 7.09 11.0525 ;
        RECT  7.025 13.6775 7.09 13.7425 ;
        RECT  7.025 16.3675 7.09 16.4325 ;
        RECT  6.955 7.535 7.02 7.6 ;
        RECT  7.1975 7.535 7.2625 7.6 ;
        RECT  6.955 6.83 7.02 6.895 ;
        RECT  7.4025 6.83 7.4675 6.895 ;
        RECT  6.955 6.125 7.02 6.19 ;
        RECT  7.6075 6.125 7.6725 6.19 ;
        RECT  6.955 5.42 7.02 5.485 ;
        RECT  7.8125 5.42 7.8775 5.485 ;
        RECT  6.955 7.8875 7.02 7.9525 ;
        RECT  8.2875 7.8875 8.3525 7.9525 ;
        RECT  6.955 7.1825 7.02 7.2475 ;
        RECT  8.2875 7.1825 8.3525 7.2475 ;
        RECT  6.955 6.4775 7.02 6.5425 ;
        RECT  8.2875 6.4775 8.3525 6.5425 ;
        RECT  6.955 5.7725 7.02 5.8375 ;
        RECT  8.2875 5.7725 8.3525 5.8375 ;
        RECT  6.955 5.0675 7.02 5.1325 ;
        RECT  8.2875 5.0675 8.3525 5.1325 ;
        RECT  9.425 3.795 9.49 3.86 ;
        RECT  9.015 1.61 9.08 1.675 ;
        RECT  9.22 3.1575 9.285 3.2225 ;
        RECT  9.425 41.395 9.49 41.46 ;
        RECT  9.63 10.2975 9.695 10.3625 ;
        RECT  9.835 14.3225 9.9 14.3875 ;
        RECT  8.81 8.125 8.875 8.19 ;
        RECT  4.6325 40.7825 4.6975 40.8475 ;
        RECT  8.81 40.815 8.875 40.88 ;
        RECT  8.5025 3.0275 8.5675 3.0925 ;
        RECT  8.5025 14.4525 8.5675 14.5175 ;
        RECT  8.5025 3.955 8.5675 4.02 ;
        RECT  8.5025 11.23 8.5675 11.295 ;
        RECT  -3.845 24.9675 -3.78 25.0325 ;
        RECT  -3.3375 19.79 -3.2725 19.855 ;
        RECT  -3.48 23.8725 -3.415 23.9375 ;
        RECT  -3.4775 22.265 -3.4125 22.33 ;
        RECT  -3.4775 20.8675 -3.4125 20.9325 ;
        RECT  -4.0425 19.65 -3.9775 19.715 ;
        RECT  -3.3375 22.7275 -3.2725 22.7925 ;
        RECT  -3.8425 21.5325 -3.7775 21.5975 ;
        RECT  -3.4775 25.225 -3.4125 25.29 ;
        RECT  -3.655 24.715 -3.59 24.78 ;
        RECT  -3.3375 24.3025 -3.2725 24.3675 ;
        RECT  -3.3375 19.6 -3.2725 19.665 ;
        RECT  -3.3375 21.3425 -3.2725 21.4075 ;
        RECT  -3.8425 21.1425 -3.7775 21.2075 ;
        RECT  -3.655 21.1425 -3.59 21.2075 ;
        RECT  -3.655 21.755 -3.59 21.82 ;
        RECT  -3.845 24.1025 -3.78 24.1675 ;
        RECT  -3.655 24.1025 -3.59 24.1675 ;
        RECT  -2.83 24.9675 -2.765 25.0325 ;
        RECT  -3.3375 19.79 -3.2725 19.855 ;
        RECT  -3.195 23.8725 -3.13 23.9375 ;
        RECT  -3.1975 22.265 -3.1325 22.33 ;
        RECT  -3.1975 20.8675 -3.1325 20.9325 ;
        RECT  -2.6325 19.65 -2.5675 19.715 ;
        RECT  -3.3375 22.7275 -3.2725 22.7925 ;
        RECT  -2.8325 21.5325 -2.7675 21.5975 ;
        RECT  -3.1975 25.225 -3.1325 25.29 ;
        RECT  -3.02 24.715 -2.955 24.78 ;
        RECT  -3.3375 24.3025 -3.2725 24.3675 ;
        RECT  -3.3375 19.6 -3.2725 19.665 ;
        RECT  -3.3375 21.3425 -3.2725 21.4075 ;
        RECT  -2.8325 21.1425 -2.7675 21.2075 ;
        RECT  -3.02 21.1425 -2.955 21.2075 ;
        RECT  -3.02 21.755 -2.955 21.82 ;
        RECT  -2.83 24.1025 -2.765 24.1675 ;
        RECT  -3.02 24.1025 -2.955 24.1675 ;
        RECT  -2.435 24.9675 -2.37 25.0325 ;
        RECT  -1.9275 19.79 -1.8625 19.855 ;
        RECT  -2.07 23.8725 -2.005 23.9375 ;
        RECT  -2.0675 22.265 -2.0025 22.33 ;
        RECT  -2.0675 20.8675 -2.0025 20.9325 ;
        RECT  -2.6325 19.65 -2.5675 19.715 ;
        RECT  -1.9275 22.7275 -1.8625 22.7925 ;
        RECT  -2.4325 21.5325 -2.3675 21.5975 ;
        RECT  -2.0675 25.225 -2.0025 25.29 ;
        RECT  -2.245 24.715 -2.18 24.78 ;
        RECT  -1.9275 24.3025 -1.8625 24.3675 ;
        RECT  -1.9275 19.6 -1.8625 19.665 ;
        RECT  -1.9275 21.3425 -1.8625 21.4075 ;
        RECT  -2.4325 21.1425 -2.3675 21.2075 ;
        RECT  -2.245 21.1425 -2.18 21.2075 ;
        RECT  -2.245 21.755 -2.18 21.82 ;
        RECT  -2.435 24.1025 -2.37 24.1675 ;
        RECT  -2.245 24.1025 -2.18 24.1675 ;
        RECT  -1.3025 28.8825 -1.2375 28.9475 ;
        RECT  -1.3025 29.2625 -1.2375 29.3275 ;
        RECT  -1.9825 29.1075 -1.9175 29.1725 ;
        RECT  -2.515 29.1075 -2.45 29.1725 ;
        RECT  -3.9925 29.4425 -3.9275 29.5075 ;
        RECT  -3.9925 29.8225 -3.9275 29.8875 ;
        RECT  -3.845 25.705 -3.78 25.77 ;
        RECT  -3.69 25.705 -3.625 25.77 ;
        RECT  -2.83 25.705 -2.765 25.77 ;
        RECT  -2.435 25.705 -2.37 25.77 ;
        RECT  -0.7575 34.635 -0.6925 34.7 ;
        RECT  -0.7575 34.075 -0.6925 34.14 ;
        RECT  -2.2775 33.65 -2.2125 33.715 ;
        RECT  -2.2775 34.21 -2.2125 34.275 ;
        RECT  -0.7575 34.3125 -0.6925 34.3775 ;
        RECT  -0.7575 33.7525 -0.6925 33.8175 ;
        RECT  -2.2775 33.9725 -2.2125 34.0375 ;
        RECT  -3.2725 34.6975 -3.2075 34.7625 ;
        RECT  -3.9775 35.1725 -3.9125 35.2375 ;
        RECT  -3.2725 35.1725 -3.2075 35.2375 ;
        RECT  -3.725 34.6925 -3.66 34.7575 ;
        RECT  -3.525 34.6975 -3.46 34.7625 ;
        RECT  -3.9775 34.3675 -3.9125 34.4325 ;
        RECT  -3.2725 34.3675 -3.2075 34.4325 ;
        RECT  -3.9775 33.55 -3.9125 33.615 ;
        RECT  -3.9775 33.55 -3.9125 33.615 ;
        RECT  -3.9775 33.55 -3.9125 33.615 ;
        RECT  -3.9775 33.55 -3.9125 33.615 ;
        RECT  -3.9775 33.55 -3.9125 33.615 ;
        RECT  -3.9775 33.55 -3.9125 33.615 ;
        RECT  -3.2725 34.3675 -3.2075 34.4325 ;
        RECT  -3.9775 34.3675 -3.9125 34.4325 ;
        RECT  -3.9775 33.55 -3.9125 33.615 ;
        RECT  -3.9775 33.55 -3.9125 33.615 ;
        RECT  -3.9775 33.55 -3.9125 33.615 ;
        RECT  -3.9775 33.55 -3.9125 33.615 ;
        RECT  -3.9775 33.55 -3.9125 33.615 ;
        RECT  -3.9775 33.55 -3.9125 33.615 ;
        RECT  -3.9775 33.55 -3.9125 33.615 ;
        RECT  -3.9775 33.55 -3.9125 33.615 ;
        RECT  -3.5275 34.0425 -3.4625 34.1075 ;
        RECT  -3.2725 33.55 -3.2075 33.615 ;
        RECT  -3.2725 33.55 -3.2075 33.615 ;
        RECT  -3.2725 33.55 -3.2075 33.615 ;
        RECT  -3.2725 33.55 -3.2075 33.615 ;
        RECT  -3.2725 33.55 -3.2075 33.615 ;
        RECT  -3.2725 33.55 -3.2075 33.615 ;
        RECT  -3.9775 33.55 -3.9125 33.615 ;
        RECT  -3.9775 33.55 -3.9125 33.615 ;
        RECT  -3.9775 33.55 -3.9125 33.615 ;
        RECT  -3.9775 33.55 -3.9125 33.615 ;
        RECT  -3.7225 34.0425 -3.6575 34.1075 ;
        RECT  -3.9775 34.3675 -3.9125 34.4325 ;
        RECT  -3.9775 34.3675 -3.9125 34.4325 ;
        RECT  -3.9775 34.3675 -3.9125 34.4325 ;
        RECT  -3.9775 33.55 -3.9125 33.615 ;
        RECT  -3.9775 33.55 -3.9125 33.615 ;
        RECT  -3.9775 33.55 -3.9125 33.615 ;
        RECT  -3.9775 33.55 -3.9125 33.615 ;
        RECT  -3.9775 33.55 -3.9125 33.615 ;
        RECT  -3.9775 33.55 -3.9125 33.615 ;
        RECT  -3.2725 34.3675 -3.2075 34.4325 ;
        RECT  -3.9775 32.495 -3.9125 32.56 ;
        RECT  -3.9775 32.495 -3.9125 32.56 ;
        RECT  -3.9775 32.495 -3.9125 32.56 ;
        RECT  -3.9775 32.495 -3.9125 32.56 ;
        RECT  -3.9775 32.495 -3.9125 32.56 ;
        RECT  -3.9775 32.495 -3.9125 32.56 ;
        RECT  -3.2725 31.6775 -3.2075 31.7425 ;
        RECT  -3.9775 31.6775 -3.9125 31.7425 ;
        RECT  -3.9775 32.495 -3.9125 32.56 ;
        RECT  -3.9775 32.495 -3.9125 32.56 ;
        RECT  -3.9775 32.495 -3.9125 32.56 ;
        RECT  -3.9775 32.495 -3.9125 32.56 ;
        RECT  -3.9775 32.495 -3.9125 32.56 ;
        RECT  -3.9775 32.495 -3.9125 32.56 ;
        RECT  -3.9775 32.495 -3.9125 32.56 ;
        RECT  -3.9775 32.495 -3.9125 32.56 ;
        RECT  -3.5275 32.0025 -3.4625 32.0675 ;
        RECT  -3.2725 32.495 -3.2075 32.56 ;
        RECT  -3.2725 32.495 -3.2075 32.56 ;
        RECT  -3.2725 32.495 -3.2075 32.56 ;
        RECT  -3.2725 32.495 -3.2075 32.56 ;
        RECT  -3.2725 32.495 -3.2075 32.56 ;
        RECT  -3.2725 32.495 -3.2075 32.56 ;
        RECT  -3.9775 32.495 -3.9125 32.56 ;
        RECT  -3.9775 32.495 -3.9125 32.56 ;
        RECT  -3.9775 32.495 -3.9125 32.56 ;
        RECT  -3.9775 32.495 -3.9125 32.56 ;
        RECT  -3.7225 32.0025 -3.6575 32.0675 ;
        RECT  -3.9775 31.6775 -3.9125 31.7425 ;
        RECT  -3.9775 31.6775 -3.9125 31.7425 ;
        RECT  -3.9775 31.6775 -3.9125 31.7425 ;
        RECT  -3.9775 32.495 -3.9125 32.56 ;
        RECT  -3.9775 32.495 -3.9125 32.56 ;
        RECT  -3.9775 32.495 -3.9125 32.56 ;
        RECT  -3.9775 32.495 -3.9125 32.56 ;
        RECT  -3.9775 32.495 -3.9125 32.56 ;
        RECT  -3.9775 32.495 -3.9125 32.56 ;
        RECT  -3.2725 31.6775 -3.2075 31.7425 ;
        RECT  -2.8625 34.4075 -2.7975 34.4725 ;
        RECT  -2.8625 36.8175 -2.7975 36.8825 ;
        RECT  -2.8625 34.635 -2.7975 34.7 ;
        RECT  -2.8625 32.26 -2.7975 32.325 ;
        RECT  -2.8625 37.2925 -2.7975 37.3575 ;
        RECT  -3.2725 37.2925 -3.2075 37.3575 ;
        RECT  -3.035 33.1575 -2.97 33.2225 ;
        RECT  -3.035 32.56 -2.97 32.625 ;
        RECT  -3.4575 32.56 -3.3925 32.625 ;
        RECT  -0.755 26.6175 -0.69 26.6825 ;
        RECT  -0.755 23.035 -0.69 23.1 ;
        RECT  -1.7225 19.435 -1.6575 19.5 ;
        RECT  -2.445 26.6175 -2.38 26.6825 ;
        RECT  -2.305 27.0275 -2.24 27.0925 ;
        RECT  -1.92 29.67 -1.855 29.735 ;
        RECT  -2.45 29.67 -2.385 29.735 ;
        RECT  -1.055 28.0525 -0.99 28.1175 ;
        RECT  -0.92 27.8475 -0.855 27.9125 ;
        RECT  -0.785 27.2325 -0.72 27.2975 ;
        RECT  -3.745 28.0525 -3.68 28.1175 ;
        RECT  -3.61 27.4375 -3.545 27.5025 ;
        RECT  -3.475 27.2325 -3.41 27.2975 ;
        RECT  -2.445 29.445 -2.38 29.51 ;
        RECT  -2.2325 30.42 -2.1675 30.485 ;
        RECT  -3.445 31.885 -3.38 31.95 ;
        RECT  -2.28 30.645 -2.215 30.71 ;
        RECT  -0.1725 26.8225 -0.1075 26.8875 ;
        RECT  -1.5175 27.6425 -1.4525 27.7075 ;
        RECT  -2.8625 26.8225 -2.7975 26.8875 ;
        RECT  -4.2075 27.6425 -4.1425 27.7075 ;
        RECT  0.1425 27.6425 0.2075 27.7075 ;
        LAYER  metal2 ;
        RECT  9.8325 30.44 9.9025 30.645 ;
        RECT  9.6275 31.68 9.6975 31.885 ;
        RECT  9.2175 29.24 9.2875 29.445 ;
        RECT  9.0125 30.215 9.0825 30.42 ;
        RECT  9.4225 27.88 9.4925 28.085 ;
        RECT  8.8075 26.445 8.8775 26.65 ;
        RECT  -0.14 27.64 0.175 27.71 ;
        RECT  8.3925 26.65 8.4625 26.855 ;
        RECT  10.6625 0.0 10.7325 0.14 ;
        RECT  11.3675 0.0 11.4375 0.14 ;
        RECT  8.2525 0.0 8.6025 42.02 ;
        RECT  8.8075 0.0 8.8775 42.02 ;
        RECT  9.0125 0.0 9.0825 42.02 ;
        RECT  9.2175 0.0 9.2875 42.02 ;
        RECT  9.4225 0.0 9.4925 42.02 ;
        RECT  9.6275 0.0 9.6975 42.02 ;
        RECT  9.8325 0.0 9.9025 42.02 ;
        RECT  7.2275 4.69 7.2975 19.09 ;
        RECT  7.4325 4.69 7.5025 19.09 ;
        RECT  7.6375 4.69 7.7075 19.09 ;
        RECT  7.8425 4.69 7.9125 19.09 ;
        RECT  10.495 40.71 10.565 41.06 ;
        RECT  10.83 40.71 10.9 41.06 ;
        RECT  11.2 40.71 11.27 41.06 ;
        RECT  11.535 40.71 11.605 41.06 ;
        RECT  10.6625 0.44 10.7325 0.51 ;
        RECT  10.4875 0.44 10.6975 0.51 ;
        RECT  10.6625 0.475 10.7325 0.615 ;
        RECT  11.3675 0.44 11.4375 0.51 ;
        RECT  11.1925 0.44 11.4025 0.51 ;
        RECT  11.3675 0.475 11.4375 0.615 ;
        RECT  4.63 40.61 4.7 40.815 ;
        RECT  10.6625 0.0 10.7325 0.14 ;
        RECT  11.3675 0.0 11.4375 0.14 ;
        RECT  9.6275 0.0 9.6975 42.02 ;
        RECT  9.4225 0.0 9.4925 42.02 ;
        RECT  8.8075 0.0 8.8775 42.02 ;
        RECT  9.8325 0.0 9.9025 42.02 ;
        RECT  9.0125 0.0 9.0825 42.02 ;
        RECT  8.2525 0.0 8.6025 42.02 ;
        RECT  9.2175 0.0 9.2875 42.02 ;
        RECT  10.83 18.99 10.9 40.71 ;
        RECT  11.2 18.99 11.27 40.71 ;
        RECT  11.535 18.99 11.605 40.71 ;
        RECT  10.495 18.99 10.565 40.71 ;
        RECT  10.31 18.99 10.38 40.71 ;
        RECT  11.015 18.99 11.085 40.71 ;
        RECT  11.015 19.84 11.085 19.975 ;
        RECT  11.015 19.84 11.085 19.975 ;
        RECT  11.015 19.84 11.085 19.975 ;
        RECT  11.015 19.84 11.085 19.975 ;
        RECT  11.015 19.84 11.085 19.975 ;
        RECT  11.015 19.84 11.085 19.975 ;
        RECT  10.2775 19.055 10.4125 19.125 ;
        RECT  10.9825 19.055 11.1175 19.125 ;
        RECT  11.015 19.84 11.085 19.975 ;
        RECT  11.015 19.84 11.085 19.975 ;
        RECT  11.015 19.84 11.085 19.975 ;
        RECT  11.015 19.84 11.085 19.975 ;
        RECT  11.015 19.84 11.085 19.975 ;
        RECT  11.015 19.84 11.085 19.975 ;
        RECT  11.015 19.84 11.085 19.975 ;
        RECT  11.015 19.84 11.085 19.975 ;
        RECT  10.565 19.3475 10.635 19.4825 ;
        RECT  10.31 19.84 10.38 19.975 ;
        RECT  10.31 19.84 10.38 19.975 ;
        RECT  10.31 19.84 10.38 19.975 ;
        RECT  10.31 19.84 10.38 19.975 ;
        RECT  10.31 19.84 10.38 19.975 ;
        RECT  10.31 19.84 10.38 19.975 ;
        RECT  11.015 19.84 11.085 19.975 ;
        RECT  11.015 19.84 11.085 19.975 ;
        RECT  11.015 19.84 11.085 19.975 ;
        RECT  11.015 19.84 11.085 19.975 ;
        RECT  10.76 19.3475 10.83 19.4825 ;
        RECT  10.9825 19.055 11.1175 19.125 ;
        RECT  10.9825 19.055 11.1175 19.125 ;
        RECT  10.9825 19.055 11.1175 19.125 ;
        RECT  11.015 19.84 11.085 19.975 ;
        RECT  11.015 19.84 11.085 19.975 ;
        RECT  11.015 19.84 11.085 19.975 ;
        RECT  11.015 19.84 11.085 19.975 ;
        RECT  11.015 19.84 11.085 19.975 ;
        RECT  11.015 19.84 11.085 19.975 ;
        RECT  10.2775 19.055 10.4125 19.125 ;
        RECT  11.015 19.0575 11.085 20.4675 ;
        RECT  10.315 19.06 10.375 19.1175 ;
        RECT  10.5025 19.065 10.5575 19.1175 ;
        RECT  10.8375 19.0575 10.895 19.1175 ;
        RECT  11.02 19.065 11.08 19.1225 ;
        RECT  10.83 18.99 10.9 20.535 ;
        RECT  10.495 18.99 10.565 20.535 ;
        RECT  10.31 18.99 10.38 20.535 ;
        RECT  11.015 18.99 11.085 20.535 ;
        RECT  10.495 18.99 10.565 20.535 ;
        RECT  10.31 18.99 10.38 20.535 ;
        RECT  11.015 18.99 11.085 20.535 ;
        RECT  10.83 18.99 10.9 20.535 ;
        RECT  11.015 20.895 11.085 21.03 ;
        RECT  11.015 20.895 11.085 21.03 ;
        RECT  11.015 20.895 11.085 21.03 ;
        RECT  11.015 20.895 11.085 21.03 ;
        RECT  11.015 20.895 11.085 21.03 ;
        RECT  11.015 20.895 11.085 21.03 ;
        RECT  10.2775 21.745 10.4125 21.815 ;
        RECT  10.9825 21.745 11.1175 21.815 ;
        RECT  11.015 20.895 11.085 21.03 ;
        RECT  11.015 20.895 11.085 21.03 ;
        RECT  11.015 20.895 11.085 21.03 ;
        RECT  11.015 20.895 11.085 21.03 ;
        RECT  11.015 20.895 11.085 21.03 ;
        RECT  11.015 20.895 11.085 21.03 ;
        RECT  11.015 20.895 11.085 21.03 ;
        RECT  11.015 20.895 11.085 21.03 ;
        RECT  10.565 21.3875 10.635 21.5225 ;
        RECT  10.31 20.895 10.38 21.03 ;
        RECT  10.31 20.895 10.38 21.03 ;
        RECT  10.31 20.895 10.38 21.03 ;
        RECT  10.31 20.895 10.38 21.03 ;
        RECT  10.31 20.895 10.38 21.03 ;
        RECT  10.31 20.895 10.38 21.03 ;
        RECT  11.015 20.895 11.085 21.03 ;
        RECT  11.015 20.895 11.085 21.03 ;
        RECT  11.015 20.895 11.085 21.03 ;
        RECT  11.015 20.895 11.085 21.03 ;
        RECT  10.76 21.3875 10.83 21.5225 ;
        RECT  10.9825 21.745 11.1175 21.815 ;
        RECT  10.9825 21.745 11.1175 21.815 ;
        RECT  10.9825 21.745 11.1175 21.815 ;
        RECT  11.015 20.895 11.085 21.03 ;
        RECT  11.015 20.895 11.085 21.03 ;
        RECT  11.015 20.895 11.085 21.03 ;
        RECT  11.015 20.895 11.085 21.03 ;
        RECT  11.015 20.895 11.085 21.03 ;
        RECT  11.015 20.895 11.085 21.03 ;
        RECT  10.2775 21.745 10.4125 21.815 ;
        RECT  11.015 20.4025 11.085 21.8125 ;
        RECT  10.315 21.7525 10.375 21.81 ;
        RECT  10.5025 21.7525 10.5575 21.805 ;
        RECT  10.8375 21.7525 10.895 21.8125 ;
        RECT  11.02 21.7475 11.08 21.805 ;
        RECT  10.83 20.335 10.9 21.88 ;
        RECT  10.495 20.335 10.565 21.88 ;
        RECT  10.31 20.335 10.38 21.88 ;
        RECT  11.015 20.335 11.085 21.88 ;
        RECT  10.495 20.335 10.565 21.88 ;
        RECT  10.31 20.335 10.38 21.88 ;
        RECT  11.015 20.335 11.085 21.88 ;
        RECT  10.83 20.335 10.9 21.88 ;
        RECT  11.015 22.53 11.085 22.665 ;
        RECT  11.015 22.53 11.085 22.665 ;
        RECT  11.015 22.53 11.085 22.665 ;
        RECT  11.015 22.53 11.085 22.665 ;
        RECT  11.015 22.53 11.085 22.665 ;
        RECT  11.015 22.53 11.085 22.665 ;
        RECT  10.2775 21.745 10.4125 21.815 ;
        RECT  10.9825 21.745 11.1175 21.815 ;
        RECT  11.015 22.53 11.085 22.665 ;
        RECT  11.015 22.53 11.085 22.665 ;
        RECT  11.015 22.53 11.085 22.665 ;
        RECT  11.015 22.53 11.085 22.665 ;
        RECT  11.015 22.53 11.085 22.665 ;
        RECT  11.015 22.53 11.085 22.665 ;
        RECT  11.015 22.53 11.085 22.665 ;
        RECT  11.015 22.53 11.085 22.665 ;
        RECT  10.565 22.0375 10.635 22.1725 ;
        RECT  10.31 22.53 10.38 22.665 ;
        RECT  10.31 22.53 10.38 22.665 ;
        RECT  10.31 22.53 10.38 22.665 ;
        RECT  10.31 22.53 10.38 22.665 ;
        RECT  10.31 22.53 10.38 22.665 ;
        RECT  10.31 22.53 10.38 22.665 ;
        RECT  11.015 22.53 11.085 22.665 ;
        RECT  11.015 22.53 11.085 22.665 ;
        RECT  11.015 22.53 11.085 22.665 ;
        RECT  11.015 22.53 11.085 22.665 ;
        RECT  10.76 22.0375 10.83 22.1725 ;
        RECT  10.9825 21.745 11.1175 21.815 ;
        RECT  10.9825 21.745 11.1175 21.815 ;
        RECT  10.9825 21.745 11.1175 21.815 ;
        RECT  11.015 22.53 11.085 22.665 ;
        RECT  11.015 22.53 11.085 22.665 ;
        RECT  11.015 22.53 11.085 22.665 ;
        RECT  11.015 22.53 11.085 22.665 ;
        RECT  11.015 22.53 11.085 22.665 ;
        RECT  11.015 22.53 11.085 22.665 ;
        RECT  10.2775 21.745 10.4125 21.815 ;
        RECT  11.015 21.7475 11.085 23.1575 ;
        RECT  10.315 21.75 10.375 21.8075 ;
        RECT  10.5025 21.755 10.5575 21.8075 ;
        RECT  10.8375 21.7475 10.895 21.8075 ;
        RECT  11.02 21.755 11.08 21.8125 ;
        RECT  10.83 21.68 10.9 23.225 ;
        RECT  10.495 21.68 10.565 23.225 ;
        RECT  10.31 21.68 10.38 23.225 ;
        RECT  11.015 21.68 11.085 23.225 ;
        RECT  10.495 21.68 10.565 23.225 ;
        RECT  10.31 21.68 10.38 23.225 ;
        RECT  11.015 21.68 11.085 23.225 ;
        RECT  10.83 21.68 10.9 23.225 ;
        RECT  11.015 23.585 11.085 23.72 ;
        RECT  11.015 23.585 11.085 23.72 ;
        RECT  11.015 23.585 11.085 23.72 ;
        RECT  11.015 23.585 11.085 23.72 ;
        RECT  11.015 23.585 11.085 23.72 ;
        RECT  11.015 23.585 11.085 23.72 ;
        RECT  10.2775 24.435 10.4125 24.505 ;
        RECT  10.9825 24.435 11.1175 24.505 ;
        RECT  11.015 23.585 11.085 23.72 ;
        RECT  11.015 23.585 11.085 23.72 ;
        RECT  11.015 23.585 11.085 23.72 ;
        RECT  11.015 23.585 11.085 23.72 ;
        RECT  11.015 23.585 11.085 23.72 ;
        RECT  11.015 23.585 11.085 23.72 ;
        RECT  11.015 23.585 11.085 23.72 ;
        RECT  11.015 23.585 11.085 23.72 ;
        RECT  10.565 24.0775 10.635 24.2125 ;
        RECT  10.31 23.585 10.38 23.72 ;
        RECT  10.31 23.585 10.38 23.72 ;
        RECT  10.31 23.585 10.38 23.72 ;
        RECT  10.31 23.585 10.38 23.72 ;
        RECT  10.31 23.585 10.38 23.72 ;
        RECT  10.31 23.585 10.38 23.72 ;
        RECT  11.015 23.585 11.085 23.72 ;
        RECT  11.015 23.585 11.085 23.72 ;
        RECT  11.015 23.585 11.085 23.72 ;
        RECT  11.015 23.585 11.085 23.72 ;
        RECT  10.76 24.0775 10.83 24.2125 ;
        RECT  10.9825 24.435 11.1175 24.505 ;
        RECT  10.9825 24.435 11.1175 24.505 ;
        RECT  10.9825 24.435 11.1175 24.505 ;
        RECT  11.015 23.585 11.085 23.72 ;
        RECT  11.015 23.585 11.085 23.72 ;
        RECT  11.015 23.585 11.085 23.72 ;
        RECT  11.015 23.585 11.085 23.72 ;
        RECT  11.015 23.585 11.085 23.72 ;
        RECT  11.015 23.585 11.085 23.72 ;
        RECT  10.2775 24.435 10.4125 24.505 ;
        RECT  11.015 23.0925 11.085 24.5025 ;
        RECT  10.315 24.4425 10.375 24.5 ;
        RECT  10.5025 24.4425 10.5575 24.495 ;
        RECT  10.8375 24.4425 10.895 24.5025 ;
        RECT  11.02 24.4375 11.08 24.495 ;
        RECT  10.83 23.025 10.9 24.57 ;
        RECT  10.495 23.025 10.565 24.57 ;
        RECT  10.31 23.025 10.38 24.57 ;
        RECT  11.015 23.025 11.085 24.57 ;
        RECT  10.495 23.025 10.565 24.57 ;
        RECT  10.31 23.025 10.38 24.57 ;
        RECT  11.015 23.025 11.085 24.57 ;
        RECT  10.83 23.025 10.9 24.57 ;
        RECT  11.015 25.22 11.085 25.355 ;
        RECT  11.015 25.22 11.085 25.355 ;
        RECT  11.015 25.22 11.085 25.355 ;
        RECT  11.015 25.22 11.085 25.355 ;
        RECT  11.015 25.22 11.085 25.355 ;
        RECT  11.015 25.22 11.085 25.355 ;
        RECT  10.2775 24.435 10.4125 24.505 ;
        RECT  10.9825 24.435 11.1175 24.505 ;
        RECT  11.015 25.22 11.085 25.355 ;
        RECT  11.015 25.22 11.085 25.355 ;
        RECT  11.015 25.22 11.085 25.355 ;
        RECT  11.015 25.22 11.085 25.355 ;
        RECT  11.015 25.22 11.085 25.355 ;
        RECT  11.015 25.22 11.085 25.355 ;
        RECT  11.015 25.22 11.085 25.355 ;
        RECT  11.015 25.22 11.085 25.355 ;
        RECT  10.565 24.7275 10.635 24.8625 ;
        RECT  10.31 25.22 10.38 25.355 ;
        RECT  10.31 25.22 10.38 25.355 ;
        RECT  10.31 25.22 10.38 25.355 ;
        RECT  10.31 25.22 10.38 25.355 ;
        RECT  10.31 25.22 10.38 25.355 ;
        RECT  10.31 25.22 10.38 25.355 ;
        RECT  11.015 25.22 11.085 25.355 ;
        RECT  11.015 25.22 11.085 25.355 ;
        RECT  11.015 25.22 11.085 25.355 ;
        RECT  11.015 25.22 11.085 25.355 ;
        RECT  10.76 24.7275 10.83 24.8625 ;
        RECT  10.9825 24.435 11.1175 24.505 ;
        RECT  10.9825 24.435 11.1175 24.505 ;
        RECT  10.9825 24.435 11.1175 24.505 ;
        RECT  11.015 25.22 11.085 25.355 ;
        RECT  11.015 25.22 11.085 25.355 ;
        RECT  11.015 25.22 11.085 25.355 ;
        RECT  11.015 25.22 11.085 25.355 ;
        RECT  11.015 25.22 11.085 25.355 ;
        RECT  11.015 25.22 11.085 25.355 ;
        RECT  10.2775 24.435 10.4125 24.505 ;
        RECT  11.015 24.4375 11.085 25.8475 ;
        RECT  10.315 24.44 10.375 24.4975 ;
        RECT  10.5025 24.445 10.5575 24.4975 ;
        RECT  10.8375 24.4375 10.895 24.4975 ;
        RECT  11.02 24.445 11.08 24.5025 ;
        RECT  10.83 24.37 10.9 25.915 ;
        RECT  10.495 24.37 10.565 25.915 ;
        RECT  10.31 24.37 10.38 25.915 ;
        RECT  11.015 24.37 11.085 25.915 ;
        RECT  10.495 24.37 10.565 25.915 ;
        RECT  10.31 24.37 10.38 25.915 ;
        RECT  11.015 24.37 11.085 25.915 ;
        RECT  10.83 24.37 10.9 25.915 ;
        RECT  11.015 26.275 11.085 26.41 ;
        RECT  11.015 26.275 11.085 26.41 ;
        RECT  11.015 26.275 11.085 26.41 ;
        RECT  11.015 26.275 11.085 26.41 ;
        RECT  11.015 26.275 11.085 26.41 ;
        RECT  11.015 26.275 11.085 26.41 ;
        RECT  10.2775 27.125 10.4125 27.195 ;
        RECT  10.9825 27.125 11.1175 27.195 ;
        RECT  11.015 26.275 11.085 26.41 ;
        RECT  11.015 26.275 11.085 26.41 ;
        RECT  11.015 26.275 11.085 26.41 ;
        RECT  11.015 26.275 11.085 26.41 ;
        RECT  11.015 26.275 11.085 26.41 ;
        RECT  11.015 26.275 11.085 26.41 ;
        RECT  11.015 26.275 11.085 26.41 ;
        RECT  11.015 26.275 11.085 26.41 ;
        RECT  10.565 26.7675 10.635 26.9025 ;
        RECT  10.31 26.275 10.38 26.41 ;
        RECT  10.31 26.275 10.38 26.41 ;
        RECT  10.31 26.275 10.38 26.41 ;
        RECT  10.31 26.275 10.38 26.41 ;
        RECT  10.31 26.275 10.38 26.41 ;
        RECT  10.31 26.275 10.38 26.41 ;
        RECT  11.015 26.275 11.085 26.41 ;
        RECT  11.015 26.275 11.085 26.41 ;
        RECT  11.015 26.275 11.085 26.41 ;
        RECT  11.015 26.275 11.085 26.41 ;
        RECT  10.76 26.7675 10.83 26.9025 ;
        RECT  10.9825 27.125 11.1175 27.195 ;
        RECT  10.9825 27.125 11.1175 27.195 ;
        RECT  10.9825 27.125 11.1175 27.195 ;
        RECT  11.015 26.275 11.085 26.41 ;
        RECT  11.015 26.275 11.085 26.41 ;
        RECT  11.015 26.275 11.085 26.41 ;
        RECT  11.015 26.275 11.085 26.41 ;
        RECT  11.015 26.275 11.085 26.41 ;
        RECT  11.015 26.275 11.085 26.41 ;
        RECT  10.2775 27.125 10.4125 27.195 ;
        RECT  11.015 25.7825 11.085 27.1925 ;
        RECT  10.315 27.1325 10.375 27.19 ;
        RECT  10.5025 27.1325 10.5575 27.185 ;
        RECT  10.8375 27.1325 10.895 27.1925 ;
        RECT  11.02 27.1275 11.08 27.185 ;
        RECT  10.83 25.715 10.9 27.26 ;
        RECT  10.495 25.715 10.565 27.26 ;
        RECT  10.31 25.715 10.38 27.26 ;
        RECT  11.015 25.715 11.085 27.26 ;
        RECT  10.495 25.715 10.565 27.26 ;
        RECT  10.31 25.715 10.38 27.26 ;
        RECT  11.015 25.715 11.085 27.26 ;
        RECT  10.83 25.715 10.9 27.26 ;
        RECT  11.015 27.91 11.085 28.045 ;
        RECT  11.015 27.91 11.085 28.045 ;
        RECT  11.015 27.91 11.085 28.045 ;
        RECT  11.015 27.91 11.085 28.045 ;
        RECT  11.015 27.91 11.085 28.045 ;
        RECT  11.015 27.91 11.085 28.045 ;
        RECT  10.2775 27.125 10.4125 27.195 ;
        RECT  10.9825 27.125 11.1175 27.195 ;
        RECT  11.015 27.91 11.085 28.045 ;
        RECT  11.015 27.91 11.085 28.045 ;
        RECT  11.015 27.91 11.085 28.045 ;
        RECT  11.015 27.91 11.085 28.045 ;
        RECT  11.015 27.91 11.085 28.045 ;
        RECT  11.015 27.91 11.085 28.045 ;
        RECT  11.015 27.91 11.085 28.045 ;
        RECT  11.015 27.91 11.085 28.045 ;
        RECT  10.565 27.4175 10.635 27.5525 ;
        RECT  10.31 27.91 10.38 28.045 ;
        RECT  10.31 27.91 10.38 28.045 ;
        RECT  10.31 27.91 10.38 28.045 ;
        RECT  10.31 27.91 10.38 28.045 ;
        RECT  10.31 27.91 10.38 28.045 ;
        RECT  10.31 27.91 10.38 28.045 ;
        RECT  11.015 27.91 11.085 28.045 ;
        RECT  11.015 27.91 11.085 28.045 ;
        RECT  11.015 27.91 11.085 28.045 ;
        RECT  11.015 27.91 11.085 28.045 ;
        RECT  10.76 27.4175 10.83 27.5525 ;
        RECT  10.9825 27.125 11.1175 27.195 ;
        RECT  10.9825 27.125 11.1175 27.195 ;
        RECT  10.9825 27.125 11.1175 27.195 ;
        RECT  11.015 27.91 11.085 28.045 ;
        RECT  11.015 27.91 11.085 28.045 ;
        RECT  11.015 27.91 11.085 28.045 ;
        RECT  11.015 27.91 11.085 28.045 ;
        RECT  11.015 27.91 11.085 28.045 ;
        RECT  11.015 27.91 11.085 28.045 ;
        RECT  10.2775 27.125 10.4125 27.195 ;
        RECT  11.015 27.1275 11.085 28.5375 ;
        RECT  10.315 27.13 10.375 27.1875 ;
        RECT  10.5025 27.135 10.5575 27.1875 ;
        RECT  10.8375 27.1275 10.895 27.1875 ;
        RECT  11.02 27.135 11.08 27.1925 ;
        RECT  10.83 27.06 10.9 28.605 ;
        RECT  10.495 27.06 10.565 28.605 ;
        RECT  10.31 27.06 10.38 28.605 ;
        RECT  11.015 27.06 11.085 28.605 ;
        RECT  10.495 27.06 10.565 28.605 ;
        RECT  10.31 27.06 10.38 28.605 ;
        RECT  11.015 27.06 11.085 28.605 ;
        RECT  10.83 27.06 10.9 28.605 ;
        RECT  11.015 28.965 11.085 29.1 ;
        RECT  11.015 28.965 11.085 29.1 ;
        RECT  11.015 28.965 11.085 29.1 ;
        RECT  11.015 28.965 11.085 29.1 ;
        RECT  11.015 28.965 11.085 29.1 ;
        RECT  11.015 28.965 11.085 29.1 ;
        RECT  10.2775 29.815 10.4125 29.885 ;
        RECT  10.9825 29.815 11.1175 29.885 ;
        RECT  11.015 28.965 11.085 29.1 ;
        RECT  11.015 28.965 11.085 29.1 ;
        RECT  11.015 28.965 11.085 29.1 ;
        RECT  11.015 28.965 11.085 29.1 ;
        RECT  11.015 28.965 11.085 29.1 ;
        RECT  11.015 28.965 11.085 29.1 ;
        RECT  11.015 28.965 11.085 29.1 ;
        RECT  11.015 28.965 11.085 29.1 ;
        RECT  10.565 29.4575 10.635 29.5925 ;
        RECT  10.31 28.965 10.38 29.1 ;
        RECT  10.31 28.965 10.38 29.1 ;
        RECT  10.31 28.965 10.38 29.1 ;
        RECT  10.31 28.965 10.38 29.1 ;
        RECT  10.31 28.965 10.38 29.1 ;
        RECT  10.31 28.965 10.38 29.1 ;
        RECT  11.015 28.965 11.085 29.1 ;
        RECT  11.015 28.965 11.085 29.1 ;
        RECT  11.015 28.965 11.085 29.1 ;
        RECT  11.015 28.965 11.085 29.1 ;
        RECT  10.76 29.4575 10.83 29.5925 ;
        RECT  10.9825 29.815 11.1175 29.885 ;
        RECT  10.9825 29.815 11.1175 29.885 ;
        RECT  10.9825 29.815 11.1175 29.885 ;
        RECT  11.015 28.965 11.085 29.1 ;
        RECT  11.015 28.965 11.085 29.1 ;
        RECT  11.015 28.965 11.085 29.1 ;
        RECT  11.015 28.965 11.085 29.1 ;
        RECT  11.015 28.965 11.085 29.1 ;
        RECT  11.015 28.965 11.085 29.1 ;
        RECT  10.2775 29.815 10.4125 29.885 ;
        RECT  11.015 28.4725 11.085 29.8825 ;
        RECT  10.315 29.8225 10.375 29.88 ;
        RECT  10.5025 29.8225 10.5575 29.875 ;
        RECT  10.8375 29.8225 10.895 29.8825 ;
        RECT  11.02 29.8175 11.08 29.875 ;
        RECT  10.83 28.405 10.9 29.95 ;
        RECT  10.495 28.405 10.565 29.95 ;
        RECT  10.31 28.405 10.38 29.95 ;
        RECT  11.015 28.405 11.085 29.95 ;
        RECT  10.495 28.405 10.565 29.95 ;
        RECT  10.31 28.405 10.38 29.95 ;
        RECT  11.015 28.405 11.085 29.95 ;
        RECT  10.83 28.405 10.9 29.95 ;
        RECT  11.015 30.6 11.085 30.735 ;
        RECT  11.015 30.6 11.085 30.735 ;
        RECT  11.015 30.6 11.085 30.735 ;
        RECT  11.015 30.6 11.085 30.735 ;
        RECT  11.015 30.6 11.085 30.735 ;
        RECT  11.015 30.6 11.085 30.735 ;
        RECT  10.2775 29.815 10.4125 29.885 ;
        RECT  10.9825 29.815 11.1175 29.885 ;
        RECT  11.015 30.6 11.085 30.735 ;
        RECT  11.015 30.6 11.085 30.735 ;
        RECT  11.015 30.6 11.085 30.735 ;
        RECT  11.015 30.6 11.085 30.735 ;
        RECT  11.015 30.6 11.085 30.735 ;
        RECT  11.015 30.6 11.085 30.735 ;
        RECT  11.015 30.6 11.085 30.735 ;
        RECT  11.015 30.6 11.085 30.735 ;
        RECT  10.565 30.1075 10.635 30.2425 ;
        RECT  10.31 30.6 10.38 30.735 ;
        RECT  10.31 30.6 10.38 30.735 ;
        RECT  10.31 30.6 10.38 30.735 ;
        RECT  10.31 30.6 10.38 30.735 ;
        RECT  10.31 30.6 10.38 30.735 ;
        RECT  10.31 30.6 10.38 30.735 ;
        RECT  11.015 30.6 11.085 30.735 ;
        RECT  11.015 30.6 11.085 30.735 ;
        RECT  11.015 30.6 11.085 30.735 ;
        RECT  11.015 30.6 11.085 30.735 ;
        RECT  10.76 30.1075 10.83 30.2425 ;
        RECT  10.9825 29.815 11.1175 29.885 ;
        RECT  10.9825 29.815 11.1175 29.885 ;
        RECT  10.9825 29.815 11.1175 29.885 ;
        RECT  11.015 30.6 11.085 30.735 ;
        RECT  11.015 30.6 11.085 30.735 ;
        RECT  11.015 30.6 11.085 30.735 ;
        RECT  11.015 30.6 11.085 30.735 ;
        RECT  11.015 30.6 11.085 30.735 ;
        RECT  11.015 30.6 11.085 30.735 ;
        RECT  10.2775 29.815 10.4125 29.885 ;
        RECT  11.015 29.8175 11.085 31.2275 ;
        RECT  10.315 29.82 10.375 29.8775 ;
        RECT  10.5025 29.825 10.5575 29.8775 ;
        RECT  10.8375 29.8175 10.895 29.8775 ;
        RECT  11.02 29.825 11.08 29.8825 ;
        RECT  10.83 29.75 10.9 31.295 ;
        RECT  10.495 29.75 10.565 31.295 ;
        RECT  10.31 29.75 10.38 31.295 ;
        RECT  11.015 29.75 11.085 31.295 ;
        RECT  10.495 29.75 10.565 31.295 ;
        RECT  10.31 29.75 10.38 31.295 ;
        RECT  11.015 29.75 11.085 31.295 ;
        RECT  10.83 29.75 10.9 31.295 ;
        RECT  11.015 31.655 11.085 31.79 ;
        RECT  11.015 31.655 11.085 31.79 ;
        RECT  11.015 31.655 11.085 31.79 ;
        RECT  11.015 31.655 11.085 31.79 ;
        RECT  11.015 31.655 11.085 31.79 ;
        RECT  11.015 31.655 11.085 31.79 ;
        RECT  10.2775 32.505 10.4125 32.575 ;
        RECT  10.9825 32.505 11.1175 32.575 ;
        RECT  11.015 31.655 11.085 31.79 ;
        RECT  11.015 31.655 11.085 31.79 ;
        RECT  11.015 31.655 11.085 31.79 ;
        RECT  11.015 31.655 11.085 31.79 ;
        RECT  11.015 31.655 11.085 31.79 ;
        RECT  11.015 31.655 11.085 31.79 ;
        RECT  11.015 31.655 11.085 31.79 ;
        RECT  11.015 31.655 11.085 31.79 ;
        RECT  10.565 32.1475 10.635 32.2825 ;
        RECT  10.31 31.655 10.38 31.79 ;
        RECT  10.31 31.655 10.38 31.79 ;
        RECT  10.31 31.655 10.38 31.79 ;
        RECT  10.31 31.655 10.38 31.79 ;
        RECT  10.31 31.655 10.38 31.79 ;
        RECT  10.31 31.655 10.38 31.79 ;
        RECT  11.015 31.655 11.085 31.79 ;
        RECT  11.015 31.655 11.085 31.79 ;
        RECT  11.015 31.655 11.085 31.79 ;
        RECT  11.015 31.655 11.085 31.79 ;
        RECT  10.76 32.1475 10.83 32.2825 ;
        RECT  10.9825 32.505 11.1175 32.575 ;
        RECT  10.9825 32.505 11.1175 32.575 ;
        RECT  10.9825 32.505 11.1175 32.575 ;
        RECT  11.015 31.655 11.085 31.79 ;
        RECT  11.015 31.655 11.085 31.79 ;
        RECT  11.015 31.655 11.085 31.79 ;
        RECT  11.015 31.655 11.085 31.79 ;
        RECT  11.015 31.655 11.085 31.79 ;
        RECT  11.015 31.655 11.085 31.79 ;
        RECT  10.2775 32.505 10.4125 32.575 ;
        RECT  11.015 31.1625 11.085 32.5725 ;
        RECT  10.315 32.5125 10.375 32.57 ;
        RECT  10.5025 32.5125 10.5575 32.565 ;
        RECT  10.8375 32.5125 10.895 32.5725 ;
        RECT  11.02 32.5075 11.08 32.565 ;
        RECT  10.83 31.095 10.9 32.64 ;
        RECT  10.495 31.095 10.565 32.64 ;
        RECT  10.31 31.095 10.38 32.64 ;
        RECT  11.015 31.095 11.085 32.64 ;
        RECT  10.495 31.095 10.565 32.64 ;
        RECT  10.31 31.095 10.38 32.64 ;
        RECT  11.015 31.095 11.085 32.64 ;
        RECT  10.83 31.095 10.9 32.64 ;
        RECT  11.015 33.29 11.085 33.425 ;
        RECT  11.015 33.29 11.085 33.425 ;
        RECT  11.015 33.29 11.085 33.425 ;
        RECT  11.015 33.29 11.085 33.425 ;
        RECT  11.015 33.29 11.085 33.425 ;
        RECT  11.015 33.29 11.085 33.425 ;
        RECT  10.2775 32.505 10.4125 32.575 ;
        RECT  10.9825 32.505 11.1175 32.575 ;
        RECT  11.015 33.29 11.085 33.425 ;
        RECT  11.015 33.29 11.085 33.425 ;
        RECT  11.015 33.29 11.085 33.425 ;
        RECT  11.015 33.29 11.085 33.425 ;
        RECT  11.015 33.29 11.085 33.425 ;
        RECT  11.015 33.29 11.085 33.425 ;
        RECT  11.015 33.29 11.085 33.425 ;
        RECT  11.015 33.29 11.085 33.425 ;
        RECT  10.565 32.7975 10.635 32.9325 ;
        RECT  10.31 33.29 10.38 33.425 ;
        RECT  10.31 33.29 10.38 33.425 ;
        RECT  10.31 33.29 10.38 33.425 ;
        RECT  10.31 33.29 10.38 33.425 ;
        RECT  10.31 33.29 10.38 33.425 ;
        RECT  10.31 33.29 10.38 33.425 ;
        RECT  11.015 33.29 11.085 33.425 ;
        RECT  11.015 33.29 11.085 33.425 ;
        RECT  11.015 33.29 11.085 33.425 ;
        RECT  11.015 33.29 11.085 33.425 ;
        RECT  10.76 32.7975 10.83 32.9325 ;
        RECT  10.9825 32.505 11.1175 32.575 ;
        RECT  10.9825 32.505 11.1175 32.575 ;
        RECT  10.9825 32.505 11.1175 32.575 ;
        RECT  11.015 33.29 11.085 33.425 ;
        RECT  11.015 33.29 11.085 33.425 ;
        RECT  11.015 33.29 11.085 33.425 ;
        RECT  11.015 33.29 11.085 33.425 ;
        RECT  11.015 33.29 11.085 33.425 ;
        RECT  11.015 33.29 11.085 33.425 ;
        RECT  10.2775 32.505 10.4125 32.575 ;
        RECT  11.015 32.5075 11.085 33.9175 ;
        RECT  10.315 32.51 10.375 32.5675 ;
        RECT  10.5025 32.515 10.5575 32.5675 ;
        RECT  10.8375 32.5075 10.895 32.5675 ;
        RECT  11.02 32.515 11.08 32.5725 ;
        RECT  10.83 32.44 10.9 33.985 ;
        RECT  10.495 32.44 10.565 33.985 ;
        RECT  10.31 32.44 10.38 33.985 ;
        RECT  11.015 32.44 11.085 33.985 ;
        RECT  10.495 32.44 10.565 33.985 ;
        RECT  10.31 32.44 10.38 33.985 ;
        RECT  11.015 32.44 11.085 33.985 ;
        RECT  10.83 32.44 10.9 33.985 ;
        RECT  11.015 34.345 11.085 34.48 ;
        RECT  11.015 34.345 11.085 34.48 ;
        RECT  11.015 34.345 11.085 34.48 ;
        RECT  11.015 34.345 11.085 34.48 ;
        RECT  11.015 34.345 11.085 34.48 ;
        RECT  11.015 34.345 11.085 34.48 ;
        RECT  10.2775 35.195 10.4125 35.265 ;
        RECT  10.9825 35.195 11.1175 35.265 ;
        RECT  11.015 34.345 11.085 34.48 ;
        RECT  11.015 34.345 11.085 34.48 ;
        RECT  11.015 34.345 11.085 34.48 ;
        RECT  11.015 34.345 11.085 34.48 ;
        RECT  11.015 34.345 11.085 34.48 ;
        RECT  11.015 34.345 11.085 34.48 ;
        RECT  11.015 34.345 11.085 34.48 ;
        RECT  11.015 34.345 11.085 34.48 ;
        RECT  10.565 34.8375 10.635 34.9725 ;
        RECT  10.31 34.345 10.38 34.48 ;
        RECT  10.31 34.345 10.38 34.48 ;
        RECT  10.31 34.345 10.38 34.48 ;
        RECT  10.31 34.345 10.38 34.48 ;
        RECT  10.31 34.345 10.38 34.48 ;
        RECT  10.31 34.345 10.38 34.48 ;
        RECT  11.015 34.345 11.085 34.48 ;
        RECT  11.015 34.345 11.085 34.48 ;
        RECT  11.015 34.345 11.085 34.48 ;
        RECT  11.015 34.345 11.085 34.48 ;
        RECT  10.76 34.8375 10.83 34.9725 ;
        RECT  10.9825 35.195 11.1175 35.265 ;
        RECT  10.9825 35.195 11.1175 35.265 ;
        RECT  10.9825 35.195 11.1175 35.265 ;
        RECT  11.015 34.345 11.085 34.48 ;
        RECT  11.015 34.345 11.085 34.48 ;
        RECT  11.015 34.345 11.085 34.48 ;
        RECT  11.015 34.345 11.085 34.48 ;
        RECT  11.015 34.345 11.085 34.48 ;
        RECT  11.015 34.345 11.085 34.48 ;
        RECT  10.2775 35.195 10.4125 35.265 ;
        RECT  11.015 33.8525 11.085 35.2625 ;
        RECT  10.315 35.2025 10.375 35.26 ;
        RECT  10.5025 35.2025 10.5575 35.255 ;
        RECT  10.8375 35.2025 10.895 35.2625 ;
        RECT  11.02 35.1975 11.08 35.255 ;
        RECT  10.83 33.785 10.9 35.33 ;
        RECT  10.495 33.785 10.565 35.33 ;
        RECT  10.31 33.785 10.38 35.33 ;
        RECT  11.015 33.785 11.085 35.33 ;
        RECT  10.495 33.785 10.565 35.33 ;
        RECT  10.31 33.785 10.38 35.33 ;
        RECT  11.015 33.785 11.085 35.33 ;
        RECT  10.83 33.785 10.9 35.33 ;
        RECT  11.015 35.98 11.085 36.115 ;
        RECT  11.015 35.98 11.085 36.115 ;
        RECT  11.015 35.98 11.085 36.115 ;
        RECT  11.015 35.98 11.085 36.115 ;
        RECT  11.015 35.98 11.085 36.115 ;
        RECT  11.015 35.98 11.085 36.115 ;
        RECT  10.2775 35.195 10.4125 35.265 ;
        RECT  10.9825 35.195 11.1175 35.265 ;
        RECT  11.015 35.98 11.085 36.115 ;
        RECT  11.015 35.98 11.085 36.115 ;
        RECT  11.015 35.98 11.085 36.115 ;
        RECT  11.015 35.98 11.085 36.115 ;
        RECT  11.015 35.98 11.085 36.115 ;
        RECT  11.015 35.98 11.085 36.115 ;
        RECT  11.015 35.98 11.085 36.115 ;
        RECT  11.015 35.98 11.085 36.115 ;
        RECT  10.565 35.4875 10.635 35.6225 ;
        RECT  10.31 35.98 10.38 36.115 ;
        RECT  10.31 35.98 10.38 36.115 ;
        RECT  10.31 35.98 10.38 36.115 ;
        RECT  10.31 35.98 10.38 36.115 ;
        RECT  10.31 35.98 10.38 36.115 ;
        RECT  10.31 35.98 10.38 36.115 ;
        RECT  11.015 35.98 11.085 36.115 ;
        RECT  11.015 35.98 11.085 36.115 ;
        RECT  11.015 35.98 11.085 36.115 ;
        RECT  11.015 35.98 11.085 36.115 ;
        RECT  10.76 35.4875 10.83 35.6225 ;
        RECT  10.9825 35.195 11.1175 35.265 ;
        RECT  10.9825 35.195 11.1175 35.265 ;
        RECT  10.9825 35.195 11.1175 35.265 ;
        RECT  11.015 35.98 11.085 36.115 ;
        RECT  11.015 35.98 11.085 36.115 ;
        RECT  11.015 35.98 11.085 36.115 ;
        RECT  11.015 35.98 11.085 36.115 ;
        RECT  11.015 35.98 11.085 36.115 ;
        RECT  11.015 35.98 11.085 36.115 ;
        RECT  10.2775 35.195 10.4125 35.265 ;
        RECT  11.015 35.1975 11.085 36.6075 ;
        RECT  10.315 35.2 10.375 35.2575 ;
        RECT  10.5025 35.205 10.5575 35.2575 ;
        RECT  10.8375 35.1975 10.895 35.2575 ;
        RECT  11.02 35.205 11.08 35.2625 ;
        RECT  10.83 35.13 10.9 36.675 ;
        RECT  10.495 35.13 10.565 36.675 ;
        RECT  10.31 35.13 10.38 36.675 ;
        RECT  11.015 35.13 11.085 36.675 ;
        RECT  10.495 35.13 10.565 36.675 ;
        RECT  10.31 35.13 10.38 36.675 ;
        RECT  11.015 35.13 11.085 36.675 ;
        RECT  10.83 35.13 10.9 36.675 ;
        RECT  11.015 37.035 11.085 37.17 ;
        RECT  11.015 37.035 11.085 37.17 ;
        RECT  11.015 37.035 11.085 37.17 ;
        RECT  11.015 37.035 11.085 37.17 ;
        RECT  11.015 37.035 11.085 37.17 ;
        RECT  11.015 37.035 11.085 37.17 ;
        RECT  10.2775 37.885 10.4125 37.955 ;
        RECT  10.9825 37.885 11.1175 37.955 ;
        RECT  11.015 37.035 11.085 37.17 ;
        RECT  11.015 37.035 11.085 37.17 ;
        RECT  11.015 37.035 11.085 37.17 ;
        RECT  11.015 37.035 11.085 37.17 ;
        RECT  11.015 37.035 11.085 37.17 ;
        RECT  11.015 37.035 11.085 37.17 ;
        RECT  11.015 37.035 11.085 37.17 ;
        RECT  11.015 37.035 11.085 37.17 ;
        RECT  10.565 37.5275 10.635 37.6625 ;
        RECT  10.31 37.035 10.38 37.17 ;
        RECT  10.31 37.035 10.38 37.17 ;
        RECT  10.31 37.035 10.38 37.17 ;
        RECT  10.31 37.035 10.38 37.17 ;
        RECT  10.31 37.035 10.38 37.17 ;
        RECT  10.31 37.035 10.38 37.17 ;
        RECT  11.015 37.035 11.085 37.17 ;
        RECT  11.015 37.035 11.085 37.17 ;
        RECT  11.015 37.035 11.085 37.17 ;
        RECT  11.015 37.035 11.085 37.17 ;
        RECT  10.76 37.5275 10.83 37.6625 ;
        RECT  10.9825 37.885 11.1175 37.955 ;
        RECT  10.9825 37.885 11.1175 37.955 ;
        RECT  10.9825 37.885 11.1175 37.955 ;
        RECT  11.015 37.035 11.085 37.17 ;
        RECT  11.015 37.035 11.085 37.17 ;
        RECT  11.015 37.035 11.085 37.17 ;
        RECT  11.015 37.035 11.085 37.17 ;
        RECT  11.015 37.035 11.085 37.17 ;
        RECT  11.015 37.035 11.085 37.17 ;
        RECT  10.2775 37.885 10.4125 37.955 ;
        RECT  11.015 36.5425 11.085 37.9525 ;
        RECT  10.315 37.8925 10.375 37.95 ;
        RECT  10.5025 37.8925 10.5575 37.945 ;
        RECT  10.8375 37.8925 10.895 37.9525 ;
        RECT  11.02 37.8875 11.08 37.945 ;
        RECT  10.83 36.475 10.9 38.02 ;
        RECT  10.495 36.475 10.565 38.02 ;
        RECT  10.31 36.475 10.38 38.02 ;
        RECT  11.015 36.475 11.085 38.02 ;
        RECT  10.495 36.475 10.565 38.02 ;
        RECT  10.31 36.475 10.38 38.02 ;
        RECT  11.015 36.475 11.085 38.02 ;
        RECT  10.83 36.475 10.9 38.02 ;
        RECT  11.015 38.67 11.085 38.805 ;
        RECT  11.015 38.67 11.085 38.805 ;
        RECT  11.015 38.67 11.085 38.805 ;
        RECT  11.015 38.67 11.085 38.805 ;
        RECT  11.015 38.67 11.085 38.805 ;
        RECT  11.015 38.67 11.085 38.805 ;
        RECT  10.2775 37.885 10.4125 37.955 ;
        RECT  10.9825 37.885 11.1175 37.955 ;
        RECT  11.015 38.67 11.085 38.805 ;
        RECT  11.015 38.67 11.085 38.805 ;
        RECT  11.015 38.67 11.085 38.805 ;
        RECT  11.015 38.67 11.085 38.805 ;
        RECT  11.015 38.67 11.085 38.805 ;
        RECT  11.015 38.67 11.085 38.805 ;
        RECT  11.015 38.67 11.085 38.805 ;
        RECT  11.015 38.67 11.085 38.805 ;
        RECT  10.565 38.1775 10.635 38.3125 ;
        RECT  10.31 38.67 10.38 38.805 ;
        RECT  10.31 38.67 10.38 38.805 ;
        RECT  10.31 38.67 10.38 38.805 ;
        RECT  10.31 38.67 10.38 38.805 ;
        RECT  10.31 38.67 10.38 38.805 ;
        RECT  10.31 38.67 10.38 38.805 ;
        RECT  11.015 38.67 11.085 38.805 ;
        RECT  11.015 38.67 11.085 38.805 ;
        RECT  11.015 38.67 11.085 38.805 ;
        RECT  11.015 38.67 11.085 38.805 ;
        RECT  10.76 38.1775 10.83 38.3125 ;
        RECT  10.9825 37.885 11.1175 37.955 ;
        RECT  10.9825 37.885 11.1175 37.955 ;
        RECT  10.9825 37.885 11.1175 37.955 ;
        RECT  11.015 38.67 11.085 38.805 ;
        RECT  11.015 38.67 11.085 38.805 ;
        RECT  11.015 38.67 11.085 38.805 ;
        RECT  11.015 38.67 11.085 38.805 ;
        RECT  11.015 38.67 11.085 38.805 ;
        RECT  11.015 38.67 11.085 38.805 ;
        RECT  10.2775 37.885 10.4125 37.955 ;
        RECT  11.015 37.8875 11.085 39.2975 ;
        RECT  10.315 37.89 10.375 37.9475 ;
        RECT  10.5025 37.895 10.5575 37.9475 ;
        RECT  10.8375 37.8875 10.895 37.9475 ;
        RECT  11.02 37.895 11.08 37.9525 ;
        RECT  10.83 37.82 10.9 39.365 ;
        RECT  10.495 37.82 10.565 39.365 ;
        RECT  10.31 37.82 10.38 39.365 ;
        RECT  11.015 37.82 11.085 39.365 ;
        RECT  10.495 37.82 10.565 39.365 ;
        RECT  10.31 37.82 10.38 39.365 ;
        RECT  11.015 37.82 11.085 39.365 ;
        RECT  10.83 37.82 10.9 39.365 ;
        RECT  11.015 39.725 11.085 39.86 ;
        RECT  11.015 39.725 11.085 39.86 ;
        RECT  11.015 39.725 11.085 39.86 ;
        RECT  11.015 39.725 11.085 39.86 ;
        RECT  11.015 39.725 11.085 39.86 ;
        RECT  11.015 39.725 11.085 39.86 ;
        RECT  10.2775 40.575 10.4125 40.645 ;
        RECT  10.9825 40.575 11.1175 40.645 ;
        RECT  11.015 39.725 11.085 39.86 ;
        RECT  11.015 39.725 11.085 39.86 ;
        RECT  11.015 39.725 11.085 39.86 ;
        RECT  11.015 39.725 11.085 39.86 ;
        RECT  11.015 39.725 11.085 39.86 ;
        RECT  11.015 39.725 11.085 39.86 ;
        RECT  11.015 39.725 11.085 39.86 ;
        RECT  11.015 39.725 11.085 39.86 ;
        RECT  10.565 40.2175 10.635 40.3525 ;
        RECT  10.31 39.725 10.38 39.86 ;
        RECT  10.31 39.725 10.38 39.86 ;
        RECT  10.31 39.725 10.38 39.86 ;
        RECT  10.31 39.725 10.38 39.86 ;
        RECT  10.31 39.725 10.38 39.86 ;
        RECT  10.31 39.725 10.38 39.86 ;
        RECT  11.015 39.725 11.085 39.86 ;
        RECT  11.015 39.725 11.085 39.86 ;
        RECT  11.015 39.725 11.085 39.86 ;
        RECT  11.015 39.725 11.085 39.86 ;
        RECT  10.76 40.2175 10.83 40.3525 ;
        RECT  10.9825 40.575 11.1175 40.645 ;
        RECT  10.9825 40.575 11.1175 40.645 ;
        RECT  10.9825 40.575 11.1175 40.645 ;
        RECT  11.015 39.725 11.085 39.86 ;
        RECT  11.015 39.725 11.085 39.86 ;
        RECT  11.015 39.725 11.085 39.86 ;
        RECT  11.015 39.725 11.085 39.86 ;
        RECT  11.015 39.725 11.085 39.86 ;
        RECT  11.015 39.725 11.085 39.86 ;
        RECT  10.2775 40.575 10.4125 40.645 ;
        RECT  11.015 39.2325 11.085 40.6425 ;
        RECT  10.315 40.5825 10.375 40.64 ;
        RECT  10.5025 40.5825 10.5575 40.635 ;
        RECT  10.8375 40.5825 10.895 40.6425 ;
        RECT  11.02 40.5775 11.08 40.635 ;
        RECT  10.83 39.165 10.9 40.71 ;
        RECT  10.495 39.165 10.565 40.71 ;
        RECT  10.31 39.165 10.38 40.71 ;
        RECT  11.015 39.165 11.085 40.71 ;
        RECT  10.495 39.165 10.565 40.71 ;
        RECT  10.31 39.165 10.38 40.71 ;
        RECT  11.015 39.165 11.085 40.71 ;
        RECT  10.83 39.165 10.9 40.71 ;
        RECT  11.72 19.84 11.79 19.975 ;
        RECT  11.72 19.84 11.79 19.975 ;
        RECT  11.72 19.84 11.79 19.975 ;
        RECT  11.72 19.84 11.79 19.975 ;
        RECT  11.72 19.84 11.79 19.975 ;
        RECT  11.72 19.84 11.79 19.975 ;
        RECT  10.9825 19.055 11.1175 19.125 ;
        RECT  11.6875 19.055 11.8225 19.125 ;
        RECT  11.72 19.84 11.79 19.975 ;
        RECT  11.72 19.84 11.79 19.975 ;
        RECT  11.72 19.84 11.79 19.975 ;
        RECT  11.72 19.84 11.79 19.975 ;
        RECT  11.72 19.84 11.79 19.975 ;
        RECT  11.72 19.84 11.79 19.975 ;
        RECT  11.72 19.84 11.79 19.975 ;
        RECT  11.72 19.84 11.79 19.975 ;
        RECT  11.27 19.3475 11.34 19.4825 ;
        RECT  11.015 19.84 11.085 19.975 ;
        RECT  11.015 19.84 11.085 19.975 ;
        RECT  11.015 19.84 11.085 19.975 ;
        RECT  11.015 19.84 11.085 19.975 ;
        RECT  11.015 19.84 11.085 19.975 ;
        RECT  11.015 19.84 11.085 19.975 ;
        RECT  11.72 19.84 11.79 19.975 ;
        RECT  11.72 19.84 11.79 19.975 ;
        RECT  11.72 19.84 11.79 19.975 ;
        RECT  11.72 19.84 11.79 19.975 ;
        RECT  11.465 19.3475 11.535 19.4825 ;
        RECT  11.6875 19.055 11.8225 19.125 ;
        RECT  11.6875 19.055 11.8225 19.125 ;
        RECT  11.6875 19.055 11.8225 19.125 ;
        RECT  11.72 19.84 11.79 19.975 ;
        RECT  11.72 19.84 11.79 19.975 ;
        RECT  11.72 19.84 11.79 19.975 ;
        RECT  11.72 19.84 11.79 19.975 ;
        RECT  11.72 19.84 11.79 19.975 ;
        RECT  11.72 19.84 11.79 19.975 ;
        RECT  10.9825 19.055 11.1175 19.125 ;
        RECT  11.72 19.0575 11.79 20.4675 ;
        RECT  11.02 19.06 11.08 19.1175 ;
        RECT  11.2075 19.065 11.2625 19.1175 ;
        RECT  11.5425 19.0575 11.6 19.1175 ;
        RECT  11.725 19.065 11.785 19.1225 ;
        RECT  11.535 18.99 11.605 20.535 ;
        RECT  11.2 18.99 11.27 20.535 ;
        RECT  11.015 18.99 11.085 20.535 ;
        RECT  11.72 18.99 11.79 20.535 ;
        RECT  11.2 18.99 11.27 20.535 ;
        RECT  11.015 18.99 11.085 20.535 ;
        RECT  11.72 18.99 11.79 20.535 ;
        RECT  11.535 18.99 11.605 20.535 ;
        RECT  11.72 20.895 11.79 21.03 ;
        RECT  11.72 20.895 11.79 21.03 ;
        RECT  11.72 20.895 11.79 21.03 ;
        RECT  11.72 20.895 11.79 21.03 ;
        RECT  11.72 20.895 11.79 21.03 ;
        RECT  11.72 20.895 11.79 21.03 ;
        RECT  10.9825 21.745 11.1175 21.815 ;
        RECT  11.6875 21.745 11.8225 21.815 ;
        RECT  11.72 20.895 11.79 21.03 ;
        RECT  11.72 20.895 11.79 21.03 ;
        RECT  11.72 20.895 11.79 21.03 ;
        RECT  11.72 20.895 11.79 21.03 ;
        RECT  11.72 20.895 11.79 21.03 ;
        RECT  11.72 20.895 11.79 21.03 ;
        RECT  11.72 20.895 11.79 21.03 ;
        RECT  11.72 20.895 11.79 21.03 ;
        RECT  11.27 21.3875 11.34 21.5225 ;
        RECT  11.015 20.895 11.085 21.03 ;
        RECT  11.015 20.895 11.085 21.03 ;
        RECT  11.015 20.895 11.085 21.03 ;
        RECT  11.015 20.895 11.085 21.03 ;
        RECT  11.015 20.895 11.085 21.03 ;
        RECT  11.015 20.895 11.085 21.03 ;
        RECT  11.72 20.895 11.79 21.03 ;
        RECT  11.72 20.895 11.79 21.03 ;
        RECT  11.72 20.895 11.79 21.03 ;
        RECT  11.72 20.895 11.79 21.03 ;
        RECT  11.465 21.3875 11.535 21.5225 ;
        RECT  11.6875 21.745 11.8225 21.815 ;
        RECT  11.6875 21.745 11.8225 21.815 ;
        RECT  11.6875 21.745 11.8225 21.815 ;
        RECT  11.72 20.895 11.79 21.03 ;
        RECT  11.72 20.895 11.79 21.03 ;
        RECT  11.72 20.895 11.79 21.03 ;
        RECT  11.72 20.895 11.79 21.03 ;
        RECT  11.72 20.895 11.79 21.03 ;
        RECT  11.72 20.895 11.79 21.03 ;
        RECT  10.9825 21.745 11.1175 21.815 ;
        RECT  11.72 20.4025 11.79 21.8125 ;
        RECT  11.02 21.7525 11.08 21.81 ;
        RECT  11.2075 21.7525 11.2625 21.805 ;
        RECT  11.5425 21.7525 11.6 21.8125 ;
        RECT  11.725 21.7475 11.785 21.805 ;
        RECT  11.535 20.335 11.605 21.88 ;
        RECT  11.2 20.335 11.27 21.88 ;
        RECT  11.015 20.335 11.085 21.88 ;
        RECT  11.72 20.335 11.79 21.88 ;
        RECT  11.2 20.335 11.27 21.88 ;
        RECT  11.015 20.335 11.085 21.88 ;
        RECT  11.72 20.335 11.79 21.88 ;
        RECT  11.535 20.335 11.605 21.88 ;
        RECT  11.72 22.53 11.79 22.665 ;
        RECT  11.72 22.53 11.79 22.665 ;
        RECT  11.72 22.53 11.79 22.665 ;
        RECT  11.72 22.53 11.79 22.665 ;
        RECT  11.72 22.53 11.79 22.665 ;
        RECT  11.72 22.53 11.79 22.665 ;
        RECT  10.9825 21.745 11.1175 21.815 ;
        RECT  11.6875 21.745 11.8225 21.815 ;
        RECT  11.72 22.53 11.79 22.665 ;
        RECT  11.72 22.53 11.79 22.665 ;
        RECT  11.72 22.53 11.79 22.665 ;
        RECT  11.72 22.53 11.79 22.665 ;
        RECT  11.72 22.53 11.79 22.665 ;
        RECT  11.72 22.53 11.79 22.665 ;
        RECT  11.72 22.53 11.79 22.665 ;
        RECT  11.72 22.53 11.79 22.665 ;
        RECT  11.27 22.0375 11.34 22.1725 ;
        RECT  11.015 22.53 11.085 22.665 ;
        RECT  11.015 22.53 11.085 22.665 ;
        RECT  11.015 22.53 11.085 22.665 ;
        RECT  11.015 22.53 11.085 22.665 ;
        RECT  11.015 22.53 11.085 22.665 ;
        RECT  11.015 22.53 11.085 22.665 ;
        RECT  11.72 22.53 11.79 22.665 ;
        RECT  11.72 22.53 11.79 22.665 ;
        RECT  11.72 22.53 11.79 22.665 ;
        RECT  11.72 22.53 11.79 22.665 ;
        RECT  11.465 22.0375 11.535 22.1725 ;
        RECT  11.6875 21.745 11.8225 21.815 ;
        RECT  11.6875 21.745 11.8225 21.815 ;
        RECT  11.6875 21.745 11.8225 21.815 ;
        RECT  11.72 22.53 11.79 22.665 ;
        RECT  11.72 22.53 11.79 22.665 ;
        RECT  11.72 22.53 11.79 22.665 ;
        RECT  11.72 22.53 11.79 22.665 ;
        RECT  11.72 22.53 11.79 22.665 ;
        RECT  11.72 22.53 11.79 22.665 ;
        RECT  10.9825 21.745 11.1175 21.815 ;
        RECT  11.72 21.7475 11.79 23.1575 ;
        RECT  11.02 21.75 11.08 21.8075 ;
        RECT  11.2075 21.755 11.2625 21.8075 ;
        RECT  11.5425 21.7475 11.6 21.8075 ;
        RECT  11.725 21.755 11.785 21.8125 ;
        RECT  11.535 21.68 11.605 23.225 ;
        RECT  11.2 21.68 11.27 23.225 ;
        RECT  11.015 21.68 11.085 23.225 ;
        RECT  11.72 21.68 11.79 23.225 ;
        RECT  11.2 21.68 11.27 23.225 ;
        RECT  11.015 21.68 11.085 23.225 ;
        RECT  11.72 21.68 11.79 23.225 ;
        RECT  11.535 21.68 11.605 23.225 ;
        RECT  11.72 23.585 11.79 23.72 ;
        RECT  11.72 23.585 11.79 23.72 ;
        RECT  11.72 23.585 11.79 23.72 ;
        RECT  11.72 23.585 11.79 23.72 ;
        RECT  11.72 23.585 11.79 23.72 ;
        RECT  11.72 23.585 11.79 23.72 ;
        RECT  10.9825 24.435 11.1175 24.505 ;
        RECT  11.6875 24.435 11.8225 24.505 ;
        RECT  11.72 23.585 11.79 23.72 ;
        RECT  11.72 23.585 11.79 23.72 ;
        RECT  11.72 23.585 11.79 23.72 ;
        RECT  11.72 23.585 11.79 23.72 ;
        RECT  11.72 23.585 11.79 23.72 ;
        RECT  11.72 23.585 11.79 23.72 ;
        RECT  11.72 23.585 11.79 23.72 ;
        RECT  11.72 23.585 11.79 23.72 ;
        RECT  11.27 24.0775 11.34 24.2125 ;
        RECT  11.015 23.585 11.085 23.72 ;
        RECT  11.015 23.585 11.085 23.72 ;
        RECT  11.015 23.585 11.085 23.72 ;
        RECT  11.015 23.585 11.085 23.72 ;
        RECT  11.015 23.585 11.085 23.72 ;
        RECT  11.015 23.585 11.085 23.72 ;
        RECT  11.72 23.585 11.79 23.72 ;
        RECT  11.72 23.585 11.79 23.72 ;
        RECT  11.72 23.585 11.79 23.72 ;
        RECT  11.72 23.585 11.79 23.72 ;
        RECT  11.465 24.0775 11.535 24.2125 ;
        RECT  11.6875 24.435 11.8225 24.505 ;
        RECT  11.6875 24.435 11.8225 24.505 ;
        RECT  11.6875 24.435 11.8225 24.505 ;
        RECT  11.72 23.585 11.79 23.72 ;
        RECT  11.72 23.585 11.79 23.72 ;
        RECT  11.72 23.585 11.79 23.72 ;
        RECT  11.72 23.585 11.79 23.72 ;
        RECT  11.72 23.585 11.79 23.72 ;
        RECT  11.72 23.585 11.79 23.72 ;
        RECT  10.9825 24.435 11.1175 24.505 ;
        RECT  11.72 23.0925 11.79 24.5025 ;
        RECT  11.02 24.4425 11.08 24.5 ;
        RECT  11.2075 24.4425 11.2625 24.495 ;
        RECT  11.5425 24.4425 11.6 24.5025 ;
        RECT  11.725 24.4375 11.785 24.495 ;
        RECT  11.535 23.025 11.605 24.57 ;
        RECT  11.2 23.025 11.27 24.57 ;
        RECT  11.015 23.025 11.085 24.57 ;
        RECT  11.72 23.025 11.79 24.57 ;
        RECT  11.2 23.025 11.27 24.57 ;
        RECT  11.015 23.025 11.085 24.57 ;
        RECT  11.72 23.025 11.79 24.57 ;
        RECT  11.535 23.025 11.605 24.57 ;
        RECT  11.72 25.22 11.79 25.355 ;
        RECT  11.72 25.22 11.79 25.355 ;
        RECT  11.72 25.22 11.79 25.355 ;
        RECT  11.72 25.22 11.79 25.355 ;
        RECT  11.72 25.22 11.79 25.355 ;
        RECT  11.72 25.22 11.79 25.355 ;
        RECT  10.9825 24.435 11.1175 24.505 ;
        RECT  11.6875 24.435 11.8225 24.505 ;
        RECT  11.72 25.22 11.79 25.355 ;
        RECT  11.72 25.22 11.79 25.355 ;
        RECT  11.72 25.22 11.79 25.355 ;
        RECT  11.72 25.22 11.79 25.355 ;
        RECT  11.72 25.22 11.79 25.355 ;
        RECT  11.72 25.22 11.79 25.355 ;
        RECT  11.72 25.22 11.79 25.355 ;
        RECT  11.72 25.22 11.79 25.355 ;
        RECT  11.27 24.7275 11.34 24.8625 ;
        RECT  11.015 25.22 11.085 25.355 ;
        RECT  11.015 25.22 11.085 25.355 ;
        RECT  11.015 25.22 11.085 25.355 ;
        RECT  11.015 25.22 11.085 25.355 ;
        RECT  11.015 25.22 11.085 25.355 ;
        RECT  11.015 25.22 11.085 25.355 ;
        RECT  11.72 25.22 11.79 25.355 ;
        RECT  11.72 25.22 11.79 25.355 ;
        RECT  11.72 25.22 11.79 25.355 ;
        RECT  11.72 25.22 11.79 25.355 ;
        RECT  11.465 24.7275 11.535 24.8625 ;
        RECT  11.6875 24.435 11.8225 24.505 ;
        RECT  11.6875 24.435 11.8225 24.505 ;
        RECT  11.6875 24.435 11.8225 24.505 ;
        RECT  11.72 25.22 11.79 25.355 ;
        RECT  11.72 25.22 11.79 25.355 ;
        RECT  11.72 25.22 11.79 25.355 ;
        RECT  11.72 25.22 11.79 25.355 ;
        RECT  11.72 25.22 11.79 25.355 ;
        RECT  11.72 25.22 11.79 25.355 ;
        RECT  10.9825 24.435 11.1175 24.505 ;
        RECT  11.72 24.4375 11.79 25.8475 ;
        RECT  11.02 24.44 11.08 24.4975 ;
        RECT  11.2075 24.445 11.2625 24.4975 ;
        RECT  11.5425 24.4375 11.6 24.4975 ;
        RECT  11.725 24.445 11.785 24.5025 ;
        RECT  11.535 24.37 11.605 25.915 ;
        RECT  11.2 24.37 11.27 25.915 ;
        RECT  11.015 24.37 11.085 25.915 ;
        RECT  11.72 24.37 11.79 25.915 ;
        RECT  11.2 24.37 11.27 25.915 ;
        RECT  11.015 24.37 11.085 25.915 ;
        RECT  11.72 24.37 11.79 25.915 ;
        RECT  11.535 24.37 11.605 25.915 ;
        RECT  11.72 26.275 11.79 26.41 ;
        RECT  11.72 26.275 11.79 26.41 ;
        RECT  11.72 26.275 11.79 26.41 ;
        RECT  11.72 26.275 11.79 26.41 ;
        RECT  11.72 26.275 11.79 26.41 ;
        RECT  11.72 26.275 11.79 26.41 ;
        RECT  10.9825 27.125 11.1175 27.195 ;
        RECT  11.6875 27.125 11.8225 27.195 ;
        RECT  11.72 26.275 11.79 26.41 ;
        RECT  11.72 26.275 11.79 26.41 ;
        RECT  11.72 26.275 11.79 26.41 ;
        RECT  11.72 26.275 11.79 26.41 ;
        RECT  11.72 26.275 11.79 26.41 ;
        RECT  11.72 26.275 11.79 26.41 ;
        RECT  11.72 26.275 11.79 26.41 ;
        RECT  11.72 26.275 11.79 26.41 ;
        RECT  11.27 26.7675 11.34 26.9025 ;
        RECT  11.015 26.275 11.085 26.41 ;
        RECT  11.015 26.275 11.085 26.41 ;
        RECT  11.015 26.275 11.085 26.41 ;
        RECT  11.015 26.275 11.085 26.41 ;
        RECT  11.015 26.275 11.085 26.41 ;
        RECT  11.015 26.275 11.085 26.41 ;
        RECT  11.72 26.275 11.79 26.41 ;
        RECT  11.72 26.275 11.79 26.41 ;
        RECT  11.72 26.275 11.79 26.41 ;
        RECT  11.72 26.275 11.79 26.41 ;
        RECT  11.465 26.7675 11.535 26.9025 ;
        RECT  11.6875 27.125 11.8225 27.195 ;
        RECT  11.6875 27.125 11.8225 27.195 ;
        RECT  11.6875 27.125 11.8225 27.195 ;
        RECT  11.72 26.275 11.79 26.41 ;
        RECT  11.72 26.275 11.79 26.41 ;
        RECT  11.72 26.275 11.79 26.41 ;
        RECT  11.72 26.275 11.79 26.41 ;
        RECT  11.72 26.275 11.79 26.41 ;
        RECT  11.72 26.275 11.79 26.41 ;
        RECT  10.9825 27.125 11.1175 27.195 ;
        RECT  11.72 25.7825 11.79 27.1925 ;
        RECT  11.02 27.1325 11.08 27.19 ;
        RECT  11.2075 27.1325 11.2625 27.185 ;
        RECT  11.5425 27.1325 11.6 27.1925 ;
        RECT  11.725 27.1275 11.785 27.185 ;
        RECT  11.535 25.715 11.605 27.26 ;
        RECT  11.2 25.715 11.27 27.26 ;
        RECT  11.015 25.715 11.085 27.26 ;
        RECT  11.72 25.715 11.79 27.26 ;
        RECT  11.2 25.715 11.27 27.26 ;
        RECT  11.015 25.715 11.085 27.26 ;
        RECT  11.72 25.715 11.79 27.26 ;
        RECT  11.535 25.715 11.605 27.26 ;
        RECT  11.72 27.91 11.79 28.045 ;
        RECT  11.72 27.91 11.79 28.045 ;
        RECT  11.72 27.91 11.79 28.045 ;
        RECT  11.72 27.91 11.79 28.045 ;
        RECT  11.72 27.91 11.79 28.045 ;
        RECT  11.72 27.91 11.79 28.045 ;
        RECT  10.9825 27.125 11.1175 27.195 ;
        RECT  11.6875 27.125 11.8225 27.195 ;
        RECT  11.72 27.91 11.79 28.045 ;
        RECT  11.72 27.91 11.79 28.045 ;
        RECT  11.72 27.91 11.79 28.045 ;
        RECT  11.72 27.91 11.79 28.045 ;
        RECT  11.72 27.91 11.79 28.045 ;
        RECT  11.72 27.91 11.79 28.045 ;
        RECT  11.72 27.91 11.79 28.045 ;
        RECT  11.72 27.91 11.79 28.045 ;
        RECT  11.27 27.4175 11.34 27.5525 ;
        RECT  11.015 27.91 11.085 28.045 ;
        RECT  11.015 27.91 11.085 28.045 ;
        RECT  11.015 27.91 11.085 28.045 ;
        RECT  11.015 27.91 11.085 28.045 ;
        RECT  11.015 27.91 11.085 28.045 ;
        RECT  11.015 27.91 11.085 28.045 ;
        RECT  11.72 27.91 11.79 28.045 ;
        RECT  11.72 27.91 11.79 28.045 ;
        RECT  11.72 27.91 11.79 28.045 ;
        RECT  11.72 27.91 11.79 28.045 ;
        RECT  11.465 27.4175 11.535 27.5525 ;
        RECT  11.6875 27.125 11.8225 27.195 ;
        RECT  11.6875 27.125 11.8225 27.195 ;
        RECT  11.6875 27.125 11.8225 27.195 ;
        RECT  11.72 27.91 11.79 28.045 ;
        RECT  11.72 27.91 11.79 28.045 ;
        RECT  11.72 27.91 11.79 28.045 ;
        RECT  11.72 27.91 11.79 28.045 ;
        RECT  11.72 27.91 11.79 28.045 ;
        RECT  11.72 27.91 11.79 28.045 ;
        RECT  10.9825 27.125 11.1175 27.195 ;
        RECT  11.72 27.1275 11.79 28.5375 ;
        RECT  11.02 27.13 11.08 27.1875 ;
        RECT  11.2075 27.135 11.2625 27.1875 ;
        RECT  11.5425 27.1275 11.6 27.1875 ;
        RECT  11.725 27.135 11.785 27.1925 ;
        RECT  11.535 27.06 11.605 28.605 ;
        RECT  11.2 27.06 11.27 28.605 ;
        RECT  11.015 27.06 11.085 28.605 ;
        RECT  11.72 27.06 11.79 28.605 ;
        RECT  11.2 27.06 11.27 28.605 ;
        RECT  11.015 27.06 11.085 28.605 ;
        RECT  11.72 27.06 11.79 28.605 ;
        RECT  11.535 27.06 11.605 28.605 ;
        RECT  11.72 28.965 11.79 29.1 ;
        RECT  11.72 28.965 11.79 29.1 ;
        RECT  11.72 28.965 11.79 29.1 ;
        RECT  11.72 28.965 11.79 29.1 ;
        RECT  11.72 28.965 11.79 29.1 ;
        RECT  11.72 28.965 11.79 29.1 ;
        RECT  10.9825 29.815 11.1175 29.885 ;
        RECT  11.6875 29.815 11.8225 29.885 ;
        RECT  11.72 28.965 11.79 29.1 ;
        RECT  11.72 28.965 11.79 29.1 ;
        RECT  11.72 28.965 11.79 29.1 ;
        RECT  11.72 28.965 11.79 29.1 ;
        RECT  11.72 28.965 11.79 29.1 ;
        RECT  11.72 28.965 11.79 29.1 ;
        RECT  11.72 28.965 11.79 29.1 ;
        RECT  11.72 28.965 11.79 29.1 ;
        RECT  11.27 29.4575 11.34 29.5925 ;
        RECT  11.015 28.965 11.085 29.1 ;
        RECT  11.015 28.965 11.085 29.1 ;
        RECT  11.015 28.965 11.085 29.1 ;
        RECT  11.015 28.965 11.085 29.1 ;
        RECT  11.015 28.965 11.085 29.1 ;
        RECT  11.015 28.965 11.085 29.1 ;
        RECT  11.72 28.965 11.79 29.1 ;
        RECT  11.72 28.965 11.79 29.1 ;
        RECT  11.72 28.965 11.79 29.1 ;
        RECT  11.72 28.965 11.79 29.1 ;
        RECT  11.465 29.4575 11.535 29.5925 ;
        RECT  11.6875 29.815 11.8225 29.885 ;
        RECT  11.6875 29.815 11.8225 29.885 ;
        RECT  11.6875 29.815 11.8225 29.885 ;
        RECT  11.72 28.965 11.79 29.1 ;
        RECT  11.72 28.965 11.79 29.1 ;
        RECT  11.72 28.965 11.79 29.1 ;
        RECT  11.72 28.965 11.79 29.1 ;
        RECT  11.72 28.965 11.79 29.1 ;
        RECT  11.72 28.965 11.79 29.1 ;
        RECT  10.9825 29.815 11.1175 29.885 ;
        RECT  11.72 28.4725 11.79 29.8825 ;
        RECT  11.02 29.8225 11.08 29.88 ;
        RECT  11.2075 29.8225 11.2625 29.875 ;
        RECT  11.5425 29.8225 11.6 29.8825 ;
        RECT  11.725 29.8175 11.785 29.875 ;
        RECT  11.535 28.405 11.605 29.95 ;
        RECT  11.2 28.405 11.27 29.95 ;
        RECT  11.015 28.405 11.085 29.95 ;
        RECT  11.72 28.405 11.79 29.95 ;
        RECT  11.2 28.405 11.27 29.95 ;
        RECT  11.015 28.405 11.085 29.95 ;
        RECT  11.72 28.405 11.79 29.95 ;
        RECT  11.535 28.405 11.605 29.95 ;
        RECT  11.72 30.6 11.79 30.735 ;
        RECT  11.72 30.6 11.79 30.735 ;
        RECT  11.72 30.6 11.79 30.735 ;
        RECT  11.72 30.6 11.79 30.735 ;
        RECT  11.72 30.6 11.79 30.735 ;
        RECT  11.72 30.6 11.79 30.735 ;
        RECT  10.9825 29.815 11.1175 29.885 ;
        RECT  11.6875 29.815 11.8225 29.885 ;
        RECT  11.72 30.6 11.79 30.735 ;
        RECT  11.72 30.6 11.79 30.735 ;
        RECT  11.72 30.6 11.79 30.735 ;
        RECT  11.72 30.6 11.79 30.735 ;
        RECT  11.72 30.6 11.79 30.735 ;
        RECT  11.72 30.6 11.79 30.735 ;
        RECT  11.72 30.6 11.79 30.735 ;
        RECT  11.72 30.6 11.79 30.735 ;
        RECT  11.27 30.1075 11.34 30.2425 ;
        RECT  11.015 30.6 11.085 30.735 ;
        RECT  11.015 30.6 11.085 30.735 ;
        RECT  11.015 30.6 11.085 30.735 ;
        RECT  11.015 30.6 11.085 30.735 ;
        RECT  11.015 30.6 11.085 30.735 ;
        RECT  11.015 30.6 11.085 30.735 ;
        RECT  11.72 30.6 11.79 30.735 ;
        RECT  11.72 30.6 11.79 30.735 ;
        RECT  11.72 30.6 11.79 30.735 ;
        RECT  11.72 30.6 11.79 30.735 ;
        RECT  11.465 30.1075 11.535 30.2425 ;
        RECT  11.6875 29.815 11.8225 29.885 ;
        RECT  11.6875 29.815 11.8225 29.885 ;
        RECT  11.6875 29.815 11.8225 29.885 ;
        RECT  11.72 30.6 11.79 30.735 ;
        RECT  11.72 30.6 11.79 30.735 ;
        RECT  11.72 30.6 11.79 30.735 ;
        RECT  11.72 30.6 11.79 30.735 ;
        RECT  11.72 30.6 11.79 30.735 ;
        RECT  11.72 30.6 11.79 30.735 ;
        RECT  10.9825 29.815 11.1175 29.885 ;
        RECT  11.72 29.8175 11.79 31.2275 ;
        RECT  11.02 29.82 11.08 29.8775 ;
        RECT  11.2075 29.825 11.2625 29.8775 ;
        RECT  11.5425 29.8175 11.6 29.8775 ;
        RECT  11.725 29.825 11.785 29.8825 ;
        RECT  11.535 29.75 11.605 31.295 ;
        RECT  11.2 29.75 11.27 31.295 ;
        RECT  11.015 29.75 11.085 31.295 ;
        RECT  11.72 29.75 11.79 31.295 ;
        RECT  11.2 29.75 11.27 31.295 ;
        RECT  11.015 29.75 11.085 31.295 ;
        RECT  11.72 29.75 11.79 31.295 ;
        RECT  11.535 29.75 11.605 31.295 ;
        RECT  11.72 31.655 11.79 31.79 ;
        RECT  11.72 31.655 11.79 31.79 ;
        RECT  11.72 31.655 11.79 31.79 ;
        RECT  11.72 31.655 11.79 31.79 ;
        RECT  11.72 31.655 11.79 31.79 ;
        RECT  11.72 31.655 11.79 31.79 ;
        RECT  10.9825 32.505 11.1175 32.575 ;
        RECT  11.6875 32.505 11.8225 32.575 ;
        RECT  11.72 31.655 11.79 31.79 ;
        RECT  11.72 31.655 11.79 31.79 ;
        RECT  11.72 31.655 11.79 31.79 ;
        RECT  11.72 31.655 11.79 31.79 ;
        RECT  11.72 31.655 11.79 31.79 ;
        RECT  11.72 31.655 11.79 31.79 ;
        RECT  11.72 31.655 11.79 31.79 ;
        RECT  11.72 31.655 11.79 31.79 ;
        RECT  11.27 32.1475 11.34 32.2825 ;
        RECT  11.015 31.655 11.085 31.79 ;
        RECT  11.015 31.655 11.085 31.79 ;
        RECT  11.015 31.655 11.085 31.79 ;
        RECT  11.015 31.655 11.085 31.79 ;
        RECT  11.015 31.655 11.085 31.79 ;
        RECT  11.015 31.655 11.085 31.79 ;
        RECT  11.72 31.655 11.79 31.79 ;
        RECT  11.72 31.655 11.79 31.79 ;
        RECT  11.72 31.655 11.79 31.79 ;
        RECT  11.72 31.655 11.79 31.79 ;
        RECT  11.465 32.1475 11.535 32.2825 ;
        RECT  11.6875 32.505 11.8225 32.575 ;
        RECT  11.6875 32.505 11.8225 32.575 ;
        RECT  11.6875 32.505 11.8225 32.575 ;
        RECT  11.72 31.655 11.79 31.79 ;
        RECT  11.72 31.655 11.79 31.79 ;
        RECT  11.72 31.655 11.79 31.79 ;
        RECT  11.72 31.655 11.79 31.79 ;
        RECT  11.72 31.655 11.79 31.79 ;
        RECT  11.72 31.655 11.79 31.79 ;
        RECT  10.9825 32.505 11.1175 32.575 ;
        RECT  11.72 31.1625 11.79 32.5725 ;
        RECT  11.02 32.5125 11.08 32.57 ;
        RECT  11.2075 32.5125 11.2625 32.565 ;
        RECT  11.5425 32.5125 11.6 32.5725 ;
        RECT  11.725 32.5075 11.785 32.565 ;
        RECT  11.535 31.095 11.605 32.64 ;
        RECT  11.2 31.095 11.27 32.64 ;
        RECT  11.015 31.095 11.085 32.64 ;
        RECT  11.72 31.095 11.79 32.64 ;
        RECT  11.2 31.095 11.27 32.64 ;
        RECT  11.015 31.095 11.085 32.64 ;
        RECT  11.72 31.095 11.79 32.64 ;
        RECT  11.535 31.095 11.605 32.64 ;
        RECT  11.72 33.29 11.79 33.425 ;
        RECT  11.72 33.29 11.79 33.425 ;
        RECT  11.72 33.29 11.79 33.425 ;
        RECT  11.72 33.29 11.79 33.425 ;
        RECT  11.72 33.29 11.79 33.425 ;
        RECT  11.72 33.29 11.79 33.425 ;
        RECT  10.9825 32.505 11.1175 32.575 ;
        RECT  11.6875 32.505 11.8225 32.575 ;
        RECT  11.72 33.29 11.79 33.425 ;
        RECT  11.72 33.29 11.79 33.425 ;
        RECT  11.72 33.29 11.79 33.425 ;
        RECT  11.72 33.29 11.79 33.425 ;
        RECT  11.72 33.29 11.79 33.425 ;
        RECT  11.72 33.29 11.79 33.425 ;
        RECT  11.72 33.29 11.79 33.425 ;
        RECT  11.72 33.29 11.79 33.425 ;
        RECT  11.27 32.7975 11.34 32.9325 ;
        RECT  11.015 33.29 11.085 33.425 ;
        RECT  11.015 33.29 11.085 33.425 ;
        RECT  11.015 33.29 11.085 33.425 ;
        RECT  11.015 33.29 11.085 33.425 ;
        RECT  11.015 33.29 11.085 33.425 ;
        RECT  11.015 33.29 11.085 33.425 ;
        RECT  11.72 33.29 11.79 33.425 ;
        RECT  11.72 33.29 11.79 33.425 ;
        RECT  11.72 33.29 11.79 33.425 ;
        RECT  11.72 33.29 11.79 33.425 ;
        RECT  11.465 32.7975 11.535 32.9325 ;
        RECT  11.6875 32.505 11.8225 32.575 ;
        RECT  11.6875 32.505 11.8225 32.575 ;
        RECT  11.6875 32.505 11.8225 32.575 ;
        RECT  11.72 33.29 11.79 33.425 ;
        RECT  11.72 33.29 11.79 33.425 ;
        RECT  11.72 33.29 11.79 33.425 ;
        RECT  11.72 33.29 11.79 33.425 ;
        RECT  11.72 33.29 11.79 33.425 ;
        RECT  11.72 33.29 11.79 33.425 ;
        RECT  10.9825 32.505 11.1175 32.575 ;
        RECT  11.72 32.5075 11.79 33.9175 ;
        RECT  11.02 32.51 11.08 32.5675 ;
        RECT  11.2075 32.515 11.2625 32.5675 ;
        RECT  11.5425 32.5075 11.6 32.5675 ;
        RECT  11.725 32.515 11.785 32.5725 ;
        RECT  11.535 32.44 11.605 33.985 ;
        RECT  11.2 32.44 11.27 33.985 ;
        RECT  11.015 32.44 11.085 33.985 ;
        RECT  11.72 32.44 11.79 33.985 ;
        RECT  11.2 32.44 11.27 33.985 ;
        RECT  11.015 32.44 11.085 33.985 ;
        RECT  11.72 32.44 11.79 33.985 ;
        RECT  11.535 32.44 11.605 33.985 ;
        RECT  11.72 34.345 11.79 34.48 ;
        RECT  11.72 34.345 11.79 34.48 ;
        RECT  11.72 34.345 11.79 34.48 ;
        RECT  11.72 34.345 11.79 34.48 ;
        RECT  11.72 34.345 11.79 34.48 ;
        RECT  11.72 34.345 11.79 34.48 ;
        RECT  10.9825 35.195 11.1175 35.265 ;
        RECT  11.6875 35.195 11.8225 35.265 ;
        RECT  11.72 34.345 11.79 34.48 ;
        RECT  11.72 34.345 11.79 34.48 ;
        RECT  11.72 34.345 11.79 34.48 ;
        RECT  11.72 34.345 11.79 34.48 ;
        RECT  11.72 34.345 11.79 34.48 ;
        RECT  11.72 34.345 11.79 34.48 ;
        RECT  11.72 34.345 11.79 34.48 ;
        RECT  11.72 34.345 11.79 34.48 ;
        RECT  11.27 34.8375 11.34 34.9725 ;
        RECT  11.015 34.345 11.085 34.48 ;
        RECT  11.015 34.345 11.085 34.48 ;
        RECT  11.015 34.345 11.085 34.48 ;
        RECT  11.015 34.345 11.085 34.48 ;
        RECT  11.015 34.345 11.085 34.48 ;
        RECT  11.015 34.345 11.085 34.48 ;
        RECT  11.72 34.345 11.79 34.48 ;
        RECT  11.72 34.345 11.79 34.48 ;
        RECT  11.72 34.345 11.79 34.48 ;
        RECT  11.72 34.345 11.79 34.48 ;
        RECT  11.465 34.8375 11.535 34.9725 ;
        RECT  11.6875 35.195 11.8225 35.265 ;
        RECT  11.6875 35.195 11.8225 35.265 ;
        RECT  11.6875 35.195 11.8225 35.265 ;
        RECT  11.72 34.345 11.79 34.48 ;
        RECT  11.72 34.345 11.79 34.48 ;
        RECT  11.72 34.345 11.79 34.48 ;
        RECT  11.72 34.345 11.79 34.48 ;
        RECT  11.72 34.345 11.79 34.48 ;
        RECT  11.72 34.345 11.79 34.48 ;
        RECT  10.9825 35.195 11.1175 35.265 ;
        RECT  11.72 33.8525 11.79 35.2625 ;
        RECT  11.02 35.2025 11.08 35.26 ;
        RECT  11.2075 35.2025 11.2625 35.255 ;
        RECT  11.5425 35.2025 11.6 35.2625 ;
        RECT  11.725 35.1975 11.785 35.255 ;
        RECT  11.535 33.785 11.605 35.33 ;
        RECT  11.2 33.785 11.27 35.33 ;
        RECT  11.015 33.785 11.085 35.33 ;
        RECT  11.72 33.785 11.79 35.33 ;
        RECT  11.2 33.785 11.27 35.33 ;
        RECT  11.015 33.785 11.085 35.33 ;
        RECT  11.72 33.785 11.79 35.33 ;
        RECT  11.535 33.785 11.605 35.33 ;
        RECT  11.72 35.98 11.79 36.115 ;
        RECT  11.72 35.98 11.79 36.115 ;
        RECT  11.72 35.98 11.79 36.115 ;
        RECT  11.72 35.98 11.79 36.115 ;
        RECT  11.72 35.98 11.79 36.115 ;
        RECT  11.72 35.98 11.79 36.115 ;
        RECT  10.9825 35.195 11.1175 35.265 ;
        RECT  11.6875 35.195 11.8225 35.265 ;
        RECT  11.72 35.98 11.79 36.115 ;
        RECT  11.72 35.98 11.79 36.115 ;
        RECT  11.72 35.98 11.79 36.115 ;
        RECT  11.72 35.98 11.79 36.115 ;
        RECT  11.72 35.98 11.79 36.115 ;
        RECT  11.72 35.98 11.79 36.115 ;
        RECT  11.72 35.98 11.79 36.115 ;
        RECT  11.72 35.98 11.79 36.115 ;
        RECT  11.27 35.4875 11.34 35.6225 ;
        RECT  11.015 35.98 11.085 36.115 ;
        RECT  11.015 35.98 11.085 36.115 ;
        RECT  11.015 35.98 11.085 36.115 ;
        RECT  11.015 35.98 11.085 36.115 ;
        RECT  11.015 35.98 11.085 36.115 ;
        RECT  11.015 35.98 11.085 36.115 ;
        RECT  11.72 35.98 11.79 36.115 ;
        RECT  11.72 35.98 11.79 36.115 ;
        RECT  11.72 35.98 11.79 36.115 ;
        RECT  11.72 35.98 11.79 36.115 ;
        RECT  11.465 35.4875 11.535 35.6225 ;
        RECT  11.6875 35.195 11.8225 35.265 ;
        RECT  11.6875 35.195 11.8225 35.265 ;
        RECT  11.6875 35.195 11.8225 35.265 ;
        RECT  11.72 35.98 11.79 36.115 ;
        RECT  11.72 35.98 11.79 36.115 ;
        RECT  11.72 35.98 11.79 36.115 ;
        RECT  11.72 35.98 11.79 36.115 ;
        RECT  11.72 35.98 11.79 36.115 ;
        RECT  11.72 35.98 11.79 36.115 ;
        RECT  10.9825 35.195 11.1175 35.265 ;
        RECT  11.72 35.1975 11.79 36.6075 ;
        RECT  11.02 35.2 11.08 35.2575 ;
        RECT  11.2075 35.205 11.2625 35.2575 ;
        RECT  11.5425 35.1975 11.6 35.2575 ;
        RECT  11.725 35.205 11.785 35.2625 ;
        RECT  11.535 35.13 11.605 36.675 ;
        RECT  11.2 35.13 11.27 36.675 ;
        RECT  11.015 35.13 11.085 36.675 ;
        RECT  11.72 35.13 11.79 36.675 ;
        RECT  11.2 35.13 11.27 36.675 ;
        RECT  11.015 35.13 11.085 36.675 ;
        RECT  11.72 35.13 11.79 36.675 ;
        RECT  11.535 35.13 11.605 36.675 ;
        RECT  11.72 37.035 11.79 37.17 ;
        RECT  11.72 37.035 11.79 37.17 ;
        RECT  11.72 37.035 11.79 37.17 ;
        RECT  11.72 37.035 11.79 37.17 ;
        RECT  11.72 37.035 11.79 37.17 ;
        RECT  11.72 37.035 11.79 37.17 ;
        RECT  10.9825 37.885 11.1175 37.955 ;
        RECT  11.6875 37.885 11.8225 37.955 ;
        RECT  11.72 37.035 11.79 37.17 ;
        RECT  11.72 37.035 11.79 37.17 ;
        RECT  11.72 37.035 11.79 37.17 ;
        RECT  11.72 37.035 11.79 37.17 ;
        RECT  11.72 37.035 11.79 37.17 ;
        RECT  11.72 37.035 11.79 37.17 ;
        RECT  11.72 37.035 11.79 37.17 ;
        RECT  11.72 37.035 11.79 37.17 ;
        RECT  11.27 37.5275 11.34 37.6625 ;
        RECT  11.015 37.035 11.085 37.17 ;
        RECT  11.015 37.035 11.085 37.17 ;
        RECT  11.015 37.035 11.085 37.17 ;
        RECT  11.015 37.035 11.085 37.17 ;
        RECT  11.015 37.035 11.085 37.17 ;
        RECT  11.015 37.035 11.085 37.17 ;
        RECT  11.72 37.035 11.79 37.17 ;
        RECT  11.72 37.035 11.79 37.17 ;
        RECT  11.72 37.035 11.79 37.17 ;
        RECT  11.72 37.035 11.79 37.17 ;
        RECT  11.465 37.5275 11.535 37.6625 ;
        RECT  11.6875 37.885 11.8225 37.955 ;
        RECT  11.6875 37.885 11.8225 37.955 ;
        RECT  11.6875 37.885 11.8225 37.955 ;
        RECT  11.72 37.035 11.79 37.17 ;
        RECT  11.72 37.035 11.79 37.17 ;
        RECT  11.72 37.035 11.79 37.17 ;
        RECT  11.72 37.035 11.79 37.17 ;
        RECT  11.72 37.035 11.79 37.17 ;
        RECT  11.72 37.035 11.79 37.17 ;
        RECT  10.9825 37.885 11.1175 37.955 ;
        RECT  11.72 36.5425 11.79 37.9525 ;
        RECT  11.02 37.8925 11.08 37.95 ;
        RECT  11.2075 37.8925 11.2625 37.945 ;
        RECT  11.5425 37.8925 11.6 37.9525 ;
        RECT  11.725 37.8875 11.785 37.945 ;
        RECT  11.535 36.475 11.605 38.02 ;
        RECT  11.2 36.475 11.27 38.02 ;
        RECT  11.015 36.475 11.085 38.02 ;
        RECT  11.72 36.475 11.79 38.02 ;
        RECT  11.2 36.475 11.27 38.02 ;
        RECT  11.015 36.475 11.085 38.02 ;
        RECT  11.72 36.475 11.79 38.02 ;
        RECT  11.535 36.475 11.605 38.02 ;
        RECT  11.72 38.67 11.79 38.805 ;
        RECT  11.72 38.67 11.79 38.805 ;
        RECT  11.72 38.67 11.79 38.805 ;
        RECT  11.72 38.67 11.79 38.805 ;
        RECT  11.72 38.67 11.79 38.805 ;
        RECT  11.72 38.67 11.79 38.805 ;
        RECT  10.9825 37.885 11.1175 37.955 ;
        RECT  11.6875 37.885 11.8225 37.955 ;
        RECT  11.72 38.67 11.79 38.805 ;
        RECT  11.72 38.67 11.79 38.805 ;
        RECT  11.72 38.67 11.79 38.805 ;
        RECT  11.72 38.67 11.79 38.805 ;
        RECT  11.72 38.67 11.79 38.805 ;
        RECT  11.72 38.67 11.79 38.805 ;
        RECT  11.72 38.67 11.79 38.805 ;
        RECT  11.72 38.67 11.79 38.805 ;
        RECT  11.27 38.1775 11.34 38.3125 ;
        RECT  11.015 38.67 11.085 38.805 ;
        RECT  11.015 38.67 11.085 38.805 ;
        RECT  11.015 38.67 11.085 38.805 ;
        RECT  11.015 38.67 11.085 38.805 ;
        RECT  11.015 38.67 11.085 38.805 ;
        RECT  11.015 38.67 11.085 38.805 ;
        RECT  11.72 38.67 11.79 38.805 ;
        RECT  11.72 38.67 11.79 38.805 ;
        RECT  11.72 38.67 11.79 38.805 ;
        RECT  11.72 38.67 11.79 38.805 ;
        RECT  11.465 38.1775 11.535 38.3125 ;
        RECT  11.6875 37.885 11.8225 37.955 ;
        RECT  11.6875 37.885 11.8225 37.955 ;
        RECT  11.6875 37.885 11.8225 37.955 ;
        RECT  11.72 38.67 11.79 38.805 ;
        RECT  11.72 38.67 11.79 38.805 ;
        RECT  11.72 38.67 11.79 38.805 ;
        RECT  11.72 38.67 11.79 38.805 ;
        RECT  11.72 38.67 11.79 38.805 ;
        RECT  11.72 38.67 11.79 38.805 ;
        RECT  10.9825 37.885 11.1175 37.955 ;
        RECT  11.72 37.8875 11.79 39.2975 ;
        RECT  11.02 37.89 11.08 37.9475 ;
        RECT  11.2075 37.895 11.2625 37.9475 ;
        RECT  11.5425 37.8875 11.6 37.9475 ;
        RECT  11.725 37.895 11.785 37.9525 ;
        RECT  11.535 37.82 11.605 39.365 ;
        RECT  11.2 37.82 11.27 39.365 ;
        RECT  11.015 37.82 11.085 39.365 ;
        RECT  11.72 37.82 11.79 39.365 ;
        RECT  11.2 37.82 11.27 39.365 ;
        RECT  11.015 37.82 11.085 39.365 ;
        RECT  11.72 37.82 11.79 39.365 ;
        RECT  11.535 37.82 11.605 39.365 ;
        RECT  11.72 39.725 11.79 39.86 ;
        RECT  11.72 39.725 11.79 39.86 ;
        RECT  11.72 39.725 11.79 39.86 ;
        RECT  11.72 39.725 11.79 39.86 ;
        RECT  11.72 39.725 11.79 39.86 ;
        RECT  11.72 39.725 11.79 39.86 ;
        RECT  10.9825 40.575 11.1175 40.645 ;
        RECT  11.6875 40.575 11.8225 40.645 ;
        RECT  11.72 39.725 11.79 39.86 ;
        RECT  11.72 39.725 11.79 39.86 ;
        RECT  11.72 39.725 11.79 39.86 ;
        RECT  11.72 39.725 11.79 39.86 ;
        RECT  11.72 39.725 11.79 39.86 ;
        RECT  11.72 39.725 11.79 39.86 ;
        RECT  11.72 39.725 11.79 39.86 ;
        RECT  11.72 39.725 11.79 39.86 ;
        RECT  11.27 40.2175 11.34 40.3525 ;
        RECT  11.015 39.725 11.085 39.86 ;
        RECT  11.015 39.725 11.085 39.86 ;
        RECT  11.015 39.725 11.085 39.86 ;
        RECT  11.015 39.725 11.085 39.86 ;
        RECT  11.015 39.725 11.085 39.86 ;
        RECT  11.015 39.725 11.085 39.86 ;
        RECT  11.72 39.725 11.79 39.86 ;
        RECT  11.72 39.725 11.79 39.86 ;
        RECT  11.72 39.725 11.79 39.86 ;
        RECT  11.72 39.725 11.79 39.86 ;
        RECT  11.465 40.2175 11.535 40.3525 ;
        RECT  11.6875 40.575 11.8225 40.645 ;
        RECT  11.6875 40.575 11.8225 40.645 ;
        RECT  11.6875 40.575 11.8225 40.645 ;
        RECT  11.72 39.725 11.79 39.86 ;
        RECT  11.72 39.725 11.79 39.86 ;
        RECT  11.72 39.725 11.79 39.86 ;
        RECT  11.72 39.725 11.79 39.86 ;
        RECT  11.72 39.725 11.79 39.86 ;
        RECT  11.72 39.725 11.79 39.86 ;
        RECT  10.9825 40.575 11.1175 40.645 ;
        RECT  11.72 39.2325 11.79 40.6425 ;
        RECT  11.02 40.5825 11.08 40.64 ;
        RECT  11.2075 40.5825 11.2625 40.635 ;
        RECT  11.5425 40.5825 11.6 40.6425 ;
        RECT  11.725 40.5775 11.785 40.635 ;
        RECT  11.535 39.165 11.605 40.71 ;
        RECT  11.2 39.165 11.27 40.71 ;
        RECT  11.015 39.165 11.085 40.71 ;
        RECT  11.72 39.165 11.79 40.71 ;
        RECT  11.2 39.165 11.27 40.71 ;
        RECT  11.015 39.165 11.085 40.71 ;
        RECT  11.72 39.165 11.79 40.71 ;
        RECT  11.535 39.165 11.605 40.71 ;
        RECT  11.2 41.06 11.27 42.02 ;
        RECT  10.495 41.06 10.565 42.02 ;
        RECT  11.535 41.06 11.605 42.02 ;
        RECT  10.83 41.06 10.9 42.02 ;
        RECT  10.53 41.6075 10.5725 41.7425 ;
        RECT  10.83 41.6075 10.9175 41.7425 ;
        RECT  10.53 41.1575 10.575 41.2925 ;
        RECT  10.73 41.1575 10.83 41.2925 ;
        RECT  10.495 41.06 10.565 42.02 ;
        RECT  10.83 41.06 10.9 42.02 ;
        RECT  10.5375 41.6075 10.6075 41.7425 ;
        RECT  10.9175 41.6075 10.9875 41.7425 ;
        RECT  10.5375 41.1575 10.6075 41.2925 ;
        RECT  10.7275 41.1575 10.7975 41.2925 ;
        RECT  11.235 41.6075 11.2775 41.7425 ;
        RECT  11.535 41.6075 11.6225 41.7425 ;
        RECT  11.235 41.1575 11.28 41.2925 ;
        RECT  11.435 41.1575 11.535 41.2925 ;
        RECT  11.2 41.06 11.27 42.02 ;
        RECT  11.535 41.06 11.605 42.02 ;
        RECT  11.2425 41.6075 11.3125 41.7425 ;
        RECT  11.6225 41.6075 11.6925 41.7425 ;
        RECT  11.2425 41.1575 11.3125 41.2925 ;
        RECT  11.4325 41.1575 11.5025 41.2925 ;
        RECT  11.2 14.205 11.27 19.09 ;
        RECT  10.495 14.205 10.565 19.09 ;
        RECT  11.535 14.205 11.605 18.29 ;
        RECT  10.83 14.205 10.9 18.29 ;
        RECT  10.31 14.205 10.38 19.09 ;
        RECT  10.495 14.205 10.565 19.09 ;
        RECT  10.83 14.205 10.9 17.75 ;
        RECT  10.6625 16.48 10.7325 18.49 ;
        RECT  10.83 15.005 10.9 19.09 ;
        RECT  11.015 14.205 11.085 19.09 ;
        RECT  10.835 19.04 10.895 19.09 ;
        RECT  10.495 19.03 10.565 19.09 ;
        RECT  10.6575 19.035 10.7275 19.09 ;
        RECT  10.6575 18.6925 10.7275 19.09 ;
        RECT  10.6625 16.345 10.7325 16.48 ;
        RECT  10.6625 18.4875 10.7325 18.6225 ;
        RECT  10.47 17.645 10.54 17.78 ;
        RECT  10.8525 17.235 10.9225 17.37 ;
        RECT  10.31 14.4525 10.38 14.5875 ;
        RECT  11.015 14.4525 11.085 14.5875 ;
        RECT  10.6575 18.6925 10.7275 18.8275 ;
        RECT  10.6575 18.95 10.7275 19.09 ;
        RECT  10.83 15.005 10.9 19.09 ;
        RECT  10.495 14.205 10.565 19.09 ;
        RECT  11.015 14.205 11.085 19.09 ;
        RECT  11.2 14.205 11.27 19.09 ;
        RECT  11.535 14.205 11.605 17.75 ;
        RECT  11.3675 16.48 11.4375 18.49 ;
        RECT  11.535 15.005 11.605 19.09 ;
        RECT  11.72 14.205 11.79 19.09 ;
        RECT  11.54 19.04 11.6 19.09 ;
        RECT  11.2 19.03 11.27 19.09 ;
        RECT  11.3625 19.035 11.4325 19.09 ;
        RECT  11.3625 18.6925 11.4325 19.09 ;
        RECT  11.3675 16.345 11.4375 16.48 ;
        RECT  11.3675 18.4875 11.4375 18.6225 ;
        RECT  11.175 17.645 11.245 17.78 ;
        RECT  11.5575 17.235 11.6275 17.37 ;
        RECT  11.015 14.4525 11.085 14.5875 ;
        RECT  11.72 14.4525 11.79 14.5875 ;
        RECT  11.3625 18.6925 11.4325 18.8275 ;
        RECT  11.3625 18.95 11.4325 19.09 ;
        RECT  11.535 15.005 11.605 19.09 ;
        RECT  11.2 14.205 11.27 19.09 ;
        RECT  10.6625 10.03 10.7325 10.17 ;
        RECT  11.3675 10.03 11.4375 10.17 ;
        RECT  10.495 13.905 10.565 14.205 ;
        RECT  11.2 13.905 11.27 14.205 ;
        RECT  11.535 11.765 11.605 14.205 ;
        RECT  10.83 11.765 10.9 14.205 ;
        RECT  10.5525 10.1625 10.6875 10.2325 ;
        RECT  11.015 11.765 11.085 11.9 ;
        RECT  11.015 11.195 11.085 11.33 ;
        RECT  10.31 11.195 10.38 11.33 ;
        RECT  10.73 11.4 10.8 11.535 ;
        RECT  11.015 13.6925 11.085 13.8275 ;
        RECT  10.73 10.99 10.8 11.125 ;
        RECT  10.59 10.99 10.66 11.125 ;
        RECT  11.015 11.4 11.085 11.535 ;
        RECT  10.31 11.4 10.38 11.535 ;
        RECT  10.45 10.425 10.585 10.495 ;
        RECT  10.59 13.37 10.66 13.505 ;
        RECT  10.76 11.765 10.83 11.9 ;
        RECT  10.45 12.68 10.52 12.815 ;
        RECT  10.59 11.4 10.66 11.535 ;
        RECT  10.31 11.765 10.38 11.9 ;
        RECT  10.76 12.28 10.83 12.415 ;
        RECT  10.495 13.9025 10.565 14.0375 ;
        RECT  10.31 13.6925 10.38 13.8275 ;
        RECT  10.495 13.905 10.565 14.205 ;
        RECT  10.495 14.14 10.565 14.205 ;
        RECT  10.8325 14.145 10.8975 14.205 ;
        RECT  10.665 10.035 10.73 10.0975 ;
        RECT  11.015 10.03 11.085 14.205 ;
        RECT  10.31 10.03 10.38 14.205 ;
        RECT  10.83 11.765 10.9 14.205 ;
        RECT  10.54 10.1625 10.7325 10.2325 ;
        RECT  10.73 11.125 10.8 11.4 ;
        RECT  10.45 10.495 10.52 12.815 ;
        RECT  10.59 11.125 10.66 11.4 ;
        RECT  10.59 11.4 10.66 13.4975 ;
        RECT  10.6625 10.03 10.7325 10.17 ;
        RECT  10.6625 10.03 10.7325 10.17 ;
        RECT  10.83 11.765 10.9 14.205 ;
        RECT  10.495 13.905 10.565 14.205 ;
        RECT  11.2575 10.1625 11.3925 10.2325 ;
        RECT  11.72 11.765 11.79 11.9 ;
        RECT  11.72 11.195 11.79 11.33 ;
        RECT  11.015 11.195 11.085 11.33 ;
        RECT  11.435 11.4 11.505 11.535 ;
        RECT  11.72 13.6925 11.79 13.8275 ;
        RECT  11.435 10.99 11.505 11.125 ;
        RECT  11.295 10.99 11.365 11.125 ;
        RECT  11.72 11.4 11.79 11.535 ;
        RECT  11.015 11.4 11.085 11.535 ;
        RECT  11.155 10.425 11.29 10.495 ;
        RECT  11.295 13.37 11.365 13.505 ;
        RECT  11.465 11.765 11.535 11.9 ;
        RECT  11.155 12.68 11.225 12.815 ;
        RECT  11.295 11.4 11.365 11.535 ;
        RECT  11.015 11.765 11.085 11.9 ;
        RECT  11.465 12.28 11.535 12.415 ;
        RECT  11.2 13.9025 11.27 14.0375 ;
        RECT  11.015 13.6925 11.085 13.8275 ;
        RECT  11.2 13.905 11.27 14.205 ;
        RECT  11.2 14.14 11.27 14.205 ;
        RECT  11.5375 14.145 11.6025 14.205 ;
        RECT  11.37 10.035 11.435 10.0975 ;
        RECT  11.72 10.03 11.79 14.205 ;
        RECT  11.015 10.03 11.085 14.205 ;
        RECT  11.535 11.765 11.605 14.205 ;
        RECT  11.245 10.1625 11.4375 10.2325 ;
        RECT  11.435 11.125 11.505 11.4 ;
        RECT  11.155 10.495 11.225 12.815 ;
        RECT  11.295 11.125 11.365 11.4 ;
        RECT  11.295 11.4 11.365 13.4975 ;
        RECT  11.3675 10.03 11.4375 10.17 ;
        RECT  11.3675 10.03 11.4375 10.17 ;
        RECT  11.535 11.765 11.605 14.205 ;
        RECT  11.2 13.905 11.27 14.205 ;
        RECT  11.5225 9.3425 11.5925 10.03 ;
        RECT  11.3675 3.59 11.4375 3.735 ;
        RECT  10.6625 3.59 10.7325 3.735 ;
        RECT  10.31 3.59 10.38 10.03 ;
        RECT  11.015 3.59 11.085 10.03 ;
        RECT  11.72 3.59 11.79 10.03 ;
        RECT  10.5075 9.3425 10.5775 10.03 ;
        RECT  10.6625 9.76 10.7325 10.03 ;
        RECT  11.3675 9.76 11.4375 10.03 ;
        RECT  10.5075 9.2925 10.5775 9.4275 ;
        RECT  11.015 4.115 11.085 4.25 ;
        RECT  10.8725 8.1975 10.9425 8.3325 ;
        RECT  10.875 6.59 10.945 6.725 ;
        RECT  10.875 5.1925 10.945 5.3275 ;
        RECT  10.31 3.975 10.38 4.11 ;
        RECT  10.6625 3.59 10.7325 3.73 ;
        RECT  11.015 7.0525 11.085 7.1875 ;
        RECT  10.51 5.8575 10.58 5.9925 ;
        RECT  10.875 9.55 10.945 9.685 ;
        RECT  10.6975 9.04 10.7675 9.175 ;
        RECT  11.015 8.6275 11.085 8.7625 ;
        RECT  11.015 3.925 11.085 4.06 ;
        RECT  11.015 5.6675 11.085 5.8025 ;
        RECT  10.51 5.4675 10.58 5.6025 ;
        RECT  10.6975 5.4675 10.7675 5.6025 ;
        RECT  10.6975 6.08 10.7675 6.215 ;
        RECT  10.5075 8.4275 10.5775 8.5625 ;
        RECT  10.6975 8.4275 10.7675 8.5625 ;
        RECT  10.7325 9.76 10.875 9.83 ;
        RECT  10.6625 3.59 10.7325 3.735 ;
        RECT  10.7275 3.665 10.875 3.735 ;
        RECT  10.6625 9.76 10.7325 10.03 ;
        RECT  10.3125 9.5525 10.375 9.6125 ;
        RECT  10.31 3.59 10.38 10.03 ;
        RECT  10.665 9.965 10.73 10.025 ;
        RECT  10.875 9.55 10.945 9.83 ;
        RECT  10.875 3.665 10.945 5.3275 ;
        RECT  10.5075 9.3425 10.5775 10.03 ;
        RECT  10.875 6.725 10.945 8.3325 ;
        RECT  10.6975 8.4275 10.7675 9.145 ;
        RECT  10.51 5.4675 10.58 5.9925 ;
        RECT  10.5125 9.8925 10.575 9.9525 ;
        RECT  10.5075 8.4275 10.5775 9.3675 ;
        RECT  10.6625 3.595 10.73 3.66 ;
        RECT  11.015 3.59 11.085 10.03 ;
        RECT  10.6975 5.4675 10.7675 6.185 ;
        RECT  10.6625 3.59 10.7325 3.735 ;
        RECT  10.6625 9.76 10.7325 10.03 ;
        RECT  10.5075 9.3425 10.5775 10.03 ;
        RECT  10.31 3.59 10.38 10.03 ;
        RECT  11.015 3.59 11.085 10.03 ;
        RECT  11.5225 9.2925 11.5925 9.4275 ;
        RECT  11.015 4.115 11.085 4.25 ;
        RECT  11.1575 8.1975 11.2275 8.3325 ;
        RECT  11.155 6.59 11.225 6.725 ;
        RECT  11.155 5.1925 11.225 5.3275 ;
        RECT  11.72 3.975 11.79 4.11 ;
        RECT  11.3675 3.59 11.4375 3.73 ;
        RECT  11.015 7.0525 11.085 7.1875 ;
        RECT  11.52 5.8575 11.59 5.9925 ;
        RECT  11.155 9.55 11.225 9.685 ;
        RECT  11.3325 9.04 11.4025 9.175 ;
        RECT  11.015 8.6275 11.085 8.7625 ;
        RECT  11.015 3.925 11.085 4.06 ;
        RECT  11.015 5.6675 11.085 5.8025 ;
        RECT  11.52 5.4675 11.59 5.6025 ;
        RECT  11.3325 5.4675 11.4025 5.6025 ;
        RECT  11.3325 6.08 11.4025 6.215 ;
        RECT  11.5225 8.4275 11.5925 8.5625 ;
        RECT  11.3325 8.4275 11.4025 8.5625 ;
        RECT  11.225 9.76 11.3675 9.83 ;
        RECT  11.3675 3.59 11.4375 3.735 ;
        RECT  11.225 3.665 11.3725 3.735 ;
        RECT  11.3675 9.76 11.4375 10.03 ;
        RECT  11.725 9.5525 11.7875 9.6125 ;
        RECT  11.72 3.59 11.79 10.03 ;
        RECT  11.37 9.965 11.435 10.025 ;
        RECT  11.155 9.55 11.225 9.83 ;
        RECT  11.155 3.665 11.225 5.3275 ;
        RECT  11.5225 9.3425 11.5925 10.03 ;
        RECT  11.155 6.725 11.225 8.3325 ;
        RECT  11.3325 8.4275 11.4025 9.145 ;
        RECT  11.52 5.4675 11.59 5.9925 ;
        RECT  11.525 9.8925 11.5875 9.9525 ;
        RECT  11.5225 8.4275 11.5925 9.3675 ;
        RECT  11.37 3.595 11.4375 3.66 ;
        RECT  11.015 3.59 11.085 10.03 ;
        RECT  11.3325 5.4675 11.4025 6.185 ;
        RECT  11.3675 3.59 11.4375 3.735 ;
        RECT  11.3675 9.76 11.4375 10.03 ;
        RECT  11.5225 9.3425 11.5925 10.03 ;
        RECT  11.72 3.59 11.79 10.03 ;
        RECT  11.015 3.59 11.085 10.03 ;
        RECT  10.6625 0.615 10.7325 0.855 ;
        RECT  10.6625 3.24 10.7325 3.59 ;
        RECT  11.3675 3.24 11.4375 3.59 ;
        RECT  11.3675 0.615 11.4375 0.855 ;
        RECT  10.45 3.87 10.52 4.24 ;
        RECT  10.5225 4.505 10.7625 4.575 ;
        RECT  10.7625 4.505 10.8975 4.575 ;
        RECT  11.015 4.1625 11.085 4.22 ;
        RECT  11.015 3.59 11.085 6.565 ;
        RECT  10.695 5.4425 10.765 5.68 ;
        RECT  10.835 6.0125 10.905 6.395 ;
        RECT  10.4525 4.505 10.5225 6.0925 ;
        RECT  10.6625 3.745 10.7325 3.8075 ;
        RECT  10.6625 6.5075 10.7325 6.56 ;
        RECT  10.6625 6.325 10.7325 6.565 ;
        RECT  10.7325 6.325 10.835 6.395 ;
        RECT  10.6625 3.59 10.7325 3.94 ;
        RECT  10.45 3.87 10.6625 3.94 ;
        RECT  10.695 5.68 10.765 5.815 ;
        RECT  10.4875 5.9575 10.5575 6.0925 ;
        RECT  11.015 6.1475 11.085 6.2825 ;
        RECT  10.7625 6.0125 10.8975 6.0825 ;
        RECT  10.6625 3.7425 10.7325 3.8825 ;
        RECT  11.015 4.0875 11.085 4.2225 ;
        RECT  10.63 5.3725 10.765 5.4425 ;
        RECT  11.015 3.59 11.085 6.565 ;
        RECT  10.6625 6.325 10.7325 6.565 ;
        RECT  10.6625 3.59 10.7325 3.94 ;
        RECT  10.45 4.24 10.52 4.375 ;
        RECT  11.155 3.87 11.225 4.24 ;
        RECT  11.2275 4.505 11.4675 4.575 ;
        RECT  11.4675 4.505 11.6025 4.575 ;
        RECT  11.72 4.1625 11.79 4.22 ;
        RECT  11.72 3.59 11.79 6.565 ;
        RECT  11.4 5.4425 11.47 5.68 ;
        RECT  11.54 6.0125 11.61 6.395 ;
        RECT  11.1575 4.505 11.2275 6.0925 ;
        RECT  11.3675 3.745 11.4375 3.8075 ;
        RECT  11.3675 6.5075 11.4375 6.56 ;
        RECT  11.3675 6.325 11.4375 6.565 ;
        RECT  11.4375 6.325 11.54 6.395 ;
        RECT  11.3675 3.59 11.4375 3.94 ;
        RECT  11.155 3.87 11.3675 3.94 ;
        RECT  11.4 5.68 11.47 5.815 ;
        RECT  11.1925 5.9575 11.2625 6.0925 ;
        RECT  11.72 6.1475 11.79 6.2825 ;
        RECT  11.4675 6.0125 11.6025 6.0825 ;
        RECT  11.3675 3.7425 11.4375 3.8825 ;
        RECT  11.72 4.0875 11.79 4.2225 ;
        RECT  11.335 5.3725 11.47 5.4425 ;
        RECT  11.72 3.59 11.79 6.565 ;
        RECT  11.3675 6.325 11.4375 6.565 ;
        RECT  11.3675 3.59 11.4375 3.94 ;
        RECT  11.155 4.24 11.225 4.375 ;
        RECT  1.725 8.33 1.795 40.61 ;
        RECT  1.9 8.33 1.97 40.61 ;
        RECT  2.075 8.33 2.145 40.61 ;
        RECT  2.25 8.33 2.32 40.61 ;
        RECT  2.425 8.33 2.495 40.61 ;
        RECT  2.6 8.33 2.67 40.61 ;
        RECT  2.775 8.33 2.845 40.61 ;
        RECT  2.95 8.33 3.02 40.61 ;
        RECT  6.575 13.71 6.645 19.02 ;
        RECT  6.575 8.33 6.645 13.64 ;
        RECT  6.85 8.33 6.92 13.64 ;
        RECT  6.85 13.71 6.92 19.02 ;
        RECT  4.915 8.33 4.985 13.64 ;
        RECT  4.64 8.33 4.71 13.64 ;
        RECT  5.465 8.33 5.535 13.64 ;
        RECT  5.19 8.33 5.26 13.64 ;
        RECT  6.85 8.33 6.92 13.64 ;
        RECT  6.575 8.33 6.645 13.64 ;
        RECT  5.435 9.4075 5.57 9.4775 ;
        RECT  6.82 8.8075 6.955 8.8775 ;
        RECT  5.16 10.7525 5.295 10.8225 ;
        RECT  6.545 10.3325 6.68 10.4025 ;
        RECT  6.82 11.0775 6.955 11.1475 ;
        RECT  4.885 11.0775 5.02 11.1475 ;
        RECT  6.545 12.4225 6.68 12.4925 ;
        RECT  4.61 12.4225 4.745 12.4925 ;
        RECT  5.435 9.1675 5.57 9.2375 ;
        RECT  5.16 8.6375 5.295 8.7075 ;
        RECT  4.885 9.9725 5.02 10.0425 ;
        RECT  5.16 10.5025 5.295 10.5725 ;
        RECT  5.435 11.8575 5.57 11.9275 ;
        RECT  4.61 11.3275 4.745 11.3975 ;
        RECT  4.885 12.6625 5.02 12.7325 ;
        RECT  4.61 13.1925 4.745 13.2625 ;
        RECT  4.915 13.71 4.985 19.02 ;
        RECT  4.64 13.71 4.71 19.02 ;
        RECT  5.465 13.71 5.535 19.02 ;
        RECT  5.19 13.71 5.26 19.02 ;
        RECT  6.85 13.71 6.92 19.02 ;
        RECT  6.575 13.71 6.645 19.02 ;
        RECT  5.435 14.7875 5.57 14.8575 ;
        RECT  6.82 14.1875 6.955 14.2575 ;
        RECT  5.16 16.1325 5.295 16.2025 ;
        RECT  6.545 15.7125 6.68 15.7825 ;
        RECT  6.82 16.4575 6.955 16.5275 ;
        RECT  4.885 16.4575 5.02 16.5275 ;
        RECT  6.545 17.8025 6.68 17.8725 ;
        RECT  4.61 17.8025 4.745 17.8725 ;
        RECT  5.435 14.5475 5.57 14.6175 ;
        RECT  5.16 14.0175 5.295 14.0875 ;
        RECT  4.885 15.3525 5.02 15.4225 ;
        RECT  5.16 15.8825 5.295 15.9525 ;
        RECT  5.435 17.2375 5.57 17.3075 ;
        RECT  4.61 16.7075 4.745 16.7775 ;
        RECT  4.885 18.0425 5.02 18.1125 ;
        RECT  4.61 18.5725 4.745 18.6425 ;
        RECT  1.695 8.8775 1.83 8.9475 ;
        RECT  1.87 10.4025 2.005 10.4725 ;
        RECT  2.045 11.5675 2.18 11.6375 ;
        RECT  2.22 13.0925 2.355 13.1625 ;
        RECT  2.395 14.2575 2.53 14.3275 ;
        RECT  2.57 15.7825 2.705 15.8525 ;
        RECT  2.745 16.9475 2.88 17.0175 ;
        RECT  2.92 18.4725 3.055 18.5425 ;
        RECT  1.695 19.9975 1.83 20.0675 ;
        RECT  2.395 19.4675 2.53 19.5375 ;
        RECT  1.695 20.8025 1.83 20.8725 ;
        RECT  2.57 21.3325 2.705 21.4025 ;
        RECT  1.695 22.6875 1.83 22.7575 ;
        RECT  2.745 22.1575 2.88 22.2275 ;
        RECT  1.695 23.4925 1.83 23.5625 ;
        RECT  2.92 24.0225 3.055 24.0925 ;
        RECT  1.87 25.3775 2.005 25.4475 ;
        RECT  2.395 24.8475 2.53 24.9175 ;
        RECT  1.87 26.1825 2.005 26.2525 ;
        RECT  2.57 26.7125 2.705 26.7825 ;
        RECT  1.87 28.0675 2.005 28.1375 ;
        RECT  2.745 27.5375 2.88 27.6075 ;
        RECT  1.87 28.8725 2.005 28.9425 ;
        RECT  2.92 29.4025 3.055 29.4725 ;
        RECT  2.045 30.7575 2.18 30.8275 ;
        RECT  2.395 30.2275 2.53 30.2975 ;
        RECT  2.045 31.5625 2.18 31.6325 ;
        RECT  2.57 32.0925 2.705 32.1625 ;
        RECT  2.045 33.4475 2.18 33.5175 ;
        RECT  2.745 32.9175 2.88 32.9875 ;
        RECT  2.045 34.2525 2.18 34.3225 ;
        RECT  2.92 34.7825 3.055 34.8525 ;
        RECT  2.22 36.1375 2.355 36.2075 ;
        RECT  2.395 35.6075 2.53 35.6775 ;
        RECT  2.22 36.9425 2.355 37.0125 ;
        RECT  2.57 37.4725 2.705 37.5425 ;
        RECT  2.22 38.8275 2.355 38.8975 ;
        RECT  2.745 38.2975 2.88 38.3675 ;
        RECT  2.22 39.6325 2.355 39.7025 ;
        RECT  2.92 40.1625 3.055 40.2325 ;
        RECT  4.805 19.9975 5.45 20.0675 ;
        RECT  4.805 20.8025 5.45 20.8725 ;
        RECT  4.805 22.6875 5.45 22.7575 ;
        RECT  4.805 23.4925 5.45 23.5625 ;
        RECT  4.805 25.3775 5.45 25.4475 ;
        RECT  4.805 26.1825 5.45 26.2525 ;
        RECT  4.805 28.0675 5.45 28.1375 ;
        RECT  4.805 28.8725 5.45 28.9425 ;
        RECT  4.805 30.7575 5.45 30.8275 ;
        RECT  4.805 31.5625 5.45 31.6325 ;
        RECT  4.805 33.4475 5.45 33.5175 ;
        RECT  4.805 34.2525 5.45 34.3225 ;
        RECT  4.805 36.1375 5.45 36.2075 ;
        RECT  4.805 36.9425 5.45 37.0125 ;
        RECT  4.805 38.8275 5.45 38.8975 ;
        RECT  4.805 39.6325 5.45 39.7025 ;
        RECT  4.63 19.09 4.7 40.61 ;
        RECT  4.63 19.605 4.7 19.74 ;
        RECT  4.77 19.965 4.84 20.1 ;
        RECT  5.45 19.9975 5.585 20.0675 ;
        RECT  4.63 21.13 4.7 21.265 ;
        RECT  4.77 20.77 4.84 20.905 ;
        RECT  5.45 20.8025 5.585 20.8725 ;
        RECT  4.63 22.295 4.7 22.43 ;
        RECT  4.77 22.655 4.84 22.79 ;
        RECT  5.45 22.6875 5.585 22.7575 ;
        RECT  4.63 23.82 4.7 23.955 ;
        RECT  4.77 23.46 4.84 23.595 ;
        RECT  5.45 23.4925 5.585 23.5625 ;
        RECT  4.63 24.985 4.7 25.12 ;
        RECT  4.77 25.345 4.84 25.48 ;
        RECT  5.45 25.3775 5.585 25.4475 ;
        RECT  4.63 26.51 4.7 26.645 ;
        RECT  4.77 26.15 4.84 26.285 ;
        RECT  5.45 26.1825 5.585 26.2525 ;
        RECT  4.63 27.675 4.7 27.81 ;
        RECT  4.77 28.035 4.84 28.17 ;
        RECT  5.45 28.0675 5.585 28.1375 ;
        RECT  4.63 29.2 4.7 29.335 ;
        RECT  4.77 28.84 4.84 28.975 ;
        RECT  5.45 28.8725 5.585 28.9425 ;
        RECT  4.63 30.365 4.7 30.5 ;
        RECT  4.77 30.725 4.84 30.86 ;
        RECT  5.45 30.7575 5.585 30.8275 ;
        RECT  4.63 31.89 4.7 32.025 ;
        RECT  4.77 31.53 4.84 31.665 ;
        RECT  5.45 31.5625 5.585 31.6325 ;
        RECT  4.63 33.055 4.7 33.19 ;
        RECT  4.77 33.415 4.84 33.55 ;
        RECT  5.45 33.4475 5.585 33.5175 ;
        RECT  4.63 34.58 4.7 34.715 ;
        RECT  4.77 34.22 4.84 34.355 ;
        RECT  5.45 34.2525 5.585 34.3225 ;
        RECT  4.63 35.745 4.7 35.88 ;
        RECT  4.77 36.105 4.84 36.24 ;
        RECT  5.45 36.1375 5.585 36.2075 ;
        RECT  4.63 37.27 4.7 37.405 ;
        RECT  4.77 36.91 4.84 37.045 ;
        RECT  5.45 36.9425 5.585 37.0125 ;
        RECT  4.63 38.435 4.7 38.57 ;
        RECT  4.77 38.795 4.84 38.93 ;
        RECT  5.45 38.8275 5.585 38.8975 ;
        RECT  4.63 39.96 4.7 40.095 ;
        RECT  4.77 39.6 4.84 39.735 ;
        RECT  5.45 39.6325 5.585 39.7025 ;
        RECT  6.2325 6.6725 6.92 6.7425 ;
        RECT  0.48 5.4175 0.625 5.4875 ;
        RECT  6.2325 6.2775 6.92 6.3475 ;
        RECT  6.2325 5.2625 6.92 5.3325 ;
        RECT  0.48 6.8275 0.625 6.8975 ;
        RECT  0.48 7.5325 0.625 7.6025 ;
        RECT  0.48 6.1225 0.625 6.1925 ;
        RECT  0.48 7.885 6.92 7.955 ;
        RECT  0.48 7.18 6.92 7.25 ;
        RECT  0.48 6.475 6.92 6.545 ;
        RECT  0.48 5.77 6.92 5.84 ;
        RECT  0.48 5.065 6.92 5.135 ;
        RECT  6.2325 7.6875 6.92 7.7575 ;
        RECT  6.65 7.5325 6.92 7.6025 ;
        RECT  6.65 6.8275 6.92 6.8975 ;
        RECT  6.65 5.4175 6.92 5.4875 ;
        RECT  6.65 6.1225 6.92 6.1925 ;
        RECT  6.1825 7.6875 6.3175 7.7575 ;
        RECT  1.005 7.18 1.14 7.25 ;
        RECT  5.0875 7.3225 5.2225 7.3925 ;
        RECT  3.48 7.32 3.615 7.39 ;
        RECT  2.0825 7.32 2.2175 7.39 ;
        RECT  0.865 7.885 1.0 7.955 ;
        RECT  0.48 7.5325 0.62 7.6025 ;
        RECT  3.9425 7.18 4.0775 7.25 ;
        RECT  2.7475 7.685 2.8825 7.755 ;
        RECT  6.44 7.32 6.575 7.39 ;
        RECT  5.93 7.4975 6.065 7.5675 ;
        RECT  5.5175 7.18 5.6525 7.25 ;
        RECT  0.815 7.18 0.95 7.25 ;
        RECT  2.5575 7.18 2.6925 7.25 ;
        RECT  2.3575 7.685 2.4925 7.755 ;
        RECT  2.3575 7.4975 2.4925 7.5675 ;
        RECT  2.97 7.4975 3.105 7.5675 ;
        RECT  5.3175 7.6875 5.4525 7.7575 ;
        RECT  5.3175 7.4975 5.4525 7.5675 ;
        RECT  6.65 7.39 6.72 7.5325 ;
        RECT  0.48 7.5325 0.625 7.6025 ;
        RECT  0.555 7.39 0.625 7.5375 ;
        RECT  6.65 7.5325 6.92 7.6025 ;
        RECT  6.4425 7.89 6.5025 7.9525 ;
        RECT  0.48 7.885 6.92 7.955 ;
        RECT  6.855 7.535 6.915 7.6 ;
        RECT  6.44 7.32 6.72 7.39 ;
        RECT  0.555 7.32 2.2175 7.39 ;
        RECT  6.2325 7.6875 6.92 7.7575 ;
        RECT  3.615 7.32 5.2225 7.39 ;
        RECT  5.3175 7.4975 6.035 7.5675 ;
        RECT  2.3575 7.685 2.8825 7.755 ;
        RECT  6.7825 7.69 6.8425 7.7525 ;
        RECT  5.3175 7.6875 6.2575 7.7575 ;
        RECT  0.485 7.535 0.55 7.6025 ;
        RECT  0.48 7.18 6.92 7.25 ;
        RECT  2.3575 7.4975 3.075 7.5675 ;
        RECT  0.48 7.5325 0.625 7.6025 ;
        RECT  6.65 7.5325 6.92 7.6025 ;
        RECT  6.2325 7.6875 6.92 7.7575 ;
        RECT  0.48 7.885 6.92 7.955 ;
        RECT  0.48 7.18 6.92 7.25 ;
        RECT  6.1825 6.6725 6.3175 6.7425 ;
        RECT  1.005 7.18 1.14 7.25 ;
        RECT  5.0875 7.0375 5.2225 7.1075 ;
        RECT  3.48 7.04 3.615 7.11 ;
        RECT  2.0825 7.04 2.2175 7.11 ;
        RECT  0.865 6.475 1.0 6.545 ;
        RECT  0.48 6.8275 0.62 6.8975 ;
        RECT  3.9425 7.18 4.0775 7.25 ;
        RECT  2.7475 6.675 2.8825 6.745 ;
        RECT  6.44 7.04 6.575 7.11 ;
        RECT  5.93 6.8625 6.065 6.9325 ;
        RECT  5.5175 7.18 5.6525 7.25 ;
        RECT  0.815 7.18 0.95 7.25 ;
        RECT  2.5575 7.18 2.6925 7.25 ;
        RECT  2.3575 6.675 2.4925 6.745 ;
        RECT  2.3575 6.8625 2.4925 6.9325 ;
        RECT  2.97 6.8625 3.105 6.9325 ;
        RECT  5.3175 6.6725 5.4525 6.7425 ;
        RECT  5.3175 6.8625 5.4525 6.9325 ;
        RECT  6.65 6.8975 6.72 7.04 ;
        RECT  0.48 6.8275 0.625 6.8975 ;
        RECT  0.555 6.8925 0.625 7.04 ;
        RECT  6.65 6.8275 6.92 6.8975 ;
        RECT  6.4425 6.4775 6.5025 6.54 ;
        RECT  0.48 6.475 6.92 6.545 ;
        RECT  6.855 6.83 6.915 6.895 ;
        RECT  6.44 7.04 6.72 7.11 ;
        RECT  0.555 7.04 2.2175 7.11 ;
        RECT  6.2325 6.6725 6.92 6.7425 ;
        RECT  3.615 7.04 5.2225 7.11 ;
        RECT  5.3175 6.8625 6.035 6.9325 ;
        RECT  2.3575 6.675 2.8825 6.745 ;
        RECT  6.7825 6.6775 6.8425 6.74 ;
        RECT  5.3175 6.6725 6.2575 6.7425 ;
        RECT  0.485 6.8275 0.55 6.895 ;
        RECT  0.48 7.18 6.92 7.25 ;
        RECT  2.3575 6.8625 3.075 6.9325 ;
        RECT  0.48 6.8275 0.625 6.8975 ;
        RECT  6.65 6.8275 6.92 6.8975 ;
        RECT  6.2325 6.6725 6.92 6.7425 ;
        RECT  0.48 6.475 6.92 6.545 ;
        RECT  0.48 7.18 6.92 7.25 ;
        RECT  6.1825 6.2775 6.3175 6.3475 ;
        RECT  1.005 5.77 1.14 5.84 ;
        RECT  5.0875 5.9125 5.2225 5.9825 ;
        RECT  3.48 5.91 3.615 5.98 ;
        RECT  2.0825 5.91 2.2175 5.98 ;
        RECT  0.865 6.475 1.0 6.545 ;
        RECT  0.48 6.1225 0.62 6.1925 ;
        RECT  3.9425 5.77 4.0775 5.84 ;
        RECT  2.7475 6.275 2.8825 6.345 ;
        RECT  6.44 5.91 6.575 5.98 ;
        RECT  5.93 6.0875 6.065 6.1575 ;
        RECT  5.5175 5.77 5.6525 5.84 ;
        RECT  0.815 5.77 0.95 5.84 ;
        RECT  2.5575 5.77 2.6925 5.84 ;
        RECT  2.3575 6.275 2.4925 6.345 ;
        RECT  2.3575 6.0875 2.4925 6.1575 ;
        RECT  2.97 6.0875 3.105 6.1575 ;
        RECT  5.3175 6.2775 5.4525 6.3475 ;
        RECT  5.3175 6.0875 5.4525 6.1575 ;
        RECT  6.65 5.98 6.72 6.1225 ;
        RECT  0.48 6.1225 0.625 6.1925 ;
        RECT  0.555 5.98 0.625 6.1275 ;
        RECT  6.65 6.1225 6.92 6.1925 ;
        RECT  6.4425 6.48 6.5025 6.5425 ;
        RECT  0.48 6.475 6.92 6.545 ;
        RECT  6.855 6.125 6.915 6.19 ;
        RECT  6.44 5.91 6.72 5.98 ;
        RECT  0.555 5.91 2.2175 5.98 ;
        RECT  6.2325 6.2775 6.92 6.3475 ;
        RECT  3.615 5.91 5.2225 5.98 ;
        RECT  5.3175 6.0875 6.035 6.1575 ;
        RECT  2.3575 6.275 2.8825 6.345 ;
        RECT  6.7825 6.28 6.8425 6.3425 ;
        RECT  5.3175 6.2775 6.2575 6.3475 ;
        RECT  0.485 6.125 0.55 6.1925 ;
        RECT  0.48 5.77 6.92 5.84 ;
        RECT  2.3575 6.0875 3.075 6.1575 ;
        RECT  0.48 6.1225 0.625 6.1925 ;
        RECT  6.65 6.1225 6.92 6.1925 ;
        RECT  6.2325 6.2775 6.92 6.3475 ;
        RECT  0.48 6.475 6.92 6.545 ;
        RECT  0.48 5.77 6.92 5.84 ;
        RECT  6.1825 5.2625 6.3175 5.3325 ;
        RECT  1.005 5.77 1.14 5.84 ;
        RECT  5.0875 5.6275 5.2225 5.6975 ;
        RECT  3.48 5.63 3.615 5.7 ;
        RECT  2.0825 5.63 2.2175 5.7 ;
        RECT  0.865 5.065 1.0 5.135 ;
        RECT  0.48 5.4175 0.62 5.4875 ;
        RECT  3.9425 5.77 4.0775 5.84 ;
        RECT  2.7475 5.265 2.8825 5.335 ;
        RECT  6.44 5.63 6.575 5.7 ;
        RECT  5.93 5.4525 6.065 5.5225 ;
        RECT  5.5175 5.77 5.6525 5.84 ;
        RECT  0.815 5.77 0.95 5.84 ;
        RECT  2.5575 5.77 2.6925 5.84 ;
        RECT  2.3575 5.265 2.4925 5.335 ;
        RECT  2.3575 5.4525 2.4925 5.5225 ;
        RECT  2.97 5.4525 3.105 5.5225 ;
        RECT  5.3175 5.2625 5.4525 5.3325 ;
        RECT  5.3175 5.4525 5.4525 5.5225 ;
        RECT  6.65 5.4875 6.72 5.63 ;
        RECT  0.48 5.4175 0.625 5.4875 ;
        RECT  0.555 5.4825 0.625 5.63 ;
        RECT  6.65 5.4175 6.92 5.4875 ;
        RECT  6.4425 5.0675 6.5025 5.13 ;
        RECT  0.48 5.065 6.92 5.135 ;
        RECT  6.855 5.42 6.915 5.485 ;
        RECT  6.44 5.63 6.72 5.7 ;
        RECT  0.555 5.63 2.2175 5.7 ;
        RECT  6.2325 5.2625 6.92 5.3325 ;
        RECT  3.615 5.63 5.2225 5.7 ;
        RECT  5.3175 5.4525 6.035 5.5225 ;
        RECT  2.3575 5.265 2.8825 5.335 ;
        RECT  6.7825 5.2675 6.8425 5.33 ;
        RECT  5.3175 5.2625 6.2575 5.3325 ;
        RECT  0.485 5.4175 0.55 5.485 ;
        RECT  0.48 5.77 6.92 5.84 ;
        RECT  2.3575 5.4525 3.075 5.5225 ;
        RECT  0.48 5.4175 0.625 5.4875 ;
        RECT  6.65 5.4175 6.92 5.4875 ;
        RECT  6.2325 5.2625 6.92 5.3325 ;
        RECT  0.48 5.065 6.92 5.135 ;
        RECT  0.48 5.77 6.92 5.84 ;
        RECT  10.4525 0.44 10.5225 0.575 ;
        RECT  11.1575 0.44 11.2275 0.575 ;
        RECT  10.6625 0.0 10.7325 0.135 ;
        RECT  11.3675 0.0 11.4375 0.135 ;
        RECT  8.2525 19.055 8.3875 19.125 ;
        RECT  8.2525 21.745 8.3875 21.815 ;
        RECT  8.2525 24.435 8.3875 24.505 ;
        RECT  8.2525 27.125 8.3875 27.195 ;
        RECT  8.2525 29.815 8.3875 29.885 ;
        RECT  8.2525 32.505 8.3875 32.575 ;
        RECT  8.2525 35.195 8.3875 35.265 ;
        RECT  8.2525 37.885 8.3875 37.955 ;
        RECT  8.2525 40.575 8.3875 40.645 ;
        RECT  6.785 8.5 6.92 8.57 ;
        RECT  7.1625 8.5 7.2975 8.57 ;
        RECT  6.51 9.845 6.645 9.915 ;
        RECT  7.3675 9.845 7.5025 9.915 ;
        RECT  6.785 13.88 6.92 13.95 ;
        RECT  7.5725 13.88 7.7075 13.95 ;
        RECT  6.51 15.225 6.645 15.295 ;
        RECT  7.7775 15.225 7.9125 15.295 ;
        RECT  6.99 8.295 7.125 8.365 ;
        RECT  6.99 8.295 7.125 8.365 ;
        RECT  8.185 8.295 8.32 8.365 ;
        RECT  6.99 10.985 7.125 11.055 ;
        RECT  6.99 10.985 7.125 11.055 ;
        RECT  8.185 10.985 8.32 11.055 ;
        RECT  6.99 13.675 7.125 13.745 ;
        RECT  6.99 13.675 7.125 13.745 ;
        RECT  8.185 13.675 8.32 13.745 ;
        RECT  6.99 16.365 7.125 16.435 ;
        RECT  6.99 16.365 7.125 16.435 ;
        RECT  8.185 16.365 8.32 16.435 ;
        RECT  6.92 7.5325 7.055 7.6025 ;
        RECT  7.1625 7.5325 7.2975 7.6025 ;
        RECT  6.92 6.8275 7.055 6.8975 ;
        RECT  7.3675 6.8275 7.5025 6.8975 ;
        RECT  6.92 6.1225 7.055 6.1925 ;
        RECT  7.5725 6.1225 7.7075 6.1925 ;
        RECT  6.92 5.4175 7.055 5.4875 ;
        RECT  7.7775 5.4175 7.9125 5.4875 ;
        RECT  6.92 7.885 7.055 7.955 ;
        RECT  8.2525 7.885 8.3875 7.955 ;
        RECT  6.92 7.18 7.055 7.25 ;
        RECT  8.2525 7.18 8.3875 7.25 ;
        RECT  6.92 6.475 7.055 6.545 ;
        RECT  8.2525 6.475 8.3875 6.545 ;
        RECT  6.92 5.77 7.055 5.84 ;
        RECT  8.2525 5.77 8.3875 5.84 ;
        RECT  6.92 5.065 7.055 5.135 ;
        RECT  8.2525 5.065 8.3875 5.135 ;
        RECT  9.39 3.7925 9.525 3.8625 ;
        RECT  8.98 1.6075 9.115 1.6775 ;
        RECT  9.185 3.155 9.32 3.225 ;
        RECT  9.39 41.3925 9.525 41.4625 ;
        RECT  9.595 10.295 9.73 10.365 ;
        RECT  9.8 14.32 9.935 14.39 ;
        RECT  8.8075 8.09 8.8775 8.225 ;
        RECT  4.5975 40.78 4.7325 40.85 ;
        RECT  8.8075 40.78 8.8775 40.915 ;
        RECT  8.4675 3.025 8.6025 3.095 ;
        RECT  8.4675 14.45 8.6025 14.52 ;
        RECT  8.4675 3.9525 8.6025 4.0225 ;
        RECT  8.4675 11.2275 8.6025 11.2975 ;
        RECT  -4.175 27.025 -0.14 27.095 ;
        RECT  -4.175 27.23 -0.14 27.3 ;
        RECT  -4.175 27.435 -0.14 27.505 ;
        RECT  -4.175 27.845 -0.14 27.915 ;
        RECT  -3.8125 27.845 -3.6075 27.915 ;
        RECT  -3.6575 27.025 -3.4525 27.095 ;
        RECT  -2.7975 27.23 -2.5925 27.3 ;
        RECT  -2.4025 27.435 -2.1975 27.505 ;
        RECT  -4.01 26.82 -3.805 26.89 ;
        RECT  -3.305 26.82 -3.1 26.89 ;
        RECT  -2.6 26.82 -2.395 26.89 ;
        RECT  -1.895 26.82 -1.69 26.89 ;
        RECT  -0.7225 26.615 -0.5175 26.685 ;
        RECT  -0.7225 28.05 -0.5175 28.12 ;
        RECT  -1.725 19.4675 -1.655 26.65 ;
        RECT  -2.4125 26.615 -2.2075 26.685 ;
        RECT  -2.2725 27.025 -2.0675 27.095 ;
        RECT  -1.8875 28.05 -1.6825 28.12 ;
        RECT  -2.4175 27.845 -2.2125 27.915 ;
        RECT  -1.0225 28.05 -0.8175 28.12 ;
        RECT  -0.8875 27.845 -0.6825 27.915 ;
        RECT  -0.7525 27.23 -0.5475 27.3 ;
        RECT  -3.7125 28.05 -3.5075 28.12 ;
        RECT  -3.5775 27.435 -3.3725 27.505 ;
        RECT  -3.4425 27.23 -3.2375 27.3 ;
        RECT  -0.345 26.82 -0.14 26.89 ;
        RECT  -1.485 27.64 -1.28 27.71 ;
        RECT  -2.83 26.82 -2.625 26.89 ;
        RECT  -4.175 27.64 -3.97 27.71 ;
        RECT  -4.175 28.05 -0.14 28.12 ;
        RECT  -3.445 31.85 -0.14 31.92 ;
        RECT  -4.175 26.615 -0.14 26.685 ;
        RECT  -2.2325 30.385 -0.14 30.455 ;
        RECT  -4.175 27.64 -0.14 27.71 ;
        RECT  -4.175 26.82 -0.14 26.89 ;
        RECT  -2.28 30.61 -0.14 30.68 ;
        RECT  -2.445 29.41 -0.14 29.48 ;
        RECT  -2.8325 24.9825 -2.7625 25.67 ;
        RECT  -2.4375 24.9825 -2.3675 25.67 ;
        RECT  -2.9875 19.23 -2.9175 19.375 ;
        RECT  -3.6925 19.23 -3.6225 19.375 ;
        RECT  -2.2825 19.23 -2.2125 19.375 ;
        RECT  -4.045 19.23 -3.975 25.67 ;
        RECT  -3.34 19.23 -3.27 25.67 ;
        RECT  -2.635 19.23 -2.565 25.67 ;
        RECT  -1.93 19.23 -1.86 25.67 ;
        RECT  -3.8475 24.9825 -3.7775 25.67 ;
        RECT  -3.6925 25.4 -3.6225 25.67 ;
        RECT  -2.9875 25.4 -2.9175 25.67 ;
        RECT  -2.2825 25.4 -2.2125 25.67 ;
        RECT  -3.8475 24.9325 -3.7775 25.0675 ;
        RECT  -3.34 19.755 -3.27 19.89 ;
        RECT  -3.4825 23.8375 -3.4125 23.9725 ;
        RECT  -3.48 22.23 -3.41 22.365 ;
        RECT  -3.48 20.8325 -3.41 20.9675 ;
        RECT  -4.045 19.615 -3.975 19.75 ;
        RECT  -3.6925 19.23 -3.6225 19.37 ;
        RECT  -3.34 22.6925 -3.27 22.8275 ;
        RECT  -3.845 21.4975 -3.775 21.6325 ;
        RECT  -3.48 25.19 -3.41 25.325 ;
        RECT  -3.6575 24.68 -3.5875 24.815 ;
        RECT  -3.34 24.2675 -3.27 24.4025 ;
        RECT  -3.34 19.565 -3.27 19.7 ;
        RECT  -3.34 21.3075 -3.27 21.4425 ;
        RECT  -3.845 21.1075 -3.775 21.2425 ;
        RECT  -3.6575 21.1075 -3.5875 21.2425 ;
        RECT  -3.6575 21.72 -3.5875 21.855 ;
        RECT  -3.8475 24.0675 -3.7775 24.2025 ;
        RECT  -3.6575 24.0675 -3.5875 24.2025 ;
        RECT  -3.6225 25.4 -3.48 25.47 ;
        RECT  -3.6925 19.23 -3.6225 19.375 ;
        RECT  -3.6275 19.305 -3.48 19.375 ;
        RECT  -3.6925 25.4 -3.6225 25.67 ;
        RECT  -4.0425 25.1925 -3.98 25.2525 ;
        RECT  -4.045 19.23 -3.975 25.67 ;
        RECT  -3.69 25.605 -3.625 25.665 ;
        RECT  -3.48 25.19 -3.41 25.47 ;
        RECT  -3.48 19.305 -3.41 20.9675 ;
        RECT  -3.8475 24.9825 -3.7775 25.67 ;
        RECT  -3.48 22.365 -3.41 23.9725 ;
        RECT  -3.6575 24.0675 -3.5875 24.785 ;
        RECT  -3.845 21.1075 -3.775 21.6325 ;
        RECT  -3.8425 25.5325 -3.78 25.5925 ;
        RECT  -3.8475 24.0675 -3.7775 25.0075 ;
        RECT  -3.6925 19.235 -3.625 19.3 ;
        RECT  -3.34 19.23 -3.27 25.67 ;
        RECT  -3.6575 21.1075 -3.5875 21.825 ;
        RECT  -3.6925 19.23 -3.6225 19.375 ;
        RECT  -3.6925 25.4 -3.6225 25.67 ;
        RECT  -3.8475 24.9825 -3.7775 25.67 ;
        RECT  -4.045 19.23 -3.975 25.67 ;
        RECT  -3.34 19.23 -3.27 25.67 ;
        RECT  -2.8325 24.9325 -2.7625 25.0675 ;
        RECT  -3.34 19.755 -3.27 19.89 ;
        RECT  -3.1975 23.8375 -3.1275 23.9725 ;
        RECT  -3.2 22.23 -3.13 22.365 ;
        RECT  -3.2 20.8325 -3.13 20.9675 ;
        RECT  -2.635 19.615 -2.565 19.75 ;
        RECT  -2.9875 19.23 -2.9175 19.37 ;
        RECT  -3.34 22.6925 -3.27 22.8275 ;
        RECT  -2.835 21.4975 -2.765 21.6325 ;
        RECT  -3.2 25.19 -3.13 25.325 ;
        RECT  -3.0225 24.68 -2.9525 24.815 ;
        RECT  -3.34 24.2675 -3.27 24.4025 ;
        RECT  -3.34 19.565 -3.27 19.7 ;
        RECT  -3.34 21.3075 -3.27 21.4425 ;
        RECT  -2.835 21.1075 -2.765 21.2425 ;
        RECT  -3.0225 21.1075 -2.9525 21.2425 ;
        RECT  -3.0225 21.72 -2.9525 21.855 ;
        RECT  -2.8325 24.0675 -2.7625 24.2025 ;
        RECT  -3.0225 24.0675 -2.9525 24.2025 ;
        RECT  -3.13 25.4 -2.9875 25.47 ;
        RECT  -2.9875 19.23 -2.9175 19.375 ;
        RECT  -3.13 19.305 -2.9825 19.375 ;
        RECT  -2.9875 25.4 -2.9175 25.67 ;
        RECT  -2.63 25.1925 -2.5675 25.2525 ;
        RECT  -2.635 19.23 -2.565 25.67 ;
        RECT  -2.985 25.605 -2.92 25.665 ;
        RECT  -3.2 25.19 -3.13 25.47 ;
        RECT  -3.2 19.305 -3.13 20.9675 ;
        RECT  -2.8325 24.9825 -2.7625 25.67 ;
        RECT  -3.2 22.365 -3.13 23.9725 ;
        RECT  -3.0225 24.0675 -2.9525 24.785 ;
        RECT  -2.835 21.1075 -2.765 21.6325 ;
        RECT  -2.83 25.5325 -2.7675 25.5925 ;
        RECT  -2.8325 24.0675 -2.7625 25.0075 ;
        RECT  -2.985 19.235 -2.9175 19.3 ;
        RECT  -3.34 19.23 -3.27 25.67 ;
        RECT  -3.0225 21.1075 -2.9525 21.825 ;
        RECT  -2.9875 19.23 -2.9175 19.375 ;
        RECT  -2.9875 25.4 -2.9175 25.67 ;
        RECT  -2.8325 24.9825 -2.7625 25.67 ;
        RECT  -2.635 19.23 -2.565 25.67 ;
        RECT  -3.34 19.23 -3.27 25.67 ;
        RECT  -2.4375 24.9325 -2.3675 25.0675 ;
        RECT  -1.93 19.755 -1.86 19.89 ;
        RECT  -2.0725 23.8375 -2.0025 23.9725 ;
        RECT  -2.07 22.23 -2.0 22.365 ;
        RECT  -2.07 20.8325 -2.0 20.9675 ;
        RECT  -2.635 19.615 -2.565 19.75 ;
        RECT  -2.2825 19.23 -2.2125 19.37 ;
        RECT  -1.93 22.6925 -1.86 22.8275 ;
        RECT  -2.435 21.4975 -2.365 21.6325 ;
        RECT  -2.07 25.19 -2.0 25.325 ;
        RECT  -2.2475 24.68 -2.1775 24.815 ;
        RECT  -1.93 24.2675 -1.86 24.4025 ;
        RECT  -1.93 19.565 -1.86 19.7 ;
        RECT  -1.93 21.3075 -1.86 21.4425 ;
        RECT  -2.435 21.1075 -2.365 21.2425 ;
        RECT  -2.2475 21.1075 -2.1775 21.2425 ;
        RECT  -2.2475 21.72 -2.1775 21.855 ;
        RECT  -2.4375 24.0675 -2.3675 24.2025 ;
        RECT  -2.2475 24.0675 -2.1775 24.2025 ;
        RECT  -2.2125 25.4 -2.07 25.47 ;
        RECT  -2.2825 19.23 -2.2125 19.375 ;
        RECT  -2.2175 19.305 -2.07 19.375 ;
        RECT  -2.2825 25.4 -2.2125 25.67 ;
        RECT  -2.6325 25.1925 -2.57 25.2525 ;
        RECT  -2.635 19.23 -2.565 25.67 ;
        RECT  -2.28 25.605 -2.215 25.665 ;
        RECT  -2.07 25.19 -2.0 25.47 ;
        RECT  -2.07 19.305 -2.0 20.9675 ;
        RECT  -2.4375 24.9825 -2.3675 25.67 ;
        RECT  -2.07 22.365 -2.0 23.9725 ;
        RECT  -2.2475 24.0675 -2.1775 24.785 ;
        RECT  -2.435 21.1075 -2.365 21.6325 ;
        RECT  -2.4325 25.5325 -2.37 25.5925 ;
        RECT  -2.4375 24.0675 -2.3675 25.0075 ;
        RECT  -2.2825 19.235 -2.215 19.3 ;
        RECT  -1.93 19.23 -1.86 25.67 ;
        RECT  -2.2475 21.1075 -2.1775 21.825 ;
        RECT  -2.2825 19.23 -2.2125 19.375 ;
        RECT  -2.2825 25.4 -2.2125 25.67 ;
        RECT  -2.4375 24.9825 -2.3675 25.67 ;
        RECT  -2.635 19.23 -2.565 25.67 ;
        RECT  -1.93 19.23 -1.86 25.67 ;
        RECT  -1.2725 28.88 -1.2025 29.33 ;
        RECT  -1.3375 28.88 -1.2025 28.95 ;
        RECT  -1.3375 29.26 -1.2025 29.33 ;
        RECT  -2.4125 29.105 -1.8825 29.175 ;
        RECT  -2.0175 29.105 -1.8825 29.175 ;
        RECT  -2.5175 29.0725 -2.4475 29.2075 ;
        RECT  -3.9625 29.44 -3.8925 29.89 ;
        RECT  -4.0275 29.44 -3.8925 29.51 ;
        RECT  -4.0275 29.82 -3.8925 29.89 ;
        RECT  -3.8475 27.8125 -3.7775 27.9475 ;
        RECT  -3.8475 25.67 -3.7775 25.805 ;
        RECT  -3.8475 25.67 -3.7775 25.805 ;
        RECT  -3.6925 26.9925 -3.6225 27.1275 ;
        RECT  -3.6925 25.67 -3.6225 25.805 ;
        RECT  -3.6925 25.67 -3.6225 25.805 ;
        RECT  -2.8325 27.1975 -2.7625 27.3325 ;
        RECT  -2.8325 25.67 -2.7625 25.805 ;
        RECT  -2.8325 25.67 -2.7625 25.805 ;
        RECT  -2.4375 27.4025 -2.3675 27.5375 ;
        RECT  -2.4375 25.67 -2.3675 25.805 ;
        RECT  -2.4375 25.67 -2.3675 25.805 ;
        RECT  -4.045 26.7875 -3.975 26.9225 ;
        RECT  -4.045 25.67 -3.975 25.805 ;
        RECT  -3.34 26.7875 -3.27 26.9225 ;
        RECT  -3.34 25.67 -3.27 25.805 ;
        RECT  -2.635 26.7875 -2.565 26.9225 ;
        RECT  -2.635 25.67 -2.565 25.805 ;
        RECT  -1.93 26.7875 -1.86 26.9225 ;
        RECT  -1.93 25.67 -1.86 25.805 ;
        RECT  -2.865 32.495 -2.795 37.295 ;
        RECT  -2.865 33.055 -2.795 33.26 ;
        RECT  -2.865 33.26 -2.795 37.395 ;
        RECT  -3.275 37.19 -3.205 37.395 ;
        RECT  -3.0375 32.6625 -2.9675 33.26 ;
        RECT  -3.46 32.6625 -3.39 32.9425 ;
        RECT  -0.76 34.175 -0.69 34.4125 ;
        RECT  -0.76 33.65 -0.69 33.8525 ;
        RECT  -2.28 33.615 -2.21 33.65 ;
        RECT  -2.28 33.9375 -2.21 34.175 ;
        RECT  -0.76 34.6 -0.69 34.735 ;
        RECT  -0.76 34.04 -0.69 34.175 ;
        RECT  -2.28 33.615 -2.21 33.75 ;
        RECT  -2.28 34.175 -2.21 34.31 ;
        RECT  -0.76 34.2775 -0.69 34.4125 ;
        RECT  -0.76 33.7175 -0.69 33.8525 ;
        RECT  -0.76 33.5825 -0.69 33.7175 ;
        RECT  -2.28 33.5825 -2.21 33.7175 ;
        RECT  -2.28 33.9375 -2.21 34.0725 ;
        RECT  -3.275 34.6625 -3.205 34.7975 ;
        RECT  -3.98 35.1375 -3.91 35.2725 ;
        RECT  -3.275 35.1375 -3.205 35.2725 ;
        RECT  -3.7275 34.6575 -3.6575 34.7925 ;
        RECT  -3.5275 34.6625 -3.4575 34.7975 ;
        RECT  -4.0125 34.365 -3.8775 34.435 ;
        RECT  -3.3075 34.365 -3.1725 34.435 ;
        RECT  -3.795 34.3675 -3.725 34.4325 ;
        RECT  -3.46 34.3675 -3.39 34.4325 ;
        RECT  -3.275 34.365 -3.205 34.435 ;
        RECT  -3.46 34.3 -3.39 35.8575 ;
        RECT  -3.795 34.3 -3.725 35.865 ;
        RECT  -3.98 34.3 -3.91 35.8675 ;
        RECT  -3.275 34.3 -3.205 35.845 ;
        RECT  -3.46 34.3 -3.39 35.8575 ;
        RECT  -3.275 34.3 -3.205 35.845 ;
        RECT  -3.795 34.3 -3.725 35.865 ;
        RECT  -3.46 31.61 -3.39 34.5 ;
        RECT  -3.275 31.61 -3.205 34.5 ;
        RECT  -3.98 31.61 -3.91 34.5 ;
        RECT  -3.795 31.61 -3.725 34.5 ;
        RECT  -3.98 33.515 -3.91 33.65 ;
        RECT  -3.98 33.515 -3.91 33.65 ;
        RECT  -3.98 33.515 -3.91 33.65 ;
        RECT  -3.98 33.515 -3.91 33.65 ;
        RECT  -3.98 33.515 -3.91 33.65 ;
        RECT  -3.98 33.515 -3.91 33.65 ;
        RECT  -3.3075 34.365 -3.1725 34.435 ;
        RECT  -4.0125 34.365 -3.8775 34.435 ;
        RECT  -3.98 33.515 -3.91 33.65 ;
        RECT  -3.98 33.515 -3.91 33.65 ;
        RECT  -3.98 33.515 -3.91 33.65 ;
        RECT  -3.98 33.515 -3.91 33.65 ;
        RECT  -3.98 33.515 -3.91 33.65 ;
        RECT  -3.98 33.515 -3.91 33.65 ;
        RECT  -3.98 33.515 -3.91 33.65 ;
        RECT  -3.98 33.515 -3.91 33.65 ;
        RECT  -3.53 34.0075 -3.46 34.1425 ;
        RECT  -3.275 33.515 -3.205 33.65 ;
        RECT  -3.275 33.515 -3.205 33.65 ;
        RECT  -3.275 33.515 -3.205 33.65 ;
        RECT  -3.275 33.515 -3.205 33.65 ;
        RECT  -3.275 33.515 -3.205 33.65 ;
        RECT  -3.275 33.515 -3.205 33.65 ;
        RECT  -3.98 33.515 -3.91 33.65 ;
        RECT  -3.98 33.515 -3.91 33.65 ;
        RECT  -3.98 33.515 -3.91 33.65 ;
        RECT  -3.98 33.515 -3.91 33.65 ;
        RECT  -3.725 34.0075 -3.655 34.1425 ;
        RECT  -4.0125 34.365 -3.8775 34.435 ;
        RECT  -4.0125 34.365 -3.8775 34.435 ;
        RECT  -4.0125 34.365 -3.8775 34.435 ;
        RECT  -3.98 33.515 -3.91 33.65 ;
        RECT  -3.98 33.515 -3.91 33.65 ;
        RECT  -3.98 33.515 -3.91 33.65 ;
        RECT  -3.98 33.515 -3.91 33.65 ;
        RECT  -3.98 33.515 -3.91 33.65 ;
        RECT  -3.98 33.515 -3.91 33.65 ;
        RECT  -3.3075 34.365 -3.1725 34.435 ;
        RECT  -3.98 33.0225 -3.91 34.4325 ;
        RECT  -3.27 34.3725 -3.21 34.43 ;
        RECT  -3.4525 34.3725 -3.3975 34.425 ;
        RECT  -3.79 34.3725 -3.7325 34.4325 ;
        RECT  -3.975 34.3675 -3.915 34.425 ;
        RECT  -3.795 32.955 -3.725 34.5 ;
        RECT  -3.46 32.955 -3.39 34.5 ;
        RECT  -3.275 32.955 -3.205 34.5 ;
        RECT  -3.98 32.955 -3.91 34.5 ;
        RECT  -3.46 32.955 -3.39 34.5 ;
        RECT  -3.275 32.955 -3.205 34.5 ;
        RECT  -3.98 32.955 -3.91 34.5 ;
        RECT  -3.795 32.955 -3.725 34.5 ;
        RECT  -3.98 32.46 -3.91 32.595 ;
        RECT  -3.98 32.46 -3.91 32.595 ;
        RECT  -3.98 32.46 -3.91 32.595 ;
        RECT  -3.98 32.46 -3.91 32.595 ;
        RECT  -3.98 32.46 -3.91 32.595 ;
        RECT  -3.98 32.46 -3.91 32.595 ;
        RECT  -3.3075 31.675 -3.1725 31.745 ;
        RECT  -4.0125 31.675 -3.8775 31.745 ;
        RECT  -3.98 32.46 -3.91 32.595 ;
        RECT  -3.98 32.46 -3.91 32.595 ;
        RECT  -3.98 32.46 -3.91 32.595 ;
        RECT  -3.98 32.46 -3.91 32.595 ;
        RECT  -3.98 32.46 -3.91 32.595 ;
        RECT  -3.98 32.46 -3.91 32.595 ;
        RECT  -3.98 32.46 -3.91 32.595 ;
        RECT  -3.98 32.46 -3.91 32.595 ;
        RECT  -3.53 31.9675 -3.46 32.1025 ;
        RECT  -3.275 32.46 -3.205 32.595 ;
        RECT  -3.275 32.46 -3.205 32.595 ;
        RECT  -3.275 32.46 -3.205 32.595 ;
        RECT  -3.275 32.46 -3.205 32.595 ;
        RECT  -3.275 32.46 -3.205 32.595 ;
        RECT  -3.275 32.46 -3.205 32.595 ;
        RECT  -3.98 32.46 -3.91 32.595 ;
        RECT  -3.98 32.46 -3.91 32.595 ;
        RECT  -3.98 32.46 -3.91 32.595 ;
        RECT  -3.98 32.46 -3.91 32.595 ;
        RECT  -3.725 31.9675 -3.655 32.1025 ;
        RECT  -4.0125 31.675 -3.8775 31.745 ;
        RECT  -4.0125 31.675 -3.8775 31.745 ;
        RECT  -4.0125 31.675 -3.8775 31.745 ;
        RECT  -3.98 32.46 -3.91 32.595 ;
        RECT  -3.98 32.46 -3.91 32.595 ;
        RECT  -3.98 32.46 -3.91 32.595 ;
        RECT  -3.98 32.46 -3.91 32.595 ;
        RECT  -3.98 32.46 -3.91 32.595 ;
        RECT  -3.98 32.46 -3.91 32.595 ;
        RECT  -3.3075 31.675 -3.1725 31.745 ;
        RECT  -3.98 31.6775 -3.91 33.0875 ;
        RECT  -3.27 31.68 -3.21 31.7375 ;
        RECT  -3.4525 31.685 -3.3975 31.7375 ;
        RECT  -3.79 31.6775 -3.7325 31.7375 ;
        RECT  -3.975 31.685 -3.915 31.7425 ;
        RECT  -3.795 31.61 -3.725 33.155 ;
        RECT  -3.46 31.61 -3.39 33.155 ;
        RECT  -3.275 31.61 -3.205 33.155 ;
        RECT  -3.98 31.61 -3.91 33.155 ;
        RECT  -3.46 31.61 -3.39 33.155 ;
        RECT  -3.275 31.61 -3.205 33.155 ;
        RECT  -3.98 31.61 -3.91 33.155 ;
        RECT  -3.795 31.61 -3.725 33.155 ;
        RECT  -2.865 34.3725 -2.795 34.5075 ;
        RECT  -2.865 36.7825 -2.795 36.9175 ;
        RECT  -2.865 34.6 -2.795 34.735 ;
        RECT  -2.865 32.225 -2.795 32.36 ;
        RECT  -2.8975 37.29 -2.7625 37.36 ;
        RECT  -3.3075 37.29 -3.1725 37.36 ;
        RECT  -3.07 33.155 -2.935 33.225 ;
        RECT  -3.07 32.5575 -2.935 32.6275 ;
        RECT  -3.4925 32.5575 -3.3575 32.6275 ;
        RECT  -0.7575 26.5825 -0.6875 26.7175 ;
        RECT  -0.7575 28.0175 -0.6875 28.1525 ;
        RECT  -0.7575 23.0 -0.6875 23.135 ;
        RECT  -0.7575 23.0 -0.6875 23.135 ;
        RECT  -1.725 19.4 -1.655 19.535 ;
        RECT  -2.4475 26.5825 -2.3775 26.7175 ;
        RECT  -2.3075 26.9925 -2.2375 27.1275 ;
        RECT  -1.9225 28.0175 -1.8525 28.1525 ;
        RECT  -1.9225 29.635 -1.8525 29.77 ;
        RECT  -1.9225 29.635 -1.8525 29.77 ;
        RECT  -2.4525 27.8125 -2.3825 27.9475 ;
        RECT  -2.4525 29.635 -2.3825 29.77 ;
        RECT  -2.4525 29.635 -2.3825 29.77 ;
        RECT  -1.0575 28.0175 -0.9875 28.1525 ;
        RECT  -0.9225 27.8125 -0.8525 27.9475 ;
        RECT  -0.7875 27.1975 -0.7175 27.3325 ;
        RECT  -3.7475 28.0175 -3.6775 28.1525 ;
        RECT  -3.6125 27.4025 -3.5425 27.5375 ;
        RECT  -3.4775 27.1975 -3.4075 27.3325 ;
        RECT  -2.4475 29.41 -2.3775 29.545 ;
        RECT  -2.235 30.385 -2.165 30.52 ;
        RECT  -3.4475 31.85 -3.3775 31.985 ;
        RECT  -2.2825 30.61 -2.2125 30.745 ;
        RECT  -0.175 26.7875 -0.105 26.9225 ;
        RECT  -1.52 27.6075 -1.45 27.7425 ;
        RECT  -2.865 26.7875 -2.795 26.9225 ;
        RECT  -4.21 27.6075 -4.14 27.7425 ;
        RECT  9.8 30.61 9.935 30.68 ;
        RECT  -0.275 30.61 -0.14 30.68 ;
        RECT  9.595 31.85 9.73 31.92 ;
        RECT  -0.275 31.85 -0.14 31.92 ;
        RECT  9.185 29.41 9.32 29.48 ;
        RECT  -0.275 29.41 -0.14 29.48 ;
        RECT  8.98 30.385 9.115 30.455 ;
        RECT  -0.275 30.385 -0.14 30.455 ;
        RECT  9.39 28.05 9.525 28.12 ;
        RECT  -0.275 28.05 -0.14 28.12 ;
        RECT  8.775 26.615 8.91 26.685 ;
        RECT  -0.275 26.615 -0.14 26.685 ;
        RECT  0.1075 27.64 0.2425 27.71 ;
        RECT  8.36 26.82 8.495 26.89 ;
        RECT  -0.275 26.82 -0.14 26.89 ;
        LAYER  via2 ;
        RECT  10.6575 18.985 10.7275 19.055 ;
        RECT  11.3625 18.985 11.4325 19.055 ;
        RECT  10.6625 3.625 10.7325 3.695 ;
        RECT  11.3675 3.625 11.4375 3.695 ;
        RECT  10.6625 3.7775 10.7325 3.8475 ;
        RECT  11.3675 3.7775 11.4375 3.8475 ;
        RECT  0.515 7.5325 0.585 7.6025 ;
        RECT  0.515 6.8275 0.585 6.8975 ;
        RECT  0.515 6.1225 0.585 6.1925 ;
        RECT  0.515 5.4175 0.585 5.4875 ;
        RECT  10.455 0.475 10.52 0.54 ;
        RECT  11.16 0.475 11.225 0.54 ;
        RECT  10.665 0.035 10.73 0.1 ;
        RECT  11.37 0.035 11.435 0.1 ;
        RECT  7.025 8.2975 7.09 8.3625 ;
        RECT  8.22 8.2975 8.285 8.3625 ;
        RECT  7.025 10.9875 7.09 11.0525 ;
        RECT  8.22 10.9875 8.285 11.0525 ;
        RECT  7.025 13.6775 7.09 13.7425 ;
        RECT  8.22 13.6775 8.285 13.7425 ;
        RECT  7.025 16.3675 7.09 16.4325 ;
        RECT  8.22 16.3675 8.285 16.4325 ;
        RECT  -3.6925 19.265 -3.6225 19.335 ;
        RECT  -2.9875 19.265 -2.9175 19.335 ;
        RECT  -2.2825 19.265 -2.2125 19.335 ;
        RECT  -3.845 27.8475 -3.78 27.9125 ;
        RECT  -3.845 25.705 -3.78 25.77 ;
        RECT  -3.69 27.0275 -3.625 27.0925 ;
        RECT  -3.69 25.705 -3.625 25.77 ;
        RECT  -2.83 27.2325 -2.765 27.2975 ;
        RECT  -2.83 25.705 -2.765 25.77 ;
        RECT  -2.435 27.4375 -2.37 27.5025 ;
        RECT  -2.435 25.705 -2.37 25.77 ;
        RECT  -4.0425 26.8225 -3.9775 26.8875 ;
        RECT  -4.0425 25.705 -3.9775 25.77 ;
        RECT  -3.3375 26.8225 -3.2725 26.8875 ;
        RECT  -3.3375 25.705 -3.2725 25.77 ;
        RECT  -2.6325 26.8225 -2.5675 26.8875 ;
        RECT  -2.6325 25.705 -2.5675 25.77 ;
        RECT  -1.9275 26.8225 -1.8625 26.8875 ;
        RECT  -1.9275 25.705 -1.8625 25.77 ;
        RECT  -0.7575 33.6175 -0.6925 33.6825 ;
        RECT  -2.2775 33.6175 -2.2125 33.6825 ;
        RECT  -0.755 28.0525 -0.69 28.1175 ;
        RECT  -0.755 23.035 -0.69 23.1 ;
        RECT  -1.92 28.0525 -1.855 28.1175 ;
        RECT  -1.92 29.67 -1.855 29.735 ;
        RECT  -2.45 27.8475 -2.385 27.9125 ;
        RECT  -2.45 29.67 -2.385 29.735 ;
        RECT  9.835 30.6125 9.9 30.6775 ;
        RECT  -0.24 30.6125 -0.175 30.6775 ;
        RECT  9.63 31.8525 9.695 31.9175 ;
        RECT  -0.24 31.8525 -0.175 31.9175 ;
        RECT  9.22 29.4125 9.285 29.4775 ;
        RECT  -0.24 29.4125 -0.175 29.4775 ;
        RECT  9.015 30.3875 9.08 30.4525 ;
        RECT  -0.24 30.3875 -0.175 30.4525 ;
        RECT  9.425 28.0525 9.49 28.1175 ;
        RECT  -0.24 28.0525 -0.175 28.1175 ;
        RECT  8.81 26.6175 8.875 26.6825 ;
        RECT  -0.24 26.6175 -0.175 26.6825 ;
        RECT  8.395 26.8225 8.46 26.8875 ;
        RECT  -0.24 26.8225 -0.175 26.8875 ;
        LAYER  metal3 ;
        RECT  -0.14 30.61 9.8675 30.68 ;
        RECT  -0.14 31.85 9.6625 31.92 ;
        RECT  -0.14 29.41 9.2525 29.48 ;
        RECT  -0.14 30.385 9.0475 30.455 ;
        RECT  -0.14 28.05 9.4575 28.12 ;
        RECT  -0.14 26.615 8.8425 26.685 ;
        RECT  -0.14 26.82 8.4275 26.89 ;
        RECT  -2.2825 19.23 -2.2125 19.37 ;
        RECT  0.0 5.4175 0.48 5.4875 ;
        RECT  -2.9875 19.23 -2.9175 19.37 ;
        RECT  0.0 6.8275 0.48 6.8975 ;
        RECT  0.0 7.5325 0.48 7.6025 ;
        RECT  0.0 6.1225 0.48 6.1925 ;
        RECT  -3.6925 19.23 -3.6225 19.37 ;
        RECT  10.4525 18.985 10.5225 19.055 ;
        RECT  10.4525 0.475 10.5225 19.02 ;
        RECT  10.4875 18.985 10.6575 19.055 ;
        RECT  11.1575 18.985 11.2275 19.055 ;
        RECT  11.1575 0.475 11.2275 19.02 ;
        RECT  11.1925 18.985 11.3625 19.055 ;
        RECT  10.6625 0.0 10.7325 3.59 ;
        RECT  11.3675 0.0 11.4375 3.59 ;
        RECT  7.0575 8.295 8.2525 8.365 ;
        RECT  7.0575 10.985 8.2525 11.055 ;
        RECT  7.0575 13.675 8.2525 13.745 ;
        RECT  7.0575 16.365 8.2525 16.435 ;
        RECT  0.0 5.4175 0.48 5.4875 ;
        RECT  0.0 6.8275 0.48 6.8975 ;
        RECT  0.0 7.5325 0.48 7.6025 ;
        RECT  0.0 6.1225 0.48 6.1925 ;
        RECT  10.6575 18.95 10.7275 19.09 ;
        RECT  11.3625 18.95 11.4325 19.09 ;
        RECT  10.6575 18.95 10.7275 19.09 ;
        RECT  10.6575 18.95 10.7275 19.09 ;
        RECT  11.3625 18.95 11.4325 19.09 ;
        RECT  11.3625 18.95 11.4325 19.09 ;
        RECT  11.3675 3.59 11.4375 3.73 ;
        RECT  10.6625 3.59 10.7325 3.73 ;
        RECT  10.6625 3.59 10.7325 3.73 ;
        RECT  10.6625 3.59 10.7325 3.73 ;
        RECT  11.3675 3.59 11.4375 3.73 ;
        RECT  11.3675 3.59 11.4375 3.73 ;
        RECT  10.6625 3.7425 10.7325 3.8825 ;
        RECT  11.3675 3.7425 11.4375 3.8825 ;
        RECT  0.48 5.4175 0.62 5.4875 ;
        RECT  0.48 6.8275 0.62 6.8975 ;
        RECT  0.48 7.5325 0.62 7.6025 ;
        RECT  0.48 6.1225 0.62 6.1925 ;
        RECT  0.48 7.5325 0.62 7.6025 ;
        RECT  0.48 7.5325 0.62 7.6025 ;
        RECT  0.48 6.8275 0.62 6.8975 ;
        RECT  0.48 6.8275 0.62 6.8975 ;
        RECT  0.48 6.1225 0.62 6.1925 ;
        RECT  0.48 6.1225 0.62 6.1925 ;
        RECT  0.48 5.4175 0.62 5.4875 ;
        RECT  0.48 5.4175 0.62 5.4875 ;
        RECT  10.4525 0.44 10.5225 0.575 ;
        RECT  11.1575 0.44 11.2275 0.575 ;
        RECT  10.6625 0.0 10.7325 0.135 ;
        RECT  11.3675 0.0 11.4375 0.135 ;
        RECT  6.99 8.295 7.125 8.365 ;
        RECT  8.185 8.295 8.32 8.365 ;
        RECT  6.99 10.985 7.125 11.055 ;
        RECT  8.185 10.985 8.32 11.055 ;
        RECT  6.99 13.675 7.125 13.745 ;
        RECT  8.185 13.675 8.32 13.745 ;
        RECT  6.99 16.365 7.125 16.435 ;
        RECT  8.185 16.365 8.32 16.435 ;
        RECT  -3.8475 25.67 -3.7775 27.88 ;
        RECT  -3.6925 25.67 -3.6225 27.06 ;
        RECT  -2.8325 25.67 -2.7625 27.265 ;
        RECT  -2.4375 25.67 -2.3675 27.47 ;
        RECT  -4.045 25.67 -3.975 26.855 ;
        RECT  -3.34 25.67 -3.27 26.855 ;
        RECT  -2.635 25.67 -2.565 26.855 ;
        RECT  -1.93 25.67 -1.86 26.855 ;
        RECT  -0.7575 23.0 -0.6875 28.085 ;
        RECT  -1.9225 28.085 -1.8525 29.635 ;
        RECT  -2.4525 27.88 -2.3825 29.635 ;
        RECT  -2.2825 19.23 -2.2125 19.37 ;
        RECT  -2.9875 19.23 -2.9175 19.37 ;
        RECT  -3.6925 19.23 -3.6225 19.37 ;
        RECT  -2.9875 19.23 -2.9175 19.37 ;
        RECT  -3.6925 19.23 -3.6225 19.37 ;
        RECT  -2.2825 19.23 -2.2125 19.37 ;
        RECT  -3.6925 19.23 -3.6225 19.37 ;
        RECT  -3.6925 19.23 -3.6225 19.37 ;
        RECT  -2.9875 19.23 -2.9175 19.37 ;
        RECT  -2.9875 19.23 -2.9175 19.37 ;
        RECT  -2.2825 19.23 -2.2125 19.37 ;
        RECT  -2.2825 19.23 -2.2125 19.37 ;
        RECT  -3.8475 27.8125 -3.7775 27.9475 ;
        RECT  -3.8475 25.67 -3.7775 25.805 ;
        RECT  -3.6925 26.9925 -3.6225 27.1275 ;
        RECT  -3.6925 25.67 -3.6225 25.805 ;
        RECT  -2.8325 27.1975 -2.7625 27.3325 ;
        RECT  -2.8325 25.67 -2.7625 25.805 ;
        RECT  -2.4375 27.4025 -2.3675 27.5375 ;
        RECT  -2.4375 25.67 -2.3675 25.805 ;
        RECT  -4.045 26.7875 -3.975 26.9225 ;
        RECT  -4.045 25.67 -3.975 25.805 ;
        RECT  -3.34 26.7875 -3.27 26.9225 ;
        RECT  -3.34 25.67 -3.27 25.805 ;
        RECT  -2.635 26.7875 -2.565 26.9225 ;
        RECT  -2.635 25.67 -2.565 25.805 ;
        RECT  -1.93 26.7875 -1.86 26.9225 ;
        RECT  -1.93 25.67 -1.86 25.805 ;
        RECT  -2.245 33.615 -0.725 33.685 ;
        RECT  -0.76 33.5825 -0.69 33.7175 ;
        RECT  -2.28 33.5825 -2.21 33.7175 ;
        RECT  -0.7575 28.0175 -0.6875 28.1525 ;
        RECT  -0.7575 23.0 -0.6875 23.135 ;
        RECT  -1.9225 28.0175 -1.8525 28.1525 ;
        RECT  -1.9225 29.635 -1.8525 29.77 ;
        RECT  -2.4525 27.8125 -2.3825 27.9475 ;
        RECT  -2.4525 29.635 -2.3825 29.77 ;
        RECT  9.8 30.61 9.935 30.68 ;
        RECT  -0.275 30.61 -0.14 30.68 ;
        RECT  9.595 31.85 9.73 31.92 ;
        RECT  -0.275 31.85 -0.14 31.92 ;
        RECT  9.185 29.41 9.32 29.48 ;
        RECT  -0.275 29.41 -0.14 29.48 ;
        RECT  8.98 30.385 9.115 30.455 ;
        RECT  -0.275 30.385 -0.14 30.455 ;
        RECT  9.39 28.05 9.525 28.12 ;
        RECT  -0.275 28.05 -0.14 28.12 ;
        RECT  8.775 26.615 8.91 26.685 ;
        RECT  -0.275 26.615 -0.14 26.685 ;
        RECT  8.36 26.82 8.495 26.89 ;
        RECT  -0.275 26.82 -0.14 26.89 ;
    END
END    sram_2_16_1_freepdk45
END    LIBRARY
