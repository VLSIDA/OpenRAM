magic
tech sky130A
magscale 1 2
timestamp 1595931502
<< checkpaint >>
rect -1260 -1316 8744 7665
<< locali >>
rect 5475 6185 5538 6219
rect 5504 6038 5538 6185
rect 7438 6156 7466 6190
rect 5504 6004 5607 6038
rect 5504 5812 5607 5846
rect 5504 5723 5538 5812
rect 5475 5689 5538 5723
rect 7438 5660 7466 5694
rect 5475 5395 5538 5429
rect 5504 5248 5538 5395
rect 7438 5366 7466 5400
rect 5504 5214 5607 5248
rect 5504 5022 5607 5056
rect 5504 4933 5538 5022
rect 5475 4899 5538 4933
rect 7438 4870 7466 4904
rect 5475 4605 5538 4639
rect 5504 4458 5538 4605
rect 7438 4576 7466 4610
rect 5504 4424 5607 4458
rect 5504 4232 5607 4266
rect 5504 4143 5538 4232
rect 5475 4109 5538 4143
rect 7438 4080 7466 4114
rect 5475 3815 5538 3849
rect 5504 3668 5538 3815
rect 7438 3786 7466 3820
rect 5504 3634 5607 3668
rect 5504 3442 5607 3476
rect 5504 3353 5538 3442
rect 5475 3319 5538 3353
rect 7438 3290 7466 3324
rect 5475 3025 5538 3059
rect 5504 2878 5538 3025
rect 7438 2996 7466 3030
rect 5504 2844 5607 2878
rect 5504 2652 5607 2686
rect 5504 2563 5538 2652
rect 5475 2529 5538 2563
rect 7438 2500 7466 2534
rect 5475 2235 5538 2269
rect 5504 2088 5538 2235
rect 7438 2206 7466 2240
rect 5504 2054 5607 2088
rect 5504 1862 5607 1896
rect 5504 1773 5538 1862
rect 5475 1739 5538 1773
rect 7438 1710 7466 1744
rect 5475 1445 5538 1479
rect 5504 1298 5538 1445
rect 7438 1416 7466 1450
rect 5504 1264 5607 1298
rect 5504 1072 5607 1106
rect 5504 983 5538 1072
rect 5475 949 5538 983
rect 7438 920 7466 954
rect 5475 655 5538 689
rect 5504 508 5538 655
rect 7438 626 7466 660
rect 5504 474 5607 508
rect 5504 282 5607 316
rect 5504 193 5538 282
rect 5475 159 5538 193
rect 7438 130 7466 164
<< metal1 >>
rect 18 29 46 3979
rect 98 29 126 3979
rect 178 29 206 3979
rect 258 29 286 3979
<< metal2 >>
rect 5590 0 5618 6320
rect 5762 3121 5818 3169
rect 6187 3120 6243 3168
rect 6604 3136 6660 3184
rect 7102 3136 7158 3184
<< metal3 >>
rect 4219 5912 4317 6010
rect 4644 5912 4742 6010
rect 5023 5905 5121 6003
rect 5295 5905 5393 6003
rect 4219 5540 4317 5638
rect 4644 5542 4742 5640
rect 5023 5510 5121 5608
rect 5295 5510 5393 5608
rect 4219 5122 4317 5220
rect 4644 5122 4742 5220
rect 5023 5115 5121 5213
rect 5295 5115 5393 5213
rect 4219 4750 4317 4848
rect 4644 4752 4742 4850
rect 5023 4720 5121 4818
rect 5295 4720 5393 4818
rect 4219 4332 4317 4430
rect 4644 4332 4742 4430
rect 5023 4325 5121 4423
rect 5295 4325 5393 4423
rect 4219 3960 4317 4058
rect 4644 3962 4742 4060
rect 5023 3930 5121 4028
rect 5295 3930 5393 4028
rect 2005 3542 2103 3640
rect 2430 3542 2528 3640
rect 2809 3535 2907 3633
rect 3081 3535 3179 3633
rect 4219 3542 4317 3640
rect 4644 3542 4742 3640
rect 5023 3535 5121 3633
rect 5295 3535 5393 3633
rect 4219 3170 4317 3268
rect 4644 3172 4742 3270
rect 5023 3140 5121 3238
rect 5295 3140 5393 3238
rect 5741 3096 5839 3194
rect 6166 3095 6264 3193
rect 6583 3111 6681 3209
rect 7081 3111 7179 3209
rect 835 2745 933 2843
rect 1107 2745 1205 2843
rect 2005 2752 2103 2850
rect 2430 2752 2528 2850
rect 2809 2745 2907 2843
rect 3081 2745 3179 2843
rect 4219 2752 4317 2850
rect 4644 2752 4742 2850
rect 5023 2745 5121 2843
rect 5295 2745 5393 2843
rect 4219 2380 4317 2478
rect 4644 2382 4742 2480
rect 5023 2350 5121 2448
rect 5295 2350 5393 2448
rect 4219 1962 4317 2060
rect 4644 1962 4742 2060
rect 5023 1955 5121 2053
rect 5295 1955 5393 2053
rect 4219 1590 4317 1688
rect 4644 1592 4742 1690
rect 5023 1560 5121 1658
rect 5295 1560 5393 1658
rect 2005 1172 2103 1270
rect 2430 1172 2528 1270
rect 2809 1165 2907 1263
rect 3081 1165 3179 1263
rect 4219 1172 4317 1270
rect 4644 1172 4742 1270
rect 5023 1165 5121 1263
rect 5295 1165 5393 1263
rect 4219 800 4317 898
rect 4644 802 4742 900
rect 5023 770 5121 868
rect 5295 770 5393 868
rect 835 375 933 473
rect 1107 375 1205 473
rect 2005 382 2103 480
rect 2430 382 2528 480
rect 2809 375 2907 473
rect 3081 375 3179 473
rect 4219 382 4317 480
rect 4644 382 4742 480
rect 5023 375 5121 473
rect 5295 375 5393 473
use wordline_driver_array  wordline_driver_array_0
timestamp 1595931502
transform 1 0 5520 0 1 0
box 70 -56 1964 6376
use contact_9  contact_9_3
timestamp 1595931502
transform 1 0 7097 0 1 3123
box 0 0 66 74
use contact_9  contact_9_2
timestamp 1595931502
transform 1 0 6182 0 1 3107
box 0 0 66 74
use contact_9  contact_9_1
timestamp 1595931502
transform 1 0 6599 0 1 3123
box 0 0 66 74
use contact_9  contact_9_0
timestamp 1595931502
transform 1 0 5757 0 1 3108
box 0 0 66 74
use hierarchical_decoder  hierarchical_decoder_0
timestamp 1595931502
transform 1 0 0 0 1 0
box 0 -27 5510 6405
use contact_8  contact_8_3
timestamp 1595931502
transform 1 0 7098 0 1 3128
box 0 0 64 64
use contact_8  contact_8_2
timestamp 1595931502
transform 1 0 6183 0 1 3112
box 0 0 64 64
use contact_8  contact_8_1
timestamp 1595931502
transform 1 0 6600 0 1 3128
box 0 0 64 64
use contact_8  contact_8_0
timestamp 1595931502
transform 1 0 5758 0 1 3113
box 0 0 64 64
<< labels >>
rlabel corelocali s 7452 147 7452 147 4 wl_0
rlabel corelocali s 7452 937 7452 937 4 wl_2
rlabel corelocali s 7452 4097 7452 4097 4 wl_10
rlabel corelocali s 7452 1433 7452 1433 4 wl_3
rlabel metal1 s 32 2004 32 2004 4 addr_0
rlabel corelocali s 7452 5383 7452 5383 4 wl_13
rlabel corelocali s 7452 3307 7452 3307 4 wl_8
rlabel corelocali s 7452 4593 7452 4593 4 wl_11
rlabel metal1 s 192 2004 192 2004 4 addr_2
rlabel metal1 s 112 2004 112 2004 4 addr_1
rlabel metal3 s 5072 3189 5072 3189 4 gnd
rlabel metal3 s 5790 3145 5790 3145 4 gnd
rlabel metal3 s 5072 424 5072 424 4 gnd
rlabel metal3 s 4268 3219 4268 3219 4 gnd
rlabel metal3 s 4268 4799 4268 4799 4 gnd
rlabel metal3 s 2858 3584 2858 3584 4 gnd
rlabel metal3 s 5072 819 5072 819 4 gnd
rlabel metal3 s 2858 1214 2858 1214 4 gnd
rlabel metal3 s 4268 1221 4268 1221 4 gnd
rlabel metal3 s 4268 2801 4268 2801 4 gnd
rlabel metal3 s 5072 5559 5072 5559 4 gnd
rlabel metal3 s 4268 431 4268 431 4 gnd
rlabel metal3 s 5072 5954 5072 5954 4 gnd
rlabel metal3 s 4268 1639 4268 1639 4 gnd
rlabel metal3 s 2054 3591 2054 3591 4 gnd
rlabel metal3 s 4268 849 4268 849 4 gnd
rlabel metal3 s 884 424 884 424 4 gnd
rlabel metal3 s 2858 2794 2858 2794 4 gnd
rlabel metal3 s 4268 5589 4268 5589 4 gnd
rlabel metal3 s 4268 4381 4268 4381 4 gnd
rlabel metal3 s 884 2794 884 2794 4 gnd
rlabel metal3 s 5072 3979 5072 3979 4 gnd
rlabel metal3 s 5072 5164 5072 5164 4 gnd
rlabel metal3 s 2054 1221 2054 1221 4 gnd
rlabel metal3 s 2054 2801 2054 2801 4 gnd
rlabel metal3 s 5072 4374 5072 4374 4 gnd
rlabel metal3 s 2858 424 2858 424 4 gnd
rlabel metal3 s 5072 2399 5072 2399 4 gnd
rlabel metal3 s 5072 3584 5072 3584 4 gnd
rlabel metal3 s 4268 3591 4268 3591 4 gnd
rlabel metal3 s 5072 4769 5072 4769 4 gnd
rlabel metal3 s 4268 5171 4268 5171 4 gnd
rlabel metal3 s 4268 2429 4268 2429 4 gnd
rlabel metal3 s 4268 4009 4268 4009 4 gnd
rlabel metal3 s 2054 431 2054 431 4 gnd
rlabel metal3 s 6632 3160 6632 3160 4 gnd
rlabel metal3 s 4268 2011 4268 2011 4 gnd
rlabel metal3 s 4268 5961 4268 5961 4 gnd
rlabel metal3 s 5072 1214 5072 1214 4 gnd
rlabel metal3 s 5072 1609 5072 1609 4 gnd
rlabel metal3 s 5072 2794 5072 2794 4 gnd
rlabel metal3 s 5072 2004 5072 2004 4 gnd
rlabel corelocali s 7452 4887 7452 4887 4 wl_12
rlabel corelocali s 7452 2517 7452 2517 4 wl_6
rlabel corelocali s 7452 3803 7452 3803 4 wl_9
rlabel corelocali s 7452 3013 7452 3013 4 wl_7
rlabel metal1 s 272 2004 272 2004 4 addr_3
rlabel corelocali s 7452 1727 7452 1727 4 wl_4
rlabel corelocali s 7452 5677 7452 5677 4 wl_14
rlabel corelocali s 7452 6173 7452 6173 4 wl_15
rlabel corelocali s 7452 643 7452 643 4 wl_1
rlabel corelocali s 7452 2223 7452 2223 4 wl_5
rlabel metal3 s 4693 2431 4693 2431 4 vdd
rlabel metal3 s 4693 431 4693 431 4 vdd
rlabel metal3 s 5344 1609 5344 1609 4 vdd
rlabel metal3 s 5344 5954 5344 5954 4 vdd
rlabel metal3 s 4693 3221 4693 3221 4 vdd
rlabel metal3 s 2479 3591 2479 3591 4 vdd
rlabel metal3 s 5344 3584 5344 3584 4 vdd
rlabel metal3 s 1156 424 1156 424 4 vdd
rlabel metal3 s 4693 4801 4693 4801 4 vdd
rlabel metal3 s 5344 1214 5344 1214 4 vdd
rlabel metal3 s 1156 2794 1156 2794 4 vdd
rlabel metal3 s 5344 3979 5344 3979 4 vdd
rlabel metal3 s 3130 3584 3130 3584 4 vdd
rlabel metal3 s 3130 1214 3130 1214 4 vdd
rlabel metal3 s 4693 2011 4693 2011 4 vdd
rlabel metal3 s 2479 1221 2479 1221 4 vdd
rlabel metal3 s 5344 2794 5344 2794 4 vdd
rlabel metal3 s 5344 2399 5344 2399 4 vdd
rlabel metal3 s 4693 4381 4693 4381 4 vdd
rlabel metal3 s 5344 5559 5344 5559 4 vdd
rlabel metal3 s 6215 3144 6215 3144 4 vdd
rlabel metal3 s 2479 431 2479 431 4 vdd
rlabel metal3 s 7130 3160 7130 3160 4 vdd
rlabel metal3 s 2479 2801 2479 2801 4 vdd
rlabel metal3 s 4693 5591 4693 5591 4 vdd
rlabel metal3 s 4693 3591 4693 3591 4 vdd
rlabel metal3 s 4693 851 4693 851 4 vdd
rlabel metal3 s 5344 5164 5344 5164 4 vdd
rlabel metal3 s 5344 424 5344 424 4 vdd
rlabel metal3 s 4693 5961 4693 5961 4 vdd
rlabel metal3 s 5344 4769 5344 4769 4 vdd
rlabel metal3 s 4693 4011 4693 4011 4 vdd
rlabel metal3 s 5344 2004 5344 2004 4 vdd
rlabel metal3 s 4693 5171 4693 5171 4 vdd
rlabel metal3 s 4693 1641 4693 1641 4 vdd
rlabel metal3 s 5344 3189 5344 3189 4 vdd
rlabel metal3 s 3130 424 3130 424 4 vdd
rlabel metal3 s 3130 2794 3130 2794 4 vdd
rlabel metal3 s 5344 819 5344 819 4 vdd
rlabel metal3 s 4693 1221 4693 1221 4 vdd
rlabel metal3 s 4693 2801 4693 2801 4 vdd
rlabel metal3 s 5344 4374 5344 4374 4 vdd
rlabel metal2 s 5604 3160 5604 3160 4 wl_en
<< properties >>
string FIXED_BBOX 0 0 7502 6348
<< end >>
