*********************************************
* Transistor Models
* Note: These models are approximate 
*       and should be substituted with actual
*       models from MOSIS or SCN3ME
*********************************************

.MODEL n NMOS (LEVEL=49 VTO=0.669845 KP=113.7771E-6
+ NSUB=6E16 U0=459 GAMMA=0.5705 TOX=13.9n)

