magic
tech gf180mcuD
magscale 1 10
timestamp 1694481086
<< nwell >>
rect 620 0 1222 620
<< nmos >>
rect 156 340 326 400
rect 156 230 326 290
<< pmos >>
rect 710 370 1051 430
rect 710 200 1051 260
<< ndiff >>
rect 156 478 326 500
rect 156 432 218 478
rect 264 432 326 478
rect 156 400 326 432
rect 156 290 326 340
rect 156 198 326 230
rect 156 152 218 198
rect 264 152 326 198
rect 156 130 326 152
<< pdiff >>
rect 710 508 1051 530
rect 710 462 763 508
rect 997 462 1051 508
rect 710 430 1051 462
rect 710 338 1051 370
rect 710 292 763 338
rect 997 292 1051 338
rect 710 260 1051 292
rect 710 168 1051 200
rect 710 122 763 168
rect 997 122 1051 168
rect 710 100 1051 122
<< ndiffc >>
rect 218 432 264 478
rect 218 152 264 198
<< pdiffc >>
rect 763 462 997 508
rect 763 292 997 338
rect 763 122 997 168
<< psubdiff >>
rect 19 63 126 80
rect 19 17 59 63
rect 105 17 126 63
rect 19 0 126 17
<< nsubdiff >>
rect 1117 147 1197 184
rect 1117 101 1134 147
rect 1180 101 1197 147
rect 1117 77 1197 101
<< psubdiffcont >>
rect 59 17 105 63
<< nsubdiffcont >>
rect 1134 101 1180 147
<< polysilicon >>
rect 33 413 116 440
rect 33 367 49 413
rect 95 400 116 413
rect 376 400 710 430
rect 95 367 156 400
rect 33 340 156 367
rect 326 370 710 400
rect 1051 370 1101 430
rect 326 340 416 370
rect 33 274 156 290
rect 33 228 49 274
rect 95 230 156 274
rect 326 260 416 290
rect 326 230 710 260
rect 95 228 116 230
rect 33 190 116 228
rect 376 200 710 230
rect 1051 200 1101 260
<< polycontact >>
rect 49 367 95 413
rect 49 228 95 274
<< metal1 >>
rect 156 478 396 480
rect 46 413 98 465
rect 156 432 218 478
rect 264 432 396 478
rect 752 462 763 508
rect 997 462 1009 508
rect 848 456 860 462
rect 912 456 924 462
rect 156 430 396 432
rect 46 367 49 413
rect 95 367 98 413
rect 46 353 98 367
rect 346 340 396 430
rect 1075 340 1127 503
rect 346 338 1127 340
rect 346 292 763 338
rect 997 292 1127 338
rect 346 290 1127 292
rect 46 274 98 288
rect 46 228 49 274
rect 95 228 98 274
rect 46 169 98 228
rect 186 146 218 198
rect 270 146 293 198
rect 848 168 860 174
rect 912 168 924 174
rect 186 140 293 146
rect 752 122 763 168
rect 997 122 1009 168
rect 1084 98 1131 150
rect 1183 98 1195 150
rect 25 66 124 76
rect 25 14 56 66
rect 108 14 124 66
rect 25 6 124 14
<< via1 >>
rect 860 462 912 508
rect 860 456 912 462
rect 218 152 264 198
rect 264 152 270 198
rect 218 146 270 152
rect 860 168 912 174
rect 860 122 912 168
rect 1131 147 1183 150
rect 1131 101 1134 147
rect 1134 101 1180 147
rect 1180 101 1183 147
rect 1131 98 1183 101
rect 56 63 108 66
rect 56 17 59 63
rect 59 17 105 63
rect 105 17 108 63
rect 56 14 108 17
<< metal2 >>
rect 216 198 272 560
rect 216 146 218 198
rect 270 146 272 198
rect 216 68 272 146
rect 34 66 272 68
rect 34 14 56 66
rect 108 14 272 66
rect 858 508 914 560
rect 858 456 860 508
rect 912 456 914 508
rect 858 174 914 456
rect 858 122 860 174
rect 912 152 914 174
rect 912 150 1195 152
rect 912 122 1131 150
rect 858 98 1131 122
rect 1183 98 1195 150
rect 858 96 1195 98
rect 858 48 914 96
rect 34 12 272 14
<< labels >>
rlabel metal1 s 73 390 73 390 4 B
rlabel metal1 s 73 251 73 251 4 A
rlabel metal2 s 886 73 886 73 4 VDD
rlabel metal2 s 245 96 245 96 4 GND
rlabel metal1 1101 479 1101 479 1 Y
<< properties >>
string FIXED_BBOX 0 0 1339 620
string GDS_END 11704
string GDS_START 6968
<< end >>
