magic
tech sky130A
magscale 1 2
timestamp 1595931502
<< checkpaint >>
rect -1268 -1309 2436 6965
<< metal1 >>
rect 552 5630 616 5682
rect 552 4216 616 4268
rect 552 2802 616 2854
rect 552 1388 616 1440
rect 552 -26 616 26
<< metal2 >>
rect 137 5066 203 5118
rect 137 3366 203 3418
rect 137 2238 203 2290
rect 137 538 203 590
rect 369 0 397 5656
rect 556 5632 612 5680
rect 1082 4995 1148 5047
rect 556 4218 612 4266
rect 1082 3437 1148 3489
rect 556 2804 612 2852
rect 1082 2167 1148 2219
rect 556 1390 612 1438
rect 1082 609 1148 661
rect 556 -24 612 24
<< metal3 >>
rect 535 5607 633 5705
rect 535 4193 633 4291
rect 535 2779 633 2877
rect 535 1365 633 1463
rect 0 278 1168 338
rect 535 -49 633 49
use contact_9  contact_9_8
timestamp 1595931502
transform 1 0 551 0 1 1377
box 0 0 66 74
use contact_9  contact_9_7
timestamp 1595931502
transform 1 0 551 0 1 -37
box 0 0 66 74
use contact_9  contact_9_6
timestamp 1595931502
transform 1 0 551 0 1 1377
box 0 0 66 74
use contact_9  contact_9_5
timestamp 1595931502
transform 1 0 551 0 1 2791
box 0 0 66 74
use contact_9  contact_9_4
timestamp 1595931502
transform 1 0 551 0 1 4205
box 0 0 66 74
use contact_9  contact_9_3
timestamp 1595931502
transform 1 0 551 0 1 2791
box 0 0 66 74
use contact_9  contact_9_2
timestamp 1595931502
transform 1 0 551 0 1 4205
box 0 0 66 74
use contact_9  contact_9_1
timestamp 1595931502
transform 1 0 551 0 1 5619
box 0 0 66 74
use contact_9  contact_9_0
timestamp 1595931502
transform 1 0 363 0 1 271
box 0 0 66 74
use contact_8  contact_8_0
timestamp 1595931502
transform 1 0 552 0 1 5624
box 0 0 64 64
use contact_7  contact_7_0
timestamp 1595931502
transform 1 0 555 0 1 5623
box 0 0 58 66
use contact_8  contact_8_1
timestamp 1595931502
transform 1 0 552 0 1 4210
box 0 0 64 64
use contact_7  contact_7_1
timestamp 1595931502
transform 1 0 555 0 1 4209
box 0 0 58 66
use contact_8  contact_8_2
timestamp 1595931502
transform 1 0 552 0 1 2796
box 0 0 64 64
use contact_7  contact_7_2
timestamp 1595931502
transform 1 0 555 0 1 2795
box 0 0 58 66
use contact_8  contact_8_3
timestamp 1595931502
transform 1 0 552 0 1 4210
box 0 0 64 64
use contact_7  contact_7_3
timestamp 1595931502
transform 1 0 555 0 1 4209
box 0 0 58 66
use contact_8  contact_8_4
timestamp 1595931502
transform 1 0 552 0 1 2796
box 0 0 64 64
use contact_7  contact_7_4
timestamp 1595931502
transform 1 0 555 0 1 2795
box 0 0 58 66
use contact_8  contact_8_5
timestamp 1595931502
transform 1 0 552 0 1 1382
box 0 0 64 64
use contact_7  contact_7_5
timestamp 1595931502
transform 1 0 555 0 1 1381
box 0 0 58 66
use contact_8  contact_8_6
timestamp 1595931502
transform 1 0 552 0 1 -32
box 0 0 64 64
use contact_7  contact_7_6
timestamp 1595931502
transform 1 0 555 0 1 -33
box 0 0 58 66
use contact_8  contact_8_7
timestamp 1595931502
transform 1 0 552 0 1 1382
box 0 0 64 64
use contact_7  contact_7_7
timestamp 1595931502
transform 1 0 555 0 1 1381
box 0 0 58 66
use dff  dff_0
timestamp 1595931502
transform 1 0 0 0 -1 5656
box -8 -20 1176 1467
use dff  dff_1
timestamp 1595931502
transform 1 0 0 0 1 2828
box -8 -20 1176 1467
use dff  dff_2
timestamp 1595931502
transform 1 0 0 0 -1 2828
box -8 -20 1176 1467
use dff  dff_3
timestamp 1595931502
transform 1 0 0 0 1 0
box -8 -20 1176 1467
<< labels >>
rlabel metal3 s 584 0 584 0 4 gnd
rlabel metal3 s 584 5656 584 5656 4 gnd
rlabel metal3 s 584 2828 584 2828 4 gnd
rlabel metal2 s 1115 3463 1115 3463 4 dout_2
rlabel metal2 s 1115 635 1115 635 4 dout_0
rlabel metal2 s 1115 2193 1115 2193 4 dout_1
rlabel metal2 s 170 564 170 564 4 din_0
rlabel metal3 s 584 4242 584 4242 4 vdd
rlabel metal3 s 584 1414 584 1414 4 vdd
rlabel metal2 s 1115 5021 1115 5021 4 dout_3
rlabel metal3 s 584 308 584 308 4 clk
rlabel metal2 s 170 3392 170 3392 4 din_2
rlabel metal2 s 170 5092 170 5092 4 din_3
rlabel metal2 s 170 2264 170 2264 4 din_1
<< properties >>
string FIXED_BBOX 0 0 1168 5656
<< end >>
