magic
tech sky130A
timestamp 1595931502
<< checkpaint >>
rect -630 -630 663 663
<< poly >>
rect 0 25 33 33
rect 0 8 8 25
rect 25 8 33 25
rect 0 0 33 8
<< polycont >>
rect 8 8 25 25
<< locali >>
rect 8 25 25 33
rect 8 0 25 8
<< properties >>
string FIXED_BBOX -10 -10 43 43
<< end >>
