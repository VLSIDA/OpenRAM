MACRO sram_2_16_1_freepdk45
    CLASS RING ;
    ORIGIN 5.765 0.0 ;
    FOREIGN  sram 0.0 0.0 ;
    SIZE 19.165 BY 41.725 ;
    SYMMETRY X Y R90 ;
    PIN vdd
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  0.0325 0.0 0.7325 41.725 ;
        RECT  12.7675 0.0 13.4675 41.725 ;
        END
    END vdd
    PIN gnd
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal2 ;
        RECT  8.9225 0.0 9.6225 41.725 ;
        END
    END gnd
    PIN DATA[0]
        DIRECTION INOUT ;
        PORT
        LAYER metal3 ;
        RECT  11.48 0.0 11.55 3.22 ;
        RECT  11.48 0.0 11.55 0.135 ;
        END
    END DATA[0]
    PIN DATA[1]
        DIRECTION INOUT ;
        PORT
        LAYER metal3 ;
        RECT  12.185 0.0 12.255 3.22 ;
        RECT  12.185 0.0 12.255 0.135 ;
        END
    END DATA[1]
    PIN ADDR[0]
        DIRECTION INPUT ;
        PORT
        LAYER metal3 ;
        RECT  0.0325 7.4525 1.015 7.5225 ;
        END
    END ADDR[0]
    PIN ADDR[1]
        DIRECTION INPUT ;
        PORT
        LAYER metal3 ;
        RECT  0.0325 6.7475 1.015 6.8175 ;
        END
    END ADDR[1]
    PIN ADDR[2]
        DIRECTION INPUT ;
        PORT
        LAYER metal3 ;
        RECT  0.0325 6.0425 1.015 6.1125 ;
        END
    END ADDR[2]
    PIN ADDR[3]
        DIRECTION INPUT ;
        PORT
        LAYER metal3 ;
        RECT  0.0325 5.3375 1.015 5.4075 ;
        END
    END ADDR[3]
    PIN CSb
        DIRECTION INPUT ;
        PORT
        LAYER metal3 ;
        RECT  -5.4125 8.275 -5.3425 8.415 ;
        END
    END CSb
    PIN OEb
        DIRECTION INPUT ;
        PORT
        LAYER metal3 ;
        RECT  -4.0025 8.275 -3.9325 8.415 ;
        END
    END OEb
    PIN WEb
        DIRECTION INPUT ;
        PORT
        LAYER metal3 ;
        RECT  -4.7075 8.275 -4.6375 8.415 ;
        END
    END WEb
    PIN clk
        DIRECTION INPUT ;
        PORT
        LAYER metal3 ;
        RECT  -2.0525 8.275 9.7625 8.345 ;
        RECT  -2.085 8.275 -2.015 8.41 ;
        END
    END clk
    OBS
        LAYER  metal1 ;
        RECT  -0.545 26.2975 0.0325 26.3625 ;
        RECT  12.7675 0.0 13.4675 41.725 ;
        RECT  0.0325 0.0 0.7325 41.725 ;
        RECT  5.5625 19.49 5.6275 19.87 ;
        RECT  7.8875 19.0025 7.9525 19.0675 ;
        RECT  7.92 19.0025 11.195 19.0675 ;
        RECT  7.8875 19.035 7.9525 19.575 ;
        RECT  5.5625 20.61 5.6275 20.99 ;
        RECT  7.8875 21.4125 7.9525 21.4775 ;
        RECT  7.92 21.4125 11.195 21.4775 ;
        RECT  7.8875 20.905 7.9525 21.445 ;
        RECT  5.5625 22.18 5.6275 22.56 ;
        RECT  7.8875 21.6925 7.9525 21.7575 ;
        RECT  7.92 21.6925 11.195 21.7575 ;
        RECT  7.8875 21.725 7.9525 22.265 ;
        RECT  5.5625 23.3 5.6275 23.68 ;
        RECT  7.8875 24.1025 7.9525 24.1675 ;
        RECT  7.92 24.1025 11.195 24.1675 ;
        RECT  7.8875 23.595 7.9525 24.135 ;
        RECT  5.5625 24.87 5.6275 25.25 ;
        RECT  7.8875 24.3825 7.9525 24.4475 ;
        RECT  7.92 24.3825 11.195 24.4475 ;
        RECT  7.8875 24.415 7.9525 24.955 ;
        RECT  5.5625 25.99 5.6275 26.37 ;
        RECT  7.8875 26.7925 7.9525 26.8575 ;
        RECT  7.92 26.7925 11.195 26.8575 ;
        RECT  7.8875 26.285 7.9525 26.825 ;
        RECT  5.5625 27.56 5.6275 27.94 ;
        RECT  7.8875 27.0725 7.9525 27.1375 ;
        RECT  7.92 27.0725 11.195 27.1375 ;
        RECT  7.8875 27.105 7.9525 27.645 ;
        RECT  5.5625 28.68 5.6275 29.06 ;
        RECT  7.8875 29.4825 7.9525 29.5475 ;
        RECT  7.92 29.4825 11.195 29.5475 ;
        RECT  7.8875 28.975 7.9525 29.515 ;
        RECT  5.5625 30.25 5.6275 30.63 ;
        RECT  7.8875 29.7625 7.9525 29.8275 ;
        RECT  7.92 29.7625 11.195 29.8275 ;
        RECT  7.8875 29.795 7.9525 30.335 ;
        RECT  5.5625 31.37 5.6275 31.75 ;
        RECT  7.8875 32.1725 7.9525 32.2375 ;
        RECT  7.92 32.1725 11.195 32.2375 ;
        RECT  7.8875 31.665 7.9525 32.205 ;
        RECT  5.5625 32.94 5.6275 33.32 ;
        RECT  7.8875 32.4525 7.9525 32.5175 ;
        RECT  7.92 32.4525 11.195 32.5175 ;
        RECT  7.8875 32.485 7.9525 33.025 ;
        RECT  5.5625 34.06 5.6275 34.44 ;
        RECT  7.8875 34.8625 7.9525 34.9275 ;
        RECT  7.92 34.8625 11.195 34.9275 ;
        RECT  7.8875 34.355 7.9525 34.895 ;
        RECT  5.5625 35.63 5.6275 36.01 ;
        RECT  7.8875 35.1425 7.9525 35.2075 ;
        RECT  7.92 35.1425 11.195 35.2075 ;
        RECT  7.8875 35.175 7.9525 35.715 ;
        RECT  5.5625 36.75 5.6275 37.13 ;
        RECT  7.8875 37.5525 7.9525 37.6175 ;
        RECT  7.92 37.5525 11.195 37.6175 ;
        RECT  7.8875 37.045 7.9525 37.585 ;
        RECT  5.5625 38.32 5.6275 38.7 ;
        RECT  7.8875 37.8325 7.9525 37.8975 ;
        RECT  7.92 37.8325 11.195 37.8975 ;
        RECT  7.8875 37.865 7.9525 38.405 ;
        RECT  5.5625 39.44 5.6275 39.82 ;
        RECT  7.8875 40.2425 7.9525 40.3075 ;
        RECT  7.92 40.2425 11.195 40.3075 ;
        RECT  7.8875 39.735 7.9525 40.275 ;
        RECT  7.8875 20.2075 11.1625 20.2725 ;
        RECT  7.8875 22.8975 11.1625 22.9625 ;
        RECT  7.8875 25.5875 11.1625 25.6525 ;
        RECT  7.8875 28.2775 11.1625 28.3425 ;
        RECT  7.8875 30.9675 11.1625 31.0325 ;
        RECT  7.8875 33.6575 11.1625 33.7225 ;
        RECT  7.8875 36.3475 11.1625 36.4125 ;
        RECT  7.8875 39.0375 11.1625 39.1025 ;
        RECT  7.2775 8.73 8.6425 8.795 ;
        RECT  7.2775 10.165 8.4325 10.23 ;
        RECT  7.2775 14.11 8.2225 14.175 ;
        RECT  7.2775 15.545 8.0125 15.61 ;
        RECT  10.3925 3.6 11.515 3.665 ;
        RECT  9.9725 1.415 11.5325 1.48 ;
        RECT  10.1825 2.9625 11.5325 3.0275 ;
        RECT  10.3925 41.1 11.1625 41.165 ;
        RECT  10.6025 10.1025 11.1625 10.1675 ;
        RECT  10.8125 14.1275 11.1625 14.1925 ;
        RECT  5.7575 41.53 5.8225 41.595 ;
        RECT  5.7575 40.415 5.8225 41.5625 ;
        RECT  5.79 41.53 9.8275 41.595 ;
        RECT  11.1625 20.2075 12.7675 20.2725 ;
        RECT  11.1625 22.8975 12.7675 22.9625 ;
        RECT  11.1625 25.5875 12.7675 25.6525 ;
        RECT  11.1625 28.2775 12.7675 28.3425 ;
        RECT  11.1625 30.9675 12.7675 31.0325 ;
        RECT  11.1625 33.6575 12.7675 33.7225 ;
        RECT  11.1625 36.3475 12.7675 36.4125 ;
        RECT  11.1625 39.0375 12.7675 39.1025 ;
        RECT  11.1625 41.66 12.7675 41.725 ;
        RECT  11.1625 18.7 12.7675 18.765 ;
        RECT  11.1625 10.2325 12.7675 10.2975 ;
        RECT  11.1625 9.565 12.7675 9.63 ;
        RECT  11.5325 1.545 12.7675 1.61 ;
        RECT  12.2025 1.545 12.7675 1.61 ;
        RECT  0.0325 20.2075 4.2525 20.2725 ;
        RECT  0.0325 22.8975 4.2525 22.9625 ;
        RECT  0.0325 25.5875 4.2525 25.6525 ;
        RECT  0.0325 28.2775 4.2525 28.3425 ;
        RECT  0.0325 30.9675 4.2525 31.0325 ;
        RECT  0.0325 33.6575 4.2525 33.7225 ;
        RECT  0.0325 36.3475 4.2525 36.4125 ;
        RECT  0.0325 39.0375 4.2525 39.1025 ;
        RECT  0.0325 12.1375 4.2525 12.2025 ;
        RECT  0.0325 17.5175 4.2525 17.5825 ;
        RECT  0.0 4.825 0.065 4.89 ;
        RECT  7.1125 4.825 7.1775 4.89 ;
        RECT  0.0 4.825 0.065 4.8575 ;
        RECT  0.0325 4.825 7.145 4.89 ;
        RECT  7.1125 4.8575 7.1775 5.02 ;
        RECT  8.9225 40.545 12.5725 40.61 ;
        RECT  9.4175 0.355 12.5725 0.42 ;
        RECT  4.2525 13.4825 8.9225 13.5475 ;
        RECT  4.2525 18.8625 8.9225 18.9275 ;
        RECT  7.3825 7.8075 8.9225 7.8725 ;
        RECT  7.3825 6.3975 8.9225 6.4625 ;
        RECT  7.3825 6.3975 8.9225 6.4625 ;
        RECT  7.3825 4.9875 8.9225 5.0525 ;
        RECT  11.8325 20.0075 11.8975 20.1425 ;
        RECT  11.6475 20.0075 11.7125 20.1425 ;
        RECT  11.1325 20.0075 11.1975 20.1425 ;
        RECT  11.3175 20.0075 11.3825 20.1425 ;
        RECT  11.6475 19.5425 11.7125 19.6775 ;
        RECT  11.8325 19.5425 11.8975 19.6775 ;
        RECT  11.3175 19.5425 11.3825 19.6775 ;
        RECT  11.1325 19.5425 11.1975 19.6775 ;
        RECT  11.7525 19.1525 11.8175 19.2875 ;
        RECT  11.5675 19.1525 11.6325 19.2875 ;
        RECT  11.3975 19.1525 11.4625 19.2875 ;
        RECT  11.2125 19.1525 11.2775 19.2875 ;
        RECT  11.835 19.645 11.9 19.78 ;
        RECT  11.835 19.645 11.9 19.78 ;
        RECT  11.835 19.645 11.9 19.78 ;
        RECT  11.835 19.645 11.9 19.78 ;
        RECT  11.835 19.645 11.9 19.78 ;
        RECT  11.835 19.645 11.9 19.78 ;
        RECT  11.4425 20.2075 11.5775 20.2725 ;
        RECT  11.095 18.8625 11.23 18.9275 ;
        RECT  11.8 18.8625 11.935 18.9275 ;
        RECT  11.43 19.0025 11.565 19.0675 ;
        RECT  11.835 19.645 11.9 19.78 ;
        RECT  11.835 19.645 11.9 19.78 ;
        RECT  11.835 19.645 11.9 19.78 ;
        RECT  11.835 19.645 11.9 19.78 ;
        RECT  11.335 19.8925 11.47 19.9575 ;
        RECT  11.335 19.8925 11.47 19.9575 ;
        RECT  11.56 19.7425 11.695 19.8075 ;
        RECT  11.56 19.7425 11.695 19.8075 ;
        RECT  11.835 19.645 11.9 19.78 ;
        RECT  11.835 19.645 11.9 19.78 ;
        RECT  11.835 19.645 11.9 19.78 ;
        RECT  11.835 19.645 11.9 19.78 ;
        RECT  11.385 19.1525 11.45 19.2875 ;
        RECT  11.13 19.645 11.195 19.78 ;
        RECT  11.13 19.645 11.195 19.78 ;
        RECT  11.13 19.645 11.195 19.78 ;
        RECT  11.13 19.645 11.195 19.78 ;
        RECT  11.13 19.645 11.195 19.78 ;
        RECT  11.13 19.645 11.195 19.78 ;
        RECT  11.835 19.645 11.9 19.78 ;
        RECT  11.835 19.645 11.9 19.78 ;
        RECT  11.835 19.645 11.9 19.78 ;
        RECT  11.835 19.645 11.9 19.78 ;
        RECT  11.58 19.1525 11.645 19.2875 ;
        RECT  11.4475 18.8625 11.5825 18.9275 ;
        RECT  11.4475 18.8625 11.5825 18.9275 ;
        RECT  11.8 18.8625 11.935 18.9275 ;
        RECT  11.4425 20.2075 11.5775 20.2725 ;
        RECT  11.8 18.8625 11.935 18.9275 ;
        RECT  11.8 18.8625 11.935 18.9275 ;
        RECT  11.835 19.645 11.9 19.78 ;
        RECT  11.835 19.645 11.9 19.78 ;
        RECT  11.835 19.645 11.9 19.78 ;
        RECT  11.835 19.645 11.9 19.78 ;
        RECT  11.835 19.645 11.9 19.78 ;
        RECT  11.835 19.645 11.9 19.78 ;
        RECT  11.095 18.8625 11.23 18.9275 ;
        RECT  11.455 20.2075 11.555 20.27 ;
        RECT  11.455 20.21 11.555 20.2725 ;
        RECT  11.7825 19.005 11.835 19.0675 ;
        RECT  11.455 20.2075 11.555 20.27 ;
        RECT  11.8325 20.0075 11.9025 20.2075 ;
        RECT  11.8325 19.5425 11.9025 19.6775 ;
        RECT  11.8325 19.5425 11.9025 19.6775 ;
        RECT  11.0725 18.8625 11.9575 18.9275 ;
        RECT  11.6475 19.3775 11.8225 19.4425 ;
        RECT  11.1275 19.5425 11.1975 19.6775 ;
        RECT  11.3175 19.3775 11.3825 20.1175 ;
        RECT  11.455 20.21 11.555 20.2725 ;
        RECT  11.0775 19.005 11.13 19.0675 ;
        RECT  11.8325 19.5425 11.9025 19.6775 ;
        RECT  11.0725 20.2075 11.9575 20.2725 ;
        RECT  11.6475 19.3775 11.7125 20.0075 ;
        RECT  11.8325 19.5425 11.9025 19.6775 ;
        RECT  11.8325 19.5425 11.9025 19.6775 ;
        RECT  11.2125 19.1525 11.2825 19.4425 ;
        RECT  11.1275 19.5425 11.1975 19.6775 ;
        RECT  11.0725 19.0025 11.9575 19.0675 ;
        RECT  11.8325 19.5425 11.9025 19.6775 ;
        RECT  11.8325 20.0075 11.9025 20.2075 ;
        RECT  11.1275 20.0075 11.1975 20.2075 ;
        RECT  11.7525 19.1525 11.8225 19.4425 ;
        RECT  11.2125 19.3775 11.3825 19.4425 ;
        RECT  11.8325 20.3375 11.8975 20.4725 ;
        RECT  11.6475 20.3375 11.7125 20.4725 ;
        RECT  11.1325 20.3375 11.1975 20.4725 ;
        RECT  11.3175 20.3375 11.3825 20.4725 ;
        RECT  11.6475 20.8025 11.7125 20.9375 ;
        RECT  11.8325 20.8025 11.8975 20.9375 ;
        RECT  11.3175 20.8025 11.3825 20.9375 ;
        RECT  11.1325 20.8025 11.1975 20.9375 ;
        RECT  11.7525 21.1925 11.8175 21.3275 ;
        RECT  11.5675 21.1925 11.6325 21.3275 ;
        RECT  11.3975 21.1925 11.4625 21.3275 ;
        RECT  11.2125 21.1925 11.2775 21.3275 ;
        RECT  11.835 20.7 11.9 20.835 ;
        RECT  11.835 20.7 11.9 20.835 ;
        RECT  11.835 20.7 11.9 20.835 ;
        RECT  11.835 20.7 11.9 20.835 ;
        RECT  11.835 20.7 11.9 20.835 ;
        RECT  11.835 20.7 11.9 20.835 ;
        RECT  11.4425 20.2075 11.5775 20.2725 ;
        RECT  11.095 21.5525 11.23 21.6175 ;
        RECT  11.8 21.5525 11.935 21.6175 ;
        RECT  11.43 21.4125 11.565 21.4775 ;
        RECT  11.835 20.7 11.9 20.835 ;
        RECT  11.835 20.7 11.9 20.835 ;
        RECT  11.835 20.7 11.9 20.835 ;
        RECT  11.835 20.7 11.9 20.835 ;
        RECT  11.335 20.5225 11.47 20.5875 ;
        RECT  11.335 20.5225 11.47 20.5875 ;
        RECT  11.56 20.6725 11.695 20.7375 ;
        RECT  11.56 20.6725 11.695 20.7375 ;
        RECT  11.835 20.7 11.9 20.835 ;
        RECT  11.835 20.7 11.9 20.835 ;
        RECT  11.835 20.7 11.9 20.835 ;
        RECT  11.835 20.7 11.9 20.835 ;
        RECT  11.385 21.1925 11.45 21.3275 ;
        RECT  11.13 20.7 11.195 20.835 ;
        RECT  11.13 20.7 11.195 20.835 ;
        RECT  11.13 20.7 11.195 20.835 ;
        RECT  11.13 20.7 11.195 20.835 ;
        RECT  11.13 20.7 11.195 20.835 ;
        RECT  11.13 20.7 11.195 20.835 ;
        RECT  11.835 20.7 11.9 20.835 ;
        RECT  11.835 20.7 11.9 20.835 ;
        RECT  11.835 20.7 11.9 20.835 ;
        RECT  11.835 20.7 11.9 20.835 ;
        RECT  11.58 21.1925 11.645 21.3275 ;
        RECT  11.4475 21.5525 11.5825 21.6175 ;
        RECT  11.4475 21.5525 11.5825 21.6175 ;
        RECT  11.8 21.5525 11.935 21.6175 ;
        RECT  11.4425 20.2075 11.5775 20.2725 ;
        RECT  11.8 21.5525 11.935 21.6175 ;
        RECT  11.8 21.5525 11.935 21.6175 ;
        RECT  11.835 20.7 11.9 20.835 ;
        RECT  11.835 20.7 11.9 20.835 ;
        RECT  11.835 20.7 11.9 20.835 ;
        RECT  11.835 20.7 11.9 20.835 ;
        RECT  11.835 20.7 11.9 20.835 ;
        RECT  11.835 20.7 11.9 20.835 ;
        RECT  11.095 21.5525 11.23 21.6175 ;
        RECT  11.455 20.21 11.555 20.2725 ;
        RECT  11.455 20.2075 11.555 20.27 ;
        RECT  11.7825 21.4125 11.835 21.475 ;
        RECT  11.455 20.21 11.555 20.2725 ;
        RECT  11.8325 20.2725 11.9025 20.4725 ;
        RECT  11.8325 20.8025 11.9025 20.9375 ;
        RECT  11.8325 20.8025 11.9025 20.9375 ;
        RECT  11.0725 21.5525 11.9575 21.6175 ;
        RECT  11.6475 21.0375 11.8225 21.1025 ;
        RECT  11.1275 20.8025 11.1975 20.9375 ;
        RECT  11.3175 20.3625 11.3825 21.1025 ;
        RECT  11.455 20.2075 11.555 20.27 ;
        RECT  11.0775 21.4125 11.13 21.475 ;
        RECT  11.8325 20.8025 11.9025 20.9375 ;
        RECT  11.0725 20.2075 11.9575 20.2725 ;
        RECT  11.6475 20.4725 11.7125 21.1025 ;
        RECT  11.8325 20.8025 11.9025 20.9375 ;
        RECT  11.8325 20.8025 11.9025 20.9375 ;
        RECT  11.2125 21.0375 11.2825 21.3275 ;
        RECT  11.1275 20.8025 11.1975 20.9375 ;
        RECT  11.0725 21.4125 11.9575 21.4775 ;
        RECT  11.8325 20.8025 11.9025 20.9375 ;
        RECT  11.8325 20.2725 11.9025 20.4725 ;
        RECT  11.1275 20.2725 11.1975 20.4725 ;
        RECT  11.7525 21.0375 11.8225 21.3275 ;
        RECT  11.2125 21.0375 11.3825 21.1025 ;
        RECT  11.8325 22.6975 11.8975 22.8325 ;
        RECT  11.6475 22.6975 11.7125 22.8325 ;
        RECT  11.1325 22.6975 11.1975 22.8325 ;
        RECT  11.3175 22.6975 11.3825 22.8325 ;
        RECT  11.6475 22.2325 11.7125 22.3675 ;
        RECT  11.8325 22.2325 11.8975 22.3675 ;
        RECT  11.3175 22.2325 11.3825 22.3675 ;
        RECT  11.1325 22.2325 11.1975 22.3675 ;
        RECT  11.7525 21.8425 11.8175 21.9775 ;
        RECT  11.5675 21.8425 11.6325 21.9775 ;
        RECT  11.3975 21.8425 11.4625 21.9775 ;
        RECT  11.2125 21.8425 11.2775 21.9775 ;
        RECT  11.835 22.335 11.9 22.47 ;
        RECT  11.835 22.335 11.9 22.47 ;
        RECT  11.835 22.335 11.9 22.47 ;
        RECT  11.835 22.335 11.9 22.47 ;
        RECT  11.835 22.335 11.9 22.47 ;
        RECT  11.835 22.335 11.9 22.47 ;
        RECT  11.4425 22.8975 11.5775 22.9625 ;
        RECT  11.095 21.5525 11.23 21.6175 ;
        RECT  11.8 21.5525 11.935 21.6175 ;
        RECT  11.43 21.6925 11.565 21.7575 ;
        RECT  11.835 22.335 11.9 22.47 ;
        RECT  11.835 22.335 11.9 22.47 ;
        RECT  11.835 22.335 11.9 22.47 ;
        RECT  11.835 22.335 11.9 22.47 ;
        RECT  11.335 22.5825 11.47 22.6475 ;
        RECT  11.335 22.5825 11.47 22.6475 ;
        RECT  11.56 22.4325 11.695 22.4975 ;
        RECT  11.56 22.4325 11.695 22.4975 ;
        RECT  11.835 22.335 11.9 22.47 ;
        RECT  11.835 22.335 11.9 22.47 ;
        RECT  11.835 22.335 11.9 22.47 ;
        RECT  11.835 22.335 11.9 22.47 ;
        RECT  11.385 21.8425 11.45 21.9775 ;
        RECT  11.13 22.335 11.195 22.47 ;
        RECT  11.13 22.335 11.195 22.47 ;
        RECT  11.13 22.335 11.195 22.47 ;
        RECT  11.13 22.335 11.195 22.47 ;
        RECT  11.13 22.335 11.195 22.47 ;
        RECT  11.13 22.335 11.195 22.47 ;
        RECT  11.835 22.335 11.9 22.47 ;
        RECT  11.835 22.335 11.9 22.47 ;
        RECT  11.835 22.335 11.9 22.47 ;
        RECT  11.835 22.335 11.9 22.47 ;
        RECT  11.58 21.8425 11.645 21.9775 ;
        RECT  11.4475 21.5525 11.5825 21.6175 ;
        RECT  11.4475 21.5525 11.5825 21.6175 ;
        RECT  11.8 21.5525 11.935 21.6175 ;
        RECT  11.4425 22.8975 11.5775 22.9625 ;
        RECT  11.8 21.5525 11.935 21.6175 ;
        RECT  11.8 21.5525 11.935 21.6175 ;
        RECT  11.835 22.335 11.9 22.47 ;
        RECT  11.835 22.335 11.9 22.47 ;
        RECT  11.835 22.335 11.9 22.47 ;
        RECT  11.835 22.335 11.9 22.47 ;
        RECT  11.835 22.335 11.9 22.47 ;
        RECT  11.835 22.335 11.9 22.47 ;
        RECT  11.095 21.5525 11.23 21.6175 ;
        RECT  11.455 22.8975 11.555 22.96 ;
        RECT  11.455 22.9 11.555 22.9625 ;
        RECT  11.7825 21.695 11.835 21.7575 ;
        RECT  11.455 22.8975 11.555 22.96 ;
        RECT  11.8325 22.6975 11.9025 22.8975 ;
        RECT  11.8325 22.2325 11.9025 22.3675 ;
        RECT  11.8325 22.2325 11.9025 22.3675 ;
        RECT  11.0725 21.5525 11.9575 21.6175 ;
        RECT  11.6475 22.0675 11.8225 22.1325 ;
        RECT  11.1275 22.2325 11.1975 22.3675 ;
        RECT  11.3175 22.0675 11.3825 22.8075 ;
        RECT  11.455 22.9 11.555 22.9625 ;
        RECT  11.0775 21.695 11.13 21.7575 ;
        RECT  11.8325 22.2325 11.9025 22.3675 ;
        RECT  11.0725 22.8975 11.9575 22.9625 ;
        RECT  11.6475 22.0675 11.7125 22.6975 ;
        RECT  11.8325 22.2325 11.9025 22.3675 ;
        RECT  11.8325 22.2325 11.9025 22.3675 ;
        RECT  11.2125 21.8425 11.2825 22.1325 ;
        RECT  11.1275 22.2325 11.1975 22.3675 ;
        RECT  11.0725 21.6925 11.9575 21.7575 ;
        RECT  11.8325 22.2325 11.9025 22.3675 ;
        RECT  11.8325 22.6975 11.9025 22.8975 ;
        RECT  11.1275 22.6975 11.1975 22.8975 ;
        RECT  11.7525 21.8425 11.8225 22.1325 ;
        RECT  11.2125 22.0675 11.3825 22.1325 ;
        RECT  11.8325 23.0275 11.8975 23.1625 ;
        RECT  11.6475 23.0275 11.7125 23.1625 ;
        RECT  11.1325 23.0275 11.1975 23.1625 ;
        RECT  11.3175 23.0275 11.3825 23.1625 ;
        RECT  11.6475 23.4925 11.7125 23.6275 ;
        RECT  11.8325 23.4925 11.8975 23.6275 ;
        RECT  11.3175 23.4925 11.3825 23.6275 ;
        RECT  11.1325 23.4925 11.1975 23.6275 ;
        RECT  11.7525 23.8825 11.8175 24.0175 ;
        RECT  11.5675 23.8825 11.6325 24.0175 ;
        RECT  11.3975 23.8825 11.4625 24.0175 ;
        RECT  11.2125 23.8825 11.2775 24.0175 ;
        RECT  11.835 23.39 11.9 23.525 ;
        RECT  11.835 23.39 11.9 23.525 ;
        RECT  11.835 23.39 11.9 23.525 ;
        RECT  11.835 23.39 11.9 23.525 ;
        RECT  11.835 23.39 11.9 23.525 ;
        RECT  11.835 23.39 11.9 23.525 ;
        RECT  11.4425 22.8975 11.5775 22.9625 ;
        RECT  11.095 24.2425 11.23 24.3075 ;
        RECT  11.8 24.2425 11.935 24.3075 ;
        RECT  11.43 24.1025 11.565 24.1675 ;
        RECT  11.835 23.39 11.9 23.525 ;
        RECT  11.835 23.39 11.9 23.525 ;
        RECT  11.835 23.39 11.9 23.525 ;
        RECT  11.835 23.39 11.9 23.525 ;
        RECT  11.335 23.2125 11.47 23.2775 ;
        RECT  11.335 23.2125 11.47 23.2775 ;
        RECT  11.56 23.3625 11.695 23.4275 ;
        RECT  11.56 23.3625 11.695 23.4275 ;
        RECT  11.835 23.39 11.9 23.525 ;
        RECT  11.835 23.39 11.9 23.525 ;
        RECT  11.835 23.39 11.9 23.525 ;
        RECT  11.835 23.39 11.9 23.525 ;
        RECT  11.385 23.8825 11.45 24.0175 ;
        RECT  11.13 23.39 11.195 23.525 ;
        RECT  11.13 23.39 11.195 23.525 ;
        RECT  11.13 23.39 11.195 23.525 ;
        RECT  11.13 23.39 11.195 23.525 ;
        RECT  11.13 23.39 11.195 23.525 ;
        RECT  11.13 23.39 11.195 23.525 ;
        RECT  11.835 23.39 11.9 23.525 ;
        RECT  11.835 23.39 11.9 23.525 ;
        RECT  11.835 23.39 11.9 23.525 ;
        RECT  11.835 23.39 11.9 23.525 ;
        RECT  11.58 23.8825 11.645 24.0175 ;
        RECT  11.4475 24.2425 11.5825 24.3075 ;
        RECT  11.4475 24.2425 11.5825 24.3075 ;
        RECT  11.8 24.2425 11.935 24.3075 ;
        RECT  11.4425 22.8975 11.5775 22.9625 ;
        RECT  11.8 24.2425 11.935 24.3075 ;
        RECT  11.8 24.2425 11.935 24.3075 ;
        RECT  11.835 23.39 11.9 23.525 ;
        RECT  11.835 23.39 11.9 23.525 ;
        RECT  11.835 23.39 11.9 23.525 ;
        RECT  11.835 23.39 11.9 23.525 ;
        RECT  11.835 23.39 11.9 23.525 ;
        RECT  11.835 23.39 11.9 23.525 ;
        RECT  11.095 24.2425 11.23 24.3075 ;
        RECT  11.455 22.9 11.555 22.9625 ;
        RECT  11.455 22.8975 11.555 22.96 ;
        RECT  11.7825 24.1025 11.835 24.165 ;
        RECT  11.455 22.9 11.555 22.9625 ;
        RECT  11.8325 22.9625 11.9025 23.1625 ;
        RECT  11.8325 23.4925 11.9025 23.6275 ;
        RECT  11.8325 23.4925 11.9025 23.6275 ;
        RECT  11.0725 24.2425 11.9575 24.3075 ;
        RECT  11.6475 23.7275 11.8225 23.7925 ;
        RECT  11.1275 23.4925 11.1975 23.6275 ;
        RECT  11.3175 23.0525 11.3825 23.7925 ;
        RECT  11.455 22.8975 11.555 22.96 ;
        RECT  11.0775 24.1025 11.13 24.165 ;
        RECT  11.8325 23.4925 11.9025 23.6275 ;
        RECT  11.0725 22.8975 11.9575 22.9625 ;
        RECT  11.6475 23.1625 11.7125 23.7925 ;
        RECT  11.8325 23.4925 11.9025 23.6275 ;
        RECT  11.8325 23.4925 11.9025 23.6275 ;
        RECT  11.2125 23.7275 11.2825 24.0175 ;
        RECT  11.1275 23.4925 11.1975 23.6275 ;
        RECT  11.0725 24.1025 11.9575 24.1675 ;
        RECT  11.8325 23.4925 11.9025 23.6275 ;
        RECT  11.8325 22.9625 11.9025 23.1625 ;
        RECT  11.1275 22.9625 11.1975 23.1625 ;
        RECT  11.7525 23.7275 11.8225 24.0175 ;
        RECT  11.2125 23.7275 11.3825 23.7925 ;
        RECT  11.8325 25.3875 11.8975 25.5225 ;
        RECT  11.6475 25.3875 11.7125 25.5225 ;
        RECT  11.1325 25.3875 11.1975 25.5225 ;
        RECT  11.3175 25.3875 11.3825 25.5225 ;
        RECT  11.6475 24.9225 11.7125 25.0575 ;
        RECT  11.8325 24.9225 11.8975 25.0575 ;
        RECT  11.3175 24.9225 11.3825 25.0575 ;
        RECT  11.1325 24.9225 11.1975 25.0575 ;
        RECT  11.7525 24.5325 11.8175 24.6675 ;
        RECT  11.5675 24.5325 11.6325 24.6675 ;
        RECT  11.3975 24.5325 11.4625 24.6675 ;
        RECT  11.2125 24.5325 11.2775 24.6675 ;
        RECT  11.835 25.025 11.9 25.16 ;
        RECT  11.835 25.025 11.9 25.16 ;
        RECT  11.835 25.025 11.9 25.16 ;
        RECT  11.835 25.025 11.9 25.16 ;
        RECT  11.835 25.025 11.9 25.16 ;
        RECT  11.835 25.025 11.9 25.16 ;
        RECT  11.4425 25.5875 11.5775 25.6525 ;
        RECT  11.095 24.2425 11.23 24.3075 ;
        RECT  11.8 24.2425 11.935 24.3075 ;
        RECT  11.43 24.3825 11.565 24.4475 ;
        RECT  11.835 25.025 11.9 25.16 ;
        RECT  11.835 25.025 11.9 25.16 ;
        RECT  11.835 25.025 11.9 25.16 ;
        RECT  11.835 25.025 11.9 25.16 ;
        RECT  11.335 25.2725 11.47 25.3375 ;
        RECT  11.335 25.2725 11.47 25.3375 ;
        RECT  11.56 25.1225 11.695 25.1875 ;
        RECT  11.56 25.1225 11.695 25.1875 ;
        RECT  11.835 25.025 11.9 25.16 ;
        RECT  11.835 25.025 11.9 25.16 ;
        RECT  11.835 25.025 11.9 25.16 ;
        RECT  11.835 25.025 11.9 25.16 ;
        RECT  11.385 24.5325 11.45 24.6675 ;
        RECT  11.13 25.025 11.195 25.16 ;
        RECT  11.13 25.025 11.195 25.16 ;
        RECT  11.13 25.025 11.195 25.16 ;
        RECT  11.13 25.025 11.195 25.16 ;
        RECT  11.13 25.025 11.195 25.16 ;
        RECT  11.13 25.025 11.195 25.16 ;
        RECT  11.835 25.025 11.9 25.16 ;
        RECT  11.835 25.025 11.9 25.16 ;
        RECT  11.835 25.025 11.9 25.16 ;
        RECT  11.835 25.025 11.9 25.16 ;
        RECT  11.58 24.5325 11.645 24.6675 ;
        RECT  11.4475 24.2425 11.5825 24.3075 ;
        RECT  11.4475 24.2425 11.5825 24.3075 ;
        RECT  11.8 24.2425 11.935 24.3075 ;
        RECT  11.4425 25.5875 11.5775 25.6525 ;
        RECT  11.8 24.2425 11.935 24.3075 ;
        RECT  11.8 24.2425 11.935 24.3075 ;
        RECT  11.835 25.025 11.9 25.16 ;
        RECT  11.835 25.025 11.9 25.16 ;
        RECT  11.835 25.025 11.9 25.16 ;
        RECT  11.835 25.025 11.9 25.16 ;
        RECT  11.835 25.025 11.9 25.16 ;
        RECT  11.835 25.025 11.9 25.16 ;
        RECT  11.095 24.2425 11.23 24.3075 ;
        RECT  11.455 25.5875 11.555 25.65 ;
        RECT  11.455 25.59 11.555 25.6525 ;
        RECT  11.7825 24.385 11.835 24.4475 ;
        RECT  11.455 25.5875 11.555 25.65 ;
        RECT  11.8325 25.3875 11.9025 25.5875 ;
        RECT  11.8325 24.9225 11.9025 25.0575 ;
        RECT  11.8325 24.9225 11.9025 25.0575 ;
        RECT  11.0725 24.2425 11.9575 24.3075 ;
        RECT  11.6475 24.7575 11.8225 24.8225 ;
        RECT  11.1275 24.9225 11.1975 25.0575 ;
        RECT  11.3175 24.7575 11.3825 25.4975 ;
        RECT  11.455 25.59 11.555 25.6525 ;
        RECT  11.0775 24.385 11.13 24.4475 ;
        RECT  11.8325 24.9225 11.9025 25.0575 ;
        RECT  11.0725 25.5875 11.9575 25.6525 ;
        RECT  11.6475 24.7575 11.7125 25.3875 ;
        RECT  11.8325 24.9225 11.9025 25.0575 ;
        RECT  11.8325 24.9225 11.9025 25.0575 ;
        RECT  11.2125 24.5325 11.2825 24.8225 ;
        RECT  11.1275 24.9225 11.1975 25.0575 ;
        RECT  11.0725 24.3825 11.9575 24.4475 ;
        RECT  11.8325 24.9225 11.9025 25.0575 ;
        RECT  11.8325 25.3875 11.9025 25.5875 ;
        RECT  11.1275 25.3875 11.1975 25.5875 ;
        RECT  11.7525 24.5325 11.8225 24.8225 ;
        RECT  11.2125 24.7575 11.3825 24.8225 ;
        RECT  11.8325 25.7175 11.8975 25.8525 ;
        RECT  11.6475 25.7175 11.7125 25.8525 ;
        RECT  11.1325 25.7175 11.1975 25.8525 ;
        RECT  11.3175 25.7175 11.3825 25.8525 ;
        RECT  11.6475 26.1825 11.7125 26.3175 ;
        RECT  11.8325 26.1825 11.8975 26.3175 ;
        RECT  11.3175 26.1825 11.3825 26.3175 ;
        RECT  11.1325 26.1825 11.1975 26.3175 ;
        RECT  11.7525 26.5725 11.8175 26.7075 ;
        RECT  11.5675 26.5725 11.6325 26.7075 ;
        RECT  11.3975 26.5725 11.4625 26.7075 ;
        RECT  11.2125 26.5725 11.2775 26.7075 ;
        RECT  11.835 26.08 11.9 26.215 ;
        RECT  11.835 26.08 11.9 26.215 ;
        RECT  11.835 26.08 11.9 26.215 ;
        RECT  11.835 26.08 11.9 26.215 ;
        RECT  11.835 26.08 11.9 26.215 ;
        RECT  11.835 26.08 11.9 26.215 ;
        RECT  11.4425 25.5875 11.5775 25.6525 ;
        RECT  11.095 26.9325 11.23 26.9975 ;
        RECT  11.8 26.9325 11.935 26.9975 ;
        RECT  11.43 26.7925 11.565 26.8575 ;
        RECT  11.835 26.08 11.9 26.215 ;
        RECT  11.835 26.08 11.9 26.215 ;
        RECT  11.835 26.08 11.9 26.215 ;
        RECT  11.835 26.08 11.9 26.215 ;
        RECT  11.335 25.9025 11.47 25.9675 ;
        RECT  11.335 25.9025 11.47 25.9675 ;
        RECT  11.56 26.0525 11.695 26.1175 ;
        RECT  11.56 26.0525 11.695 26.1175 ;
        RECT  11.835 26.08 11.9 26.215 ;
        RECT  11.835 26.08 11.9 26.215 ;
        RECT  11.835 26.08 11.9 26.215 ;
        RECT  11.835 26.08 11.9 26.215 ;
        RECT  11.385 26.5725 11.45 26.7075 ;
        RECT  11.13 26.08 11.195 26.215 ;
        RECT  11.13 26.08 11.195 26.215 ;
        RECT  11.13 26.08 11.195 26.215 ;
        RECT  11.13 26.08 11.195 26.215 ;
        RECT  11.13 26.08 11.195 26.215 ;
        RECT  11.13 26.08 11.195 26.215 ;
        RECT  11.835 26.08 11.9 26.215 ;
        RECT  11.835 26.08 11.9 26.215 ;
        RECT  11.835 26.08 11.9 26.215 ;
        RECT  11.835 26.08 11.9 26.215 ;
        RECT  11.58 26.5725 11.645 26.7075 ;
        RECT  11.4475 26.9325 11.5825 26.9975 ;
        RECT  11.4475 26.9325 11.5825 26.9975 ;
        RECT  11.8 26.9325 11.935 26.9975 ;
        RECT  11.4425 25.5875 11.5775 25.6525 ;
        RECT  11.8 26.9325 11.935 26.9975 ;
        RECT  11.8 26.9325 11.935 26.9975 ;
        RECT  11.835 26.08 11.9 26.215 ;
        RECT  11.835 26.08 11.9 26.215 ;
        RECT  11.835 26.08 11.9 26.215 ;
        RECT  11.835 26.08 11.9 26.215 ;
        RECT  11.835 26.08 11.9 26.215 ;
        RECT  11.835 26.08 11.9 26.215 ;
        RECT  11.095 26.9325 11.23 26.9975 ;
        RECT  11.455 25.59 11.555 25.6525 ;
        RECT  11.455 25.5875 11.555 25.65 ;
        RECT  11.7825 26.7925 11.835 26.855 ;
        RECT  11.455 25.59 11.555 25.6525 ;
        RECT  11.8325 25.6525 11.9025 25.8525 ;
        RECT  11.8325 26.1825 11.9025 26.3175 ;
        RECT  11.8325 26.1825 11.9025 26.3175 ;
        RECT  11.0725 26.9325 11.9575 26.9975 ;
        RECT  11.6475 26.4175 11.8225 26.4825 ;
        RECT  11.1275 26.1825 11.1975 26.3175 ;
        RECT  11.3175 25.7425 11.3825 26.4825 ;
        RECT  11.455 25.5875 11.555 25.65 ;
        RECT  11.0775 26.7925 11.13 26.855 ;
        RECT  11.8325 26.1825 11.9025 26.3175 ;
        RECT  11.0725 25.5875 11.9575 25.6525 ;
        RECT  11.6475 25.8525 11.7125 26.4825 ;
        RECT  11.8325 26.1825 11.9025 26.3175 ;
        RECT  11.8325 26.1825 11.9025 26.3175 ;
        RECT  11.2125 26.4175 11.2825 26.7075 ;
        RECT  11.1275 26.1825 11.1975 26.3175 ;
        RECT  11.0725 26.7925 11.9575 26.8575 ;
        RECT  11.8325 26.1825 11.9025 26.3175 ;
        RECT  11.8325 25.6525 11.9025 25.8525 ;
        RECT  11.1275 25.6525 11.1975 25.8525 ;
        RECT  11.7525 26.4175 11.8225 26.7075 ;
        RECT  11.2125 26.4175 11.3825 26.4825 ;
        RECT  11.8325 28.0775 11.8975 28.2125 ;
        RECT  11.6475 28.0775 11.7125 28.2125 ;
        RECT  11.1325 28.0775 11.1975 28.2125 ;
        RECT  11.3175 28.0775 11.3825 28.2125 ;
        RECT  11.6475 27.6125 11.7125 27.7475 ;
        RECT  11.8325 27.6125 11.8975 27.7475 ;
        RECT  11.3175 27.6125 11.3825 27.7475 ;
        RECT  11.1325 27.6125 11.1975 27.7475 ;
        RECT  11.7525 27.2225 11.8175 27.3575 ;
        RECT  11.5675 27.2225 11.6325 27.3575 ;
        RECT  11.3975 27.2225 11.4625 27.3575 ;
        RECT  11.2125 27.2225 11.2775 27.3575 ;
        RECT  11.835 27.715 11.9 27.85 ;
        RECT  11.835 27.715 11.9 27.85 ;
        RECT  11.835 27.715 11.9 27.85 ;
        RECT  11.835 27.715 11.9 27.85 ;
        RECT  11.835 27.715 11.9 27.85 ;
        RECT  11.835 27.715 11.9 27.85 ;
        RECT  11.4425 28.2775 11.5775 28.3425 ;
        RECT  11.095 26.9325 11.23 26.9975 ;
        RECT  11.8 26.9325 11.935 26.9975 ;
        RECT  11.43 27.0725 11.565 27.1375 ;
        RECT  11.835 27.715 11.9 27.85 ;
        RECT  11.835 27.715 11.9 27.85 ;
        RECT  11.835 27.715 11.9 27.85 ;
        RECT  11.835 27.715 11.9 27.85 ;
        RECT  11.335 27.9625 11.47 28.0275 ;
        RECT  11.335 27.9625 11.47 28.0275 ;
        RECT  11.56 27.8125 11.695 27.8775 ;
        RECT  11.56 27.8125 11.695 27.8775 ;
        RECT  11.835 27.715 11.9 27.85 ;
        RECT  11.835 27.715 11.9 27.85 ;
        RECT  11.835 27.715 11.9 27.85 ;
        RECT  11.835 27.715 11.9 27.85 ;
        RECT  11.385 27.2225 11.45 27.3575 ;
        RECT  11.13 27.715 11.195 27.85 ;
        RECT  11.13 27.715 11.195 27.85 ;
        RECT  11.13 27.715 11.195 27.85 ;
        RECT  11.13 27.715 11.195 27.85 ;
        RECT  11.13 27.715 11.195 27.85 ;
        RECT  11.13 27.715 11.195 27.85 ;
        RECT  11.835 27.715 11.9 27.85 ;
        RECT  11.835 27.715 11.9 27.85 ;
        RECT  11.835 27.715 11.9 27.85 ;
        RECT  11.835 27.715 11.9 27.85 ;
        RECT  11.58 27.2225 11.645 27.3575 ;
        RECT  11.4475 26.9325 11.5825 26.9975 ;
        RECT  11.4475 26.9325 11.5825 26.9975 ;
        RECT  11.8 26.9325 11.935 26.9975 ;
        RECT  11.4425 28.2775 11.5775 28.3425 ;
        RECT  11.8 26.9325 11.935 26.9975 ;
        RECT  11.8 26.9325 11.935 26.9975 ;
        RECT  11.835 27.715 11.9 27.85 ;
        RECT  11.835 27.715 11.9 27.85 ;
        RECT  11.835 27.715 11.9 27.85 ;
        RECT  11.835 27.715 11.9 27.85 ;
        RECT  11.835 27.715 11.9 27.85 ;
        RECT  11.835 27.715 11.9 27.85 ;
        RECT  11.095 26.9325 11.23 26.9975 ;
        RECT  11.455 28.2775 11.555 28.34 ;
        RECT  11.455 28.28 11.555 28.3425 ;
        RECT  11.7825 27.075 11.835 27.1375 ;
        RECT  11.455 28.2775 11.555 28.34 ;
        RECT  11.8325 28.0775 11.9025 28.2775 ;
        RECT  11.8325 27.6125 11.9025 27.7475 ;
        RECT  11.8325 27.6125 11.9025 27.7475 ;
        RECT  11.0725 26.9325 11.9575 26.9975 ;
        RECT  11.6475 27.4475 11.8225 27.5125 ;
        RECT  11.1275 27.6125 11.1975 27.7475 ;
        RECT  11.3175 27.4475 11.3825 28.1875 ;
        RECT  11.455 28.28 11.555 28.3425 ;
        RECT  11.0775 27.075 11.13 27.1375 ;
        RECT  11.8325 27.6125 11.9025 27.7475 ;
        RECT  11.0725 28.2775 11.9575 28.3425 ;
        RECT  11.6475 27.4475 11.7125 28.0775 ;
        RECT  11.8325 27.6125 11.9025 27.7475 ;
        RECT  11.8325 27.6125 11.9025 27.7475 ;
        RECT  11.2125 27.2225 11.2825 27.5125 ;
        RECT  11.1275 27.6125 11.1975 27.7475 ;
        RECT  11.0725 27.0725 11.9575 27.1375 ;
        RECT  11.8325 27.6125 11.9025 27.7475 ;
        RECT  11.8325 28.0775 11.9025 28.2775 ;
        RECT  11.1275 28.0775 11.1975 28.2775 ;
        RECT  11.7525 27.2225 11.8225 27.5125 ;
        RECT  11.2125 27.4475 11.3825 27.5125 ;
        RECT  11.8325 28.4075 11.8975 28.5425 ;
        RECT  11.6475 28.4075 11.7125 28.5425 ;
        RECT  11.1325 28.4075 11.1975 28.5425 ;
        RECT  11.3175 28.4075 11.3825 28.5425 ;
        RECT  11.6475 28.8725 11.7125 29.0075 ;
        RECT  11.8325 28.8725 11.8975 29.0075 ;
        RECT  11.3175 28.8725 11.3825 29.0075 ;
        RECT  11.1325 28.8725 11.1975 29.0075 ;
        RECT  11.7525 29.2625 11.8175 29.3975 ;
        RECT  11.5675 29.2625 11.6325 29.3975 ;
        RECT  11.3975 29.2625 11.4625 29.3975 ;
        RECT  11.2125 29.2625 11.2775 29.3975 ;
        RECT  11.835 28.77 11.9 28.905 ;
        RECT  11.835 28.77 11.9 28.905 ;
        RECT  11.835 28.77 11.9 28.905 ;
        RECT  11.835 28.77 11.9 28.905 ;
        RECT  11.835 28.77 11.9 28.905 ;
        RECT  11.835 28.77 11.9 28.905 ;
        RECT  11.4425 28.2775 11.5775 28.3425 ;
        RECT  11.095 29.6225 11.23 29.6875 ;
        RECT  11.8 29.6225 11.935 29.6875 ;
        RECT  11.43 29.4825 11.565 29.5475 ;
        RECT  11.835 28.77 11.9 28.905 ;
        RECT  11.835 28.77 11.9 28.905 ;
        RECT  11.835 28.77 11.9 28.905 ;
        RECT  11.835 28.77 11.9 28.905 ;
        RECT  11.335 28.5925 11.47 28.6575 ;
        RECT  11.335 28.5925 11.47 28.6575 ;
        RECT  11.56 28.7425 11.695 28.8075 ;
        RECT  11.56 28.7425 11.695 28.8075 ;
        RECT  11.835 28.77 11.9 28.905 ;
        RECT  11.835 28.77 11.9 28.905 ;
        RECT  11.835 28.77 11.9 28.905 ;
        RECT  11.835 28.77 11.9 28.905 ;
        RECT  11.385 29.2625 11.45 29.3975 ;
        RECT  11.13 28.77 11.195 28.905 ;
        RECT  11.13 28.77 11.195 28.905 ;
        RECT  11.13 28.77 11.195 28.905 ;
        RECT  11.13 28.77 11.195 28.905 ;
        RECT  11.13 28.77 11.195 28.905 ;
        RECT  11.13 28.77 11.195 28.905 ;
        RECT  11.835 28.77 11.9 28.905 ;
        RECT  11.835 28.77 11.9 28.905 ;
        RECT  11.835 28.77 11.9 28.905 ;
        RECT  11.835 28.77 11.9 28.905 ;
        RECT  11.58 29.2625 11.645 29.3975 ;
        RECT  11.4475 29.6225 11.5825 29.6875 ;
        RECT  11.4475 29.6225 11.5825 29.6875 ;
        RECT  11.8 29.6225 11.935 29.6875 ;
        RECT  11.4425 28.2775 11.5775 28.3425 ;
        RECT  11.8 29.6225 11.935 29.6875 ;
        RECT  11.8 29.6225 11.935 29.6875 ;
        RECT  11.835 28.77 11.9 28.905 ;
        RECT  11.835 28.77 11.9 28.905 ;
        RECT  11.835 28.77 11.9 28.905 ;
        RECT  11.835 28.77 11.9 28.905 ;
        RECT  11.835 28.77 11.9 28.905 ;
        RECT  11.835 28.77 11.9 28.905 ;
        RECT  11.095 29.6225 11.23 29.6875 ;
        RECT  11.455 28.28 11.555 28.3425 ;
        RECT  11.455 28.2775 11.555 28.34 ;
        RECT  11.7825 29.4825 11.835 29.545 ;
        RECT  11.455 28.28 11.555 28.3425 ;
        RECT  11.8325 28.3425 11.9025 28.5425 ;
        RECT  11.8325 28.8725 11.9025 29.0075 ;
        RECT  11.8325 28.8725 11.9025 29.0075 ;
        RECT  11.0725 29.6225 11.9575 29.6875 ;
        RECT  11.6475 29.1075 11.8225 29.1725 ;
        RECT  11.1275 28.8725 11.1975 29.0075 ;
        RECT  11.3175 28.4325 11.3825 29.1725 ;
        RECT  11.455 28.2775 11.555 28.34 ;
        RECT  11.0775 29.4825 11.13 29.545 ;
        RECT  11.8325 28.8725 11.9025 29.0075 ;
        RECT  11.0725 28.2775 11.9575 28.3425 ;
        RECT  11.6475 28.5425 11.7125 29.1725 ;
        RECT  11.8325 28.8725 11.9025 29.0075 ;
        RECT  11.8325 28.8725 11.9025 29.0075 ;
        RECT  11.2125 29.1075 11.2825 29.3975 ;
        RECT  11.1275 28.8725 11.1975 29.0075 ;
        RECT  11.0725 29.4825 11.9575 29.5475 ;
        RECT  11.8325 28.8725 11.9025 29.0075 ;
        RECT  11.8325 28.3425 11.9025 28.5425 ;
        RECT  11.1275 28.3425 11.1975 28.5425 ;
        RECT  11.7525 29.1075 11.8225 29.3975 ;
        RECT  11.2125 29.1075 11.3825 29.1725 ;
        RECT  11.8325 30.7675 11.8975 30.9025 ;
        RECT  11.6475 30.7675 11.7125 30.9025 ;
        RECT  11.1325 30.7675 11.1975 30.9025 ;
        RECT  11.3175 30.7675 11.3825 30.9025 ;
        RECT  11.6475 30.3025 11.7125 30.4375 ;
        RECT  11.8325 30.3025 11.8975 30.4375 ;
        RECT  11.3175 30.3025 11.3825 30.4375 ;
        RECT  11.1325 30.3025 11.1975 30.4375 ;
        RECT  11.7525 29.9125 11.8175 30.0475 ;
        RECT  11.5675 29.9125 11.6325 30.0475 ;
        RECT  11.3975 29.9125 11.4625 30.0475 ;
        RECT  11.2125 29.9125 11.2775 30.0475 ;
        RECT  11.835 30.405 11.9 30.54 ;
        RECT  11.835 30.405 11.9 30.54 ;
        RECT  11.835 30.405 11.9 30.54 ;
        RECT  11.835 30.405 11.9 30.54 ;
        RECT  11.835 30.405 11.9 30.54 ;
        RECT  11.835 30.405 11.9 30.54 ;
        RECT  11.4425 30.9675 11.5775 31.0325 ;
        RECT  11.095 29.6225 11.23 29.6875 ;
        RECT  11.8 29.6225 11.935 29.6875 ;
        RECT  11.43 29.7625 11.565 29.8275 ;
        RECT  11.835 30.405 11.9 30.54 ;
        RECT  11.835 30.405 11.9 30.54 ;
        RECT  11.835 30.405 11.9 30.54 ;
        RECT  11.835 30.405 11.9 30.54 ;
        RECT  11.335 30.6525 11.47 30.7175 ;
        RECT  11.335 30.6525 11.47 30.7175 ;
        RECT  11.56 30.5025 11.695 30.5675 ;
        RECT  11.56 30.5025 11.695 30.5675 ;
        RECT  11.835 30.405 11.9 30.54 ;
        RECT  11.835 30.405 11.9 30.54 ;
        RECT  11.835 30.405 11.9 30.54 ;
        RECT  11.835 30.405 11.9 30.54 ;
        RECT  11.385 29.9125 11.45 30.0475 ;
        RECT  11.13 30.405 11.195 30.54 ;
        RECT  11.13 30.405 11.195 30.54 ;
        RECT  11.13 30.405 11.195 30.54 ;
        RECT  11.13 30.405 11.195 30.54 ;
        RECT  11.13 30.405 11.195 30.54 ;
        RECT  11.13 30.405 11.195 30.54 ;
        RECT  11.835 30.405 11.9 30.54 ;
        RECT  11.835 30.405 11.9 30.54 ;
        RECT  11.835 30.405 11.9 30.54 ;
        RECT  11.835 30.405 11.9 30.54 ;
        RECT  11.58 29.9125 11.645 30.0475 ;
        RECT  11.4475 29.6225 11.5825 29.6875 ;
        RECT  11.4475 29.6225 11.5825 29.6875 ;
        RECT  11.8 29.6225 11.935 29.6875 ;
        RECT  11.4425 30.9675 11.5775 31.0325 ;
        RECT  11.8 29.6225 11.935 29.6875 ;
        RECT  11.8 29.6225 11.935 29.6875 ;
        RECT  11.835 30.405 11.9 30.54 ;
        RECT  11.835 30.405 11.9 30.54 ;
        RECT  11.835 30.405 11.9 30.54 ;
        RECT  11.835 30.405 11.9 30.54 ;
        RECT  11.835 30.405 11.9 30.54 ;
        RECT  11.835 30.405 11.9 30.54 ;
        RECT  11.095 29.6225 11.23 29.6875 ;
        RECT  11.455 30.9675 11.555 31.03 ;
        RECT  11.455 30.97 11.555 31.0325 ;
        RECT  11.7825 29.765 11.835 29.8275 ;
        RECT  11.455 30.9675 11.555 31.03 ;
        RECT  11.8325 30.7675 11.9025 30.9675 ;
        RECT  11.8325 30.3025 11.9025 30.4375 ;
        RECT  11.8325 30.3025 11.9025 30.4375 ;
        RECT  11.0725 29.6225 11.9575 29.6875 ;
        RECT  11.6475 30.1375 11.8225 30.2025 ;
        RECT  11.1275 30.3025 11.1975 30.4375 ;
        RECT  11.3175 30.1375 11.3825 30.8775 ;
        RECT  11.455 30.97 11.555 31.0325 ;
        RECT  11.0775 29.765 11.13 29.8275 ;
        RECT  11.8325 30.3025 11.9025 30.4375 ;
        RECT  11.0725 30.9675 11.9575 31.0325 ;
        RECT  11.6475 30.1375 11.7125 30.7675 ;
        RECT  11.8325 30.3025 11.9025 30.4375 ;
        RECT  11.8325 30.3025 11.9025 30.4375 ;
        RECT  11.2125 29.9125 11.2825 30.2025 ;
        RECT  11.1275 30.3025 11.1975 30.4375 ;
        RECT  11.0725 29.7625 11.9575 29.8275 ;
        RECT  11.8325 30.3025 11.9025 30.4375 ;
        RECT  11.8325 30.7675 11.9025 30.9675 ;
        RECT  11.1275 30.7675 11.1975 30.9675 ;
        RECT  11.7525 29.9125 11.8225 30.2025 ;
        RECT  11.2125 30.1375 11.3825 30.2025 ;
        RECT  11.8325 31.0975 11.8975 31.2325 ;
        RECT  11.6475 31.0975 11.7125 31.2325 ;
        RECT  11.1325 31.0975 11.1975 31.2325 ;
        RECT  11.3175 31.0975 11.3825 31.2325 ;
        RECT  11.6475 31.5625 11.7125 31.6975 ;
        RECT  11.8325 31.5625 11.8975 31.6975 ;
        RECT  11.3175 31.5625 11.3825 31.6975 ;
        RECT  11.1325 31.5625 11.1975 31.6975 ;
        RECT  11.7525 31.9525 11.8175 32.0875 ;
        RECT  11.5675 31.9525 11.6325 32.0875 ;
        RECT  11.3975 31.9525 11.4625 32.0875 ;
        RECT  11.2125 31.9525 11.2775 32.0875 ;
        RECT  11.835 31.46 11.9 31.595 ;
        RECT  11.835 31.46 11.9 31.595 ;
        RECT  11.835 31.46 11.9 31.595 ;
        RECT  11.835 31.46 11.9 31.595 ;
        RECT  11.835 31.46 11.9 31.595 ;
        RECT  11.835 31.46 11.9 31.595 ;
        RECT  11.4425 30.9675 11.5775 31.0325 ;
        RECT  11.095 32.3125 11.23 32.3775 ;
        RECT  11.8 32.3125 11.935 32.3775 ;
        RECT  11.43 32.1725 11.565 32.2375 ;
        RECT  11.835 31.46 11.9 31.595 ;
        RECT  11.835 31.46 11.9 31.595 ;
        RECT  11.835 31.46 11.9 31.595 ;
        RECT  11.835 31.46 11.9 31.595 ;
        RECT  11.335 31.2825 11.47 31.3475 ;
        RECT  11.335 31.2825 11.47 31.3475 ;
        RECT  11.56 31.4325 11.695 31.4975 ;
        RECT  11.56 31.4325 11.695 31.4975 ;
        RECT  11.835 31.46 11.9 31.595 ;
        RECT  11.835 31.46 11.9 31.595 ;
        RECT  11.835 31.46 11.9 31.595 ;
        RECT  11.835 31.46 11.9 31.595 ;
        RECT  11.385 31.9525 11.45 32.0875 ;
        RECT  11.13 31.46 11.195 31.595 ;
        RECT  11.13 31.46 11.195 31.595 ;
        RECT  11.13 31.46 11.195 31.595 ;
        RECT  11.13 31.46 11.195 31.595 ;
        RECT  11.13 31.46 11.195 31.595 ;
        RECT  11.13 31.46 11.195 31.595 ;
        RECT  11.835 31.46 11.9 31.595 ;
        RECT  11.835 31.46 11.9 31.595 ;
        RECT  11.835 31.46 11.9 31.595 ;
        RECT  11.835 31.46 11.9 31.595 ;
        RECT  11.58 31.9525 11.645 32.0875 ;
        RECT  11.4475 32.3125 11.5825 32.3775 ;
        RECT  11.4475 32.3125 11.5825 32.3775 ;
        RECT  11.8 32.3125 11.935 32.3775 ;
        RECT  11.4425 30.9675 11.5775 31.0325 ;
        RECT  11.8 32.3125 11.935 32.3775 ;
        RECT  11.8 32.3125 11.935 32.3775 ;
        RECT  11.835 31.46 11.9 31.595 ;
        RECT  11.835 31.46 11.9 31.595 ;
        RECT  11.835 31.46 11.9 31.595 ;
        RECT  11.835 31.46 11.9 31.595 ;
        RECT  11.835 31.46 11.9 31.595 ;
        RECT  11.835 31.46 11.9 31.595 ;
        RECT  11.095 32.3125 11.23 32.3775 ;
        RECT  11.455 30.97 11.555 31.0325 ;
        RECT  11.455 30.9675 11.555 31.03 ;
        RECT  11.7825 32.1725 11.835 32.235 ;
        RECT  11.455 30.97 11.555 31.0325 ;
        RECT  11.8325 31.0325 11.9025 31.2325 ;
        RECT  11.8325 31.5625 11.9025 31.6975 ;
        RECT  11.8325 31.5625 11.9025 31.6975 ;
        RECT  11.0725 32.3125 11.9575 32.3775 ;
        RECT  11.6475 31.7975 11.8225 31.8625 ;
        RECT  11.1275 31.5625 11.1975 31.6975 ;
        RECT  11.3175 31.1225 11.3825 31.8625 ;
        RECT  11.455 30.9675 11.555 31.03 ;
        RECT  11.0775 32.1725 11.13 32.235 ;
        RECT  11.8325 31.5625 11.9025 31.6975 ;
        RECT  11.0725 30.9675 11.9575 31.0325 ;
        RECT  11.6475 31.2325 11.7125 31.8625 ;
        RECT  11.8325 31.5625 11.9025 31.6975 ;
        RECT  11.8325 31.5625 11.9025 31.6975 ;
        RECT  11.2125 31.7975 11.2825 32.0875 ;
        RECT  11.1275 31.5625 11.1975 31.6975 ;
        RECT  11.0725 32.1725 11.9575 32.2375 ;
        RECT  11.8325 31.5625 11.9025 31.6975 ;
        RECT  11.8325 31.0325 11.9025 31.2325 ;
        RECT  11.1275 31.0325 11.1975 31.2325 ;
        RECT  11.7525 31.7975 11.8225 32.0875 ;
        RECT  11.2125 31.7975 11.3825 31.8625 ;
        RECT  11.8325 33.4575 11.8975 33.5925 ;
        RECT  11.6475 33.4575 11.7125 33.5925 ;
        RECT  11.1325 33.4575 11.1975 33.5925 ;
        RECT  11.3175 33.4575 11.3825 33.5925 ;
        RECT  11.6475 32.9925 11.7125 33.1275 ;
        RECT  11.8325 32.9925 11.8975 33.1275 ;
        RECT  11.3175 32.9925 11.3825 33.1275 ;
        RECT  11.1325 32.9925 11.1975 33.1275 ;
        RECT  11.7525 32.6025 11.8175 32.7375 ;
        RECT  11.5675 32.6025 11.6325 32.7375 ;
        RECT  11.3975 32.6025 11.4625 32.7375 ;
        RECT  11.2125 32.6025 11.2775 32.7375 ;
        RECT  11.835 33.095 11.9 33.23 ;
        RECT  11.835 33.095 11.9 33.23 ;
        RECT  11.835 33.095 11.9 33.23 ;
        RECT  11.835 33.095 11.9 33.23 ;
        RECT  11.835 33.095 11.9 33.23 ;
        RECT  11.835 33.095 11.9 33.23 ;
        RECT  11.4425 33.6575 11.5775 33.7225 ;
        RECT  11.095 32.3125 11.23 32.3775 ;
        RECT  11.8 32.3125 11.935 32.3775 ;
        RECT  11.43 32.4525 11.565 32.5175 ;
        RECT  11.835 33.095 11.9 33.23 ;
        RECT  11.835 33.095 11.9 33.23 ;
        RECT  11.835 33.095 11.9 33.23 ;
        RECT  11.835 33.095 11.9 33.23 ;
        RECT  11.335 33.3425 11.47 33.4075 ;
        RECT  11.335 33.3425 11.47 33.4075 ;
        RECT  11.56 33.1925 11.695 33.2575 ;
        RECT  11.56 33.1925 11.695 33.2575 ;
        RECT  11.835 33.095 11.9 33.23 ;
        RECT  11.835 33.095 11.9 33.23 ;
        RECT  11.835 33.095 11.9 33.23 ;
        RECT  11.835 33.095 11.9 33.23 ;
        RECT  11.385 32.6025 11.45 32.7375 ;
        RECT  11.13 33.095 11.195 33.23 ;
        RECT  11.13 33.095 11.195 33.23 ;
        RECT  11.13 33.095 11.195 33.23 ;
        RECT  11.13 33.095 11.195 33.23 ;
        RECT  11.13 33.095 11.195 33.23 ;
        RECT  11.13 33.095 11.195 33.23 ;
        RECT  11.835 33.095 11.9 33.23 ;
        RECT  11.835 33.095 11.9 33.23 ;
        RECT  11.835 33.095 11.9 33.23 ;
        RECT  11.835 33.095 11.9 33.23 ;
        RECT  11.58 32.6025 11.645 32.7375 ;
        RECT  11.4475 32.3125 11.5825 32.3775 ;
        RECT  11.4475 32.3125 11.5825 32.3775 ;
        RECT  11.8 32.3125 11.935 32.3775 ;
        RECT  11.4425 33.6575 11.5775 33.7225 ;
        RECT  11.8 32.3125 11.935 32.3775 ;
        RECT  11.8 32.3125 11.935 32.3775 ;
        RECT  11.835 33.095 11.9 33.23 ;
        RECT  11.835 33.095 11.9 33.23 ;
        RECT  11.835 33.095 11.9 33.23 ;
        RECT  11.835 33.095 11.9 33.23 ;
        RECT  11.835 33.095 11.9 33.23 ;
        RECT  11.835 33.095 11.9 33.23 ;
        RECT  11.095 32.3125 11.23 32.3775 ;
        RECT  11.455 33.6575 11.555 33.72 ;
        RECT  11.455 33.66 11.555 33.7225 ;
        RECT  11.7825 32.455 11.835 32.5175 ;
        RECT  11.455 33.6575 11.555 33.72 ;
        RECT  11.8325 33.4575 11.9025 33.6575 ;
        RECT  11.8325 32.9925 11.9025 33.1275 ;
        RECT  11.8325 32.9925 11.9025 33.1275 ;
        RECT  11.0725 32.3125 11.9575 32.3775 ;
        RECT  11.6475 32.8275 11.8225 32.8925 ;
        RECT  11.1275 32.9925 11.1975 33.1275 ;
        RECT  11.3175 32.8275 11.3825 33.5675 ;
        RECT  11.455 33.66 11.555 33.7225 ;
        RECT  11.0775 32.455 11.13 32.5175 ;
        RECT  11.8325 32.9925 11.9025 33.1275 ;
        RECT  11.0725 33.6575 11.9575 33.7225 ;
        RECT  11.6475 32.8275 11.7125 33.4575 ;
        RECT  11.8325 32.9925 11.9025 33.1275 ;
        RECT  11.8325 32.9925 11.9025 33.1275 ;
        RECT  11.2125 32.6025 11.2825 32.8925 ;
        RECT  11.1275 32.9925 11.1975 33.1275 ;
        RECT  11.0725 32.4525 11.9575 32.5175 ;
        RECT  11.8325 32.9925 11.9025 33.1275 ;
        RECT  11.8325 33.4575 11.9025 33.6575 ;
        RECT  11.1275 33.4575 11.1975 33.6575 ;
        RECT  11.7525 32.6025 11.8225 32.8925 ;
        RECT  11.2125 32.8275 11.3825 32.8925 ;
        RECT  11.8325 33.7875 11.8975 33.9225 ;
        RECT  11.6475 33.7875 11.7125 33.9225 ;
        RECT  11.1325 33.7875 11.1975 33.9225 ;
        RECT  11.3175 33.7875 11.3825 33.9225 ;
        RECT  11.6475 34.2525 11.7125 34.3875 ;
        RECT  11.8325 34.2525 11.8975 34.3875 ;
        RECT  11.3175 34.2525 11.3825 34.3875 ;
        RECT  11.1325 34.2525 11.1975 34.3875 ;
        RECT  11.7525 34.6425 11.8175 34.7775 ;
        RECT  11.5675 34.6425 11.6325 34.7775 ;
        RECT  11.3975 34.6425 11.4625 34.7775 ;
        RECT  11.2125 34.6425 11.2775 34.7775 ;
        RECT  11.835 34.15 11.9 34.285 ;
        RECT  11.835 34.15 11.9 34.285 ;
        RECT  11.835 34.15 11.9 34.285 ;
        RECT  11.835 34.15 11.9 34.285 ;
        RECT  11.835 34.15 11.9 34.285 ;
        RECT  11.835 34.15 11.9 34.285 ;
        RECT  11.4425 33.6575 11.5775 33.7225 ;
        RECT  11.095 35.0025 11.23 35.0675 ;
        RECT  11.8 35.0025 11.935 35.0675 ;
        RECT  11.43 34.8625 11.565 34.9275 ;
        RECT  11.835 34.15 11.9 34.285 ;
        RECT  11.835 34.15 11.9 34.285 ;
        RECT  11.835 34.15 11.9 34.285 ;
        RECT  11.835 34.15 11.9 34.285 ;
        RECT  11.335 33.9725 11.47 34.0375 ;
        RECT  11.335 33.9725 11.47 34.0375 ;
        RECT  11.56 34.1225 11.695 34.1875 ;
        RECT  11.56 34.1225 11.695 34.1875 ;
        RECT  11.835 34.15 11.9 34.285 ;
        RECT  11.835 34.15 11.9 34.285 ;
        RECT  11.835 34.15 11.9 34.285 ;
        RECT  11.835 34.15 11.9 34.285 ;
        RECT  11.385 34.6425 11.45 34.7775 ;
        RECT  11.13 34.15 11.195 34.285 ;
        RECT  11.13 34.15 11.195 34.285 ;
        RECT  11.13 34.15 11.195 34.285 ;
        RECT  11.13 34.15 11.195 34.285 ;
        RECT  11.13 34.15 11.195 34.285 ;
        RECT  11.13 34.15 11.195 34.285 ;
        RECT  11.835 34.15 11.9 34.285 ;
        RECT  11.835 34.15 11.9 34.285 ;
        RECT  11.835 34.15 11.9 34.285 ;
        RECT  11.835 34.15 11.9 34.285 ;
        RECT  11.58 34.6425 11.645 34.7775 ;
        RECT  11.4475 35.0025 11.5825 35.0675 ;
        RECT  11.4475 35.0025 11.5825 35.0675 ;
        RECT  11.8 35.0025 11.935 35.0675 ;
        RECT  11.4425 33.6575 11.5775 33.7225 ;
        RECT  11.8 35.0025 11.935 35.0675 ;
        RECT  11.8 35.0025 11.935 35.0675 ;
        RECT  11.835 34.15 11.9 34.285 ;
        RECT  11.835 34.15 11.9 34.285 ;
        RECT  11.835 34.15 11.9 34.285 ;
        RECT  11.835 34.15 11.9 34.285 ;
        RECT  11.835 34.15 11.9 34.285 ;
        RECT  11.835 34.15 11.9 34.285 ;
        RECT  11.095 35.0025 11.23 35.0675 ;
        RECT  11.455 33.66 11.555 33.7225 ;
        RECT  11.455 33.6575 11.555 33.72 ;
        RECT  11.7825 34.8625 11.835 34.925 ;
        RECT  11.455 33.66 11.555 33.7225 ;
        RECT  11.8325 33.7225 11.9025 33.9225 ;
        RECT  11.8325 34.2525 11.9025 34.3875 ;
        RECT  11.8325 34.2525 11.9025 34.3875 ;
        RECT  11.0725 35.0025 11.9575 35.0675 ;
        RECT  11.6475 34.4875 11.8225 34.5525 ;
        RECT  11.1275 34.2525 11.1975 34.3875 ;
        RECT  11.3175 33.8125 11.3825 34.5525 ;
        RECT  11.455 33.6575 11.555 33.72 ;
        RECT  11.0775 34.8625 11.13 34.925 ;
        RECT  11.8325 34.2525 11.9025 34.3875 ;
        RECT  11.0725 33.6575 11.9575 33.7225 ;
        RECT  11.6475 33.9225 11.7125 34.5525 ;
        RECT  11.8325 34.2525 11.9025 34.3875 ;
        RECT  11.8325 34.2525 11.9025 34.3875 ;
        RECT  11.2125 34.4875 11.2825 34.7775 ;
        RECT  11.1275 34.2525 11.1975 34.3875 ;
        RECT  11.0725 34.8625 11.9575 34.9275 ;
        RECT  11.8325 34.2525 11.9025 34.3875 ;
        RECT  11.8325 33.7225 11.9025 33.9225 ;
        RECT  11.1275 33.7225 11.1975 33.9225 ;
        RECT  11.7525 34.4875 11.8225 34.7775 ;
        RECT  11.2125 34.4875 11.3825 34.5525 ;
        RECT  11.8325 36.1475 11.8975 36.2825 ;
        RECT  11.6475 36.1475 11.7125 36.2825 ;
        RECT  11.1325 36.1475 11.1975 36.2825 ;
        RECT  11.3175 36.1475 11.3825 36.2825 ;
        RECT  11.6475 35.6825 11.7125 35.8175 ;
        RECT  11.8325 35.6825 11.8975 35.8175 ;
        RECT  11.3175 35.6825 11.3825 35.8175 ;
        RECT  11.1325 35.6825 11.1975 35.8175 ;
        RECT  11.7525 35.2925 11.8175 35.4275 ;
        RECT  11.5675 35.2925 11.6325 35.4275 ;
        RECT  11.3975 35.2925 11.4625 35.4275 ;
        RECT  11.2125 35.2925 11.2775 35.4275 ;
        RECT  11.835 35.785 11.9 35.92 ;
        RECT  11.835 35.785 11.9 35.92 ;
        RECT  11.835 35.785 11.9 35.92 ;
        RECT  11.835 35.785 11.9 35.92 ;
        RECT  11.835 35.785 11.9 35.92 ;
        RECT  11.835 35.785 11.9 35.92 ;
        RECT  11.4425 36.3475 11.5775 36.4125 ;
        RECT  11.095 35.0025 11.23 35.0675 ;
        RECT  11.8 35.0025 11.935 35.0675 ;
        RECT  11.43 35.1425 11.565 35.2075 ;
        RECT  11.835 35.785 11.9 35.92 ;
        RECT  11.835 35.785 11.9 35.92 ;
        RECT  11.835 35.785 11.9 35.92 ;
        RECT  11.835 35.785 11.9 35.92 ;
        RECT  11.335 36.0325 11.47 36.0975 ;
        RECT  11.335 36.0325 11.47 36.0975 ;
        RECT  11.56 35.8825 11.695 35.9475 ;
        RECT  11.56 35.8825 11.695 35.9475 ;
        RECT  11.835 35.785 11.9 35.92 ;
        RECT  11.835 35.785 11.9 35.92 ;
        RECT  11.835 35.785 11.9 35.92 ;
        RECT  11.835 35.785 11.9 35.92 ;
        RECT  11.385 35.2925 11.45 35.4275 ;
        RECT  11.13 35.785 11.195 35.92 ;
        RECT  11.13 35.785 11.195 35.92 ;
        RECT  11.13 35.785 11.195 35.92 ;
        RECT  11.13 35.785 11.195 35.92 ;
        RECT  11.13 35.785 11.195 35.92 ;
        RECT  11.13 35.785 11.195 35.92 ;
        RECT  11.835 35.785 11.9 35.92 ;
        RECT  11.835 35.785 11.9 35.92 ;
        RECT  11.835 35.785 11.9 35.92 ;
        RECT  11.835 35.785 11.9 35.92 ;
        RECT  11.58 35.2925 11.645 35.4275 ;
        RECT  11.4475 35.0025 11.5825 35.0675 ;
        RECT  11.4475 35.0025 11.5825 35.0675 ;
        RECT  11.8 35.0025 11.935 35.0675 ;
        RECT  11.4425 36.3475 11.5775 36.4125 ;
        RECT  11.8 35.0025 11.935 35.0675 ;
        RECT  11.8 35.0025 11.935 35.0675 ;
        RECT  11.835 35.785 11.9 35.92 ;
        RECT  11.835 35.785 11.9 35.92 ;
        RECT  11.835 35.785 11.9 35.92 ;
        RECT  11.835 35.785 11.9 35.92 ;
        RECT  11.835 35.785 11.9 35.92 ;
        RECT  11.835 35.785 11.9 35.92 ;
        RECT  11.095 35.0025 11.23 35.0675 ;
        RECT  11.455 36.3475 11.555 36.41 ;
        RECT  11.455 36.35 11.555 36.4125 ;
        RECT  11.7825 35.145 11.835 35.2075 ;
        RECT  11.455 36.3475 11.555 36.41 ;
        RECT  11.8325 36.1475 11.9025 36.3475 ;
        RECT  11.8325 35.6825 11.9025 35.8175 ;
        RECT  11.8325 35.6825 11.9025 35.8175 ;
        RECT  11.0725 35.0025 11.9575 35.0675 ;
        RECT  11.6475 35.5175 11.8225 35.5825 ;
        RECT  11.1275 35.6825 11.1975 35.8175 ;
        RECT  11.3175 35.5175 11.3825 36.2575 ;
        RECT  11.455 36.35 11.555 36.4125 ;
        RECT  11.0775 35.145 11.13 35.2075 ;
        RECT  11.8325 35.6825 11.9025 35.8175 ;
        RECT  11.0725 36.3475 11.9575 36.4125 ;
        RECT  11.6475 35.5175 11.7125 36.1475 ;
        RECT  11.8325 35.6825 11.9025 35.8175 ;
        RECT  11.8325 35.6825 11.9025 35.8175 ;
        RECT  11.2125 35.2925 11.2825 35.5825 ;
        RECT  11.1275 35.6825 11.1975 35.8175 ;
        RECT  11.0725 35.1425 11.9575 35.2075 ;
        RECT  11.8325 35.6825 11.9025 35.8175 ;
        RECT  11.8325 36.1475 11.9025 36.3475 ;
        RECT  11.1275 36.1475 11.1975 36.3475 ;
        RECT  11.7525 35.2925 11.8225 35.5825 ;
        RECT  11.2125 35.5175 11.3825 35.5825 ;
        RECT  11.8325 36.4775 11.8975 36.6125 ;
        RECT  11.6475 36.4775 11.7125 36.6125 ;
        RECT  11.1325 36.4775 11.1975 36.6125 ;
        RECT  11.3175 36.4775 11.3825 36.6125 ;
        RECT  11.6475 36.9425 11.7125 37.0775 ;
        RECT  11.8325 36.9425 11.8975 37.0775 ;
        RECT  11.3175 36.9425 11.3825 37.0775 ;
        RECT  11.1325 36.9425 11.1975 37.0775 ;
        RECT  11.7525 37.3325 11.8175 37.4675 ;
        RECT  11.5675 37.3325 11.6325 37.4675 ;
        RECT  11.3975 37.3325 11.4625 37.4675 ;
        RECT  11.2125 37.3325 11.2775 37.4675 ;
        RECT  11.835 36.84 11.9 36.975 ;
        RECT  11.835 36.84 11.9 36.975 ;
        RECT  11.835 36.84 11.9 36.975 ;
        RECT  11.835 36.84 11.9 36.975 ;
        RECT  11.835 36.84 11.9 36.975 ;
        RECT  11.835 36.84 11.9 36.975 ;
        RECT  11.4425 36.3475 11.5775 36.4125 ;
        RECT  11.095 37.6925 11.23 37.7575 ;
        RECT  11.8 37.6925 11.935 37.7575 ;
        RECT  11.43 37.5525 11.565 37.6175 ;
        RECT  11.835 36.84 11.9 36.975 ;
        RECT  11.835 36.84 11.9 36.975 ;
        RECT  11.835 36.84 11.9 36.975 ;
        RECT  11.835 36.84 11.9 36.975 ;
        RECT  11.335 36.6625 11.47 36.7275 ;
        RECT  11.335 36.6625 11.47 36.7275 ;
        RECT  11.56 36.8125 11.695 36.8775 ;
        RECT  11.56 36.8125 11.695 36.8775 ;
        RECT  11.835 36.84 11.9 36.975 ;
        RECT  11.835 36.84 11.9 36.975 ;
        RECT  11.835 36.84 11.9 36.975 ;
        RECT  11.835 36.84 11.9 36.975 ;
        RECT  11.385 37.3325 11.45 37.4675 ;
        RECT  11.13 36.84 11.195 36.975 ;
        RECT  11.13 36.84 11.195 36.975 ;
        RECT  11.13 36.84 11.195 36.975 ;
        RECT  11.13 36.84 11.195 36.975 ;
        RECT  11.13 36.84 11.195 36.975 ;
        RECT  11.13 36.84 11.195 36.975 ;
        RECT  11.835 36.84 11.9 36.975 ;
        RECT  11.835 36.84 11.9 36.975 ;
        RECT  11.835 36.84 11.9 36.975 ;
        RECT  11.835 36.84 11.9 36.975 ;
        RECT  11.58 37.3325 11.645 37.4675 ;
        RECT  11.4475 37.6925 11.5825 37.7575 ;
        RECT  11.4475 37.6925 11.5825 37.7575 ;
        RECT  11.8 37.6925 11.935 37.7575 ;
        RECT  11.4425 36.3475 11.5775 36.4125 ;
        RECT  11.8 37.6925 11.935 37.7575 ;
        RECT  11.8 37.6925 11.935 37.7575 ;
        RECT  11.835 36.84 11.9 36.975 ;
        RECT  11.835 36.84 11.9 36.975 ;
        RECT  11.835 36.84 11.9 36.975 ;
        RECT  11.835 36.84 11.9 36.975 ;
        RECT  11.835 36.84 11.9 36.975 ;
        RECT  11.835 36.84 11.9 36.975 ;
        RECT  11.095 37.6925 11.23 37.7575 ;
        RECT  11.455 36.35 11.555 36.4125 ;
        RECT  11.455 36.3475 11.555 36.41 ;
        RECT  11.7825 37.5525 11.835 37.615 ;
        RECT  11.455 36.35 11.555 36.4125 ;
        RECT  11.8325 36.4125 11.9025 36.6125 ;
        RECT  11.8325 36.9425 11.9025 37.0775 ;
        RECT  11.8325 36.9425 11.9025 37.0775 ;
        RECT  11.0725 37.6925 11.9575 37.7575 ;
        RECT  11.6475 37.1775 11.8225 37.2425 ;
        RECT  11.1275 36.9425 11.1975 37.0775 ;
        RECT  11.3175 36.5025 11.3825 37.2425 ;
        RECT  11.455 36.3475 11.555 36.41 ;
        RECT  11.0775 37.5525 11.13 37.615 ;
        RECT  11.8325 36.9425 11.9025 37.0775 ;
        RECT  11.0725 36.3475 11.9575 36.4125 ;
        RECT  11.6475 36.6125 11.7125 37.2425 ;
        RECT  11.8325 36.9425 11.9025 37.0775 ;
        RECT  11.8325 36.9425 11.9025 37.0775 ;
        RECT  11.2125 37.1775 11.2825 37.4675 ;
        RECT  11.1275 36.9425 11.1975 37.0775 ;
        RECT  11.0725 37.5525 11.9575 37.6175 ;
        RECT  11.8325 36.9425 11.9025 37.0775 ;
        RECT  11.8325 36.4125 11.9025 36.6125 ;
        RECT  11.1275 36.4125 11.1975 36.6125 ;
        RECT  11.7525 37.1775 11.8225 37.4675 ;
        RECT  11.2125 37.1775 11.3825 37.2425 ;
        RECT  11.8325 38.8375 11.8975 38.9725 ;
        RECT  11.6475 38.8375 11.7125 38.9725 ;
        RECT  11.1325 38.8375 11.1975 38.9725 ;
        RECT  11.3175 38.8375 11.3825 38.9725 ;
        RECT  11.6475 38.3725 11.7125 38.5075 ;
        RECT  11.8325 38.3725 11.8975 38.5075 ;
        RECT  11.3175 38.3725 11.3825 38.5075 ;
        RECT  11.1325 38.3725 11.1975 38.5075 ;
        RECT  11.7525 37.9825 11.8175 38.1175 ;
        RECT  11.5675 37.9825 11.6325 38.1175 ;
        RECT  11.3975 37.9825 11.4625 38.1175 ;
        RECT  11.2125 37.9825 11.2775 38.1175 ;
        RECT  11.835 38.475 11.9 38.61 ;
        RECT  11.835 38.475 11.9 38.61 ;
        RECT  11.835 38.475 11.9 38.61 ;
        RECT  11.835 38.475 11.9 38.61 ;
        RECT  11.835 38.475 11.9 38.61 ;
        RECT  11.835 38.475 11.9 38.61 ;
        RECT  11.4425 39.0375 11.5775 39.1025 ;
        RECT  11.095 37.6925 11.23 37.7575 ;
        RECT  11.8 37.6925 11.935 37.7575 ;
        RECT  11.43 37.8325 11.565 37.8975 ;
        RECT  11.835 38.475 11.9 38.61 ;
        RECT  11.835 38.475 11.9 38.61 ;
        RECT  11.835 38.475 11.9 38.61 ;
        RECT  11.835 38.475 11.9 38.61 ;
        RECT  11.335 38.7225 11.47 38.7875 ;
        RECT  11.335 38.7225 11.47 38.7875 ;
        RECT  11.56 38.5725 11.695 38.6375 ;
        RECT  11.56 38.5725 11.695 38.6375 ;
        RECT  11.835 38.475 11.9 38.61 ;
        RECT  11.835 38.475 11.9 38.61 ;
        RECT  11.835 38.475 11.9 38.61 ;
        RECT  11.835 38.475 11.9 38.61 ;
        RECT  11.385 37.9825 11.45 38.1175 ;
        RECT  11.13 38.475 11.195 38.61 ;
        RECT  11.13 38.475 11.195 38.61 ;
        RECT  11.13 38.475 11.195 38.61 ;
        RECT  11.13 38.475 11.195 38.61 ;
        RECT  11.13 38.475 11.195 38.61 ;
        RECT  11.13 38.475 11.195 38.61 ;
        RECT  11.835 38.475 11.9 38.61 ;
        RECT  11.835 38.475 11.9 38.61 ;
        RECT  11.835 38.475 11.9 38.61 ;
        RECT  11.835 38.475 11.9 38.61 ;
        RECT  11.58 37.9825 11.645 38.1175 ;
        RECT  11.4475 37.6925 11.5825 37.7575 ;
        RECT  11.4475 37.6925 11.5825 37.7575 ;
        RECT  11.8 37.6925 11.935 37.7575 ;
        RECT  11.4425 39.0375 11.5775 39.1025 ;
        RECT  11.8 37.6925 11.935 37.7575 ;
        RECT  11.8 37.6925 11.935 37.7575 ;
        RECT  11.835 38.475 11.9 38.61 ;
        RECT  11.835 38.475 11.9 38.61 ;
        RECT  11.835 38.475 11.9 38.61 ;
        RECT  11.835 38.475 11.9 38.61 ;
        RECT  11.835 38.475 11.9 38.61 ;
        RECT  11.835 38.475 11.9 38.61 ;
        RECT  11.095 37.6925 11.23 37.7575 ;
        RECT  11.455 39.0375 11.555 39.1 ;
        RECT  11.455 39.04 11.555 39.1025 ;
        RECT  11.7825 37.835 11.835 37.8975 ;
        RECT  11.455 39.0375 11.555 39.1 ;
        RECT  11.8325 38.8375 11.9025 39.0375 ;
        RECT  11.8325 38.3725 11.9025 38.5075 ;
        RECT  11.8325 38.3725 11.9025 38.5075 ;
        RECT  11.0725 37.6925 11.9575 37.7575 ;
        RECT  11.6475 38.2075 11.8225 38.2725 ;
        RECT  11.1275 38.3725 11.1975 38.5075 ;
        RECT  11.3175 38.2075 11.3825 38.9475 ;
        RECT  11.455 39.04 11.555 39.1025 ;
        RECT  11.0775 37.835 11.13 37.8975 ;
        RECT  11.8325 38.3725 11.9025 38.5075 ;
        RECT  11.0725 39.0375 11.9575 39.1025 ;
        RECT  11.6475 38.2075 11.7125 38.8375 ;
        RECT  11.8325 38.3725 11.9025 38.5075 ;
        RECT  11.8325 38.3725 11.9025 38.5075 ;
        RECT  11.2125 37.9825 11.2825 38.2725 ;
        RECT  11.1275 38.3725 11.1975 38.5075 ;
        RECT  11.0725 37.8325 11.9575 37.8975 ;
        RECT  11.8325 38.3725 11.9025 38.5075 ;
        RECT  11.8325 38.8375 11.9025 39.0375 ;
        RECT  11.1275 38.8375 11.1975 39.0375 ;
        RECT  11.7525 37.9825 11.8225 38.2725 ;
        RECT  11.2125 38.2075 11.3825 38.2725 ;
        RECT  11.8325 39.1675 11.8975 39.3025 ;
        RECT  11.6475 39.1675 11.7125 39.3025 ;
        RECT  11.1325 39.1675 11.1975 39.3025 ;
        RECT  11.3175 39.1675 11.3825 39.3025 ;
        RECT  11.6475 39.6325 11.7125 39.7675 ;
        RECT  11.8325 39.6325 11.8975 39.7675 ;
        RECT  11.3175 39.6325 11.3825 39.7675 ;
        RECT  11.1325 39.6325 11.1975 39.7675 ;
        RECT  11.7525 40.0225 11.8175 40.1575 ;
        RECT  11.5675 40.0225 11.6325 40.1575 ;
        RECT  11.3975 40.0225 11.4625 40.1575 ;
        RECT  11.2125 40.0225 11.2775 40.1575 ;
        RECT  11.835 39.53 11.9 39.665 ;
        RECT  11.835 39.53 11.9 39.665 ;
        RECT  11.835 39.53 11.9 39.665 ;
        RECT  11.835 39.53 11.9 39.665 ;
        RECT  11.835 39.53 11.9 39.665 ;
        RECT  11.835 39.53 11.9 39.665 ;
        RECT  11.4425 39.0375 11.5775 39.1025 ;
        RECT  11.095 40.3825 11.23 40.4475 ;
        RECT  11.8 40.3825 11.935 40.4475 ;
        RECT  11.43 40.2425 11.565 40.3075 ;
        RECT  11.835 39.53 11.9 39.665 ;
        RECT  11.835 39.53 11.9 39.665 ;
        RECT  11.835 39.53 11.9 39.665 ;
        RECT  11.835 39.53 11.9 39.665 ;
        RECT  11.335 39.3525 11.47 39.4175 ;
        RECT  11.335 39.3525 11.47 39.4175 ;
        RECT  11.56 39.5025 11.695 39.5675 ;
        RECT  11.56 39.5025 11.695 39.5675 ;
        RECT  11.835 39.53 11.9 39.665 ;
        RECT  11.835 39.53 11.9 39.665 ;
        RECT  11.835 39.53 11.9 39.665 ;
        RECT  11.835 39.53 11.9 39.665 ;
        RECT  11.385 40.0225 11.45 40.1575 ;
        RECT  11.13 39.53 11.195 39.665 ;
        RECT  11.13 39.53 11.195 39.665 ;
        RECT  11.13 39.53 11.195 39.665 ;
        RECT  11.13 39.53 11.195 39.665 ;
        RECT  11.13 39.53 11.195 39.665 ;
        RECT  11.13 39.53 11.195 39.665 ;
        RECT  11.835 39.53 11.9 39.665 ;
        RECT  11.835 39.53 11.9 39.665 ;
        RECT  11.835 39.53 11.9 39.665 ;
        RECT  11.835 39.53 11.9 39.665 ;
        RECT  11.58 40.0225 11.645 40.1575 ;
        RECT  11.4475 40.3825 11.5825 40.4475 ;
        RECT  11.4475 40.3825 11.5825 40.4475 ;
        RECT  11.8 40.3825 11.935 40.4475 ;
        RECT  11.4425 39.0375 11.5775 39.1025 ;
        RECT  11.8 40.3825 11.935 40.4475 ;
        RECT  11.8 40.3825 11.935 40.4475 ;
        RECT  11.835 39.53 11.9 39.665 ;
        RECT  11.835 39.53 11.9 39.665 ;
        RECT  11.835 39.53 11.9 39.665 ;
        RECT  11.835 39.53 11.9 39.665 ;
        RECT  11.835 39.53 11.9 39.665 ;
        RECT  11.835 39.53 11.9 39.665 ;
        RECT  11.095 40.3825 11.23 40.4475 ;
        RECT  11.455 39.04 11.555 39.1025 ;
        RECT  11.455 39.0375 11.555 39.1 ;
        RECT  11.7825 40.2425 11.835 40.305 ;
        RECT  11.455 39.04 11.555 39.1025 ;
        RECT  11.8325 39.1025 11.9025 39.3025 ;
        RECT  11.8325 39.6325 11.9025 39.7675 ;
        RECT  11.8325 39.6325 11.9025 39.7675 ;
        RECT  11.0725 40.3825 11.9575 40.4475 ;
        RECT  11.6475 39.8675 11.8225 39.9325 ;
        RECT  11.1275 39.6325 11.1975 39.7675 ;
        RECT  11.3175 39.1925 11.3825 39.9325 ;
        RECT  11.455 39.0375 11.555 39.1 ;
        RECT  11.0775 40.2425 11.13 40.305 ;
        RECT  11.8325 39.6325 11.9025 39.7675 ;
        RECT  11.0725 39.0375 11.9575 39.1025 ;
        RECT  11.6475 39.3025 11.7125 39.9325 ;
        RECT  11.8325 39.6325 11.9025 39.7675 ;
        RECT  11.8325 39.6325 11.9025 39.7675 ;
        RECT  11.2125 39.8675 11.2825 40.1575 ;
        RECT  11.1275 39.6325 11.1975 39.7675 ;
        RECT  11.0725 40.2425 11.9575 40.3075 ;
        RECT  11.8325 39.6325 11.9025 39.7675 ;
        RECT  11.8325 39.1025 11.9025 39.3025 ;
        RECT  11.1275 39.1025 11.1975 39.3025 ;
        RECT  11.7525 39.8675 11.8225 40.1575 ;
        RECT  11.2125 39.8675 11.3825 39.9325 ;
        RECT  12.5375 20.0075 12.6025 20.1425 ;
        RECT  12.3525 20.0075 12.4175 20.1425 ;
        RECT  11.8375 20.0075 11.9025 20.1425 ;
        RECT  12.0225 20.0075 12.0875 20.1425 ;
        RECT  12.3525 19.5425 12.4175 19.6775 ;
        RECT  12.5375 19.5425 12.6025 19.6775 ;
        RECT  12.0225 19.5425 12.0875 19.6775 ;
        RECT  11.8375 19.5425 11.9025 19.6775 ;
        RECT  12.4575 19.1525 12.5225 19.2875 ;
        RECT  12.2725 19.1525 12.3375 19.2875 ;
        RECT  12.1025 19.1525 12.1675 19.2875 ;
        RECT  11.9175 19.1525 11.9825 19.2875 ;
        RECT  12.54 19.645 12.605 19.78 ;
        RECT  12.54 19.645 12.605 19.78 ;
        RECT  12.54 19.645 12.605 19.78 ;
        RECT  12.54 19.645 12.605 19.78 ;
        RECT  12.54 19.645 12.605 19.78 ;
        RECT  12.54 19.645 12.605 19.78 ;
        RECT  12.1475 20.2075 12.2825 20.2725 ;
        RECT  11.8 18.8625 11.935 18.9275 ;
        RECT  12.505 18.8625 12.64 18.9275 ;
        RECT  12.135 19.0025 12.27 19.0675 ;
        RECT  12.54 19.645 12.605 19.78 ;
        RECT  12.54 19.645 12.605 19.78 ;
        RECT  12.54 19.645 12.605 19.78 ;
        RECT  12.54 19.645 12.605 19.78 ;
        RECT  12.04 19.8925 12.175 19.9575 ;
        RECT  12.04 19.8925 12.175 19.9575 ;
        RECT  12.265 19.7425 12.4 19.8075 ;
        RECT  12.265 19.7425 12.4 19.8075 ;
        RECT  12.54 19.645 12.605 19.78 ;
        RECT  12.54 19.645 12.605 19.78 ;
        RECT  12.54 19.645 12.605 19.78 ;
        RECT  12.54 19.645 12.605 19.78 ;
        RECT  12.09 19.1525 12.155 19.2875 ;
        RECT  11.835 19.645 11.9 19.78 ;
        RECT  11.835 19.645 11.9 19.78 ;
        RECT  11.835 19.645 11.9 19.78 ;
        RECT  11.835 19.645 11.9 19.78 ;
        RECT  11.835 19.645 11.9 19.78 ;
        RECT  11.835 19.645 11.9 19.78 ;
        RECT  12.54 19.645 12.605 19.78 ;
        RECT  12.54 19.645 12.605 19.78 ;
        RECT  12.54 19.645 12.605 19.78 ;
        RECT  12.54 19.645 12.605 19.78 ;
        RECT  12.285 19.1525 12.35 19.2875 ;
        RECT  12.1525 18.8625 12.2875 18.9275 ;
        RECT  12.1525 18.8625 12.2875 18.9275 ;
        RECT  12.505 18.8625 12.64 18.9275 ;
        RECT  12.1475 20.2075 12.2825 20.2725 ;
        RECT  12.505 18.8625 12.64 18.9275 ;
        RECT  12.505 18.8625 12.64 18.9275 ;
        RECT  12.54 19.645 12.605 19.78 ;
        RECT  12.54 19.645 12.605 19.78 ;
        RECT  12.54 19.645 12.605 19.78 ;
        RECT  12.54 19.645 12.605 19.78 ;
        RECT  12.54 19.645 12.605 19.78 ;
        RECT  12.54 19.645 12.605 19.78 ;
        RECT  11.8 18.8625 11.935 18.9275 ;
        RECT  12.16 20.2075 12.26 20.27 ;
        RECT  12.16 20.21 12.26 20.2725 ;
        RECT  12.4875 19.005 12.54 19.0675 ;
        RECT  12.16 20.2075 12.26 20.27 ;
        RECT  12.5375 20.0075 12.6075 20.2075 ;
        RECT  12.5375 19.5425 12.6075 19.6775 ;
        RECT  12.5375 19.5425 12.6075 19.6775 ;
        RECT  11.7775 18.8625 12.6625 18.9275 ;
        RECT  12.3525 19.3775 12.5275 19.4425 ;
        RECT  11.8325 19.5425 11.9025 19.6775 ;
        RECT  12.0225 19.3775 12.0875 20.1175 ;
        RECT  12.16 20.21 12.26 20.2725 ;
        RECT  11.7825 19.005 11.835 19.0675 ;
        RECT  12.5375 19.5425 12.6075 19.6775 ;
        RECT  11.7775 20.2075 12.6625 20.2725 ;
        RECT  12.3525 19.3775 12.4175 20.0075 ;
        RECT  12.5375 19.5425 12.6075 19.6775 ;
        RECT  12.5375 19.5425 12.6075 19.6775 ;
        RECT  11.9175 19.1525 11.9875 19.4425 ;
        RECT  11.8325 19.5425 11.9025 19.6775 ;
        RECT  11.7775 19.0025 12.6625 19.0675 ;
        RECT  12.5375 19.5425 12.6075 19.6775 ;
        RECT  12.5375 20.0075 12.6075 20.2075 ;
        RECT  11.8325 20.0075 11.9025 20.2075 ;
        RECT  12.4575 19.1525 12.5275 19.4425 ;
        RECT  11.9175 19.3775 12.0875 19.4425 ;
        RECT  12.5375 20.3375 12.6025 20.4725 ;
        RECT  12.3525 20.3375 12.4175 20.4725 ;
        RECT  11.8375 20.3375 11.9025 20.4725 ;
        RECT  12.0225 20.3375 12.0875 20.4725 ;
        RECT  12.3525 20.8025 12.4175 20.9375 ;
        RECT  12.5375 20.8025 12.6025 20.9375 ;
        RECT  12.0225 20.8025 12.0875 20.9375 ;
        RECT  11.8375 20.8025 11.9025 20.9375 ;
        RECT  12.4575 21.1925 12.5225 21.3275 ;
        RECT  12.2725 21.1925 12.3375 21.3275 ;
        RECT  12.1025 21.1925 12.1675 21.3275 ;
        RECT  11.9175 21.1925 11.9825 21.3275 ;
        RECT  12.54 20.7 12.605 20.835 ;
        RECT  12.54 20.7 12.605 20.835 ;
        RECT  12.54 20.7 12.605 20.835 ;
        RECT  12.54 20.7 12.605 20.835 ;
        RECT  12.54 20.7 12.605 20.835 ;
        RECT  12.54 20.7 12.605 20.835 ;
        RECT  12.1475 20.2075 12.2825 20.2725 ;
        RECT  11.8 21.5525 11.935 21.6175 ;
        RECT  12.505 21.5525 12.64 21.6175 ;
        RECT  12.135 21.4125 12.27 21.4775 ;
        RECT  12.54 20.7 12.605 20.835 ;
        RECT  12.54 20.7 12.605 20.835 ;
        RECT  12.54 20.7 12.605 20.835 ;
        RECT  12.54 20.7 12.605 20.835 ;
        RECT  12.04 20.5225 12.175 20.5875 ;
        RECT  12.04 20.5225 12.175 20.5875 ;
        RECT  12.265 20.6725 12.4 20.7375 ;
        RECT  12.265 20.6725 12.4 20.7375 ;
        RECT  12.54 20.7 12.605 20.835 ;
        RECT  12.54 20.7 12.605 20.835 ;
        RECT  12.54 20.7 12.605 20.835 ;
        RECT  12.54 20.7 12.605 20.835 ;
        RECT  12.09 21.1925 12.155 21.3275 ;
        RECT  11.835 20.7 11.9 20.835 ;
        RECT  11.835 20.7 11.9 20.835 ;
        RECT  11.835 20.7 11.9 20.835 ;
        RECT  11.835 20.7 11.9 20.835 ;
        RECT  11.835 20.7 11.9 20.835 ;
        RECT  11.835 20.7 11.9 20.835 ;
        RECT  12.54 20.7 12.605 20.835 ;
        RECT  12.54 20.7 12.605 20.835 ;
        RECT  12.54 20.7 12.605 20.835 ;
        RECT  12.54 20.7 12.605 20.835 ;
        RECT  12.285 21.1925 12.35 21.3275 ;
        RECT  12.1525 21.5525 12.2875 21.6175 ;
        RECT  12.1525 21.5525 12.2875 21.6175 ;
        RECT  12.505 21.5525 12.64 21.6175 ;
        RECT  12.1475 20.2075 12.2825 20.2725 ;
        RECT  12.505 21.5525 12.64 21.6175 ;
        RECT  12.505 21.5525 12.64 21.6175 ;
        RECT  12.54 20.7 12.605 20.835 ;
        RECT  12.54 20.7 12.605 20.835 ;
        RECT  12.54 20.7 12.605 20.835 ;
        RECT  12.54 20.7 12.605 20.835 ;
        RECT  12.54 20.7 12.605 20.835 ;
        RECT  12.54 20.7 12.605 20.835 ;
        RECT  11.8 21.5525 11.935 21.6175 ;
        RECT  12.16 20.21 12.26 20.2725 ;
        RECT  12.16 20.2075 12.26 20.27 ;
        RECT  12.4875 21.4125 12.54 21.475 ;
        RECT  12.16 20.21 12.26 20.2725 ;
        RECT  12.5375 20.2725 12.6075 20.4725 ;
        RECT  12.5375 20.8025 12.6075 20.9375 ;
        RECT  12.5375 20.8025 12.6075 20.9375 ;
        RECT  11.7775 21.5525 12.6625 21.6175 ;
        RECT  12.3525 21.0375 12.5275 21.1025 ;
        RECT  11.8325 20.8025 11.9025 20.9375 ;
        RECT  12.0225 20.3625 12.0875 21.1025 ;
        RECT  12.16 20.2075 12.26 20.27 ;
        RECT  11.7825 21.4125 11.835 21.475 ;
        RECT  12.5375 20.8025 12.6075 20.9375 ;
        RECT  11.7775 20.2075 12.6625 20.2725 ;
        RECT  12.3525 20.4725 12.4175 21.1025 ;
        RECT  12.5375 20.8025 12.6075 20.9375 ;
        RECT  12.5375 20.8025 12.6075 20.9375 ;
        RECT  11.9175 21.0375 11.9875 21.3275 ;
        RECT  11.8325 20.8025 11.9025 20.9375 ;
        RECT  11.7775 21.4125 12.6625 21.4775 ;
        RECT  12.5375 20.8025 12.6075 20.9375 ;
        RECT  12.5375 20.2725 12.6075 20.4725 ;
        RECT  11.8325 20.2725 11.9025 20.4725 ;
        RECT  12.4575 21.0375 12.5275 21.3275 ;
        RECT  11.9175 21.0375 12.0875 21.1025 ;
        RECT  12.5375 22.6975 12.6025 22.8325 ;
        RECT  12.3525 22.6975 12.4175 22.8325 ;
        RECT  11.8375 22.6975 11.9025 22.8325 ;
        RECT  12.0225 22.6975 12.0875 22.8325 ;
        RECT  12.3525 22.2325 12.4175 22.3675 ;
        RECT  12.5375 22.2325 12.6025 22.3675 ;
        RECT  12.0225 22.2325 12.0875 22.3675 ;
        RECT  11.8375 22.2325 11.9025 22.3675 ;
        RECT  12.4575 21.8425 12.5225 21.9775 ;
        RECT  12.2725 21.8425 12.3375 21.9775 ;
        RECT  12.1025 21.8425 12.1675 21.9775 ;
        RECT  11.9175 21.8425 11.9825 21.9775 ;
        RECT  12.54 22.335 12.605 22.47 ;
        RECT  12.54 22.335 12.605 22.47 ;
        RECT  12.54 22.335 12.605 22.47 ;
        RECT  12.54 22.335 12.605 22.47 ;
        RECT  12.54 22.335 12.605 22.47 ;
        RECT  12.54 22.335 12.605 22.47 ;
        RECT  12.1475 22.8975 12.2825 22.9625 ;
        RECT  11.8 21.5525 11.935 21.6175 ;
        RECT  12.505 21.5525 12.64 21.6175 ;
        RECT  12.135 21.6925 12.27 21.7575 ;
        RECT  12.54 22.335 12.605 22.47 ;
        RECT  12.54 22.335 12.605 22.47 ;
        RECT  12.54 22.335 12.605 22.47 ;
        RECT  12.54 22.335 12.605 22.47 ;
        RECT  12.04 22.5825 12.175 22.6475 ;
        RECT  12.04 22.5825 12.175 22.6475 ;
        RECT  12.265 22.4325 12.4 22.4975 ;
        RECT  12.265 22.4325 12.4 22.4975 ;
        RECT  12.54 22.335 12.605 22.47 ;
        RECT  12.54 22.335 12.605 22.47 ;
        RECT  12.54 22.335 12.605 22.47 ;
        RECT  12.54 22.335 12.605 22.47 ;
        RECT  12.09 21.8425 12.155 21.9775 ;
        RECT  11.835 22.335 11.9 22.47 ;
        RECT  11.835 22.335 11.9 22.47 ;
        RECT  11.835 22.335 11.9 22.47 ;
        RECT  11.835 22.335 11.9 22.47 ;
        RECT  11.835 22.335 11.9 22.47 ;
        RECT  11.835 22.335 11.9 22.47 ;
        RECT  12.54 22.335 12.605 22.47 ;
        RECT  12.54 22.335 12.605 22.47 ;
        RECT  12.54 22.335 12.605 22.47 ;
        RECT  12.54 22.335 12.605 22.47 ;
        RECT  12.285 21.8425 12.35 21.9775 ;
        RECT  12.1525 21.5525 12.2875 21.6175 ;
        RECT  12.1525 21.5525 12.2875 21.6175 ;
        RECT  12.505 21.5525 12.64 21.6175 ;
        RECT  12.1475 22.8975 12.2825 22.9625 ;
        RECT  12.505 21.5525 12.64 21.6175 ;
        RECT  12.505 21.5525 12.64 21.6175 ;
        RECT  12.54 22.335 12.605 22.47 ;
        RECT  12.54 22.335 12.605 22.47 ;
        RECT  12.54 22.335 12.605 22.47 ;
        RECT  12.54 22.335 12.605 22.47 ;
        RECT  12.54 22.335 12.605 22.47 ;
        RECT  12.54 22.335 12.605 22.47 ;
        RECT  11.8 21.5525 11.935 21.6175 ;
        RECT  12.16 22.8975 12.26 22.96 ;
        RECT  12.16 22.9 12.26 22.9625 ;
        RECT  12.4875 21.695 12.54 21.7575 ;
        RECT  12.16 22.8975 12.26 22.96 ;
        RECT  12.5375 22.6975 12.6075 22.8975 ;
        RECT  12.5375 22.2325 12.6075 22.3675 ;
        RECT  12.5375 22.2325 12.6075 22.3675 ;
        RECT  11.7775 21.5525 12.6625 21.6175 ;
        RECT  12.3525 22.0675 12.5275 22.1325 ;
        RECT  11.8325 22.2325 11.9025 22.3675 ;
        RECT  12.0225 22.0675 12.0875 22.8075 ;
        RECT  12.16 22.9 12.26 22.9625 ;
        RECT  11.7825 21.695 11.835 21.7575 ;
        RECT  12.5375 22.2325 12.6075 22.3675 ;
        RECT  11.7775 22.8975 12.6625 22.9625 ;
        RECT  12.3525 22.0675 12.4175 22.6975 ;
        RECT  12.5375 22.2325 12.6075 22.3675 ;
        RECT  12.5375 22.2325 12.6075 22.3675 ;
        RECT  11.9175 21.8425 11.9875 22.1325 ;
        RECT  11.8325 22.2325 11.9025 22.3675 ;
        RECT  11.7775 21.6925 12.6625 21.7575 ;
        RECT  12.5375 22.2325 12.6075 22.3675 ;
        RECT  12.5375 22.6975 12.6075 22.8975 ;
        RECT  11.8325 22.6975 11.9025 22.8975 ;
        RECT  12.4575 21.8425 12.5275 22.1325 ;
        RECT  11.9175 22.0675 12.0875 22.1325 ;
        RECT  12.5375 23.0275 12.6025 23.1625 ;
        RECT  12.3525 23.0275 12.4175 23.1625 ;
        RECT  11.8375 23.0275 11.9025 23.1625 ;
        RECT  12.0225 23.0275 12.0875 23.1625 ;
        RECT  12.3525 23.4925 12.4175 23.6275 ;
        RECT  12.5375 23.4925 12.6025 23.6275 ;
        RECT  12.0225 23.4925 12.0875 23.6275 ;
        RECT  11.8375 23.4925 11.9025 23.6275 ;
        RECT  12.4575 23.8825 12.5225 24.0175 ;
        RECT  12.2725 23.8825 12.3375 24.0175 ;
        RECT  12.1025 23.8825 12.1675 24.0175 ;
        RECT  11.9175 23.8825 11.9825 24.0175 ;
        RECT  12.54 23.39 12.605 23.525 ;
        RECT  12.54 23.39 12.605 23.525 ;
        RECT  12.54 23.39 12.605 23.525 ;
        RECT  12.54 23.39 12.605 23.525 ;
        RECT  12.54 23.39 12.605 23.525 ;
        RECT  12.54 23.39 12.605 23.525 ;
        RECT  12.1475 22.8975 12.2825 22.9625 ;
        RECT  11.8 24.2425 11.935 24.3075 ;
        RECT  12.505 24.2425 12.64 24.3075 ;
        RECT  12.135 24.1025 12.27 24.1675 ;
        RECT  12.54 23.39 12.605 23.525 ;
        RECT  12.54 23.39 12.605 23.525 ;
        RECT  12.54 23.39 12.605 23.525 ;
        RECT  12.54 23.39 12.605 23.525 ;
        RECT  12.04 23.2125 12.175 23.2775 ;
        RECT  12.04 23.2125 12.175 23.2775 ;
        RECT  12.265 23.3625 12.4 23.4275 ;
        RECT  12.265 23.3625 12.4 23.4275 ;
        RECT  12.54 23.39 12.605 23.525 ;
        RECT  12.54 23.39 12.605 23.525 ;
        RECT  12.54 23.39 12.605 23.525 ;
        RECT  12.54 23.39 12.605 23.525 ;
        RECT  12.09 23.8825 12.155 24.0175 ;
        RECT  11.835 23.39 11.9 23.525 ;
        RECT  11.835 23.39 11.9 23.525 ;
        RECT  11.835 23.39 11.9 23.525 ;
        RECT  11.835 23.39 11.9 23.525 ;
        RECT  11.835 23.39 11.9 23.525 ;
        RECT  11.835 23.39 11.9 23.525 ;
        RECT  12.54 23.39 12.605 23.525 ;
        RECT  12.54 23.39 12.605 23.525 ;
        RECT  12.54 23.39 12.605 23.525 ;
        RECT  12.54 23.39 12.605 23.525 ;
        RECT  12.285 23.8825 12.35 24.0175 ;
        RECT  12.1525 24.2425 12.2875 24.3075 ;
        RECT  12.1525 24.2425 12.2875 24.3075 ;
        RECT  12.505 24.2425 12.64 24.3075 ;
        RECT  12.1475 22.8975 12.2825 22.9625 ;
        RECT  12.505 24.2425 12.64 24.3075 ;
        RECT  12.505 24.2425 12.64 24.3075 ;
        RECT  12.54 23.39 12.605 23.525 ;
        RECT  12.54 23.39 12.605 23.525 ;
        RECT  12.54 23.39 12.605 23.525 ;
        RECT  12.54 23.39 12.605 23.525 ;
        RECT  12.54 23.39 12.605 23.525 ;
        RECT  12.54 23.39 12.605 23.525 ;
        RECT  11.8 24.2425 11.935 24.3075 ;
        RECT  12.16 22.9 12.26 22.9625 ;
        RECT  12.16 22.8975 12.26 22.96 ;
        RECT  12.4875 24.1025 12.54 24.165 ;
        RECT  12.16 22.9 12.26 22.9625 ;
        RECT  12.5375 22.9625 12.6075 23.1625 ;
        RECT  12.5375 23.4925 12.6075 23.6275 ;
        RECT  12.5375 23.4925 12.6075 23.6275 ;
        RECT  11.7775 24.2425 12.6625 24.3075 ;
        RECT  12.3525 23.7275 12.5275 23.7925 ;
        RECT  11.8325 23.4925 11.9025 23.6275 ;
        RECT  12.0225 23.0525 12.0875 23.7925 ;
        RECT  12.16 22.8975 12.26 22.96 ;
        RECT  11.7825 24.1025 11.835 24.165 ;
        RECT  12.5375 23.4925 12.6075 23.6275 ;
        RECT  11.7775 22.8975 12.6625 22.9625 ;
        RECT  12.3525 23.1625 12.4175 23.7925 ;
        RECT  12.5375 23.4925 12.6075 23.6275 ;
        RECT  12.5375 23.4925 12.6075 23.6275 ;
        RECT  11.9175 23.7275 11.9875 24.0175 ;
        RECT  11.8325 23.4925 11.9025 23.6275 ;
        RECT  11.7775 24.1025 12.6625 24.1675 ;
        RECT  12.5375 23.4925 12.6075 23.6275 ;
        RECT  12.5375 22.9625 12.6075 23.1625 ;
        RECT  11.8325 22.9625 11.9025 23.1625 ;
        RECT  12.4575 23.7275 12.5275 24.0175 ;
        RECT  11.9175 23.7275 12.0875 23.7925 ;
        RECT  12.5375 25.3875 12.6025 25.5225 ;
        RECT  12.3525 25.3875 12.4175 25.5225 ;
        RECT  11.8375 25.3875 11.9025 25.5225 ;
        RECT  12.0225 25.3875 12.0875 25.5225 ;
        RECT  12.3525 24.9225 12.4175 25.0575 ;
        RECT  12.5375 24.9225 12.6025 25.0575 ;
        RECT  12.0225 24.9225 12.0875 25.0575 ;
        RECT  11.8375 24.9225 11.9025 25.0575 ;
        RECT  12.4575 24.5325 12.5225 24.6675 ;
        RECT  12.2725 24.5325 12.3375 24.6675 ;
        RECT  12.1025 24.5325 12.1675 24.6675 ;
        RECT  11.9175 24.5325 11.9825 24.6675 ;
        RECT  12.54 25.025 12.605 25.16 ;
        RECT  12.54 25.025 12.605 25.16 ;
        RECT  12.54 25.025 12.605 25.16 ;
        RECT  12.54 25.025 12.605 25.16 ;
        RECT  12.54 25.025 12.605 25.16 ;
        RECT  12.54 25.025 12.605 25.16 ;
        RECT  12.1475 25.5875 12.2825 25.6525 ;
        RECT  11.8 24.2425 11.935 24.3075 ;
        RECT  12.505 24.2425 12.64 24.3075 ;
        RECT  12.135 24.3825 12.27 24.4475 ;
        RECT  12.54 25.025 12.605 25.16 ;
        RECT  12.54 25.025 12.605 25.16 ;
        RECT  12.54 25.025 12.605 25.16 ;
        RECT  12.54 25.025 12.605 25.16 ;
        RECT  12.04 25.2725 12.175 25.3375 ;
        RECT  12.04 25.2725 12.175 25.3375 ;
        RECT  12.265 25.1225 12.4 25.1875 ;
        RECT  12.265 25.1225 12.4 25.1875 ;
        RECT  12.54 25.025 12.605 25.16 ;
        RECT  12.54 25.025 12.605 25.16 ;
        RECT  12.54 25.025 12.605 25.16 ;
        RECT  12.54 25.025 12.605 25.16 ;
        RECT  12.09 24.5325 12.155 24.6675 ;
        RECT  11.835 25.025 11.9 25.16 ;
        RECT  11.835 25.025 11.9 25.16 ;
        RECT  11.835 25.025 11.9 25.16 ;
        RECT  11.835 25.025 11.9 25.16 ;
        RECT  11.835 25.025 11.9 25.16 ;
        RECT  11.835 25.025 11.9 25.16 ;
        RECT  12.54 25.025 12.605 25.16 ;
        RECT  12.54 25.025 12.605 25.16 ;
        RECT  12.54 25.025 12.605 25.16 ;
        RECT  12.54 25.025 12.605 25.16 ;
        RECT  12.285 24.5325 12.35 24.6675 ;
        RECT  12.1525 24.2425 12.2875 24.3075 ;
        RECT  12.1525 24.2425 12.2875 24.3075 ;
        RECT  12.505 24.2425 12.64 24.3075 ;
        RECT  12.1475 25.5875 12.2825 25.6525 ;
        RECT  12.505 24.2425 12.64 24.3075 ;
        RECT  12.505 24.2425 12.64 24.3075 ;
        RECT  12.54 25.025 12.605 25.16 ;
        RECT  12.54 25.025 12.605 25.16 ;
        RECT  12.54 25.025 12.605 25.16 ;
        RECT  12.54 25.025 12.605 25.16 ;
        RECT  12.54 25.025 12.605 25.16 ;
        RECT  12.54 25.025 12.605 25.16 ;
        RECT  11.8 24.2425 11.935 24.3075 ;
        RECT  12.16 25.5875 12.26 25.65 ;
        RECT  12.16 25.59 12.26 25.6525 ;
        RECT  12.4875 24.385 12.54 24.4475 ;
        RECT  12.16 25.5875 12.26 25.65 ;
        RECT  12.5375 25.3875 12.6075 25.5875 ;
        RECT  12.5375 24.9225 12.6075 25.0575 ;
        RECT  12.5375 24.9225 12.6075 25.0575 ;
        RECT  11.7775 24.2425 12.6625 24.3075 ;
        RECT  12.3525 24.7575 12.5275 24.8225 ;
        RECT  11.8325 24.9225 11.9025 25.0575 ;
        RECT  12.0225 24.7575 12.0875 25.4975 ;
        RECT  12.16 25.59 12.26 25.6525 ;
        RECT  11.7825 24.385 11.835 24.4475 ;
        RECT  12.5375 24.9225 12.6075 25.0575 ;
        RECT  11.7775 25.5875 12.6625 25.6525 ;
        RECT  12.3525 24.7575 12.4175 25.3875 ;
        RECT  12.5375 24.9225 12.6075 25.0575 ;
        RECT  12.5375 24.9225 12.6075 25.0575 ;
        RECT  11.9175 24.5325 11.9875 24.8225 ;
        RECT  11.8325 24.9225 11.9025 25.0575 ;
        RECT  11.7775 24.3825 12.6625 24.4475 ;
        RECT  12.5375 24.9225 12.6075 25.0575 ;
        RECT  12.5375 25.3875 12.6075 25.5875 ;
        RECT  11.8325 25.3875 11.9025 25.5875 ;
        RECT  12.4575 24.5325 12.5275 24.8225 ;
        RECT  11.9175 24.7575 12.0875 24.8225 ;
        RECT  12.5375 25.7175 12.6025 25.8525 ;
        RECT  12.3525 25.7175 12.4175 25.8525 ;
        RECT  11.8375 25.7175 11.9025 25.8525 ;
        RECT  12.0225 25.7175 12.0875 25.8525 ;
        RECT  12.3525 26.1825 12.4175 26.3175 ;
        RECT  12.5375 26.1825 12.6025 26.3175 ;
        RECT  12.0225 26.1825 12.0875 26.3175 ;
        RECT  11.8375 26.1825 11.9025 26.3175 ;
        RECT  12.4575 26.5725 12.5225 26.7075 ;
        RECT  12.2725 26.5725 12.3375 26.7075 ;
        RECT  12.1025 26.5725 12.1675 26.7075 ;
        RECT  11.9175 26.5725 11.9825 26.7075 ;
        RECT  12.54 26.08 12.605 26.215 ;
        RECT  12.54 26.08 12.605 26.215 ;
        RECT  12.54 26.08 12.605 26.215 ;
        RECT  12.54 26.08 12.605 26.215 ;
        RECT  12.54 26.08 12.605 26.215 ;
        RECT  12.54 26.08 12.605 26.215 ;
        RECT  12.1475 25.5875 12.2825 25.6525 ;
        RECT  11.8 26.9325 11.935 26.9975 ;
        RECT  12.505 26.9325 12.64 26.9975 ;
        RECT  12.135 26.7925 12.27 26.8575 ;
        RECT  12.54 26.08 12.605 26.215 ;
        RECT  12.54 26.08 12.605 26.215 ;
        RECT  12.54 26.08 12.605 26.215 ;
        RECT  12.54 26.08 12.605 26.215 ;
        RECT  12.04 25.9025 12.175 25.9675 ;
        RECT  12.04 25.9025 12.175 25.9675 ;
        RECT  12.265 26.0525 12.4 26.1175 ;
        RECT  12.265 26.0525 12.4 26.1175 ;
        RECT  12.54 26.08 12.605 26.215 ;
        RECT  12.54 26.08 12.605 26.215 ;
        RECT  12.54 26.08 12.605 26.215 ;
        RECT  12.54 26.08 12.605 26.215 ;
        RECT  12.09 26.5725 12.155 26.7075 ;
        RECT  11.835 26.08 11.9 26.215 ;
        RECT  11.835 26.08 11.9 26.215 ;
        RECT  11.835 26.08 11.9 26.215 ;
        RECT  11.835 26.08 11.9 26.215 ;
        RECT  11.835 26.08 11.9 26.215 ;
        RECT  11.835 26.08 11.9 26.215 ;
        RECT  12.54 26.08 12.605 26.215 ;
        RECT  12.54 26.08 12.605 26.215 ;
        RECT  12.54 26.08 12.605 26.215 ;
        RECT  12.54 26.08 12.605 26.215 ;
        RECT  12.285 26.5725 12.35 26.7075 ;
        RECT  12.1525 26.9325 12.2875 26.9975 ;
        RECT  12.1525 26.9325 12.2875 26.9975 ;
        RECT  12.505 26.9325 12.64 26.9975 ;
        RECT  12.1475 25.5875 12.2825 25.6525 ;
        RECT  12.505 26.9325 12.64 26.9975 ;
        RECT  12.505 26.9325 12.64 26.9975 ;
        RECT  12.54 26.08 12.605 26.215 ;
        RECT  12.54 26.08 12.605 26.215 ;
        RECT  12.54 26.08 12.605 26.215 ;
        RECT  12.54 26.08 12.605 26.215 ;
        RECT  12.54 26.08 12.605 26.215 ;
        RECT  12.54 26.08 12.605 26.215 ;
        RECT  11.8 26.9325 11.935 26.9975 ;
        RECT  12.16 25.59 12.26 25.6525 ;
        RECT  12.16 25.5875 12.26 25.65 ;
        RECT  12.4875 26.7925 12.54 26.855 ;
        RECT  12.16 25.59 12.26 25.6525 ;
        RECT  12.5375 25.6525 12.6075 25.8525 ;
        RECT  12.5375 26.1825 12.6075 26.3175 ;
        RECT  12.5375 26.1825 12.6075 26.3175 ;
        RECT  11.7775 26.9325 12.6625 26.9975 ;
        RECT  12.3525 26.4175 12.5275 26.4825 ;
        RECT  11.8325 26.1825 11.9025 26.3175 ;
        RECT  12.0225 25.7425 12.0875 26.4825 ;
        RECT  12.16 25.5875 12.26 25.65 ;
        RECT  11.7825 26.7925 11.835 26.855 ;
        RECT  12.5375 26.1825 12.6075 26.3175 ;
        RECT  11.7775 25.5875 12.6625 25.6525 ;
        RECT  12.3525 25.8525 12.4175 26.4825 ;
        RECT  12.5375 26.1825 12.6075 26.3175 ;
        RECT  12.5375 26.1825 12.6075 26.3175 ;
        RECT  11.9175 26.4175 11.9875 26.7075 ;
        RECT  11.8325 26.1825 11.9025 26.3175 ;
        RECT  11.7775 26.7925 12.6625 26.8575 ;
        RECT  12.5375 26.1825 12.6075 26.3175 ;
        RECT  12.5375 25.6525 12.6075 25.8525 ;
        RECT  11.8325 25.6525 11.9025 25.8525 ;
        RECT  12.4575 26.4175 12.5275 26.7075 ;
        RECT  11.9175 26.4175 12.0875 26.4825 ;
        RECT  12.5375 28.0775 12.6025 28.2125 ;
        RECT  12.3525 28.0775 12.4175 28.2125 ;
        RECT  11.8375 28.0775 11.9025 28.2125 ;
        RECT  12.0225 28.0775 12.0875 28.2125 ;
        RECT  12.3525 27.6125 12.4175 27.7475 ;
        RECT  12.5375 27.6125 12.6025 27.7475 ;
        RECT  12.0225 27.6125 12.0875 27.7475 ;
        RECT  11.8375 27.6125 11.9025 27.7475 ;
        RECT  12.4575 27.2225 12.5225 27.3575 ;
        RECT  12.2725 27.2225 12.3375 27.3575 ;
        RECT  12.1025 27.2225 12.1675 27.3575 ;
        RECT  11.9175 27.2225 11.9825 27.3575 ;
        RECT  12.54 27.715 12.605 27.85 ;
        RECT  12.54 27.715 12.605 27.85 ;
        RECT  12.54 27.715 12.605 27.85 ;
        RECT  12.54 27.715 12.605 27.85 ;
        RECT  12.54 27.715 12.605 27.85 ;
        RECT  12.54 27.715 12.605 27.85 ;
        RECT  12.1475 28.2775 12.2825 28.3425 ;
        RECT  11.8 26.9325 11.935 26.9975 ;
        RECT  12.505 26.9325 12.64 26.9975 ;
        RECT  12.135 27.0725 12.27 27.1375 ;
        RECT  12.54 27.715 12.605 27.85 ;
        RECT  12.54 27.715 12.605 27.85 ;
        RECT  12.54 27.715 12.605 27.85 ;
        RECT  12.54 27.715 12.605 27.85 ;
        RECT  12.04 27.9625 12.175 28.0275 ;
        RECT  12.04 27.9625 12.175 28.0275 ;
        RECT  12.265 27.8125 12.4 27.8775 ;
        RECT  12.265 27.8125 12.4 27.8775 ;
        RECT  12.54 27.715 12.605 27.85 ;
        RECT  12.54 27.715 12.605 27.85 ;
        RECT  12.54 27.715 12.605 27.85 ;
        RECT  12.54 27.715 12.605 27.85 ;
        RECT  12.09 27.2225 12.155 27.3575 ;
        RECT  11.835 27.715 11.9 27.85 ;
        RECT  11.835 27.715 11.9 27.85 ;
        RECT  11.835 27.715 11.9 27.85 ;
        RECT  11.835 27.715 11.9 27.85 ;
        RECT  11.835 27.715 11.9 27.85 ;
        RECT  11.835 27.715 11.9 27.85 ;
        RECT  12.54 27.715 12.605 27.85 ;
        RECT  12.54 27.715 12.605 27.85 ;
        RECT  12.54 27.715 12.605 27.85 ;
        RECT  12.54 27.715 12.605 27.85 ;
        RECT  12.285 27.2225 12.35 27.3575 ;
        RECT  12.1525 26.9325 12.2875 26.9975 ;
        RECT  12.1525 26.9325 12.2875 26.9975 ;
        RECT  12.505 26.9325 12.64 26.9975 ;
        RECT  12.1475 28.2775 12.2825 28.3425 ;
        RECT  12.505 26.9325 12.64 26.9975 ;
        RECT  12.505 26.9325 12.64 26.9975 ;
        RECT  12.54 27.715 12.605 27.85 ;
        RECT  12.54 27.715 12.605 27.85 ;
        RECT  12.54 27.715 12.605 27.85 ;
        RECT  12.54 27.715 12.605 27.85 ;
        RECT  12.54 27.715 12.605 27.85 ;
        RECT  12.54 27.715 12.605 27.85 ;
        RECT  11.8 26.9325 11.935 26.9975 ;
        RECT  12.16 28.2775 12.26 28.34 ;
        RECT  12.16 28.28 12.26 28.3425 ;
        RECT  12.4875 27.075 12.54 27.1375 ;
        RECT  12.16 28.2775 12.26 28.34 ;
        RECT  12.5375 28.0775 12.6075 28.2775 ;
        RECT  12.5375 27.6125 12.6075 27.7475 ;
        RECT  12.5375 27.6125 12.6075 27.7475 ;
        RECT  11.7775 26.9325 12.6625 26.9975 ;
        RECT  12.3525 27.4475 12.5275 27.5125 ;
        RECT  11.8325 27.6125 11.9025 27.7475 ;
        RECT  12.0225 27.4475 12.0875 28.1875 ;
        RECT  12.16 28.28 12.26 28.3425 ;
        RECT  11.7825 27.075 11.835 27.1375 ;
        RECT  12.5375 27.6125 12.6075 27.7475 ;
        RECT  11.7775 28.2775 12.6625 28.3425 ;
        RECT  12.3525 27.4475 12.4175 28.0775 ;
        RECT  12.5375 27.6125 12.6075 27.7475 ;
        RECT  12.5375 27.6125 12.6075 27.7475 ;
        RECT  11.9175 27.2225 11.9875 27.5125 ;
        RECT  11.8325 27.6125 11.9025 27.7475 ;
        RECT  11.7775 27.0725 12.6625 27.1375 ;
        RECT  12.5375 27.6125 12.6075 27.7475 ;
        RECT  12.5375 28.0775 12.6075 28.2775 ;
        RECT  11.8325 28.0775 11.9025 28.2775 ;
        RECT  12.4575 27.2225 12.5275 27.5125 ;
        RECT  11.9175 27.4475 12.0875 27.5125 ;
        RECT  12.5375 28.4075 12.6025 28.5425 ;
        RECT  12.3525 28.4075 12.4175 28.5425 ;
        RECT  11.8375 28.4075 11.9025 28.5425 ;
        RECT  12.0225 28.4075 12.0875 28.5425 ;
        RECT  12.3525 28.8725 12.4175 29.0075 ;
        RECT  12.5375 28.8725 12.6025 29.0075 ;
        RECT  12.0225 28.8725 12.0875 29.0075 ;
        RECT  11.8375 28.8725 11.9025 29.0075 ;
        RECT  12.4575 29.2625 12.5225 29.3975 ;
        RECT  12.2725 29.2625 12.3375 29.3975 ;
        RECT  12.1025 29.2625 12.1675 29.3975 ;
        RECT  11.9175 29.2625 11.9825 29.3975 ;
        RECT  12.54 28.77 12.605 28.905 ;
        RECT  12.54 28.77 12.605 28.905 ;
        RECT  12.54 28.77 12.605 28.905 ;
        RECT  12.54 28.77 12.605 28.905 ;
        RECT  12.54 28.77 12.605 28.905 ;
        RECT  12.54 28.77 12.605 28.905 ;
        RECT  12.1475 28.2775 12.2825 28.3425 ;
        RECT  11.8 29.6225 11.935 29.6875 ;
        RECT  12.505 29.6225 12.64 29.6875 ;
        RECT  12.135 29.4825 12.27 29.5475 ;
        RECT  12.54 28.77 12.605 28.905 ;
        RECT  12.54 28.77 12.605 28.905 ;
        RECT  12.54 28.77 12.605 28.905 ;
        RECT  12.54 28.77 12.605 28.905 ;
        RECT  12.04 28.5925 12.175 28.6575 ;
        RECT  12.04 28.5925 12.175 28.6575 ;
        RECT  12.265 28.7425 12.4 28.8075 ;
        RECT  12.265 28.7425 12.4 28.8075 ;
        RECT  12.54 28.77 12.605 28.905 ;
        RECT  12.54 28.77 12.605 28.905 ;
        RECT  12.54 28.77 12.605 28.905 ;
        RECT  12.54 28.77 12.605 28.905 ;
        RECT  12.09 29.2625 12.155 29.3975 ;
        RECT  11.835 28.77 11.9 28.905 ;
        RECT  11.835 28.77 11.9 28.905 ;
        RECT  11.835 28.77 11.9 28.905 ;
        RECT  11.835 28.77 11.9 28.905 ;
        RECT  11.835 28.77 11.9 28.905 ;
        RECT  11.835 28.77 11.9 28.905 ;
        RECT  12.54 28.77 12.605 28.905 ;
        RECT  12.54 28.77 12.605 28.905 ;
        RECT  12.54 28.77 12.605 28.905 ;
        RECT  12.54 28.77 12.605 28.905 ;
        RECT  12.285 29.2625 12.35 29.3975 ;
        RECT  12.1525 29.6225 12.2875 29.6875 ;
        RECT  12.1525 29.6225 12.2875 29.6875 ;
        RECT  12.505 29.6225 12.64 29.6875 ;
        RECT  12.1475 28.2775 12.2825 28.3425 ;
        RECT  12.505 29.6225 12.64 29.6875 ;
        RECT  12.505 29.6225 12.64 29.6875 ;
        RECT  12.54 28.77 12.605 28.905 ;
        RECT  12.54 28.77 12.605 28.905 ;
        RECT  12.54 28.77 12.605 28.905 ;
        RECT  12.54 28.77 12.605 28.905 ;
        RECT  12.54 28.77 12.605 28.905 ;
        RECT  12.54 28.77 12.605 28.905 ;
        RECT  11.8 29.6225 11.935 29.6875 ;
        RECT  12.16 28.28 12.26 28.3425 ;
        RECT  12.16 28.2775 12.26 28.34 ;
        RECT  12.4875 29.4825 12.54 29.545 ;
        RECT  12.16 28.28 12.26 28.3425 ;
        RECT  12.5375 28.3425 12.6075 28.5425 ;
        RECT  12.5375 28.8725 12.6075 29.0075 ;
        RECT  12.5375 28.8725 12.6075 29.0075 ;
        RECT  11.7775 29.6225 12.6625 29.6875 ;
        RECT  12.3525 29.1075 12.5275 29.1725 ;
        RECT  11.8325 28.8725 11.9025 29.0075 ;
        RECT  12.0225 28.4325 12.0875 29.1725 ;
        RECT  12.16 28.2775 12.26 28.34 ;
        RECT  11.7825 29.4825 11.835 29.545 ;
        RECT  12.5375 28.8725 12.6075 29.0075 ;
        RECT  11.7775 28.2775 12.6625 28.3425 ;
        RECT  12.3525 28.5425 12.4175 29.1725 ;
        RECT  12.5375 28.8725 12.6075 29.0075 ;
        RECT  12.5375 28.8725 12.6075 29.0075 ;
        RECT  11.9175 29.1075 11.9875 29.3975 ;
        RECT  11.8325 28.8725 11.9025 29.0075 ;
        RECT  11.7775 29.4825 12.6625 29.5475 ;
        RECT  12.5375 28.8725 12.6075 29.0075 ;
        RECT  12.5375 28.3425 12.6075 28.5425 ;
        RECT  11.8325 28.3425 11.9025 28.5425 ;
        RECT  12.4575 29.1075 12.5275 29.3975 ;
        RECT  11.9175 29.1075 12.0875 29.1725 ;
        RECT  12.5375 30.7675 12.6025 30.9025 ;
        RECT  12.3525 30.7675 12.4175 30.9025 ;
        RECT  11.8375 30.7675 11.9025 30.9025 ;
        RECT  12.0225 30.7675 12.0875 30.9025 ;
        RECT  12.3525 30.3025 12.4175 30.4375 ;
        RECT  12.5375 30.3025 12.6025 30.4375 ;
        RECT  12.0225 30.3025 12.0875 30.4375 ;
        RECT  11.8375 30.3025 11.9025 30.4375 ;
        RECT  12.4575 29.9125 12.5225 30.0475 ;
        RECT  12.2725 29.9125 12.3375 30.0475 ;
        RECT  12.1025 29.9125 12.1675 30.0475 ;
        RECT  11.9175 29.9125 11.9825 30.0475 ;
        RECT  12.54 30.405 12.605 30.54 ;
        RECT  12.54 30.405 12.605 30.54 ;
        RECT  12.54 30.405 12.605 30.54 ;
        RECT  12.54 30.405 12.605 30.54 ;
        RECT  12.54 30.405 12.605 30.54 ;
        RECT  12.54 30.405 12.605 30.54 ;
        RECT  12.1475 30.9675 12.2825 31.0325 ;
        RECT  11.8 29.6225 11.935 29.6875 ;
        RECT  12.505 29.6225 12.64 29.6875 ;
        RECT  12.135 29.7625 12.27 29.8275 ;
        RECT  12.54 30.405 12.605 30.54 ;
        RECT  12.54 30.405 12.605 30.54 ;
        RECT  12.54 30.405 12.605 30.54 ;
        RECT  12.54 30.405 12.605 30.54 ;
        RECT  12.04 30.6525 12.175 30.7175 ;
        RECT  12.04 30.6525 12.175 30.7175 ;
        RECT  12.265 30.5025 12.4 30.5675 ;
        RECT  12.265 30.5025 12.4 30.5675 ;
        RECT  12.54 30.405 12.605 30.54 ;
        RECT  12.54 30.405 12.605 30.54 ;
        RECT  12.54 30.405 12.605 30.54 ;
        RECT  12.54 30.405 12.605 30.54 ;
        RECT  12.09 29.9125 12.155 30.0475 ;
        RECT  11.835 30.405 11.9 30.54 ;
        RECT  11.835 30.405 11.9 30.54 ;
        RECT  11.835 30.405 11.9 30.54 ;
        RECT  11.835 30.405 11.9 30.54 ;
        RECT  11.835 30.405 11.9 30.54 ;
        RECT  11.835 30.405 11.9 30.54 ;
        RECT  12.54 30.405 12.605 30.54 ;
        RECT  12.54 30.405 12.605 30.54 ;
        RECT  12.54 30.405 12.605 30.54 ;
        RECT  12.54 30.405 12.605 30.54 ;
        RECT  12.285 29.9125 12.35 30.0475 ;
        RECT  12.1525 29.6225 12.2875 29.6875 ;
        RECT  12.1525 29.6225 12.2875 29.6875 ;
        RECT  12.505 29.6225 12.64 29.6875 ;
        RECT  12.1475 30.9675 12.2825 31.0325 ;
        RECT  12.505 29.6225 12.64 29.6875 ;
        RECT  12.505 29.6225 12.64 29.6875 ;
        RECT  12.54 30.405 12.605 30.54 ;
        RECT  12.54 30.405 12.605 30.54 ;
        RECT  12.54 30.405 12.605 30.54 ;
        RECT  12.54 30.405 12.605 30.54 ;
        RECT  12.54 30.405 12.605 30.54 ;
        RECT  12.54 30.405 12.605 30.54 ;
        RECT  11.8 29.6225 11.935 29.6875 ;
        RECT  12.16 30.9675 12.26 31.03 ;
        RECT  12.16 30.97 12.26 31.0325 ;
        RECT  12.4875 29.765 12.54 29.8275 ;
        RECT  12.16 30.9675 12.26 31.03 ;
        RECT  12.5375 30.7675 12.6075 30.9675 ;
        RECT  12.5375 30.3025 12.6075 30.4375 ;
        RECT  12.5375 30.3025 12.6075 30.4375 ;
        RECT  11.7775 29.6225 12.6625 29.6875 ;
        RECT  12.3525 30.1375 12.5275 30.2025 ;
        RECT  11.8325 30.3025 11.9025 30.4375 ;
        RECT  12.0225 30.1375 12.0875 30.8775 ;
        RECT  12.16 30.97 12.26 31.0325 ;
        RECT  11.7825 29.765 11.835 29.8275 ;
        RECT  12.5375 30.3025 12.6075 30.4375 ;
        RECT  11.7775 30.9675 12.6625 31.0325 ;
        RECT  12.3525 30.1375 12.4175 30.7675 ;
        RECT  12.5375 30.3025 12.6075 30.4375 ;
        RECT  12.5375 30.3025 12.6075 30.4375 ;
        RECT  11.9175 29.9125 11.9875 30.2025 ;
        RECT  11.8325 30.3025 11.9025 30.4375 ;
        RECT  11.7775 29.7625 12.6625 29.8275 ;
        RECT  12.5375 30.3025 12.6075 30.4375 ;
        RECT  12.5375 30.7675 12.6075 30.9675 ;
        RECT  11.8325 30.7675 11.9025 30.9675 ;
        RECT  12.4575 29.9125 12.5275 30.2025 ;
        RECT  11.9175 30.1375 12.0875 30.2025 ;
        RECT  12.5375 31.0975 12.6025 31.2325 ;
        RECT  12.3525 31.0975 12.4175 31.2325 ;
        RECT  11.8375 31.0975 11.9025 31.2325 ;
        RECT  12.0225 31.0975 12.0875 31.2325 ;
        RECT  12.3525 31.5625 12.4175 31.6975 ;
        RECT  12.5375 31.5625 12.6025 31.6975 ;
        RECT  12.0225 31.5625 12.0875 31.6975 ;
        RECT  11.8375 31.5625 11.9025 31.6975 ;
        RECT  12.4575 31.9525 12.5225 32.0875 ;
        RECT  12.2725 31.9525 12.3375 32.0875 ;
        RECT  12.1025 31.9525 12.1675 32.0875 ;
        RECT  11.9175 31.9525 11.9825 32.0875 ;
        RECT  12.54 31.46 12.605 31.595 ;
        RECT  12.54 31.46 12.605 31.595 ;
        RECT  12.54 31.46 12.605 31.595 ;
        RECT  12.54 31.46 12.605 31.595 ;
        RECT  12.54 31.46 12.605 31.595 ;
        RECT  12.54 31.46 12.605 31.595 ;
        RECT  12.1475 30.9675 12.2825 31.0325 ;
        RECT  11.8 32.3125 11.935 32.3775 ;
        RECT  12.505 32.3125 12.64 32.3775 ;
        RECT  12.135 32.1725 12.27 32.2375 ;
        RECT  12.54 31.46 12.605 31.595 ;
        RECT  12.54 31.46 12.605 31.595 ;
        RECT  12.54 31.46 12.605 31.595 ;
        RECT  12.54 31.46 12.605 31.595 ;
        RECT  12.04 31.2825 12.175 31.3475 ;
        RECT  12.04 31.2825 12.175 31.3475 ;
        RECT  12.265 31.4325 12.4 31.4975 ;
        RECT  12.265 31.4325 12.4 31.4975 ;
        RECT  12.54 31.46 12.605 31.595 ;
        RECT  12.54 31.46 12.605 31.595 ;
        RECT  12.54 31.46 12.605 31.595 ;
        RECT  12.54 31.46 12.605 31.595 ;
        RECT  12.09 31.9525 12.155 32.0875 ;
        RECT  11.835 31.46 11.9 31.595 ;
        RECT  11.835 31.46 11.9 31.595 ;
        RECT  11.835 31.46 11.9 31.595 ;
        RECT  11.835 31.46 11.9 31.595 ;
        RECT  11.835 31.46 11.9 31.595 ;
        RECT  11.835 31.46 11.9 31.595 ;
        RECT  12.54 31.46 12.605 31.595 ;
        RECT  12.54 31.46 12.605 31.595 ;
        RECT  12.54 31.46 12.605 31.595 ;
        RECT  12.54 31.46 12.605 31.595 ;
        RECT  12.285 31.9525 12.35 32.0875 ;
        RECT  12.1525 32.3125 12.2875 32.3775 ;
        RECT  12.1525 32.3125 12.2875 32.3775 ;
        RECT  12.505 32.3125 12.64 32.3775 ;
        RECT  12.1475 30.9675 12.2825 31.0325 ;
        RECT  12.505 32.3125 12.64 32.3775 ;
        RECT  12.505 32.3125 12.64 32.3775 ;
        RECT  12.54 31.46 12.605 31.595 ;
        RECT  12.54 31.46 12.605 31.595 ;
        RECT  12.54 31.46 12.605 31.595 ;
        RECT  12.54 31.46 12.605 31.595 ;
        RECT  12.54 31.46 12.605 31.595 ;
        RECT  12.54 31.46 12.605 31.595 ;
        RECT  11.8 32.3125 11.935 32.3775 ;
        RECT  12.16 30.97 12.26 31.0325 ;
        RECT  12.16 30.9675 12.26 31.03 ;
        RECT  12.4875 32.1725 12.54 32.235 ;
        RECT  12.16 30.97 12.26 31.0325 ;
        RECT  12.5375 31.0325 12.6075 31.2325 ;
        RECT  12.5375 31.5625 12.6075 31.6975 ;
        RECT  12.5375 31.5625 12.6075 31.6975 ;
        RECT  11.7775 32.3125 12.6625 32.3775 ;
        RECT  12.3525 31.7975 12.5275 31.8625 ;
        RECT  11.8325 31.5625 11.9025 31.6975 ;
        RECT  12.0225 31.1225 12.0875 31.8625 ;
        RECT  12.16 30.9675 12.26 31.03 ;
        RECT  11.7825 32.1725 11.835 32.235 ;
        RECT  12.5375 31.5625 12.6075 31.6975 ;
        RECT  11.7775 30.9675 12.6625 31.0325 ;
        RECT  12.3525 31.2325 12.4175 31.8625 ;
        RECT  12.5375 31.5625 12.6075 31.6975 ;
        RECT  12.5375 31.5625 12.6075 31.6975 ;
        RECT  11.9175 31.7975 11.9875 32.0875 ;
        RECT  11.8325 31.5625 11.9025 31.6975 ;
        RECT  11.7775 32.1725 12.6625 32.2375 ;
        RECT  12.5375 31.5625 12.6075 31.6975 ;
        RECT  12.5375 31.0325 12.6075 31.2325 ;
        RECT  11.8325 31.0325 11.9025 31.2325 ;
        RECT  12.4575 31.7975 12.5275 32.0875 ;
        RECT  11.9175 31.7975 12.0875 31.8625 ;
        RECT  12.5375 33.4575 12.6025 33.5925 ;
        RECT  12.3525 33.4575 12.4175 33.5925 ;
        RECT  11.8375 33.4575 11.9025 33.5925 ;
        RECT  12.0225 33.4575 12.0875 33.5925 ;
        RECT  12.3525 32.9925 12.4175 33.1275 ;
        RECT  12.5375 32.9925 12.6025 33.1275 ;
        RECT  12.0225 32.9925 12.0875 33.1275 ;
        RECT  11.8375 32.9925 11.9025 33.1275 ;
        RECT  12.4575 32.6025 12.5225 32.7375 ;
        RECT  12.2725 32.6025 12.3375 32.7375 ;
        RECT  12.1025 32.6025 12.1675 32.7375 ;
        RECT  11.9175 32.6025 11.9825 32.7375 ;
        RECT  12.54 33.095 12.605 33.23 ;
        RECT  12.54 33.095 12.605 33.23 ;
        RECT  12.54 33.095 12.605 33.23 ;
        RECT  12.54 33.095 12.605 33.23 ;
        RECT  12.54 33.095 12.605 33.23 ;
        RECT  12.54 33.095 12.605 33.23 ;
        RECT  12.1475 33.6575 12.2825 33.7225 ;
        RECT  11.8 32.3125 11.935 32.3775 ;
        RECT  12.505 32.3125 12.64 32.3775 ;
        RECT  12.135 32.4525 12.27 32.5175 ;
        RECT  12.54 33.095 12.605 33.23 ;
        RECT  12.54 33.095 12.605 33.23 ;
        RECT  12.54 33.095 12.605 33.23 ;
        RECT  12.54 33.095 12.605 33.23 ;
        RECT  12.04 33.3425 12.175 33.4075 ;
        RECT  12.04 33.3425 12.175 33.4075 ;
        RECT  12.265 33.1925 12.4 33.2575 ;
        RECT  12.265 33.1925 12.4 33.2575 ;
        RECT  12.54 33.095 12.605 33.23 ;
        RECT  12.54 33.095 12.605 33.23 ;
        RECT  12.54 33.095 12.605 33.23 ;
        RECT  12.54 33.095 12.605 33.23 ;
        RECT  12.09 32.6025 12.155 32.7375 ;
        RECT  11.835 33.095 11.9 33.23 ;
        RECT  11.835 33.095 11.9 33.23 ;
        RECT  11.835 33.095 11.9 33.23 ;
        RECT  11.835 33.095 11.9 33.23 ;
        RECT  11.835 33.095 11.9 33.23 ;
        RECT  11.835 33.095 11.9 33.23 ;
        RECT  12.54 33.095 12.605 33.23 ;
        RECT  12.54 33.095 12.605 33.23 ;
        RECT  12.54 33.095 12.605 33.23 ;
        RECT  12.54 33.095 12.605 33.23 ;
        RECT  12.285 32.6025 12.35 32.7375 ;
        RECT  12.1525 32.3125 12.2875 32.3775 ;
        RECT  12.1525 32.3125 12.2875 32.3775 ;
        RECT  12.505 32.3125 12.64 32.3775 ;
        RECT  12.1475 33.6575 12.2825 33.7225 ;
        RECT  12.505 32.3125 12.64 32.3775 ;
        RECT  12.505 32.3125 12.64 32.3775 ;
        RECT  12.54 33.095 12.605 33.23 ;
        RECT  12.54 33.095 12.605 33.23 ;
        RECT  12.54 33.095 12.605 33.23 ;
        RECT  12.54 33.095 12.605 33.23 ;
        RECT  12.54 33.095 12.605 33.23 ;
        RECT  12.54 33.095 12.605 33.23 ;
        RECT  11.8 32.3125 11.935 32.3775 ;
        RECT  12.16 33.6575 12.26 33.72 ;
        RECT  12.16 33.66 12.26 33.7225 ;
        RECT  12.4875 32.455 12.54 32.5175 ;
        RECT  12.16 33.6575 12.26 33.72 ;
        RECT  12.5375 33.4575 12.6075 33.6575 ;
        RECT  12.5375 32.9925 12.6075 33.1275 ;
        RECT  12.5375 32.9925 12.6075 33.1275 ;
        RECT  11.7775 32.3125 12.6625 32.3775 ;
        RECT  12.3525 32.8275 12.5275 32.8925 ;
        RECT  11.8325 32.9925 11.9025 33.1275 ;
        RECT  12.0225 32.8275 12.0875 33.5675 ;
        RECT  12.16 33.66 12.26 33.7225 ;
        RECT  11.7825 32.455 11.835 32.5175 ;
        RECT  12.5375 32.9925 12.6075 33.1275 ;
        RECT  11.7775 33.6575 12.6625 33.7225 ;
        RECT  12.3525 32.8275 12.4175 33.4575 ;
        RECT  12.5375 32.9925 12.6075 33.1275 ;
        RECT  12.5375 32.9925 12.6075 33.1275 ;
        RECT  11.9175 32.6025 11.9875 32.8925 ;
        RECT  11.8325 32.9925 11.9025 33.1275 ;
        RECT  11.7775 32.4525 12.6625 32.5175 ;
        RECT  12.5375 32.9925 12.6075 33.1275 ;
        RECT  12.5375 33.4575 12.6075 33.6575 ;
        RECT  11.8325 33.4575 11.9025 33.6575 ;
        RECT  12.4575 32.6025 12.5275 32.8925 ;
        RECT  11.9175 32.8275 12.0875 32.8925 ;
        RECT  12.5375 33.7875 12.6025 33.9225 ;
        RECT  12.3525 33.7875 12.4175 33.9225 ;
        RECT  11.8375 33.7875 11.9025 33.9225 ;
        RECT  12.0225 33.7875 12.0875 33.9225 ;
        RECT  12.3525 34.2525 12.4175 34.3875 ;
        RECT  12.5375 34.2525 12.6025 34.3875 ;
        RECT  12.0225 34.2525 12.0875 34.3875 ;
        RECT  11.8375 34.2525 11.9025 34.3875 ;
        RECT  12.4575 34.6425 12.5225 34.7775 ;
        RECT  12.2725 34.6425 12.3375 34.7775 ;
        RECT  12.1025 34.6425 12.1675 34.7775 ;
        RECT  11.9175 34.6425 11.9825 34.7775 ;
        RECT  12.54 34.15 12.605 34.285 ;
        RECT  12.54 34.15 12.605 34.285 ;
        RECT  12.54 34.15 12.605 34.285 ;
        RECT  12.54 34.15 12.605 34.285 ;
        RECT  12.54 34.15 12.605 34.285 ;
        RECT  12.54 34.15 12.605 34.285 ;
        RECT  12.1475 33.6575 12.2825 33.7225 ;
        RECT  11.8 35.0025 11.935 35.0675 ;
        RECT  12.505 35.0025 12.64 35.0675 ;
        RECT  12.135 34.8625 12.27 34.9275 ;
        RECT  12.54 34.15 12.605 34.285 ;
        RECT  12.54 34.15 12.605 34.285 ;
        RECT  12.54 34.15 12.605 34.285 ;
        RECT  12.54 34.15 12.605 34.285 ;
        RECT  12.04 33.9725 12.175 34.0375 ;
        RECT  12.04 33.9725 12.175 34.0375 ;
        RECT  12.265 34.1225 12.4 34.1875 ;
        RECT  12.265 34.1225 12.4 34.1875 ;
        RECT  12.54 34.15 12.605 34.285 ;
        RECT  12.54 34.15 12.605 34.285 ;
        RECT  12.54 34.15 12.605 34.285 ;
        RECT  12.54 34.15 12.605 34.285 ;
        RECT  12.09 34.6425 12.155 34.7775 ;
        RECT  11.835 34.15 11.9 34.285 ;
        RECT  11.835 34.15 11.9 34.285 ;
        RECT  11.835 34.15 11.9 34.285 ;
        RECT  11.835 34.15 11.9 34.285 ;
        RECT  11.835 34.15 11.9 34.285 ;
        RECT  11.835 34.15 11.9 34.285 ;
        RECT  12.54 34.15 12.605 34.285 ;
        RECT  12.54 34.15 12.605 34.285 ;
        RECT  12.54 34.15 12.605 34.285 ;
        RECT  12.54 34.15 12.605 34.285 ;
        RECT  12.285 34.6425 12.35 34.7775 ;
        RECT  12.1525 35.0025 12.2875 35.0675 ;
        RECT  12.1525 35.0025 12.2875 35.0675 ;
        RECT  12.505 35.0025 12.64 35.0675 ;
        RECT  12.1475 33.6575 12.2825 33.7225 ;
        RECT  12.505 35.0025 12.64 35.0675 ;
        RECT  12.505 35.0025 12.64 35.0675 ;
        RECT  12.54 34.15 12.605 34.285 ;
        RECT  12.54 34.15 12.605 34.285 ;
        RECT  12.54 34.15 12.605 34.285 ;
        RECT  12.54 34.15 12.605 34.285 ;
        RECT  12.54 34.15 12.605 34.285 ;
        RECT  12.54 34.15 12.605 34.285 ;
        RECT  11.8 35.0025 11.935 35.0675 ;
        RECT  12.16 33.66 12.26 33.7225 ;
        RECT  12.16 33.6575 12.26 33.72 ;
        RECT  12.4875 34.8625 12.54 34.925 ;
        RECT  12.16 33.66 12.26 33.7225 ;
        RECT  12.5375 33.7225 12.6075 33.9225 ;
        RECT  12.5375 34.2525 12.6075 34.3875 ;
        RECT  12.5375 34.2525 12.6075 34.3875 ;
        RECT  11.7775 35.0025 12.6625 35.0675 ;
        RECT  12.3525 34.4875 12.5275 34.5525 ;
        RECT  11.8325 34.2525 11.9025 34.3875 ;
        RECT  12.0225 33.8125 12.0875 34.5525 ;
        RECT  12.16 33.6575 12.26 33.72 ;
        RECT  11.7825 34.8625 11.835 34.925 ;
        RECT  12.5375 34.2525 12.6075 34.3875 ;
        RECT  11.7775 33.6575 12.6625 33.7225 ;
        RECT  12.3525 33.9225 12.4175 34.5525 ;
        RECT  12.5375 34.2525 12.6075 34.3875 ;
        RECT  12.5375 34.2525 12.6075 34.3875 ;
        RECT  11.9175 34.4875 11.9875 34.7775 ;
        RECT  11.8325 34.2525 11.9025 34.3875 ;
        RECT  11.7775 34.8625 12.6625 34.9275 ;
        RECT  12.5375 34.2525 12.6075 34.3875 ;
        RECT  12.5375 33.7225 12.6075 33.9225 ;
        RECT  11.8325 33.7225 11.9025 33.9225 ;
        RECT  12.4575 34.4875 12.5275 34.7775 ;
        RECT  11.9175 34.4875 12.0875 34.5525 ;
        RECT  12.5375 36.1475 12.6025 36.2825 ;
        RECT  12.3525 36.1475 12.4175 36.2825 ;
        RECT  11.8375 36.1475 11.9025 36.2825 ;
        RECT  12.0225 36.1475 12.0875 36.2825 ;
        RECT  12.3525 35.6825 12.4175 35.8175 ;
        RECT  12.5375 35.6825 12.6025 35.8175 ;
        RECT  12.0225 35.6825 12.0875 35.8175 ;
        RECT  11.8375 35.6825 11.9025 35.8175 ;
        RECT  12.4575 35.2925 12.5225 35.4275 ;
        RECT  12.2725 35.2925 12.3375 35.4275 ;
        RECT  12.1025 35.2925 12.1675 35.4275 ;
        RECT  11.9175 35.2925 11.9825 35.4275 ;
        RECT  12.54 35.785 12.605 35.92 ;
        RECT  12.54 35.785 12.605 35.92 ;
        RECT  12.54 35.785 12.605 35.92 ;
        RECT  12.54 35.785 12.605 35.92 ;
        RECT  12.54 35.785 12.605 35.92 ;
        RECT  12.54 35.785 12.605 35.92 ;
        RECT  12.1475 36.3475 12.2825 36.4125 ;
        RECT  11.8 35.0025 11.935 35.0675 ;
        RECT  12.505 35.0025 12.64 35.0675 ;
        RECT  12.135 35.1425 12.27 35.2075 ;
        RECT  12.54 35.785 12.605 35.92 ;
        RECT  12.54 35.785 12.605 35.92 ;
        RECT  12.54 35.785 12.605 35.92 ;
        RECT  12.54 35.785 12.605 35.92 ;
        RECT  12.04 36.0325 12.175 36.0975 ;
        RECT  12.04 36.0325 12.175 36.0975 ;
        RECT  12.265 35.8825 12.4 35.9475 ;
        RECT  12.265 35.8825 12.4 35.9475 ;
        RECT  12.54 35.785 12.605 35.92 ;
        RECT  12.54 35.785 12.605 35.92 ;
        RECT  12.54 35.785 12.605 35.92 ;
        RECT  12.54 35.785 12.605 35.92 ;
        RECT  12.09 35.2925 12.155 35.4275 ;
        RECT  11.835 35.785 11.9 35.92 ;
        RECT  11.835 35.785 11.9 35.92 ;
        RECT  11.835 35.785 11.9 35.92 ;
        RECT  11.835 35.785 11.9 35.92 ;
        RECT  11.835 35.785 11.9 35.92 ;
        RECT  11.835 35.785 11.9 35.92 ;
        RECT  12.54 35.785 12.605 35.92 ;
        RECT  12.54 35.785 12.605 35.92 ;
        RECT  12.54 35.785 12.605 35.92 ;
        RECT  12.54 35.785 12.605 35.92 ;
        RECT  12.285 35.2925 12.35 35.4275 ;
        RECT  12.1525 35.0025 12.2875 35.0675 ;
        RECT  12.1525 35.0025 12.2875 35.0675 ;
        RECT  12.505 35.0025 12.64 35.0675 ;
        RECT  12.1475 36.3475 12.2825 36.4125 ;
        RECT  12.505 35.0025 12.64 35.0675 ;
        RECT  12.505 35.0025 12.64 35.0675 ;
        RECT  12.54 35.785 12.605 35.92 ;
        RECT  12.54 35.785 12.605 35.92 ;
        RECT  12.54 35.785 12.605 35.92 ;
        RECT  12.54 35.785 12.605 35.92 ;
        RECT  12.54 35.785 12.605 35.92 ;
        RECT  12.54 35.785 12.605 35.92 ;
        RECT  11.8 35.0025 11.935 35.0675 ;
        RECT  12.16 36.3475 12.26 36.41 ;
        RECT  12.16 36.35 12.26 36.4125 ;
        RECT  12.4875 35.145 12.54 35.2075 ;
        RECT  12.16 36.3475 12.26 36.41 ;
        RECT  12.5375 36.1475 12.6075 36.3475 ;
        RECT  12.5375 35.6825 12.6075 35.8175 ;
        RECT  12.5375 35.6825 12.6075 35.8175 ;
        RECT  11.7775 35.0025 12.6625 35.0675 ;
        RECT  12.3525 35.5175 12.5275 35.5825 ;
        RECT  11.8325 35.6825 11.9025 35.8175 ;
        RECT  12.0225 35.5175 12.0875 36.2575 ;
        RECT  12.16 36.35 12.26 36.4125 ;
        RECT  11.7825 35.145 11.835 35.2075 ;
        RECT  12.5375 35.6825 12.6075 35.8175 ;
        RECT  11.7775 36.3475 12.6625 36.4125 ;
        RECT  12.3525 35.5175 12.4175 36.1475 ;
        RECT  12.5375 35.6825 12.6075 35.8175 ;
        RECT  12.5375 35.6825 12.6075 35.8175 ;
        RECT  11.9175 35.2925 11.9875 35.5825 ;
        RECT  11.8325 35.6825 11.9025 35.8175 ;
        RECT  11.7775 35.1425 12.6625 35.2075 ;
        RECT  12.5375 35.6825 12.6075 35.8175 ;
        RECT  12.5375 36.1475 12.6075 36.3475 ;
        RECT  11.8325 36.1475 11.9025 36.3475 ;
        RECT  12.4575 35.2925 12.5275 35.5825 ;
        RECT  11.9175 35.5175 12.0875 35.5825 ;
        RECT  12.5375 36.4775 12.6025 36.6125 ;
        RECT  12.3525 36.4775 12.4175 36.6125 ;
        RECT  11.8375 36.4775 11.9025 36.6125 ;
        RECT  12.0225 36.4775 12.0875 36.6125 ;
        RECT  12.3525 36.9425 12.4175 37.0775 ;
        RECT  12.5375 36.9425 12.6025 37.0775 ;
        RECT  12.0225 36.9425 12.0875 37.0775 ;
        RECT  11.8375 36.9425 11.9025 37.0775 ;
        RECT  12.4575 37.3325 12.5225 37.4675 ;
        RECT  12.2725 37.3325 12.3375 37.4675 ;
        RECT  12.1025 37.3325 12.1675 37.4675 ;
        RECT  11.9175 37.3325 11.9825 37.4675 ;
        RECT  12.54 36.84 12.605 36.975 ;
        RECT  12.54 36.84 12.605 36.975 ;
        RECT  12.54 36.84 12.605 36.975 ;
        RECT  12.54 36.84 12.605 36.975 ;
        RECT  12.54 36.84 12.605 36.975 ;
        RECT  12.54 36.84 12.605 36.975 ;
        RECT  12.1475 36.3475 12.2825 36.4125 ;
        RECT  11.8 37.6925 11.935 37.7575 ;
        RECT  12.505 37.6925 12.64 37.7575 ;
        RECT  12.135 37.5525 12.27 37.6175 ;
        RECT  12.54 36.84 12.605 36.975 ;
        RECT  12.54 36.84 12.605 36.975 ;
        RECT  12.54 36.84 12.605 36.975 ;
        RECT  12.54 36.84 12.605 36.975 ;
        RECT  12.04 36.6625 12.175 36.7275 ;
        RECT  12.04 36.6625 12.175 36.7275 ;
        RECT  12.265 36.8125 12.4 36.8775 ;
        RECT  12.265 36.8125 12.4 36.8775 ;
        RECT  12.54 36.84 12.605 36.975 ;
        RECT  12.54 36.84 12.605 36.975 ;
        RECT  12.54 36.84 12.605 36.975 ;
        RECT  12.54 36.84 12.605 36.975 ;
        RECT  12.09 37.3325 12.155 37.4675 ;
        RECT  11.835 36.84 11.9 36.975 ;
        RECT  11.835 36.84 11.9 36.975 ;
        RECT  11.835 36.84 11.9 36.975 ;
        RECT  11.835 36.84 11.9 36.975 ;
        RECT  11.835 36.84 11.9 36.975 ;
        RECT  11.835 36.84 11.9 36.975 ;
        RECT  12.54 36.84 12.605 36.975 ;
        RECT  12.54 36.84 12.605 36.975 ;
        RECT  12.54 36.84 12.605 36.975 ;
        RECT  12.54 36.84 12.605 36.975 ;
        RECT  12.285 37.3325 12.35 37.4675 ;
        RECT  12.1525 37.6925 12.2875 37.7575 ;
        RECT  12.1525 37.6925 12.2875 37.7575 ;
        RECT  12.505 37.6925 12.64 37.7575 ;
        RECT  12.1475 36.3475 12.2825 36.4125 ;
        RECT  12.505 37.6925 12.64 37.7575 ;
        RECT  12.505 37.6925 12.64 37.7575 ;
        RECT  12.54 36.84 12.605 36.975 ;
        RECT  12.54 36.84 12.605 36.975 ;
        RECT  12.54 36.84 12.605 36.975 ;
        RECT  12.54 36.84 12.605 36.975 ;
        RECT  12.54 36.84 12.605 36.975 ;
        RECT  12.54 36.84 12.605 36.975 ;
        RECT  11.8 37.6925 11.935 37.7575 ;
        RECT  12.16 36.35 12.26 36.4125 ;
        RECT  12.16 36.3475 12.26 36.41 ;
        RECT  12.4875 37.5525 12.54 37.615 ;
        RECT  12.16 36.35 12.26 36.4125 ;
        RECT  12.5375 36.4125 12.6075 36.6125 ;
        RECT  12.5375 36.9425 12.6075 37.0775 ;
        RECT  12.5375 36.9425 12.6075 37.0775 ;
        RECT  11.7775 37.6925 12.6625 37.7575 ;
        RECT  12.3525 37.1775 12.5275 37.2425 ;
        RECT  11.8325 36.9425 11.9025 37.0775 ;
        RECT  12.0225 36.5025 12.0875 37.2425 ;
        RECT  12.16 36.3475 12.26 36.41 ;
        RECT  11.7825 37.5525 11.835 37.615 ;
        RECT  12.5375 36.9425 12.6075 37.0775 ;
        RECT  11.7775 36.3475 12.6625 36.4125 ;
        RECT  12.3525 36.6125 12.4175 37.2425 ;
        RECT  12.5375 36.9425 12.6075 37.0775 ;
        RECT  12.5375 36.9425 12.6075 37.0775 ;
        RECT  11.9175 37.1775 11.9875 37.4675 ;
        RECT  11.8325 36.9425 11.9025 37.0775 ;
        RECT  11.7775 37.5525 12.6625 37.6175 ;
        RECT  12.5375 36.9425 12.6075 37.0775 ;
        RECT  12.5375 36.4125 12.6075 36.6125 ;
        RECT  11.8325 36.4125 11.9025 36.6125 ;
        RECT  12.4575 37.1775 12.5275 37.4675 ;
        RECT  11.9175 37.1775 12.0875 37.2425 ;
        RECT  12.5375 38.8375 12.6025 38.9725 ;
        RECT  12.3525 38.8375 12.4175 38.9725 ;
        RECT  11.8375 38.8375 11.9025 38.9725 ;
        RECT  12.0225 38.8375 12.0875 38.9725 ;
        RECT  12.3525 38.3725 12.4175 38.5075 ;
        RECT  12.5375 38.3725 12.6025 38.5075 ;
        RECT  12.0225 38.3725 12.0875 38.5075 ;
        RECT  11.8375 38.3725 11.9025 38.5075 ;
        RECT  12.4575 37.9825 12.5225 38.1175 ;
        RECT  12.2725 37.9825 12.3375 38.1175 ;
        RECT  12.1025 37.9825 12.1675 38.1175 ;
        RECT  11.9175 37.9825 11.9825 38.1175 ;
        RECT  12.54 38.475 12.605 38.61 ;
        RECT  12.54 38.475 12.605 38.61 ;
        RECT  12.54 38.475 12.605 38.61 ;
        RECT  12.54 38.475 12.605 38.61 ;
        RECT  12.54 38.475 12.605 38.61 ;
        RECT  12.54 38.475 12.605 38.61 ;
        RECT  12.1475 39.0375 12.2825 39.1025 ;
        RECT  11.8 37.6925 11.935 37.7575 ;
        RECT  12.505 37.6925 12.64 37.7575 ;
        RECT  12.135 37.8325 12.27 37.8975 ;
        RECT  12.54 38.475 12.605 38.61 ;
        RECT  12.54 38.475 12.605 38.61 ;
        RECT  12.54 38.475 12.605 38.61 ;
        RECT  12.54 38.475 12.605 38.61 ;
        RECT  12.04 38.7225 12.175 38.7875 ;
        RECT  12.04 38.7225 12.175 38.7875 ;
        RECT  12.265 38.5725 12.4 38.6375 ;
        RECT  12.265 38.5725 12.4 38.6375 ;
        RECT  12.54 38.475 12.605 38.61 ;
        RECT  12.54 38.475 12.605 38.61 ;
        RECT  12.54 38.475 12.605 38.61 ;
        RECT  12.54 38.475 12.605 38.61 ;
        RECT  12.09 37.9825 12.155 38.1175 ;
        RECT  11.835 38.475 11.9 38.61 ;
        RECT  11.835 38.475 11.9 38.61 ;
        RECT  11.835 38.475 11.9 38.61 ;
        RECT  11.835 38.475 11.9 38.61 ;
        RECT  11.835 38.475 11.9 38.61 ;
        RECT  11.835 38.475 11.9 38.61 ;
        RECT  12.54 38.475 12.605 38.61 ;
        RECT  12.54 38.475 12.605 38.61 ;
        RECT  12.54 38.475 12.605 38.61 ;
        RECT  12.54 38.475 12.605 38.61 ;
        RECT  12.285 37.9825 12.35 38.1175 ;
        RECT  12.1525 37.6925 12.2875 37.7575 ;
        RECT  12.1525 37.6925 12.2875 37.7575 ;
        RECT  12.505 37.6925 12.64 37.7575 ;
        RECT  12.1475 39.0375 12.2825 39.1025 ;
        RECT  12.505 37.6925 12.64 37.7575 ;
        RECT  12.505 37.6925 12.64 37.7575 ;
        RECT  12.54 38.475 12.605 38.61 ;
        RECT  12.54 38.475 12.605 38.61 ;
        RECT  12.54 38.475 12.605 38.61 ;
        RECT  12.54 38.475 12.605 38.61 ;
        RECT  12.54 38.475 12.605 38.61 ;
        RECT  12.54 38.475 12.605 38.61 ;
        RECT  11.8 37.6925 11.935 37.7575 ;
        RECT  12.16 39.0375 12.26 39.1 ;
        RECT  12.16 39.04 12.26 39.1025 ;
        RECT  12.4875 37.835 12.54 37.8975 ;
        RECT  12.16 39.0375 12.26 39.1 ;
        RECT  12.5375 38.8375 12.6075 39.0375 ;
        RECT  12.5375 38.3725 12.6075 38.5075 ;
        RECT  12.5375 38.3725 12.6075 38.5075 ;
        RECT  11.7775 37.6925 12.6625 37.7575 ;
        RECT  12.3525 38.2075 12.5275 38.2725 ;
        RECT  11.8325 38.3725 11.9025 38.5075 ;
        RECT  12.0225 38.2075 12.0875 38.9475 ;
        RECT  12.16 39.04 12.26 39.1025 ;
        RECT  11.7825 37.835 11.835 37.8975 ;
        RECT  12.5375 38.3725 12.6075 38.5075 ;
        RECT  11.7775 39.0375 12.6625 39.1025 ;
        RECT  12.3525 38.2075 12.4175 38.8375 ;
        RECT  12.5375 38.3725 12.6075 38.5075 ;
        RECT  12.5375 38.3725 12.6075 38.5075 ;
        RECT  11.9175 37.9825 11.9875 38.2725 ;
        RECT  11.8325 38.3725 11.9025 38.5075 ;
        RECT  11.7775 37.8325 12.6625 37.8975 ;
        RECT  12.5375 38.3725 12.6075 38.5075 ;
        RECT  12.5375 38.8375 12.6075 39.0375 ;
        RECT  11.8325 38.8375 11.9025 39.0375 ;
        RECT  12.4575 37.9825 12.5275 38.2725 ;
        RECT  11.9175 38.2075 12.0875 38.2725 ;
        RECT  12.5375 39.1675 12.6025 39.3025 ;
        RECT  12.3525 39.1675 12.4175 39.3025 ;
        RECT  11.8375 39.1675 11.9025 39.3025 ;
        RECT  12.0225 39.1675 12.0875 39.3025 ;
        RECT  12.3525 39.6325 12.4175 39.7675 ;
        RECT  12.5375 39.6325 12.6025 39.7675 ;
        RECT  12.0225 39.6325 12.0875 39.7675 ;
        RECT  11.8375 39.6325 11.9025 39.7675 ;
        RECT  12.4575 40.0225 12.5225 40.1575 ;
        RECT  12.2725 40.0225 12.3375 40.1575 ;
        RECT  12.1025 40.0225 12.1675 40.1575 ;
        RECT  11.9175 40.0225 11.9825 40.1575 ;
        RECT  12.54 39.53 12.605 39.665 ;
        RECT  12.54 39.53 12.605 39.665 ;
        RECT  12.54 39.53 12.605 39.665 ;
        RECT  12.54 39.53 12.605 39.665 ;
        RECT  12.54 39.53 12.605 39.665 ;
        RECT  12.54 39.53 12.605 39.665 ;
        RECT  12.1475 39.0375 12.2825 39.1025 ;
        RECT  11.8 40.3825 11.935 40.4475 ;
        RECT  12.505 40.3825 12.64 40.4475 ;
        RECT  12.135 40.2425 12.27 40.3075 ;
        RECT  12.54 39.53 12.605 39.665 ;
        RECT  12.54 39.53 12.605 39.665 ;
        RECT  12.54 39.53 12.605 39.665 ;
        RECT  12.54 39.53 12.605 39.665 ;
        RECT  12.04 39.3525 12.175 39.4175 ;
        RECT  12.04 39.3525 12.175 39.4175 ;
        RECT  12.265 39.5025 12.4 39.5675 ;
        RECT  12.265 39.5025 12.4 39.5675 ;
        RECT  12.54 39.53 12.605 39.665 ;
        RECT  12.54 39.53 12.605 39.665 ;
        RECT  12.54 39.53 12.605 39.665 ;
        RECT  12.54 39.53 12.605 39.665 ;
        RECT  12.09 40.0225 12.155 40.1575 ;
        RECT  11.835 39.53 11.9 39.665 ;
        RECT  11.835 39.53 11.9 39.665 ;
        RECT  11.835 39.53 11.9 39.665 ;
        RECT  11.835 39.53 11.9 39.665 ;
        RECT  11.835 39.53 11.9 39.665 ;
        RECT  11.835 39.53 11.9 39.665 ;
        RECT  12.54 39.53 12.605 39.665 ;
        RECT  12.54 39.53 12.605 39.665 ;
        RECT  12.54 39.53 12.605 39.665 ;
        RECT  12.54 39.53 12.605 39.665 ;
        RECT  12.285 40.0225 12.35 40.1575 ;
        RECT  12.1525 40.3825 12.2875 40.4475 ;
        RECT  12.1525 40.3825 12.2875 40.4475 ;
        RECT  12.505 40.3825 12.64 40.4475 ;
        RECT  12.1475 39.0375 12.2825 39.1025 ;
        RECT  12.505 40.3825 12.64 40.4475 ;
        RECT  12.505 40.3825 12.64 40.4475 ;
        RECT  12.54 39.53 12.605 39.665 ;
        RECT  12.54 39.53 12.605 39.665 ;
        RECT  12.54 39.53 12.605 39.665 ;
        RECT  12.54 39.53 12.605 39.665 ;
        RECT  12.54 39.53 12.605 39.665 ;
        RECT  12.54 39.53 12.605 39.665 ;
        RECT  11.8 40.3825 11.935 40.4475 ;
        RECT  12.16 39.04 12.26 39.1025 ;
        RECT  12.16 39.0375 12.26 39.1 ;
        RECT  12.4875 40.2425 12.54 40.305 ;
        RECT  12.16 39.04 12.26 39.1025 ;
        RECT  12.5375 39.1025 12.6075 39.3025 ;
        RECT  12.5375 39.6325 12.6075 39.7675 ;
        RECT  12.5375 39.6325 12.6075 39.7675 ;
        RECT  11.7775 40.3825 12.6625 40.4475 ;
        RECT  12.3525 39.8675 12.5275 39.9325 ;
        RECT  11.8325 39.6325 11.9025 39.7675 ;
        RECT  12.0225 39.1925 12.0875 39.9325 ;
        RECT  12.16 39.0375 12.26 39.1 ;
        RECT  11.7825 40.2425 11.835 40.305 ;
        RECT  12.5375 39.6325 12.6075 39.7675 ;
        RECT  11.7775 39.0375 12.6625 39.1025 ;
        RECT  12.3525 39.3025 12.4175 39.9325 ;
        RECT  12.5375 39.6325 12.6075 39.7675 ;
        RECT  12.5375 39.6325 12.6075 39.7675 ;
        RECT  11.9175 39.8675 11.9875 40.1575 ;
        RECT  11.8325 39.6325 11.9025 39.7675 ;
        RECT  11.7775 40.2425 12.6625 40.3075 ;
        RECT  12.5375 39.6325 12.6075 39.7675 ;
        RECT  12.5375 39.1025 12.6075 39.3025 ;
        RECT  11.8325 39.1025 11.9025 39.3025 ;
        RECT  12.4575 39.8675 12.5275 40.1575 ;
        RECT  11.9175 39.8675 12.0875 39.9325 ;
        RECT  11.1625 41.66 12.5725 41.725 ;
        RECT  11.1625 41.1 12.5725 41.165 ;
        RECT  11.1625 41.1 11.8675 41.165 ;
        RECT  11.1625 41.66 11.8675 41.725 ;
        RECT  11.5475 41.3125 11.6125 41.725 ;
        RECT  11.3575 40.8625 11.4225 40.9975 ;
        RECT  11.5475 40.8625 11.6125 40.9975 ;
        RECT  11.3575 41.3125 11.4225 41.4475 ;
        RECT  11.5475 41.3125 11.6125 41.4475 ;
        RECT  11.5475 41.3125 11.6125 41.4475 ;
        RECT  11.7375 41.3125 11.8025 41.4475 ;
        RECT  11.3925 41.1 11.5275 41.165 ;
        RECT  11.5475 41.5575 11.6125 41.6925 ;
        RECT  11.3575 41.3125 11.4225 41.4475 ;
        RECT  11.7375 41.3125 11.8025 41.4475 ;
        RECT  11.3575 40.8625 11.4225 40.9975 ;
        RECT  11.5475 40.8625 11.6125 40.9975 ;
        RECT  11.8675 41.1 12.5725 41.165 ;
        RECT  11.8675 41.66 12.5725 41.725 ;
        RECT  12.2525 41.3125 12.3175 41.725 ;
        RECT  12.0625 40.8625 12.1275 40.9975 ;
        RECT  12.2525 40.8625 12.3175 40.9975 ;
        RECT  12.0625 41.3125 12.1275 41.4475 ;
        RECT  12.2525 41.3125 12.3175 41.4475 ;
        RECT  12.2525 41.3125 12.3175 41.4475 ;
        RECT  12.4425 41.3125 12.5075 41.4475 ;
        RECT  12.0975 41.1 12.2325 41.165 ;
        RECT  12.2525 41.5575 12.3175 41.6925 ;
        RECT  12.0625 41.3125 12.1275 41.4475 ;
        RECT  12.4425 41.3125 12.5075 41.4475 ;
        RECT  12.0625 40.8625 12.1275 40.9975 ;
        RECT  12.2525 40.8625 12.3175 40.9975 ;
        RECT  11.1625 18.7 12.5725 18.765 ;
        RECT  11.1625 14.2575 12.5725 14.3225 ;
        RECT  11.1625 14.1275 12.5725 14.1925 ;
        RECT  11.67 14.9225 11.735 15.1975 ;
        RECT  11.485 14.9225 11.55 15.1975 ;
        RECT  11.48 14.9225 11.545 15.1975 ;
        RECT  11.295 14.9225 11.36 15.1975 ;
        RECT  11.58 14.465 11.645 14.74 ;
        RECT  11.395 14.465 11.46 14.74 ;
        RECT  11.48 15.6675 11.545 16.2225 ;
        RECT  11.295 15.6675 11.36 16.2225 ;
        RECT  11.67 15.6675 11.735 16.2225 ;
        RECT  11.485 15.6675 11.55 16.2225 ;
        RECT  11.48 17.45 11.545 18.145 ;
        RECT  11.295 17.45 11.36 18.145 ;
        RECT  11.67 16.48 11.735 17.175 ;
        RECT  11.485 16.48 11.55 17.175 ;
        RECT  11.4775 18.4975 11.5425 18.6325 ;
        RECT  11.4525 14.1275 11.5875 14.1925 ;
        RECT  11.835 14.2575 11.9 14.3925 ;
        RECT  11.13 14.2575 11.195 14.3925 ;
        RECT  11.6725 17.04 11.7375 17.175 ;
        RECT  11.755 14.4875 11.82 14.6225 ;
        RECT  11.29 17.45 11.355 17.585 ;
        RECT  11.4475 18.3625 11.5825 18.4275 ;
        RECT  11.4825 18.2925 11.5475 18.4275 ;
        RECT  11.4825 16.15 11.5475 16.285 ;
        RECT  11.425 15.4625 11.49 15.5975 ;
        RECT  11.54 15.2625 11.605 15.3975 ;
        RECT  11.4325 14.2575 11.4925 14.3225 ;
        RECT  11.3925 14.1275 11.4575 14.1925 ;
        RECT  11.82 14.3225 11.835 14.3925 ;
        RECT  11.225 18.4275 11.2925 18.765 ;
        RECT  11.225 18.3625 11.5825 18.4275 ;
        RECT  11.7275 17.32 11.7925 18.5675 ;
        RECT  11.225 18.7 11.2925 18.765 ;
        RECT  11.58 14.3225 11.645 14.475 ;
        RECT  11.755 14.2575 11.82 14.4875 ;
        RECT  11.475 18.4975 11.7925 18.5675 ;
        RECT  11.4825 17.32 11.5475 17.5175 ;
        RECT  11.295 17.32 11.7925 17.385 ;
        RECT  11.485 16.35 11.55 16.545 ;
        RECT  11.485 16.35 11.735 16.415 ;
        RECT  11.445 14.6525 11.515 14.98 ;
        RECT  11.1275 14.2575 11.9025 14.3225 ;
        RECT  11.67 16.22 11.735 16.415 ;
        RECT  11.295 16.2225 11.36 17.32 ;
        RECT  11.1275 18.7 11.9025 18.765 ;
        RECT  11.445 15.4975 11.735 15.5625 ;
        RECT  11.295 15.2975 11.585 15.3625 ;
        RECT  11.295 15.1925 11.36 16.06 ;
        RECT  11.67 15.1975 11.735 16.06 ;
        RECT  11.1275 14.1275 11.9025 14.1925 ;
        RECT  12.375 14.9225 12.44 15.1975 ;
        RECT  12.19 14.9225 12.255 15.1975 ;
        RECT  12.185 14.9225 12.25 15.1975 ;
        RECT  12.0 14.9225 12.065 15.1975 ;
        RECT  12.285 14.465 12.35 14.74 ;
        RECT  12.1 14.465 12.165 14.74 ;
        RECT  12.185 15.6675 12.25 16.2225 ;
        RECT  12.0 15.6675 12.065 16.2225 ;
        RECT  12.375 15.6675 12.44 16.2225 ;
        RECT  12.19 15.6675 12.255 16.2225 ;
        RECT  12.185 17.45 12.25 18.145 ;
        RECT  12.0 17.45 12.065 18.145 ;
        RECT  12.375 16.48 12.44 17.175 ;
        RECT  12.19 16.48 12.255 17.175 ;
        RECT  12.1825 18.4975 12.2475 18.6325 ;
        RECT  12.1575 14.1275 12.2925 14.1925 ;
        RECT  12.54 14.2575 12.605 14.3925 ;
        RECT  11.835 14.2575 11.9 14.3925 ;
        RECT  12.3775 17.04 12.4425 17.175 ;
        RECT  12.46 14.4875 12.525 14.6225 ;
        RECT  11.995 17.45 12.06 17.585 ;
        RECT  12.1525 18.3625 12.2875 18.4275 ;
        RECT  12.1875 18.2925 12.2525 18.4275 ;
        RECT  12.1875 16.15 12.2525 16.285 ;
        RECT  12.13 15.4625 12.195 15.5975 ;
        RECT  12.245 15.2625 12.31 15.3975 ;
        RECT  12.1375 14.2575 12.1975 14.3225 ;
        RECT  12.0975 14.1275 12.1625 14.1925 ;
        RECT  12.525 14.3225 12.54 14.3925 ;
        RECT  11.93 18.4275 11.9975 18.765 ;
        RECT  11.93 18.3625 12.2875 18.4275 ;
        RECT  12.4325 17.32 12.4975 18.5675 ;
        RECT  11.93 18.7 11.9975 18.765 ;
        RECT  12.285 14.3225 12.35 14.475 ;
        RECT  12.46 14.2575 12.525 14.4875 ;
        RECT  12.18 18.4975 12.4975 18.5675 ;
        RECT  12.1875 17.32 12.2525 17.5175 ;
        RECT  12.0 17.32 12.4975 17.385 ;
        RECT  12.19 16.35 12.255 16.545 ;
        RECT  12.19 16.35 12.44 16.415 ;
        RECT  12.15 14.6525 12.22 14.98 ;
        RECT  11.8325 14.2575 12.6075 14.3225 ;
        RECT  12.375 16.22 12.44 16.415 ;
        RECT  12.0 16.2225 12.065 17.32 ;
        RECT  11.8325 18.7 12.6075 18.765 ;
        RECT  12.15 15.4975 12.44 15.5625 ;
        RECT  12.0 15.2975 12.29 15.3625 ;
        RECT  12.0 15.1925 12.065 16.06 ;
        RECT  12.375 15.1975 12.44 16.06 ;
        RECT  11.8325 14.1275 12.6075 14.1925 ;
        RECT  11.1625 10.1025 12.5725 10.1675 ;
        RECT  11.1625 10.2325 12.5725 10.2975 ;
        RECT  11.1625 11.035 12.5725 11.1 ;
        RECT  11.5825 13.4975 11.6475 13.6325 ;
        RECT  11.2075 13.4975 11.2725 13.6325 ;
        RECT  11.2075 11.57 11.2725 11.705 ;
        RECT  11.5825 11.57 11.6475 11.705 ;
        RECT  11.5825 12.7025 11.6475 13.1175 ;
        RECT  11.2075 12.7025 11.2725 13.1175 ;
        RECT  11.2075 12.085 11.2725 12.5 ;
        RECT  11.5825 12.085 11.6475 12.5 ;
        RECT  11.3925 10.515 11.4575 10.93 ;
        RECT  11.2075 10.515 11.2725 10.93 ;
        RECT  11.5475 10.515 11.6125 10.93 ;
        RECT  11.7325 10.515 11.7975 10.93 ;
        RECT  11.3925 11.205 11.4575 11.34 ;
        RECT  11.2075 11.205 11.2725 11.34 ;
        RECT  11.5475 11.205 11.6125 11.34 ;
        RECT  11.7325 11.205 11.7975 11.34 ;
        RECT  11.37 9.97 11.505 10.035 ;
        RECT  11.445 11.925 11.51 12.06 ;
        RECT  11.835 11.57 11.9 11.705 ;
        RECT  11.7475 11.57 11.8125 11.705 ;
        RECT  11.13 12.5325 11.195 12.6675 ;
        RECT  11.835 11.0 11.9 11.135 ;
        RECT  11.13 11.0 11.195 11.135 ;
        RECT  11.55 11.205 11.615 11.34 ;
        RECT  11.835 13.4975 11.9 13.6325 ;
        RECT  11.75 13.4975 11.815 13.6325 ;
        RECT  11.55 10.795 11.615 10.93 ;
        RECT  11.41 10.795 11.475 10.93 ;
        RECT  11.4325 10.3825 11.5675 10.4475 ;
        RECT  11.265 9.9725 11.4 10.0375 ;
        RECT  11.605 10.1025 11.74 10.1675 ;
        RECT  11.835 11.205 11.9 11.34 ;
        RECT  11.13 11.205 11.195 11.34 ;
        RECT  11.2675 10.2325 11.4025 10.2975 ;
        RECT  11.41 13.175 11.475 13.31 ;
        RECT  11.58 11.57 11.645 11.705 ;
        RECT  11.27 12.485 11.335 12.62 ;
        RECT  11.41 11.205 11.475 11.34 ;
        RECT  11.3475 13.175 11.4125 13.31 ;
        RECT  11.13 11.57 11.195 11.705 ;
        RECT  11.58 12.085 11.645 12.22 ;
        RECT  11.315 13.7075 11.38 13.8425 ;
        RECT  11.13 13.4975 11.195 13.6325 ;
        RECT  11.815 13.4975 11.835 13.6325 ;
        RECT  11.8125 11.57 11.835 11.705 ;
        RECT  11.4825 11.0375 11.54 11.0975 ;
        RECT  11.4575 10.1025 11.53 10.1675 ;
        RECT  11.46 10.2325 11.53 10.2975 ;
        RECT  11.19 13.4975 11.2025 13.6325 ;
        RECT  11.195 12.5325 11.3375 12.6675 ;
        RECT  11.1275 11.035 11.9025 11.1 ;
        RECT  11.465 10.2975 11.53 10.4475 ;
        RECT  11.7925 11.205 11.835 11.34 ;
        RECT  11.7325 10.2975 11.7975 10.515 ;
        RECT  11.2075 10.2975 11.2725 10.515 ;
        RECT  11.1275 10.2325 11.9025 10.2975 ;
        RECT  11.1275 10.1025 11.9025 10.1675 ;
        RECT  11.19 11.205 11.2025 11.34 ;
        RECT  11.2575 12.485 11.2725 12.62 ;
        RECT  11.19 11.57 11.2025 11.705 ;
        RECT  11.2075 12.5 11.2725 12.7025 ;
        RECT  11.5825 13.6325 11.6475 13.7075 ;
        RECT  11.445 11.4125 11.6075 11.4775 ;
        RECT  11.1975 13.4975 11.2075 13.6325 ;
        RECT  11.1975 11.57 11.2075 11.705 ;
        RECT  11.5425 11.2875 11.6075 11.4125 ;
        RECT  11.445 11.4125 11.51 12.01 ;
        RECT  11.5825 13.1175 11.6475 13.4975 ;
        RECT  11.3125 13.7075 11.6475 13.7725 ;
        RECT  11.1975 11.205 11.2075 11.34 ;
        RECT  12.2875 13.4975 12.3525 13.6325 ;
        RECT  11.9125 13.4975 11.9775 13.6325 ;
        RECT  11.9125 11.57 11.9775 11.705 ;
        RECT  12.2875 11.57 12.3525 11.705 ;
        RECT  12.2875 12.7025 12.3525 13.1175 ;
        RECT  11.9125 12.7025 11.9775 13.1175 ;
        RECT  11.9125 12.085 11.9775 12.5 ;
        RECT  12.2875 12.085 12.3525 12.5 ;
        RECT  12.0975 10.515 12.1625 10.93 ;
        RECT  11.9125 10.515 11.9775 10.93 ;
        RECT  12.2525 10.515 12.3175 10.93 ;
        RECT  12.4375 10.515 12.5025 10.93 ;
        RECT  12.0975 11.205 12.1625 11.34 ;
        RECT  11.9125 11.205 11.9775 11.34 ;
        RECT  12.2525 11.205 12.3175 11.34 ;
        RECT  12.4375 11.205 12.5025 11.34 ;
        RECT  12.075 9.97 12.21 10.035 ;
        RECT  12.15 11.925 12.215 12.06 ;
        RECT  12.54 11.57 12.605 11.705 ;
        RECT  12.4525 11.57 12.5175 11.705 ;
        RECT  11.835 12.5325 11.9 12.6675 ;
        RECT  12.54 11.0 12.605 11.135 ;
        RECT  11.835 11.0 11.9 11.135 ;
        RECT  12.255 11.205 12.32 11.34 ;
        RECT  12.54 13.4975 12.605 13.6325 ;
        RECT  12.455 13.4975 12.52 13.6325 ;
        RECT  12.255 10.795 12.32 10.93 ;
        RECT  12.115 10.795 12.18 10.93 ;
        RECT  12.1375 10.3825 12.2725 10.4475 ;
        RECT  11.97 9.9725 12.105 10.0375 ;
        RECT  12.31 10.1025 12.445 10.1675 ;
        RECT  12.54 11.205 12.605 11.34 ;
        RECT  11.835 11.205 11.9 11.34 ;
        RECT  11.9725 10.2325 12.1075 10.2975 ;
        RECT  12.115 13.175 12.18 13.31 ;
        RECT  12.285 11.57 12.35 11.705 ;
        RECT  11.975 12.485 12.04 12.62 ;
        RECT  12.115 11.205 12.18 11.34 ;
        RECT  12.0525 13.175 12.1175 13.31 ;
        RECT  11.835 11.57 11.9 11.705 ;
        RECT  12.285 12.085 12.35 12.22 ;
        RECT  12.02 13.7075 12.085 13.8425 ;
        RECT  11.835 13.4975 11.9 13.6325 ;
        RECT  12.52 13.4975 12.54 13.6325 ;
        RECT  12.5175 11.57 12.54 11.705 ;
        RECT  12.1875 11.0375 12.245 11.0975 ;
        RECT  12.1625 10.1025 12.235 10.1675 ;
        RECT  12.165 10.2325 12.235 10.2975 ;
        RECT  11.895 13.4975 11.9075 13.6325 ;
        RECT  11.9 12.5325 12.0425 12.6675 ;
        RECT  11.8325 11.035 12.6075 11.1 ;
        RECT  12.17 10.2975 12.235 10.4475 ;
        RECT  12.4975 11.205 12.54 11.34 ;
        RECT  12.4375 10.2975 12.5025 10.515 ;
        RECT  11.9125 10.2975 11.9775 10.515 ;
        RECT  11.8325 10.2325 12.6075 10.2975 ;
        RECT  11.8325 10.1025 12.6075 10.1675 ;
        RECT  11.895 11.205 11.9075 11.34 ;
        RECT  11.9625 12.485 11.9775 12.62 ;
        RECT  11.895 11.57 11.9075 11.705 ;
        RECT  11.9125 12.5 11.9775 12.7025 ;
        RECT  12.2875 13.6325 12.3525 13.7075 ;
        RECT  12.15 11.4125 12.3125 11.4775 ;
        RECT  11.9025 13.4975 11.9125 13.6325 ;
        RECT  11.9025 11.57 11.9125 11.705 ;
        RECT  12.2475 11.2875 12.3125 11.4125 ;
        RECT  12.15 11.4125 12.215 12.01 ;
        RECT  12.2875 13.1175 12.3525 13.4975 ;
        RECT  12.0175 13.7075 12.3525 13.7725 ;
        RECT  11.9025 11.205 11.9125 11.34 ;
        RECT  11.1625 3.5675 12.5725 3.6325 ;
        RECT  11.1625 9.565 12.5725 9.63 ;
        RECT  11.7025 6.085 11.7675 6.22 ;
        RECT  11.5175 6.085 11.5825 6.22 ;
        RECT  11.7025 4.85 11.7675 4.985 ;
        RECT  11.5175 4.85 11.5825 4.985 ;
        RECT  11.5125 6.085 11.5775 6.22 ;
        RECT  11.3275 6.085 11.3925 6.22 ;
        RECT  11.5125 9.045 11.5775 9.18 ;
        RECT  11.3275 9.045 11.3925 9.18 ;
        RECT  11.5125 4.85 11.5775 4.985 ;
        RECT  11.3275 4.85 11.3925 4.985 ;
        RECT  11.7025 9.045 11.7675 9.18 ;
        RECT  11.5175 9.045 11.5825 9.18 ;
        RECT  11.5125 4.315 11.5775 4.45 ;
        RECT  11.3275 4.315 11.3925 4.45 ;
        RECT  11.6525 7.275 11.7175 7.41 ;
        RECT  11.4675 7.275 11.5325 7.41 ;
        RECT  11.7025 7.81 11.7675 7.945 ;
        RECT  11.5175 7.81 11.5825 7.945 ;
        RECT  11.5125 7.81 11.5775 7.945 ;
        RECT  11.3275 7.81 11.3925 7.945 ;
        RECT  11.7025 8.235 11.7675 8.37 ;
        RECT  11.5175 8.235 11.5825 8.37 ;
        RECT  11.7025 5.275 11.7675 5.41 ;
        RECT  11.5175 5.275 11.5825 5.41 ;
        RECT  11.7025 8.62 11.7675 8.755 ;
        RECT  11.5175 8.62 11.5825 8.755 ;
        RECT  11.5125 8.62 11.5775 8.755 ;
        RECT  11.3275 8.62 11.3925 8.755 ;
        RECT  11.5125 5.275 11.5775 5.41 ;
        RECT  11.3275 5.275 11.3925 5.41 ;
        RECT  11.5125 8.235 11.5775 8.37 ;
        RECT  11.3275 8.235 11.3925 8.37 ;
        RECT  11.5125 5.66 11.5775 5.795 ;
        RECT  11.3275 5.66 11.3925 5.795 ;
        RECT  11.7025 5.66 11.7675 5.795 ;
        RECT  11.5175 5.66 11.5825 5.795 ;
        RECT  11.5125 3.89 11.5775 4.025 ;
        RECT  11.3275 3.89 11.3925 4.025 ;
        RECT  11.5875 6.865 11.6525 7.0 ;
        RECT  11.4025 6.865 11.4675 7.0 ;
        RECT  11.39 3.6 11.525 3.665 ;
        RECT  11.3275 9.0975 11.3925 9.2325 ;
        RECT  11.2175 7.2825 11.2825 7.4175 ;
        RECT  11.3275 6.3825 11.3925 6.5175 ;
        RECT  11.75 6.8575 11.815 6.9925 ;
        RECT  11.3275 9.4625 11.3925 9.5975 ;
        RECT  11.835 3.92 11.9 4.055 ;
        RECT  11.6925 8.0025 11.7575 8.1375 ;
        RECT  11.695 6.395 11.76 6.53 ;
        RECT  11.695 4.9975 11.76 5.1325 ;
        RECT  11.13 3.78 11.195 3.915 ;
        RECT  11.705 3.8975 11.77 4.0325 ;
        RECT  11.705 5.5075 11.84 5.5725 ;
        RECT  11.745 4.4225 11.81 4.5575 ;
        RECT  11.705 8.4675 11.84 8.5325 ;
        RECT  11.6525 9.355 11.7175 9.49 ;
        RECT  11.5725 5.885 11.6375 6.02 ;
        RECT  11.5625 8.845 11.6275 8.98 ;
        RECT  11.33 7.155 11.465 7.22 ;
        RECT  11.835 6.8575 11.9 6.9925 ;
        RECT  11.22 4.15 11.355 4.215 ;
        RECT  11.33 5.6625 11.395 5.7975 ;
        RECT  11.695 9.355 11.76 9.49 ;
        RECT  11.5175 8.845 11.5825 8.98 ;
        RECT  11.835 8.4325 11.9 8.5675 ;
        RECT  11.835 3.73 11.9 3.865 ;
        RECT  11.695 6.395 11.76 6.53 ;
        RECT  11.835 5.4725 11.9 5.6075 ;
        RECT  11.33 5.2725 11.395 5.4075 ;
        RECT  11.5175 5.2725 11.5825 5.4075 ;
        RECT  11.5175 5.885 11.5825 6.02 ;
        RECT  11.3275 8.2325 11.3925 8.3675 ;
        RECT  11.5175 8.2325 11.5825 8.3675 ;
        RECT  11.1275 3.6 11.9025 3.665 ;
        RECT  11.1975 6.67 11.2625 9.565 ;
        RECT  11.7025 9.18 11.7675 9.49 ;
        RECT  11.3275 8.755 11.3925 9.045 ;
        RECT  11.3275 7.945 11.3925 8.235 ;
        RECT  11.4675 9.5675 11.54 9.63 ;
        RECT  11.5125 9.18 11.5825 9.565 ;
        RECT  11.5125 7.945 11.5825 8.235 ;
        RECT  11.5125 8.465 11.5825 8.6225 ;
        RECT  11.7025 8.755 11.7675 9.045 ;
        RECT  11.7025 7.945 11.7675 8.235 ;
        RECT  11.5125 8.465 11.8975 8.535 ;
        RECT  11.1275 9.565 11.9025 9.63 ;
        RECT  11.1275 7.575 11.9025 7.64 ;
        RECT  11.1975 4.68 11.2625 6.605 ;
        RECT  11.7025 6.22 11.7675 6.53 ;
        RECT  11.3275 5.795 11.3925 6.085 ;
        RECT  11.4025 6.96 11.4675 7.41 ;
        RECT  11.5125 6.22 11.5825 6.605 ;
        RECT  11.5125 5.505 11.5825 5.6625 ;
        RECT  11.3275 6.5175 11.3925 6.605 ;
        RECT  11.7025 5.795 11.7675 6.085 ;
        RECT  11.5875 6.735 11.8325 6.8 ;
        RECT  11.75 6.735 11.8325 6.8575 ;
        RECT  11.77 6.8575 11.8375 6.9925 ;
        RECT  11.1275 6.605 11.9025 6.67 ;
        RECT  11.3275 4.985 11.3925 5.275 ;
        RECT  11.5125 4.4475 11.5775 4.615 ;
        RECT  11.5775 3.955 11.835 4.025 ;
        RECT  11.3275 3.89 11.3925 4.315 ;
        RECT  11.5125 4.985 11.5825 5.275 ;
        RECT  11.22 4.145 11.3925 4.22 ;
        RECT  11.7025 4.985 11.7675 5.275 ;
        RECT  11.705 3.825 11.77 3.8975 ;
        RECT  11.5125 5.505 11.8975 5.575 ;
        RECT  11.745 4.535 11.81 4.65 ;
        RECT  11.1275 3.76 11.9025 3.825 ;
        RECT  11.1275 4.615 11.9025 4.68 ;
        RECT  11.2675 3.605 11.3325 3.6625 ;
        RECT  11.835 3.845 11.9 3.9675 ;
        RECT  11.6525 7.4075 11.7175 7.575 ;
        RECT  11.5875 6.8 11.655 6.9025 ;
        RECT  11.9675 6.085 12.0325 6.22 ;
        RECT  12.1525 6.085 12.2175 6.22 ;
        RECT  11.9675 4.85 12.0325 4.985 ;
        RECT  12.1525 4.85 12.2175 4.985 ;
        RECT  12.1575 6.085 12.2225 6.22 ;
        RECT  12.3425 6.085 12.4075 6.22 ;
        RECT  12.1575 9.045 12.2225 9.18 ;
        RECT  12.3425 9.045 12.4075 9.18 ;
        RECT  12.1575 4.85 12.2225 4.985 ;
        RECT  12.3425 4.85 12.4075 4.985 ;
        RECT  11.9675 9.045 12.0325 9.18 ;
        RECT  12.1525 9.045 12.2175 9.18 ;
        RECT  12.1575 4.315 12.2225 4.45 ;
        RECT  12.3425 4.315 12.4075 4.45 ;
        RECT  12.0175 7.275 12.0825 7.41 ;
        RECT  12.2025 7.275 12.2675 7.41 ;
        RECT  11.9675 7.81 12.0325 7.945 ;
        RECT  12.1525 7.81 12.2175 7.945 ;
        RECT  12.1575 7.81 12.2225 7.945 ;
        RECT  12.3425 7.81 12.4075 7.945 ;
        RECT  11.9675 8.235 12.0325 8.37 ;
        RECT  12.1525 8.235 12.2175 8.37 ;
        RECT  11.9675 5.275 12.0325 5.41 ;
        RECT  12.1525 5.275 12.2175 5.41 ;
        RECT  11.9675 8.62 12.0325 8.755 ;
        RECT  12.1525 8.62 12.2175 8.755 ;
        RECT  12.1575 8.62 12.2225 8.755 ;
        RECT  12.3425 8.62 12.4075 8.755 ;
        RECT  12.1575 5.275 12.2225 5.41 ;
        RECT  12.3425 5.275 12.4075 5.41 ;
        RECT  12.1575 8.235 12.2225 8.37 ;
        RECT  12.3425 8.235 12.4075 8.37 ;
        RECT  12.1575 5.66 12.2225 5.795 ;
        RECT  12.3425 5.66 12.4075 5.795 ;
        RECT  11.9675 5.66 12.0325 5.795 ;
        RECT  12.1525 5.66 12.2175 5.795 ;
        RECT  12.1575 3.89 12.2225 4.025 ;
        RECT  12.3425 3.89 12.4075 4.025 ;
        RECT  12.0825 6.865 12.1475 7.0 ;
        RECT  12.2675 6.865 12.3325 7.0 ;
        RECT  12.21 3.6 12.345 3.665 ;
        RECT  12.3425 9.0975 12.4075 9.2325 ;
        RECT  12.4525 7.2825 12.5175 7.4175 ;
        RECT  12.3425 6.3825 12.4075 6.5175 ;
        RECT  11.92 6.8575 11.985 6.9925 ;
        RECT  12.3425 9.4625 12.4075 9.5975 ;
        RECT  11.835 3.92 11.9 4.055 ;
        RECT  11.9775 8.0025 12.0425 8.1375 ;
        RECT  11.975 6.395 12.04 6.53 ;
        RECT  11.975 4.9975 12.04 5.1325 ;
        RECT  12.54 3.78 12.605 3.915 ;
        RECT  11.965 3.8975 12.03 4.0325 ;
        RECT  11.895 5.5075 12.03 5.5725 ;
        RECT  11.925 4.4225 11.99 4.5575 ;
        RECT  11.895 8.4675 12.03 8.5325 ;
        RECT  12.0175 9.355 12.0825 9.49 ;
        RECT  12.0975 5.885 12.1625 6.02 ;
        RECT  12.1075 8.845 12.1725 8.98 ;
        RECT  12.27 7.155 12.405 7.22 ;
        RECT  11.835 6.8575 11.9 6.9925 ;
        RECT  12.38 4.15 12.515 4.215 ;
        RECT  12.34 5.6625 12.405 5.7975 ;
        RECT  11.975 9.355 12.04 9.49 ;
        RECT  12.1525 8.845 12.2175 8.98 ;
        RECT  11.835 8.4325 11.9 8.5675 ;
        RECT  11.835 3.73 11.9 3.865 ;
        RECT  11.975 6.395 12.04 6.53 ;
        RECT  11.835 5.4725 11.9 5.6075 ;
        RECT  12.34 5.2725 12.405 5.4075 ;
        RECT  12.1525 5.2725 12.2175 5.4075 ;
        RECT  12.1525 5.885 12.2175 6.02 ;
        RECT  12.3425 8.2325 12.4075 8.3675 ;
        RECT  12.1525 8.2325 12.2175 8.3675 ;
        RECT  11.8325 3.6 12.6075 3.665 ;
        RECT  12.4725 6.67 12.5375 9.565 ;
        RECT  11.9675 9.18 12.0325 9.49 ;
        RECT  12.3425 8.755 12.4075 9.045 ;
        RECT  12.3425 7.945 12.4075 8.235 ;
        RECT  12.195 9.5675 12.2675 9.63 ;
        RECT  12.1525 9.18 12.2225 9.565 ;
        RECT  12.1525 7.945 12.2225 8.235 ;
        RECT  12.1525 8.465 12.2225 8.6225 ;
        RECT  11.9675 8.755 12.0325 9.045 ;
        RECT  11.9675 7.945 12.0325 8.235 ;
        RECT  11.8375 8.465 12.2225 8.535 ;
        RECT  11.8325 9.565 12.6075 9.63 ;
        RECT  11.8325 7.575 12.6075 7.64 ;
        RECT  12.4725 4.68 12.5375 6.605 ;
        RECT  11.9675 6.22 12.0325 6.53 ;
        RECT  12.3425 5.795 12.4075 6.085 ;
        RECT  12.2675 6.96 12.3325 7.41 ;
        RECT  12.1525 6.22 12.2225 6.605 ;
        RECT  12.1525 5.505 12.2225 5.6625 ;
        RECT  12.3425 6.5175 12.4075 6.605 ;
        RECT  11.9675 5.795 12.0325 6.085 ;
        RECT  11.9025 6.735 12.1475 6.8 ;
        RECT  11.9025 6.735 11.985 6.8575 ;
        RECT  11.8975 6.8575 11.965 6.9925 ;
        RECT  11.8325 6.605 12.6075 6.67 ;
        RECT  12.3425 4.985 12.4075 5.275 ;
        RECT  12.1575 4.4475 12.2225 4.615 ;
        RECT  11.9 3.955 12.1575 4.025 ;
        RECT  12.3425 3.89 12.4075 4.315 ;
        RECT  12.1525 4.985 12.2225 5.275 ;
        RECT  12.3425 4.145 12.515 4.22 ;
        RECT  11.9675 4.985 12.0325 5.275 ;
        RECT  11.965 3.825 12.03 3.8975 ;
        RECT  11.8375 5.505 12.2225 5.575 ;
        RECT  11.925 4.535 11.99 4.65 ;
        RECT  11.8325 3.76 12.6075 3.825 ;
        RECT  11.8325 4.615 12.6075 4.68 ;
        RECT  12.4025 3.605 12.4675 3.6625 ;
        RECT  11.835 3.845 11.9 3.9675 ;
        RECT  12.0175 7.4075 12.0825 7.575 ;
        RECT  12.08 6.8 12.1475 6.9025 ;
        RECT  11.1625 2.9625 12.5725 3.0275 ;
        RECT  11.1625 1.415 12.5725 1.48 ;
        RECT  11.1625 1.545 12.5725 1.61 ;
        RECT  11.5175 5.44 11.5825 5.575 ;
        RECT  11.3325 5.44 11.3975 5.575 ;
        RECT  11.5175 5.955 11.5825 6.09 ;
        RECT  11.3325 5.955 11.3975 6.09 ;
        RECT  11.645 4.045 11.71 4.18 ;
        RECT  11.27 4.045 11.335 4.18 ;
        RECT  11.645 4.6725 11.71 5.0875 ;
        RECT  11.27 4.6725 11.335 5.0875 ;
        RECT  11.66 4.3125 11.795 4.3775 ;
        RECT  11.6825 5.9625 11.7475 6.0975 ;
        RECT  11.4475 5.18 11.5825 5.245 ;
        RECT  11.6025 3.8925 11.7375 3.9575 ;
        RECT  11.835 3.8925 11.9 4.0275 ;
        RECT  11.22 5.31 11.355 5.375 ;
        RECT  11.325 3.7625 11.46 3.8275 ;
        RECT  11.58 5.82 11.715 5.885 ;
        RECT  11.835 5.9525 11.9 6.0875 ;
        RECT  11.58 5.78 11.715 5.845 ;
        RECT  11.6025 5.18 11.7375 5.245 ;
        RECT  11.3075 5.7625 11.3725 5.8975 ;
        RECT  11.515 5.485 11.58 5.62 ;
        RECT  11.4875 3.7625 11.545 3.8275 ;
        RECT  11.44 5.31 11.5025 5.375 ;
        RECT  11.3325 5.57 11.3975 6.09 ;
        RECT  11.27 4.1575 11.335 4.6725 ;
        RECT  11.58 4.3125 11.715 4.3775 ;
        RECT  11.1625 3.7625 11.9025 3.8275 ;
        RECT  11.1625 3.8925 11.9025 3.9575 ;
        RECT  11.645 3.9575 11.71 4.045 ;
        RECT  11.5375 5.9525 11.835 6.0875 ;
        RECT  11.1625 5.31 11.9025 5.375 ;
        RECT  11.1625 5.18 11.9025 5.245 ;
        RECT  11.645 5.0875 11.71 5.18 ;
        RECT  11.305 5.18 11.37 5.245 ;
        RECT  11.27 4.045 11.335 4.18 ;
        RECT  12.1525 5.44 12.2175 5.575 ;
        RECT  12.3375 5.44 12.4025 5.575 ;
        RECT  12.1525 5.955 12.2175 6.09 ;
        RECT  12.3375 5.955 12.4025 6.09 ;
        RECT  12.025 4.045 12.09 4.18 ;
        RECT  12.4 4.045 12.465 4.18 ;
        RECT  12.025 4.6725 12.09 5.0875 ;
        RECT  12.4 4.6725 12.465 5.0875 ;
        RECT  11.94 4.3125 12.075 4.3775 ;
        RECT  11.9875 5.9625 12.0525 6.0975 ;
        RECT  12.1525 5.18 12.2875 5.245 ;
        RECT  11.9975 3.8925 12.1325 3.9575 ;
        RECT  11.835 3.8925 11.9 4.0275 ;
        RECT  12.38 5.31 12.515 5.375 ;
        RECT  12.275 3.7625 12.41 3.8275 ;
        RECT  12.02 5.82 12.155 5.885 ;
        RECT  11.835 5.9525 11.9 6.0875 ;
        RECT  12.02 5.78 12.155 5.845 ;
        RECT  11.9975 5.18 12.1325 5.245 ;
        RECT  12.3625 5.7625 12.4275 5.8975 ;
        RECT  12.155 5.485 12.22 5.62 ;
        RECT  12.19 3.7625 12.2475 3.8275 ;
        RECT  12.2325 5.31 12.295 5.375 ;
        RECT  12.3375 5.57 12.4025 6.09 ;
        RECT  12.4 4.1575 12.465 4.6725 ;
        RECT  12.02 4.3125 12.155 4.3775 ;
        RECT  11.8325 3.7625 12.5725 3.8275 ;
        RECT  11.8325 3.8925 12.5725 3.9575 ;
        RECT  12.025 3.9575 12.09 4.045 ;
        RECT  11.9 5.9525 12.1975 6.0875 ;
        RECT  11.8325 5.31 12.5725 5.375 ;
        RECT  11.8325 5.18 12.5725 5.245 ;
        RECT  12.025 5.0875 12.09 5.18 ;
        RECT  12.365 5.18 12.43 5.245 ;
        RECT  12.4 4.045 12.465 4.18 ;
        RECT  5.0025 19.4925 5.0675 19.5575 ;
        RECT  5.0025 20.9225 5.0675 20.9875 ;
        RECT  5.0025 22.1825 5.0675 22.2475 ;
        RECT  5.0025 23.6125 5.0675 23.6775 ;
        RECT  5.0025 24.8725 5.0675 24.9375 ;
        RECT  5.0025 26.3025 5.0675 26.3675 ;
        RECT  5.0025 27.5625 5.0675 27.6275 ;
        RECT  5.0025 28.9925 5.0675 29.0575 ;
        RECT  5.0025 30.2525 5.0675 30.3175 ;
        RECT  5.0025 31.6825 5.0675 31.7475 ;
        RECT  5.0025 32.9425 5.0675 33.0075 ;
        RECT  5.0025 34.3725 5.0675 34.4375 ;
        RECT  5.0025 35.6325 5.0675 35.6975 ;
        RECT  5.0025 37.0625 5.0675 37.1275 ;
        RECT  5.0025 38.3225 5.0675 38.3875 ;
        RECT  5.0025 39.7525 5.0675 39.8175 ;
        RECT  2.8525 8.73 4.2525 8.795 ;
        RECT  3.0275 10.165 4.2525 10.23 ;
        RECT  3.2025 11.42 4.2525 11.485 ;
        RECT  3.3775 12.855 4.2525 12.92 ;
        RECT  3.5525 14.11 4.2525 14.175 ;
        RECT  3.7275 15.545 4.2525 15.61 ;
        RECT  3.9025 16.8 4.2525 16.865 ;
        RECT  4.0775 18.235 4.2525 18.3 ;
        RECT  2.8525 19.805 4.2525 19.87 ;
        RECT  3.5525 19.275 4.2525 19.34 ;
        RECT  2.8525 20.61 4.2525 20.675 ;
        RECT  3.7275 21.14 4.2525 21.205 ;
        RECT  2.8525 22.495 4.2525 22.56 ;
        RECT  3.9025 21.965 4.2525 22.03 ;
        RECT  2.8525 23.3 4.2525 23.365 ;
        RECT  4.0775 23.83 4.2525 23.895 ;
        RECT  3.0275 25.185 4.2525 25.25 ;
        RECT  3.5525 24.655 4.2525 24.72 ;
        RECT  3.0275 25.99 4.2525 26.055 ;
        RECT  3.7275 26.52 4.2525 26.585 ;
        RECT  3.0275 27.875 4.2525 27.94 ;
        RECT  3.9025 27.345 4.2525 27.41 ;
        RECT  3.0275 28.68 4.2525 28.745 ;
        RECT  4.0775 29.21 4.2525 29.275 ;
        RECT  3.2025 30.565 4.2525 30.63 ;
        RECT  3.5525 30.035 4.2525 30.1 ;
        RECT  3.2025 31.37 4.2525 31.435 ;
        RECT  3.7275 31.9 4.2525 31.965 ;
        RECT  3.2025 33.255 4.2525 33.32 ;
        RECT  3.9025 32.725 4.2525 32.79 ;
        RECT  3.2025 34.06 4.2525 34.125 ;
        RECT  4.0775 34.59 4.2525 34.655 ;
        RECT  3.3775 35.945 4.2525 36.01 ;
        RECT  3.5525 35.415 4.2525 35.48 ;
        RECT  3.3775 36.75 4.2525 36.815 ;
        RECT  3.7275 37.28 4.2525 37.345 ;
        RECT  3.3775 38.635 4.2525 38.7 ;
        RECT  3.9025 38.105 4.2525 38.17 ;
        RECT  3.3775 39.44 4.2525 39.505 ;
        RECT  4.0775 39.97 4.2525 40.035 ;
        RECT  4.7475 8.7325 4.8125 8.7975 ;
        RECT  4.7475 10.1625 4.8125 10.2275 ;
        RECT  4.7475 11.4225 4.8125 11.4875 ;
        RECT  4.7475 12.8525 4.8125 12.9175 ;
        RECT  6.6525 8.73 6.7175 9.3175 ;
        RECT  6.1925 9.2525 6.7175 9.3175 ;
        RECT  7.2075 8.73 7.6275 8.795 ;
        RECT  6.5425 9.4475 7.2775 9.5125 ;
        RECT  6.3675 8.1025 7.2775 8.1675 ;
        RECT  6.6525 9.6425 6.7175 10.23 ;
        RECT  6.0175 9.6425 6.7175 9.7075 ;
        RECT  7.2075 10.165 7.4525 10.23 ;
        RECT  6.5425 9.4475 7.2775 9.5125 ;
        RECT  6.3675 10.7925 7.2775 10.8575 ;
        RECT  5.5625 9.045 6.2625 9.11 ;
        RECT  5.5625 8.515 6.0875 8.58 ;
        RECT  5.5625 9.85 5.9125 9.915 ;
        RECT  5.5625 10.38 6.0875 10.445 ;
        RECT  5.5625 11.735 6.2625 11.8 ;
        RECT  5.5625 11.205 5.7375 11.27 ;
        RECT  5.5625 12.54 5.9125 12.605 ;
        RECT  5.5625 12.54 7.6275 12.605 ;
        RECT  5.5625 13.07 5.7375 13.135 ;
        RECT  5.5625 13.07 7.4525 13.135 ;
        RECT  5.5625 8.1025 6.4375 8.1675 ;
        RECT  5.5625 9.4475 6.6125 9.5125 ;
        RECT  5.5625 10.7925 6.4375 10.8575 ;
        RECT  5.5625 12.1375 6.6125 12.2025 ;
        RECT  5.5625 13.4825 6.4375 13.5475 ;
        RECT  6.3725 13.305 6.4375 13.4825 ;
        RECT  6.7175 8.1025 7.2775 8.1675 ;
        RECT  6.7175 6.7575 7.2775 6.8225 ;
        RECT  6.785 6.8225 6.85 7.0725 ;
        RECT  6.785 7.9675 6.85 8.1025 ;
        RECT  7.145 8.0325 7.21 8.1025 ;
        RECT  7.145 6.8225 7.21 6.9375 ;
        RECT  6.955 6.9375 7.02 8.0 ;
        RECT  7.2425 7.475 7.2775 7.54 ;
        RECT  6.7175 7.475 6.955 7.54 ;
        RECT  7.145 7.7625 7.21 7.8975 ;
        RECT  6.955 7.7625 7.02 7.8975 ;
        RECT  7.145 6.9375 7.21 7.0725 ;
        RECT  6.955 6.9375 7.02 7.0725 ;
        RECT  6.785 6.9375 6.85 7.0725 ;
        RECT  6.785 7.8975 6.85 8.0325 ;
        RECT  7.1075 7.475 7.2425 7.54 ;
        RECT  6.7175 10.7925 7.2775 10.8575 ;
        RECT  6.7175 12.1375 7.2775 12.2025 ;
        RECT  6.785 11.8875 6.85 12.1375 ;
        RECT  6.785 10.8575 6.85 10.9925 ;
        RECT  7.145 10.8575 7.21 10.9275 ;
        RECT  7.145 12.0225 7.21 12.1375 ;
        RECT  6.955 10.96 7.02 12.0225 ;
        RECT  7.2425 11.42 7.2775 11.485 ;
        RECT  6.7175 11.42 6.955 11.485 ;
        RECT  7.145 10.9925 7.21 11.1275 ;
        RECT  6.955 10.9925 7.02 11.1275 ;
        RECT  7.145 11.5975 7.21 11.7325 ;
        RECT  6.955 11.5975 7.02 11.7325 ;
        RECT  6.785 11.7525 6.85 11.8875 ;
        RECT  6.785 10.7925 6.85 10.9275 ;
        RECT  7.1075 11.345 7.2425 11.41 ;
        RECT  4.2525 8.1025 4.8125 8.1675 ;
        RECT  4.2525 6.7575 4.8125 6.8225 ;
        RECT  4.32 6.8225 4.385 7.0725 ;
        RECT  4.32 7.9675 4.385 8.1025 ;
        RECT  4.68 8.0325 4.745 8.1025 ;
        RECT  4.68 6.8225 4.745 6.9375 ;
        RECT  4.49 6.9375 4.555 8.0 ;
        RECT  4.7775 7.475 4.8125 7.54 ;
        RECT  4.2525 7.475 4.49 7.54 ;
        RECT  4.68 7.7625 4.745 7.8975 ;
        RECT  4.49 7.7625 4.555 7.8975 ;
        RECT  4.68 6.9375 4.745 7.0725 ;
        RECT  4.49 6.9375 4.555 7.0725 ;
        RECT  4.32 6.9375 4.385 7.0725 ;
        RECT  4.32 7.8975 4.385 8.0325 ;
        RECT  4.6425 7.475 4.7775 7.54 ;
        RECT  4.2525 10.7925 4.8125 10.8575 ;
        RECT  4.2525 12.1375 4.8125 12.2025 ;
        RECT  4.32 11.8875 4.385 12.1375 ;
        RECT  4.32 10.8575 4.385 10.9925 ;
        RECT  4.68 10.8575 4.745 10.9275 ;
        RECT  4.68 12.0225 4.745 12.1375 ;
        RECT  4.49 10.96 4.555 12.0225 ;
        RECT  4.7775 11.42 4.8125 11.485 ;
        RECT  4.2525 11.42 4.49 11.485 ;
        RECT  4.68 10.9925 4.745 11.1275 ;
        RECT  4.49 10.9925 4.555 11.1275 ;
        RECT  4.68 11.5975 4.745 11.7325 ;
        RECT  4.49 11.5975 4.555 11.7325 ;
        RECT  4.32 11.7525 4.385 11.8875 ;
        RECT  4.32 10.7925 4.385 10.9275 ;
        RECT  4.6425 11.345 4.7775 11.41 ;
        RECT  4.2525 10.7925 4.8125 10.8575 ;
        RECT  4.2525 9.4475 4.8125 9.5125 ;
        RECT  4.32 9.5125 4.385 9.7625 ;
        RECT  4.32 10.6575 4.385 10.7925 ;
        RECT  4.68 10.7225 4.745 10.7925 ;
        RECT  4.68 9.5125 4.745 9.6275 ;
        RECT  4.49 9.6275 4.555 10.69 ;
        RECT  4.7775 10.165 4.8125 10.23 ;
        RECT  4.2525 10.165 4.49 10.23 ;
        RECT  4.68 10.4525 4.745 10.5875 ;
        RECT  4.49 10.4525 4.555 10.5875 ;
        RECT  4.68 9.6275 4.745 9.7625 ;
        RECT  4.49 9.6275 4.555 9.7625 ;
        RECT  4.32 9.6275 4.385 9.7625 ;
        RECT  4.32 10.5875 4.385 10.7225 ;
        RECT  4.6425 10.165 4.7775 10.23 ;
        RECT  4.2525 13.4825 4.8125 13.5475 ;
        RECT  4.2525 14.8275 4.8125 14.8925 ;
        RECT  4.32 14.5775 4.385 14.8275 ;
        RECT  4.32 13.5475 4.385 13.6825 ;
        RECT  4.68 13.5475 4.745 13.6175 ;
        RECT  4.68 14.7125 4.745 14.8275 ;
        RECT  4.49 13.65 4.555 14.7125 ;
        RECT  4.7775 14.11 4.8125 14.175 ;
        RECT  4.2525 14.11 4.49 14.175 ;
        RECT  4.68 13.6825 4.745 13.8175 ;
        RECT  4.49 13.6825 4.555 13.8175 ;
        RECT  4.68 14.2875 4.745 14.4225 ;
        RECT  4.49 14.2875 4.555 14.4225 ;
        RECT  4.32 14.4425 4.385 14.5775 ;
        RECT  4.32 13.4825 4.385 13.6175 ;
        RECT  4.6425 14.035 4.7775 14.1 ;
        RECT  4.8125 8.1025 5.5625 8.1675 ;
        RECT  4.8125 6.7575 5.5625 6.8225 ;
        RECT  4.88 6.79 4.945 7.0725 ;
        RECT  4.88 7.955 4.945 8.135 ;
        RECT  5.43 6.79 5.495 7.0725 ;
        RECT  5.05 6.79 5.115 7.0725 ;
        RECT  5.43 7.8525 5.495 8.135 ;
        RECT  5.0175 7.175 5.0825 7.24 ;
        RECT  5.24 7.175 5.305 7.24 ;
        RECT  5.0175 7.2075 5.0825 7.9875 ;
        RECT  5.05 7.175 5.2725 7.24 ;
        RECT  5.24 7.0725 5.305 7.2075 ;
        RECT  5.5275 7.16 5.5625 7.225 ;
        RECT  5.2875 7.69 5.5625 7.755 ;
        RECT  4.8125 7.4725 5.05 7.5375 ;
        RECT  5.43 7.7175 5.495 7.8525 ;
        RECT  5.24 7.7175 5.305 7.8525 ;
        RECT  5.24 7.7175 5.305 7.8525 ;
        RECT  5.05 7.7175 5.115 7.8525 ;
        RECT  5.43 6.9375 5.495 7.0725 ;
        RECT  5.24 6.9375 5.305 7.0725 ;
        RECT  5.24 6.9375 5.305 7.0725 ;
        RECT  5.05 6.9375 5.115 7.0725 ;
        RECT  4.88 6.9375 4.945 7.0725 ;
        RECT  4.88 7.8525 4.945 7.9875 ;
        RECT  5.3925 7.16 5.5275 7.225 ;
        RECT  5.1525 7.69 5.2875 7.755 ;
        RECT  4.8125 10.7925 5.5625 10.8575 ;
        RECT  4.8125 12.1375 5.5625 12.2025 ;
        RECT  4.88 11.8875 4.945 12.17 ;
        RECT  4.88 10.825 4.945 11.005 ;
        RECT  5.43 11.8875 5.495 12.17 ;
        RECT  5.05 11.8875 5.115 12.17 ;
        RECT  5.43 10.825 5.495 11.1075 ;
        RECT  5.0175 11.72 5.0825 11.785 ;
        RECT  5.24 11.72 5.305 11.785 ;
        RECT  5.0175 10.9725 5.0825 11.7525 ;
        RECT  5.05 11.72 5.2725 11.785 ;
        RECT  5.24 11.7525 5.305 11.8875 ;
        RECT  5.5275 11.735 5.5625 11.8 ;
        RECT  5.2875 11.205 5.5625 11.27 ;
        RECT  4.8125 11.4225 5.05 11.4875 ;
        RECT  5.43 11.1275 5.495 11.2625 ;
        RECT  5.24 11.1275 5.305 11.2625 ;
        RECT  5.24 11.1275 5.305 11.2625 ;
        RECT  5.05 11.1275 5.115 11.2625 ;
        RECT  5.43 11.5975 5.495 11.7325 ;
        RECT  5.24 11.5975 5.305 11.7325 ;
        RECT  5.24 11.5975 5.305 11.7325 ;
        RECT  5.05 11.5975 5.115 11.7325 ;
        RECT  4.88 11.7525 4.945 11.8875 ;
        RECT  4.88 10.8375 4.945 10.9725 ;
        RECT  5.3925 11.66 5.5275 11.725 ;
        RECT  5.1525 11.13 5.2875 11.195 ;
        RECT  4.8125 10.7925 5.5625 10.8575 ;
        RECT  4.8125 9.4475 5.5625 9.5125 ;
        RECT  4.88 9.48 4.945 9.7625 ;
        RECT  4.88 10.645 4.945 10.825 ;
        RECT  5.43 9.48 5.495 9.7625 ;
        RECT  5.05 9.48 5.115 9.7625 ;
        RECT  5.43 10.5425 5.495 10.825 ;
        RECT  5.0175 9.865 5.0825 9.93 ;
        RECT  5.24 9.865 5.305 9.93 ;
        RECT  5.0175 9.8975 5.0825 10.6775 ;
        RECT  5.05 9.865 5.2725 9.93 ;
        RECT  5.24 9.7625 5.305 9.8975 ;
        RECT  5.5275 9.85 5.5625 9.915 ;
        RECT  5.2875 10.38 5.5625 10.445 ;
        RECT  4.8125 10.1625 5.05 10.2275 ;
        RECT  5.43 10.4075 5.495 10.5425 ;
        RECT  5.24 10.4075 5.305 10.5425 ;
        RECT  5.24 10.4075 5.305 10.5425 ;
        RECT  5.05 10.4075 5.115 10.5425 ;
        RECT  5.43 9.6275 5.495 9.7625 ;
        RECT  5.24 9.6275 5.305 9.7625 ;
        RECT  5.24 9.6275 5.305 9.7625 ;
        RECT  5.05 9.6275 5.115 9.7625 ;
        RECT  4.88 9.6275 4.945 9.7625 ;
        RECT  4.88 10.5425 4.945 10.6775 ;
        RECT  5.3925 9.85 5.5275 9.915 ;
        RECT  5.1525 10.38 5.2875 10.445 ;
        RECT  4.8125 13.4825 5.5625 13.5475 ;
        RECT  4.8125 14.8275 5.5625 14.8925 ;
        RECT  4.88 14.5775 4.945 14.86 ;
        RECT  4.88 13.515 4.945 13.695 ;
        RECT  5.43 14.5775 5.495 14.86 ;
        RECT  5.05 14.5775 5.115 14.86 ;
        RECT  5.43 13.515 5.495 13.7975 ;
        RECT  5.0175 14.41 5.0825 14.475 ;
        RECT  5.24 14.41 5.305 14.475 ;
        RECT  5.0175 13.6625 5.0825 14.4425 ;
        RECT  5.05 14.41 5.2725 14.475 ;
        RECT  5.24 14.4425 5.305 14.5775 ;
        RECT  5.5275 14.425 5.5625 14.49 ;
        RECT  5.2875 13.895 5.5625 13.96 ;
        RECT  4.8125 14.1125 5.05 14.1775 ;
        RECT  5.43 13.8175 5.495 13.9525 ;
        RECT  5.24 13.8175 5.305 13.9525 ;
        RECT  5.24 13.8175 5.305 13.9525 ;
        RECT  5.05 13.8175 5.115 13.9525 ;
        RECT  5.43 14.2875 5.495 14.4225 ;
        RECT  5.24 14.2875 5.305 14.4225 ;
        RECT  5.24 14.2875 5.305 14.4225 ;
        RECT  5.05 14.2875 5.115 14.4225 ;
        RECT  4.88 14.4425 4.945 14.5775 ;
        RECT  4.88 13.5275 4.945 13.6625 ;
        RECT  5.3925 14.35 5.5275 14.415 ;
        RECT  5.1525 13.82 5.2875 13.885 ;
        RECT  6.1575 9.1825 6.2925 9.2475 ;
        RECT  7.5225 8.66 7.6575 8.725 ;
        RECT  5.9825 9.5725 6.1175 9.6375 ;
        RECT  7.3475 10.095 7.4825 10.16 ;
        RECT  6.1575 8.975 6.2925 9.04 ;
        RECT  5.9825 8.445 6.1175 8.51 ;
        RECT  5.8075 9.78 5.9425 9.845 ;
        RECT  5.9825 10.31 6.1175 10.375 ;
        RECT  6.1575 11.665 6.2925 11.73 ;
        RECT  5.6325 11.135 5.7675 11.2 ;
        RECT  5.8075 12.47 5.9425 12.535 ;
        RECT  7.5225 12.47 7.6575 12.535 ;
        RECT  5.6325 13.0 5.7675 13.065 ;
        RECT  7.3475 13.0 7.4825 13.065 ;
        RECT  6.3325 8.0325 6.4675 8.0975 ;
        RECT  6.5075 9.3775 6.6425 9.4425 ;
        RECT  6.3325 10.7225 6.4675 10.7875 ;
        RECT  6.5075 12.0675 6.6425 12.1325 ;
        RECT  6.3325 13.235 6.4675 13.3 ;
        RECT  4.7475 14.1125 4.8125 14.1775 ;
        RECT  4.7475 15.5425 4.8125 15.6075 ;
        RECT  4.7475 16.8025 4.8125 16.8675 ;
        RECT  4.7475 18.2325 4.8125 18.2975 ;
        RECT  6.6525 14.11 6.7175 14.6975 ;
        RECT  6.1925 14.6325 6.7175 14.6975 ;
        RECT  7.2075 14.11 7.6275 14.175 ;
        RECT  6.5425 14.8275 7.2775 14.8925 ;
        RECT  6.3675 13.4825 7.2775 13.5475 ;
        RECT  6.6525 15.0225 6.7175 15.61 ;
        RECT  6.0175 15.0225 6.7175 15.0875 ;
        RECT  7.2075 15.545 7.4525 15.61 ;
        RECT  6.5425 14.8275 7.2775 14.8925 ;
        RECT  6.3675 16.1725 7.2775 16.2375 ;
        RECT  5.5625 14.425 6.2625 14.49 ;
        RECT  5.5625 13.895 6.0875 13.96 ;
        RECT  5.5625 15.23 5.9125 15.295 ;
        RECT  5.5625 15.76 6.0875 15.825 ;
        RECT  5.5625 17.115 6.2625 17.18 ;
        RECT  5.5625 16.585 5.7375 16.65 ;
        RECT  5.5625 17.92 5.9125 17.985 ;
        RECT  5.5625 17.92 7.6275 17.985 ;
        RECT  5.5625 18.45 5.7375 18.515 ;
        RECT  5.5625 18.45 7.4525 18.515 ;
        RECT  5.5625 13.4825 6.4375 13.5475 ;
        RECT  5.5625 14.8275 6.6125 14.8925 ;
        RECT  5.5625 16.1725 6.4375 16.2375 ;
        RECT  5.5625 17.5175 6.6125 17.5825 ;
        RECT  5.5625 18.8625 6.4375 18.9275 ;
        RECT  6.3725 18.685 6.4375 18.8625 ;
        RECT  6.7175 13.4825 7.2775 13.5475 ;
        RECT  6.7175 12.1375 7.2775 12.2025 ;
        RECT  6.785 12.2025 6.85 12.4525 ;
        RECT  6.785 13.3475 6.85 13.4825 ;
        RECT  7.145 13.4125 7.21 13.4825 ;
        RECT  7.145 12.2025 7.21 12.3175 ;
        RECT  6.955 12.3175 7.02 13.38 ;
        RECT  7.2425 12.855 7.2775 12.92 ;
        RECT  6.7175 12.855 6.955 12.92 ;
        RECT  7.145 13.1425 7.21 13.2775 ;
        RECT  6.955 13.1425 7.02 13.2775 ;
        RECT  7.145 12.3175 7.21 12.4525 ;
        RECT  6.955 12.3175 7.02 12.4525 ;
        RECT  6.785 12.3175 6.85 12.4525 ;
        RECT  6.785 13.2775 6.85 13.4125 ;
        RECT  7.1075 12.855 7.2425 12.92 ;
        RECT  6.7175 16.1725 7.2775 16.2375 ;
        RECT  6.7175 17.5175 7.2775 17.5825 ;
        RECT  6.785 17.2675 6.85 17.5175 ;
        RECT  6.785 16.2375 6.85 16.3725 ;
        RECT  7.145 16.2375 7.21 16.3075 ;
        RECT  7.145 17.4025 7.21 17.5175 ;
        RECT  6.955 16.34 7.02 17.4025 ;
        RECT  7.2425 16.8 7.2775 16.865 ;
        RECT  6.7175 16.8 6.955 16.865 ;
        RECT  7.145 16.3725 7.21 16.5075 ;
        RECT  6.955 16.3725 7.02 16.5075 ;
        RECT  7.145 16.9775 7.21 17.1125 ;
        RECT  6.955 16.9775 7.02 17.1125 ;
        RECT  6.785 17.1325 6.85 17.2675 ;
        RECT  6.785 16.1725 6.85 16.3075 ;
        RECT  7.1075 16.725 7.2425 16.79 ;
        RECT  4.2525 13.4825 4.8125 13.5475 ;
        RECT  4.2525 12.1375 4.8125 12.2025 ;
        RECT  4.32 12.2025 4.385 12.4525 ;
        RECT  4.32 13.3475 4.385 13.4825 ;
        RECT  4.68 13.4125 4.745 13.4825 ;
        RECT  4.68 12.2025 4.745 12.3175 ;
        RECT  4.49 12.3175 4.555 13.38 ;
        RECT  4.7775 12.855 4.8125 12.92 ;
        RECT  4.2525 12.855 4.49 12.92 ;
        RECT  4.68 13.1425 4.745 13.2775 ;
        RECT  4.49 13.1425 4.555 13.2775 ;
        RECT  4.68 12.3175 4.745 12.4525 ;
        RECT  4.49 12.3175 4.555 12.4525 ;
        RECT  4.32 12.3175 4.385 12.4525 ;
        RECT  4.32 13.2775 4.385 13.4125 ;
        RECT  4.6425 12.855 4.7775 12.92 ;
        RECT  4.2525 16.1725 4.8125 16.2375 ;
        RECT  4.2525 17.5175 4.8125 17.5825 ;
        RECT  4.32 17.2675 4.385 17.5175 ;
        RECT  4.32 16.2375 4.385 16.3725 ;
        RECT  4.68 16.2375 4.745 16.3075 ;
        RECT  4.68 17.4025 4.745 17.5175 ;
        RECT  4.49 16.34 4.555 17.4025 ;
        RECT  4.7775 16.8 4.8125 16.865 ;
        RECT  4.2525 16.8 4.49 16.865 ;
        RECT  4.68 16.3725 4.745 16.5075 ;
        RECT  4.49 16.3725 4.555 16.5075 ;
        RECT  4.68 16.9775 4.745 17.1125 ;
        RECT  4.49 16.9775 4.555 17.1125 ;
        RECT  4.32 17.1325 4.385 17.2675 ;
        RECT  4.32 16.1725 4.385 16.3075 ;
        RECT  4.6425 16.725 4.7775 16.79 ;
        RECT  4.2525 16.1725 4.8125 16.2375 ;
        RECT  4.2525 14.8275 4.8125 14.8925 ;
        RECT  4.32 14.8925 4.385 15.1425 ;
        RECT  4.32 16.0375 4.385 16.1725 ;
        RECT  4.68 16.1025 4.745 16.1725 ;
        RECT  4.68 14.8925 4.745 15.0075 ;
        RECT  4.49 15.0075 4.555 16.07 ;
        RECT  4.7775 15.545 4.8125 15.61 ;
        RECT  4.2525 15.545 4.49 15.61 ;
        RECT  4.68 15.8325 4.745 15.9675 ;
        RECT  4.49 15.8325 4.555 15.9675 ;
        RECT  4.68 15.0075 4.745 15.1425 ;
        RECT  4.49 15.0075 4.555 15.1425 ;
        RECT  4.32 15.0075 4.385 15.1425 ;
        RECT  4.32 15.9675 4.385 16.1025 ;
        RECT  4.6425 15.545 4.7775 15.61 ;
        RECT  4.2525 18.8625 4.8125 18.9275 ;
        RECT  4.2525 20.2075 4.8125 20.2725 ;
        RECT  4.32 19.9575 4.385 20.2075 ;
        RECT  4.32 18.9275 4.385 19.0625 ;
        RECT  4.68 18.9275 4.745 18.9975 ;
        RECT  4.68 20.0925 4.745 20.2075 ;
        RECT  4.49 19.03 4.555 20.0925 ;
        RECT  4.7775 19.49 4.8125 19.555 ;
        RECT  4.2525 19.49 4.49 19.555 ;
        RECT  4.68 19.0625 4.745 19.1975 ;
        RECT  4.49 19.0625 4.555 19.1975 ;
        RECT  4.68 19.6675 4.745 19.8025 ;
        RECT  4.49 19.6675 4.555 19.8025 ;
        RECT  4.32 19.8225 4.385 19.9575 ;
        RECT  4.32 18.8625 4.385 18.9975 ;
        RECT  4.6425 19.415 4.7775 19.48 ;
        RECT  4.8125 13.4825 5.5625 13.5475 ;
        RECT  4.8125 12.1375 5.5625 12.2025 ;
        RECT  4.88 12.17 4.945 12.4525 ;
        RECT  4.88 13.335 4.945 13.515 ;
        RECT  5.43 12.17 5.495 12.4525 ;
        RECT  5.05 12.17 5.115 12.4525 ;
        RECT  5.43 13.2325 5.495 13.515 ;
        RECT  5.0175 12.555 5.0825 12.62 ;
        RECT  5.24 12.555 5.305 12.62 ;
        RECT  5.0175 12.5875 5.0825 13.3675 ;
        RECT  5.05 12.555 5.2725 12.62 ;
        RECT  5.24 12.4525 5.305 12.5875 ;
        RECT  5.5275 12.54 5.5625 12.605 ;
        RECT  5.2875 13.07 5.5625 13.135 ;
        RECT  4.8125 12.8525 5.05 12.9175 ;
        RECT  5.43 13.0975 5.495 13.2325 ;
        RECT  5.24 13.0975 5.305 13.2325 ;
        RECT  5.24 13.0975 5.305 13.2325 ;
        RECT  5.05 13.0975 5.115 13.2325 ;
        RECT  5.43 12.3175 5.495 12.4525 ;
        RECT  5.24 12.3175 5.305 12.4525 ;
        RECT  5.24 12.3175 5.305 12.4525 ;
        RECT  5.05 12.3175 5.115 12.4525 ;
        RECT  4.88 12.3175 4.945 12.4525 ;
        RECT  4.88 13.2325 4.945 13.3675 ;
        RECT  5.3925 12.54 5.5275 12.605 ;
        RECT  5.1525 13.07 5.2875 13.135 ;
        RECT  4.8125 16.1725 5.5625 16.2375 ;
        RECT  4.8125 17.5175 5.5625 17.5825 ;
        RECT  4.88 17.2675 4.945 17.55 ;
        RECT  4.88 16.205 4.945 16.385 ;
        RECT  5.43 17.2675 5.495 17.55 ;
        RECT  5.05 17.2675 5.115 17.55 ;
        RECT  5.43 16.205 5.495 16.4875 ;
        RECT  5.0175 17.1 5.0825 17.165 ;
        RECT  5.24 17.1 5.305 17.165 ;
        RECT  5.0175 16.3525 5.0825 17.1325 ;
        RECT  5.05 17.1 5.2725 17.165 ;
        RECT  5.24 17.1325 5.305 17.2675 ;
        RECT  5.5275 17.115 5.5625 17.18 ;
        RECT  5.2875 16.585 5.5625 16.65 ;
        RECT  4.8125 16.8025 5.05 16.8675 ;
        RECT  5.43 16.5075 5.495 16.6425 ;
        RECT  5.24 16.5075 5.305 16.6425 ;
        RECT  5.24 16.5075 5.305 16.6425 ;
        RECT  5.05 16.5075 5.115 16.6425 ;
        RECT  5.43 16.9775 5.495 17.1125 ;
        RECT  5.24 16.9775 5.305 17.1125 ;
        RECT  5.24 16.9775 5.305 17.1125 ;
        RECT  5.05 16.9775 5.115 17.1125 ;
        RECT  4.88 17.1325 4.945 17.2675 ;
        RECT  4.88 16.2175 4.945 16.3525 ;
        RECT  5.3925 17.04 5.5275 17.105 ;
        RECT  5.1525 16.51 5.2875 16.575 ;
        RECT  4.8125 16.1725 5.5625 16.2375 ;
        RECT  4.8125 14.8275 5.5625 14.8925 ;
        RECT  4.88 14.86 4.945 15.1425 ;
        RECT  4.88 16.025 4.945 16.205 ;
        RECT  5.43 14.86 5.495 15.1425 ;
        RECT  5.05 14.86 5.115 15.1425 ;
        RECT  5.43 15.9225 5.495 16.205 ;
        RECT  5.0175 15.245 5.0825 15.31 ;
        RECT  5.24 15.245 5.305 15.31 ;
        RECT  5.0175 15.2775 5.0825 16.0575 ;
        RECT  5.05 15.245 5.2725 15.31 ;
        RECT  5.24 15.1425 5.305 15.2775 ;
        RECT  5.5275 15.23 5.5625 15.295 ;
        RECT  5.2875 15.76 5.5625 15.825 ;
        RECT  4.8125 15.5425 5.05 15.6075 ;
        RECT  5.43 15.7875 5.495 15.9225 ;
        RECT  5.24 15.7875 5.305 15.9225 ;
        RECT  5.24 15.7875 5.305 15.9225 ;
        RECT  5.05 15.7875 5.115 15.9225 ;
        RECT  5.43 15.0075 5.495 15.1425 ;
        RECT  5.24 15.0075 5.305 15.1425 ;
        RECT  5.24 15.0075 5.305 15.1425 ;
        RECT  5.05 15.0075 5.115 15.1425 ;
        RECT  4.88 15.0075 4.945 15.1425 ;
        RECT  4.88 15.9225 4.945 16.0575 ;
        RECT  5.3925 15.23 5.5275 15.295 ;
        RECT  5.1525 15.76 5.2875 15.825 ;
        RECT  4.8125 18.8625 5.5625 18.9275 ;
        RECT  4.8125 20.2075 5.5625 20.2725 ;
        RECT  4.88 19.9575 4.945 20.24 ;
        RECT  4.88 18.895 4.945 19.075 ;
        RECT  5.43 19.9575 5.495 20.24 ;
        RECT  5.05 19.9575 5.115 20.24 ;
        RECT  5.43 18.895 5.495 19.1775 ;
        RECT  5.0175 19.79 5.0825 19.855 ;
        RECT  5.24 19.79 5.305 19.855 ;
        RECT  5.0175 19.0425 5.0825 19.8225 ;
        RECT  5.05 19.79 5.2725 19.855 ;
        RECT  5.24 19.8225 5.305 19.9575 ;
        RECT  5.5275 19.805 5.5625 19.87 ;
        RECT  5.2875 19.275 5.5625 19.34 ;
        RECT  4.8125 19.4925 5.05 19.5575 ;
        RECT  5.43 19.1975 5.495 19.3325 ;
        RECT  5.24 19.1975 5.305 19.3325 ;
        RECT  5.24 19.1975 5.305 19.3325 ;
        RECT  5.05 19.1975 5.115 19.3325 ;
        RECT  5.43 19.6675 5.495 19.8025 ;
        RECT  5.24 19.6675 5.305 19.8025 ;
        RECT  5.24 19.6675 5.305 19.8025 ;
        RECT  5.05 19.6675 5.115 19.8025 ;
        RECT  4.88 19.8225 4.945 19.9575 ;
        RECT  4.88 18.9075 4.945 19.0425 ;
        RECT  5.3925 19.73 5.5275 19.795 ;
        RECT  5.1525 19.2 5.2875 19.265 ;
        RECT  6.1575 14.5625 6.2925 14.6275 ;
        RECT  7.5225 14.04 7.6575 14.105 ;
        RECT  5.9825 14.9525 6.1175 15.0175 ;
        RECT  7.3475 15.475 7.4825 15.54 ;
        RECT  6.1575 14.355 6.2925 14.42 ;
        RECT  5.9825 13.825 6.1175 13.89 ;
        RECT  5.8075 15.16 5.9425 15.225 ;
        RECT  5.9825 15.69 6.1175 15.755 ;
        RECT  6.1575 17.045 6.2925 17.11 ;
        RECT  5.6325 16.515 5.7675 16.58 ;
        RECT  5.8075 17.85 5.9425 17.915 ;
        RECT  7.5225 17.85 7.6575 17.915 ;
        RECT  5.6325 18.38 5.7675 18.445 ;
        RECT  7.3475 18.38 7.4825 18.445 ;
        RECT  6.3325 13.4125 6.4675 13.4775 ;
        RECT  6.5075 14.7575 6.6425 14.8225 ;
        RECT  6.3325 16.1025 6.4675 16.1675 ;
        RECT  6.5075 17.4475 6.6425 17.5125 ;
        RECT  6.3325 18.615 6.4675 18.68 ;
        RECT  4.2525 18.8625 5.0025 18.9275 ;
        RECT  4.2525 20.2075 5.0025 20.2725 ;
        RECT  4.87 19.9575 4.935 20.24 ;
        RECT  4.87 18.895 4.935 19.075 ;
        RECT  4.32 19.9575 4.385 20.24 ;
        RECT  4.7 19.9575 4.765 20.24 ;
        RECT  4.32 18.895 4.385 19.1775 ;
        RECT  4.7325 19.79 4.7975 19.855 ;
        RECT  4.51 19.79 4.575 19.855 ;
        RECT  4.7325 19.0425 4.7975 19.8225 ;
        RECT  4.5425 19.79 4.765 19.855 ;
        RECT  4.51 19.8225 4.575 19.9575 ;
        RECT  4.2525 19.805 4.2875 19.87 ;
        RECT  4.2525 19.275 4.5275 19.34 ;
        RECT  4.765 19.4925 5.0025 19.5575 ;
        RECT  4.32 19.1775 4.385 19.3125 ;
        RECT  4.51 19.1775 4.575 19.3125 ;
        RECT  4.51 19.1775 4.575 19.3125 ;
        RECT  4.7 19.1775 4.765 19.3125 ;
        RECT  4.32 19.9575 4.385 20.0925 ;
        RECT  4.51 19.9575 4.575 20.0925 ;
        RECT  4.51 19.9575 4.575 20.0925 ;
        RECT  4.7 19.9575 4.765 20.0925 ;
        RECT  4.87 19.9575 4.935 20.0925 ;
        RECT  4.87 19.0425 4.935 19.1775 ;
        RECT  4.2875 19.805 4.4225 19.87 ;
        RECT  4.5275 19.275 4.6625 19.34 ;
        RECT  4.2525 21.5525 5.0025 21.6175 ;
        RECT  4.2525 20.2075 5.0025 20.2725 ;
        RECT  4.87 20.24 4.935 20.5225 ;
        RECT  4.87 21.405 4.935 21.585 ;
        RECT  4.32 20.24 4.385 20.5225 ;
        RECT  4.7 20.24 4.765 20.5225 ;
        RECT  4.32 21.3025 4.385 21.585 ;
        RECT  4.7325 20.625 4.7975 20.69 ;
        RECT  4.51 20.625 4.575 20.69 ;
        RECT  4.7325 20.6575 4.7975 21.4375 ;
        RECT  4.5425 20.625 4.765 20.69 ;
        RECT  4.51 20.5225 4.575 20.6575 ;
        RECT  4.2525 20.61 4.2875 20.675 ;
        RECT  4.2525 21.14 4.5275 21.205 ;
        RECT  4.765 20.9225 5.0025 20.9875 ;
        RECT  4.32 21.1475 4.385 21.2825 ;
        RECT  4.51 21.1475 4.575 21.2825 ;
        RECT  4.51 21.1475 4.575 21.2825 ;
        RECT  4.7 21.1475 4.765 21.2825 ;
        RECT  4.32 20.6775 4.385 20.8125 ;
        RECT  4.51 20.6775 4.575 20.8125 ;
        RECT  4.51 20.6775 4.575 20.8125 ;
        RECT  4.7 20.6775 4.765 20.8125 ;
        RECT  4.87 20.5225 4.935 20.6575 ;
        RECT  4.87 21.4375 4.935 21.5725 ;
        RECT  4.2875 20.685 4.4225 20.75 ;
        RECT  4.5275 21.215 4.6625 21.28 ;
        RECT  4.2525 21.5525 5.0025 21.6175 ;
        RECT  4.2525 22.8975 5.0025 22.9625 ;
        RECT  4.87 22.6475 4.935 22.93 ;
        RECT  4.87 21.585 4.935 21.765 ;
        RECT  4.32 22.6475 4.385 22.93 ;
        RECT  4.7 22.6475 4.765 22.93 ;
        RECT  4.32 21.585 4.385 21.8675 ;
        RECT  4.7325 22.48 4.7975 22.545 ;
        RECT  4.51 22.48 4.575 22.545 ;
        RECT  4.7325 21.7325 4.7975 22.5125 ;
        RECT  4.5425 22.48 4.765 22.545 ;
        RECT  4.51 22.5125 4.575 22.6475 ;
        RECT  4.2525 22.495 4.2875 22.56 ;
        RECT  4.2525 21.965 4.5275 22.03 ;
        RECT  4.765 22.1825 5.0025 22.2475 ;
        RECT  4.32 21.8675 4.385 22.0025 ;
        RECT  4.51 21.8675 4.575 22.0025 ;
        RECT  4.51 21.8675 4.575 22.0025 ;
        RECT  4.7 21.8675 4.765 22.0025 ;
        RECT  4.32 22.6475 4.385 22.7825 ;
        RECT  4.51 22.6475 4.575 22.7825 ;
        RECT  4.51 22.6475 4.575 22.7825 ;
        RECT  4.7 22.6475 4.765 22.7825 ;
        RECT  4.87 22.6475 4.935 22.7825 ;
        RECT  4.87 21.7325 4.935 21.8675 ;
        RECT  4.2875 22.495 4.4225 22.56 ;
        RECT  4.5275 21.965 4.6625 22.03 ;
        RECT  4.2525 24.2425 5.0025 24.3075 ;
        RECT  4.2525 22.8975 5.0025 22.9625 ;
        RECT  4.87 22.93 4.935 23.2125 ;
        RECT  4.87 24.095 4.935 24.275 ;
        RECT  4.32 22.93 4.385 23.2125 ;
        RECT  4.7 22.93 4.765 23.2125 ;
        RECT  4.32 23.9925 4.385 24.275 ;
        RECT  4.7325 23.315 4.7975 23.38 ;
        RECT  4.51 23.315 4.575 23.38 ;
        RECT  4.7325 23.3475 4.7975 24.1275 ;
        RECT  4.5425 23.315 4.765 23.38 ;
        RECT  4.51 23.2125 4.575 23.3475 ;
        RECT  4.2525 23.3 4.2875 23.365 ;
        RECT  4.2525 23.83 4.5275 23.895 ;
        RECT  4.765 23.6125 5.0025 23.6775 ;
        RECT  4.32 23.8375 4.385 23.9725 ;
        RECT  4.51 23.8375 4.575 23.9725 ;
        RECT  4.51 23.8375 4.575 23.9725 ;
        RECT  4.7 23.8375 4.765 23.9725 ;
        RECT  4.32 23.3675 4.385 23.5025 ;
        RECT  4.51 23.3675 4.575 23.5025 ;
        RECT  4.51 23.3675 4.575 23.5025 ;
        RECT  4.7 23.3675 4.765 23.5025 ;
        RECT  4.87 23.2125 4.935 23.3475 ;
        RECT  4.87 24.1275 4.935 24.2625 ;
        RECT  4.2875 23.375 4.4225 23.44 ;
        RECT  4.5275 23.905 4.6625 23.97 ;
        RECT  4.2525 24.2425 5.0025 24.3075 ;
        RECT  4.2525 25.5875 5.0025 25.6525 ;
        RECT  4.87 25.3375 4.935 25.62 ;
        RECT  4.87 24.275 4.935 24.455 ;
        RECT  4.32 25.3375 4.385 25.62 ;
        RECT  4.7 25.3375 4.765 25.62 ;
        RECT  4.32 24.275 4.385 24.5575 ;
        RECT  4.7325 25.17 4.7975 25.235 ;
        RECT  4.51 25.17 4.575 25.235 ;
        RECT  4.7325 24.4225 4.7975 25.2025 ;
        RECT  4.5425 25.17 4.765 25.235 ;
        RECT  4.51 25.2025 4.575 25.3375 ;
        RECT  4.2525 25.185 4.2875 25.25 ;
        RECT  4.2525 24.655 4.5275 24.72 ;
        RECT  4.765 24.8725 5.0025 24.9375 ;
        RECT  4.32 24.5575 4.385 24.6925 ;
        RECT  4.51 24.5575 4.575 24.6925 ;
        RECT  4.51 24.5575 4.575 24.6925 ;
        RECT  4.7 24.5575 4.765 24.6925 ;
        RECT  4.32 25.3375 4.385 25.4725 ;
        RECT  4.51 25.3375 4.575 25.4725 ;
        RECT  4.51 25.3375 4.575 25.4725 ;
        RECT  4.7 25.3375 4.765 25.4725 ;
        RECT  4.87 25.3375 4.935 25.4725 ;
        RECT  4.87 24.4225 4.935 24.5575 ;
        RECT  4.2875 25.185 4.4225 25.25 ;
        RECT  4.5275 24.655 4.6625 24.72 ;
        RECT  4.2525 26.9325 5.0025 26.9975 ;
        RECT  4.2525 25.5875 5.0025 25.6525 ;
        RECT  4.87 25.62 4.935 25.9025 ;
        RECT  4.87 26.785 4.935 26.965 ;
        RECT  4.32 25.62 4.385 25.9025 ;
        RECT  4.7 25.62 4.765 25.9025 ;
        RECT  4.32 26.6825 4.385 26.965 ;
        RECT  4.7325 26.005 4.7975 26.07 ;
        RECT  4.51 26.005 4.575 26.07 ;
        RECT  4.7325 26.0375 4.7975 26.8175 ;
        RECT  4.5425 26.005 4.765 26.07 ;
        RECT  4.51 25.9025 4.575 26.0375 ;
        RECT  4.2525 25.99 4.2875 26.055 ;
        RECT  4.2525 26.52 4.5275 26.585 ;
        RECT  4.765 26.3025 5.0025 26.3675 ;
        RECT  4.32 26.5275 4.385 26.6625 ;
        RECT  4.51 26.5275 4.575 26.6625 ;
        RECT  4.51 26.5275 4.575 26.6625 ;
        RECT  4.7 26.5275 4.765 26.6625 ;
        RECT  4.32 26.0575 4.385 26.1925 ;
        RECT  4.51 26.0575 4.575 26.1925 ;
        RECT  4.51 26.0575 4.575 26.1925 ;
        RECT  4.7 26.0575 4.765 26.1925 ;
        RECT  4.87 25.9025 4.935 26.0375 ;
        RECT  4.87 26.8175 4.935 26.9525 ;
        RECT  4.2875 26.065 4.4225 26.13 ;
        RECT  4.5275 26.595 4.6625 26.66 ;
        RECT  4.2525 26.9325 5.0025 26.9975 ;
        RECT  4.2525 28.2775 5.0025 28.3425 ;
        RECT  4.87 28.0275 4.935 28.31 ;
        RECT  4.87 26.965 4.935 27.145 ;
        RECT  4.32 28.0275 4.385 28.31 ;
        RECT  4.7 28.0275 4.765 28.31 ;
        RECT  4.32 26.965 4.385 27.2475 ;
        RECT  4.7325 27.86 4.7975 27.925 ;
        RECT  4.51 27.86 4.575 27.925 ;
        RECT  4.7325 27.1125 4.7975 27.8925 ;
        RECT  4.5425 27.86 4.765 27.925 ;
        RECT  4.51 27.8925 4.575 28.0275 ;
        RECT  4.2525 27.875 4.2875 27.94 ;
        RECT  4.2525 27.345 4.5275 27.41 ;
        RECT  4.765 27.5625 5.0025 27.6275 ;
        RECT  4.32 27.2475 4.385 27.3825 ;
        RECT  4.51 27.2475 4.575 27.3825 ;
        RECT  4.51 27.2475 4.575 27.3825 ;
        RECT  4.7 27.2475 4.765 27.3825 ;
        RECT  4.32 28.0275 4.385 28.1625 ;
        RECT  4.51 28.0275 4.575 28.1625 ;
        RECT  4.51 28.0275 4.575 28.1625 ;
        RECT  4.7 28.0275 4.765 28.1625 ;
        RECT  4.87 28.0275 4.935 28.1625 ;
        RECT  4.87 27.1125 4.935 27.2475 ;
        RECT  4.2875 27.875 4.4225 27.94 ;
        RECT  4.5275 27.345 4.6625 27.41 ;
        RECT  4.2525 29.6225 5.0025 29.6875 ;
        RECT  4.2525 28.2775 5.0025 28.3425 ;
        RECT  4.87 28.31 4.935 28.5925 ;
        RECT  4.87 29.475 4.935 29.655 ;
        RECT  4.32 28.31 4.385 28.5925 ;
        RECT  4.7 28.31 4.765 28.5925 ;
        RECT  4.32 29.3725 4.385 29.655 ;
        RECT  4.7325 28.695 4.7975 28.76 ;
        RECT  4.51 28.695 4.575 28.76 ;
        RECT  4.7325 28.7275 4.7975 29.5075 ;
        RECT  4.5425 28.695 4.765 28.76 ;
        RECT  4.51 28.5925 4.575 28.7275 ;
        RECT  4.2525 28.68 4.2875 28.745 ;
        RECT  4.2525 29.21 4.5275 29.275 ;
        RECT  4.765 28.9925 5.0025 29.0575 ;
        RECT  4.32 29.2175 4.385 29.3525 ;
        RECT  4.51 29.2175 4.575 29.3525 ;
        RECT  4.51 29.2175 4.575 29.3525 ;
        RECT  4.7 29.2175 4.765 29.3525 ;
        RECT  4.32 28.7475 4.385 28.8825 ;
        RECT  4.51 28.7475 4.575 28.8825 ;
        RECT  4.51 28.7475 4.575 28.8825 ;
        RECT  4.7 28.7475 4.765 28.8825 ;
        RECT  4.87 28.5925 4.935 28.7275 ;
        RECT  4.87 29.5075 4.935 29.6425 ;
        RECT  4.2875 28.755 4.4225 28.82 ;
        RECT  4.5275 29.285 4.6625 29.35 ;
        RECT  4.2525 29.6225 5.0025 29.6875 ;
        RECT  4.2525 30.9675 5.0025 31.0325 ;
        RECT  4.87 30.7175 4.935 31.0 ;
        RECT  4.87 29.655 4.935 29.835 ;
        RECT  4.32 30.7175 4.385 31.0 ;
        RECT  4.7 30.7175 4.765 31.0 ;
        RECT  4.32 29.655 4.385 29.9375 ;
        RECT  4.7325 30.55 4.7975 30.615 ;
        RECT  4.51 30.55 4.575 30.615 ;
        RECT  4.7325 29.8025 4.7975 30.5825 ;
        RECT  4.5425 30.55 4.765 30.615 ;
        RECT  4.51 30.5825 4.575 30.7175 ;
        RECT  4.2525 30.565 4.2875 30.63 ;
        RECT  4.2525 30.035 4.5275 30.1 ;
        RECT  4.765 30.2525 5.0025 30.3175 ;
        RECT  4.32 29.9375 4.385 30.0725 ;
        RECT  4.51 29.9375 4.575 30.0725 ;
        RECT  4.51 29.9375 4.575 30.0725 ;
        RECT  4.7 29.9375 4.765 30.0725 ;
        RECT  4.32 30.7175 4.385 30.8525 ;
        RECT  4.51 30.7175 4.575 30.8525 ;
        RECT  4.51 30.7175 4.575 30.8525 ;
        RECT  4.7 30.7175 4.765 30.8525 ;
        RECT  4.87 30.7175 4.935 30.8525 ;
        RECT  4.87 29.8025 4.935 29.9375 ;
        RECT  4.2875 30.565 4.4225 30.63 ;
        RECT  4.5275 30.035 4.6625 30.1 ;
        RECT  4.2525 32.3125 5.0025 32.3775 ;
        RECT  4.2525 30.9675 5.0025 31.0325 ;
        RECT  4.87 31.0 4.935 31.2825 ;
        RECT  4.87 32.165 4.935 32.345 ;
        RECT  4.32 31.0 4.385 31.2825 ;
        RECT  4.7 31.0 4.765 31.2825 ;
        RECT  4.32 32.0625 4.385 32.345 ;
        RECT  4.7325 31.385 4.7975 31.45 ;
        RECT  4.51 31.385 4.575 31.45 ;
        RECT  4.7325 31.4175 4.7975 32.1975 ;
        RECT  4.5425 31.385 4.765 31.45 ;
        RECT  4.51 31.2825 4.575 31.4175 ;
        RECT  4.2525 31.37 4.2875 31.435 ;
        RECT  4.2525 31.9 4.5275 31.965 ;
        RECT  4.765 31.6825 5.0025 31.7475 ;
        RECT  4.32 31.9075 4.385 32.0425 ;
        RECT  4.51 31.9075 4.575 32.0425 ;
        RECT  4.51 31.9075 4.575 32.0425 ;
        RECT  4.7 31.9075 4.765 32.0425 ;
        RECT  4.32 31.4375 4.385 31.5725 ;
        RECT  4.51 31.4375 4.575 31.5725 ;
        RECT  4.51 31.4375 4.575 31.5725 ;
        RECT  4.7 31.4375 4.765 31.5725 ;
        RECT  4.87 31.2825 4.935 31.4175 ;
        RECT  4.87 32.1975 4.935 32.3325 ;
        RECT  4.2875 31.445 4.4225 31.51 ;
        RECT  4.5275 31.975 4.6625 32.04 ;
        RECT  4.2525 32.3125 5.0025 32.3775 ;
        RECT  4.2525 33.6575 5.0025 33.7225 ;
        RECT  4.87 33.4075 4.935 33.69 ;
        RECT  4.87 32.345 4.935 32.525 ;
        RECT  4.32 33.4075 4.385 33.69 ;
        RECT  4.7 33.4075 4.765 33.69 ;
        RECT  4.32 32.345 4.385 32.6275 ;
        RECT  4.7325 33.24 4.7975 33.305 ;
        RECT  4.51 33.24 4.575 33.305 ;
        RECT  4.7325 32.4925 4.7975 33.2725 ;
        RECT  4.5425 33.24 4.765 33.305 ;
        RECT  4.51 33.2725 4.575 33.4075 ;
        RECT  4.2525 33.255 4.2875 33.32 ;
        RECT  4.2525 32.725 4.5275 32.79 ;
        RECT  4.765 32.9425 5.0025 33.0075 ;
        RECT  4.32 32.6275 4.385 32.7625 ;
        RECT  4.51 32.6275 4.575 32.7625 ;
        RECT  4.51 32.6275 4.575 32.7625 ;
        RECT  4.7 32.6275 4.765 32.7625 ;
        RECT  4.32 33.4075 4.385 33.5425 ;
        RECT  4.51 33.4075 4.575 33.5425 ;
        RECT  4.51 33.4075 4.575 33.5425 ;
        RECT  4.7 33.4075 4.765 33.5425 ;
        RECT  4.87 33.4075 4.935 33.5425 ;
        RECT  4.87 32.4925 4.935 32.6275 ;
        RECT  4.2875 33.255 4.4225 33.32 ;
        RECT  4.5275 32.725 4.6625 32.79 ;
        RECT  4.2525 35.0025 5.0025 35.0675 ;
        RECT  4.2525 33.6575 5.0025 33.7225 ;
        RECT  4.87 33.69 4.935 33.9725 ;
        RECT  4.87 34.855 4.935 35.035 ;
        RECT  4.32 33.69 4.385 33.9725 ;
        RECT  4.7 33.69 4.765 33.9725 ;
        RECT  4.32 34.7525 4.385 35.035 ;
        RECT  4.7325 34.075 4.7975 34.14 ;
        RECT  4.51 34.075 4.575 34.14 ;
        RECT  4.7325 34.1075 4.7975 34.8875 ;
        RECT  4.5425 34.075 4.765 34.14 ;
        RECT  4.51 33.9725 4.575 34.1075 ;
        RECT  4.2525 34.06 4.2875 34.125 ;
        RECT  4.2525 34.59 4.5275 34.655 ;
        RECT  4.765 34.3725 5.0025 34.4375 ;
        RECT  4.32 34.5975 4.385 34.7325 ;
        RECT  4.51 34.5975 4.575 34.7325 ;
        RECT  4.51 34.5975 4.575 34.7325 ;
        RECT  4.7 34.5975 4.765 34.7325 ;
        RECT  4.32 34.1275 4.385 34.2625 ;
        RECT  4.51 34.1275 4.575 34.2625 ;
        RECT  4.51 34.1275 4.575 34.2625 ;
        RECT  4.7 34.1275 4.765 34.2625 ;
        RECT  4.87 33.9725 4.935 34.1075 ;
        RECT  4.87 34.8875 4.935 35.0225 ;
        RECT  4.2875 34.135 4.4225 34.2 ;
        RECT  4.5275 34.665 4.6625 34.73 ;
        RECT  4.2525 35.0025 5.0025 35.0675 ;
        RECT  4.2525 36.3475 5.0025 36.4125 ;
        RECT  4.87 36.0975 4.935 36.38 ;
        RECT  4.87 35.035 4.935 35.215 ;
        RECT  4.32 36.0975 4.385 36.38 ;
        RECT  4.7 36.0975 4.765 36.38 ;
        RECT  4.32 35.035 4.385 35.3175 ;
        RECT  4.7325 35.93 4.7975 35.995 ;
        RECT  4.51 35.93 4.575 35.995 ;
        RECT  4.7325 35.1825 4.7975 35.9625 ;
        RECT  4.5425 35.93 4.765 35.995 ;
        RECT  4.51 35.9625 4.575 36.0975 ;
        RECT  4.2525 35.945 4.2875 36.01 ;
        RECT  4.2525 35.415 4.5275 35.48 ;
        RECT  4.765 35.6325 5.0025 35.6975 ;
        RECT  4.32 35.3175 4.385 35.4525 ;
        RECT  4.51 35.3175 4.575 35.4525 ;
        RECT  4.51 35.3175 4.575 35.4525 ;
        RECT  4.7 35.3175 4.765 35.4525 ;
        RECT  4.32 36.0975 4.385 36.2325 ;
        RECT  4.51 36.0975 4.575 36.2325 ;
        RECT  4.51 36.0975 4.575 36.2325 ;
        RECT  4.7 36.0975 4.765 36.2325 ;
        RECT  4.87 36.0975 4.935 36.2325 ;
        RECT  4.87 35.1825 4.935 35.3175 ;
        RECT  4.2875 35.945 4.4225 36.01 ;
        RECT  4.5275 35.415 4.6625 35.48 ;
        RECT  4.2525 37.6925 5.0025 37.7575 ;
        RECT  4.2525 36.3475 5.0025 36.4125 ;
        RECT  4.87 36.38 4.935 36.6625 ;
        RECT  4.87 37.545 4.935 37.725 ;
        RECT  4.32 36.38 4.385 36.6625 ;
        RECT  4.7 36.38 4.765 36.6625 ;
        RECT  4.32 37.4425 4.385 37.725 ;
        RECT  4.7325 36.765 4.7975 36.83 ;
        RECT  4.51 36.765 4.575 36.83 ;
        RECT  4.7325 36.7975 4.7975 37.5775 ;
        RECT  4.5425 36.765 4.765 36.83 ;
        RECT  4.51 36.6625 4.575 36.7975 ;
        RECT  4.2525 36.75 4.2875 36.815 ;
        RECT  4.2525 37.28 4.5275 37.345 ;
        RECT  4.765 37.0625 5.0025 37.1275 ;
        RECT  4.32 37.2875 4.385 37.4225 ;
        RECT  4.51 37.2875 4.575 37.4225 ;
        RECT  4.51 37.2875 4.575 37.4225 ;
        RECT  4.7 37.2875 4.765 37.4225 ;
        RECT  4.32 36.8175 4.385 36.9525 ;
        RECT  4.51 36.8175 4.575 36.9525 ;
        RECT  4.51 36.8175 4.575 36.9525 ;
        RECT  4.7 36.8175 4.765 36.9525 ;
        RECT  4.87 36.6625 4.935 36.7975 ;
        RECT  4.87 37.5775 4.935 37.7125 ;
        RECT  4.2875 36.825 4.4225 36.89 ;
        RECT  4.5275 37.355 4.6625 37.42 ;
        RECT  4.2525 37.6925 5.0025 37.7575 ;
        RECT  4.2525 39.0375 5.0025 39.1025 ;
        RECT  4.87 38.7875 4.935 39.07 ;
        RECT  4.87 37.725 4.935 37.905 ;
        RECT  4.32 38.7875 4.385 39.07 ;
        RECT  4.7 38.7875 4.765 39.07 ;
        RECT  4.32 37.725 4.385 38.0075 ;
        RECT  4.7325 38.62 4.7975 38.685 ;
        RECT  4.51 38.62 4.575 38.685 ;
        RECT  4.7325 37.8725 4.7975 38.6525 ;
        RECT  4.5425 38.62 4.765 38.685 ;
        RECT  4.51 38.6525 4.575 38.7875 ;
        RECT  4.2525 38.635 4.2875 38.7 ;
        RECT  4.2525 38.105 4.5275 38.17 ;
        RECT  4.765 38.3225 5.0025 38.3875 ;
        RECT  4.32 38.0075 4.385 38.1425 ;
        RECT  4.51 38.0075 4.575 38.1425 ;
        RECT  4.51 38.0075 4.575 38.1425 ;
        RECT  4.7 38.0075 4.765 38.1425 ;
        RECT  4.32 38.7875 4.385 38.9225 ;
        RECT  4.51 38.7875 4.575 38.9225 ;
        RECT  4.51 38.7875 4.575 38.9225 ;
        RECT  4.7 38.7875 4.765 38.9225 ;
        RECT  4.87 38.7875 4.935 38.9225 ;
        RECT  4.87 37.8725 4.935 38.0075 ;
        RECT  4.2875 38.635 4.4225 38.7 ;
        RECT  4.5275 38.105 4.6625 38.17 ;
        RECT  4.2525 40.3825 5.0025 40.4475 ;
        RECT  4.2525 39.0375 5.0025 39.1025 ;
        RECT  4.87 39.07 4.935 39.3525 ;
        RECT  4.87 40.235 4.935 40.415 ;
        RECT  4.32 39.07 4.385 39.3525 ;
        RECT  4.7 39.07 4.765 39.3525 ;
        RECT  4.32 40.1325 4.385 40.415 ;
        RECT  4.7325 39.455 4.7975 39.52 ;
        RECT  4.51 39.455 4.575 39.52 ;
        RECT  4.7325 39.4875 4.7975 40.2675 ;
        RECT  4.5425 39.455 4.765 39.52 ;
        RECT  4.51 39.3525 4.575 39.4875 ;
        RECT  4.2525 39.44 4.2875 39.505 ;
        RECT  4.2525 39.97 4.5275 40.035 ;
        RECT  4.765 39.7525 5.0025 39.8175 ;
        RECT  4.32 39.9775 4.385 40.1125 ;
        RECT  4.51 39.9775 4.575 40.1125 ;
        RECT  4.51 39.9775 4.575 40.1125 ;
        RECT  4.7 39.9775 4.765 40.1125 ;
        RECT  4.32 39.5075 4.385 39.6425 ;
        RECT  4.51 39.5075 4.575 39.6425 ;
        RECT  4.51 39.5075 4.575 39.6425 ;
        RECT  4.7 39.5075 4.765 39.6425 ;
        RECT  4.87 39.3525 4.935 39.4875 ;
        RECT  4.87 40.2675 4.935 40.4025 ;
        RECT  4.2875 39.515 4.4225 39.58 ;
        RECT  4.5275 40.045 4.6625 40.11 ;
        RECT  5.0025 18.8625 5.5625 18.9275 ;
        RECT  5.0025 20.2075 5.5625 20.2725 ;
        RECT  5.43 19.9575 5.495 20.2075 ;
        RECT  5.43 18.9275 5.495 19.0625 ;
        RECT  5.07 18.9275 5.135 18.9975 ;
        RECT  5.07 20.0925 5.135 20.2075 ;
        RECT  5.26 19.03 5.325 20.0925 ;
        RECT  5.0025 19.49 5.0375 19.555 ;
        RECT  5.325 19.49 5.5625 19.555 ;
        RECT  5.07 19.1325 5.135 19.2675 ;
        RECT  5.26 19.1325 5.325 19.2675 ;
        RECT  5.07 19.9575 5.135 20.0925 ;
        RECT  5.26 19.9575 5.325 20.0925 ;
        RECT  5.43 19.9575 5.495 20.0925 ;
        RECT  5.43 18.9975 5.495 19.1325 ;
        RECT  5.0375 19.49 5.1725 19.555 ;
        RECT  5.0025 21.5525 5.5625 21.6175 ;
        RECT  5.0025 20.2075 5.5625 20.2725 ;
        RECT  5.43 20.2725 5.495 20.5225 ;
        RECT  5.43 21.4175 5.495 21.5525 ;
        RECT  5.07 21.4825 5.135 21.5525 ;
        RECT  5.07 20.2725 5.135 20.3875 ;
        RECT  5.26 20.3875 5.325 21.45 ;
        RECT  5.0025 20.925 5.0375 20.99 ;
        RECT  5.325 20.925 5.5625 20.99 ;
        RECT  5.07 21.2825 5.135 21.4175 ;
        RECT  5.26 21.2825 5.325 21.4175 ;
        RECT  5.07 20.6775 5.135 20.8125 ;
        RECT  5.26 20.6775 5.325 20.8125 ;
        RECT  5.43 20.5225 5.495 20.6575 ;
        RECT  5.43 21.4825 5.495 21.6175 ;
        RECT  5.0375 21.0 5.1725 21.065 ;
        RECT  5.0025 21.5525 5.5625 21.6175 ;
        RECT  5.0025 22.8975 5.5625 22.9625 ;
        RECT  5.43 22.6475 5.495 22.8975 ;
        RECT  5.43 21.6175 5.495 21.7525 ;
        RECT  5.07 21.6175 5.135 21.6875 ;
        RECT  5.07 22.7825 5.135 22.8975 ;
        RECT  5.26 21.72 5.325 22.7825 ;
        RECT  5.0025 22.18 5.0375 22.245 ;
        RECT  5.325 22.18 5.5625 22.245 ;
        RECT  5.07 21.8225 5.135 21.9575 ;
        RECT  5.26 21.8225 5.325 21.9575 ;
        RECT  5.07 22.6475 5.135 22.7825 ;
        RECT  5.26 22.6475 5.325 22.7825 ;
        RECT  5.43 22.6475 5.495 22.7825 ;
        RECT  5.43 21.6875 5.495 21.8225 ;
        RECT  5.0375 22.18 5.1725 22.245 ;
        RECT  5.0025 24.2425 5.5625 24.3075 ;
        RECT  5.0025 22.8975 5.5625 22.9625 ;
        RECT  5.43 22.9625 5.495 23.2125 ;
        RECT  5.43 24.1075 5.495 24.2425 ;
        RECT  5.07 24.1725 5.135 24.2425 ;
        RECT  5.07 22.9625 5.135 23.0775 ;
        RECT  5.26 23.0775 5.325 24.14 ;
        RECT  5.0025 23.615 5.0375 23.68 ;
        RECT  5.325 23.615 5.5625 23.68 ;
        RECT  5.07 23.9725 5.135 24.1075 ;
        RECT  5.26 23.9725 5.325 24.1075 ;
        RECT  5.07 23.3675 5.135 23.5025 ;
        RECT  5.26 23.3675 5.325 23.5025 ;
        RECT  5.43 23.2125 5.495 23.3475 ;
        RECT  5.43 24.1725 5.495 24.3075 ;
        RECT  5.0375 23.69 5.1725 23.755 ;
        RECT  5.0025 24.2425 5.5625 24.3075 ;
        RECT  5.0025 25.5875 5.5625 25.6525 ;
        RECT  5.43 25.3375 5.495 25.5875 ;
        RECT  5.43 24.3075 5.495 24.4425 ;
        RECT  5.07 24.3075 5.135 24.3775 ;
        RECT  5.07 25.4725 5.135 25.5875 ;
        RECT  5.26 24.41 5.325 25.4725 ;
        RECT  5.0025 24.87 5.0375 24.935 ;
        RECT  5.325 24.87 5.5625 24.935 ;
        RECT  5.07 24.5125 5.135 24.6475 ;
        RECT  5.26 24.5125 5.325 24.6475 ;
        RECT  5.07 25.3375 5.135 25.4725 ;
        RECT  5.26 25.3375 5.325 25.4725 ;
        RECT  5.43 25.3375 5.495 25.4725 ;
        RECT  5.43 24.3775 5.495 24.5125 ;
        RECT  5.0375 24.87 5.1725 24.935 ;
        RECT  5.0025 26.9325 5.5625 26.9975 ;
        RECT  5.0025 25.5875 5.5625 25.6525 ;
        RECT  5.43 25.6525 5.495 25.9025 ;
        RECT  5.43 26.7975 5.495 26.9325 ;
        RECT  5.07 26.8625 5.135 26.9325 ;
        RECT  5.07 25.6525 5.135 25.7675 ;
        RECT  5.26 25.7675 5.325 26.83 ;
        RECT  5.0025 26.305 5.0375 26.37 ;
        RECT  5.325 26.305 5.5625 26.37 ;
        RECT  5.07 26.6625 5.135 26.7975 ;
        RECT  5.26 26.6625 5.325 26.7975 ;
        RECT  5.07 26.0575 5.135 26.1925 ;
        RECT  5.26 26.0575 5.325 26.1925 ;
        RECT  5.43 25.9025 5.495 26.0375 ;
        RECT  5.43 26.8625 5.495 26.9975 ;
        RECT  5.0375 26.38 5.1725 26.445 ;
        RECT  5.0025 26.9325 5.5625 26.9975 ;
        RECT  5.0025 28.2775 5.5625 28.3425 ;
        RECT  5.43 28.0275 5.495 28.2775 ;
        RECT  5.43 26.9975 5.495 27.1325 ;
        RECT  5.07 26.9975 5.135 27.0675 ;
        RECT  5.07 28.1625 5.135 28.2775 ;
        RECT  5.26 27.1 5.325 28.1625 ;
        RECT  5.0025 27.56 5.0375 27.625 ;
        RECT  5.325 27.56 5.5625 27.625 ;
        RECT  5.07 27.2025 5.135 27.3375 ;
        RECT  5.26 27.2025 5.325 27.3375 ;
        RECT  5.07 28.0275 5.135 28.1625 ;
        RECT  5.26 28.0275 5.325 28.1625 ;
        RECT  5.43 28.0275 5.495 28.1625 ;
        RECT  5.43 27.0675 5.495 27.2025 ;
        RECT  5.0375 27.56 5.1725 27.625 ;
        RECT  5.0025 29.6225 5.5625 29.6875 ;
        RECT  5.0025 28.2775 5.5625 28.3425 ;
        RECT  5.43 28.3425 5.495 28.5925 ;
        RECT  5.43 29.4875 5.495 29.6225 ;
        RECT  5.07 29.5525 5.135 29.6225 ;
        RECT  5.07 28.3425 5.135 28.4575 ;
        RECT  5.26 28.4575 5.325 29.52 ;
        RECT  5.0025 28.995 5.0375 29.06 ;
        RECT  5.325 28.995 5.5625 29.06 ;
        RECT  5.07 29.3525 5.135 29.4875 ;
        RECT  5.26 29.3525 5.325 29.4875 ;
        RECT  5.07 28.7475 5.135 28.8825 ;
        RECT  5.26 28.7475 5.325 28.8825 ;
        RECT  5.43 28.5925 5.495 28.7275 ;
        RECT  5.43 29.5525 5.495 29.6875 ;
        RECT  5.0375 29.07 5.1725 29.135 ;
        RECT  5.0025 29.6225 5.5625 29.6875 ;
        RECT  5.0025 30.9675 5.5625 31.0325 ;
        RECT  5.43 30.7175 5.495 30.9675 ;
        RECT  5.43 29.6875 5.495 29.8225 ;
        RECT  5.07 29.6875 5.135 29.7575 ;
        RECT  5.07 30.8525 5.135 30.9675 ;
        RECT  5.26 29.79 5.325 30.8525 ;
        RECT  5.0025 30.25 5.0375 30.315 ;
        RECT  5.325 30.25 5.5625 30.315 ;
        RECT  5.07 29.8925 5.135 30.0275 ;
        RECT  5.26 29.8925 5.325 30.0275 ;
        RECT  5.07 30.7175 5.135 30.8525 ;
        RECT  5.26 30.7175 5.325 30.8525 ;
        RECT  5.43 30.7175 5.495 30.8525 ;
        RECT  5.43 29.7575 5.495 29.8925 ;
        RECT  5.0375 30.25 5.1725 30.315 ;
        RECT  5.0025 32.3125 5.5625 32.3775 ;
        RECT  5.0025 30.9675 5.5625 31.0325 ;
        RECT  5.43 31.0325 5.495 31.2825 ;
        RECT  5.43 32.1775 5.495 32.3125 ;
        RECT  5.07 32.2425 5.135 32.3125 ;
        RECT  5.07 31.0325 5.135 31.1475 ;
        RECT  5.26 31.1475 5.325 32.21 ;
        RECT  5.0025 31.685 5.0375 31.75 ;
        RECT  5.325 31.685 5.5625 31.75 ;
        RECT  5.07 32.0425 5.135 32.1775 ;
        RECT  5.26 32.0425 5.325 32.1775 ;
        RECT  5.07 31.4375 5.135 31.5725 ;
        RECT  5.26 31.4375 5.325 31.5725 ;
        RECT  5.43 31.2825 5.495 31.4175 ;
        RECT  5.43 32.2425 5.495 32.3775 ;
        RECT  5.0375 31.76 5.1725 31.825 ;
        RECT  5.0025 32.3125 5.5625 32.3775 ;
        RECT  5.0025 33.6575 5.5625 33.7225 ;
        RECT  5.43 33.4075 5.495 33.6575 ;
        RECT  5.43 32.3775 5.495 32.5125 ;
        RECT  5.07 32.3775 5.135 32.4475 ;
        RECT  5.07 33.5425 5.135 33.6575 ;
        RECT  5.26 32.48 5.325 33.5425 ;
        RECT  5.0025 32.94 5.0375 33.005 ;
        RECT  5.325 32.94 5.5625 33.005 ;
        RECT  5.07 32.5825 5.135 32.7175 ;
        RECT  5.26 32.5825 5.325 32.7175 ;
        RECT  5.07 33.4075 5.135 33.5425 ;
        RECT  5.26 33.4075 5.325 33.5425 ;
        RECT  5.43 33.4075 5.495 33.5425 ;
        RECT  5.43 32.4475 5.495 32.5825 ;
        RECT  5.0375 32.94 5.1725 33.005 ;
        RECT  5.0025 35.0025 5.5625 35.0675 ;
        RECT  5.0025 33.6575 5.5625 33.7225 ;
        RECT  5.43 33.7225 5.495 33.9725 ;
        RECT  5.43 34.8675 5.495 35.0025 ;
        RECT  5.07 34.9325 5.135 35.0025 ;
        RECT  5.07 33.7225 5.135 33.8375 ;
        RECT  5.26 33.8375 5.325 34.9 ;
        RECT  5.0025 34.375 5.0375 34.44 ;
        RECT  5.325 34.375 5.5625 34.44 ;
        RECT  5.07 34.7325 5.135 34.8675 ;
        RECT  5.26 34.7325 5.325 34.8675 ;
        RECT  5.07 34.1275 5.135 34.2625 ;
        RECT  5.26 34.1275 5.325 34.2625 ;
        RECT  5.43 33.9725 5.495 34.1075 ;
        RECT  5.43 34.9325 5.495 35.0675 ;
        RECT  5.0375 34.45 5.1725 34.515 ;
        RECT  5.0025 35.0025 5.5625 35.0675 ;
        RECT  5.0025 36.3475 5.5625 36.4125 ;
        RECT  5.43 36.0975 5.495 36.3475 ;
        RECT  5.43 35.0675 5.495 35.2025 ;
        RECT  5.07 35.0675 5.135 35.1375 ;
        RECT  5.07 36.2325 5.135 36.3475 ;
        RECT  5.26 35.17 5.325 36.2325 ;
        RECT  5.0025 35.63 5.0375 35.695 ;
        RECT  5.325 35.63 5.5625 35.695 ;
        RECT  5.07 35.2725 5.135 35.4075 ;
        RECT  5.26 35.2725 5.325 35.4075 ;
        RECT  5.07 36.0975 5.135 36.2325 ;
        RECT  5.26 36.0975 5.325 36.2325 ;
        RECT  5.43 36.0975 5.495 36.2325 ;
        RECT  5.43 35.1375 5.495 35.2725 ;
        RECT  5.0375 35.63 5.1725 35.695 ;
        RECT  5.0025 37.6925 5.5625 37.7575 ;
        RECT  5.0025 36.3475 5.5625 36.4125 ;
        RECT  5.43 36.4125 5.495 36.6625 ;
        RECT  5.43 37.5575 5.495 37.6925 ;
        RECT  5.07 37.6225 5.135 37.6925 ;
        RECT  5.07 36.4125 5.135 36.5275 ;
        RECT  5.26 36.5275 5.325 37.59 ;
        RECT  5.0025 37.065 5.0375 37.13 ;
        RECT  5.325 37.065 5.5625 37.13 ;
        RECT  5.07 37.4225 5.135 37.5575 ;
        RECT  5.26 37.4225 5.325 37.5575 ;
        RECT  5.07 36.8175 5.135 36.9525 ;
        RECT  5.26 36.8175 5.325 36.9525 ;
        RECT  5.43 36.6625 5.495 36.7975 ;
        RECT  5.43 37.6225 5.495 37.7575 ;
        RECT  5.0375 37.14 5.1725 37.205 ;
        RECT  5.0025 37.6925 5.5625 37.7575 ;
        RECT  5.0025 39.0375 5.5625 39.1025 ;
        RECT  5.43 38.7875 5.495 39.0375 ;
        RECT  5.43 37.7575 5.495 37.8925 ;
        RECT  5.07 37.7575 5.135 37.8275 ;
        RECT  5.07 38.9225 5.135 39.0375 ;
        RECT  5.26 37.86 5.325 38.9225 ;
        RECT  5.0025 38.32 5.0375 38.385 ;
        RECT  5.325 38.32 5.5625 38.385 ;
        RECT  5.07 37.9625 5.135 38.0975 ;
        RECT  5.26 37.9625 5.325 38.0975 ;
        RECT  5.07 38.7875 5.135 38.9225 ;
        RECT  5.26 38.7875 5.325 38.9225 ;
        RECT  5.43 38.7875 5.495 38.9225 ;
        RECT  5.43 37.8275 5.495 37.9625 ;
        RECT  5.0375 38.32 5.1725 38.385 ;
        RECT  5.0025 40.3825 5.5625 40.4475 ;
        RECT  5.0025 39.0375 5.5625 39.1025 ;
        RECT  5.43 39.1025 5.495 39.3525 ;
        RECT  5.43 40.2475 5.495 40.3825 ;
        RECT  5.07 40.3125 5.135 40.3825 ;
        RECT  5.07 39.1025 5.135 39.2175 ;
        RECT  5.26 39.2175 5.325 40.28 ;
        RECT  5.0025 39.755 5.0375 39.82 ;
        RECT  5.325 39.755 5.5625 39.82 ;
        RECT  5.07 40.1125 5.135 40.2475 ;
        RECT  5.26 40.1125 5.325 40.2475 ;
        RECT  5.07 39.5075 5.135 39.6425 ;
        RECT  5.26 39.5075 5.325 39.6425 ;
        RECT  5.43 39.3525 5.495 39.4875 ;
        RECT  5.43 40.3125 5.495 40.4475 ;
        RECT  5.0375 39.83 5.1725 39.895 ;
        RECT  2.8225 8.73 2.9575 8.795 ;
        RECT  2.9975 10.165 3.1325 10.23 ;
        RECT  3.1725 11.42 3.3075 11.485 ;
        RECT  3.3475 12.855 3.4825 12.92 ;
        RECT  3.5225 14.11 3.6575 14.175 ;
        RECT  3.6975 15.545 3.8325 15.61 ;
        RECT  3.8725 16.8 4.0075 16.865 ;
        RECT  4.0475 18.235 4.1825 18.3 ;
        RECT  2.8225 19.805 2.9575 19.87 ;
        RECT  3.5225 19.275 3.6575 19.34 ;
        RECT  2.8225 20.61 2.9575 20.675 ;
        RECT  3.6975 21.14 3.8325 21.205 ;
        RECT  2.8225 22.495 2.9575 22.56 ;
        RECT  3.8725 21.965 4.0075 22.03 ;
        RECT  2.8225 23.3 2.9575 23.365 ;
        RECT  4.0475 23.83 4.1825 23.895 ;
        RECT  2.9975 25.185 3.1325 25.25 ;
        RECT  3.5225 24.655 3.6575 24.72 ;
        RECT  2.9975 25.99 3.1325 26.055 ;
        RECT  3.6975 26.52 3.8325 26.585 ;
        RECT  2.9975 27.875 3.1325 27.94 ;
        RECT  3.8725 27.345 4.0075 27.41 ;
        RECT  2.9975 28.68 3.1325 28.745 ;
        RECT  4.0475 29.21 4.1825 29.275 ;
        RECT  3.1725 30.565 3.3075 30.63 ;
        RECT  3.5225 30.035 3.6575 30.1 ;
        RECT  3.1725 31.37 3.3075 31.435 ;
        RECT  3.6975 31.9 3.8325 31.965 ;
        RECT  3.1725 33.255 3.3075 33.32 ;
        RECT  3.8725 32.725 4.0075 32.79 ;
        RECT  3.1725 34.06 3.3075 34.125 ;
        RECT  4.0475 34.59 4.1825 34.655 ;
        RECT  3.3475 35.945 3.4825 36.01 ;
        RECT  3.5225 35.415 3.6575 35.48 ;
        RECT  3.3475 36.75 3.4825 36.815 ;
        RECT  3.6975 37.28 3.8325 37.345 ;
        RECT  3.3475 38.635 3.4825 38.7 ;
        RECT  3.8725 38.105 4.0075 38.17 ;
        RECT  3.3475 39.44 3.4825 39.505 ;
        RECT  4.0475 39.97 4.1825 40.035 ;
        RECT  5.7575 19.025 5.8225 40.805 ;
        RECT  5.7575 19.445 6.0825 19.51 ;
        RECT  6.5125 19.275 6.5775 19.51 ;
        RECT  7.3275 19.4925 7.3925 19.5575 ;
        RECT  7.8875 19.445 7.9525 19.51 ;
        RECT  5.7575 20.97 6.0825 21.035 ;
        RECT  6.5125 20.97 6.5775 21.205 ;
        RECT  7.3275 20.9225 7.3925 20.9875 ;
        RECT  7.8225 20.97 7.8875 21.035 ;
        RECT  5.7575 22.135 6.0825 22.2 ;
        RECT  6.5125 21.965 6.5775 22.2 ;
        RECT  7.3275 22.1825 7.3925 22.2475 ;
        RECT  7.8875 22.135 7.9525 22.2 ;
        RECT  5.7575 23.66 6.0825 23.725 ;
        RECT  6.5125 23.66 6.5775 23.895 ;
        RECT  7.3275 23.6125 7.3925 23.6775 ;
        RECT  7.8225 23.66 7.8875 23.725 ;
        RECT  5.7575 24.825 6.0825 24.89 ;
        RECT  6.5125 24.655 6.5775 24.89 ;
        RECT  7.3275 24.8725 7.3925 24.9375 ;
        RECT  7.8875 24.825 7.9525 24.89 ;
        RECT  5.7575 26.35 6.0825 26.415 ;
        RECT  6.5125 26.35 6.5775 26.585 ;
        RECT  7.3275 26.3025 7.3925 26.3675 ;
        RECT  7.8225 26.35 7.8875 26.415 ;
        RECT  5.7575 27.515 6.0825 27.58 ;
        RECT  6.5125 27.345 6.5775 27.58 ;
        RECT  7.3275 27.5625 7.3925 27.6275 ;
        RECT  7.8875 27.515 7.9525 27.58 ;
        RECT  5.7575 29.04 6.0825 29.105 ;
        RECT  6.5125 29.04 6.5775 29.275 ;
        RECT  7.3275 28.9925 7.3925 29.0575 ;
        RECT  7.8225 29.04 7.8875 29.105 ;
        RECT  5.7575 30.205 6.0825 30.27 ;
        RECT  6.5125 30.035 6.5775 30.27 ;
        RECT  7.3275 30.2525 7.3925 30.3175 ;
        RECT  7.8875 30.205 7.9525 30.27 ;
        RECT  5.7575 31.73 6.0825 31.795 ;
        RECT  6.5125 31.73 6.5775 31.965 ;
        RECT  7.3275 31.6825 7.3925 31.7475 ;
        RECT  7.8225 31.73 7.8875 31.795 ;
        RECT  5.7575 32.895 6.0825 32.96 ;
        RECT  6.5125 32.725 6.5775 32.96 ;
        RECT  7.3275 32.9425 7.3925 33.0075 ;
        RECT  7.8875 32.895 7.9525 32.96 ;
        RECT  5.7575 34.42 6.0825 34.485 ;
        RECT  6.5125 34.42 6.5775 34.655 ;
        RECT  7.3275 34.3725 7.3925 34.4375 ;
        RECT  7.8225 34.42 7.8875 34.485 ;
        RECT  5.7575 35.585 6.0825 35.65 ;
        RECT  6.5125 35.415 6.5775 35.65 ;
        RECT  7.3275 35.6325 7.3925 35.6975 ;
        RECT  7.8875 35.585 7.9525 35.65 ;
        RECT  5.7575 37.11 6.0825 37.175 ;
        RECT  6.5125 37.11 6.5775 37.345 ;
        RECT  7.3275 37.0625 7.3925 37.1275 ;
        RECT  7.8225 37.11 7.8875 37.175 ;
        RECT  5.7575 38.275 6.0825 38.34 ;
        RECT  6.5125 38.105 6.5775 38.34 ;
        RECT  7.3275 38.3225 7.3925 38.3875 ;
        RECT  7.8875 38.275 7.9525 38.34 ;
        RECT  5.7575 39.8 6.0825 39.865 ;
        RECT  6.5125 39.8 6.5775 40.035 ;
        RECT  7.3275 39.7525 7.3925 39.8175 ;
        RECT  7.8225 39.8 7.8875 39.865 ;
        RECT  5.4925 20.2075 5.6275 20.2725 ;
        RECT  5.9475 20.2075 6.0825 20.2725 ;
        RECT  6.0175 18.8625 6.5775 18.9275 ;
        RECT  6.0175 20.2075 6.5775 20.2725 ;
        RECT  6.445 19.8425 6.51 20.2075 ;
        RECT  6.445 18.9275 6.51 19.0625 ;
        RECT  6.085 18.9275 6.15 18.9975 ;
        RECT  6.085 20.1175 6.15 20.2075 ;
        RECT  6.275 19.03 6.34 19.9775 ;
        RECT  6.0175 19.445 6.0525 19.51 ;
        RECT  6.34 19.445 6.5775 19.51 ;
        RECT  6.085 19.1325 6.15 19.2675 ;
        RECT  6.275 19.1325 6.34 19.2675 ;
        RECT  6.085 19.8425 6.15 20.1175 ;
        RECT  6.275 19.8425 6.34 20.1175 ;
        RECT  6.445 19.8425 6.51 20.1175 ;
        RECT  6.445 18.9975 6.51 19.1325 ;
        RECT  6.0525 19.445 6.1875 19.51 ;
        RECT  6.5775 18.8625 7.3275 18.9275 ;
        RECT  6.5775 20.2075 7.3275 20.2725 ;
        RECT  7.195 19.9575 7.26 20.24 ;
        RECT  7.195 18.895 7.26 19.075 ;
        RECT  6.645 19.9575 6.71 20.24 ;
        RECT  7.025 19.9575 7.09 20.24 ;
        RECT  6.645 18.895 6.71 19.1775 ;
        RECT  7.0575 19.79 7.1225 19.855 ;
        RECT  6.835 19.79 6.9 19.855 ;
        RECT  7.0575 19.0425 7.1225 19.8225 ;
        RECT  6.8675 19.79 7.09 19.855 ;
        RECT  6.835 19.8225 6.9 19.9575 ;
        RECT  6.5775 19.805 6.6125 19.87 ;
        RECT  6.5775 19.275 6.8525 19.34 ;
        RECT  7.09 19.4925 7.3275 19.5575 ;
        RECT  6.645 19.1775 6.71 19.3125 ;
        RECT  6.835 19.1775 6.9 19.3125 ;
        RECT  6.835 19.1775 6.9 19.3125 ;
        RECT  7.025 19.1775 7.09 19.3125 ;
        RECT  6.645 19.9575 6.71 20.0925 ;
        RECT  6.835 19.9575 6.9 20.0925 ;
        RECT  6.835 19.9575 6.9 20.0925 ;
        RECT  7.025 19.9575 7.09 20.0925 ;
        RECT  7.195 19.9575 7.26 20.0925 ;
        RECT  7.195 19.0425 7.26 19.1775 ;
        RECT  6.6125 19.805 6.7475 19.87 ;
        RECT  6.8525 19.275 6.9875 19.34 ;
        RECT  7.3275 18.8625 7.8875 18.9275 ;
        RECT  7.3275 20.2075 7.8875 20.2725 ;
        RECT  7.755 19.8425 7.82 20.2075 ;
        RECT  7.755 18.9275 7.82 19.0625 ;
        RECT  7.395 18.9275 7.46 18.9975 ;
        RECT  7.395 20.1175 7.46 20.2075 ;
        RECT  7.585 19.03 7.65 19.9775 ;
        RECT  7.3275 19.445 7.3625 19.51 ;
        RECT  7.65 19.445 7.8875 19.51 ;
        RECT  7.395 19.1325 7.46 19.2675 ;
        RECT  7.585 19.1325 7.65 19.2675 ;
        RECT  7.395 19.8425 7.46 20.1175 ;
        RECT  7.585 19.8425 7.65 20.1175 ;
        RECT  7.755 19.8425 7.82 20.1175 ;
        RECT  7.755 18.9975 7.82 19.1325 ;
        RECT  7.3625 19.445 7.4975 19.51 ;
        RECT  6.5775 19.8075 6.7125 19.8725 ;
        RECT  5.565 19.805 5.63 19.94 ;
        RECT  5.4925 21.5525 5.6275 21.6175 ;
        RECT  5.9475 21.5525 6.0825 21.6175 ;
        RECT  6.0175 21.5525 6.5775 21.6175 ;
        RECT  6.0175 20.2075 6.5775 20.2725 ;
        RECT  6.445 20.2725 6.51 20.6375 ;
        RECT  6.445 21.4175 6.51 21.5525 ;
        RECT  6.085 21.4825 6.15 21.5525 ;
        RECT  6.085 20.2725 6.15 20.3625 ;
        RECT  6.275 20.5025 6.34 21.45 ;
        RECT  6.0175 20.97 6.0525 21.035 ;
        RECT  6.34 20.97 6.5775 21.035 ;
        RECT  6.085 21.2825 6.15 21.4175 ;
        RECT  6.275 21.2825 6.34 21.4175 ;
        RECT  6.085 20.7425 6.15 21.0175 ;
        RECT  6.275 20.7425 6.34 21.0175 ;
        RECT  6.445 20.6375 6.51 20.9125 ;
        RECT  6.445 21.4825 6.51 21.6175 ;
        RECT  6.0525 21.045 6.1875 21.11 ;
        RECT  6.5775 21.5525 7.3275 21.6175 ;
        RECT  6.5775 20.2075 7.3275 20.2725 ;
        RECT  7.195 20.24 7.26 20.5225 ;
        RECT  7.195 21.405 7.26 21.585 ;
        RECT  6.645 20.24 6.71 20.5225 ;
        RECT  7.025 20.24 7.09 20.5225 ;
        RECT  6.645 21.3025 6.71 21.585 ;
        RECT  7.0575 20.625 7.1225 20.69 ;
        RECT  6.835 20.625 6.9 20.69 ;
        RECT  7.0575 20.6575 7.1225 21.4375 ;
        RECT  6.8675 20.625 7.09 20.69 ;
        RECT  6.835 20.5225 6.9 20.6575 ;
        RECT  6.5775 20.61 6.6125 20.675 ;
        RECT  6.5775 21.14 6.8525 21.205 ;
        RECT  7.09 20.9225 7.3275 20.9875 ;
        RECT  6.645 21.1475 6.71 21.2825 ;
        RECT  6.835 21.1475 6.9 21.2825 ;
        RECT  6.835 21.1475 6.9 21.2825 ;
        RECT  7.025 21.1475 7.09 21.2825 ;
        RECT  6.645 20.6775 6.71 20.8125 ;
        RECT  6.835 20.6775 6.9 20.8125 ;
        RECT  6.835 20.6775 6.9 20.8125 ;
        RECT  7.025 20.6775 7.09 20.8125 ;
        RECT  7.195 20.5225 7.26 20.6575 ;
        RECT  7.195 21.4375 7.26 21.5725 ;
        RECT  6.6125 20.685 6.7475 20.75 ;
        RECT  6.8525 21.215 6.9875 21.28 ;
        RECT  7.3275 21.5525 7.8875 21.6175 ;
        RECT  7.3275 20.2075 7.8875 20.2725 ;
        RECT  7.755 20.2725 7.82 20.6375 ;
        RECT  7.755 21.4175 7.82 21.5525 ;
        RECT  7.395 21.4825 7.46 21.5525 ;
        RECT  7.395 20.2725 7.46 20.3625 ;
        RECT  7.585 20.5025 7.65 21.45 ;
        RECT  7.3275 20.97 7.3625 21.035 ;
        RECT  7.65 20.97 7.8875 21.035 ;
        RECT  7.395 21.2825 7.46 21.4175 ;
        RECT  7.585 21.2825 7.65 21.4175 ;
        RECT  7.395 20.7425 7.46 21.0175 ;
        RECT  7.585 20.7425 7.65 21.0175 ;
        RECT  7.755 20.6375 7.82 20.9125 ;
        RECT  7.755 21.4825 7.82 21.6175 ;
        RECT  7.3625 21.045 7.4975 21.11 ;
        RECT  6.5775 20.6075 6.7125 20.6725 ;
        RECT  5.565 20.54 5.63 20.675 ;
        RECT  5.4925 22.8975 5.6275 22.9625 ;
        RECT  5.9475 22.8975 6.0825 22.9625 ;
        RECT  6.0175 21.5525 6.5775 21.6175 ;
        RECT  6.0175 22.8975 6.5775 22.9625 ;
        RECT  6.445 22.5325 6.51 22.8975 ;
        RECT  6.445 21.6175 6.51 21.7525 ;
        RECT  6.085 21.6175 6.15 21.6875 ;
        RECT  6.085 22.8075 6.15 22.8975 ;
        RECT  6.275 21.72 6.34 22.6675 ;
        RECT  6.0175 22.135 6.0525 22.2 ;
        RECT  6.34 22.135 6.5775 22.2 ;
        RECT  6.085 21.8225 6.15 21.9575 ;
        RECT  6.275 21.8225 6.34 21.9575 ;
        RECT  6.085 22.5325 6.15 22.8075 ;
        RECT  6.275 22.5325 6.34 22.8075 ;
        RECT  6.445 22.5325 6.51 22.8075 ;
        RECT  6.445 21.6875 6.51 21.8225 ;
        RECT  6.0525 22.135 6.1875 22.2 ;
        RECT  6.5775 21.5525 7.3275 21.6175 ;
        RECT  6.5775 22.8975 7.3275 22.9625 ;
        RECT  7.195 22.6475 7.26 22.93 ;
        RECT  7.195 21.585 7.26 21.765 ;
        RECT  6.645 22.6475 6.71 22.93 ;
        RECT  7.025 22.6475 7.09 22.93 ;
        RECT  6.645 21.585 6.71 21.8675 ;
        RECT  7.0575 22.48 7.1225 22.545 ;
        RECT  6.835 22.48 6.9 22.545 ;
        RECT  7.0575 21.7325 7.1225 22.5125 ;
        RECT  6.8675 22.48 7.09 22.545 ;
        RECT  6.835 22.5125 6.9 22.6475 ;
        RECT  6.5775 22.495 6.6125 22.56 ;
        RECT  6.5775 21.965 6.8525 22.03 ;
        RECT  7.09 22.1825 7.3275 22.2475 ;
        RECT  6.645 21.8675 6.71 22.0025 ;
        RECT  6.835 21.8675 6.9 22.0025 ;
        RECT  6.835 21.8675 6.9 22.0025 ;
        RECT  7.025 21.8675 7.09 22.0025 ;
        RECT  6.645 22.6475 6.71 22.7825 ;
        RECT  6.835 22.6475 6.9 22.7825 ;
        RECT  6.835 22.6475 6.9 22.7825 ;
        RECT  7.025 22.6475 7.09 22.7825 ;
        RECT  7.195 22.6475 7.26 22.7825 ;
        RECT  7.195 21.7325 7.26 21.8675 ;
        RECT  6.6125 22.495 6.7475 22.56 ;
        RECT  6.8525 21.965 6.9875 22.03 ;
        RECT  7.3275 21.5525 7.8875 21.6175 ;
        RECT  7.3275 22.8975 7.8875 22.9625 ;
        RECT  7.755 22.5325 7.82 22.8975 ;
        RECT  7.755 21.6175 7.82 21.7525 ;
        RECT  7.395 21.6175 7.46 21.6875 ;
        RECT  7.395 22.8075 7.46 22.8975 ;
        RECT  7.585 21.72 7.65 22.6675 ;
        RECT  7.3275 22.135 7.3625 22.2 ;
        RECT  7.65 22.135 7.8875 22.2 ;
        RECT  7.395 21.8225 7.46 21.9575 ;
        RECT  7.585 21.8225 7.65 21.9575 ;
        RECT  7.395 22.5325 7.46 22.8075 ;
        RECT  7.585 22.5325 7.65 22.8075 ;
        RECT  7.755 22.5325 7.82 22.8075 ;
        RECT  7.755 21.6875 7.82 21.8225 ;
        RECT  7.3625 22.135 7.4975 22.2 ;
        RECT  6.5775 22.4975 6.7125 22.5625 ;
        RECT  5.565 22.495 5.63 22.63 ;
        RECT  5.4925 24.2425 5.6275 24.3075 ;
        RECT  5.9475 24.2425 6.0825 24.3075 ;
        RECT  6.0175 24.2425 6.5775 24.3075 ;
        RECT  6.0175 22.8975 6.5775 22.9625 ;
        RECT  6.445 22.9625 6.51 23.3275 ;
        RECT  6.445 24.1075 6.51 24.2425 ;
        RECT  6.085 24.1725 6.15 24.2425 ;
        RECT  6.085 22.9625 6.15 23.0525 ;
        RECT  6.275 23.1925 6.34 24.14 ;
        RECT  6.0175 23.66 6.0525 23.725 ;
        RECT  6.34 23.66 6.5775 23.725 ;
        RECT  6.085 23.9725 6.15 24.1075 ;
        RECT  6.275 23.9725 6.34 24.1075 ;
        RECT  6.085 23.4325 6.15 23.7075 ;
        RECT  6.275 23.4325 6.34 23.7075 ;
        RECT  6.445 23.3275 6.51 23.6025 ;
        RECT  6.445 24.1725 6.51 24.3075 ;
        RECT  6.0525 23.735 6.1875 23.8 ;
        RECT  6.5775 24.2425 7.3275 24.3075 ;
        RECT  6.5775 22.8975 7.3275 22.9625 ;
        RECT  7.195 22.93 7.26 23.2125 ;
        RECT  7.195 24.095 7.26 24.275 ;
        RECT  6.645 22.93 6.71 23.2125 ;
        RECT  7.025 22.93 7.09 23.2125 ;
        RECT  6.645 23.9925 6.71 24.275 ;
        RECT  7.0575 23.315 7.1225 23.38 ;
        RECT  6.835 23.315 6.9 23.38 ;
        RECT  7.0575 23.3475 7.1225 24.1275 ;
        RECT  6.8675 23.315 7.09 23.38 ;
        RECT  6.835 23.2125 6.9 23.3475 ;
        RECT  6.5775 23.3 6.6125 23.365 ;
        RECT  6.5775 23.83 6.8525 23.895 ;
        RECT  7.09 23.6125 7.3275 23.6775 ;
        RECT  6.645 23.8375 6.71 23.9725 ;
        RECT  6.835 23.8375 6.9 23.9725 ;
        RECT  6.835 23.8375 6.9 23.9725 ;
        RECT  7.025 23.8375 7.09 23.9725 ;
        RECT  6.645 23.3675 6.71 23.5025 ;
        RECT  6.835 23.3675 6.9 23.5025 ;
        RECT  6.835 23.3675 6.9 23.5025 ;
        RECT  7.025 23.3675 7.09 23.5025 ;
        RECT  7.195 23.2125 7.26 23.3475 ;
        RECT  7.195 24.1275 7.26 24.2625 ;
        RECT  6.6125 23.375 6.7475 23.44 ;
        RECT  6.8525 23.905 6.9875 23.97 ;
        RECT  7.3275 24.2425 7.8875 24.3075 ;
        RECT  7.3275 22.8975 7.8875 22.9625 ;
        RECT  7.755 22.9625 7.82 23.3275 ;
        RECT  7.755 24.1075 7.82 24.2425 ;
        RECT  7.395 24.1725 7.46 24.2425 ;
        RECT  7.395 22.9625 7.46 23.0525 ;
        RECT  7.585 23.1925 7.65 24.14 ;
        RECT  7.3275 23.66 7.3625 23.725 ;
        RECT  7.65 23.66 7.8875 23.725 ;
        RECT  7.395 23.9725 7.46 24.1075 ;
        RECT  7.585 23.9725 7.65 24.1075 ;
        RECT  7.395 23.4325 7.46 23.7075 ;
        RECT  7.585 23.4325 7.65 23.7075 ;
        RECT  7.755 23.3275 7.82 23.6025 ;
        RECT  7.755 24.1725 7.82 24.3075 ;
        RECT  7.3625 23.735 7.4975 23.8 ;
        RECT  6.5775 23.2975 6.7125 23.3625 ;
        RECT  5.565 23.23 5.63 23.365 ;
        RECT  5.4925 25.5875 5.6275 25.6525 ;
        RECT  5.9475 25.5875 6.0825 25.6525 ;
        RECT  6.0175 24.2425 6.5775 24.3075 ;
        RECT  6.0175 25.5875 6.5775 25.6525 ;
        RECT  6.445 25.2225 6.51 25.5875 ;
        RECT  6.445 24.3075 6.51 24.4425 ;
        RECT  6.085 24.3075 6.15 24.3775 ;
        RECT  6.085 25.4975 6.15 25.5875 ;
        RECT  6.275 24.41 6.34 25.3575 ;
        RECT  6.0175 24.825 6.0525 24.89 ;
        RECT  6.34 24.825 6.5775 24.89 ;
        RECT  6.085 24.5125 6.15 24.6475 ;
        RECT  6.275 24.5125 6.34 24.6475 ;
        RECT  6.085 25.2225 6.15 25.4975 ;
        RECT  6.275 25.2225 6.34 25.4975 ;
        RECT  6.445 25.2225 6.51 25.4975 ;
        RECT  6.445 24.3775 6.51 24.5125 ;
        RECT  6.0525 24.825 6.1875 24.89 ;
        RECT  6.5775 24.2425 7.3275 24.3075 ;
        RECT  6.5775 25.5875 7.3275 25.6525 ;
        RECT  7.195 25.3375 7.26 25.62 ;
        RECT  7.195 24.275 7.26 24.455 ;
        RECT  6.645 25.3375 6.71 25.62 ;
        RECT  7.025 25.3375 7.09 25.62 ;
        RECT  6.645 24.275 6.71 24.5575 ;
        RECT  7.0575 25.17 7.1225 25.235 ;
        RECT  6.835 25.17 6.9 25.235 ;
        RECT  7.0575 24.4225 7.1225 25.2025 ;
        RECT  6.8675 25.17 7.09 25.235 ;
        RECT  6.835 25.2025 6.9 25.3375 ;
        RECT  6.5775 25.185 6.6125 25.25 ;
        RECT  6.5775 24.655 6.8525 24.72 ;
        RECT  7.09 24.8725 7.3275 24.9375 ;
        RECT  6.645 24.5575 6.71 24.6925 ;
        RECT  6.835 24.5575 6.9 24.6925 ;
        RECT  6.835 24.5575 6.9 24.6925 ;
        RECT  7.025 24.5575 7.09 24.6925 ;
        RECT  6.645 25.3375 6.71 25.4725 ;
        RECT  6.835 25.3375 6.9 25.4725 ;
        RECT  6.835 25.3375 6.9 25.4725 ;
        RECT  7.025 25.3375 7.09 25.4725 ;
        RECT  7.195 25.3375 7.26 25.4725 ;
        RECT  7.195 24.4225 7.26 24.5575 ;
        RECT  6.6125 25.185 6.7475 25.25 ;
        RECT  6.8525 24.655 6.9875 24.72 ;
        RECT  7.3275 24.2425 7.8875 24.3075 ;
        RECT  7.3275 25.5875 7.8875 25.6525 ;
        RECT  7.755 25.2225 7.82 25.5875 ;
        RECT  7.755 24.3075 7.82 24.4425 ;
        RECT  7.395 24.3075 7.46 24.3775 ;
        RECT  7.395 25.4975 7.46 25.5875 ;
        RECT  7.585 24.41 7.65 25.3575 ;
        RECT  7.3275 24.825 7.3625 24.89 ;
        RECT  7.65 24.825 7.8875 24.89 ;
        RECT  7.395 24.5125 7.46 24.6475 ;
        RECT  7.585 24.5125 7.65 24.6475 ;
        RECT  7.395 25.2225 7.46 25.4975 ;
        RECT  7.585 25.2225 7.65 25.4975 ;
        RECT  7.755 25.2225 7.82 25.4975 ;
        RECT  7.755 24.3775 7.82 24.5125 ;
        RECT  7.3625 24.825 7.4975 24.89 ;
        RECT  6.5775 25.1875 6.7125 25.2525 ;
        RECT  5.565 25.185 5.63 25.32 ;
        RECT  5.4925 26.9325 5.6275 26.9975 ;
        RECT  5.9475 26.9325 6.0825 26.9975 ;
        RECT  6.0175 26.9325 6.5775 26.9975 ;
        RECT  6.0175 25.5875 6.5775 25.6525 ;
        RECT  6.445 25.6525 6.51 26.0175 ;
        RECT  6.445 26.7975 6.51 26.9325 ;
        RECT  6.085 26.8625 6.15 26.9325 ;
        RECT  6.085 25.6525 6.15 25.7425 ;
        RECT  6.275 25.8825 6.34 26.83 ;
        RECT  6.0175 26.35 6.0525 26.415 ;
        RECT  6.34 26.35 6.5775 26.415 ;
        RECT  6.085 26.6625 6.15 26.7975 ;
        RECT  6.275 26.6625 6.34 26.7975 ;
        RECT  6.085 26.1225 6.15 26.3975 ;
        RECT  6.275 26.1225 6.34 26.3975 ;
        RECT  6.445 26.0175 6.51 26.2925 ;
        RECT  6.445 26.8625 6.51 26.9975 ;
        RECT  6.0525 26.425 6.1875 26.49 ;
        RECT  6.5775 26.9325 7.3275 26.9975 ;
        RECT  6.5775 25.5875 7.3275 25.6525 ;
        RECT  7.195 25.62 7.26 25.9025 ;
        RECT  7.195 26.785 7.26 26.965 ;
        RECT  6.645 25.62 6.71 25.9025 ;
        RECT  7.025 25.62 7.09 25.9025 ;
        RECT  6.645 26.6825 6.71 26.965 ;
        RECT  7.0575 26.005 7.1225 26.07 ;
        RECT  6.835 26.005 6.9 26.07 ;
        RECT  7.0575 26.0375 7.1225 26.8175 ;
        RECT  6.8675 26.005 7.09 26.07 ;
        RECT  6.835 25.9025 6.9 26.0375 ;
        RECT  6.5775 25.99 6.6125 26.055 ;
        RECT  6.5775 26.52 6.8525 26.585 ;
        RECT  7.09 26.3025 7.3275 26.3675 ;
        RECT  6.645 26.5275 6.71 26.6625 ;
        RECT  6.835 26.5275 6.9 26.6625 ;
        RECT  6.835 26.5275 6.9 26.6625 ;
        RECT  7.025 26.5275 7.09 26.6625 ;
        RECT  6.645 26.0575 6.71 26.1925 ;
        RECT  6.835 26.0575 6.9 26.1925 ;
        RECT  6.835 26.0575 6.9 26.1925 ;
        RECT  7.025 26.0575 7.09 26.1925 ;
        RECT  7.195 25.9025 7.26 26.0375 ;
        RECT  7.195 26.8175 7.26 26.9525 ;
        RECT  6.6125 26.065 6.7475 26.13 ;
        RECT  6.8525 26.595 6.9875 26.66 ;
        RECT  7.3275 26.9325 7.8875 26.9975 ;
        RECT  7.3275 25.5875 7.8875 25.6525 ;
        RECT  7.755 25.6525 7.82 26.0175 ;
        RECT  7.755 26.7975 7.82 26.9325 ;
        RECT  7.395 26.8625 7.46 26.9325 ;
        RECT  7.395 25.6525 7.46 25.7425 ;
        RECT  7.585 25.8825 7.65 26.83 ;
        RECT  7.3275 26.35 7.3625 26.415 ;
        RECT  7.65 26.35 7.8875 26.415 ;
        RECT  7.395 26.6625 7.46 26.7975 ;
        RECT  7.585 26.6625 7.65 26.7975 ;
        RECT  7.395 26.1225 7.46 26.3975 ;
        RECT  7.585 26.1225 7.65 26.3975 ;
        RECT  7.755 26.0175 7.82 26.2925 ;
        RECT  7.755 26.8625 7.82 26.9975 ;
        RECT  7.3625 26.425 7.4975 26.49 ;
        RECT  6.5775 25.9875 6.7125 26.0525 ;
        RECT  5.565 25.92 5.63 26.055 ;
        RECT  5.4925 28.2775 5.6275 28.3425 ;
        RECT  5.9475 28.2775 6.0825 28.3425 ;
        RECT  6.0175 26.9325 6.5775 26.9975 ;
        RECT  6.0175 28.2775 6.5775 28.3425 ;
        RECT  6.445 27.9125 6.51 28.2775 ;
        RECT  6.445 26.9975 6.51 27.1325 ;
        RECT  6.085 26.9975 6.15 27.0675 ;
        RECT  6.085 28.1875 6.15 28.2775 ;
        RECT  6.275 27.1 6.34 28.0475 ;
        RECT  6.0175 27.515 6.0525 27.58 ;
        RECT  6.34 27.515 6.5775 27.58 ;
        RECT  6.085 27.2025 6.15 27.3375 ;
        RECT  6.275 27.2025 6.34 27.3375 ;
        RECT  6.085 27.9125 6.15 28.1875 ;
        RECT  6.275 27.9125 6.34 28.1875 ;
        RECT  6.445 27.9125 6.51 28.1875 ;
        RECT  6.445 27.0675 6.51 27.2025 ;
        RECT  6.0525 27.515 6.1875 27.58 ;
        RECT  6.5775 26.9325 7.3275 26.9975 ;
        RECT  6.5775 28.2775 7.3275 28.3425 ;
        RECT  7.195 28.0275 7.26 28.31 ;
        RECT  7.195 26.965 7.26 27.145 ;
        RECT  6.645 28.0275 6.71 28.31 ;
        RECT  7.025 28.0275 7.09 28.31 ;
        RECT  6.645 26.965 6.71 27.2475 ;
        RECT  7.0575 27.86 7.1225 27.925 ;
        RECT  6.835 27.86 6.9 27.925 ;
        RECT  7.0575 27.1125 7.1225 27.8925 ;
        RECT  6.8675 27.86 7.09 27.925 ;
        RECT  6.835 27.8925 6.9 28.0275 ;
        RECT  6.5775 27.875 6.6125 27.94 ;
        RECT  6.5775 27.345 6.8525 27.41 ;
        RECT  7.09 27.5625 7.3275 27.6275 ;
        RECT  6.645 27.2475 6.71 27.3825 ;
        RECT  6.835 27.2475 6.9 27.3825 ;
        RECT  6.835 27.2475 6.9 27.3825 ;
        RECT  7.025 27.2475 7.09 27.3825 ;
        RECT  6.645 28.0275 6.71 28.1625 ;
        RECT  6.835 28.0275 6.9 28.1625 ;
        RECT  6.835 28.0275 6.9 28.1625 ;
        RECT  7.025 28.0275 7.09 28.1625 ;
        RECT  7.195 28.0275 7.26 28.1625 ;
        RECT  7.195 27.1125 7.26 27.2475 ;
        RECT  6.6125 27.875 6.7475 27.94 ;
        RECT  6.8525 27.345 6.9875 27.41 ;
        RECT  7.3275 26.9325 7.8875 26.9975 ;
        RECT  7.3275 28.2775 7.8875 28.3425 ;
        RECT  7.755 27.9125 7.82 28.2775 ;
        RECT  7.755 26.9975 7.82 27.1325 ;
        RECT  7.395 26.9975 7.46 27.0675 ;
        RECT  7.395 28.1875 7.46 28.2775 ;
        RECT  7.585 27.1 7.65 28.0475 ;
        RECT  7.3275 27.515 7.3625 27.58 ;
        RECT  7.65 27.515 7.8875 27.58 ;
        RECT  7.395 27.2025 7.46 27.3375 ;
        RECT  7.585 27.2025 7.65 27.3375 ;
        RECT  7.395 27.9125 7.46 28.1875 ;
        RECT  7.585 27.9125 7.65 28.1875 ;
        RECT  7.755 27.9125 7.82 28.1875 ;
        RECT  7.755 27.0675 7.82 27.2025 ;
        RECT  7.3625 27.515 7.4975 27.58 ;
        RECT  6.5775 27.8775 6.7125 27.9425 ;
        RECT  5.565 27.875 5.63 28.01 ;
        RECT  5.4925 29.6225 5.6275 29.6875 ;
        RECT  5.9475 29.6225 6.0825 29.6875 ;
        RECT  6.0175 29.6225 6.5775 29.6875 ;
        RECT  6.0175 28.2775 6.5775 28.3425 ;
        RECT  6.445 28.3425 6.51 28.7075 ;
        RECT  6.445 29.4875 6.51 29.6225 ;
        RECT  6.085 29.5525 6.15 29.6225 ;
        RECT  6.085 28.3425 6.15 28.4325 ;
        RECT  6.275 28.5725 6.34 29.52 ;
        RECT  6.0175 29.04 6.0525 29.105 ;
        RECT  6.34 29.04 6.5775 29.105 ;
        RECT  6.085 29.3525 6.15 29.4875 ;
        RECT  6.275 29.3525 6.34 29.4875 ;
        RECT  6.085 28.8125 6.15 29.0875 ;
        RECT  6.275 28.8125 6.34 29.0875 ;
        RECT  6.445 28.7075 6.51 28.9825 ;
        RECT  6.445 29.5525 6.51 29.6875 ;
        RECT  6.0525 29.115 6.1875 29.18 ;
        RECT  6.5775 29.6225 7.3275 29.6875 ;
        RECT  6.5775 28.2775 7.3275 28.3425 ;
        RECT  7.195 28.31 7.26 28.5925 ;
        RECT  7.195 29.475 7.26 29.655 ;
        RECT  6.645 28.31 6.71 28.5925 ;
        RECT  7.025 28.31 7.09 28.5925 ;
        RECT  6.645 29.3725 6.71 29.655 ;
        RECT  7.0575 28.695 7.1225 28.76 ;
        RECT  6.835 28.695 6.9 28.76 ;
        RECT  7.0575 28.7275 7.1225 29.5075 ;
        RECT  6.8675 28.695 7.09 28.76 ;
        RECT  6.835 28.5925 6.9 28.7275 ;
        RECT  6.5775 28.68 6.6125 28.745 ;
        RECT  6.5775 29.21 6.8525 29.275 ;
        RECT  7.09 28.9925 7.3275 29.0575 ;
        RECT  6.645 29.2175 6.71 29.3525 ;
        RECT  6.835 29.2175 6.9 29.3525 ;
        RECT  6.835 29.2175 6.9 29.3525 ;
        RECT  7.025 29.2175 7.09 29.3525 ;
        RECT  6.645 28.7475 6.71 28.8825 ;
        RECT  6.835 28.7475 6.9 28.8825 ;
        RECT  6.835 28.7475 6.9 28.8825 ;
        RECT  7.025 28.7475 7.09 28.8825 ;
        RECT  7.195 28.5925 7.26 28.7275 ;
        RECT  7.195 29.5075 7.26 29.6425 ;
        RECT  6.6125 28.755 6.7475 28.82 ;
        RECT  6.8525 29.285 6.9875 29.35 ;
        RECT  7.3275 29.6225 7.8875 29.6875 ;
        RECT  7.3275 28.2775 7.8875 28.3425 ;
        RECT  7.755 28.3425 7.82 28.7075 ;
        RECT  7.755 29.4875 7.82 29.6225 ;
        RECT  7.395 29.5525 7.46 29.6225 ;
        RECT  7.395 28.3425 7.46 28.4325 ;
        RECT  7.585 28.5725 7.65 29.52 ;
        RECT  7.3275 29.04 7.3625 29.105 ;
        RECT  7.65 29.04 7.8875 29.105 ;
        RECT  7.395 29.3525 7.46 29.4875 ;
        RECT  7.585 29.3525 7.65 29.4875 ;
        RECT  7.395 28.8125 7.46 29.0875 ;
        RECT  7.585 28.8125 7.65 29.0875 ;
        RECT  7.755 28.7075 7.82 28.9825 ;
        RECT  7.755 29.5525 7.82 29.6875 ;
        RECT  7.3625 29.115 7.4975 29.18 ;
        RECT  6.5775 28.6775 6.7125 28.7425 ;
        RECT  5.565 28.61 5.63 28.745 ;
        RECT  5.4925 30.9675 5.6275 31.0325 ;
        RECT  5.9475 30.9675 6.0825 31.0325 ;
        RECT  6.0175 29.6225 6.5775 29.6875 ;
        RECT  6.0175 30.9675 6.5775 31.0325 ;
        RECT  6.445 30.6025 6.51 30.9675 ;
        RECT  6.445 29.6875 6.51 29.8225 ;
        RECT  6.085 29.6875 6.15 29.7575 ;
        RECT  6.085 30.8775 6.15 30.9675 ;
        RECT  6.275 29.79 6.34 30.7375 ;
        RECT  6.0175 30.205 6.0525 30.27 ;
        RECT  6.34 30.205 6.5775 30.27 ;
        RECT  6.085 29.8925 6.15 30.0275 ;
        RECT  6.275 29.8925 6.34 30.0275 ;
        RECT  6.085 30.6025 6.15 30.8775 ;
        RECT  6.275 30.6025 6.34 30.8775 ;
        RECT  6.445 30.6025 6.51 30.8775 ;
        RECT  6.445 29.7575 6.51 29.8925 ;
        RECT  6.0525 30.205 6.1875 30.27 ;
        RECT  6.5775 29.6225 7.3275 29.6875 ;
        RECT  6.5775 30.9675 7.3275 31.0325 ;
        RECT  7.195 30.7175 7.26 31.0 ;
        RECT  7.195 29.655 7.26 29.835 ;
        RECT  6.645 30.7175 6.71 31.0 ;
        RECT  7.025 30.7175 7.09 31.0 ;
        RECT  6.645 29.655 6.71 29.9375 ;
        RECT  7.0575 30.55 7.1225 30.615 ;
        RECT  6.835 30.55 6.9 30.615 ;
        RECT  7.0575 29.8025 7.1225 30.5825 ;
        RECT  6.8675 30.55 7.09 30.615 ;
        RECT  6.835 30.5825 6.9 30.7175 ;
        RECT  6.5775 30.565 6.6125 30.63 ;
        RECT  6.5775 30.035 6.8525 30.1 ;
        RECT  7.09 30.2525 7.3275 30.3175 ;
        RECT  6.645 29.9375 6.71 30.0725 ;
        RECT  6.835 29.9375 6.9 30.0725 ;
        RECT  6.835 29.9375 6.9 30.0725 ;
        RECT  7.025 29.9375 7.09 30.0725 ;
        RECT  6.645 30.7175 6.71 30.8525 ;
        RECT  6.835 30.7175 6.9 30.8525 ;
        RECT  6.835 30.7175 6.9 30.8525 ;
        RECT  7.025 30.7175 7.09 30.8525 ;
        RECT  7.195 30.7175 7.26 30.8525 ;
        RECT  7.195 29.8025 7.26 29.9375 ;
        RECT  6.6125 30.565 6.7475 30.63 ;
        RECT  6.8525 30.035 6.9875 30.1 ;
        RECT  7.3275 29.6225 7.8875 29.6875 ;
        RECT  7.3275 30.9675 7.8875 31.0325 ;
        RECT  7.755 30.6025 7.82 30.9675 ;
        RECT  7.755 29.6875 7.82 29.8225 ;
        RECT  7.395 29.6875 7.46 29.7575 ;
        RECT  7.395 30.8775 7.46 30.9675 ;
        RECT  7.585 29.79 7.65 30.7375 ;
        RECT  7.3275 30.205 7.3625 30.27 ;
        RECT  7.65 30.205 7.8875 30.27 ;
        RECT  7.395 29.8925 7.46 30.0275 ;
        RECT  7.585 29.8925 7.65 30.0275 ;
        RECT  7.395 30.6025 7.46 30.8775 ;
        RECT  7.585 30.6025 7.65 30.8775 ;
        RECT  7.755 30.6025 7.82 30.8775 ;
        RECT  7.755 29.7575 7.82 29.8925 ;
        RECT  7.3625 30.205 7.4975 30.27 ;
        RECT  6.5775 30.5675 6.7125 30.6325 ;
        RECT  5.565 30.565 5.63 30.7 ;
        RECT  5.4925 32.3125 5.6275 32.3775 ;
        RECT  5.9475 32.3125 6.0825 32.3775 ;
        RECT  6.0175 32.3125 6.5775 32.3775 ;
        RECT  6.0175 30.9675 6.5775 31.0325 ;
        RECT  6.445 31.0325 6.51 31.3975 ;
        RECT  6.445 32.1775 6.51 32.3125 ;
        RECT  6.085 32.2425 6.15 32.3125 ;
        RECT  6.085 31.0325 6.15 31.1225 ;
        RECT  6.275 31.2625 6.34 32.21 ;
        RECT  6.0175 31.73 6.0525 31.795 ;
        RECT  6.34 31.73 6.5775 31.795 ;
        RECT  6.085 32.0425 6.15 32.1775 ;
        RECT  6.275 32.0425 6.34 32.1775 ;
        RECT  6.085 31.5025 6.15 31.7775 ;
        RECT  6.275 31.5025 6.34 31.7775 ;
        RECT  6.445 31.3975 6.51 31.6725 ;
        RECT  6.445 32.2425 6.51 32.3775 ;
        RECT  6.0525 31.805 6.1875 31.87 ;
        RECT  6.5775 32.3125 7.3275 32.3775 ;
        RECT  6.5775 30.9675 7.3275 31.0325 ;
        RECT  7.195 31.0 7.26 31.2825 ;
        RECT  7.195 32.165 7.26 32.345 ;
        RECT  6.645 31.0 6.71 31.2825 ;
        RECT  7.025 31.0 7.09 31.2825 ;
        RECT  6.645 32.0625 6.71 32.345 ;
        RECT  7.0575 31.385 7.1225 31.45 ;
        RECT  6.835 31.385 6.9 31.45 ;
        RECT  7.0575 31.4175 7.1225 32.1975 ;
        RECT  6.8675 31.385 7.09 31.45 ;
        RECT  6.835 31.2825 6.9 31.4175 ;
        RECT  6.5775 31.37 6.6125 31.435 ;
        RECT  6.5775 31.9 6.8525 31.965 ;
        RECT  7.09 31.6825 7.3275 31.7475 ;
        RECT  6.645 31.9075 6.71 32.0425 ;
        RECT  6.835 31.9075 6.9 32.0425 ;
        RECT  6.835 31.9075 6.9 32.0425 ;
        RECT  7.025 31.9075 7.09 32.0425 ;
        RECT  6.645 31.4375 6.71 31.5725 ;
        RECT  6.835 31.4375 6.9 31.5725 ;
        RECT  6.835 31.4375 6.9 31.5725 ;
        RECT  7.025 31.4375 7.09 31.5725 ;
        RECT  7.195 31.2825 7.26 31.4175 ;
        RECT  7.195 32.1975 7.26 32.3325 ;
        RECT  6.6125 31.445 6.7475 31.51 ;
        RECT  6.8525 31.975 6.9875 32.04 ;
        RECT  7.3275 32.3125 7.8875 32.3775 ;
        RECT  7.3275 30.9675 7.8875 31.0325 ;
        RECT  7.755 31.0325 7.82 31.3975 ;
        RECT  7.755 32.1775 7.82 32.3125 ;
        RECT  7.395 32.2425 7.46 32.3125 ;
        RECT  7.395 31.0325 7.46 31.1225 ;
        RECT  7.585 31.2625 7.65 32.21 ;
        RECT  7.3275 31.73 7.3625 31.795 ;
        RECT  7.65 31.73 7.8875 31.795 ;
        RECT  7.395 32.0425 7.46 32.1775 ;
        RECT  7.585 32.0425 7.65 32.1775 ;
        RECT  7.395 31.5025 7.46 31.7775 ;
        RECT  7.585 31.5025 7.65 31.7775 ;
        RECT  7.755 31.3975 7.82 31.6725 ;
        RECT  7.755 32.2425 7.82 32.3775 ;
        RECT  7.3625 31.805 7.4975 31.87 ;
        RECT  6.5775 31.3675 6.7125 31.4325 ;
        RECT  5.565 31.3 5.63 31.435 ;
        RECT  5.4925 33.6575 5.6275 33.7225 ;
        RECT  5.9475 33.6575 6.0825 33.7225 ;
        RECT  6.0175 32.3125 6.5775 32.3775 ;
        RECT  6.0175 33.6575 6.5775 33.7225 ;
        RECT  6.445 33.2925 6.51 33.6575 ;
        RECT  6.445 32.3775 6.51 32.5125 ;
        RECT  6.085 32.3775 6.15 32.4475 ;
        RECT  6.085 33.5675 6.15 33.6575 ;
        RECT  6.275 32.48 6.34 33.4275 ;
        RECT  6.0175 32.895 6.0525 32.96 ;
        RECT  6.34 32.895 6.5775 32.96 ;
        RECT  6.085 32.5825 6.15 32.7175 ;
        RECT  6.275 32.5825 6.34 32.7175 ;
        RECT  6.085 33.2925 6.15 33.5675 ;
        RECT  6.275 33.2925 6.34 33.5675 ;
        RECT  6.445 33.2925 6.51 33.5675 ;
        RECT  6.445 32.4475 6.51 32.5825 ;
        RECT  6.0525 32.895 6.1875 32.96 ;
        RECT  6.5775 32.3125 7.3275 32.3775 ;
        RECT  6.5775 33.6575 7.3275 33.7225 ;
        RECT  7.195 33.4075 7.26 33.69 ;
        RECT  7.195 32.345 7.26 32.525 ;
        RECT  6.645 33.4075 6.71 33.69 ;
        RECT  7.025 33.4075 7.09 33.69 ;
        RECT  6.645 32.345 6.71 32.6275 ;
        RECT  7.0575 33.24 7.1225 33.305 ;
        RECT  6.835 33.24 6.9 33.305 ;
        RECT  7.0575 32.4925 7.1225 33.2725 ;
        RECT  6.8675 33.24 7.09 33.305 ;
        RECT  6.835 33.2725 6.9 33.4075 ;
        RECT  6.5775 33.255 6.6125 33.32 ;
        RECT  6.5775 32.725 6.8525 32.79 ;
        RECT  7.09 32.9425 7.3275 33.0075 ;
        RECT  6.645 32.6275 6.71 32.7625 ;
        RECT  6.835 32.6275 6.9 32.7625 ;
        RECT  6.835 32.6275 6.9 32.7625 ;
        RECT  7.025 32.6275 7.09 32.7625 ;
        RECT  6.645 33.4075 6.71 33.5425 ;
        RECT  6.835 33.4075 6.9 33.5425 ;
        RECT  6.835 33.4075 6.9 33.5425 ;
        RECT  7.025 33.4075 7.09 33.5425 ;
        RECT  7.195 33.4075 7.26 33.5425 ;
        RECT  7.195 32.4925 7.26 32.6275 ;
        RECT  6.6125 33.255 6.7475 33.32 ;
        RECT  6.8525 32.725 6.9875 32.79 ;
        RECT  7.3275 32.3125 7.8875 32.3775 ;
        RECT  7.3275 33.6575 7.8875 33.7225 ;
        RECT  7.755 33.2925 7.82 33.6575 ;
        RECT  7.755 32.3775 7.82 32.5125 ;
        RECT  7.395 32.3775 7.46 32.4475 ;
        RECT  7.395 33.5675 7.46 33.6575 ;
        RECT  7.585 32.48 7.65 33.4275 ;
        RECT  7.3275 32.895 7.3625 32.96 ;
        RECT  7.65 32.895 7.8875 32.96 ;
        RECT  7.395 32.5825 7.46 32.7175 ;
        RECT  7.585 32.5825 7.65 32.7175 ;
        RECT  7.395 33.2925 7.46 33.5675 ;
        RECT  7.585 33.2925 7.65 33.5675 ;
        RECT  7.755 33.2925 7.82 33.5675 ;
        RECT  7.755 32.4475 7.82 32.5825 ;
        RECT  7.3625 32.895 7.4975 32.96 ;
        RECT  6.5775 33.2575 6.7125 33.3225 ;
        RECT  5.565 33.255 5.63 33.39 ;
        RECT  5.4925 35.0025 5.6275 35.0675 ;
        RECT  5.9475 35.0025 6.0825 35.0675 ;
        RECT  6.0175 35.0025 6.5775 35.0675 ;
        RECT  6.0175 33.6575 6.5775 33.7225 ;
        RECT  6.445 33.7225 6.51 34.0875 ;
        RECT  6.445 34.8675 6.51 35.0025 ;
        RECT  6.085 34.9325 6.15 35.0025 ;
        RECT  6.085 33.7225 6.15 33.8125 ;
        RECT  6.275 33.9525 6.34 34.9 ;
        RECT  6.0175 34.42 6.0525 34.485 ;
        RECT  6.34 34.42 6.5775 34.485 ;
        RECT  6.085 34.7325 6.15 34.8675 ;
        RECT  6.275 34.7325 6.34 34.8675 ;
        RECT  6.085 34.1925 6.15 34.4675 ;
        RECT  6.275 34.1925 6.34 34.4675 ;
        RECT  6.445 34.0875 6.51 34.3625 ;
        RECT  6.445 34.9325 6.51 35.0675 ;
        RECT  6.0525 34.495 6.1875 34.56 ;
        RECT  6.5775 35.0025 7.3275 35.0675 ;
        RECT  6.5775 33.6575 7.3275 33.7225 ;
        RECT  7.195 33.69 7.26 33.9725 ;
        RECT  7.195 34.855 7.26 35.035 ;
        RECT  6.645 33.69 6.71 33.9725 ;
        RECT  7.025 33.69 7.09 33.9725 ;
        RECT  6.645 34.7525 6.71 35.035 ;
        RECT  7.0575 34.075 7.1225 34.14 ;
        RECT  6.835 34.075 6.9 34.14 ;
        RECT  7.0575 34.1075 7.1225 34.8875 ;
        RECT  6.8675 34.075 7.09 34.14 ;
        RECT  6.835 33.9725 6.9 34.1075 ;
        RECT  6.5775 34.06 6.6125 34.125 ;
        RECT  6.5775 34.59 6.8525 34.655 ;
        RECT  7.09 34.3725 7.3275 34.4375 ;
        RECT  6.645 34.5975 6.71 34.7325 ;
        RECT  6.835 34.5975 6.9 34.7325 ;
        RECT  6.835 34.5975 6.9 34.7325 ;
        RECT  7.025 34.5975 7.09 34.7325 ;
        RECT  6.645 34.1275 6.71 34.2625 ;
        RECT  6.835 34.1275 6.9 34.2625 ;
        RECT  6.835 34.1275 6.9 34.2625 ;
        RECT  7.025 34.1275 7.09 34.2625 ;
        RECT  7.195 33.9725 7.26 34.1075 ;
        RECT  7.195 34.8875 7.26 35.0225 ;
        RECT  6.6125 34.135 6.7475 34.2 ;
        RECT  6.8525 34.665 6.9875 34.73 ;
        RECT  7.3275 35.0025 7.8875 35.0675 ;
        RECT  7.3275 33.6575 7.8875 33.7225 ;
        RECT  7.755 33.7225 7.82 34.0875 ;
        RECT  7.755 34.8675 7.82 35.0025 ;
        RECT  7.395 34.9325 7.46 35.0025 ;
        RECT  7.395 33.7225 7.46 33.8125 ;
        RECT  7.585 33.9525 7.65 34.9 ;
        RECT  7.3275 34.42 7.3625 34.485 ;
        RECT  7.65 34.42 7.8875 34.485 ;
        RECT  7.395 34.7325 7.46 34.8675 ;
        RECT  7.585 34.7325 7.65 34.8675 ;
        RECT  7.395 34.1925 7.46 34.4675 ;
        RECT  7.585 34.1925 7.65 34.4675 ;
        RECT  7.755 34.0875 7.82 34.3625 ;
        RECT  7.755 34.9325 7.82 35.0675 ;
        RECT  7.3625 34.495 7.4975 34.56 ;
        RECT  6.5775 34.0575 6.7125 34.1225 ;
        RECT  5.565 33.99 5.63 34.125 ;
        RECT  5.4925 36.3475 5.6275 36.4125 ;
        RECT  5.9475 36.3475 6.0825 36.4125 ;
        RECT  6.0175 35.0025 6.5775 35.0675 ;
        RECT  6.0175 36.3475 6.5775 36.4125 ;
        RECT  6.445 35.9825 6.51 36.3475 ;
        RECT  6.445 35.0675 6.51 35.2025 ;
        RECT  6.085 35.0675 6.15 35.1375 ;
        RECT  6.085 36.2575 6.15 36.3475 ;
        RECT  6.275 35.17 6.34 36.1175 ;
        RECT  6.0175 35.585 6.0525 35.65 ;
        RECT  6.34 35.585 6.5775 35.65 ;
        RECT  6.085 35.2725 6.15 35.4075 ;
        RECT  6.275 35.2725 6.34 35.4075 ;
        RECT  6.085 35.9825 6.15 36.2575 ;
        RECT  6.275 35.9825 6.34 36.2575 ;
        RECT  6.445 35.9825 6.51 36.2575 ;
        RECT  6.445 35.1375 6.51 35.2725 ;
        RECT  6.0525 35.585 6.1875 35.65 ;
        RECT  6.5775 35.0025 7.3275 35.0675 ;
        RECT  6.5775 36.3475 7.3275 36.4125 ;
        RECT  7.195 36.0975 7.26 36.38 ;
        RECT  7.195 35.035 7.26 35.215 ;
        RECT  6.645 36.0975 6.71 36.38 ;
        RECT  7.025 36.0975 7.09 36.38 ;
        RECT  6.645 35.035 6.71 35.3175 ;
        RECT  7.0575 35.93 7.1225 35.995 ;
        RECT  6.835 35.93 6.9 35.995 ;
        RECT  7.0575 35.1825 7.1225 35.9625 ;
        RECT  6.8675 35.93 7.09 35.995 ;
        RECT  6.835 35.9625 6.9 36.0975 ;
        RECT  6.5775 35.945 6.6125 36.01 ;
        RECT  6.5775 35.415 6.8525 35.48 ;
        RECT  7.09 35.6325 7.3275 35.6975 ;
        RECT  6.645 35.3175 6.71 35.4525 ;
        RECT  6.835 35.3175 6.9 35.4525 ;
        RECT  6.835 35.3175 6.9 35.4525 ;
        RECT  7.025 35.3175 7.09 35.4525 ;
        RECT  6.645 36.0975 6.71 36.2325 ;
        RECT  6.835 36.0975 6.9 36.2325 ;
        RECT  6.835 36.0975 6.9 36.2325 ;
        RECT  7.025 36.0975 7.09 36.2325 ;
        RECT  7.195 36.0975 7.26 36.2325 ;
        RECT  7.195 35.1825 7.26 35.3175 ;
        RECT  6.6125 35.945 6.7475 36.01 ;
        RECT  6.8525 35.415 6.9875 35.48 ;
        RECT  7.3275 35.0025 7.8875 35.0675 ;
        RECT  7.3275 36.3475 7.8875 36.4125 ;
        RECT  7.755 35.9825 7.82 36.3475 ;
        RECT  7.755 35.0675 7.82 35.2025 ;
        RECT  7.395 35.0675 7.46 35.1375 ;
        RECT  7.395 36.2575 7.46 36.3475 ;
        RECT  7.585 35.17 7.65 36.1175 ;
        RECT  7.3275 35.585 7.3625 35.65 ;
        RECT  7.65 35.585 7.8875 35.65 ;
        RECT  7.395 35.2725 7.46 35.4075 ;
        RECT  7.585 35.2725 7.65 35.4075 ;
        RECT  7.395 35.9825 7.46 36.2575 ;
        RECT  7.585 35.9825 7.65 36.2575 ;
        RECT  7.755 35.9825 7.82 36.2575 ;
        RECT  7.755 35.1375 7.82 35.2725 ;
        RECT  7.3625 35.585 7.4975 35.65 ;
        RECT  6.5775 35.9475 6.7125 36.0125 ;
        RECT  5.565 35.945 5.63 36.08 ;
        RECT  5.4925 37.6925 5.6275 37.7575 ;
        RECT  5.9475 37.6925 6.0825 37.7575 ;
        RECT  6.0175 37.6925 6.5775 37.7575 ;
        RECT  6.0175 36.3475 6.5775 36.4125 ;
        RECT  6.445 36.4125 6.51 36.7775 ;
        RECT  6.445 37.5575 6.51 37.6925 ;
        RECT  6.085 37.6225 6.15 37.6925 ;
        RECT  6.085 36.4125 6.15 36.5025 ;
        RECT  6.275 36.6425 6.34 37.59 ;
        RECT  6.0175 37.11 6.0525 37.175 ;
        RECT  6.34 37.11 6.5775 37.175 ;
        RECT  6.085 37.4225 6.15 37.5575 ;
        RECT  6.275 37.4225 6.34 37.5575 ;
        RECT  6.085 36.8825 6.15 37.1575 ;
        RECT  6.275 36.8825 6.34 37.1575 ;
        RECT  6.445 36.7775 6.51 37.0525 ;
        RECT  6.445 37.6225 6.51 37.7575 ;
        RECT  6.0525 37.185 6.1875 37.25 ;
        RECT  6.5775 37.6925 7.3275 37.7575 ;
        RECT  6.5775 36.3475 7.3275 36.4125 ;
        RECT  7.195 36.38 7.26 36.6625 ;
        RECT  7.195 37.545 7.26 37.725 ;
        RECT  6.645 36.38 6.71 36.6625 ;
        RECT  7.025 36.38 7.09 36.6625 ;
        RECT  6.645 37.4425 6.71 37.725 ;
        RECT  7.0575 36.765 7.1225 36.83 ;
        RECT  6.835 36.765 6.9 36.83 ;
        RECT  7.0575 36.7975 7.1225 37.5775 ;
        RECT  6.8675 36.765 7.09 36.83 ;
        RECT  6.835 36.6625 6.9 36.7975 ;
        RECT  6.5775 36.75 6.6125 36.815 ;
        RECT  6.5775 37.28 6.8525 37.345 ;
        RECT  7.09 37.0625 7.3275 37.1275 ;
        RECT  6.645 37.2875 6.71 37.4225 ;
        RECT  6.835 37.2875 6.9 37.4225 ;
        RECT  6.835 37.2875 6.9 37.4225 ;
        RECT  7.025 37.2875 7.09 37.4225 ;
        RECT  6.645 36.8175 6.71 36.9525 ;
        RECT  6.835 36.8175 6.9 36.9525 ;
        RECT  6.835 36.8175 6.9 36.9525 ;
        RECT  7.025 36.8175 7.09 36.9525 ;
        RECT  7.195 36.6625 7.26 36.7975 ;
        RECT  7.195 37.5775 7.26 37.7125 ;
        RECT  6.6125 36.825 6.7475 36.89 ;
        RECT  6.8525 37.355 6.9875 37.42 ;
        RECT  7.3275 37.6925 7.8875 37.7575 ;
        RECT  7.3275 36.3475 7.8875 36.4125 ;
        RECT  7.755 36.4125 7.82 36.7775 ;
        RECT  7.755 37.5575 7.82 37.6925 ;
        RECT  7.395 37.6225 7.46 37.6925 ;
        RECT  7.395 36.4125 7.46 36.5025 ;
        RECT  7.585 36.6425 7.65 37.59 ;
        RECT  7.3275 37.11 7.3625 37.175 ;
        RECT  7.65 37.11 7.8875 37.175 ;
        RECT  7.395 37.4225 7.46 37.5575 ;
        RECT  7.585 37.4225 7.65 37.5575 ;
        RECT  7.395 36.8825 7.46 37.1575 ;
        RECT  7.585 36.8825 7.65 37.1575 ;
        RECT  7.755 36.7775 7.82 37.0525 ;
        RECT  7.755 37.6225 7.82 37.7575 ;
        RECT  7.3625 37.185 7.4975 37.25 ;
        RECT  6.5775 36.7475 6.7125 36.8125 ;
        RECT  5.565 36.68 5.63 36.815 ;
        RECT  5.4925 39.0375 5.6275 39.1025 ;
        RECT  5.9475 39.0375 6.0825 39.1025 ;
        RECT  6.0175 37.6925 6.5775 37.7575 ;
        RECT  6.0175 39.0375 6.5775 39.1025 ;
        RECT  6.445 38.6725 6.51 39.0375 ;
        RECT  6.445 37.7575 6.51 37.8925 ;
        RECT  6.085 37.7575 6.15 37.8275 ;
        RECT  6.085 38.9475 6.15 39.0375 ;
        RECT  6.275 37.86 6.34 38.8075 ;
        RECT  6.0175 38.275 6.0525 38.34 ;
        RECT  6.34 38.275 6.5775 38.34 ;
        RECT  6.085 37.9625 6.15 38.0975 ;
        RECT  6.275 37.9625 6.34 38.0975 ;
        RECT  6.085 38.6725 6.15 38.9475 ;
        RECT  6.275 38.6725 6.34 38.9475 ;
        RECT  6.445 38.6725 6.51 38.9475 ;
        RECT  6.445 37.8275 6.51 37.9625 ;
        RECT  6.0525 38.275 6.1875 38.34 ;
        RECT  6.5775 37.6925 7.3275 37.7575 ;
        RECT  6.5775 39.0375 7.3275 39.1025 ;
        RECT  7.195 38.7875 7.26 39.07 ;
        RECT  7.195 37.725 7.26 37.905 ;
        RECT  6.645 38.7875 6.71 39.07 ;
        RECT  7.025 38.7875 7.09 39.07 ;
        RECT  6.645 37.725 6.71 38.0075 ;
        RECT  7.0575 38.62 7.1225 38.685 ;
        RECT  6.835 38.62 6.9 38.685 ;
        RECT  7.0575 37.8725 7.1225 38.6525 ;
        RECT  6.8675 38.62 7.09 38.685 ;
        RECT  6.835 38.6525 6.9 38.7875 ;
        RECT  6.5775 38.635 6.6125 38.7 ;
        RECT  6.5775 38.105 6.8525 38.17 ;
        RECT  7.09 38.3225 7.3275 38.3875 ;
        RECT  6.645 38.0075 6.71 38.1425 ;
        RECT  6.835 38.0075 6.9 38.1425 ;
        RECT  6.835 38.0075 6.9 38.1425 ;
        RECT  7.025 38.0075 7.09 38.1425 ;
        RECT  6.645 38.7875 6.71 38.9225 ;
        RECT  6.835 38.7875 6.9 38.9225 ;
        RECT  6.835 38.7875 6.9 38.9225 ;
        RECT  7.025 38.7875 7.09 38.9225 ;
        RECT  7.195 38.7875 7.26 38.9225 ;
        RECT  7.195 37.8725 7.26 38.0075 ;
        RECT  6.6125 38.635 6.7475 38.7 ;
        RECT  6.8525 38.105 6.9875 38.17 ;
        RECT  7.3275 37.6925 7.8875 37.7575 ;
        RECT  7.3275 39.0375 7.8875 39.1025 ;
        RECT  7.755 38.6725 7.82 39.0375 ;
        RECT  7.755 37.7575 7.82 37.8925 ;
        RECT  7.395 37.7575 7.46 37.8275 ;
        RECT  7.395 38.9475 7.46 39.0375 ;
        RECT  7.585 37.86 7.65 38.8075 ;
        RECT  7.3275 38.275 7.3625 38.34 ;
        RECT  7.65 38.275 7.8875 38.34 ;
        RECT  7.395 37.9625 7.46 38.0975 ;
        RECT  7.585 37.9625 7.65 38.0975 ;
        RECT  7.395 38.6725 7.46 38.9475 ;
        RECT  7.585 38.6725 7.65 38.9475 ;
        RECT  7.755 38.6725 7.82 38.9475 ;
        RECT  7.755 37.8275 7.82 37.9625 ;
        RECT  7.3625 38.275 7.4975 38.34 ;
        RECT  6.5775 38.6375 6.7125 38.7025 ;
        RECT  5.565 38.635 5.63 38.77 ;
        RECT  5.4925 40.3825 5.6275 40.4475 ;
        RECT  5.9475 40.3825 6.0825 40.4475 ;
        RECT  6.0175 40.3825 6.5775 40.4475 ;
        RECT  6.0175 39.0375 6.5775 39.1025 ;
        RECT  6.445 39.1025 6.51 39.4675 ;
        RECT  6.445 40.2475 6.51 40.3825 ;
        RECT  6.085 40.3125 6.15 40.3825 ;
        RECT  6.085 39.1025 6.15 39.1925 ;
        RECT  6.275 39.3325 6.34 40.28 ;
        RECT  6.0175 39.8 6.0525 39.865 ;
        RECT  6.34 39.8 6.5775 39.865 ;
        RECT  6.085 40.1125 6.15 40.2475 ;
        RECT  6.275 40.1125 6.34 40.2475 ;
        RECT  6.085 39.5725 6.15 39.8475 ;
        RECT  6.275 39.5725 6.34 39.8475 ;
        RECT  6.445 39.4675 6.51 39.7425 ;
        RECT  6.445 40.3125 6.51 40.4475 ;
        RECT  6.0525 39.875 6.1875 39.94 ;
        RECT  6.5775 40.3825 7.3275 40.4475 ;
        RECT  6.5775 39.0375 7.3275 39.1025 ;
        RECT  7.195 39.07 7.26 39.3525 ;
        RECT  7.195 40.235 7.26 40.415 ;
        RECT  6.645 39.07 6.71 39.3525 ;
        RECT  7.025 39.07 7.09 39.3525 ;
        RECT  6.645 40.1325 6.71 40.415 ;
        RECT  7.0575 39.455 7.1225 39.52 ;
        RECT  6.835 39.455 6.9 39.52 ;
        RECT  7.0575 39.4875 7.1225 40.2675 ;
        RECT  6.8675 39.455 7.09 39.52 ;
        RECT  6.835 39.3525 6.9 39.4875 ;
        RECT  6.5775 39.44 6.6125 39.505 ;
        RECT  6.5775 39.97 6.8525 40.035 ;
        RECT  7.09 39.7525 7.3275 39.8175 ;
        RECT  6.645 39.9775 6.71 40.1125 ;
        RECT  6.835 39.9775 6.9 40.1125 ;
        RECT  6.835 39.9775 6.9 40.1125 ;
        RECT  7.025 39.9775 7.09 40.1125 ;
        RECT  6.645 39.5075 6.71 39.6425 ;
        RECT  6.835 39.5075 6.9 39.6425 ;
        RECT  6.835 39.5075 6.9 39.6425 ;
        RECT  7.025 39.5075 7.09 39.6425 ;
        RECT  7.195 39.3525 7.26 39.4875 ;
        RECT  7.195 40.2675 7.26 40.4025 ;
        RECT  6.6125 39.515 6.7475 39.58 ;
        RECT  6.8525 40.045 6.9875 40.11 ;
        RECT  7.3275 40.3825 7.8875 40.4475 ;
        RECT  7.3275 39.0375 7.8875 39.1025 ;
        RECT  7.755 39.1025 7.82 39.4675 ;
        RECT  7.755 40.2475 7.82 40.3825 ;
        RECT  7.395 40.3125 7.46 40.3825 ;
        RECT  7.395 39.1025 7.46 39.1925 ;
        RECT  7.585 39.3325 7.65 40.28 ;
        RECT  7.3275 39.8 7.3625 39.865 ;
        RECT  7.65 39.8 7.8875 39.865 ;
        RECT  7.395 40.1125 7.46 40.2475 ;
        RECT  7.585 40.1125 7.65 40.2475 ;
        RECT  7.395 39.5725 7.46 39.8475 ;
        RECT  7.585 39.5725 7.65 39.8475 ;
        RECT  7.755 39.4675 7.82 39.7425 ;
        RECT  7.755 40.3125 7.82 40.4475 ;
        RECT  7.3625 39.875 7.4975 39.94 ;
        RECT  6.5775 39.4375 6.7125 39.5025 ;
        RECT  5.565 39.37 5.63 39.505 ;
        RECT  1.115 5.02 1.18 7.84 ;
        RECT  7.1125 5.02 7.1775 7.84 ;
        RECT  3.6325 7.235 3.7675 7.3 ;
        RECT  3.6325 7.42 3.7675 7.485 ;
        RECT  2.3975 7.235 2.5325 7.3 ;
        RECT  2.3975 7.42 2.5325 7.485 ;
        RECT  3.6325 7.425 3.7675 7.49 ;
        RECT  3.6325 7.61 3.7675 7.675 ;
        RECT  6.5925 7.425 6.7275 7.49 ;
        RECT  6.5925 7.61 6.7275 7.675 ;
        RECT  2.3975 7.425 2.5325 7.49 ;
        RECT  2.3975 7.61 2.5325 7.675 ;
        RECT  6.5925 7.235 6.7275 7.3 ;
        RECT  6.5925 7.42 6.7275 7.485 ;
        RECT  1.8625 7.425 1.9975 7.49 ;
        RECT  1.8625 7.61 1.9975 7.675 ;
        RECT  4.8225 7.285 4.9575 7.35 ;
        RECT  4.8225 7.47 4.9575 7.535 ;
        RECT  5.3575 7.235 5.4925 7.3 ;
        RECT  5.3575 7.42 5.4925 7.485 ;
        RECT  5.3575 7.425 5.4925 7.49 ;
        RECT  5.3575 7.61 5.4925 7.675 ;
        RECT  5.7825 7.235 5.9175 7.3 ;
        RECT  5.7825 7.42 5.9175 7.485 ;
        RECT  2.8225 7.235 2.9575 7.3 ;
        RECT  2.8225 7.42 2.9575 7.485 ;
        RECT  6.1675 7.235 6.3025 7.3 ;
        RECT  6.1675 7.42 6.3025 7.485 ;
        RECT  6.1675 7.425 6.3025 7.49 ;
        RECT  6.1675 7.61 6.3025 7.675 ;
        RECT  2.8225 7.425 2.9575 7.49 ;
        RECT  2.8225 7.61 2.9575 7.675 ;
        RECT  5.7825 7.425 5.9175 7.49 ;
        RECT  5.7825 7.61 5.9175 7.675 ;
        RECT  3.2075 7.425 3.3425 7.49 ;
        RECT  3.2075 7.61 3.3425 7.675 ;
        RECT  3.2075 7.235 3.3425 7.3 ;
        RECT  3.2075 7.42 3.3425 7.485 ;
        RECT  1.4375 7.425 1.5725 7.49 ;
        RECT  1.4375 7.61 1.5725 7.675 ;
        RECT  4.4125 7.35 4.5475 7.415 ;
        RECT  4.4125 7.535 4.5475 7.6 ;
        RECT  1.1475 7.4775 1.2125 7.6125 ;
        RECT  6.645 7.61 6.78 7.675 ;
        RECT  4.83 7.72 4.965 7.785 ;
        RECT  3.93 7.61 4.065 7.675 ;
        RECT  4.405 7.1875 4.54 7.2525 ;
        RECT  7.01 7.61 7.145 7.675 ;
        RECT  1.4675 7.1025 1.6025 7.1675 ;
        RECT  5.55 7.245 5.685 7.31 ;
        RECT  3.9425 7.2425 4.0775 7.3075 ;
        RECT  2.545 7.2425 2.68 7.3075 ;
        RECT  1.3275 7.8075 1.4625 7.8725 ;
        RECT  1.445 7.2325 1.58 7.2975 ;
        RECT  3.055 7.1625 3.12 7.2975 ;
        RECT  1.97 7.1925 2.105 7.2575 ;
        RECT  6.015 7.1625 6.08 7.2975 ;
        RECT  6.9025 7.285 7.0375 7.35 ;
        RECT  3.4325 7.365 3.5675 7.43 ;
        RECT  6.3925 7.375 6.5275 7.44 ;
        RECT  4.7025 7.5375 4.7675 7.6725 ;
        RECT  4.405 7.1025 4.54 7.1675 ;
        RECT  1.6975 7.6475 1.7625 7.7825 ;
        RECT  3.21 7.6075 3.345 7.6725 ;
        RECT  6.9025 7.2425 7.0375 7.3075 ;
        RECT  6.3925 7.42 6.5275 7.485 ;
        RECT  5.98 7.1025 6.115 7.1675 ;
        RECT  1.2775 7.1025 1.4125 7.1675 ;
        RECT  3.9425 7.2425 4.0775 7.3075 ;
        RECT  3.02 7.1025 3.155 7.1675 ;
        RECT  2.82 7.6075 2.955 7.6725 ;
        RECT  2.82 7.42 2.955 7.485 ;
        RECT  3.4325 7.42 3.5675 7.485 ;
        RECT  5.78 7.61 5.915 7.675 ;
        RECT  5.78 7.42 5.915 7.485 ;
        RECT  1.1475 7.1 1.2125 7.875 ;
        RECT  4.2175 7.74 7.1125 7.805 ;
        RECT  6.7275 7.235 7.0375 7.3 ;
        RECT  6.3025 7.61 6.5925 7.675 ;
        RECT  5.4925 7.61 5.7825 7.675 ;
        RECT  7.115 7.4625 7.1775 7.535 ;
        RECT  6.7275 7.42 7.1125 7.49 ;
        RECT  5.4925 7.42 5.7825 7.49 ;
        RECT  6.0125 7.42 6.17 7.49 ;
        RECT  6.3025 7.235 6.5925 7.3 ;
        RECT  5.4925 7.235 5.7825 7.3 ;
        RECT  6.0125 7.105 6.0825 7.49 ;
        RECT  7.1125 7.1 7.1775 7.875 ;
        RECT  5.1225 7.1 5.1875 7.875 ;
        RECT  2.2275 7.74 4.1525 7.805 ;
        RECT  3.7675 7.235 4.0775 7.3 ;
        RECT  3.3425 7.61 3.6325 7.675 ;
        RECT  4.5075 7.535 4.9575 7.6 ;
        RECT  3.7675 7.42 4.1525 7.49 ;
        RECT  3.0525 7.42 3.21 7.49 ;
        RECT  4.065 7.61 4.1525 7.675 ;
        RECT  3.3425 7.235 3.6325 7.3 ;
        RECT  4.2825 7.17 4.3475 7.415 ;
        RECT  4.2825 7.17 4.405 7.2525 ;
        RECT  4.405 7.165 4.54 7.2325 ;
        RECT  4.1525 7.1 4.2175 7.875 ;
        RECT  2.5325 7.61 2.8225 7.675 ;
        RECT  1.995 7.425 2.1625 7.49 ;
        RECT  1.5025 7.1675 1.5725 7.425 ;
        RECT  1.4375 7.61 1.8625 7.675 ;
        RECT  2.5325 7.42 2.8225 7.49 ;
        RECT  1.6925 7.61 1.7675 7.7825 ;
        RECT  2.5325 7.235 2.8225 7.3 ;
        RECT  1.3725 7.2325 1.445 7.2975 ;
        RECT  3.0525 7.105 3.1225 7.49 ;
        RECT  2.0825 7.1925 2.1975 7.2575 ;
        RECT  1.3075 7.1 1.3725 7.875 ;
        RECT  2.1625 7.1 2.2275 7.875 ;
        RECT  1.1525 7.67 1.21 7.735 ;
        RECT  1.3925 7.1025 1.515 7.1675 ;
        RECT  4.955 7.285 5.1225 7.35 ;
        RECT  4.3475 7.3475 4.45 7.415 ;
        RECT  3.6325 6.97 3.7675 7.035 ;
        RECT  3.6325 6.785 3.7675 6.85 ;
        RECT  2.3975 6.97 2.5325 7.035 ;
        RECT  2.3975 6.785 2.5325 6.85 ;
        RECT  3.6325 6.78 3.7675 6.845 ;
        RECT  3.6325 6.595 3.7675 6.66 ;
        RECT  6.5925 6.78 6.7275 6.845 ;
        RECT  6.5925 6.595 6.7275 6.66 ;
        RECT  2.3975 6.78 2.5325 6.845 ;
        RECT  2.3975 6.595 2.5325 6.66 ;
        RECT  6.5925 6.97 6.7275 7.035 ;
        RECT  6.5925 6.785 6.7275 6.85 ;
        RECT  1.8625 6.78 1.9975 6.845 ;
        RECT  1.8625 6.595 1.9975 6.66 ;
        RECT  4.8225 6.92 4.9575 6.985 ;
        RECT  4.8225 6.735 4.9575 6.8 ;
        RECT  5.3575 6.97 5.4925 7.035 ;
        RECT  5.3575 6.785 5.4925 6.85 ;
        RECT  5.3575 6.78 5.4925 6.845 ;
        RECT  5.3575 6.595 5.4925 6.66 ;
        RECT  5.7825 6.97 5.9175 7.035 ;
        RECT  5.7825 6.785 5.9175 6.85 ;
        RECT  2.8225 6.97 2.9575 7.035 ;
        RECT  2.8225 6.785 2.9575 6.85 ;
        RECT  6.1675 6.97 6.3025 7.035 ;
        RECT  6.1675 6.785 6.3025 6.85 ;
        RECT  6.1675 6.78 6.3025 6.845 ;
        RECT  6.1675 6.595 6.3025 6.66 ;
        RECT  2.8225 6.78 2.9575 6.845 ;
        RECT  2.8225 6.595 2.9575 6.66 ;
        RECT  5.7825 6.78 5.9175 6.845 ;
        RECT  5.7825 6.595 5.9175 6.66 ;
        RECT  3.2075 6.78 3.3425 6.845 ;
        RECT  3.2075 6.595 3.3425 6.66 ;
        RECT  3.2075 6.97 3.3425 7.035 ;
        RECT  3.2075 6.785 3.3425 6.85 ;
        RECT  1.4375 6.78 1.5725 6.845 ;
        RECT  1.4375 6.595 1.5725 6.66 ;
        RECT  4.4125 6.855 4.5475 6.92 ;
        RECT  4.4125 6.67 4.5475 6.735 ;
        RECT  1.1475 6.6575 1.2125 6.7925 ;
        RECT  6.645 6.595 6.78 6.66 ;
        RECT  4.83 6.485 4.965 6.55 ;
        RECT  3.93 6.595 4.065 6.66 ;
        RECT  4.405 7.0175 4.54 7.0825 ;
        RECT  7.01 6.595 7.145 6.66 ;
        RECT  1.4675 7.1025 1.6025 7.1675 ;
        RECT  5.55 6.96 5.685 7.025 ;
        RECT  3.9425 6.9625 4.0775 7.0275 ;
        RECT  2.545 6.9625 2.68 7.0275 ;
        RECT  1.3275 6.3975 1.4625 6.4625 ;
        RECT  1.445 6.9725 1.58 7.0375 ;
        RECT  3.055 6.9725 3.12 7.1075 ;
        RECT  1.97 7.0125 2.105 7.0775 ;
        RECT  6.015 6.9725 6.08 7.1075 ;
        RECT  6.9025 6.92 7.0375 6.985 ;
        RECT  3.4325 6.84 3.5675 6.905 ;
        RECT  6.3925 6.83 6.5275 6.895 ;
        RECT  4.7025 6.5975 4.7675 6.7325 ;
        RECT  4.405 7.1025 4.54 7.1675 ;
        RECT  1.6975 6.4875 1.7625 6.6225 ;
        RECT  3.21 6.5975 3.345 6.6625 ;
        RECT  6.9025 6.9625 7.0375 7.0275 ;
        RECT  6.3925 6.785 6.5275 6.85 ;
        RECT  5.98 7.1025 6.115 7.1675 ;
        RECT  1.2775 7.1025 1.4125 7.1675 ;
        RECT  3.9425 6.9625 4.0775 7.0275 ;
        RECT  3.02 7.1025 3.155 7.1675 ;
        RECT  2.82 6.5975 2.955 6.6625 ;
        RECT  2.82 6.785 2.955 6.85 ;
        RECT  3.4325 6.785 3.5675 6.85 ;
        RECT  5.78 6.595 5.915 6.66 ;
        RECT  5.78 6.785 5.915 6.85 ;
        RECT  1.1475 6.395 1.2125 7.17 ;
        RECT  4.2175 6.465 7.1125 6.53 ;
        RECT  6.7275 6.97 7.0375 7.035 ;
        RECT  6.3025 6.595 6.5925 6.66 ;
        RECT  5.4925 6.595 5.7825 6.66 ;
        RECT  7.115 6.735 7.1775 6.8075 ;
        RECT  6.7275 6.78 7.1125 6.85 ;
        RECT  5.4925 6.78 5.7825 6.85 ;
        RECT  6.0125 6.78 6.17 6.85 ;
        RECT  6.3025 6.97 6.5925 7.035 ;
        RECT  5.4925 6.97 5.7825 7.035 ;
        RECT  6.0125 6.78 6.0825 7.165 ;
        RECT  7.1125 6.395 7.1775 7.17 ;
        RECT  5.1225 6.395 5.1875 7.17 ;
        RECT  2.2275 6.465 4.1525 6.53 ;
        RECT  3.7675 6.97 4.0775 7.035 ;
        RECT  3.3425 6.595 3.6325 6.66 ;
        RECT  4.5075 6.67 4.9575 6.735 ;
        RECT  3.7675 6.78 4.1525 6.85 ;
        RECT  3.0525 6.78 3.21 6.85 ;
        RECT  4.065 6.595 4.1525 6.66 ;
        RECT  3.3425 6.97 3.6325 7.035 ;
        RECT  4.2825 6.855 4.3475 7.1 ;
        RECT  4.2825 7.0175 4.405 7.1 ;
        RECT  4.405 7.0375 4.54 7.105 ;
        RECT  4.1525 6.395 4.2175 7.17 ;
        RECT  2.5325 6.595 2.8225 6.66 ;
        RECT  1.995 6.78 2.1625 6.845 ;
        RECT  1.5025 6.845 1.5725 7.1025 ;
        RECT  1.4375 6.595 1.8625 6.66 ;
        RECT  2.5325 6.78 2.8225 6.85 ;
        RECT  1.6925 6.4875 1.7675 6.66 ;
        RECT  2.5325 6.97 2.8225 7.035 ;
        RECT  1.3725 6.9725 1.445 7.0375 ;
        RECT  3.0525 6.78 3.1225 7.165 ;
        RECT  2.0825 7.0125 2.1975 7.0775 ;
        RECT  1.3075 6.395 1.3725 7.17 ;
        RECT  2.1625 6.395 2.2275 7.17 ;
        RECT  1.1525 6.535 1.21 6.6 ;
        RECT  1.3925 7.1025 1.515 7.1675 ;
        RECT  4.955 6.92 5.1225 6.985 ;
        RECT  4.3475 6.855 4.45 6.9225 ;
        RECT  3.6325 5.825 3.7675 5.89 ;
        RECT  3.6325 6.01 3.7675 6.075 ;
        RECT  2.3975 5.825 2.5325 5.89 ;
        RECT  2.3975 6.01 2.5325 6.075 ;
        RECT  3.6325 6.015 3.7675 6.08 ;
        RECT  3.6325 6.2 3.7675 6.265 ;
        RECT  6.5925 6.015 6.7275 6.08 ;
        RECT  6.5925 6.2 6.7275 6.265 ;
        RECT  2.3975 6.015 2.5325 6.08 ;
        RECT  2.3975 6.2 2.5325 6.265 ;
        RECT  6.5925 5.825 6.7275 5.89 ;
        RECT  6.5925 6.01 6.7275 6.075 ;
        RECT  1.8625 6.015 1.9975 6.08 ;
        RECT  1.8625 6.2 1.9975 6.265 ;
        RECT  4.8225 5.875 4.9575 5.94 ;
        RECT  4.8225 6.06 4.9575 6.125 ;
        RECT  5.3575 5.825 5.4925 5.89 ;
        RECT  5.3575 6.01 5.4925 6.075 ;
        RECT  5.3575 6.015 5.4925 6.08 ;
        RECT  5.3575 6.2 5.4925 6.265 ;
        RECT  5.7825 5.825 5.9175 5.89 ;
        RECT  5.7825 6.01 5.9175 6.075 ;
        RECT  2.8225 5.825 2.9575 5.89 ;
        RECT  2.8225 6.01 2.9575 6.075 ;
        RECT  6.1675 5.825 6.3025 5.89 ;
        RECT  6.1675 6.01 6.3025 6.075 ;
        RECT  6.1675 6.015 6.3025 6.08 ;
        RECT  6.1675 6.2 6.3025 6.265 ;
        RECT  2.8225 6.015 2.9575 6.08 ;
        RECT  2.8225 6.2 2.9575 6.265 ;
        RECT  5.7825 6.015 5.9175 6.08 ;
        RECT  5.7825 6.2 5.9175 6.265 ;
        RECT  3.2075 6.015 3.3425 6.08 ;
        RECT  3.2075 6.2 3.3425 6.265 ;
        RECT  3.2075 5.825 3.3425 5.89 ;
        RECT  3.2075 6.01 3.3425 6.075 ;
        RECT  1.4375 6.015 1.5725 6.08 ;
        RECT  1.4375 6.2 1.5725 6.265 ;
        RECT  4.4125 5.94 4.5475 6.005 ;
        RECT  4.4125 6.125 4.5475 6.19 ;
        RECT  1.1475 6.0675 1.2125 6.2025 ;
        RECT  6.645 6.2 6.78 6.265 ;
        RECT  4.83 6.31 4.965 6.375 ;
        RECT  3.93 6.2 4.065 6.265 ;
        RECT  4.405 5.7775 4.54 5.8425 ;
        RECT  7.01 6.2 7.145 6.265 ;
        RECT  1.4675 5.6925 1.6025 5.7575 ;
        RECT  5.55 5.835 5.685 5.9 ;
        RECT  3.9425 5.8325 4.0775 5.8975 ;
        RECT  2.545 5.8325 2.68 5.8975 ;
        RECT  1.3275 6.3975 1.4625 6.4625 ;
        RECT  1.445 5.8225 1.58 5.8875 ;
        RECT  3.055 5.7525 3.12 5.8875 ;
        RECT  1.97 5.7825 2.105 5.8475 ;
        RECT  6.015 5.7525 6.08 5.8875 ;
        RECT  6.9025 5.875 7.0375 5.94 ;
        RECT  3.4325 5.955 3.5675 6.02 ;
        RECT  6.3925 5.965 6.5275 6.03 ;
        RECT  4.7025 6.1275 4.7675 6.2625 ;
        RECT  4.405 5.6925 4.54 5.7575 ;
        RECT  1.6975 6.2375 1.7625 6.3725 ;
        RECT  3.21 6.1975 3.345 6.2625 ;
        RECT  6.9025 5.8325 7.0375 5.8975 ;
        RECT  6.3925 6.01 6.5275 6.075 ;
        RECT  5.98 5.6925 6.115 5.7575 ;
        RECT  1.2775 5.6925 1.4125 5.7575 ;
        RECT  3.9425 5.8325 4.0775 5.8975 ;
        RECT  3.02 5.6925 3.155 5.7575 ;
        RECT  2.82 6.1975 2.955 6.2625 ;
        RECT  2.82 6.01 2.955 6.075 ;
        RECT  3.4325 6.01 3.5675 6.075 ;
        RECT  5.78 6.2 5.915 6.265 ;
        RECT  5.78 6.01 5.915 6.075 ;
        RECT  1.1475 5.69 1.2125 6.465 ;
        RECT  4.2175 6.33 7.1125 6.395 ;
        RECT  6.7275 5.825 7.0375 5.89 ;
        RECT  6.3025 6.2 6.5925 6.265 ;
        RECT  5.4925 6.2 5.7825 6.265 ;
        RECT  7.115 6.0525 7.1775 6.125 ;
        RECT  6.7275 6.01 7.1125 6.08 ;
        RECT  5.4925 6.01 5.7825 6.08 ;
        RECT  6.0125 6.01 6.17 6.08 ;
        RECT  6.3025 5.825 6.5925 5.89 ;
        RECT  5.4925 5.825 5.7825 5.89 ;
        RECT  6.0125 5.695 6.0825 6.08 ;
        RECT  7.1125 5.69 7.1775 6.465 ;
        RECT  5.1225 5.69 5.1875 6.465 ;
        RECT  2.2275 6.33 4.1525 6.395 ;
        RECT  3.7675 5.825 4.0775 5.89 ;
        RECT  3.3425 6.2 3.6325 6.265 ;
        RECT  4.5075 6.125 4.9575 6.19 ;
        RECT  3.7675 6.01 4.1525 6.08 ;
        RECT  3.0525 6.01 3.21 6.08 ;
        RECT  4.065 6.2 4.1525 6.265 ;
        RECT  3.3425 5.825 3.6325 5.89 ;
        RECT  4.2825 5.76 4.3475 6.005 ;
        RECT  4.2825 5.76 4.405 5.8425 ;
        RECT  4.405 5.755 4.54 5.8225 ;
        RECT  4.1525 5.69 4.2175 6.465 ;
        RECT  2.5325 6.2 2.8225 6.265 ;
        RECT  1.995 6.015 2.1625 6.08 ;
        RECT  1.5025 5.7575 1.5725 6.015 ;
        RECT  1.4375 6.2 1.8625 6.265 ;
        RECT  2.5325 6.01 2.8225 6.08 ;
        RECT  1.6925 6.2 1.7675 6.3725 ;
        RECT  2.5325 5.825 2.8225 5.89 ;
        RECT  1.3725 5.8225 1.445 5.8875 ;
        RECT  3.0525 5.695 3.1225 6.08 ;
        RECT  2.0825 5.7825 2.1975 5.8475 ;
        RECT  1.3075 5.69 1.3725 6.465 ;
        RECT  2.1625 5.69 2.2275 6.465 ;
        RECT  1.1525 6.26 1.21 6.325 ;
        RECT  1.3925 5.6925 1.515 5.7575 ;
        RECT  4.955 5.875 5.1225 5.94 ;
        RECT  4.3475 5.9375 4.45 6.005 ;
        RECT  3.6325 5.56 3.7675 5.625 ;
        RECT  3.6325 5.375 3.7675 5.44 ;
        RECT  2.3975 5.56 2.5325 5.625 ;
        RECT  2.3975 5.375 2.5325 5.44 ;
        RECT  3.6325 5.37 3.7675 5.435 ;
        RECT  3.6325 5.185 3.7675 5.25 ;
        RECT  6.5925 5.37 6.7275 5.435 ;
        RECT  6.5925 5.185 6.7275 5.25 ;
        RECT  2.3975 5.37 2.5325 5.435 ;
        RECT  2.3975 5.185 2.5325 5.25 ;
        RECT  6.5925 5.56 6.7275 5.625 ;
        RECT  6.5925 5.375 6.7275 5.44 ;
        RECT  1.8625 5.37 1.9975 5.435 ;
        RECT  1.8625 5.185 1.9975 5.25 ;
        RECT  4.8225 5.51 4.9575 5.575 ;
        RECT  4.8225 5.325 4.9575 5.39 ;
        RECT  5.3575 5.56 5.4925 5.625 ;
        RECT  5.3575 5.375 5.4925 5.44 ;
        RECT  5.3575 5.37 5.4925 5.435 ;
        RECT  5.3575 5.185 5.4925 5.25 ;
        RECT  5.7825 5.56 5.9175 5.625 ;
        RECT  5.7825 5.375 5.9175 5.44 ;
        RECT  2.8225 5.56 2.9575 5.625 ;
        RECT  2.8225 5.375 2.9575 5.44 ;
        RECT  6.1675 5.56 6.3025 5.625 ;
        RECT  6.1675 5.375 6.3025 5.44 ;
        RECT  6.1675 5.37 6.3025 5.435 ;
        RECT  6.1675 5.185 6.3025 5.25 ;
        RECT  2.8225 5.37 2.9575 5.435 ;
        RECT  2.8225 5.185 2.9575 5.25 ;
        RECT  5.7825 5.37 5.9175 5.435 ;
        RECT  5.7825 5.185 5.9175 5.25 ;
        RECT  3.2075 5.37 3.3425 5.435 ;
        RECT  3.2075 5.185 3.3425 5.25 ;
        RECT  3.2075 5.56 3.3425 5.625 ;
        RECT  3.2075 5.375 3.3425 5.44 ;
        RECT  1.4375 5.37 1.5725 5.435 ;
        RECT  1.4375 5.185 1.5725 5.25 ;
        RECT  4.4125 5.445 4.5475 5.51 ;
        RECT  4.4125 5.26 4.5475 5.325 ;
        RECT  1.1475 5.2475 1.2125 5.3825 ;
        RECT  6.645 5.185 6.78 5.25 ;
        RECT  4.83 5.075 4.965 5.14 ;
        RECT  3.93 5.185 4.065 5.25 ;
        RECT  4.405 5.6075 4.54 5.6725 ;
        RECT  7.01 5.185 7.145 5.25 ;
        RECT  1.4675 5.6925 1.6025 5.7575 ;
        RECT  5.55 5.55 5.685 5.615 ;
        RECT  3.9425 5.5525 4.0775 5.6175 ;
        RECT  2.545 5.5525 2.68 5.6175 ;
        RECT  1.3275 4.9875 1.4625 5.0525 ;
        RECT  1.445 5.5625 1.58 5.6275 ;
        RECT  3.055 5.5625 3.12 5.6975 ;
        RECT  1.97 5.6025 2.105 5.6675 ;
        RECT  6.015 5.5625 6.08 5.6975 ;
        RECT  6.9025 5.51 7.0375 5.575 ;
        RECT  3.4325 5.43 3.5675 5.495 ;
        RECT  6.3925 5.42 6.5275 5.485 ;
        RECT  4.7025 5.1875 4.7675 5.3225 ;
        RECT  4.405 5.6925 4.54 5.7575 ;
        RECT  1.6975 5.0775 1.7625 5.2125 ;
        RECT  3.21 5.1875 3.345 5.2525 ;
        RECT  6.9025 5.5525 7.0375 5.6175 ;
        RECT  6.3925 5.375 6.5275 5.44 ;
        RECT  5.98 5.6925 6.115 5.7575 ;
        RECT  1.2775 5.6925 1.4125 5.7575 ;
        RECT  3.9425 5.5525 4.0775 5.6175 ;
        RECT  3.02 5.6925 3.155 5.7575 ;
        RECT  2.82 5.1875 2.955 5.2525 ;
        RECT  2.82 5.375 2.955 5.44 ;
        RECT  3.4325 5.375 3.5675 5.44 ;
        RECT  5.78 5.185 5.915 5.25 ;
        RECT  5.78 5.375 5.915 5.44 ;
        RECT  1.1475 4.985 1.2125 5.76 ;
        RECT  4.2175 5.055 7.1125 5.12 ;
        RECT  6.7275 5.56 7.0375 5.625 ;
        RECT  6.3025 5.185 6.5925 5.25 ;
        RECT  5.4925 5.185 5.7825 5.25 ;
        RECT  7.115 5.325 7.1775 5.3975 ;
        RECT  6.7275 5.37 7.1125 5.44 ;
        RECT  5.4925 5.37 5.7825 5.44 ;
        RECT  6.0125 5.37 6.17 5.44 ;
        RECT  6.3025 5.56 6.5925 5.625 ;
        RECT  5.4925 5.56 5.7825 5.625 ;
        RECT  6.0125 5.37 6.0825 5.755 ;
        RECT  7.1125 4.985 7.1775 5.76 ;
        RECT  5.1225 4.985 5.1875 5.76 ;
        RECT  2.2275 5.055 4.1525 5.12 ;
        RECT  3.7675 5.56 4.0775 5.625 ;
        RECT  3.3425 5.185 3.6325 5.25 ;
        RECT  4.5075 5.26 4.9575 5.325 ;
        RECT  3.7675 5.37 4.1525 5.44 ;
        RECT  3.0525 5.37 3.21 5.44 ;
        RECT  4.065 5.185 4.1525 5.25 ;
        RECT  3.3425 5.56 3.6325 5.625 ;
        RECT  4.2825 5.445 4.3475 5.69 ;
        RECT  4.2825 5.6075 4.405 5.69 ;
        RECT  4.405 5.6275 4.54 5.695 ;
        RECT  4.1525 4.985 4.2175 5.76 ;
        RECT  2.5325 5.185 2.8225 5.25 ;
        RECT  1.995 5.37 2.1625 5.435 ;
        RECT  1.5025 5.435 1.5725 5.6925 ;
        RECT  1.4375 5.185 1.8625 5.25 ;
        RECT  2.5325 5.37 2.8225 5.44 ;
        RECT  1.6925 5.0775 1.7675 5.25 ;
        RECT  2.5325 5.56 2.8225 5.625 ;
        RECT  1.3725 5.5625 1.445 5.6275 ;
        RECT  3.0525 5.37 3.1225 5.755 ;
        RECT  2.0825 5.6025 2.1975 5.6675 ;
        RECT  1.3075 4.985 1.3725 5.76 ;
        RECT  2.1625 4.985 2.2275 5.76 ;
        RECT  1.1525 5.125 1.21 5.19 ;
        RECT  1.3925 5.6925 1.515 5.7575 ;
        RECT  4.955 5.51 5.1225 5.575 ;
        RECT  4.3475 5.445 4.45 5.5125 ;
        RECT  8.575 8.73 8.64 8.865 ;
        RECT  8.365 10.165 8.43 10.3 ;
        RECT  8.155 14.11 8.22 14.245 ;
        RECT  7.945 15.545 8.01 15.68 ;
        RECT  10.395 3.6 10.46 3.735 ;
        RECT  9.975 1.415 10.04 1.55 ;
        RECT  10.185 2.9625 10.25 3.0975 ;
        RECT  10.395 41.1 10.46 41.235 ;
        RECT  10.605 10.1025 10.67 10.2375 ;
        RECT  10.815 14.1275 10.88 14.2625 ;
        RECT  1.0125 7.63 1.1475 7.695 ;
        RECT  9.765 41.53 9.83 41.665 ;
        RECT  8.9225 40.545 9.1275 40.68 ;
        RECT  11.8025 40.5475 11.9375 40.6125 ;
        RECT  12.5075 40.5475 12.6425 40.6125 ;
        RECT  11.0275 40.5475 11.1625 40.6125 ;
        RECT  9.4175 0.355 9.6225 0.49 ;
        RECT  11.835 0.355 11.9 0.49 ;
        RECT  11.835 0.355 11.9 0.49 ;
        RECT  7.7875 21.555 7.9225 21.62 ;
        RECT  7.7875 24.245 7.9225 24.31 ;
        RECT  7.7875 26.935 7.9225 27.0 ;
        RECT  7.7875 29.625 7.9225 29.69 ;
        RECT  7.7875 32.315 7.9225 32.38 ;
        RECT  7.7875 35.005 7.9225 35.07 ;
        RECT  7.7875 37.695 7.9225 37.76 ;
        RECT  7.7875 40.385 7.9225 40.45 ;
        RECT  8.9225 13.4125 9.1275 13.5475 ;
        RECT  8.9225 18.7925 9.1275 18.9275 ;
        RECT  7.3125 7.81 7.4475 7.875 ;
        RECT  8.9225 7.8075 9.1275 7.9425 ;
        RECT  7.3125 6.4 7.4475 6.465 ;
        RECT  8.9225 6.3975 9.1275 6.5325 ;
        RECT  7.3125 6.4 7.4475 6.465 ;
        RECT  8.9225 6.3975 9.1275 6.5325 ;
        RECT  7.3125 4.99 7.4475 5.055 ;
        RECT  8.9225 4.9875 9.1275 5.1225 ;
        RECT  -2.49 17.335 -2.3225 17.4 ;
        RECT  -3.7575 17.335 -3.59 17.4 ;
        RECT  -3.9975 14.715 -3.9325 15.205 ;
        RECT  -4.1525 14.715 -4.0875 15.415 ;
        RECT  -5.5625 14.715 -5.4975 15.625 ;
        RECT  -4.5475 14.715 -4.4825 15.835 ;
        RECT  -1.325 15.345 -1.26 16.185 ;
        RECT  -0.795 15.975 -0.73 16.185 ;
        RECT  -2.12 15.975 -2.055 16.185 ;
        RECT  -2.6425 15.345 -2.5775 16.185 ;
        RECT  -2.7825 15.555 -2.7175 16.185 ;
        RECT  -4.025 15.975 -3.96 16.185 ;
        RECT  -3.5025 15.765 -3.4375 16.185 ;
        RECT  -3.3625 15.555 -3.2975 16.185 ;
        RECT  -0.9975 9.745 -0.9325 9.885 ;
        RECT  -0.22 9.885 -0.155 15.17 ;
        RECT  -0.965 14.7525 -0.9 14.8175 ;
        RECT  -0.795 14.7525 -0.73 14.8175 ;
        RECT  -0.965 14.715 -0.9 14.785 ;
        RECT  -0.9325 14.7525 -0.7625 14.8175 ;
        RECT  -0.795 14.785 -0.73 16.185 ;
        RECT  -2.49 17.895 -2.425 19.505 ;
        RECT  -3.655 19.015 -3.59 19.295 ;
        RECT  -0.965 18.455 -0.9 19.715 ;
        RECT  -0.205 19.47 -0.14 23.825 ;
        RECT  -0.385 23.7925 -0.14 23.8575 ;
        RECT  -1.7275 8.415 -1.6625 20.065 ;
        RECT  -4.4175 17.335 -4.3525 19.925 ;
        RECT  -5.73 14.4425 -1.6625 14.5075 ;
        RECT  -0.3825 8.415 -0.3175 20.835 ;
        RECT  -3.0725 17.335 -3.0075 20.76 ;
        RECT  -0.965 13.445 -0.9 13.585 ;
        RECT  -2.085 8.275 -2.02 13.445 ;
        RECT  -5.3775 8.4775 -2.0525 8.5425 ;
        RECT  -0.965 13.2025 -0.9 13.2675 ;
        RECT  -0.8675 13.2025 -0.8025 13.2675 ;
        RECT  -0.965 13.235 -0.9 13.445 ;
        RECT  -0.9325 13.2025 -0.835 13.2675 ;
        RECT  -0.8675 9.745 -0.8025 13.235 ;
        RECT  -5.73 8.4475 -3.615 8.5125 ;
        RECT  -5.73 14.445 -3.615 14.51 ;
        RECT  -5.19 10.965 -5.125 11.1 ;
        RECT  -5.375 10.965 -5.31 11.1 ;
        RECT  -5.19 9.73 -5.125 9.865 ;
        RECT  -5.375 9.73 -5.31 9.865 ;
        RECT  -5.38 10.965 -5.315 11.1 ;
        RECT  -5.565 10.965 -5.5 11.1 ;
        RECT  -5.38 13.925 -5.315 14.06 ;
        RECT  -5.565 13.925 -5.5 14.06 ;
        RECT  -5.38 9.73 -5.315 9.865 ;
        RECT  -5.565 9.73 -5.5 9.865 ;
        RECT  -5.19 13.925 -5.125 14.06 ;
        RECT  -5.375 13.925 -5.31 14.06 ;
        RECT  -5.38 9.195 -5.315 9.33 ;
        RECT  -5.565 9.195 -5.5 9.33 ;
        RECT  -5.24 12.155 -5.175 12.29 ;
        RECT  -5.425 12.155 -5.36 12.29 ;
        RECT  -5.19 12.69 -5.125 12.825 ;
        RECT  -5.375 12.69 -5.31 12.825 ;
        RECT  -5.38 12.69 -5.315 12.825 ;
        RECT  -5.565 12.69 -5.5 12.825 ;
        RECT  -5.19 13.115 -5.125 13.25 ;
        RECT  -5.375 13.115 -5.31 13.25 ;
        RECT  -5.19 10.155 -5.125 10.29 ;
        RECT  -5.375 10.155 -5.31 10.29 ;
        RECT  -5.19 13.5 -5.125 13.635 ;
        RECT  -5.375 13.5 -5.31 13.635 ;
        RECT  -5.38 13.5 -5.315 13.635 ;
        RECT  -5.565 13.5 -5.5 13.635 ;
        RECT  -5.38 10.155 -5.315 10.29 ;
        RECT  -5.565 10.155 -5.5 10.29 ;
        RECT  -5.38 13.115 -5.315 13.25 ;
        RECT  -5.565 13.115 -5.5 13.25 ;
        RECT  -5.38 10.54 -5.315 10.675 ;
        RECT  -5.565 10.54 -5.5 10.675 ;
        RECT  -5.19 10.54 -5.125 10.675 ;
        RECT  -5.375 10.54 -5.31 10.675 ;
        RECT  -5.38 8.77 -5.315 8.905 ;
        RECT  -5.565 8.77 -5.5 8.905 ;
        RECT  -5.305 11.745 -5.24 11.88 ;
        RECT  -5.49 11.745 -5.425 11.88 ;
        RECT  -5.5025 8.48 -5.3675 8.545 ;
        RECT  -5.565 13.9775 -5.5 14.1125 ;
        RECT  -5.675 12.1625 -5.61 12.2975 ;
        RECT  -5.565 11.2625 -5.5 11.3975 ;
        RECT  -5.1425 11.7375 -5.0775 11.8725 ;
        RECT  -5.565 14.3425 -5.5 14.4775 ;
        RECT  -5.0575 8.8 -4.9925 8.935 ;
        RECT  -5.2 12.8825 -5.135 13.0175 ;
        RECT  -5.1975 11.275 -5.1325 11.41 ;
        RECT  -5.1975 9.8775 -5.1325 10.0125 ;
        RECT  -5.7625 8.66 -5.6975 8.795 ;
        RECT  -5.1875 8.7775 -5.1225 8.9125 ;
        RECT  -5.1875 10.3875 -5.0525 10.4525 ;
        RECT  -5.1475 9.3025 -5.0825 9.4375 ;
        RECT  -5.1875 13.3475 -5.0525 13.4125 ;
        RECT  -5.24 14.235 -5.175 14.37 ;
        RECT  -5.32 10.765 -5.255 10.9 ;
        RECT  -5.33 13.725 -5.265 13.86 ;
        RECT  -5.5625 12.035 -5.4275 12.1 ;
        RECT  -5.0575 11.7375 -4.9925 11.8725 ;
        RECT  -5.6725 9.03 -5.5375 9.095 ;
        RECT  -5.5625 10.5425 -5.4975 10.6775 ;
        RECT  -5.1975 14.235 -5.1325 14.37 ;
        RECT  -5.375 13.725 -5.31 13.86 ;
        RECT  -5.0575 13.3125 -4.9925 13.4475 ;
        RECT  -5.0575 8.61 -4.9925 8.745 ;
        RECT  -5.1975 11.275 -5.1325 11.41 ;
        RECT  -5.0575 10.3525 -4.9925 10.4875 ;
        RECT  -5.5625 10.1525 -5.4975 10.2875 ;
        RECT  -5.375 10.1525 -5.31 10.2875 ;
        RECT  -5.375 10.765 -5.31 10.9 ;
        RECT  -5.565 13.1125 -5.5 13.2475 ;
        RECT  -5.375 13.1125 -5.31 13.2475 ;
        RECT  -5.765 8.48 -4.99 8.545 ;
        RECT  -5.695 11.55 -5.63 14.445 ;
        RECT  -5.19 14.06 -5.125 14.37 ;
        RECT  -5.565 13.635 -5.5 13.925 ;
        RECT  -5.565 12.825 -5.5 13.115 ;
        RECT  -5.425 14.4475 -5.3525 14.51 ;
        RECT  -5.38 14.06 -5.31 14.445 ;
        RECT  -5.38 12.825 -5.31 13.115 ;
        RECT  -5.38 13.345 -5.31 13.5025 ;
        RECT  -5.19 13.635 -5.125 13.925 ;
        RECT  -5.19 12.825 -5.125 13.115 ;
        RECT  -5.38 13.345 -4.995 13.415 ;
        RECT  -5.765 14.445 -4.99 14.51 ;
        RECT  -5.765 12.455 -4.99 12.52 ;
        RECT  -5.695 9.56 -5.63 11.485 ;
        RECT  -5.19 11.1 -5.125 11.41 ;
        RECT  -5.565 10.675 -5.5 10.965 ;
        RECT  -5.49 11.84 -5.425 12.29 ;
        RECT  -5.38 11.1 -5.31 11.485 ;
        RECT  -5.38 10.385 -5.31 10.5425 ;
        RECT  -5.565 11.3975 -5.5 11.485 ;
        RECT  -5.19 10.675 -5.125 10.965 ;
        RECT  -5.305 11.615 -5.06 11.68 ;
        RECT  -5.1425 11.615 -5.06 11.7375 ;
        RECT  -5.1225 11.7375 -5.055 11.8725 ;
        RECT  -5.765 11.485 -4.99 11.55 ;
        RECT  -5.565 9.865 -5.5 10.155 ;
        RECT  -5.38 9.3275 -5.315 9.495 ;
        RECT  -5.315 8.835 -5.0575 8.905 ;
        RECT  -5.565 8.77 -5.5 9.195 ;
        RECT  -5.38 9.865 -5.31 10.155 ;
        RECT  -5.6725 9.025 -5.5 9.1 ;
        RECT  -5.19 9.865 -5.125 10.155 ;
        RECT  -5.1875 8.705 -5.1225 8.7775 ;
        RECT  -5.38 10.385 -4.995 10.455 ;
        RECT  -5.1475 9.415 -5.0825 9.53 ;
        RECT  -5.765 8.64 -4.99 8.705 ;
        RECT  -5.765 9.495 -4.99 9.56 ;
        RECT  -5.625 8.485 -5.56 8.5425 ;
        RECT  -5.0575 8.725 -4.9925 8.8475 ;
        RECT  -5.24 12.2875 -5.175 12.455 ;
        RECT  -5.305 11.68 -5.2375 11.7825 ;
        RECT  -4.925 10.965 -4.86 11.1 ;
        RECT  -4.74 10.965 -4.675 11.1 ;
        RECT  -4.925 9.73 -4.86 9.865 ;
        RECT  -4.74 9.73 -4.675 9.865 ;
        RECT  -4.735 10.965 -4.67 11.1 ;
        RECT  -4.55 10.965 -4.485 11.1 ;
        RECT  -4.735 13.925 -4.67 14.06 ;
        RECT  -4.55 13.925 -4.485 14.06 ;
        RECT  -4.735 9.73 -4.67 9.865 ;
        RECT  -4.55 9.73 -4.485 9.865 ;
        RECT  -4.925 13.925 -4.86 14.06 ;
        RECT  -4.74 13.925 -4.675 14.06 ;
        RECT  -4.735 9.195 -4.67 9.33 ;
        RECT  -4.55 9.195 -4.485 9.33 ;
        RECT  -4.875 12.155 -4.81 12.29 ;
        RECT  -4.69 12.155 -4.625 12.29 ;
        RECT  -4.925 12.69 -4.86 12.825 ;
        RECT  -4.74 12.69 -4.675 12.825 ;
        RECT  -4.735 12.69 -4.67 12.825 ;
        RECT  -4.55 12.69 -4.485 12.825 ;
        RECT  -4.925 13.115 -4.86 13.25 ;
        RECT  -4.74 13.115 -4.675 13.25 ;
        RECT  -4.925 10.155 -4.86 10.29 ;
        RECT  -4.74 10.155 -4.675 10.29 ;
        RECT  -4.925 13.5 -4.86 13.635 ;
        RECT  -4.74 13.5 -4.675 13.635 ;
        RECT  -4.735 13.5 -4.67 13.635 ;
        RECT  -4.55 13.5 -4.485 13.635 ;
        RECT  -4.735 10.155 -4.67 10.29 ;
        RECT  -4.55 10.155 -4.485 10.29 ;
        RECT  -4.735 13.115 -4.67 13.25 ;
        RECT  -4.55 13.115 -4.485 13.25 ;
        RECT  -4.735 10.54 -4.67 10.675 ;
        RECT  -4.55 10.54 -4.485 10.675 ;
        RECT  -4.925 10.54 -4.86 10.675 ;
        RECT  -4.74 10.54 -4.675 10.675 ;
        RECT  -4.735 8.77 -4.67 8.905 ;
        RECT  -4.55 8.77 -4.485 8.905 ;
        RECT  -4.81 11.745 -4.745 11.88 ;
        RECT  -4.625 11.745 -4.56 11.88 ;
        RECT  -4.6825 8.48 -4.5475 8.545 ;
        RECT  -4.55 13.9775 -4.485 14.1125 ;
        RECT  -4.44 12.1625 -4.375 12.2975 ;
        RECT  -4.55 11.2625 -4.485 11.3975 ;
        RECT  -4.9725 11.7375 -4.9075 11.8725 ;
        RECT  -4.55 14.3425 -4.485 14.4775 ;
        RECT  -5.0575 8.8 -4.9925 8.935 ;
        RECT  -4.915 12.8825 -4.85 13.0175 ;
        RECT  -4.9175 11.275 -4.8525 11.41 ;
        RECT  -4.9175 9.8775 -4.8525 10.0125 ;
        RECT  -4.3525 8.66 -4.2875 8.795 ;
        RECT  -4.9275 8.7775 -4.8625 8.9125 ;
        RECT  -4.9975 10.3875 -4.8625 10.4525 ;
        RECT  -4.9675 9.3025 -4.9025 9.4375 ;
        RECT  -4.9975 13.3475 -4.8625 13.4125 ;
        RECT  -4.875 14.235 -4.81 14.37 ;
        RECT  -4.795 10.765 -4.73 10.9 ;
        RECT  -4.785 13.725 -4.72 13.86 ;
        RECT  -4.6225 12.035 -4.4875 12.1 ;
        RECT  -5.0575 11.7375 -4.9925 11.8725 ;
        RECT  -4.5125 9.03 -4.3775 9.095 ;
        RECT  -4.5525 10.5425 -4.4875 10.6775 ;
        RECT  -4.9175 14.235 -4.8525 14.37 ;
        RECT  -4.74 13.725 -4.675 13.86 ;
        RECT  -5.0575 13.3125 -4.9925 13.4475 ;
        RECT  -5.0575 8.61 -4.9925 8.745 ;
        RECT  -4.9175 11.275 -4.8525 11.41 ;
        RECT  -5.0575 10.3525 -4.9925 10.4875 ;
        RECT  -4.5525 10.1525 -4.4875 10.2875 ;
        RECT  -4.74 10.1525 -4.675 10.2875 ;
        RECT  -4.74 10.765 -4.675 10.9 ;
        RECT  -4.55 13.1125 -4.485 13.2475 ;
        RECT  -4.74 13.1125 -4.675 13.2475 ;
        RECT  -5.06 8.48 -4.285 8.545 ;
        RECT  -4.42 11.55 -4.355 14.445 ;
        RECT  -4.925 14.06 -4.86 14.37 ;
        RECT  -4.55 13.635 -4.485 13.925 ;
        RECT  -4.55 12.825 -4.485 13.115 ;
        RECT  -4.6975 14.4475 -4.625 14.51 ;
        RECT  -4.74 14.06 -4.67 14.445 ;
        RECT  -4.74 12.825 -4.67 13.115 ;
        RECT  -4.74 13.345 -4.67 13.5025 ;
        RECT  -4.925 13.635 -4.86 13.925 ;
        RECT  -4.925 12.825 -4.86 13.115 ;
        RECT  -5.055 13.345 -4.67 13.415 ;
        RECT  -5.06 14.445 -4.285 14.51 ;
        RECT  -5.06 12.455 -4.285 12.52 ;
        RECT  -4.42 9.56 -4.355 11.485 ;
        RECT  -4.925 11.1 -4.86 11.41 ;
        RECT  -4.55 10.675 -4.485 10.965 ;
        RECT  -4.625 11.84 -4.56 12.29 ;
        RECT  -4.74 11.1 -4.67 11.485 ;
        RECT  -4.74 10.385 -4.67 10.5425 ;
        RECT  -4.55 11.3975 -4.485 11.485 ;
        RECT  -4.925 10.675 -4.86 10.965 ;
        RECT  -4.99 11.615 -4.745 11.68 ;
        RECT  -4.99 11.615 -4.9075 11.7375 ;
        RECT  -4.995 11.7375 -4.9275 11.8725 ;
        RECT  -5.06 11.485 -4.285 11.55 ;
        RECT  -4.55 9.865 -4.485 10.155 ;
        RECT  -4.735 9.3275 -4.67 9.495 ;
        RECT  -4.9925 8.835 -4.735 8.905 ;
        RECT  -4.55 8.77 -4.485 9.195 ;
        RECT  -4.74 9.865 -4.67 10.155 ;
        RECT  -4.55 9.025 -4.3775 9.1 ;
        RECT  -4.925 9.865 -4.86 10.155 ;
        RECT  -4.9275 8.705 -4.8625 8.7775 ;
        RECT  -5.055 10.385 -4.67 10.455 ;
        RECT  -4.9675 9.415 -4.9025 9.53 ;
        RECT  -5.06 8.64 -4.285 8.705 ;
        RECT  -5.06 9.495 -4.285 9.56 ;
        RECT  -4.49 8.485 -4.425 8.5425 ;
        RECT  -5.0575 8.725 -4.9925 8.8475 ;
        RECT  -4.875 12.2875 -4.81 12.455 ;
        RECT  -4.8125 11.68 -4.745 11.7825 ;
        RECT  -3.78 10.965 -3.715 11.1 ;
        RECT  -3.965 10.965 -3.9 11.1 ;
        RECT  -3.78 9.73 -3.715 9.865 ;
        RECT  -3.965 9.73 -3.9 9.865 ;
        RECT  -3.97 10.965 -3.905 11.1 ;
        RECT  -4.155 10.965 -4.09 11.1 ;
        RECT  -3.97 13.925 -3.905 14.06 ;
        RECT  -4.155 13.925 -4.09 14.06 ;
        RECT  -3.97 9.73 -3.905 9.865 ;
        RECT  -4.155 9.73 -4.09 9.865 ;
        RECT  -3.78 13.925 -3.715 14.06 ;
        RECT  -3.965 13.925 -3.9 14.06 ;
        RECT  -3.97 9.195 -3.905 9.33 ;
        RECT  -4.155 9.195 -4.09 9.33 ;
        RECT  -3.83 12.155 -3.765 12.29 ;
        RECT  -4.015 12.155 -3.95 12.29 ;
        RECT  -3.78 12.69 -3.715 12.825 ;
        RECT  -3.965 12.69 -3.9 12.825 ;
        RECT  -3.97 12.69 -3.905 12.825 ;
        RECT  -4.155 12.69 -4.09 12.825 ;
        RECT  -3.78 13.115 -3.715 13.25 ;
        RECT  -3.965 13.115 -3.9 13.25 ;
        RECT  -3.78 10.155 -3.715 10.29 ;
        RECT  -3.965 10.155 -3.9 10.29 ;
        RECT  -3.78 13.5 -3.715 13.635 ;
        RECT  -3.965 13.5 -3.9 13.635 ;
        RECT  -3.97 13.5 -3.905 13.635 ;
        RECT  -4.155 13.5 -4.09 13.635 ;
        RECT  -3.97 10.155 -3.905 10.29 ;
        RECT  -4.155 10.155 -4.09 10.29 ;
        RECT  -3.97 13.115 -3.905 13.25 ;
        RECT  -4.155 13.115 -4.09 13.25 ;
        RECT  -3.97 10.54 -3.905 10.675 ;
        RECT  -4.155 10.54 -4.09 10.675 ;
        RECT  -3.78 10.54 -3.715 10.675 ;
        RECT  -3.965 10.54 -3.9 10.675 ;
        RECT  -3.97 8.77 -3.905 8.905 ;
        RECT  -4.155 8.77 -4.09 8.905 ;
        RECT  -3.895 11.745 -3.83 11.88 ;
        RECT  -4.08 11.745 -4.015 11.88 ;
        RECT  -4.0925 8.48 -3.9575 8.545 ;
        RECT  -4.155 13.9775 -4.09 14.1125 ;
        RECT  -4.265 12.1625 -4.2 12.2975 ;
        RECT  -4.155 11.2625 -4.09 11.3975 ;
        RECT  -3.7325 11.7375 -3.6675 11.8725 ;
        RECT  -4.155 14.3425 -4.09 14.4775 ;
        RECT  -3.6475 8.8 -3.5825 8.935 ;
        RECT  -3.79 12.8825 -3.725 13.0175 ;
        RECT  -3.7875 11.275 -3.7225 11.41 ;
        RECT  -3.7875 9.8775 -3.7225 10.0125 ;
        RECT  -4.3525 8.66 -4.2875 8.795 ;
        RECT  -3.7775 8.7775 -3.7125 8.9125 ;
        RECT  -3.7775 10.3875 -3.6425 10.4525 ;
        RECT  -3.7375 9.3025 -3.6725 9.4375 ;
        RECT  -3.7775 13.3475 -3.6425 13.4125 ;
        RECT  -3.83 14.235 -3.765 14.37 ;
        RECT  -3.91 10.765 -3.845 10.9 ;
        RECT  -3.92 13.725 -3.855 13.86 ;
        RECT  -4.1525 12.035 -4.0175 12.1 ;
        RECT  -3.6475 11.7375 -3.5825 11.8725 ;
        RECT  -4.2625 9.03 -4.1275 9.095 ;
        RECT  -4.1525 10.5425 -4.0875 10.6775 ;
        RECT  -3.7875 14.235 -3.7225 14.37 ;
        RECT  -3.965 13.725 -3.9 13.86 ;
        RECT  -3.6475 13.3125 -3.5825 13.4475 ;
        RECT  -3.6475 8.61 -3.5825 8.745 ;
        RECT  -3.7875 11.275 -3.7225 11.41 ;
        RECT  -3.6475 10.3525 -3.5825 10.4875 ;
        RECT  -4.1525 10.1525 -4.0875 10.2875 ;
        RECT  -3.965 10.1525 -3.9 10.2875 ;
        RECT  -3.965 10.765 -3.9 10.9 ;
        RECT  -4.155 13.1125 -4.09 13.2475 ;
        RECT  -3.965 13.1125 -3.9 13.2475 ;
        RECT  -4.355 8.48 -3.58 8.545 ;
        RECT  -4.285 11.55 -4.22 14.445 ;
        RECT  -3.78 14.06 -3.715 14.37 ;
        RECT  -4.155 13.635 -4.09 13.925 ;
        RECT  -4.155 12.825 -4.09 13.115 ;
        RECT  -4.015 14.4475 -3.9425 14.51 ;
        RECT  -3.97 14.06 -3.9 14.445 ;
        RECT  -3.97 12.825 -3.9 13.115 ;
        RECT  -3.97 13.345 -3.9 13.5025 ;
        RECT  -3.78 13.635 -3.715 13.925 ;
        RECT  -3.78 12.825 -3.715 13.115 ;
        RECT  -3.97 13.345 -3.585 13.415 ;
        RECT  -4.355 14.445 -3.58 14.51 ;
        RECT  -4.355 12.455 -3.58 12.52 ;
        RECT  -4.285 9.56 -4.22 11.485 ;
        RECT  -3.78 11.1 -3.715 11.41 ;
        RECT  -4.155 10.675 -4.09 10.965 ;
        RECT  -4.08 11.84 -4.015 12.29 ;
        RECT  -3.97 11.1 -3.9 11.485 ;
        RECT  -3.97 10.385 -3.9 10.5425 ;
        RECT  -4.155 11.3975 -4.09 11.485 ;
        RECT  -3.78 10.675 -3.715 10.965 ;
        RECT  -3.895 11.615 -3.65 11.68 ;
        RECT  -3.7325 11.615 -3.65 11.7375 ;
        RECT  -3.7125 11.7375 -3.645 11.8725 ;
        RECT  -4.355 11.485 -3.58 11.55 ;
        RECT  -4.155 9.865 -4.09 10.155 ;
        RECT  -3.97 9.3275 -3.905 9.495 ;
        RECT  -3.905 8.835 -3.6475 8.905 ;
        RECT  -4.155 8.77 -4.09 9.195 ;
        RECT  -3.97 9.865 -3.9 10.155 ;
        RECT  -4.2625 9.025 -4.09 9.1 ;
        RECT  -3.78 9.865 -3.715 10.155 ;
        RECT  -3.7775 8.705 -3.7125 8.7775 ;
        RECT  -3.97 10.385 -3.585 10.455 ;
        RECT  -3.7375 9.415 -3.6725 9.53 ;
        RECT  -4.355 8.64 -3.58 8.705 ;
        RECT  -4.355 9.495 -3.58 9.56 ;
        RECT  -4.215 8.485 -4.15 8.5425 ;
        RECT  -3.6475 8.725 -3.5825 8.8475 ;
        RECT  -3.83 12.2875 -3.765 12.455 ;
        RECT  -3.895 11.68 -3.8275 11.7825 ;
        RECT  -0.3825 13.585 -0.3175 14.715 ;
        RECT  -1.7275 13.585 -1.6625 14.715 ;
        RECT  -1.6625 14.5825 -1.2975 14.6475 ;
        RECT  -0.5175 14.5825 -0.3825 14.6475 ;
        RECT  -1.4325 13.8425 -0.485 13.9075 ;
        RECT  -1.4325 14.2225 -0.485 14.2875 ;
        RECT  -0.965 13.585 -0.9 13.62 ;
        RECT  -0.965 14.2875 -0.9 14.715 ;
        RECT  -0.385 13.6525 -0.32 13.7175 ;
        RECT  -0.385 14.0325 -0.32 14.0975 ;
        RECT  -0.385 14.0325 -0.32 14.0975 ;
        RECT  -0.385 14.4125 -0.32 14.4775 ;
        RECT  -0.5875 13.6525 -0.3875 13.7175 ;
        RECT  -0.3875 13.6525 -0.3525 13.7175 ;
        RECT  -0.385 13.685 -0.32 14.065 ;
        RECT  -0.5875 14.0325 -0.3525 14.0975 ;
        RECT  -0.5875 14.0325 -0.3875 14.0975 ;
        RECT  -0.3875 14.0325 -0.3525 14.0975 ;
        RECT  -0.385 14.065 -0.32 14.445 ;
        RECT  -0.5875 14.4125 -0.3525 14.4775 ;
        RECT  -0.7175 13.8425 -0.6525 13.9075 ;
        RECT  -0.7175 14.2225 -0.6525 14.2875 ;
        RECT  -0.6525 13.8425 -0.5875 13.9075 ;
        RECT  -0.685 13.8425 -0.6525 13.9075 ;
        RECT  -0.7175 13.875 -0.6525 14.255 ;
        RECT  -0.685 14.2225 -0.5875 14.2875 ;
        RECT  -0.7225 13.6525 -0.5875 13.7175 ;
        RECT  -0.7225 13.8425 -0.5875 13.9075 ;
        RECT  -0.7225 14.0325 -0.5875 14.0975 ;
        RECT  -0.7225 14.2225 -0.5875 14.2875 ;
        RECT  -0.7225 14.4125 -0.5875 14.4775 ;
        RECT  -1.705 13.6525 -1.64 13.7175 ;
        RECT  -1.705 14.0325 -1.64 14.0975 ;
        RECT  -1.705 14.0325 -1.64 14.0975 ;
        RECT  -1.705 14.4125 -1.64 14.4775 ;
        RECT  -1.6375 13.6525 -1.3675 13.7175 ;
        RECT  -1.6725 13.6525 -1.6375 13.7175 ;
        RECT  -1.705 13.685 -1.64 14.065 ;
        RECT  -1.6725 14.0325 -1.3675 14.0975 ;
        RECT  -1.6375 14.0325 -1.3675 14.0975 ;
        RECT  -1.6725 14.0325 -1.6375 14.0975 ;
        RECT  -1.705 14.065 -1.64 14.445 ;
        RECT  -1.6725 14.4125 -1.3675 14.4775 ;
        RECT  -1.2325 13.8425 -1.1675 13.9075 ;
        RECT  -1.2325 14.2225 -1.1675 14.2875 ;
        RECT  -1.3675 13.8425 -1.2325 13.9075 ;
        RECT  -1.2325 13.8425 -1.2 13.9075 ;
        RECT  -1.2325 13.875 -1.1675 14.255 ;
        RECT  -1.3675 14.2225 -1.2 14.2875 ;
        RECT  -1.5725 13.6525 -1.2975 13.7175 ;
        RECT  -1.5725 13.8425 -1.2975 13.9075 ;
        RECT  -1.5725 14.0325 -1.2975 14.0975 ;
        RECT  -1.5725 14.2225 -1.2975 14.2875 ;
        RECT  -1.5725 14.4125 -1.2975 14.4775 ;
        RECT  -1.5725 14.5825 -1.2975 14.6475 ;
        RECT  -0.5875 14.5825 -0.4525 14.6475 ;
        RECT  -0.965 13.62 -0.9 13.755 ;
        RECT  -0.3825 8.415 -0.3175 9.745 ;
        RECT  -1.7275 8.415 -1.6625 9.745 ;
        RECT  -0.8675 9.575 -0.8025 9.745 ;
        RECT  -0.9975 8.995 -0.9325 9.745 ;
        RECT  -0.8675 9.4225 -0.8025 9.4875 ;
        RECT  -0.8675 8.415 -0.8025 9.455 ;
        RECT  -0.835 9.4225 -0.4525 9.4875 ;
        RECT  -0.8675 8.415 -0.8025 8.875 ;
        RECT  -1.695 8.4825 -1.4125 8.5475 ;
        RECT  -0.4525 9.0625 -0.35 9.1275 ;
        RECT  -1.6625 9.6125 -1.4125 9.6775 ;
        RECT  -1.1275 9.4225 -1.0625 9.4875 ;
        RECT  -1.4125 9.4225 -1.095 9.4875 ;
        RECT  -1.1275 9.165 -1.0625 9.455 ;
        RECT  -1.6625 9.2325 -1.4125 9.2975 ;
        RECT  -1.1275 9.0325 -1.0625 9.0975 ;
        RECT  -1.4125 9.0325 -1.095 9.0975 ;
        RECT  -1.1275 9.065 -1.0625 9.165 ;
        RECT  -1.1275 8.6525 -1.0625 8.7175 ;
        RECT  -1.4125 8.6525 -1.095 8.7175 ;
        RECT  -1.1275 8.685 -1.0625 9.165 ;
        RECT  -0.4525 9.6125 -0.3175 9.6775 ;
        RECT  -0.4525 9.2325 -0.3175 9.2975 ;
        RECT  -0.6525 9.6125 -0.5175 9.6775 ;
        RECT  -0.6525 9.4225 -0.5175 9.4875 ;
        RECT  -0.6525 9.4225 -0.5175 9.4875 ;
        RECT  -0.6525 9.2325 -0.5175 9.2975 ;
        RECT  -1.2575 9.6125 -1.1225 9.6775 ;
        RECT  -1.2575 9.4225 -1.1225 9.4875 ;
        RECT  -1.2575 9.2325 -1.1225 9.2975 ;
        RECT  -1.2575 9.0325 -1.1225 9.0975 ;
        RECT  -1.2575 8.8425 -1.1225 8.9075 ;
        RECT  -1.2575 8.6525 -1.1225 8.7175 ;
        RECT  -1.4125 8.4825 -1.2775 8.5475 ;
        RECT  -0.4525 9.0625 -0.3175 9.1275 ;
        RECT  -0.7925 9.575 -0.7275 9.71 ;
        RECT  -0.9225 8.995 -0.8575 9.13 ;
        RECT  -1.4125 8.8425 -1.2775 8.9075 ;
        RECT  -0.7975 8.8075 -0.7325 8.9425 ;
        RECT  -0.3825 16.185 -0.3175 16.935 ;
        RECT  -1.7275 16.185 -1.6625 16.935 ;
        RECT  -1.695 16.8025 -1.4125 16.8675 ;
        RECT  -0.53 16.8025 -0.35 16.8675 ;
        RECT  -1.695 16.2525 -1.4125 16.3175 ;
        RECT  -1.695 16.6325 -1.4125 16.6975 ;
        RECT  -0.6325 16.2525 -0.35 16.3175 ;
        RECT  -1.31 16.665 -1.245 16.73 ;
        RECT  -1.31 16.4425 -1.245 16.5075 ;
        RECT  -1.2775 16.665 -0.4975 16.73 ;
        RECT  -1.31 16.475 -1.245 16.6975 ;
        RECT  -1.4125 16.4425 -1.2775 16.5075 ;
        RECT  -1.325 16.185 -1.26 16.22 ;
        RECT  -0.795 16.185 -0.73 16.46 ;
        RECT  -1.0125 16.6975 -0.9475 16.935 ;
        RECT  -0.7675 16.2525 -0.6325 16.3175 ;
        RECT  -0.7675 16.4425 -0.6325 16.5075 ;
        RECT  -0.7675 16.4425 -0.6325 16.5075 ;
        RECT  -0.7675 16.6325 -0.6325 16.6975 ;
        RECT  -1.5475 16.2525 -1.4125 16.3175 ;
        RECT  -1.5475 16.4425 -1.4125 16.5075 ;
        RECT  -1.5475 16.4425 -1.4125 16.5075 ;
        RECT  -1.5475 16.6325 -1.4125 16.6975 ;
        RECT  -1.5475 16.8025 -1.4125 16.8675 ;
        RECT  -0.6325 16.8025 -0.4975 16.8675 ;
        RECT  -1.325 16.22 -1.26 16.355 ;
        RECT  -0.795 16.46 -0.73 16.595 ;
        RECT  -1.98 21.28 -1.91 21.415 ;
        RECT  -1.0 23.7925 -0.935 23.8575 ;
        RECT  -0.9675 23.7925 -0.385 23.8575 ;
        RECT  -1.0 23.825 -0.935 23.965 ;
        RECT  -1.3825 21.1725 -1.3175 21.3125 ;
        RECT  -2.1375 21.1725 -2.0725 21.2 ;
        RECT  -2.1375 21.1675 -2.0725 21.2325 ;
        RECT  -4.38 21.1675 -2.105 21.2325 ;
        RECT  -2.525 23.5125 -0.6175 23.5775 ;
        RECT  -4.195 22.6025 -3.9625 22.6675 ;
        RECT  -0.9425 22.0425 -0.8775 22.1075 ;
        RECT  -0.9425 21.6925 -0.8775 22.075 ;
        RECT  -1.35 22.0425 -0.91 22.1075 ;
        RECT  -3.705 22.0425 -1.35 22.1075 ;
        RECT  -0.9425 21.28 -0.8775 21.345 ;
        RECT  -0.9425 21.3125 -0.8775 21.5025 ;
        RECT  -1.35 21.28 -0.91 21.345 ;
        RECT  -4.905 26.2675 -0.385 26.3325 ;
        RECT  -1.7625 23.8025 -1.6975 23.8675 ;
        RECT  -1.7625 23.835 -1.6975 23.965 ;
        RECT  -3.705 23.8025 -1.73 23.8675 ;
        RECT  -3.705 23.8025 -1.73 23.8675 ;
        RECT  -1.35 20.6975 -0.385 20.7625 ;
        RECT  -3.075 25.1925 -0.385 25.2575 ;
        RECT  -0.4175 24.105 -0.3525 25.225 ;
        RECT  -3.1075 24.105 -3.0425 25.225 ;
        RECT  -3.495 23.965 -3.0425 24.03 ;
        RECT  -4.195 22.8825 -3.495 22.9475 ;
        RECT  -4.195 24.0875 -3.705 24.1525 ;
        RECT  -3.495 23.965 -3.0425 24.03 ;
        RECT  -4.195 25.2925 -3.495 25.3575 ;
        RECT  -4.5475 21.3975 -3.705 21.4625 ;
        RECT  -4.9 20.6975 -0.79 20.7625 ;
        RECT  -4.195 20.6975 -0.79 20.7625 ;
        RECT  -1.91 20.6975 -1.35 20.7625 ;
        RECT  -1.91 19.3525 -1.35 19.4175 ;
        RECT  -1.8425 19.4175 -1.7775 19.7825 ;
        RECT  -1.8425 20.5625 -1.7775 20.6975 ;
        RECT  -1.4825 20.6275 -1.4175 20.6975 ;
        RECT  -1.4825 19.4175 -1.4175 19.5075 ;
        RECT  -1.6725 19.6475 -1.6075 20.595 ;
        RECT  -1.385 20.115 -1.35 20.18 ;
        RECT  -1.91 20.115 -1.6725 20.18 ;
        RECT  -1.4825 20.3575 -1.4175 20.4925 ;
        RECT  -1.6725 20.3575 -1.6075 20.4925 ;
        RECT  -1.4825 19.5075 -1.4175 19.7825 ;
        RECT  -1.6725 19.5075 -1.6075 19.7825 ;
        RECT  -1.8425 19.5075 -1.7775 19.7825 ;
        RECT  -1.8425 20.4925 -1.7775 20.6275 ;
        RECT  -1.52 20.115 -1.385 20.18 ;
        RECT  -0.9425 21.27 -0.8075 21.335 ;
        RECT  -0.9425 21.08 -0.8075 21.145 ;
        RECT  -1.0025 23.83 -0.9375 23.965 ;
        RECT  -0.4175 23.405 -0.3525 23.965 ;
        RECT  -1.7625 23.405 -1.6975 23.965 ;
        RECT  -1.6975 23.4725 -1.3325 23.5375 ;
        RECT  -0.5525 23.4725 -0.4175 23.5375 ;
        RECT  -0.4875 23.8325 -0.4175 23.8975 ;
        RECT  -1.6975 23.8325 -1.6075 23.8975 ;
        RECT  -1.4675 23.6425 -0.52 23.7075 ;
        RECT  -1.0 23.93 -0.935 23.965 ;
        RECT  -0.6875 23.8325 -0.5525 23.8975 ;
        RECT  -0.6875 23.6425 -0.5525 23.7075 ;
        RECT  -1.2275 23.8325 -0.9525 23.8975 ;
        RECT  -1.2275 23.6425 -0.9525 23.7075 ;
        RECT  -1.3325 23.4725 -1.0575 23.5375 ;
        RECT  -0.4875 23.4725 -0.3525 23.5375 ;
        RECT  -0.925 23.795 -0.86 23.93 ;
        RECT  -1.0025 23.27 -0.9375 23.405 ;
        RECT  -0.4175 22.845 -0.3525 23.405 ;
        RECT  -1.7625 22.845 -1.6975 23.405 ;
        RECT  -1.6975 22.9125 -1.3325 22.9775 ;
        RECT  -0.5525 22.9125 -0.4175 22.9775 ;
        RECT  -0.4875 23.2725 -0.4175 23.3375 ;
        RECT  -1.6975 23.2725 -1.6075 23.3375 ;
        RECT  -1.4675 23.0825 -0.52 23.1475 ;
        RECT  -1.0 23.37 -0.935 23.405 ;
        RECT  -0.6875 23.2725 -0.5525 23.3375 ;
        RECT  -0.6875 23.0825 -0.5525 23.1475 ;
        RECT  -1.2275 23.2725 -0.9525 23.3375 ;
        RECT  -1.2275 23.0825 -0.9525 23.1475 ;
        RECT  -1.3325 22.9125 -1.0575 22.9775 ;
        RECT  -0.4875 22.9125 -0.3525 22.9775 ;
        RECT  -0.925 23.235 -0.86 23.37 ;
        RECT  -2.5225 22.845 -2.4575 22.98 ;
        RECT  -3.1075 22.845 -3.0425 23.405 ;
        RECT  -1.7625 22.845 -1.6975 23.405 ;
        RECT  -2.1275 23.2725 -1.7625 23.3375 ;
        RECT  -3.0425 23.2725 -2.9075 23.3375 ;
        RECT  -3.0425 22.9125 -2.9725 22.9775 ;
        RECT  -1.8525 22.9125 -1.7625 22.9775 ;
        RECT  -2.94 23.1025 -1.9925 23.1675 ;
        RECT  -2.525 22.845 -2.46 22.88 ;
        RECT  -2.9075 22.9125 -2.7725 22.9775 ;
        RECT  -2.9075 23.1025 -2.7725 23.1675 ;
        RECT  -2.5075 22.9125 -2.2325 22.9775 ;
        RECT  -2.5075 23.1025 -2.2325 23.1675 ;
        RECT  -2.4025 23.2725 -2.1275 23.3375 ;
        RECT  -3.1075 23.2725 -2.9725 23.3375 ;
        RECT  -2.6 22.88 -2.535 23.015 ;
        RECT  -2.5225 23.405 -2.4575 23.54 ;
        RECT  -3.1075 23.405 -3.0425 23.965 ;
        RECT  -1.7625 23.405 -1.6975 23.965 ;
        RECT  -2.1275 23.8325 -1.7625 23.8975 ;
        RECT  -3.0425 23.8325 -2.9075 23.8975 ;
        RECT  -3.0425 23.4725 -2.9725 23.5375 ;
        RECT  -1.8525 23.4725 -1.7625 23.5375 ;
        RECT  -2.94 23.6625 -1.9925 23.7275 ;
        RECT  -2.525 23.405 -2.46 23.44 ;
        RECT  -2.9075 23.4725 -2.7725 23.5375 ;
        RECT  -2.9075 23.6625 -2.7725 23.7275 ;
        RECT  -2.5075 23.4725 -2.2325 23.5375 ;
        RECT  -2.5075 23.6625 -2.2325 23.7275 ;
        RECT  -2.4025 23.8325 -2.1275 23.8975 ;
        RECT  -3.1075 23.8325 -2.9725 23.8975 ;
        RECT  -2.6 23.44 -2.535 23.575 ;
        RECT  -1.0025 23.5075 -0.9375 23.6425 ;
        RECT  -1.0025 22.9475 -0.9375 23.0825 ;
        RECT  -2.5225 23.1675 -2.4575 23.3025 ;
        RECT  -4.85 23.0325 -4.785 23.1675 ;
        RECT  -4.665 23.0325 -4.6 23.1675 ;
        RECT  -4.495 23.0375 -4.43 23.1725 ;
        RECT  -4.31 23.0375 -4.245 23.1725 ;
        RECT  -4.93 23.4225 -4.865 23.5575 ;
        RECT  -4.745 23.4225 -4.68 23.5575 ;
        RECT  -4.415 23.4225 -4.35 23.5575 ;
        RECT  -4.23 23.4225 -4.165 23.5575 ;
        RECT  -4.93 23.8875 -4.865 24.0225 ;
        RECT  -4.745 23.8875 -4.68 24.0225 ;
        RECT  -4.415 23.8875 -4.35 24.0225 ;
        RECT  -4.23 23.8875 -4.165 24.0225 ;
        RECT  -4.2275 23.0375 -4.1625 23.1725 ;
        RECT  -4.9325 23.5125 -4.8675 23.6475 ;
        RECT  -4.2275 23.5125 -4.1625 23.6475 ;
        RECT  -4.68 23.0325 -4.615 23.1675 ;
        RECT  -4.48 23.0375 -4.415 23.1725 ;
        RECT  -4.7275 23.6275 -4.5925 23.6925 ;
        RECT  -4.5025 23.7775 -4.3675 23.8425 ;
        RECT  -4.605 22.8825 -4.47 22.9475 ;
        RECT  -4.6125 24.0875 -4.4775 24.1525 ;
        RECT  -4.61 22.7425 -4.475 22.8075 ;
        RECT  -4.9675 22.7425 -4.8325 22.8075 ;
        RECT  -4.2475 23.0375 -4.195 23.1725 ;
        RECT  -4.2625 22.7425 -4.1275 22.8075 ;
        RECT  -4.5775 24.0875 -4.5125 24.1525 ;
        RECT  -4.23 22.8825 -4.16 22.9475 ;
        RECT  -4.785 23.2575 -4.68 23.3225 ;
        RECT  -4.745 23.3225 -4.68 23.4225 ;
        RECT  -4.85 23.1675 -4.785 23.3225 ;
        RECT  -4.415 23.2575 -4.31 23.3225 ;
        RECT  -4.415 23.3225 -4.35 23.4225 ;
        RECT  -4.31 23.1725 -4.245 23.3225 ;
        RECT  -4.93 24.0225 -4.865 24.0875 ;
        RECT  -4.23 24.0225 -4.165 24.0875 ;
        RECT  -4.745 23.4225 -4.68 23.9125 ;
        RECT  -4.415 23.4225 -4.35 23.9125 ;
        RECT  -4.99 22.8825 -4.105 22.9475 ;
        RECT  -4.99 24.0875 -4.105 24.1525 ;
        RECT  -4.99 22.7425 -4.105 22.8075 ;
        RECT  -4.93 21.5275 -4.865 21.6625 ;
        RECT  -4.745 21.5275 -4.68 21.6625 ;
        RECT  -4.23 21.5275 -4.165 21.6625 ;
        RECT  -4.415 21.5275 -4.35 21.6625 ;
        RECT  -4.745 21.9925 -4.68 22.1275 ;
        RECT  -4.93 21.9925 -4.865 22.1275 ;
        RECT  -4.415 21.9925 -4.35 22.1275 ;
        RECT  -4.23 21.9925 -4.165 22.1275 ;
        RECT  -4.85 22.3825 -4.785 22.5175 ;
        RECT  -4.665 22.3825 -4.6 22.5175 ;
        RECT  -4.495 22.3825 -4.43 22.5175 ;
        RECT  -4.31 22.3825 -4.245 22.5175 ;
        RECT  -4.9325 21.89 -4.8675 22.025 ;
        RECT  -4.9325 21.89 -4.8675 22.025 ;
        RECT  -4.9325 21.89 -4.8675 22.025 ;
        RECT  -4.9325 21.89 -4.8675 22.025 ;
        RECT  -4.9325 21.89 -4.8675 22.025 ;
        RECT  -4.9325 21.89 -4.8675 22.025 ;
        RECT  -4.61 21.3975 -4.475 21.4625 ;
        RECT  -4.2625 22.7425 -4.1275 22.8075 ;
        RECT  -4.9675 22.7425 -4.8325 22.8075 ;
        RECT  -4.5975 22.6025 -4.4625 22.6675 ;
        RECT  -4.9325 21.89 -4.8675 22.025 ;
        RECT  -4.9325 21.89 -4.8675 22.025 ;
        RECT  -4.9325 21.89 -4.8675 22.025 ;
        RECT  -4.9325 21.89 -4.8675 22.025 ;
        RECT  -4.5025 21.7125 -4.3675 21.7775 ;
        RECT  -4.5025 21.7125 -4.3675 21.7775 ;
        RECT  -4.7275 21.8625 -4.5925 21.9275 ;
        RECT  -4.7275 21.8625 -4.5925 21.9275 ;
        RECT  -4.9325 21.89 -4.8675 22.025 ;
        RECT  -4.9325 21.89 -4.8675 22.025 ;
        RECT  -4.9325 21.89 -4.8675 22.025 ;
        RECT  -4.9325 21.89 -4.8675 22.025 ;
        RECT  -4.4825 22.3825 -4.4175 22.5175 ;
        RECT  -4.2275 21.89 -4.1625 22.025 ;
        RECT  -4.2275 21.89 -4.1625 22.025 ;
        RECT  -4.2275 21.89 -4.1625 22.025 ;
        RECT  -4.2275 21.89 -4.1625 22.025 ;
        RECT  -4.2275 21.89 -4.1625 22.025 ;
        RECT  -4.2275 21.89 -4.1625 22.025 ;
        RECT  -4.9325 21.89 -4.8675 22.025 ;
        RECT  -4.9325 21.89 -4.8675 22.025 ;
        RECT  -4.9325 21.89 -4.8675 22.025 ;
        RECT  -4.9325 21.89 -4.8675 22.025 ;
        RECT  -4.6775 22.3825 -4.6125 22.5175 ;
        RECT  -4.615 22.7425 -4.48 22.8075 ;
        RECT  -4.615 22.7425 -4.48 22.8075 ;
        RECT  -4.9675 22.7425 -4.8325 22.8075 ;
        RECT  -4.61 21.3975 -4.475 21.4625 ;
        RECT  -4.9675 22.7425 -4.8325 22.8075 ;
        RECT  -4.9675 22.7425 -4.8325 22.8075 ;
        RECT  -4.9325 21.89 -4.8675 22.025 ;
        RECT  -4.9325 21.89 -4.8675 22.025 ;
        RECT  -4.9325 21.89 -4.8675 22.025 ;
        RECT  -4.9325 21.89 -4.8675 22.025 ;
        RECT  -4.9325 21.89 -4.8675 22.025 ;
        RECT  -4.9325 21.89 -4.8675 22.025 ;
        RECT  -4.2625 22.7425 -4.1275 22.8075 ;
        RECT  -4.5875 21.4 -4.4875 21.4625 ;
        RECT  -4.5875 21.3975 -4.4875 21.46 ;
        RECT  -4.8675 22.6025 -4.815 22.665 ;
        RECT  -4.5875 21.4 -4.4875 21.4625 ;
        RECT  -4.935 21.4625 -4.865 21.6625 ;
        RECT  -4.935 21.9925 -4.865 22.1275 ;
        RECT  -4.935 21.9925 -4.865 22.1275 ;
        RECT  -4.99 22.7425 -4.105 22.8075 ;
        RECT  -4.855 22.2275 -4.68 22.2925 ;
        RECT  -4.23 21.9925 -4.16 22.1275 ;
        RECT  -4.415 21.5525 -4.35 22.2925 ;
        RECT  -4.5875 21.3975 -4.4875 21.46 ;
        RECT  -4.1625 22.6025 -4.11 22.665 ;
        RECT  -4.935 21.9925 -4.865 22.1275 ;
        RECT  -4.99 21.3975 -4.105 21.4625 ;
        RECT  -4.745 21.6625 -4.68 22.2925 ;
        RECT  -4.935 21.9925 -4.865 22.1275 ;
        RECT  -4.935 21.9925 -4.865 22.1275 ;
        RECT  -4.315 22.2275 -4.245 22.5175 ;
        RECT  -4.23 21.9925 -4.16 22.1275 ;
        RECT  -4.99 22.6025 -4.105 22.6675 ;
        RECT  -4.935 21.9925 -4.865 22.1275 ;
        RECT  -4.935 21.4625 -4.865 21.6625 ;
        RECT  -4.23 21.4625 -4.16 21.6625 ;
        RECT  -4.855 22.2275 -4.785 22.5175 ;
        RECT  -4.415 22.2275 -4.245 22.2925 ;
        RECT  -4.93 21.1975 -4.865 21.3325 ;
        RECT  -4.745 21.1975 -4.68 21.3325 ;
        RECT  -4.23 21.1975 -4.165 21.3325 ;
        RECT  -4.415 21.1975 -4.35 21.3325 ;
        RECT  -4.745 20.7325 -4.68 20.8675 ;
        RECT  -4.93 20.7325 -4.865 20.8675 ;
        RECT  -4.415 20.7325 -4.35 20.8675 ;
        RECT  -4.23 20.7325 -4.165 20.8675 ;
        RECT  -4.85 20.3425 -4.785 20.4775 ;
        RECT  -4.665 20.3425 -4.6 20.4775 ;
        RECT  -4.495 20.3425 -4.43 20.4775 ;
        RECT  -4.31 20.3425 -4.245 20.4775 ;
        RECT  -4.9325 20.835 -4.8675 20.97 ;
        RECT  -4.9325 20.835 -4.8675 20.97 ;
        RECT  -4.9325 20.835 -4.8675 20.97 ;
        RECT  -4.9325 20.835 -4.8675 20.97 ;
        RECT  -4.9325 20.835 -4.8675 20.97 ;
        RECT  -4.9325 20.835 -4.8675 20.97 ;
        RECT  -4.61 21.3975 -4.475 21.4625 ;
        RECT  -4.2625 20.0525 -4.1275 20.1175 ;
        RECT  -4.9675 20.0525 -4.8325 20.1175 ;
        RECT  -4.5975 20.1925 -4.4625 20.2575 ;
        RECT  -4.9325 20.835 -4.8675 20.97 ;
        RECT  -4.9325 20.835 -4.8675 20.97 ;
        RECT  -4.9325 20.835 -4.8675 20.97 ;
        RECT  -4.9325 20.835 -4.8675 20.97 ;
        RECT  -4.5025 21.0825 -4.3675 21.1475 ;
        RECT  -4.5025 21.0825 -4.3675 21.1475 ;
        RECT  -4.7275 20.9325 -4.5925 20.9975 ;
        RECT  -4.7275 20.9325 -4.5925 20.9975 ;
        RECT  -4.9325 20.835 -4.8675 20.97 ;
        RECT  -4.9325 20.835 -4.8675 20.97 ;
        RECT  -4.9325 20.835 -4.8675 20.97 ;
        RECT  -4.9325 20.835 -4.8675 20.97 ;
        RECT  -4.4825 20.3425 -4.4175 20.4775 ;
        RECT  -4.2275 20.835 -4.1625 20.97 ;
        RECT  -4.2275 20.835 -4.1625 20.97 ;
        RECT  -4.2275 20.835 -4.1625 20.97 ;
        RECT  -4.2275 20.835 -4.1625 20.97 ;
        RECT  -4.2275 20.835 -4.1625 20.97 ;
        RECT  -4.2275 20.835 -4.1625 20.97 ;
        RECT  -4.9325 20.835 -4.8675 20.97 ;
        RECT  -4.9325 20.835 -4.8675 20.97 ;
        RECT  -4.9325 20.835 -4.8675 20.97 ;
        RECT  -4.9325 20.835 -4.8675 20.97 ;
        RECT  -4.6775 20.3425 -4.6125 20.4775 ;
        RECT  -4.615 20.0525 -4.48 20.1175 ;
        RECT  -4.615 20.0525 -4.48 20.1175 ;
        RECT  -4.9675 20.0525 -4.8325 20.1175 ;
        RECT  -4.61 21.3975 -4.475 21.4625 ;
        RECT  -4.9675 20.0525 -4.8325 20.1175 ;
        RECT  -4.9675 20.0525 -4.8325 20.1175 ;
        RECT  -4.9325 20.835 -4.8675 20.97 ;
        RECT  -4.9325 20.835 -4.8675 20.97 ;
        RECT  -4.9325 20.835 -4.8675 20.97 ;
        RECT  -4.9325 20.835 -4.8675 20.97 ;
        RECT  -4.9325 20.835 -4.8675 20.97 ;
        RECT  -4.9325 20.835 -4.8675 20.97 ;
        RECT  -4.2625 20.0525 -4.1275 20.1175 ;
        RECT  -4.5875 21.3975 -4.4875 21.46 ;
        RECT  -4.5875 21.4 -4.4875 21.4625 ;
        RECT  -4.8675 20.195 -4.815 20.2575 ;
        RECT  -4.5875 21.3975 -4.4875 21.46 ;
        RECT  -4.935 21.1975 -4.865 21.3975 ;
        RECT  -4.935 20.7325 -4.865 20.8675 ;
        RECT  -4.935 20.7325 -4.865 20.8675 ;
        RECT  -4.99 20.0525 -4.105 20.1175 ;
        RECT  -4.855 20.5675 -4.68 20.6325 ;
        RECT  -4.23 20.7325 -4.16 20.8675 ;
        RECT  -4.415 20.5675 -4.35 21.3075 ;
        RECT  -4.5875 21.4 -4.4875 21.4625 ;
        RECT  -4.1625 20.195 -4.11 20.2575 ;
        RECT  -4.935 20.7325 -4.865 20.8675 ;
        RECT  -4.99 21.3975 -4.105 21.4625 ;
        RECT  -4.745 20.5675 -4.68 21.1975 ;
        RECT  -4.935 20.7325 -4.865 20.8675 ;
        RECT  -4.935 20.7325 -4.865 20.8675 ;
        RECT  -4.315 20.3425 -4.245 20.6325 ;
        RECT  -4.23 20.7325 -4.16 20.8675 ;
        RECT  -4.99 20.1925 -4.105 20.2575 ;
        RECT  -4.935 20.7325 -4.865 20.8675 ;
        RECT  -4.935 21.1975 -4.865 21.3975 ;
        RECT  -4.23 21.1975 -4.16 21.3975 ;
        RECT  -4.855 20.3425 -4.785 20.6325 ;
        RECT  -4.415 20.5675 -4.245 20.6325 ;
        RECT  -1.9775 21.1775 -1.9125 21.3125 ;
        RECT  -1.4175 21.07 -1.2825 21.135 ;
        RECT  -2.1725 21.07 -2.0375 21.135 ;
        RECT  -4.4475 21.0975 -4.3125 21.1625 ;
        RECT  -0.655 21.395 -0.59 21.53 ;
        RECT  -0.685 23.4425 -0.55 23.5075 ;
        RECT  -2.5925 23.4425 -2.4575 23.5075 ;
        RECT  -2.5925 24.2025 -2.5275 24.3375 ;
        RECT  -0.65 21.365 -0.585 21.5 ;
        RECT  -4.0275 22.4325 -3.9625 22.5675 ;
        RECT  -3.7725 21.9725 -3.6375 22.0375 ;
        RECT  -3.7725 23.7325 -3.6375 23.7975 ;
        RECT  -0.4525 20.6275 -0.3175 20.6925 ;
        RECT  -0.4525 25.1225 -0.3175 25.1875 ;
        RECT  -3.1425 25.1225 -3.0075 25.1875 ;
        RECT  -3.7725 26.2675 -3.7075 26.4025 ;
        RECT  -3.5625 23.895 -3.4275 23.96 ;
        RECT  -3.5625 22.8125 -3.4275 22.8775 ;
        RECT  -3.7725 24.0175 -3.6375 24.0825 ;
        RECT  -3.5625 23.895 -3.4275 23.96 ;
        RECT  -3.5625 25.2225 -3.4275 25.2875 ;
        RECT  -3.7725 21.3275 -3.6375 21.3925 ;
        RECT  -4.9675 20.6275 -4.8325 20.6925 ;
        RECT  -4.2625 20.6275 -4.1275 20.6925 ;
        RECT  -0.3825 17.335 -0.3175 17.895 ;
        RECT  -1.7275 17.335 -1.6625 17.895 ;
        RECT  -1.6625 17.4025 -1.2975 17.4675 ;
        RECT  -0.5175 17.4025 -0.3825 17.4675 ;
        RECT  -0.4525 17.7625 -0.3825 17.8275 ;
        RECT  -1.6625 17.7625 -1.5725 17.8275 ;
        RECT  -1.4325 17.5725 -0.485 17.6375 ;
        RECT  -0.965 17.86 -0.9 17.895 ;
        RECT  -0.965 17.335 -0.9 17.5725 ;
        RECT  -0.6525 17.7625 -0.5175 17.8275 ;
        RECT  -0.6525 17.5725 -0.5175 17.6375 ;
        RECT  -1.1925 17.7625 -0.9175 17.8275 ;
        RECT  -1.1925 17.5725 -0.9175 17.6375 ;
        RECT  -1.2975 17.4025 -1.0225 17.4675 ;
        RECT  -0.4525 17.4025 -0.3175 17.4675 ;
        RECT  -0.89 17.725 -0.825 17.86 ;
        RECT  -0.3825 17.895 -0.3175 18.455 ;
        RECT  -1.7275 17.895 -1.6625 18.455 ;
        RECT  -1.6625 17.9625 -1.2975 18.0275 ;
        RECT  -0.5175 17.9625 -0.3825 18.0275 ;
        RECT  -0.4525 18.3225 -0.3825 18.3875 ;
        RECT  -1.6625 18.3225 -1.5725 18.3875 ;
        RECT  -1.4325 18.1325 -0.485 18.1975 ;
        RECT  -0.965 18.42 -0.9 18.455 ;
        RECT  -0.965 17.895 -0.9 18.1325 ;
        RECT  -0.6525 18.3225 -0.5175 18.3875 ;
        RECT  -0.6525 18.1325 -0.5175 18.1975 ;
        RECT  -1.1925 18.3225 -0.9175 18.3875 ;
        RECT  -1.1925 18.1325 -0.9175 18.1975 ;
        RECT  -1.2975 17.9625 -1.0225 18.0275 ;
        RECT  -0.4525 17.9625 -0.3175 18.0275 ;
        RECT  -0.89 18.285 -0.825 18.42 ;
        RECT  -3.0725 16.185 -3.0075 17.335 ;
        RECT  -1.7275 16.185 -1.6625 17.335 ;
        RECT  -2.91 17.02 -1.825 17.085 ;
        RECT  -1.9775 17.1575 -1.695 17.2225 ;
        RECT  -3.04 17.1575 -2.77 17.2225 ;
        RECT  -1.9775 16.4175 -1.695 16.4825 ;
        RECT  -1.9775 16.7975 -1.695 16.8625 ;
        RECT  -3.04 16.4175 -2.7575 16.4825 ;
        RECT  -2.12 16.185 -2.055 16.495 ;
        RECT  -2.6425 16.185 -2.5775 16.35 ;
        RECT  -2.7825 16.185 -2.7175 16.35 ;
        RECT  -2.3875 17.02 -2.3225 17.335 ;
        RECT  -2.8125 16.4175 -2.5375 16.4825 ;
        RECT  -2.8125 16.6075 -2.5375 16.6725 ;
        RECT  -2.8125 16.6075 -2.5375 16.6725 ;
        RECT  -2.8125 16.7975 -2.5375 16.8625 ;
        RECT  -2.8125 16.7975 -2.5375 16.8625 ;
        RECT  -2.8125 16.9875 -2.5375 17.0525 ;
        RECT  -2.2675 16.4175 -2.1325 16.4825 ;
        RECT  -2.2675 16.6075 -2.1325 16.6725 ;
        RECT  -2.2675 16.6075 -2.1325 16.6725 ;
        RECT  -2.2675 16.7975 -2.1325 16.8625 ;
        RECT  -2.2675 16.7975 -2.1325 16.8625 ;
        RECT  -2.2675 16.9875 -2.1325 17.0525 ;
        RECT  -2.1125 17.1575 -1.9775 17.2225 ;
        RECT  -3.1925 17.1575 -2.9175 17.2225 ;
        RECT  -2.1125 16.6075 -1.9775 16.6725 ;
        RECT  -2.1125 16.9875 -1.9775 17.0525 ;
        RECT  -2.2 16.36 -2.135 16.495 ;
        RECT  -2.7125 16.665 -2.5775 16.73 ;
        RECT  -2.7125 16.6625 -2.5775 16.7275 ;
        RECT  -2.715 16.215 -2.65 16.35 ;
        RECT  -2.7125 16.855 -2.5775 16.92 ;
        RECT  -2.7125 16.8525 -2.5775 16.9175 ;
        RECT  -2.855 16.215 -2.79 16.35 ;
        RECT  -3.0725 16.185 -3.0075 17.335 ;
        RECT  -4.4175 16.185 -4.3525 17.335 ;
        RECT  -4.255 17.02 -3.17 17.085 ;
        RECT  -4.385 17.1575 -4.1025 17.2225 ;
        RECT  -3.31 17.1575 -3.04 17.2225 ;
        RECT  -4.385 16.4175 -4.1025 16.4825 ;
        RECT  -4.385 16.7975 -4.1025 16.8625 ;
        RECT  -3.3225 16.4175 -3.04 16.4825 ;
        RECT  -4.025 16.185 -3.96 16.495 ;
        RECT  -3.5025 16.185 -3.4375 16.35 ;
        RECT  -3.3625 16.185 -3.2975 16.35 ;
        RECT  -3.7575 17.02 -3.6925 17.335 ;
        RECT  -3.7125 16.4175 -3.4375 16.4825 ;
        RECT  -3.7125 16.6075 -3.4375 16.6725 ;
        RECT  -3.7125 16.6075 -3.4375 16.6725 ;
        RECT  -3.7125 16.7975 -3.4375 16.8625 ;
        RECT  -3.7125 16.7975 -3.4375 16.8625 ;
        RECT  -3.7125 16.9875 -3.4375 17.0525 ;
        RECT  -4.2375 16.4175 -4.1025 16.4825 ;
        RECT  -4.2375 16.6075 -4.1025 16.6725 ;
        RECT  -4.2375 16.6075 -4.1025 16.6725 ;
        RECT  -4.2375 16.7975 -4.1025 16.8625 ;
        RECT  -4.2375 16.7975 -4.1025 16.8625 ;
        RECT  -4.2375 16.9875 -4.1025 17.0525 ;
        RECT  -4.2375 17.1575 -4.1025 17.2225 ;
        RECT  -3.4375 17.1575 -3.1625 17.2225 ;
        RECT  -4.2375 16.6075 -4.1025 16.6725 ;
        RECT  -4.2375 16.9875 -4.1025 17.0525 ;
        RECT  -4.02 16.36 -3.955 16.495 ;
        RECT  -3.6375 16.665 -3.5025 16.73 ;
        RECT  -3.6375 16.6625 -3.5025 16.7275 ;
        RECT  -3.5 16.215 -3.435 16.35 ;
        RECT  -3.6375 16.855 -3.5025 16.92 ;
        RECT  -3.6375 16.8525 -3.5025 16.9175 ;
        RECT  -3.36 16.215 -3.295 16.35 ;
        RECT  -3.0725 17.335 -3.0075 17.895 ;
        RECT  -1.7275 17.335 -1.6625 17.895 ;
        RECT  -2.0925 17.7625 -1.7275 17.8275 ;
        RECT  -3.0075 17.7625 -2.8725 17.8275 ;
        RECT  -3.0075 17.4025 -2.9375 17.4675 ;
        RECT  -1.8175 17.4025 -1.7275 17.4675 ;
        RECT  -2.905 17.5925 -1.9575 17.6575 ;
        RECT  -2.49 17.335 -2.425 17.37 ;
        RECT  -2.49 17.6575 -2.425 17.895 ;
        RECT  -2.8725 17.4025 -2.7375 17.4675 ;
        RECT  -2.8725 17.5925 -2.7375 17.6575 ;
        RECT  -2.4725 17.4025 -2.1975 17.4675 ;
        RECT  -2.4725 17.5925 -2.1975 17.6575 ;
        RECT  -2.3675 17.7625 -2.0925 17.8275 ;
        RECT  -3.0725 17.7625 -2.9375 17.8275 ;
        RECT  -2.565 17.37 -2.5 17.505 ;
        RECT  -3.0725 17.335 -3.0075 17.895 ;
        RECT  -4.4175 17.335 -4.3525 17.895 ;
        RECT  -4.3525 17.7625 -3.9875 17.8275 ;
        RECT  -3.2075 17.7625 -3.0725 17.8275 ;
        RECT  -3.1425 17.4025 -3.0725 17.4675 ;
        RECT  -4.3525 17.4025 -4.2625 17.4675 ;
        RECT  -4.1225 17.5925 -3.175 17.6575 ;
        RECT  -3.655 17.335 -3.59 17.37 ;
        RECT  -3.655 17.6575 -3.59 17.895 ;
        RECT  -3.4125 17.4025 -3.2775 17.4675 ;
        RECT  -3.4125 17.5925 -3.2775 17.6575 ;
        RECT  -4.2625 17.4025 -3.9875 17.4675 ;
        RECT  -4.2625 17.5925 -3.9875 17.6575 ;
        RECT  -4.2625 17.7625 -3.9875 17.8275 ;
        RECT  -3.2775 17.7625 -3.1425 17.8275 ;
        RECT  -3.655 17.37 -3.59 17.505 ;
        RECT  -3.0725 17.895 -3.0075 18.455 ;
        RECT  -4.4175 17.895 -4.3525 18.455 ;
        RECT  -4.3525 18.3225 -3.9875 18.3875 ;
        RECT  -3.2075 18.3225 -3.0725 18.3875 ;
        RECT  -3.1425 17.9625 -3.0725 18.0275 ;
        RECT  -4.3525 17.9625 -4.2625 18.0275 ;
        RECT  -4.1225 18.1525 -3.175 18.2175 ;
        RECT  -3.655 17.895 -3.59 17.93 ;
        RECT  -3.655 18.2175 -3.59 18.455 ;
        RECT  -3.4125 17.9625 -3.2775 18.0275 ;
        RECT  -3.4125 18.1525 -3.2775 18.2175 ;
        RECT  -4.2625 17.9625 -3.9875 18.0275 ;
        RECT  -4.2625 18.1525 -3.9875 18.2175 ;
        RECT  -4.2625 18.3225 -3.9875 18.3875 ;
        RECT  -3.2775 18.3225 -3.1425 18.3875 ;
        RECT  -3.655 17.93 -3.59 18.065 ;
        RECT  -3.0725 18.455 -3.0075 19.015 ;
        RECT  -4.4175 18.455 -4.3525 19.015 ;
        RECT  -4.3525 18.8825 -3.9875 18.9475 ;
        RECT  -3.2075 18.8825 -3.0725 18.9475 ;
        RECT  -3.1425 18.5225 -3.0725 18.5875 ;
        RECT  -4.3525 18.5225 -4.2625 18.5875 ;
        RECT  -4.1225 18.7125 -3.175 18.7775 ;
        RECT  -3.655 18.455 -3.59 18.49 ;
        RECT  -3.655 18.7775 -3.59 19.015 ;
        RECT  -3.4125 18.5225 -3.2775 18.5875 ;
        RECT  -3.4125 18.7125 -3.2775 18.7775 ;
        RECT  -4.2625 18.5225 -3.9875 18.5875 ;
        RECT  -4.2625 18.7125 -3.9875 18.7775 ;
        RECT  -4.2625 18.8825 -3.9875 18.9475 ;
        RECT  -3.2775 18.8825 -3.1425 18.9475 ;
        RECT  -3.655 18.49 -3.59 18.625 ;
        RECT  -3.9975 14.615 -3.9325 14.75 ;
        RECT  -3.9975 15.105 -3.9325 15.24 ;
        RECT  -4.1525 14.615 -4.0875 14.75 ;
        RECT  -4.1525 15.315 -4.0875 15.45 ;
        RECT  -5.5625 14.615 -5.4975 14.75 ;
        RECT  -5.5625 15.525 -5.4975 15.66 ;
        RECT  -4.5475 14.615 -4.4825 14.75 ;
        RECT  -4.5475 15.735 -4.4825 15.87 ;
        RECT  -1.325 15.315 -1.26 15.45 ;
        RECT  -0.795 15.945 -0.73 16.08 ;
        RECT  -2.12 15.945 -2.055 16.08 ;
        RECT  -2.6425 15.315 -2.5775 15.45 ;
        RECT  -2.7825 15.525 -2.7175 15.66 ;
        RECT  -4.025 15.945 -3.96 16.08 ;
        RECT  -3.5025 15.735 -3.4375 15.87 ;
        RECT  -3.3625 15.525 -3.2975 15.66 ;
        RECT  -0.9975 9.8175 -0.9325 9.9525 ;
        RECT  -0.22 9.8175 -0.155 9.9525 ;
        RECT  -0.22 15.1025 -0.155 15.2375 ;
        RECT  -2.49 19.405 -2.425 19.54 ;
        RECT  -3.655 19.195 -3.59 19.33 ;
        RECT  -0.965 19.615 -0.9 19.75 ;
        RECT  -0.205 19.4025 -0.14 19.5375 ;
        RECT  -1.7275 19.825 -1.6625 19.96 ;
        RECT  -4.4175 19.825 -4.3525 19.96 ;
        RECT  -0.3825 14.895 -0.3175 15.03 ;
        RECT  -0.965 13.3775 -0.9 13.5125 ;
        RECT  -2.085 13.3775 -2.02 13.5125 ;
        RECT  -2.0825 8.275 -2.0175 8.41 ;
        RECT  -0.865 8.415 -0.8 8.55 ;
        RECT  -1.0825 16.8675 -0.9475 16.9325 ;
        RECT  -1.035 17.3375 -0.9 17.4025 ;
        RECT  0.0325 19.855 0.2375 19.99 ;
        LAYER  via1 ;
        RECT  11.835 19.68 11.9 19.745 ;
        RECT  11.835 19.68 11.9 19.745 ;
        RECT  11.835 19.68 11.9 19.745 ;
        RECT  11.835 19.68 11.9 19.745 ;
        RECT  11.835 19.68 11.9 19.745 ;
        RECT  11.835 19.68 11.9 19.745 ;
        RECT  11.13 18.8625 11.195 18.9275 ;
        RECT  11.835 18.8625 11.9 18.9275 ;
        RECT  11.835 19.68 11.9 19.745 ;
        RECT  11.835 19.68 11.9 19.745 ;
        RECT  11.835 19.68 11.9 19.745 ;
        RECT  11.835 19.68 11.9 19.745 ;
        RECT  11.835 19.68 11.9 19.745 ;
        RECT  11.835 19.68 11.9 19.745 ;
        RECT  11.835 19.68 11.9 19.745 ;
        RECT  11.835 19.68 11.9 19.745 ;
        RECT  11.385 19.1875 11.45 19.2525 ;
        RECT  11.13 19.68 11.195 19.745 ;
        RECT  11.13 19.68 11.195 19.745 ;
        RECT  11.13 19.68 11.195 19.745 ;
        RECT  11.13 19.68 11.195 19.745 ;
        RECT  11.13 19.68 11.195 19.745 ;
        RECT  11.13 19.68 11.195 19.745 ;
        RECT  11.835 19.68 11.9 19.745 ;
        RECT  11.835 19.68 11.9 19.745 ;
        RECT  11.835 19.68 11.9 19.745 ;
        RECT  11.835 19.68 11.9 19.745 ;
        RECT  11.58 19.1875 11.645 19.2525 ;
        RECT  11.835 18.8625 11.9 18.9275 ;
        RECT  11.835 18.8625 11.9 18.9275 ;
        RECT  11.835 18.8625 11.9 18.9275 ;
        RECT  11.835 19.68 11.9 19.745 ;
        RECT  11.835 19.68 11.9 19.745 ;
        RECT  11.835 19.68 11.9 19.745 ;
        RECT  11.835 19.68 11.9 19.745 ;
        RECT  11.835 19.68 11.9 19.745 ;
        RECT  11.835 19.68 11.9 19.745 ;
        RECT  11.13 18.8625 11.195 18.9275 ;
        RECT  11.835 20.735 11.9 20.8 ;
        RECT  11.835 20.735 11.9 20.8 ;
        RECT  11.835 20.735 11.9 20.8 ;
        RECT  11.835 20.735 11.9 20.8 ;
        RECT  11.835 20.735 11.9 20.8 ;
        RECT  11.835 20.735 11.9 20.8 ;
        RECT  11.13 21.5525 11.195 21.6175 ;
        RECT  11.835 21.5525 11.9 21.6175 ;
        RECT  11.835 20.735 11.9 20.8 ;
        RECT  11.835 20.735 11.9 20.8 ;
        RECT  11.835 20.735 11.9 20.8 ;
        RECT  11.835 20.735 11.9 20.8 ;
        RECT  11.835 20.735 11.9 20.8 ;
        RECT  11.835 20.735 11.9 20.8 ;
        RECT  11.835 20.735 11.9 20.8 ;
        RECT  11.835 20.735 11.9 20.8 ;
        RECT  11.385 21.2275 11.45 21.2925 ;
        RECT  11.13 20.735 11.195 20.8 ;
        RECT  11.13 20.735 11.195 20.8 ;
        RECT  11.13 20.735 11.195 20.8 ;
        RECT  11.13 20.735 11.195 20.8 ;
        RECT  11.13 20.735 11.195 20.8 ;
        RECT  11.13 20.735 11.195 20.8 ;
        RECT  11.835 20.735 11.9 20.8 ;
        RECT  11.835 20.735 11.9 20.8 ;
        RECT  11.835 20.735 11.9 20.8 ;
        RECT  11.835 20.735 11.9 20.8 ;
        RECT  11.58 21.2275 11.645 21.2925 ;
        RECT  11.835 21.5525 11.9 21.6175 ;
        RECT  11.835 21.5525 11.9 21.6175 ;
        RECT  11.835 21.5525 11.9 21.6175 ;
        RECT  11.835 20.735 11.9 20.8 ;
        RECT  11.835 20.735 11.9 20.8 ;
        RECT  11.835 20.735 11.9 20.8 ;
        RECT  11.835 20.735 11.9 20.8 ;
        RECT  11.835 20.735 11.9 20.8 ;
        RECT  11.835 20.735 11.9 20.8 ;
        RECT  11.13 21.5525 11.195 21.6175 ;
        RECT  11.835 22.37 11.9 22.435 ;
        RECT  11.835 22.37 11.9 22.435 ;
        RECT  11.835 22.37 11.9 22.435 ;
        RECT  11.835 22.37 11.9 22.435 ;
        RECT  11.835 22.37 11.9 22.435 ;
        RECT  11.835 22.37 11.9 22.435 ;
        RECT  11.13 21.5525 11.195 21.6175 ;
        RECT  11.835 21.5525 11.9 21.6175 ;
        RECT  11.835 22.37 11.9 22.435 ;
        RECT  11.835 22.37 11.9 22.435 ;
        RECT  11.835 22.37 11.9 22.435 ;
        RECT  11.835 22.37 11.9 22.435 ;
        RECT  11.835 22.37 11.9 22.435 ;
        RECT  11.835 22.37 11.9 22.435 ;
        RECT  11.835 22.37 11.9 22.435 ;
        RECT  11.835 22.37 11.9 22.435 ;
        RECT  11.385 21.8775 11.45 21.9425 ;
        RECT  11.13 22.37 11.195 22.435 ;
        RECT  11.13 22.37 11.195 22.435 ;
        RECT  11.13 22.37 11.195 22.435 ;
        RECT  11.13 22.37 11.195 22.435 ;
        RECT  11.13 22.37 11.195 22.435 ;
        RECT  11.13 22.37 11.195 22.435 ;
        RECT  11.835 22.37 11.9 22.435 ;
        RECT  11.835 22.37 11.9 22.435 ;
        RECT  11.835 22.37 11.9 22.435 ;
        RECT  11.835 22.37 11.9 22.435 ;
        RECT  11.58 21.8775 11.645 21.9425 ;
        RECT  11.835 21.5525 11.9 21.6175 ;
        RECT  11.835 21.5525 11.9 21.6175 ;
        RECT  11.835 21.5525 11.9 21.6175 ;
        RECT  11.835 22.37 11.9 22.435 ;
        RECT  11.835 22.37 11.9 22.435 ;
        RECT  11.835 22.37 11.9 22.435 ;
        RECT  11.835 22.37 11.9 22.435 ;
        RECT  11.835 22.37 11.9 22.435 ;
        RECT  11.835 22.37 11.9 22.435 ;
        RECT  11.13 21.5525 11.195 21.6175 ;
        RECT  11.835 23.425 11.9 23.49 ;
        RECT  11.835 23.425 11.9 23.49 ;
        RECT  11.835 23.425 11.9 23.49 ;
        RECT  11.835 23.425 11.9 23.49 ;
        RECT  11.835 23.425 11.9 23.49 ;
        RECT  11.835 23.425 11.9 23.49 ;
        RECT  11.13 24.2425 11.195 24.3075 ;
        RECT  11.835 24.2425 11.9 24.3075 ;
        RECT  11.835 23.425 11.9 23.49 ;
        RECT  11.835 23.425 11.9 23.49 ;
        RECT  11.835 23.425 11.9 23.49 ;
        RECT  11.835 23.425 11.9 23.49 ;
        RECT  11.835 23.425 11.9 23.49 ;
        RECT  11.835 23.425 11.9 23.49 ;
        RECT  11.835 23.425 11.9 23.49 ;
        RECT  11.835 23.425 11.9 23.49 ;
        RECT  11.385 23.9175 11.45 23.9825 ;
        RECT  11.13 23.425 11.195 23.49 ;
        RECT  11.13 23.425 11.195 23.49 ;
        RECT  11.13 23.425 11.195 23.49 ;
        RECT  11.13 23.425 11.195 23.49 ;
        RECT  11.13 23.425 11.195 23.49 ;
        RECT  11.13 23.425 11.195 23.49 ;
        RECT  11.835 23.425 11.9 23.49 ;
        RECT  11.835 23.425 11.9 23.49 ;
        RECT  11.835 23.425 11.9 23.49 ;
        RECT  11.835 23.425 11.9 23.49 ;
        RECT  11.58 23.9175 11.645 23.9825 ;
        RECT  11.835 24.2425 11.9 24.3075 ;
        RECT  11.835 24.2425 11.9 24.3075 ;
        RECT  11.835 24.2425 11.9 24.3075 ;
        RECT  11.835 23.425 11.9 23.49 ;
        RECT  11.835 23.425 11.9 23.49 ;
        RECT  11.835 23.425 11.9 23.49 ;
        RECT  11.835 23.425 11.9 23.49 ;
        RECT  11.835 23.425 11.9 23.49 ;
        RECT  11.835 23.425 11.9 23.49 ;
        RECT  11.13 24.2425 11.195 24.3075 ;
        RECT  11.835 25.06 11.9 25.125 ;
        RECT  11.835 25.06 11.9 25.125 ;
        RECT  11.835 25.06 11.9 25.125 ;
        RECT  11.835 25.06 11.9 25.125 ;
        RECT  11.835 25.06 11.9 25.125 ;
        RECT  11.835 25.06 11.9 25.125 ;
        RECT  11.13 24.2425 11.195 24.3075 ;
        RECT  11.835 24.2425 11.9 24.3075 ;
        RECT  11.835 25.06 11.9 25.125 ;
        RECT  11.835 25.06 11.9 25.125 ;
        RECT  11.835 25.06 11.9 25.125 ;
        RECT  11.835 25.06 11.9 25.125 ;
        RECT  11.835 25.06 11.9 25.125 ;
        RECT  11.835 25.06 11.9 25.125 ;
        RECT  11.835 25.06 11.9 25.125 ;
        RECT  11.835 25.06 11.9 25.125 ;
        RECT  11.385 24.5675 11.45 24.6325 ;
        RECT  11.13 25.06 11.195 25.125 ;
        RECT  11.13 25.06 11.195 25.125 ;
        RECT  11.13 25.06 11.195 25.125 ;
        RECT  11.13 25.06 11.195 25.125 ;
        RECT  11.13 25.06 11.195 25.125 ;
        RECT  11.13 25.06 11.195 25.125 ;
        RECT  11.835 25.06 11.9 25.125 ;
        RECT  11.835 25.06 11.9 25.125 ;
        RECT  11.835 25.06 11.9 25.125 ;
        RECT  11.835 25.06 11.9 25.125 ;
        RECT  11.58 24.5675 11.645 24.6325 ;
        RECT  11.835 24.2425 11.9 24.3075 ;
        RECT  11.835 24.2425 11.9 24.3075 ;
        RECT  11.835 24.2425 11.9 24.3075 ;
        RECT  11.835 25.06 11.9 25.125 ;
        RECT  11.835 25.06 11.9 25.125 ;
        RECT  11.835 25.06 11.9 25.125 ;
        RECT  11.835 25.06 11.9 25.125 ;
        RECT  11.835 25.06 11.9 25.125 ;
        RECT  11.835 25.06 11.9 25.125 ;
        RECT  11.13 24.2425 11.195 24.3075 ;
        RECT  11.835 26.115 11.9 26.18 ;
        RECT  11.835 26.115 11.9 26.18 ;
        RECT  11.835 26.115 11.9 26.18 ;
        RECT  11.835 26.115 11.9 26.18 ;
        RECT  11.835 26.115 11.9 26.18 ;
        RECT  11.835 26.115 11.9 26.18 ;
        RECT  11.13 26.9325 11.195 26.9975 ;
        RECT  11.835 26.9325 11.9 26.9975 ;
        RECT  11.835 26.115 11.9 26.18 ;
        RECT  11.835 26.115 11.9 26.18 ;
        RECT  11.835 26.115 11.9 26.18 ;
        RECT  11.835 26.115 11.9 26.18 ;
        RECT  11.835 26.115 11.9 26.18 ;
        RECT  11.835 26.115 11.9 26.18 ;
        RECT  11.835 26.115 11.9 26.18 ;
        RECT  11.835 26.115 11.9 26.18 ;
        RECT  11.385 26.6075 11.45 26.6725 ;
        RECT  11.13 26.115 11.195 26.18 ;
        RECT  11.13 26.115 11.195 26.18 ;
        RECT  11.13 26.115 11.195 26.18 ;
        RECT  11.13 26.115 11.195 26.18 ;
        RECT  11.13 26.115 11.195 26.18 ;
        RECT  11.13 26.115 11.195 26.18 ;
        RECT  11.835 26.115 11.9 26.18 ;
        RECT  11.835 26.115 11.9 26.18 ;
        RECT  11.835 26.115 11.9 26.18 ;
        RECT  11.835 26.115 11.9 26.18 ;
        RECT  11.58 26.6075 11.645 26.6725 ;
        RECT  11.835 26.9325 11.9 26.9975 ;
        RECT  11.835 26.9325 11.9 26.9975 ;
        RECT  11.835 26.9325 11.9 26.9975 ;
        RECT  11.835 26.115 11.9 26.18 ;
        RECT  11.835 26.115 11.9 26.18 ;
        RECT  11.835 26.115 11.9 26.18 ;
        RECT  11.835 26.115 11.9 26.18 ;
        RECT  11.835 26.115 11.9 26.18 ;
        RECT  11.835 26.115 11.9 26.18 ;
        RECT  11.13 26.9325 11.195 26.9975 ;
        RECT  11.835 27.75 11.9 27.815 ;
        RECT  11.835 27.75 11.9 27.815 ;
        RECT  11.835 27.75 11.9 27.815 ;
        RECT  11.835 27.75 11.9 27.815 ;
        RECT  11.835 27.75 11.9 27.815 ;
        RECT  11.835 27.75 11.9 27.815 ;
        RECT  11.13 26.9325 11.195 26.9975 ;
        RECT  11.835 26.9325 11.9 26.9975 ;
        RECT  11.835 27.75 11.9 27.815 ;
        RECT  11.835 27.75 11.9 27.815 ;
        RECT  11.835 27.75 11.9 27.815 ;
        RECT  11.835 27.75 11.9 27.815 ;
        RECT  11.835 27.75 11.9 27.815 ;
        RECT  11.835 27.75 11.9 27.815 ;
        RECT  11.835 27.75 11.9 27.815 ;
        RECT  11.835 27.75 11.9 27.815 ;
        RECT  11.385 27.2575 11.45 27.3225 ;
        RECT  11.13 27.75 11.195 27.815 ;
        RECT  11.13 27.75 11.195 27.815 ;
        RECT  11.13 27.75 11.195 27.815 ;
        RECT  11.13 27.75 11.195 27.815 ;
        RECT  11.13 27.75 11.195 27.815 ;
        RECT  11.13 27.75 11.195 27.815 ;
        RECT  11.835 27.75 11.9 27.815 ;
        RECT  11.835 27.75 11.9 27.815 ;
        RECT  11.835 27.75 11.9 27.815 ;
        RECT  11.835 27.75 11.9 27.815 ;
        RECT  11.58 27.2575 11.645 27.3225 ;
        RECT  11.835 26.9325 11.9 26.9975 ;
        RECT  11.835 26.9325 11.9 26.9975 ;
        RECT  11.835 26.9325 11.9 26.9975 ;
        RECT  11.835 27.75 11.9 27.815 ;
        RECT  11.835 27.75 11.9 27.815 ;
        RECT  11.835 27.75 11.9 27.815 ;
        RECT  11.835 27.75 11.9 27.815 ;
        RECT  11.835 27.75 11.9 27.815 ;
        RECT  11.835 27.75 11.9 27.815 ;
        RECT  11.13 26.9325 11.195 26.9975 ;
        RECT  11.835 28.805 11.9 28.87 ;
        RECT  11.835 28.805 11.9 28.87 ;
        RECT  11.835 28.805 11.9 28.87 ;
        RECT  11.835 28.805 11.9 28.87 ;
        RECT  11.835 28.805 11.9 28.87 ;
        RECT  11.835 28.805 11.9 28.87 ;
        RECT  11.13 29.6225 11.195 29.6875 ;
        RECT  11.835 29.6225 11.9 29.6875 ;
        RECT  11.835 28.805 11.9 28.87 ;
        RECT  11.835 28.805 11.9 28.87 ;
        RECT  11.835 28.805 11.9 28.87 ;
        RECT  11.835 28.805 11.9 28.87 ;
        RECT  11.835 28.805 11.9 28.87 ;
        RECT  11.835 28.805 11.9 28.87 ;
        RECT  11.835 28.805 11.9 28.87 ;
        RECT  11.835 28.805 11.9 28.87 ;
        RECT  11.385 29.2975 11.45 29.3625 ;
        RECT  11.13 28.805 11.195 28.87 ;
        RECT  11.13 28.805 11.195 28.87 ;
        RECT  11.13 28.805 11.195 28.87 ;
        RECT  11.13 28.805 11.195 28.87 ;
        RECT  11.13 28.805 11.195 28.87 ;
        RECT  11.13 28.805 11.195 28.87 ;
        RECT  11.835 28.805 11.9 28.87 ;
        RECT  11.835 28.805 11.9 28.87 ;
        RECT  11.835 28.805 11.9 28.87 ;
        RECT  11.835 28.805 11.9 28.87 ;
        RECT  11.58 29.2975 11.645 29.3625 ;
        RECT  11.835 29.6225 11.9 29.6875 ;
        RECT  11.835 29.6225 11.9 29.6875 ;
        RECT  11.835 29.6225 11.9 29.6875 ;
        RECT  11.835 28.805 11.9 28.87 ;
        RECT  11.835 28.805 11.9 28.87 ;
        RECT  11.835 28.805 11.9 28.87 ;
        RECT  11.835 28.805 11.9 28.87 ;
        RECT  11.835 28.805 11.9 28.87 ;
        RECT  11.835 28.805 11.9 28.87 ;
        RECT  11.13 29.6225 11.195 29.6875 ;
        RECT  11.835 30.44 11.9 30.505 ;
        RECT  11.835 30.44 11.9 30.505 ;
        RECT  11.835 30.44 11.9 30.505 ;
        RECT  11.835 30.44 11.9 30.505 ;
        RECT  11.835 30.44 11.9 30.505 ;
        RECT  11.835 30.44 11.9 30.505 ;
        RECT  11.13 29.6225 11.195 29.6875 ;
        RECT  11.835 29.6225 11.9 29.6875 ;
        RECT  11.835 30.44 11.9 30.505 ;
        RECT  11.835 30.44 11.9 30.505 ;
        RECT  11.835 30.44 11.9 30.505 ;
        RECT  11.835 30.44 11.9 30.505 ;
        RECT  11.835 30.44 11.9 30.505 ;
        RECT  11.835 30.44 11.9 30.505 ;
        RECT  11.835 30.44 11.9 30.505 ;
        RECT  11.835 30.44 11.9 30.505 ;
        RECT  11.385 29.9475 11.45 30.0125 ;
        RECT  11.13 30.44 11.195 30.505 ;
        RECT  11.13 30.44 11.195 30.505 ;
        RECT  11.13 30.44 11.195 30.505 ;
        RECT  11.13 30.44 11.195 30.505 ;
        RECT  11.13 30.44 11.195 30.505 ;
        RECT  11.13 30.44 11.195 30.505 ;
        RECT  11.835 30.44 11.9 30.505 ;
        RECT  11.835 30.44 11.9 30.505 ;
        RECT  11.835 30.44 11.9 30.505 ;
        RECT  11.835 30.44 11.9 30.505 ;
        RECT  11.58 29.9475 11.645 30.0125 ;
        RECT  11.835 29.6225 11.9 29.6875 ;
        RECT  11.835 29.6225 11.9 29.6875 ;
        RECT  11.835 29.6225 11.9 29.6875 ;
        RECT  11.835 30.44 11.9 30.505 ;
        RECT  11.835 30.44 11.9 30.505 ;
        RECT  11.835 30.44 11.9 30.505 ;
        RECT  11.835 30.44 11.9 30.505 ;
        RECT  11.835 30.44 11.9 30.505 ;
        RECT  11.835 30.44 11.9 30.505 ;
        RECT  11.13 29.6225 11.195 29.6875 ;
        RECT  11.835 31.495 11.9 31.56 ;
        RECT  11.835 31.495 11.9 31.56 ;
        RECT  11.835 31.495 11.9 31.56 ;
        RECT  11.835 31.495 11.9 31.56 ;
        RECT  11.835 31.495 11.9 31.56 ;
        RECT  11.835 31.495 11.9 31.56 ;
        RECT  11.13 32.3125 11.195 32.3775 ;
        RECT  11.835 32.3125 11.9 32.3775 ;
        RECT  11.835 31.495 11.9 31.56 ;
        RECT  11.835 31.495 11.9 31.56 ;
        RECT  11.835 31.495 11.9 31.56 ;
        RECT  11.835 31.495 11.9 31.56 ;
        RECT  11.835 31.495 11.9 31.56 ;
        RECT  11.835 31.495 11.9 31.56 ;
        RECT  11.835 31.495 11.9 31.56 ;
        RECT  11.835 31.495 11.9 31.56 ;
        RECT  11.385 31.9875 11.45 32.0525 ;
        RECT  11.13 31.495 11.195 31.56 ;
        RECT  11.13 31.495 11.195 31.56 ;
        RECT  11.13 31.495 11.195 31.56 ;
        RECT  11.13 31.495 11.195 31.56 ;
        RECT  11.13 31.495 11.195 31.56 ;
        RECT  11.13 31.495 11.195 31.56 ;
        RECT  11.835 31.495 11.9 31.56 ;
        RECT  11.835 31.495 11.9 31.56 ;
        RECT  11.835 31.495 11.9 31.56 ;
        RECT  11.835 31.495 11.9 31.56 ;
        RECT  11.58 31.9875 11.645 32.0525 ;
        RECT  11.835 32.3125 11.9 32.3775 ;
        RECT  11.835 32.3125 11.9 32.3775 ;
        RECT  11.835 32.3125 11.9 32.3775 ;
        RECT  11.835 31.495 11.9 31.56 ;
        RECT  11.835 31.495 11.9 31.56 ;
        RECT  11.835 31.495 11.9 31.56 ;
        RECT  11.835 31.495 11.9 31.56 ;
        RECT  11.835 31.495 11.9 31.56 ;
        RECT  11.835 31.495 11.9 31.56 ;
        RECT  11.13 32.3125 11.195 32.3775 ;
        RECT  11.835 33.13 11.9 33.195 ;
        RECT  11.835 33.13 11.9 33.195 ;
        RECT  11.835 33.13 11.9 33.195 ;
        RECT  11.835 33.13 11.9 33.195 ;
        RECT  11.835 33.13 11.9 33.195 ;
        RECT  11.835 33.13 11.9 33.195 ;
        RECT  11.13 32.3125 11.195 32.3775 ;
        RECT  11.835 32.3125 11.9 32.3775 ;
        RECT  11.835 33.13 11.9 33.195 ;
        RECT  11.835 33.13 11.9 33.195 ;
        RECT  11.835 33.13 11.9 33.195 ;
        RECT  11.835 33.13 11.9 33.195 ;
        RECT  11.835 33.13 11.9 33.195 ;
        RECT  11.835 33.13 11.9 33.195 ;
        RECT  11.835 33.13 11.9 33.195 ;
        RECT  11.835 33.13 11.9 33.195 ;
        RECT  11.385 32.6375 11.45 32.7025 ;
        RECT  11.13 33.13 11.195 33.195 ;
        RECT  11.13 33.13 11.195 33.195 ;
        RECT  11.13 33.13 11.195 33.195 ;
        RECT  11.13 33.13 11.195 33.195 ;
        RECT  11.13 33.13 11.195 33.195 ;
        RECT  11.13 33.13 11.195 33.195 ;
        RECT  11.835 33.13 11.9 33.195 ;
        RECT  11.835 33.13 11.9 33.195 ;
        RECT  11.835 33.13 11.9 33.195 ;
        RECT  11.835 33.13 11.9 33.195 ;
        RECT  11.58 32.6375 11.645 32.7025 ;
        RECT  11.835 32.3125 11.9 32.3775 ;
        RECT  11.835 32.3125 11.9 32.3775 ;
        RECT  11.835 32.3125 11.9 32.3775 ;
        RECT  11.835 33.13 11.9 33.195 ;
        RECT  11.835 33.13 11.9 33.195 ;
        RECT  11.835 33.13 11.9 33.195 ;
        RECT  11.835 33.13 11.9 33.195 ;
        RECT  11.835 33.13 11.9 33.195 ;
        RECT  11.835 33.13 11.9 33.195 ;
        RECT  11.13 32.3125 11.195 32.3775 ;
        RECT  11.835 34.185 11.9 34.25 ;
        RECT  11.835 34.185 11.9 34.25 ;
        RECT  11.835 34.185 11.9 34.25 ;
        RECT  11.835 34.185 11.9 34.25 ;
        RECT  11.835 34.185 11.9 34.25 ;
        RECT  11.835 34.185 11.9 34.25 ;
        RECT  11.13 35.0025 11.195 35.0675 ;
        RECT  11.835 35.0025 11.9 35.0675 ;
        RECT  11.835 34.185 11.9 34.25 ;
        RECT  11.835 34.185 11.9 34.25 ;
        RECT  11.835 34.185 11.9 34.25 ;
        RECT  11.835 34.185 11.9 34.25 ;
        RECT  11.835 34.185 11.9 34.25 ;
        RECT  11.835 34.185 11.9 34.25 ;
        RECT  11.835 34.185 11.9 34.25 ;
        RECT  11.835 34.185 11.9 34.25 ;
        RECT  11.385 34.6775 11.45 34.7425 ;
        RECT  11.13 34.185 11.195 34.25 ;
        RECT  11.13 34.185 11.195 34.25 ;
        RECT  11.13 34.185 11.195 34.25 ;
        RECT  11.13 34.185 11.195 34.25 ;
        RECT  11.13 34.185 11.195 34.25 ;
        RECT  11.13 34.185 11.195 34.25 ;
        RECT  11.835 34.185 11.9 34.25 ;
        RECT  11.835 34.185 11.9 34.25 ;
        RECT  11.835 34.185 11.9 34.25 ;
        RECT  11.835 34.185 11.9 34.25 ;
        RECT  11.58 34.6775 11.645 34.7425 ;
        RECT  11.835 35.0025 11.9 35.0675 ;
        RECT  11.835 35.0025 11.9 35.0675 ;
        RECT  11.835 35.0025 11.9 35.0675 ;
        RECT  11.835 34.185 11.9 34.25 ;
        RECT  11.835 34.185 11.9 34.25 ;
        RECT  11.835 34.185 11.9 34.25 ;
        RECT  11.835 34.185 11.9 34.25 ;
        RECT  11.835 34.185 11.9 34.25 ;
        RECT  11.835 34.185 11.9 34.25 ;
        RECT  11.13 35.0025 11.195 35.0675 ;
        RECT  11.835 35.82 11.9 35.885 ;
        RECT  11.835 35.82 11.9 35.885 ;
        RECT  11.835 35.82 11.9 35.885 ;
        RECT  11.835 35.82 11.9 35.885 ;
        RECT  11.835 35.82 11.9 35.885 ;
        RECT  11.835 35.82 11.9 35.885 ;
        RECT  11.13 35.0025 11.195 35.0675 ;
        RECT  11.835 35.0025 11.9 35.0675 ;
        RECT  11.835 35.82 11.9 35.885 ;
        RECT  11.835 35.82 11.9 35.885 ;
        RECT  11.835 35.82 11.9 35.885 ;
        RECT  11.835 35.82 11.9 35.885 ;
        RECT  11.835 35.82 11.9 35.885 ;
        RECT  11.835 35.82 11.9 35.885 ;
        RECT  11.835 35.82 11.9 35.885 ;
        RECT  11.835 35.82 11.9 35.885 ;
        RECT  11.385 35.3275 11.45 35.3925 ;
        RECT  11.13 35.82 11.195 35.885 ;
        RECT  11.13 35.82 11.195 35.885 ;
        RECT  11.13 35.82 11.195 35.885 ;
        RECT  11.13 35.82 11.195 35.885 ;
        RECT  11.13 35.82 11.195 35.885 ;
        RECT  11.13 35.82 11.195 35.885 ;
        RECT  11.835 35.82 11.9 35.885 ;
        RECT  11.835 35.82 11.9 35.885 ;
        RECT  11.835 35.82 11.9 35.885 ;
        RECT  11.835 35.82 11.9 35.885 ;
        RECT  11.58 35.3275 11.645 35.3925 ;
        RECT  11.835 35.0025 11.9 35.0675 ;
        RECT  11.835 35.0025 11.9 35.0675 ;
        RECT  11.835 35.0025 11.9 35.0675 ;
        RECT  11.835 35.82 11.9 35.885 ;
        RECT  11.835 35.82 11.9 35.885 ;
        RECT  11.835 35.82 11.9 35.885 ;
        RECT  11.835 35.82 11.9 35.885 ;
        RECT  11.835 35.82 11.9 35.885 ;
        RECT  11.835 35.82 11.9 35.885 ;
        RECT  11.13 35.0025 11.195 35.0675 ;
        RECT  11.835 36.875 11.9 36.94 ;
        RECT  11.835 36.875 11.9 36.94 ;
        RECT  11.835 36.875 11.9 36.94 ;
        RECT  11.835 36.875 11.9 36.94 ;
        RECT  11.835 36.875 11.9 36.94 ;
        RECT  11.835 36.875 11.9 36.94 ;
        RECT  11.13 37.6925 11.195 37.7575 ;
        RECT  11.835 37.6925 11.9 37.7575 ;
        RECT  11.835 36.875 11.9 36.94 ;
        RECT  11.835 36.875 11.9 36.94 ;
        RECT  11.835 36.875 11.9 36.94 ;
        RECT  11.835 36.875 11.9 36.94 ;
        RECT  11.835 36.875 11.9 36.94 ;
        RECT  11.835 36.875 11.9 36.94 ;
        RECT  11.835 36.875 11.9 36.94 ;
        RECT  11.835 36.875 11.9 36.94 ;
        RECT  11.385 37.3675 11.45 37.4325 ;
        RECT  11.13 36.875 11.195 36.94 ;
        RECT  11.13 36.875 11.195 36.94 ;
        RECT  11.13 36.875 11.195 36.94 ;
        RECT  11.13 36.875 11.195 36.94 ;
        RECT  11.13 36.875 11.195 36.94 ;
        RECT  11.13 36.875 11.195 36.94 ;
        RECT  11.835 36.875 11.9 36.94 ;
        RECT  11.835 36.875 11.9 36.94 ;
        RECT  11.835 36.875 11.9 36.94 ;
        RECT  11.835 36.875 11.9 36.94 ;
        RECT  11.58 37.3675 11.645 37.4325 ;
        RECT  11.835 37.6925 11.9 37.7575 ;
        RECT  11.835 37.6925 11.9 37.7575 ;
        RECT  11.835 37.6925 11.9 37.7575 ;
        RECT  11.835 36.875 11.9 36.94 ;
        RECT  11.835 36.875 11.9 36.94 ;
        RECT  11.835 36.875 11.9 36.94 ;
        RECT  11.835 36.875 11.9 36.94 ;
        RECT  11.835 36.875 11.9 36.94 ;
        RECT  11.835 36.875 11.9 36.94 ;
        RECT  11.13 37.6925 11.195 37.7575 ;
        RECT  11.835 38.51 11.9 38.575 ;
        RECT  11.835 38.51 11.9 38.575 ;
        RECT  11.835 38.51 11.9 38.575 ;
        RECT  11.835 38.51 11.9 38.575 ;
        RECT  11.835 38.51 11.9 38.575 ;
        RECT  11.835 38.51 11.9 38.575 ;
        RECT  11.13 37.6925 11.195 37.7575 ;
        RECT  11.835 37.6925 11.9 37.7575 ;
        RECT  11.835 38.51 11.9 38.575 ;
        RECT  11.835 38.51 11.9 38.575 ;
        RECT  11.835 38.51 11.9 38.575 ;
        RECT  11.835 38.51 11.9 38.575 ;
        RECT  11.835 38.51 11.9 38.575 ;
        RECT  11.835 38.51 11.9 38.575 ;
        RECT  11.835 38.51 11.9 38.575 ;
        RECT  11.835 38.51 11.9 38.575 ;
        RECT  11.385 38.0175 11.45 38.0825 ;
        RECT  11.13 38.51 11.195 38.575 ;
        RECT  11.13 38.51 11.195 38.575 ;
        RECT  11.13 38.51 11.195 38.575 ;
        RECT  11.13 38.51 11.195 38.575 ;
        RECT  11.13 38.51 11.195 38.575 ;
        RECT  11.13 38.51 11.195 38.575 ;
        RECT  11.835 38.51 11.9 38.575 ;
        RECT  11.835 38.51 11.9 38.575 ;
        RECT  11.835 38.51 11.9 38.575 ;
        RECT  11.835 38.51 11.9 38.575 ;
        RECT  11.58 38.0175 11.645 38.0825 ;
        RECT  11.835 37.6925 11.9 37.7575 ;
        RECT  11.835 37.6925 11.9 37.7575 ;
        RECT  11.835 37.6925 11.9 37.7575 ;
        RECT  11.835 38.51 11.9 38.575 ;
        RECT  11.835 38.51 11.9 38.575 ;
        RECT  11.835 38.51 11.9 38.575 ;
        RECT  11.835 38.51 11.9 38.575 ;
        RECT  11.835 38.51 11.9 38.575 ;
        RECT  11.835 38.51 11.9 38.575 ;
        RECT  11.13 37.6925 11.195 37.7575 ;
        RECT  11.835 39.565 11.9 39.63 ;
        RECT  11.835 39.565 11.9 39.63 ;
        RECT  11.835 39.565 11.9 39.63 ;
        RECT  11.835 39.565 11.9 39.63 ;
        RECT  11.835 39.565 11.9 39.63 ;
        RECT  11.835 39.565 11.9 39.63 ;
        RECT  11.13 40.3825 11.195 40.4475 ;
        RECT  11.835 40.3825 11.9 40.4475 ;
        RECT  11.835 39.565 11.9 39.63 ;
        RECT  11.835 39.565 11.9 39.63 ;
        RECT  11.835 39.565 11.9 39.63 ;
        RECT  11.835 39.565 11.9 39.63 ;
        RECT  11.835 39.565 11.9 39.63 ;
        RECT  11.835 39.565 11.9 39.63 ;
        RECT  11.835 39.565 11.9 39.63 ;
        RECT  11.835 39.565 11.9 39.63 ;
        RECT  11.385 40.0575 11.45 40.1225 ;
        RECT  11.13 39.565 11.195 39.63 ;
        RECT  11.13 39.565 11.195 39.63 ;
        RECT  11.13 39.565 11.195 39.63 ;
        RECT  11.13 39.565 11.195 39.63 ;
        RECT  11.13 39.565 11.195 39.63 ;
        RECT  11.13 39.565 11.195 39.63 ;
        RECT  11.835 39.565 11.9 39.63 ;
        RECT  11.835 39.565 11.9 39.63 ;
        RECT  11.835 39.565 11.9 39.63 ;
        RECT  11.835 39.565 11.9 39.63 ;
        RECT  11.58 40.0575 11.645 40.1225 ;
        RECT  11.835 40.3825 11.9 40.4475 ;
        RECT  11.835 40.3825 11.9 40.4475 ;
        RECT  11.835 40.3825 11.9 40.4475 ;
        RECT  11.835 39.565 11.9 39.63 ;
        RECT  11.835 39.565 11.9 39.63 ;
        RECT  11.835 39.565 11.9 39.63 ;
        RECT  11.835 39.565 11.9 39.63 ;
        RECT  11.835 39.565 11.9 39.63 ;
        RECT  11.835 39.565 11.9 39.63 ;
        RECT  11.13 40.3825 11.195 40.4475 ;
        RECT  12.54 19.68 12.605 19.745 ;
        RECT  12.54 19.68 12.605 19.745 ;
        RECT  12.54 19.68 12.605 19.745 ;
        RECT  12.54 19.68 12.605 19.745 ;
        RECT  12.54 19.68 12.605 19.745 ;
        RECT  12.54 19.68 12.605 19.745 ;
        RECT  11.835 18.8625 11.9 18.9275 ;
        RECT  12.54 18.8625 12.605 18.9275 ;
        RECT  12.54 19.68 12.605 19.745 ;
        RECT  12.54 19.68 12.605 19.745 ;
        RECT  12.54 19.68 12.605 19.745 ;
        RECT  12.54 19.68 12.605 19.745 ;
        RECT  12.54 19.68 12.605 19.745 ;
        RECT  12.54 19.68 12.605 19.745 ;
        RECT  12.54 19.68 12.605 19.745 ;
        RECT  12.54 19.68 12.605 19.745 ;
        RECT  12.09 19.1875 12.155 19.2525 ;
        RECT  11.835 19.68 11.9 19.745 ;
        RECT  11.835 19.68 11.9 19.745 ;
        RECT  11.835 19.68 11.9 19.745 ;
        RECT  11.835 19.68 11.9 19.745 ;
        RECT  11.835 19.68 11.9 19.745 ;
        RECT  11.835 19.68 11.9 19.745 ;
        RECT  12.54 19.68 12.605 19.745 ;
        RECT  12.54 19.68 12.605 19.745 ;
        RECT  12.54 19.68 12.605 19.745 ;
        RECT  12.54 19.68 12.605 19.745 ;
        RECT  12.285 19.1875 12.35 19.2525 ;
        RECT  12.54 18.8625 12.605 18.9275 ;
        RECT  12.54 18.8625 12.605 18.9275 ;
        RECT  12.54 18.8625 12.605 18.9275 ;
        RECT  12.54 19.68 12.605 19.745 ;
        RECT  12.54 19.68 12.605 19.745 ;
        RECT  12.54 19.68 12.605 19.745 ;
        RECT  12.54 19.68 12.605 19.745 ;
        RECT  12.54 19.68 12.605 19.745 ;
        RECT  12.54 19.68 12.605 19.745 ;
        RECT  11.835 18.8625 11.9 18.9275 ;
        RECT  12.54 20.735 12.605 20.8 ;
        RECT  12.54 20.735 12.605 20.8 ;
        RECT  12.54 20.735 12.605 20.8 ;
        RECT  12.54 20.735 12.605 20.8 ;
        RECT  12.54 20.735 12.605 20.8 ;
        RECT  12.54 20.735 12.605 20.8 ;
        RECT  11.835 21.5525 11.9 21.6175 ;
        RECT  12.54 21.5525 12.605 21.6175 ;
        RECT  12.54 20.735 12.605 20.8 ;
        RECT  12.54 20.735 12.605 20.8 ;
        RECT  12.54 20.735 12.605 20.8 ;
        RECT  12.54 20.735 12.605 20.8 ;
        RECT  12.54 20.735 12.605 20.8 ;
        RECT  12.54 20.735 12.605 20.8 ;
        RECT  12.54 20.735 12.605 20.8 ;
        RECT  12.54 20.735 12.605 20.8 ;
        RECT  12.09 21.2275 12.155 21.2925 ;
        RECT  11.835 20.735 11.9 20.8 ;
        RECT  11.835 20.735 11.9 20.8 ;
        RECT  11.835 20.735 11.9 20.8 ;
        RECT  11.835 20.735 11.9 20.8 ;
        RECT  11.835 20.735 11.9 20.8 ;
        RECT  11.835 20.735 11.9 20.8 ;
        RECT  12.54 20.735 12.605 20.8 ;
        RECT  12.54 20.735 12.605 20.8 ;
        RECT  12.54 20.735 12.605 20.8 ;
        RECT  12.54 20.735 12.605 20.8 ;
        RECT  12.285 21.2275 12.35 21.2925 ;
        RECT  12.54 21.5525 12.605 21.6175 ;
        RECT  12.54 21.5525 12.605 21.6175 ;
        RECT  12.54 21.5525 12.605 21.6175 ;
        RECT  12.54 20.735 12.605 20.8 ;
        RECT  12.54 20.735 12.605 20.8 ;
        RECT  12.54 20.735 12.605 20.8 ;
        RECT  12.54 20.735 12.605 20.8 ;
        RECT  12.54 20.735 12.605 20.8 ;
        RECT  12.54 20.735 12.605 20.8 ;
        RECT  11.835 21.5525 11.9 21.6175 ;
        RECT  12.54 22.37 12.605 22.435 ;
        RECT  12.54 22.37 12.605 22.435 ;
        RECT  12.54 22.37 12.605 22.435 ;
        RECT  12.54 22.37 12.605 22.435 ;
        RECT  12.54 22.37 12.605 22.435 ;
        RECT  12.54 22.37 12.605 22.435 ;
        RECT  11.835 21.5525 11.9 21.6175 ;
        RECT  12.54 21.5525 12.605 21.6175 ;
        RECT  12.54 22.37 12.605 22.435 ;
        RECT  12.54 22.37 12.605 22.435 ;
        RECT  12.54 22.37 12.605 22.435 ;
        RECT  12.54 22.37 12.605 22.435 ;
        RECT  12.54 22.37 12.605 22.435 ;
        RECT  12.54 22.37 12.605 22.435 ;
        RECT  12.54 22.37 12.605 22.435 ;
        RECT  12.54 22.37 12.605 22.435 ;
        RECT  12.09 21.8775 12.155 21.9425 ;
        RECT  11.835 22.37 11.9 22.435 ;
        RECT  11.835 22.37 11.9 22.435 ;
        RECT  11.835 22.37 11.9 22.435 ;
        RECT  11.835 22.37 11.9 22.435 ;
        RECT  11.835 22.37 11.9 22.435 ;
        RECT  11.835 22.37 11.9 22.435 ;
        RECT  12.54 22.37 12.605 22.435 ;
        RECT  12.54 22.37 12.605 22.435 ;
        RECT  12.54 22.37 12.605 22.435 ;
        RECT  12.54 22.37 12.605 22.435 ;
        RECT  12.285 21.8775 12.35 21.9425 ;
        RECT  12.54 21.5525 12.605 21.6175 ;
        RECT  12.54 21.5525 12.605 21.6175 ;
        RECT  12.54 21.5525 12.605 21.6175 ;
        RECT  12.54 22.37 12.605 22.435 ;
        RECT  12.54 22.37 12.605 22.435 ;
        RECT  12.54 22.37 12.605 22.435 ;
        RECT  12.54 22.37 12.605 22.435 ;
        RECT  12.54 22.37 12.605 22.435 ;
        RECT  12.54 22.37 12.605 22.435 ;
        RECT  11.835 21.5525 11.9 21.6175 ;
        RECT  12.54 23.425 12.605 23.49 ;
        RECT  12.54 23.425 12.605 23.49 ;
        RECT  12.54 23.425 12.605 23.49 ;
        RECT  12.54 23.425 12.605 23.49 ;
        RECT  12.54 23.425 12.605 23.49 ;
        RECT  12.54 23.425 12.605 23.49 ;
        RECT  11.835 24.2425 11.9 24.3075 ;
        RECT  12.54 24.2425 12.605 24.3075 ;
        RECT  12.54 23.425 12.605 23.49 ;
        RECT  12.54 23.425 12.605 23.49 ;
        RECT  12.54 23.425 12.605 23.49 ;
        RECT  12.54 23.425 12.605 23.49 ;
        RECT  12.54 23.425 12.605 23.49 ;
        RECT  12.54 23.425 12.605 23.49 ;
        RECT  12.54 23.425 12.605 23.49 ;
        RECT  12.54 23.425 12.605 23.49 ;
        RECT  12.09 23.9175 12.155 23.9825 ;
        RECT  11.835 23.425 11.9 23.49 ;
        RECT  11.835 23.425 11.9 23.49 ;
        RECT  11.835 23.425 11.9 23.49 ;
        RECT  11.835 23.425 11.9 23.49 ;
        RECT  11.835 23.425 11.9 23.49 ;
        RECT  11.835 23.425 11.9 23.49 ;
        RECT  12.54 23.425 12.605 23.49 ;
        RECT  12.54 23.425 12.605 23.49 ;
        RECT  12.54 23.425 12.605 23.49 ;
        RECT  12.54 23.425 12.605 23.49 ;
        RECT  12.285 23.9175 12.35 23.9825 ;
        RECT  12.54 24.2425 12.605 24.3075 ;
        RECT  12.54 24.2425 12.605 24.3075 ;
        RECT  12.54 24.2425 12.605 24.3075 ;
        RECT  12.54 23.425 12.605 23.49 ;
        RECT  12.54 23.425 12.605 23.49 ;
        RECT  12.54 23.425 12.605 23.49 ;
        RECT  12.54 23.425 12.605 23.49 ;
        RECT  12.54 23.425 12.605 23.49 ;
        RECT  12.54 23.425 12.605 23.49 ;
        RECT  11.835 24.2425 11.9 24.3075 ;
        RECT  12.54 25.06 12.605 25.125 ;
        RECT  12.54 25.06 12.605 25.125 ;
        RECT  12.54 25.06 12.605 25.125 ;
        RECT  12.54 25.06 12.605 25.125 ;
        RECT  12.54 25.06 12.605 25.125 ;
        RECT  12.54 25.06 12.605 25.125 ;
        RECT  11.835 24.2425 11.9 24.3075 ;
        RECT  12.54 24.2425 12.605 24.3075 ;
        RECT  12.54 25.06 12.605 25.125 ;
        RECT  12.54 25.06 12.605 25.125 ;
        RECT  12.54 25.06 12.605 25.125 ;
        RECT  12.54 25.06 12.605 25.125 ;
        RECT  12.54 25.06 12.605 25.125 ;
        RECT  12.54 25.06 12.605 25.125 ;
        RECT  12.54 25.06 12.605 25.125 ;
        RECT  12.54 25.06 12.605 25.125 ;
        RECT  12.09 24.5675 12.155 24.6325 ;
        RECT  11.835 25.06 11.9 25.125 ;
        RECT  11.835 25.06 11.9 25.125 ;
        RECT  11.835 25.06 11.9 25.125 ;
        RECT  11.835 25.06 11.9 25.125 ;
        RECT  11.835 25.06 11.9 25.125 ;
        RECT  11.835 25.06 11.9 25.125 ;
        RECT  12.54 25.06 12.605 25.125 ;
        RECT  12.54 25.06 12.605 25.125 ;
        RECT  12.54 25.06 12.605 25.125 ;
        RECT  12.54 25.06 12.605 25.125 ;
        RECT  12.285 24.5675 12.35 24.6325 ;
        RECT  12.54 24.2425 12.605 24.3075 ;
        RECT  12.54 24.2425 12.605 24.3075 ;
        RECT  12.54 24.2425 12.605 24.3075 ;
        RECT  12.54 25.06 12.605 25.125 ;
        RECT  12.54 25.06 12.605 25.125 ;
        RECT  12.54 25.06 12.605 25.125 ;
        RECT  12.54 25.06 12.605 25.125 ;
        RECT  12.54 25.06 12.605 25.125 ;
        RECT  12.54 25.06 12.605 25.125 ;
        RECT  11.835 24.2425 11.9 24.3075 ;
        RECT  12.54 26.115 12.605 26.18 ;
        RECT  12.54 26.115 12.605 26.18 ;
        RECT  12.54 26.115 12.605 26.18 ;
        RECT  12.54 26.115 12.605 26.18 ;
        RECT  12.54 26.115 12.605 26.18 ;
        RECT  12.54 26.115 12.605 26.18 ;
        RECT  11.835 26.9325 11.9 26.9975 ;
        RECT  12.54 26.9325 12.605 26.9975 ;
        RECT  12.54 26.115 12.605 26.18 ;
        RECT  12.54 26.115 12.605 26.18 ;
        RECT  12.54 26.115 12.605 26.18 ;
        RECT  12.54 26.115 12.605 26.18 ;
        RECT  12.54 26.115 12.605 26.18 ;
        RECT  12.54 26.115 12.605 26.18 ;
        RECT  12.54 26.115 12.605 26.18 ;
        RECT  12.54 26.115 12.605 26.18 ;
        RECT  12.09 26.6075 12.155 26.6725 ;
        RECT  11.835 26.115 11.9 26.18 ;
        RECT  11.835 26.115 11.9 26.18 ;
        RECT  11.835 26.115 11.9 26.18 ;
        RECT  11.835 26.115 11.9 26.18 ;
        RECT  11.835 26.115 11.9 26.18 ;
        RECT  11.835 26.115 11.9 26.18 ;
        RECT  12.54 26.115 12.605 26.18 ;
        RECT  12.54 26.115 12.605 26.18 ;
        RECT  12.54 26.115 12.605 26.18 ;
        RECT  12.54 26.115 12.605 26.18 ;
        RECT  12.285 26.6075 12.35 26.6725 ;
        RECT  12.54 26.9325 12.605 26.9975 ;
        RECT  12.54 26.9325 12.605 26.9975 ;
        RECT  12.54 26.9325 12.605 26.9975 ;
        RECT  12.54 26.115 12.605 26.18 ;
        RECT  12.54 26.115 12.605 26.18 ;
        RECT  12.54 26.115 12.605 26.18 ;
        RECT  12.54 26.115 12.605 26.18 ;
        RECT  12.54 26.115 12.605 26.18 ;
        RECT  12.54 26.115 12.605 26.18 ;
        RECT  11.835 26.9325 11.9 26.9975 ;
        RECT  12.54 27.75 12.605 27.815 ;
        RECT  12.54 27.75 12.605 27.815 ;
        RECT  12.54 27.75 12.605 27.815 ;
        RECT  12.54 27.75 12.605 27.815 ;
        RECT  12.54 27.75 12.605 27.815 ;
        RECT  12.54 27.75 12.605 27.815 ;
        RECT  11.835 26.9325 11.9 26.9975 ;
        RECT  12.54 26.9325 12.605 26.9975 ;
        RECT  12.54 27.75 12.605 27.815 ;
        RECT  12.54 27.75 12.605 27.815 ;
        RECT  12.54 27.75 12.605 27.815 ;
        RECT  12.54 27.75 12.605 27.815 ;
        RECT  12.54 27.75 12.605 27.815 ;
        RECT  12.54 27.75 12.605 27.815 ;
        RECT  12.54 27.75 12.605 27.815 ;
        RECT  12.54 27.75 12.605 27.815 ;
        RECT  12.09 27.2575 12.155 27.3225 ;
        RECT  11.835 27.75 11.9 27.815 ;
        RECT  11.835 27.75 11.9 27.815 ;
        RECT  11.835 27.75 11.9 27.815 ;
        RECT  11.835 27.75 11.9 27.815 ;
        RECT  11.835 27.75 11.9 27.815 ;
        RECT  11.835 27.75 11.9 27.815 ;
        RECT  12.54 27.75 12.605 27.815 ;
        RECT  12.54 27.75 12.605 27.815 ;
        RECT  12.54 27.75 12.605 27.815 ;
        RECT  12.54 27.75 12.605 27.815 ;
        RECT  12.285 27.2575 12.35 27.3225 ;
        RECT  12.54 26.9325 12.605 26.9975 ;
        RECT  12.54 26.9325 12.605 26.9975 ;
        RECT  12.54 26.9325 12.605 26.9975 ;
        RECT  12.54 27.75 12.605 27.815 ;
        RECT  12.54 27.75 12.605 27.815 ;
        RECT  12.54 27.75 12.605 27.815 ;
        RECT  12.54 27.75 12.605 27.815 ;
        RECT  12.54 27.75 12.605 27.815 ;
        RECT  12.54 27.75 12.605 27.815 ;
        RECT  11.835 26.9325 11.9 26.9975 ;
        RECT  12.54 28.805 12.605 28.87 ;
        RECT  12.54 28.805 12.605 28.87 ;
        RECT  12.54 28.805 12.605 28.87 ;
        RECT  12.54 28.805 12.605 28.87 ;
        RECT  12.54 28.805 12.605 28.87 ;
        RECT  12.54 28.805 12.605 28.87 ;
        RECT  11.835 29.6225 11.9 29.6875 ;
        RECT  12.54 29.6225 12.605 29.6875 ;
        RECT  12.54 28.805 12.605 28.87 ;
        RECT  12.54 28.805 12.605 28.87 ;
        RECT  12.54 28.805 12.605 28.87 ;
        RECT  12.54 28.805 12.605 28.87 ;
        RECT  12.54 28.805 12.605 28.87 ;
        RECT  12.54 28.805 12.605 28.87 ;
        RECT  12.54 28.805 12.605 28.87 ;
        RECT  12.54 28.805 12.605 28.87 ;
        RECT  12.09 29.2975 12.155 29.3625 ;
        RECT  11.835 28.805 11.9 28.87 ;
        RECT  11.835 28.805 11.9 28.87 ;
        RECT  11.835 28.805 11.9 28.87 ;
        RECT  11.835 28.805 11.9 28.87 ;
        RECT  11.835 28.805 11.9 28.87 ;
        RECT  11.835 28.805 11.9 28.87 ;
        RECT  12.54 28.805 12.605 28.87 ;
        RECT  12.54 28.805 12.605 28.87 ;
        RECT  12.54 28.805 12.605 28.87 ;
        RECT  12.54 28.805 12.605 28.87 ;
        RECT  12.285 29.2975 12.35 29.3625 ;
        RECT  12.54 29.6225 12.605 29.6875 ;
        RECT  12.54 29.6225 12.605 29.6875 ;
        RECT  12.54 29.6225 12.605 29.6875 ;
        RECT  12.54 28.805 12.605 28.87 ;
        RECT  12.54 28.805 12.605 28.87 ;
        RECT  12.54 28.805 12.605 28.87 ;
        RECT  12.54 28.805 12.605 28.87 ;
        RECT  12.54 28.805 12.605 28.87 ;
        RECT  12.54 28.805 12.605 28.87 ;
        RECT  11.835 29.6225 11.9 29.6875 ;
        RECT  12.54 30.44 12.605 30.505 ;
        RECT  12.54 30.44 12.605 30.505 ;
        RECT  12.54 30.44 12.605 30.505 ;
        RECT  12.54 30.44 12.605 30.505 ;
        RECT  12.54 30.44 12.605 30.505 ;
        RECT  12.54 30.44 12.605 30.505 ;
        RECT  11.835 29.6225 11.9 29.6875 ;
        RECT  12.54 29.6225 12.605 29.6875 ;
        RECT  12.54 30.44 12.605 30.505 ;
        RECT  12.54 30.44 12.605 30.505 ;
        RECT  12.54 30.44 12.605 30.505 ;
        RECT  12.54 30.44 12.605 30.505 ;
        RECT  12.54 30.44 12.605 30.505 ;
        RECT  12.54 30.44 12.605 30.505 ;
        RECT  12.54 30.44 12.605 30.505 ;
        RECT  12.54 30.44 12.605 30.505 ;
        RECT  12.09 29.9475 12.155 30.0125 ;
        RECT  11.835 30.44 11.9 30.505 ;
        RECT  11.835 30.44 11.9 30.505 ;
        RECT  11.835 30.44 11.9 30.505 ;
        RECT  11.835 30.44 11.9 30.505 ;
        RECT  11.835 30.44 11.9 30.505 ;
        RECT  11.835 30.44 11.9 30.505 ;
        RECT  12.54 30.44 12.605 30.505 ;
        RECT  12.54 30.44 12.605 30.505 ;
        RECT  12.54 30.44 12.605 30.505 ;
        RECT  12.54 30.44 12.605 30.505 ;
        RECT  12.285 29.9475 12.35 30.0125 ;
        RECT  12.54 29.6225 12.605 29.6875 ;
        RECT  12.54 29.6225 12.605 29.6875 ;
        RECT  12.54 29.6225 12.605 29.6875 ;
        RECT  12.54 30.44 12.605 30.505 ;
        RECT  12.54 30.44 12.605 30.505 ;
        RECT  12.54 30.44 12.605 30.505 ;
        RECT  12.54 30.44 12.605 30.505 ;
        RECT  12.54 30.44 12.605 30.505 ;
        RECT  12.54 30.44 12.605 30.505 ;
        RECT  11.835 29.6225 11.9 29.6875 ;
        RECT  12.54 31.495 12.605 31.56 ;
        RECT  12.54 31.495 12.605 31.56 ;
        RECT  12.54 31.495 12.605 31.56 ;
        RECT  12.54 31.495 12.605 31.56 ;
        RECT  12.54 31.495 12.605 31.56 ;
        RECT  12.54 31.495 12.605 31.56 ;
        RECT  11.835 32.3125 11.9 32.3775 ;
        RECT  12.54 32.3125 12.605 32.3775 ;
        RECT  12.54 31.495 12.605 31.56 ;
        RECT  12.54 31.495 12.605 31.56 ;
        RECT  12.54 31.495 12.605 31.56 ;
        RECT  12.54 31.495 12.605 31.56 ;
        RECT  12.54 31.495 12.605 31.56 ;
        RECT  12.54 31.495 12.605 31.56 ;
        RECT  12.54 31.495 12.605 31.56 ;
        RECT  12.54 31.495 12.605 31.56 ;
        RECT  12.09 31.9875 12.155 32.0525 ;
        RECT  11.835 31.495 11.9 31.56 ;
        RECT  11.835 31.495 11.9 31.56 ;
        RECT  11.835 31.495 11.9 31.56 ;
        RECT  11.835 31.495 11.9 31.56 ;
        RECT  11.835 31.495 11.9 31.56 ;
        RECT  11.835 31.495 11.9 31.56 ;
        RECT  12.54 31.495 12.605 31.56 ;
        RECT  12.54 31.495 12.605 31.56 ;
        RECT  12.54 31.495 12.605 31.56 ;
        RECT  12.54 31.495 12.605 31.56 ;
        RECT  12.285 31.9875 12.35 32.0525 ;
        RECT  12.54 32.3125 12.605 32.3775 ;
        RECT  12.54 32.3125 12.605 32.3775 ;
        RECT  12.54 32.3125 12.605 32.3775 ;
        RECT  12.54 31.495 12.605 31.56 ;
        RECT  12.54 31.495 12.605 31.56 ;
        RECT  12.54 31.495 12.605 31.56 ;
        RECT  12.54 31.495 12.605 31.56 ;
        RECT  12.54 31.495 12.605 31.56 ;
        RECT  12.54 31.495 12.605 31.56 ;
        RECT  11.835 32.3125 11.9 32.3775 ;
        RECT  12.54 33.13 12.605 33.195 ;
        RECT  12.54 33.13 12.605 33.195 ;
        RECT  12.54 33.13 12.605 33.195 ;
        RECT  12.54 33.13 12.605 33.195 ;
        RECT  12.54 33.13 12.605 33.195 ;
        RECT  12.54 33.13 12.605 33.195 ;
        RECT  11.835 32.3125 11.9 32.3775 ;
        RECT  12.54 32.3125 12.605 32.3775 ;
        RECT  12.54 33.13 12.605 33.195 ;
        RECT  12.54 33.13 12.605 33.195 ;
        RECT  12.54 33.13 12.605 33.195 ;
        RECT  12.54 33.13 12.605 33.195 ;
        RECT  12.54 33.13 12.605 33.195 ;
        RECT  12.54 33.13 12.605 33.195 ;
        RECT  12.54 33.13 12.605 33.195 ;
        RECT  12.54 33.13 12.605 33.195 ;
        RECT  12.09 32.6375 12.155 32.7025 ;
        RECT  11.835 33.13 11.9 33.195 ;
        RECT  11.835 33.13 11.9 33.195 ;
        RECT  11.835 33.13 11.9 33.195 ;
        RECT  11.835 33.13 11.9 33.195 ;
        RECT  11.835 33.13 11.9 33.195 ;
        RECT  11.835 33.13 11.9 33.195 ;
        RECT  12.54 33.13 12.605 33.195 ;
        RECT  12.54 33.13 12.605 33.195 ;
        RECT  12.54 33.13 12.605 33.195 ;
        RECT  12.54 33.13 12.605 33.195 ;
        RECT  12.285 32.6375 12.35 32.7025 ;
        RECT  12.54 32.3125 12.605 32.3775 ;
        RECT  12.54 32.3125 12.605 32.3775 ;
        RECT  12.54 32.3125 12.605 32.3775 ;
        RECT  12.54 33.13 12.605 33.195 ;
        RECT  12.54 33.13 12.605 33.195 ;
        RECT  12.54 33.13 12.605 33.195 ;
        RECT  12.54 33.13 12.605 33.195 ;
        RECT  12.54 33.13 12.605 33.195 ;
        RECT  12.54 33.13 12.605 33.195 ;
        RECT  11.835 32.3125 11.9 32.3775 ;
        RECT  12.54 34.185 12.605 34.25 ;
        RECT  12.54 34.185 12.605 34.25 ;
        RECT  12.54 34.185 12.605 34.25 ;
        RECT  12.54 34.185 12.605 34.25 ;
        RECT  12.54 34.185 12.605 34.25 ;
        RECT  12.54 34.185 12.605 34.25 ;
        RECT  11.835 35.0025 11.9 35.0675 ;
        RECT  12.54 35.0025 12.605 35.0675 ;
        RECT  12.54 34.185 12.605 34.25 ;
        RECT  12.54 34.185 12.605 34.25 ;
        RECT  12.54 34.185 12.605 34.25 ;
        RECT  12.54 34.185 12.605 34.25 ;
        RECT  12.54 34.185 12.605 34.25 ;
        RECT  12.54 34.185 12.605 34.25 ;
        RECT  12.54 34.185 12.605 34.25 ;
        RECT  12.54 34.185 12.605 34.25 ;
        RECT  12.09 34.6775 12.155 34.7425 ;
        RECT  11.835 34.185 11.9 34.25 ;
        RECT  11.835 34.185 11.9 34.25 ;
        RECT  11.835 34.185 11.9 34.25 ;
        RECT  11.835 34.185 11.9 34.25 ;
        RECT  11.835 34.185 11.9 34.25 ;
        RECT  11.835 34.185 11.9 34.25 ;
        RECT  12.54 34.185 12.605 34.25 ;
        RECT  12.54 34.185 12.605 34.25 ;
        RECT  12.54 34.185 12.605 34.25 ;
        RECT  12.54 34.185 12.605 34.25 ;
        RECT  12.285 34.6775 12.35 34.7425 ;
        RECT  12.54 35.0025 12.605 35.0675 ;
        RECT  12.54 35.0025 12.605 35.0675 ;
        RECT  12.54 35.0025 12.605 35.0675 ;
        RECT  12.54 34.185 12.605 34.25 ;
        RECT  12.54 34.185 12.605 34.25 ;
        RECT  12.54 34.185 12.605 34.25 ;
        RECT  12.54 34.185 12.605 34.25 ;
        RECT  12.54 34.185 12.605 34.25 ;
        RECT  12.54 34.185 12.605 34.25 ;
        RECT  11.835 35.0025 11.9 35.0675 ;
        RECT  12.54 35.82 12.605 35.885 ;
        RECT  12.54 35.82 12.605 35.885 ;
        RECT  12.54 35.82 12.605 35.885 ;
        RECT  12.54 35.82 12.605 35.885 ;
        RECT  12.54 35.82 12.605 35.885 ;
        RECT  12.54 35.82 12.605 35.885 ;
        RECT  11.835 35.0025 11.9 35.0675 ;
        RECT  12.54 35.0025 12.605 35.0675 ;
        RECT  12.54 35.82 12.605 35.885 ;
        RECT  12.54 35.82 12.605 35.885 ;
        RECT  12.54 35.82 12.605 35.885 ;
        RECT  12.54 35.82 12.605 35.885 ;
        RECT  12.54 35.82 12.605 35.885 ;
        RECT  12.54 35.82 12.605 35.885 ;
        RECT  12.54 35.82 12.605 35.885 ;
        RECT  12.54 35.82 12.605 35.885 ;
        RECT  12.09 35.3275 12.155 35.3925 ;
        RECT  11.835 35.82 11.9 35.885 ;
        RECT  11.835 35.82 11.9 35.885 ;
        RECT  11.835 35.82 11.9 35.885 ;
        RECT  11.835 35.82 11.9 35.885 ;
        RECT  11.835 35.82 11.9 35.885 ;
        RECT  11.835 35.82 11.9 35.885 ;
        RECT  12.54 35.82 12.605 35.885 ;
        RECT  12.54 35.82 12.605 35.885 ;
        RECT  12.54 35.82 12.605 35.885 ;
        RECT  12.54 35.82 12.605 35.885 ;
        RECT  12.285 35.3275 12.35 35.3925 ;
        RECT  12.54 35.0025 12.605 35.0675 ;
        RECT  12.54 35.0025 12.605 35.0675 ;
        RECT  12.54 35.0025 12.605 35.0675 ;
        RECT  12.54 35.82 12.605 35.885 ;
        RECT  12.54 35.82 12.605 35.885 ;
        RECT  12.54 35.82 12.605 35.885 ;
        RECT  12.54 35.82 12.605 35.885 ;
        RECT  12.54 35.82 12.605 35.885 ;
        RECT  12.54 35.82 12.605 35.885 ;
        RECT  11.835 35.0025 11.9 35.0675 ;
        RECT  12.54 36.875 12.605 36.94 ;
        RECT  12.54 36.875 12.605 36.94 ;
        RECT  12.54 36.875 12.605 36.94 ;
        RECT  12.54 36.875 12.605 36.94 ;
        RECT  12.54 36.875 12.605 36.94 ;
        RECT  12.54 36.875 12.605 36.94 ;
        RECT  11.835 37.6925 11.9 37.7575 ;
        RECT  12.54 37.6925 12.605 37.7575 ;
        RECT  12.54 36.875 12.605 36.94 ;
        RECT  12.54 36.875 12.605 36.94 ;
        RECT  12.54 36.875 12.605 36.94 ;
        RECT  12.54 36.875 12.605 36.94 ;
        RECT  12.54 36.875 12.605 36.94 ;
        RECT  12.54 36.875 12.605 36.94 ;
        RECT  12.54 36.875 12.605 36.94 ;
        RECT  12.54 36.875 12.605 36.94 ;
        RECT  12.09 37.3675 12.155 37.4325 ;
        RECT  11.835 36.875 11.9 36.94 ;
        RECT  11.835 36.875 11.9 36.94 ;
        RECT  11.835 36.875 11.9 36.94 ;
        RECT  11.835 36.875 11.9 36.94 ;
        RECT  11.835 36.875 11.9 36.94 ;
        RECT  11.835 36.875 11.9 36.94 ;
        RECT  12.54 36.875 12.605 36.94 ;
        RECT  12.54 36.875 12.605 36.94 ;
        RECT  12.54 36.875 12.605 36.94 ;
        RECT  12.54 36.875 12.605 36.94 ;
        RECT  12.285 37.3675 12.35 37.4325 ;
        RECT  12.54 37.6925 12.605 37.7575 ;
        RECT  12.54 37.6925 12.605 37.7575 ;
        RECT  12.54 37.6925 12.605 37.7575 ;
        RECT  12.54 36.875 12.605 36.94 ;
        RECT  12.54 36.875 12.605 36.94 ;
        RECT  12.54 36.875 12.605 36.94 ;
        RECT  12.54 36.875 12.605 36.94 ;
        RECT  12.54 36.875 12.605 36.94 ;
        RECT  12.54 36.875 12.605 36.94 ;
        RECT  11.835 37.6925 11.9 37.7575 ;
        RECT  12.54 38.51 12.605 38.575 ;
        RECT  12.54 38.51 12.605 38.575 ;
        RECT  12.54 38.51 12.605 38.575 ;
        RECT  12.54 38.51 12.605 38.575 ;
        RECT  12.54 38.51 12.605 38.575 ;
        RECT  12.54 38.51 12.605 38.575 ;
        RECT  11.835 37.6925 11.9 37.7575 ;
        RECT  12.54 37.6925 12.605 37.7575 ;
        RECT  12.54 38.51 12.605 38.575 ;
        RECT  12.54 38.51 12.605 38.575 ;
        RECT  12.54 38.51 12.605 38.575 ;
        RECT  12.54 38.51 12.605 38.575 ;
        RECT  12.54 38.51 12.605 38.575 ;
        RECT  12.54 38.51 12.605 38.575 ;
        RECT  12.54 38.51 12.605 38.575 ;
        RECT  12.54 38.51 12.605 38.575 ;
        RECT  12.09 38.0175 12.155 38.0825 ;
        RECT  11.835 38.51 11.9 38.575 ;
        RECT  11.835 38.51 11.9 38.575 ;
        RECT  11.835 38.51 11.9 38.575 ;
        RECT  11.835 38.51 11.9 38.575 ;
        RECT  11.835 38.51 11.9 38.575 ;
        RECT  11.835 38.51 11.9 38.575 ;
        RECT  12.54 38.51 12.605 38.575 ;
        RECT  12.54 38.51 12.605 38.575 ;
        RECT  12.54 38.51 12.605 38.575 ;
        RECT  12.54 38.51 12.605 38.575 ;
        RECT  12.285 38.0175 12.35 38.0825 ;
        RECT  12.54 37.6925 12.605 37.7575 ;
        RECT  12.54 37.6925 12.605 37.7575 ;
        RECT  12.54 37.6925 12.605 37.7575 ;
        RECT  12.54 38.51 12.605 38.575 ;
        RECT  12.54 38.51 12.605 38.575 ;
        RECT  12.54 38.51 12.605 38.575 ;
        RECT  12.54 38.51 12.605 38.575 ;
        RECT  12.54 38.51 12.605 38.575 ;
        RECT  12.54 38.51 12.605 38.575 ;
        RECT  11.835 37.6925 11.9 37.7575 ;
        RECT  12.54 39.565 12.605 39.63 ;
        RECT  12.54 39.565 12.605 39.63 ;
        RECT  12.54 39.565 12.605 39.63 ;
        RECT  12.54 39.565 12.605 39.63 ;
        RECT  12.54 39.565 12.605 39.63 ;
        RECT  12.54 39.565 12.605 39.63 ;
        RECT  11.835 40.3825 11.9 40.4475 ;
        RECT  12.54 40.3825 12.605 40.4475 ;
        RECT  12.54 39.565 12.605 39.63 ;
        RECT  12.54 39.565 12.605 39.63 ;
        RECT  12.54 39.565 12.605 39.63 ;
        RECT  12.54 39.565 12.605 39.63 ;
        RECT  12.54 39.565 12.605 39.63 ;
        RECT  12.54 39.565 12.605 39.63 ;
        RECT  12.54 39.565 12.605 39.63 ;
        RECT  12.54 39.565 12.605 39.63 ;
        RECT  12.09 40.0575 12.155 40.1225 ;
        RECT  11.835 39.565 11.9 39.63 ;
        RECT  11.835 39.565 11.9 39.63 ;
        RECT  11.835 39.565 11.9 39.63 ;
        RECT  11.835 39.565 11.9 39.63 ;
        RECT  11.835 39.565 11.9 39.63 ;
        RECT  11.835 39.565 11.9 39.63 ;
        RECT  12.54 39.565 12.605 39.63 ;
        RECT  12.54 39.565 12.605 39.63 ;
        RECT  12.54 39.565 12.605 39.63 ;
        RECT  12.54 39.565 12.605 39.63 ;
        RECT  12.285 40.0575 12.35 40.1225 ;
        RECT  12.54 40.3825 12.605 40.4475 ;
        RECT  12.54 40.3825 12.605 40.4475 ;
        RECT  12.54 40.3825 12.605 40.4475 ;
        RECT  12.54 39.565 12.605 39.63 ;
        RECT  12.54 39.565 12.605 39.63 ;
        RECT  12.54 39.565 12.605 39.63 ;
        RECT  12.54 39.565 12.605 39.63 ;
        RECT  12.54 39.565 12.605 39.63 ;
        RECT  12.54 39.565 12.605 39.63 ;
        RECT  11.835 40.3825 11.9 40.4475 ;
        RECT  11.3575 41.3475 11.4225 41.4125 ;
        RECT  11.7375 41.3475 11.8025 41.4125 ;
        RECT  11.3575 40.8975 11.4225 40.9625 ;
        RECT  11.5475 40.8975 11.6125 40.9625 ;
        RECT  12.0625 41.3475 12.1275 41.4125 ;
        RECT  12.4425 41.3475 12.5075 41.4125 ;
        RECT  12.0625 40.8975 12.1275 40.9625 ;
        RECT  12.2525 40.8975 12.3175 40.9625 ;
        RECT  11.4775 18.5325 11.5425 18.5975 ;
        RECT  11.835 14.2925 11.9 14.3575 ;
        RECT  11.13 14.2925 11.195 14.3575 ;
        RECT  11.6725 17.075 11.7375 17.14 ;
        RECT  11.29 17.485 11.355 17.55 ;
        RECT  11.4825 18.3275 11.5475 18.3925 ;
        RECT  11.4825 16.185 11.5475 16.25 ;
        RECT  12.1825 18.5325 12.2475 18.5975 ;
        RECT  12.54 14.2925 12.605 14.3575 ;
        RECT  11.835 14.2925 11.9 14.3575 ;
        RECT  12.3775 17.075 12.4425 17.14 ;
        RECT  11.995 17.485 12.06 17.55 ;
        RECT  12.1875 18.3275 12.2525 18.3925 ;
        RECT  12.1875 16.185 12.2525 16.25 ;
        RECT  11.405 9.97 11.47 10.035 ;
        RECT  11.835 11.605 11.9 11.67 ;
        RECT  11.835 11.035 11.9 11.1 ;
        RECT  11.13 11.035 11.195 11.1 ;
        RECT  11.55 11.24 11.615 11.305 ;
        RECT  11.835 13.5325 11.9 13.5975 ;
        RECT  11.55 10.83 11.615 10.895 ;
        RECT  11.41 10.83 11.475 10.895 ;
        RECT  11.835 11.24 11.9 11.305 ;
        RECT  11.13 11.24 11.195 11.305 ;
        RECT  11.3025 10.2325 11.3675 10.2975 ;
        RECT  11.41 13.21 11.475 13.275 ;
        RECT  11.58 11.605 11.645 11.67 ;
        RECT  11.27 12.52 11.335 12.585 ;
        RECT  11.41 11.24 11.475 11.305 ;
        RECT  11.13 11.605 11.195 11.67 ;
        RECT  11.58 12.12 11.645 12.185 ;
        RECT  11.315 13.7425 11.38 13.8075 ;
        RECT  11.13 13.5325 11.195 13.5975 ;
        RECT  12.11 9.97 12.175 10.035 ;
        RECT  12.54 11.605 12.605 11.67 ;
        RECT  12.54 11.035 12.605 11.1 ;
        RECT  11.835 11.035 11.9 11.1 ;
        RECT  12.255 11.24 12.32 11.305 ;
        RECT  12.54 13.5325 12.605 13.5975 ;
        RECT  12.255 10.83 12.32 10.895 ;
        RECT  12.115 10.83 12.18 10.895 ;
        RECT  12.54 11.24 12.605 11.305 ;
        RECT  11.835 11.24 11.9 11.305 ;
        RECT  12.0075 10.2325 12.0725 10.2975 ;
        RECT  12.115 13.21 12.18 13.275 ;
        RECT  12.285 11.605 12.35 11.67 ;
        RECT  11.975 12.52 12.04 12.585 ;
        RECT  12.115 11.24 12.18 11.305 ;
        RECT  11.835 11.605 11.9 11.67 ;
        RECT  12.285 12.12 12.35 12.185 ;
        RECT  12.02 13.7425 12.085 13.8075 ;
        RECT  11.835 13.5325 11.9 13.5975 ;
        RECT  11.3275 9.1325 11.3925 9.1975 ;
        RECT  11.835 3.955 11.9 4.02 ;
        RECT  11.6925 8.0375 11.7575 8.1025 ;
        RECT  11.695 6.43 11.76 6.495 ;
        RECT  11.695 5.0325 11.76 5.0975 ;
        RECT  11.13 3.815 11.195 3.88 ;
        RECT  11.835 6.8925 11.9 6.9575 ;
        RECT  11.33 5.6975 11.395 5.7625 ;
        RECT  11.695 9.39 11.76 9.455 ;
        RECT  11.5175 8.88 11.5825 8.945 ;
        RECT  11.835 8.4675 11.9 8.5325 ;
        RECT  11.835 3.765 11.9 3.83 ;
        RECT  11.835 5.5075 11.9 5.5725 ;
        RECT  11.33 5.3075 11.395 5.3725 ;
        RECT  11.5175 5.3075 11.5825 5.3725 ;
        RECT  11.5175 5.92 11.5825 5.985 ;
        RECT  11.3275 8.2675 11.3925 8.3325 ;
        RECT  11.5175 8.2675 11.5825 8.3325 ;
        RECT  12.3425 9.1325 12.4075 9.1975 ;
        RECT  11.835 3.955 11.9 4.02 ;
        RECT  11.9775 8.0375 12.0425 8.1025 ;
        RECT  11.975 6.43 12.04 6.495 ;
        RECT  11.975 5.0325 12.04 5.0975 ;
        RECT  12.54 3.815 12.605 3.88 ;
        RECT  11.835 6.8925 11.9 6.9575 ;
        RECT  12.34 5.6975 12.405 5.7625 ;
        RECT  11.975 9.39 12.04 9.455 ;
        RECT  12.1525 8.88 12.2175 8.945 ;
        RECT  11.835 8.4675 11.9 8.5325 ;
        RECT  11.835 3.765 11.9 3.83 ;
        RECT  11.835 5.5075 11.9 5.5725 ;
        RECT  12.34 5.3075 12.405 5.3725 ;
        RECT  12.1525 5.3075 12.2175 5.3725 ;
        RECT  12.1525 5.92 12.2175 5.985 ;
        RECT  12.3425 8.2675 12.4075 8.3325 ;
        RECT  12.1525 8.2675 12.2175 8.3325 ;
        RECT  11.4825 5.18 11.5475 5.245 ;
        RECT  11.835 3.9275 11.9 3.9925 ;
        RECT  11.615 5.82 11.68 5.885 ;
        RECT  11.835 5.9875 11.9 6.0525 ;
        RECT  11.3075 5.7975 11.3725 5.8625 ;
        RECT  11.515 5.52 11.58 5.585 ;
        RECT  11.615 4.3125 11.68 4.3775 ;
        RECT  11.27 4.08 11.335 4.145 ;
        RECT  12.1875 5.18 12.2525 5.245 ;
        RECT  11.835 3.9275 11.9 3.9925 ;
        RECT  12.055 5.82 12.12 5.885 ;
        RECT  11.835 5.9875 11.9 6.0525 ;
        RECT  12.3625 5.7975 12.4275 5.8625 ;
        RECT  12.155 5.52 12.22 5.585 ;
        RECT  12.055 4.3125 12.12 4.3775 ;
        RECT  12.4 4.08 12.465 4.145 ;
        RECT  6.1925 9.1825 6.2575 9.2475 ;
        RECT  7.5575 8.66 7.6225 8.725 ;
        RECT  6.0175 9.5725 6.0825 9.6375 ;
        RECT  7.3825 10.095 7.4475 10.16 ;
        RECT  6.1925 8.975 6.2575 9.04 ;
        RECT  6.0175 8.445 6.0825 8.51 ;
        RECT  5.8425 9.78 5.9075 9.845 ;
        RECT  6.0175 10.31 6.0825 10.375 ;
        RECT  6.1925 11.665 6.2575 11.73 ;
        RECT  5.6675 11.135 5.7325 11.2 ;
        RECT  5.8425 12.47 5.9075 12.535 ;
        RECT  7.5575 12.47 7.6225 12.535 ;
        RECT  5.6675 13.0 5.7325 13.065 ;
        RECT  7.3825 13.0 7.4475 13.065 ;
        RECT  6.3675 8.0325 6.4325 8.0975 ;
        RECT  6.5425 9.3775 6.6075 9.4425 ;
        RECT  6.3675 10.7225 6.4325 10.7875 ;
        RECT  6.5425 12.0675 6.6075 12.1325 ;
        RECT  6.3675 13.235 6.4325 13.3 ;
        RECT  6.1925 14.5625 6.2575 14.6275 ;
        RECT  7.5575 14.04 7.6225 14.105 ;
        RECT  6.0175 14.9525 6.0825 15.0175 ;
        RECT  7.3825 15.475 7.4475 15.54 ;
        RECT  6.1925 14.355 6.2575 14.42 ;
        RECT  6.0175 13.825 6.0825 13.89 ;
        RECT  5.8425 15.16 5.9075 15.225 ;
        RECT  6.0175 15.69 6.0825 15.755 ;
        RECT  6.1925 17.045 6.2575 17.11 ;
        RECT  5.6675 16.515 5.7325 16.58 ;
        RECT  5.8425 17.85 5.9075 17.915 ;
        RECT  7.5575 17.85 7.6225 17.915 ;
        RECT  5.6675 18.38 5.7325 18.445 ;
        RECT  7.3825 18.38 7.4475 18.445 ;
        RECT  6.3675 13.4125 6.4325 13.4775 ;
        RECT  6.5425 14.7575 6.6075 14.8225 ;
        RECT  6.3675 16.1025 6.4325 16.1675 ;
        RECT  6.5425 17.4475 6.6075 17.5125 ;
        RECT  6.3675 18.615 6.4325 18.68 ;
        RECT  2.8575 8.73 2.9225 8.795 ;
        RECT  3.0325 10.165 3.0975 10.23 ;
        RECT  3.2075 11.42 3.2725 11.485 ;
        RECT  3.3825 12.855 3.4475 12.92 ;
        RECT  3.5575 14.11 3.6225 14.175 ;
        RECT  3.7325 15.545 3.7975 15.61 ;
        RECT  3.9075 16.8 3.9725 16.865 ;
        RECT  4.0825 18.235 4.1475 18.3 ;
        RECT  2.8575 19.805 2.9225 19.87 ;
        RECT  3.5575 19.275 3.6225 19.34 ;
        RECT  2.8575 20.61 2.9225 20.675 ;
        RECT  3.7325 21.14 3.7975 21.205 ;
        RECT  2.8575 22.495 2.9225 22.56 ;
        RECT  3.9075 21.965 3.9725 22.03 ;
        RECT  2.8575 23.3 2.9225 23.365 ;
        RECT  4.0825 23.83 4.1475 23.895 ;
        RECT  3.0325 25.185 3.0975 25.25 ;
        RECT  3.5575 24.655 3.6225 24.72 ;
        RECT  3.0325 25.99 3.0975 26.055 ;
        RECT  3.7325 26.52 3.7975 26.585 ;
        RECT  3.0325 27.875 3.0975 27.94 ;
        RECT  3.9075 27.345 3.9725 27.41 ;
        RECT  3.0325 28.68 3.0975 28.745 ;
        RECT  4.0825 29.21 4.1475 29.275 ;
        RECT  3.2075 30.565 3.2725 30.63 ;
        RECT  3.5575 30.035 3.6225 30.1 ;
        RECT  3.2075 31.37 3.2725 31.435 ;
        RECT  3.7325 31.9 3.7975 31.965 ;
        RECT  3.2075 33.255 3.2725 33.32 ;
        RECT  3.9075 32.725 3.9725 32.79 ;
        RECT  3.2075 34.06 3.2725 34.125 ;
        RECT  4.0825 34.59 4.1475 34.655 ;
        RECT  3.3825 35.945 3.4475 36.01 ;
        RECT  3.5575 35.415 3.6225 35.48 ;
        RECT  3.3825 36.75 3.4475 36.815 ;
        RECT  3.7325 37.28 3.7975 37.345 ;
        RECT  3.3825 38.635 3.4475 38.7 ;
        RECT  3.9075 38.105 3.9725 38.17 ;
        RECT  3.3825 39.44 3.4475 39.505 ;
        RECT  4.0825 39.97 4.1475 40.035 ;
        RECT  5.5275 20.2075 5.5925 20.2725 ;
        RECT  5.9825 20.2075 6.0475 20.2725 ;
        RECT  6.6125 19.8075 6.6775 19.8725 ;
        RECT  5.565 19.84 5.63 19.905 ;
        RECT  5.5275 21.5525 5.5925 21.6175 ;
        RECT  5.9825 21.5525 6.0475 21.6175 ;
        RECT  6.6125 20.6075 6.6775 20.6725 ;
        RECT  5.565 20.575 5.63 20.64 ;
        RECT  5.5275 22.8975 5.5925 22.9625 ;
        RECT  5.9825 22.8975 6.0475 22.9625 ;
        RECT  6.6125 22.4975 6.6775 22.5625 ;
        RECT  5.565 22.53 5.63 22.595 ;
        RECT  5.5275 24.2425 5.5925 24.3075 ;
        RECT  5.9825 24.2425 6.0475 24.3075 ;
        RECT  6.6125 23.2975 6.6775 23.3625 ;
        RECT  5.565 23.265 5.63 23.33 ;
        RECT  5.5275 25.5875 5.5925 25.6525 ;
        RECT  5.9825 25.5875 6.0475 25.6525 ;
        RECT  6.6125 25.1875 6.6775 25.2525 ;
        RECT  5.565 25.22 5.63 25.285 ;
        RECT  5.5275 26.9325 5.5925 26.9975 ;
        RECT  5.9825 26.9325 6.0475 26.9975 ;
        RECT  6.6125 25.9875 6.6775 26.0525 ;
        RECT  5.565 25.955 5.63 26.02 ;
        RECT  5.5275 28.2775 5.5925 28.3425 ;
        RECT  5.9825 28.2775 6.0475 28.3425 ;
        RECT  6.6125 27.8775 6.6775 27.9425 ;
        RECT  5.565 27.91 5.63 27.975 ;
        RECT  5.5275 29.6225 5.5925 29.6875 ;
        RECT  5.9825 29.6225 6.0475 29.6875 ;
        RECT  6.6125 28.6775 6.6775 28.7425 ;
        RECT  5.565 28.645 5.63 28.71 ;
        RECT  5.5275 30.9675 5.5925 31.0325 ;
        RECT  5.9825 30.9675 6.0475 31.0325 ;
        RECT  6.6125 30.5675 6.6775 30.6325 ;
        RECT  5.565 30.6 5.63 30.665 ;
        RECT  5.5275 32.3125 5.5925 32.3775 ;
        RECT  5.9825 32.3125 6.0475 32.3775 ;
        RECT  6.6125 31.3675 6.6775 31.4325 ;
        RECT  5.565 31.335 5.63 31.4 ;
        RECT  5.5275 33.6575 5.5925 33.7225 ;
        RECT  5.9825 33.6575 6.0475 33.7225 ;
        RECT  6.6125 33.2575 6.6775 33.3225 ;
        RECT  5.565 33.29 5.63 33.355 ;
        RECT  5.5275 35.0025 5.5925 35.0675 ;
        RECT  5.9825 35.0025 6.0475 35.0675 ;
        RECT  6.6125 34.0575 6.6775 34.1225 ;
        RECT  5.565 34.025 5.63 34.09 ;
        RECT  5.5275 36.3475 5.5925 36.4125 ;
        RECT  5.9825 36.3475 6.0475 36.4125 ;
        RECT  6.6125 35.9475 6.6775 36.0125 ;
        RECT  5.565 35.98 5.63 36.045 ;
        RECT  5.5275 37.6925 5.5925 37.7575 ;
        RECT  5.9825 37.6925 6.0475 37.7575 ;
        RECT  6.6125 36.7475 6.6775 36.8125 ;
        RECT  5.565 36.715 5.63 36.78 ;
        RECT  5.5275 39.0375 5.5925 39.1025 ;
        RECT  5.9825 39.0375 6.0475 39.1025 ;
        RECT  6.6125 38.6375 6.6775 38.7025 ;
        RECT  5.565 38.67 5.63 38.735 ;
        RECT  5.5275 40.3825 5.5925 40.4475 ;
        RECT  5.9825 40.3825 6.0475 40.4475 ;
        RECT  6.6125 39.4375 6.6775 39.5025 ;
        RECT  5.565 39.405 5.63 39.47 ;
        RECT  6.68 7.61 6.745 7.675 ;
        RECT  1.5025 7.1025 1.5675 7.1675 ;
        RECT  5.585 7.245 5.65 7.31 ;
        RECT  3.9775 7.2425 4.0425 7.3075 ;
        RECT  2.58 7.2425 2.645 7.3075 ;
        RECT  1.3625 7.8075 1.4275 7.8725 ;
        RECT  4.44 7.1025 4.505 7.1675 ;
        RECT  3.245 7.6075 3.31 7.6725 ;
        RECT  6.9375 7.2425 7.0025 7.3075 ;
        RECT  6.4275 7.42 6.4925 7.485 ;
        RECT  6.015 7.1025 6.08 7.1675 ;
        RECT  1.3125 7.1025 1.3775 7.1675 ;
        RECT  3.055 7.1025 3.12 7.1675 ;
        RECT  2.855 7.6075 2.92 7.6725 ;
        RECT  2.855 7.42 2.92 7.485 ;
        RECT  3.4675 7.42 3.5325 7.485 ;
        RECT  5.815 7.61 5.88 7.675 ;
        RECT  5.815 7.42 5.88 7.485 ;
        RECT  6.68 6.595 6.745 6.66 ;
        RECT  1.5025 7.1025 1.5675 7.1675 ;
        RECT  5.585 6.96 5.65 7.025 ;
        RECT  3.9775 6.9625 4.0425 7.0275 ;
        RECT  2.58 6.9625 2.645 7.0275 ;
        RECT  1.3625 6.3975 1.4275 6.4625 ;
        RECT  4.44 7.1025 4.505 7.1675 ;
        RECT  3.245 6.5975 3.31 6.6625 ;
        RECT  6.9375 6.9625 7.0025 7.0275 ;
        RECT  6.4275 6.785 6.4925 6.85 ;
        RECT  6.015 7.1025 6.08 7.1675 ;
        RECT  1.3125 7.1025 1.3775 7.1675 ;
        RECT  3.055 7.1025 3.12 7.1675 ;
        RECT  2.855 6.5975 2.92 6.6625 ;
        RECT  2.855 6.785 2.92 6.85 ;
        RECT  3.4675 6.785 3.5325 6.85 ;
        RECT  5.815 6.595 5.88 6.66 ;
        RECT  5.815 6.785 5.88 6.85 ;
        RECT  6.68 6.2 6.745 6.265 ;
        RECT  1.5025 5.6925 1.5675 5.7575 ;
        RECT  5.585 5.835 5.65 5.9 ;
        RECT  3.9775 5.8325 4.0425 5.8975 ;
        RECT  2.58 5.8325 2.645 5.8975 ;
        RECT  1.3625 6.3975 1.4275 6.4625 ;
        RECT  4.44 5.6925 4.505 5.7575 ;
        RECT  3.245 6.1975 3.31 6.2625 ;
        RECT  6.9375 5.8325 7.0025 5.8975 ;
        RECT  6.4275 6.01 6.4925 6.075 ;
        RECT  6.015 5.6925 6.08 5.7575 ;
        RECT  1.3125 5.6925 1.3775 5.7575 ;
        RECT  3.055 5.6925 3.12 5.7575 ;
        RECT  2.855 6.1975 2.92 6.2625 ;
        RECT  2.855 6.01 2.92 6.075 ;
        RECT  3.4675 6.01 3.5325 6.075 ;
        RECT  5.815 6.2 5.88 6.265 ;
        RECT  5.815 6.01 5.88 6.075 ;
        RECT  6.68 5.185 6.745 5.25 ;
        RECT  1.5025 5.6925 1.5675 5.7575 ;
        RECT  5.585 5.55 5.65 5.615 ;
        RECT  3.9775 5.5525 4.0425 5.6175 ;
        RECT  2.58 5.5525 2.645 5.6175 ;
        RECT  1.3625 4.9875 1.4275 5.0525 ;
        RECT  4.44 5.6925 4.505 5.7575 ;
        RECT  3.245 5.1875 3.31 5.2525 ;
        RECT  6.9375 5.5525 7.0025 5.6175 ;
        RECT  6.4275 5.375 6.4925 5.44 ;
        RECT  6.015 5.6925 6.08 5.7575 ;
        RECT  1.3125 5.6925 1.3775 5.7575 ;
        RECT  3.055 5.6925 3.12 5.7575 ;
        RECT  2.855 5.1875 2.92 5.2525 ;
        RECT  2.855 5.375 2.92 5.44 ;
        RECT  3.4675 5.375 3.5325 5.44 ;
        RECT  5.815 5.185 5.88 5.25 ;
        RECT  5.815 5.375 5.88 5.44 ;
        RECT  8.575 8.765 8.64 8.83 ;
        RECT  8.365 10.2 8.43 10.265 ;
        RECT  8.155 14.145 8.22 14.21 ;
        RECT  7.945 15.58 8.01 15.645 ;
        RECT  10.395 3.635 10.46 3.7 ;
        RECT  9.975 1.45 10.04 1.515 ;
        RECT  10.185 2.9975 10.25 3.0625 ;
        RECT  10.395 41.135 10.46 41.2 ;
        RECT  10.605 10.1375 10.67 10.2025 ;
        RECT  10.815 14.1625 10.88 14.2275 ;
        RECT  1.0475 7.63 1.1125 7.695 ;
        RECT  9.765 41.565 9.83 41.63 ;
        RECT  8.9225 40.58 8.9875 40.645 ;
        RECT  9.0625 40.58 9.1275 40.645 ;
        RECT  11.8375 40.5475 11.9025 40.6125 ;
        RECT  12.5425 40.5475 12.6075 40.6125 ;
        RECT  11.0625 40.5475 11.1275 40.6125 ;
        RECT  9.4175 0.39 9.4825 0.455 ;
        RECT  9.5575 0.39 9.6225 0.455 ;
        RECT  11.835 0.39 11.9 0.455 ;
        RECT  11.835 0.39 11.9 0.455 ;
        RECT  7.8225 21.555 7.8875 21.62 ;
        RECT  7.8225 24.245 7.8875 24.31 ;
        RECT  7.8225 26.935 7.8875 27.0 ;
        RECT  7.8225 29.625 7.8875 29.69 ;
        RECT  7.8225 32.315 7.8875 32.38 ;
        RECT  7.8225 35.005 7.8875 35.07 ;
        RECT  7.8225 37.695 7.8875 37.76 ;
        RECT  7.8225 40.385 7.8875 40.45 ;
        RECT  8.9225 13.4475 8.9875 13.5125 ;
        RECT  9.0625 13.4475 9.1275 13.5125 ;
        RECT  8.9225 18.8275 8.9875 18.8925 ;
        RECT  9.0625 18.8275 9.1275 18.8925 ;
        RECT  7.3475 7.81 7.4125 7.875 ;
        RECT  8.9225 7.8425 8.9875 7.9075 ;
        RECT  9.0625 7.8425 9.1275 7.9075 ;
        RECT  7.3475 6.4 7.4125 6.465 ;
        RECT  8.9225 6.4325 8.9875 6.4975 ;
        RECT  9.0625 6.4325 9.1275 6.4975 ;
        RECT  7.3475 6.4 7.4125 6.465 ;
        RECT  8.9225 6.4325 8.9875 6.4975 ;
        RECT  9.0625 6.4325 9.1275 6.4975 ;
        RECT  7.3475 4.99 7.4125 5.055 ;
        RECT  8.9225 5.0225 8.9875 5.0875 ;
        RECT  9.0625 5.0225 9.1275 5.0875 ;
        RECT  -5.565 14.0125 -5.5 14.0775 ;
        RECT  -5.0575 8.835 -4.9925 8.9 ;
        RECT  -5.2 12.9175 -5.135 12.9825 ;
        RECT  -5.1975 11.31 -5.1325 11.375 ;
        RECT  -5.1975 9.9125 -5.1325 9.9775 ;
        RECT  -5.7625 8.695 -5.6975 8.76 ;
        RECT  -5.0575 11.7725 -4.9925 11.8375 ;
        RECT  -5.5625 10.5775 -5.4975 10.6425 ;
        RECT  -5.1975 14.27 -5.1325 14.335 ;
        RECT  -5.375 13.76 -5.31 13.825 ;
        RECT  -5.0575 13.3475 -4.9925 13.4125 ;
        RECT  -5.0575 8.645 -4.9925 8.71 ;
        RECT  -5.0575 10.3875 -4.9925 10.4525 ;
        RECT  -5.5625 10.1875 -5.4975 10.2525 ;
        RECT  -5.375 10.1875 -5.31 10.2525 ;
        RECT  -5.375 10.8 -5.31 10.865 ;
        RECT  -5.565 13.1475 -5.5 13.2125 ;
        RECT  -5.375 13.1475 -5.31 13.2125 ;
        RECT  -4.55 14.0125 -4.485 14.0775 ;
        RECT  -5.0575 8.835 -4.9925 8.9 ;
        RECT  -4.915 12.9175 -4.85 12.9825 ;
        RECT  -4.9175 11.31 -4.8525 11.375 ;
        RECT  -4.9175 9.9125 -4.8525 9.9775 ;
        RECT  -4.3525 8.695 -4.2875 8.76 ;
        RECT  -5.0575 11.7725 -4.9925 11.8375 ;
        RECT  -4.5525 10.5775 -4.4875 10.6425 ;
        RECT  -4.9175 14.27 -4.8525 14.335 ;
        RECT  -4.74 13.76 -4.675 13.825 ;
        RECT  -5.0575 13.3475 -4.9925 13.4125 ;
        RECT  -5.0575 8.645 -4.9925 8.71 ;
        RECT  -5.0575 10.3875 -4.9925 10.4525 ;
        RECT  -4.5525 10.1875 -4.4875 10.2525 ;
        RECT  -4.74 10.1875 -4.675 10.2525 ;
        RECT  -4.74 10.8 -4.675 10.865 ;
        RECT  -4.55 13.1475 -4.485 13.2125 ;
        RECT  -4.74 13.1475 -4.675 13.2125 ;
        RECT  -4.155 14.0125 -4.09 14.0775 ;
        RECT  -3.6475 8.835 -3.5825 8.9 ;
        RECT  -3.79 12.9175 -3.725 12.9825 ;
        RECT  -3.7875 11.31 -3.7225 11.375 ;
        RECT  -3.7875 9.9125 -3.7225 9.9775 ;
        RECT  -4.3525 8.695 -4.2875 8.76 ;
        RECT  -3.6475 11.7725 -3.5825 11.8375 ;
        RECT  -4.1525 10.5775 -4.0875 10.6425 ;
        RECT  -3.7875 14.27 -3.7225 14.335 ;
        RECT  -3.965 13.76 -3.9 13.825 ;
        RECT  -3.6475 13.3475 -3.5825 13.4125 ;
        RECT  -3.6475 8.645 -3.5825 8.71 ;
        RECT  -3.6475 10.3875 -3.5825 10.4525 ;
        RECT  -4.1525 10.1875 -4.0875 10.2525 ;
        RECT  -3.965 10.1875 -3.9 10.2525 ;
        RECT  -3.965 10.8 -3.9 10.865 ;
        RECT  -4.155 13.1475 -4.09 13.2125 ;
        RECT  -3.965 13.1475 -3.9 13.2125 ;
        RECT  -1.3775 8.8425 -1.3125 8.9075 ;
        RECT  -0.7975 8.8425 -0.7325 8.9075 ;
        RECT  -1.0025 23.865 -0.9375 23.93 ;
        RECT  -1.0025 23.305 -0.9375 23.37 ;
        RECT  -2.5225 22.88 -2.4575 22.945 ;
        RECT  -2.5225 23.44 -2.4575 23.505 ;
        RECT  -1.0025 23.5425 -0.9375 23.6075 ;
        RECT  -1.0025 22.9825 -0.9375 23.0475 ;
        RECT  -2.5225 23.2025 -2.4575 23.2675 ;
        RECT  -4.2275 23.0725 -4.1625 23.1375 ;
        RECT  -4.9325 23.5475 -4.8675 23.6125 ;
        RECT  -4.2275 23.5475 -4.1625 23.6125 ;
        RECT  -4.68 23.0675 -4.615 23.1325 ;
        RECT  -4.48 23.0725 -4.415 23.1375 ;
        RECT  -4.9325 22.7425 -4.8675 22.8075 ;
        RECT  -4.2275 22.7425 -4.1625 22.8075 ;
        RECT  -4.9325 21.925 -4.8675 21.99 ;
        RECT  -4.9325 21.925 -4.8675 21.99 ;
        RECT  -4.9325 21.925 -4.8675 21.99 ;
        RECT  -4.9325 21.925 -4.8675 21.99 ;
        RECT  -4.9325 21.925 -4.8675 21.99 ;
        RECT  -4.9325 21.925 -4.8675 21.99 ;
        RECT  -4.2275 22.7425 -4.1625 22.8075 ;
        RECT  -4.9325 22.7425 -4.8675 22.8075 ;
        RECT  -4.9325 21.925 -4.8675 21.99 ;
        RECT  -4.9325 21.925 -4.8675 21.99 ;
        RECT  -4.9325 21.925 -4.8675 21.99 ;
        RECT  -4.9325 21.925 -4.8675 21.99 ;
        RECT  -4.9325 21.925 -4.8675 21.99 ;
        RECT  -4.9325 21.925 -4.8675 21.99 ;
        RECT  -4.9325 21.925 -4.8675 21.99 ;
        RECT  -4.9325 21.925 -4.8675 21.99 ;
        RECT  -4.4825 22.4175 -4.4175 22.4825 ;
        RECT  -4.2275 21.925 -4.1625 21.99 ;
        RECT  -4.2275 21.925 -4.1625 21.99 ;
        RECT  -4.2275 21.925 -4.1625 21.99 ;
        RECT  -4.2275 21.925 -4.1625 21.99 ;
        RECT  -4.2275 21.925 -4.1625 21.99 ;
        RECT  -4.2275 21.925 -4.1625 21.99 ;
        RECT  -4.9325 21.925 -4.8675 21.99 ;
        RECT  -4.9325 21.925 -4.8675 21.99 ;
        RECT  -4.9325 21.925 -4.8675 21.99 ;
        RECT  -4.9325 21.925 -4.8675 21.99 ;
        RECT  -4.6775 22.4175 -4.6125 22.4825 ;
        RECT  -4.9325 22.7425 -4.8675 22.8075 ;
        RECT  -4.9325 22.7425 -4.8675 22.8075 ;
        RECT  -4.9325 22.7425 -4.8675 22.8075 ;
        RECT  -4.9325 21.925 -4.8675 21.99 ;
        RECT  -4.9325 21.925 -4.8675 21.99 ;
        RECT  -4.9325 21.925 -4.8675 21.99 ;
        RECT  -4.9325 21.925 -4.8675 21.99 ;
        RECT  -4.9325 21.925 -4.8675 21.99 ;
        RECT  -4.9325 21.925 -4.8675 21.99 ;
        RECT  -4.2275 22.7425 -4.1625 22.8075 ;
        RECT  -4.9325 20.87 -4.8675 20.935 ;
        RECT  -4.9325 20.87 -4.8675 20.935 ;
        RECT  -4.9325 20.87 -4.8675 20.935 ;
        RECT  -4.9325 20.87 -4.8675 20.935 ;
        RECT  -4.9325 20.87 -4.8675 20.935 ;
        RECT  -4.9325 20.87 -4.8675 20.935 ;
        RECT  -4.2275 20.0525 -4.1625 20.1175 ;
        RECT  -4.9325 20.0525 -4.8675 20.1175 ;
        RECT  -4.9325 20.87 -4.8675 20.935 ;
        RECT  -4.9325 20.87 -4.8675 20.935 ;
        RECT  -4.9325 20.87 -4.8675 20.935 ;
        RECT  -4.9325 20.87 -4.8675 20.935 ;
        RECT  -4.9325 20.87 -4.8675 20.935 ;
        RECT  -4.9325 20.87 -4.8675 20.935 ;
        RECT  -4.9325 20.87 -4.8675 20.935 ;
        RECT  -4.9325 20.87 -4.8675 20.935 ;
        RECT  -4.4825 20.3775 -4.4175 20.4425 ;
        RECT  -4.2275 20.87 -4.1625 20.935 ;
        RECT  -4.2275 20.87 -4.1625 20.935 ;
        RECT  -4.2275 20.87 -4.1625 20.935 ;
        RECT  -4.2275 20.87 -4.1625 20.935 ;
        RECT  -4.2275 20.87 -4.1625 20.935 ;
        RECT  -4.2275 20.87 -4.1625 20.935 ;
        RECT  -4.9325 20.87 -4.8675 20.935 ;
        RECT  -4.9325 20.87 -4.8675 20.935 ;
        RECT  -4.9325 20.87 -4.8675 20.935 ;
        RECT  -4.9325 20.87 -4.8675 20.935 ;
        RECT  -4.6775 20.3775 -4.6125 20.4425 ;
        RECT  -4.9325 20.0525 -4.8675 20.1175 ;
        RECT  -4.9325 20.0525 -4.8675 20.1175 ;
        RECT  -4.9325 20.0525 -4.8675 20.1175 ;
        RECT  -4.9325 20.87 -4.8675 20.935 ;
        RECT  -4.9325 20.87 -4.8675 20.935 ;
        RECT  -4.9325 20.87 -4.8675 20.935 ;
        RECT  -4.9325 20.87 -4.8675 20.935 ;
        RECT  -4.9325 20.87 -4.8675 20.935 ;
        RECT  -4.9325 20.87 -4.8675 20.935 ;
        RECT  -4.2275 20.0525 -4.1625 20.1175 ;
        RECT  -1.9775 21.2125 -1.9125 21.2775 ;
        RECT  -1.3825 21.07 -1.3175 21.135 ;
        RECT  -2.1375 21.07 -2.0725 21.135 ;
        RECT  -4.4125 21.0975 -4.3475 21.1625 ;
        RECT  -0.65 23.4425 -0.585 23.5075 ;
        RECT  -2.5575 23.4425 -2.4925 23.5075 ;
        RECT  -2.5925 24.2375 -2.5275 24.3025 ;
        RECT  -0.65 21.4 -0.585 21.465 ;
        RECT  -4.0275 22.4675 -3.9625 22.5325 ;
        RECT  -3.7375 21.9725 -3.6725 22.0375 ;
        RECT  -3.7375 23.7325 -3.6725 23.7975 ;
        RECT  -0.4175 20.6275 -0.3525 20.6925 ;
        RECT  -0.4175 25.1225 -0.3525 25.1875 ;
        RECT  -3.1075 25.1225 -3.0425 25.1875 ;
        RECT  -3.7725 26.3025 -3.7075 26.3675 ;
        RECT  -3.5275 23.895 -3.4625 23.96 ;
        RECT  -3.5275 22.8125 -3.4625 22.8775 ;
        RECT  -3.7375 24.0175 -3.6725 24.0825 ;
        RECT  -3.5275 23.895 -3.4625 23.96 ;
        RECT  -3.5275 25.2225 -3.4625 25.2875 ;
        RECT  -3.7375 21.3275 -3.6725 21.3925 ;
        RECT  -4.9325 20.6275 -4.8675 20.6925 ;
        RECT  -4.2275 20.6275 -4.1625 20.6925 ;
        RECT  -2.0775 16.6075 -2.0125 16.6725 ;
        RECT  -2.0775 16.9875 -2.0125 17.0525 ;
        RECT  -2.6775 16.6625 -2.6125 16.7275 ;
        RECT  -2.715 16.25 -2.65 16.315 ;
        RECT  -2.6775 16.8525 -2.6125 16.9175 ;
        RECT  -2.855 16.25 -2.79 16.315 ;
        RECT  -4.2025 16.6075 -4.1375 16.6725 ;
        RECT  -4.2025 16.9875 -4.1375 17.0525 ;
        RECT  -3.6025 16.6625 -3.5375 16.7275 ;
        RECT  -3.5 16.25 -3.435 16.315 ;
        RECT  -3.6025 16.8525 -3.5375 16.9175 ;
        RECT  -3.36 16.25 -3.295 16.315 ;
        RECT  -3.9975 14.65 -3.9325 14.715 ;
        RECT  -3.9975 15.14 -3.9325 15.205 ;
        RECT  -4.1525 14.65 -4.0875 14.715 ;
        RECT  -4.1525 15.35 -4.0875 15.415 ;
        RECT  -5.5625 14.65 -5.4975 14.715 ;
        RECT  -5.5625 15.56 -5.4975 15.625 ;
        RECT  -4.5475 14.65 -4.4825 14.715 ;
        RECT  -4.5475 15.77 -4.4825 15.835 ;
        RECT  -1.325 15.35 -1.26 15.415 ;
        RECT  -0.795 15.98 -0.73 16.045 ;
        RECT  -2.12 15.98 -2.055 16.045 ;
        RECT  -2.6425 15.35 -2.5775 15.415 ;
        RECT  -2.7825 15.56 -2.7175 15.625 ;
        RECT  -4.025 15.98 -3.96 16.045 ;
        RECT  -3.5025 15.77 -3.4375 15.835 ;
        RECT  -3.3625 15.56 -3.2975 15.625 ;
        RECT  -0.9975 9.8525 -0.9325 9.9175 ;
        RECT  -0.22 9.8525 -0.155 9.9175 ;
        RECT  -0.22 15.1375 -0.155 15.2025 ;
        RECT  -2.49 19.44 -2.425 19.505 ;
        RECT  -3.655 19.23 -3.59 19.295 ;
        RECT  -0.965 19.65 -0.9 19.715 ;
        RECT  -0.205 19.4375 -0.14 19.5025 ;
        RECT  -1.7275 19.86 -1.6625 19.925 ;
        RECT  -4.4175 19.86 -4.3525 19.925 ;
        RECT  -0.3825 14.93 -0.3175 14.995 ;
        RECT  -0.965 13.4125 -0.9 13.4775 ;
        RECT  -2.085 13.4125 -2.02 13.4775 ;
        RECT  -2.0825 8.31 -2.0175 8.375 ;
        RECT  -0.865 8.45 -0.8 8.515 ;
        RECT  -1.0475 16.8675 -0.9825 16.9325 ;
        RECT  -1.0 17.3375 -0.935 17.4025 ;
        RECT  0.0325 19.89 0.0975 19.955 ;
        RECT  0.1725 19.89 0.2375 19.955 ;
        LAYER  metal2 ;
        RECT  -0.35 19.855 0.0325 19.925 ;
        RECT  8.9225 0.0 9.6225 41.725 ;
        RECT  10.8125 0.0 10.8825 41.725 ;
        RECT  10.6025 0.0 10.6725 41.725 ;
        RECT  10.3925 0.0 10.4625 41.725 ;
        RECT  10.1825 0.0 10.2525 41.725 ;
        RECT  9.9725 0.0 10.0425 41.725 ;
        RECT  9.7625 0.0 9.8325 41.725 ;
        RECT  8.5725 5.02 8.6425 18.615 ;
        RECT  8.3625 5.02 8.4325 18.615 ;
        RECT  8.1525 5.02 8.2225 18.615 ;
        RECT  7.9425 5.02 8.0125 18.615 ;
        RECT  11.3125 40.415 11.3825 40.765 ;
        RECT  11.6475 40.415 11.7175 40.765 ;
        RECT  12.0175 40.415 12.0875 40.765 ;
        RECT  12.3525 40.415 12.4225 40.765 ;
        RECT  11.48 0.2775 11.55 0.3475 ;
        RECT  11.305 0.2775 11.515 0.3475 ;
        RECT  11.48 0.3125 11.55 0.54 ;
        RECT  12.185 0.2775 12.255 0.3475 ;
        RECT  12.01 0.2775 12.22 0.3475 ;
        RECT  12.185 0.3125 12.255 0.54 ;
        RECT  10.3925 18.895 10.4625 41.24 ;
        RECT  11.8325 40.415 11.9025 40.61 ;
        RECT  12.5375 40.415 12.6075 40.61 ;
        RECT  11.0925 18.895 11.1625 40.61 ;
        RECT  7.8875 21.5525 8.9225 21.6225 ;
        RECT  7.8875 24.2425 8.9225 24.3125 ;
        RECT  7.8875 26.9325 8.9225 27.0025 ;
        RECT  7.8875 29.6225 8.9225 29.6925 ;
        RECT  7.8875 32.3125 8.9225 32.3825 ;
        RECT  7.8875 35.0025 8.9225 35.0725 ;
        RECT  7.8875 37.6925 8.9225 37.7625 ;
        RECT  7.8875 40.3825 8.9225 40.4525 ;
        RECT  11.8325 19.645 11.9025 19.78 ;
        RECT  11.8325 19.645 11.9025 19.78 ;
        RECT  11.8325 19.645 11.9025 19.78 ;
        RECT  11.8325 19.645 11.9025 19.78 ;
        RECT  11.8325 19.645 11.9025 19.78 ;
        RECT  11.8325 19.645 11.9025 19.78 ;
        RECT  11.095 18.86 11.23 18.93 ;
        RECT  11.8 18.86 11.935 18.93 ;
        RECT  11.8325 19.645 11.9025 19.78 ;
        RECT  11.8325 19.645 11.9025 19.78 ;
        RECT  11.8325 19.645 11.9025 19.78 ;
        RECT  11.8325 19.645 11.9025 19.78 ;
        RECT  11.8325 19.645 11.9025 19.78 ;
        RECT  11.8325 19.645 11.9025 19.78 ;
        RECT  11.8325 19.645 11.9025 19.78 ;
        RECT  11.8325 19.645 11.9025 19.78 ;
        RECT  11.3825 19.1525 11.4525 19.2875 ;
        RECT  11.1275 19.645 11.1975 19.78 ;
        RECT  11.1275 19.645 11.1975 19.78 ;
        RECT  11.1275 19.645 11.1975 19.78 ;
        RECT  11.1275 19.645 11.1975 19.78 ;
        RECT  11.1275 19.645 11.1975 19.78 ;
        RECT  11.1275 19.645 11.1975 19.78 ;
        RECT  11.8325 19.645 11.9025 19.78 ;
        RECT  11.8325 19.645 11.9025 19.78 ;
        RECT  11.8325 19.645 11.9025 19.78 ;
        RECT  11.8325 19.645 11.9025 19.78 ;
        RECT  11.5775 19.1525 11.6475 19.2875 ;
        RECT  11.8 18.86 11.935 18.93 ;
        RECT  11.8 18.86 11.935 18.93 ;
        RECT  11.8 18.86 11.935 18.93 ;
        RECT  11.8325 19.645 11.9025 19.78 ;
        RECT  11.8325 19.645 11.9025 19.78 ;
        RECT  11.8325 19.645 11.9025 19.78 ;
        RECT  11.8325 19.645 11.9025 19.78 ;
        RECT  11.8325 19.645 11.9025 19.78 ;
        RECT  11.8325 19.645 11.9025 19.78 ;
        RECT  11.095 18.86 11.23 18.93 ;
        RECT  11.8325 18.8625 11.9025 20.2725 ;
        RECT  11.1325 18.865 11.1925 18.9225 ;
        RECT  11.32 18.87 11.375 18.9225 ;
        RECT  11.655 18.8625 11.7125 18.9225 ;
        RECT  11.8375 18.87 11.8975 18.9275 ;
        RECT  11.6475 18.795 11.7175 20.34 ;
        RECT  11.3125 18.795 11.3825 20.34 ;
        RECT  11.1275 18.795 11.1975 20.34 ;
        RECT  11.8325 18.795 11.9025 20.34 ;
        RECT  11.8325 20.7 11.9025 20.835 ;
        RECT  11.8325 20.7 11.9025 20.835 ;
        RECT  11.8325 20.7 11.9025 20.835 ;
        RECT  11.8325 20.7 11.9025 20.835 ;
        RECT  11.8325 20.7 11.9025 20.835 ;
        RECT  11.8325 20.7 11.9025 20.835 ;
        RECT  11.095 21.55 11.23 21.62 ;
        RECT  11.8 21.55 11.935 21.62 ;
        RECT  11.8325 20.7 11.9025 20.835 ;
        RECT  11.8325 20.7 11.9025 20.835 ;
        RECT  11.8325 20.7 11.9025 20.835 ;
        RECT  11.8325 20.7 11.9025 20.835 ;
        RECT  11.8325 20.7 11.9025 20.835 ;
        RECT  11.8325 20.7 11.9025 20.835 ;
        RECT  11.8325 20.7 11.9025 20.835 ;
        RECT  11.8325 20.7 11.9025 20.835 ;
        RECT  11.3825 21.1925 11.4525 21.3275 ;
        RECT  11.1275 20.7 11.1975 20.835 ;
        RECT  11.1275 20.7 11.1975 20.835 ;
        RECT  11.1275 20.7 11.1975 20.835 ;
        RECT  11.1275 20.7 11.1975 20.835 ;
        RECT  11.1275 20.7 11.1975 20.835 ;
        RECT  11.1275 20.7 11.1975 20.835 ;
        RECT  11.8325 20.7 11.9025 20.835 ;
        RECT  11.8325 20.7 11.9025 20.835 ;
        RECT  11.8325 20.7 11.9025 20.835 ;
        RECT  11.8325 20.7 11.9025 20.835 ;
        RECT  11.5775 21.1925 11.6475 21.3275 ;
        RECT  11.8 21.55 11.935 21.62 ;
        RECT  11.8 21.55 11.935 21.62 ;
        RECT  11.8 21.55 11.935 21.62 ;
        RECT  11.8325 20.7 11.9025 20.835 ;
        RECT  11.8325 20.7 11.9025 20.835 ;
        RECT  11.8325 20.7 11.9025 20.835 ;
        RECT  11.8325 20.7 11.9025 20.835 ;
        RECT  11.8325 20.7 11.9025 20.835 ;
        RECT  11.8325 20.7 11.9025 20.835 ;
        RECT  11.095 21.55 11.23 21.62 ;
        RECT  11.8325 20.2075 11.9025 21.6175 ;
        RECT  11.1325 21.5575 11.1925 21.615 ;
        RECT  11.32 21.5575 11.375 21.61 ;
        RECT  11.655 21.5575 11.7125 21.6175 ;
        RECT  11.8375 21.5525 11.8975 21.61 ;
        RECT  11.6475 20.14 11.7175 21.685 ;
        RECT  11.3125 20.14 11.3825 21.685 ;
        RECT  11.1275 20.14 11.1975 21.685 ;
        RECT  11.8325 20.14 11.9025 21.685 ;
        RECT  11.8325 22.335 11.9025 22.47 ;
        RECT  11.8325 22.335 11.9025 22.47 ;
        RECT  11.8325 22.335 11.9025 22.47 ;
        RECT  11.8325 22.335 11.9025 22.47 ;
        RECT  11.8325 22.335 11.9025 22.47 ;
        RECT  11.8325 22.335 11.9025 22.47 ;
        RECT  11.095 21.55 11.23 21.62 ;
        RECT  11.8 21.55 11.935 21.62 ;
        RECT  11.8325 22.335 11.9025 22.47 ;
        RECT  11.8325 22.335 11.9025 22.47 ;
        RECT  11.8325 22.335 11.9025 22.47 ;
        RECT  11.8325 22.335 11.9025 22.47 ;
        RECT  11.8325 22.335 11.9025 22.47 ;
        RECT  11.8325 22.335 11.9025 22.47 ;
        RECT  11.8325 22.335 11.9025 22.47 ;
        RECT  11.8325 22.335 11.9025 22.47 ;
        RECT  11.3825 21.8425 11.4525 21.9775 ;
        RECT  11.1275 22.335 11.1975 22.47 ;
        RECT  11.1275 22.335 11.1975 22.47 ;
        RECT  11.1275 22.335 11.1975 22.47 ;
        RECT  11.1275 22.335 11.1975 22.47 ;
        RECT  11.1275 22.335 11.1975 22.47 ;
        RECT  11.1275 22.335 11.1975 22.47 ;
        RECT  11.8325 22.335 11.9025 22.47 ;
        RECT  11.8325 22.335 11.9025 22.47 ;
        RECT  11.8325 22.335 11.9025 22.47 ;
        RECT  11.8325 22.335 11.9025 22.47 ;
        RECT  11.5775 21.8425 11.6475 21.9775 ;
        RECT  11.8 21.55 11.935 21.62 ;
        RECT  11.8 21.55 11.935 21.62 ;
        RECT  11.8 21.55 11.935 21.62 ;
        RECT  11.8325 22.335 11.9025 22.47 ;
        RECT  11.8325 22.335 11.9025 22.47 ;
        RECT  11.8325 22.335 11.9025 22.47 ;
        RECT  11.8325 22.335 11.9025 22.47 ;
        RECT  11.8325 22.335 11.9025 22.47 ;
        RECT  11.8325 22.335 11.9025 22.47 ;
        RECT  11.095 21.55 11.23 21.62 ;
        RECT  11.8325 21.5525 11.9025 22.9625 ;
        RECT  11.1325 21.555 11.1925 21.6125 ;
        RECT  11.32 21.56 11.375 21.6125 ;
        RECT  11.655 21.5525 11.7125 21.6125 ;
        RECT  11.8375 21.56 11.8975 21.6175 ;
        RECT  11.6475 21.485 11.7175 23.03 ;
        RECT  11.3125 21.485 11.3825 23.03 ;
        RECT  11.1275 21.485 11.1975 23.03 ;
        RECT  11.8325 21.485 11.9025 23.03 ;
        RECT  11.8325 23.39 11.9025 23.525 ;
        RECT  11.8325 23.39 11.9025 23.525 ;
        RECT  11.8325 23.39 11.9025 23.525 ;
        RECT  11.8325 23.39 11.9025 23.525 ;
        RECT  11.8325 23.39 11.9025 23.525 ;
        RECT  11.8325 23.39 11.9025 23.525 ;
        RECT  11.095 24.24 11.23 24.31 ;
        RECT  11.8 24.24 11.935 24.31 ;
        RECT  11.8325 23.39 11.9025 23.525 ;
        RECT  11.8325 23.39 11.9025 23.525 ;
        RECT  11.8325 23.39 11.9025 23.525 ;
        RECT  11.8325 23.39 11.9025 23.525 ;
        RECT  11.8325 23.39 11.9025 23.525 ;
        RECT  11.8325 23.39 11.9025 23.525 ;
        RECT  11.8325 23.39 11.9025 23.525 ;
        RECT  11.8325 23.39 11.9025 23.525 ;
        RECT  11.3825 23.8825 11.4525 24.0175 ;
        RECT  11.1275 23.39 11.1975 23.525 ;
        RECT  11.1275 23.39 11.1975 23.525 ;
        RECT  11.1275 23.39 11.1975 23.525 ;
        RECT  11.1275 23.39 11.1975 23.525 ;
        RECT  11.1275 23.39 11.1975 23.525 ;
        RECT  11.1275 23.39 11.1975 23.525 ;
        RECT  11.8325 23.39 11.9025 23.525 ;
        RECT  11.8325 23.39 11.9025 23.525 ;
        RECT  11.8325 23.39 11.9025 23.525 ;
        RECT  11.8325 23.39 11.9025 23.525 ;
        RECT  11.5775 23.8825 11.6475 24.0175 ;
        RECT  11.8 24.24 11.935 24.31 ;
        RECT  11.8 24.24 11.935 24.31 ;
        RECT  11.8 24.24 11.935 24.31 ;
        RECT  11.8325 23.39 11.9025 23.525 ;
        RECT  11.8325 23.39 11.9025 23.525 ;
        RECT  11.8325 23.39 11.9025 23.525 ;
        RECT  11.8325 23.39 11.9025 23.525 ;
        RECT  11.8325 23.39 11.9025 23.525 ;
        RECT  11.8325 23.39 11.9025 23.525 ;
        RECT  11.095 24.24 11.23 24.31 ;
        RECT  11.8325 22.8975 11.9025 24.3075 ;
        RECT  11.1325 24.2475 11.1925 24.305 ;
        RECT  11.32 24.2475 11.375 24.3 ;
        RECT  11.655 24.2475 11.7125 24.3075 ;
        RECT  11.8375 24.2425 11.8975 24.3 ;
        RECT  11.6475 22.83 11.7175 24.375 ;
        RECT  11.3125 22.83 11.3825 24.375 ;
        RECT  11.1275 22.83 11.1975 24.375 ;
        RECT  11.8325 22.83 11.9025 24.375 ;
        RECT  11.8325 25.025 11.9025 25.16 ;
        RECT  11.8325 25.025 11.9025 25.16 ;
        RECT  11.8325 25.025 11.9025 25.16 ;
        RECT  11.8325 25.025 11.9025 25.16 ;
        RECT  11.8325 25.025 11.9025 25.16 ;
        RECT  11.8325 25.025 11.9025 25.16 ;
        RECT  11.095 24.24 11.23 24.31 ;
        RECT  11.8 24.24 11.935 24.31 ;
        RECT  11.8325 25.025 11.9025 25.16 ;
        RECT  11.8325 25.025 11.9025 25.16 ;
        RECT  11.8325 25.025 11.9025 25.16 ;
        RECT  11.8325 25.025 11.9025 25.16 ;
        RECT  11.8325 25.025 11.9025 25.16 ;
        RECT  11.8325 25.025 11.9025 25.16 ;
        RECT  11.8325 25.025 11.9025 25.16 ;
        RECT  11.8325 25.025 11.9025 25.16 ;
        RECT  11.3825 24.5325 11.4525 24.6675 ;
        RECT  11.1275 25.025 11.1975 25.16 ;
        RECT  11.1275 25.025 11.1975 25.16 ;
        RECT  11.1275 25.025 11.1975 25.16 ;
        RECT  11.1275 25.025 11.1975 25.16 ;
        RECT  11.1275 25.025 11.1975 25.16 ;
        RECT  11.1275 25.025 11.1975 25.16 ;
        RECT  11.8325 25.025 11.9025 25.16 ;
        RECT  11.8325 25.025 11.9025 25.16 ;
        RECT  11.8325 25.025 11.9025 25.16 ;
        RECT  11.8325 25.025 11.9025 25.16 ;
        RECT  11.5775 24.5325 11.6475 24.6675 ;
        RECT  11.8 24.24 11.935 24.31 ;
        RECT  11.8 24.24 11.935 24.31 ;
        RECT  11.8 24.24 11.935 24.31 ;
        RECT  11.8325 25.025 11.9025 25.16 ;
        RECT  11.8325 25.025 11.9025 25.16 ;
        RECT  11.8325 25.025 11.9025 25.16 ;
        RECT  11.8325 25.025 11.9025 25.16 ;
        RECT  11.8325 25.025 11.9025 25.16 ;
        RECT  11.8325 25.025 11.9025 25.16 ;
        RECT  11.095 24.24 11.23 24.31 ;
        RECT  11.8325 24.2425 11.9025 25.6525 ;
        RECT  11.1325 24.245 11.1925 24.3025 ;
        RECT  11.32 24.25 11.375 24.3025 ;
        RECT  11.655 24.2425 11.7125 24.3025 ;
        RECT  11.8375 24.25 11.8975 24.3075 ;
        RECT  11.6475 24.175 11.7175 25.72 ;
        RECT  11.3125 24.175 11.3825 25.72 ;
        RECT  11.1275 24.175 11.1975 25.72 ;
        RECT  11.8325 24.175 11.9025 25.72 ;
        RECT  11.8325 26.08 11.9025 26.215 ;
        RECT  11.8325 26.08 11.9025 26.215 ;
        RECT  11.8325 26.08 11.9025 26.215 ;
        RECT  11.8325 26.08 11.9025 26.215 ;
        RECT  11.8325 26.08 11.9025 26.215 ;
        RECT  11.8325 26.08 11.9025 26.215 ;
        RECT  11.095 26.93 11.23 27.0 ;
        RECT  11.8 26.93 11.935 27.0 ;
        RECT  11.8325 26.08 11.9025 26.215 ;
        RECT  11.8325 26.08 11.9025 26.215 ;
        RECT  11.8325 26.08 11.9025 26.215 ;
        RECT  11.8325 26.08 11.9025 26.215 ;
        RECT  11.8325 26.08 11.9025 26.215 ;
        RECT  11.8325 26.08 11.9025 26.215 ;
        RECT  11.8325 26.08 11.9025 26.215 ;
        RECT  11.8325 26.08 11.9025 26.215 ;
        RECT  11.3825 26.5725 11.4525 26.7075 ;
        RECT  11.1275 26.08 11.1975 26.215 ;
        RECT  11.1275 26.08 11.1975 26.215 ;
        RECT  11.1275 26.08 11.1975 26.215 ;
        RECT  11.1275 26.08 11.1975 26.215 ;
        RECT  11.1275 26.08 11.1975 26.215 ;
        RECT  11.1275 26.08 11.1975 26.215 ;
        RECT  11.8325 26.08 11.9025 26.215 ;
        RECT  11.8325 26.08 11.9025 26.215 ;
        RECT  11.8325 26.08 11.9025 26.215 ;
        RECT  11.8325 26.08 11.9025 26.215 ;
        RECT  11.5775 26.5725 11.6475 26.7075 ;
        RECT  11.8 26.93 11.935 27.0 ;
        RECT  11.8 26.93 11.935 27.0 ;
        RECT  11.8 26.93 11.935 27.0 ;
        RECT  11.8325 26.08 11.9025 26.215 ;
        RECT  11.8325 26.08 11.9025 26.215 ;
        RECT  11.8325 26.08 11.9025 26.215 ;
        RECT  11.8325 26.08 11.9025 26.215 ;
        RECT  11.8325 26.08 11.9025 26.215 ;
        RECT  11.8325 26.08 11.9025 26.215 ;
        RECT  11.095 26.93 11.23 27.0 ;
        RECT  11.8325 25.5875 11.9025 26.9975 ;
        RECT  11.1325 26.9375 11.1925 26.995 ;
        RECT  11.32 26.9375 11.375 26.99 ;
        RECT  11.655 26.9375 11.7125 26.9975 ;
        RECT  11.8375 26.9325 11.8975 26.99 ;
        RECT  11.6475 25.52 11.7175 27.065 ;
        RECT  11.3125 25.52 11.3825 27.065 ;
        RECT  11.1275 25.52 11.1975 27.065 ;
        RECT  11.8325 25.52 11.9025 27.065 ;
        RECT  11.8325 27.715 11.9025 27.85 ;
        RECT  11.8325 27.715 11.9025 27.85 ;
        RECT  11.8325 27.715 11.9025 27.85 ;
        RECT  11.8325 27.715 11.9025 27.85 ;
        RECT  11.8325 27.715 11.9025 27.85 ;
        RECT  11.8325 27.715 11.9025 27.85 ;
        RECT  11.095 26.93 11.23 27.0 ;
        RECT  11.8 26.93 11.935 27.0 ;
        RECT  11.8325 27.715 11.9025 27.85 ;
        RECT  11.8325 27.715 11.9025 27.85 ;
        RECT  11.8325 27.715 11.9025 27.85 ;
        RECT  11.8325 27.715 11.9025 27.85 ;
        RECT  11.8325 27.715 11.9025 27.85 ;
        RECT  11.8325 27.715 11.9025 27.85 ;
        RECT  11.8325 27.715 11.9025 27.85 ;
        RECT  11.8325 27.715 11.9025 27.85 ;
        RECT  11.3825 27.2225 11.4525 27.3575 ;
        RECT  11.1275 27.715 11.1975 27.85 ;
        RECT  11.1275 27.715 11.1975 27.85 ;
        RECT  11.1275 27.715 11.1975 27.85 ;
        RECT  11.1275 27.715 11.1975 27.85 ;
        RECT  11.1275 27.715 11.1975 27.85 ;
        RECT  11.1275 27.715 11.1975 27.85 ;
        RECT  11.8325 27.715 11.9025 27.85 ;
        RECT  11.8325 27.715 11.9025 27.85 ;
        RECT  11.8325 27.715 11.9025 27.85 ;
        RECT  11.8325 27.715 11.9025 27.85 ;
        RECT  11.5775 27.2225 11.6475 27.3575 ;
        RECT  11.8 26.93 11.935 27.0 ;
        RECT  11.8 26.93 11.935 27.0 ;
        RECT  11.8 26.93 11.935 27.0 ;
        RECT  11.8325 27.715 11.9025 27.85 ;
        RECT  11.8325 27.715 11.9025 27.85 ;
        RECT  11.8325 27.715 11.9025 27.85 ;
        RECT  11.8325 27.715 11.9025 27.85 ;
        RECT  11.8325 27.715 11.9025 27.85 ;
        RECT  11.8325 27.715 11.9025 27.85 ;
        RECT  11.095 26.93 11.23 27.0 ;
        RECT  11.8325 26.9325 11.9025 28.3425 ;
        RECT  11.1325 26.935 11.1925 26.9925 ;
        RECT  11.32 26.94 11.375 26.9925 ;
        RECT  11.655 26.9325 11.7125 26.9925 ;
        RECT  11.8375 26.94 11.8975 26.9975 ;
        RECT  11.6475 26.865 11.7175 28.41 ;
        RECT  11.3125 26.865 11.3825 28.41 ;
        RECT  11.1275 26.865 11.1975 28.41 ;
        RECT  11.8325 26.865 11.9025 28.41 ;
        RECT  11.8325 28.77 11.9025 28.905 ;
        RECT  11.8325 28.77 11.9025 28.905 ;
        RECT  11.8325 28.77 11.9025 28.905 ;
        RECT  11.8325 28.77 11.9025 28.905 ;
        RECT  11.8325 28.77 11.9025 28.905 ;
        RECT  11.8325 28.77 11.9025 28.905 ;
        RECT  11.095 29.62 11.23 29.69 ;
        RECT  11.8 29.62 11.935 29.69 ;
        RECT  11.8325 28.77 11.9025 28.905 ;
        RECT  11.8325 28.77 11.9025 28.905 ;
        RECT  11.8325 28.77 11.9025 28.905 ;
        RECT  11.8325 28.77 11.9025 28.905 ;
        RECT  11.8325 28.77 11.9025 28.905 ;
        RECT  11.8325 28.77 11.9025 28.905 ;
        RECT  11.8325 28.77 11.9025 28.905 ;
        RECT  11.8325 28.77 11.9025 28.905 ;
        RECT  11.3825 29.2625 11.4525 29.3975 ;
        RECT  11.1275 28.77 11.1975 28.905 ;
        RECT  11.1275 28.77 11.1975 28.905 ;
        RECT  11.1275 28.77 11.1975 28.905 ;
        RECT  11.1275 28.77 11.1975 28.905 ;
        RECT  11.1275 28.77 11.1975 28.905 ;
        RECT  11.1275 28.77 11.1975 28.905 ;
        RECT  11.8325 28.77 11.9025 28.905 ;
        RECT  11.8325 28.77 11.9025 28.905 ;
        RECT  11.8325 28.77 11.9025 28.905 ;
        RECT  11.8325 28.77 11.9025 28.905 ;
        RECT  11.5775 29.2625 11.6475 29.3975 ;
        RECT  11.8 29.62 11.935 29.69 ;
        RECT  11.8 29.62 11.935 29.69 ;
        RECT  11.8 29.62 11.935 29.69 ;
        RECT  11.8325 28.77 11.9025 28.905 ;
        RECT  11.8325 28.77 11.9025 28.905 ;
        RECT  11.8325 28.77 11.9025 28.905 ;
        RECT  11.8325 28.77 11.9025 28.905 ;
        RECT  11.8325 28.77 11.9025 28.905 ;
        RECT  11.8325 28.77 11.9025 28.905 ;
        RECT  11.095 29.62 11.23 29.69 ;
        RECT  11.8325 28.2775 11.9025 29.6875 ;
        RECT  11.1325 29.6275 11.1925 29.685 ;
        RECT  11.32 29.6275 11.375 29.68 ;
        RECT  11.655 29.6275 11.7125 29.6875 ;
        RECT  11.8375 29.6225 11.8975 29.68 ;
        RECT  11.6475 28.21 11.7175 29.755 ;
        RECT  11.3125 28.21 11.3825 29.755 ;
        RECT  11.1275 28.21 11.1975 29.755 ;
        RECT  11.8325 28.21 11.9025 29.755 ;
        RECT  11.8325 30.405 11.9025 30.54 ;
        RECT  11.8325 30.405 11.9025 30.54 ;
        RECT  11.8325 30.405 11.9025 30.54 ;
        RECT  11.8325 30.405 11.9025 30.54 ;
        RECT  11.8325 30.405 11.9025 30.54 ;
        RECT  11.8325 30.405 11.9025 30.54 ;
        RECT  11.095 29.62 11.23 29.69 ;
        RECT  11.8 29.62 11.935 29.69 ;
        RECT  11.8325 30.405 11.9025 30.54 ;
        RECT  11.8325 30.405 11.9025 30.54 ;
        RECT  11.8325 30.405 11.9025 30.54 ;
        RECT  11.8325 30.405 11.9025 30.54 ;
        RECT  11.8325 30.405 11.9025 30.54 ;
        RECT  11.8325 30.405 11.9025 30.54 ;
        RECT  11.8325 30.405 11.9025 30.54 ;
        RECT  11.8325 30.405 11.9025 30.54 ;
        RECT  11.3825 29.9125 11.4525 30.0475 ;
        RECT  11.1275 30.405 11.1975 30.54 ;
        RECT  11.1275 30.405 11.1975 30.54 ;
        RECT  11.1275 30.405 11.1975 30.54 ;
        RECT  11.1275 30.405 11.1975 30.54 ;
        RECT  11.1275 30.405 11.1975 30.54 ;
        RECT  11.1275 30.405 11.1975 30.54 ;
        RECT  11.8325 30.405 11.9025 30.54 ;
        RECT  11.8325 30.405 11.9025 30.54 ;
        RECT  11.8325 30.405 11.9025 30.54 ;
        RECT  11.8325 30.405 11.9025 30.54 ;
        RECT  11.5775 29.9125 11.6475 30.0475 ;
        RECT  11.8 29.62 11.935 29.69 ;
        RECT  11.8 29.62 11.935 29.69 ;
        RECT  11.8 29.62 11.935 29.69 ;
        RECT  11.8325 30.405 11.9025 30.54 ;
        RECT  11.8325 30.405 11.9025 30.54 ;
        RECT  11.8325 30.405 11.9025 30.54 ;
        RECT  11.8325 30.405 11.9025 30.54 ;
        RECT  11.8325 30.405 11.9025 30.54 ;
        RECT  11.8325 30.405 11.9025 30.54 ;
        RECT  11.095 29.62 11.23 29.69 ;
        RECT  11.8325 29.6225 11.9025 31.0325 ;
        RECT  11.1325 29.625 11.1925 29.6825 ;
        RECT  11.32 29.63 11.375 29.6825 ;
        RECT  11.655 29.6225 11.7125 29.6825 ;
        RECT  11.8375 29.63 11.8975 29.6875 ;
        RECT  11.6475 29.555 11.7175 31.1 ;
        RECT  11.3125 29.555 11.3825 31.1 ;
        RECT  11.1275 29.555 11.1975 31.1 ;
        RECT  11.8325 29.555 11.9025 31.1 ;
        RECT  11.8325 31.46 11.9025 31.595 ;
        RECT  11.8325 31.46 11.9025 31.595 ;
        RECT  11.8325 31.46 11.9025 31.595 ;
        RECT  11.8325 31.46 11.9025 31.595 ;
        RECT  11.8325 31.46 11.9025 31.595 ;
        RECT  11.8325 31.46 11.9025 31.595 ;
        RECT  11.095 32.31 11.23 32.38 ;
        RECT  11.8 32.31 11.935 32.38 ;
        RECT  11.8325 31.46 11.9025 31.595 ;
        RECT  11.8325 31.46 11.9025 31.595 ;
        RECT  11.8325 31.46 11.9025 31.595 ;
        RECT  11.8325 31.46 11.9025 31.595 ;
        RECT  11.8325 31.46 11.9025 31.595 ;
        RECT  11.8325 31.46 11.9025 31.595 ;
        RECT  11.8325 31.46 11.9025 31.595 ;
        RECT  11.8325 31.46 11.9025 31.595 ;
        RECT  11.3825 31.9525 11.4525 32.0875 ;
        RECT  11.1275 31.46 11.1975 31.595 ;
        RECT  11.1275 31.46 11.1975 31.595 ;
        RECT  11.1275 31.46 11.1975 31.595 ;
        RECT  11.1275 31.46 11.1975 31.595 ;
        RECT  11.1275 31.46 11.1975 31.595 ;
        RECT  11.1275 31.46 11.1975 31.595 ;
        RECT  11.8325 31.46 11.9025 31.595 ;
        RECT  11.8325 31.46 11.9025 31.595 ;
        RECT  11.8325 31.46 11.9025 31.595 ;
        RECT  11.8325 31.46 11.9025 31.595 ;
        RECT  11.5775 31.9525 11.6475 32.0875 ;
        RECT  11.8 32.31 11.935 32.38 ;
        RECT  11.8 32.31 11.935 32.38 ;
        RECT  11.8 32.31 11.935 32.38 ;
        RECT  11.8325 31.46 11.9025 31.595 ;
        RECT  11.8325 31.46 11.9025 31.595 ;
        RECT  11.8325 31.46 11.9025 31.595 ;
        RECT  11.8325 31.46 11.9025 31.595 ;
        RECT  11.8325 31.46 11.9025 31.595 ;
        RECT  11.8325 31.46 11.9025 31.595 ;
        RECT  11.095 32.31 11.23 32.38 ;
        RECT  11.8325 30.9675 11.9025 32.3775 ;
        RECT  11.1325 32.3175 11.1925 32.375 ;
        RECT  11.32 32.3175 11.375 32.37 ;
        RECT  11.655 32.3175 11.7125 32.3775 ;
        RECT  11.8375 32.3125 11.8975 32.37 ;
        RECT  11.6475 30.9 11.7175 32.445 ;
        RECT  11.3125 30.9 11.3825 32.445 ;
        RECT  11.1275 30.9 11.1975 32.445 ;
        RECT  11.8325 30.9 11.9025 32.445 ;
        RECT  11.8325 33.095 11.9025 33.23 ;
        RECT  11.8325 33.095 11.9025 33.23 ;
        RECT  11.8325 33.095 11.9025 33.23 ;
        RECT  11.8325 33.095 11.9025 33.23 ;
        RECT  11.8325 33.095 11.9025 33.23 ;
        RECT  11.8325 33.095 11.9025 33.23 ;
        RECT  11.095 32.31 11.23 32.38 ;
        RECT  11.8 32.31 11.935 32.38 ;
        RECT  11.8325 33.095 11.9025 33.23 ;
        RECT  11.8325 33.095 11.9025 33.23 ;
        RECT  11.8325 33.095 11.9025 33.23 ;
        RECT  11.8325 33.095 11.9025 33.23 ;
        RECT  11.8325 33.095 11.9025 33.23 ;
        RECT  11.8325 33.095 11.9025 33.23 ;
        RECT  11.8325 33.095 11.9025 33.23 ;
        RECT  11.8325 33.095 11.9025 33.23 ;
        RECT  11.3825 32.6025 11.4525 32.7375 ;
        RECT  11.1275 33.095 11.1975 33.23 ;
        RECT  11.1275 33.095 11.1975 33.23 ;
        RECT  11.1275 33.095 11.1975 33.23 ;
        RECT  11.1275 33.095 11.1975 33.23 ;
        RECT  11.1275 33.095 11.1975 33.23 ;
        RECT  11.1275 33.095 11.1975 33.23 ;
        RECT  11.8325 33.095 11.9025 33.23 ;
        RECT  11.8325 33.095 11.9025 33.23 ;
        RECT  11.8325 33.095 11.9025 33.23 ;
        RECT  11.8325 33.095 11.9025 33.23 ;
        RECT  11.5775 32.6025 11.6475 32.7375 ;
        RECT  11.8 32.31 11.935 32.38 ;
        RECT  11.8 32.31 11.935 32.38 ;
        RECT  11.8 32.31 11.935 32.38 ;
        RECT  11.8325 33.095 11.9025 33.23 ;
        RECT  11.8325 33.095 11.9025 33.23 ;
        RECT  11.8325 33.095 11.9025 33.23 ;
        RECT  11.8325 33.095 11.9025 33.23 ;
        RECT  11.8325 33.095 11.9025 33.23 ;
        RECT  11.8325 33.095 11.9025 33.23 ;
        RECT  11.095 32.31 11.23 32.38 ;
        RECT  11.8325 32.3125 11.9025 33.7225 ;
        RECT  11.1325 32.315 11.1925 32.3725 ;
        RECT  11.32 32.32 11.375 32.3725 ;
        RECT  11.655 32.3125 11.7125 32.3725 ;
        RECT  11.8375 32.32 11.8975 32.3775 ;
        RECT  11.6475 32.245 11.7175 33.79 ;
        RECT  11.3125 32.245 11.3825 33.79 ;
        RECT  11.1275 32.245 11.1975 33.79 ;
        RECT  11.8325 32.245 11.9025 33.79 ;
        RECT  11.8325 34.15 11.9025 34.285 ;
        RECT  11.8325 34.15 11.9025 34.285 ;
        RECT  11.8325 34.15 11.9025 34.285 ;
        RECT  11.8325 34.15 11.9025 34.285 ;
        RECT  11.8325 34.15 11.9025 34.285 ;
        RECT  11.8325 34.15 11.9025 34.285 ;
        RECT  11.095 35.0 11.23 35.07 ;
        RECT  11.8 35.0 11.935 35.07 ;
        RECT  11.8325 34.15 11.9025 34.285 ;
        RECT  11.8325 34.15 11.9025 34.285 ;
        RECT  11.8325 34.15 11.9025 34.285 ;
        RECT  11.8325 34.15 11.9025 34.285 ;
        RECT  11.8325 34.15 11.9025 34.285 ;
        RECT  11.8325 34.15 11.9025 34.285 ;
        RECT  11.8325 34.15 11.9025 34.285 ;
        RECT  11.8325 34.15 11.9025 34.285 ;
        RECT  11.3825 34.6425 11.4525 34.7775 ;
        RECT  11.1275 34.15 11.1975 34.285 ;
        RECT  11.1275 34.15 11.1975 34.285 ;
        RECT  11.1275 34.15 11.1975 34.285 ;
        RECT  11.1275 34.15 11.1975 34.285 ;
        RECT  11.1275 34.15 11.1975 34.285 ;
        RECT  11.1275 34.15 11.1975 34.285 ;
        RECT  11.8325 34.15 11.9025 34.285 ;
        RECT  11.8325 34.15 11.9025 34.285 ;
        RECT  11.8325 34.15 11.9025 34.285 ;
        RECT  11.8325 34.15 11.9025 34.285 ;
        RECT  11.5775 34.6425 11.6475 34.7775 ;
        RECT  11.8 35.0 11.935 35.07 ;
        RECT  11.8 35.0 11.935 35.07 ;
        RECT  11.8 35.0 11.935 35.07 ;
        RECT  11.8325 34.15 11.9025 34.285 ;
        RECT  11.8325 34.15 11.9025 34.285 ;
        RECT  11.8325 34.15 11.9025 34.285 ;
        RECT  11.8325 34.15 11.9025 34.285 ;
        RECT  11.8325 34.15 11.9025 34.285 ;
        RECT  11.8325 34.15 11.9025 34.285 ;
        RECT  11.095 35.0 11.23 35.07 ;
        RECT  11.8325 33.6575 11.9025 35.0675 ;
        RECT  11.1325 35.0075 11.1925 35.065 ;
        RECT  11.32 35.0075 11.375 35.06 ;
        RECT  11.655 35.0075 11.7125 35.0675 ;
        RECT  11.8375 35.0025 11.8975 35.06 ;
        RECT  11.6475 33.59 11.7175 35.135 ;
        RECT  11.3125 33.59 11.3825 35.135 ;
        RECT  11.1275 33.59 11.1975 35.135 ;
        RECT  11.8325 33.59 11.9025 35.135 ;
        RECT  11.8325 35.785 11.9025 35.92 ;
        RECT  11.8325 35.785 11.9025 35.92 ;
        RECT  11.8325 35.785 11.9025 35.92 ;
        RECT  11.8325 35.785 11.9025 35.92 ;
        RECT  11.8325 35.785 11.9025 35.92 ;
        RECT  11.8325 35.785 11.9025 35.92 ;
        RECT  11.095 35.0 11.23 35.07 ;
        RECT  11.8 35.0 11.935 35.07 ;
        RECT  11.8325 35.785 11.9025 35.92 ;
        RECT  11.8325 35.785 11.9025 35.92 ;
        RECT  11.8325 35.785 11.9025 35.92 ;
        RECT  11.8325 35.785 11.9025 35.92 ;
        RECT  11.8325 35.785 11.9025 35.92 ;
        RECT  11.8325 35.785 11.9025 35.92 ;
        RECT  11.8325 35.785 11.9025 35.92 ;
        RECT  11.8325 35.785 11.9025 35.92 ;
        RECT  11.3825 35.2925 11.4525 35.4275 ;
        RECT  11.1275 35.785 11.1975 35.92 ;
        RECT  11.1275 35.785 11.1975 35.92 ;
        RECT  11.1275 35.785 11.1975 35.92 ;
        RECT  11.1275 35.785 11.1975 35.92 ;
        RECT  11.1275 35.785 11.1975 35.92 ;
        RECT  11.1275 35.785 11.1975 35.92 ;
        RECT  11.8325 35.785 11.9025 35.92 ;
        RECT  11.8325 35.785 11.9025 35.92 ;
        RECT  11.8325 35.785 11.9025 35.92 ;
        RECT  11.8325 35.785 11.9025 35.92 ;
        RECT  11.5775 35.2925 11.6475 35.4275 ;
        RECT  11.8 35.0 11.935 35.07 ;
        RECT  11.8 35.0 11.935 35.07 ;
        RECT  11.8 35.0 11.935 35.07 ;
        RECT  11.8325 35.785 11.9025 35.92 ;
        RECT  11.8325 35.785 11.9025 35.92 ;
        RECT  11.8325 35.785 11.9025 35.92 ;
        RECT  11.8325 35.785 11.9025 35.92 ;
        RECT  11.8325 35.785 11.9025 35.92 ;
        RECT  11.8325 35.785 11.9025 35.92 ;
        RECT  11.095 35.0 11.23 35.07 ;
        RECT  11.8325 35.0025 11.9025 36.4125 ;
        RECT  11.1325 35.005 11.1925 35.0625 ;
        RECT  11.32 35.01 11.375 35.0625 ;
        RECT  11.655 35.0025 11.7125 35.0625 ;
        RECT  11.8375 35.01 11.8975 35.0675 ;
        RECT  11.6475 34.935 11.7175 36.48 ;
        RECT  11.3125 34.935 11.3825 36.48 ;
        RECT  11.1275 34.935 11.1975 36.48 ;
        RECT  11.8325 34.935 11.9025 36.48 ;
        RECT  11.8325 36.84 11.9025 36.975 ;
        RECT  11.8325 36.84 11.9025 36.975 ;
        RECT  11.8325 36.84 11.9025 36.975 ;
        RECT  11.8325 36.84 11.9025 36.975 ;
        RECT  11.8325 36.84 11.9025 36.975 ;
        RECT  11.8325 36.84 11.9025 36.975 ;
        RECT  11.095 37.69 11.23 37.76 ;
        RECT  11.8 37.69 11.935 37.76 ;
        RECT  11.8325 36.84 11.9025 36.975 ;
        RECT  11.8325 36.84 11.9025 36.975 ;
        RECT  11.8325 36.84 11.9025 36.975 ;
        RECT  11.8325 36.84 11.9025 36.975 ;
        RECT  11.8325 36.84 11.9025 36.975 ;
        RECT  11.8325 36.84 11.9025 36.975 ;
        RECT  11.8325 36.84 11.9025 36.975 ;
        RECT  11.8325 36.84 11.9025 36.975 ;
        RECT  11.3825 37.3325 11.4525 37.4675 ;
        RECT  11.1275 36.84 11.1975 36.975 ;
        RECT  11.1275 36.84 11.1975 36.975 ;
        RECT  11.1275 36.84 11.1975 36.975 ;
        RECT  11.1275 36.84 11.1975 36.975 ;
        RECT  11.1275 36.84 11.1975 36.975 ;
        RECT  11.1275 36.84 11.1975 36.975 ;
        RECT  11.8325 36.84 11.9025 36.975 ;
        RECT  11.8325 36.84 11.9025 36.975 ;
        RECT  11.8325 36.84 11.9025 36.975 ;
        RECT  11.8325 36.84 11.9025 36.975 ;
        RECT  11.5775 37.3325 11.6475 37.4675 ;
        RECT  11.8 37.69 11.935 37.76 ;
        RECT  11.8 37.69 11.935 37.76 ;
        RECT  11.8 37.69 11.935 37.76 ;
        RECT  11.8325 36.84 11.9025 36.975 ;
        RECT  11.8325 36.84 11.9025 36.975 ;
        RECT  11.8325 36.84 11.9025 36.975 ;
        RECT  11.8325 36.84 11.9025 36.975 ;
        RECT  11.8325 36.84 11.9025 36.975 ;
        RECT  11.8325 36.84 11.9025 36.975 ;
        RECT  11.095 37.69 11.23 37.76 ;
        RECT  11.8325 36.3475 11.9025 37.7575 ;
        RECT  11.1325 37.6975 11.1925 37.755 ;
        RECT  11.32 37.6975 11.375 37.75 ;
        RECT  11.655 37.6975 11.7125 37.7575 ;
        RECT  11.8375 37.6925 11.8975 37.75 ;
        RECT  11.6475 36.28 11.7175 37.825 ;
        RECT  11.3125 36.28 11.3825 37.825 ;
        RECT  11.1275 36.28 11.1975 37.825 ;
        RECT  11.8325 36.28 11.9025 37.825 ;
        RECT  11.8325 38.475 11.9025 38.61 ;
        RECT  11.8325 38.475 11.9025 38.61 ;
        RECT  11.8325 38.475 11.9025 38.61 ;
        RECT  11.8325 38.475 11.9025 38.61 ;
        RECT  11.8325 38.475 11.9025 38.61 ;
        RECT  11.8325 38.475 11.9025 38.61 ;
        RECT  11.095 37.69 11.23 37.76 ;
        RECT  11.8 37.69 11.935 37.76 ;
        RECT  11.8325 38.475 11.9025 38.61 ;
        RECT  11.8325 38.475 11.9025 38.61 ;
        RECT  11.8325 38.475 11.9025 38.61 ;
        RECT  11.8325 38.475 11.9025 38.61 ;
        RECT  11.8325 38.475 11.9025 38.61 ;
        RECT  11.8325 38.475 11.9025 38.61 ;
        RECT  11.8325 38.475 11.9025 38.61 ;
        RECT  11.8325 38.475 11.9025 38.61 ;
        RECT  11.3825 37.9825 11.4525 38.1175 ;
        RECT  11.1275 38.475 11.1975 38.61 ;
        RECT  11.1275 38.475 11.1975 38.61 ;
        RECT  11.1275 38.475 11.1975 38.61 ;
        RECT  11.1275 38.475 11.1975 38.61 ;
        RECT  11.1275 38.475 11.1975 38.61 ;
        RECT  11.1275 38.475 11.1975 38.61 ;
        RECT  11.8325 38.475 11.9025 38.61 ;
        RECT  11.8325 38.475 11.9025 38.61 ;
        RECT  11.8325 38.475 11.9025 38.61 ;
        RECT  11.8325 38.475 11.9025 38.61 ;
        RECT  11.5775 37.9825 11.6475 38.1175 ;
        RECT  11.8 37.69 11.935 37.76 ;
        RECT  11.8 37.69 11.935 37.76 ;
        RECT  11.8 37.69 11.935 37.76 ;
        RECT  11.8325 38.475 11.9025 38.61 ;
        RECT  11.8325 38.475 11.9025 38.61 ;
        RECT  11.8325 38.475 11.9025 38.61 ;
        RECT  11.8325 38.475 11.9025 38.61 ;
        RECT  11.8325 38.475 11.9025 38.61 ;
        RECT  11.8325 38.475 11.9025 38.61 ;
        RECT  11.095 37.69 11.23 37.76 ;
        RECT  11.8325 37.6925 11.9025 39.1025 ;
        RECT  11.1325 37.695 11.1925 37.7525 ;
        RECT  11.32 37.7 11.375 37.7525 ;
        RECT  11.655 37.6925 11.7125 37.7525 ;
        RECT  11.8375 37.7 11.8975 37.7575 ;
        RECT  11.6475 37.625 11.7175 39.17 ;
        RECT  11.3125 37.625 11.3825 39.17 ;
        RECT  11.1275 37.625 11.1975 39.17 ;
        RECT  11.8325 37.625 11.9025 39.17 ;
        RECT  11.8325 39.53 11.9025 39.665 ;
        RECT  11.8325 39.53 11.9025 39.665 ;
        RECT  11.8325 39.53 11.9025 39.665 ;
        RECT  11.8325 39.53 11.9025 39.665 ;
        RECT  11.8325 39.53 11.9025 39.665 ;
        RECT  11.8325 39.53 11.9025 39.665 ;
        RECT  11.095 40.38 11.23 40.45 ;
        RECT  11.8 40.38 11.935 40.45 ;
        RECT  11.8325 39.53 11.9025 39.665 ;
        RECT  11.8325 39.53 11.9025 39.665 ;
        RECT  11.8325 39.53 11.9025 39.665 ;
        RECT  11.8325 39.53 11.9025 39.665 ;
        RECT  11.8325 39.53 11.9025 39.665 ;
        RECT  11.8325 39.53 11.9025 39.665 ;
        RECT  11.8325 39.53 11.9025 39.665 ;
        RECT  11.8325 39.53 11.9025 39.665 ;
        RECT  11.3825 40.0225 11.4525 40.1575 ;
        RECT  11.1275 39.53 11.1975 39.665 ;
        RECT  11.1275 39.53 11.1975 39.665 ;
        RECT  11.1275 39.53 11.1975 39.665 ;
        RECT  11.1275 39.53 11.1975 39.665 ;
        RECT  11.1275 39.53 11.1975 39.665 ;
        RECT  11.1275 39.53 11.1975 39.665 ;
        RECT  11.8325 39.53 11.9025 39.665 ;
        RECT  11.8325 39.53 11.9025 39.665 ;
        RECT  11.8325 39.53 11.9025 39.665 ;
        RECT  11.8325 39.53 11.9025 39.665 ;
        RECT  11.5775 40.0225 11.6475 40.1575 ;
        RECT  11.8 40.38 11.935 40.45 ;
        RECT  11.8 40.38 11.935 40.45 ;
        RECT  11.8 40.38 11.935 40.45 ;
        RECT  11.8325 39.53 11.9025 39.665 ;
        RECT  11.8325 39.53 11.9025 39.665 ;
        RECT  11.8325 39.53 11.9025 39.665 ;
        RECT  11.8325 39.53 11.9025 39.665 ;
        RECT  11.8325 39.53 11.9025 39.665 ;
        RECT  11.8325 39.53 11.9025 39.665 ;
        RECT  11.095 40.38 11.23 40.45 ;
        RECT  11.8325 39.0375 11.9025 40.4475 ;
        RECT  11.1325 40.3875 11.1925 40.445 ;
        RECT  11.32 40.3875 11.375 40.44 ;
        RECT  11.655 40.3875 11.7125 40.4475 ;
        RECT  11.8375 40.3825 11.8975 40.44 ;
        RECT  11.6475 38.97 11.7175 40.515 ;
        RECT  11.3125 38.97 11.3825 40.515 ;
        RECT  11.1275 38.97 11.1975 40.515 ;
        RECT  11.8325 38.97 11.9025 40.515 ;
        RECT  12.5375 19.645 12.6075 19.78 ;
        RECT  12.5375 19.645 12.6075 19.78 ;
        RECT  12.5375 19.645 12.6075 19.78 ;
        RECT  12.5375 19.645 12.6075 19.78 ;
        RECT  12.5375 19.645 12.6075 19.78 ;
        RECT  12.5375 19.645 12.6075 19.78 ;
        RECT  11.8 18.86 11.935 18.93 ;
        RECT  12.505 18.86 12.64 18.93 ;
        RECT  12.5375 19.645 12.6075 19.78 ;
        RECT  12.5375 19.645 12.6075 19.78 ;
        RECT  12.5375 19.645 12.6075 19.78 ;
        RECT  12.5375 19.645 12.6075 19.78 ;
        RECT  12.5375 19.645 12.6075 19.78 ;
        RECT  12.5375 19.645 12.6075 19.78 ;
        RECT  12.5375 19.645 12.6075 19.78 ;
        RECT  12.5375 19.645 12.6075 19.78 ;
        RECT  12.0875 19.1525 12.1575 19.2875 ;
        RECT  11.8325 19.645 11.9025 19.78 ;
        RECT  11.8325 19.645 11.9025 19.78 ;
        RECT  11.8325 19.645 11.9025 19.78 ;
        RECT  11.8325 19.645 11.9025 19.78 ;
        RECT  11.8325 19.645 11.9025 19.78 ;
        RECT  11.8325 19.645 11.9025 19.78 ;
        RECT  12.5375 19.645 12.6075 19.78 ;
        RECT  12.5375 19.645 12.6075 19.78 ;
        RECT  12.5375 19.645 12.6075 19.78 ;
        RECT  12.5375 19.645 12.6075 19.78 ;
        RECT  12.2825 19.1525 12.3525 19.2875 ;
        RECT  12.505 18.86 12.64 18.93 ;
        RECT  12.505 18.86 12.64 18.93 ;
        RECT  12.505 18.86 12.64 18.93 ;
        RECT  12.5375 19.645 12.6075 19.78 ;
        RECT  12.5375 19.645 12.6075 19.78 ;
        RECT  12.5375 19.645 12.6075 19.78 ;
        RECT  12.5375 19.645 12.6075 19.78 ;
        RECT  12.5375 19.645 12.6075 19.78 ;
        RECT  12.5375 19.645 12.6075 19.78 ;
        RECT  11.8 18.86 11.935 18.93 ;
        RECT  12.5375 18.8625 12.6075 20.2725 ;
        RECT  11.8375 18.865 11.8975 18.9225 ;
        RECT  12.025 18.87 12.08 18.9225 ;
        RECT  12.36 18.8625 12.4175 18.9225 ;
        RECT  12.5425 18.87 12.6025 18.9275 ;
        RECT  12.3525 18.795 12.4225 20.34 ;
        RECT  12.0175 18.795 12.0875 20.34 ;
        RECT  11.8325 18.795 11.9025 20.34 ;
        RECT  12.5375 18.795 12.6075 20.34 ;
        RECT  12.5375 20.7 12.6075 20.835 ;
        RECT  12.5375 20.7 12.6075 20.835 ;
        RECT  12.5375 20.7 12.6075 20.835 ;
        RECT  12.5375 20.7 12.6075 20.835 ;
        RECT  12.5375 20.7 12.6075 20.835 ;
        RECT  12.5375 20.7 12.6075 20.835 ;
        RECT  11.8 21.55 11.935 21.62 ;
        RECT  12.505 21.55 12.64 21.62 ;
        RECT  12.5375 20.7 12.6075 20.835 ;
        RECT  12.5375 20.7 12.6075 20.835 ;
        RECT  12.5375 20.7 12.6075 20.835 ;
        RECT  12.5375 20.7 12.6075 20.835 ;
        RECT  12.5375 20.7 12.6075 20.835 ;
        RECT  12.5375 20.7 12.6075 20.835 ;
        RECT  12.5375 20.7 12.6075 20.835 ;
        RECT  12.5375 20.7 12.6075 20.835 ;
        RECT  12.0875 21.1925 12.1575 21.3275 ;
        RECT  11.8325 20.7 11.9025 20.835 ;
        RECT  11.8325 20.7 11.9025 20.835 ;
        RECT  11.8325 20.7 11.9025 20.835 ;
        RECT  11.8325 20.7 11.9025 20.835 ;
        RECT  11.8325 20.7 11.9025 20.835 ;
        RECT  11.8325 20.7 11.9025 20.835 ;
        RECT  12.5375 20.7 12.6075 20.835 ;
        RECT  12.5375 20.7 12.6075 20.835 ;
        RECT  12.5375 20.7 12.6075 20.835 ;
        RECT  12.5375 20.7 12.6075 20.835 ;
        RECT  12.2825 21.1925 12.3525 21.3275 ;
        RECT  12.505 21.55 12.64 21.62 ;
        RECT  12.505 21.55 12.64 21.62 ;
        RECT  12.505 21.55 12.64 21.62 ;
        RECT  12.5375 20.7 12.6075 20.835 ;
        RECT  12.5375 20.7 12.6075 20.835 ;
        RECT  12.5375 20.7 12.6075 20.835 ;
        RECT  12.5375 20.7 12.6075 20.835 ;
        RECT  12.5375 20.7 12.6075 20.835 ;
        RECT  12.5375 20.7 12.6075 20.835 ;
        RECT  11.8 21.55 11.935 21.62 ;
        RECT  12.5375 20.2075 12.6075 21.6175 ;
        RECT  11.8375 21.5575 11.8975 21.615 ;
        RECT  12.025 21.5575 12.08 21.61 ;
        RECT  12.36 21.5575 12.4175 21.6175 ;
        RECT  12.5425 21.5525 12.6025 21.61 ;
        RECT  12.3525 20.14 12.4225 21.685 ;
        RECT  12.0175 20.14 12.0875 21.685 ;
        RECT  11.8325 20.14 11.9025 21.685 ;
        RECT  12.5375 20.14 12.6075 21.685 ;
        RECT  12.5375 22.335 12.6075 22.47 ;
        RECT  12.5375 22.335 12.6075 22.47 ;
        RECT  12.5375 22.335 12.6075 22.47 ;
        RECT  12.5375 22.335 12.6075 22.47 ;
        RECT  12.5375 22.335 12.6075 22.47 ;
        RECT  12.5375 22.335 12.6075 22.47 ;
        RECT  11.8 21.55 11.935 21.62 ;
        RECT  12.505 21.55 12.64 21.62 ;
        RECT  12.5375 22.335 12.6075 22.47 ;
        RECT  12.5375 22.335 12.6075 22.47 ;
        RECT  12.5375 22.335 12.6075 22.47 ;
        RECT  12.5375 22.335 12.6075 22.47 ;
        RECT  12.5375 22.335 12.6075 22.47 ;
        RECT  12.5375 22.335 12.6075 22.47 ;
        RECT  12.5375 22.335 12.6075 22.47 ;
        RECT  12.5375 22.335 12.6075 22.47 ;
        RECT  12.0875 21.8425 12.1575 21.9775 ;
        RECT  11.8325 22.335 11.9025 22.47 ;
        RECT  11.8325 22.335 11.9025 22.47 ;
        RECT  11.8325 22.335 11.9025 22.47 ;
        RECT  11.8325 22.335 11.9025 22.47 ;
        RECT  11.8325 22.335 11.9025 22.47 ;
        RECT  11.8325 22.335 11.9025 22.47 ;
        RECT  12.5375 22.335 12.6075 22.47 ;
        RECT  12.5375 22.335 12.6075 22.47 ;
        RECT  12.5375 22.335 12.6075 22.47 ;
        RECT  12.5375 22.335 12.6075 22.47 ;
        RECT  12.2825 21.8425 12.3525 21.9775 ;
        RECT  12.505 21.55 12.64 21.62 ;
        RECT  12.505 21.55 12.64 21.62 ;
        RECT  12.505 21.55 12.64 21.62 ;
        RECT  12.5375 22.335 12.6075 22.47 ;
        RECT  12.5375 22.335 12.6075 22.47 ;
        RECT  12.5375 22.335 12.6075 22.47 ;
        RECT  12.5375 22.335 12.6075 22.47 ;
        RECT  12.5375 22.335 12.6075 22.47 ;
        RECT  12.5375 22.335 12.6075 22.47 ;
        RECT  11.8 21.55 11.935 21.62 ;
        RECT  12.5375 21.5525 12.6075 22.9625 ;
        RECT  11.8375 21.555 11.8975 21.6125 ;
        RECT  12.025 21.56 12.08 21.6125 ;
        RECT  12.36 21.5525 12.4175 21.6125 ;
        RECT  12.5425 21.56 12.6025 21.6175 ;
        RECT  12.3525 21.485 12.4225 23.03 ;
        RECT  12.0175 21.485 12.0875 23.03 ;
        RECT  11.8325 21.485 11.9025 23.03 ;
        RECT  12.5375 21.485 12.6075 23.03 ;
        RECT  12.5375 23.39 12.6075 23.525 ;
        RECT  12.5375 23.39 12.6075 23.525 ;
        RECT  12.5375 23.39 12.6075 23.525 ;
        RECT  12.5375 23.39 12.6075 23.525 ;
        RECT  12.5375 23.39 12.6075 23.525 ;
        RECT  12.5375 23.39 12.6075 23.525 ;
        RECT  11.8 24.24 11.935 24.31 ;
        RECT  12.505 24.24 12.64 24.31 ;
        RECT  12.5375 23.39 12.6075 23.525 ;
        RECT  12.5375 23.39 12.6075 23.525 ;
        RECT  12.5375 23.39 12.6075 23.525 ;
        RECT  12.5375 23.39 12.6075 23.525 ;
        RECT  12.5375 23.39 12.6075 23.525 ;
        RECT  12.5375 23.39 12.6075 23.525 ;
        RECT  12.5375 23.39 12.6075 23.525 ;
        RECT  12.5375 23.39 12.6075 23.525 ;
        RECT  12.0875 23.8825 12.1575 24.0175 ;
        RECT  11.8325 23.39 11.9025 23.525 ;
        RECT  11.8325 23.39 11.9025 23.525 ;
        RECT  11.8325 23.39 11.9025 23.525 ;
        RECT  11.8325 23.39 11.9025 23.525 ;
        RECT  11.8325 23.39 11.9025 23.525 ;
        RECT  11.8325 23.39 11.9025 23.525 ;
        RECT  12.5375 23.39 12.6075 23.525 ;
        RECT  12.5375 23.39 12.6075 23.525 ;
        RECT  12.5375 23.39 12.6075 23.525 ;
        RECT  12.5375 23.39 12.6075 23.525 ;
        RECT  12.2825 23.8825 12.3525 24.0175 ;
        RECT  12.505 24.24 12.64 24.31 ;
        RECT  12.505 24.24 12.64 24.31 ;
        RECT  12.505 24.24 12.64 24.31 ;
        RECT  12.5375 23.39 12.6075 23.525 ;
        RECT  12.5375 23.39 12.6075 23.525 ;
        RECT  12.5375 23.39 12.6075 23.525 ;
        RECT  12.5375 23.39 12.6075 23.525 ;
        RECT  12.5375 23.39 12.6075 23.525 ;
        RECT  12.5375 23.39 12.6075 23.525 ;
        RECT  11.8 24.24 11.935 24.31 ;
        RECT  12.5375 22.8975 12.6075 24.3075 ;
        RECT  11.8375 24.2475 11.8975 24.305 ;
        RECT  12.025 24.2475 12.08 24.3 ;
        RECT  12.36 24.2475 12.4175 24.3075 ;
        RECT  12.5425 24.2425 12.6025 24.3 ;
        RECT  12.3525 22.83 12.4225 24.375 ;
        RECT  12.0175 22.83 12.0875 24.375 ;
        RECT  11.8325 22.83 11.9025 24.375 ;
        RECT  12.5375 22.83 12.6075 24.375 ;
        RECT  12.5375 25.025 12.6075 25.16 ;
        RECT  12.5375 25.025 12.6075 25.16 ;
        RECT  12.5375 25.025 12.6075 25.16 ;
        RECT  12.5375 25.025 12.6075 25.16 ;
        RECT  12.5375 25.025 12.6075 25.16 ;
        RECT  12.5375 25.025 12.6075 25.16 ;
        RECT  11.8 24.24 11.935 24.31 ;
        RECT  12.505 24.24 12.64 24.31 ;
        RECT  12.5375 25.025 12.6075 25.16 ;
        RECT  12.5375 25.025 12.6075 25.16 ;
        RECT  12.5375 25.025 12.6075 25.16 ;
        RECT  12.5375 25.025 12.6075 25.16 ;
        RECT  12.5375 25.025 12.6075 25.16 ;
        RECT  12.5375 25.025 12.6075 25.16 ;
        RECT  12.5375 25.025 12.6075 25.16 ;
        RECT  12.5375 25.025 12.6075 25.16 ;
        RECT  12.0875 24.5325 12.1575 24.6675 ;
        RECT  11.8325 25.025 11.9025 25.16 ;
        RECT  11.8325 25.025 11.9025 25.16 ;
        RECT  11.8325 25.025 11.9025 25.16 ;
        RECT  11.8325 25.025 11.9025 25.16 ;
        RECT  11.8325 25.025 11.9025 25.16 ;
        RECT  11.8325 25.025 11.9025 25.16 ;
        RECT  12.5375 25.025 12.6075 25.16 ;
        RECT  12.5375 25.025 12.6075 25.16 ;
        RECT  12.5375 25.025 12.6075 25.16 ;
        RECT  12.5375 25.025 12.6075 25.16 ;
        RECT  12.2825 24.5325 12.3525 24.6675 ;
        RECT  12.505 24.24 12.64 24.31 ;
        RECT  12.505 24.24 12.64 24.31 ;
        RECT  12.505 24.24 12.64 24.31 ;
        RECT  12.5375 25.025 12.6075 25.16 ;
        RECT  12.5375 25.025 12.6075 25.16 ;
        RECT  12.5375 25.025 12.6075 25.16 ;
        RECT  12.5375 25.025 12.6075 25.16 ;
        RECT  12.5375 25.025 12.6075 25.16 ;
        RECT  12.5375 25.025 12.6075 25.16 ;
        RECT  11.8 24.24 11.935 24.31 ;
        RECT  12.5375 24.2425 12.6075 25.6525 ;
        RECT  11.8375 24.245 11.8975 24.3025 ;
        RECT  12.025 24.25 12.08 24.3025 ;
        RECT  12.36 24.2425 12.4175 24.3025 ;
        RECT  12.5425 24.25 12.6025 24.3075 ;
        RECT  12.3525 24.175 12.4225 25.72 ;
        RECT  12.0175 24.175 12.0875 25.72 ;
        RECT  11.8325 24.175 11.9025 25.72 ;
        RECT  12.5375 24.175 12.6075 25.72 ;
        RECT  12.5375 26.08 12.6075 26.215 ;
        RECT  12.5375 26.08 12.6075 26.215 ;
        RECT  12.5375 26.08 12.6075 26.215 ;
        RECT  12.5375 26.08 12.6075 26.215 ;
        RECT  12.5375 26.08 12.6075 26.215 ;
        RECT  12.5375 26.08 12.6075 26.215 ;
        RECT  11.8 26.93 11.935 27.0 ;
        RECT  12.505 26.93 12.64 27.0 ;
        RECT  12.5375 26.08 12.6075 26.215 ;
        RECT  12.5375 26.08 12.6075 26.215 ;
        RECT  12.5375 26.08 12.6075 26.215 ;
        RECT  12.5375 26.08 12.6075 26.215 ;
        RECT  12.5375 26.08 12.6075 26.215 ;
        RECT  12.5375 26.08 12.6075 26.215 ;
        RECT  12.5375 26.08 12.6075 26.215 ;
        RECT  12.5375 26.08 12.6075 26.215 ;
        RECT  12.0875 26.5725 12.1575 26.7075 ;
        RECT  11.8325 26.08 11.9025 26.215 ;
        RECT  11.8325 26.08 11.9025 26.215 ;
        RECT  11.8325 26.08 11.9025 26.215 ;
        RECT  11.8325 26.08 11.9025 26.215 ;
        RECT  11.8325 26.08 11.9025 26.215 ;
        RECT  11.8325 26.08 11.9025 26.215 ;
        RECT  12.5375 26.08 12.6075 26.215 ;
        RECT  12.5375 26.08 12.6075 26.215 ;
        RECT  12.5375 26.08 12.6075 26.215 ;
        RECT  12.5375 26.08 12.6075 26.215 ;
        RECT  12.2825 26.5725 12.3525 26.7075 ;
        RECT  12.505 26.93 12.64 27.0 ;
        RECT  12.505 26.93 12.64 27.0 ;
        RECT  12.505 26.93 12.64 27.0 ;
        RECT  12.5375 26.08 12.6075 26.215 ;
        RECT  12.5375 26.08 12.6075 26.215 ;
        RECT  12.5375 26.08 12.6075 26.215 ;
        RECT  12.5375 26.08 12.6075 26.215 ;
        RECT  12.5375 26.08 12.6075 26.215 ;
        RECT  12.5375 26.08 12.6075 26.215 ;
        RECT  11.8 26.93 11.935 27.0 ;
        RECT  12.5375 25.5875 12.6075 26.9975 ;
        RECT  11.8375 26.9375 11.8975 26.995 ;
        RECT  12.025 26.9375 12.08 26.99 ;
        RECT  12.36 26.9375 12.4175 26.9975 ;
        RECT  12.5425 26.9325 12.6025 26.99 ;
        RECT  12.3525 25.52 12.4225 27.065 ;
        RECT  12.0175 25.52 12.0875 27.065 ;
        RECT  11.8325 25.52 11.9025 27.065 ;
        RECT  12.5375 25.52 12.6075 27.065 ;
        RECT  12.5375 27.715 12.6075 27.85 ;
        RECT  12.5375 27.715 12.6075 27.85 ;
        RECT  12.5375 27.715 12.6075 27.85 ;
        RECT  12.5375 27.715 12.6075 27.85 ;
        RECT  12.5375 27.715 12.6075 27.85 ;
        RECT  12.5375 27.715 12.6075 27.85 ;
        RECT  11.8 26.93 11.935 27.0 ;
        RECT  12.505 26.93 12.64 27.0 ;
        RECT  12.5375 27.715 12.6075 27.85 ;
        RECT  12.5375 27.715 12.6075 27.85 ;
        RECT  12.5375 27.715 12.6075 27.85 ;
        RECT  12.5375 27.715 12.6075 27.85 ;
        RECT  12.5375 27.715 12.6075 27.85 ;
        RECT  12.5375 27.715 12.6075 27.85 ;
        RECT  12.5375 27.715 12.6075 27.85 ;
        RECT  12.5375 27.715 12.6075 27.85 ;
        RECT  12.0875 27.2225 12.1575 27.3575 ;
        RECT  11.8325 27.715 11.9025 27.85 ;
        RECT  11.8325 27.715 11.9025 27.85 ;
        RECT  11.8325 27.715 11.9025 27.85 ;
        RECT  11.8325 27.715 11.9025 27.85 ;
        RECT  11.8325 27.715 11.9025 27.85 ;
        RECT  11.8325 27.715 11.9025 27.85 ;
        RECT  12.5375 27.715 12.6075 27.85 ;
        RECT  12.5375 27.715 12.6075 27.85 ;
        RECT  12.5375 27.715 12.6075 27.85 ;
        RECT  12.5375 27.715 12.6075 27.85 ;
        RECT  12.2825 27.2225 12.3525 27.3575 ;
        RECT  12.505 26.93 12.64 27.0 ;
        RECT  12.505 26.93 12.64 27.0 ;
        RECT  12.505 26.93 12.64 27.0 ;
        RECT  12.5375 27.715 12.6075 27.85 ;
        RECT  12.5375 27.715 12.6075 27.85 ;
        RECT  12.5375 27.715 12.6075 27.85 ;
        RECT  12.5375 27.715 12.6075 27.85 ;
        RECT  12.5375 27.715 12.6075 27.85 ;
        RECT  12.5375 27.715 12.6075 27.85 ;
        RECT  11.8 26.93 11.935 27.0 ;
        RECT  12.5375 26.9325 12.6075 28.3425 ;
        RECT  11.8375 26.935 11.8975 26.9925 ;
        RECT  12.025 26.94 12.08 26.9925 ;
        RECT  12.36 26.9325 12.4175 26.9925 ;
        RECT  12.5425 26.94 12.6025 26.9975 ;
        RECT  12.3525 26.865 12.4225 28.41 ;
        RECT  12.0175 26.865 12.0875 28.41 ;
        RECT  11.8325 26.865 11.9025 28.41 ;
        RECT  12.5375 26.865 12.6075 28.41 ;
        RECT  12.5375 28.77 12.6075 28.905 ;
        RECT  12.5375 28.77 12.6075 28.905 ;
        RECT  12.5375 28.77 12.6075 28.905 ;
        RECT  12.5375 28.77 12.6075 28.905 ;
        RECT  12.5375 28.77 12.6075 28.905 ;
        RECT  12.5375 28.77 12.6075 28.905 ;
        RECT  11.8 29.62 11.935 29.69 ;
        RECT  12.505 29.62 12.64 29.69 ;
        RECT  12.5375 28.77 12.6075 28.905 ;
        RECT  12.5375 28.77 12.6075 28.905 ;
        RECT  12.5375 28.77 12.6075 28.905 ;
        RECT  12.5375 28.77 12.6075 28.905 ;
        RECT  12.5375 28.77 12.6075 28.905 ;
        RECT  12.5375 28.77 12.6075 28.905 ;
        RECT  12.5375 28.77 12.6075 28.905 ;
        RECT  12.5375 28.77 12.6075 28.905 ;
        RECT  12.0875 29.2625 12.1575 29.3975 ;
        RECT  11.8325 28.77 11.9025 28.905 ;
        RECT  11.8325 28.77 11.9025 28.905 ;
        RECT  11.8325 28.77 11.9025 28.905 ;
        RECT  11.8325 28.77 11.9025 28.905 ;
        RECT  11.8325 28.77 11.9025 28.905 ;
        RECT  11.8325 28.77 11.9025 28.905 ;
        RECT  12.5375 28.77 12.6075 28.905 ;
        RECT  12.5375 28.77 12.6075 28.905 ;
        RECT  12.5375 28.77 12.6075 28.905 ;
        RECT  12.5375 28.77 12.6075 28.905 ;
        RECT  12.2825 29.2625 12.3525 29.3975 ;
        RECT  12.505 29.62 12.64 29.69 ;
        RECT  12.505 29.62 12.64 29.69 ;
        RECT  12.505 29.62 12.64 29.69 ;
        RECT  12.5375 28.77 12.6075 28.905 ;
        RECT  12.5375 28.77 12.6075 28.905 ;
        RECT  12.5375 28.77 12.6075 28.905 ;
        RECT  12.5375 28.77 12.6075 28.905 ;
        RECT  12.5375 28.77 12.6075 28.905 ;
        RECT  12.5375 28.77 12.6075 28.905 ;
        RECT  11.8 29.62 11.935 29.69 ;
        RECT  12.5375 28.2775 12.6075 29.6875 ;
        RECT  11.8375 29.6275 11.8975 29.685 ;
        RECT  12.025 29.6275 12.08 29.68 ;
        RECT  12.36 29.6275 12.4175 29.6875 ;
        RECT  12.5425 29.6225 12.6025 29.68 ;
        RECT  12.3525 28.21 12.4225 29.755 ;
        RECT  12.0175 28.21 12.0875 29.755 ;
        RECT  11.8325 28.21 11.9025 29.755 ;
        RECT  12.5375 28.21 12.6075 29.755 ;
        RECT  12.5375 30.405 12.6075 30.54 ;
        RECT  12.5375 30.405 12.6075 30.54 ;
        RECT  12.5375 30.405 12.6075 30.54 ;
        RECT  12.5375 30.405 12.6075 30.54 ;
        RECT  12.5375 30.405 12.6075 30.54 ;
        RECT  12.5375 30.405 12.6075 30.54 ;
        RECT  11.8 29.62 11.935 29.69 ;
        RECT  12.505 29.62 12.64 29.69 ;
        RECT  12.5375 30.405 12.6075 30.54 ;
        RECT  12.5375 30.405 12.6075 30.54 ;
        RECT  12.5375 30.405 12.6075 30.54 ;
        RECT  12.5375 30.405 12.6075 30.54 ;
        RECT  12.5375 30.405 12.6075 30.54 ;
        RECT  12.5375 30.405 12.6075 30.54 ;
        RECT  12.5375 30.405 12.6075 30.54 ;
        RECT  12.5375 30.405 12.6075 30.54 ;
        RECT  12.0875 29.9125 12.1575 30.0475 ;
        RECT  11.8325 30.405 11.9025 30.54 ;
        RECT  11.8325 30.405 11.9025 30.54 ;
        RECT  11.8325 30.405 11.9025 30.54 ;
        RECT  11.8325 30.405 11.9025 30.54 ;
        RECT  11.8325 30.405 11.9025 30.54 ;
        RECT  11.8325 30.405 11.9025 30.54 ;
        RECT  12.5375 30.405 12.6075 30.54 ;
        RECT  12.5375 30.405 12.6075 30.54 ;
        RECT  12.5375 30.405 12.6075 30.54 ;
        RECT  12.5375 30.405 12.6075 30.54 ;
        RECT  12.2825 29.9125 12.3525 30.0475 ;
        RECT  12.505 29.62 12.64 29.69 ;
        RECT  12.505 29.62 12.64 29.69 ;
        RECT  12.505 29.62 12.64 29.69 ;
        RECT  12.5375 30.405 12.6075 30.54 ;
        RECT  12.5375 30.405 12.6075 30.54 ;
        RECT  12.5375 30.405 12.6075 30.54 ;
        RECT  12.5375 30.405 12.6075 30.54 ;
        RECT  12.5375 30.405 12.6075 30.54 ;
        RECT  12.5375 30.405 12.6075 30.54 ;
        RECT  11.8 29.62 11.935 29.69 ;
        RECT  12.5375 29.6225 12.6075 31.0325 ;
        RECT  11.8375 29.625 11.8975 29.6825 ;
        RECT  12.025 29.63 12.08 29.6825 ;
        RECT  12.36 29.6225 12.4175 29.6825 ;
        RECT  12.5425 29.63 12.6025 29.6875 ;
        RECT  12.3525 29.555 12.4225 31.1 ;
        RECT  12.0175 29.555 12.0875 31.1 ;
        RECT  11.8325 29.555 11.9025 31.1 ;
        RECT  12.5375 29.555 12.6075 31.1 ;
        RECT  12.5375 31.46 12.6075 31.595 ;
        RECT  12.5375 31.46 12.6075 31.595 ;
        RECT  12.5375 31.46 12.6075 31.595 ;
        RECT  12.5375 31.46 12.6075 31.595 ;
        RECT  12.5375 31.46 12.6075 31.595 ;
        RECT  12.5375 31.46 12.6075 31.595 ;
        RECT  11.8 32.31 11.935 32.38 ;
        RECT  12.505 32.31 12.64 32.38 ;
        RECT  12.5375 31.46 12.6075 31.595 ;
        RECT  12.5375 31.46 12.6075 31.595 ;
        RECT  12.5375 31.46 12.6075 31.595 ;
        RECT  12.5375 31.46 12.6075 31.595 ;
        RECT  12.5375 31.46 12.6075 31.595 ;
        RECT  12.5375 31.46 12.6075 31.595 ;
        RECT  12.5375 31.46 12.6075 31.595 ;
        RECT  12.5375 31.46 12.6075 31.595 ;
        RECT  12.0875 31.9525 12.1575 32.0875 ;
        RECT  11.8325 31.46 11.9025 31.595 ;
        RECT  11.8325 31.46 11.9025 31.595 ;
        RECT  11.8325 31.46 11.9025 31.595 ;
        RECT  11.8325 31.46 11.9025 31.595 ;
        RECT  11.8325 31.46 11.9025 31.595 ;
        RECT  11.8325 31.46 11.9025 31.595 ;
        RECT  12.5375 31.46 12.6075 31.595 ;
        RECT  12.5375 31.46 12.6075 31.595 ;
        RECT  12.5375 31.46 12.6075 31.595 ;
        RECT  12.5375 31.46 12.6075 31.595 ;
        RECT  12.2825 31.9525 12.3525 32.0875 ;
        RECT  12.505 32.31 12.64 32.38 ;
        RECT  12.505 32.31 12.64 32.38 ;
        RECT  12.505 32.31 12.64 32.38 ;
        RECT  12.5375 31.46 12.6075 31.595 ;
        RECT  12.5375 31.46 12.6075 31.595 ;
        RECT  12.5375 31.46 12.6075 31.595 ;
        RECT  12.5375 31.46 12.6075 31.595 ;
        RECT  12.5375 31.46 12.6075 31.595 ;
        RECT  12.5375 31.46 12.6075 31.595 ;
        RECT  11.8 32.31 11.935 32.38 ;
        RECT  12.5375 30.9675 12.6075 32.3775 ;
        RECT  11.8375 32.3175 11.8975 32.375 ;
        RECT  12.025 32.3175 12.08 32.37 ;
        RECT  12.36 32.3175 12.4175 32.3775 ;
        RECT  12.5425 32.3125 12.6025 32.37 ;
        RECT  12.3525 30.9 12.4225 32.445 ;
        RECT  12.0175 30.9 12.0875 32.445 ;
        RECT  11.8325 30.9 11.9025 32.445 ;
        RECT  12.5375 30.9 12.6075 32.445 ;
        RECT  12.5375 33.095 12.6075 33.23 ;
        RECT  12.5375 33.095 12.6075 33.23 ;
        RECT  12.5375 33.095 12.6075 33.23 ;
        RECT  12.5375 33.095 12.6075 33.23 ;
        RECT  12.5375 33.095 12.6075 33.23 ;
        RECT  12.5375 33.095 12.6075 33.23 ;
        RECT  11.8 32.31 11.935 32.38 ;
        RECT  12.505 32.31 12.64 32.38 ;
        RECT  12.5375 33.095 12.6075 33.23 ;
        RECT  12.5375 33.095 12.6075 33.23 ;
        RECT  12.5375 33.095 12.6075 33.23 ;
        RECT  12.5375 33.095 12.6075 33.23 ;
        RECT  12.5375 33.095 12.6075 33.23 ;
        RECT  12.5375 33.095 12.6075 33.23 ;
        RECT  12.5375 33.095 12.6075 33.23 ;
        RECT  12.5375 33.095 12.6075 33.23 ;
        RECT  12.0875 32.6025 12.1575 32.7375 ;
        RECT  11.8325 33.095 11.9025 33.23 ;
        RECT  11.8325 33.095 11.9025 33.23 ;
        RECT  11.8325 33.095 11.9025 33.23 ;
        RECT  11.8325 33.095 11.9025 33.23 ;
        RECT  11.8325 33.095 11.9025 33.23 ;
        RECT  11.8325 33.095 11.9025 33.23 ;
        RECT  12.5375 33.095 12.6075 33.23 ;
        RECT  12.5375 33.095 12.6075 33.23 ;
        RECT  12.5375 33.095 12.6075 33.23 ;
        RECT  12.5375 33.095 12.6075 33.23 ;
        RECT  12.2825 32.6025 12.3525 32.7375 ;
        RECT  12.505 32.31 12.64 32.38 ;
        RECT  12.505 32.31 12.64 32.38 ;
        RECT  12.505 32.31 12.64 32.38 ;
        RECT  12.5375 33.095 12.6075 33.23 ;
        RECT  12.5375 33.095 12.6075 33.23 ;
        RECT  12.5375 33.095 12.6075 33.23 ;
        RECT  12.5375 33.095 12.6075 33.23 ;
        RECT  12.5375 33.095 12.6075 33.23 ;
        RECT  12.5375 33.095 12.6075 33.23 ;
        RECT  11.8 32.31 11.935 32.38 ;
        RECT  12.5375 32.3125 12.6075 33.7225 ;
        RECT  11.8375 32.315 11.8975 32.3725 ;
        RECT  12.025 32.32 12.08 32.3725 ;
        RECT  12.36 32.3125 12.4175 32.3725 ;
        RECT  12.5425 32.32 12.6025 32.3775 ;
        RECT  12.3525 32.245 12.4225 33.79 ;
        RECT  12.0175 32.245 12.0875 33.79 ;
        RECT  11.8325 32.245 11.9025 33.79 ;
        RECT  12.5375 32.245 12.6075 33.79 ;
        RECT  12.5375 34.15 12.6075 34.285 ;
        RECT  12.5375 34.15 12.6075 34.285 ;
        RECT  12.5375 34.15 12.6075 34.285 ;
        RECT  12.5375 34.15 12.6075 34.285 ;
        RECT  12.5375 34.15 12.6075 34.285 ;
        RECT  12.5375 34.15 12.6075 34.285 ;
        RECT  11.8 35.0 11.935 35.07 ;
        RECT  12.505 35.0 12.64 35.07 ;
        RECT  12.5375 34.15 12.6075 34.285 ;
        RECT  12.5375 34.15 12.6075 34.285 ;
        RECT  12.5375 34.15 12.6075 34.285 ;
        RECT  12.5375 34.15 12.6075 34.285 ;
        RECT  12.5375 34.15 12.6075 34.285 ;
        RECT  12.5375 34.15 12.6075 34.285 ;
        RECT  12.5375 34.15 12.6075 34.285 ;
        RECT  12.5375 34.15 12.6075 34.285 ;
        RECT  12.0875 34.6425 12.1575 34.7775 ;
        RECT  11.8325 34.15 11.9025 34.285 ;
        RECT  11.8325 34.15 11.9025 34.285 ;
        RECT  11.8325 34.15 11.9025 34.285 ;
        RECT  11.8325 34.15 11.9025 34.285 ;
        RECT  11.8325 34.15 11.9025 34.285 ;
        RECT  11.8325 34.15 11.9025 34.285 ;
        RECT  12.5375 34.15 12.6075 34.285 ;
        RECT  12.5375 34.15 12.6075 34.285 ;
        RECT  12.5375 34.15 12.6075 34.285 ;
        RECT  12.5375 34.15 12.6075 34.285 ;
        RECT  12.2825 34.6425 12.3525 34.7775 ;
        RECT  12.505 35.0 12.64 35.07 ;
        RECT  12.505 35.0 12.64 35.07 ;
        RECT  12.505 35.0 12.64 35.07 ;
        RECT  12.5375 34.15 12.6075 34.285 ;
        RECT  12.5375 34.15 12.6075 34.285 ;
        RECT  12.5375 34.15 12.6075 34.285 ;
        RECT  12.5375 34.15 12.6075 34.285 ;
        RECT  12.5375 34.15 12.6075 34.285 ;
        RECT  12.5375 34.15 12.6075 34.285 ;
        RECT  11.8 35.0 11.935 35.07 ;
        RECT  12.5375 33.6575 12.6075 35.0675 ;
        RECT  11.8375 35.0075 11.8975 35.065 ;
        RECT  12.025 35.0075 12.08 35.06 ;
        RECT  12.36 35.0075 12.4175 35.0675 ;
        RECT  12.5425 35.0025 12.6025 35.06 ;
        RECT  12.3525 33.59 12.4225 35.135 ;
        RECT  12.0175 33.59 12.0875 35.135 ;
        RECT  11.8325 33.59 11.9025 35.135 ;
        RECT  12.5375 33.59 12.6075 35.135 ;
        RECT  12.5375 35.785 12.6075 35.92 ;
        RECT  12.5375 35.785 12.6075 35.92 ;
        RECT  12.5375 35.785 12.6075 35.92 ;
        RECT  12.5375 35.785 12.6075 35.92 ;
        RECT  12.5375 35.785 12.6075 35.92 ;
        RECT  12.5375 35.785 12.6075 35.92 ;
        RECT  11.8 35.0 11.935 35.07 ;
        RECT  12.505 35.0 12.64 35.07 ;
        RECT  12.5375 35.785 12.6075 35.92 ;
        RECT  12.5375 35.785 12.6075 35.92 ;
        RECT  12.5375 35.785 12.6075 35.92 ;
        RECT  12.5375 35.785 12.6075 35.92 ;
        RECT  12.5375 35.785 12.6075 35.92 ;
        RECT  12.5375 35.785 12.6075 35.92 ;
        RECT  12.5375 35.785 12.6075 35.92 ;
        RECT  12.5375 35.785 12.6075 35.92 ;
        RECT  12.0875 35.2925 12.1575 35.4275 ;
        RECT  11.8325 35.785 11.9025 35.92 ;
        RECT  11.8325 35.785 11.9025 35.92 ;
        RECT  11.8325 35.785 11.9025 35.92 ;
        RECT  11.8325 35.785 11.9025 35.92 ;
        RECT  11.8325 35.785 11.9025 35.92 ;
        RECT  11.8325 35.785 11.9025 35.92 ;
        RECT  12.5375 35.785 12.6075 35.92 ;
        RECT  12.5375 35.785 12.6075 35.92 ;
        RECT  12.5375 35.785 12.6075 35.92 ;
        RECT  12.5375 35.785 12.6075 35.92 ;
        RECT  12.2825 35.2925 12.3525 35.4275 ;
        RECT  12.505 35.0 12.64 35.07 ;
        RECT  12.505 35.0 12.64 35.07 ;
        RECT  12.505 35.0 12.64 35.07 ;
        RECT  12.5375 35.785 12.6075 35.92 ;
        RECT  12.5375 35.785 12.6075 35.92 ;
        RECT  12.5375 35.785 12.6075 35.92 ;
        RECT  12.5375 35.785 12.6075 35.92 ;
        RECT  12.5375 35.785 12.6075 35.92 ;
        RECT  12.5375 35.785 12.6075 35.92 ;
        RECT  11.8 35.0 11.935 35.07 ;
        RECT  12.5375 35.0025 12.6075 36.4125 ;
        RECT  11.8375 35.005 11.8975 35.0625 ;
        RECT  12.025 35.01 12.08 35.0625 ;
        RECT  12.36 35.0025 12.4175 35.0625 ;
        RECT  12.5425 35.01 12.6025 35.0675 ;
        RECT  12.3525 34.935 12.4225 36.48 ;
        RECT  12.0175 34.935 12.0875 36.48 ;
        RECT  11.8325 34.935 11.9025 36.48 ;
        RECT  12.5375 34.935 12.6075 36.48 ;
        RECT  12.5375 36.84 12.6075 36.975 ;
        RECT  12.5375 36.84 12.6075 36.975 ;
        RECT  12.5375 36.84 12.6075 36.975 ;
        RECT  12.5375 36.84 12.6075 36.975 ;
        RECT  12.5375 36.84 12.6075 36.975 ;
        RECT  12.5375 36.84 12.6075 36.975 ;
        RECT  11.8 37.69 11.935 37.76 ;
        RECT  12.505 37.69 12.64 37.76 ;
        RECT  12.5375 36.84 12.6075 36.975 ;
        RECT  12.5375 36.84 12.6075 36.975 ;
        RECT  12.5375 36.84 12.6075 36.975 ;
        RECT  12.5375 36.84 12.6075 36.975 ;
        RECT  12.5375 36.84 12.6075 36.975 ;
        RECT  12.5375 36.84 12.6075 36.975 ;
        RECT  12.5375 36.84 12.6075 36.975 ;
        RECT  12.5375 36.84 12.6075 36.975 ;
        RECT  12.0875 37.3325 12.1575 37.4675 ;
        RECT  11.8325 36.84 11.9025 36.975 ;
        RECT  11.8325 36.84 11.9025 36.975 ;
        RECT  11.8325 36.84 11.9025 36.975 ;
        RECT  11.8325 36.84 11.9025 36.975 ;
        RECT  11.8325 36.84 11.9025 36.975 ;
        RECT  11.8325 36.84 11.9025 36.975 ;
        RECT  12.5375 36.84 12.6075 36.975 ;
        RECT  12.5375 36.84 12.6075 36.975 ;
        RECT  12.5375 36.84 12.6075 36.975 ;
        RECT  12.5375 36.84 12.6075 36.975 ;
        RECT  12.2825 37.3325 12.3525 37.4675 ;
        RECT  12.505 37.69 12.64 37.76 ;
        RECT  12.505 37.69 12.64 37.76 ;
        RECT  12.505 37.69 12.64 37.76 ;
        RECT  12.5375 36.84 12.6075 36.975 ;
        RECT  12.5375 36.84 12.6075 36.975 ;
        RECT  12.5375 36.84 12.6075 36.975 ;
        RECT  12.5375 36.84 12.6075 36.975 ;
        RECT  12.5375 36.84 12.6075 36.975 ;
        RECT  12.5375 36.84 12.6075 36.975 ;
        RECT  11.8 37.69 11.935 37.76 ;
        RECT  12.5375 36.3475 12.6075 37.7575 ;
        RECT  11.8375 37.6975 11.8975 37.755 ;
        RECT  12.025 37.6975 12.08 37.75 ;
        RECT  12.36 37.6975 12.4175 37.7575 ;
        RECT  12.5425 37.6925 12.6025 37.75 ;
        RECT  12.3525 36.28 12.4225 37.825 ;
        RECT  12.0175 36.28 12.0875 37.825 ;
        RECT  11.8325 36.28 11.9025 37.825 ;
        RECT  12.5375 36.28 12.6075 37.825 ;
        RECT  12.5375 38.475 12.6075 38.61 ;
        RECT  12.5375 38.475 12.6075 38.61 ;
        RECT  12.5375 38.475 12.6075 38.61 ;
        RECT  12.5375 38.475 12.6075 38.61 ;
        RECT  12.5375 38.475 12.6075 38.61 ;
        RECT  12.5375 38.475 12.6075 38.61 ;
        RECT  11.8 37.69 11.935 37.76 ;
        RECT  12.505 37.69 12.64 37.76 ;
        RECT  12.5375 38.475 12.6075 38.61 ;
        RECT  12.5375 38.475 12.6075 38.61 ;
        RECT  12.5375 38.475 12.6075 38.61 ;
        RECT  12.5375 38.475 12.6075 38.61 ;
        RECT  12.5375 38.475 12.6075 38.61 ;
        RECT  12.5375 38.475 12.6075 38.61 ;
        RECT  12.5375 38.475 12.6075 38.61 ;
        RECT  12.5375 38.475 12.6075 38.61 ;
        RECT  12.0875 37.9825 12.1575 38.1175 ;
        RECT  11.8325 38.475 11.9025 38.61 ;
        RECT  11.8325 38.475 11.9025 38.61 ;
        RECT  11.8325 38.475 11.9025 38.61 ;
        RECT  11.8325 38.475 11.9025 38.61 ;
        RECT  11.8325 38.475 11.9025 38.61 ;
        RECT  11.8325 38.475 11.9025 38.61 ;
        RECT  12.5375 38.475 12.6075 38.61 ;
        RECT  12.5375 38.475 12.6075 38.61 ;
        RECT  12.5375 38.475 12.6075 38.61 ;
        RECT  12.5375 38.475 12.6075 38.61 ;
        RECT  12.2825 37.9825 12.3525 38.1175 ;
        RECT  12.505 37.69 12.64 37.76 ;
        RECT  12.505 37.69 12.64 37.76 ;
        RECT  12.505 37.69 12.64 37.76 ;
        RECT  12.5375 38.475 12.6075 38.61 ;
        RECT  12.5375 38.475 12.6075 38.61 ;
        RECT  12.5375 38.475 12.6075 38.61 ;
        RECT  12.5375 38.475 12.6075 38.61 ;
        RECT  12.5375 38.475 12.6075 38.61 ;
        RECT  12.5375 38.475 12.6075 38.61 ;
        RECT  11.8 37.69 11.935 37.76 ;
        RECT  12.5375 37.6925 12.6075 39.1025 ;
        RECT  11.8375 37.695 11.8975 37.7525 ;
        RECT  12.025 37.7 12.08 37.7525 ;
        RECT  12.36 37.6925 12.4175 37.7525 ;
        RECT  12.5425 37.7 12.6025 37.7575 ;
        RECT  12.3525 37.625 12.4225 39.17 ;
        RECT  12.0175 37.625 12.0875 39.17 ;
        RECT  11.8325 37.625 11.9025 39.17 ;
        RECT  12.5375 37.625 12.6075 39.17 ;
        RECT  12.5375 39.53 12.6075 39.665 ;
        RECT  12.5375 39.53 12.6075 39.665 ;
        RECT  12.5375 39.53 12.6075 39.665 ;
        RECT  12.5375 39.53 12.6075 39.665 ;
        RECT  12.5375 39.53 12.6075 39.665 ;
        RECT  12.5375 39.53 12.6075 39.665 ;
        RECT  11.8 40.38 11.935 40.45 ;
        RECT  12.505 40.38 12.64 40.45 ;
        RECT  12.5375 39.53 12.6075 39.665 ;
        RECT  12.5375 39.53 12.6075 39.665 ;
        RECT  12.5375 39.53 12.6075 39.665 ;
        RECT  12.5375 39.53 12.6075 39.665 ;
        RECT  12.5375 39.53 12.6075 39.665 ;
        RECT  12.5375 39.53 12.6075 39.665 ;
        RECT  12.5375 39.53 12.6075 39.665 ;
        RECT  12.5375 39.53 12.6075 39.665 ;
        RECT  12.0875 40.0225 12.1575 40.1575 ;
        RECT  11.8325 39.53 11.9025 39.665 ;
        RECT  11.8325 39.53 11.9025 39.665 ;
        RECT  11.8325 39.53 11.9025 39.665 ;
        RECT  11.8325 39.53 11.9025 39.665 ;
        RECT  11.8325 39.53 11.9025 39.665 ;
        RECT  11.8325 39.53 11.9025 39.665 ;
        RECT  12.5375 39.53 12.6075 39.665 ;
        RECT  12.5375 39.53 12.6075 39.665 ;
        RECT  12.5375 39.53 12.6075 39.665 ;
        RECT  12.5375 39.53 12.6075 39.665 ;
        RECT  12.2825 40.0225 12.3525 40.1575 ;
        RECT  12.505 40.38 12.64 40.45 ;
        RECT  12.505 40.38 12.64 40.45 ;
        RECT  12.505 40.38 12.64 40.45 ;
        RECT  12.5375 39.53 12.6075 39.665 ;
        RECT  12.5375 39.53 12.6075 39.665 ;
        RECT  12.5375 39.53 12.6075 39.665 ;
        RECT  12.5375 39.53 12.6075 39.665 ;
        RECT  12.5375 39.53 12.6075 39.665 ;
        RECT  12.5375 39.53 12.6075 39.665 ;
        RECT  11.8 40.38 11.935 40.45 ;
        RECT  12.5375 39.0375 12.6075 40.4475 ;
        RECT  11.8375 40.3875 11.8975 40.445 ;
        RECT  12.025 40.3875 12.08 40.44 ;
        RECT  12.36 40.3875 12.4175 40.4475 ;
        RECT  12.5425 40.3825 12.6025 40.44 ;
        RECT  12.3525 38.97 12.4225 40.515 ;
        RECT  12.0175 38.97 12.0875 40.515 ;
        RECT  11.8325 38.97 11.9025 40.515 ;
        RECT  12.5375 38.97 12.6075 40.515 ;
        RECT  11.3125 40.765 11.3825 41.725 ;
        RECT  11.6475 40.765 11.7175 41.725 ;
        RECT  11.3475 41.3125 11.39 41.4475 ;
        RECT  11.6475 41.3125 11.735 41.4475 ;
        RECT  11.3475 40.8625 11.3925 40.9975 ;
        RECT  11.5475 40.8625 11.6475 40.9975 ;
        RECT  11.355 41.3125 11.425 41.4475 ;
        RECT  11.735 41.3125 11.805 41.4475 ;
        RECT  11.355 40.8625 11.425 40.9975 ;
        RECT  11.545 40.8625 11.615 40.9975 ;
        RECT  12.0175 40.765 12.0875 41.725 ;
        RECT  12.3525 40.765 12.4225 41.725 ;
        RECT  12.0525 41.3125 12.095 41.4475 ;
        RECT  12.3525 41.3125 12.44 41.4475 ;
        RECT  12.0525 40.8625 12.0975 40.9975 ;
        RECT  12.2525 40.8625 12.3525 40.9975 ;
        RECT  12.06 41.3125 12.13 41.4475 ;
        RECT  12.44 41.3125 12.51 41.4475 ;
        RECT  12.06 40.8625 12.13 40.9975 ;
        RECT  12.25 40.8625 12.32 40.9975 ;
        RECT  11.475 18.755 11.545 18.895 ;
        RECT  11.475 18.4975 11.545 18.6325 ;
        RECT  11.8325 14.2575 11.9025 14.3925 ;
        RECT  11.1275 14.2575 11.1975 14.3925 ;
        RECT  11.67 17.04 11.74 17.175 ;
        RECT  11.2875 17.45 11.3575 17.585 ;
        RECT  11.48 18.2925 11.55 18.4275 ;
        RECT  11.48 16.15 11.55 16.285 ;
        RECT  11.475 18.4975 11.545 18.895 ;
        RECT  11.475 18.84 11.545 18.895 ;
        RECT  11.3125 18.835 11.3825 18.895 ;
        RECT  11.6525 18.845 11.7125 18.895 ;
        RECT  11.8325 14.01 11.9025 18.895 ;
        RECT  11.6475 14.81 11.7175 18.895 ;
        RECT  11.48 16.285 11.55 18.295 ;
        RECT  11.6475 14.01 11.7175 17.555 ;
        RECT  11.3125 14.01 11.3825 18.895 ;
        RECT  11.1275 14.01 11.1975 18.895 ;
        RECT  12.18 18.755 12.25 18.895 ;
        RECT  12.18 18.4975 12.25 18.6325 ;
        RECT  12.5375 14.2575 12.6075 14.3925 ;
        RECT  11.8325 14.2575 11.9025 14.3925 ;
        RECT  12.375 17.04 12.445 17.175 ;
        RECT  11.9925 17.45 12.0625 17.585 ;
        RECT  12.185 18.2925 12.255 18.4275 ;
        RECT  12.185 16.15 12.255 16.285 ;
        RECT  12.18 18.4975 12.25 18.895 ;
        RECT  12.18 18.84 12.25 18.895 ;
        RECT  12.0175 18.835 12.0875 18.895 ;
        RECT  12.3575 18.845 12.4175 18.895 ;
        RECT  12.5375 14.01 12.6075 18.895 ;
        RECT  12.3525 14.81 12.4225 18.895 ;
        RECT  12.185 16.285 12.255 18.295 ;
        RECT  12.3525 14.01 12.4225 17.555 ;
        RECT  12.0175 14.01 12.0875 18.895 ;
        RECT  11.8325 14.01 11.9025 18.895 ;
        RECT  11.37 9.9675 11.505 10.0375 ;
        RECT  11.48 9.835 11.55 9.975 ;
        RECT  11.8325 11.57 11.9025 11.705 ;
        RECT  11.8325 11.0 11.9025 11.135 ;
        RECT  11.1275 11.0 11.1975 11.135 ;
        RECT  11.5475 11.205 11.6175 11.34 ;
        RECT  11.8325 13.4975 11.9025 13.6325 ;
        RECT  11.5475 10.795 11.6175 10.93 ;
        RECT  11.4075 10.795 11.4775 10.93 ;
        RECT  11.8325 11.205 11.9025 11.34 ;
        RECT  11.1275 11.205 11.1975 11.34 ;
        RECT  11.2675 10.23 11.4025 10.3 ;
        RECT  11.4075 13.175 11.4775 13.31 ;
        RECT  11.5775 11.57 11.6475 11.705 ;
        RECT  11.2675 12.485 11.3375 12.62 ;
        RECT  11.4075 11.205 11.4775 11.34 ;
        RECT  11.1275 11.57 11.1975 11.705 ;
        RECT  11.5775 12.085 11.6475 12.22 ;
        RECT  11.3125 13.7075 11.3825 13.8425 ;
        RECT  11.1275 13.4975 11.1975 13.6325 ;
        RECT  11.3125 13.71 11.3825 14.01 ;
        RECT  11.3125 13.945 11.3825 14.01 ;
        RECT  11.65 13.95 11.715 14.01 ;
        RECT  11.4825 9.84 11.5475 9.9025 ;
        RECT  11.8325 9.835 11.9025 14.01 ;
        RECT  11.1275 9.835 11.1975 14.01 ;
        RECT  11.6475 11.57 11.7175 14.01 ;
        RECT  11.3575 9.9675 11.55 10.0375 ;
        RECT  11.5475 10.93 11.6175 11.205 ;
        RECT  11.2675 10.3 11.3375 12.62 ;
        RECT  11.4075 10.93 11.4775 11.205 ;
        RECT  11.4075 11.205 11.4775 13.3025 ;
        RECT  12.075 9.9675 12.21 10.0375 ;
        RECT  12.185 9.835 12.255 9.975 ;
        RECT  12.5375 11.57 12.6075 11.705 ;
        RECT  12.5375 11.0 12.6075 11.135 ;
        RECT  11.8325 11.0 11.9025 11.135 ;
        RECT  12.2525 11.205 12.3225 11.34 ;
        RECT  12.5375 13.4975 12.6075 13.6325 ;
        RECT  12.2525 10.795 12.3225 10.93 ;
        RECT  12.1125 10.795 12.1825 10.93 ;
        RECT  12.5375 11.205 12.6075 11.34 ;
        RECT  11.8325 11.205 11.9025 11.34 ;
        RECT  11.9725 10.23 12.1075 10.3 ;
        RECT  12.1125 13.175 12.1825 13.31 ;
        RECT  12.2825 11.57 12.3525 11.705 ;
        RECT  11.9725 12.485 12.0425 12.62 ;
        RECT  12.1125 11.205 12.1825 11.34 ;
        RECT  11.8325 11.57 11.9025 11.705 ;
        RECT  12.2825 12.085 12.3525 12.22 ;
        RECT  12.0175 13.7075 12.0875 13.8425 ;
        RECT  11.8325 13.4975 11.9025 13.6325 ;
        RECT  12.0175 13.71 12.0875 14.01 ;
        RECT  12.0175 13.945 12.0875 14.01 ;
        RECT  12.355 13.95 12.42 14.01 ;
        RECT  12.1875 9.84 12.2525 9.9025 ;
        RECT  12.5375 9.835 12.6075 14.01 ;
        RECT  11.8325 9.835 11.9025 14.01 ;
        RECT  12.3525 11.57 12.4225 14.01 ;
        RECT  12.0625 9.9675 12.255 10.0375 ;
        RECT  12.2525 10.93 12.3225 11.205 ;
        RECT  11.9725 10.3 12.0425 12.62 ;
        RECT  12.1125 10.93 12.1825 11.205 ;
        RECT  12.1125 11.205 12.1825 13.3025 ;
        RECT  11.325 9.0975 11.395 9.2325 ;
        RECT  11.8325 3.92 11.9025 4.055 ;
        RECT  11.69 8.0025 11.76 8.1375 ;
        RECT  11.6925 6.395 11.7625 6.53 ;
        RECT  11.6925 4.9975 11.7625 5.1325 ;
        RECT  11.1275 3.78 11.1975 3.915 ;
        RECT  11.48 3.395 11.55 3.535 ;
        RECT  11.8325 6.8575 11.9025 6.9925 ;
        RECT  11.3275 5.6625 11.3975 5.7975 ;
        RECT  11.6925 9.355 11.7625 9.49 ;
        RECT  11.515 8.845 11.585 8.98 ;
        RECT  11.8325 8.4325 11.9025 8.5675 ;
        RECT  11.8325 3.73 11.9025 3.865 ;
        RECT  11.8325 5.4725 11.9025 5.6075 ;
        RECT  11.3275 5.2725 11.3975 5.4075 ;
        RECT  11.515 5.2725 11.585 5.4075 ;
        RECT  11.515 5.885 11.585 6.02 ;
        RECT  11.325 8.2325 11.395 8.3675 ;
        RECT  11.515 8.2325 11.585 8.3675 ;
        RECT  11.55 9.565 11.6925 9.635 ;
        RECT  11.48 3.395 11.55 3.54 ;
        RECT  11.545 3.47 11.6925 3.54 ;
        RECT  11.48 9.565 11.55 9.835 ;
        RECT  11.13 9.3575 11.1925 9.4175 ;
        RECT  11.1275 3.395 11.1975 9.835 ;
        RECT  11.4825 9.77 11.5475 9.83 ;
        RECT  11.6925 9.355 11.7625 9.635 ;
        RECT  11.6925 3.47 11.7625 5.1325 ;
        RECT  11.325 9.1475 11.395 9.835 ;
        RECT  11.6925 6.53 11.7625 8.1375 ;
        RECT  11.515 8.2325 11.585 8.95 ;
        RECT  11.3275 5.2725 11.3975 5.7975 ;
        RECT  11.33 9.6975 11.3925 9.7575 ;
        RECT  11.325 8.2325 11.395 9.1725 ;
        RECT  11.48 3.4 11.5475 3.465 ;
        RECT  11.8325 3.395 11.9025 9.835 ;
        RECT  11.515 5.2725 11.585 5.99 ;
        RECT  12.34 9.0975 12.41 9.2325 ;
        RECT  11.8325 3.92 11.9025 4.055 ;
        RECT  11.975 8.0025 12.045 8.1375 ;
        RECT  11.9725 6.395 12.0425 6.53 ;
        RECT  11.9725 4.9975 12.0425 5.1325 ;
        RECT  12.5375 3.78 12.6075 3.915 ;
        RECT  12.185 3.395 12.255 3.535 ;
        RECT  11.8325 6.8575 11.9025 6.9925 ;
        RECT  12.3375 5.6625 12.4075 5.7975 ;
        RECT  11.9725 9.355 12.0425 9.49 ;
        RECT  12.15 8.845 12.22 8.98 ;
        RECT  11.8325 8.4325 11.9025 8.5675 ;
        RECT  11.8325 3.73 11.9025 3.865 ;
        RECT  11.8325 5.4725 11.9025 5.6075 ;
        RECT  12.3375 5.2725 12.4075 5.4075 ;
        RECT  12.15 5.2725 12.22 5.4075 ;
        RECT  12.15 5.885 12.22 6.02 ;
        RECT  12.34 8.2325 12.41 8.3675 ;
        RECT  12.15 8.2325 12.22 8.3675 ;
        RECT  12.0425 9.565 12.185 9.635 ;
        RECT  12.185 3.395 12.255 3.54 ;
        RECT  12.0425 3.47 12.19 3.54 ;
        RECT  12.185 9.565 12.255 9.835 ;
        RECT  12.5425 9.3575 12.605 9.4175 ;
        RECT  12.5375 3.395 12.6075 9.835 ;
        RECT  12.1875 9.77 12.2525 9.83 ;
        RECT  11.9725 9.355 12.0425 9.635 ;
        RECT  11.9725 3.47 12.0425 5.1325 ;
        RECT  12.34 9.1475 12.41 9.835 ;
        RECT  11.9725 6.53 12.0425 8.1375 ;
        RECT  12.15 8.2325 12.22 8.95 ;
        RECT  12.3375 5.2725 12.4075 5.7975 ;
        RECT  12.3425 9.6975 12.405 9.7575 ;
        RECT  12.34 8.2325 12.41 9.1725 ;
        RECT  12.1875 3.4 12.255 3.465 ;
        RECT  11.8325 3.395 11.9025 9.835 ;
        RECT  12.15 5.2725 12.22 5.99 ;
        RECT  11.4475 5.1775 11.5825 5.2475 ;
        RECT  11.8325 3.8925 11.9025 4.0275 ;
        RECT  11.48 3.5475 11.55 3.6875 ;
        RECT  11.58 5.8175 11.715 5.8875 ;
        RECT  11.8325 5.9525 11.9025 6.0875 ;
        RECT  11.305 5.7625 11.375 5.8975 ;
        RECT  11.5125 5.485 11.5825 5.62 ;
        RECT  11.2675 3.675 11.48 3.745 ;
        RECT  11.48 3.395 11.55 3.745 ;
        RECT  11.55 6.13 11.6525 6.2 ;
        RECT  11.48 6.13 11.55 6.37 ;
        RECT  11.48 6.3125 11.55 6.365 ;
        RECT  11.48 3.55 11.55 3.6125 ;
        RECT  11.27 4.31 11.34 5.8975 ;
        RECT  11.6525 5.8175 11.7225 6.2 ;
        RECT  11.5125 5.2475 11.5825 5.485 ;
        RECT  11.8325 3.395 11.9025 6.37 ;
        RECT  11.8325 3.9675 11.9025 4.025 ;
        RECT  11.58 4.31 11.715 4.38 ;
        RECT  11.34 4.31 11.58 4.38 ;
        RECT  11.2675 3.675 11.3375 4.045 ;
        RECT  11.2675 4.045 11.3375 4.18 ;
        RECT  12.1525 5.1775 12.2875 5.2475 ;
        RECT  11.8325 3.8925 11.9025 4.0275 ;
        RECT  12.185 3.5475 12.255 3.6875 ;
        RECT  12.02 5.8175 12.155 5.8875 ;
        RECT  11.8325 5.9525 11.9025 6.0875 ;
        RECT  12.36 5.7625 12.43 5.8975 ;
        RECT  12.1525 5.485 12.2225 5.62 ;
        RECT  12.255 3.675 12.4675 3.745 ;
        RECT  12.185 3.395 12.255 3.745 ;
        RECT  12.0825 6.13 12.185 6.2 ;
        RECT  12.185 6.13 12.255 6.37 ;
        RECT  12.185 6.3125 12.255 6.365 ;
        RECT  12.185 3.55 12.255 3.6125 ;
        RECT  12.395 4.31 12.465 5.8975 ;
        RECT  12.0125 5.8175 12.0825 6.2 ;
        RECT  12.1525 5.2475 12.2225 5.485 ;
        RECT  11.8325 3.395 11.9025 6.37 ;
        RECT  11.8325 3.9675 11.9025 4.025 ;
        RECT  12.02 4.31 12.155 4.38 ;
        RECT  12.155 4.31 12.395 4.38 ;
        RECT  12.3975 3.675 12.4675 4.045 ;
        RECT  12.3975 4.045 12.4675 4.18 ;
        RECT  4.0775 8.135 4.1475 40.415 ;
        RECT  3.9025 8.135 3.9725 40.415 ;
        RECT  3.7275 8.135 3.7975 40.415 ;
        RECT  3.5525 8.135 3.6225 40.415 ;
        RECT  3.3775 8.135 3.4475 40.415 ;
        RECT  3.2025 8.135 3.2725 40.415 ;
        RECT  3.0275 8.135 3.0975 40.415 ;
        RECT  2.8525 8.135 2.9225 40.415 ;
        RECT  7.5575 8.135 7.6275 13.305 ;
        RECT  7.3825 8.135 7.4525 13.305 ;
        RECT  6.5425 8.135 6.6125 13.305 ;
        RECT  6.3675 8.135 6.4375 13.305 ;
        RECT  6.1925 8.135 6.2625 13.305 ;
        RECT  6.0175 8.135 6.0875 13.305 ;
        RECT  5.8425 8.135 5.9125 13.305 ;
        RECT  5.6675 8.135 5.7375 13.305 ;
        RECT  6.1575 9.18 6.2925 9.25 ;
        RECT  7.5225 8.6575 7.6575 8.7275 ;
        RECT  5.9825 9.57 6.1175 9.64 ;
        RECT  7.3475 10.0925 7.4825 10.1625 ;
        RECT  6.1575 8.9725 6.2925 9.0425 ;
        RECT  5.9825 8.4425 6.1175 8.5125 ;
        RECT  5.8075 9.7775 5.9425 9.8475 ;
        RECT  5.9825 10.3075 6.1175 10.3775 ;
        RECT  6.1575 11.6625 6.2925 11.7325 ;
        RECT  5.6325 11.1325 5.7675 11.2025 ;
        RECT  5.8075 12.4675 5.9425 12.5375 ;
        RECT  7.5225 12.4675 7.6575 12.5375 ;
        RECT  5.6325 12.9975 5.7675 13.0675 ;
        RECT  7.3475 12.9975 7.4825 13.0675 ;
        RECT  6.3325 8.03 6.4675 8.1 ;
        RECT  6.5075 9.375 6.6425 9.445 ;
        RECT  6.3325 10.72 6.4675 10.79 ;
        RECT  6.5075 12.065 6.6425 12.135 ;
        RECT  6.3325 13.2325 6.4675 13.3025 ;
        RECT  7.5575 13.515 7.6275 18.685 ;
        RECT  7.3825 13.515 7.4525 18.685 ;
        RECT  6.5425 13.515 6.6125 18.685 ;
        RECT  6.3675 13.515 6.4375 18.685 ;
        RECT  6.1925 13.515 6.2625 18.685 ;
        RECT  6.0175 13.515 6.0875 18.685 ;
        RECT  5.8425 13.515 5.9125 18.685 ;
        RECT  5.6675 13.515 5.7375 18.685 ;
        RECT  6.1575 14.56 6.2925 14.63 ;
        RECT  7.5225 14.0375 7.6575 14.1075 ;
        RECT  5.9825 14.95 6.1175 15.02 ;
        RECT  7.3475 15.4725 7.4825 15.5425 ;
        RECT  6.1575 14.3525 6.2925 14.4225 ;
        RECT  5.9825 13.8225 6.1175 13.8925 ;
        RECT  5.8075 15.1575 5.9425 15.2275 ;
        RECT  5.9825 15.6875 6.1175 15.7575 ;
        RECT  6.1575 17.0425 6.2925 17.1125 ;
        RECT  5.6325 16.5125 5.7675 16.5825 ;
        RECT  5.8075 17.8475 5.9425 17.9175 ;
        RECT  7.5225 17.8475 7.6575 17.9175 ;
        RECT  5.6325 18.3775 5.7675 18.4475 ;
        RECT  7.3475 18.3775 7.4825 18.4475 ;
        RECT  6.3325 13.41 6.4675 13.48 ;
        RECT  6.5075 14.755 6.6425 14.825 ;
        RECT  6.3325 16.1 6.4675 16.17 ;
        RECT  6.5075 17.445 6.6425 17.515 ;
        RECT  6.3325 18.6125 6.4675 18.6825 ;
        RECT  2.8225 8.7275 2.9575 8.7975 ;
        RECT  2.9975 10.1625 3.1325 10.2325 ;
        RECT  3.1725 11.4175 3.3075 11.4875 ;
        RECT  3.3475 12.8525 3.4825 12.9225 ;
        RECT  3.5225 14.1075 3.6575 14.1775 ;
        RECT  3.6975 15.5425 3.8325 15.6125 ;
        RECT  3.8725 16.7975 4.0075 16.8675 ;
        RECT  4.0475 18.2325 4.1825 18.3025 ;
        RECT  2.8225 19.8025 2.9575 19.8725 ;
        RECT  3.5225 19.2725 3.6575 19.3425 ;
        RECT  2.8225 20.6075 2.9575 20.6775 ;
        RECT  3.6975 21.1375 3.8325 21.2075 ;
        RECT  2.8225 22.4925 2.9575 22.5625 ;
        RECT  3.8725 21.9625 4.0075 22.0325 ;
        RECT  2.8225 23.2975 2.9575 23.3675 ;
        RECT  4.0475 23.8275 4.1825 23.8975 ;
        RECT  2.9975 25.1825 3.1325 25.2525 ;
        RECT  3.5225 24.6525 3.6575 24.7225 ;
        RECT  2.9975 25.9875 3.1325 26.0575 ;
        RECT  3.6975 26.5175 3.8325 26.5875 ;
        RECT  2.9975 27.8725 3.1325 27.9425 ;
        RECT  3.8725 27.3425 4.0075 27.4125 ;
        RECT  2.9975 28.6775 3.1325 28.7475 ;
        RECT  4.0475 29.2075 4.1825 29.2775 ;
        RECT  3.1725 30.5625 3.3075 30.6325 ;
        RECT  3.5225 30.0325 3.6575 30.1025 ;
        RECT  3.1725 31.3675 3.3075 31.4375 ;
        RECT  3.6975 31.8975 3.8325 31.9675 ;
        RECT  3.1725 33.2525 3.3075 33.3225 ;
        RECT  3.8725 32.7225 4.0075 32.7925 ;
        RECT  3.1725 34.0575 3.3075 34.1275 ;
        RECT  4.0475 34.5875 4.1825 34.6575 ;
        RECT  3.3475 35.9425 3.4825 36.0125 ;
        RECT  3.5225 35.4125 3.6575 35.4825 ;
        RECT  3.3475 36.7475 3.4825 36.8175 ;
        RECT  3.6975 37.2775 3.8325 37.3475 ;
        RECT  3.3475 38.6325 3.4825 38.7025 ;
        RECT  3.8725 38.1025 4.0075 38.1725 ;
        RECT  3.3475 39.4375 3.4825 39.5075 ;
        RECT  4.0475 39.9675 4.1825 40.0375 ;
        RECT  5.5625 20.205 6.0175 20.275 ;
        RECT  5.5625 19.805 6.5775 19.875 ;
        RECT  5.5625 21.55 6.0175 21.62 ;
        RECT  5.5625 20.605 6.5775 20.675 ;
        RECT  5.5625 22.895 6.0175 22.965 ;
        RECT  5.5625 22.495 6.5775 22.565 ;
        RECT  5.5625 24.24 6.0175 24.31 ;
        RECT  5.5625 23.295 6.5775 23.365 ;
        RECT  5.5625 25.585 6.0175 25.655 ;
        RECT  5.5625 25.185 6.5775 25.255 ;
        RECT  5.5625 26.93 6.0175 27.0 ;
        RECT  5.5625 25.985 6.5775 26.055 ;
        RECT  5.5625 28.275 6.0175 28.345 ;
        RECT  5.5625 27.875 6.5775 27.945 ;
        RECT  5.5625 29.62 6.0175 29.69 ;
        RECT  5.5625 28.675 6.5775 28.745 ;
        RECT  5.5625 30.965 6.0175 31.035 ;
        RECT  5.5625 30.565 6.5775 30.635 ;
        RECT  5.5625 32.31 6.0175 32.38 ;
        RECT  5.5625 31.365 6.5775 31.435 ;
        RECT  5.5625 33.655 6.0175 33.725 ;
        RECT  5.5625 33.255 6.5775 33.325 ;
        RECT  5.5625 35.0 6.0175 35.07 ;
        RECT  5.5625 34.055 6.5775 34.125 ;
        RECT  5.5625 36.345 6.0175 36.415 ;
        RECT  5.5625 35.945 6.5775 36.015 ;
        RECT  5.5625 37.69 6.0175 37.76 ;
        RECT  5.5625 36.745 6.5775 36.815 ;
        RECT  5.5625 39.035 6.0175 39.105 ;
        RECT  5.5625 38.635 6.5775 38.705 ;
        RECT  5.5625 40.38 6.0175 40.45 ;
        RECT  5.5625 39.435 6.5775 39.505 ;
        RECT  5.4925 20.205 5.6275 20.275 ;
        RECT  5.9475 20.205 6.0825 20.275 ;
        RECT  6.5775 19.805 6.7125 19.875 ;
        RECT  5.5625 19.805 5.6325 19.94 ;
        RECT  5.4925 21.55 5.6275 21.62 ;
        RECT  5.9475 21.55 6.0825 21.62 ;
        RECT  6.5775 20.605 6.7125 20.675 ;
        RECT  5.5625 20.54 5.6325 20.675 ;
        RECT  5.4925 22.895 5.6275 22.965 ;
        RECT  5.9475 22.895 6.0825 22.965 ;
        RECT  6.5775 22.495 6.7125 22.565 ;
        RECT  5.5625 22.495 5.6325 22.63 ;
        RECT  5.4925 24.24 5.6275 24.31 ;
        RECT  5.9475 24.24 6.0825 24.31 ;
        RECT  6.5775 23.295 6.7125 23.365 ;
        RECT  5.5625 23.23 5.6325 23.365 ;
        RECT  5.4925 25.585 5.6275 25.655 ;
        RECT  5.9475 25.585 6.0825 25.655 ;
        RECT  6.5775 25.185 6.7125 25.255 ;
        RECT  5.5625 25.185 5.6325 25.32 ;
        RECT  5.4925 26.93 5.6275 27.0 ;
        RECT  5.9475 26.93 6.0825 27.0 ;
        RECT  6.5775 25.985 6.7125 26.055 ;
        RECT  5.5625 25.92 5.6325 26.055 ;
        RECT  5.4925 28.275 5.6275 28.345 ;
        RECT  5.9475 28.275 6.0825 28.345 ;
        RECT  6.5775 27.875 6.7125 27.945 ;
        RECT  5.5625 27.875 5.6325 28.01 ;
        RECT  5.4925 29.62 5.6275 29.69 ;
        RECT  5.9475 29.62 6.0825 29.69 ;
        RECT  6.5775 28.675 6.7125 28.745 ;
        RECT  5.5625 28.61 5.6325 28.745 ;
        RECT  5.4925 30.965 5.6275 31.035 ;
        RECT  5.9475 30.965 6.0825 31.035 ;
        RECT  6.5775 30.565 6.7125 30.635 ;
        RECT  5.5625 30.565 5.6325 30.7 ;
        RECT  5.4925 32.31 5.6275 32.38 ;
        RECT  5.9475 32.31 6.0825 32.38 ;
        RECT  6.5775 31.365 6.7125 31.435 ;
        RECT  5.5625 31.3 5.6325 31.435 ;
        RECT  5.4925 33.655 5.6275 33.725 ;
        RECT  5.9475 33.655 6.0825 33.725 ;
        RECT  6.5775 33.255 6.7125 33.325 ;
        RECT  5.5625 33.255 5.6325 33.39 ;
        RECT  5.4925 35.0 5.6275 35.07 ;
        RECT  5.9475 35.0 6.0825 35.07 ;
        RECT  6.5775 34.055 6.7125 34.125 ;
        RECT  5.5625 33.99 5.6325 34.125 ;
        RECT  5.4925 36.345 5.6275 36.415 ;
        RECT  5.9475 36.345 6.0825 36.415 ;
        RECT  6.5775 35.945 6.7125 36.015 ;
        RECT  5.5625 35.945 5.6325 36.08 ;
        RECT  5.4925 37.69 5.6275 37.76 ;
        RECT  5.9475 37.69 6.0825 37.76 ;
        RECT  6.5775 36.745 6.7125 36.815 ;
        RECT  5.5625 36.68 5.6325 36.815 ;
        RECT  5.4925 39.035 5.6275 39.105 ;
        RECT  5.9475 39.035 6.0825 39.105 ;
        RECT  6.5775 38.635 6.7125 38.705 ;
        RECT  5.5625 38.635 5.6325 38.77 ;
        RECT  5.4925 40.38 5.6275 40.45 ;
        RECT  5.9475 40.38 6.0825 40.45 ;
        RECT  6.5775 39.435 6.7125 39.505 ;
        RECT  5.5625 39.37 5.6325 39.505 ;
        RECT  6.645 7.6075 6.78 7.6775 ;
        RECT  1.4675 7.1 1.6025 7.17 ;
        RECT  5.55 7.2425 5.685 7.3125 ;
        RECT  3.9425 7.24 4.0775 7.31 ;
        RECT  2.545 7.24 2.68 7.31 ;
        RECT  1.3275 7.805 1.4625 7.875 ;
        RECT  0.9425 7.4525 1.0825 7.5225 ;
        RECT  4.405 7.1 4.54 7.17 ;
        RECT  3.21 7.605 3.345 7.675 ;
        RECT  6.9025 7.24 7.0375 7.31 ;
        RECT  6.3925 7.4175 6.5275 7.4875 ;
        RECT  5.98 7.1 6.115 7.17 ;
        RECT  1.2775 7.1 1.4125 7.17 ;
        RECT  3.02 7.1 3.155 7.17 ;
        RECT  2.82 7.605 2.955 7.675 ;
        RECT  2.82 7.4175 2.955 7.4875 ;
        RECT  3.4325 7.4175 3.5675 7.4875 ;
        RECT  5.78 7.6075 5.915 7.6775 ;
        RECT  5.78 7.4175 5.915 7.4875 ;
        RECT  7.1125 7.31 7.1825 7.4525 ;
        RECT  0.9425 7.4525 1.0875 7.5225 ;
        RECT  1.0175 7.31 1.0875 7.4575 ;
        RECT  7.1125 7.4525 7.3825 7.5225 ;
        RECT  6.905 7.81 6.965 7.8725 ;
        RECT  0.9425 7.805 7.3825 7.875 ;
        RECT  7.3175 7.455 7.3775 7.52 ;
        RECT  6.9025 7.24 7.1825 7.31 ;
        RECT  1.0175 7.24 2.68 7.31 ;
        RECT  6.695 7.6075 7.3825 7.6775 ;
        RECT  4.0775 7.24 5.685 7.31 ;
        RECT  5.78 7.4175 6.4975 7.4875 ;
        RECT  2.82 7.605 3.345 7.675 ;
        RECT  7.245 7.61 7.305 7.6725 ;
        RECT  5.78 7.6075 6.72 7.6775 ;
        RECT  0.9475 7.455 1.0125 7.5225 ;
        RECT  0.9425 7.1 7.3825 7.17 ;
        RECT  2.82 7.4175 3.5375 7.4875 ;
        RECT  6.645 6.5925 6.78 6.6625 ;
        RECT  1.4675 7.1 1.6025 7.17 ;
        RECT  5.55 6.9575 5.685 7.0275 ;
        RECT  3.9425 6.96 4.0775 7.03 ;
        RECT  2.545 6.96 2.68 7.03 ;
        RECT  1.3275 6.395 1.4625 6.465 ;
        RECT  0.9425 6.7475 1.0825 6.8175 ;
        RECT  4.405 7.1 4.54 7.17 ;
        RECT  3.21 6.595 3.345 6.665 ;
        RECT  6.9025 6.96 7.0375 7.03 ;
        RECT  6.3925 6.7825 6.5275 6.8525 ;
        RECT  5.98 7.1 6.115 7.17 ;
        RECT  1.2775 7.1 1.4125 7.17 ;
        RECT  3.02 7.1 3.155 7.17 ;
        RECT  2.82 6.595 2.955 6.665 ;
        RECT  2.82 6.7825 2.955 6.8525 ;
        RECT  3.4325 6.7825 3.5675 6.8525 ;
        RECT  5.78 6.5925 5.915 6.6625 ;
        RECT  5.78 6.7825 5.915 6.8525 ;
        RECT  7.1125 6.8175 7.1825 6.96 ;
        RECT  0.9425 6.7475 1.0875 6.8175 ;
        RECT  1.0175 6.8125 1.0875 6.96 ;
        RECT  7.1125 6.7475 7.3825 6.8175 ;
        RECT  6.905 6.3975 6.965 6.46 ;
        RECT  0.9425 6.395 7.3825 6.465 ;
        RECT  7.3175 6.75 7.3775 6.815 ;
        RECT  6.9025 6.96 7.1825 7.03 ;
        RECT  1.0175 6.96 2.68 7.03 ;
        RECT  6.695 6.5925 7.3825 6.6625 ;
        RECT  4.0775 6.96 5.685 7.03 ;
        RECT  5.78 6.7825 6.4975 6.8525 ;
        RECT  2.82 6.595 3.345 6.665 ;
        RECT  7.245 6.5975 7.305 6.66 ;
        RECT  5.78 6.5925 6.72 6.6625 ;
        RECT  0.9475 6.7475 1.0125 6.815 ;
        RECT  0.9425 7.1 7.3825 7.17 ;
        RECT  2.82 6.7825 3.5375 6.8525 ;
        RECT  6.645 6.1975 6.78 6.2675 ;
        RECT  1.4675 5.69 1.6025 5.76 ;
        RECT  5.55 5.8325 5.685 5.9025 ;
        RECT  3.9425 5.83 4.0775 5.9 ;
        RECT  2.545 5.83 2.68 5.9 ;
        RECT  1.3275 6.395 1.4625 6.465 ;
        RECT  0.9425 6.0425 1.0825 6.1125 ;
        RECT  4.405 5.69 4.54 5.76 ;
        RECT  3.21 6.195 3.345 6.265 ;
        RECT  6.9025 5.83 7.0375 5.9 ;
        RECT  6.3925 6.0075 6.5275 6.0775 ;
        RECT  5.98 5.69 6.115 5.76 ;
        RECT  1.2775 5.69 1.4125 5.76 ;
        RECT  3.02 5.69 3.155 5.76 ;
        RECT  2.82 6.195 2.955 6.265 ;
        RECT  2.82 6.0075 2.955 6.0775 ;
        RECT  3.4325 6.0075 3.5675 6.0775 ;
        RECT  5.78 6.1975 5.915 6.2675 ;
        RECT  5.78 6.0075 5.915 6.0775 ;
        RECT  7.1125 5.9 7.1825 6.0425 ;
        RECT  0.9425 6.0425 1.0875 6.1125 ;
        RECT  1.0175 5.9 1.0875 6.0475 ;
        RECT  7.1125 6.0425 7.3825 6.1125 ;
        RECT  6.905 6.4 6.965 6.4625 ;
        RECT  0.9425 6.395 7.3825 6.465 ;
        RECT  7.3175 6.045 7.3775 6.11 ;
        RECT  6.9025 5.83 7.1825 5.9 ;
        RECT  1.0175 5.83 2.68 5.9 ;
        RECT  6.695 6.1975 7.3825 6.2675 ;
        RECT  4.0775 5.83 5.685 5.9 ;
        RECT  5.78 6.0075 6.4975 6.0775 ;
        RECT  2.82 6.195 3.345 6.265 ;
        RECT  7.245 6.2 7.305 6.2625 ;
        RECT  5.78 6.1975 6.72 6.2675 ;
        RECT  0.9475 6.045 1.0125 6.1125 ;
        RECT  0.9425 5.69 7.3825 5.76 ;
        RECT  2.82 6.0075 3.5375 6.0775 ;
        RECT  6.645 5.1825 6.78 5.2525 ;
        RECT  1.4675 5.69 1.6025 5.76 ;
        RECT  5.55 5.5475 5.685 5.6175 ;
        RECT  3.9425 5.55 4.0775 5.62 ;
        RECT  2.545 5.55 2.68 5.62 ;
        RECT  1.3275 4.985 1.4625 5.055 ;
        RECT  0.9425 5.3375 1.0825 5.4075 ;
        RECT  4.405 5.69 4.54 5.76 ;
        RECT  3.21 5.185 3.345 5.255 ;
        RECT  6.9025 5.55 7.0375 5.62 ;
        RECT  6.3925 5.3725 6.5275 5.4425 ;
        RECT  5.98 5.69 6.115 5.76 ;
        RECT  1.2775 5.69 1.4125 5.76 ;
        RECT  3.02 5.69 3.155 5.76 ;
        RECT  2.82 5.185 2.955 5.255 ;
        RECT  2.82 5.3725 2.955 5.4425 ;
        RECT  3.4325 5.3725 3.5675 5.4425 ;
        RECT  5.78 5.1825 5.915 5.2525 ;
        RECT  5.78 5.3725 5.915 5.4425 ;
        RECT  7.1125 5.4075 7.1825 5.55 ;
        RECT  0.9425 5.3375 1.0875 5.4075 ;
        RECT  1.0175 5.4025 1.0875 5.55 ;
        RECT  7.1125 5.3375 7.3825 5.4075 ;
        RECT  6.905 4.9875 6.965 5.05 ;
        RECT  0.9425 4.985 7.3825 5.055 ;
        RECT  7.3175 5.34 7.3775 5.405 ;
        RECT  6.9025 5.55 7.1825 5.62 ;
        RECT  1.0175 5.55 2.68 5.62 ;
        RECT  6.695 5.1825 7.3825 5.2525 ;
        RECT  4.0775 5.55 5.685 5.62 ;
        RECT  5.78 5.3725 6.4975 5.4425 ;
        RECT  2.82 5.185 3.345 5.255 ;
        RECT  7.245 5.1875 7.305 5.25 ;
        RECT  5.78 5.1825 6.72 5.2525 ;
        RECT  0.9475 5.3375 1.0125 5.405 ;
        RECT  0.9425 5.69 7.3825 5.76 ;
        RECT  2.82 5.3725 3.5375 5.4425 ;
        RECT  11.27 0.2775 11.34 0.4125 ;
        RECT  11.975 0.2775 12.045 0.4125 ;
        RECT  11.48 0.0 11.55 0.135 ;
        RECT  12.185 0.0 12.255 0.135 ;
        RECT  8.5725 8.73 8.6425 8.865 ;
        RECT  8.5725 7.4525 8.6425 7.5875 ;
        RECT  7.1125 7.4525 7.2475 7.5225 ;
        RECT  8.3625 10.165 8.4325 10.3 ;
        RECT  8.3625 6.7475 8.4325 6.8825 ;
        RECT  7.1125 6.7475 7.2475 6.8175 ;
        RECT  8.1525 14.11 8.2225 14.245 ;
        RECT  8.1525 6.0425 8.2225 6.1775 ;
        RECT  7.1125 6.0425 7.2475 6.1125 ;
        RECT  7.9425 15.545 8.0125 15.68 ;
        RECT  7.9425 5.3375 8.0125 5.4725 ;
        RECT  7.1125 5.3375 7.2475 5.4075 ;
        RECT  10.3925 3.6 10.4625 3.735 ;
        RECT  9.9725 1.415 10.0425 1.55 ;
        RECT  10.1825 2.9625 10.2525 3.0975 ;
        RECT  10.3925 41.1 10.4625 41.235 ;
        RECT  10.6025 10.1025 10.6725 10.2375 ;
        RECT  10.8125 14.1275 10.8825 14.2625 ;
        RECT  1.0125 7.6275 1.1475 7.6975 ;
        RECT  1.0125 7.6275 1.1475 7.6975 ;
        RECT  9.7625 7.98 9.8325 8.115 ;
        RECT  9.7625 41.53 9.8325 41.665 ;
        RECT  8.9225 40.545 9.1275 40.68 ;
        RECT  11.8025 40.545 11.9375 40.615 ;
        RECT  12.5075 40.545 12.6425 40.615 ;
        RECT  11.0275 40.545 11.1625 40.615 ;
        RECT  9.4175 0.355 9.6225 0.49 ;
        RECT  11.8325 0.355 11.9025 0.49 ;
        RECT  11.8325 0.355 11.9025 0.49 ;
        RECT  7.7875 21.5525 7.9225 21.6225 ;
        RECT  7.7875 24.2425 7.9225 24.3125 ;
        RECT  7.7875 26.9325 7.9225 27.0025 ;
        RECT  7.7875 29.6225 7.9225 29.6925 ;
        RECT  7.7875 32.3125 7.9225 32.3825 ;
        RECT  7.7875 35.0025 7.9225 35.0725 ;
        RECT  7.7875 37.6925 7.9225 37.7625 ;
        RECT  7.7875 40.3825 7.9225 40.4525 ;
        RECT  8.9225 13.4125 9.1275 13.5475 ;
        RECT  8.9225 18.7925 9.1275 18.9275 ;
        RECT  7.3125 7.8075 7.4475 7.8775 ;
        RECT  8.9225 7.8075 9.1275 7.9425 ;
        RECT  7.3125 6.3975 7.4475 6.4675 ;
        RECT  8.9225 6.3975 9.1275 6.5325 ;
        RECT  7.3125 6.3975 7.4475 6.4675 ;
        RECT  8.9225 6.3975 9.1275 6.5325 ;
        RECT  7.3125 4.9875 7.4475 5.0575 ;
        RECT  8.9225 4.9875 9.1275 5.1225 ;
        RECT  -5.73 14.925 -0.35 14.995 ;
        RECT  -5.73 15.135 -0.35 15.205 ;
        RECT  -5.73 15.345 -0.35 15.415 ;
        RECT  -5.73 15.555 -0.35 15.625 ;
        RECT  -5.73 15.765 -0.35 15.835 ;
        RECT  -5.73 15.975 -0.35 16.045 ;
        RECT  -5.73 19.225 -0.35 19.295 ;
        RECT  -5.73 19.435 -0.35 19.505 ;
        RECT  -5.73 19.645 -0.35 19.715 ;
        RECT  -5.73 19.855 -0.35 19.925 ;
        RECT  -0.965 9.85 -0.1875 9.92 ;
        RECT  -0.35 15.135 -0.1875 15.205 ;
        RECT  -0.35 19.435 -0.1725 19.505 ;
        RECT  -5.765 14.715 -5.695 14.995 ;
        RECT  -4.355 14.715 -4.285 14.995 ;
        RECT  -4.355 14.715 -4.285 14.995 ;
        RECT  -2.0525 13.41 -0.9325 13.48 ;
        RECT  -0.35 15.975 -0.14 16.045 ;
        RECT  -0.8675 8.415 -0.14 8.485 ;
        RECT  -1.0125 16.865 -0.14 16.935 ;
        RECT  -0.35 19.225 -0.14 19.295 ;
        RECT  -0.965 17.335 -0.14 17.405 ;
        RECT  -5.5675 13.9775 -5.4975 14.1125 ;
        RECT  -5.06 8.8 -4.99 8.935 ;
        RECT  -5.2025 12.8825 -5.1325 13.0175 ;
        RECT  -5.2 11.275 -5.13 11.41 ;
        RECT  -5.2 9.8775 -5.13 10.0125 ;
        RECT  -5.765 8.66 -5.695 8.795 ;
        RECT  -5.4125 8.275 -5.3425 8.415 ;
        RECT  -5.06 11.7375 -4.99 11.8725 ;
        RECT  -5.565 10.5425 -5.495 10.6775 ;
        RECT  -5.2 14.235 -5.13 14.37 ;
        RECT  -5.3775 13.725 -5.3075 13.86 ;
        RECT  -5.06 13.3125 -4.99 13.4475 ;
        RECT  -5.06 8.61 -4.99 8.745 ;
        RECT  -5.06 10.3525 -4.99 10.4875 ;
        RECT  -5.565 10.1525 -5.495 10.2875 ;
        RECT  -5.3775 10.1525 -5.3075 10.2875 ;
        RECT  -5.3775 10.765 -5.3075 10.9 ;
        RECT  -5.5675 13.1125 -5.4975 13.2475 ;
        RECT  -5.3775 13.1125 -5.3075 13.2475 ;
        RECT  -5.3425 14.445 -5.2 14.515 ;
        RECT  -5.4125 8.275 -5.3425 8.42 ;
        RECT  -5.3475 8.35 -5.2 8.42 ;
        RECT  -5.4125 14.445 -5.3425 14.715 ;
        RECT  -5.7625 14.2375 -5.7 14.2975 ;
        RECT  -5.765 8.275 -5.695 14.715 ;
        RECT  -5.41 14.65 -5.345 14.71 ;
        RECT  -5.2 14.235 -5.13 14.515 ;
        RECT  -5.2 8.35 -5.13 10.0125 ;
        RECT  -5.5675 14.0275 -5.4975 14.715 ;
        RECT  -5.2 11.41 -5.13 13.0175 ;
        RECT  -5.3775 13.1125 -5.3075 13.83 ;
        RECT  -5.565 10.1525 -5.495 10.6775 ;
        RECT  -5.5625 14.5775 -5.5 14.6375 ;
        RECT  -5.5675 13.1125 -5.4975 14.0525 ;
        RECT  -5.4125 8.28 -5.345 8.345 ;
        RECT  -5.06 8.275 -4.99 14.715 ;
        RECT  -5.3775 10.1525 -5.3075 10.87 ;
        RECT  -4.5525 13.9775 -4.4825 14.1125 ;
        RECT  -5.06 8.8 -4.99 8.935 ;
        RECT  -4.9175 12.8825 -4.8475 13.0175 ;
        RECT  -4.92 11.275 -4.85 11.41 ;
        RECT  -4.92 9.8775 -4.85 10.0125 ;
        RECT  -4.355 8.66 -4.285 8.795 ;
        RECT  -4.7075 8.275 -4.6375 8.415 ;
        RECT  -5.06 11.7375 -4.99 11.8725 ;
        RECT  -4.555 10.5425 -4.485 10.6775 ;
        RECT  -4.92 14.235 -4.85 14.37 ;
        RECT  -4.7425 13.725 -4.6725 13.86 ;
        RECT  -5.06 13.3125 -4.99 13.4475 ;
        RECT  -5.06 8.61 -4.99 8.745 ;
        RECT  -5.06 10.3525 -4.99 10.4875 ;
        RECT  -4.555 10.1525 -4.485 10.2875 ;
        RECT  -4.7425 10.1525 -4.6725 10.2875 ;
        RECT  -4.7425 10.765 -4.6725 10.9 ;
        RECT  -4.5525 13.1125 -4.4825 13.2475 ;
        RECT  -4.7425 13.1125 -4.6725 13.2475 ;
        RECT  -4.85 14.445 -4.7075 14.515 ;
        RECT  -4.7075 8.275 -4.6375 8.42 ;
        RECT  -4.85 8.35 -4.7025 8.42 ;
        RECT  -4.7075 14.445 -4.6375 14.715 ;
        RECT  -4.35 14.2375 -4.2875 14.2975 ;
        RECT  -4.355 8.275 -4.285 14.715 ;
        RECT  -4.705 14.65 -4.64 14.71 ;
        RECT  -4.92 14.235 -4.85 14.515 ;
        RECT  -4.92 8.35 -4.85 10.0125 ;
        RECT  -4.5525 14.0275 -4.4825 14.715 ;
        RECT  -4.92 11.41 -4.85 13.0175 ;
        RECT  -4.7425 13.1125 -4.6725 13.83 ;
        RECT  -4.555 10.1525 -4.485 10.6775 ;
        RECT  -4.55 14.5775 -4.4875 14.6375 ;
        RECT  -4.5525 13.1125 -4.4825 14.0525 ;
        RECT  -4.705 8.28 -4.6375 8.345 ;
        RECT  -5.06 8.275 -4.99 14.715 ;
        RECT  -4.7425 10.1525 -4.6725 10.87 ;
        RECT  -4.1575 13.9775 -4.0875 14.1125 ;
        RECT  -3.65 8.8 -3.58 8.935 ;
        RECT  -3.7925 12.8825 -3.7225 13.0175 ;
        RECT  -3.79 11.275 -3.72 11.41 ;
        RECT  -3.79 9.8775 -3.72 10.0125 ;
        RECT  -4.355 8.66 -4.285 8.795 ;
        RECT  -4.0025 8.275 -3.9325 8.415 ;
        RECT  -3.65 11.7375 -3.58 11.8725 ;
        RECT  -4.155 10.5425 -4.085 10.6775 ;
        RECT  -3.79 14.235 -3.72 14.37 ;
        RECT  -3.9675 13.725 -3.8975 13.86 ;
        RECT  -3.65 13.3125 -3.58 13.4475 ;
        RECT  -3.65 8.61 -3.58 8.745 ;
        RECT  -3.65 10.3525 -3.58 10.4875 ;
        RECT  -4.155 10.1525 -4.085 10.2875 ;
        RECT  -3.9675 10.1525 -3.8975 10.2875 ;
        RECT  -3.9675 10.765 -3.8975 10.9 ;
        RECT  -4.1575 13.1125 -4.0875 13.2475 ;
        RECT  -3.9675 13.1125 -3.8975 13.2475 ;
        RECT  -3.9325 14.445 -3.79 14.515 ;
        RECT  -4.0025 8.275 -3.9325 8.42 ;
        RECT  -3.9375 8.35 -3.79 8.42 ;
        RECT  -4.0025 14.445 -3.9325 14.715 ;
        RECT  -4.3525 14.2375 -4.29 14.2975 ;
        RECT  -4.355 8.275 -4.285 14.715 ;
        RECT  -4.0 14.65 -3.935 14.71 ;
        RECT  -3.79 14.235 -3.72 14.515 ;
        RECT  -3.79 8.35 -3.72 10.0125 ;
        RECT  -4.1575 14.0275 -4.0875 14.715 ;
        RECT  -3.79 11.41 -3.72 13.0175 ;
        RECT  -3.9675 13.1125 -3.8975 13.83 ;
        RECT  -4.155 10.1525 -4.085 10.6775 ;
        RECT  -4.1525 14.5775 -4.09 14.6375 ;
        RECT  -4.1575 13.1125 -4.0875 14.0525 ;
        RECT  -4.0025 8.28 -3.935 8.345 ;
        RECT  -3.65 8.275 -3.58 14.715 ;
        RECT  -3.9675 10.1525 -3.8975 10.87 ;
        RECT  -1.4125 8.84 -0.835 8.91 ;
        RECT  -1.4125 8.84 -1.2775 8.91 ;
        RECT  -0.8 8.8075 -0.73 8.9425 ;
        RECT  -1.98 21.28 -1.91 21.415 ;
        RECT  -2.105 21.1375 -1.35 21.2075 ;
        RECT  -4.415 21.2 -4.345 22.775 ;
        RECT  -0.6525 21.5675 -0.5825 23.545 ;
        RECT  -2.56 23.545 -2.49 24.2025 ;
        RECT  -0.6525 20.695 -0.5825 20.765 ;
        RECT  -4.03 20.695 -3.96 20.765 ;
        RECT  -0.6525 20.73 -0.5825 21.5675 ;
        RECT  -2.105 20.695 -0.6175 20.765 ;
        RECT  -3.995 20.695 -2.105 20.765 ;
        RECT  -4.03 20.73 -3.96 22.635 ;
        RECT  -3.74 22.075 -3.67 26.2675 ;
        RECT  -3.74 23.835 -3.67 26.2675 ;
        RECT  -0.42 20.73 -0.35 25.225 ;
        RECT  -3.11 23.965 -3.04 25.225 ;
        RECT  -3.53 22.915 -3.46 23.9975 ;
        RECT  -3.74 24.12 -3.67 26.2675 ;
        RECT  -3.53 23.9975 -3.46 25.325 ;
        RECT  -3.74 21.43 -3.67 26.2675 ;
        RECT  -4.935 20.73 -4.865 25.465 ;
        RECT  -4.23 20.73 -4.16 25.465 ;
        RECT  -1.005 23.405 -0.935 23.6425 ;
        RECT  -1.005 22.88 -0.935 23.0825 ;
        RECT  -2.525 22.845 -2.455 22.88 ;
        RECT  -2.525 23.1675 -2.455 23.405 ;
        RECT  -1.005 23.83 -0.935 23.965 ;
        RECT  -1.005 23.27 -0.935 23.405 ;
        RECT  -2.525 22.845 -2.455 22.98 ;
        RECT  -2.525 23.405 -2.455 23.54 ;
        RECT  -1.005 23.5075 -0.935 23.6425 ;
        RECT  -1.005 22.9475 -0.935 23.0825 ;
        RECT  -1.005 22.8125 -0.935 22.9475 ;
        RECT  -2.525 22.8125 -2.455 22.9475 ;
        RECT  -2.525 23.1675 -2.455 23.3025 ;
        RECT  -4.23 23.0375 -4.16 23.1725 ;
        RECT  -4.935 23.5125 -4.865 23.6475 ;
        RECT  -4.23 23.5125 -4.16 23.6475 ;
        RECT  -4.6825 23.0325 -4.6125 23.1675 ;
        RECT  -4.4825 23.0375 -4.4125 23.1725 ;
        RECT  -4.9675 22.74 -4.8325 22.81 ;
        RECT  -4.2625 22.74 -4.1275 22.81 ;
        RECT  -4.75 22.7425 -4.68 22.8075 ;
        RECT  -4.415 22.7425 -4.345 22.8075 ;
        RECT  -4.23 22.74 -4.16 22.81 ;
        RECT  -4.415 22.675 -4.345 24.2325 ;
        RECT  -4.75 22.675 -4.68 24.24 ;
        RECT  -4.935 22.675 -4.865 24.2425 ;
        RECT  -4.23 22.675 -4.16 24.22 ;
        RECT  -4.935 21.89 -4.865 22.025 ;
        RECT  -4.935 21.89 -4.865 22.025 ;
        RECT  -4.935 21.89 -4.865 22.025 ;
        RECT  -4.935 21.89 -4.865 22.025 ;
        RECT  -4.935 21.89 -4.865 22.025 ;
        RECT  -4.935 21.89 -4.865 22.025 ;
        RECT  -4.2625 22.74 -4.1275 22.81 ;
        RECT  -4.9675 22.74 -4.8325 22.81 ;
        RECT  -4.935 21.89 -4.865 22.025 ;
        RECT  -4.935 21.89 -4.865 22.025 ;
        RECT  -4.935 21.89 -4.865 22.025 ;
        RECT  -4.935 21.89 -4.865 22.025 ;
        RECT  -4.935 21.89 -4.865 22.025 ;
        RECT  -4.935 21.89 -4.865 22.025 ;
        RECT  -4.935 21.89 -4.865 22.025 ;
        RECT  -4.935 21.89 -4.865 22.025 ;
        RECT  -4.485 22.3825 -4.415 22.5175 ;
        RECT  -4.23 21.89 -4.16 22.025 ;
        RECT  -4.23 21.89 -4.16 22.025 ;
        RECT  -4.23 21.89 -4.16 22.025 ;
        RECT  -4.23 21.89 -4.16 22.025 ;
        RECT  -4.23 21.89 -4.16 22.025 ;
        RECT  -4.23 21.89 -4.16 22.025 ;
        RECT  -4.935 21.89 -4.865 22.025 ;
        RECT  -4.935 21.89 -4.865 22.025 ;
        RECT  -4.935 21.89 -4.865 22.025 ;
        RECT  -4.935 21.89 -4.865 22.025 ;
        RECT  -4.68 22.3825 -4.61 22.5175 ;
        RECT  -4.9675 22.74 -4.8325 22.81 ;
        RECT  -4.9675 22.74 -4.8325 22.81 ;
        RECT  -4.9675 22.74 -4.8325 22.81 ;
        RECT  -4.935 21.89 -4.865 22.025 ;
        RECT  -4.935 21.89 -4.865 22.025 ;
        RECT  -4.935 21.89 -4.865 22.025 ;
        RECT  -4.935 21.89 -4.865 22.025 ;
        RECT  -4.935 21.89 -4.865 22.025 ;
        RECT  -4.935 21.89 -4.865 22.025 ;
        RECT  -4.2625 22.74 -4.1275 22.81 ;
        RECT  -4.935 21.3975 -4.865 22.8075 ;
        RECT  -4.225 22.7475 -4.165 22.805 ;
        RECT  -4.4075 22.7475 -4.3525 22.8 ;
        RECT  -4.745 22.7475 -4.6875 22.8075 ;
        RECT  -4.93 22.7425 -4.87 22.8 ;
        RECT  -4.75 21.33 -4.68 22.875 ;
        RECT  -4.415 21.33 -4.345 22.875 ;
        RECT  -4.23 21.33 -4.16 22.875 ;
        RECT  -4.935 21.33 -4.865 22.875 ;
        RECT  -4.935 20.835 -4.865 20.97 ;
        RECT  -4.935 20.835 -4.865 20.97 ;
        RECT  -4.935 20.835 -4.865 20.97 ;
        RECT  -4.935 20.835 -4.865 20.97 ;
        RECT  -4.935 20.835 -4.865 20.97 ;
        RECT  -4.935 20.835 -4.865 20.97 ;
        RECT  -4.2625 20.05 -4.1275 20.12 ;
        RECT  -4.9675 20.05 -4.8325 20.12 ;
        RECT  -4.935 20.835 -4.865 20.97 ;
        RECT  -4.935 20.835 -4.865 20.97 ;
        RECT  -4.935 20.835 -4.865 20.97 ;
        RECT  -4.935 20.835 -4.865 20.97 ;
        RECT  -4.935 20.835 -4.865 20.97 ;
        RECT  -4.935 20.835 -4.865 20.97 ;
        RECT  -4.935 20.835 -4.865 20.97 ;
        RECT  -4.935 20.835 -4.865 20.97 ;
        RECT  -4.485 20.3425 -4.415 20.4775 ;
        RECT  -4.23 20.835 -4.16 20.97 ;
        RECT  -4.23 20.835 -4.16 20.97 ;
        RECT  -4.23 20.835 -4.16 20.97 ;
        RECT  -4.23 20.835 -4.16 20.97 ;
        RECT  -4.23 20.835 -4.16 20.97 ;
        RECT  -4.23 20.835 -4.16 20.97 ;
        RECT  -4.935 20.835 -4.865 20.97 ;
        RECT  -4.935 20.835 -4.865 20.97 ;
        RECT  -4.935 20.835 -4.865 20.97 ;
        RECT  -4.935 20.835 -4.865 20.97 ;
        RECT  -4.68 20.3425 -4.61 20.4775 ;
        RECT  -4.9675 20.05 -4.8325 20.12 ;
        RECT  -4.9675 20.05 -4.8325 20.12 ;
        RECT  -4.9675 20.05 -4.8325 20.12 ;
        RECT  -4.935 20.835 -4.865 20.97 ;
        RECT  -4.935 20.835 -4.865 20.97 ;
        RECT  -4.935 20.835 -4.865 20.97 ;
        RECT  -4.935 20.835 -4.865 20.97 ;
        RECT  -4.935 20.835 -4.865 20.97 ;
        RECT  -4.935 20.835 -4.865 20.97 ;
        RECT  -4.2625 20.05 -4.1275 20.12 ;
        RECT  -4.935 20.0525 -4.865 21.4625 ;
        RECT  -4.225 20.055 -4.165 20.1125 ;
        RECT  -4.4075 20.06 -4.3525 20.1125 ;
        RECT  -4.745 20.0525 -4.6875 20.1125 ;
        RECT  -4.93 20.06 -4.87 20.1175 ;
        RECT  -4.75 19.985 -4.68 21.53 ;
        RECT  -4.415 19.985 -4.345 21.53 ;
        RECT  -4.23 19.985 -4.16 21.53 ;
        RECT  -4.935 19.985 -4.865 21.53 ;
        RECT  -1.98 21.1775 -1.91 21.3125 ;
        RECT  -1.4175 21.0675 -1.2825 21.1375 ;
        RECT  -2.1725 21.0675 -2.0375 21.1375 ;
        RECT  -4.4475 21.095 -4.3125 21.165 ;
        RECT  -0.685 23.44 -0.55 23.51 ;
        RECT  -2.5925 23.44 -2.4575 23.51 ;
        RECT  -2.595 24.2025 -2.525 24.3375 ;
        RECT  -0.6525 21.365 -0.5825 21.5 ;
        RECT  -4.03 22.4325 -3.96 22.5675 ;
        RECT  -3.7725 21.97 -3.6375 22.04 ;
        RECT  -3.7725 23.73 -3.6375 23.8 ;
        RECT  -0.4525 20.625 -0.3175 20.695 ;
        RECT  -0.4525 25.12 -0.3175 25.19 ;
        RECT  -3.1425 25.12 -3.0075 25.19 ;
        RECT  -3.775 26.2675 -3.705 26.4025 ;
        RECT  -3.5625 23.8925 -3.4275 23.9625 ;
        RECT  -3.5625 22.81 -3.4275 22.88 ;
        RECT  -3.7725 24.015 -3.6375 24.085 ;
        RECT  -3.5625 23.8925 -3.4275 23.9625 ;
        RECT  -3.5625 25.22 -3.4275 25.29 ;
        RECT  -3.7725 21.325 -3.6375 21.395 ;
        RECT  -4.9675 20.625 -4.8325 20.695 ;
        RECT  -4.2625 20.625 -4.1275 20.695 ;
        RECT  -1.9775 16.605 -1.9075 17.055 ;
        RECT  -2.6475 16.255 -2.5775 16.73 ;
        RECT  -2.7875 16.255 -2.7175 16.92 ;
        RECT  -2.7175 16.85 -2.5775 16.92 ;
        RECT  -2.1125 16.605 -1.9775 16.675 ;
        RECT  -2.1125 16.985 -1.9775 17.055 ;
        RECT  -2.7125 16.66 -2.5775 16.73 ;
        RECT  -2.7175 16.215 -2.6475 16.35 ;
        RECT  -2.7125 16.85 -2.5775 16.92 ;
        RECT  -2.8575 16.215 -2.7875 16.35 ;
        RECT  -4.1725 16.605 -4.1025 17.055 ;
        RECT  -3.5025 16.255 -3.4325 16.73 ;
        RECT  -3.3625 16.255 -3.2925 16.92 ;
        RECT  -3.5025 16.85 -3.3625 16.92 ;
        RECT  -4.2375 16.605 -4.1025 16.675 ;
        RECT  -4.2375 16.985 -4.1025 17.055 ;
        RECT  -3.6375 16.66 -3.5025 16.73 ;
        RECT  -3.5025 16.215 -3.4325 16.35 ;
        RECT  -3.6375 16.85 -3.5025 16.92 ;
        RECT  -3.3625 16.215 -3.2925 16.35 ;
        RECT  -4.0 14.615 -3.93 14.75 ;
        RECT  -4.0 15.105 -3.93 15.24 ;
        RECT  -4.155 14.615 -4.085 14.75 ;
        RECT  -4.155 15.315 -4.085 15.45 ;
        RECT  -5.565 14.615 -5.495 14.75 ;
        RECT  -5.565 15.525 -5.495 15.66 ;
        RECT  -4.55 14.615 -4.48 14.75 ;
        RECT  -4.55 15.735 -4.48 15.87 ;
        RECT  -1.3275 15.315 -1.2575 15.45 ;
        RECT  -0.7975 15.945 -0.7275 16.08 ;
        RECT  -2.1225 15.945 -2.0525 16.08 ;
        RECT  -2.645 15.315 -2.575 15.45 ;
        RECT  -2.785 15.525 -2.715 15.66 ;
        RECT  -4.0275 15.945 -3.9575 16.08 ;
        RECT  -3.505 15.735 -3.435 15.87 ;
        RECT  -3.365 15.525 -3.295 15.66 ;
        RECT  -1.0 9.8175 -0.93 9.9525 ;
        RECT  -0.2225 9.8175 -0.1525 9.9525 ;
        RECT  -0.2225 15.1025 -0.1525 15.2375 ;
        RECT  -2.4925 19.405 -2.4225 19.54 ;
        RECT  -3.6575 19.195 -3.5875 19.33 ;
        RECT  -0.9675 19.615 -0.8975 19.75 ;
        RECT  -0.2075 19.4025 -0.1375 19.5375 ;
        RECT  -2.045 19.645 -1.91 19.715 ;
        RECT  -2.045 21.28 -1.91 21.35 ;
        RECT  -1.73 19.825 -1.66 19.96 ;
        RECT  -4.42 19.825 -4.35 19.96 ;
        RECT  -0.385 14.895 -0.315 15.03 ;
        RECT  -0.9675 13.3775 -0.8975 13.5125 ;
        RECT  -2.0875 13.3775 -2.0175 13.5125 ;
        RECT  -2.085 8.275 -2.015 8.41 ;
        RECT  -2.085 8.275 -2.015 8.41 ;
        RECT  -0.275 15.975 -0.14 16.045 ;
        RECT  -0.8675 8.415 -0.7975 8.55 ;
        RECT  -0.275 8.415 -0.14 8.485 ;
        RECT  -1.0825 16.865 -0.9475 16.935 ;
        RECT  -0.275 16.865 -0.14 16.935 ;
        RECT  -0.275 19.225 -0.14 19.295 ;
        RECT  -1.035 17.335 -0.9 17.405 ;
        RECT  -0.275 17.335 -0.14 17.405 ;
        RECT  9.6975 8.275 9.8325 8.345 ;
        RECT  10.3275 15.975 10.4625 16.045 ;
        RECT  10.1175 8.415 10.2525 8.485 ;
        RECT  9.9075 16.865 10.0425 16.935 ;
        RECT  10.5375 19.225 10.6725 19.295 ;
        RECT  10.7475 17.335 10.8825 17.405 ;
        RECT  0.0325 19.855 0.2375 19.99 ;
        RECT  8.9225 20.695 9.1275 20.83 ;
        RECT  -0.415 20.695 -0.28 20.765 ;
        LAYER  via2 ;
        RECT  11.475 18.79 11.545 18.86 ;
        RECT  12.18 18.79 12.25 18.86 ;
        RECT  11.48 9.87 11.55 9.94 ;
        RECT  12.185 9.87 12.255 9.94 ;
        RECT  11.48 3.43 11.55 3.5 ;
        RECT  12.185 3.43 12.255 3.5 ;
        RECT  11.48 3.5825 11.55 3.6525 ;
        RECT  12.185 3.5825 12.255 3.6525 ;
        RECT  0.9775 7.4525 1.0475 7.5225 ;
        RECT  0.9775 6.7475 1.0475 6.8175 ;
        RECT  0.9775 6.0425 1.0475 6.1125 ;
        RECT  0.9775 5.3375 1.0475 5.4075 ;
        RECT  11.2725 0.3125 11.3375 0.3775 ;
        RECT  11.9775 0.3125 12.0425 0.3775 ;
        RECT  11.4825 0.035 11.5475 0.1 ;
        RECT  12.1875 0.035 12.2525 0.1 ;
        RECT  8.575 7.4875 8.64 7.5525 ;
        RECT  7.1475 7.455 7.2125 7.52 ;
        RECT  8.365 6.7825 8.43 6.8475 ;
        RECT  7.1475 6.75 7.2125 6.815 ;
        RECT  8.155 6.0775 8.22 6.1425 ;
        RECT  7.1475 6.045 7.2125 6.11 ;
        RECT  7.945 5.3725 8.01 5.4375 ;
        RECT  7.1475 5.34 7.2125 5.405 ;
        RECT  1.0475 7.63 1.1125 7.695 ;
        RECT  9.765 8.015 9.83 8.08 ;
        RECT  -5.4125 8.31 -5.3425 8.38 ;
        RECT  -4.7075 8.31 -4.6375 8.38 ;
        RECT  -4.0025 8.31 -3.9325 8.38 ;
        RECT  -1.0025 22.8475 -0.9375 22.9125 ;
        RECT  -2.5225 22.8475 -2.4575 22.9125 ;
        RECT  -2.01 19.6475 -1.945 19.7125 ;
        RECT  -2.01 21.2825 -1.945 21.3475 ;
        RECT  -2.0825 8.31 -2.0175 8.375 ;
        RECT  -0.24 15.9775 -0.175 16.0425 ;
        RECT  -0.24 8.4175 -0.175 8.4825 ;
        RECT  -0.24 16.8675 -0.175 16.9325 ;
        RECT  -0.24 19.2275 -0.175 19.2925 ;
        RECT  -0.24 17.3375 -0.175 17.4025 ;
        RECT  9.7325 8.2775 9.7975 8.3425 ;
        RECT  10.3625 15.9775 10.4275 16.0425 ;
        RECT  10.1525 8.4175 10.2175 8.4825 ;
        RECT  9.9425 16.8675 10.0075 16.9325 ;
        RECT  10.5725 19.2275 10.6375 19.2925 ;
        RECT  10.7825 17.3375 10.8475 17.4025 ;
        RECT  8.9225 20.73 8.9875 20.795 ;
        RECT  9.0625 20.73 9.1275 20.795 ;
        RECT  -0.38 20.6975 -0.315 20.7625 ;
        LAYER  metal3 ;
        RECT  -2.0525 8.275 9.7625 8.345 ;
        RECT  -0.14 15.975 10.3925 16.045 ;
        RECT  -0.14 8.415 10.1825 8.485 ;
        RECT  -0.14 16.865 9.9725 16.935 ;
        RECT  -0.14 19.225 10.6025 19.295 ;
        RECT  -0.14 17.335 10.8125 17.405 ;
        RECT  -0.28 20.695 8.9225 20.765 ;
        RECT  11.27 18.73 11.34 18.8 ;
        RECT  11.27 0.3125 11.34 18.7675 ;
        RECT  11.305 18.73 11.545 18.8 ;
        RECT  11.975 18.73 12.045 18.8 ;
        RECT  11.975 0.3125 12.045 18.7675 ;
        RECT  12.01 18.73 12.25 18.8 ;
        RECT  11.48 0.0 11.55 3.22 ;
        RECT  12.185 0.0 12.255 3.22 ;
        RECT  7.2475 7.4525 8.6425 7.5225 ;
        RECT  7.2475 6.7475 8.4325 6.8175 ;
        RECT  7.2475 6.0425 8.2225 6.1125 ;
        RECT  7.2475 5.3375 8.0125 5.4075 ;
        RECT  0.0325 7.4525 1.015 7.5225 ;
        RECT  0.0325 6.7475 1.015 6.8175 ;
        RECT  0.0325 6.0425 1.015 6.1125 ;
        RECT  0.0325 5.3375 1.015 5.4075 ;
        RECT  1.1125 7.98 1.1825 8.05 ;
        RECT  1.1125 7.6275 1.1825 8.015 ;
        RECT  1.1475 7.98 9.765 8.05 ;
        RECT  11.475 18.755 11.545 18.895 ;
        RECT  12.18 18.755 12.25 18.895 ;
        RECT  11.48 9.835 11.55 9.975 ;
        RECT  12.185 9.835 12.255 9.975 ;
        RECT  11.48 3.395 11.55 3.535 ;
        RECT  12.185 3.395 12.255 3.535 ;
        RECT  11.48 3.5475 11.55 3.6875 ;
        RECT  12.185 3.5475 12.255 3.6875 ;
        RECT  0.9425 7.4525 1.0825 7.5225 ;
        RECT  0.9425 6.7475 1.0825 6.8175 ;
        RECT  0.9425 6.0425 1.0825 6.1125 ;
        RECT  0.9425 5.3375 1.0825 5.4075 ;
        RECT  11.27 0.2775 11.34 0.4125 ;
        RECT  11.975 0.2775 12.045 0.4125 ;
        RECT  11.48 0.0 11.55 0.135 ;
        RECT  12.185 0.0 12.255 0.135 ;
        RECT  8.5725 7.4525 8.6425 7.5875 ;
        RECT  7.1125 7.4525 7.2475 7.5225 ;
        RECT  8.3625 6.7475 8.4325 6.8825 ;
        RECT  7.1125 6.7475 7.2475 6.8175 ;
        RECT  8.1525 6.0425 8.2225 6.1775 ;
        RECT  7.1125 6.0425 7.2475 6.1125 ;
        RECT  7.9425 5.3375 8.0125 5.4725 ;
        RECT  7.1125 5.3375 7.2475 5.4075 ;
        RECT  1.0125 7.6275 1.1475 7.6975 ;
        RECT  9.7625 7.98 9.8325 8.115 ;
        RECT  -1.98 19.645 -1.91 21.3125 ;
        RECT  -5.4125 8.275 -5.3425 8.415 ;
        RECT  -4.7075 8.275 -4.6375 8.415 ;
        RECT  -4.0025 8.275 -3.9325 8.415 ;
        RECT  -2.49 22.845 -0.97 22.915 ;
        RECT  -1.005 22.8125 -0.935 22.9475 ;
        RECT  -2.525 22.8125 -2.455 22.9475 ;
        RECT  -2.045 19.645 -1.91 19.715 ;
        RECT  -2.045 21.28 -1.91 21.35 ;
        RECT  -2.085 8.275 -2.015 8.41 ;
        RECT  -0.275 15.975 -0.14 16.045 ;
        RECT  -0.275 8.415 -0.14 8.485 ;
        RECT  -0.275 16.865 -0.14 16.935 ;
        RECT  -0.275 19.225 -0.14 19.295 ;
        RECT  -0.275 17.335 -0.14 17.405 ;
        RECT  9.6975 8.275 9.8325 8.345 ;
        RECT  10.3275 15.975 10.4625 16.045 ;
        RECT  10.1175 8.415 10.2525 8.485 ;
        RECT  9.9075 16.865 10.0425 16.935 ;
        RECT  10.5375 19.225 10.6725 19.295 ;
        RECT  10.7475 17.335 10.8825 17.405 ;
        RECT  8.9225 20.695 9.1275 20.83 ;
        RECT  -0.415 20.695 -0.28 20.765 ;
    END
END    sram_2_16_1_freepdk45
END    LIBRARY
