magic
tech sky130A
magscale 1 2
timestamp 1595931502
<< checkpaint >>
rect -1190 -1316 2772 1750
<< locali >>
rect 70 282 136 316
rect 549 314 970 348
rect 70 174 136 208
rect 936 197 970 314
rect 1041 130 1494 164
<< metal1 >>
rect 246 -30 294 402
rect 670 -32 720 402
rect 1060 0 1088 395
rect 1332 0 1360 395
use pinv_dec  pinv_dec_0
timestamp 1595931502
transform 1 0 876 0 1 0
box 44 0 636 490
use nand2_dec  nand2_dec_0
timestamp 1595931502
transform 1 0 0 0 1 0
box 70 -56 888 476
<< labels >>
rlabel metal1 s 270 186 270 186 4 gnd
rlabel metal1 s 1074 197 1074 197 4 gnd
rlabel corelocali s 103 191 103 191 4 B
rlabel corelocali s 1267 147 1267 147 4 Z
rlabel metal1 s 695 185 695 185 4 vdd
rlabel metal1 s 1346 197 1346 197 4 vdd
rlabel corelocali s 103 299 103 299 4 A
<< properties >>
string FIXED_BBOX 0 0 1494 395
<< end >>
