magic
tech sky130A
magscale 1 2
timestamp 1593453062
<< nwell >>
rect -160 524 682 1614
rect -160 264 684 524
<< nmos >>
rect 242 2005 272 2135
rect 154 1689 184 1819
rect 242 1689 272 1819
rect 156 66 186 196
<< pmos >>
rect 154 1324 184 1576
rect 242 1324 272 1576
rect 154 702 184 1102
rect 346 702 376 1102
rect 156 302 186 554
<< ndiff >>
rect 184 2126 242 2135
rect 184 2013 196 2126
rect 230 2013 242 2126
rect 184 2005 242 2013
rect 272 2126 330 2135
rect 272 2017 284 2126
rect 318 2017 330 2126
rect 272 2005 330 2017
rect 96 1811 154 1819
rect 96 1701 108 1811
rect 142 1701 154 1811
rect 96 1689 154 1701
rect 184 1811 242 1819
rect 184 1701 196 1811
rect 230 1701 242 1811
rect 184 1689 242 1701
rect 272 1811 330 1819
rect 272 1701 284 1811
rect 318 1701 330 1811
rect 272 1689 330 1701
rect 98 184 156 196
rect 98 78 110 184
rect 144 78 156 184
rect 98 66 156 78
rect 186 184 242 196
rect 186 78 198 184
rect 232 78 242 184
rect 186 66 242 78
<< pdiff >>
rect 100 1564 154 1576
rect 100 1336 108 1564
rect 142 1336 154 1564
rect 100 1324 154 1336
rect 184 1564 242 1576
rect 184 1336 196 1564
rect 230 1336 242 1564
rect 184 1324 242 1336
rect 272 1564 326 1576
rect 272 1336 284 1564
rect 318 1336 326 1564
rect 272 1324 326 1336
rect 100 1090 154 1102
rect 100 714 108 1090
rect 142 714 154 1090
rect 100 702 154 714
rect 184 1090 238 1102
rect 184 714 196 1090
rect 230 714 238 1090
rect 184 702 238 714
rect 292 1090 346 1102
rect 292 714 300 1090
rect 334 714 346 1090
rect 292 702 346 714
rect 376 1090 430 1102
rect 376 714 388 1090
rect 422 714 430 1090
rect 376 702 430 714
rect 98 542 156 554
rect 98 314 110 542
rect 144 314 156 542
rect 98 302 156 314
rect 186 542 240 554
rect 186 314 198 542
rect 232 314 240 542
rect 186 302 240 314
<< ndiffc >>
rect 196 2013 230 2126
rect 284 2017 318 2126
rect 108 1701 142 1811
rect 196 1701 230 1811
rect 284 1701 318 1811
rect 110 78 144 184
rect 198 78 232 184
<< pdiffc >>
rect 108 1336 142 1564
rect 196 1336 230 1564
rect 284 1336 318 1564
rect 108 714 142 1090
rect 196 714 230 1090
rect 300 714 334 1090
rect 388 714 422 1090
rect 110 314 144 542
rect 198 314 232 542
<< psubdiff >>
rect 434 2085 468 2109
rect 434 2017 468 2051
rect 364 151 398 175
rect 364 83 398 117
<< nsubdiff >>
rect 388 1348 422 1372
rect 388 1290 422 1314
<< psubdiffcont >>
rect 434 2051 468 2085
rect 364 117 398 151
<< nsubdiffcont >>
rect 388 1314 422 1348
<< poly >>
rect 240 2220 274 2226
rect 230 2210 284 2220
rect 230 2176 240 2210
rect 274 2176 284 2210
rect 230 2166 284 2176
rect 240 2160 274 2166
rect 242 2135 272 2160
rect 242 1989 272 2005
rect 26 1959 272 1989
rect 26 1148 56 1959
rect 306 1917 372 1927
rect 154 1887 322 1917
rect 154 1819 184 1887
rect 306 1883 322 1887
rect 356 1883 372 1917
rect 306 1873 372 1883
rect 342 1862 372 1873
rect 242 1819 272 1845
rect 342 1828 376 1862
rect 154 1576 184 1689
rect 242 1576 272 1689
rect 345 1676 375 1828
rect 342 1642 376 1676
rect 154 1298 184 1324
rect 242 1256 272 1324
rect 98 1240 272 1256
rect 98 1206 108 1240
rect 142 1226 272 1240
rect 342 1232 372 1642
rect 142 1206 152 1226
rect 98 1196 152 1206
rect 342 1206 474 1232
rect 342 1202 430 1206
rect 108 1190 142 1196
rect 420 1172 430 1202
rect 464 1172 474 1206
rect 420 1158 474 1172
rect 430 1156 474 1158
rect 26 1118 184 1148
rect 154 1102 184 1118
rect 346 1102 376 1128
rect 154 686 184 702
rect 346 686 376 702
rect 154 656 376 686
rect 156 598 432 614
rect 156 584 388 598
rect 156 554 186 584
rect 378 564 388 584
rect 422 564 432 598
rect 378 548 432 564
rect 156 196 186 302
rect 156 36 186 66
<< polycont >>
rect 240 2176 274 2210
rect 322 1883 356 1917
rect 108 1206 142 1240
rect 430 1172 464 1206
rect 388 564 422 598
<< locali >>
rect 140 2176 240 2210
rect 274 2176 290 2210
rect 196 2126 230 2142
rect 108 1811 142 1830
rect 108 1564 142 1701
rect 196 1811 230 2013
rect 284 2126 318 2142
rect 434 2085 468 2101
rect 318 2051 434 2085
rect 284 2001 318 2017
rect 196 1685 230 1701
rect 284 1883 322 1917
rect 356 1883 374 1917
rect 284 1811 318 1883
rect 108 1240 142 1336
rect 196 1564 230 1580
rect 196 1286 230 1336
rect 284 1564 318 1701
rect 284 1320 318 1336
rect 352 1314 388 1348
rect 422 1314 438 1348
rect 352 1286 386 1314
rect 196 1252 352 1286
rect 108 1090 142 1206
rect 420 1206 474 1222
rect 420 1190 430 1206
rect 388 1172 430 1190
rect 464 1172 474 1206
rect 388 1156 474 1172
rect 108 656 142 714
rect 196 694 230 714
rect 300 1090 334 1096
rect 300 698 334 714
rect 388 1090 422 1156
rect 388 598 422 714
rect 110 542 144 558
rect 110 242 144 314
rect 198 542 232 558
rect 388 548 422 564
rect 232 412 364 446
rect 198 298 232 314
rect 110 184 144 208
rect 110 60 144 78
rect 196 184 232 200
rect 196 78 198 184
rect 364 152 398 167
rect 232 151 398 152
rect 232 116 364 151
rect 196 60 232 78
<< viali >>
rect 106 2176 140 2212
rect 434 2017 468 2051
rect 352 1252 386 1286
rect 196 1090 230 1124
rect 300 1096 334 1130
rect 364 412 398 446
rect 110 208 144 242
rect 364 83 398 117
<< metal1 >>
rect 94 2212 152 2224
rect 94 2176 106 2212
rect 140 2176 152 2212
rect 94 2164 152 2176
rect 196 1130 230 2256
rect 272 1142 300 2256
rect 428 2051 474 2079
rect 428 2017 434 2051
rect 468 2017 474 2051
rect 428 2005 474 2017
rect 338 1286 400 1302
rect 338 1252 352 1286
rect 386 1252 400 1286
rect 338 1234 400 1252
rect 272 1130 340 1142
rect 184 1124 242 1130
rect 184 1090 196 1124
rect 230 1090 242 1124
rect 184 1084 242 1090
rect 272 1096 300 1130
rect 334 1096 340 1130
rect 272 1084 340 1096
rect 104 242 150 254
rect 104 208 110 242
rect 144 208 150 242
rect 104 0 150 208
rect 196 0 230 1084
rect 272 0 300 1084
rect 358 446 404 468
rect 358 412 364 446
rect 398 412 404 446
rect 358 392 404 412
rect 358 117 404 145
rect 358 83 364 117
rect 398 83 404 117
rect 358 71 404 83
<< labels >>
rlabel metal1 394 1268 394 1268 1 vdd
rlabel metal1 450 2011 450 2011 1 gnd
rlabel metal1 214 2248 214 2248 1 bl
rlabel metal1 286 2246 286 2246 1 br
rlabel metal1 122 28 124 28 1 dout
rlabel metal1 380 77 380 77 1 gnd
rlabel metal1 378 400 378 400 1 vdd
rlabel metal1 100 2190 100 2190 1 en
<< properties >>
string FIXED_BBOX 0 0 500 2256
<< end >>
