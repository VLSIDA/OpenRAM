VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 1000 ;
END UNITS
SITE  MacroSite
   CLASS Core ;
   SIZE 24385.0 by 72042.5 ;
END  MacroSite
MACRO sram_2_16_1_freepdk45
   CLASS BLOCK ;
   SIZE 24385.0 BY 72042.5 ;
   SYMMETRY X Y R90 ;
   SITE MacroSite ;
   PIN DATA[0]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  16402.5 35.0 16472.5 175.0 ;
      END
   END DATA[0]
   PIN DATA[1]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  19222.5 35.0 19292.5 175.0 ;
      END
   END DATA[1]
   PIN ADDR[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  4175.0 10372.5 4655.0 10442.5 ;
      END
   END ADDR[0]
   PIN ADDR[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  4175.0 9667.5 4655.0 9737.5 ;
      END
   END ADDR[1]
   PIN ADDR[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  4175.0 8962.5 4655.0 9032.5 ;
      END
   END ADDR[2]
   PIN ADDR[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  4175.0 8257.5 4655.0 8327.5 ;
      END
   END ADDR[3]
   PIN ADDR[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  4175.0 7552.5 4655.0 7622.5 ;
      END
   END ADDR[4]
   PIN ADDR[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  4175.0 6847.5 4655.0 6917.5 ;
      END
   END ADDR[5]
   PIN ADDR[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  4175.0 6142.5 4655.0 6212.5 ;
      END
   END ADDR[6]
   PIN CSb
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1187.5 27450.0 1257.5 27590.0 ;
      END
   END CSb
   PIN WEb
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1892.5 27450.0 1962.5 27590.0 ;
      END
   END WEb
   PIN OEb
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  482.5 27450.0 552.5 27590.0 ;
      END
   END OEb
   PIN clk
      DIRECTION INPUT ;
      PORT
         LAYER metal1 ;
         RECT  3340.0 27450.0 3475.0 27640.0 ;
      END
   END clk
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal1 ;
         RECT  21920.0 35.0 22270.0 72077.5 ;
         LAYER metal1 ;
         RECT  4175.0 35.0 4525.0 72077.5 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal2 ;
         RECT  13992.5 35.0 14342.5 72077.5 ;
      END
   END gnd
   OBS
   LAYER  metal1 ;
      RECT  4317.5 35155.0 4382.5 35360.0 ;
      RECT  8100.0 27905.0 8165.0 27970.0 ;
      RECT  8100.0 27632.5 8165.0 27697.5 ;
      RECT  8030.0 27905.0 8132.5 27970.0 ;
      RECT  8100.0 27665.0 8165.0 27937.5 ;
      RECT  8132.5 27632.5 8235.0 27697.5 ;
      RECT  13227.5 27905.0 13292.5 27970.0 ;
      RECT  13227.5 27417.5 13292.5 27482.5 ;
      RECT  10525.0 27905.0 13260.0 27970.0 ;
      RECT  13227.5 27450.0 13292.5 27937.5 ;
      RECT  13260.0 27417.5 15995.0 27482.5 ;
      RECT  8100.0 29340.0 8165.0 29405.0 ;
      RECT  8100.0 29612.5 8165.0 29677.5 ;
      RECT  8030.0 29340.0 8132.5 29405.0 ;
      RECT  8100.0 29372.5 8165.0 29645.0 ;
      RECT  8132.5 29612.5 8235.0 29677.5 ;
      RECT  13227.5 29340.0 13292.5 29405.0 ;
      RECT  13227.5 29827.5 13292.5 29892.5 ;
      RECT  10525.0 29340.0 13260.0 29405.0 ;
      RECT  13227.5 29372.5 13292.5 29860.0 ;
      RECT  13260.0 29827.5 15995.0 29892.5 ;
      RECT  8100.0 30595.0 8165.0 30660.0 ;
      RECT  8100.0 30322.5 8165.0 30387.5 ;
      RECT  8030.0 30595.0 8132.5 30660.0 ;
      RECT  8100.0 30355.0 8165.0 30627.5 ;
      RECT  8132.5 30322.5 8235.0 30387.5 ;
      RECT  13227.5 30595.0 13292.5 30660.0 ;
      RECT  13227.5 30107.5 13292.5 30172.5 ;
      RECT  10525.0 30595.0 13260.0 30660.0 ;
      RECT  13227.5 30140.0 13292.5 30627.5 ;
      RECT  13260.0 30107.5 15995.0 30172.5 ;
      RECT  8100.0 32030.0 8165.0 32095.0 ;
      RECT  8100.0 32302.5 8165.0 32367.5 ;
      RECT  8030.0 32030.0 8132.5 32095.0 ;
      RECT  8100.0 32062.5 8165.0 32335.0 ;
      RECT  8132.5 32302.5 8235.0 32367.5 ;
      RECT  13227.5 32030.0 13292.5 32095.0 ;
      RECT  13227.5 32517.5 13292.5 32582.5 ;
      RECT  10525.0 32030.0 13260.0 32095.0 ;
      RECT  13227.5 32062.5 13292.5 32550.0 ;
      RECT  13260.0 32517.5 15995.0 32582.5 ;
      RECT  8100.0 33285.0 8165.0 33350.0 ;
      RECT  8100.0 33012.5 8165.0 33077.5 ;
      RECT  8030.0 33285.0 8132.5 33350.0 ;
      RECT  8100.0 33045.0 8165.0 33317.5 ;
      RECT  8132.5 33012.5 8235.0 33077.5 ;
      RECT  13227.5 33285.0 13292.5 33350.0 ;
      RECT  13227.5 32797.5 13292.5 32862.5 ;
      RECT  10525.0 33285.0 13260.0 33350.0 ;
      RECT  13227.5 32830.0 13292.5 33317.5 ;
      RECT  13260.0 32797.5 15995.0 32862.5 ;
      RECT  8100.0 34720.0 8165.0 34785.0 ;
      RECT  8100.0 34992.5 8165.0 35057.5 ;
      RECT  8030.0 34720.0 8132.5 34785.0 ;
      RECT  8100.0 34752.5 8165.0 35025.0 ;
      RECT  8132.5 34992.5 8235.0 35057.5 ;
      RECT  13227.5 34720.0 13292.5 34785.0 ;
      RECT  13227.5 35207.5 13292.5 35272.5 ;
      RECT  10525.0 34720.0 13260.0 34785.0 ;
      RECT  13227.5 34752.5 13292.5 35240.0 ;
      RECT  13260.0 35207.5 15995.0 35272.5 ;
      RECT  8100.0 35975.0 8165.0 36040.0 ;
      RECT  8100.0 35702.5 8165.0 35767.5 ;
      RECT  8030.0 35975.0 8132.5 36040.0 ;
      RECT  8100.0 35735.0 8165.0 36007.5 ;
      RECT  8132.5 35702.5 8235.0 35767.5 ;
      RECT  13227.5 35975.0 13292.5 36040.0 ;
      RECT  13227.5 35487.5 13292.5 35552.5 ;
      RECT  10525.0 35975.0 13260.0 36040.0 ;
      RECT  13227.5 35520.0 13292.5 36007.5 ;
      RECT  13260.0 35487.5 15995.0 35552.5 ;
      RECT  8100.0 37410.0 8165.0 37475.0 ;
      RECT  8100.0 37682.5 8165.0 37747.5 ;
      RECT  8030.0 37410.0 8132.5 37475.0 ;
      RECT  8100.0 37442.5 8165.0 37715.0 ;
      RECT  8132.5 37682.5 8235.0 37747.5 ;
      RECT  13227.5 37410.0 13292.5 37475.0 ;
      RECT  13227.5 37897.5 13292.5 37962.5 ;
      RECT  10525.0 37410.0 13260.0 37475.0 ;
      RECT  13227.5 37442.5 13292.5 37930.0 ;
      RECT  13260.0 37897.5 15995.0 37962.5 ;
      RECT  8100.0 38665.0 8165.0 38730.0 ;
      RECT  8100.0 38392.5 8165.0 38457.5 ;
      RECT  8030.0 38665.0 8132.5 38730.0 ;
      RECT  8100.0 38425.0 8165.0 38697.5 ;
      RECT  8132.5 38392.5 8235.0 38457.5 ;
      RECT  13227.5 38665.0 13292.5 38730.0 ;
      RECT  13227.5 38177.5 13292.5 38242.5 ;
      RECT  10525.0 38665.0 13260.0 38730.0 ;
      RECT  13227.5 38210.0 13292.5 38697.5 ;
      RECT  13260.0 38177.5 15995.0 38242.5 ;
      RECT  8100.0 40100.0 8165.0 40165.0 ;
      RECT  8100.0 40372.5 8165.0 40437.5 ;
      RECT  8030.0 40100.0 8132.5 40165.0 ;
      RECT  8100.0 40132.5 8165.0 40405.0 ;
      RECT  8132.5 40372.5 8235.0 40437.5 ;
      RECT  13227.5 40100.0 13292.5 40165.0 ;
      RECT  13227.5 40587.5 13292.5 40652.5 ;
      RECT  10525.0 40100.0 13260.0 40165.0 ;
      RECT  13227.5 40132.5 13292.5 40620.0 ;
      RECT  13260.0 40587.5 15995.0 40652.5 ;
      RECT  8100.0 41355.0 8165.0 41420.0 ;
      RECT  8100.0 41082.5 8165.0 41147.5 ;
      RECT  8030.0 41355.0 8132.5 41420.0 ;
      RECT  8100.0 41115.0 8165.0 41387.5 ;
      RECT  8132.5 41082.5 8235.0 41147.5 ;
      RECT  13227.5 41355.0 13292.5 41420.0 ;
      RECT  13227.5 40867.5 13292.5 40932.5 ;
      RECT  10525.0 41355.0 13260.0 41420.0 ;
      RECT  13227.5 40900.0 13292.5 41387.5 ;
      RECT  13260.0 40867.5 15995.0 40932.5 ;
      RECT  8100.0 42790.0 8165.0 42855.0 ;
      RECT  8100.0 43062.5 8165.0 43127.5 ;
      RECT  8030.0 42790.0 8132.5 42855.0 ;
      RECT  8100.0 42822.5 8165.0 43095.0 ;
      RECT  8132.5 43062.5 8235.0 43127.5 ;
      RECT  13227.5 42790.0 13292.5 42855.0 ;
      RECT  13227.5 43277.5 13292.5 43342.5 ;
      RECT  10525.0 42790.0 13260.0 42855.0 ;
      RECT  13227.5 42822.5 13292.5 43310.0 ;
      RECT  13260.0 43277.5 15995.0 43342.5 ;
      RECT  8100.0 44045.0 8165.0 44110.0 ;
      RECT  8100.0 43772.5 8165.0 43837.5 ;
      RECT  8030.0 44045.0 8132.5 44110.0 ;
      RECT  8100.0 43805.0 8165.0 44077.5 ;
      RECT  8132.5 43772.5 8235.0 43837.5 ;
      RECT  13227.5 44045.0 13292.5 44110.0 ;
      RECT  13227.5 43557.5 13292.5 43622.5 ;
      RECT  10525.0 44045.0 13260.0 44110.0 ;
      RECT  13227.5 43590.0 13292.5 44077.5 ;
      RECT  13260.0 43557.5 15995.0 43622.5 ;
      RECT  8100.0 45480.0 8165.0 45545.0 ;
      RECT  8100.0 45752.5 8165.0 45817.5 ;
      RECT  8030.0 45480.0 8132.5 45545.0 ;
      RECT  8100.0 45512.5 8165.0 45785.0 ;
      RECT  8132.5 45752.5 8235.0 45817.5 ;
      RECT  13227.5 45480.0 13292.5 45545.0 ;
      RECT  13227.5 45967.5 13292.5 46032.5 ;
      RECT  10525.0 45480.0 13260.0 45545.0 ;
      RECT  13227.5 45512.5 13292.5 46000.0 ;
      RECT  13260.0 45967.5 15995.0 46032.5 ;
      RECT  8100.0 46735.0 8165.0 46800.0 ;
      RECT  8100.0 46462.5 8165.0 46527.5 ;
      RECT  8030.0 46735.0 8132.5 46800.0 ;
      RECT  8100.0 46495.0 8165.0 46767.5 ;
      RECT  8132.5 46462.5 8235.0 46527.5 ;
      RECT  13227.5 46735.0 13292.5 46800.0 ;
      RECT  13227.5 46247.5 13292.5 46312.5 ;
      RECT  10525.0 46735.0 13260.0 46800.0 ;
      RECT  13227.5 46280.0 13292.5 46767.5 ;
      RECT  13260.0 46247.5 15995.0 46312.5 ;
      RECT  8100.0 48170.0 8165.0 48235.0 ;
      RECT  8100.0 48442.5 8165.0 48507.5 ;
      RECT  8030.0 48170.0 8132.5 48235.0 ;
      RECT  8100.0 48202.5 8165.0 48475.0 ;
      RECT  8132.5 48442.5 8235.0 48507.5 ;
      RECT  13227.5 48170.0 13292.5 48235.0 ;
      RECT  13227.5 48657.5 13292.5 48722.5 ;
      RECT  10525.0 48170.0 13260.0 48235.0 ;
      RECT  13227.5 48202.5 13292.5 48690.0 ;
      RECT  13260.0 48657.5 15995.0 48722.5 ;
      RECT  8100.0 49425.0 8165.0 49490.0 ;
      RECT  8100.0 49152.5 8165.0 49217.5 ;
      RECT  8030.0 49425.0 8132.5 49490.0 ;
      RECT  8100.0 49185.0 8165.0 49457.5 ;
      RECT  8132.5 49152.5 8235.0 49217.5 ;
      RECT  13227.5 49425.0 13292.5 49490.0 ;
      RECT  13227.5 48937.5 13292.5 49002.5 ;
      RECT  10525.0 49425.0 13260.0 49490.0 ;
      RECT  13227.5 48970.0 13292.5 49457.5 ;
      RECT  13260.0 48937.5 15995.0 49002.5 ;
      RECT  8100.0 50860.0 8165.0 50925.0 ;
      RECT  8100.0 51132.5 8165.0 51197.5 ;
      RECT  8030.0 50860.0 8132.5 50925.0 ;
      RECT  8100.0 50892.5 8165.0 51165.0 ;
      RECT  8132.5 51132.5 8235.0 51197.5 ;
      RECT  13227.5 50860.0 13292.5 50925.0 ;
      RECT  13227.5 51347.5 13292.5 51412.5 ;
      RECT  10525.0 50860.0 13260.0 50925.0 ;
      RECT  13227.5 50892.5 13292.5 51380.0 ;
      RECT  13260.0 51347.5 15995.0 51412.5 ;
      RECT  8100.0 52115.0 8165.0 52180.0 ;
      RECT  8100.0 51842.5 8165.0 51907.5 ;
      RECT  8030.0 52115.0 8132.5 52180.0 ;
      RECT  8100.0 51875.0 8165.0 52147.5 ;
      RECT  8132.5 51842.5 8235.0 51907.5 ;
      RECT  13227.5 52115.0 13292.5 52180.0 ;
      RECT  13227.5 51627.5 13292.5 51692.5 ;
      RECT  10525.0 52115.0 13260.0 52180.0 ;
      RECT  13227.5 51660.0 13292.5 52147.5 ;
      RECT  13260.0 51627.5 15995.0 51692.5 ;
      RECT  8100.0 53550.0 8165.0 53615.0 ;
      RECT  8100.0 53822.5 8165.0 53887.5 ;
      RECT  8030.0 53550.0 8132.5 53615.0 ;
      RECT  8100.0 53582.5 8165.0 53855.0 ;
      RECT  8132.5 53822.5 8235.0 53887.5 ;
      RECT  13227.5 53550.0 13292.5 53615.0 ;
      RECT  13227.5 54037.5 13292.5 54102.5 ;
      RECT  10525.0 53550.0 13260.0 53615.0 ;
      RECT  13227.5 53582.5 13292.5 54070.0 ;
      RECT  13260.0 54037.5 15995.0 54102.5 ;
      RECT  8100.0 54805.0 8165.0 54870.0 ;
      RECT  8100.0 54532.5 8165.0 54597.5 ;
      RECT  8030.0 54805.0 8132.5 54870.0 ;
      RECT  8100.0 54565.0 8165.0 54837.5 ;
      RECT  8132.5 54532.5 8235.0 54597.5 ;
      RECT  13227.5 54805.0 13292.5 54870.0 ;
      RECT  13227.5 54317.5 13292.5 54382.5 ;
      RECT  10525.0 54805.0 13260.0 54870.0 ;
      RECT  13227.5 54350.0 13292.5 54837.5 ;
      RECT  13260.0 54317.5 15995.0 54382.5 ;
      RECT  8100.0 56240.0 8165.0 56305.0 ;
      RECT  8100.0 56512.5 8165.0 56577.5 ;
      RECT  8030.0 56240.0 8132.5 56305.0 ;
      RECT  8100.0 56272.5 8165.0 56545.0 ;
      RECT  8132.5 56512.5 8235.0 56577.5 ;
      RECT  13227.5 56240.0 13292.5 56305.0 ;
      RECT  13227.5 56727.5 13292.5 56792.5 ;
      RECT  10525.0 56240.0 13260.0 56305.0 ;
      RECT  13227.5 56272.5 13292.5 56760.0 ;
      RECT  13260.0 56727.5 15995.0 56792.5 ;
      RECT  8100.0 57495.0 8165.0 57560.0 ;
      RECT  8100.0 57222.5 8165.0 57287.5 ;
      RECT  8030.0 57495.0 8132.5 57560.0 ;
      RECT  8100.0 57255.0 8165.0 57527.5 ;
      RECT  8132.5 57222.5 8235.0 57287.5 ;
      RECT  13227.5 57495.0 13292.5 57560.0 ;
      RECT  13227.5 57007.5 13292.5 57072.5 ;
      RECT  10525.0 57495.0 13260.0 57560.0 ;
      RECT  13227.5 57040.0 13292.5 57527.5 ;
      RECT  13260.0 57007.5 15995.0 57072.5 ;
      RECT  8100.0 58930.0 8165.0 58995.0 ;
      RECT  8100.0 59202.5 8165.0 59267.5 ;
      RECT  8030.0 58930.0 8132.5 58995.0 ;
      RECT  8100.0 58962.5 8165.0 59235.0 ;
      RECT  8132.5 59202.5 8235.0 59267.5 ;
      RECT  13227.5 58930.0 13292.5 58995.0 ;
      RECT  13227.5 59417.5 13292.5 59482.5 ;
      RECT  10525.0 58930.0 13260.0 58995.0 ;
      RECT  13227.5 58962.5 13292.5 59450.0 ;
      RECT  13260.0 59417.5 15995.0 59482.5 ;
      RECT  8100.0 60185.0 8165.0 60250.0 ;
      RECT  8100.0 59912.5 8165.0 59977.5 ;
      RECT  8030.0 60185.0 8132.5 60250.0 ;
      RECT  8100.0 59945.0 8165.0 60217.5 ;
      RECT  8132.5 59912.5 8235.0 59977.5 ;
      RECT  13227.5 60185.0 13292.5 60250.0 ;
      RECT  13227.5 59697.5 13292.5 59762.5 ;
      RECT  10525.0 60185.0 13260.0 60250.0 ;
      RECT  13227.5 59730.0 13292.5 60217.5 ;
      RECT  13260.0 59697.5 15995.0 59762.5 ;
      RECT  8100.0 61620.0 8165.0 61685.0 ;
      RECT  8100.0 61892.5 8165.0 61957.5 ;
      RECT  8030.0 61620.0 8132.5 61685.0 ;
      RECT  8100.0 61652.5 8165.0 61925.0 ;
      RECT  8132.5 61892.5 8235.0 61957.5 ;
      RECT  13227.5 61620.0 13292.5 61685.0 ;
      RECT  13227.5 62107.5 13292.5 62172.5 ;
      RECT  10525.0 61620.0 13260.0 61685.0 ;
      RECT  13227.5 61652.5 13292.5 62140.0 ;
      RECT  13260.0 62107.5 15995.0 62172.5 ;
      RECT  8100.0 62875.0 8165.0 62940.0 ;
      RECT  8100.0 62602.5 8165.0 62667.5 ;
      RECT  8030.0 62875.0 8132.5 62940.0 ;
      RECT  8100.0 62635.0 8165.0 62907.5 ;
      RECT  8132.5 62602.5 8235.0 62667.5 ;
      RECT  13227.5 62875.0 13292.5 62940.0 ;
      RECT  13227.5 62387.5 13292.5 62452.5 ;
      RECT  10525.0 62875.0 13260.0 62940.0 ;
      RECT  13227.5 62420.0 13292.5 62907.5 ;
      RECT  13260.0 62387.5 15995.0 62452.5 ;
      RECT  8100.0 64310.0 8165.0 64375.0 ;
      RECT  8100.0 64582.5 8165.0 64647.5 ;
      RECT  8030.0 64310.0 8132.5 64375.0 ;
      RECT  8100.0 64342.5 8165.0 64615.0 ;
      RECT  8132.5 64582.5 8235.0 64647.5 ;
      RECT  13227.5 64310.0 13292.5 64375.0 ;
      RECT  13227.5 64797.5 13292.5 64862.5 ;
      RECT  10525.0 64310.0 13260.0 64375.0 ;
      RECT  13227.5 64342.5 13292.5 64830.0 ;
      RECT  13260.0 64797.5 15995.0 64862.5 ;
      RECT  8100.0 65565.0 8165.0 65630.0 ;
      RECT  8100.0 65292.5 8165.0 65357.5 ;
      RECT  8030.0 65565.0 8132.5 65630.0 ;
      RECT  8100.0 65325.0 8165.0 65597.5 ;
      RECT  8132.5 65292.5 8235.0 65357.5 ;
      RECT  13227.5 65565.0 13292.5 65630.0 ;
      RECT  13227.5 65077.5 13292.5 65142.5 ;
      RECT  10525.0 65565.0 13260.0 65630.0 ;
      RECT  13227.5 65110.0 13292.5 65597.5 ;
      RECT  13260.0 65077.5 15995.0 65142.5 ;
      RECT  8100.0 67000.0 8165.0 67065.0 ;
      RECT  8100.0 67272.5 8165.0 67337.5 ;
      RECT  8030.0 67000.0 8132.5 67065.0 ;
      RECT  8100.0 67032.5 8165.0 67305.0 ;
      RECT  8132.5 67272.5 8235.0 67337.5 ;
      RECT  13227.5 67000.0 13292.5 67065.0 ;
      RECT  13227.5 67487.5 13292.5 67552.5 ;
      RECT  10525.0 67000.0 13260.0 67065.0 ;
      RECT  13227.5 67032.5 13292.5 67520.0 ;
      RECT  13260.0 67487.5 15995.0 67552.5 ;
      RECT  8100.0 68255.0 8165.0 68320.0 ;
      RECT  8100.0 67982.5 8165.0 68047.5 ;
      RECT  8030.0 68255.0 8132.5 68320.0 ;
      RECT  8100.0 68015.0 8165.0 68287.5 ;
      RECT  8132.5 67982.5 8235.0 68047.5 ;
      RECT  13227.5 68255.0 13292.5 68320.0 ;
      RECT  13227.5 67767.5 13292.5 67832.5 ;
      RECT  10525.0 68255.0 13260.0 68320.0 ;
      RECT  13227.5 67800.0 13292.5 68287.5 ;
      RECT  13260.0 67767.5 15995.0 67832.5 ;
      RECT  8100.0 69690.0 8165.0 69755.0 ;
      RECT  8100.0 69962.5 8165.0 70027.5 ;
      RECT  8030.0 69690.0 8132.5 69755.0 ;
      RECT  8100.0 69722.5 8165.0 69995.0 ;
      RECT  8132.5 69962.5 8235.0 70027.5 ;
      RECT  13227.5 69690.0 13292.5 69755.0 ;
      RECT  13227.5 70177.5 13292.5 70242.5 ;
      RECT  10525.0 69690.0 13260.0 69755.0 ;
      RECT  13227.5 69722.5 13292.5 70210.0 ;
      RECT  13260.0 70177.5 15995.0 70242.5 ;
      RECT  8690.0 27277.5 16085.0 27342.5 ;
      RECT  8690.0 29967.5 16085.0 30032.5 ;
      RECT  8690.0 32657.5 16085.0 32722.5 ;
      RECT  8690.0 35347.5 16085.0 35412.5 ;
      RECT  8690.0 38037.5 16085.0 38102.5 ;
      RECT  8690.0 40727.5 16085.0 40792.5 ;
      RECT  8690.0 43417.5 16085.0 43482.5 ;
      RECT  8690.0 46107.5 16085.0 46172.5 ;
      RECT  8690.0 48797.5 16085.0 48862.5 ;
      RECT  8690.0 51487.5 16085.0 51552.5 ;
      RECT  8690.0 54177.5 16085.0 54242.5 ;
      RECT  8690.0 56867.5 16085.0 56932.5 ;
      RECT  8690.0 59557.5 16085.0 59622.5 ;
      RECT  8690.0 62247.5 16085.0 62312.5 ;
      RECT  8690.0 64937.5 16085.0 65002.5 ;
      RECT  8690.0 67627.5 16085.0 67692.5 ;
      RECT  8690.0 70317.5 16085.0 70382.5 ;
      RECT  4175.0 28622.5 22270.0 28687.5 ;
      RECT  4175.0 31312.5 22270.0 31377.5 ;
      RECT  4175.0 34002.5 22270.0 34067.5 ;
      RECT  4175.0 36692.5 22270.0 36757.5 ;
      RECT  4175.0 39382.5 22270.0 39447.5 ;
      RECT  4175.0 42072.5 22270.0 42137.5 ;
      RECT  4175.0 44762.5 22270.0 44827.5 ;
      RECT  4175.0 47452.5 22270.0 47517.5 ;
      RECT  4175.0 50142.5 22270.0 50207.5 ;
      RECT  4175.0 52832.5 22270.0 52897.5 ;
      RECT  4175.0 55522.5 22270.0 55587.5 ;
      RECT  4175.0 58212.5 22270.0 58277.5 ;
      RECT  4175.0 60902.5 22270.0 60967.5 ;
      RECT  4175.0 63592.5 22270.0 63657.5 ;
      RECT  4175.0 66282.5 22270.0 66347.5 ;
      RECT  4175.0 68972.5 22270.0 69037.5 ;
      RECT  10720.0 11342.5 11977.5 11407.5 ;
      RECT  10445.0 12687.5 12182.5 12752.5 ;
      RECT  11635.0 16722.5 12387.5 16787.5 ;
      RECT  11360.0 18067.5 12592.5 18132.5 ;
      RECT  11085.0 19412.5 12797.5 19477.5 ;
      RECT  11635.0 11137.5 11772.5 11202.5 ;
      RECT  11635.0 13827.5 11772.5 13892.5 ;
      RECT  11635.0 16517.5 11772.5 16582.5 ;
      RECT  11635.0 19207.5 11772.5 19272.5 ;
      RECT  11635.0 21897.5 11772.5 21962.5 ;
      RECT  11635.0 24587.5 11772.5 24652.5 ;
      RECT  4175.0 12482.5 11635.0 12547.5 ;
      RECT  4175.0 15172.5 11635.0 15237.5 ;
      RECT  4175.0 17862.5 11635.0 17927.5 ;
      RECT  4175.0 20552.5 11635.0 20617.5 ;
      RECT  4175.0 23242.5 11635.0 23307.5 ;
      RECT  4175.0 25932.5 11635.0 25997.5 ;
      RECT  13002.5 25307.5 16085.0 25372.5 ;
      RECT  13207.5 25167.5 16085.0 25232.5 ;
      RECT  13412.5 25027.5 16085.0 25092.5 ;
      RECT  13617.5 24887.5 16085.0 24952.5 ;
      RECT  11225.0 630.0 13002.5 695.0 ;
      RECT  11225.0 2065.0 13207.5 2130.0 ;
      RECT  11225.0 3320.0 13412.5 3385.0 ;
      RECT  11225.0 4755.0 13617.5 4820.0 ;
      RECT  11225.0 2.5 13992.5 67.5 ;
      RECT  11225.0 2692.5 13992.5 2757.5 ;
      RECT  11225.0 5382.5 13992.5 5447.5 ;
      RECT  4175.0 1347.5 13992.5 1412.5 ;
      RECT  4175.0 4037.5 13992.5 4102.5 ;
      RECT  11095.0 10375.0 11977.5 10440.0 ;
      RECT  11095.0 9670.0 12182.5 9735.0 ;
      RECT  11095.0 8965.0 12387.5 9030.0 ;
      RECT  11095.0 8260.0 12592.5 8325.0 ;
      RECT  11095.0 7555.0 12797.5 7620.0 ;
      RECT  11095.0 10727.5 14127.5 10792.5 ;
      RECT  11095.0 10022.5 14127.5 10087.5 ;
      RECT  11095.0 9317.5 14127.5 9382.5 ;
      RECT  11095.0 8612.5 14127.5 8677.5 ;
      RECT  11095.0 7907.5 14127.5 7972.5 ;
      RECT  11095.0 7202.5 14127.5 7267.5 ;
      RECT  11095.0 6497.5 14127.5 6562.5 ;
      RECT  11095.0 5792.5 14127.5 5857.5 ;
      RECT  7865.0 5587.5 7930.0 5652.5 ;
      RECT  7865.0 5620.0 7930.0 5825.0 ;
      RECT  4175.0 5587.5 7897.5 5652.5 ;
      RECT  10825.0 5587.5 10890.0 5652.5 ;
      RECT  10825.0 5620.0 10890.0 5825.0 ;
      RECT  4175.0 5587.5 10857.5 5652.5 ;
      RECT  5875.0 5587.5 5940.0 5652.5 ;
      RECT  5875.0 5620.0 5940.0 5825.0 ;
      RECT  4175.0 5587.5 5907.5 5652.5 ;
      RECT  8835.0 5587.5 8900.0 5652.5 ;
      RECT  8835.0 5620.0 8900.0 5825.0 ;
      RECT  4175.0 5587.5 8867.5 5652.5 ;
      RECT  15197.5 9170.0 16085.0 9235.0 ;
      RECT  14787.5 6985.0 16085.0 7050.0 ;
      RECT  14992.5 8532.5 16085.0 8597.5 ;
      RECT  15197.5 71327.5 16085.0 71392.5 ;
      RECT  15402.5 15672.5 16085.0 15737.5 ;
      RECT  15607.5 19697.5 16085.0 19762.5 ;
      RECT  4860.0 10932.5 4925.0 10997.5 ;
      RECT  4860.0 10760.0 4925.0 10965.0 ;
      RECT  4892.5 10932.5 14582.5 10997.5 ;
      RECT  8465.0 70522.5 14647.5 70587.5 ;
      RECT  16085.0 72012.5 21920.0 72077.5 ;
      RECT  16085.0 24270.0 21920.0 24335.0 ;
      RECT  16085.0 15802.5 21920.0 15867.5 ;
      RECT  16085.0 12175.0 21920.0 12240.0 ;
      RECT  16085.0 15135.0 21920.0 15200.0 ;
      RECT  16085.0 10185.0 21920.0 10250.0 ;
      RECT  16085.0 13145.0 21920.0 13210.0 ;
      RECT  16085.0 7115.0 21920.0 7180.0 ;
      RECT  14342.5 8402.5 16085.0 8467.5 ;
      RECT  14342.5 19827.5 16085.0 19892.5 ;
      RECT  14342.5 9330.0 16085.0 9395.0 ;
      RECT  14342.5 16605.0 16085.0 16670.0 ;
      RECT  16085.0 27310.0 16790.0 28655.0 ;
      RECT  16085.0 30000.0 16790.0 28655.0 ;
      RECT  16085.0 30000.0 16790.0 31345.0 ;
      RECT  16085.0 32690.0 16790.0 31345.0 ;
      RECT  16085.0 32690.0 16790.0 34035.0 ;
      RECT  16085.0 35380.0 16790.0 34035.0 ;
      RECT  16085.0 35380.0 16790.0 36725.0 ;
      RECT  16085.0 38070.0 16790.0 36725.0 ;
      RECT  16085.0 38070.0 16790.0 39415.0 ;
      RECT  16085.0 40760.0 16790.0 39415.0 ;
      RECT  16085.0 40760.0 16790.0 42105.0 ;
      RECT  16085.0 43450.0 16790.0 42105.0 ;
      RECT  16085.0 43450.0 16790.0 44795.0 ;
      RECT  16085.0 46140.0 16790.0 44795.0 ;
      RECT  16085.0 46140.0 16790.0 47485.0 ;
      RECT  16085.0 48830.0 16790.0 47485.0 ;
      RECT  16085.0 48830.0 16790.0 50175.0 ;
      RECT  16085.0 51520.0 16790.0 50175.0 ;
      RECT  16085.0 51520.0 16790.0 52865.0 ;
      RECT  16085.0 54210.0 16790.0 52865.0 ;
      RECT  16085.0 54210.0 16790.0 55555.0 ;
      RECT  16085.0 56900.0 16790.0 55555.0 ;
      RECT  16085.0 56900.0 16790.0 58245.0 ;
      RECT  16085.0 59590.0 16790.0 58245.0 ;
      RECT  16085.0 59590.0 16790.0 60935.0 ;
      RECT  16085.0 62280.0 16790.0 60935.0 ;
      RECT  16085.0 62280.0 16790.0 63625.0 ;
      RECT  16085.0 64970.0 16790.0 63625.0 ;
      RECT  16085.0 64970.0 16790.0 66315.0 ;
      RECT  16085.0 67660.0 16790.0 66315.0 ;
      RECT  16085.0 67660.0 16790.0 69005.0 ;
      RECT  16085.0 70350.0 16790.0 69005.0 ;
      RECT  16790.0 27310.0 17495.0 28655.0 ;
      RECT  16790.0 30000.0 17495.0 28655.0 ;
      RECT  16790.0 30000.0 17495.0 31345.0 ;
      RECT  16790.0 32690.0 17495.0 31345.0 ;
      RECT  16790.0 32690.0 17495.0 34035.0 ;
      RECT  16790.0 35380.0 17495.0 34035.0 ;
      RECT  16790.0 35380.0 17495.0 36725.0 ;
      RECT  16790.0 38070.0 17495.0 36725.0 ;
      RECT  16790.0 38070.0 17495.0 39415.0 ;
      RECT  16790.0 40760.0 17495.0 39415.0 ;
      RECT  16790.0 40760.0 17495.0 42105.0 ;
      RECT  16790.0 43450.0 17495.0 42105.0 ;
      RECT  16790.0 43450.0 17495.0 44795.0 ;
      RECT  16790.0 46140.0 17495.0 44795.0 ;
      RECT  16790.0 46140.0 17495.0 47485.0 ;
      RECT  16790.0 48830.0 17495.0 47485.0 ;
      RECT  16790.0 48830.0 17495.0 50175.0 ;
      RECT  16790.0 51520.0 17495.0 50175.0 ;
      RECT  16790.0 51520.0 17495.0 52865.0 ;
      RECT  16790.0 54210.0 17495.0 52865.0 ;
      RECT  16790.0 54210.0 17495.0 55555.0 ;
      RECT  16790.0 56900.0 17495.0 55555.0 ;
      RECT  16790.0 56900.0 17495.0 58245.0 ;
      RECT  16790.0 59590.0 17495.0 58245.0 ;
      RECT  16790.0 59590.0 17495.0 60935.0 ;
      RECT  16790.0 62280.0 17495.0 60935.0 ;
      RECT  16790.0 62280.0 17495.0 63625.0 ;
      RECT  16790.0 64970.0 17495.0 63625.0 ;
      RECT  16790.0 64970.0 17495.0 66315.0 ;
      RECT  16790.0 67660.0 17495.0 66315.0 ;
      RECT  16790.0 67660.0 17495.0 69005.0 ;
      RECT  16790.0 70350.0 17495.0 69005.0 ;
      RECT  17495.0 27310.0 18200.0 28655.0 ;
      RECT  17495.0 30000.0 18200.0 28655.0 ;
      RECT  17495.0 30000.0 18200.0 31345.0 ;
      RECT  17495.0 32690.0 18200.0 31345.0 ;
      RECT  17495.0 32690.0 18200.0 34035.0 ;
      RECT  17495.0 35380.0 18200.0 34035.0 ;
      RECT  17495.0 35380.0 18200.0 36725.0 ;
      RECT  17495.0 38070.0 18200.0 36725.0 ;
      RECT  17495.0 38070.0 18200.0 39415.0 ;
      RECT  17495.0 40760.0 18200.0 39415.0 ;
      RECT  17495.0 40760.0 18200.0 42105.0 ;
      RECT  17495.0 43450.0 18200.0 42105.0 ;
      RECT  17495.0 43450.0 18200.0 44795.0 ;
      RECT  17495.0 46140.0 18200.0 44795.0 ;
      RECT  17495.0 46140.0 18200.0 47485.0 ;
      RECT  17495.0 48830.0 18200.0 47485.0 ;
      RECT  17495.0 48830.0 18200.0 50175.0 ;
      RECT  17495.0 51520.0 18200.0 50175.0 ;
      RECT  17495.0 51520.0 18200.0 52865.0 ;
      RECT  17495.0 54210.0 18200.0 52865.0 ;
      RECT  17495.0 54210.0 18200.0 55555.0 ;
      RECT  17495.0 56900.0 18200.0 55555.0 ;
      RECT  17495.0 56900.0 18200.0 58245.0 ;
      RECT  17495.0 59590.0 18200.0 58245.0 ;
      RECT  17495.0 59590.0 18200.0 60935.0 ;
      RECT  17495.0 62280.0 18200.0 60935.0 ;
      RECT  17495.0 62280.0 18200.0 63625.0 ;
      RECT  17495.0 64970.0 18200.0 63625.0 ;
      RECT  17495.0 64970.0 18200.0 66315.0 ;
      RECT  17495.0 67660.0 18200.0 66315.0 ;
      RECT  17495.0 67660.0 18200.0 69005.0 ;
      RECT  17495.0 70350.0 18200.0 69005.0 ;
      RECT  18200.0 27310.0 18905.0 28655.0 ;
      RECT  18200.0 30000.0 18905.0 28655.0 ;
      RECT  18200.0 30000.0 18905.0 31345.0 ;
      RECT  18200.0 32690.0 18905.0 31345.0 ;
      RECT  18200.0 32690.0 18905.0 34035.0 ;
      RECT  18200.0 35380.0 18905.0 34035.0 ;
      RECT  18200.0 35380.0 18905.0 36725.0 ;
      RECT  18200.0 38070.0 18905.0 36725.0 ;
      RECT  18200.0 38070.0 18905.0 39415.0 ;
      RECT  18200.0 40760.0 18905.0 39415.0 ;
      RECT  18200.0 40760.0 18905.0 42105.0 ;
      RECT  18200.0 43450.0 18905.0 42105.0 ;
      RECT  18200.0 43450.0 18905.0 44795.0 ;
      RECT  18200.0 46140.0 18905.0 44795.0 ;
      RECT  18200.0 46140.0 18905.0 47485.0 ;
      RECT  18200.0 48830.0 18905.0 47485.0 ;
      RECT  18200.0 48830.0 18905.0 50175.0 ;
      RECT  18200.0 51520.0 18905.0 50175.0 ;
      RECT  18200.0 51520.0 18905.0 52865.0 ;
      RECT  18200.0 54210.0 18905.0 52865.0 ;
      RECT  18200.0 54210.0 18905.0 55555.0 ;
      RECT  18200.0 56900.0 18905.0 55555.0 ;
      RECT  18200.0 56900.0 18905.0 58245.0 ;
      RECT  18200.0 59590.0 18905.0 58245.0 ;
      RECT  18200.0 59590.0 18905.0 60935.0 ;
      RECT  18200.0 62280.0 18905.0 60935.0 ;
      RECT  18200.0 62280.0 18905.0 63625.0 ;
      RECT  18200.0 64970.0 18905.0 63625.0 ;
      RECT  18200.0 64970.0 18905.0 66315.0 ;
      RECT  18200.0 67660.0 18905.0 66315.0 ;
      RECT  18200.0 67660.0 18905.0 69005.0 ;
      RECT  18200.0 70350.0 18905.0 69005.0 ;
      RECT  18905.0 27310.0 19610.0 28655.0 ;
      RECT  18905.0 30000.0 19610.0 28655.0 ;
      RECT  18905.0 30000.0 19610.0 31345.0 ;
      RECT  18905.0 32690.0 19610.0 31345.0 ;
      RECT  18905.0 32690.0 19610.0 34035.0 ;
      RECT  18905.0 35380.0 19610.0 34035.0 ;
      RECT  18905.0 35380.0 19610.0 36725.0 ;
      RECT  18905.0 38070.0 19610.0 36725.0 ;
      RECT  18905.0 38070.0 19610.0 39415.0 ;
      RECT  18905.0 40760.0 19610.0 39415.0 ;
      RECT  18905.0 40760.0 19610.0 42105.0 ;
      RECT  18905.0 43450.0 19610.0 42105.0 ;
      RECT  18905.0 43450.0 19610.0 44795.0 ;
      RECT  18905.0 46140.0 19610.0 44795.0 ;
      RECT  18905.0 46140.0 19610.0 47485.0 ;
      RECT  18905.0 48830.0 19610.0 47485.0 ;
      RECT  18905.0 48830.0 19610.0 50175.0 ;
      RECT  18905.0 51520.0 19610.0 50175.0 ;
      RECT  18905.0 51520.0 19610.0 52865.0 ;
      RECT  18905.0 54210.0 19610.0 52865.0 ;
      RECT  18905.0 54210.0 19610.0 55555.0 ;
      RECT  18905.0 56900.0 19610.0 55555.0 ;
      RECT  18905.0 56900.0 19610.0 58245.0 ;
      RECT  18905.0 59590.0 19610.0 58245.0 ;
      RECT  18905.0 59590.0 19610.0 60935.0 ;
      RECT  18905.0 62280.0 19610.0 60935.0 ;
      RECT  18905.0 62280.0 19610.0 63625.0 ;
      RECT  18905.0 64970.0 19610.0 63625.0 ;
      RECT  18905.0 64970.0 19610.0 66315.0 ;
      RECT  18905.0 67660.0 19610.0 66315.0 ;
      RECT  18905.0 67660.0 19610.0 69005.0 ;
      RECT  18905.0 70350.0 19610.0 69005.0 ;
      RECT  19610.0 27310.0 20315.0 28655.0 ;
      RECT  19610.0 30000.0 20315.0 28655.0 ;
      RECT  19610.0 30000.0 20315.0 31345.0 ;
      RECT  19610.0 32690.0 20315.0 31345.0 ;
      RECT  19610.0 32690.0 20315.0 34035.0 ;
      RECT  19610.0 35380.0 20315.0 34035.0 ;
      RECT  19610.0 35380.0 20315.0 36725.0 ;
      RECT  19610.0 38070.0 20315.0 36725.0 ;
      RECT  19610.0 38070.0 20315.0 39415.0 ;
      RECT  19610.0 40760.0 20315.0 39415.0 ;
      RECT  19610.0 40760.0 20315.0 42105.0 ;
      RECT  19610.0 43450.0 20315.0 42105.0 ;
      RECT  19610.0 43450.0 20315.0 44795.0 ;
      RECT  19610.0 46140.0 20315.0 44795.0 ;
      RECT  19610.0 46140.0 20315.0 47485.0 ;
      RECT  19610.0 48830.0 20315.0 47485.0 ;
      RECT  19610.0 48830.0 20315.0 50175.0 ;
      RECT  19610.0 51520.0 20315.0 50175.0 ;
      RECT  19610.0 51520.0 20315.0 52865.0 ;
      RECT  19610.0 54210.0 20315.0 52865.0 ;
      RECT  19610.0 54210.0 20315.0 55555.0 ;
      RECT  19610.0 56900.0 20315.0 55555.0 ;
      RECT  19610.0 56900.0 20315.0 58245.0 ;
      RECT  19610.0 59590.0 20315.0 58245.0 ;
      RECT  19610.0 59590.0 20315.0 60935.0 ;
      RECT  19610.0 62280.0 20315.0 60935.0 ;
      RECT  19610.0 62280.0 20315.0 63625.0 ;
      RECT  19610.0 64970.0 20315.0 63625.0 ;
      RECT  19610.0 64970.0 20315.0 66315.0 ;
      RECT  19610.0 67660.0 20315.0 66315.0 ;
      RECT  19610.0 67660.0 20315.0 69005.0 ;
      RECT  19610.0 70350.0 20315.0 69005.0 ;
      RECT  20315.0 27310.0 21020.0 28655.0 ;
      RECT  20315.0 30000.0 21020.0 28655.0 ;
      RECT  20315.0 30000.0 21020.0 31345.0 ;
      RECT  20315.0 32690.0 21020.0 31345.0 ;
      RECT  20315.0 32690.0 21020.0 34035.0 ;
      RECT  20315.0 35380.0 21020.0 34035.0 ;
      RECT  20315.0 35380.0 21020.0 36725.0 ;
      RECT  20315.0 38070.0 21020.0 36725.0 ;
      RECT  20315.0 38070.0 21020.0 39415.0 ;
      RECT  20315.0 40760.0 21020.0 39415.0 ;
      RECT  20315.0 40760.0 21020.0 42105.0 ;
      RECT  20315.0 43450.0 21020.0 42105.0 ;
      RECT  20315.0 43450.0 21020.0 44795.0 ;
      RECT  20315.0 46140.0 21020.0 44795.0 ;
      RECT  20315.0 46140.0 21020.0 47485.0 ;
      RECT  20315.0 48830.0 21020.0 47485.0 ;
      RECT  20315.0 48830.0 21020.0 50175.0 ;
      RECT  20315.0 51520.0 21020.0 50175.0 ;
      RECT  20315.0 51520.0 21020.0 52865.0 ;
      RECT  20315.0 54210.0 21020.0 52865.0 ;
      RECT  20315.0 54210.0 21020.0 55555.0 ;
      RECT  20315.0 56900.0 21020.0 55555.0 ;
      RECT  20315.0 56900.0 21020.0 58245.0 ;
      RECT  20315.0 59590.0 21020.0 58245.0 ;
      RECT  20315.0 59590.0 21020.0 60935.0 ;
      RECT  20315.0 62280.0 21020.0 60935.0 ;
      RECT  20315.0 62280.0 21020.0 63625.0 ;
      RECT  20315.0 64970.0 21020.0 63625.0 ;
      RECT  20315.0 64970.0 21020.0 66315.0 ;
      RECT  20315.0 67660.0 21020.0 66315.0 ;
      RECT  20315.0 67660.0 21020.0 69005.0 ;
      RECT  20315.0 70350.0 21020.0 69005.0 ;
      RECT  21020.0 27310.0 21725.0 28655.0 ;
      RECT  21020.0 30000.0 21725.0 28655.0 ;
      RECT  21020.0 30000.0 21725.0 31345.0 ;
      RECT  21020.0 32690.0 21725.0 31345.0 ;
      RECT  21020.0 32690.0 21725.0 34035.0 ;
      RECT  21020.0 35380.0 21725.0 34035.0 ;
      RECT  21020.0 35380.0 21725.0 36725.0 ;
      RECT  21020.0 38070.0 21725.0 36725.0 ;
      RECT  21020.0 38070.0 21725.0 39415.0 ;
      RECT  21020.0 40760.0 21725.0 39415.0 ;
      RECT  21020.0 40760.0 21725.0 42105.0 ;
      RECT  21020.0 43450.0 21725.0 42105.0 ;
      RECT  21020.0 43450.0 21725.0 44795.0 ;
      RECT  21020.0 46140.0 21725.0 44795.0 ;
      RECT  21020.0 46140.0 21725.0 47485.0 ;
      RECT  21020.0 48830.0 21725.0 47485.0 ;
      RECT  21020.0 48830.0 21725.0 50175.0 ;
      RECT  21020.0 51520.0 21725.0 50175.0 ;
      RECT  21020.0 51520.0 21725.0 52865.0 ;
      RECT  21020.0 54210.0 21725.0 52865.0 ;
      RECT  21020.0 54210.0 21725.0 55555.0 ;
      RECT  21020.0 56900.0 21725.0 55555.0 ;
      RECT  21020.0 56900.0 21725.0 58245.0 ;
      RECT  21020.0 59590.0 21725.0 58245.0 ;
      RECT  21020.0 59590.0 21725.0 60935.0 ;
      RECT  21020.0 62280.0 21725.0 60935.0 ;
      RECT  21020.0 62280.0 21725.0 63625.0 ;
      RECT  21020.0 64970.0 21725.0 63625.0 ;
      RECT  21020.0 64970.0 21725.0 66315.0 ;
      RECT  21020.0 67660.0 21725.0 66315.0 ;
      RECT  21020.0 67660.0 21725.0 69005.0 ;
      RECT  21020.0 70350.0 21725.0 69005.0 ;
      RECT  15995.0 27417.5 21815.0 27482.5 ;
      RECT  15995.0 29827.5 21815.0 29892.5 ;
      RECT  15995.0 30107.5 21815.0 30172.5 ;
      RECT  15995.0 32517.5 21815.0 32582.5 ;
      RECT  15995.0 32797.5 21815.0 32862.5 ;
      RECT  15995.0 35207.5 21815.0 35272.5 ;
      RECT  15995.0 35487.5 21815.0 35552.5 ;
      RECT  15995.0 37897.5 21815.0 37962.5 ;
      RECT  15995.0 38177.5 21815.0 38242.5 ;
      RECT  15995.0 40587.5 21815.0 40652.5 ;
      RECT  15995.0 40867.5 21815.0 40932.5 ;
      RECT  15995.0 43277.5 21815.0 43342.5 ;
      RECT  15995.0 43557.5 21815.0 43622.5 ;
      RECT  15995.0 45967.5 21815.0 46032.5 ;
      RECT  15995.0 46247.5 21815.0 46312.5 ;
      RECT  15995.0 48657.5 21815.0 48722.5 ;
      RECT  15995.0 48937.5 21815.0 49002.5 ;
      RECT  15995.0 51347.5 21815.0 51412.5 ;
      RECT  15995.0 51627.5 21815.0 51692.5 ;
      RECT  15995.0 54037.5 21815.0 54102.5 ;
      RECT  15995.0 54317.5 21815.0 54382.5 ;
      RECT  15995.0 56727.5 21815.0 56792.5 ;
      RECT  15995.0 57007.5 21815.0 57072.5 ;
      RECT  15995.0 59417.5 21815.0 59482.5 ;
      RECT  15995.0 59697.5 21815.0 59762.5 ;
      RECT  15995.0 62107.5 21815.0 62172.5 ;
      RECT  15995.0 62387.5 21815.0 62452.5 ;
      RECT  15995.0 64797.5 21815.0 64862.5 ;
      RECT  15995.0 65077.5 21815.0 65142.5 ;
      RECT  15995.0 67487.5 21815.0 67552.5 ;
      RECT  15995.0 67767.5 21815.0 67832.5 ;
      RECT  15995.0 70177.5 21815.0 70242.5 ;
      RECT  15995.0 28622.5 21815.0 28687.5 ;
      RECT  15995.0 31312.5 21815.0 31377.5 ;
      RECT  15995.0 34002.5 21815.0 34067.5 ;
      RECT  15995.0 36692.5 21815.0 36757.5 ;
      RECT  15995.0 39382.5 21815.0 39447.5 ;
      RECT  15995.0 42072.5 21815.0 42137.5 ;
      RECT  15995.0 44762.5 21815.0 44827.5 ;
      RECT  15995.0 47452.5 21815.0 47517.5 ;
      RECT  15995.0 50142.5 21815.0 50207.5 ;
      RECT  15995.0 52832.5 21815.0 52897.5 ;
      RECT  15995.0 55522.5 21815.0 55587.5 ;
      RECT  15995.0 58212.5 21815.0 58277.5 ;
      RECT  15995.0 60902.5 21815.0 60967.5 ;
      RECT  15995.0 63592.5 21815.0 63657.5 ;
      RECT  15995.0 66282.5 21815.0 66347.5 ;
      RECT  15995.0 68972.5 21815.0 69037.5 ;
      RECT  15995.0 27277.5 21815.0 27342.5 ;
      RECT  15995.0 29967.5 21815.0 30032.5 ;
      RECT  15995.0 32657.5 21815.0 32722.5 ;
      RECT  15995.0 35347.5 21815.0 35412.5 ;
      RECT  15995.0 38037.5 21815.0 38102.5 ;
      RECT  15995.0 40727.5 21815.0 40792.5 ;
      RECT  15995.0 43417.5 21815.0 43482.5 ;
      RECT  15995.0 46107.5 21815.0 46172.5 ;
      RECT  15995.0 48797.5 21815.0 48862.5 ;
      RECT  15995.0 51487.5 21815.0 51552.5 ;
      RECT  15995.0 54177.5 21815.0 54242.5 ;
      RECT  15995.0 56867.5 21815.0 56932.5 ;
      RECT  15995.0 59557.5 21815.0 59622.5 ;
      RECT  15995.0 62247.5 21815.0 62312.5 ;
      RECT  15995.0 64937.5 21815.0 65002.5 ;
      RECT  15995.0 67627.5 21815.0 67692.5 ;
      RECT  15995.0 70317.5 21815.0 70382.5 ;
      RECT  16437.5 71562.5 16502.5 72077.5 ;
      RECT  16247.5 71032.5 16312.5 71167.5 ;
      RECT  16437.5 71032.5 16502.5 71167.5 ;
      RECT  16437.5 71032.5 16502.5 71167.5 ;
      RECT  16247.5 71032.5 16312.5 71167.5 ;
      RECT  16247.5 71562.5 16312.5 71697.5 ;
      RECT  16437.5 71562.5 16502.5 71697.5 ;
      RECT  16437.5 71562.5 16502.5 71697.5 ;
      RECT  16247.5 71562.5 16312.5 71697.5 ;
      RECT  16437.5 71562.5 16502.5 71697.5 ;
      RECT  16627.5 71562.5 16692.5 71697.5 ;
      RECT  16627.5 71562.5 16692.5 71697.5 ;
      RECT  16437.5 71562.5 16502.5 71697.5 ;
      RECT  16417.5 71327.5 16282.5 71392.5 ;
      RECT  16437.5 71875.0 16502.5 72010.0 ;
      RECT  16247.5 71032.5 16312.5 71167.5 ;
      RECT  16437.5 71032.5 16502.5 71167.5 ;
      RECT  16247.5 71562.5 16312.5 71697.5 ;
      RECT  16627.5 71562.5 16692.5 71697.5 ;
      RECT  16085.0 71327.5 16790.0 71392.5 ;
      RECT  16085.0 72012.5 16790.0 72077.5 ;
      RECT  17142.5 71562.5 17207.5 72077.5 ;
      RECT  16952.5 71032.5 17017.5 71167.5 ;
      RECT  17142.5 71032.5 17207.5 71167.5 ;
      RECT  17142.5 71032.5 17207.5 71167.5 ;
      RECT  16952.5 71032.5 17017.5 71167.5 ;
      RECT  16952.5 71562.5 17017.5 71697.5 ;
      RECT  17142.5 71562.5 17207.5 71697.5 ;
      RECT  17142.5 71562.5 17207.5 71697.5 ;
      RECT  16952.5 71562.5 17017.5 71697.5 ;
      RECT  17142.5 71562.5 17207.5 71697.5 ;
      RECT  17332.5 71562.5 17397.5 71697.5 ;
      RECT  17332.5 71562.5 17397.5 71697.5 ;
      RECT  17142.5 71562.5 17207.5 71697.5 ;
      RECT  17122.5 71327.5 16987.5 71392.5 ;
      RECT  17142.5 71875.0 17207.5 72010.0 ;
      RECT  16952.5 71032.5 17017.5 71167.5 ;
      RECT  17142.5 71032.5 17207.5 71167.5 ;
      RECT  16952.5 71562.5 17017.5 71697.5 ;
      RECT  17332.5 71562.5 17397.5 71697.5 ;
      RECT  16790.0 71327.5 17495.0 71392.5 ;
      RECT  16790.0 72012.5 17495.0 72077.5 ;
      RECT  17847.5 71562.5 17912.5 72077.5 ;
      RECT  17657.5 71032.5 17722.5 71167.5 ;
      RECT  17847.5 71032.5 17912.5 71167.5 ;
      RECT  17847.5 71032.5 17912.5 71167.5 ;
      RECT  17657.5 71032.5 17722.5 71167.5 ;
      RECT  17657.5 71562.5 17722.5 71697.5 ;
      RECT  17847.5 71562.5 17912.5 71697.5 ;
      RECT  17847.5 71562.5 17912.5 71697.5 ;
      RECT  17657.5 71562.5 17722.5 71697.5 ;
      RECT  17847.5 71562.5 17912.5 71697.5 ;
      RECT  18037.5 71562.5 18102.5 71697.5 ;
      RECT  18037.5 71562.5 18102.5 71697.5 ;
      RECT  17847.5 71562.5 17912.5 71697.5 ;
      RECT  17827.5 71327.5 17692.5 71392.5 ;
      RECT  17847.5 71875.0 17912.5 72010.0 ;
      RECT  17657.5 71032.5 17722.5 71167.5 ;
      RECT  17847.5 71032.5 17912.5 71167.5 ;
      RECT  17657.5 71562.5 17722.5 71697.5 ;
      RECT  18037.5 71562.5 18102.5 71697.5 ;
      RECT  17495.0 71327.5 18200.0 71392.5 ;
      RECT  17495.0 72012.5 18200.0 72077.5 ;
      RECT  18552.5 71562.5 18617.5 72077.5 ;
      RECT  18362.5 71032.5 18427.5 71167.5 ;
      RECT  18552.5 71032.5 18617.5 71167.5 ;
      RECT  18552.5 71032.5 18617.5 71167.5 ;
      RECT  18362.5 71032.5 18427.5 71167.5 ;
      RECT  18362.5 71562.5 18427.5 71697.5 ;
      RECT  18552.5 71562.5 18617.5 71697.5 ;
      RECT  18552.5 71562.5 18617.5 71697.5 ;
      RECT  18362.5 71562.5 18427.5 71697.5 ;
      RECT  18552.5 71562.5 18617.5 71697.5 ;
      RECT  18742.5 71562.5 18807.5 71697.5 ;
      RECT  18742.5 71562.5 18807.5 71697.5 ;
      RECT  18552.5 71562.5 18617.5 71697.5 ;
      RECT  18532.5 71327.5 18397.5 71392.5 ;
      RECT  18552.5 71875.0 18617.5 72010.0 ;
      RECT  18362.5 71032.5 18427.5 71167.5 ;
      RECT  18552.5 71032.5 18617.5 71167.5 ;
      RECT  18362.5 71562.5 18427.5 71697.5 ;
      RECT  18742.5 71562.5 18807.5 71697.5 ;
      RECT  18200.0 71327.5 18905.0 71392.5 ;
      RECT  18200.0 72012.5 18905.0 72077.5 ;
      RECT  19257.5 71562.5 19322.5 72077.5 ;
      RECT  19067.5 71032.5 19132.5 71167.5 ;
      RECT  19257.5 71032.5 19322.5 71167.5 ;
      RECT  19257.5 71032.5 19322.5 71167.5 ;
      RECT  19067.5 71032.5 19132.5 71167.5 ;
      RECT  19067.5 71562.5 19132.5 71697.5 ;
      RECT  19257.5 71562.5 19322.5 71697.5 ;
      RECT  19257.5 71562.5 19322.5 71697.5 ;
      RECT  19067.5 71562.5 19132.5 71697.5 ;
      RECT  19257.5 71562.5 19322.5 71697.5 ;
      RECT  19447.5 71562.5 19512.5 71697.5 ;
      RECT  19447.5 71562.5 19512.5 71697.5 ;
      RECT  19257.5 71562.5 19322.5 71697.5 ;
      RECT  19237.5 71327.5 19102.5 71392.5 ;
      RECT  19257.5 71875.0 19322.5 72010.0 ;
      RECT  19067.5 71032.5 19132.5 71167.5 ;
      RECT  19257.5 71032.5 19322.5 71167.5 ;
      RECT  19067.5 71562.5 19132.5 71697.5 ;
      RECT  19447.5 71562.5 19512.5 71697.5 ;
      RECT  18905.0 71327.5 19610.0 71392.5 ;
      RECT  18905.0 72012.5 19610.0 72077.5 ;
      RECT  19962.5 71562.5 20027.5 72077.5 ;
      RECT  19772.5 71032.5 19837.5 71167.5 ;
      RECT  19962.5 71032.5 20027.5 71167.5 ;
      RECT  19962.5 71032.5 20027.5 71167.5 ;
      RECT  19772.5 71032.5 19837.5 71167.5 ;
      RECT  19772.5 71562.5 19837.5 71697.5 ;
      RECT  19962.5 71562.5 20027.5 71697.5 ;
      RECT  19962.5 71562.5 20027.5 71697.5 ;
      RECT  19772.5 71562.5 19837.5 71697.5 ;
      RECT  19962.5 71562.5 20027.5 71697.5 ;
      RECT  20152.5 71562.5 20217.5 71697.5 ;
      RECT  20152.5 71562.5 20217.5 71697.5 ;
      RECT  19962.5 71562.5 20027.5 71697.5 ;
      RECT  19942.5 71327.5 19807.5 71392.5 ;
      RECT  19962.5 71875.0 20027.5 72010.0 ;
      RECT  19772.5 71032.5 19837.5 71167.5 ;
      RECT  19962.5 71032.5 20027.5 71167.5 ;
      RECT  19772.5 71562.5 19837.5 71697.5 ;
      RECT  20152.5 71562.5 20217.5 71697.5 ;
      RECT  19610.0 71327.5 20315.0 71392.5 ;
      RECT  19610.0 72012.5 20315.0 72077.5 ;
      RECT  20667.5 71562.5 20732.5 72077.5 ;
      RECT  20477.5 71032.5 20542.5 71167.5 ;
      RECT  20667.5 71032.5 20732.5 71167.5 ;
      RECT  20667.5 71032.5 20732.5 71167.5 ;
      RECT  20477.5 71032.5 20542.5 71167.5 ;
      RECT  20477.5 71562.5 20542.5 71697.5 ;
      RECT  20667.5 71562.5 20732.5 71697.5 ;
      RECT  20667.5 71562.5 20732.5 71697.5 ;
      RECT  20477.5 71562.5 20542.5 71697.5 ;
      RECT  20667.5 71562.5 20732.5 71697.5 ;
      RECT  20857.5 71562.5 20922.5 71697.5 ;
      RECT  20857.5 71562.5 20922.5 71697.5 ;
      RECT  20667.5 71562.5 20732.5 71697.5 ;
      RECT  20647.5 71327.5 20512.5 71392.5 ;
      RECT  20667.5 71875.0 20732.5 72010.0 ;
      RECT  20477.5 71032.5 20542.5 71167.5 ;
      RECT  20667.5 71032.5 20732.5 71167.5 ;
      RECT  20477.5 71562.5 20542.5 71697.5 ;
      RECT  20857.5 71562.5 20922.5 71697.5 ;
      RECT  20315.0 71327.5 21020.0 71392.5 ;
      RECT  20315.0 72012.5 21020.0 72077.5 ;
      RECT  21372.5 71562.5 21437.5 72077.5 ;
      RECT  21182.5 71032.5 21247.5 71167.5 ;
      RECT  21372.5 71032.5 21437.5 71167.5 ;
      RECT  21372.5 71032.5 21437.5 71167.5 ;
      RECT  21182.5 71032.5 21247.5 71167.5 ;
      RECT  21182.5 71562.5 21247.5 71697.5 ;
      RECT  21372.5 71562.5 21437.5 71697.5 ;
      RECT  21372.5 71562.5 21437.5 71697.5 ;
      RECT  21182.5 71562.5 21247.5 71697.5 ;
      RECT  21372.5 71562.5 21437.5 71697.5 ;
      RECT  21562.5 71562.5 21627.5 71697.5 ;
      RECT  21562.5 71562.5 21627.5 71697.5 ;
      RECT  21372.5 71562.5 21437.5 71697.5 ;
      RECT  21352.5 71327.5 21217.5 71392.5 ;
      RECT  21372.5 71875.0 21437.5 72010.0 ;
      RECT  21182.5 71032.5 21247.5 71167.5 ;
      RECT  21372.5 71032.5 21437.5 71167.5 ;
      RECT  21182.5 71562.5 21247.5 71697.5 ;
      RECT  21562.5 71562.5 21627.5 71697.5 ;
      RECT  21020.0 71327.5 21725.0 71392.5 ;
      RECT  21020.0 72012.5 21725.0 72077.5 ;
      RECT  16085.0 71327.5 21725.0 71392.5 ;
      RECT  16085.0 72012.5 21725.0 72077.5 ;
      RECT  16235.0 24745.0 18420.0 24815.0 ;
      RECT  16570.0 24605.0 18755.0 24675.0 ;
      RECT  19055.0 24745.0 21240.0 24815.0 ;
      RECT  19390.0 24605.0 21575.0 24675.0 ;
      RECT  16500.0 27102.5 16565.0 27167.5 ;
      RECT  16235.0 27102.5 16532.5 27167.5 ;
      RECT  16500.0 26720.0 16565.0 27135.0 ;
      RECT  16310.0 25552.5 16375.0 25617.5 ;
      RECT  16342.5 25552.5 16605.0 25617.5 ;
      RECT  16310.0 25585.0 16375.0 25860.0 ;
      RECT  16310.0 25792.5 16375.0 25927.5 ;
      RECT  16500.0 25792.5 16565.0 25927.5 ;
      RECT  16500.0 25792.5 16565.0 25927.5 ;
      RECT  16310.0 25792.5 16375.0 25927.5 ;
      RECT  16310.0 26652.5 16375.0 26787.5 ;
      RECT  16500.0 26652.5 16565.0 26787.5 ;
      RECT  16500.0 26652.5 16565.0 26787.5 ;
      RECT  16310.0 26652.5 16375.0 26787.5 ;
      RECT  16237.5 27067.5 16302.5 27202.5 ;
      RECT  16572.5 25517.5 16637.5 25652.5 ;
      RECT  16310.0 26652.5 16375.0 26787.5 ;
      RECT  16500.0 25792.5 16565.0 25927.5 ;
      RECT  16757.5 25692.5 16822.5 25827.5 ;
      RECT  16757.5 25692.5 16822.5 25827.5 ;
      RECT  17205.0 27102.5 17270.0 27167.5 ;
      RECT  16940.0 27102.5 17237.5 27167.5 ;
      RECT  17205.0 26720.0 17270.0 27135.0 ;
      RECT  17015.0 25552.5 17080.0 25617.5 ;
      RECT  17047.5 25552.5 17310.0 25617.5 ;
      RECT  17015.0 25585.0 17080.0 25860.0 ;
      RECT  17015.0 25792.5 17080.0 25927.5 ;
      RECT  17205.0 25792.5 17270.0 25927.5 ;
      RECT  17205.0 25792.5 17270.0 25927.5 ;
      RECT  17015.0 25792.5 17080.0 25927.5 ;
      RECT  17015.0 26652.5 17080.0 26787.5 ;
      RECT  17205.0 26652.5 17270.0 26787.5 ;
      RECT  17205.0 26652.5 17270.0 26787.5 ;
      RECT  17015.0 26652.5 17080.0 26787.5 ;
      RECT  16942.5 27067.5 17007.5 27202.5 ;
      RECT  17277.5 25517.5 17342.5 25652.5 ;
      RECT  17015.0 26652.5 17080.0 26787.5 ;
      RECT  17205.0 25792.5 17270.0 25927.5 ;
      RECT  17462.5 25692.5 17527.5 25827.5 ;
      RECT  17462.5 25692.5 17527.5 25827.5 ;
      RECT  17910.0 27102.5 17975.0 27167.5 ;
      RECT  17645.0 27102.5 17942.5 27167.5 ;
      RECT  17910.0 26720.0 17975.0 27135.0 ;
      RECT  17720.0 25552.5 17785.0 25617.5 ;
      RECT  17752.5 25552.5 18015.0 25617.5 ;
      RECT  17720.0 25585.0 17785.0 25860.0 ;
      RECT  17720.0 25792.5 17785.0 25927.5 ;
      RECT  17910.0 25792.5 17975.0 25927.5 ;
      RECT  17910.0 25792.5 17975.0 25927.5 ;
      RECT  17720.0 25792.5 17785.0 25927.5 ;
      RECT  17720.0 26652.5 17785.0 26787.5 ;
      RECT  17910.0 26652.5 17975.0 26787.5 ;
      RECT  17910.0 26652.5 17975.0 26787.5 ;
      RECT  17720.0 26652.5 17785.0 26787.5 ;
      RECT  17647.5 27067.5 17712.5 27202.5 ;
      RECT  17982.5 25517.5 18047.5 25652.5 ;
      RECT  17720.0 26652.5 17785.0 26787.5 ;
      RECT  17910.0 25792.5 17975.0 25927.5 ;
      RECT  18167.5 25692.5 18232.5 25827.5 ;
      RECT  18167.5 25692.5 18232.5 25827.5 ;
      RECT  18615.0 27102.5 18680.0 27167.5 ;
      RECT  18350.0 27102.5 18647.5 27167.5 ;
      RECT  18615.0 26720.0 18680.0 27135.0 ;
      RECT  18425.0 25552.5 18490.0 25617.5 ;
      RECT  18457.5 25552.5 18720.0 25617.5 ;
      RECT  18425.0 25585.0 18490.0 25860.0 ;
      RECT  18425.0 25792.5 18490.0 25927.5 ;
      RECT  18615.0 25792.5 18680.0 25927.5 ;
      RECT  18615.0 25792.5 18680.0 25927.5 ;
      RECT  18425.0 25792.5 18490.0 25927.5 ;
      RECT  18425.0 26652.5 18490.0 26787.5 ;
      RECT  18615.0 26652.5 18680.0 26787.5 ;
      RECT  18615.0 26652.5 18680.0 26787.5 ;
      RECT  18425.0 26652.5 18490.0 26787.5 ;
      RECT  18352.5 27067.5 18417.5 27202.5 ;
      RECT  18687.5 25517.5 18752.5 25652.5 ;
      RECT  18425.0 26652.5 18490.0 26787.5 ;
      RECT  18615.0 25792.5 18680.0 25927.5 ;
      RECT  18872.5 25692.5 18937.5 25827.5 ;
      RECT  18872.5 25692.5 18937.5 25827.5 ;
      RECT  19320.0 27102.5 19385.0 27167.5 ;
      RECT  19055.0 27102.5 19352.5 27167.5 ;
      RECT  19320.0 26720.0 19385.0 27135.0 ;
      RECT  19130.0 25552.5 19195.0 25617.5 ;
      RECT  19162.5 25552.5 19425.0 25617.5 ;
      RECT  19130.0 25585.0 19195.0 25860.0 ;
      RECT  19130.0 25792.5 19195.0 25927.5 ;
      RECT  19320.0 25792.5 19385.0 25927.5 ;
      RECT  19320.0 25792.5 19385.0 25927.5 ;
      RECT  19130.0 25792.5 19195.0 25927.5 ;
      RECT  19130.0 26652.5 19195.0 26787.5 ;
      RECT  19320.0 26652.5 19385.0 26787.5 ;
      RECT  19320.0 26652.5 19385.0 26787.5 ;
      RECT  19130.0 26652.5 19195.0 26787.5 ;
      RECT  19057.5 27067.5 19122.5 27202.5 ;
      RECT  19392.5 25517.5 19457.5 25652.5 ;
      RECT  19130.0 26652.5 19195.0 26787.5 ;
      RECT  19320.0 25792.5 19385.0 25927.5 ;
      RECT  19577.5 25692.5 19642.5 25827.5 ;
      RECT  19577.5 25692.5 19642.5 25827.5 ;
      RECT  20025.0 27102.5 20090.0 27167.5 ;
      RECT  19760.0 27102.5 20057.5 27167.5 ;
      RECT  20025.0 26720.0 20090.0 27135.0 ;
      RECT  19835.0 25552.5 19900.0 25617.5 ;
      RECT  19867.5 25552.5 20130.0 25617.5 ;
      RECT  19835.0 25585.0 19900.0 25860.0 ;
      RECT  19835.0 25792.5 19900.0 25927.5 ;
      RECT  20025.0 25792.5 20090.0 25927.5 ;
      RECT  20025.0 25792.5 20090.0 25927.5 ;
      RECT  19835.0 25792.5 19900.0 25927.5 ;
      RECT  19835.0 26652.5 19900.0 26787.5 ;
      RECT  20025.0 26652.5 20090.0 26787.5 ;
      RECT  20025.0 26652.5 20090.0 26787.5 ;
      RECT  19835.0 26652.5 19900.0 26787.5 ;
      RECT  19762.5 27067.5 19827.5 27202.5 ;
      RECT  20097.5 25517.5 20162.5 25652.5 ;
      RECT  19835.0 26652.5 19900.0 26787.5 ;
      RECT  20025.0 25792.5 20090.0 25927.5 ;
      RECT  20282.5 25692.5 20347.5 25827.5 ;
      RECT  20282.5 25692.5 20347.5 25827.5 ;
      RECT  20730.0 27102.5 20795.0 27167.5 ;
      RECT  20465.0 27102.5 20762.5 27167.5 ;
      RECT  20730.0 26720.0 20795.0 27135.0 ;
      RECT  20540.0 25552.5 20605.0 25617.5 ;
      RECT  20572.5 25552.5 20835.0 25617.5 ;
      RECT  20540.0 25585.0 20605.0 25860.0 ;
      RECT  20540.0 25792.5 20605.0 25927.5 ;
      RECT  20730.0 25792.5 20795.0 25927.5 ;
      RECT  20730.0 25792.5 20795.0 25927.5 ;
      RECT  20540.0 25792.5 20605.0 25927.5 ;
      RECT  20540.0 26652.5 20605.0 26787.5 ;
      RECT  20730.0 26652.5 20795.0 26787.5 ;
      RECT  20730.0 26652.5 20795.0 26787.5 ;
      RECT  20540.0 26652.5 20605.0 26787.5 ;
      RECT  20467.5 27067.5 20532.5 27202.5 ;
      RECT  20802.5 25517.5 20867.5 25652.5 ;
      RECT  20540.0 26652.5 20605.0 26787.5 ;
      RECT  20730.0 25792.5 20795.0 25927.5 ;
      RECT  20987.5 25692.5 21052.5 25827.5 ;
      RECT  20987.5 25692.5 21052.5 25827.5 ;
      RECT  21435.0 27102.5 21500.0 27167.5 ;
      RECT  21170.0 27102.5 21467.5 27167.5 ;
      RECT  21435.0 26720.0 21500.0 27135.0 ;
      RECT  21245.0 25552.5 21310.0 25617.5 ;
      RECT  21277.5 25552.5 21540.0 25617.5 ;
      RECT  21245.0 25585.0 21310.0 25860.0 ;
      RECT  21245.0 25792.5 21310.0 25927.5 ;
      RECT  21435.0 25792.5 21500.0 25927.5 ;
      RECT  21435.0 25792.5 21500.0 25927.5 ;
      RECT  21245.0 25792.5 21310.0 25927.5 ;
      RECT  21245.0 26652.5 21310.0 26787.5 ;
      RECT  21435.0 26652.5 21500.0 26787.5 ;
      RECT  21435.0 26652.5 21500.0 26787.5 ;
      RECT  21245.0 26652.5 21310.0 26787.5 ;
      RECT  21172.5 27067.5 21237.5 27202.5 ;
      RECT  21507.5 25517.5 21572.5 25652.5 ;
      RECT  21245.0 26652.5 21310.0 26787.5 ;
      RECT  21435.0 25792.5 21500.0 25927.5 ;
      RECT  21692.5 25692.5 21757.5 25827.5 ;
      RECT  21692.5 25692.5 21757.5 25827.5 ;
      RECT  16505.0 25307.5 16370.0 25372.5 ;
      RECT  17210.0 25167.5 17075.0 25232.5 ;
      RECT  17915.0 25027.5 17780.0 25092.5 ;
      RECT  18620.0 24887.5 18485.0 24952.5 ;
      RECT  19325.0 25307.5 19190.0 25372.5 ;
      RECT  20030.0 25167.5 19895.0 25232.5 ;
      RECT  20735.0 25027.5 20600.0 25092.5 ;
      RECT  21440.0 24887.5 21305.0 24952.5 ;
      RECT  16370.0 24747.5 16235.0 24812.5 ;
      RECT  16570.0 24607.5 16435.0 24672.5 ;
      RECT  17075.0 24747.5 16940.0 24812.5 ;
      RECT  17275.0 24607.5 17140.0 24672.5 ;
      RECT  17780.0 24747.5 17645.0 24812.5 ;
      RECT  17980.0 24607.5 17845.0 24672.5 ;
      RECT  18485.0 24747.5 18350.0 24812.5 ;
      RECT  18685.0 24607.5 18550.0 24672.5 ;
      RECT  19190.0 24747.5 19055.0 24812.5 ;
      RECT  19390.0 24607.5 19255.0 24672.5 ;
      RECT  19895.0 24747.5 19760.0 24812.5 ;
      RECT  20095.0 24607.5 19960.0 24672.5 ;
      RECT  20600.0 24747.5 20465.0 24812.5 ;
      RECT  20800.0 24607.5 20665.0 24672.5 ;
      RECT  21305.0 24747.5 21170.0 24812.5 ;
      RECT  21505.0 24607.5 21370.0 24672.5 ;
      RECT  16085.0 25305.0 21725.0 25375.0 ;
      RECT  16085.0 25165.0 21725.0 25235.0 ;
      RECT  16085.0 25025.0 21725.0 25095.0 ;
      RECT  16085.0 24885.0 21725.0 24955.0 ;
      RECT  8402.5 630.0 8467.5 695.0 ;
      RECT  8402.5 1152.5 8467.5 1217.5 ;
      RECT  8165.0 630.0 8435.0 695.0 ;
      RECT  8402.5 662.5 8467.5 1185.0 ;
      RECT  8435.0 1152.5 8680.0 1217.5 ;
      RECT  7295.0 630.0 7935.0 695.0 ;
      RECT  8402.5 2065.0 8467.5 2130.0 ;
      RECT  8402.5 2497.5 8467.5 2562.5 ;
      RECT  8165.0 2065.0 8435.0 2130.0 ;
      RECT  8402.5 2097.5 8467.5 2530.0 ;
      RECT  8435.0 2497.5 8955.0 2562.5 ;
      RECT  7570.0 2065.0 7935.0 2130.0 ;
      RECT  7295.0 2827.5 9230.0 2892.5 ;
      RECT  7570.0 4172.5 9505.0 4237.5 ;
      RECT  8680.0 642.5 9805.0 707.5 ;
      RECT  8955.0 427.5 10062.5 492.5 ;
      RECT  9230.0 2052.5 9805.0 2117.5 ;
      RECT  8955.0 2267.5 10062.5 2332.5 ;
      RECT  8680.0 3332.5 9805.0 3397.5 ;
      RECT  9505.0 3117.5 10062.5 3182.5 ;
      RECT  9230.0 4742.5 9805.0 4807.5 ;
      RECT  9505.0 4957.5 10062.5 5022.5 ;
      RECT  10510.0 642.5 10575.0 707.5 ;
      RECT  10510.0 630.0 10575.0 695.0 ;
      RECT  10292.5 642.5 10542.5 707.5 ;
      RECT  10510.0 662.5 10575.0 675.0 ;
      RECT  10542.5 630.0 10790.0 695.0 ;
      RECT  10510.0 2052.5 10575.0 2117.5 ;
      RECT  10510.0 2065.0 10575.0 2130.0 ;
      RECT  10292.5 2052.5 10542.5 2117.5 ;
      RECT  10510.0 2085.0 10575.0 2097.5 ;
      RECT  10542.5 2065.0 10790.0 2130.0 ;
      RECT  10510.0 3332.5 10575.0 3397.5 ;
      RECT  10510.0 3320.0 10575.0 3385.0 ;
      RECT  10292.5 3332.5 10542.5 3397.5 ;
      RECT  10510.0 3352.5 10575.0 3365.0 ;
      RECT  10542.5 3320.0 10790.0 3385.0 ;
      RECT  10510.0 4742.5 10575.0 4807.5 ;
      RECT  10510.0 4755.0 10575.0 4820.0 ;
      RECT  10292.5 4742.5 10542.5 4807.5 ;
      RECT  10510.0 4775.0 10575.0 4787.5 ;
      RECT  10542.5 4755.0 10790.0 4820.0 ;
      RECT  8237.5 1195.0 8302.5 1380.0 ;
      RECT  8237.5 35.0 8302.5 220.0 ;
      RECT  7877.5 152.5 7942.5 2.5 ;
      RECT  7877.5 1037.5 7942.5 1412.5 ;
      RECT  8067.5 152.5 8132.5 1037.5 ;
      RECT  7877.5 1037.5 7942.5 1172.5 ;
      RECT  8067.5 1037.5 8132.5 1172.5 ;
      RECT  8067.5 1037.5 8132.5 1172.5 ;
      RECT  7877.5 1037.5 7942.5 1172.5 ;
      RECT  7877.5 152.5 7942.5 287.5 ;
      RECT  8067.5 152.5 8132.5 287.5 ;
      RECT  8067.5 152.5 8132.5 287.5 ;
      RECT  7877.5 152.5 7942.5 287.5 ;
      RECT  8237.5 1127.5 8302.5 1262.5 ;
      RECT  8237.5 152.5 8302.5 287.5 ;
      RECT  7935.0 595.0 8000.0 730.0 ;
      RECT  7935.0 595.0 8000.0 730.0 ;
      RECT  8100.0 630.0 8165.0 695.0 ;
      RECT  7810.0 1347.5 8370.0 1412.5 ;
      RECT  7810.0 2.5 8370.0 67.5 ;
      RECT  8237.5 1565.0 8302.5 1380.0 ;
      RECT  8237.5 2725.0 8302.5 2540.0 ;
      RECT  7877.5 2607.5 7942.5 2757.5 ;
      RECT  7877.5 1722.5 7942.5 1347.5 ;
      RECT  8067.5 2607.5 8132.5 1722.5 ;
      RECT  7877.5 1722.5 7942.5 1587.5 ;
      RECT  8067.5 1722.5 8132.5 1587.5 ;
      RECT  8067.5 1722.5 8132.5 1587.5 ;
      RECT  7877.5 1722.5 7942.5 1587.5 ;
      RECT  7877.5 2607.5 7942.5 2472.5 ;
      RECT  8067.5 2607.5 8132.5 2472.5 ;
      RECT  8067.5 2607.5 8132.5 2472.5 ;
      RECT  7877.5 2607.5 7942.5 2472.5 ;
      RECT  8237.5 1632.5 8302.5 1497.5 ;
      RECT  8237.5 2607.5 8302.5 2472.5 ;
      RECT  7935.0 2165.0 8000.0 2030.0 ;
      RECT  7935.0 2165.0 8000.0 2030.0 ;
      RECT  8100.0 2130.0 8165.0 2065.0 ;
      RECT  7810.0 1412.5 8370.0 1347.5 ;
      RECT  7810.0 2757.5 8370.0 2692.5 ;
      RECT  11092.5 1195.0 11157.5 1380.0 ;
      RECT  11092.5 35.0 11157.5 220.0 ;
      RECT  10732.5 152.5 10797.5 2.5 ;
      RECT  10732.5 1037.5 10797.5 1412.5 ;
      RECT  10922.5 152.5 10987.5 1037.5 ;
      RECT  10732.5 1037.5 10797.5 1172.5 ;
      RECT  10922.5 1037.5 10987.5 1172.5 ;
      RECT  10922.5 1037.5 10987.5 1172.5 ;
      RECT  10732.5 1037.5 10797.5 1172.5 ;
      RECT  10732.5 152.5 10797.5 287.5 ;
      RECT  10922.5 152.5 10987.5 287.5 ;
      RECT  10922.5 152.5 10987.5 287.5 ;
      RECT  10732.5 152.5 10797.5 287.5 ;
      RECT  11092.5 1127.5 11157.5 1262.5 ;
      RECT  11092.5 152.5 11157.5 287.5 ;
      RECT  10790.0 595.0 10855.0 730.0 ;
      RECT  10790.0 595.0 10855.0 730.0 ;
      RECT  10955.0 630.0 11020.0 695.0 ;
      RECT  10665.0 1347.5 11225.0 1412.5 ;
      RECT  10665.0 2.5 11225.0 67.5 ;
      RECT  11092.5 1565.0 11157.5 1380.0 ;
      RECT  11092.5 2725.0 11157.5 2540.0 ;
      RECT  10732.5 2607.5 10797.5 2757.5 ;
      RECT  10732.5 1722.5 10797.5 1347.5 ;
      RECT  10922.5 2607.5 10987.5 1722.5 ;
      RECT  10732.5 1722.5 10797.5 1587.5 ;
      RECT  10922.5 1722.5 10987.5 1587.5 ;
      RECT  10922.5 1722.5 10987.5 1587.5 ;
      RECT  10732.5 1722.5 10797.5 1587.5 ;
      RECT  10732.5 2607.5 10797.5 2472.5 ;
      RECT  10922.5 2607.5 10987.5 2472.5 ;
      RECT  10922.5 2607.5 10987.5 2472.5 ;
      RECT  10732.5 2607.5 10797.5 2472.5 ;
      RECT  11092.5 1632.5 11157.5 1497.5 ;
      RECT  11092.5 2607.5 11157.5 2472.5 ;
      RECT  10790.0 2165.0 10855.0 2030.0 ;
      RECT  10790.0 2165.0 10855.0 2030.0 ;
      RECT  10955.0 2130.0 11020.0 2065.0 ;
      RECT  10665.0 1412.5 11225.0 1347.5 ;
      RECT  10665.0 2757.5 11225.0 2692.5 ;
      RECT  11092.5 3885.0 11157.5 4070.0 ;
      RECT  11092.5 2725.0 11157.5 2910.0 ;
      RECT  10732.5 2842.5 10797.5 2692.5 ;
      RECT  10732.5 3727.5 10797.5 4102.5 ;
      RECT  10922.5 2842.5 10987.5 3727.5 ;
      RECT  10732.5 3727.5 10797.5 3862.5 ;
      RECT  10922.5 3727.5 10987.5 3862.5 ;
      RECT  10922.5 3727.5 10987.5 3862.5 ;
      RECT  10732.5 3727.5 10797.5 3862.5 ;
      RECT  10732.5 2842.5 10797.5 2977.5 ;
      RECT  10922.5 2842.5 10987.5 2977.5 ;
      RECT  10922.5 2842.5 10987.5 2977.5 ;
      RECT  10732.5 2842.5 10797.5 2977.5 ;
      RECT  11092.5 3817.5 11157.5 3952.5 ;
      RECT  11092.5 2842.5 11157.5 2977.5 ;
      RECT  10790.0 3285.0 10855.0 3420.0 ;
      RECT  10790.0 3285.0 10855.0 3420.0 ;
      RECT  10955.0 3320.0 11020.0 3385.0 ;
      RECT  10665.0 4037.5 11225.0 4102.5 ;
      RECT  10665.0 2692.5 11225.0 2757.5 ;
      RECT  11092.5 4255.0 11157.5 4070.0 ;
      RECT  11092.5 5415.0 11157.5 5230.0 ;
      RECT  10732.5 5297.5 10797.5 5447.5 ;
      RECT  10732.5 4412.5 10797.5 4037.5 ;
      RECT  10922.5 5297.5 10987.5 4412.5 ;
      RECT  10732.5 4412.5 10797.5 4277.5 ;
      RECT  10922.5 4412.5 10987.5 4277.5 ;
      RECT  10922.5 4412.5 10987.5 4277.5 ;
      RECT  10732.5 4412.5 10797.5 4277.5 ;
      RECT  10732.5 5297.5 10797.5 5162.5 ;
      RECT  10922.5 5297.5 10987.5 5162.5 ;
      RECT  10922.5 5297.5 10987.5 5162.5 ;
      RECT  10732.5 5297.5 10797.5 5162.5 ;
      RECT  11092.5 4322.5 11157.5 4187.5 ;
      RECT  11092.5 5297.5 11157.5 5162.5 ;
      RECT  10790.0 4855.0 10855.0 4720.0 ;
      RECT  10790.0 4855.0 10855.0 4720.0 ;
      RECT  10955.0 4820.0 11020.0 4755.0 ;
      RECT  10665.0 4102.5 11225.0 4037.5 ;
      RECT  10665.0 5447.5 11225.0 5382.5 ;
      RECT  9812.5 197.5 9877.5 2.5 ;
      RECT  9812.5 1037.5 9877.5 1412.5 ;
      RECT  10192.5 1037.5 10257.5 1412.5 ;
      RECT  10362.5 1195.0 10427.5 1380.0 ;
      RECT  10362.5 35.0 10427.5 220.0 ;
      RECT  9812.5 1037.5 9877.5 1172.5 ;
      RECT  10002.5 1037.5 10067.5 1172.5 ;
      RECT  10002.5 1037.5 10067.5 1172.5 ;
      RECT  9812.5 1037.5 9877.5 1172.5 ;
      RECT  10002.5 1037.5 10067.5 1172.5 ;
      RECT  10192.5 1037.5 10257.5 1172.5 ;
      RECT  10192.5 1037.5 10257.5 1172.5 ;
      RECT  10002.5 1037.5 10067.5 1172.5 ;
      RECT  9812.5 197.5 9877.5 332.5 ;
      RECT  10002.5 197.5 10067.5 332.5 ;
      RECT  10002.5 197.5 10067.5 332.5 ;
      RECT  9812.5 197.5 9877.5 332.5 ;
      RECT  10002.5 197.5 10067.5 332.5 ;
      RECT  10192.5 197.5 10257.5 332.5 ;
      RECT  10192.5 197.5 10257.5 332.5 ;
      RECT  10002.5 197.5 10067.5 332.5 ;
      RECT  10362.5 1127.5 10427.5 1262.5 ;
      RECT  10362.5 152.5 10427.5 287.5 ;
      RECT  10197.5 427.5 10062.5 492.5 ;
      RECT  9940.0 642.5 9805.0 707.5 ;
      RECT  10002.5 1037.5 10067.5 1172.5 ;
      RECT  10192.5 197.5 10257.5 332.5 ;
      RECT  10292.5 642.5 10157.5 707.5 ;
      RECT  9805.0 642.5 9940.0 707.5 ;
      RECT  10062.5 427.5 10197.5 492.5 ;
      RECT  10157.5 642.5 10292.5 707.5 ;
      RECT  9745.0 1347.5 10665.0 1412.5 ;
      RECT  9745.0 2.5 10665.0 67.5 ;
      RECT  9812.5 2562.5 9877.5 2757.5 ;
      RECT  9812.5 1722.5 9877.5 1347.5 ;
      RECT  10192.5 1722.5 10257.5 1347.5 ;
      RECT  10362.5 1565.0 10427.5 1380.0 ;
      RECT  10362.5 2725.0 10427.5 2540.0 ;
      RECT  9812.5 1722.5 9877.5 1587.5 ;
      RECT  10002.5 1722.5 10067.5 1587.5 ;
      RECT  10002.5 1722.5 10067.5 1587.5 ;
      RECT  9812.5 1722.5 9877.5 1587.5 ;
      RECT  10002.5 1722.5 10067.5 1587.5 ;
      RECT  10192.5 1722.5 10257.5 1587.5 ;
      RECT  10192.5 1722.5 10257.5 1587.5 ;
      RECT  10002.5 1722.5 10067.5 1587.5 ;
      RECT  9812.5 2562.5 9877.5 2427.5 ;
      RECT  10002.5 2562.5 10067.5 2427.5 ;
      RECT  10002.5 2562.5 10067.5 2427.5 ;
      RECT  9812.5 2562.5 9877.5 2427.5 ;
      RECT  10002.5 2562.5 10067.5 2427.5 ;
      RECT  10192.5 2562.5 10257.5 2427.5 ;
      RECT  10192.5 2562.5 10257.5 2427.5 ;
      RECT  10002.5 2562.5 10067.5 2427.5 ;
      RECT  10362.5 1632.5 10427.5 1497.5 ;
      RECT  10362.5 2607.5 10427.5 2472.5 ;
      RECT  10197.5 2332.5 10062.5 2267.5 ;
      RECT  9940.0 2117.5 9805.0 2052.5 ;
      RECT  10002.5 1722.5 10067.5 1587.5 ;
      RECT  10192.5 2562.5 10257.5 2427.5 ;
      RECT  10292.5 2117.5 10157.5 2052.5 ;
      RECT  9805.0 2117.5 9940.0 2052.5 ;
      RECT  10062.5 2332.5 10197.5 2267.5 ;
      RECT  10157.5 2117.5 10292.5 2052.5 ;
      RECT  9745.0 1412.5 10665.0 1347.5 ;
      RECT  9745.0 2757.5 10665.0 2692.5 ;
      RECT  9812.5 2887.5 9877.5 2692.5 ;
      RECT  9812.5 3727.5 9877.5 4102.5 ;
      RECT  10192.5 3727.5 10257.5 4102.5 ;
      RECT  10362.5 3885.0 10427.5 4070.0 ;
      RECT  10362.5 2725.0 10427.5 2910.0 ;
      RECT  9812.5 3727.5 9877.5 3862.5 ;
      RECT  10002.5 3727.5 10067.5 3862.5 ;
      RECT  10002.5 3727.5 10067.5 3862.5 ;
      RECT  9812.5 3727.5 9877.5 3862.5 ;
      RECT  10002.5 3727.5 10067.5 3862.5 ;
      RECT  10192.5 3727.5 10257.5 3862.5 ;
      RECT  10192.5 3727.5 10257.5 3862.5 ;
      RECT  10002.5 3727.5 10067.5 3862.5 ;
      RECT  9812.5 2887.5 9877.5 3022.5 ;
      RECT  10002.5 2887.5 10067.5 3022.5 ;
      RECT  10002.5 2887.5 10067.5 3022.5 ;
      RECT  9812.5 2887.5 9877.5 3022.5 ;
      RECT  10002.5 2887.5 10067.5 3022.5 ;
      RECT  10192.5 2887.5 10257.5 3022.5 ;
      RECT  10192.5 2887.5 10257.5 3022.5 ;
      RECT  10002.5 2887.5 10067.5 3022.5 ;
      RECT  10362.5 3817.5 10427.5 3952.5 ;
      RECT  10362.5 2842.5 10427.5 2977.5 ;
      RECT  10197.5 3117.5 10062.5 3182.5 ;
      RECT  9940.0 3332.5 9805.0 3397.5 ;
      RECT  10002.5 3727.5 10067.5 3862.5 ;
      RECT  10192.5 2887.5 10257.5 3022.5 ;
      RECT  10292.5 3332.5 10157.5 3397.5 ;
      RECT  9805.0 3332.5 9940.0 3397.5 ;
      RECT  10062.5 3117.5 10197.5 3182.5 ;
      RECT  10157.5 3332.5 10292.5 3397.5 ;
      RECT  9745.0 4037.5 10665.0 4102.5 ;
      RECT  9745.0 2692.5 10665.0 2757.5 ;
      RECT  9812.5 5252.5 9877.5 5447.5 ;
      RECT  9812.5 4412.5 9877.5 4037.5 ;
      RECT  10192.5 4412.5 10257.5 4037.5 ;
      RECT  10362.5 4255.0 10427.5 4070.0 ;
      RECT  10362.5 5415.0 10427.5 5230.0 ;
      RECT  9812.5 4412.5 9877.5 4277.5 ;
      RECT  10002.5 4412.5 10067.5 4277.5 ;
      RECT  10002.5 4412.5 10067.5 4277.5 ;
      RECT  9812.5 4412.5 9877.5 4277.5 ;
      RECT  10002.5 4412.5 10067.5 4277.5 ;
      RECT  10192.5 4412.5 10257.5 4277.5 ;
      RECT  10192.5 4412.5 10257.5 4277.5 ;
      RECT  10002.5 4412.5 10067.5 4277.5 ;
      RECT  9812.5 5252.5 9877.5 5117.5 ;
      RECT  10002.5 5252.5 10067.5 5117.5 ;
      RECT  10002.5 5252.5 10067.5 5117.5 ;
      RECT  9812.5 5252.5 9877.5 5117.5 ;
      RECT  10002.5 5252.5 10067.5 5117.5 ;
      RECT  10192.5 5252.5 10257.5 5117.5 ;
      RECT  10192.5 5252.5 10257.5 5117.5 ;
      RECT  10002.5 5252.5 10067.5 5117.5 ;
      RECT  10362.5 4322.5 10427.5 4187.5 ;
      RECT  10362.5 5297.5 10427.5 5162.5 ;
      RECT  10197.5 5022.5 10062.5 4957.5 ;
      RECT  9940.0 4807.5 9805.0 4742.5 ;
      RECT  10002.5 4412.5 10067.5 4277.5 ;
      RECT  10192.5 5252.5 10257.5 5117.5 ;
      RECT  10292.5 4807.5 10157.5 4742.5 ;
      RECT  9805.0 4807.5 9940.0 4742.5 ;
      RECT  10062.5 5022.5 10197.5 4957.5 ;
      RECT  10157.5 4807.5 10292.5 4742.5 ;
      RECT  9745.0 4102.5 10665.0 4037.5 ;
      RECT  9745.0 5447.5 10665.0 5382.5 ;
      RECT  8747.5 1152.5 8612.5 1217.5 ;
      RECT  7362.5 630.0 7227.5 695.0 ;
      RECT  9022.5 2497.5 8887.5 2562.5 ;
      RECT  7637.5 2065.0 7502.5 2130.0 ;
      RECT  7362.5 2827.5 7227.5 2892.5 ;
      RECT  9297.5 2827.5 9162.5 2892.5 ;
      RECT  7637.5 4172.5 7502.5 4237.5 ;
      RECT  9572.5 4172.5 9437.5 4237.5 ;
      RECT  8747.5 642.5 8612.5 707.5 ;
      RECT  9022.5 427.5 8887.5 492.5 ;
      RECT  9297.5 2052.5 9162.5 2117.5 ;
      RECT  9022.5 2267.5 8887.5 2332.5 ;
      RECT  8747.5 3332.5 8612.5 3397.5 ;
      RECT  9572.5 3117.5 9437.5 3182.5 ;
      RECT  9297.5 4742.5 9162.5 4807.5 ;
      RECT  9572.5 4957.5 9437.5 5022.5 ;
      RECT  11020.0 630.0 11225.0 695.0 ;
      RECT  11020.0 2065.0 11225.0 2130.0 ;
      RECT  11020.0 3320.0 11225.0 3385.0 ;
      RECT  11020.0 4755.0 11225.0 4820.0 ;
      RECT  7260.0 1347.5 11225.0 1412.5 ;
      RECT  7260.0 4037.5 11225.0 4102.5 ;
      RECT  7260.0 2.5 11225.0 67.5 ;
      RECT  7260.0 2692.5 11225.0 2757.5 ;
      RECT  7260.0 5382.5 11225.0 5447.5 ;
      RECT  16085.0 19580.0 16790.0 24465.0 ;
      RECT  18905.0 19580.0 19610.0 24465.0 ;
      RECT  16085.0 19697.5 21725.0 19762.5 ;
      RECT  16085.0 24270.0 21725.0 24335.0 ;
      RECT  16085.0 19827.5 21725.0 19892.5 ;
      RECT  16085.0 15405.0 16790.0 19580.0 ;
      RECT  18905.0 15405.0 19610.0 19580.0 ;
      RECT  16085.0 15672.5 21725.0 15737.5 ;
      RECT  16085.0 15802.5 21725.0 15867.5 ;
      RECT  16085.0 16605.0 21725.0 16670.0 ;
      RECT  16085.0 8965.0 16790.0 15405.0 ;
      RECT  18905.0 8965.0 19610.0 15405.0 ;
      RECT  16085.0 9170.0 21725.0 9235.0 ;
      RECT  16085.0 12175.0 21725.0 12240.0 ;
      RECT  16085.0 15135.0 21725.0 15200.0 ;
      RECT  16085.0 10185.0 21725.0 10250.0 ;
      RECT  16085.0 13145.0 21725.0 13210.0 ;
      RECT  16085.0 9330.0 21725.0 9395.0 ;
      RECT  16085.0 8965.0 16790.0 5990.0 ;
      RECT  18905.0 8965.0 19610.0 5990.0 ;
      RECT  16085.0 8597.5 19610.0 8532.5 ;
      RECT  16085.0 7050.0 19610.0 6985.0 ;
      RECT  16085.0 7180.0 19610.0 7115.0 ;
      RECT  16085.0 8467.5 19610.0 8402.5 ;
      RECT  7520.0 27917.5 7585.0 27982.5 ;
      RECT  7520.0 27905.0 7585.0 27970.0 ;
      RECT  7302.5 27917.5 7552.5 27982.5 ;
      RECT  7520.0 27937.5 7585.0 27950.0 ;
      RECT  7552.5 27905.0 7800.0 27970.0 ;
      RECT  7520.0 29327.5 7585.0 29392.5 ;
      RECT  7520.0 29340.0 7585.0 29405.0 ;
      RECT  7302.5 29327.5 7552.5 29392.5 ;
      RECT  7520.0 29360.0 7585.0 29372.5 ;
      RECT  7552.5 29340.0 7800.0 29405.0 ;
      RECT  7520.0 30607.5 7585.0 30672.5 ;
      RECT  7520.0 30595.0 7585.0 30660.0 ;
      RECT  7302.5 30607.5 7552.5 30672.5 ;
      RECT  7520.0 30627.5 7585.0 30640.0 ;
      RECT  7552.5 30595.0 7800.0 30660.0 ;
      RECT  7520.0 32017.5 7585.0 32082.5 ;
      RECT  7520.0 32030.0 7585.0 32095.0 ;
      RECT  7302.5 32017.5 7552.5 32082.5 ;
      RECT  7520.0 32050.0 7585.0 32062.5 ;
      RECT  7552.5 32030.0 7800.0 32095.0 ;
      RECT  7520.0 33297.5 7585.0 33362.5 ;
      RECT  7520.0 33285.0 7585.0 33350.0 ;
      RECT  7302.5 33297.5 7552.5 33362.5 ;
      RECT  7520.0 33317.5 7585.0 33330.0 ;
      RECT  7552.5 33285.0 7800.0 33350.0 ;
      RECT  7520.0 34707.5 7585.0 34772.5 ;
      RECT  7520.0 34720.0 7585.0 34785.0 ;
      RECT  7302.5 34707.5 7552.5 34772.5 ;
      RECT  7520.0 34740.0 7585.0 34752.5 ;
      RECT  7552.5 34720.0 7800.0 34785.0 ;
      RECT  7520.0 35987.5 7585.0 36052.5 ;
      RECT  7520.0 35975.0 7585.0 36040.0 ;
      RECT  7302.5 35987.5 7552.5 36052.5 ;
      RECT  7520.0 36007.5 7585.0 36020.0 ;
      RECT  7552.5 35975.0 7800.0 36040.0 ;
      RECT  7520.0 37397.5 7585.0 37462.5 ;
      RECT  7520.0 37410.0 7585.0 37475.0 ;
      RECT  7302.5 37397.5 7552.5 37462.5 ;
      RECT  7520.0 37430.0 7585.0 37442.5 ;
      RECT  7552.5 37410.0 7800.0 37475.0 ;
      RECT  7520.0 38677.5 7585.0 38742.5 ;
      RECT  7520.0 38665.0 7585.0 38730.0 ;
      RECT  7302.5 38677.5 7552.5 38742.5 ;
      RECT  7520.0 38697.5 7585.0 38710.0 ;
      RECT  7552.5 38665.0 7800.0 38730.0 ;
      RECT  7520.0 40087.5 7585.0 40152.5 ;
      RECT  7520.0 40100.0 7585.0 40165.0 ;
      RECT  7302.5 40087.5 7552.5 40152.5 ;
      RECT  7520.0 40120.0 7585.0 40132.5 ;
      RECT  7552.5 40100.0 7800.0 40165.0 ;
      RECT  7520.0 41367.5 7585.0 41432.5 ;
      RECT  7520.0 41355.0 7585.0 41420.0 ;
      RECT  7302.5 41367.5 7552.5 41432.5 ;
      RECT  7520.0 41387.5 7585.0 41400.0 ;
      RECT  7552.5 41355.0 7800.0 41420.0 ;
      RECT  7520.0 42777.5 7585.0 42842.5 ;
      RECT  7520.0 42790.0 7585.0 42855.0 ;
      RECT  7302.5 42777.5 7552.5 42842.5 ;
      RECT  7520.0 42810.0 7585.0 42822.5 ;
      RECT  7552.5 42790.0 7800.0 42855.0 ;
      RECT  7520.0 44057.5 7585.0 44122.5 ;
      RECT  7520.0 44045.0 7585.0 44110.0 ;
      RECT  7302.5 44057.5 7552.5 44122.5 ;
      RECT  7520.0 44077.5 7585.0 44090.0 ;
      RECT  7552.5 44045.0 7800.0 44110.0 ;
      RECT  7520.0 45467.5 7585.0 45532.5 ;
      RECT  7520.0 45480.0 7585.0 45545.0 ;
      RECT  7302.5 45467.5 7552.5 45532.5 ;
      RECT  7520.0 45500.0 7585.0 45512.5 ;
      RECT  7552.5 45480.0 7800.0 45545.0 ;
      RECT  7520.0 46747.5 7585.0 46812.5 ;
      RECT  7520.0 46735.0 7585.0 46800.0 ;
      RECT  7302.5 46747.5 7552.5 46812.5 ;
      RECT  7520.0 46767.5 7585.0 46780.0 ;
      RECT  7552.5 46735.0 7800.0 46800.0 ;
      RECT  7520.0 48157.5 7585.0 48222.5 ;
      RECT  7520.0 48170.0 7585.0 48235.0 ;
      RECT  7302.5 48157.5 7552.5 48222.5 ;
      RECT  7520.0 48190.0 7585.0 48202.5 ;
      RECT  7552.5 48170.0 7800.0 48235.0 ;
      RECT  7520.0 49437.5 7585.0 49502.5 ;
      RECT  7520.0 49425.0 7585.0 49490.0 ;
      RECT  7302.5 49437.5 7552.5 49502.5 ;
      RECT  7520.0 49457.5 7585.0 49470.0 ;
      RECT  7552.5 49425.0 7800.0 49490.0 ;
      RECT  7520.0 50847.5 7585.0 50912.5 ;
      RECT  7520.0 50860.0 7585.0 50925.0 ;
      RECT  7302.5 50847.5 7552.5 50912.5 ;
      RECT  7520.0 50880.0 7585.0 50892.5 ;
      RECT  7552.5 50860.0 7800.0 50925.0 ;
      RECT  7520.0 52127.5 7585.0 52192.5 ;
      RECT  7520.0 52115.0 7585.0 52180.0 ;
      RECT  7302.5 52127.5 7552.5 52192.5 ;
      RECT  7520.0 52147.5 7585.0 52160.0 ;
      RECT  7552.5 52115.0 7800.0 52180.0 ;
      RECT  7520.0 53537.5 7585.0 53602.5 ;
      RECT  7520.0 53550.0 7585.0 53615.0 ;
      RECT  7302.5 53537.5 7552.5 53602.5 ;
      RECT  7520.0 53570.0 7585.0 53582.5 ;
      RECT  7552.5 53550.0 7800.0 53615.0 ;
      RECT  7520.0 54817.5 7585.0 54882.5 ;
      RECT  7520.0 54805.0 7585.0 54870.0 ;
      RECT  7302.5 54817.5 7552.5 54882.5 ;
      RECT  7520.0 54837.5 7585.0 54850.0 ;
      RECT  7552.5 54805.0 7800.0 54870.0 ;
      RECT  7520.0 56227.5 7585.0 56292.5 ;
      RECT  7520.0 56240.0 7585.0 56305.0 ;
      RECT  7302.5 56227.5 7552.5 56292.5 ;
      RECT  7520.0 56260.0 7585.0 56272.5 ;
      RECT  7552.5 56240.0 7800.0 56305.0 ;
      RECT  7520.0 57507.5 7585.0 57572.5 ;
      RECT  7520.0 57495.0 7585.0 57560.0 ;
      RECT  7302.5 57507.5 7552.5 57572.5 ;
      RECT  7520.0 57527.5 7585.0 57540.0 ;
      RECT  7552.5 57495.0 7800.0 57560.0 ;
      RECT  7520.0 58917.5 7585.0 58982.5 ;
      RECT  7520.0 58930.0 7585.0 58995.0 ;
      RECT  7302.5 58917.5 7552.5 58982.5 ;
      RECT  7520.0 58950.0 7585.0 58962.5 ;
      RECT  7552.5 58930.0 7800.0 58995.0 ;
      RECT  7520.0 60197.5 7585.0 60262.5 ;
      RECT  7520.0 60185.0 7585.0 60250.0 ;
      RECT  7302.5 60197.5 7552.5 60262.5 ;
      RECT  7520.0 60217.5 7585.0 60230.0 ;
      RECT  7552.5 60185.0 7800.0 60250.0 ;
      RECT  7520.0 61607.5 7585.0 61672.5 ;
      RECT  7520.0 61620.0 7585.0 61685.0 ;
      RECT  7302.5 61607.5 7552.5 61672.5 ;
      RECT  7520.0 61640.0 7585.0 61652.5 ;
      RECT  7552.5 61620.0 7800.0 61685.0 ;
      RECT  7520.0 62887.5 7585.0 62952.5 ;
      RECT  7520.0 62875.0 7585.0 62940.0 ;
      RECT  7302.5 62887.5 7552.5 62952.5 ;
      RECT  7520.0 62907.5 7585.0 62920.0 ;
      RECT  7552.5 62875.0 7800.0 62940.0 ;
      RECT  7520.0 64297.5 7585.0 64362.5 ;
      RECT  7520.0 64310.0 7585.0 64375.0 ;
      RECT  7302.5 64297.5 7552.5 64362.5 ;
      RECT  7520.0 64330.0 7585.0 64342.5 ;
      RECT  7552.5 64310.0 7800.0 64375.0 ;
      RECT  7520.0 65577.5 7585.0 65642.5 ;
      RECT  7520.0 65565.0 7585.0 65630.0 ;
      RECT  7302.5 65577.5 7552.5 65642.5 ;
      RECT  7520.0 65597.5 7585.0 65610.0 ;
      RECT  7552.5 65565.0 7800.0 65630.0 ;
      RECT  7520.0 66987.5 7585.0 67052.5 ;
      RECT  7520.0 67000.0 7585.0 67065.0 ;
      RECT  7302.5 66987.5 7552.5 67052.5 ;
      RECT  7520.0 67020.0 7585.0 67032.5 ;
      RECT  7552.5 67000.0 7800.0 67065.0 ;
      RECT  7520.0 68267.5 7585.0 68332.5 ;
      RECT  7520.0 68255.0 7585.0 68320.0 ;
      RECT  7302.5 68267.5 7552.5 68332.5 ;
      RECT  7520.0 68287.5 7585.0 68300.0 ;
      RECT  7552.5 68255.0 7800.0 68320.0 ;
      RECT  7520.0 69677.5 7585.0 69742.5 ;
      RECT  7520.0 69690.0 7585.0 69755.0 ;
      RECT  7302.5 69677.5 7552.5 69742.5 ;
      RECT  7520.0 69710.0 7585.0 69722.5 ;
      RECT  7552.5 69690.0 7800.0 69755.0 ;
      RECT  4690.0 11765.0 6755.0 11830.0 ;
      RECT  4865.0 13200.0 6755.0 13265.0 ;
      RECT  5040.0 14455.0 6755.0 14520.0 ;
      RECT  5215.0 15890.0 6755.0 15955.0 ;
      RECT  5390.0 17145.0 6755.0 17210.0 ;
      RECT  5565.0 18580.0 6755.0 18645.0 ;
      RECT  5740.0 19835.0 6755.0 19900.0 ;
      RECT  5915.0 21270.0 6755.0 21335.0 ;
      RECT  6090.0 22525.0 6755.0 22590.0 ;
      RECT  6265.0 23960.0 6755.0 24025.0 ;
      RECT  6440.0 25215.0 6755.0 25280.0 ;
      RECT  6615.0 26650.0 6755.0 26715.0 ;
      RECT  4690.0 27917.5 6815.0 27982.5 ;
      RECT  5390.0 27702.5 7072.5 27767.5 ;
      RECT  4690.0 29327.5 6815.0 29392.5 ;
      RECT  5565.0 29542.5 7072.5 29607.5 ;
      RECT  4690.0 30607.5 6815.0 30672.5 ;
      RECT  5740.0 30392.5 7072.5 30457.5 ;
      RECT  4690.0 32017.5 6815.0 32082.5 ;
      RECT  5915.0 32232.5 7072.5 32297.5 ;
      RECT  4690.0 33297.5 6815.0 33362.5 ;
      RECT  6090.0 33082.5 7072.5 33147.5 ;
      RECT  4690.0 34707.5 6815.0 34772.5 ;
      RECT  6265.0 34922.5 7072.5 34987.5 ;
      RECT  4690.0 35987.5 6815.0 36052.5 ;
      RECT  6440.0 35772.5 7072.5 35837.5 ;
      RECT  4690.0 37397.5 6815.0 37462.5 ;
      RECT  6615.0 37612.5 7072.5 37677.5 ;
      RECT  4865.0 38677.5 6815.0 38742.5 ;
      RECT  5390.0 38462.5 7072.5 38527.5 ;
      RECT  4865.0 40087.5 6815.0 40152.5 ;
      RECT  5565.0 40302.5 7072.5 40367.5 ;
      RECT  4865.0 41367.5 6815.0 41432.5 ;
      RECT  5740.0 41152.5 7072.5 41217.5 ;
      RECT  4865.0 42777.5 6815.0 42842.5 ;
      RECT  5915.0 42992.5 7072.5 43057.5 ;
      RECT  4865.0 44057.5 6815.0 44122.5 ;
      RECT  6090.0 43842.5 7072.5 43907.5 ;
      RECT  4865.0 45467.5 6815.0 45532.5 ;
      RECT  6265.0 45682.5 7072.5 45747.5 ;
      RECT  4865.0 46747.5 6815.0 46812.5 ;
      RECT  6440.0 46532.5 7072.5 46597.5 ;
      RECT  4865.0 48157.5 6815.0 48222.5 ;
      RECT  6615.0 48372.5 7072.5 48437.5 ;
      RECT  5040.0 49437.5 6815.0 49502.5 ;
      RECT  5390.0 49222.5 7072.5 49287.5 ;
      RECT  5040.0 50847.5 6815.0 50912.5 ;
      RECT  5565.0 51062.5 7072.5 51127.5 ;
      RECT  5040.0 52127.5 6815.0 52192.5 ;
      RECT  5740.0 51912.5 7072.5 51977.5 ;
      RECT  5040.0 53537.5 6815.0 53602.5 ;
      RECT  5915.0 53752.5 7072.5 53817.5 ;
      RECT  5040.0 54817.5 6815.0 54882.5 ;
      RECT  6090.0 54602.5 7072.5 54667.5 ;
      RECT  5040.0 56227.5 6815.0 56292.5 ;
      RECT  6265.0 56442.5 7072.5 56507.5 ;
      RECT  5040.0 57507.5 6815.0 57572.5 ;
      RECT  6440.0 57292.5 7072.5 57357.5 ;
      RECT  5040.0 58917.5 6815.0 58982.5 ;
      RECT  6615.0 59132.5 7072.5 59197.5 ;
      RECT  5215.0 60197.5 6815.0 60262.5 ;
      RECT  5390.0 59982.5 7072.5 60047.5 ;
      RECT  5215.0 61607.5 6815.0 61672.5 ;
      RECT  5565.0 61822.5 7072.5 61887.5 ;
      RECT  5215.0 62887.5 6815.0 62952.5 ;
      RECT  5740.0 62672.5 7072.5 62737.5 ;
      RECT  5215.0 64297.5 6815.0 64362.5 ;
      RECT  5915.0 64512.5 7072.5 64577.5 ;
      RECT  5215.0 65577.5 6815.0 65642.5 ;
      RECT  6090.0 65362.5 7072.5 65427.5 ;
      RECT  5215.0 66987.5 6815.0 67052.5 ;
      RECT  6265.0 67202.5 7072.5 67267.5 ;
      RECT  5215.0 68267.5 6815.0 68332.5 ;
      RECT  6440.0 68052.5 7072.5 68117.5 ;
      RECT  5215.0 69677.5 6815.0 69742.5 ;
      RECT  6615.0 69892.5 7072.5 69957.5 ;
      RECT  9577.5 11765.0 9512.5 11830.0 ;
      RECT  9577.5 12287.5 9512.5 12352.5 ;
      RECT  9815.0 11765.0 9545.0 11830.0 ;
      RECT  9577.5 11797.5 9512.5 12320.0 ;
      RECT  9545.0 12287.5 9300.0 12352.5 ;
      RECT  10685.0 11765.0 10045.0 11830.0 ;
      RECT  9577.5 13200.0 9512.5 13265.0 ;
      RECT  9577.5 13632.5 9512.5 13697.5 ;
      RECT  9815.0 13200.0 9545.0 13265.0 ;
      RECT  9577.5 13232.5 9512.5 13665.0 ;
      RECT  9545.0 13632.5 9025.0 13697.5 ;
      RECT  10410.0 13200.0 10045.0 13265.0 ;
      RECT  10685.0 13962.5 8750.0 14027.5 ;
      RECT  10410.0 15307.5 8475.0 15372.5 ;
      RECT  9300.0 11777.5 8175.0 11842.5 ;
      RECT  9025.0 11562.5 7917.5 11627.5 ;
      RECT  8750.0 13187.5 8175.0 13252.5 ;
      RECT  9025.0 13402.5 7917.5 13467.5 ;
      RECT  9300.0 14467.5 8175.0 14532.5 ;
      RECT  8475.0 14252.5 7917.5 14317.5 ;
      RECT  8750.0 15877.5 8175.0 15942.5 ;
      RECT  8475.0 16092.5 7917.5 16157.5 ;
      RECT  7470.0 11777.5 7405.0 11842.5 ;
      RECT  7470.0 11765.0 7405.0 11830.0 ;
      RECT  7687.5 11777.5 7437.5 11842.5 ;
      RECT  7470.0 11797.5 7405.0 11810.0 ;
      RECT  7437.5 11765.0 7190.0 11830.0 ;
      RECT  7470.0 13187.5 7405.0 13252.5 ;
      RECT  7470.0 13200.0 7405.0 13265.0 ;
      RECT  7687.5 13187.5 7437.5 13252.5 ;
      RECT  7470.0 13220.0 7405.0 13232.5 ;
      RECT  7437.5 13200.0 7190.0 13265.0 ;
      RECT  7470.0 14467.5 7405.0 14532.5 ;
      RECT  7470.0 14455.0 7405.0 14520.0 ;
      RECT  7687.5 14467.5 7437.5 14532.5 ;
      RECT  7470.0 14487.5 7405.0 14500.0 ;
      RECT  7437.5 14455.0 7190.0 14520.0 ;
      RECT  7470.0 15877.5 7405.0 15942.5 ;
      RECT  7470.0 15890.0 7405.0 15955.0 ;
      RECT  7687.5 15877.5 7437.5 15942.5 ;
      RECT  7470.0 15910.0 7405.0 15922.5 ;
      RECT  7437.5 15890.0 7190.0 15955.0 ;
      RECT  9742.5 12330.0 9677.5 12515.0 ;
      RECT  9742.5 11170.0 9677.5 11355.0 ;
      RECT  10102.5 11287.5 10037.5 11137.5 ;
      RECT  10102.5 12172.5 10037.5 12547.5 ;
      RECT  9912.5 11287.5 9847.5 12172.5 ;
      RECT  10102.5 12172.5 10037.5 12307.5 ;
      RECT  9912.5 12172.5 9847.5 12307.5 ;
      RECT  9912.5 12172.5 9847.5 12307.5 ;
      RECT  10102.5 12172.5 10037.5 12307.5 ;
      RECT  10102.5 11287.5 10037.5 11422.5 ;
      RECT  9912.5 11287.5 9847.5 11422.5 ;
      RECT  9912.5 11287.5 9847.5 11422.5 ;
      RECT  10102.5 11287.5 10037.5 11422.5 ;
      RECT  9742.5 12262.5 9677.5 12397.5 ;
      RECT  9742.5 11287.5 9677.5 11422.5 ;
      RECT  10045.0 11730.0 9980.0 11865.0 ;
      RECT  10045.0 11730.0 9980.0 11865.0 ;
      RECT  9880.0 11765.0 9815.0 11830.0 ;
      RECT  10170.0 12482.5 9610.0 12547.5 ;
      RECT  10170.0 11137.5 9610.0 11202.5 ;
      RECT  9742.5 12700.0 9677.5 12515.0 ;
      RECT  9742.5 13860.0 9677.5 13675.0 ;
      RECT  10102.5 13742.5 10037.5 13892.5 ;
      RECT  10102.5 12857.5 10037.5 12482.5 ;
      RECT  9912.5 13742.5 9847.5 12857.5 ;
      RECT  10102.5 12857.5 10037.5 12722.5 ;
      RECT  9912.5 12857.5 9847.5 12722.5 ;
      RECT  9912.5 12857.5 9847.5 12722.5 ;
      RECT  10102.5 12857.5 10037.5 12722.5 ;
      RECT  10102.5 13742.5 10037.5 13607.5 ;
      RECT  9912.5 13742.5 9847.5 13607.5 ;
      RECT  9912.5 13742.5 9847.5 13607.5 ;
      RECT  10102.5 13742.5 10037.5 13607.5 ;
      RECT  9742.5 12767.5 9677.5 12632.5 ;
      RECT  9742.5 13742.5 9677.5 13607.5 ;
      RECT  10045.0 13300.0 9980.0 13165.0 ;
      RECT  10045.0 13300.0 9980.0 13165.0 ;
      RECT  9880.0 13265.0 9815.0 13200.0 ;
      RECT  10170.0 12547.5 9610.0 12482.5 ;
      RECT  10170.0 13892.5 9610.0 13827.5 ;
      RECT  6887.5 12330.0 6822.5 12515.0 ;
      RECT  6887.5 11170.0 6822.5 11355.0 ;
      RECT  7247.5 11287.5 7182.5 11137.5 ;
      RECT  7247.5 12172.5 7182.5 12547.5 ;
      RECT  7057.5 11287.5 6992.5 12172.5 ;
      RECT  7247.5 12172.5 7182.5 12307.5 ;
      RECT  7057.5 12172.5 6992.5 12307.5 ;
      RECT  7057.5 12172.5 6992.5 12307.5 ;
      RECT  7247.5 12172.5 7182.5 12307.5 ;
      RECT  7247.5 11287.5 7182.5 11422.5 ;
      RECT  7057.5 11287.5 6992.5 11422.5 ;
      RECT  7057.5 11287.5 6992.5 11422.5 ;
      RECT  7247.5 11287.5 7182.5 11422.5 ;
      RECT  6887.5 12262.5 6822.5 12397.5 ;
      RECT  6887.5 11287.5 6822.5 11422.5 ;
      RECT  7190.0 11730.0 7125.0 11865.0 ;
      RECT  7190.0 11730.0 7125.0 11865.0 ;
      RECT  7025.0 11765.0 6960.0 11830.0 ;
      RECT  7315.0 12482.5 6755.0 12547.5 ;
      RECT  7315.0 11137.5 6755.0 11202.5 ;
      RECT  6887.5 12700.0 6822.5 12515.0 ;
      RECT  6887.5 13860.0 6822.5 13675.0 ;
      RECT  7247.5 13742.5 7182.5 13892.5 ;
      RECT  7247.5 12857.5 7182.5 12482.5 ;
      RECT  7057.5 13742.5 6992.5 12857.5 ;
      RECT  7247.5 12857.5 7182.5 12722.5 ;
      RECT  7057.5 12857.5 6992.5 12722.5 ;
      RECT  7057.5 12857.5 6992.5 12722.5 ;
      RECT  7247.5 12857.5 7182.5 12722.5 ;
      RECT  7247.5 13742.5 7182.5 13607.5 ;
      RECT  7057.5 13742.5 6992.5 13607.5 ;
      RECT  7057.5 13742.5 6992.5 13607.5 ;
      RECT  7247.5 13742.5 7182.5 13607.5 ;
      RECT  6887.5 12767.5 6822.5 12632.5 ;
      RECT  6887.5 13742.5 6822.5 13607.5 ;
      RECT  7190.0 13300.0 7125.0 13165.0 ;
      RECT  7190.0 13300.0 7125.0 13165.0 ;
      RECT  7025.0 13265.0 6960.0 13200.0 ;
      RECT  7315.0 12547.5 6755.0 12482.5 ;
      RECT  7315.0 13892.5 6755.0 13827.5 ;
      RECT  6887.5 15020.0 6822.5 15205.0 ;
      RECT  6887.5 13860.0 6822.5 14045.0 ;
      RECT  7247.5 13977.5 7182.5 13827.5 ;
      RECT  7247.5 14862.5 7182.5 15237.5 ;
      RECT  7057.5 13977.5 6992.5 14862.5 ;
      RECT  7247.5 14862.5 7182.5 14997.5 ;
      RECT  7057.5 14862.5 6992.5 14997.5 ;
      RECT  7057.5 14862.5 6992.5 14997.5 ;
      RECT  7247.5 14862.5 7182.5 14997.5 ;
      RECT  7247.5 13977.5 7182.5 14112.5 ;
      RECT  7057.5 13977.5 6992.5 14112.5 ;
      RECT  7057.5 13977.5 6992.5 14112.5 ;
      RECT  7247.5 13977.5 7182.5 14112.5 ;
      RECT  6887.5 14952.5 6822.5 15087.5 ;
      RECT  6887.5 13977.5 6822.5 14112.5 ;
      RECT  7190.0 14420.0 7125.0 14555.0 ;
      RECT  7190.0 14420.0 7125.0 14555.0 ;
      RECT  7025.0 14455.0 6960.0 14520.0 ;
      RECT  7315.0 15172.5 6755.0 15237.5 ;
      RECT  7315.0 13827.5 6755.0 13892.5 ;
      RECT  6887.5 15390.0 6822.5 15205.0 ;
      RECT  6887.5 16550.0 6822.5 16365.0 ;
      RECT  7247.5 16432.5 7182.5 16582.5 ;
      RECT  7247.5 15547.5 7182.5 15172.5 ;
      RECT  7057.5 16432.5 6992.5 15547.5 ;
      RECT  7247.5 15547.5 7182.5 15412.5 ;
      RECT  7057.5 15547.5 6992.5 15412.5 ;
      RECT  7057.5 15547.5 6992.5 15412.5 ;
      RECT  7247.5 15547.5 7182.5 15412.5 ;
      RECT  7247.5 16432.5 7182.5 16297.5 ;
      RECT  7057.5 16432.5 6992.5 16297.5 ;
      RECT  7057.5 16432.5 6992.5 16297.5 ;
      RECT  7247.5 16432.5 7182.5 16297.5 ;
      RECT  6887.5 15457.5 6822.5 15322.5 ;
      RECT  6887.5 16432.5 6822.5 16297.5 ;
      RECT  7190.0 15990.0 7125.0 15855.0 ;
      RECT  7190.0 15990.0 7125.0 15855.0 ;
      RECT  7025.0 15955.0 6960.0 15890.0 ;
      RECT  7315.0 15237.5 6755.0 15172.5 ;
      RECT  7315.0 16582.5 6755.0 16517.5 ;
      RECT  8167.5 11332.5 8102.5 11137.5 ;
      RECT  8167.5 12172.5 8102.5 12547.5 ;
      RECT  7787.5 12172.5 7722.5 12547.5 ;
      RECT  7617.5 12330.0 7552.5 12515.0 ;
      RECT  7617.5 11170.0 7552.5 11355.0 ;
      RECT  8167.5 12172.5 8102.5 12307.5 ;
      RECT  7977.5 12172.5 7912.5 12307.5 ;
      RECT  7977.5 12172.5 7912.5 12307.5 ;
      RECT  8167.5 12172.5 8102.5 12307.5 ;
      RECT  7977.5 12172.5 7912.5 12307.5 ;
      RECT  7787.5 12172.5 7722.5 12307.5 ;
      RECT  7787.5 12172.5 7722.5 12307.5 ;
      RECT  7977.5 12172.5 7912.5 12307.5 ;
      RECT  8167.5 11332.5 8102.5 11467.5 ;
      RECT  7977.5 11332.5 7912.5 11467.5 ;
      RECT  7977.5 11332.5 7912.5 11467.5 ;
      RECT  8167.5 11332.5 8102.5 11467.5 ;
      RECT  7977.5 11332.5 7912.5 11467.5 ;
      RECT  7787.5 11332.5 7722.5 11467.5 ;
      RECT  7787.5 11332.5 7722.5 11467.5 ;
      RECT  7977.5 11332.5 7912.5 11467.5 ;
      RECT  7617.5 12262.5 7552.5 12397.5 ;
      RECT  7617.5 11287.5 7552.5 11422.5 ;
      RECT  7782.5 11562.5 7917.5 11627.5 ;
      RECT  8040.0 11777.5 8175.0 11842.5 ;
      RECT  7977.5 12172.5 7912.5 12307.5 ;
      RECT  7787.5 11332.5 7722.5 11467.5 ;
      RECT  7687.5 11777.5 7822.5 11842.5 ;
      RECT  8175.0 11777.5 8040.0 11842.5 ;
      RECT  7917.5 11562.5 7782.5 11627.5 ;
      RECT  7822.5 11777.5 7687.5 11842.5 ;
      RECT  8235.0 12482.5 7315.0 12547.5 ;
      RECT  8235.0 11137.5 7315.0 11202.5 ;
      RECT  8167.5 13697.5 8102.5 13892.5 ;
      RECT  8167.5 12857.5 8102.5 12482.5 ;
      RECT  7787.5 12857.5 7722.5 12482.5 ;
      RECT  7617.5 12700.0 7552.5 12515.0 ;
      RECT  7617.5 13860.0 7552.5 13675.0 ;
      RECT  8167.5 12857.5 8102.5 12722.5 ;
      RECT  7977.5 12857.5 7912.5 12722.5 ;
      RECT  7977.5 12857.5 7912.5 12722.5 ;
      RECT  8167.5 12857.5 8102.5 12722.5 ;
      RECT  7977.5 12857.5 7912.5 12722.5 ;
      RECT  7787.5 12857.5 7722.5 12722.5 ;
      RECT  7787.5 12857.5 7722.5 12722.5 ;
      RECT  7977.5 12857.5 7912.5 12722.5 ;
      RECT  8167.5 13697.5 8102.5 13562.5 ;
      RECT  7977.5 13697.5 7912.5 13562.5 ;
      RECT  7977.5 13697.5 7912.5 13562.5 ;
      RECT  8167.5 13697.5 8102.5 13562.5 ;
      RECT  7977.5 13697.5 7912.5 13562.5 ;
      RECT  7787.5 13697.5 7722.5 13562.5 ;
      RECT  7787.5 13697.5 7722.5 13562.5 ;
      RECT  7977.5 13697.5 7912.5 13562.5 ;
      RECT  7617.5 12767.5 7552.5 12632.5 ;
      RECT  7617.5 13742.5 7552.5 13607.5 ;
      RECT  7782.5 13467.5 7917.5 13402.5 ;
      RECT  8040.0 13252.5 8175.0 13187.5 ;
      RECT  7977.5 12857.5 7912.5 12722.5 ;
      RECT  7787.5 13697.5 7722.5 13562.5 ;
      RECT  7687.5 13252.5 7822.5 13187.5 ;
      RECT  8175.0 13252.5 8040.0 13187.5 ;
      RECT  7917.5 13467.5 7782.5 13402.5 ;
      RECT  7822.5 13252.5 7687.5 13187.5 ;
      RECT  8235.0 12547.5 7315.0 12482.5 ;
      RECT  8235.0 13892.5 7315.0 13827.5 ;
      RECT  8167.5 14022.5 8102.5 13827.5 ;
      RECT  8167.5 14862.5 8102.5 15237.5 ;
      RECT  7787.5 14862.5 7722.5 15237.5 ;
      RECT  7617.5 15020.0 7552.5 15205.0 ;
      RECT  7617.5 13860.0 7552.5 14045.0 ;
      RECT  8167.5 14862.5 8102.5 14997.5 ;
      RECT  7977.5 14862.5 7912.5 14997.5 ;
      RECT  7977.5 14862.5 7912.5 14997.5 ;
      RECT  8167.5 14862.5 8102.5 14997.5 ;
      RECT  7977.5 14862.5 7912.5 14997.5 ;
      RECT  7787.5 14862.5 7722.5 14997.5 ;
      RECT  7787.5 14862.5 7722.5 14997.5 ;
      RECT  7977.5 14862.5 7912.5 14997.5 ;
      RECT  8167.5 14022.5 8102.5 14157.5 ;
      RECT  7977.5 14022.5 7912.5 14157.5 ;
      RECT  7977.5 14022.5 7912.5 14157.5 ;
      RECT  8167.5 14022.5 8102.5 14157.5 ;
      RECT  7977.5 14022.5 7912.5 14157.5 ;
      RECT  7787.5 14022.5 7722.5 14157.5 ;
      RECT  7787.5 14022.5 7722.5 14157.5 ;
      RECT  7977.5 14022.5 7912.5 14157.5 ;
      RECT  7617.5 14952.5 7552.5 15087.5 ;
      RECT  7617.5 13977.5 7552.5 14112.5 ;
      RECT  7782.5 14252.5 7917.5 14317.5 ;
      RECT  8040.0 14467.5 8175.0 14532.5 ;
      RECT  7977.5 14862.5 7912.5 14997.5 ;
      RECT  7787.5 14022.5 7722.5 14157.5 ;
      RECT  7687.5 14467.5 7822.5 14532.5 ;
      RECT  8175.0 14467.5 8040.0 14532.5 ;
      RECT  7917.5 14252.5 7782.5 14317.5 ;
      RECT  7822.5 14467.5 7687.5 14532.5 ;
      RECT  8235.0 15172.5 7315.0 15237.5 ;
      RECT  8235.0 13827.5 7315.0 13892.5 ;
      RECT  8167.5 16387.5 8102.5 16582.5 ;
      RECT  8167.5 15547.5 8102.5 15172.5 ;
      RECT  7787.5 15547.5 7722.5 15172.5 ;
      RECT  7617.5 15390.0 7552.5 15205.0 ;
      RECT  7617.5 16550.0 7552.5 16365.0 ;
      RECT  8167.5 15547.5 8102.5 15412.5 ;
      RECT  7977.5 15547.5 7912.5 15412.5 ;
      RECT  7977.5 15547.5 7912.5 15412.5 ;
      RECT  8167.5 15547.5 8102.5 15412.5 ;
      RECT  7977.5 15547.5 7912.5 15412.5 ;
      RECT  7787.5 15547.5 7722.5 15412.5 ;
      RECT  7787.5 15547.5 7722.5 15412.5 ;
      RECT  7977.5 15547.5 7912.5 15412.5 ;
      RECT  8167.5 16387.5 8102.5 16252.5 ;
      RECT  7977.5 16387.5 7912.5 16252.5 ;
      RECT  7977.5 16387.5 7912.5 16252.5 ;
      RECT  8167.5 16387.5 8102.5 16252.5 ;
      RECT  7977.5 16387.5 7912.5 16252.5 ;
      RECT  7787.5 16387.5 7722.5 16252.5 ;
      RECT  7787.5 16387.5 7722.5 16252.5 ;
      RECT  7977.5 16387.5 7912.5 16252.5 ;
      RECT  7617.5 15457.5 7552.5 15322.5 ;
      RECT  7617.5 16432.5 7552.5 16297.5 ;
      RECT  7782.5 16157.5 7917.5 16092.5 ;
      RECT  8040.0 15942.5 8175.0 15877.5 ;
      RECT  7977.5 15547.5 7912.5 15412.5 ;
      RECT  7787.5 16387.5 7722.5 16252.5 ;
      RECT  7687.5 15942.5 7822.5 15877.5 ;
      RECT  8175.0 15942.5 8040.0 15877.5 ;
      RECT  7917.5 16157.5 7782.5 16092.5 ;
      RECT  7822.5 15942.5 7687.5 15877.5 ;
      RECT  8235.0 15237.5 7315.0 15172.5 ;
      RECT  8235.0 16582.5 7315.0 16517.5 ;
      RECT  9232.5 12287.5 9367.5 12352.5 ;
      RECT  10617.5 11765.0 10752.5 11830.0 ;
      RECT  8957.5 13632.5 9092.5 13697.5 ;
      RECT  10342.5 13200.0 10477.5 13265.0 ;
      RECT  10617.5 13962.5 10752.5 14027.5 ;
      RECT  8682.5 13962.5 8817.5 14027.5 ;
      RECT  10342.5 15307.5 10477.5 15372.5 ;
      RECT  8407.5 15307.5 8542.5 15372.5 ;
      RECT  9232.5 11777.5 9367.5 11842.5 ;
      RECT  8957.5 11562.5 9092.5 11627.5 ;
      RECT  8682.5 13187.5 8817.5 13252.5 ;
      RECT  8957.5 13402.5 9092.5 13467.5 ;
      RECT  9232.5 14467.5 9367.5 14532.5 ;
      RECT  8407.5 14252.5 8542.5 14317.5 ;
      RECT  8682.5 15877.5 8817.5 15942.5 ;
      RECT  8407.5 16092.5 8542.5 16157.5 ;
      RECT  6960.0 11765.0 6755.0 11830.0 ;
      RECT  6960.0 13200.0 6755.0 13265.0 ;
      RECT  6960.0 14455.0 6755.0 14520.0 ;
      RECT  6960.0 15890.0 6755.0 15955.0 ;
      RECT  10720.0 12482.5 6755.0 12547.5 ;
      RECT  10720.0 15172.5 6755.0 15237.5 ;
      RECT  10720.0 11137.5 6755.0 11202.5 ;
      RECT  10720.0 13827.5 6755.0 13892.5 ;
      RECT  10720.0 16517.5 6755.0 16582.5 ;
      RECT  10217.5 17145.0 10152.5 17210.0 ;
      RECT  10217.5 17667.5 10152.5 17732.5 ;
      RECT  10455.0 17145.0 10185.0 17210.0 ;
      RECT  10217.5 17177.5 10152.5 17700.0 ;
      RECT  10185.0 17667.5 9940.0 17732.5 ;
      RECT  11600.0 17145.0 10685.0 17210.0 ;
      RECT  10217.5 18580.0 10152.5 18645.0 ;
      RECT  10217.5 19012.5 10152.5 19077.5 ;
      RECT  10455.0 18580.0 10185.0 18645.0 ;
      RECT  10217.5 18612.5 10152.5 19045.0 ;
      RECT  10185.0 19012.5 9665.0 19077.5 ;
      RECT  11325.0 18580.0 10685.0 18645.0 ;
      RECT  10217.5 19835.0 10152.5 19900.0 ;
      RECT  10217.5 20357.5 10152.5 20422.5 ;
      RECT  10455.0 19835.0 10185.0 19900.0 ;
      RECT  10217.5 19867.5 10152.5 20390.0 ;
      RECT  10185.0 20357.5 9390.0 20422.5 ;
      RECT  11050.0 19835.0 10685.0 19900.0 ;
      RECT  11600.0 20687.5 9115.0 20752.5 ;
      RECT  11325.0 22032.5 8840.0 22097.5 ;
      RECT  11050.0 23377.5 8565.0 23442.5 ;
      RECT  9940.0 17205.0 8197.5 17270.0 ;
      RECT  9665.0 17065.0 8007.5 17130.0 ;
      RECT  9390.0 16925.0 7817.5 16990.0 ;
      RECT  9115.0 18520.0 8197.5 18585.0 ;
      RECT  9665.0 18660.0 8007.5 18725.0 ;
      RECT  9390.0 18800.0 7817.5 18865.0 ;
      RECT  9940.0 19895.0 8197.5 19960.0 ;
      RECT  8840.0 19755.0 8007.5 19820.0 ;
      RECT  9390.0 19615.0 7817.5 19680.0 ;
      RECT  9115.0 21210.0 8197.5 21275.0 ;
      RECT  8840.0 21350.0 8007.5 21415.0 ;
      RECT  9390.0 21490.0 7817.5 21555.0 ;
      RECT  9940.0 22585.0 8197.5 22650.0 ;
      RECT  9665.0 22445.0 8007.5 22510.0 ;
      RECT  8565.0 22305.0 7817.5 22370.0 ;
      RECT  9115.0 23900.0 8197.5 23965.0 ;
      RECT  9665.0 24040.0 8007.5 24105.0 ;
      RECT  8565.0 24180.0 7817.5 24245.0 ;
      RECT  9940.0 25275.0 8197.5 25340.0 ;
      RECT  8840.0 25135.0 8007.5 25200.0 ;
      RECT  8565.0 24995.0 7817.5 25060.0 ;
      RECT  9115.0 26590.0 8197.5 26655.0 ;
      RECT  8840.0 26730.0 8007.5 26795.0 ;
      RECT  8565.0 26870.0 7817.5 26935.0 ;
      RECT  7437.5 17205.0 7372.5 17270.0 ;
      RECT  7437.5 17145.0 7372.5 17210.0 ;
      RECT  7622.5 17205.0 7405.0 17270.0 ;
      RECT  7437.5 17177.5 7372.5 17237.5 ;
      RECT  7405.0 17145.0 7190.0 17210.0 ;
      RECT  7437.5 18520.0 7372.5 18585.0 ;
      RECT  7437.5 18580.0 7372.5 18645.0 ;
      RECT  7622.5 18520.0 7405.0 18585.0 ;
      RECT  7437.5 18552.5 7372.5 18612.5 ;
      RECT  7405.0 18580.0 7190.0 18645.0 ;
      RECT  7437.5 19895.0 7372.5 19960.0 ;
      RECT  7437.5 19835.0 7372.5 19900.0 ;
      RECT  7622.5 19895.0 7405.0 19960.0 ;
      RECT  7437.5 19867.5 7372.5 19927.5 ;
      RECT  7405.0 19835.0 7190.0 19900.0 ;
      RECT  7437.5 21210.0 7372.5 21275.0 ;
      RECT  7437.5 21270.0 7372.5 21335.0 ;
      RECT  7622.5 21210.0 7405.0 21275.0 ;
      RECT  7437.5 21242.5 7372.5 21302.5 ;
      RECT  7405.0 21270.0 7190.0 21335.0 ;
      RECT  7437.5 22585.0 7372.5 22650.0 ;
      RECT  7437.5 22525.0 7372.5 22590.0 ;
      RECT  7622.5 22585.0 7405.0 22650.0 ;
      RECT  7437.5 22557.5 7372.5 22617.5 ;
      RECT  7405.0 22525.0 7190.0 22590.0 ;
      RECT  7437.5 23900.0 7372.5 23965.0 ;
      RECT  7437.5 23960.0 7372.5 24025.0 ;
      RECT  7622.5 23900.0 7405.0 23965.0 ;
      RECT  7437.5 23932.5 7372.5 23992.5 ;
      RECT  7405.0 23960.0 7190.0 24025.0 ;
      RECT  7437.5 25275.0 7372.5 25340.0 ;
      RECT  7437.5 25215.0 7372.5 25280.0 ;
      RECT  7622.5 25275.0 7405.0 25340.0 ;
      RECT  7437.5 25247.5 7372.5 25307.5 ;
      RECT  7405.0 25215.0 7190.0 25280.0 ;
      RECT  7437.5 26590.0 7372.5 26655.0 ;
      RECT  7437.5 26650.0 7372.5 26715.0 ;
      RECT  7622.5 26590.0 7405.0 26655.0 ;
      RECT  7437.5 26622.5 7372.5 26682.5 ;
      RECT  7405.0 26650.0 7190.0 26715.0 ;
      RECT  10382.5 17710.0 10317.5 17895.0 ;
      RECT  10382.5 16550.0 10317.5 16735.0 ;
      RECT  10742.5 16667.5 10677.5 16517.5 ;
      RECT  10742.5 17552.5 10677.5 17927.5 ;
      RECT  10552.5 16667.5 10487.5 17552.5 ;
      RECT  10742.5 17552.5 10677.5 17687.5 ;
      RECT  10552.5 17552.5 10487.5 17687.5 ;
      RECT  10552.5 17552.5 10487.5 17687.5 ;
      RECT  10742.5 17552.5 10677.5 17687.5 ;
      RECT  10742.5 16667.5 10677.5 16802.5 ;
      RECT  10552.5 16667.5 10487.5 16802.5 ;
      RECT  10552.5 16667.5 10487.5 16802.5 ;
      RECT  10742.5 16667.5 10677.5 16802.5 ;
      RECT  10382.5 17642.5 10317.5 17777.5 ;
      RECT  10382.5 16667.5 10317.5 16802.5 ;
      RECT  10685.0 17110.0 10620.0 17245.0 ;
      RECT  10685.0 17110.0 10620.0 17245.0 ;
      RECT  10520.0 17145.0 10455.0 17210.0 ;
      RECT  10810.0 17862.5 10250.0 17927.5 ;
      RECT  10810.0 16517.5 10250.0 16582.5 ;
      RECT  10382.5 18080.0 10317.5 17895.0 ;
      RECT  10382.5 19240.0 10317.5 19055.0 ;
      RECT  10742.5 19122.5 10677.5 19272.5 ;
      RECT  10742.5 18237.5 10677.5 17862.5 ;
      RECT  10552.5 19122.5 10487.5 18237.5 ;
      RECT  10742.5 18237.5 10677.5 18102.5 ;
      RECT  10552.5 18237.5 10487.5 18102.5 ;
      RECT  10552.5 18237.5 10487.5 18102.5 ;
      RECT  10742.5 18237.5 10677.5 18102.5 ;
      RECT  10742.5 19122.5 10677.5 18987.5 ;
      RECT  10552.5 19122.5 10487.5 18987.5 ;
      RECT  10552.5 19122.5 10487.5 18987.5 ;
      RECT  10742.5 19122.5 10677.5 18987.5 ;
      RECT  10382.5 18147.5 10317.5 18012.5 ;
      RECT  10382.5 19122.5 10317.5 18987.5 ;
      RECT  10685.0 18680.0 10620.0 18545.0 ;
      RECT  10685.0 18680.0 10620.0 18545.0 ;
      RECT  10520.0 18645.0 10455.0 18580.0 ;
      RECT  10810.0 17927.5 10250.0 17862.5 ;
      RECT  10810.0 19272.5 10250.0 19207.5 ;
      RECT  10382.5 20400.0 10317.5 20585.0 ;
      RECT  10382.5 19240.0 10317.5 19425.0 ;
      RECT  10742.5 19357.5 10677.5 19207.5 ;
      RECT  10742.5 20242.5 10677.5 20617.5 ;
      RECT  10552.5 19357.5 10487.5 20242.5 ;
      RECT  10742.5 20242.5 10677.5 20377.5 ;
      RECT  10552.5 20242.5 10487.5 20377.5 ;
      RECT  10552.5 20242.5 10487.5 20377.5 ;
      RECT  10742.5 20242.5 10677.5 20377.5 ;
      RECT  10742.5 19357.5 10677.5 19492.5 ;
      RECT  10552.5 19357.5 10487.5 19492.5 ;
      RECT  10552.5 19357.5 10487.5 19492.5 ;
      RECT  10742.5 19357.5 10677.5 19492.5 ;
      RECT  10382.5 20332.5 10317.5 20467.5 ;
      RECT  10382.5 19357.5 10317.5 19492.5 ;
      RECT  10685.0 19800.0 10620.0 19935.0 ;
      RECT  10685.0 19800.0 10620.0 19935.0 ;
      RECT  10520.0 19835.0 10455.0 19900.0 ;
      RECT  10810.0 20552.5 10250.0 20617.5 ;
      RECT  10810.0 19207.5 10250.0 19272.5 ;
      RECT  6887.5 17710.0 6822.5 17895.0 ;
      RECT  6887.5 16550.0 6822.5 16735.0 ;
      RECT  7247.5 16667.5 7182.5 16517.5 ;
      RECT  7247.5 17552.5 7182.5 17927.5 ;
      RECT  7057.5 16667.5 6992.5 17552.5 ;
      RECT  7247.5 17552.5 7182.5 17687.5 ;
      RECT  7057.5 17552.5 6992.5 17687.5 ;
      RECT  7057.5 17552.5 6992.5 17687.5 ;
      RECT  7247.5 17552.5 7182.5 17687.5 ;
      RECT  7247.5 16667.5 7182.5 16802.5 ;
      RECT  7057.5 16667.5 6992.5 16802.5 ;
      RECT  7057.5 16667.5 6992.5 16802.5 ;
      RECT  7247.5 16667.5 7182.5 16802.5 ;
      RECT  6887.5 17642.5 6822.5 17777.5 ;
      RECT  6887.5 16667.5 6822.5 16802.5 ;
      RECT  7190.0 17110.0 7125.0 17245.0 ;
      RECT  7190.0 17110.0 7125.0 17245.0 ;
      RECT  7025.0 17145.0 6960.0 17210.0 ;
      RECT  7315.0 17862.5 6755.0 17927.5 ;
      RECT  7315.0 16517.5 6755.0 16582.5 ;
      RECT  6887.5 18080.0 6822.5 17895.0 ;
      RECT  6887.5 19240.0 6822.5 19055.0 ;
      RECT  7247.5 19122.5 7182.5 19272.5 ;
      RECT  7247.5 18237.5 7182.5 17862.5 ;
      RECT  7057.5 19122.5 6992.5 18237.5 ;
      RECT  7247.5 18237.5 7182.5 18102.5 ;
      RECT  7057.5 18237.5 6992.5 18102.5 ;
      RECT  7057.5 18237.5 6992.5 18102.5 ;
      RECT  7247.5 18237.5 7182.5 18102.5 ;
      RECT  7247.5 19122.5 7182.5 18987.5 ;
      RECT  7057.5 19122.5 6992.5 18987.5 ;
      RECT  7057.5 19122.5 6992.5 18987.5 ;
      RECT  7247.5 19122.5 7182.5 18987.5 ;
      RECT  6887.5 18147.5 6822.5 18012.5 ;
      RECT  6887.5 19122.5 6822.5 18987.5 ;
      RECT  7190.0 18680.0 7125.0 18545.0 ;
      RECT  7190.0 18680.0 7125.0 18545.0 ;
      RECT  7025.0 18645.0 6960.0 18580.0 ;
      RECT  7315.0 17927.5 6755.0 17862.5 ;
      RECT  7315.0 19272.5 6755.0 19207.5 ;
      RECT  6887.5 20400.0 6822.5 20585.0 ;
      RECT  6887.5 19240.0 6822.5 19425.0 ;
      RECT  7247.5 19357.5 7182.5 19207.5 ;
      RECT  7247.5 20242.5 7182.5 20617.5 ;
      RECT  7057.5 19357.5 6992.5 20242.5 ;
      RECT  7247.5 20242.5 7182.5 20377.5 ;
      RECT  7057.5 20242.5 6992.5 20377.5 ;
      RECT  7057.5 20242.5 6992.5 20377.5 ;
      RECT  7247.5 20242.5 7182.5 20377.5 ;
      RECT  7247.5 19357.5 7182.5 19492.5 ;
      RECT  7057.5 19357.5 6992.5 19492.5 ;
      RECT  7057.5 19357.5 6992.5 19492.5 ;
      RECT  7247.5 19357.5 7182.5 19492.5 ;
      RECT  6887.5 20332.5 6822.5 20467.5 ;
      RECT  6887.5 19357.5 6822.5 19492.5 ;
      RECT  7190.0 19800.0 7125.0 19935.0 ;
      RECT  7190.0 19800.0 7125.0 19935.0 ;
      RECT  7025.0 19835.0 6960.0 19900.0 ;
      RECT  7315.0 20552.5 6755.0 20617.5 ;
      RECT  7315.0 19207.5 6755.0 19272.5 ;
      RECT  6887.5 20770.0 6822.5 20585.0 ;
      RECT  6887.5 21930.0 6822.5 21745.0 ;
      RECT  7247.5 21812.5 7182.5 21962.5 ;
      RECT  7247.5 20927.5 7182.5 20552.5 ;
      RECT  7057.5 21812.5 6992.5 20927.5 ;
      RECT  7247.5 20927.5 7182.5 20792.5 ;
      RECT  7057.5 20927.5 6992.5 20792.5 ;
      RECT  7057.5 20927.5 6992.5 20792.5 ;
      RECT  7247.5 20927.5 7182.5 20792.5 ;
      RECT  7247.5 21812.5 7182.5 21677.5 ;
      RECT  7057.5 21812.5 6992.5 21677.5 ;
      RECT  7057.5 21812.5 6992.5 21677.5 ;
      RECT  7247.5 21812.5 7182.5 21677.5 ;
      RECT  6887.5 20837.5 6822.5 20702.5 ;
      RECT  6887.5 21812.5 6822.5 21677.5 ;
      RECT  7190.0 21370.0 7125.0 21235.0 ;
      RECT  7190.0 21370.0 7125.0 21235.0 ;
      RECT  7025.0 21335.0 6960.0 21270.0 ;
      RECT  7315.0 20617.5 6755.0 20552.5 ;
      RECT  7315.0 21962.5 6755.0 21897.5 ;
      RECT  6887.5 23090.0 6822.5 23275.0 ;
      RECT  6887.5 21930.0 6822.5 22115.0 ;
      RECT  7247.5 22047.5 7182.5 21897.5 ;
      RECT  7247.5 22932.5 7182.5 23307.5 ;
      RECT  7057.5 22047.5 6992.5 22932.5 ;
      RECT  7247.5 22932.5 7182.5 23067.5 ;
      RECT  7057.5 22932.5 6992.5 23067.5 ;
      RECT  7057.5 22932.5 6992.5 23067.5 ;
      RECT  7247.5 22932.5 7182.5 23067.5 ;
      RECT  7247.5 22047.5 7182.5 22182.5 ;
      RECT  7057.5 22047.5 6992.5 22182.5 ;
      RECT  7057.5 22047.5 6992.5 22182.5 ;
      RECT  7247.5 22047.5 7182.5 22182.5 ;
      RECT  6887.5 23022.5 6822.5 23157.5 ;
      RECT  6887.5 22047.5 6822.5 22182.5 ;
      RECT  7190.0 22490.0 7125.0 22625.0 ;
      RECT  7190.0 22490.0 7125.0 22625.0 ;
      RECT  7025.0 22525.0 6960.0 22590.0 ;
      RECT  7315.0 23242.5 6755.0 23307.5 ;
      RECT  7315.0 21897.5 6755.0 21962.5 ;
      RECT  6887.5 23460.0 6822.5 23275.0 ;
      RECT  6887.5 24620.0 6822.5 24435.0 ;
      RECT  7247.5 24502.5 7182.5 24652.5 ;
      RECT  7247.5 23617.5 7182.5 23242.5 ;
      RECT  7057.5 24502.5 6992.5 23617.5 ;
      RECT  7247.5 23617.5 7182.5 23482.5 ;
      RECT  7057.5 23617.5 6992.5 23482.5 ;
      RECT  7057.5 23617.5 6992.5 23482.5 ;
      RECT  7247.5 23617.5 7182.5 23482.5 ;
      RECT  7247.5 24502.5 7182.5 24367.5 ;
      RECT  7057.5 24502.5 6992.5 24367.5 ;
      RECT  7057.5 24502.5 6992.5 24367.5 ;
      RECT  7247.5 24502.5 7182.5 24367.5 ;
      RECT  6887.5 23527.5 6822.5 23392.5 ;
      RECT  6887.5 24502.5 6822.5 24367.5 ;
      RECT  7190.0 24060.0 7125.0 23925.0 ;
      RECT  7190.0 24060.0 7125.0 23925.0 ;
      RECT  7025.0 24025.0 6960.0 23960.0 ;
      RECT  7315.0 23307.5 6755.0 23242.5 ;
      RECT  7315.0 24652.5 6755.0 24587.5 ;
      RECT  6887.5 25780.0 6822.5 25965.0 ;
      RECT  6887.5 24620.0 6822.5 24805.0 ;
      RECT  7247.5 24737.5 7182.5 24587.5 ;
      RECT  7247.5 25622.5 7182.5 25997.5 ;
      RECT  7057.5 24737.5 6992.5 25622.5 ;
      RECT  7247.5 25622.5 7182.5 25757.5 ;
      RECT  7057.5 25622.5 6992.5 25757.5 ;
      RECT  7057.5 25622.5 6992.5 25757.5 ;
      RECT  7247.5 25622.5 7182.5 25757.5 ;
      RECT  7247.5 24737.5 7182.5 24872.5 ;
      RECT  7057.5 24737.5 6992.5 24872.5 ;
      RECT  7057.5 24737.5 6992.5 24872.5 ;
      RECT  7247.5 24737.5 7182.5 24872.5 ;
      RECT  6887.5 25712.5 6822.5 25847.5 ;
      RECT  6887.5 24737.5 6822.5 24872.5 ;
      RECT  7190.0 25180.0 7125.0 25315.0 ;
      RECT  7190.0 25180.0 7125.0 25315.0 ;
      RECT  7025.0 25215.0 6960.0 25280.0 ;
      RECT  7315.0 25932.5 6755.0 25997.5 ;
      RECT  7315.0 24587.5 6755.0 24652.5 ;
      RECT  6887.5 26150.0 6822.5 25965.0 ;
      RECT  6887.5 27310.0 6822.5 27125.0 ;
      RECT  7247.5 27192.5 7182.5 27342.5 ;
      RECT  7247.5 26307.5 7182.5 25932.5 ;
      RECT  7057.5 27192.5 6992.5 26307.5 ;
      RECT  7247.5 26307.5 7182.5 26172.5 ;
      RECT  7057.5 26307.5 6992.5 26172.5 ;
      RECT  7057.5 26307.5 6992.5 26172.5 ;
      RECT  7247.5 26307.5 7182.5 26172.5 ;
      RECT  7247.5 27192.5 7182.5 27057.5 ;
      RECT  7057.5 27192.5 6992.5 27057.5 ;
      RECT  7057.5 27192.5 6992.5 27057.5 ;
      RECT  7247.5 27192.5 7182.5 27057.5 ;
      RECT  6887.5 26217.5 6822.5 26082.5 ;
      RECT  6887.5 27192.5 6822.5 27057.5 ;
      RECT  7190.0 26750.0 7125.0 26615.0 ;
      RECT  7190.0 26750.0 7125.0 26615.0 ;
      RECT  7025.0 26715.0 6960.0 26650.0 ;
      RECT  7315.0 25997.5 6755.0 25932.5 ;
      RECT  7315.0 27342.5 6755.0 27277.5 ;
      RECT  8257.5 16712.5 8192.5 16517.5 ;
      RECT  8257.5 17552.5 8192.5 17927.5 ;
      RECT  7877.5 17552.5 7812.5 17927.5 ;
      RECT  7517.5 17710.0 7452.5 17895.0 ;
      RECT  7517.5 16550.0 7452.5 16735.0 ;
      RECT  8257.5 17552.5 8192.5 17687.5 ;
      RECT  8067.5 17552.5 8002.5 17687.5 ;
      RECT  8067.5 17552.5 8002.5 17687.5 ;
      RECT  8257.5 17552.5 8192.5 17687.5 ;
      RECT  8067.5 17552.5 8002.5 17687.5 ;
      RECT  7877.5 17552.5 7812.5 17687.5 ;
      RECT  7877.5 17552.5 7812.5 17687.5 ;
      RECT  8067.5 17552.5 8002.5 17687.5 ;
      RECT  7877.5 17552.5 7812.5 17687.5 ;
      RECT  7687.5 17552.5 7622.5 17687.5 ;
      RECT  7687.5 17552.5 7622.5 17687.5 ;
      RECT  7877.5 17552.5 7812.5 17687.5 ;
      RECT  8257.5 16712.5 8192.5 16847.5 ;
      RECT  8067.5 16712.5 8002.5 16847.5 ;
      RECT  8067.5 16712.5 8002.5 16847.5 ;
      RECT  8257.5 16712.5 8192.5 16847.5 ;
      RECT  8067.5 16712.5 8002.5 16847.5 ;
      RECT  7877.5 16712.5 7812.5 16847.5 ;
      RECT  7877.5 16712.5 7812.5 16847.5 ;
      RECT  8067.5 16712.5 8002.5 16847.5 ;
      RECT  7877.5 16712.5 7812.5 16847.5 ;
      RECT  7687.5 16712.5 7622.5 16847.5 ;
      RECT  7687.5 16712.5 7622.5 16847.5 ;
      RECT  7877.5 16712.5 7812.5 16847.5 ;
      RECT  7517.5 17642.5 7452.5 17777.5 ;
      RECT  7517.5 16667.5 7452.5 16802.5 ;
      RECT  7682.5 16925.0 7817.5 16990.0 ;
      RECT  7872.5 17065.0 8007.5 17130.0 ;
      RECT  8062.5 17205.0 8197.5 17270.0 ;
      RECT  8067.5 17552.5 8002.5 17687.5 ;
      RECT  7687.5 17552.5 7622.5 17687.5 ;
      RECT  7687.5 16712.5 7622.5 16847.5 ;
      RECT  7687.5 17170.0 7622.5 17305.0 ;
      RECT  8197.5 17205.0 8062.5 17270.0 ;
      RECT  8007.5 17065.0 7872.5 17130.0 ;
      RECT  7817.5 16925.0 7682.5 16990.0 ;
      RECT  7687.5 17170.0 7622.5 17305.0 ;
      RECT  8325.0 17862.5 7315.0 17927.5 ;
      RECT  8325.0 16517.5 7315.0 16582.5 ;
      RECT  8257.5 19077.5 8192.5 19272.5 ;
      RECT  8257.5 18237.5 8192.5 17862.5 ;
      RECT  7877.5 18237.5 7812.5 17862.5 ;
      RECT  7517.5 18080.0 7452.5 17895.0 ;
      RECT  7517.5 19240.0 7452.5 19055.0 ;
      RECT  8257.5 18237.5 8192.5 18102.5 ;
      RECT  8067.5 18237.5 8002.5 18102.5 ;
      RECT  8067.5 18237.5 8002.5 18102.5 ;
      RECT  8257.5 18237.5 8192.5 18102.5 ;
      RECT  8067.5 18237.5 8002.5 18102.5 ;
      RECT  7877.5 18237.5 7812.5 18102.5 ;
      RECT  7877.5 18237.5 7812.5 18102.5 ;
      RECT  8067.5 18237.5 8002.5 18102.5 ;
      RECT  7877.5 18237.5 7812.5 18102.5 ;
      RECT  7687.5 18237.5 7622.5 18102.5 ;
      RECT  7687.5 18237.5 7622.5 18102.5 ;
      RECT  7877.5 18237.5 7812.5 18102.5 ;
      RECT  8257.5 19077.5 8192.5 18942.5 ;
      RECT  8067.5 19077.5 8002.5 18942.5 ;
      RECT  8067.5 19077.5 8002.5 18942.5 ;
      RECT  8257.5 19077.5 8192.5 18942.5 ;
      RECT  8067.5 19077.5 8002.5 18942.5 ;
      RECT  7877.5 19077.5 7812.5 18942.5 ;
      RECT  7877.5 19077.5 7812.5 18942.5 ;
      RECT  8067.5 19077.5 8002.5 18942.5 ;
      RECT  7877.5 19077.5 7812.5 18942.5 ;
      RECT  7687.5 19077.5 7622.5 18942.5 ;
      RECT  7687.5 19077.5 7622.5 18942.5 ;
      RECT  7877.5 19077.5 7812.5 18942.5 ;
      RECT  7517.5 18147.5 7452.5 18012.5 ;
      RECT  7517.5 19122.5 7452.5 18987.5 ;
      RECT  7682.5 18865.0 7817.5 18800.0 ;
      RECT  7872.5 18725.0 8007.5 18660.0 ;
      RECT  8062.5 18585.0 8197.5 18520.0 ;
      RECT  8067.5 18237.5 8002.5 18102.5 ;
      RECT  7687.5 18237.5 7622.5 18102.5 ;
      RECT  7687.5 19077.5 7622.5 18942.5 ;
      RECT  7687.5 18620.0 7622.5 18485.0 ;
      RECT  8197.5 18585.0 8062.5 18520.0 ;
      RECT  8007.5 18725.0 7872.5 18660.0 ;
      RECT  7817.5 18865.0 7682.5 18800.0 ;
      RECT  7687.5 18620.0 7622.5 18485.0 ;
      RECT  8325.0 17927.5 7315.0 17862.5 ;
      RECT  8325.0 19272.5 7315.0 19207.5 ;
      RECT  8257.5 19402.5 8192.5 19207.5 ;
      RECT  8257.5 20242.5 8192.5 20617.5 ;
      RECT  7877.5 20242.5 7812.5 20617.5 ;
      RECT  7517.5 20400.0 7452.5 20585.0 ;
      RECT  7517.5 19240.0 7452.5 19425.0 ;
      RECT  8257.5 20242.5 8192.5 20377.5 ;
      RECT  8067.5 20242.5 8002.5 20377.5 ;
      RECT  8067.5 20242.5 8002.5 20377.5 ;
      RECT  8257.5 20242.5 8192.5 20377.5 ;
      RECT  8067.5 20242.5 8002.5 20377.5 ;
      RECT  7877.5 20242.5 7812.5 20377.5 ;
      RECT  7877.5 20242.5 7812.5 20377.5 ;
      RECT  8067.5 20242.5 8002.5 20377.5 ;
      RECT  7877.5 20242.5 7812.5 20377.5 ;
      RECT  7687.5 20242.5 7622.5 20377.5 ;
      RECT  7687.5 20242.5 7622.5 20377.5 ;
      RECT  7877.5 20242.5 7812.5 20377.5 ;
      RECT  8257.5 19402.5 8192.5 19537.5 ;
      RECT  8067.5 19402.5 8002.5 19537.5 ;
      RECT  8067.5 19402.5 8002.5 19537.5 ;
      RECT  8257.5 19402.5 8192.5 19537.5 ;
      RECT  8067.5 19402.5 8002.5 19537.5 ;
      RECT  7877.5 19402.5 7812.5 19537.5 ;
      RECT  7877.5 19402.5 7812.5 19537.5 ;
      RECT  8067.5 19402.5 8002.5 19537.5 ;
      RECT  7877.5 19402.5 7812.5 19537.5 ;
      RECT  7687.5 19402.5 7622.5 19537.5 ;
      RECT  7687.5 19402.5 7622.5 19537.5 ;
      RECT  7877.5 19402.5 7812.5 19537.5 ;
      RECT  7517.5 20332.5 7452.5 20467.5 ;
      RECT  7517.5 19357.5 7452.5 19492.5 ;
      RECT  7682.5 19615.0 7817.5 19680.0 ;
      RECT  7872.5 19755.0 8007.5 19820.0 ;
      RECT  8062.5 19895.0 8197.5 19960.0 ;
      RECT  8067.5 20242.5 8002.5 20377.5 ;
      RECT  7687.5 20242.5 7622.5 20377.5 ;
      RECT  7687.5 19402.5 7622.5 19537.5 ;
      RECT  7687.5 19860.0 7622.5 19995.0 ;
      RECT  8197.5 19895.0 8062.5 19960.0 ;
      RECT  8007.5 19755.0 7872.5 19820.0 ;
      RECT  7817.5 19615.0 7682.5 19680.0 ;
      RECT  7687.5 19860.0 7622.5 19995.0 ;
      RECT  8325.0 20552.5 7315.0 20617.5 ;
      RECT  8325.0 19207.5 7315.0 19272.5 ;
      RECT  8257.5 21767.5 8192.5 21962.5 ;
      RECT  8257.5 20927.5 8192.5 20552.5 ;
      RECT  7877.5 20927.5 7812.5 20552.5 ;
      RECT  7517.5 20770.0 7452.5 20585.0 ;
      RECT  7517.5 21930.0 7452.5 21745.0 ;
      RECT  8257.5 20927.5 8192.5 20792.5 ;
      RECT  8067.5 20927.5 8002.5 20792.5 ;
      RECT  8067.5 20927.5 8002.5 20792.5 ;
      RECT  8257.5 20927.5 8192.5 20792.5 ;
      RECT  8067.5 20927.5 8002.5 20792.5 ;
      RECT  7877.5 20927.5 7812.5 20792.5 ;
      RECT  7877.5 20927.5 7812.5 20792.5 ;
      RECT  8067.5 20927.5 8002.5 20792.5 ;
      RECT  7877.5 20927.5 7812.5 20792.5 ;
      RECT  7687.5 20927.5 7622.5 20792.5 ;
      RECT  7687.5 20927.5 7622.5 20792.5 ;
      RECT  7877.5 20927.5 7812.5 20792.5 ;
      RECT  8257.5 21767.5 8192.5 21632.5 ;
      RECT  8067.5 21767.5 8002.5 21632.5 ;
      RECT  8067.5 21767.5 8002.5 21632.5 ;
      RECT  8257.5 21767.5 8192.5 21632.5 ;
      RECT  8067.5 21767.5 8002.5 21632.5 ;
      RECT  7877.5 21767.5 7812.5 21632.5 ;
      RECT  7877.5 21767.5 7812.5 21632.5 ;
      RECT  8067.5 21767.5 8002.5 21632.5 ;
      RECT  7877.5 21767.5 7812.5 21632.5 ;
      RECT  7687.5 21767.5 7622.5 21632.5 ;
      RECT  7687.5 21767.5 7622.5 21632.5 ;
      RECT  7877.5 21767.5 7812.5 21632.5 ;
      RECT  7517.5 20837.5 7452.5 20702.5 ;
      RECT  7517.5 21812.5 7452.5 21677.5 ;
      RECT  7682.5 21555.0 7817.5 21490.0 ;
      RECT  7872.5 21415.0 8007.5 21350.0 ;
      RECT  8062.5 21275.0 8197.5 21210.0 ;
      RECT  8067.5 20927.5 8002.5 20792.5 ;
      RECT  7687.5 20927.5 7622.5 20792.5 ;
      RECT  7687.5 21767.5 7622.5 21632.5 ;
      RECT  7687.5 21310.0 7622.5 21175.0 ;
      RECT  8197.5 21275.0 8062.5 21210.0 ;
      RECT  8007.5 21415.0 7872.5 21350.0 ;
      RECT  7817.5 21555.0 7682.5 21490.0 ;
      RECT  7687.5 21310.0 7622.5 21175.0 ;
      RECT  8325.0 20617.5 7315.0 20552.5 ;
      RECT  8325.0 21962.5 7315.0 21897.5 ;
      RECT  8257.5 22092.5 8192.5 21897.5 ;
      RECT  8257.5 22932.5 8192.5 23307.5 ;
      RECT  7877.5 22932.5 7812.5 23307.5 ;
      RECT  7517.5 23090.0 7452.5 23275.0 ;
      RECT  7517.5 21930.0 7452.5 22115.0 ;
      RECT  8257.5 22932.5 8192.5 23067.5 ;
      RECT  8067.5 22932.5 8002.5 23067.5 ;
      RECT  8067.5 22932.5 8002.5 23067.5 ;
      RECT  8257.5 22932.5 8192.5 23067.5 ;
      RECT  8067.5 22932.5 8002.5 23067.5 ;
      RECT  7877.5 22932.5 7812.5 23067.5 ;
      RECT  7877.5 22932.5 7812.5 23067.5 ;
      RECT  8067.5 22932.5 8002.5 23067.5 ;
      RECT  7877.5 22932.5 7812.5 23067.5 ;
      RECT  7687.5 22932.5 7622.5 23067.5 ;
      RECT  7687.5 22932.5 7622.5 23067.5 ;
      RECT  7877.5 22932.5 7812.5 23067.5 ;
      RECT  8257.5 22092.5 8192.5 22227.5 ;
      RECT  8067.5 22092.5 8002.5 22227.5 ;
      RECT  8067.5 22092.5 8002.5 22227.5 ;
      RECT  8257.5 22092.5 8192.5 22227.5 ;
      RECT  8067.5 22092.5 8002.5 22227.5 ;
      RECT  7877.5 22092.5 7812.5 22227.5 ;
      RECT  7877.5 22092.5 7812.5 22227.5 ;
      RECT  8067.5 22092.5 8002.5 22227.5 ;
      RECT  7877.5 22092.5 7812.5 22227.5 ;
      RECT  7687.5 22092.5 7622.5 22227.5 ;
      RECT  7687.5 22092.5 7622.5 22227.5 ;
      RECT  7877.5 22092.5 7812.5 22227.5 ;
      RECT  7517.5 23022.5 7452.5 23157.5 ;
      RECT  7517.5 22047.5 7452.5 22182.5 ;
      RECT  7682.5 22305.0 7817.5 22370.0 ;
      RECT  7872.5 22445.0 8007.5 22510.0 ;
      RECT  8062.5 22585.0 8197.5 22650.0 ;
      RECT  8067.5 22932.5 8002.5 23067.5 ;
      RECT  7687.5 22932.5 7622.5 23067.5 ;
      RECT  7687.5 22092.5 7622.5 22227.5 ;
      RECT  7687.5 22550.0 7622.5 22685.0 ;
      RECT  8197.5 22585.0 8062.5 22650.0 ;
      RECT  8007.5 22445.0 7872.5 22510.0 ;
      RECT  7817.5 22305.0 7682.5 22370.0 ;
      RECT  7687.5 22550.0 7622.5 22685.0 ;
      RECT  8325.0 23242.5 7315.0 23307.5 ;
      RECT  8325.0 21897.5 7315.0 21962.5 ;
      RECT  8257.5 24457.5 8192.5 24652.5 ;
      RECT  8257.5 23617.5 8192.5 23242.5 ;
      RECT  7877.5 23617.5 7812.5 23242.5 ;
      RECT  7517.5 23460.0 7452.5 23275.0 ;
      RECT  7517.5 24620.0 7452.5 24435.0 ;
      RECT  8257.5 23617.5 8192.5 23482.5 ;
      RECT  8067.5 23617.5 8002.5 23482.5 ;
      RECT  8067.5 23617.5 8002.5 23482.5 ;
      RECT  8257.5 23617.5 8192.5 23482.5 ;
      RECT  8067.5 23617.5 8002.5 23482.5 ;
      RECT  7877.5 23617.5 7812.5 23482.5 ;
      RECT  7877.5 23617.5 7812.5 23482.5 ;
      RECT  8067.5 23617.5 8002.5 23482.5 ;
      RECT  7877.5 23617.5 7812.5 23482.5 ;
      RECT  7687.5 23617.5 7622.5 23482.5 ;
      RECT  7687.5 23617.5 7622.5 23482.5 ;
      RECT  7877.5 23617.5 7812.5 23482.5 ;
      RECT  8257.5 24457.5 8192.5 24322.5 ;
      RECT  8067.5 24457.5 8002.5 24322.5 ;
      RECT  8067.5 24457.5 8002.5 24322.5 ;
      RECT  8257.5 24457.5 8192.5 24322.5 ;
      RECT  8067.5 24457.5 8002.5 24322.5 ;
      RECT  7877.5 24457.5 7812.5 24322.5 ;
      RECT  7877.5 24457.5 7812.5 24322.5 ;
      RECT  8067.5 24457.5 8002.5 24322.5 ;
      RECT  7877.5 24457.5 7812.5 24322.5 ;
      RECT  7687.5 24457.5 7622.5 24322.5 ;
      RECT  7687.5 24457.5 7622.5 24322.5 ;
      RECT  7877.5 24457.5 7812.5 24322.5 ;
      RECT  7517.5 23527.5 7452.5 23392.5 ;
      RECT  7517.5 24502.5 7452.5 24367.5 ;
      RECT  7682.5 24245.0 7817.5 24180.0 ;
      RECT  7872.5 24105.0 8007.5 24040.0 ;
      RECT  8062.5 23965.0 8197.5 23900.0 ;
      RECT  8067.5 23617.5 8002.5 23482.5 ;
      RECT  7687.5 23617.5 7622.5 23482.5 ;
      RECT  7687.5 24457.5 7622.5 24322.5 ;
      RECT  7687.5 24000.0 7622.5 23865.0 ;
      RECT  8197.5 23965.0 8062.5 23900.0 ;
      RECT  8007.5 24105.0 7872.5 24040.0 ;
      RECT  7817.5 24245.0 7682.5 24180.0 ;
      RECT  7687.5 24000.0 7622.5 23865.0 ;
      RECT  8325.0 23307.5 7315.0 23242.5 ;
      RECT  8325.0 24652.5 7315.0 24587.5 ;
      RECT  8257.5 24782.5 8192.5 24587.5 ;
      RECT  8257.5 25622.5 8192.5 25997.5 ;
      RECT  7877.5 25622.5 7812.5 25997.5 ;
      RECT  7517.5 25780.0 7452.5 25965.0 ;
      RECT  7517.5 24620.0 7452.5 24805.0 ;
      RECT  8257.5 25622.5 8192.5 25757.5 ;
      RECT  8067.5 25622.5 8002.5 25757.5 ;
      RECT  8067.5 25622.5 8002.5 25757.5 ;
      RECT  8257.5 25622.5 8192.5 25757.5 ;
      RECT  8067.5 25622.5 8002.5 25757.5 ;
      RECT  7877.5 25622.5 7812.5 25757.5 ;
      RECT  7877.5 25622.5 7812.5 25757.5 ;
      RECT  8067.5 25622.5 8002.5 25757.5 ;
      RECT  7877.5 25622.5 7812.5 25757.5 ;
      RECT  7687.5 25622.5 7622.5 25757.5 ;
      RECT  7687.5 25622.5 7622.5 25757.5 ;
      RECT  7877.5 25622.5 7812.5 25757.5 ;
      RECT  8257.5 24782.5 8192.5 24917.5 ;
      RECT  8067.5 24782.5 8002.5 24917.5 ;
      RECT  8067.5 24782.5 8002.5 24917.5 ;
      RECT  8257.5 24782.5 8192.5 24917.5 ;
      RECT  8067.5 24782.5 8002.5 24917.5 ;
      RECT  7877.5 24782.5 7812.5 24917.5 ;
      RECT  7877.5 24782.5 7812.5 24917.5 ;
      RECT  8067.5 24782.5 8002.5 24917.5 ;
      RECT  7877.5 24782.5 7812.5 24917.5 ;
      RECT  7687.5 24782.5 7622.5 24917.5 ;
      RECT  7687.5 24782.5 7622.5 24917.5 ;
      RECT  7877.5 24782.5 7812.5 24917.5 ;
      RECT  7517.5 25712.5 7452.5 25847.5 ;
      RECT  7517.5 24737.5 7452.5 24872.5 ;
      RECT  7682.5 24995.0 7817.5 25060.0 ;
      RECT  7872.5 25135.0 8007.5 25200.0 ;
      RECT  8062.5 25275.0 8197.5 25340.0 ;
      RECT  8067.5 25622.5 8002.5 25757.5 ;
      RECT  7687.5 25622.5 7622.5 25757.5 ;
      RECT  7687.5 24782.5 7622.5 24917.5 ;
      RECT  7687.5 25240.0 7622.5 25375.0 ;
      RECT  8197.5 25275.0 8062.5 25340.0 ;
      RECT  8007.5 25135.0 7872.5 25200.0 ;
      RECT  7817.5 24995.0 7682.5 25060.0 ;
      RECT  7687.5 25240.0 7622.5 25375.0 ;
      RECT  8325.0 25932.5 7315.0 25997.5 ;
      RECT  8325.0 24587.5 7315.0 24652.5 ;
      RECT  8257.5 27147.5 8192.5 27342.5 ;
      RECT  8257.5 26307.5 8192.5 25932.5 ;
      RECT  7877.5 26307.5 7812.5 25932.5 ;
      RECT  7517.5 26150.0 7452.5 25965.0 ;
      RECT  7517.5 27310.0 7452.5 27125.0 ;
      RECT  8257.5 26307.5 8192.5 26172.5 ;
      RECT  8067.5 26307.5 8002.5 26172.5 ;
      RECT  8067.5 26307.5 8002.5 26172.5 ;
      RECT  8257.5 26307.5 8192.5 26172.5 ;
      RECT  8067.5 26307.5 8002.5 26172.5 ;
      RECT  7877.5 26307.5 7812.5 26172.5 ;
      RECT  7877.5 26307.5 7812.5 26172.5 ;
      RECT  8067.5 26307.5 8002.5 26172.5 ;
      RECT  7877.5 26307.5 7812.5 26172.5 ;
      RECT  7687.5 26307.5 7622.5 26172.5 ;
      RECT  7687.5 26307.5 7622.5 26172.5 ;
      RECT  7877.5 26307.5 7812.5 26172.5 ;
      RECT  8257.5 27147.5 8192.5 27012.5 ;
      RECT  8067.5 27147.5 8002.5 27012.5 ;
      RECT  8067.5 27147.5 8002.5 27012.5 ;
      RECT  8257.5 27147.5 8192.5 27012.5 ;
      RECT  8067.5 27147.5 8002.5 27012.5 ;
      RECT  7877.5 27147.5 7812.5 27012.5 ;
      RECT  7877.5 27147.5 7812.5 27012.5 ;
      RECT  8067.5 27147.5 8002.5 27012.5 ;
      RECT  7877.5 27147.5 7812.5 27012.5 ;
      RECT  7687.5 27147.5 7622.5 27012.5 ;
      RECT  7687.5 27147.5 7622.5 27012.5 ;
      RECT  7877.5 27147.5 7812.5 27012.5 ;
      RECT  7517.5 26217.5 7452.5 26082.5 ;
      RECT  7517.5 27192.5 7452.5 27057.5 ;
      RECT  7682.5 26935.0 7817.5 26870.0 ;
      RECT  7872.5 26795.0 8007.5 26730.0 ;
      RECT  8062.5 26655.0 8197.5 26590.0 ;
      RECT  8067.5 26307.5 8002.5 26172.5 ;
      RECT  7687.5 26307.5 7622.5 26172.5 ;
      RECT  7687.5 27147.5 7622.5 27012.5 ;
      RECT  7687.5 26690.0 7622.5 26555.0 ;
      RECT  8197.5 26655.0 8062.5 26590.0 ;
      RECT  8007.5 26795.0 7872.5 26730.0 ;
      RECT  7817.5 26935.0 7682.5 26870.0 ;
      RECT  7687.5 26690.0 7622.5 26555.0 ;
      RECT  8325.0 25997.5 7315.0 25932.5 ;
      RECT  8325.0 27342.5 7315.0 27277.5 ;
      RECT  9872.5 17667.5 10007.5 17732.5 ;
      RECT  11532.5 17145.0 11667.5 17210.0 ;
      RECT  9597.5 19012.5 9732.5 19077.5 ;
      RECT  11257.5 18580.0 11392.5 18645.0 ;
      RECT  9322.5 20357.5 9457.5 20422.5 ;
      RECT  10982.5 19835.0 11117.5 19900.0 ;
      RECT  11532.5 20687.5 11667.5 20752.5 ;
      RECT  9047.5 20687.5 9182.5 20752.5 ;
      RECT  11257.5 22032.5 11392.5 22097.5 ;
      RECT  8772.5 22032.5 8907.5 22097.5 ;
      RECT  10982.5 23377.5 11117.5 23442.5 ;
      RECT  8497.5 23377.5 8632.5 23442.5 ;
      RECT  9872.5 17205.0 10007.5 17270.0 ;
      RECT  9597.5 17065.0 9732.5 17130.0 ;
      RECT  9322.5 16925.0 9457.5 16990.0 ;
      RECT  9047.5 18520.0 9182.5 18585.0 ;
      RECT  9597.5 18660.0 9732.5 18725.0 ;
      RECT  9322.5 18800.0 9457.5 18865.0 ;
      RECT  9872.5 19895.0 10007.5 19960.0 ;
      RECT  8772.5 19755.0 8907.5 19820.0 ;
      RECT  9322.5 19615.0 9457.5 19680.0 ;
      RECT  9047.5 21210.0 9182.5 21275.0 ;
      RECT  8772.5 21350.0 8907.5 21415.0 ;
      RECT  9322.5 21490.0 9457.5 21555.0 ;
      RECT  9872.5 22585.0 10007.5 22650.0 ;
      RECT  9597.5 22445.0 9732.5 22510.0 ;
      RECT  8497.5 22305.0 8632.5 22370.0 ;
      RECT  9047.5 23900.0 9182.5 23965.0 ;
      RECT  9597.5 24040.0 9732.5 24105.0 ;
      RECT  8497.5 24180.0 8632.5 24245.0 ;
      RECT  9872.5 25275.0 10007.5 25340.0 ;
      RECT  8772.5 25135.0 8907.5 25200.0 ;
      RECT  8497.5 24995.0 8632.5 25060.0 ;
      RECT  9047.5 26590.0 9182.5 26655.0 ;
      RECT  8772.5 26730.0 8907.5 26795.0 ;
      RECT  8497.5 26870.0 8632.5 26935.0 ;
      RECT  6960.0 17145.0 6755.0 17210.0 ;
      RECT  6960.0 18580.0 6755.0 18645.0 ;
      RECT  6960.0 19835.0 6755.0 19900.0 ;
      RECT  6960.0 21270.0 6755.0 21335.0 ;
      RECT  6960.0 22525.0 6755.0 22590.0 ;
      RECT  6960.0 23960.0 6755.0 24025.0 ;
      RECT  6960.0 25215.0 6755.0 25280.0 ;
      RECT  6960.0 26650.0 6755.0 26715.0 ;
      RECT  11635.0 17862.5 6755.0 17927.5 ;
      RECT  11635.0 20552.5 6755.0 20617.5 ;
      RECT  11635.0 23242.5 6755.0 23307.5 ;
      RECT  11635.0 25932.5 6755.0 25997.5 ;
      RECT  11635.0 16517.5 6755.0 16582.5 ;
      RECT  11635.0 19207.5 6755.0 19272.5 ;
      RECT  11635.0 21897.5 6755.0 21962.5 ;
      RECT  11635.0 24587.5 6755.0 24652.5 ;
      RECT  11635.0 27277.5 6755.0 27342.5 ;
      RECT  6822.5 27472.5 6887.5 27277.5 ;
      RECT  6822.5 28312.5 6887.5 28687.5 ;
      RECT  7202.5 28312.5 7267.5 28687.5 ;
      RECT  7372.5 28470.0 7437.5 28655.0 ;
      RECT  7372.5 27310.0 7437.5 27495.0 ;
      RECT  6822.5 28312.5 6887.5 28447.5 ;
      RECT  7012.5 28312.5 7077.5 28447.5 ;
      RECT  7012.5 28312.5 7077.5 28447.5 ;
      RECT  6822.5 28312.5 6887.5 28447.5 ;
      RECT  7012.5 28312.5 7077.5 28447.5 ;
      RECT  7202.5 28312.5 7267.5 28447.5 ;
      RECT  7202.5 28312.5 7267.5 28447.5 ;
      RECT  7012.5 28312.5 7077.5 28447.5 ;
      RECT  6822.5 27472.5 6887.5 27607.5 ;
      RECT  7012.5 27472.5 7077.5 27607.5 ;
      RECT  7012.5 27472.5 7077.5 27607.5 ;
      RECT  6822.5 27472.5 6887.5 27607.5 ;
      RECT  7012.5 27472.5 7077.5 27607.5 ;
      RECT  7202.5 27472.5 7267.5 27607.5 ;
      RECT  7202.5 27472.5 7267.5 27607.5 ;
      RECT  7012.5 27472.5 7077.5 27607.5 ;
      RECT  7372.5 28402.5 7437.5 28537.5 ;
      RECT  7372.5 27427.5 7437.5 27562.5 ;
      RECT  7207.5 27702.5 7072.5 27767.5 ;
      RECT  6950.0 27917.5 6815.0 27982.5 ;
      RECT  7012.5 28312.5 7077.5 28447.5 ;
      RECT  7202.5 27472.5 7267.5 27607.5 ;
      RECT  7302.5 27917.5 7167.5 27982.5 ;
      RECT  6815.0 27917.5 6950.0 27982.5 ;
      RECT  7072.5 27702.5 7207.5 27767.5 ;
      RECT  7167.5 27917.5 7302.5 27982.5 ;
      RECT  6755.0 28622.5 7675.0 28687.5 ;
      RECT  6755.0 27277.5 7675.0 27342.5 ;
      RECT  6822.5 29837.5 6887.5 30032.5 ;
      RECT  6822.5 28997.5 6887.5 28622.5 ;
      RECT  7202.5 28997.5 7267.5 28622.5 ;
      RECT  7372.5 28840.0 7437.5 28655.0 ;
      RECT  7372.5 30000.0 7437.5 29815.0 ;
      RECT  6822.5 28997.5 6887.5 28862.5 ;
      RECT  7012.5 28997.5 7077.5 28862.5 ;
      RECT  7012.5 28997.5 7077.5 28862.5 ;
      RECT  6822.5 28997.5 6887.5 28862.5 ;
      RECT  7012.5 28997.5 7077.5 28862.5 ;
      RECT  7202.5 28997.5 7267.5 28862.5 ;
      RECT  7202.5 28997.5 7267.5 28862.5 ;
      RECT  7012.5 28997.5 7077.5 28862.5 ;
      RECT  6822.5 29837.5 6887.5 29702.5 ;
      RECT  7012.5 29837.5 7077.5 29702.5 ;
      RECT  7012.5 29837.5 7077.5 29702.5 ;
      RECT  6822.5 29837.5 6887.5 29702.5 ;
      RECT  7012.5 29837.5 7077.5 29702.5 ;
      RECT  7202.5 29837.5 7267.5 29702.5 ;
      RECT  7202.5 29837.5 7267.5 29702.5 ;
      RECT  7012.5 29837.5 7077.5 29702.5 ;
      RECT  7372.5 28907.5 7437.5 28772.5 ;
      RECT  7372.5 29882.5 7437.5 29747.5 ;
      RECT  7207.5 29607.5 7072.5 29542.5 ;
      RECT  6950.0 29392.5 6815.0 29327.5 ;
      RECT  7012.5 28997.5 7077.5 28862.5 ;
      RECT  7202.5 29837.5 7267.5 29702.5 ;
      RECT  7302.5 29392.5 7167.5 29327.5 ;
      RECT  6815.0 29392.5 6950.0 29327.5 ;
      RECT  7072.5 29607.5 7207.5 29542.5 ;
      RECT  7167.5 29392.5 7302.5 29327.5 ;
      RECT  6755.0 28687.5 7675.0 28622.5 ;
      RECT  6755.0 30032.5 7675.0 29967.5 ;
      RECT  6822.5 30162.5 6887.5 29967.5 ;
      RECT  6822.5 31002.5 6887.5 31377.5 ;
      RECT  7202.5 31002.5 7267.5 31377.5 ;
      RECT  7372.5 31160.0 7437.5 31345.0 ;
      RECT  7372.5 30000.0 7437.5 30185.0 ;
      RECT  6822.5 31002.5 6887.5 31137.5 ;
      RECT  7012.5 31002.5 7077.5 31137.5 ;
      RECT  7012.5 31002.5 7077.5 31137.5 ;
      RECT  6822.5 31002.5 6887.5 31137.5 ;
      RECT  7012.5 31002.5 7077.5 31137.5 ;
      RECT  7202.5 31002.5 7267.5 31137.5 ;
      RECT  7202.5 31002.5 7267.5 31137.5 ;
      RECT  7012.5 31002.5 7077.5 31137.5 ;
      RECT  6822.5 30162.5 6887.5 30297.5 ;
      RECT  7012.5 30162.5 7077.5 30297.5 ;
      RECT  7012.5 30162.5 7077.5 30297.5 ;
      RECT  6822.5 30162.5 6887.5 30297.5 ;
      RECT  7012.5 30162.5 7077.5 30297.5 ;
      RECT  7202.5 30162.5 7267.5 30297.5 ;
      RECT  7202.5 30162.5 7267.5 30297.5 ;
      RECT  7012.5 30162.5 7077.5 30297.5 ;
      RECT  7372.5 31092.5 7437.5 31227.5 ;
      RECT  7372.5 30117.5 7437.5 30252.5 ;
      RECT  7207.5 30392.5 7072.5 30457.5 ;
      RECT  6950.0 30607.5 6815.0 30672.5 ;
      RECT  7012.5 31002.5 7077.5 31137.5 ;
      RECT  7202.5 30162.5 7267.5 30297.5 ;
      RECT  7302.5 30607.5 7167.5 30672.5 ;
      RECT  6815.0 30607.5 6950.0 30672.5 ;
      RECT  7072.5 30392.5 7207.5 30457.5 ;
      RECT  7167.5 30607.5 7302.5 30672.5 ;
      RECT  6755.0 31312.5 7675.0 31377.5 ;
      RECT  6755.0 29967.5 7675.0 30032.5 ;
      RECT  6822.5 32527.5 6887.5 32722.5 ;
      RECT  6822.5 31687.5 6887.5 31312.5 ;
      RECT  7202.5 31687.5 7267.5 31312.5 ;
      RECT  7372.5 31530.0 7437.5 31345.0 ;
      RECT  7372.5 32690.0 7437.5 32505.0 ;
      RECT  6822.5 31687.5 6887.5 31552.5 ;
      RECT  7012.5 31687.5 7077.5 31552.5 ;
      RECT  7012.5 31687.5 7077.5 31552.5 ;
      RECT  6822.5 31687.5 6887.5 31552.5 ;
      RECT  7012.5 31687.5 7077.5 31552.5 ;
      RECT  7202.5 31687.5 7267.5 31552.5 ;
      RECT  7202.5 31687.5 7267.5 31552.5 ;
      RECT  7012.5 31687.5 7077.5 31552.5 ;
      RECT  6822.5 32527.5 6887.5 32392.5 ;
      RECT  7012.5 32527.5 7077.5 32392.5 ;
      RECT  7012.5 32527.5 7077.5 32392.5 ;
      RECT  6822.5 32527.5 6887.5 32392.5 ;
      RECT  7012.5 32527.5 7077.5 32392.5 ;
      RECT  7202.5 32527.5 7267.5 32392.5 ;
      RECT  7202.5 32527.5 7267.5 32392.5 ;
      RECT  7012.5 32527.5 7077.5 32392.5 ;
      RECT  7372.5 31597.5 7437.5 31462.5 ;
      RECT  7372.5 32572.5 7437.5 32437.5 ;
      RECT  7207.5 32297.5 7072.5 32232.5 ;
      RECT  6950.0 32082.5 6815.0 32017.5 ;
      RECT  7012.5 31687.5 7077.5 31552.5 ;
      RECT  7202.5 32527.5 7267.5 32392.5 ;
      RECT  7302.5 32082.5 7167.5 32017.5 ;
      RECT  6815.0 32082.5 6950.0 32017.5 ;
      RECT  7072.5 32297.5 7207.5 32232.5 ;
      RECT  7167.5 32082.5 7302.5 32017.5 ;
      RECT  6755.0 31377.5 7675.0 31312.5 ;
      RECT  6755.0 32722.5 7675.0 32657.5 ;
      RECT  6822.5 32852.5 6887.5 32657.5 ;
      RECT  6822.5 33692.5 6887.5 34067.5 ;
      RECT  7202.5 33692.5 7267.5 34067.5 ;
      RECT  7372.5 33850.0 7437.5 34035.0 ;
      RECT  7372.5 32690.0 7437.5 32875.0 ;
      RECT  6822.5 33692.5 6887.5 33827.5 ;
      RECT  7012.5 33692.5 7077.5 33827.5 ;
      RECT  7012.5 33692.5 7077.5 33827.5 ;
      RECT  6822.5 33692.5 6887.5 33827.5 ;
      RECT  7012.5 33692.5 7077.5 33827.5 ;
      RECT  7202.5 33692.5 7267.5 33827.5 ;
      RECT  7202.5 33692.5 7267.5 33827.5 ;
      RECT  7012.5 33692.5 7077.5 33827.5 ;
      RECT  6822.5 32852.5 6887.5 32987.5 ;
      RECT  7012.5 32852.5 7077.5 32987.5 ;
      RECT  7012.5 32852.5 7077.5 32987.5 ;
      RECT  6822.5 32852.5 6887.5 32987.5 ;
      RECT  7012.5 32852.5 7077.5 32987.5 ;
      RECT  7202.5 32852.5 7267.5 32987.5 ;
      RECT  7202.5 32852.5 7267.5 32987.5 ;
      RECT  7012.5 32852.5 7077.5 32987.5 ;
      RECT  7372.5 33782.5 7437.5 33917.5 ;
      RECT  7372.5 32807.5 7437.5 32942.5 ;
      RECT  7207.5 33082.5 7072.5 33147.5 ;
      RECT  6950.0 33297.5 6815.0 33362.5 ;
      RECT  7012.5 33692.5 7077.5 33827.5 ;
      RECT  7202.5 32852.5 7267.5 32987.5 ;
      RECT  7302.5 33297.5 7167.5 33362.5 ;
      RECT  6815.0 33297.5 6950.0 33362.5 ;
      RECT  7072.5 33082.5 7207.5 33147.5 ;
      RECT  7167.5 33297.5 7302.5 33362.5 ;
      RECT  6755.0 34002.5 7675.0 34067.5 ;
      RECT  6755.0 32657.5 7675.0 32722.5 ;
      RECT  6822.5 35217.5 6887.5 35412.5 ;
      RECT  6822.5 34377.5 6887.5 34002.5 ;
      RECT  7202.5 34377.5 7267.5 34002.5 ;
      RECT  7372.5 34220.0 7437.5 34035.0 ;
      RECT  7372.5 35380.0 7437.5 35195.0 ;
      RECT  6822.5 34377.5 6887.5 34242.5 ;
      RECT  7012.5 34377.5 7077.5 34242.5 ;
      RECT  7012.5 34377.5 7077.5 34242.5 ;
      RECT  6822.5 34377.5 6887.5 34242.5 ;
      RECT  7012.5 34377.5 7077.5 34242.5 ;
      RECT  7202.5 34377.5 7267.5 34242.5 ;
      RECT  7202.5 34377.5 7267.5 34242.5 ;
      RECT  7012.5 34377.5 7077.5 34242.5 ;
      RECT  6822.5 35217.5 6887.5 35082.5 ;
      RECT  7012.5 35217.5 7077.5 35082.5 ;
      RECT  7012.5 35217.5 7077.5 35082.5 ;
      RECT  6822.5 35217.5 6887.5 35082.5 ;
      RECT  7012.5 35217.5 7077.5 35082.5 ;
      RECT  7202.5 35217.5 7267.5 35082.5 ;
      RECT  7202.5 35217.5 7267.5 35082.5 ;
      RECT  7012.5 35217.5 7077.5 35082.5 ;
      RECT  7372.5 34287.5 7437.5 34152.5 ;
      RECT  7372.5 35262.5 7437.5 35127.5 ;
      RECT  7207.5 34987.5 7072.5 34922.5 ;
      RECT  6950.0 34772.5 6815.0 34707.5 ;
      RECT  7012.5 34377.5 7077.5 34242.5 ;
      RECT  7202.5 35217.5 7267.5 35082.5 ;
      RECT  7302.5 34772.5 7167.5 34707.5 ;
      RECT  6815.0 34772.5 6950.0 34707.5 ;
      RECT  7072.5 34987.5 7207.5 34922.5 ;
      RECT  7167.5 34772.5 7302.5 34707.5 ;
      RECT  6755.0 34067.5 7675.0 34002.5 ;
      RECT  6755.0 35412.5 7675.0 35347.5 ;
      RECT  6822.5 35542.5 6887.5 35347.5 ;
      RECT  6822.5 36382.5 6887.5 36757.5 ;
      RECT  7202.5 36382.5 7267.5 36757.5 ;
      RECT  7372.5 36540.0 7437.5 36725.0 ;
      RECT  7372.5 35380.0 7437.5 35565.0 ;
      RECT  6822.5 36382.5 6887.5 36517.5 ;
      RECT  7012.5 36382.5 7077.5 36517.5 ;
      RECT  7012.5 36382.5 7077.5 36517.5 ;
      RECT  6822.5 36382.5 6887.5 36517.5 ;
      RECT  7012.5 36382.5 7077.5 36517.5 ;
      RECT  7202.5 36382.5 7267.5 36517.5 ;
      RECT  7202.5 36382.5 7267.5 36517.5 ;
      RECT  7012.5 36382.5 7077.5 36517.5 ;
      RECT  6822.5 35542.5 6887.5 35677.5 ;
      RECT  7012.5 35542.5 7077.5 35677.5 ;
      RECT  7012.5 35542.5 7077.5 35677.5 ;
      RECT  6822.5 35542.5 6887.5 35677.5 ;
      RECT  7012.5 35542.5 7077.5 35677.5 ;
      RECT  7202.5 35542.5 7267.5 35677.5 ;
      RECT  7202.5 35542.5 7267.5 35677.5 ;
      RECT  7012.5 35542.5 7077.5 35677.5 ;
      RECT  7372.5 36472.5 7437.5 36607.5 ;
      RECT  7372.5 35497.5 7437.5 35632.5 ;
      RECT  7207.5 35772.5 7072.5 35837.5 ;
      RECT  6950.0 35987.5 6815.0 36052.5 ;
      RECT  7012.5 36382.5 7077.5 36517.5 ;
      RECT  7202.5 35542.5 7267.5 35677.5 ;
      RECT  7302.5 35987.5 7167.5 36052.5 ;
      RECT  6815.0 35987.5 6950.0 36052.5 ;
      RECT  7072.5 35772.5 7207.5 35837.5 ;
      RECT  7167.5 35987.5 7302.5 36052.5 ;
      RECT  6755.0 36692.5 7675.0 36757.5 ;
      RECT  6755.0 35347.5 7675.0 35412.5 ;
      RECT  6822.5 37907.5 6887.5 38102.5 ;
      RECT  6822.5 37067.5 6887.5 36692.5 ;
      RECT  7202.5 37067.5 7267.5 36692.5 ;
      RECT  7372.5 36910.0 7437.5 36725.0 ;
      RECT  7372.5 38070.0 7437.5 37885.0 ;
      RECT  6822.5 37067.5 6887.5 36932.5 ;
      RECT  7012.5 37067.5 7077.5 36932.5 ;
      RECT  7012.5 37067.5 7077.5 36932.5 ;
      RECT  6822.5 37067.5 6887.5 36932.5 ;
      RECT  7012.5 37067.5 7077.5 36932.5 ;
      RECT  7202.5 37067.5 7267.5 36932.5 ;
      RECT  7202.5 37067.5 7267.5 36932.5 ;
      RECT  7012.5 37067.5 7077.5 36932.5 ;
      RECT  6822.5 37907.5 6887.5 37772.5 ;
      RECT  7012.5 37907.5 7077.5 37772.5 ;
      RECT  7012.5 37907.5 7077.5 37772.5 ;
      RECT  6822.5 37907.5 6887.5 37772.5 ;
      RECT  7012.5 37907.5 7077.5 37772.5 ;
      RECT  7202.5 37907.5 7267.5 37772.5 ;
      RECT  7202.5 37907.5 7267.5 37772.5 ;
      RECT  7012.5 37907.5 7077.5 37772.5 ;
      RECT  7372.5 36977.5 7437.5 36842.5 ;
      RECT  7372.5 37952.5 7437.5 37817.5 ;
      RECT  7207.5 37677.5 7072.5 37612.5 ;
      RECT  6950.0 37462.5 6815.0 37397.5 ;
      RECT  7012.5 37067.5 7077.5 36932.5 ;
      RECT  7202.5 37907.5 7267.5 37772.5 ;
      RECT  7302.5 37462.5 7167.5 37397.5 ;
      RECT  6815.0 37462.5 6950.0 37397.5 ;
      RECT  7072.5 37677.5 7207.5 37612.5 ;
      RECT  7167.5 37462.5 7302.5 37397.5 ;
      RECT  6755.0 36757.5 7675.0 36692.5 ;
      RECT  6755.0 38102.5 7675.0 38037.5 ;
      RECT  6822.5 38232.5 6887.5 38037.5 ;
      RECT  6822.5 39072.5 6887.5 39447.5 ;
      RECT  7202.5 39072.5 7267.5 39447.5 ;
      RECT  7372.5 39230.0 7437.5 39415.0 ;
      RECT  7372.5 38070.0 7437.5 38255.0 ;
      RECT  6822.5 39072.5 6887.5 39207.5 ;
      RECT  7012.5 39072.5 7077.5 39207.5 ;
      RECT  7012.5 39072.5 7077.5 39207.5 ;
      RECT  6822.5 39072.5 6887.5 39207.5 ;
      RECT  7012.5 39072.5 7077.5 39207.5 ;
      RECT  7202.5 39072.5 7267.5 39207.5 ;
      RECT  7202.5 39072.5 7267.5 39207.5 ;
      RECT  7012.5 39072.5 7077.5 39207.5 ;
      RECT  6822.5 38232.5 6887.5 38367.5 ;
      RECT  7012.5 38232.5 7077.5 38367.5 ;
      RECT  7012.5 38232.5 7077.5 38367.5 ;
      RECT  6822.5 38232.5 6887.5 38367.5 ;
      RECT  7012.5 38232.5 7077.5 38367.5 ;
      RECT  7202.5 38232.5 7267.5 38367.5 ;
      RECT  7202.5 38232.5 7267.5 38367.5 ;
      RECT  7012.5 38232.5 7077.5 38367.5 ;
      RECT  7372.5 39162.5 7437.5 39297.5 ;
      RECT  7372.5 38187.5 7437.5 38322.5 ;
      RECT  7207.5 38462.5 7072.5 38527.5 ;
      RECT  6950.0 38677.5 6815.0 38742.5 ;
      RECT  7012.5 39072.5 7077.5 39207.5 ;
      RECT  7202.5 38232.5 7267.5 38367.5 ;
      RECT  7302.5 38677.5 7167.5 38742.5 ;
      RECT  6815.0 38677.5 6950.0 38742.5 ;
      RECT  7072.5 38462.5 7207.5 38527.5 ;
      RECT  7167.5 38677.5 7302.5 38742.5 ;
      RECT  6755.0 39382.5 7675.0 39447.5 ;
      RECT  6755.0 38037.5 7675.0 38102.5 ;
      RECT  6822.5 40597.5 6887.5 40792.5 ;
      RECT  6822.5 39757.5 6887.5 39382.5 ;
      RECT  7202.5 39757.5 7267.5 39382.5 ;
      RECT  7372.5 39600.0 7437.5 39415.0 ;
      RECT  7372.5 40760.0 7437.5 40575.0 ;
      RECT  6822.5 39757.5 6887.5 39622.5 ;
      RECT  7012.5 39757.5 7077.5 39622.5 ;
      RECT  7012.5 39757.5 7077.5 39622.5 ;
      RECT  6822.5 39757.5 6887.5 39622.5 ;
      RECT  7012.5 39757.5 7077.5 39622.5 ;
      RECT  7202.5 39757.5 7267.5 39622.5 ;
      RECT  7202.5 39757.5 7267.5 39622.5 ;
      RECT  7012.5 39757.5 7077.5 39622.5 ;
      RECT  6822.5 40597.5 6887.5 40462.5 ;
      RECT  7012.5 40597.5 7077.5 40462.5 ;
      RECT  7012.5 40597.5 7077.5 40462.5 ;
      RECT  6822.5 40597.5 6887.5 40462.5 ;
      RECT  7012.5 40597.5 7077.5 40462.5 ;
      RECT  7202.5 40597.5 7267.5 40462.5 ;
      RECT  7202.5 40597.5 7267.5 40462.5 ;
      RECT  7012.5 40597.5 7077.5 40462.5 ;
      RECT  7372.5 39667.5 7437.5 39532.5 ;
      RECT  7372.5 40642.5 7437.5 40507.5 ;
      RECT  7207.5 40367.5 7072.5 40302.5 ;
      RECT  6950.0 40152.5 6815.0 40087.5 ;
      RECT  7012.5 39757.5 7077.5 39622.5 ;
      RECT  7202.5 40597.5 7267.5 40462.5 ;
      RECT  7302.5 40152.5 7167.5 40087.5 ;
      RECT  6815.0 40152.5 6950.0 40087.5 ;
      RECT  7072.5 40367.5 7207.5 40302.5 ;
      RECT  7167.5 40152.5 7302.5 40087.5 ;
      RECT  6755.0 39447.5 7675.0 39382.5 ;
      RECT  6755.0 40792.5 7675.0 40727.5 ;
      RECT  6822.5 40922.5 6887.5 40727.5 ;
      RECT  6822.5 41762.5 6887.5 42137.5 ;
      RECT  7202.5 41762.5 7267.5 42137.5 ;
      RECT  7372.5 41920.0 7437.5 42105.0 ;
      RECT  7372.5 40760.0 7437.5 40945.0 ;
      RECT  6822.5 41762.5 6887.5 41897.5 ;
      RECT  7012.5 41762.5 7077.5 41897.5 ;
      RECT  7012.5 41762.5 7077.5 41897.5 ;
      RECT  6822.5 41762.5 6887.5 41897.5 ;
      RECT  7012.5 41762.5 7077.5 41897.5 ;
      RECT  7202.5 41762.5 7267.5 41897.5 ;
      RECT  7202.5 41762.5 7267.5 41897.5 ;
      RECT  7012.5 41762.5 7077.5 41897.5 ;
      RECT  6822.5 40922.5 6887.5 41057.5 ;
      RECT  7012.5 40922.5 7077.5 41057.5 ;
      RECT  7012.5 40922.5 7077.5 41057.5 ;
      RECT  6822.5 40922.5 6887.5 41057.5 ;
      RECT  7012.5 40922.5 7077.5 41057.5 ;
      RECT  7202.5 40922.5 7267.5 41057.5 ;
      RECT  7202.5 40922.5 7267.5 41057.5 ;
      RECT  7012.5 40922.5 7077.5 41057.5 ;
      RECT  7372.5 41852.5 7437.5 41987.5 ;
      RECT  7372.5 40877.5 7437.5 41012.5 ;
      RECT  7207.5 41152.5 7072.5 41217.5 ;
      RECT  6950.0 41367.5 6815.0 41432.5 ;
      RECT  7012.5 41762.5 7077.5 41897.5 ;
      RECT  7202.5 40922.5 7267.5 41057.5 ;
      RECT  7302.5 41367.5 7167.5 41432.5 ;
      RECT  6815.0 41367.5 6950.0 41432.5 ;
      RECT  7072.5 41152.5 7207.5 41217.5 ;
      RECT  7167.5 41367.5 7302.5 41432.5 ;
      RECT  6755.0 42072.5 7675.0 42137.5 ;
      RECT  6755.0 40727.5 7675.0 40792.5 ;
      RECT  6822.5 43287.5 6887.5 43482.5 ;
      RECT  6822.5 42447.5 6887.5 42072.5 ;
      RECT  7202.5 42447.5 7267.5 42072.5 ;
      RECT  7372.5 42290.0 7437.5 42105.0 ;
      RECT  7372.5 43450.0 7437.5 43265.0 ;
      RECT  6822.5 42447.5 6887.5 42312.5 ;
      RECT  7012.5 42447.5 7077.5 42312.5 ;
      RECT  7012.5 42447.5 7077.5 42312.5 ;
      RECT  6822.5 42447.5 6887.5 42312.5 ;
      RECT  7012.5 42447.5 7077.5 42312.5 ;
      RECT  7202.5 42447.5 7267.5 42312.5 ;
      RECT  7202.5 42447.5 7267.5 42312.5 ;
      RECT  7012.5 42447.5 7077.5 42312.5 ;
      RECT  6822.5 43287.5 6887.5 43152.5 ;
      RECT  7012.5 43287.5 7077.5 43152.5 ;
      RECT  7012.5 43287.5 7077.5 43152.5 ;
      RECT  6822.5 43287.5 6887.5 43152.5 ;
      RECT  7012.5 43287.5 7077.5 43152.5 ;
      RECT  7202.5 43287.5 7267.5 43152.5 ;
      RECT  7202.5 43287.5 7267.5 43152.5 ;
      RECT  7012.5 43287.5 7077.5 43152.5 ;
      RECT  7372.5 42357.5 7437.5 42222.5 ;
      RECT  7372.5 43332.5 7437.5 43197.5 ;
      RECT  7207.5 43057.5 7072.5 42992.5 ;
      RECT  6950.0 42842.5 6815.0 42777.5 ;
      RECT  7012.5 42447.5 7077.5 42312.5 ;
      RECT  7202.5 43287.5 7267.5 43152.5 ;
      RECT  7302.5 42842.5 7167.5 42777.5 ;
      RECT  6815.0 42842.5 6950.0 42777.5 ;
      RECT  7072.5 43057.5 7207.5 42992.5 ;
      RECT  7167.5 42842.5 7302.5 42777.5 ;
      RECT  6755.0 42137.5 7675.0 42072.5 ;
      RECT  6755.0 43482.5 7675.0 43417.5 ;
      RECT  6822.5 43612.5 6887.5 43417.5 ;
      RECT  6822.5 44452.5 6887.5 44827.5 ;
      RECT  7202.5 44452.5 7267.5 44827.5 ;
      RECT  7372.5 44610.0 7437.5 44795.0 ;
      RECT  7372.5 43450.0 7437.5 43635.0 ;
      RECT  6822.5 44452.5 6887.5 44587.5 ;
      RECT  7012.5 44452.5 7077.5 44587.5 ;
      RECT  7012.5 44452.5 7077.5 44587.5 ;
      RECT  6822.5 44452.5 6887.5 44587.5 ;
      RECT  7012.5 44452.5 7077.5 44587.5 ;
      RECT  7202.5 44452.5 7267.5 44587.5 ;
      RECT  7202.5 44452.5 7267.5 44587.5 ;
      RECT  7012.5 44452.5 7077.5 44587.5 ;
      RECT  6822.5 43612.5 6887.5 43747.5 ;
      RECT  7012.5 43612.5 7077.5 43747.5 ;
      RECT  7012.5 43612.5 7077.5 43747.5 ;
      RECT  6822.5 43612.5 6887.5 43747.5 ;
      RECT  7012.5 43612.5 7077.5 43747.5 ;
      RECT  7202.5 43612.5 7267.5 43747.5 ;
      RECT  7202.5 43612.5 7267.5 43747.5 ;
      RECT  7012.5 43612.5 7077.5 43747.5 ;
      RECT  7372.5 44542.5 7437.5 44677.5 ;
      RECT  7372.5 43567.5 7437.5 43702.5 ;
      RECT  7207.5 43842.5 7072.5 43907.5 ;
      RECT  6950.0 44057.5 6815.0 44122.5 ;
      RECT  7012.5 44452.5 7077.5 44587.5 ;
      RECT  7202.5 43612.5 7267.5 43747.5 ;
      RECT  7302.5 44057.5 7167.5 44122.5 ;
      RECT  6815.0 44057.5 6950.0 44122.5 ;
      RECT  7072.5 43842.5 7207.5 43907.5 ;
      RECT  7167.5 44057.5 7302.5 44122.5 ;
      RECT  6755.0 44762.5 7675.0 44827.5 ;
      RECT  6755.0 43417.5 7675.0 43482.5 ;
      RECT  6822.5 45977.5 6887.5 46172.5 ;
      RECT  6822.5 45137.5 6887.5 44762.5 ;
      RECT  7202.5 45137.5 7267.5 44762.5 ;
      RECT  7372.5 44980.0 7437.5 44795.0 ;
      RECT  7372.5 46140.0 7437.5 45955.0 ;
      RECT  6822.5 45137.5 6887.5 45002.5 ;
      RECT  7012.5 45137.5 7077.5 45002.5 ;
      RECT  7012.5 45137.5 7077.5 45002.5 ;
      RECT  6822.5 45137.5 6887.5 45002.5 ;
      RECT  7012.5 45137.5 7077.5 45002.5 ;
      RECT  7202.5 45137.5 7267.5 45002.5 ;
      RECT  7202.5 45137.5 7267.5 45002.5 ;
      RECT  7012.5 45137.5 7077.5 45002.5 ;
      RECT  6822.5 45977.5 6887.5 45842.5 ;
      RECT  7012.5 45977.5 7077.5 45842.5 ;
      RECT  7012.5 45977.5 7077.5 45842.5 ;
      RECT  6822.5 45977.5 6887.5 45842.5 ;
      RECT  7012.5 45977.5 7077.5 45842.5 ;
      RECT  7202.5 45977.5 7267.5 45842.5 ;
      RECT  7202.5 45977.5 7267.5 45842.5 ;
      RECT  7012.5 45977.5 7077.5 45842.5 ;
      RECT  7372.5 45047.5 7437.5 44912.5 ;
      RECT  7372.5 46022.5 7437.5 45887.5 ;
      RECT  7207.5 45747.5 7072.5 45682.5 ;
      RECT  6950.0 45532.5 6815.0 45467.5 ;
      RECT  7012.5 45137.5 7077.5 45002.5 ;
      RECT  7202.5 45977.5 7267.5 45842.5 ;
      RECT  7302.5 45532.5 7167.5 45467.5 ;
      RECT  6815.0 45532.5 6950.0 45467.5 ;
      RECT  7072.5 45747.5 7207.5 45682.5 ;
      RECT  7167.5 45532.5 7302.5 45467.5 ;
      RECT  6755.0 44827.5 7675.0 44762.5 ;
      RECT  6755.0 46172.5 7675.0 46107.5 ;
      RECT  6822.5 46302.5 6887.5 46107.5 ;
      RECT  6822.5 47142.5 6887.5 47517.5 ;
      RECT  7202.5 47142.5 7267.5 47517.5 ;
      RECT  7372.5 47300.0 7437.5 47485.0 ;
      RECT  7372.5 46140.0 7437.5 46325.0 ;
      RECT  6822.5 47142.5 6887.5 47277.5 ;
      RECT  7012.5 47142.5 7077.5 47277.5 ;
      RECT  7012.5 47142.5 7077.5 47277.5 ;
      RECT  6822.5 47142.5 6887.5 47277.5 ;
      RECT  7012.5 47142.5 7077.5 47277.5 ;
      RECT  7202.5 47142.5 7267.5 47277.5 ;
      RECT  7202.5 47142.5 7267.5 47277.5 ;
      RECT  7012.5 47142.5 7077.5 47277.5 ;
      RECT  6822.5 46302.5 6887.5 46437.5 ;
      RECT  7012.5 46302.5 7077.5 46437.5 ;
      RECT  7012.5 46302.5 7077.5 46437.5 ;
      RECT  6822.5 46302.5 6887.5 46437.5 ;
      RECT  7012.5 46302.5 7077.5 46437.5 ;
      RECT  7202.5 46302.5 7267.5 46437.5 ;
      RECT  7202.5 46302.5 7267.5 46437.5 ;
      RECT  7012.5 46302.5 7077.5 46437.5 ;
      RECT  7372.5 47232.5 7437.5 47367.5 ;
      RECT  7372.5 46257.5 7437.5 46392.5 ;
      RECT  7207.5 46532.5 7072.5 46597.5 ;
      RECT  6950.0 46747.5 6815.0 46812.5 ;
      RECT  7012.5 47142.5 7077.5 47277.5 ;
      RECT  7202.5 46302.5 7267.5 46437.5 ;
      RECT  7302.5 46747.5 7167.5 46812.5 ;
      RECT  6815.0 46747.5 6950.0 46812.5 ;
      RECT  7072.5 46532.5 7207.5 46597.5 ;
      RECT  7167.5 46747.5 7302.5 46812.5 ;
      RECT  6755.0 47452.5 7675.0 47517.5 ;
      RECT  6755.0 46107.5 7675.0 46172.5 ;
      RECT  6822.5 48667.5 6887.5 48862.5 ;
      RECT  6822.5 47827.5 6887.5 47452.5 ;
      RECT  7202.5 47827.5 7267.5 47452.5 ;
      RECT  7372.5 47670.0 7437.5 47485.0 ;
      RECT  7372.5 48830.0 7437.5 48645.0 ;
      RECT  6822.5 47827.5 6887.5 47692.5 ;
      RECT  7012.5 47827.5 7077.5 47692.5 ;
      RECT  7012.5 47827.5 7077.5 47692.5 ;
      RECT  6822.5 47827.5 6887.5 47692.5 ;
      RECT  7012.5 47827.5 7077.5 47692.5 ;
      RECT  7202.5 47827.5 7267.5 47692.5 ;
      RECT  7202.5 47827.5 7267.5 47692.5 ;
      RECT  7012.5 47827.5 7077.5 47692.5 ;
      RECT  6822.5 48667.5 6887.5 48532.5 ;
      RECT  7012.5 48667.5 7077.5 48532.5 ;
      RECT  7012.5 48667.5 7077.5 48532.5 ;
      RECT  6822.5 48667.5 6887.5 48532.5 ;
      RECT  7012.5 48667.5 7077.5 48532.5 ;
      RECT  7202.5 48667.5 7267.5 48532.5 ;
      RECT  7202.5 48667.5 7267.5 48532.5 ;
      RECT  7012.5 48667.5 7077.5 48532.5 ;
      RECT  7372.5 47737.5 7437.5 47602.5 ;
      RECT  7372.5 48712.5 7437.5 48577.5 ;
      RECT  7207.5 48437.5 7072.5 48372.5 ;
      RECT  6950.0 48222.5 6815.0 48157.5 ;
      RECT  7012.5 47827.5 7077.5 47692.5 ;
      RECT  7202.5 48667.5 7267.5 48532.5 ;
      RECT  7302.5 48222.5 7167.5 48157.5 ;
      RECT  6815.0 48222.5 6950.0 48157.5 ;
      RECT  7072.5 48437.5 7207.5 48372.5 ;
      RECT  7167.5 48222.5 7302.5 48157.5 ;
      RECT  6755.0 47517.5 7675.0 47452.5 ;
      RECT  6755.0 48862.5 7675.0 48797.5 ;
      RECT  6822.5 48992.5 6887.5 48797.5 ;
      RECT  6822.5 49832.5 6887.5 50207.5 ;
      RECT  7202.5 49832.5 7267.5 50207.5 ;
      RECT  7372.5 49990.0 7437.5 50175.0 ;
      RECT  7372.5 48830.0 7437.5 49015.0 ;
      RECT  6822.5 49832.5 6887.5 49967.5 ;
      RECT  7012.5 49832.5 7077.5 49967.5 ;
      RECT  7012.5 49832.5 7077.5 49967.5 ;
      RECT  6822.5 49832.5 6887.5 49967.5 ;
      RECT  7012.5 49832.5 7077.5 49967.5 ;
      RECT  7202.5 49832.5 7267.5 49967.5 ;
      RECT  7202.5 49832.5 7267.5 49967.5 ;
      RECT  7012.5 49832.5 7077.5 49967.5 ;
      RECT  6822.5 48992.5 6887.5 49127.5 ;
      RECT  7012.5 48992.5 7077.5 49127.5 ;
      RECT  7012.5 48992.5 7077.5 49127.5 ;
      RECT  6822.5 48992.5 6887.5 49127.5 ;
      RECT  7012.5 48992.5 7077.5 49127.5 ;
      RECT  7202.5 48992.5 7267.5 49127.5 ;
      RECT  7202.5 48992.5 7267.5 49127.5 ;
      RECT  7012.5 48992.5 7077.5 49127.5 ;
      RECT  7372.5 49922.5 7437.5 50057.5 ;
      RECT  7372.5 48947.5 7437.5 49082.5 ;
      RECT  7207.5 49222.5 7072.5 49287.5 ;
      RECT  6950.0 49437.5 6815.0 49502.5 ;
      RECT  7012.5 49832.5 7077.5 49967.5 ;
      RECT  7202.5 48992.5 7267.5 49127.5 ;
      RECT  7302.5 49437.5 7167.5 49502.5 ;
      RECT  6815.0 49437.5 6950.0 49502.5 ;
      RECT  7072.5 49222.5 7207.5 49287.5 ;
      RECT  7167.5 49437.5 7302.5 49502.5 ;
      RECT  6755.0 50142.5 7675.0 50207.5 ;
      RECT  6755.0 48797.5 7675.0 48862.5 ;
      RECT  6822.5 51357.5 6887.5 51552.5 ;
      RECT  6822.5 50517.5 6887.5 50142.5 ;
      RECT  7202.5 50517.5 7267.5 50142.5 ;
      RECT  7372.5 50360.0 7437.5 50175.0 ;
      RECT  7372.5 51520.0 7437.5 51335.0 ;
      RECT  6822.5 50517.5 6887.5 50382.5 ;
      RECT  7012.5 50517.5 7077.5 50382.5 ;
      RECT  7012.5 50517.5 7077.5 50382.5 ;
      RECT  6822.5 50517.5 6887.5 50382.5 ;
      RECT  7012.5 50517.5 7077.5 50382.5 ;
      RECT  7202.5 50517.5 7267.5 50382.5 ;
      RECT  7202.5 50517.5 7267.5 50382.5 ;
      RECT  7012.5 50517.5 7077.5 50382.5 ;
      RECT  6822.5 51357.5 6887.5 51222.5 ;
      RECT  7012.5 51357.5 7077.5 51222.5 ;
      RECT  7012.5 51357.5 7077.5 51222.5 ;
      RECT  6822.5 51357.5 6887.5 51222.5 ;
      RECT  7012.5 51357.5 7077.5 51222.5 ;
      RECT  7202.5 51357.5 7267.5 51222.5 ;
      RECT  7202.5 51357.5 7267.5 51222.5 ;
      RECT  7012.5 51357.5 7077.5 51222.5 ;
      RECT  7372.5 50427.5 7437.5 50292.5 ;
      RECT  7372.5 51402.5 7437.5 51267.5 ;
      RECT  7207.5 51127.5 7072.5 51062.5 ;
      RECT  6950.0 50912.5 6815.0 50847.5 ;
      RECT  7012.5 50517.5 7077.5 50382.5 ;
      RECT  7202.5 51357.5 7267.5 51222.5 ;
      RECT  7302.5 50912.5 7167.5 50847.5 ;
      RECT  6815.0 50912.5 6950.0 50847.5 ;
      RECT  7072.5 51127.5 7207.5 51062.5 ;
      RECT  7167.5 50912.5 7302.5 50847.5 ;
      RECT  6755.0 50207.5 7675.0 50142.5 ;
      RECT  6755.0 51552.5 7675.0 51487.5 ;
      RECT  6822.5 51682.5 6887.5 51487.5 ;
      RECT  6822.5 52522.5 6887.5 52897.5 ;
      RECT  7202.5 52522.5 7267.5 52897.5 ;
      RECT  7372.5 52680.0 7437.5 52865.0 ;
      RECT  7372.5 51520.0 7437.5 51705.0 ;
      RECT  6822.5 52522.5 6887.5 52657.5 ;
      RECT  7012.5 52522.5 7077.5 52657.5 ;
      RECT  7012.5 52522.5 7077.5 52657.5 ;
      RECT  6822.5 52522.5 6887.5 52657.5 ;
      RECT  7012.5 52522.5 7077.5 52657.5 ;
      RECT  7202.5 52522.5 7267.5 52657.5 ;
      RECT  7202.5 52522.5 7267.5 52657.5 ;
      RECT  7012.5 52522.5 7077.5 52657.5 ;
      RECT  6822.5 51682.5 6887.5 51817.5 ;
      RECT  7012.5 51682.5 7077.5 51817.5 ;
      RECT  7012.5 51682.5 7077.5 51817.5 ;
      RECT  6822.5 51682.5 6887.5 51817.5 ;
      RECT  7012.5 51682.5 7077.5 51817.5 ;
      RECT  7202.5 51682.5 7267.5 51817.5 ;
      RECT  7202.5 51682.5 7267.5 51817.5 ;
      RECT  7012.5 51682.5 7077.5 51817.5 ;
      RECT  7372.5 52612.5 7437.5 52747.5 ;
      RECT  7372.5 51637.5 7437.5 51772.5 ;
      RECT  7207.5 51912.5 7072.5 51977.5 ;
      RECT  6950.0 52127.5 6815.0 52192.5 ;
      RECT  7012.5 52522.5 7077.5 52657.5 ;
      RECT  7202.5 51682.5 7267.5 51817.5 ;
      RECT  7302.5 52127.5 7167.5 52192.5 ;
      RECT  6815.0 52127.5 6950.0 52192.5 ;
      RECT  7072.5 51912.5 7207.5 51977.5 ;
      RECT  7167.5 52127.5 7302.5 52192.5 ;
      RECT  6755.0 52832.5 7675.0 52897.5 ;
      RECT  6755.0 51487.5 7675.0 51552.5 ;
      RECT  6822.5 54047.5 6887.5 54242.5 ;
      RECT  6822.5 53207.5 6887.5 52832.5 ;
      RECT  7202.5 53207.5 7267.5 52832.5 ;
      RECT  7372.5 53050.0 7437.5 52865.0 ;
      RECT  7372.5 54210.0 7437.5 54025.0 ;
      RECT  6822.5 53207.5 6887.5 53072.5 ;
      RECT  7012.5 53207.5 7077.5 53072.5 ;
      RECT  7012.5 53207.5 7077.5 53072.5 ;
      RECT  6822.5 53207.5 6887.5 53072.5 ;
      RECT  7012.5 53207.5 7077.5 53072.5 ;
      RECT  7202.5 53207.5 7267.5 53072.5 ;
      RECT  7202.5 53207.5 7267.5 53072.5 ;
      RECT  7012.5 53207.5 7077.5 53072.5 ;
      RECT  6822.5 54047.5 6887.5 53912.5 ;
      RECT  7012.5 54047.5 7077.5 53912.5 ;
      RECT  7012.5 54047.5 7077.5 53912.5 ;
      RECT  6822.5 54047.5 6887.5 53912.5 ;
      RECT  7012.5 54047.5 7077.5 53912.5 ;
      RECT  7202.5 54047.5 7267.5 53912.5 ;
      RECT  7202.5 54047.5 7267.5 53912.5 ;
      RECT  7012.5 54047.5 7077.5 53912.5 ;
      RECT  7372.5 53117.5 7437.5 52982.5 ;
      RECT  7372.5 54092.5 7437.5 53957.5 ;
      RECT  7207.5 53817.5 7072.5 53752.5 ;
      RECT  6950.0 53602.5 6815.0 53537.5 ;
      RECT  7012.5 53207.5 7077.5 53072.5 ;
      RECT  7202.5 54047.5 7267.5 53912.5 ;
      RECT  7302.5 53602.5 7167.5 53537.5 ;
      RECT  6815.0 53602.5 6950.0 53537.5 ;
      RECT  7072.5 53817.5 7207.5 53752.5 ;
      RECT  7167.5 53602.5 7302.5 53537.5 ;
      RECT  6755.0 52897.5 7675.0 52832.5 ;
      RECT  6755.0 54242.5 7675.0 54177.5 ;
      RECT  6822.5 54372.5 6887.5 54177.5 ;
      RECT  6822.5 55212.5 6887.5 55587.5 ;
      RECT  7202.5 55212.5 7267.5 55587.5 ;
      RECT  7372.5 55370.0 7437.5 55555.0 ;
      RECT  7372.5 54210.0 7437.5 54395.0 ;
      RECT  6822.5 55212.5 6887.5 55347.5 ;
      RECT  7012.5 55212.5 7077.5 55347.5 ;
      RECT  7012.5 55212.5 7077.5 55347.5 ;
      RECT  6822.5 55212.5 6887.5 55347.5 ;
      RECT  7012.5 55212.5 7077.5 55347.5 ;
      RECT  7202.5 55212.5 7267.5 55347.5 ;
      RECT  7202.5 55212.5 7267.5 55347.5 ;
      RECT  7012.5 55212.5 7077.5 55347.5 ;
      RECT  6822.5 54372.5 6887.5 54507.5 ;
      RECT  7012.5 54372.5 7077.5 54507.5 ;
      RECT  7012.5 54372.5 7077.5 54507.5 ;
      RECT  6822.5 54372.5 6887.5 54507.5 ;
      RECT  7012.5 54372.5 7077.5 54507.5 ;
      RECT  7202.5 54372.5 7267.5 54507.5 ;
      RECT  7202.5 54372.5 7267.5 54507.5 ;
      RECT  7012.5 54372.5 7077.5 54507.5 ;
      RECT  7372.5 55302.5 7437.5 55437.5 ;
      RECT  7372.5 54327.5 7437.5 54462.5 ;
      RECT  7207.5 54602.5 7072.5 54667.5 ;
      RECT  6950.0 54817.5 6815.0 54882.5 ;
      RECT  7012.5 55212.5 7077.5 55347.5 ;
      RECT  7202.5 54372.5 7267.5 54507.5 ;
      RECT  7302.5 54817.5 7167.5 54882.5 ;
      RECT  6815.0 54817.5 6950.0 54882.5 ;
      RECT  7072.5 54602.5 7207.5 54667.5 ;
      RECT  7167.5 54817.5 7302.5 54882.5 ;
      RECT  6755.0 55522.5 7675.0 55587.5 ;
      RECT  6755.0 54177.5 7675.0 54242.5 ;
      RECT  6822.5 56737.5 6887.5 56932.5 ;
      RECT  6822.5 55897.5 6887.5 55522.5 ;
      RECT  7202.5 55897.5 7267.5 55522.5 ;
      RECT  7372.5 55740.0 7437.5 55555.0 ;
      RECT  7372.5 56900.0 7437.5 56715.0 ;
      RECT  6822.5 55897.5 6887.5 55762.5 ;
      RECT  7012.5 55897.5 7077.5 55762.5 ;
      RECT  7012.5 55897.5 7077.5 55762.5 ;
      RECT  6822.5 55897.5 6887.5 55762.5 ;
      RECT  7012.5 55897.5 7077.5 55762.5 ;
      RECT  7202.5 55897.5 7267.5 55762.5 ;
      RECT  7202.5 55897.5 7267.5 55762.5 ;
      RECT  7012.5 55897.5 7077.5 55762.5 ;
      RECT  6822.5 56737.5 6887.5 56602.5 ;
      RECT  7012.5 56737.5 7077.5 56602.5 ;
      RECT  7012.5 56737.5 7077.5 56602.5 ;
      RECT  6822.5 56737.5 6887.5 56602.5 ;
      RECT  7012.5 56737.5 7077.5 56602.5 ;
      RECT  7202.5 56737.5 7267.5 56602.5 ;
      RECT  7202.5 56737.5 7267.5 56602.5 ;
      RECT  7012.5 56737.5 7077.5 56602.5 ;
      RECT  7372.5 55807.5 7437.5 55672.5 ;
      RECT  7372.5 56782.5 7437.5 56647.5 ;
      RECT  7207.5 56507.5 7072.5 56442.5 ;
      RECT  6950.0 56292.5 6815.0 56227.5 ;
      RECT  7012.5 55897.5 7077.5 55762.5 ;
      RECT  7202.5 56737.5 7267.5 56602.5 ;
      RECT  7302.5 56292.5 7167.5 56227.5 ;
      RECT  6815.0 56292.5 6950.0 56227.5 ;
      RECT  7072.5 56507.5 7207.5 56442.5 ;
      RECT  7167.5 56292.5 7302.5 56227.5 ;
      RECT  6755.0 55587.5 7675.0 55522.5 ;
      RECT  6755.0 56932.5 7675.0 56867.5 ;
      RECT  6822.5 57062.5 6887.5 56867.5 ;
      RECT  6822.5 57902.5 6887.5 58277.5 ;
      RECT  7202.5 57902.5 7267.5 58277.5 ;
      RECT  7372.5 58060.0 7437.5 58245.0 ;
      RECT  7372.5 56900.0 7437.5 57085.0 ;
      RECT  6822.5 57902.5 6887.5 58037.5 ;
      RECT  7012.5 57902.5 7077.5 58037.5 ;
      RECT  7012.5 57902.5 7077.5 58037.5 ;
      RECT  6822.5 57902.5 6887.5 58037.5 ;
      RECT  7012.5 57902.5 7077.5 58037.5 ;
      RECT  7202.5 57902.5 7267.5 58037.5 ;
      RECT  7202.5 57902.5 7267.5 58037.5 ;
      RECT  7012.5 57902.5 7077.5 58037.5 ;
      RECT  6822.5 57062.5 6887.5 57197.5 ;
      RECT  7012.5 57062.5 7077.5 57197.5 ;
      RECT  7012.5 57062.5 7077.5 57197.5 ;
      RECT  6822.5 57062.5 6887.5 57197.5 ;
      RECT  7012.5 57062.5 7077.5 57197.5 ;
      RECT  7202.5 57062.5 7267.5 57197.5 ;
      RECT  7202.5 57062.5 7267.5 57197.5 ;
      RECT  7012.5 57062.5 7077.5 57197.5 ;
      RECT  7372.5 57992.5 7437.5 58127.5 ;
      RECT  7372.5 57017.5 7437.5 57152.5 ;
      RECT  7207.5 57292.5 7072.5 57357.5 ;
      RECT  6950.0 57507.5 6815.0 57572.5 ;
      RECT  7012.5 57902.5 7077.5 58037.5 ;
      RECT  7202.5 57062.5 7267.5 57197.5 ;
      RECT  7302.5 57507.5 7167.5 57572.5 ;
      RECT  6815.0 57507.5 6950.0 57572.5 ;
      RECT  7072.5 57292.5 7207.5 57357.5 ;
      RECT  7167.5 57507.5 7302.5 57572.5 ;
      RECT  6755.0 58212.5 7675.0 58277.5 ;
      RECT  6755.0 56867.5 7675.0 56932.5 ;
      RECT  6822.5 59427.5 6887.5 59622.5 ;
      RECT  6822.5 58587.5 6887.5 58212.5 ;
      RECT  7202.5 58587.5 7267.5 58212.5 ;
      RECT  7372.5 58430.0 7437.5 58245.0 ;
      RECT  7372.5 59590.0 7437.5 59405.0 ;
      RECT  6822.5 58587.5 6887.5 58452.5 ;
      RECT  7012.5 58587.5 7077.5 58452.5 ;
      RECT  7012.5 58587.5 7077.5 58452.5 ;
      RECT  6822.5 58587.5 6887.5 58452.5 ;
      RECT  7012.5 58587.5 7077.5 58452.5 ;
      RECT  7202.5 58587.5 7267.5 58452.5 ;
      RECT  7202.5 58587.5 7267.5 58452.5 ;
      RECT  7012.5 58587.5 7077.5 58452.5 ;
      RECT  6822.5 59427.5 6887.5 59292.5 ;
      RECT  7012.5 59427.5 7077.5 59292.5 ;
      RECT  7012.5 59427.5 7077.5 59292.5 ;
      RECT  6822.5 59427.5 6887.5 59292.5 ;
      RECT  7012.5 59427.5 7077.5 59292.5 ;
      RECT  7202.5 59427.5 7267.5 59292.5 ;
      RECT  7202.5 59427.5 7267.5 59292.5 ;
      RECT  7012.5 59427.5 7077.5 59292.5 ;
      RECT  7372.5 58497.5 7437.5 58362.5 ;
      RECT  7372.5 59472.5 7437.5 59337.5 ;
      RECT  7207.5 59197.5 7072.5 59132.5 ;
      RECT  6950.0 58982.5 6815.0 58917.5 ;
      RECT  7012.5 58587.5 7077.5 58452.5 ;
      RECT  7202.5 59427.5 7267.5 59292.5 ;
      RECT  7302.5 58982.5 7167.5 58917.5 ;
      RECT  6815.0 58982.5 6950.0 58917.5 ;
      RECT  7072.5 59197.5 7207.5 59132.5 ;
      RECT  7167.5 58982.5 7302.5 58917.5 ;
      RECT  6755.0 58277.5 7675.0 58212.5 ;
      RECT  6755.0 59622.5 7675.0 59557.5 ;
      RECT  6822.5 59752.5 6887.5 59557.5 ;
      RECT  6822.5 60592.5 6887.5 60967.5 ;
      RECT  7202.5 60592.5 7267.5 60967.5 ;
      RECT  7372.5 60750.0 7437.5 60935.0 ;
      RECT  7372.5 59590.0 7437.5 59775.0 ;
      RECT  6822.5 60592.5 6887.5 60727.5 ;
      RECT  7012.5 60592.5 7077.5 60727.5 ;
      RECT  7012.5 60592.5 7077.5 60727.5 ;
      RECT  6822.5 60592.5 6887.5 60727.5 ;
      RECT  7012.5 60592.5 7077.5 60727.5 ;
      RECT  7202.5 60592.5 7267.5 60727.5 ;
      RECT  7202.5 60592.5 7267.5 60727.5 ;
      RECT  7012.5 60592.5 7077.5 60727.5 ;
      RECT  6822.5 59752.5 6887.5 59887.5 ;
      RECT  7012.5 59752.5 7077.5 59887.5 ;
      RECT  7012.5 59752.5 7077.5 59887.5 ;
      RECT  6822.5 59752.5 6887.5 59887.5 ;
      RECT  7012.5 59752.5 7077.5 59887.5 ;
      RECT  7202.5 59752.5 7267.5 59887.5 ;
      RECT  7202.5 59752.5 7267.5 59887.5 ;
      RECT  7012.5 59752.5 7077.5 59887.5 ;
      RECT  7372.5 60682.5 7437.5 60817.5 ;
      RECT  7372.5 59707.5 7437.5 59842.5 ;
      RECT  7207.5 59982.5 7072.5 60047.5 ;
      RECT  6950.0 60197.5 6815.0 60262.5 ;
      RECT  7012.5 60592.5 7077.5 60727.5 ;
      RECT  7202.5 59752.5 7267.5 59887.5 ;
      RECT  7302.5 60197.5 7167.5 60262.5 ;
      RECT  6815.0 60197.5 6950.0 60262.5 ;
      RECT  7072.5 59982.5 7207.5 60047.5 ;
      RECT  7167.5 60197.5 7302.5 60262.5 ;
      RECT  6755.0 60902.5 7675.0 60967.5 ;
      RECT  6755.0 59557.5 7675.0 59622.5 ;
      RECT  6822.5 62117.5 6887.5 62312.5 ;
      RECT  6822.5 61277.5 6887.5 60902.5 ;
      RECT  7202.5 61277.5 7267.5 60902.5 ;
      RECT  7372.5 61120.0 7437.5 60935.0 ;
      RECT  7372.5 62280.0 7437.5 62095.0 ;
      RECT  6822.5 61277.5 6887.5 61142.5 ;
      RECT  7012.5 61277.5 7077.5 61142.5 ;
      RECT  7012.5 61277.5 7077.5 61142.5 ;
      RECT  6822.5 61277.5 6887.5 61142.5 ;
      RECT  7012.5 61277.5 7077.5 61142.5 ;
      RECT  7202.5 61277.5 7267.5 61142.5 ;
      RECT  7202.5 61277.5 7267.5 61142.5 ;
      RECT  7012.5 61277.5 7077.5 61142.5 ;
      RECT  6822.5 62117.5 6887.5 61982.5 ;
      RECT  7012.5 62117.5 7077.5 61982.5 ;
      RECT  7012.5 62117.5 7077.5 61982.5 ;
      RECT  6822.5 62117.5 6887.5 61982.5 ;
      RECT  7012.5 62117.5 7077.5 61982.5 ;
      RECT  7202.5 62117.5 7267.5 61982.5 ;
      RECT  7202.5 62117.5 7267.5 61982.5 ;
      RECT  7012.5 62117.5 7077.5 61982.5 ;
      RECT  7372.5 61187.5 7437.5 61052.5 ;
      RECT  7372.5 62162.5 7437.5 62027.5 ;
      RECT  7207.5 61887.5 7072.5 61822.5 ;
      RECT  6950.0 61672.5 6815.0 61607.5 ;
      RECT  7012.5 61277.5 7077.5 61142.5 ;
      RECT  7202.5 62117.5 7267.5 61982.5 ;
      RECT  7302.5 61672.5 7167.5 61607.5 ;
      RECT  6815.0 61672.5 6950.0 61607.5 ;
      RECT  7072.5 61887.5 7207.5 61822.5 ;
      RECT  7167.5 61672.5 7302.5 61607.5 ;
      RECT  6755.0 60967.5 7675.0 60902.5 ;
      RECT  6755.0 62312.5 7675.0 62247.5 ;
      RECT  6822.5 62442.5 6887.5 62247.5 ;
      RECT  6822.5 63282.5 6887.5 63657.5 ;
      RECT  7202.5 63282.5 7267.5 63657.5 ;
      RECT  7372.5 63440.0 7437.5 63625.0 ;
      RECT  7372.5 62280.0 7437.5 62465.0 ;
      RECT  6822.5 63282.5 6887.5 63417.5 ;
      RECT  7012.5 63282.5 7077.5 63417.5 ;
      RECT  7012.5 63282.5 7077.5 63417.5 ;
      RECT  6822.5 63282.5 6887.5 63417.5 ;
      RECT  7012.5 63282.5 7077.5 63417.5 ;
      RECT  7202.5 63282.5 7267.5 63417.5 ;
      RECT  7202.5 63282.5 7267.5 63417.5 ;
      RECT  7012.5 63282.5 7077.5 63417.5 ;
      RECT  6822.5 62442.5 6887.5 62577.5 ;
      RECT  7012.5 62442.5 7077.5 62577.5 ;
      RECT  7012.5 62442.5 7077.5 62577.5 ;
      RECT  6822.5 62442.5 6887.5 62577.5 ;
      RECT  7012.5 62442.5 7077.5 62577.5 ;
      RECT  7202.5 62442.5 7267.5 62577.5 ;
      RECT  7202.5 62442.5 7267.5 62577.5 ;
      RECT  7012.5 62442.5 7077.5 62577.5 ;
      RECT  7372.5 63372.5 7437.5 63507.5 ;
      RECT  7372.5 62397.5 7437.5 62532.5 ;
      RECT  7207.5 62672.5 7072.5 62737.5 ;
      RECT  6950.0 62887.5 6815.0 62952.5 ;
      RECT  7012.5 63282.5 7077.5 63417.5 ;
      RECT  7202.5 62442.5 7267.5 62577.5 ;
      RECT  7302.5 62887.5 7167.5 62952.5 ;
      RECT  6815.0 62887.5 6950.0 62952.5 ;
      RECT  7072.5 62672.5 7207.5 62737.5 ;
      RECT  7167.5 62887.5 7302.5 62952.5 ;
      RECT  6755.0 63592.5 7675.0 63657.5 ;
      RECT  6755.0 62247.5 7675.0 62312.5 ;
      RECT  6822.5 64807.5 6887.5 65002.5 ;
      RECT  6822.5 63967.5 6887.5 63592.5 ;
      RECT  7202.5 63967.5 7267.5 63592.5 ;
      RECT  7372.5 63810.0 7437.5 63625.0 ;
      RECT  7372.5 64970.0 7437.5 64785.0 ;
      RECT  6822.5 63967.5 6887.5 63832.5 ;
      RECT  7012.5 63967.5 7077.5 63832.5 ;
      RECT  7012.5 63967.5 7077.5 63832.5 ;
      RECT  6822.5 63967.5 6887.5 63832.5 ;
      RECT  7012.5 63967.5 7077.5 63832.5 ;
      RECT  7202.5 63967.5 7267.5 63832.5 ;
      RECT  7202.5 63967.5 7267.5 63832.5 ;
      RECT  7012.5 63967.5 7077.5 63832.5 ;
      RECT  6822.5 64807.5 6887.5 64672.5 ;
      RECT  7012.5 64807.5 7077.5 64672.5 ;
      RECT  7012.5 64807.5 7077.5 64672.5 ;
      RECT  6822.5 64807.5 6887.5 64672.5 ;
      RECT  7012.5 64807.5 7077.5 64672.5 ;
      RECT  7202.5 64807.5 7267.5 64672.5 ;
      RECT  7202.5 64807.5 7267.5 64672.5 ;
      RECT  7012.5 64807.5 7077.5 64672.5 ;
      RECT  7372.5 63877.5 7437.5 63742.5 ;
      RECT  7372.5 64852.5 7437.5 64717.5 ;
      RECT  7207.5 64577.5 7072.5 64512.5 ;
      RECT  6950.0 64362.5 6815.0 64297.5 ;
      RECT  7012.5 63967.5 7077.5 63832.5 ;
      RECT  7202.5 64807.5 7267.5 64672.5 ;
      RECT  7302.5 64362.5 7167.5 64297.5 ;
      RECT  6815.0 64362.5 6950.0 64297.5 ;
      RECT  7072.5 64577.5 7207.5 64512.5 ;
      RECT  7167.5 64362.5 7302.5 64297.5 ;
      RECT  6755.0 63657.5 7675.0 63592.5 ;
      RECT  6755.0 65002.5 7675.0 64937.5 ;
      RECT  6822.5 65132.5 6887.5 64937.5 ;
      RECT  6822.5 65972.5 6887.5 66347.5 ;
      RECT  7202.5 65972.5 7267.5 66347.5 ;
      RECT  7372.5 66130.0 7437.5 66315.0 ;
      RECT  7372.5 64970.0 7437.5 65155.0 ;
      RECT  6822.5 65972.5 6887.5 66107.5 ;
      RECT  7012.5 65972.5 7077.5 66107.5 ;
      RECT  7012.5 65972.5 7077.5 66107.5 ;
      RECT  6822.5 65972.5 6887.5 66107.5 ;
      RECT  7012.5 65972.5 7077.5 66107.5 ;
      RECT  7202.5 65972.5 7267.5 66107.5 ;
      RECT  7202.5 65972.5 7267.5 66107.5 ;
      RECT  7012.5 65972.5 7077.5 66107.5 ;
      RECT  6822.5 65132.5 6887.5 65267.5 ;
      RECT  7012.5 65132.5 7077.5 65267.5 ;
      RECT  7012.5 65132.5 7077.5 65267.5 ;
      RECT  6822.5 65132.5 6887.5 65267.5 ;
      RECT  7012.5 65132.5 7077.5 65267.5 ;
      RECT  7202.5 65132.5 7267.5 65267.5 ;
      RECT  7202.5 65132.5 7267.5 65267.5 ;
      RECT  7012.5 65132.5 7077.5 65267.5 ;
      RECT  7372.5 66062.5 7437.5 66197.5 ;
      RECT  7372.5 65087.5 7437.5 65222.5 ;
      RECT  7207.5 65362.5 7072.5 65427.5 ;
      RECT  6950.0 65577.5 6815.0 65642.5 ;
      RECT  7012.5 65972.5 7077.5 66107.5 ;
      RECT  7202.5 65132.5 7267.5 65267.5 ;
      RECT  7302.5 65577.5 7167.5 65642.5 ;
      RECT  6815.0 65577.5 6950.0 65642.5 ;
      RECT  7072.5 65362.5 7207.5 65427.5 ;
      RECT  7167.5 65577.5 7302.5 65642.5 ;
      RECT  6755.0 66282.5 7675.0 66347.5 ;
      RECT  6755.0 64937.5 7675.0 65002.5 ;
      RECT  6822.5 67497.5 6887.5 67692.5 ;
      RECT  6822.5 66657.5 6887.5 66282.5 ;
      RECT  7202.5 66657.5 7267.5 66282.5 ;
      RECT  7372.5 66500.0 7437.5 66315.0 ;
      RECT  7372.5 67660.0 7437.5 67475.0 ;
      RECT  6822.5 66657.5 6887.5 66522.5 ;
      RECT  7012.5 66657.5 7077.5 66522.5 ;
      RECT  7012.5 66657.5 7077.5 66522.5 ;
      RECT  6822.5 66657.5 6887.5 66522.5 ;
      RECT  7012.5 66657.5 7077.5 66522.5 ;
      RECT  7202.5 66657.5 7267.5 66522.5 ;
      RECT  7202.5 66657.5 7267.5 66522.5 ;
      RECT  7012.5 66657.5 7077.5 66522.5 ;
      RECT  6822.5 67497.5 6887.5 67362.5 ;
      RECT  7012.5 67497.5 7077.5 67362.5 ;
      RECT  7012.5 67497.5 7077.5 67362.5 ;
      RECT  6822.5 67497.5 6887.5 67362.5 ;
      RECT  7012.5 67497.5 7077.5 67362.5 ;
      RECT  7202.5 67497.5 7267.5 67362.5 ;
      RECT  7202.5 67497.5 7267.5 67362.5 ;
      RECT  7012.5 67497.5 7077.5 67362.5 ;
      RECT  7372.5 66567.5 7437.5 66432.5 ;
      RECT  7372.5 67542.5 7437.5 67407.5 ;
      RECT  7207.5 67267.5 7072.5 67202.5 ;
      RECT  6950.0 67052.5 6815.0 66987.5 ;
      RECT  7012.5 66657.5 7077.5 66522.5 ;
      RECT  7202.5 67497.5 7267.5 67362.5 ;
      RECT  7302.5 67052.5 7167.5 66987.5 ;
      RECT  6815.0 67052.5 6950.0 66987.5 ;
      RECT  7072.5 67267.5 7207.5 67202.5 ;
      RECT  7167.5 67052.5 7302.5 66987.5 ;
      RECT  6755.0 66347.5 7675.0 66282.5 ;
      RECT  6755.0 67692.5 7675.0 67627.5 ;
      RECT  6822.5 67822.5 6887.5 67627.5 ;
      RECT  6822.5 68662.5 6887.5 69037.5 ;
      RECT  7202.5 68662.5 7267.5 69037.5 ;
      RECT  7372.5 68820.0 7437.5 69005.0 ;
      RECT  7372.5 67660.0 7437.5 67845.0 ;
      RECT  6822.5 68662.5 6887.5 68797.5 ;
      RECT  7012.5 68662.5 7077.5 68797.5 ;
      RECT  7012.5 68662.5 7077.5 68797.5 ;
      RECT  6822.5 68662.5 6887.5 68797.5 ;
      RECT  7012.5 68662.5 7077.5 68797.5 ;
      RECT  7202.5 68662.5 7267.5 68797.5 ;
      RECT  7202.5 68662.5 7267.5 68797.5 ;
      RECT  7012.5 68662.5 7077.5 68797.5 ;
      RECT  6822.5 67822.5 6887.5 67957.5 ;
      RECT  7012.5 67822.5 7077.5 67957.5 ;
      RECT  7012.5 67822.5 7077.5 67957.5 ;
      RECT  6822.5 67822.5 6887.5 67957.5 ;
      RECT  7012.5 67822.5 7077.5 67957.5 ;
      RECT  7202.5 67822.5 7267.5 67957.5 ;
      RECT  7202.5 67822.5 7267.5 67957.5 ;
      RECT  7012.5 67822.5 7077.5 67957.5 ;
      RECT  7372.5 68752.5 7437.5 68887.5 ;
      RECT  7372.5 67777.5 7437.5 67912.5 ;
      RECT  7207.5 68052.5 7072.5 68117.5 ;
      RECT  6950.0 68267.5 6815.0 68332.5 ;
      RECT  7012.5 68662.5 7077.5 68797.5 ;
      RECT  7202.5 67822.5 7267.5 67957.5 ;
      RECT  7302.5 68267.5 7167.5 68332.5 ;
      RECT  6815.0 68267.5 6950.0 68332.5 ;
      RECT  7072.5 68052.5 7207.5 68117.5 ;
      RECT  7167.5 68267.5 7302.5 68332.5 ;
      RECT  6755.0 68972.5 7675.0 69037.5 ;
      RECT  6755.0 67627.5 7675.0 67692.5 ;
      RECT  6822.5 70187.5 6887.5 70382.5 ;
      RECT  6822.5 69347.5 6887.5 68972.5 ;
      RECT  7202.5 69347.5 7267.5 68972.5 ;
      RECT  7372.5 69190.0 7437.5 69005.0 ;
      RECT  7372.5 70350.0 7437.5 70165.0 ;
      RECT  6822.5 69347.5 6887.5 69212.5 ;
      RECT  7012.5 69347.5 7077.5 69212.5 ;
      RECT  7012.5 69347.5 7077.5 69212.5 ;
      RECT  6822.5 69347.5 6887.5 69212.5 ;
      RECT  7012.5 69347.5 7077.5 69212.5 ;
      RECT  7202.5 69347.5 7267.5 69212.5 ;
      RECT  7202.5 69347.5 7267.5 69212.5 ;
      RECT  7012.5 69347.5 7077.5 69212.5 ;
      RECT  6822.5 70187.5 6887.5 70052.5 ;
      RECT  7012.5 70187.5 7077.5 70052.5 ;
      RECT  7012.5 70187.5 7077.5 70052.5 ;
      RECT  6822.5 70187.5 6887.5 70052.5 ;
      RECT  7012.5 70187.5 7077.5 70052.5 ;
      RECT  7202.5 70187.5 7267.5 70052.5 ;
      RECT  7202.5 70187.5 7267.5 70052.5 ;
      RECT  7012.5 70187.5 7077.5 70052.5 ;
      RECT  7372.5 69257.5 7437.5 69122.5 ;
      RECT  7372.5 70232.5 7437.5 70097.5 ;
      RECT  7207.5 69957.5 7072.5 69892.5 ;
      RECT  6950.0 69742.5 6815.0 69677.5 ;
      RECT  7012.5 69347.5 7077.5 69212.5 ;
      RECT  7202.5 70187.5 7267.5 70052.5 ;
      RECT  7302.5 69742.5 7167.5 69677.5 ;
      RECT  6815.0 69742.5 6950.0 69677.5 ;
      RECT  7072.5 69957.5 7207.5 69892.5 ;
      RECT  7167.5 69742.5 7302.5 69677.5 ;
      RECT  6755.0 69037.5 7675.0 68972.5 ;
      RECT  6755.0 70382.5 7675.0 70317.5 ;
      RECT  8102.5 28470.0 8167.5 28655.0 ;
      RECT  8102.5 27310.0 8167.5 27495.0 ;
      RECT  7742.5 27427.5 7807.5 27277.5 ;
      RECT  7742.5 28312.5 7807.5 28687.5 ;
      RECT  7932.5 27427.5 7997.5 28312.5 ;
      RECT  7742.5 28312.5 7807.5 28447.5 ;
      RECT  7932.5 28312.5 7997.5 28447.5 ;
      RECT  7932.5 28312.5 7997.5 28447.5 ;
      RECT  7742.5 28312.5 7807.5 28447.5 ;
      RECT  7742.5 27427.5 7807.5 27562.5 ;
      RECT  7932.5 27427.5 7997.5 27562.5 ;
      RECT  7932.5 27427.5 7997.5 27562.5 ;
      RECT  7742.5 27427.5 7807.5 27562.5 ;
      RECT  8102.5 28402.5 8167.5 28537.5 ;
      RECT  8102.5 27427.5 8167.5 27562.5 ;
      RECT  7800.0 27870.0 7865.0 28005.0 ;
      RECT  7800.0 27870.0 7865.0 28005.0 ;
      RECT  7965.0 27905.0 8030.0 27970.0 ;
      RECT  7675.0 28622.5 8235.0 28687.5 ;
      RECT  7675.0 27277.5 8235.0 27342.5 ;
      RECT  8102.5 28840.0 8167.5 28655.0 ;
      RECT  8102.5 30000.0 8167.5 29815.0 ;
      RECT  7742.5 29882.5 7807.5 30032.5 ;
      RECT  7742.5 28997.5 7807.5 28622.5 ;
      RECT  7932.5 29882.5 7997.5 28997.5 ;
      RECT  7742.5 28997.5 7807.5 28862.5 ;
      RECT  7932.5 28997.5 7997.5 28862.5 ;
      RECT  7932.5 28997.5 7997.5 28862.5 ;
      RECT  7742.5 28997.5 7807.5 28862.5 ;
      RECT  7742.5 29882.5 7807.5 29747.5 ;
      RECT  7932.5 29882.5 7997.5 29747.5 ;
      RECT  7932.5 29882.5 7997.5 29747.5 ;
      RECT  7742.5 29882.5 7807.5 29747.5 ;
      RECT  8102.5 28907.5 8167.5 28772.5 ;
      RECT  8102.5 29882.5 8167.5 29747.5 ;
      RECT  7800.0 29440.0 7865.0 29305.0 ;
      RECT  7800.0 29440.0 7865.0 29305.0 ;
      RECT  7965.0 29405.0 8030.0 29340.0 ;
      RECT  7675.0 28687.5 8235.0 28622.5 ;
      RECT  7675.0 30032.5 8235.0 29967.5 ;
      RECT  8102.5 31160.0 8167.5 31345.0 ;
      RECT  8102.5 30000.0 8167.5 30185.0 ;
      RECT  7742.5 30117.5 7807.5 29967.5 ;
      RECT  7742.5 31002.5 7807.5 31377.5 ;
      RECT  7932.5 30117.5 7997.5 31002.5 ;
      RECT  7742.5 31002.5 7807.5 31137.5 ;
      RECT  7932.5 31002.5 7997.5 31137.5 ;
      RECT  7932.5 31002.5 7997.5 31137.5 ;
      RECT  7742.5 31002.5 7807.5 31137.5 ;
      RECT  7742.5 30117.5 7807.5 30252.5 ;
      RECT  7932.5 30117.5 7997.5 30252.5 ;
      RECT  7932.5 30117.5 7997.5 30252.5 ;
      RECT  7742.5 30117.5 7807.5 30252.5 ;
      RECT  8102.5 31092.5 8167.5 31227.5 ;
      RECT  8102.5 30117.5 8167.5 30252.5 ;
      RECT  7800.0 30560.0 7865.0 30695.0 ;
      RECT  7800.0 30560.0 7865.0 30695.0 ;
      RECT  7965.0 30595.0 8030.0 30660.0 ;
      RECT  7675.0 31312.5 8235.0 31377.5 ;
      RECT  7675.0 29967.5 8235.0 30032.5 ;
      RECT  8102.5 31530.0 8167.5 31345.0 ;
      RECT  8102.5 32690.0 8167.5 32505.0 ;
      RECT  7742.5 32572.5 7807.5 32722.5 ;
      RECT  7742.5 31687.5 7807.5 31312.5 ;
      RECT  7932.5 32572.5 7997.5 31687.5 ;
      RECT  7742.5 31687.5 7807.5 31552.5 ;
      RECT  7932.5 31687.5 7997.5 31552.5 ;
      RECT  7932.5 31687.5 7997.5 31552.5 ;
      RECT  7742.5 31687.5 7807.5 31552.5 ;
      RECT  7742.5 32572.5 7807.5 32437.5 ;
      RECT  7932.5 32572.5 7997.5 32437.5 ;
      RECT  7932.5 32572.5 7997.5 32437.5 ;
      RECT  7742.5 32572.5 7807.5 32437.5 ;
      RECT  8102.5 31597.5 8167.5 31462.5 ;
      RECT  8102.5 32572.5 8167.5 32437.5 ;
      RECT  7800.0 32130.0 7865.0 31995.0 ;
      RECT  7800.0 32130.0 7865.0 31995.0 ;
      RECT  7965.0 32095.0 8030.0 32030.0 ;
      RECT  7675.0 31377.5 8235.0 31312.5 ;
      RECT  7675.0 32722.5 8235.0 32657.5 ;
      RECT  8102.5 33850.0 8167.5 34035.0 ;
      RECT  8102.5 32690.0 8167.5 32875.0 ;
      RECT  7742.5 32807.5 7807.5 32657.5 ;
      RECT  7742.5 33692.5 7807.5 34067.5 ;
      RECT  7932.5 32807.5 7997.5 33692.5 ;
      RECT  7742.5 33692.5 7807.5 33827.5 ;
      RECT  7932.5 33692.5 7997.5 33827.5 ;
      RECT  7932.5 33692.5 7997.5 33827.5 ;
      RECT  7742.5 33692.5 7807.5 33827.5 ;
      RECT  7742.5 32807.5 7807.5 32942.5 ;
      RECT  7932.5 32807.5 7997.5 32942.5 ;
      RECT  7932.5 32807.5 7997.5 32942.5 ;
      RECT  7742.5 32807.5 7807.5 32942.5 ;
      RECT  8102.5 33782.5 8167.5 33917.5 ;
      RECT  8102.5 32807.5 8167.5 32942.5 ;
      RECT  7800.0 33250.0 7865.0 33385.0 ;
      RECT  7800.0 33250.0 7865.0 33385.0 ;
      RECT  7965.0 33285.0 8030.0 33350.0 ;
      RECT  7675.0 34002.5 8235.0 34067.5 ;
      RECT  7675.0 32657.5 8235.0 32722.5 ;
      RECT  8102.5 34220.0 8167.5 34035.0 ;
      RECT  8102.5 35380.0 8167.5 35195.0 ;
      RECT  7742.5 35262.5 7807.5 35412.5 ;
      RECT  7742.5 34377.5 7807.5 34002.5 ;
      RECT  7932.5 35262.5 7997.5 34377.5 ;
      RECT  7742.5 34377.5 7807.5 34242.5 ;
      RECT  7932.5 34377.5 7997.5 34242.5 ;
      RECT  7932.5 34377.5 7997.5 34242.5 ;
      RECT  7742.5 34377.5 7807.5 34242.5 ;
      RECT  7742.5 35262.5 7807.5 35127.5 ;
      RECT  7932.5 35262.5 7997.5 35127.5 ;
      RECT  7932.5 35262.5 7997.5 35127.5 ;
      RECT  7742.5 35262.5 7807.5 35127.5 ;
      RECT  8102.5 34287.5 8167.5 34152.5 ;
      RECT  8102.5 35262.5 8167.5 35127.5 ;
      RECT  7800.0 34820.0 7865.0 34685.0 ;
      RECT  7800.0 34820.0 7865.0 34685.0 ;
      RECT  7965.0 34785.0 8030.0 34720.0 ;
      RECT  7675.0 34067.5 8235.0 34002.5 ;
      RECT  7675.0 35412.5 8235.0 35347.5 ;
      RECT  8102.5 36540.0 8167.5 36725.0 ;
      RECT  8102.5 35380.0 8167.5 35565.0 ;
      RECT  7742.5 35497.5 7807.5 35347.5 ;
      RECT  7742.5 36382.5 7807.5 36757.5 ;
      RECT  7932.5 35497.5 7997.5 36382.5 ;
      RECT  7742.5 36382.5 7807.5 36517.5 ;
      RECT  7932.5 36382.5 7997.5 36517.5 ;
      RECT  7932.5 36382.5 7997.5 36517.5 ;
      RECT  7742.5 36382.5 7807.5 36517.5 ;
      RECT  7742.5 35497.5 7807.5 35632.5 ;
      RECT  7932.5 35497.5 7997.5 35632.5 ;
      RECT  7932.5 35497.5 7997.5 35632.5 ;
      RECT  7742.5 35497.5 7807.5 35632.5 ;
      RECT  8102.5 36472.5 8167.5 36607.5 ;
      RECT  8102.5 35497.5 8167.5 35632.5 ;
      RECT  7800.0 35940.0 7865.0 36075.0 ;
      RECT  7800.0 35940.0 7865.0 36075.0 ;
      RECT  7965.0 35975.0 8030.0 36040.0 ;
      RECT  7675.0 36692.5 8235.0 36757.5 ;
      RECT  7675.0 35347.5 8235.0 35412.5 ;
      RECT  8102.5 36910.0 8167.5 36725.0 ;
      RECT  8102.5 38070.0 8167.5 37885.0 ;
      RECT  7742.5 37952.5 7807.5 38102.5 ;
      RECT  7742.5 37067.5 7807.5 36692.5 ;
      RECT  7932.5 37952.5 7997.5 37067.5 ;
      RECT  7742.5 37067.5 7807.5 36932.5 ;
      RECT  7932.5 37067.5 7997.5 36932.5 ;
      RECT  7932.5 37067.5 7997.5 36932.5 ;
      RECT  7742.5 37067.5 7807.5 36932.5 ;
      RECT  7742.5 37952.5 7807.5 37817.5 ;
      RECT  7932.5 37952.5 7997.5 37817.5 ;
      RECT  7932.5 37952.5 7997.5 37817.5 ;
      RECT  7742.5 37952.5 7807.5 37817.5 ;
      RECT  8102.5 36977.5 8167.5 36842.5 ;
      RECT  8102.5 37952.5 8167.5 37817.5 ;
      RECT  7800.0 37510.0 7865.0 37375.0 ;
      RECT  7800.0 37510.0 7865.0 37375.0 ;
      RECT  7965.0 37475.0 8030.0 37410.0 ;
      RECT  7675.0 36757.5 8235.0 36692.5 ;
      RECT  7675.0 38102.5 8235.0 38037.5 ;
      RECT  8102.5 39230.0 8167.5 39415.0 ;
      RECT  8102.5 38070.0 8167.5 38255.0 ;
      RECT  7742.5 38187.5 7807.5 38037.5 ;
      RECT  7742.5 39072.5 7807.5 39447.5 ;
      RECT  7932.5 38187.5 7997.5 39072.5 ;
      RECT  7742.5 39072.5 7807.5 39207.5 ;
      RECT  7932.5 39072.5 7997.5 39207.5 ;
      RECT  7932.5 39072.5 7997.5 39207.5 ;
      RECT  7742.5 39072.5 7807.5 39207.5 ;
      RECT  7742.5 38187.5 7807.5 38322.5 ;
      RECT  7932.5 38187.5 7997.5 38322.5 ;
      RECT  7932.5 38187.5 7997.5 38322.5 ;
      RECT  7742.5 38187.5 7807.5 38322.5 ;
      RECT  8102.5 39162.5 8167.5 39297.5 ;
      RECT  8102.5 38187.5 8167.5 38322.5 ;
      RECT  7800.0 38630.0 7865.0 38765.0 ;
      RECT  7800.0 38630.0 7865.0 38765.0 ;
      RECT  7965.0 38665.0 8030.0 38730.0 ;
      RECT  7675.0 39382.5 8235.0 39447.5 ;
      RECT  7675.0 38037.5 8235.0 38102.5 ;
      RECT  8102.5 39600.0 8167.5 39415.0 ;
      RECT  8102.5 40760.0 8167.5 40575.0 ;
      RECT  7742.5 40642.5 7807.5 40792.5 ;
      RECT  7742.5 39757.5 7807.5 39382.5 ;
      RECT  7932.5 40642.5 7997.5 39757.5 ;
      RECT  7742.5 39757.5 7807.5 39622.5 ;
      RECT  7932.5 39757.5 7997.5 39622.5 ;
      RECT  7932.5 39757.5 7997.5 39622.5 ;
      RECT  7742.5 39757.5 7807.5 39622.5 ;
      RECT  7742.5 40642.5 7807.5 40507.5 ;
      RECT  7932.5 40642.5 7997.5 40507.5 ;
      RECT  7932.5 40642.5 7997.5 40507.5 ;
      RECT  7742.5 40642.5 7807.5 40507.5 ;
      RECT  8102.5 39667.5 8167.5 39532.5 ;
      RECT  8102.5 40642.5 8167.5 40507.5 ;
      RECT  7800.0 40200.0 7865.0 40065.0 ;
      RECT  7800.0 40200.0 7865.0 40065.0 ;
      RECT  7965.0 40165.0 8030.0 40100.0 ;
      RECT  7675.0 39447.5 8235.0 39382.5 ;
      RECT  7675.0 40792.5 8235.0 40727.5 ;
      RECT  8102.5 41920.0 8167.5 42105.0 ;
      RECT  8102.5 40760.0 8167.5 40945.0 ;
      RECT  7742.5 40877.5 7807.5 40727.5 ;
      RECT  7742.5 41762.5 7807.5 42137.5 ;
      RECT  7932.5 40877.5 7997.5 41762.5 ;
      RECT  7742.5 41762.5 7807.5 41897.5 ;
      RECT  7932.5 41762.5 7997.5 41897.5 ;
      RECT  7932.5 41762.5 7997.5 41897.5 ;
      RECT  7742.5 41762.5 7807.5 41897.5 ;
      RECT  7742.5 40877.5 7807.5 41012.5 ;
      RECT  7932.5 40877.5 7997.5 41012.5 ;
      RECT  7932.5 40877.5 7997.5 41012.5 ;
      RECT  7742.5 40877.5 7807.5 41012.5 ;
      RECT  8102.5 41852.5 8167.5 41987.5 ;
      RECT  8102.5 40877.5 8167.5 41012.5 ;
      RECT  7800.0 41320.0 7865.0 41455.0 ;
      RECT  7800.0 41320.0 7865.0 41455.0 ;
      RECT  7965.0 41355.0 8030.0 41420.0 ;
      RECT  7675.0 42072.5 8235.0 42137.5 ;
      RECT  7675.0 40727.5 8235.0 40792.5 ;
      RECT  8102.5 42290.0 8167.5 42105.0 ;
      RECT  8102.5 43450.0 8167.5 43265.0 ;
      RECT  7742.5 43332.5 7807.5 43482.5 ;
      RECT  7742.5 42447.5 7807.5 42072.5 ;
      RECT  7932.5 43332.5 7997.5 42447.5 ;
      RECT  7742.5 42447.5 7807.5 42312.5 ;
      RECT  7932.5 42447.5 7997.5 42312.5 ;
      RECT  7932.5 42447.5 7997.5 42312.5 ;
      RECT  7742.5 42447.5 7807.5 42312.5 ;
      RECT  7742.5 43332.5 7807.5 43197.5 ;
      RECT  7932.5 43332.5 7997.5 43197.5 ;
      RECT  7932.5 43332.5 7997.5 43197.5 ;
      RECT  7742.5 43332.5 7807.5 43197.5 ;
      RECT  8102.5 42357.5 8167.5 42222.5 ;
      RECT  8102.5 43332.5 8167.5 43197.5 ;
      RECT  7800.0 42890.0 7865.0 42755.0 ;
      RECT  7800.0 42890.0 7865.0 42755.0 ;
      RECT  7965.0 42855.0 8030.0 42790.0 ;
      RECT  7675.0 42137.5 8235.0 42072.5 ;
      RECT  7675.0 43482.5 8235.0 43417.5 ;
      RECT  8102.5 44610.0 8167.5 44795.0 ;
      RECT  8102.5 43450.0 8167.5 43635.0 ;
      RECT  7742.5 43567.5 7807.5 43417.5 ;
      RECT  7742.5 44452.5 7807.5 44827.5 ;
      RECT  7932.5 43567.5 7997.5 44452.5 ;
      RECT  7742.5 44452.5 7807.5 44587.5 ;
      RECT  7932.5 44452.5 7997.5 44587.5 ;
      RECT  7932.5 44452.5 7997.5 44587.5 ;
      RECT  7742.5 44452.5 7807.5 44587.5 ;
      RECT  7742.5 43567.5 7807.5 43702.5 ;
      RECT  7932.5 43567.5 7997.5 43702.5 ;
      RECT  7932.5 43567.5 7997.5 43702.5 ;
      RECT  7742.5 43567.5 7807.5 43702.5 ;
      RECT  8102.5 44542.5 8167.5 44677.5 ;
      RECT  8102.5 43567.5 8167.5 43702.5 ;
      RECT  7800.0 44010.0 7865.0 44145.0 ;
      RECT  7800.0 44010.0 7865.0 44145.0 ;
      RECT  7965.0 44045.0 8030.0 44110.0 ;
      RECT  7675.0 44762.5 8235.0 44827.5 ;
      RECT  7675.0 43417.5 8235.0 43482.5 ;
      RECT  8102.5 44980.0 8167.5 44795.0 ;
      RECT  8102.5 46140.0 8167.5 45955.0 ;
      RECT  7742.5 46022.5 7807.5 46172.5 ;
      RECT  7742.5 45137.5 7807.5 44762.5 ;
      RECT  7932.5 46022.5 7997.5 45137.5 ;
      RECT  7742.5 45137.5 7807.5 45002.5 ;
      RECT  7932.5 45137.5 7997.5 45002.5 ;
      RECT  7932.5 45137.5 7997.5 45002.5 ;
      RECT  7742.5 45137.5 7807.5 45002.5 ;
      RECT  7742.5 46022.5 7807.5 45887.5 ;
      RECT  7932.5 46022.5 7997.5 45887.5 ;
      RECT  7932.5 46022.5 7997.5 45887.5 ;
      RECT  7742.5 46022.5 7807.5 45887.5 ;
      RECT  8102.5 45047.5 8167.5 44912.5 ;
      RECT  8102.5 46022.5 8167.5 45887.5 ;
      RECT  7800.0 45580.0 7865.0 45445.0 ;
      RECT  7800.0 45580.0 7865.0 45445.0 ;
      RECT  7965.0 45545.0 8030.0 45480.0 ;
      RECT  7675.0 44827.5 8235.0 44762.5 ;
      RECT  7675.0 46172.5 8235.0 46107.5 ;
      RECT  8102.5 47300.0 8167.5 47485.0 ;
      RECT  8102.5 46140.0 8167.5 46325.0 ;
      RECT  7742.5 46257.5 7807.5 46107.5 ;
      RECT  7742.5 47142.5 7807.5 47517.5 ;
      RECT  7932.5 46257.5 7997.5 47142.5 ;
      RECT  7742.5 47142.5 7807.5 47277.5 ;
      RECT  7932.5 47142.5 7997.5 47277.5 ;
      RECT  7932.5 47142.5 7997.5 47277.5 ;
      RECT  7742.5 47142.5 7807.5 47277.5 ;
      RECT  7742.5 46257.5 7807.5 46392.5 ;
      RECT  7932.5 46257.5 7997.5 46392.5 ;
      RECT  7932.5 46257.5 7997.5 46392.5 ;
      RECT  7742.5 46257.5 7807.5 46392.5 ;
      RECT  8102.5 47232.5 8167.5 47367.5 ;
      RECT  8102.5 46257.5 8167.5 46392.5 ;
      RECT  7800.0 46700.0 7865.0 46835.0 ;
      RECT  7800.0 46700.0 7865.0 46835.0 ;
      RECT  7965.0 46735.0 8030.0 46800.0 ;
      RECT  7675.0 47452.5 8235.0 47517.5 ;
      RECT  7675.0 46107.5 8235.0 46172.5 ;
      RECT  8102.5 47670.0 8167.5 47485.0 ;
      RECT  8102.5 48830.0 8167.5 48645.0 ;
      RECT  7742.5 48712.5 7807.5 48862.5 ;
      RECT  7742.5 47827.5 7807.5 47452.5 ;
      RECT  7932.5 48712.5 7997.5 47827.5 ;
      RECT  7742.5 47827.5 7807.5 47692.5 ;
      RECT  7932.5 47827.5 7997.5 47692.5 ;
      RECT  7932.5 47827.5 7997.5 47692.5 ;
      RECT  7742.5 47827.5 7807.5 47692.5 ;
      RECT  7742.5 48712.5 7807.5 48577.5 ;
      RECT  7932.5 48712.5 7997.5 48577.5 ;
      RECT  7932.5 48712.5 7997.5 48577.5 ;
      RECT  7742.5 48712.5 7807.5 48577.5 ;
      RECT  8102.5 47737.5 8167.5 47602.5 ;
      RECT  8102.5 48712.5 8167.5 48577.5 ;
      RECT  7800.0 48270.0 7865.0 48135.0 ;
      RECT  7800.0 48270.0 7865.0 48135.0 ;
      RECT  7965.0 48235.0 8030.0 48170.0 ;
      RECT  7675.0 47517.5 8235.0 47452.5 ;
      RECT  7675.0 48862.5 8235.0 48797.5 ;
      RECT  8102.5 49990.0 8167.5 50175.0 ;
      RECT  8102.5 48830.0 8167.5 49015.0 ;
      RECT  7742.5 48947.5 7807.5 48797.5 ;
      RECT  7742.5 49832.5 7807.5 50207.5 ;
      RECT  7932.5 48947.5 7997.5 49832.5 ;
      RECT  7742.5 49832.5 7807.5 49967.5 ;
      RECT  7932.5 49832.5 7997.5 49967.5 ;
      RECT  7932.5 49832.5 7997.5 49967.5 ;
      RECT  7742.5 49832.5 7807.5 49967.5 ;
      RECT  7742.5 48947.5 7807.5 49082.5 ;
      RECT  7932.5 48947.5 7997.5 49082.5 ;
      RECT  7932.5 48947.5 7997.5 49082.5 ;
      RECT  7742.5 48947.5 7807.5 49082.5 ;
      RECT  8102.5 49922.5 8167.5 50057.5 ;
      RECT  8102.5 48947.5 8167.5 49082.5 ;
      RECT  7800.0 49390.0 7865.0 49525.0 ;
      RECT  7800.0 49390.0 7865.0 49525.0 ;
      RECT  7965.0 49425.0 8030.0 49490.0 ;
      RECT  7675.0 50142.5 8235.0 50207.5 ;
      RECT  7675.0 48797.5 8235.0 48862.5 ;
      RECT  8102.5 50360.0 8167.5 50175.0 ;
      RECT  8102.5 51520.0 8167.5 51335.0 ;
      RECT  7742.5 51402.5 7807.5 51552.5 ;
      RECT  7742.5 50517.5 7807.5 50142.5 ;
      RECT  7932.5 51402.5 7997.5 50517.5 ;
      RECT  7742.5 50517.5 7807.5 50382.5 ;
      RECT  7932.5 50517.5 7997.5 50382.5 ;
      RECT  7932.5 50517.5 7997.5 50382.5 ;
      RECT  7742.5 50517.5 7807.5 50382.5 ;
      RECT  7742.5 51402.5 7807.5 51267.5 ;
      RECT  7932.5 51402.5 7997.5 51267.5 ;
      RECT  7932.5 51402.5 7997.5 51267.5 ;
      RECT  7742.5 51402.5 7807.5 51267.5 ;
      RECT  8102.5 50427.5 8167.5 50292.5 ;
      RECT  8102.5 51402.5 8167.5 51267.5 ;
      RECT  7800.0 50960.0 7865.0 50825.0 ;
      RECT  7800.0 50960.0 7865.0 50825.0 ;
      RECT  7965.0 50925.0 8030.0 50860.0 ;
      RECT  7675.0 50207.5 8235.0 50142.5 ;
      RECT  7675.0 51552.5 8235.0 51487.5 ;
      RECT  8102.5 52680.0 8167.5 52865.0 ;
      RECT  8102.5 51520.0 8167.5 51705.0 ;
      RECT  7742.5 51637.5 7807.5 51487.5 ;
      RECT  7742.5 52522.5 7807.5 52897.5 ;
      RECT  7932.5 51637.5 7997.5 52522.5 ;
      RECT  7742.5 52522.5 7807.5 52657.5 ;
      RECT  7932.5 52522.5 7997.5 52657.5 ;
      RECT  7932.5 52522.5 7997.5 52657.5 ;
      RECT  7742.5 52522.5 7807.5 52657.5 ;
      RECT  7742.5 51637.5 7807.5 51772.5 ;
      RECT  7932.5 51637.5 7997.5 51772.5 ;
      RECT  7932.5 51637.5 7997.5 51772.5 ;
      RECT  7742.5 51637.5 7807.5 51772.5 ;
      RECT  8102.5 52612.5 8167.5 52747.5 ;
      RECT  8102.5 51637.5 8167.5 51772.5 ;
      RECT  7800.0 52080.0 7865.0 52215.0 ;
      RECT  7800.0 52080.0 7865.0 52215.0 ;
      RECT  7965.0 52115.0 8030.0 52180.0 ;
      RECT  7675.0 52832.5 8235.0 52897.5 ;
      RECT  7675.0 51487.5 8235.0 51552.5 ;
      RECT  8102.5 53050.0 8167.5 52865.0 ;
      RECT  8102.5 54210.0 8167.5 54025.0 ;
      RECT  7742.5 54092.5 7807.5 54242.5 ;
      RECT  7742.5 53207.5 7807.5 52832.5 ;
      RECT  7932.5 54092.5 7997.5 53207.5 ;
      RECT  7742.5 53207.5 7807.5 53072.5 ;
      RECT  7932.5 53207.5 7997.5 53072.5 ;
      RECT  7932.5 53207.5 7997.5 53072.5 ;
      RECT  7742.5 53207.5 7807.5 53072.5 ;
      RECT  7742.5 54092.5 7807.5 53957.5 ;
      RECT  7932.5 54092.5 7997.5 53957.5 ;
      RECT  7932.5 54092.5 7997.5 53957.5 ;
      RECT  7742.5 54092.5 7807.5 53957.5 ;
      RECT  8102.5 53117.5 8167.5 52982.5 ;
      RECT  8102.5 54092.5 8167.5 53957.5 ;
      RECT  7800.0 53650.0 7865.0 53515.0 ;
      RECT  7800.0 53650.0 7865.0 53515.0 ;
      RECT  7965.0 53615.0 8030.0 53550.0 ;
      RECT  7675.0 52897.5 8235.0 52832.5 ;
      RECT  7675.0 54242.5 8235.0 54177.5 ;
      RECT  8102.5 55370.0 8167.5 55555.0 ;
      RECT  8102.5 54210.0 8167.5 54395.0 ;
      RECT  7742.5 54327.5 7807.5 54177.5 ;
      RECT  7742.5 55212.5 7807.5 55587.5 ;
      RECT  7932.5 54327.5 7997.5 55212.5 ;
      RECT  7742.5 55212.5 7807.5 55347.5 ;
      RECT  7932.5 55212.5 7997.5 55347.5 ;
      RECT  7932.5 55212.5 7997.5 55347.5 ;
      RECT  7742.5 55212.5 7807.5 55347.5 ;
      RECT  7742.5 54327.5 7807.5 54462.5 ;
      RECT  7932.5 54327.5 7997.5 54462.5 ;
      RECT  7932.5 54327.5 7997.5 54462.5 ;
      RECT  7742.5 54327.5 7807.5 54462.5 ;
      RECT  8102.5 55302.5 8167.5 55437.5 ;
      RECT  8102.5 54327.5 8167.5 54462.5 ;
      RECT  7800.0 54770.0 7865.0 54905.0 ;
      RECT  7800.0 54770.0 7865.0 54905.0 ;
      RECT  7965.0 54805.0 8030.0 54870.0 ;
      RECT  7675.0 55522.5 8235.0 55587.5 ;
      RECT  7675.0 54177.5 8235.0 54242.5 ;
      RECT  8102.5 55740.0 8167.5 55555.0 ;
      RECT  8102.5 56900.0 8167.5 56715.0 ;
      RECT  7742.5 56782.5 7807.5 56932.5 ;
      RECT  7742.5 55897.5 7807.5 55522.5 ;
      RECT  7932.5 56782.5 7997.5 55897.5 ;
      RECT  7742.5 55897.5 7807.5 55762.5 ;
      RECT  7932.5 55897.5 7997.5 55762.5 ;
      RECT  7932.5 55897.5 7997.5 55762.5 ;
      RECT  7742.5 55897.5 7807.5 55762.5 ;
      RECT  7742.5 56782.5 7807.5 56647.5 ;
      RECT  7932.5 56782.5 7997.5 56647.5 ;
      RECT  7932.5 56782.5 7997.5 56647.5 ;
      RECT  7742.5 56782.5 7807.5 56647.5 ;
      RECT  8102.5 55807.5 8167.5 55672.5 ;
      RECT  8102.5 56782.5 8167.5 56647.5 ;
      RECT  7800.0 56340.0 7865.0 56205.0 ;
      RECT  7800.0 56340.0 7865.0 56205.0 ;
      RECT  7965.0 56305.0 8030.0 56240.0 ;
      RECT  7675.0 55587.5 8235.0 55522.5 ;
      RECT  7675.0 56932.5 8235.0 56867.5 ;
      RECT  8102.5 58060.0 8167.5 58245.0 ;
      RECT  8102.5 56900.0 8167.5 57085.0 ;
      RECT  7742.5 57017.5 7807.5 56867.5 ;
      RECT  7742.5 57902.5 7807.5 58277.5 ;
      RECT  7932.5 57017.5 7997.5 57902.5 ;
      RECT  7742.5 57902.5 7807.5 58037.5 ;
      RECT  7932.5 57902.5 7997.5 58037.5 ;
      RECT  7932.5 57902.5 7997.5 58037.5 ;
      RECT  7742.5 57902.5 7807.5 58037.5 ;
      RECT  7742.5 57017.5 7807.5 57152.5 ;
      RECT  7932.5 57017.5 7997.5 57152.5 ;
      RECT  7932.5 57017.5 7997.5 57152.5 ;
      RECT  7742.5 57017.5 7807.5 57152.5 ;
      RECT  8102.5 57992.5 8167.5 58127.5 ;
      RECT  8102.5 57017.5 8167.5 57152.5 ;
      RECT  7800.0 57460.0 7865.0 57595.0 ;
      RECT  7800.0 57460.0 7865.0 57595.0 ;
      RECT  7965.0 57495.0 8030.0 57560.0 ;
      RECT  7675.0 58212.5 8235.0 58277.5 ;
      RECT  7675.0 56867.5 8235.0 56932.5 ;
      RECT  8102.5 58430.0 8167.5 58245.0 ;
      RECT  8102.5 59590.0 8167.5 59405.0 ;
      RECT  7742.5 59472.5 7807.5 59622.5 ;
      RECT  7742.5 58587.5 7807.5 58212.5 ;
      RECT  7932.5 59472.5 7997.5 58587.5 ;
      RECT  7742.5 58587.5 7807.5 58452.5 ;
      RECT  7932.5 58587.5 7997.5 58452.5 ;
      RECT  7932.5 58587.5 7997.5 58452.5 ;
      RECT  7742.5 58587.5 7807.5 58452.5 ;
      RECT  7742.5 59472.5 7807.5 59337.5 ;
      RECT  7932.5 59472.5 7997.5 59337.5 ;
      RECT  7932.5 59472.5 7997.5 59337.5 ;
      RECT  7742.5 59472.5 7807.5 59337.5 ;
      RECT  8102.5 58497.5 8167.5 58362.5 ;
      RECT  8102.5 59472.5 8167.5 59337.5 ;
      RECT  7800.0 59030.0 7865.0 58895.0 ;
      RECT  7800.0 59030.0 7865.0 58895.0 ;
      RECT  7965.0 58995.0 8030.0 58930.0 ;
      RECT  7675.0 58277.5 8235.0 58212.5 ;
      RECT  7675.0 59622.5 8235.0 59557.5 ;
      RECT  8102.5 60750.0 8167.5 60935.0 ;
      RECT  8102.5 59590.0 8167.5 59775.0 ;
      RECT  7742.5 59707.5 7807.5 59557.5 ;
      RECT  7742.5 60592.5 7807.5 60967.5 ;
      RECT  7932.5 59707.5 7997.5 60592.5 ;
      RECT  7742.5 60592.5 7807.5 60727.5 ;
      RECT  7932.5 60592.5 7997.5 60727.5 ;
      RECT  7932.5 60592.5 7997.5 60727.5 ;
      RECT  7742.5 60592.5 7807.5 60727.5 ;
      RECT  7742.5 59707.5 7807.5 59842.5 ;
      RECT  7932.5 59707.5 7997.5 59842.5 ;
      RECT  7932.5 59707.5 7997.5 59842.5 ;
      RECT  7742.5 59707.5 7807.5 59842.5 ;
      RECT  8102.5 60682.5 8167.5 60817.5 ;
      RECT  8102.5 59707.5 8167.5 59842.5 ;
      RECT  7800.0 60150.0 7865.0 60285.0 ;
      RECT  7800.0 60150.0 7865.0 60285.0 ;
      RECT  7965.0 60185.0 8030.0 60250.0 ;
      RECT  7675.0 60902.5 8235.0 60967.5 ;
      RECT  7675.0 59557.5 8235.0 59622.5 ;
      RECT  8102.5 61120.0 8167.5 60935.0 ;
      RECT  8102.5 62280.0 8167.5 62095.0 ;
      RECT  7742.5 62162.5 7807.5 62312.5 ;
      RECT  7742.5 61277.5 7807.5 60902.5 ;
      RECT  7932.5 62162.5 7997.5 61277.5 ;
      RECT  7742.5 61277.5 7807.5 61142.5 ;
      RECT  7932.5 61277.5 7997.5 61142.5 ;
      RECT  7932.5 61277.5 7997.5 61142.5 ;
      RECT  7742.5 61277.5 7807.5 61142.5 ;
      RECT  7742.5 62162.5 7807.5 62027.5 ;
      RECT  7932.5 62162.5 7997.5 62027.5 ;
      RECT  7932.5 62162.5 7997.5 62027.5 ;
      RECT  7742.5 62162.5 7807.5 62027.5 ;
      RECT  8102.5 61187.5 8167.5 61052.5 ;
      RECT  8102.5 62162.5 8167.5 62027.5 ;
      RECT  7800.0 61720.0 7865.0 61585.0 ;
      RECT  7800.0 61720.0 7865.0 61585.0 ;
      RECT  7965.0 61685.0 8030.0 61620.0 ;
      RECT  7675.0 60967.5 8235.0 60902.5 ;
      RECT  7675.0 62312.5 8235.0 62247.5 ;
      RECT  8102.5 63440.0 8167.5 63625.0 ;
      RECT  8102.5 62280.0 8167.5 62465.0 ;
      RECT  7742.5 62397.5 7807.5 62247.5 ;
      RECT  7742.5 63282.5 7807.5 63657.5 ;
      RECT  7932.5 62397.5 7997.5 63282.5 ;
      RECT  7742.5 63282.5 7807.5 63417.5 ;
      RECT  7932.5 63282.5 7997.5 63417.5 ;
      RECT  7932.5 63282.5 7997.5 63417.5 ;
      RECT  7742.5 63282.5 7807.5 63417.5 ;
      RECT  7742.5 62397.5 7807.5 62532.5 ;
      RECT  7932.5 62397.5 7997.5 62532.5 ;
      RECT  7932.5 62397.5 7997.5 62532.5 ;
      RECT  7742.5 62397.5 7807.5 62532.5 ;
      RECT  8102.5 63372.5 8167.5 63507.5 ;
      RECT  8102.5 62397.5 8167.5 62532.5 ;
      RECT  7800.0 62840.0 7865.0 62975.0 ;
      RECT  7800.0 62840.0 7865.0 62975.0 ;
      RECT  7965.0 62875.0 8030.0 62940.0 ;
      RECT  7675.0 63592.5 8235.0 63657.5 ;
      RECT  7675.0 62247.5 8235.0 62312.5 ;
      RECT  8102.5 63810.0 8167.5 63625.0 ;
      RECT  8102.5 64970.0 8167.5 64785.0 ;
      RECT  7742.5 64852.5 7807.5 65002.5 ;
      RECT  7742.5 63967.5 7807.5 63592.5 ;
      RECT  7932.5 64852.5 7997.5 63967.5 ;
      RECT  7742.5 63967.5 7807.5 63832.5 ;
      RECT  7932.5 63967.5 7997.5 63832.5 ;
      RECT  7932.5 63967.5 7997.5 63832.5 ;
      RECT  7742.5 63967.5 7807.5 63832.5 ;
      RECT  7742.5 64852.5 7807.5 64717.5 ;
      RECT  7932.5 64852.5 7997.5 64717.5 ;
      RECT  7932.5 64852.5 7997.5 64717.5 ;
      RECT  7742.5 64852.5 7807.5 64717.5 ;
      RECT  8102.5 63877.5 8167.5 63742.5 ;
      RECT  8102.5 64852.5 8167.5 64717.5 ;
      RECT  7800.0 64410.0 7865.0 64275.0 ;
      RECT  7800.0 64410.0 7865.0 64275.0 ;
      RECT  7965.0 64375.0 8030.0 64310.0 ;
      RECT  7675.0 63657.5 8235.0 63592.5 ;
      RECT  7675.0 65002.5 8235.0 64937.5 ;
      RECT  8102.5 66130.0 8167.5 66315.0 ;
      RECT  8102.5 64970.0 8167.5 65155.0 ;
      RECT  7742.5 65087.5 7807.5 64937.5 ;
      RECT  7742.5 65972.5 7807.5 66347.5 ;
      RECT  7932.5 65087.5 7997.5 65972.5 ;
      RECT  7742.5 65972.5 7807.5 66107.5 ;
      RECT  7932.5 65972.5 7997.5 66107.5 ;
      RECT  7932.5 65972.5 7997.5 66107.5 ;
      RECT  7742.5 65972.5 7807.5 66107.5 ;
      RECT  7742.5 65087.5 7807.5 65222.5 ;
      RECT  7932.5 65087.5 7997.5 65222.5 ;
      RECT  7932.5 65087.5 7997.5 65222.5 ;
      RECT  7742.5 65087.5 7807.5 65222.5 ;
      RECT  8102.5 66062.5 8167.5 66197.5 ;
      RECT  8102.5 65087.5 8167.5 65222.5 ;
      RECT  7800.0 65530.0 7865.0 65665.0 ;
      RECT  7800.0 65530.0 7865.0 65665.0 ;
      RECT  7965.0 65565.0 8030.0 65630.0 ;
      RECT  7675.0 66282.5 8235.0 66347.5 ;
      RECT  7675.0 64937.5 8235.0 65002.5 ;
      RECT  8102.5 66500.0 8167.5 66315.0 ;
      RECT  8102.5 67660.0 8167.5 67475.0 ;
      RECT  7742.5 67542.5 7807.5 67692.5 ;
      RECT  7742.5 66657.5 7807.5 66282.5 ;
      RECT  7932.5 67542.5 7997.5 66657.5 ;
      RECT  7742.5 66657.5 7807.5 66522.5 ;
      RECT  7932.5 66657.5 7997.5 66522.5 ;
      RECT  7932.5 66657.5 7997.5 66522.5 ;
      RECT  7742.5 66657.5 7807.5 66522.5 ;
      RECT  7742.5 67542.5 7807.5 67407.5 ;
      RECT  7932.5 67542.5 7997.5 67407.5 ;
      RECT  7932.5 67542.5 7997.5 67407.5 ;
      RECT  7742.5 67542.5 7807.5 67407.5 ;
      RECT  8102.5 66567.5 8167.5 66432.5 ;
      RECT  8102.5 67542.5 8167.5 67407.5 ;
      RECT  7800.0 67100.0 7865.0 66965.0 ;
      RECT  7800.0 67100.0 7865.0 66965.0 ;
      RECT  7965.0 67065.0 8030.0 67000.0 ;
      RECT  7675.0 66347.5 8235.0 66282.5 ;
      RECT  7675.0 67692.5 8235.0 67627.5 ;
      RECT  8102.5 68820.0 8167.5 69005.0 ;
      RECT  8102.5 67660.0 8167.5 67845.0 ;
      RECT  7742.5 67777.5 7807.5 67627.5 ;
      RECT  7742.5 68662.5 7807.5 69037.5 ;
      RECT  7932.5 67777.5 7997.5 68662.5 ;
      RECT  7742.5 68662.5 7807.5 68797.5 ;
      RECT  7932.5 68662.5 7997.5 68797.5 ;
      RECT  7932.5 68662.5 7997.5 68797.5 ;
      RECT  7742.5 68662.5 7807.5 68797.5 ;
      RECT  7742.5 67777.5 7807.5 67912.5 ;
      RECT  7932.5 67777.5 7997.5 67912.5 ;
      RECT  7932.5 67777.5 7997.5 67912.5 ;
      RECT  7742.5 67777.5 7807.5 67912.5 ;
      RECT  8102.5 68752.5 8167.5 68887.5 ;
      RECT  8102.5 67777.5 8167.5 67912.5 ;
      RECT  7800.0 68220.0 7865.0 68355.0 ;
      RECT  7800.0 68220.0 7865.0 68355.0 ;
      RECT  7965.0 68255.0 8030.0 68320.0 ;
      RECT  7675.0 68972.5 8235.0 69037.5 ;
      RECT  7675.0 67627.5 8235.0 67692.5 ;
      RECT  8102.5 69190.0 8167.5 69005.0 ;
      RECT  8102.5 70350.0 8167.5 70165.0 ;
      RECT  7742.5 70232.5 7807.5 70382.5 ;
      RECT  7742.5 69347.5 7807.5 68972.5 ;
      RECT  7932.5 70232.5 7997.5 69347.5 ;
      RECT  7742.5 69347.5 7807.5 69212.5 ;
      RECT  7932.5 69347.5 7997.5 69212.5 ;
      RECT  7932.5 69347.5 7997.5 69212.5 ;
      RECT  7742.5 69347.5 7807.5 69212.5 ;
      RECT  7742.5 70232.5 7807.5 70097.5 ;
      RECT  7932.5 70232.5 7997.5 70097.5 ;
      RECT  7932.5 70232.5 7997.5 70097.5 ;
      RECT  7742.5 70232.5 7807.5 70097.5 ;
      RECT  8102.5 69257.5 8167.5 69122.5 ;
      RECT  8102.5 70232.5 8167.5 70097.5 ;
      RECT  7800.0 69790.0 7865.0 69655.0 ;
      RECT  7800.0 69790.0 7865.0 69655.0 ;
      RECT  7965.0 69755.0 8030.0 69690.0 ;
      RECT  7675.0 69037.5 8235.0 68972.5 ;
      RECT  7675.0 70382.5 8235.0 70317.5 ;
      RECT  4757.5 11765.0 4622.5 11830.0 ;
      RECT  4932.5 13200.0 4797.5 13265.0 ;
      RECT  5107.5 14455.0 4972.5 14520.0 ;
      RECT  5282.5 15890.0 5147.5 15955.0 ;
      RECT  5457.5 17145.0 5322.5 17210.0 ;
      RECT  5632.5 18580.0 5497.5 18645.0 ;
      RECT  5807.5 19835.0 5672.5 19900.0 ;
      RECT  5982.5 21270.0 5847.5 21335.0 ;
      RECT  6157.5 22525.0 6022.5 22590.0 ;
      RECT  6332.5 23960.0 6197.5 24025.0 ;
      RECT  6507.5 25215.0 6372.5 25280.0 ;
      RECT  6682.5 26650.0 6547.5 26715.0 ;
      RECT  4757.5 27917.5 4622.5 27982.5 ;
      RECT  5457.5 27702.5 5322.5 27767.5 ;
      RECT  4757.5 29327.5 4622.5 29392.5 ;
      RECT  5632.5 29542.5 5497.5 29607.5 ;
      RECT  4757.5 30607.5 4622.5 30672.5 ;
      RECT  5807.5 30392.5 5672.5 30457.5 ;
      RECT  4757.5 32017.5 4622.5 32082.5 ;
      RECT  5982.5 32232.5 5847.5 32297.5 ;
      RECT  4757.5 33297.5 4622.5 33362.5 ;
      RECT  6157.5 33082.5 6022.5 33147.5 ;
      RECT  4757.5 34707.5 4622.5 34772.5 ;
      RECT  6332.5 34922.5 6197.5 34987.5 ;
      RECT  4757.5 35987.5 4622.5 36052.5 ;
      RECT  6507.5 35772.5 6372.5 35837.5 ;
      RECT  4757.5 37397.5 4622.5 37462.5 ;
      RECT  6682.5 37612.5 6547.5 37677.5 ;
      RECT  4932.5 38677.5 4797.5 38742.5 ;
      RECT  5457.5 38462.5 5322.5 38527.5 ;
      RECT  4932.5 40087.5 4797.5 40152.5 ;
      RECT  5632.5 40302.5 5497.5 40367.5 ;
      RECT  4932.5 41367.5 4797.5 41432.5 ;
      RECT  5807.5 41152.5 5672.5 41217.5 ;
      RECT  4932.5 42777.5 4797.5 42842.5 ;
      RECT  5982.5 42992.5 5847.5 43057.5 ;
      RECT  4932.5 44057.5 4797.5 44122.5 ;
      RECT  6157.5 43842.5 6022.5 43907.5 ;
      RECT  4932.5 45467.5 4797.5 45532.5 ;
      RECT  6332.5 45682.5 6197.5 45747.5 ;
      RECT  4932.5 46747.5 4797.5 46812.5 ;
      RECT  6507.5 46532.5 6372.5 46597.5 ;
      RECT  4932.5 48157.5 4797.5 48222.5 ;
      RECT  6682.5 48372.5 6547.5 48437.5 ;
      RECT  5107.5 49437.5 4972.5 49502.5 ;
      RECT  5457.5 49222.5 5322.5 49287.5 ;
      RECT  5107.5 50847.5 4972.5 50912.5 ;
      RECT  5632.5 51062.5 5497.5 51127.5 ;
      RECT  5107.5 52127.5 4972.5 52192.5 ;
      RECT  5807.5 51912.5 5672.5 51977.5 ;
      RECT  5107.5 53537.5 4972.5 53602.5 ;
      RECT  5982.5 53752.5 5847.5 53817.5 ;
      RECT  5107.5 54817.5 4972.5 54882.5 ;
      RECT  6157.5 54602.5 6022.5 54667.5 ;
      RECT  5107.5 56227.5 4972.5 56292.5 ;
      RECT  6332.5 56442.5 6197.5 56507.5 ;
      RECT  5107.5 57507.5 4972.5 57572.5 ;
      RECT  6507.5 57292.5 6372.5 57357.5 ;
      RECT  5107.5 58917.5 4972.5 58982.5 ;
      RECT  6682.5 59132.5 6547.5 59197.5 ;
      RECT  5282.5 60197.5 5147.5 60262.5 ;
      RECT  5457.5 59982.5 5322.5 60047.5 ;
      RECT  5282.5 61607.5 5147.5 61672.5 ;
      RECT  5632.5 61822.5 5497.5 61887.5 ;
      RECT  5282.5 62887.5 5147.5 62952.5 ;
      RECT  5807.5 62672.5 5672.5 62737.5 ;
      RECT  5282.5 64297.5 5147.5 64362.5 ;
      RECT  5982.5 64512.5 5847.5 64577.5 ;
      RECT  5282.5 65577.5 5147.5 65642.5 ;
      RECT  6157.5 65362.5 6022.5 65427.5 ;
      RECT  5282.5 66987.5 5147.5 67052.5 ;
      RECT  6332.5 67202.5 6197.5 67267.5 ;
      RECT  5282.5 68267.5 5147.5 68332.5 ;
      RECT  6507.5 68052.5 6372.5 68117.5 ;
      RECT  5282.5 69677.5 5147.5 69742.5 ;
      RECT  6682.5 69892.5 6547.5 69957.5 ;
      RECT  7965.0 27905.0 8030.0 27970.0 ;
      RECT  7965.0 29340.0 8030.0 29405.0 ;
      RECT  7965.0 30595.0 8030.0 30660.0 ;
      RECT  7965.0 32030.0 8030.0 32095.0 ;
      RECT  7965.0 33285.0 8030.0 33350.0 ;
      RECT  7965.0 34720.0 8030.0 34785.0 ;
      RECT  7965.0 35975.0 8030.0 36040.0 ;
      RECT  7965.0 37410.0 8030.0 37475.0 ;
      RECT  7965.0 38665.0 8030.0 38730.0 ;
      RECT  7965.0 40100.0 8030.0 40165.0 ;
      RECT  7965.0 41355.0 8030.0 41420.0 ;
      RECT  7965.0 42790.0 8030.0 42855.0 ;
      RECT  7965.0 44045.0 8030.0 44110.0 ;
      RECT  7965.0 45480.0 8030.0 45545.0 ;
      RECT  7965.0 46735.0 8030.0 46800.0 ;
      RECT  7965.0 48170.0 8030.0 48235.0 ;
      RECT  7965.0 49425.0 8030.0 49490.0 ;
      RECT  7965.0 50860.0 8030.0 50925.0 ;
      RECT  7965.0 52115.0 8030.0 52180.0 ;
      RECT  7965.0 53550.0 8030.0 53615.0 ;
      RECT  7965.0 54805.0 8030.0 54870.0 ;
      RECT  7965.0 56240.0 8030.0 56305.0 ;
      RECT  7965.0 57495.0 8030.0 57560.0 ;
      RECT  7965.0 58930.0 8030.0 58995.0 ;
      RECT  7965.0 60185.0 8030.0 60250.0 ;
      RECT  7965.0 61620.0 8030.0 61685.0 ;
      RECT  7965.0 62875.0 8030.0 62940.0 ;
      RECT  7965.0 64310.0 8030.0 64375.0 ;
      RECT  7965.0 65565.0 8030.0 65630.0 ;
      RECT  7965.0 67000.0 8030.0 67065.0 ;
      RECT  7965.0 68255.0 8030.0 68320.0 ;
      RECT  7965.0 69690.0 8030.0 69755.0 ;
      RECT  4655.0 12482.5 11635.0 12547.5 ;
      RECT  4655.0 15172.5 11635.0 15237.5 ;
      RECT  4655.0 17862.5 11635.0 17927.5 ;
      RECT  4655.0 20552.5 11635.0 20617.5 ;
      RECT  4655.0 23242.5 11635.0 23307.5 ;
      RECT  4655.0 25932.5 11635.0 25997.5 ;
      RECT  4655.0 28622.5 11635.0 28687.5 ;
      RECT  4655.0 31312.5 11635.0 31377.5 ;
      RECT  4655.0 34002.5 11635.0 34067.5 ;
      RECT  4655.0 36692.5 11635.0 36757.5 ;
      RECT  4655.0 39382.5 11635.0 39447.5 ;
      RECT  4655.0 42072.5 11635.0 42137.5 ;
      RECT  4655.0 44762.5 11635.0 44827.5 ;
      RECT  4655.0 47452.5 11635.0 47517.5 ;
      RECT  4655.0 50142.5 11635.0 50207.5 ;
      RECT  4655.0 52832.5 11635.0 52897.5 ;
      RECT  4655.0 55522.5 11635.0 55587.5 ;
      RECT  4655.0 58212.5 11635.0 58277.5 ;
      RECT  4655.0 60902.5 11635.0 60967.5 ;
      RECT  4655.0 63592.5 11635.0 63657.5 ;
      RECT  4655.0 66282.5 11635.0 66347.5 ;
      RECT  4655.0 68972.5 11635.0 69037.5 ;
      RECT  4655.0 11137.5 11635.0 11202.5 ;
      RECT  4655.0 13827.5 11635.0 13892.5 ;
      RECT  4655.0 16517.5 11635.0 16582.5 ;
      RECT  4655.0 19207.5 11635.0 19272.5 ;
      RECT  4655.0 21897.5 11635.0 21962.5 ;
      RECT  4655.0 24587.5 11635.0 24652.5 ;
      RECT  4655.0 27277.5 11635.0 27342.5 ;
      RECT  4655.0 29967.5 11635.0 30032.5 ;
      RECT  4655.0 32657.5 11635.0 32722.5 ;
      RECT  4655.0 35347.5 11635.0 35412.5 ;
      RECT  4655.0 38037.5 11635.0 38102.5 ;
      RECT  4655.0 40727.5 11635.0 40792.5 ;
      RECT  4655.0 43417.5 11635.0 43482.5 ;
      RECT  4655.0 46107.5 11635.0 46172.5 ;
      RECT  4655.0 48797.5 11635.0 48862.5 ;
      RECT  4655.0 51487.5 11635.0 51552.5 ;
      RECT  4655.0 54177.5 11635.0 54242.5 ;
      RECT  4655.0 56867.5 11635.0 56932.5 ;
      RECT  4655.0 59557.5 11635.0 59622.5 ;
      RECT  4655.0 62247.5 11635.0 62312.5 ;
      RECT  4655.0 64937.5 11635.0 65002.5 ;
      RECT  4655.0 67627.5 11635.0 67692.5 ;
      RECT  4655.0 70317.5 11635.0 70382.5 ;
      RECT  8465.0 27905.0 8815.0 27970.0 ;
      RECT  8980.0 27917.5 9045.0 27982.5 ;
      RECT  8980.0 27905.0 9045.0 27970.0 ;
      RECT  8980.0 27950.0 9045.0 27970.0 ;
      RECT  9012.5 27917.5 9310.0 27982.5 ;
      RECT  9310.0 27917.5 9445.0 27982.5 ;
      RECT  10015.0 27917.5 10080.0 27982.5 ;
      RECT  10015.0 27905.0 10080.0 27970.0 ;
      RECT  9797.5 27917.5 10047.5 27982.5 ;
      RECT  10015.0 27937.5 10080.0 27950.0 ;
      RECT  10047.5 27905.0 10295.0 27970.0 ;
      RECT  8465.0 29340.0 8815.0 29405.0 ;
      RECT  8980.0 29327.5 9045.0 29392.5 ;
      RECT  8980.0 29340.0 9045.0 29405.0 ;
      RECT  8980.0 29360.0 9045.0 29405.0 ;
      RECT  9012.5 29327.5 9310.0 29392.5 ;
      RECT  9310.0 29327.5 9445.0 29392.5 ;
      RECT  10015.0 29327.5 10080.0 29392.5 ;
      RECT  10015.0 29340.0 10080.0 29405.0 ;
      RECT  9797.5 29327.5 10047.5 29392.5 ;
      RECT  10015.0 29360.0 10080.0 29372.5 ;
      RECT  10047.5 29340.0 10295.0 29405.0 ;
      RECT  8465.0 30595.0 8815.0 30660.0 ;
      RECT  8980.0 30607.5 9045.0 30672.5 ;
      RECT  8980.0 30595.0 9045.0 30660.0 ;
      RECT  8980.0 30640.0 9045.0 30660.0 ;
      RECT  9012.5 30607.5 9310.0 30672.5 ;
      RECT  9310.0 30607.5 9445.0 30672.5 ;
      RECT  10015.0 30607.5 10080.0 30672.5 ;
      RECT  10015.0 30595.0 10080.0 30660.0 ;
      RECT  9797.5 30607.5 10047.5 30672.5 ;
      RECT  10015.0 30627.5 10080.0 30640.0 ;
      RECT  10047.5 30595.0 10295.0 30660.0 ;
      RECT  8465.0 32030.0 8815.0 32095.0 ;
      RECT  8980.0 32017.5 9045.0 32082.5 ;
      RECT  8980.0 32030.0 9045.0 32095.0 ;
      RECT  8980.0 32050.0 9045.0 32095.0 ;
      RECT  9012.5 32017.5 9310.0 32082.5 ;
      RECT  9310.0 32017.5 9445.0 32082.5 ;
      RECT  10015.0 32017.5 10080.0 32082.5 ;
      RECT  10015.0 32030.0 10080.0 32095.0 ;
      RECT  9797.5 32017.5 10047.5 32082.5 ;
      RECT  10015.0 32050.0 10080.0 32062.5 ;
      RECT  10047.5 32030.0 10295.0 32095.0 ;
      RECT  8465.0 33285.0 8815.0 33350.0 ;
      RECT  8980.0 33297.5 9045.0 33362.5 ;
      RECT  8980.0 33285.0 9045.0 33350.0 ;
      RECT  8980.0 33330.0 9045.0 33350.0 ;
      RECT  9012.5 33297.5 9310.0 33362.5 ;
      RECT  9310.0 33297.5 9445.0 33362.5 ;
      RECT  10015.0 33297.5 10080.0 33362.5 ;
      RECT  10015.0 33285.0 10080.0 33350.0 ;
      RECT  9797.5 33297.5 10047.5 33362.5 ;
      RECT  10015.0 33317.5 10080.0 33330.0 ;
      RECT  10047.5 33285.0 10295.0 33350.0 ;
      RECT  8465.0 34720.0 8815.0 34785.0 ;
      RECT  8980.0 34707.5 9045.0 34772.5 ;
      RECT  8980.0 34720.0 9045.0 34785.0 ;
      RECT  8980.0 34740.0 9045.0 34785.0 ;
      RECT  9012.5 34707.5 9310.0 34772.5 ;
      RECT  9310.0 34707.5 9445.0 34772.5 ;
      RECT  10015.0 34707.5 10080.0 34772.5 ;
      RECT  10015.0 34720.0 10080.0 34785.0 ;
      RECT  9797.5 34707.5 10047.5 34772.5 ;
      RECT  10015.0 34740.0 10080.0 34752.5 ;
      RECT  10047.5 34720.0 10295.0 34785.0 ;
      RECT  8465.0 35975.0 8815.0 36040.0 ;
      RECT  8980.0 35987.5 9045.0 36052.5 ;
      RECT  8980.0 35975.0 9045.0 36040.0 ;
      RECT  8980.0 36020.0 9045.0 36040.0 ;
      RECT  9012.5 35987.5 9310.0 36052.5 ;
      RECT  9310.0 35987.5 9445.0 36052.5 ;
      RECT  10015.0 35987.5 10080.0 36052.5 ;
      RECT  10015.0 35975.0 10080.0 36040.0 ;
      RECT  9797.5 35987.5 10047.5 36052.5 ;
      RECT  10015.0 36007.5 10080.0 36020.0 ;
      RECT  10047.5 35975.0 10295.0 36040.0 ;
      RECT  8465.0 37410.0 8815.0 37475.0 ;
      RECT  8980.0 37397.5 9045.0 37462.5 ;
      RECT  8980.0 37410.0 9045.0 37475.0 ;
      RECT  8980.0 37430.0 9045.0 37475.0 ;
      RECT  9012.5 37397.5 9310.0 37462.5 ;
      RECT  9310.0 37397.5 9445.0 37462.5 ;
      RECT  10015.0 37397.5 10080.0 37462.5 ;
      RECT  10015.0 37410.0 10080.0 37475.0 ;
      RECT  9797.5 37397.5 10047.5 37462.5 ;
      RECT  10015.0 37430.0 10080.0 37442.5 ;
      RECT  10047.5 37410.0 10295.0 37475.0 ;
      RECT  8465.0 38665.0 8815.0 38730.0 ;
      RECT  8980.0 38677.5 9045.0 38742.5 ;
      RECT  8980.0 38665.0 9045.0 38730.0 ;
      RECT  8980.0 38710.0 9045.0 38730.0 ;
      RECT  9012.5 38677.5 9310.0 38742.5 ;
      RECT  9310.0 38677.5 9445.0 38742.5 ;
      RECT  10015.0 38677.5 10080.0 38742.5 ;
      RECT  10015.0 38665.0 10080.0 38730.0 ;
      RECT  9797.5 38677.5 10047.5 38742.5 ;
      RECT  10015.0 38697.5 10080.0 38710.0 ;
      RECT  10047.5 38665.0 10295.0 38730.0 ;
      RECT  8465.0 40100.0 8815.0 40165.0 ;
      RECT  8980.0 40087.5 9045.0 40152.5 ;
      RECT  8980.0 40100.0 9045.0 40165.0 ;
      RECT  8980.0 40120.0 9045.0 40165.0 ;
      RECT  9012.5 40087.5 9310.0 40152.5 ;
      RECT  9310.0 40087.5 9445.0 40152.5 ;
      RECT  10015.0 40087.5 10080.0 40152.5 ;
      RECT  10015.0 40100.0 10080.0 40165.0 ;
      RECT  9797.5 40087.5 10047.5 40152.5 ;
      RECT  10015.0 40120.0 10080.0 40132.5 ;
      RECT  10047.5 40100.0 10295.0 40165.0 ;
      RECT  8465.0 41355.0 8815.0 41420.0 ;
      RECT  8980.0 41367.5 9045.0 41432.5 ;
      RECT  8980.0 41355.0 9045.0 41420.0 ;
      RECT  8980.0 41400.0 9045.0 41420.0 ;
      RECT  9012.5 41367.5 9310.0 41432.5 ;
      RECT  9310.0 41367.5 9445.0 41432.5 ;
      RECT  10015.0 41367.5 10080.0 41432.5 ;
      RECT  10015.0 41355.0 10080.0 41420.0 ;
      RECT  9797.5 41367.5 10047.5 41432.5 ;
      RECT  10015.0 41387.5 10080.0 41400.0 ;
      RECT  10047.5 41355.0 10295.0 41420.0 ;
      RECT  8465.0 42790.0 8815.0 42855.0 ;
      RECT  8980.0 42777.5 9045.0 42842.5 ;
      RECT  8980.0 42790.0 9045.0 42855.0 ;
      RECT  8980.0 42810.0 9045.0 42855.0 ;
      RECT  9012.5 42777.5 9310.0 42842.5 ;
      RECT  9310.0 42777.5 9445.0 42842.5 ;
      RECT  10015.0 42777.5 10080.0 42842.5 ;
      RECT  10015.0 42790.0 10080.0 42855.0 ;
      RECT  9797.5 42777.5 10047.5 42842.5 ;
      RECT  10015.0 42810.0 10080.0 42822.5 ;
      RECT  10047.5 42790.0 10295.0 42855.0 ;
      RECT  8465.0 44045.0 8815.0 44110.0 ;
      RECT  8980.0 44057.5 9045.0 44122.5 ;
      RECT  8980.0 44045.0 9045.0 44110.0 ;
      RECT  8980.0 44090.0 9045.0 44110.0 ;
      RECT  9012.5 44057.5 9310.0 44122.5 ;
      RECT  9310.0 44057.5 9445.0 44122.5 ;
      RECT  10015.0 44057.5 10080.0 44122.5 ;
      RECT  10015.0 44045.0 10080.0 44110.0 ;
      RECT  9797.5 44057.5 10047.5 44122.5 ;
      RECT  10015.0 44077.5 10080.0 44090.0 ;
      RECT  10047.5 44045.0 10295.0 44110.0 ;
      RECT  8465.0 45480.0 8815.0 45545.0 ;
      RECT  8980.0 45467.5 9045.0 45532.5 ;
      RECT  8980.0 45480.0 9045.0 45545.0 ;
      RECT  8980.0 45500.0 9045.0 45545.0 ;
      RECT  9012.5 45467.5 9310.0 45532.5 ;
      RECT  9310.0 45467.5 9445.0 45532.5 ;
      RECT  10015.0 45467.5 10080.0 45532.5 ;
      RECT  10015.0 45480.0 10080.0 45545.0 ;
      RECT  9797.5 45467.5 10047.5 45532.5 ;
      RECT  10015.0 45500.0 10080.0 45512.5 ;
      RECT  10047.5 45480.0 10295.0 45545.0 ;
      RECT  8465.0 46735.0 8815.0 46800.0 ;
      RECT  8980.0 46747.5 9045.0 46812.5 ;
      RECT  8980.0 46735.0 9045.0 46800.0 ;
      RECT  8980.0 46780.0 9045.0 46800.0 ;
      RECT  9012.5 46747.5 9310.0 46812.5 ;
      RECT  9310.0 46747.5 9445.0 46812.5 ;
      RECT  10015.0 46747.5 10080.0 46812.5 ;
      RECT  10015.0 46735.0 10080.0 46800.0 ;
      RECT  9797.5 46747.5 10047.5 46812.5 ;
      RECT  10015.0 46767.5 10080.0 46780.0 ;
      RECT  10047.5 46735.0 10295.0 46800.0 ;
      RECT  8465.0 48170.0 8815.0 48235.0 ;
      RECT  8980.0 48157.5 9045.0 48222.5 ;
      RECT  8980.0 48170.0 9045.0 48235.0 ;
      RECT  8980.0 48190.0 9045.0 48235.0 ;
      RECT  9012.5 48157.5 9310.0 48222.5 ;
      RECT  9310.0 48157.5 9445.0 48222.5 ;
      RECT  10015.0 48157.5 10080.0 48222.5 ;
      RECT  10015.0 48170.0 10080.0 48235.0 ;
      RECT  9797.5 48157.5 10047.5 48222.5 ;
      RECT  10015.0 48190.0 10080.0 48202.5 ;
      RECT  10047.5 48170.0 10295.0 48235.0 ;
      RECT  8465.0 49425.0 8815.0 49490.0 ;
      RECT  8980.0 49437.5 9045.0 49502.5 ;
      RECT  8980.0 49425.0 9045.0 49490.0 ;
      RECT  8980.0 49470.0 9045.0 49490.0 ;
      RECT  9012.5 49437.5 9310.0 49502.5 ;
      RECT  9310.0 49437.5 9445.0 49502.5 ;
      RECT  10015.0 49437.5 10080.0 49502.5 ;
      RECT  10015.0 49425.0 10080.0 49490.0 ;
      RECT  9797.5 49437.5 10047.5 49502.5 ;
      RECT  10015.0 49457.5 10080.0 49470.0 ;
      RECT  10047.5 49425.0 10295.0 49490.0 ;
      RECT  8465.0 50860.0 8815.0 50925.0 ;
      RECT  8980.0 50847.5 9045.0 50912.5 ;
      RECT  8980.0 50860.0 9045.0 50925.0 ;
      RECT  8980.0 50880.0 9045.0 50925.0 ;
      RECT  9012.5 50847.5 9310.0 50912.5 ;
      RECT  9310.0 50847.5 9445.0 50912.5 ;
      RECT  10015.0 50847.5 10080.0 50912.5 ;
      RECT  10015.0 50860.0 10080.0 50925.0 ;
      RECT  9797.5 50847.5 10047.5 50912.5 ;
      RECT  10015.0 50880.0 10080.0 50892.5 ;
      RECT  10047.5 50860.0 10295.0 50925.0 ;
      RECT  8465.0 52115.0 8815.0 52180.0 ;
      RECT  8980.0 52127.5 9045.0 52192.5 ;
      RECT  8980.0 52115.0 9045.0 52180.0 ;
      RECT  8980.0 52160.0 9045.0 52180.0 ;
      RECT  9012.5 52127.5 9310.0 52192.5 ;
      RECT  9310.0 52127.5 9445.0 52192.5 ;
      RECT  10015.0 52127.5 10080.0 52192.5 ;
      RECT  10015.0 52115.0 10080.0 52180.0 ;
      RECT  9797.5 52127.5 10047.5 52192.5 ;
      RECT  10015.0 52147.5 10080.0 52160.0 ;
      RECT  10047.5 52115.0 10295.0 52180.0 ;
      RECT  8465.0 53550.0 8815.0 53615.0 ;
      RECT  8980.0 53537.5 9045.0 53602.5 ;
      RECT  8980.0 53550.0 9045.0 53615.0 ;
      RECT  8980.0 53570.0 9045.0 53615.0 ;
      RECT  9012.5 53537.5 9310.0 53602.5 ;
      RECT  9310.0 53537.5 9445.0 53602.5 ;
      RECT  10015.0 53537.5 10080.0 53602.5 ;
      RECT  10015.0 53550.0 10080.0 53615.0 ;
      RECT  9797.5 53537.5 10047.5 53602.5 ;
      RECT  10015.0 53570.0 10080.0 53582.5 ;
      RECT  10047.5 53550.0 10295.0 53615.0 ;
      RECT  8465.0 54805.0 8815.0 54870.0 ;
      RECT  8980.0 54817.5 9045.0 54882.5 ;
      RECT  8980.0 54805.0 9045.0 54870.0 ;
      RECT  8980.0 54850.0 9045.0 54870.0 ;
      RECT  9012.5 54817.5 9310.0 54882.5 ;
      RECT  9310.0 54817.5 9445.0 54882.5 ;
      RECT  10015.0 54817.5 10080.0 54882.5 ;
      RECT  10015.0 54805.0 10080.0 54870.0 ;
      RECT  9797.5 54817.5 10047.5 54882.5 ;
      RECT  10015.0 54837.5 10080.0 54850.0 ;
      RECT  10047.5 54805.0 10295.0 54870.0 ;
      RECT  8465.0 56240.0 8815.0 56305.0 ;
      RECT  8980.0 56227.5 9045.0 56292.5 ;
      RECT  8980.0 56240.0 9045.0 56305.0 ;
      RECT  8980.0 56260.0 9045.0 56305.0 ;
      RECT  9012.5 56227.5 9310.0 56292.5 ;
      RECT  9310.0 56227.5 9445.0 56292.5 ;
      RECT  10015.0 56227.5 10080.0 56292.5 ;
      RECT  10015.0 56240.0 10080.0 56305.0 ;
      RECT  9797.5 56227.5 10047.5 56292.5 ;
      RECT  10015.0 56260.0 10080.0 56272.5 ;
      RECT  10047.5 56240.0 10295.0 56305.0 ;
      RECT  8465.0 57495.0 8815.0 57560.0 ;
      RECT  8980.0 57507.5 9045.0 57572.5 ;
      RECT  8980.0 57495.0 9045.0 57560.0 ;
      RECT  8980.0 57540.0 9045.0 57560.0 ;
      RECT  9012.5 57507.5 9310.0 57572.5 ;
      RECT  9310.0 57507.5 9445.0 57572.5 ;
      RECT  10015.0 57507.5 10080.0 57572.5 ;
      RECT  10015.0 57495.0 10080.0 57560.0 ;
      RECT  9797.5 57507.5 10047.5 57572.5 ;
      RECT  10015.0 57527.5 10080.0 57540.0 ;
      RECT  10047.5 57495.0 10295.0 57560.0 ;
      RECT  8465.0 58930.0 8815.0 58995.0 ;
      RECT  8980.0 58917.5 9045.0 58982.5 ;
      RECT  8980.0 58930.0 9045.0 58995.0 ;
      RECT  8980.0 58950.0 9045.0 58995.0 ;
      RECT  9012.5 58917.5 9310.0 58982.5 ;
      RECT  9310.0 58917.5 9445.0 58982.5 ;
      RECT  10015.0 58917.5 10080.0 58982.5 ;
      RECT  10015.0 58930.0 10080.0 58995.0 ;
      RECT  9797.5 58917.5 10047.5 58982.5 ;
      RECT  10015.0 58950.0 10080.0 58962.5 ;
      RECT  10047.5 58930.0 10295.0 58995.0 ;
      RECT  8465.0 60185.0 8815.0 60250.0 ;
      RECT  8980.0 60197.5 9045.0 60262.5 ;
      RECT  8980.0 60185.0 9045.0 60250.0 ;
      RECT  8980.0 60230.0 9045.0 60250.0 ;
      RECT  9012.5 60197.5 9310.0 60262.5 ;
      RECT  9310.0 60197.5 9445.0 60262.5 ;
      RECT  10015.0 60197.5 10080.0 60262.5 ;
      RECT  10015.0 60185.0 10080.0 60250.0 ;
      RECT  9797.5 60197.5 10047.5 60262.5 ;
      RECT  10015.0 60217.5 10080.0 60230.0 ;
      RECT  10047.5 60185.0 10295.0 60250.0 ;
      RECT  8465.0 61620.0 8815.0 61685.0 ;
      RECT  8980.0 61607.5 9045.0 61672.5 ;
      RECT  8980.0 61620.0 9045.0 61685.0 ;
      RECT  8980.0 61640.0 9045.0 61685.0 ;
      RECT  9012.5 61607.5 9310.0 61672.5 ;
      RECT  9310.0 61607.5 9445.0 61672.5 ;
      RECT  10015.0 61607.5 10080.0 61672.5 ;
      RECT  10015.0 61620.0 10080.0 61685.0 ;
      RECT  9797.5 61607.5 10047.5 61672.5 ;
      RECT  10015.0 61640.0 10080.0 61652.5 ;
      RECT  10047.5 61620.0 10295.0 61685.0 ;
      RECT  8465.0 62875.0 8815.0 62940.0 ;
      RECT  8980.0 62887.5 9045.0 62952.5 ;
      RECT  8980.0 62875.0 9045.0 62940.0 ;
      RECT  8980.0 62920.0 9045.0 62940.0 ;
      RECT  9012.5 62887.5 9310.0 62952.5 ;
      RECT  9310.0 62887.5 9445.0 62952.5 ;
      RECT  10015.0 62887.5 10080.0 62952.5 ;
      RECT  10015.0 62875.0 10080.0 62940.0 ;
      RECT  9797.5 62887.5 10047.5 62952.5 ;
      RECT  10015.0 62907.5 10080.0 62920.0 ;
      RECT  10047.5 62875.0 10295.0 62940.0 ;
      RECT  8465.0 64310.0 8815.0 64375.0 ;
      RECT  8980.0 64297.5 9045.0 64362.5 ;
      RECT  8980.0 64310.0 9045.0 64375.0 ;
      RECT  8980.0 64330.0 9045.0 64375.0 ;
      RECT  9012.5 64297.5 9310.0 64362.5 ;
      RECT  9310.0 64297.5 9445.0 64362.5 ;
      RECT  10015.0 64297.5 10080.0 64362.5 ;
      RECT  10015.0 64310.0 10080.0 64375.0 ;
      RECT  9797.5 64297.5 10047.5 64362.5 ;
      RECT  10015.0 64330.0 10080.0 64342.5 ;
      RECT  10047.5 64310.0 10295.0 64375.0 ;
      RECT  8465.0 65565.0 8815.0 65630.0 ;
      RECT  8980.0 65577.5 9045.0 65642.5 ;
      RECT  8980.0 65565.0 9045.0 65630.0 ;
      RECT  8980.0 65610.0 9045.0 65630.0 ;
      RECT  9012.5 65577.5 9310.0 65642.5 ;
      RECT  9310.0 65577.5 9445.0 65642.5 ;
      RECT  10015.0 65577.5 10080.0 65642.5 ;
      RECT  10015.0 65565.0 10080.0 65630.0 ;
      RECT  9797.5 65577.5 10047.5 65642.5 ;
      RECT  10015.0 65597.5 10080.0 65610.0 ;
      RECT  10047.5 65565.0 10295.0 65630.0 ;
      RECT  8465.0 67000.0 8815.0 67065.0 ;
      RECT  8980.0 66987.5 9045.0 67052.5 ;
      RECT  8980.0 67000.0 9045.0 67065.0 ;
      RECT  8980.0 67020.0 9045.0 67065.0 ;
      RECT  9012.5 66987.5 9310.0 67052.5 ;
      RECT  9310.0 66987.5 9445.0 67052.5 ;
      RECT  10015.0 66987.5 10080.0 67052.5 ;
      RECT  10015.0 67000.0 10080.0 67065.0 ;
      RECT  9797.5 66987.5 10047.5 67052.5 ;
      RECT  10015.0 67020.0 10080.0 67032.5 ;
      RECT  10047.5 67000.0 10295.0 67065.0 ;
      RECT  8465.0 68255.0 8815.0 68320.0 ;
      RECT  8980.0 68267.5 9045.0 68332.5 ;
      RECT  8980.0 68255.0 9045.0 68320.0 ;
      RECT  8980.0 68300.0 9045.0 68320.0 ;
      RECT  9012.5 68267.5 9310.0 68332.5 ;
      RECT  9310.0 68267.5 9445.0 68332.5 ;
      RECT  10015.0 68267.5 10080.0 68332.5 ;
      RECT  10015.0 68255.0 10080.0 68320.0 ;
      RECT  9797.5 68267.5 10047.5 68332.5 ;
      RECT  10015.0 68287.5 10080.0 68300.0 ;
      RECT  10047.5 68255.0 10295.0 68320.0 ;
      RECT  8465.0 69690.0 8815.0 69755.0 ;
      RECT  8980.0 69677.5 9045.0 69742.5 ;
      RECT  8980.0 69690.0 9045.0 69755.0 ;
      RECT  8980.0 69710.0 9045.0 69755.0 ;
      RECT  9012.5 69677.5 9310.0 69742.5 ;
      RECT  9310.0 69677.5 9445.0 69742.5 ;
      RECT  10015.0 69677.5 10080.0 69742.5 ;
      RECT  10015.0 69690.0 10080.0 69755.0 ;
      RECT  9797.5 69677.5 10047.5 69742.5 ;
      RECT  10015.0 69710.0 10080.0 69722.5 ;
      RECT  10047.5 69690.0 10295.0 69755.0 ;
      RECT  9117.5 28470.0 9182.5 28655.0 ;
      RECT  9117.5 27310.0 9182.5 27495.0 ;
      RECT  8757.5 27427.5 8822.5 27277.5 ;
      RECT  8757.5 28312.5 8822.5 28687.5 ;
      RECT  8947.5 27427.5 9012.5 28312.5 ;
      RECT  8757.5 28312.5 8822.5 28447.5 ;
      RECT  8947.5 28312.5 9012.5 28447.5 ;
      RECT  8947.5 28312.5 9012.5 28447.5 ;
      RECT  8757.5 28312.5 8822.5 28447.5 ;
      RECT  8757.5 27427.5 8822.5 27562.5 ;
      RECT  8947.5 27427.5 9012.5 27562.5 ;
      RECT  8947.5 27427.5 9012.5 27562.5 ;
      RECT  8757.5 27427.5 8822.5 27562.5 ;
      RECT  9117.5 28402.5 9182.5 28537.5 ;
      RECT  9117.5 27427.5 9182.5 27562.5 ;
      RECT  8815.0 27870.0 8880.0 28005.0 ;
      RECT  8815.0 27870.0 8880.0 28005.0 ;
      RECT  8980.0 27905.0 9045.0 27970.0 ;
      RECT  8690.0 28622.5 9250.0 28687.5 ;
      RECT  8690.0 27277.5 9250.0 27342.5 ;
      RECT  9317.5 27472.5 9382.5 27277.5 ;
      RECT  9317.5 28312.5 9382.5 28687.5 ;
      RECT  9697.5 28312.5 9762.5 28687.5 ;
      RECT  9867.5 28470.0 9932.5 28655.0 ;
      RECT  9867.5 27310.0 9932.5 27495.0 ;
      RECT  9317.5 28312.5 9382.5 28447.5 ;
      RECT  9507.5 28312.5 9572.5 28447.5 ;
      RECT  9507.5 28312.5 9572.5 28447.5 ;
      RECT  9317.5 28312.5 9382.5 28447.5 ;
      RECT  9507.5 28312.5 9572.5 28447.5 ;
      RECT  9697.5 28312.5 9762.5 28447.5 ;
      RECT  9697.5 28312.5 9762.5 28447.5 ;
      RECT  9507.5 28312.5 9572.5 28447.5 ;
      RECT  9317.5 27472.5 9382.5 27607.5 ;
      RECT  9507.5 27472.5 9572.5 27607.5 ;
      RECT  9507.5 27472.5 9572.5 27607.5 ;
      RECT  9317.5 27472.5 9382.5 27607.5 ;
      RECT  9507.5 27472.5 9572.5 27607.5 ;
      RECT  9697.5 27472.5 9762.5 27607.5 ;
      RECT  9697.5 27472.5 9762.5 27607.5 ;
      RECT  9507.5 27472.5 9572.5 27607.5 ;
      RECT  9867.5 28402.5 9932.5 28537.5 ;
      RECT  9867.5 27427.5 9932.5 27562.5 ;
      RECT  9702.5 27702.5 9567.5 27767.5 ;
      RECT  9445.0 27917.5 9310.0 27982.5 ;
      RECT  9507.5 28312.5 9572.5 28447.5 ;
      RECT  9697.5 27472.5 9762.5 27607.5 ;
      RECT  9797.5 27917.5 9662.5 27982.5 ;
      RECT  9310.0 27917.5 9445.0 27982.5 ;
      RECT  9567.5 27702.5 9702.5 27767.5 ;
      RECT  9662.5 27917.5 9797.5 27982.5 ;
      RECT  9250.0 28622.5 10170.0 28687.5 ;
      RECT  9250.0 27277.5 10170.0 27342.5 ;
      RECT  10597.5 28470.0 10662.5 28655.0 ;
      RECT  10597.5 27310.0 10662.5 27495.0 ;
      RECT  10237.5 27427.5 10302.5 27277.5 ;
      RECT  10237.5 28312.5 10302.5 28687.5 ;
      RECT  10427.5 27427.5 10492.5 28312.5 ;
      RECT  10237.5 28312.5 10302.5 28447.5 ;
      RECT  10427.5 28312.5 10492.5 28447.5 ;
      RECT  10427.5 28312.5 10492.5 28447.5 ;
      RECT  10237.5 28312.5 10302.5 28447.5 ;
      RECT  10237.5 27427.5 10302.5 27562.5 ;
      RECT  10427.5 27427.5 10492.5 27562.5 ;
      RECT  10427.5 27427.5 10492.5 27562.5 ;
      RECT  10237.5 27427.5 10302.5 27562.5 ;
      RECT  10597.5 28402.5 10662.5 28537.5 ;
      RECT  10597.5 27427.5 10662.5 27562.5 ;
      RECT  10295.0 27870.0 10360.0 28005.0 ;
      RECT  10295.0 27870.0 10360.0 28005.0 ;
      RECT  10460.0 27905.0 10525.0 27970.0 ;
      RECT  10170.0 28622.5 10730.0 28687.5 ;
      RECT  10170.0 27277.5 10730.0 27342.5 ;
      RECT  8432.5 27870.0 8497.5 28005.0 ;
      RECT  8572.5 27597.5 8637.5 27732.5 ;
      RECT  9567.5 27702.5 9432.5 27767.5 ;
      RECT  9117.5 28840.0 9182.5 28655.0 ;
      RECT  9117.5 30000.0 9182.5 29815.0 ;
      RECT  8757.5 29882.5 8822.5 30032.5 ;
      RECT  8757.5 28997.5 8822.5 28622.5 ;
      RECT  8947.5 29882.5 9012.5 28997.5 ;
      RECT  8757.5 28997.5 8822.5 28862.5 ;
      RECT  8947.5 28997.5 9012.5 28862.5 ;
      RECT  8947.5 28997.5 9012.5 28862.5 ;
      RECT  8757.5 28997.5 8822.5 28862.5 ;
      RECT  8757.5 29882.5 8822.5 29747.5 ;
      RECT  8947.5 29882.5 9012.5 29747.5 ;
      RECT  8947.5 29882.5 9012.5 29747.5 ;
      RECT  8757.5 29882.5 8822.5 29747.5 ;
      RECT  9117.5 28907.5 9182.5 28772.5 ;
      RECT  9117.5 29882.5 9182.5 29747.5 ;
      RECT  8815.0 29440.0 8880.0 29305.0 ;
      RECT  8815.0 29440.0 8880.0 29305.0 ;
      RECT  8980.0 29405.0 9045.0 29340.0 ;
      RECT  8690.0 28687.5 9250.0 28622.5 ;
      RECT  8690.0 30032.5 9250.0 29967.5 ;
      RECT  9317.5 29837.5 9382.5 30032.5 ;
      RECT  9317.5 28997.5 9382.5 28622.5 ;
      RECT  9697.5 28997.5 9762.5 28622.5 ;
      RECT  9867.5 28840.0 9932.5 28655.0 ;
      RECT  9867.5 30000.0 9932.5 29815.0 ;
      RECT  9317.5 28997.5 9382.5 28862.5 ;
      RECT  9507.5 28997.5 9572.5 28862.5 ;
      RECT  9507.5 28997.5 9572.5 28862.5 ;
      RECT  9317.5 28997.5 9382.5 28862.5 ;
      RECT  9507.5 28997.5 9572.5 28862.5 ;
      RECT  9697.5 28997.5 9762.5 28862.5 ;
      RECT  9697.5 28997.5 9762.5 28862.5 ;
      RECT  9507.5 28997.5 9572.5 28862.5 ;
      RECT  9317.5 29837.5 9382.5 29702.5 ;
      RECT  9507.5 29837.5 9572.5 29702.5 ;
      RECT  9507.5 29837.5 9572.5 29702.5 ;
      RECT  9317.5 29837.5 9382.5 29702.5 ;
      RECT  9507.5 29837.5 9572.5 29702.5 ;
      RECT  9697.5 29837.5 9762.5 29702.5 ;
      RECT  9697.5 29837.5 9762.5 29702.5 ;
      RECT  9507.5 29837.5 9572.5 29702.5 ;
      RECT  9867.5 28907.5 9932.5 28772.5 ;
      RECT  9867.5 29882.5 9932.5 29747.5 ;
      RECT  9702.5 29607.5 9567.5 29542.5 ;
      RECT  9445.0 29392.5 9310.0 29327.5 ;
      RECT  9507.5 28997.5 9572.5 28862.5 ;
      RECT  9697.5 29837.5 9762.5 29702.5 ;
      RECT  9797.5 29392.5 9662.5 29327.5 ;
      RECT  9310.0 29392.5 9445.0 29327.5 ;
      RECT  9567.5 29607.5 9702.5 29542.5 ;
      RECT  9662.5 29392.5 9797.5 29327.5 ;
      RECT  9250.0 28687.5 10170.0 28622.5 ;
      RECT  9250.0 30032.5 10170.0 29967.5 ;
      RECT  10597.5 28840.0 10662.5 28655.0 ;
      RECT  10597.5 30000.0 10662.5 29815.0 ;
      RECT  10237.5 29882.5 10302.5 30032.5 ;
      RECT  10237.5 28997.5 10302.5 28622.5 ;
      RECT  10427.5 29882.5 10492.5 28997.5 ;
      RECT  10237.5 28997.5 10302.5 28862.5 ;
      RECT  10427.5 28997.5 10492.5 28862.5 ;
      RECT  10427.5 28997.5 10492.5 28862.5 ;
      RECT  10237.5 28997.5 10302.5 28862.5 ;
      RECT  10237.5 29882.5 10302.5 29747.5 ;
      RECT  10427.5 29882.5 10492.5 29747.5 ;
      RECT  10427.5 29882.5 10492.5 29747.5 ;
      RECT  10237.5 29882.5 10302.5 29747.5 ;
      RECT  10597.5 28907.5 10662.5 28772.5 ;
      RECT  10597.5 29882.5 10662.5 29747.5 ;
      RECT  10295.0 29440.0 10360.0 29305.0 ;
      RECT  10295.0 29440.0 10360.0 29305.0 ;
      RECT  10460.0 29405.0 10525.0 29340.0 ;
      RECT  10170.0 28687.5 10730.0 28622.5 ;
      RECT  10170.0 30032.5 10730.0 29967.5 ;
      RECT  8432.5 29305.0 8497.5 29440.0 ;
      RECT  8572.5 29577.5 8637.5 29712.5 ;
      RECT  9567.5 29542.5 9432.5 29607.5 ;
      RECT  9117.5 31160.0 9182.5 31345.0 ;
      RECT  9117.5 30000.0 9182.5 30185.0 ;
      RECT  8757.5 30117.5 8822.5 29967.5 ;
      RECT  8757.5 31002.5 8822.5 31377.5 ;
      RECT  8947.5 30117.5 9012.5 31002.5 ;
      RECT  8757.5 31002.5 8822.5 31137.5 ;
      RECT  8947.5 31002.5 9012.5 31137.5 ;
      RECT  8947.5 31002.5 9012.5 31137.5 ;
      RECT  8757.5 31002.5 8822.5 31137.5 ;
      RECT  8757.5 30117.5 8822.5 30252.5 ;
      RECT  8947.5 30117.5 9012.5 30252.5 ;
      RECT  8947.5 30117.5 9012.5 30252.5 ;
      RECT  8757.5 30117.5 8822.5 30252.5 ;
      RECT  9117.5 31092.5 9182.5 31227.5 ;
      RECT  9117.5 30117.5 9182.5 30252.5 ;
      RECT  8815.0 30560.0 8880.0 30695.0 ;
      RECT  8815.0 30560.0 8880.0 30695.0 ;
      RECT  8980.0 30595.0 9045.0 30660.0 ;
      RECT  8690.0 31312.5 9250.0 31377.5 ;
      RECT  8690.0 29967.5 9250.0 30032.5 ;
      RECT  9317.5 30162.5 9382.5 29967.5 ;
      RECT  9317.5 31002.5 9382.5 31377.5 ;
      RECT  9697.5 31002.5 9762.5 31377.5 ;
      RECT  9867.5 31160.0 9932.5 31345.0 ;
      RECT  9867.5 30000.0 9932.5 30185.0 ;
      RECT  9317.5 31002.5 9382.5 31137.5 ;
      RECT  9507.5 31002.5 9572.5 31137.5 ;
      RECT  9507.5 31002.5 9572.5 31137.5 ;
      RECT  9317.5 31002.5 9382.5 31137.5 ;
      RECT  9507.5 31002.5 9572.5 31137.5 ;
      RECT  9697.5 31002.5 9762.5 31137.5 ;
      RECT  9697.5 31002.5 9762.5 31137.5 ;
      RECT  9507.5 31002.5 9572.5 31137.5 ;
      RECT  9317.5 30162.5 9382.5 30297.5 ;
      RECT  9507.5 30162.5 9572.5 30297.5 ;
      RECT  9507.5 30162.5 9572.5 30297.5 ;
      RECT  9317.5 30162.5 9382.5 30297.5 ;
      RECT  9507.5 30162.5 9572.5 30297.5 ;
      RECT  9697.5 30162.5 9762.5 30297.5 ;
      RECT  9697.5 30162.5 9762.5 30297.5 ;
      RECT  9507.5 30162.5 9572.5 30297.5 ;
      RECT  9867.5 31092.5 9932.5 31227.5 ;
      RECT  9867.5 30117.5 9932.5 30252.5 ;
      RECT  9702.5 30392.5 9567.5 30457.5 ;
      RECT  9445.0 30607.5 9310.0 30672.5 ;
      RECT  9507.5 31002.5 9572.5 31137.5 ;
      RECT  9697.5 30162.5 9762.5 30297.5 ;
      RECT  9797.5 30607.5 9662.5 30672.5 ;
      RECT  9310.0 30607.5 9445.0 30672.5 ;
      RECT  9567.5 30392.5 9702.5 30457.5 ;
      RECT  9662.5 30607.5 9797.5 30672.5 ;
      RECT  9250.0 31312.5 10170.0 31377.5 ;
      RECT  9250.0 29967.5 10170.0 30032.5 ;
      RECT  10597.5 31160.0 10662.5 31345.0 ;
      RECT  10597.5 30000.0 10662.5 30185.0 ;
      RECT  10237.5 30117.5 10302.5 29967.5 ;
      RECT  10237.5 31002.5 10302.5 31377.5 ;
      RECT  10427.5 30117.5 10492.5 31002.5 ;
      RECT  10237.5 31002.5 10302.5 31137.5 ;
      RECT  10427.5 31002.5 10492.5 31137.5 ;
      RECT  10427.5 31002.5 10492.5 31137.5 ;
      RECT  10237.5 31002.5 10302.5 31137.5 ;
      RECT  10237.5 30117.5 10302.5 30252.5 ;
      RECT  10427.5 30117.5 10492.5 30252.5 ;
      RECT  10427.5 30117.5 10492.5 30252.5 ;
      RECT  10237.5 30117.5 10302.5 30252.5 ;
      RECT  10597.5 31092.5 10662.5 31227.5 ;
      RECT  10597.5 30117.5 10662.5 30252.5 ;
      RECT  10295.0 30560.0 10360.0 30695.0 ;
      RECT  10295.0 30560.0 10360.0 30695.0 ;
      RECT  10460.0 30595.0 10525.0 30660.0 ;
      RECT  10170.0 31312.5 10730.0 31377.5 ;
      RECT  10170.0 29967.5 10730.0 30032.5 ;
      RECT  8432.5 30560.0 8497.5 30695.0 ;
      RECT  8572.5 30287.5 8637.5 30422.5 ;
      RECT  9567.5 30392.5 9432.5 30457.5 ;
      RECT  9117.5 31530.0 9182.5 31345.0 ;
      RECT  9117.5 32690.0 9182.5 32505.0 ;
      RECT  8757.5 32572.5 8822.5 32722.5 ;
      RECT  8757.5 31687.5 8822.5 31312.5 ;
      RECT  8947.5 32572.5 9012.5 31687.5 ;
      RECT  8757.5 31687.5 8822.5 31552.5 ;
      RECT  8947.5 31687.5 9012.5 31552.5 ;
      RECT  8947.5 31687.5 9012.5 31552.5 ;
      RECT  8757.5 31687.5 8822.5 31552.5 ;
      RECT  8757.5 32572.5 8822.5 32437.5 ;
      RECT  8947.5 32572.5 9012.5 32437.5 ;
      RECT  8947.5 32572.5 9012.5 32437.5 ;
      RECT  8757.5 32572.5 8822.5 32437.5 ;
      RECT  9117.5 31597.5 9182.5 31462.5 ;
      RECT  9117.5 32572.5 9182.5 32437.5 ;
      RECT  8815.0 32130.0 8880.0 31995.0 ;
      RECT  8815.0 32130.0 8880.0 31995.0 ;
      RECT  8980.0 32095.0 9045.0 32030.0 ;
      RECT  8690.0 31377.5 9250.0 31312.5 ;
      RECT  8690.0 32722.5 9250.0 32657.5 ;
      RECT  9317.5 32527.5 9382.5 32722.5 ;
      RECT  9317.5 31687.5 9382.5 31312.5 ;
      RECT  9697.5 31687.5 9762.5 31312.5 ;
      RECT  9867.5 31530.0 9932.5 31345.0 ;
      RECT  9867.5 32690.0 9932.5 32505.0 ;
      RECT  9317.5 31687.5 9382.5 31552.5 ;
      RECT  9507.5 31687.5 9572.5 31552.5 ;
      RECT  9507.5 31687.5 9572.5 31552.5 ;
      RECT  9317.5 31687.5 9382.5 31552.5 ;
      RECT  9507.5 31687.5 9572.5 31552.5 ;
      RECT  9697.5 31687.5 9762.5 31552.5 ;
      RECT  9697.5 31687.5 9762.5 31552.5 ;
      RECT  9507.5 31687.5 9572.5 31552.5 ;
      RECT  9317.5 32527.5 9382.5 32392.5 ;
      RECT  9507.5 32527.5 9572.5 32392.5 ;
      RECT  9507.5 32527.5 9572.5 32392.5 ;
      RECT  9317.5 32527.5 9382.5 32392.5 ;
      RECT  9507.5 32527.5 9572.5 32392.5 ;
      RECT  9697.5 32527.5 9762.5 32392.5 ;
      RECT  9697.5 32527.5 9762.5 32392.5 ;
      RECT  9507.5 32527.5 9572.5 32392.5 ;
      RECT  9867.5 31597.5 9932.5 31462.5 ;
      RECT  9867.5 32572.5 9932.5 32437.5 ;
      RECT  9702.5 32297.5 9567.5 32232.5 ;
      RECT  9445.0 32082.5 9310.0 32017.5 ;
      RECT  9507.5 31687.5 9572.5 31552.5 ;
      RECT  9697.5 32527.5 9762.5 32392.5 ;
      RECT  9797.5 32082.5 9662.5 32017.5 ;
      RECT  9310.0 32082.5 9445.0 32017.5 ;
      RECT  9567.5 32297.5 9702.5 32232.5 ;
      RECT  9662.5 32082.5 9797.5 32017.5 ;
      RECT  9250.0 31377.5 10170.0 31312.5 ;
      RECT  9250.0 32722.5 10170.0 32657.5 ;
      RECT  10597.5 31530.0 10662.5 31345.0 ;
      RECT  10597.5 32690.0 10662.5 32505.0 ;
      RECT  10237.5 32572.5 10302.5 32722.5 ;
      RECT  10237.5 31687.5 10302.5 31312.5 ;
      RECT  10427.5 32572.5 10492.5 31687.5 ;
      RECT  10237.5 31687.5 10302.5 31552.5 ;
      RECT  10427.5 31687.5 10492.5 31552.5 ;
      RECT  10427.5 31687.5 10492.5 31552.5 ;
      RECT  10237.5 31687.5 10302.5 31552.5 ;
      RECT  10237.5 32572.5 10302.5 32437.5 ;
      RECT  10427.5 32572.5 10492.5 32437.5 ;
      RECT  10427.5 32572.5 10492.5 32437.5 ;
      RECT  10237.5 32572.5 10302.5 32437.5 ;
      RECT  10597.5 31597.5 10662.5 31462.5 ;
      RECT  10597.5 32572.5 10662.5 32437.5 ;
      RECT  10295.0 32130.0 10360.0 31995.0 ;
      RECT  10295.0 32130.0 10360.0 31995.0 ;
      RECT  10460.0 32095.0 10525.0 32030.0 ;
      RECT  10170.0 31377.5 10730.0 31312.5 ;
      RECT  10170.0 32722.5 10730.0 32657.5 ;
      RECT  8432.5 31995.0 8497.5 32130.0 ;
      RECT  8572.5 32267.5 8637.5 32402.5 ;
      RECT  9567.5 32232.5 9432.5 32297.5 ;
      RECT  9117.5 33850.0 9182.5 34035.0 ;
      RECT  9117.5 32690.0 9182.5 32875.0 ;
      RECT  8757.5 32807.5 8822.5 32657.5 ;
      RECT  8757.5 33692.5 8822.5 34067.5 ;
      RECT  8947.5 32807.5 9012.5 33692.5 ;
      RECT  8757.5 33692.5 8822.5 33827.5 ;
      RECT  8947.5 33692.5 9012.5 33827.5 ;
      RECT  8947.5 33692.5 9012.5 33827.5 ;
      RECT  8757.5 33692.5 8822.5 33827.5 ;
      RECT  8757.5 32807.5 8822.5 32942.5 ;
      RECT  8947.5 32807.5 9012.5 32942.5 ;
      RECT  8947.5 32807.5 9012.5 32942.5 ;
      RECT  8757.5 32807.5 8822.5 32942.5 ;
      RECT  9117.5 33782.5 9182.5 33917.5 ;
      RECT  9117.5 32807.5 9182.5 32942.5 ;
      RECT  8815.0 33250.0 8880.0 33385.0 ;
      RECT  8815.0 33250.0 8880.0 33385.0 ;
      RECT  8980.0 33285.0 9045.0 33350.0 ;
      RECT  8690.0 34002.5 9250.0 34067.5 ;
      RECT  8690.0 32657.5 9250.0 32722.5 ;
      RECT  9317.5 32852.5 9382.5 32657.5 ;
      RECT  9317.5 33692.5 9382.5 34067.5 ;
      RECT  9697.5 33692.5 9762.5 34067.5 ;
      RECT  9867.5 33850.0 9932.5 34035.0 ;
      RECT  9867.5 32690.0 9932.5 32875.0 ;
      RECT  9317.5 33692.5 9382.5 33827.5 ;
      RECT  9507.5 33692.5 9572.5 33827.5 ;
      RECT  9507.5 33692.5 9572.5 33827.5 ;
      RECT  9317.5 33692.5 9382.5 33827.5 ;
      RECT  9507.5 33692.5 9572.5 33827.5 ;
      RECT  9697.5 33692.5 9762.5 33827.5 ;
      RECT  9697.5 33692.5 9762.5 33827.5 ;
      RECT  9507.5 33692.5 9572.5 33827.5 ;
      RECT  9317.5 32852.5 9382.5 32987.5 ;
      RECT  9507.5 32852.5 9572.5 32987.5 ;
      RECT  9507.5 32852.5 9572.5 32987.5 ;
      RECT  9317.5 32852.5 9382.5 32987.5 ;
      RECT  9507.5 32852.5 9572.5 32987.5 ;
      RECT  9697.5 32852.5 9762.5 32987.5 ;
      RECT  9697.5 32852.5 9762.5 32987.5 ;
      RECT  9507.5 32852.5 9572.5 32987.5 ;
      RECT  9867.5 33782.5 9932.5 33917.5 ;
      RECT  9867.5 32807.5 9932.5 32942.5 ;
      RECT  9702.5 33082.5 9567.5 33147.5 ;
      RECT  9445.0 33297.5 9310.0 33362.5 ;
      RECT  9507.5 33692.5 9572.5 33827.5 ;
      RECT  9697.5 32852.5 9762.5 32987.5 ;
      RECT  9797.5 33297.5 9662.5 33362.5 ;
      RECT  9310.0 33297.5 9445.0 33362.5 ;
      RECT  9567.5 33082.5 9702.5 33147.5 ;
      RECT  9662.5 33297.5 9797.5 33362.5 ;
      RECT  9250.0 34002.5 10170.0 34067.5 ;
      RECT  9250.0 32657.5 10170.0 32722.5 ;
      RECT  10597.5 33850.0 10662.5 34035.0 ;
      RECT  10597.5 32690.0 10662.5 32875.0 ;
      RECT  10237.5 32807.5 10302.5 32657.5 ;
      RECT  10237.5 33692.5 10302.5 34067.5 ;
      RECT  10427.5 32807.5 10492.5 33692.5 ;
      RECT  10237.5 33692.5 10302.5 33827.5 ;
      RECT  10427.5 33692.5 10492.5 33827.5 ;
      RECT  10427.5 33692.5 10492.5 33827.5 ;
      RECT  10237.5 33692.5 10302.5 33827.5 ;
      RECT  10237.5 32807.5 10302.5 32942.5 ;
      RECT  10427.5 32807.5 10492.5 32942.5 ;
      RECT  10427.5 32807.5 10492.5 32942.5 ;
      RECT  10237.5 32807.5 10302.5 32942.5 ;
      RECT  10597.5 33782.5 10662.5 33917.5 ;
      RECT  10597.5 32807.5 10662.5 32942.5 ;
      RECT  10295.0 33250.0 10360.0 33385.0 ;
      RECT  10295.0 33250.0 10360.0 33385.0 ;
      RECT  10460.0 33285.0 10525.0 33350.0 ;
      RECT  10170.0 34002.5 10730.0 34067.5 ;
      RECT  10170.0 32657.5 10730.0 32722.5 ;
      RECT  8432.5 33250.0 8497.5 33385.0 ;
      RECT  8572.5 32977.5 8637.5 33112.5 ;
      RECT  9567.5 33082.5 9432.5 33147.5 ;
      RECT  9117.5 34220.0 9182.5 34035.0 ;
      RECT  9117.5 35380.0 9182.5 35195.0 ;
      RECT  8757.5 35262.5 8822.5 35412.5 ;
      RECT  8757.5 34377.5 8822.5 34002.5 ;
      RECT  8947.5 35262.5 9012.5 34377.5 ;
      RECT  8757.5 34377.5 8822.5 34242.5 ;
      RECT  8947.5 34377.5 9012.5 34242.5 ;
      RECT  8947.5 34377.5 9012.5 34242.5 ;
      RECT  8757.5 34377.5 8822.5 34242.5 ;
      RECT  8757.5 35262.5 8822.5 35127.5 ;
      RECT  8947.5 35262.5 9012.5 35127.5 ;
      RECT  8947.5 35262.5 9012.5 35127.5 ;
      RECT  8757.5 35262.5 8822.5 35127.5 ;
      RECT  9117.5 34287.5 9182.5 34152.5 ;
      RECT  9117.5 35262.5 9182.5 35127.5 ;
      RECT  8815.0 34820.0 8880.0 34685.0 ;
      RECT  8815.0 34820.0 8880.0 34685.0 ;
      RECT  8980.0 34785.0 9045.0 34720.0 ;
      RECT  8690.0 34067.5 9250.0 34002.5 ;
      RECT  8690.0 35412.5 9250.0 35347.5 ;
      RECT  9317.5 35217.5 9382.5 35412.5 ;
      RECT  9317.5 34377.5 9382.5 34002.5 ;
      RECT  9697.5 34377.5 9762.5 34002.5 ;
      RECT  9867.5 34220.0 9932.5 34035.0 ;
      RECT  9867.5 35380.0 9932.5 35195.0 ;
      RECT  9317.5 34377.5 9382.5 34242.5 ;
      RECT  9507.5 34377.5 9572.5 34242.5 ;
      RECT  9507.5 34377.5 9572.5 34242.5 ;
      RECT  9317.5 34377.5 9382.5 34242.5 ;
      RECT  9507.5 34377.5 9572.5 34242.5 ;
      RECT  9697.5 34377.5 9762.5 34242.5 ;
      RECT  9697.5 34377.5 9762.5 34242.5 ;
      RECT  9507.5 34377.5 9572.5 34242.5 ;
      RECT  9317.5 35217.5 9382.5 35082.5 ;
      RECT  9507.5 35217.5 9572.5 35082.5 ;
      RECT  9507.5 35217.5 9572.5 35082.5 ;
      RECT  9317.5 35217.5 9382.5 35082.5 ;
      RECT  9507.5 35217.5 9572.5 35082.5 ;
      RECT  9697.5 35217.5 9762.5 35082.5 ;
      RECT  9697.5 35217.5 9762.5 35082.5 ;
      RECT  9507.5 35217.5 9572.5 35082.5 ;
      RECT  9867.5 34287.5 9932.5 34152.5 ;
      RECT  9867.5 35262.5 9932.5 35127.5 ;
      RECT  9702.5 34987.5 9567.5 34922.5 ;
      RECT  9445.0 34772.5 9310.0 34707.5 ;
      RECT  9507.5 34377.5 9572.5 34242.5 ;
      RECT  9697.5 35217.5 9762.5 35082.5 ;
      RECT  9797.5 34772.5 9662.5 34707.5 ;
      RECT  9310.0 34772.5 9445.0 34707.5 ;
      RECT  9567.5 34987.5 9702.5 34922.5 ;
      RECT  9662.5 34772.5 9797.5 34707.5 ;
      RECT  9250.0 34067.5 10170.0 34002.5 ;
      RECT  9250.0 35412.5 10170.0 35347.5 ;
      RECT  10597.5 34220.0 10662.5 34035.0 ;
      RECT  10597.5 35380.0 10662.5 35195.0 ;
      RECT  10237.5 35262.5 10302.5 35412.5 ;
      RECT  10237.5 34377.5 10302.5 34002.5 ;
      RECT  10427.5 35262.5 10492.5 34377.5 ;
      RECT  10237.5 34377.5 10302.5 34242.5 ;
      RECT  10427.5 34377.5 10492.5 34242.5 ;
      RECT  10427.5 34377.5 10492.5 34242.5 ;
      RECT  10237.5 34377.5 10302.5 34242.5 ;
      RECT  10237.5 35262.5 10302.5 35127.5 ;
      RECT  10427.5 35262.5 10492.5 35127.5 ;
      RECT  10427.5 35262.5 10492.5 35127.5 ;
      RECT  10237.5 35262.5 10302.5 35127.5 ;
      RECT  10597.5 34287.5 10662.5 34152.5 ;
      RECT  10597.5 35262.5 10662.5 35127.5 ;
      RECT  10295.0 34820.0 10360.0 34685.0 ;
      RECT  10295.0 34820.0 10360.0 34685.0 ;
      RECT  10460.0 34785.0 10525.0 34720.0 ;
      RECT  10170.0 34067.5 10730.0 34002.5 ;
      RECT  10170.0 35412.5 10730.0 35347.5 ;
      RECT  8432.5 34685.0 8497.5 34820.0 ;
      RECT  8572.5 34957.5 8637.5 35092.5 ;
      RECT  9567.5 34922.5 9432.5 34987.5 ;
      RECT  9117.5 36540.0 9182.5 36725.0 ;
      RECT  9117.5 35380.0 9182.5 35565.0 ;
      RECT  8757.5 35497.5 8822.5 35347.5 ;
      RECT  8757.5 36382.5 8822.5 36757.5 ;
      RECT  8947.5 35497.5 9012.5 36382.5 ;
      RECT  8757.5 36382.5 8822.5 36517.5 ;
      RECT  8947.5 36382.5 9012.5 36517.5 ;
      RECT  8947.5 36382.5 9012.5 36517.5 ;
      RECT  8757.5 36382.5 8822.5 36517.5 ;
      RECT  8757.5 35497.5 8822.5 35632.5 ;
      RECT  8947.5 35497.5 9012.5 35632.5 ;
      RECT  8947.5 35497.5 9012.5 35632.5 ;
      RECT  8757.5 35497.5 8822.5 35632.5 ;
      RECT  9117.5 36472.5 9182.5 36607.5 ;
      RECT  9117.5 35497.5 9182.5 35632.5 ;
      RECT  8815.0 35940.0 8880.0 36075.0 ;
      RECT  8815.0 35940.0 8880.0 36075.0 ;
      RECT  8980.0 35975.0 9045.0 36040.0 ;
      RECT  8690.0 36692.5 9250.0 36757.5 ;
      RECT  8690.0 35347.5 9250.0 35412.5 ;
      RECT  9317.5 35542.5 9382.5 35347.5 ;
      RECT  9317.5 36382.5 9382.5 36757.5 ;
      RECT  9697.5 36382.5 9762.5 36757.5 ;
      RECT  9867.5 36540.0 9932.5 36725.0 ;
      RECT  9867.5 35380.0 9932.5 35565.0 ;
      RECT  9317.5 36382.5 9382.5 36517.5 ;
      RECT  9507.5 36382.5 9572.5 36517.5 ;
      RECT  9507.5 36382.5 9572.5 36517.5 ;
      RECT  9317.5 36382.5 9382.5 36517.5 ;
      RECT  9507.5 36382.5 9572.5 36517.5 ;
      RECT  9697.5 36382.5 9762.5 36517.5 ;
      RECT  9697.5 36382.5 9762.5 36517.5 ;
      RECT  9507.5 36382.5 9572.5 36517.5 ;
      RECT  9317.5 35542.5 9382.5 35677.5 ;
      RECT  9507.5 35542.5 9572.5 35677.5 ;
      RECT  9507.5 35542.5 9572.5 35677.5 ;
      RECT  9317.5 35542.5 9382.5 35677.5 ;
      RECT  9507.5 35542.5 9572.5 35677.5 ;
      RECT  9697.5 35542.5 9762.5 35677.5 ;
      RECT  9697.5 35542.5 9762.5 35677.5 ;
      RECT  9507.5 35542.5 9572.5 35677.5 ;
      RECT  9867.5 36472.5 9932.5 36607.5 ;
      RECT  9867.5 35497.5 9932.5 35632.5 ;
      RECT  9702.5 35772.5 9567.5 35837.5 ;
      RECT  9445.0 35987.5 9310.0 36052.5 ;
      RECT  9507.5 36382.5 9572.5 36517.5 ;
      RECT  9697.5 35542.5 9762.5 35677.5 ;
      RECT  9797.5 35987.5 9662.5 36052.5 ;
      RECT  9310.0 35987.5 9445.0 36052.5 ;
      RECT  9567.5 35772.5 9702.5 35837.5 ;
      RECT  9662.5 35987.5 9797.5 36052.5 ;
      RECT  9250.0 36692.5 10170.0 36757.5 ;
      RECT  9250.0 35347.5 10170.0 35412.5 ;
      RECT  10597.5 36540.0 10662.5 36725.0 ;
      RECT  10597.5 35380.0 10662.5 35565.0 ;
      RECT  10237.5 35497.5 10302.5 35347.5 ;
      RECT  10237.5 36382.5 10302.5 36757.5 ;
      RECT  10427.5 35497.5 10492.5 36382.5 ;
      RECT  10237.5 36382.5 10302.5 36517.5 ;
      RECT  10427.5 36382.5 10492.5 36517.5 ;
      RECT  10427.5 36382.5 10492.5 36517.5 ;
      RECT  10237.5 36382.5 10302.5 36517.5 ;
      RECT  10237.5 35497.5 10302.5 35632.5 ;
      RECT  10427.5 35497.5 10492.5 35632.5 ;
      RECT  10427.5 35497.5 10492.5 35632.5 ;
      RECT  10237.5 35497.5 10302.5 35632.5 ;
      RECT  10597.5 36472.5 10662.5 36607.5 ;
      RECT  10597.5 35497.5 10662.5 35632.5 ;
      RECT  10295.0 35940.0 10360.0 36075.0 ;
      RECT  10295.0 35940.0 10360.0 36075.0 ;
      RECT  10460.0 35975.0 10525.0 36040.0 ;
      RECT  10170.0 36692.5 10730.0 36757.5 ;
      RECT  10170.0 35347.5 10730.0 35412.5 ;
      RECT  8432.5 35940.0 8497.5 36075.0 ;
      RECT  8572.5 35667.5 8637.5 35802.5 ;
      RECT  9567.5 35772.5 9432.5 35837.5 ;
      RECT  9117.5 36910.0 9182.5 36725.0 ;
      RECT  9117.5 38070.0 9182.5 37885.0 ;
      RECT  8757.5 37952.5 8822.5 38102.5 ;
      RECT  8757.5 37067.5 8822.5 36692.5 ;
      RECT  8947.5 37952.5 9012.5 37067.5 ;
      RECT  8757.5 37067.5 8822.5 36932.5 ;
      RECT  8947.5 37067.5 9012.5 36932.5 ;
      RECT  8947.5 37067.5 9012.5 36932.5 ;
      RECT  8757.5 37067.5 8822.5 36932.5 ;
      RECT  8757.5 37952.5 8822.5 37817.5 ;
      RECT  8947.5 37952.5 9012.5 37817.5 ;
      RECT  8947.5 37952.5 9012.5 37817.5 ;
      RECT  8757.5 37952.5 8822.5 37817.5 ;
      RECT  9117.5 36977.5 9182.5 36842.5 ;
      RECT  9117.5 37952.5 9182.5 37817.5 ;
      RECT  8815.0 37510.0 8880.0 37375.0 ;
      RECT  8815.0 37510.0 8880.0 37375.0 ;
      RECT  8980.0 37475.0 9045.0 37410.0 ;
      RECT  8690.0 36757.5 9250.0 36692.5 ;
      RECT  8690.0 38102.5 9250.0 38037.5 ;
      RECT  9317.5 37907.5 9382.5 38102.5 ;
      RECT  9317.5 37067.5 9382.5 36692.5 ;
      RECT  9697.5 37067.5 9762.5 36692.5 ;
      RECT  9867.5 36910.0 9932.5 36725.0 ;
      RECT  9867.5 38070.0 9932.5 37885.0 ;
      RECT  9317.5 37067.5 9382.5 36932.5 ;
      RECT  9507.5 37067.5 9572.5 36932.5 ;
      RECT  9507.5 37067.5 9572.5 36932.5 ;
      RECT  9317.5 37067.5 9382.5 36932.5 ;
      RECT  9507.5 37067.5 9572.5 36932.5 ;
      RECT  9697.5 37067.5 9762.5 36932.5 ;
      RECT  9697.5 37067.5 9762.5 36932.5 ;
      RECT  9507.5 37067.5 9572.5 36932.5 ;
      RECT  9317.5 37907.5 9382.5 37772.5 ;
      RECT  9507.5 37907.5 9572.5 37772.5 ;
      RECT  9507.5 37907.5 9572.5 37772.5 ;
      RECT  9317.5 37907.5 9382.5 37772.5 ;
      RECT  9507.5 37907.5 9572.5 37772.5 ;
      RECT  9697.5 37907.5 9762.5 37772.5 ;
      RECT  9697.5 37907.5 9762.5 37772.5 ;
      RECT  9507.5 37907.5 9572.5 37772.5 ;
      RECT  9867.5 36977.5 9932.5 36842.5 ;
      RECT  9867.5 37952.5 9932.5 37817.5 ;
      RECT  9702.5 37677.5 9567.5 37612.5 ;
      RECT  9445.0 37462.5 9310.0 37397.5 ;
      RECT  9507.5 37067.5 9572.5 36932.5 ;
      RECT  9697.5 37907.5 9762.5 37772.5 ;
      RECT  9797.5 37462.5 9662.5 37397.5 ;
      RECT  9310.0 37462.5 9445.0 37397.5 ;
      RECT  9567.5 37677.5 9702.5 37612.5 ;
      RECT  9662.5 37462.5 9797.5 37397.5 ;
      RECT  9250.0 36757.5 10170.0 36692.5 ;
      RECT  9250.0 38102.5 10170.0 38037.5 ;
      RECT  10597.5 36910.0 10662.5 36725.0 ;
      RECT  10597.5 38070.0 10662.5 37885.0 ;
      RECT  10237.5 37952.5 10302.5 38102.5 ;
      RECT  10237.5 37067.5 10302.5 36692.5 ;
      RECT  10427.5 37952.5 10492.5 37067.5 ;
      RECT  10237.5 37067.5 10302.5 36932.5 ;
      RECT  10427.5 37067.5 10492.5 36932.5 ;
      RECT  10427.5 37067.5 10492.5 36932.5 ;
      RECT  10237.5 37067.5 10302.5 36932.5 ;
      RECT  10237.5 37952.5 10302.5 37817.5 ;
      RECT  10427.5 37952.5 10492.5 37817.5 ;
      RECT  10427.5 37952.5 10492.5 37817.5 ;
      RECT  10237.5 37952.5 10302.5 37817.5 ;
      RECT  10597.5 36977.5 10662.5 36842.5 ;
      RECT  10597.5 37952.5 10662.5 37817.5 ;
      RECT  10295.0 37510.0 10360.0 37375.0 ;
      RECT  10295.0 37510.0 10360.0 37375.0 ;
      RECT  10460.0 37475.0 10525.0 37410.0 ;
      RECT  10170.0 36757.5 10730.0 36692.5 ;
      RECT  10170.0 38102.5 10730.0 38037.5 ;
      RECT  8432.5 37375.0 8497.5 37510.0 ;
      RECT  8572.5 37647.5 8637.5 37782.5 ;
      RECT  9567.5 37612.5 9432.5 37677.5 ;
      RECT  9117.5 39230.0 9182.5 39415.0 ;
      RECT  9117.5 38070.0 9182.5 38255.0 ;
      RECT  8757.5 38187.5 8822.5 38037.5 ;
      RECT  8757.5 39072.5 8822.5 39447.5 ;
      RECT  8947.5 38187.5 9012.5 39072.5 ;
      RECT  8757.5 39072.5 8822.5 39207.5 ;
      RECT  8947.5 39072.5 9012.5 39207.5 ;
      RECT  8947.5 39072.5 9012.5 39207.5 ;
      RECT  8757.5 39072.5 8822.5 39207.5 ;
      RECT  8757.5 38187.5 8822.5 38322.5 ;
      RECT  8947.5 38187.5 9012.5 38322.5 ;
      RECT  8947.5 38187.5 9012.5 38322.5 ;
      RECT  8757.5 38187.5 8822.5 38322.5 ;
      RECT  9117.5 39162.5 9182.5 39297.5 ;
      RECT  9117.5 38187.5 9182.5 38322.5 ;
      RECT  8815.0 38630.0 8880.0 38765.0 ;
      RECT  8815.0 38630.0 8880.0 38765.0 ;
      RECT  8980.0 38665.0 9045.0 38730.0 ;
      RECT  8690.0 39382.5 9250.0 39447.5 ;
      RECT  8690.0 38037.5 9250.0 38102.5 ;
      RECT  9317.5 38232.5 9382.5 38037.5 ;
      RECT  9317.5 39072.5 9382.5 39447.5 ;
      RECT  9697.5 39072.5 9762.5 39447.5 ;
      RECT  9867.5 39230.0 9932.5 39415.0 ;
      RECT  9867.5 38070.0 9932.5 38255.0 ;
      RECT  9317.5 39072.5 9382.5 39207.5 ;
      RECT  9507.5 39072.5 9572.5 39207.5 ;
      RECT  9507.5 39072.5 9572.5 39207.5 ;
      RECT  9317.5 39072.5 9382.5 39207.5 ;
      RECT  9507.5 39072.5 9572.5 39207.5 ;
      RECT  9697.5 39072.5 9762.5 39207.5 ;
      RECT  9697.5 39072.5 9762.5 39207.5 ;
      RECT  9507.5 39072.5 9572.5 39207.5 ;
      RECT  9317.5 38232.5 9382.5 38367.5 ;
      RECT  9507.5 38232.5 9572.5 38367.5 ;
      RECT  9507.5 38232.5 9572.5 38367.5 ;
      RECT  9317.5 38232.5 9382.5 38367.5 ;
      RECT  9507.5 38232.5 9572.5 38367.5 ;
      RECT  9697.5 38232.5 9762.5 38367.5 ;
      RECT  9697.5 38232.5 9762.5 38367.5 ;
      RECT  9507.5 38232.5 9572.5 38367.5 ;
      RECT  9867.5 39162.5 9932.5 39297.5 ;
      RECT  9867.5 38187.5 9932.5 38322.5 ;
      RECT  9702.5 38462.5 9567.5 38527.5 ;
      RECT  9445.0 38677.5 9310.0 38742.5 ;
      RECT  9507.5 39072.5 9572.5 39207.5 ;
      RECT  9697.5 38232.5 9762.5 38367.5 ;
      RECT  9797.5 38677.5 9662.5 38742.5 ;
      RECT  9310.0 38677.5 9445.0 38742.5 ;
      RECT  9567.5 38462.5 9702.5 38527.5 ;
      RECT  9662.5 38677.5 9797.5 38742.5 ;
      RECT  9250.0 39382.5 10170.0 39447.5 ;
      RECT  9250.0 38037.5 10170.0 38102.5 ;
      RECT  10597.5 39230.0 10662.5 39415.0 ;
      RECT  10597.5 38070.0 10662.5 38255.0 ;
      RECT  10237.5 38187.5 10302.5 38037.5 ;
      RECT  10237.5 39072.5 10302.5 39447.5 ;
      RECT  10427.5 38187.5 10492.5 39072.5 ;
      RECT  10237.5 39072.5 10302.5 39207.5 ;
      RECT  10427.5 39072.5 10492.5 39207.5 ;
      RECT  10427.5 39072.5 10492.5 39207.5 ;
      RECT  10237.5 39072.5 10302.5 39207.5 ;
      RECT  10237.5 38187.5 10302.5 38322.5 ;
      RECT  10427.5 38187.5 10492.5 38322.5 ;
      RECT  10427.5 38187.5 10492.5 38322.5 ;
      RECT  10237.5 38187.5 10302.5 38322.5 ;
      RECT  10597.5 39162.5 10662.5 39297.5 ;
      RECT  10597.5 38187.5 10662.5 38322.5 ;
      RECT  10295.0 38630.0 10360.0 38765.0 ;
      RECT  10295.0 38630.0 10360.0 38765.0 ;
      RECT  10460.0 38665.0 10525.0 38730.0 ;
      RECT  10170.0 39382.5 10730.0 39447.5 ;
      RECT  10170.0 38037.5 10730.0 38102.5 ;
      RECT  8432.5 38630.0 8497.5 38765.0 ;
      RECT  8572.5 38357.5 8637.5 38492.5 ;
      RECT  9567.5 38462.5 9432.5 38527.5 ;
      RECT  9117.5 39600.0 9182.5 39415.0 ;
      RECT  9117.5 40760.0 9182.5 40575.0 ;
      RECT  8757.5 40642.5 8822.5 40792.5 ;
      RECT  8757.5 39757.5 8822.5 39382.5 ;
      RECT  8947.5 40642.5 9012.5 39757.5 ;
      RECT  8757.5 39757.5 8822.5 39622.5 ;
      RECT  8947.5 39757.5 9012.5 39622.5 ;
      RECT  8947.5 39757.5 9012.5 39622.5 ;
      RECT  8757.5 39757.5 8822.5 39622.5 ;
      RECT  8757.5 40642.5 8822.5 40507.5 ;
      RECT  8947.5 40642.5 9012.5 40507.5 ;
      RECT  8947.5 40642.5 9012.5 40507.5 ;
      RECT  8757.5 40642.5 8822.5 40507.5 ;
      RECT  9117.5 39667.5 9182.5 39532.5 ;
      RECT  9117.5 40642.5 9182.5 40507.5 ;
      RECT  8815.0 40200.0 8880.0 40065.0 ;
      RECT  8815.0 40200.0 8880.0 40065.0 ;
      RECT  8980.0 40165.0 9045.0 40100.0 ;
      RECT  8690.0 39447.5 9250.0 39382.5 ;
      RECT  8690.0 40792.5 9250.0 40727.5 ;
      RECT  9317.5 40597.5 9382.5 40792.5 ;
      RECT  9317.5 39757.5 9382.5 39382.5 ;
      RECT  9697.5 39757.5 9762.5 39382.5 ;
      RECT  9867.5 39600.0 9932.5 39415.0 ;
      RECT  9867.5 40760.0 9932.5 40575.0 ;
      RECT  9317.5 39757.5 9382.5 39622.5 ;
      RECT  9507.5 39757.5 9572.5 39622.5 ;
      RECT  9507.5 39757.5 9572.5 39622.5 ;
      RECT  9317.5 39757.5 9382.5 39622.5 ;
      RECT  9507.5 39757.5 9572.5 39622.5 ;
      RECT  9697.5 39757.5 9762.5 39622.5 ;
      RECT  9697.5 39757.5 9762.5 39622.5 ;
      RECT  9507.5 39757.5 9572.5 39622.5 ;
      RECT  9317.5 40597.5 9382.5 40462.5 ;
      RECT  9507.5 40597.5 9572.5 40462.5 ;
      RECT  9507.5 40597.5 9572.5 40462.5 ;
      RECT  9317.5 40597.5 9382.5 40462.5 ;
      RECT  9507.5 40597.5 9572.5 40462.5 ;
      RECT  9697.5 40597.5 9762.5 40462.5 ;
      RECT  9697.5 40597.5 9762.5 40462.5 ;
      RECT  9507.5 40597.5 9572.5 40462.5 ;
      RECT  9867.5 39667.5 9932.5 39532.5 ;
      RECT  9867.5 40642.5 9932.5 40507.5 ;
      RECT  9702.5 40367.5 9567.5 40302.5 ;
      RECT  9445.0 40152.5 9310.0 40087.5 ;
      RECT  9507.5 39757.5 9572.5 39622.5 ;
      RECT  9697.5 40597.5 9762.5 40462.5 ;
      RECT  9797.5 40152.5 9662.5 40087.5 ;
      RECT  9310.0 40152.5 9445.0 40087.5 ;
      RECT  9567.5 40367.5 9702.5 40302.5 ;
      RECT  9662.5 40152.5 9797.5 40087.5 ;
      RECT  9250.0 39447.5 10170.0 39382.5 ;
      RECT  9250.0 40792.5 10170.0 40727.5 ;
      RECT  10597.5 39600.0 10662.5 39415.0 ;
      RECT  10597.5 40760.0 10662.5 40575.0 ;
      RECT  10237.5 40642.5 10302.5 40792.5 ;
      RECT  10237.5 39757.5 10302.5 39382.5 ;
      RECT  10427.5 40642.5 10492.5 39757.5 ;
      RECT  10237.5 39757.5 10302.5 39622.5 ;
      RECT  10427.5 39757.5 10492.5 39622.5 ;
      RECT  10427.5 39757.5 10492.5 39622.5 ;
      RECT  10237.5 39757.5 10302.5 39622.5 ;
      RECT  10237.5 40642.5 10302.5 40507.5 ;
      RECT  10427.5 40642.5 10492.5 40507.5 ;
      RECT  10427.5 40642.5 10492.5 40507.5 ;
      RECT  10237.5 40642.5 10302.5 40507.5 ;
      RECT  10597.5 39667.5 10662.5 39532.5 ;
      RECT  10597.5 40642.5 10662.5 40507.5 ;
      RECT  10295.0 40200.0 10360.0 40065.0 ;
      RECT  10295.0 40200.0 10360.0 40065.0 ;
      RECT  10460.0 40165.0 10525.0 40100.0 ;
      RECT  10170.0 39447.5 10730.0 39382.5 ;
      RECT  10170.0 40792.5 10730.0 40727.5 ;
      RECT  8432.5 40065.0 8497.5 40200.0 ;
      RECT  8572.5 40337.5 8637.5 40472.5 ;
      RECT  9567.5 40302.5 9432.5 40367.5 ;
      RECT  9117.5 41920.0 9182.5 42105.0 ;
      RECT  9117.5 40760.0 9182.5 40945.0 ;
      RECT  8757.5 40877.5 8822.5 40727.5 ;
      RECT  8757.5 41762.5 8822.5 42137.5 ;
      RECT  8947.5 40877.5 9012.5 41762.5 ;
      RECT  8757.5 41762.5 8822.5 41897.5 ;
      RECT  8947.5 41762.5 9012.5 41897.5 ;
      RECT  8947.5 41762.5 9012.5 41897.5 ;
      RECT  8757.5 41762.5 8822.5 41897.5 ;
      RECT  8757.5 40877.5 8822.5 41012.5 ;
      RECT  8947.5 40877.5 9012.5 41012.5 ;
      RECT  8947.5 40877.5 9012.5 41012.5 ;
      RECT  8757.5 40877.5 8822.5 41012.5 ;
      RECT  9117.5 41852.5 9182.5 41987.5 ;
      RECT  9117.5 40877.5 9182.5 41012.5 ;
      RECT  8815.0 41320.0 8880.0 41455.0 ;
      RECT  8815.0 41320.0 8880.0 41455.0 ;
      RECT  8980.0 41355.0 9045.0 41420.0 ;
      RECT  8690.0 42072.5 9250.0 42137.5 ;
      RECT  8690.0 40727.5 9250.0 40792.5 ;
      RECT  9317.5 40922.5 9382.5 40727.5 ;
      RECT  9317.5 41762.5 9382.5 42137.5 ;
      RECT  9697.5 41762.5 9762.5 42137.5 ;
      RECT  9867.5 41920.0 9932.5 42105.0 ;
      RECT  9867.5 40760.0 9932.5 40945.0 ;
      RECT  9317.5 41762.5 9382.5 41897.5 ;
      RECT  9507.5 41762.5 9572.5 41897.5 ;
      RECT  9507.5 41762.5 9572.5 41897.5 ;
      RECT  9317.5 41762.5 9382.5 41897.5 ;
      RECT  9507.5 41762.5 9572.5 41897.5 ;
      RECT  9697.5 41762.5 9762.5 41897.5 ;
      RECT  9697.5 41762.5 9762.5 41897.5 ;
      RECT  9507.5 41762.5 9572.5 41897.5 ;
      RECT  9317.5 40922.5 9382.5 41057.5 ;
      RECT  9507.5 40922.5 9572.5 41057.5 ;
      RECT  9507.5 40922.5 9572.5 41057.5 ;
      RECT  9317.5 40922.5 9382.5 41057.5 ;
      RECT  9507.5 40922.5 9572.5 41057.5 ;
      RECT  9697.5 40922.5 9762.5 41057.5 ;
      RECT  9697.5 40922.5 9762.5 41057.5 ;
      RECT  9507.5 40922.5 9572.5 41057.5 ;
      RECT  9867.5 41852.5 9932.5 41987.5 ;
      RECT  9867.5 40877.5 9932.5 41012.5 ;
      RECT  9702.5 41152.5 9567.5 41217.5 ;
      RECT  9445.0 41367.5 9310.0 41432.5 ;
      RECT  9507.5 41762.5 9572.5 41897.5 ;
      RECT  9697.5 40922.5 9762.5 41057.5 ;
      RECT  9797.5 41367.5 9662.5 41432.5 ;
      RECT  9310.0 41367.5 9445.0 41432.5 ;
      RECT  9567.5 41152.5 9702.5 41217.5 ;
      RECT  9662.5 41367.5 9797.5 41432.5 ;
      RECT  9250.0 42072.5 10170.0 42137.5 ;
      RECT  9250.0 40727.5 10170.0 40792.5 ;
      RECT  10597.5 41920.0 10662.5 42105.0 ;
      RECT  10597.5 40760.0 10662.5 40945.0 ;
      RECT  10237.5 40877.5 10302.5 40727.5 ;
      RECT  10237.5 41762.5 10302.5 42137.5 ;
      RECT  10427.5 40877.5 10492.5 41762.5 ;
      RECT  10237.5 41762.5 10302.5 41897.5 ;
      RECT  10427.5 41762.5 10492.5 41897.5 ;
      RECT  10427.5 41762.5 10492.5 41897.5 ;
      RECT  10237.5 41762.5 10302.5 41897.5 ;
      RECT  10237.5 40877.5 10302.5 41012.5 ;
      RECT  10427.5 40877.5 10492.5 41012.5 ;
      RECT  10427.5 40877.5 10492.5 41012.5 ;
      RECT  10237.5 40877.5 10302.5 41012.5 ;
      RECT  10597.5 41852.5 10662.5 41987.5 ;
      RECT  10597.5 40877.5 10662.5 41012.5 ;
      RECT  10295.0 41320.0 10360.0 41455.0 ;
      RECT  10295.0 41320.0 10360.0 41455.0 ;
      RECT  10460.0 41355.0 10525.0 41420.0 ;
      RECT  10170.0 42072.5 10730.0 42137.5 ;
      RECT  10170.0 40727.5 10730.0 40792.5 ;
      RECT  8432.5 41320.0 8497.5 41455.0 ;
      RECT  8572.5 41047.5 8637.5 41182.5 ;
      RECT  9567.5 41152.5 9432.5 41217.5 ;
      RECT  9117.5 42290.0 9182.5 42105.0 ;
      RECT  9117.5 43450.0 9182.5 43265.0 ;
      RECT  8757.5 43332.5 8822.5 43482.5 ;
      RECT  8757.5 42447.5 8822.5 42072.5 ;
      RECT  8947.5 43332.5 9012.5 42447.5 ;
      RECT  8757.5 42447.5 8822.5 42312.5 ;
      RECT  8947.5 42447.5 9012.5 42312.5 ;
      RECT  8947.5 42447.5 9012.5 42312.5 ;
      RECT  8757.5 42447.5 8822.5 42312.5 ;
      RECT  8757.5 43332.5 8822.5 43197.5 ;
      RECT  8947.5 43332.5 9012.5 43197.5 ;
      RECT  8947.5 43332.5 9012.5 43197.5 ;
      RECT  8757.5 43332.5 8822.5 43197.5 ;
      RECT  9117.5 42357.5 9182.5 42222.5 ;
      RECT  9117.5 43332.5 9182.5 43197.5 ;
      RECT  8815.0 42890.0 8880.0 42755.0 ;
      RECT  8815.0 42890.0 8880.0 42755.0 ;
      RECT  8980.0 42855.0 9045.0 42790.0 ;
      RECT  8690.0 42137.5 9250.0 42072.5 ;
      RECT  8690.0 43482.5 9250.0 43417.5 ;
      RECT  9317.5 43287.5 9382.5 43482.5 ;
      RECT  9317.5 42447.5 9382.5 42072.5 ;
      RECT  9697.5 42447.5 9762.5 42072.5 ;
      RECT  9867.5 42290.0 9932.5 42105.0 ;
      RECT  9867.5 43450.0 9932.5 43265.0 ;
      RECT  9317.5 42447.5 9382.5 42312.5 ;
      RECT  9507.5 42447.5 9572.5 42312.5 ;
      RECT  9507.5 42447.5 9572.5 42312.5 ;
      RECT  9317.5 42447.5 9382.5 42312.5 ;
      RECT  9507.5 42447.5 9572.5 42312.5 ;
      RECT  9697.5 42447.5 9762.5 42312.5 ;
      RECT  9697.5 42447.5 9762.5 42312.5 ;
      RECT  9507.5 42447.5 9572.5 42312.5 ;
      RECT  9317.5 43287.5 9382.5 43152.5 ;
      RECT  9507.5 43287.5 9572.5 43152.5 ;
      RECT  9507.5 43287.5 9572.5 43152.5 ;
      RECT  9317.5 43287.5 9382.5 43152.5 ;
      RECT  9507.5 43287.5 9572.5 43152.5 ;
      RECT  9697.5 43287.5 9762.5 43152.5 ;
      RECT  9697.5 43287.5 9762.5 43152.5 ;
      RECT  9507.5 43287.5 9572.5 43152.5 ;
      RECT  9867.5 42357.5 9932.5 42222.5 ;
      RECT  9867.5 43332.5 9932.5 43197.5 ;
      RECT  9702.5 43057.5 9567.5 42992.5 ;
      RECT  9445.0 42842.5 9310.0 42777.5 ;
      RECT  9507.5 42447.5 9572.5 42312.5 ;
      RECT  9697.5 43287.5 9762.5 43152.5 ;
      RECT  9797.5 42842.5 9662.5 42777.5 ;
      RECT  9310.0 42842.5 9445.0 42777.5 ;
      RECT  9567.5 43057.5 9702.5 42992.5 ;
      RECT  9662.5 42842.5 9797.5 42777.5 ;
      RECT  9250.0 42137.5 10170.0 42072.5 ;
      RECT  9250.0 43482.5 10170.0 43417.5 ;
      RECT  10597.5 42290.0 10662.5 42105.0 ;
      RECT  10597.5 43450.0 10662.5 43265.0 ;
      RECT  10237.5 43332.5 10302.5 43482.5 ;
      RECT  10237.5 42447.5 10302.5 42072.5 ;
      RECT  10427.5 43332.5 10492.5 42447.5 ;
      RECT  10237.5 42447.5 10302.5 42312.5 ;
      RECT  10427.5 42447.5 10492.5 42312.5 ;
      RECT  10427.5 42447.5 10492.5 42312.5 ;
      RECT  10237.5 42447.5 10302.5 42312.5 ;
      RECT  10237.5 43332.5 10302.5 43197.5 ;
      RECT  10427.5 43332.5 10492.5 43197.5 ;
      RECT  10427.5 43332.5 10492.5 43197.5 ;
      RECT  10237.5 43332.5 10302.5 43197.5 ;
      RECT  10597.5 42357.5 10662.5 42222.5 ;
      RECT  10597.5 43332.5 10662.5 43197.5 ;
      RECT  10295.0 42890.0 10360.0 42755.0 ;
      RECT  10295.0 42890.0 10360.0 42755.0 ;
      RECT  10460.0 42855.0 10525.0 42790.0 ;
      RECT  10170.0 42137.5 10730.0 42072.5 ;
      RECT  10170.0 43482.5 10730.0 43417.5 ;
      RECT  8432.5 42755.0 8497.5 42890.0 ;
      RECT  8572.5 43027.5 8637.5 43162.5 ;
      RECT  9567.5 42992.5 9432.5 43057.5 ;
      RECT  9117.5 44610.0 9182.5 44795.0 ;
      RECT  9117.5 43450.0 9182.5 43635.0 ;
      RECT  8757.5 43567.5 8822.5 43417.5 ;
      RECT  8757.5 44452.5 8822.5 44827.5 ;
      RECT  8947.5 43567.5 9012.5 44452.5 ;
      RECT  8757.5 44452.5 8822.5 44587.5 ;
      RECT  8947.5 44452.5 9012.5 44587.5 ;
      RECT  8947.5 44452.5 9012.5 44587.5 ;
      RECT  8757.5 44452.5 8822.5 44587.5 ;
      RECT  8757.5 43567.5 8822.5 43702.5 ;
      RECT  8947.5 43567.5 9012.5 43702.5 ;
      RECT  8947.5 43567.5 9012.5 43702.5 ;
      RECT  8757.5 43567.5 8822.5 43702.5 ;
      RECT  9117.5 44542.5 9182.5 44677.5 ;
      RECT  9117.5 43567.5 9182.5 43702.5 ;
      RECT  8815.0 44010.0 8880.0 44145.0 ;
      RECT  8815.0 44010.0 8880.0 44145.0 ;
      RECT  8980.0 44045.0 9045.0 44110.0 ;
      RECT  8690.0 44762.5 9250.0 44827.5 ;
      RECT  8690.0 43417.5 9250.0 43482.5 ;
      RECT  9317.5 43612.5 9382.5 43417.5 ;
      RECT  9317.5 44452.5 9382.5 44827.5 ;
      RECT  9697.5 44452.5 9762.5 44827.5 ;
      RECT  9867.5 44610.0 9932.5 44795.0 ;
      RECT  9867.5 43450.0 9932.5 43635.0 ;
      RECT  9317.5 44452.5 9382.5 44587.5 ;
      RECT  9507.5 44452.5 9572.5 44587.5 ;
      RECT  9507.5 44452.5 9572.5 44587.5 ;
      RECT  9317.5 44452.5 9382.5 44587.5 ;
      RECT  9507.5 44452.5 9572.5 44587.5 ;
      RECT  9697.5 44452.5 9762.5 44587.5 ;
      RECT  9697.5 44452.5 9762.5 44587.5 ;
      RECT  9507.5 44452.5 9572.5 44587.5 ;
      RECT  9317.5 43612.5 9382.5 43747.5 ;
      RECT  9507.5 43612.5 9572.5 43747.5 ;
      RECT  9507.5 43612.5 9572.5 43747.5 ;
      RECT  9317.5 43612.5 9382.5 43747.5 ;
      RECT  9507.5 43612.5 9572.5 43747.5 ;
      RECT  9697.5 43612.5 9762.5 43747.5 ;
      RECT  9697.5 43612.5 9762.5 43747.5 ;
      RECT  9507.5 43612.5 9572.5 43747.5 ;
      RECT  9867.5 44542.5 9932.5 44677.5 ;
      RECT  9867.5 43567.5 9932.5 43702.5 ;
      RECT  9702.5 43842.5 9567.5 43907.5 ;
      RECT  9445.0 44057.5 9310.0 44122.5 ;
      RECT  9507.5 44452.5 9572.5 44587.5 ;
      RECT  9697.5 43612.5 9762.5 43747.5 ;
      RECT  9797.5 44057.5 9662.5 44122.5 ;
      RECT  9310.0 44057.5 9445.0 44122.5 ;
      RECT  9567.5 43842.5 9702.5 43907.5 ;
      RECT  9662.5 44057.5 9797.5 44122.5 ;
      RECT  9250.0 44762.5 10170.0 44827.5 ;
      RECT  9250.0 43417.5 10170.0 43482.5 ;
      RECT  10597.5 44610.0 10662.5 44795.0 ;
      RECT  10597.5 43450.0 10662.5 43635.0 ;
      RECT  10237.5 43567.5 10302.5 43417.5 ;
      RECT  10237.5 44452.5 10302.5 44827.5 ;
      RECT  10427.5 43567.5 10492.5 44452.5 ;
      RECT  10237.5 44452.5 10302.5 44587.5 ;
      RECT  10427.5 44452.5 10492.5 44587.5 ;
      RECT  10427.5 44452.5 10492.5 44587.5 ;
      RECT  10237.5 44452.5 10302.5 44587.5 ;
      RECT  10237.5 43567.5 10302.5 43702.5 ;
      RECT  10427.5 43567.5 10492.5 43702.5 ;
      RECT  10427.5 43567.5 10492.5 43702.5 ;
      RECT  10237.5 43567.5 10302.5 43702.5 ;
      RECT  10597.5 44542.5 10662.5 44677.5 ;
      RECT  10597.5 43567.5 10662.5 43702.5 ;
      RECT  10295.0 44010.0 10360.0 44145.0 ;
      RECT  10295.0 44010.0 10360.0 44145.0 ;
      RECT  10460.0 44045.0 10525.0 44110.0 ;
      RECT  10170.0 44762.5 10730.0 44827.5 ;
      RECT  10170.0 43417.5 10730.0 43482.5 ;
      RECT  8432.5 44010.0 8497.5 44145.0 ;
      RECT  8572.5 43737.5 8637.5 43872.5 ;
      RECT  9567.5 43842.5 9432.5 43907.5 ;
      RECT  9117.5 44980.0 9182.5 44795.0 ;
      RECT  9117.5 46140.0 9182.5 45955.0 ;
      RECT  8757.5 46022.5 8822.5 46172.5 ;
      RECT  8757.5 45137.5 8822.5 44762.5 ;
      RECT  8947.5 46022.5 9012.5 45137.5 ;
      RECT  8757.5 45137.5 8822.5 45002.5 ;
      RECT  8947.5 45137.5 9012.5 45002.5 ;
      RECT  8947.5 45137.5 9012.5 45002.5 ;
      RECT  8757.5 45137.5 8822.5 45002.5 ;
      RECT  8757.5 46022.5 8822.5 45887.5 ;
      RECT  8947.5 46022.5 9012.5 45887.5 ;
      RECT  8947.5 46022.5 9012.5 45887.5 ;
      RECT  8757.5 46022.5 8822.5 45887.5 ;
      RECT  9117.5 45047.5 9182.5 44912.5 ;
      RECT  9117.5 46022.5 9182.5 45887.5 ;
      RECT  8815.0 45580.0 8880.0 45445.0 ;
      RECT  8815.0 45580.0 8880.0 45445.0 ;
      RECT  8980.0 45545.0 9045.0 45480.0 ;
      RECT  8690.0 44827.5 9250.0 44762.5 ;
      RECT  8690.0 46172.5 9250.0 46107.5 ;
      RECT  9317.5 45977.5 9382.5 46172.5 ;
      RECT  9317.5 45137.5 9382.5 44762.5 ;
      RECT  9697.5 45137.5 9762.5 44762.5 ;
      RECT  9867.5 44980.0 9932.5 44795.0 ;
      RECT  9867.5 46140.0 9932.5 45955.0 ;
      RECT  9317.5 45137.5 9382.5 45002.5 ;
      RECT  9507.5 45137.5 9572.5 45002.5 ;
      RECT  9507.5 45137.5 9572.5 45002.5 ;
      RECT  9317.5 45137.5 9382.5 45002.5 ;
      RECT  9507.5 45137.5 9572.5 45002.5 ;
      RECT  9697.5 45137.5 9762.5 45002.5 ;
      RECT  9697.5 45137.5 9762.5 45002.5 ;
      RECT  9507.5 45137.5 9572.5 45002.5 ;
      RECT  9317.5 45977.5 9382.5 45842.5 ;
      RECT  9507.5 45977.5 9572.5 45842.5 ;
      RECT  9507.5 45977.5 9572.5 45842.5 ;
      RECT  9317.5 45977.5 9382.5 45842.5 ;
      RECT  9507.5 45977.5 9572.5 45842.5 ;
      RECT  9697.5 45977.5 9762.5 45842.5 ;
      RECT  9697.5 45977.5 9762.5 45842.5 ;
      RECT  9507.5 45977.5 9572.5 45842.5 ;
      RECT  9867.5 45047.5 9932.5 44912.5 ;
      RECT  9867.5 46022.5 9932.5 45887.5 ;
      RECT  9702.5 45747.5 9567.5 45682.5 ;
      RECT  9445.0 45532.5 9310.0 45467.5 ;
      RECT  9507.5 45137.5 9572.5 45002.5 ;
      RECT  9697.5 45977.5 9762.5 45842.5 ;
      RECT  9797.5 45532.5 9662.5 45467.5 ;
      RECT  9310.0 45532.5 9445.0 45467.5 ;
      RECT  9567.5 45747.5 9702.5 45682.5 ;
      RECT  9662.5 45532.5 9797.5 45467.5 ;
      RECT  9250.0 44827.5 10170.0 44762.5 ;
      RECT  9250.0 46172.5 10170.0 46107.5 ;
      RECT  10597.5 44980.0 10662.5 44795.0 ;
      RECT  10597.5 46140.0 10662.5 45955.0 ;
      RECT  10237.5 46022.5 10302.5 46172.5 ;
      RECT  10237.5 45137.5 10302.5 44762.5 ;
      RECT  10427.5 46022.5 10492.5 45137.5 ;
      RECT  10237.5 45137.5 10302.5 45002.5 ;
      RECT  10427.5 45137.5 10492.5 45002.5 ;
      RECT  10427.5 45137.5 10492.5 45002.5 ;
      RECT  10237.5 45137.5 10302.5 45002.5 ;
      RECT  10237.5 46022.5 10302.5 45887.5 ;
      RECT  10427.5 46022.5 10492.5 45887.5 ;
      RECT  10427.5 46022.5 10492.5 45887.5 ;
      RECT  10237.5 46022.5 10302.5 45887.5 ;
      RECT  10597.5 45047.5 10662.5 44912.5 ;
      RECT  10597.5 46022.5 10662.5 45887.5 ;
      RECT  10295.0 45580.0 10360.0 45445.0 ;
      RECT  10295.0 45580.0 10360.0 45445.0 ;
      RECT  10460.0 45545.0 10525.0 45480.0 ;
      RECT  10170.0 44827.5 10730.0 44762.5 ;
      RECT  10170.0 46172.5 10730.0 46107.5 ;
      RECT  8432.5 45445.0 8497.5 45580.0 ;
      RECT  8572.5 45717.5 8637.5 45852.5 ;
      RECT  9567.5 45682.5 9432.5 45747.5 ;
      RECT  9117.5 47300.0 9182.5 47485.0 ;
      RECT  9117.5 46140.0 9182.5 46325.0 ;
      RECT  8757.5 46257.5 8822.5 46107.5 ;
      RECT  8757.5 47142.5 8822.5 47517.5 ;
      RECT  8947.5 46257.5 9012.5 47142.5 ;
      RECT  8757.5 47142.5 8822.5 47277.5 ;
      RECT  8947.5 47142.5 9012.5 47277.5 ;
      RECT  8947.5 47142.5 9012.5 47277.5 ;
      RECT  8757.5 47142.5 8822.5 47277.5 ;
      RECT  8757.5 46257.5 8822.5 46392.5 ;
      RECT  8947.5 46257.5 9012.5 46392.5 ;
      RECT  8947.5 46257.5 9012.5 46392.5 ;
      RECT  8757.5 46257.5 8822.5 46392.5 ;
      RECT  9117.5 47232.5 9182.5 47367.5 ;
      RECT  9117.5 46257.5 9182.5 46392.5 ;
      RECT  8815.0 46700.0 8880.0 46835.0 ;
      RECT  8815.0 46700.0 8880.0 46835.0 ;
      RECT  8980.0 46735.0 9045.0 46800.0 ;
      RECT  8690.0 47452.5 9250.0 47517.5 ;
      RECT  8690.0 46107.5 9250.0 46172.5 ;
      RECT  9317.5 46302.5 9382.5 46107.5 ;
      RECT  9317.5 47142.5 9382.5 47517.5 ;
      RECT  9697.5 47142.5 9762.5 47517.5 ;
      RECT  9867.5 47300.0 9932.5 47485.0 ;
      RECT  9867.5 46140.0 9932.5 46325.0 ;
      RECT  9317.5 47142.5 9382.5 47277.5 ;
      RECT  9507.5 47142.5 9572.5 47277.5 ;
      RECT  9507.5 47142.5 9572.5 47277.5 ;
      RECT  9317.5 47142.5 9382.5 47277.5 ;
      RECT  9507.5 47142.5 9572.5 47277.5 ;
      RECT  9697.5 47142.5 9762.5 47277.5 ;
      RECT  9697.5 47142.5 9762.5 47277.5 ;
      RECT  9507.5 47142.5 9572.5 47277.5 ;
      RECT  9317.5 46302.5 9382.5 46437.5 ;
      RECT  9507.5 46302.5 9572.5 46437.5 ;
      RECT  9507.5 46302.5 9572.5 46437.5 ;
      RECT  9317.5 46302.5 9382.5 46437.5 ;
      RECT  9507.5 46302.5 9572.5 46437.5 ;
      RECT  9697.5 46302.5 9762.5 46437.5 ;
      RECT  9697.5 46302.5 9762.5 46437.5 ;
      RECT  9507.5 46302.5 9572.5 46437.5 ;
      RECT  9867.5 47232.5 9932.5 47367.5 ;
      RECT  9867.5 46257.5 9932.5 46392.5 ;
      RECT  9702.5 46532.5 9567.5 46597.5 ;
      RECT  9445.0 46747.5 9310.0 46812.5 ;
      RECT  9507.5 47142.5 9572.5 47277.5 ;
      RECT  9697.5 46302.5 9762.5 46437.5 ;
      RECT  9797.5 46747.5 9662.5 46812.5 ;
      RECT  9310.0 46747.5 9445.0 46812.5 ;
      RECT  9567.5 46532.5 9702.5 46597.5 ;
      RECT  9662.5 46747.5 9797.5 46812.5 ;
      RECT  9250.0 47452.5 10170.0 47517.5 ;
      RECT  9250.0 46107.5 10170.0 46172.5 ;
      RECT  10597.5 47300.0 10662.5 47485.0 ;
      RECT  10597.5 46140.0 10662.5 46325.0 ;
      RECT  10237.5 46257.5 10302.5 46107.5 ;
      RECT  10237.5 47142.5 10302.5 47517.5 ;
      RECT  10427.5 46257.5 10492.5 47142.5 ;
      RECT  10237.5 47142.5 10302.5 47277.5 ;
      RECT  10427.5 47142.5 10492.5 47277.5 ;
      RECT  10427.5 47142.5 10492.5 47277.5 ;
      RECT  10237.5 47142.5 10302.5 47277.5 ;
      RECT  10237.5 46257.5 10302.5 46392.5 ;
      RECT  10427.5 46257.5 10492.5 46392.5 ;
      RECT  10427.5 46257.5 10492.5 46392.5 ;
      RECT  10237.5 46257.5 10302.5 46392.5 ;
      RECT  10597.5 47232.5 10662.5 47367.5 ;
      RECT  10597.5 46257.5 10662.5 46392.5 ;
      RECT  10295.0 46700.0 10360.0 46835.0 ;
      RECT  10295.0 46700.0 10360.0 46835.0 ;
      RECT  10460.0 46735.0 10525.0 46800.0 ;
      RECT  10170.0 47452.5 10730.0 47517.5 ;
      RECT  10170.0 46107.5 10730.0 46172.5 ;
      RECT  8432.5 46700.0 8497.5 46835.0 ;
      RECT  8572.5 46427.5 8637.5 46562.5 ;
      RECT  9567.5 46532.5 9432.5 46597.5 ;
      RECT  9117.5 47670.0 9182.5 47485.0 ;
      RECT  9117.5 48830.0 9182.5 48645.0 ;
      RECT  8757.5 48712.5 8822.5 48862.5 ;
      RECT  8757.5 47827.5 8822.5 47452.5 ;
      RECT  8947.5 48712.5 9012.5 47827.5 ;
      RECT  8757.5 47827.5 8822.5 47692.5 ;
      RECT  8947.5 47827.5 9012.5 47692.5 ;
      RECT  8947.5 47827.5 9012.5 47692.5 ;
      RECT  8757.5 47827.5 8822.5 47692.5 ;
      RECT  8757.5 48712.5 8822.5 48577.5 ;
      RECT  8947.5 48712.5 9012.5 48577.5 ;
      RECT  8947.5 48712.5 9012.5 48577.5 ;
      RECT  8757.5 48712.5 8822.5 48577.5 ;
      RECT  9117.5 47737.5 9182.5 47602.5 ;
      RECT  9117.5 48712.5 9182.5 48577.5 ;
      RECT  8815.0 48270.0 8880.0 48135.0 ;
      RECT  8815.0 48270.0 8880.0 48135.0 ;
      RECT  8980.0 48235.0 9045.0 48170.0 ;
      RECT  8690.0 47517.5 9250.0 47452.5 ;
      RECT  8690.0 48862.5 9250.0 48797.5 ;
      RECT  9317.5 48667.5 9382.5 48862.5 ;
      RECT  9317.5 47827.5 9382.5 47452.5 ;
      RECT  9697.5 47827.5 9762.5 47452.5 ;
      RECT  9867.5 47670.0 9932.5 47485.0 ;
      RECT  9867.5 48830.0 9932.5 48645.0 ;
      RECT  9317.5 47827.5 9382.5 47692.5 ;
      RECT  9507.5 47827.5 9572.5 47692.5 ;
      RECT  9507.5 47827.5 9572.5 47692.5 ;
      RECT  9317.5 47827.5 9382.5 47692.5 ;
      RECT  9507.5 47827.5 9572.5 47692.5 ;
      RECT  9697.5 47827.5 9762.5 47692.5 ;
      RECT  9697.5 47827.5 9762.5 47692.5 ;
      RECT  9507.5 47827.5 9572.5 47692.5 ;
      RECT  9317.5 48667.5 9382.5 48532.5 ;
      RECT  9507.5 48667.5 9572.5 48532.5 ;
      RECT  9507.5 48667.5 9572.5 48532.5 ;
      RECT  9317.5 48667.5 9382.5 48532.5 ;
      RECT  9507.5 48667.5 9572.5 48532.5 ;
      RECT  9697.5 48667.5 9762.5 48532.5 ;
      RECT  9697.5 48667.5 9762.5 48532.5 ;
      RECT  9507.5 48667.5 9572.5 48532.5 ;
      RECT  9867.5 47737.5 9932.5 47602.5 ;
      RECT  9867.5 48712.5 9932.5 48577.5 ;
      RECT  9702.5 48437.5 9567.5 48372.5 ;
      RECT  9445.0 48222.5 9310.0 48157.5 ;
      RECT  9507.5 47827.5 9572.5 47692.5 ;
      RECT  9697.5 48667.5 9762.5 48532.5 ;
      RECT  9797.5 48222.5 9662.5 48157.5 ;
      RECT  9310.0 48222.5 9445.0 48157.5 ;
      RECT  9567.5 48437.5 9702.5 48372.5 ;
      RECT  9662.5 48222.5 9797.5 48157.5 ;
      RECT  9250.0 47517.5 10170.0 47452.5 ;
      RECT  9250.0 48862.5 10170.0 48797.5 ;
      RECT  10597.5 47670.0 10662.5 47485.0 ;
      RECT  10597.5 48830.0 10662.5 48645.0 ;
      RECT  10237.5 48712.5 10302.5 48862.5 ;
      RECT  10237.5 47827.5 10302.5 47452.5 ;
      RECT  10427.5 48712.5 10492.5 47827.5 ;
      RECT  10237.5 47827.5 10302.5 47692.5 ;
      RECT  10427.5 47827.5 10492.5 47692.5 ;
      RECT  10427.5 47827.5 10492.5 47692.5 ;
      RECT  10237.5 47827.5 10302.5 47692.5 ;
      RECT  10237.5 48712.5 10302.5 48577.5 ;
      RECT  10427.5 48712.5 10492.5 48577.5 ;
      RECT  10427.5 48712.5 10492.5 48577.5 ;
      RECT  10237.5 48712.5 10302.5 48577.5 ;
      RECT  10597.5 47737.5 10662.5 47602.5 ;
      RECT  10597.5 48712.5 10662.5 48577.5 ;
      RECT  10295.0 48270.0 10360.0 48135.0 ;
      RECT  10295.0 48270.0 10360.0 48135.0 ;
      RECT  10460.0 48235.0 10525.0 48170.0 ;
      RECT  10170.0 47517.5 10730.0 47452.5 ;
      RECT  10170.0 48862.5 10730.0 48797.5 ;
      RECT  8432.5 48135.0 8497.5 48270.0 ;
      RECT  8572.5 48407.5 8637.5 48542.5 ;
      RECT  9567.5 48372.5 9432.5 48437.5 ;
      RECT  9117.5 49990.0 9182.5 50175.0 ;
      RECT  9117.5 48830.0 9182.5 49015.0 ;
      RECT  8757.5 48947.5 8822.5 48797.5 ;
      RECT  8757.5 49832.5 8822.5 50207.5 ;
      RECT  8947.5 48947.5 9012.5 49832.5 ;
      RECT  8757.5 49832.5 8822.5 49967.5 ;
      RECT  8947.5 49832.5 9012.5 49967.5 ;
      RECT  8947.5 49832.5 9012.5 49967.5 ;
      RECT  8757.5 49832.5 8822.5 49967.5 ;
      RECT  8757.5 48947.5 8822.5 49082.5 ;
      RECT  8947.5 48947.5 9012.5 49082.5 ;
      RECT  8947.5 48947.5 9012.5 49082.5 ;
      RECT  8757.5 48947.5 8822.5 49082.5 ;
      RECT  9117.5 49922.5 9182.5 50057.5 ;
      RECT  9117.5 48947.5 9182.5 49082.5 ;
      RECT  8815.0 49390.0 8880.0 49525.0 ;
      RECT  8815.0 49390.0 8880.0 49525.0 ;
      RECT  8980.0 49425.0 9045.0 49490.0 ;
      RECT  8690.0 50142.5 9250.0 50207.5 ;
      RECT  8690.0 48797.5 9250.0 48862.5 ;
      RECT  9317.5 48992.5 9382.5 48797.5 ;
      RECT  9317.5 49832.5 9382.5 50207.5 ;
      RECT  9697.5 49832.5 9762.5 50207.5 ;
      RECT  9867.5 49990.0 9932.5 50175.0 ;
      RECT  9867.5 48830.0 9932.5 49015.0 ;
      RECT  9317.5 49832.5 9382.5 49967.5 ;
      RECT  9507.5 49832.5 9572.5 49967.5 ;
      RECT  9507.5 49832.5 9572.5 49967.5 ;
      RECT  9317.5 49832.5 9382.5 49967.5 ;
      RECT  9507.5 49832.5 9572.5 49967.5 ;
      RECT  9697.5 49832.5 9762.5 49967.5 ;
      RECT  9697.5 49832.5 9762.5 49967.5 ;
      RECT  9507.5 49832.5 9572.5 49967.5 ;
      RECT  9317.5 48992.5 9382.5 49127.5 ;
      RECT  9507.5 48992.5 9572.5 49127.5 ;
      RECT  9507.5 48992.5 9572.5 49127.5 ;
      RECT  9317.5 48992.5 9382.5 49127.5 ;
      RECT  9507.5 48992.5 9572.5 49127.5 ;
      RECT  9697.5 48992.5 9762.5 49127.5 ;
      RECT  9697.5 48992.5 9762.5 49127.5 ;
      RECT  9507.5 48992.5 9572.5 49127.5 ;
      RECT  9867.5 49922.5 9932.5 50057.5 ;
      RECT  9867.5 48947.5 9932.5 49082.5 ;
      RECT  9702.5 49222.5 9567.5 49287.5 ;
      RECT  9445.0 49437.5 9310.0 49502.5 ;
      RECT  9507.5 49832.5 9572.5 49967.5 ;
      RECT  9697.5 48992.5 9762.5 49127.5 ;
      RECT  9797.5 49437.5 9662.5 49502.5 ;
      RECT  9310.0 49437.5 9445.0 49502.5 ;
      RECT  9567.5 49222.5 9702.5 49287.5 ;
      RECT  9662.5 49437.5 9797.5 49502.5 ;
      RECT  9250.0 50142.5 10170.0 50207.5 ;
      RECT  9250.0 48797.5 10170.0 48862.5 ;
      RECT  10597.5 49990.0 10662.5 50175.0 ;
      RECT  10597.5 48830.0 10662.5 49015.0 ;
      RECT  10237.5 48947.5 10302.5 48797.5 ;
      RECT  10237.5 49832.5 10302.5 50207.5 ;
      RECT  10427.5 48947.5 10492.5 49832.5 ;
      RECT  10237.5 49832.5 10302.5 49967.5 ;
      RECT  10427.5 49832.5 10492.5 49967.5 ;
      RECT  10427.5 49832.5 10492.5 49967.5 ;
      RECT  10237.5 49832.5 10302.5 49967.5 ;
      RECT  10237.5 48947.5 10302.5 49082.5 ;
      RECT  10427.5 48947.5 10492.5 49082.5 ;
      RECT  10427.5 48947.5 10492.5 49082.5 ;
      RECT  10237.5 48947.5 10302.5 49082.5 ;
      RECT  10597.5 49922.5 10662.5 50057.5 ;
      RECT  10597.5 48947.5 10662.5 49082.5 ;
      RECT  10295.0 49390.0 10360.0 49525.0 ;
      RECT  10295.0 49390.0 10360.0 49525.0 ;
      RECT  10460.0 49425.0 10525.0 49490.0 ;
      RECT  10170.0 50142.5 10730.0 50207.5 ;
      RECT  10170.0 48797.5 10730.0 48862.5 ;
      RECT  8432.5 49390.0 8497.5 49525.0 ;
      RECT  8572.5 49117.5 8637.5 49252.5 ;
      RECT  9567.5 49222.5 9432.5 49287.5 ;
      RECT  9117.5 50360.0 9182.5 50175.0 ;
      RECT  9117.5 51520.0 9182.5 51335.0 ;
      RECT  8757.5 51402.5 8822.5 51552.5 ;
      RECT  8757.5 50517.5 8822.5 50142.5 ;
      RECT  8947.5 51402.5 9012.5 50517.5 ;
      RECT  8757.5 50517.5 8822.5 50382.5 ;
      RECT  8947.5 50517.5 9012.5 50382.5 ;
      RECT  8947.5 50517.5 9012.5 50382.5 ;
      RECT  8757.5 50517.5 8822.5 50382.5 ;
      RECT  8757.5 51402.5 8822.5 51267.5 ;
      RECT  8947.5 51402.5 9012.5 51267.5 ;
      RECT  8947.5 51402.5 9012.5 51267.5 ;
      RECT  8757.5 51402.5 8822.5 51267.5 ;
      RECT  9117.5 50427.5 9182.5 50292.5 ;
      RECT  9117.5 51402.5 9182.5 51267.5 ;
      RECT  8815.0 50960.0 8880.0 50825.0 ;
      RECT  8815.0 50960.0 8880.0 50825.0 ;
      RECT  8980.0 50925.0 9045.0 50860.0 ;
      RECT  8690.0 50207.5 9250.0 50142.5 ;
      RECT  8690.0 51552.5 9250.0 51487.5 ;
      RECT  9317.5 51357.5 9382.5 51552.5 ;
      RECT  9317.5 50517.5 9382.5 50142.5 ;
      RECT  9697.5 50517.5 9762.5 50142.5 ;
      RECT  9867.5 50360.0 9932.5 50175.0 ;
      RECT  9867.5 51520.0 9932.5 51335.0 ;
      RECT  9317.5 50517.5 9382.5 50382.5 ;
      RECT  9507.5 50517.5 9572.5 50382.5 ;
      RECT  9507.5 50517.5 9572.5 50382.5 ;
      RECT  9317.5 50517.5 9382.5 50382.5 ;
      RECT  9507.5 50517.5 9572.5 50382.5 ;
      RECT  9697.5 50517.5 9762.5 50382.5 ;
      RECT  9697.5 50517.5 9762.5 50382.5 ;
      RECT  9507.5 50517.5 9572.5 50382.5 ;
      RECT  9317.5 51357.5 9382.5 51222.5 ;
      RECT  9507.5 51357.5 9572.5 51222.5 ;
      RECT  9507.5 51357.5 9572.5 51222.5 ;
      RECT  9317.5 51357.5 9382.5 51222.5 ;
      RECT  9507.5 51357.5 9572.5 51222.5 ;
      RECT  9697.5 51357.5 9762.5 51222.5 ;
      RECT  9697.5 51357.5 9762.5 51222.5 ;
      RECT  9507.5 51357.5 9572.5 51222.5 ;
      RECT  9867.5 50427.5 9932.5 50292.5 ;
      RECT  9867.5 51402.5 9932.5 51267.5 ;
      RECT  9702.5 51127.5 9567.5 51062.5 ;
      RECT  9445.0 50912.5 9310.0 50847.5 ;
      RECT  9507.5 50517.5 9572.5 50382.5 ;
      RECT  9697.5 51357.5 9762.5 51222.5 ;
      RECT  9797.5 50912.5 9662.5 50847.5 ;
      RECT  9310.0 50912.5 9445.0 50847.5 ;
      RECT  9567.5 51127.5 9702.5 51062.5 ;
      RECT  9662.5 50912.5 9797.5 50847.5 ;
      RECT  9250.0 50207.5 10170.0 50142.5 ;
      RECT  9250.0 51552.5 10170.0 51487.5 ;
      RECT  10597.5 50360.0 10662.5 50175.0 ;
      RECT  10597.5 51520.0 10662.5 51335.0 ;
      RECT  10237.5 51402.5 10302.5 51552.5 ;
      RECT  10237.5 50517.5 10302.5 50142.5 ;
      RECT  10427.5 51402.5 10492.5 50517.5 ;
      RECT  10237.5 50517.5 10302.5 50382.5 ;
      RECT  10427.5 50517.5 10492.5 50382.5 ;
      RECT  10427.5 50517.5 10492.5 50382.5 ;
      RECT  10237.5 50517.5 10302.5 50382.5 ;
      RECT  10237.5 51402.5 10302.5 51267.5 ;
      RECT  10427.5 51402.5 10492.5 51267.5 ;
      RECT  10427.5 51402.5 10492.5 51267.5 ;
      RECT  10237.5 51402.5 10302.5 51267.5 ;
      RECT  10597.5 50427.5 10662.5 50292.5 ;
      RECT  10597.5 51402.5 10662.5 51267.5 ;
      RECT  10295.0 50960.0 10360.0 50825.0 ;
      RECT  10295.0 50960.0 10360.0 50825.0 ;
      RECT  10460.0 50925.0 10525.0 50860.0 ;
      RECT  10170.0 50207.5 10730.0 50142.5 ;
      RECT  10170.0 51552.5 10730.0 51487.5 ;
      RECT  8432.5 50825.0 8497.5 50960.0 ;
      RECT  8572.5 51097.5 8637.5 51232.5 ;
      RECT  9567.5 51062.5 9432.5 51127.5 ;
      RECT  9117.5 52680.0 9182.5 52865.0 ;
      RECT  9117.5 51520.0 9182.5 51705.0 ;
      RECT  8757.5 51637.5 8822.5 51487.5 ;
      RECT  8757.5 52522.5 8822.5 52897.5 ;
      RECT  8947.5 51637.5 9012.5 52522.5 ;
      RECT  8757.5 52522.5 8822.5 52657.5 ;
      RECT  8947.5 52522.5 9012.5 52657.5 ;
      RECT  8947.5 52522.5 9012.5 52657.5 ;
      RECT  8757.5 52522.5 8822.5 52657.5 ;
      RECT  8757.5 51637.5 8822.5 51772.5 ;
      RECT  8947.5 51637.5 9012.5 51772.5 ;
      RECT  8947.5 51637.5 9012.5 51772.5 ;
      RECT  8757.5 51637.5 8822.5 51772.5 ;
      RECT  9117.5 52612.5 9182.5 52747.5 ;
      RECT  9117.5 51637.5 9182.5 51772.5 ;
      RECT  8815.0 52080.0 8880.0 52215.0 ;
      RECT  8815.0 52080.0 8880.0 52215.0 ;
      RECT  8980.0 52115.0 9045.0 52180.0 ;
      RECT  8690.0 52832.5 9250.0 52897.5 ;
      RECT  8690.0 51487.5 9250.0 51552.5 ;
      RECT  9317.5 51682.5 9382.5 51487.5 ;
      RECT  9317.5 52522.5 9382.5 52897.5 ;
      RECT  9697.5 52522.5 9762.5 52897.5 ;
      RECT  9867.5 52680.0 9932.5 52865.0 ;
      RECT  9867.5 51520.0 9932.5 51705.0 ;
      RECT  9317.5 52522.5 9382.5 52657.5 ;
      RECT  9507.5 52522.5 9572.5 52657.5 ;
      RECT  9507.5 52522.5 9572.5 52657.5 ;
      RECT  9317.5 52522.5 9382.5 52657.5 ;
      RECT  9507.5 52522.5 9572.5 52657.5 ;
      RECT  9697.5 52522.5 9762.5 52657.5 ;
      RECT  9697.5 52522.5 9762.5 52657.5 ;
      RECT  9507.5 52522.5 9572.5 52657.5 ;
      RECT  9317.5 51682.5 9382.5 51817.5 ;
      RECT  9507.5 51682.5 9572.5 51817.5 ;
      RECT  9507.5 51682.5 9572.5 51817.5 ;
      RECT  9317.5 51682.5 9382.5 51817.5 ;
      RECT  9507.5 51682.5 9572.5 51817.5 ;
      RECT  9697.5 51682.5 9762.5 51817.5 ;
      RECT  9697.5 51682.5 9762.5 51817.5 ;
      RECT  9507.5 51682.5 9572.5 51817.5 ;
      RECT  9867.5 52612.5 9932.5 52747.5 ;
      RECT  9867.5 51637.5 9932.5 51772.5 ;
      RECT  9702.5 51912.5 9567.5 51977.5 ;
      RECT  9445.0 52127.5 9310.0 52192.5 ;
      RECT  9507.5 52522.5 9572.5 52657.5 ;
      RECT  9697.5 51682.5 9762.5 51817.5 ;
      RECT  9797.5 52127.5 9662.5 52192.5 ;
      RECT  9310.0 52127.5 9445.0 52192.5 ;
      RECT  9567.5 51912.5 9702.5 51977.5 ;
      RECT  9662.5 52127.5 9797.5 52192.5 ;
      RECT  9250.0 52832.5 10170.0 52897.5 ;
      RECT  9250.0 51487.5 10170.0 51552.5 ;
      RECT  10597.5 52680.0 10662.5 52865.0 ;
      RECT  10597.5 51520.0 10662.5 51705.0 ;
      RECT  10237.5 51637.5 10302.5 51487.5 ;
      RECT  10237.5 52522.5 10302.5 52897.5 ;
      RECT  10427.5 51637.5 10492.5 52522.5 ;
      RECT  10237.5 52522.5 10302.5 52657.5 ;
      RECT  10427.5 52522.5 10492.5 52657.5 ;
      RECT  10427.5 52522.5 10492.5 52657.5 ;
      RECT  10237.5 52522.5 10302.5 52657.5 ;
      RECT  10237.5 51637.5 10302.5 51772.5 ;
      RECT  10427.5 51637.5 10492.5 51772.5 ;
      RECT  10427.5 51637.5 10492.5 51772.5 ;
      RECT  10237.5 51637.5 10302.5 51772.5 ;
      RECT  10597.5 52612.5 10662.5 52747.5 ;
      RECT  10597.5 51637.5 10662.5 51772.5 ;
      RECT  10295.0 52080.0 10360.0 52215.0 ;
      RECT  10295.0 52080.0 10360.0 52215.0 ;
      RECT  10460.0 52115.0 10525.0 52180.0 ;
      RECT  10170.0 52832.5 10730.0 52897.5 ;
      RECT  10170.0 51487.5 10730.0 51552.5 ;
      RECT  8432.5 52080.0 8497.5 52215.0 ;
      RECT  8572.5 51807.5 8637.5 51942.5 ;
      RECT  9567.5 51912.5 9432.5 51977.5 ;
      RECT  9117.5 53050.0 9182.5 52865.0 ;
      RECT  9117.5 54210.0 9182.5 54025.0 ;
      RECT  8757.5 54092.5 8822.5 54242.5 ;
      RECT  8757.5 53207.5 8822.5 52832.5 ;
      RECT  8947.5 54092.5 9012.5 53207.5 ;
      RECT  8757.5 53207.5 8822.5 53072.5 ;
      RECT  8947.5 53207.5 9012.5 53072.5 ;
      RECT  8947.5 53207.5 9012.5 53072.5 ;
      RECT  8757.5 53207.5 8822.5 53072.5 ;
      RECT  8757.5 54092.5 8822.5 53957.5 ;
      RECT  8947.5 54092.5 9012.5 53957.5 ;
      RECT  8947.5 54092.5 9012.5 53957.5 ;
      RECT  8757.5 54092.5 8822.5 53957.5 ;
      RECT  9117.5 53117.5 9182.5 52982.5 ;
      RECT  9117.5 54092.5 9182.5 53957.5 ;
      RECT  8815.0 53650.0 8880.0 53515.0 ;
      RECT  8815.0 53650.0 8880.0 53515.0 ;
      RECT  8980.0 53615.0 9045.0 53550.0 ;
      RECT  8690.0 52897.5 9250.0 52832.5 ;
      RECT  8690.0 54242.5 9250.0 54177.5 ;
      RECT  9317.5 54047.5 9382.5 54242.5 ;
      RECT  9317.5 53207.5 9382.5 52832.5 ;
      RECT  9697.5 53207.5 9762.5 52832.5 ;
      RECT  9867.5 53050.0 9932.5 52865.0 ;
      RECT  9867.5 54210.0 9932.5 54025.0 ;
      RECT  9317.5 53207.5 9382.5 53072.5 ;
      RECT  9507.5 53207.5 9572.5 53072.5 ;
      RECT  9507.5 53207.5 9572.5 53072.5 ;
      RECT  9317.5 53207.5 9382.5 53072.5 ;
      RECT  9507.5 53207.5 9572.5 53072.5 ;
      RECT  9697.5 53207.5 9762.5 53072.5 ;
      RECT  9697.5 53207.5 9762.5 53072.5 ;
      RECT  9507.5 53207.5 9572.5 53072.5 ;
      RECT  9317.5 54047.5 9382.5 53912.5 ;
      RECT  9507.5 54047.5 9572.5 53912.5 ;
      RECT  9507.5 54047.5 9572.5 53912.5 ;
      RECT  9317.5 54047.5 9382.5 53912.5 ;
      RECT  9507.5 54047.5 9572.5 53912.5 ;
      RECT  9697.5 54047.5 9762.5 53912.5 ;
      RECT  9697.5 54047.5 9762.5 53912.5 ;
      RECT  9507.5 54047.5 9572.5 53912.5 ;
      RECT  9867.5 53117.5 9932.5 52982.5 ;
      RECT  9867.5 54092.5 9932.5 53957.5 ;
      RECT  9702.5 53817.5 9567.5 53752.5 ;
      RECT  9445.0 53602.5 9310.0 53537.5 ;
      RECT  9507.5 53207.5 9572.5 53072.5 ;
      RECT  9697.5 54047.5 9762.5 53912.5 ;
      RECT  9797.5 53602.5 9662.5 53537.5 ;
      RECT  9310.0 53602.5 9445.0 53537.5 ;
      RECT  9567.5 53817.5 9702.5 53752.5 ;
      RECT  9662.5 53602.5 9797.5 53537.5 ;
      RECT  9250.0 52897.5 10170.0 52832.5 ;
      RECT  9250.0 54242.5 10170.0 54177.5 ;
      RECT  10597.5 53050.0 10662.5 52865.0 ;
      RECT  10597.5 54210.0 10662.5 54025.0 ;
      RECT  10237.5 54092.5 10302.5 54242.5 ;
      RECT  10237.5 53207.5 10302.5 52832.5 ;
      RECT  10427.5 54092.5 10492.5 53207.5 ;
      RECT  10237.5 53207.5 10302.5 53072.5 ;
      RECT  10427.5 53207.5 10492.5 53072.5 ;
      RECT  10427.5 53207.5 10492.5 53072.5 ;
      RECT  10237.5 53207.5 10302.5 53072.5 ;
      RECT  10237.5 54092.5 10302.5 53957.5 ;
      RECT  10427.5 54092.5 10492.5 53957.5 ;
      RECT  10427.5 54092.5 10492.5 53957.5 ;
      RECT  10237.5 54092.5 10302.5 53957.5 ;
      RECT  10597.5 53117.5 10662.5 52982.5 ;
      RECT  10597.5 54092.5 10662.5 53957.5 ;
      RECT  10295.0 53650.0 10360.0 53515.0 ;
      RECT  10295.0 53650.0 10360.0 53515.0 ;
      RECT  10460.0 53615.0 10525.0 53550.0 ;
      RECT  10170.0 52897.5 10730.0 52832.5 ;
      RECT  10170.0 54242.5 10730.0 54177.5 ;
      RECT  8432.5 53515.0 8497.5 53650.0 ;
      RECT  8572.5 53787.5 8637.5 53922.5 ;
      RECT  9567.5 53752.5 9432.5 53817.5 ;
      RECT  9117.5 55370.0 9182.5 55555.0 ;
      RECT  9117.5 54210.0 9182.5 54395.0 ;
      RECT  8757.5 54327.5 8822.5 54177.5 ;
      RECT  8757.5 55212.5 8822.5 55587.5 ;
      RECT  8947.5 54327.5 9012.5 55212.5 ;
      RECT  8757.5 55212.5 8822.5 55347.5 ;
      RECT  8947.5 55212.5 9012.5 55347.5 ;
      RECT  8947.5 55212.5 9012.5 55347.5 ;
      RECT  8757.5 55212.5 8822.5 55347.5 ;
      RECT  8757.5 54327.5 8822.5 54462.5 ;
      RECT  8947.5 54327.5 9012.5 54462.5 ;
      RECT  8947.5 54327.5 9012.5 54462.5 ;
      RECT  8757.5 54327.5 8822.5 54462.5 ;
      RECT  9117.5 55302.5 9182.5 55437.5 ;
      RECT  9117.5 54327.5 9182.5 54462.5 ;
      RECT  8815.0 54770.0 8880.0 54905.0 ;
      RECT  8815.0 54770.0 8880.0 54905.0 ;
      RECT  8980.0 54805.0 9045.0 54870.0 ;
      RECT  8690.0 55522.5 9250.0 55587.5 ;
      RECT  8690.0 54177.5 9250.0 54242.5 ;
      RECT  9317.5 54372.5 9382.5 54177.5 ;
      RECT  9317.5 55212.5 9382.5 55587.5 ;
      RECT  9697.5 55212.5 9762.5 55587.5 ;
      RECT  9867.5 55370.0 9932.5 55555.0 ;
      RECT  9867.5 54210.0 9932.5 54395.0 ;
      RECT  9317.5 55212.5 9382.5 55347.5 ;
      RECT  9507.5 55212.5 9572.5 55347.5 ;
      RECT  9507.5 55212.5 9572.5 55347.5 ;
      RECT  9317.5 55212.5 9382.5 55347.5 ;
      RECT  9507.5 55212.5 9572.5 55347.5 ;
      RECT  9697.5 55212.5 9762.5 55347.5 ;
      RECT  9697.5 55212.5 9762.5 55347.5 ;
      RECT  9507.5 55212.5 9572.5 55347.5 ;
      RECT  9317.5 54372.5 9382.5 54507.5 ;
      RECT  9507.5 54372.5 9572.5 54507.5 ;
      RECT  9507.5 54372.5 9572.5 54507.5 ;
      RECT  9317.5 54372.5 9382.5 54507.5 ;
      RECT  9507.5 54372.5 9572.5 54507.5 ;
      RECT  9697.5 54372.5 9762.5 54507.5 ;
      RECT  9697.5 54372.5 9762.5 54507.5 ;
      RECT  9507.5 54372.5 9572.5 54507.5 ;
      RECT  9867.5 55302.5 9932.5 55437.5 ;
      RECT  9867.5 54327.5 9932.5 54462.5 ;
      RECT  9702.5 54602.5 9567.5 54667.5 ;
      RECT  9445.0 54817.5 9310.0 54882.5 ;
      RECT  9507.5 55212.5 9572.5 55347.5 ;
      RECT  9697.5 54372.5 9762.5 54507.5 ;
      RECT  9797.5 54817.5 9662.5 54882.5 ;
      RECT  9310.0 54817.5 9445.0 54882.5 ;
      RECT  9567.5 54602.5 9702.5 54667.5 ;
      RECT  9662.5 54817.5 9797.5 54882.5 ;
      RECT  9250.0 55522.5 10170.0 55587.5 ;
      RECT  9250.0 54177.5 10170.0 54242.5 ;
      RECT  10597.5 55370.0 10662.5 55555.0 ;
      RECT  10597.5 54210.0 10662.5 54395.0 ;
      RECT  10237.5 54327.5 10302.5 54177.5 ;
      RECT  10237.5 55212.5 10302.5 55587.5 ;
      RECT  10427.5 54327.5 10492.5 55212.5 ;
      RECT  10237.5 55212.5 10302.5 55347.5 ;
      RECT  10427.5 55212.5 10492.5 55347.5 ;
      RECT  10427.5 55212.5 10492.5 55347.5 ;
      RECT  10237.5 55212.5 10302.5 55347.5 ;
      RECT  10237.5 54327.5 10302.5 54462.5 ;
      RECT  10427.5 54327.5 10492.5 54462.5 ;
      RECT  10427.5 54327.5 10492.5 54462.5 ;
      RECT  10237.5 54327.5 10302.5 54462.5 ;
      RECT  10597.5 55302.5 10662.5 55437.5 ;
      RECT  10597.5 54327.5 10662.5 54462.5 ;
      RECT  10295.0 54770.0 10360.0 54905.0 ;
      RECT  10295.0 54770.0 10360.0 54905.0 ;
      RECT  10460.0 54805.0 10525.0 54870.0 ;
      RECT  10170.0 55522.5 10730.0 55587.5 ;
      RECT  10170.0 54177.5 10730.0 54242.5 ;
      RECT  8432.5 54770.0 8497.5 54905.0 ;
      RECT  8572.5 54497.5 8637.5 54632.5 ;
      RECT  9567.5 54602.5 9432.5 54667.5 ;
      RECT  9117.5 55740.0 9182.5 55555.0 ;
      RECT  9117.5 56900.0 9182.5 56715.0 ;
      RECT  8757.5 56782.5 8822.5 56932.5 ;
      RECT  8757.5 55897.5 8822.5 55522.5 ;
      RECT  8947.5 56782.5 9012.5 55897.5 ;
      RECT  8757.5 55897.5 8822.5 55762.5 ;
      RECT  8947.5 55897.5 9012.5 55762.5 ;
      RECT  8947.5 55897.5 9012.5 55762.5 ;
      RECT  8757.5 55897.5 8822.5 55762.5 ;
      RECT  8757.5 56782.5 8822.5 56647.5 ;
      RECT  8947.5 56782.5 9012.5 56647.5 ;
      RECT  8947.5 56782.5 9012.5 56647.5 ;
      RECT  8757.5 56782.5 8822.5 56647.5 ;
      RECT  9117.5 55807.5 9182.5 55672.5 ;
      RECT  9117.5 56782.5 9182.5 56647.5 ;
      RECT  8815.0 56340.0 8880.0 56205.0 ;
      RECT  8815.0 56340.0 8880.0 56205.0 ;
      RECT  8980.0 56305.0 9045.0 56240.0 ;
      RECT  8690.0 55587.5 9250.0 55522.5 ;
      RECT  8690.0 56932.5 9250.0 56867.5 ;
      RECT  9317.5 56737.5 9382.5 56932.5 ;
      RECT  9317.5 55897.5 9382.5 55522.5 ;
      RECT  9697.5 55897.5 9762.5 55522.5 ;
      RECT  9867.5 55740.0 9932.5 55555.0 ;
      RECT  9867.5 56900.0 9932.5 56715.0 ;
      RECT  9317.5 55897.5 9382.5 55762.5 ;
      RECT  9507.5 55897.5 9572.5 55762.5 ;
      RECT  9507.5 55897.5 9572.5 55762.5 ;
      RECT  9317.5 55897.5 9382.5 55762.5 ;
      RECT  9507.5 55897.5 9572.5 55762.5 ;
      RECT  9697.5 55897.5 9762.5 55762.5 ;
      RECT  9697.5 55897.5 9762.5 55762.5 ;
      RECT  9507.5 55897.5 9572.5 55762.5 ;
      RECT  9317.5 56737.5 9382.5 56602.5 ;
      RECT  9507.5 56737.5 9572.5 56602.5 ;
      RECT  9507.5 56737.5 9572.5 56602.5 ;
      RECT  9317.5 56737.5 9382.5 56602.5 ;
      RECT  9507.5 56737.5 9572.5 56602.5 ;
      RECT  9697.5 56737.5 9762.5 56602.5 ;
      RECT  9697.5 56737.5 9762.5 56602.5 ;
      RECT  9507.5 56737.5 9572.5 56602.5 ;
      RECT  9867.5 55807.5 9932.5 55672.5 ;
      RECT  9867.5 56782.5 9932.5 56647.5 ;
      RECT  9702.5 56507.5 9567.5 56442.5 ;
      RECT  9445.0 56292.5 9310.0 56227.5 ;
      RECT  9507.5 55897.5 9572.5 55762.5 ;
      RECT  9697.5 56737.5 9762.5 56602.5 ;
      RECT  9797.5 56292.5 9662.5 56227.5 ;
      RECT  9310.0 56292.5 9445.0 56227.5 ;
      RECT  9567.5 56507.5 9702.5 56442.5 ;
      RECT  9662.5 56292.5 9797.5 56227.5 ;
      RECT  9250.0 55587.5 10170.0 55522.5 ;
      RECT  9250.0 56932.5 10170.0 56867.5 ;
      RECT  10597.5 55740.0 10662.5 55555.0 ;
      RECT  10597.5 56900.0 10662.5 56715.0 ;
      RECT  10237.5 56782.5 10302.5 56932.5 ;
      RECT  10237.5 55897.5 10302.5 55522.5 ;
      RECT  10427.5 56782.5 10492.5 55897.5 ;
      RECT  10237.5 55897.5 10302.5 55762.5 ;
      RECT  10427.5 55897.5 10492.5 55762.5 ;
      RECT  10427.5 55897.5 10492.5 55762.5 ;
      RECT  10237.5 55897.5 10302.5 55762.5 ;
      RECT  10237.5 56782.5 10302.5 56647.5 ;
      RECT  10427.5 56782.5 10492.5 56647.5 ;
      RECT  10427.5 56782.5 10492.5 56647.5 ;
      RECT  10237.5 56782.5 10302.5 56647.5 ;
      RECT  10597.5 55807.5 10662.5 55672.5 ;
      RECT  10597.5 56782.5 10662.5 56647.5 ;
      RECT  10295.0 56340.0 10360.0 56205.0 ;
      RECT  10295.0 56340.0 10360.0 56205.0 ;
      RECT  10460.0 56305.0 10525.0 56240.0 ;
      RECT  10170.0 55587.5 10730.0 55522.5 ;
      RECT  10170.0 56932.5 10730.0 56867.5 ;
      RECT  8432.5 56205.0 8497.5 56340.0 ;
      RECT  8572.5 56477.5 8637.5 56612.5 ;
      RECT  9567.5 56442.5 9432.5 56507.5 ;
      RECT  9117.5 58060.0 9182.5 58245.0 ;
      RECT  9117.5 56900.0 9182.5 57085.0 ;
      RECT  8757.5 57017.5 8822.5 56867.5 ;
      RECT  8757.5 57902.5 8822.5 58277.5 ;
      RECT  8947.5 57017.5 9012.5 57902.5 ;
      RECT  8757.5 57902.5 8822.5 58037.5 ;
      RECT  8947.5 57902.5 9012.5 58037.5 ;
      RECT  8947.5 57902.5 9012.5 58037.5 ;
      RECT  8757.5 57902.5 8822.5 58037.5 ;
      RECT  8757.5 57017.5 8822.5 57152.5 ;
      RECT  8947.5 57017.5 9012.5 57152.5 ;
      RECT  8947.5 57017.5 9012.5 57152.5 ;
      RECT  8757.5 57017.5 8822.5 57152.5 ;
      RECT  9117.5 57992.5 9182.5 58127.5 ;
      RECT  9117.5 57017.5 9182.5 57152.5 ;
      RECT  8815.0 57460.0 8880.0 57595.0 ;
      RECT  8815.0 57460.0 8880.0 57595.0 ;
      RECT  8980.0 57495.0 9045.0 57560.0 ;
      RECT  8690.0 58212.5 9250.0 58277.5 ;
      RECT  8690.0 56867.5 9250.0 56932.5 ;
      RECT  9317.5 57062.5 9382.5 56867.5 ;
      RECT  9317.5 57902.5 9382.5 58277.5 ;
      RECT  9697.5 57902.5 9762.5 58277.5 ;
      RECT  9867.5 58060.0 9932.5 58245.0 ;
      RECT  9867.5 56900.0 9932.5 57085.0 ;
      RECT  9317.5 57902.5 9382.5 58037.5 ;
      RECT  9507.5 57902.5 9572.5 58037.5 ;
      RECT  9507.5 57902.5 9572.5 58037.5 ;
      RECT  9317.5 57902.5 9382.5 58037.5 ;
      RECT  9507.5 57902.5 9572.5 58037.5 ;
      RECT  9697.5 57902.5 9762.5 58037.5 ;
      RECT  9697.5 57902.5 9762.5 58037.5 ;
      RECT  9507.5 57902.5 9572.5 58037.5 ;
      RECT  9317.5 57062.5 9382.5 57197.5 ;
      RECT  9507.5 57062.5 9572.5 57197.5 ;
      RECT  9507.5 57062.5 9572.5 57197.5 ;
      RECT  9317.5 57062.5 9382.5 57197.5 ;
      RECT  9507.5 57062.5 9572.5 57197.5 ;
      RECT  9697.5 57062.5 9762.5 57197.5 ;
      RECT  9697.5 57062.5 9762.5 57197.5 ;
      RECT  9507.5 57062.5 9572.5 57197.5 ;
      RECT  9867.5 57992.5 9932.5 58127.5 ;
      RECT  9867.5 57017.5 9932.5 57152.5 ;
      RECT  9702.5 57292.5 9567.5 57357.5 ;
      RECT  9445.0 57507.5 9310.0 57572.5 ;
      RECT  9507.5 57902.5 9572.5 58037.5 ;
      RECT  9697.5 57062.5 9762.5 57197.5 ;
      RECT  9797.5 57507.5 9662.5 57572.5 ;
      RECT  9310.0 57507.5 9445.0 57572.5 ;
      RECT  9567.5 57292.5 9702.5 57357.5 ;
      RECT  9662.5 57507.5 9797.5 57572.5 ;
      RECT  9250.0 58212.5 10170.0 58277.5 ;
      RECT  9250.0 56867.5 10170.0 56932.5 ;
      RECT  10597.5 58060.0 10662.5 58245.0 ;
      RECT  10597.5 56900.0 10662.5 57085.0 ;
      RECT  10237.5 57017.5 10302.5 56867.5 ;
      RECT  10237.5 57902.5 10302.5 58277.5 ;
      RECT  10427.5 57017.5 10492.5 57902.5 ;
      RECT  10237.5 57902.5 10302.5 58037.5 ;
      RECT  10427.5 57902.5 10492.5 58037.5 ;
      RECT  10427.5 57902.5 10492.5 58037.5 ;
      RECT  10237.5 57902.5 10302.5 58037.5 ;
      RECT  10237.5 57017.5 10302.5 57152.5 ;
      RECT  10427.5 57017.5 10492.5 57152.5 ;
      RECT  10427.5 57017.5 10492.5 57152.5 ;
      RECT  10237.5 57017.5 10302.5 57152.5 ;
      RECT  10597.5 57992.5 10662.5 58127.5 ;
      RECT  10597.5 57017.5 10662.5 57152.5 ;
      RECT  10295.0 57460.0 10360.0 57595.0 ;
      RECT  10295.0 57460.0 10360.0 57595.0 ;
      RECT  10460.0 57495.0 10525.0 57560.0 ;
      RECT  10170.0 58212.5 10730.0 58277.5 ;
      RECT  10170.0 56867.5 10730.0 56932.5 ;
      RECT  8432.5 57460.0 8497.5 57595.0 ;
      RECT  8572.5 57187.5 8637.5 57322.5 ;
      RECT  9567.5 57292.5 9432.5 57357.5 ;
      RECT  9117.5 58430.0 9182.5 58245.0 ;
      RECT  9117.5 59590.0 9182.5 59405.0 ;
      RECT  8757.5 59472.5 8822.5 59622.5 ;
      RECT  8757.5 58587.5 8822.5 58212.5 ;
      RECT  8947.5 59472.5 9012.5 58587.5 ;
      RECT  8757.5 58587.5 8822.5 58452.5 ;
      RECT  8947.5 58587.5 9012.5 58452.5 ;
      RECT  8947.5 58587.5 9012.5 58452.5 ;
      RECT  8757.5 58587.5 8822.5 58452.5 ;
      RECT  8757.5 59472.5 8822.5 59337.5 ;
      RECT  8947.5 59472.5 9012.5 59337.5 ;
      RECT  8947.5 59472.5 9012.5 59337.5 ;
      RECT  8757.5 59472.5 8822.5 59337.5 ;
      RECT  9117.5 58497.5 9182.5 58362.5 ;
      RECT  9117.5 59472.5 9182.5 59337.5 ;
      RECT  8815.0 59030.0 8880.0 58895.0 ;
      RECT  8815.0 59030.0 8880.0 58895.0 ;
      RECT  8980.0 58995.0 9045.0 58930.0 ;
      RECT  8690.0 58277.5 9250.0 58212.5 ;
      RECT  8690.0 59622.5 9250.0 59557.5 ;
      RECT  9317.5 59427.5 9382.5 59622.5 ;
      RECT  9317.5 58587.5 9382.5 58212.5 ;
      RECT  9697.5 58587.5 9762.5 58212.5 ;
      RECT  9867.5 58430.0 9932.5 58245.0 ;
      RECT  9867.5 59590.0 9932.5 59405.0 ;
      RECT  9317.5 58587.5 9382.5 58452.5 ;
      RECT  9507.5 58587.5 9572.5 58452.5 ;
      RECT  9507.5 58587.5 9572.5 58452.5 ;
      RECT  9317.5 58587.5 9382.5 58452.5 ;
      RECT  9507.5 58587.5 9572.5 58452.5 ;
      RECT  9697.5 58587.5 9762.5 58452.5 ;
      RECT  9697.5 58587.5 9762.5 58452.5 ;
      RECT  9507.5 58587.5 9572.5 58452.5 ;
      RECT  9317.5 59427.5 9382.5 59292.5 ;
      RECT  9507.5 59427.5 9572.5 59292.5 ;
      RECT  9507.5 59427.5 9572.5 59292.5 ;
      RECT  9317.5 59427.5 9382.5 59292.5 ;
      RECT  9507.5 59427.5 9572.5 59292.5 ;
      RECT  9697.5 59427.5 9762.5 59292.5 ;
      RECT  9697.5 59427.5 9762.5 59292.5 ;
      RECT  9507.5 59427.5 9572.5 59292.5 ;
      RECT  9867.5 58497.5 9932.5 58362.5 ;
      RECT  9867.5 59472.5 9932.5 59337.5 ;
      RECT  9702.5 59197.5 9567.5 59132.5 ;
      RECT  9445.0 58982.5 9310.0 58917.5 ;
      RECT  9507.5 58587.5 9572.5 58452.5 ;
      RECT  9697.5 59427.5 9762.5 59292.5 ;
      RECT  9797.5 58982.5 9662.5 58917.5 ;
      RECT  9310.0 58982.5 9445.0 58917.5 ;
      RECT  9567.5 59197.5 9702.5 59132.5 ;
      RECT  9662.5 58982.5 9797.5 58917.5 ;
      RECT  9250.0 58277.5 10170.0 58212.5 ;
      RECT  9250.0 59622.5 10170.0 59557.5 ;
      RECT  10597.5 58430.0 10662.5 58245.0 ;
      RECT  10597.5 59590.0 10662.5 59405.0 ;
      RECT  10237.5 59472.5 10302.5 59622.5 ;
      RECT  10237.5 58587.5 10302.5 58212.5 ;
      RECT  10427.5 59472.5 10492.5 58587.5 ;
      RECT  10237.5 58587.5 10302.5 58452.5 ;
      RECT  10427.5 58587.5 10492.5 58452.5 ;
      RECT  10427.5 58587.5 10492.5 58452.5 ;
      RECT  10237.5 58587.5 10302.5 58452.5 ;
      RECT  10237.5 59472.5 10302.5 59337.5 ;
      RECT  10427.5 59472.5 10492.5 59337.5 ;
      RECT  10427.5 59472.5 10492.5 59337.5 ;
      RECT  10237.5 59472.5 10302.5 59337.5 ;
      RECT  10597.5 58497.5 10662.5 58362.5 ;
      RECT  10597.5 59472.5 10662.5 59337.5 ;
      RECT  10295.0 59030.0 10360.0 58895.0 ;
      RECT  10295.0 59030.0 10360.0 58895.0 ;
      RECT  10460.0 58995.0 10525.0 58930.0 ;
      RECT  10170.0 58277.5 10730.0 58212.5 ;
      RECT  10170.0 59622.5 10730.0 59557.5 ;
      RECT  8432.5 58895.0 8497.5 59030.0 ;
      RECT  8572.5 59167.5 8637.5 59302.5 ;
      RECT  9567.5 59132.5 9432.5 59197.5 ;
      RECT  9117.5 60750.0 9182.5 60935.0 ;
      RECT  9117.5 59590.0 9182.5 59775.0 ;
      RECT  8757.5 59707.5 8822.5 59557.5 ;
      RECT  8757.5 60592.5 8822.5 60967.5 ;
      RECT  8947.5 59707.5 9012.5 60592.5 ;
      RECT  8757.5 60592.5 8822.5 60727.5 ;
      RECT  8947.5 60592.5 9012.5 60727.5 ;
      RECT  8947.5 60592.5 9012.5 60727.5 ;
      RECT  8757.5 60592.5 8822.5 60727.5 ;
      RECT  8757.5 59707.5 8822.5 59842.5 ;
      RECT  8947.5 59707.5 9012.5 59842.5 ;
      RECT  8947.5 59707.5 9012.5 59842.5 ;
      RECT  8757.5 59707.5 8822.5 59842.5 ;
      RECT  9117.5 60682.5 9182.5 60817.5 ;
      RECT  9117.5 59707.5 9182.5 59842.5 ;
      RECT  8815.0 60150.0 8880.0 60285.0 ;
      RECT  8815.0 60150.0 8880.0 60285.0 ;
      RECT  8980.0 60185.0 9045.0 60250.0 ;
      RECT  8690.0 60902.5 9250.0 60967.5 ;
      RECT  8690.0 59557.5 9250.0 59622.5 ;
      RECT  9317.5 59752.5 9382.5 59557.5 ;
      RECT  9317.5 60592.5 9382.5 60967.5 ;
      RECT  9697.5 60592.5 9762.5 60967.5 ;
      RECT  9867.5 60750.0 9932.5 60935.0 ;
      RECT  9867.5 59590.0 9932.5 59775.0 ;
      RECT  9317.5 60592.5 9382.5 60727.5 ;
      RECT  9507.5 60592.5 9572.5 60727.5 ;
      RECT  9507.5 60592.5 9572.5 60727.5 ;
      RECT  9317.5 60592.5 9382.5 60727.5 ;
      RECT  9507.5 60592.5 9572.5 60727.5 ;
      RECT  9697.5 60592.5 9762.5 60727.5 ;
      RECT  9697.5 60592.5 9762.5 60727.5 ;
      RECT  9507.5 60592.5 9572.5 60727.5 ;
      RECT  9317.5 59752.5 9382.5 59887.5 ;
      RECT  9507.5 59752.5 9572.5 59887.5 ;
      RECT  9507.5 59752.5 9572.5 59887.5 ;
      RECT  9317.5 59752.5 9382.5 59887.5 ;
      RECT  9507.5 59752.5 9572.5 59887.5 ;
      RECT  9697.5 59752.5 9762.5 59887.5 ;
      RECT  9697.5 59752.5 9762.5 59887.5 ;
      RECT  9507.5 59752.5 9572.5 59887.5 ;
      RECT  9867.5 60682.5 9932.5 60817.5 ;
      RECT  9867.5 59707.5 9932.5 59842.5 ;
      RECT  9702.5 59982.5 9567.5 60047.5 ;
      RECT  9445.0 60197.5 9310.0 60262.5 ;
      RECT  9507.5 60592.5 9572.5 60727.5 ;
      RECT  9697.5 59752.5 9762.5 59887.5 ;
      RECT  9797.5 60197.5 9662.5 60262.5 ;
      RECT  9310.0 60197.5 9445.0 60262.5 ;
      RECT  9567.5 59982.5 9702.5 60047.5 ;
      RECT  9662.5 60197.5 9797.5 60262.5 ;
      RECT  9250.0 60902.5 10170.0 60967.5 ;
      RECT  9250.0 59557.5 10170.0 59622.5 ;
      RECT  10597.5 60750.0 10662.5 60935.0 ;
      RECT  10597.5 59590.0 10662.5 59775.0 ;
      RECT  10237.5 59707.5 10302.5 59557.5 ;
      RECT  10237.5 60592.5 10302.5 60967.5 ;
      RECT  10427.5 59707.5 10492.5 60592.5 ;
      RECT  10237.5 60592.5 10302.5 60727.5 ;
      RECT  10427.5 60592.5 10492.5 60727.5 ;
      RECT  10427.5 60592.5 10492.5 60727.5 ;
      RECT  10237.5 60592.5 10302.5 60727.5 ;
      RECT  10237.5 59707.5 10302.5 59842.5 ;
      RECT  10427.5 59707.5 10492.5 59842.5 ;
      RECT  10427.5 59707.5 10492.5 59842.5 ;
      RECT  10237.5 59707.5 10302.5 59842.5 ;
      RECT  10597.5 60682.5 10662.5 60817.5 ;
      RECT  10597.5 59707.5 10662.5 59842.5 ;
      RECT  10295.0 60150.0 10360.0 60285.0 ;
      RECT  10295.0 60150.0 10360.0 60285.0 ;
      RECT  10460.0 60185.0 10525.0 60250.0 ;
      RECT  10170.0 60902.5 10730.0 60967.5 ;
      RECT  10170.0 59557.5 10730.0 59622.5 ;
      RECT  8432.5 60150.0 8497.5 60285.0 ;
      RECT  8572.5 59877.5 8637.5 60012.5 ;
      RECT  9567.5 59982.5 9432.5 60047.5 ;
      RECT  9117.5 61120.0 9182.5 60935.0 ;
      RECT  9117.5 62280.0 9182.5 62095.0 ;
      RECT  8757.5 62162.5 8822.5 62312.5 ;
      RECT  8757.5 61277.5 8822.5 60902.5 ;
      RECT  8947.5 62162.5 9012.5 61277.5 ;
      RECT  8757.5 61277.5 8822.5 61142.5 ;
      RECT  8947.5 61277.5 9012.5 61142.5 ;
      RECT  8947.5 61277.5 9012.5 61142.5 ;
      RECT  8757.5 61277.5 8822.5 61142.5 ;
      RECT  8757.5 62162.5 8822.5 62027.5 ;
      RECT  8947.5 62162.5 9012.5 62027.5 ;
      RECT  8947.5 62162.5 9012.5 62027.5 ;
      RECT  8757.5 62162.5 8822.5 62027.5 ;
      RECT  9117.5 61187.5 9182.5 61052.5 ;
      RECT  9117.5 62162.5 9182.5 62027.5 ;
      RECT  8815.0 61720.0 8880.0 61585.0 ;
      RECT  8815.0 61720.0 8880.0 61585.0 ;
      RECT  8980.0 61685.0 9045.0 61620.0 ;
      RECT  8690.0 60967.5 9250.0 60902.5 ;
      RECT  8690.0 62312.5 9250.0 62247.5 ;
      RECT  9317.5 62117.5 9382.5 62312.5 ;
      RECT  9317.5 61277.5 9382.5 60902.5 ;
      RECT  9697.5 61277.5 9762.5 60902.5 ;
      RECT  9867.5 61120.0 9932.5 60935.0 ;
      RECT  9867.5 62280.0 9932.5 62095.0 ;
      RECT  9317.5 61277.5 9382.5 61142.5 ;
      RECT  9507.5 61277.5 9572.5 61142.5 ;
      RECT  9507.5 61277.5 9572.5 61142.5 ;
      RECT  9317.5 61277.5 9382.5 61142.5 ;
      RECT  9507.5 61277.5 9572.5 61142.5 ;
      RECT  9697.5 61277.5 9762.5 61142.5 ;
      RECT  9697.5 61277.5 9762.5 61142.5 ;
      RECT  9507.5 61277.5 9572.5 61142.5 ;
      RECT  9317.5 62117.5 9382.5 61982.5 ;
      RECT  9507.5 62117.5 9572.5 61982.5 ;
      RECT  9507.5 62117.5 9572.5 61982.5 ;
      RECT  9317.5 62117.5 9382.5 61982.5 ;
      RECT  9507.5 62117.5 9572.5 61982.5 ;
      RECT  9697.5 62117.5 9762.5 61982.5 ;
      RECT  9697.5 62117.5 9762.5 61982.5 ;
      RECT  9507.5 62117.5 9572.5 61982.5 ;
      RECT  9867.5 61187.5 9932.5 61052.5 ;
      RECT  9867.5 62162.5 9932.5 62027.5 ;
      RECT  9702.5 61887.5 9567.5 61822.5 ;
      RECT  9445.0 61672.5 9310.0 61607.5 ;
      RECT  9507.5 61277.5 9572.5 61142.5 ;
      RECT  9697.5 62117.5 9762.5 61982.5 ;
      RECT  9797.5 61672.5 9662.5 61607.5 ;
      RECT  9310.0 61672.5 9445.0 61607.5 ;
      RECT  9567.5 61887.5 9702.5 61822.5 ;
      RECT  9662.5 61672.5 9797.5 61607.5 ;
      RECT  9250.0 60967.5 10170.0 60902.5 ;
      RECT  9250.0 62312.5 10170.0 62247.5 ;
      RECT  10597.5 61120.0 10662.5 60935.0 ;
      RECT  10597.5 62280.0 10662.5 62095.0 ;
      RECT  10237.5 62162.5 10302.5 62312.5 ;
      RECT  10237.5 61277.5 10302.5 60902.5 ;
      RECT  10427.5 62162.5 10492.5 61277.5 ;
      RECT  10237.5 61277.5 10302.5 61142.5 ;
      RECT  10427.5 61277.5 10492.5 61142.5 ;
      RECT  10427.5 61277.5 10492.5 61142.5 ;
      RECT  10237.5 61277.5 10302.5 61142.5 ;
      RECT  10237.5 62162.5 10302.5 62027.5 ;
      RECT  10427.5 62162.5 10492.5 62027.5 ;
      RECT  10427.5 62162.5 10492.5 62027.5 ;
      RECT  10237.5 62162.5 10302.5 62027.5 ;
      RECT  10597.5 61187.5 10662.5 61052.5 ;
      RECT  10597.5 62162.5 10662.5 62027.5 ;
      RECT  10295.0 61720.0 10360.0 61585.0 ;
      RECT  10295.0 61720.0 10360.0 61585.0 ;
      RECT  10460.0 61685.0 10525.0 61620.0 ;
      RECT  10170.0 60967.5 10730.0 60902.5 ;
      RECT  10170.0 62312.5 10730.0 62247.5 ;
      RECT  8432.5 61585.0 8497.5 61720.0 ;
      RECT  8572.5 61857.5 8637.5 61992.5 ;
      RECT  9567.5 61822.5 9432.5 61887.5 ;
      RECT  9117.5 63440.0 9182.5 63625.0 ;
      RECT  9117.5 62280.0 9182.5 62465.0 ;
      RECT  8757.5 62397.5 8822.5 62247.5 ;
      RECT  8757.5 63282.5 8822.5 63657.5 ;
      RECT  8947.5 62397.5 9012.5 63282.5 ;
      RECT  8757.5 63282.5 8822.5 63417.5 ;
      RECT  8947.5 63282.5 9012.5 63417.5 ;
      RECT  8947.5 63282.5 9012.5 63417.5 ;
      RECT  8757.5 63282.5 8822.5 63417.5 ;
      RECT  8757.5 62397.5 8822.5 62532.5 ;
      RECT  8947.5 62397.5 9012.5 62532.5 ;
      RECT  8947.5 62397.5 9012.5 62532.5 ;
      RECT  8757.5 62397.5 8822.5 62532.5 ;
      RECT  9117.5 63372.5 9182.5 63507.5 ;
      RECT  9117.5 62397.5 9182.5 62532.5 ;
      RECT  8815.0 62840.0 8880.0 62975.0 ;
      RECT  8815.0 62840.0 8880.0 62975.0 ;
      RECT  8980.0 62875.0 9045.0 62940.0 ;
      RECT  8690.0 63592.5 9250.0 63657.5 ;
      RECT  8690.0 62247.5 9250.0 62312.5 ;
      RECT  9317.5 62442.5 9382.5 62247.5 ;
      RECT  9317.5 63282.5 9382.5 63657.5 ;
      RECT  9697.5 63282.5 9762.5 63657.5 ;
      RECT  9867.5 63440.0 9932.5 63625.0 ;
      RECT  9867.5 62280.0 9932.5 62465.0 ;
      RECT  9317.5 63282.5 9382.5 63417.5 ;
      RECT  9507.5 63282.5 9572.5 63417.5 ;
      RECT  9507.5 63282.5 9572.5 63417.5 ;
      RECT  9317.5 63282.5 9382.5 63417.5 ;
      RECT  9507.5 63282.5 9572.5 63417.5 ;
      RECT  9697.5 63282.5 9762.5 63417.5 ;
      RECT  9697.5 63282.5 9762.5 63417.5 ;
      RECT  9507.5 63282.5 9572.5 63417.5 ;
      RECT  9317.5 62442.5 9382.5 62577.5 ;
      RECT  9507.5 62442.5 9572.5 62577.5 ;
      RECT  9507.5 62442.5 9572.5 62577.5 ;
      RECT  9317.5 62442.5 9382.5 62577.5 ;
      RECT  9507.5 62442.5 9572.5 62577.5 ;
      RECT  9697.5 62442.5 9762.5 62577.5 ;
      RECT  9697.5 62442.5 9762.5 62577.5 ;
      RECT  9507.5 62442.5 9572.5 62577.5 ;
      RECT  9867.5 63372.5 9932.5 63507.5 ;
      RECT  9867.5 62397.5 9932.5 62532.5 ;
      RECT  9702.5 62672.5 9567.5 62737.5 ;
      RECT  9445.0 62887.5 9310.0 62952.5 ;
      RECT  9507.5 63282.5 9572.5 63417.5 ;
      RECT  9697.5 62442.5 9762.5 62577.5 ;
      RECT  9797.5 62887.5 9662.5 62952.5 ;
      RECT  9310.0 62887.5 9445.0 62952.5 ;
      RECT  9567.5 62672.5 9702.5 62737.5 ;
      RECT  9662.5 62887.5 9797.5 62952.5 ;
      RECT  9250.0 63592.5 10170.0 63657.5 ;
      RECT  9250.0 62247.5 10170.0 62312.5 ;
      RECT  10597.5 63440.0 10662.5 63625.0 ;
      RECT  10597.5 62280.0 10662.5 62465.0 ;
      RECT  10237.5 62397.5 10302.5 62247.5 ;
      RECT  10237.5 63282.5 10302.5 63657.5 ;
      RECT  10427.5 62397.5 10492.5 63282.5 ;
      RECT  10237.5 63282.5 10302.5 63417.5 ;
      RECT  10427.5 63282.5 10492.5 63417.5 ;
      RECT  10427.5 63282.5 10492.5 63417.5 ;
      RECT  10237.5 63282.5 10302.5 63417.5 ;
      RECT  10237.5 62397.5 10302.5 62532.5 ;
      RECT  10427.5 62397.5 10492.5 62532.5 ;
      RECT  10427.5 62397.5 10492.5 62532.5 ;
      RECT  10237.5 62397.5 10302.5 62532.5 ;
      RECT  10597.5 63372.5 10662.5 63507.5 ;
      RECT  10597.5 62397.5 10662.5 62532.5 ;
      RECT  10295.0 62840.0 10360.0 62975.0 ;
      RECT  10295.0 62840.0 10360.0 62975.0 ;
      RECT  10460.0 62875.0 10525.0 62940.0 ;
      RECT  10170.0 63592.5 10730.0 63657.5 ;
      RECT  10170.0 62247.5 10730.0 62312.5 ;
      RECT  8432.5 62840.0 8497.5 62975.0 ;
      RECT  8572.5 62567.5 8637.5 62702.5 ;
      RECT  9567.5 62672.5 9432.5 62737.5 ;
      RECT  9117.5 63810.0 9182.5 63625.0 ;
      RECT  9117.5 64970.0 9182.5 64785.0 ;
      RECT  8757.5 64852.5 8822.5 65002.5 ;
      RECT  8757.5 63967.5 8822.5 63592.5 ;
      RECT  8947.5 64852.5 9012.5 63967.5 ;
      RECT  8757.5 63967.5 8822.5 63832.5 ;
      RECT  8947.5 63967.5 9012.5 63832.5 ;
      RECT  8947.5 63967.5 9012.5 63832.5 ;
      RECT  8757.5 63967.5 8822.5 63832.5 ;
      RECT  8757.5 64852.5 8822.5 64717.5 ;
      RECT  8947.5 64852.5 9012.5 64717.5 ;
      RECT  8947.5 64852.5 9012.5 64717.5 ;
      RECT  8757.5 64852.5 8822.5 64717.5 ;
      RECT  9117.5 63877.5 9182.5 63742.5 ;
      RECT  9117.5 64852.5 9182.5 64717.5 ;
      RECT  8815.0 64410.0 8880.0 64275.0 ;
      RECT  8815.0 64410.0 8880.0 64275.0 ;
      RECT  8980.0 64375.0 9045.0 64310.0 ;
      RECT  8690.0 63657.5 9250.0 63592.5 ;
      RECT  8690.0 65002.5 9250.0 64937.5 ;
      RECT  9317.5 64807.5 9382.5 65002.5 ;
      RECT  9317.5 63967.5 9382.5 63592.5 ;
      RECT  9697.5 63967.5 9762.5 63592.5 ;
      RECT  9867.5 63810.0 9932.5 63625.0 ;
      RECT  9867.5 64970.0 9932.5 64785.0 ;
      RECT  9317.5 63967.5 9382.5 63832.5 ;
      RECT  9507.5 63967.5 9572.5 63832.5 ;
      RECT  9507.5 63967.5 9572.5 63832.5 ;
      RECT  9317.5 63967.5 9382.5 63832.5 ;
      RECT  9507.5 63967.5 9572.5 63832.5 ;
      RECT  9697.5 63967.5 9762.5 63832.5 ;
      RECT  9697.5 63967.5 9762.5 63832.5 ;
      RECT  9507.5 63967.5 9572.5 63832.5 ;
      RECT  9317.5 64807.5 9382.5 64672.5 ;
      RECT  9507.5 64807.5 9572.5 64672.5 ;
      RECT  9507.5 64807.5 9572.5 64672.5 ;
      RECT  9317.5 64807.5 9382.5 64672.5 ;
      RECT  9507.5 64807.5 9572.5 64672.5 ;
      RECT  9697.5 64807.5 9762.5 64672.5 ;
      RECT  9697.5 64807.5 9762.5 64672.5 ;
      RECT  9507.5 64807.5 9572.5 64672.5 ;
      RECT  9867.5 63877.5 9932.5 63742.5 ;
      RECT  9867.5 64852.5 9932.5 64717.5 ;
      RECT  9702.5 64577.5 9567.5 64512.5 ;
      RECT  9445.0 64362.5 9310.0 64297.5 ;
      RECT  9507.5 63967.5 9572.5 63832.5 ;
      RECT  9697.5 64807.5 9762.5 64672.5 ;
      RECT  9797.5 64362.5 9662.5 64297.5 ;
      RECT  9310.0 64362.5 9445.0 64297.5 ;
      RECT  9567.5 64577.5 9702.5 64512.5 ;
      RECT  9662.5 64362.5 9797.5 64297.5 ;
      RECT  9250.0 63657.5 10170.0 63592.5 ;
      RECT  9250.0 65002.5 10170.0 64937.5 ;
      RECT  10597.5 63810.0 10662.5 63625.0 ;
      RECT  10597.5 64970.0 10662.5 64785.0 ;
      RECT  10237.5 64852.5 10302.5 65002.5 ;
      RECT  10237.5 63967.5 10302.5 63592.5 ;
      RECT  10427.5 64852.5 10492.5 63967.5 ;
      RECT  10237.5 63967.5 10302.5 63832.5 ;
      RECT  10427.5 63967.5 10492.5 63832.5 ;
      RECT  10427.5 63967.5 10492.5 63832.5 ;
      RECT  10237.5 63967.5 10302.5 63832.5 ;
      RECT  10237.5 64852.5 10302.5 64717.5 ;
      RECT  10427.5 64852.5 10492.5 64717.5 ;
      RECT  10427.5 64852.5 10492.5 64717.5 ;
      RECT  10237.5 64852.5 10302.5 64717.5 ;
      RECT  10597.5 63877.5 10662.5 63742.5 ;
      RECT  10597.5 64852.5 10662.5 64717.5 ;
      RECT  10295.0 64410.0 10360.0 64275.0 ;
      RECT  10295.0 64410.0 10360.0 64275.0 ;
      RECT  10460.0 64375.0 10525.0 64310.0 ;
      RECT  10170.0 63657.5 10730.0 63592.5 ;
      RECT  10170.0 65002.5 10730.0 64937.5 ;
      RECT  8432.5 64275.0 8497.5 64410.0 ;
      RECT  8572.5 64547.5 8637.5 64682.5 ;
      RECT  9567.5 64512.5 9432.5 64577.5 ;
      RECT  9117.5 66130.0 9182.5 66315.0 ;
      RECT  9117.5 64970.0 9182.5 65155.0 ;
      RECT  8757.5 65087.5 8822.5 64937.5 ;
      RECT  8757.5 65972.5 8822.5 66347.5 ;
      RECT  8947.5 65087.5 9012.5 65972.5 ;
      RECT  8757.5 65972.5 8822.5 66107.5 ;
      RECT  8947.5 65972.5 9012.5 66107.5 ;
      RECT  8947.5 65972.5 9012.5 66107.5 ;
      RECT  8757.5 65972.5 8822.5 66107.5 ;
      RECT  8757.5 65087.5 8822.5 65222.5 ;
      RECT  8947.5 65087.5 9012.5 65222.5 ;
      RECT  8947.5 65087.5 9012.5 65222.5 ;
      RECT  8757.5 65087.5 8822.5 65222.5 ;
      RECT  9117.5 66062.5 9182.5 66197.5 ;
      RECT  9117.5 65087.5 9182.5 65222.5 ;
      RECT  8815.0 65530.0 8880.0 65665.0 ;
      RECT  8815.0 65530.0 8880.0 65665.0 ;
      RECT  8980.0 65565.0 9045.0 65630.0 ;
      RECT  8690.0 66282.5 9250.0 66347.5 ;
      RECT  8690.0 64937.5 9250.0 65002.5 ;
      RECT  9317.5 65132.5 9382.5 64937.5 ;
      RECT  9317.5 65972.5 9382.5 66347.5 ;
      RECT  9697.5 65972.5 9762.5 66347.5 ;
      RECT  9867.5 66130.0 9932.5 66315.0 ;
      RECT  9867.5 64970.0 9932.5 65155.0 ;
      RECT  9317.5 65972.5 9382.5 66107.5 ;
      RECT  9507.5 65972.5 9572.5 66107.5 ;
      RECT  9507.5 65972.5 9572.5 66107.5 ;
      RECT  9317.5 65972.5 9382.5 66107.5 ;
      RECT  9507.5 65972.5 9572.5 66107.5 ;
      RECT  9697.5 65972.5 9762.5 66107.5 ;
      RECT  9697.5 65972.5 9762.5 66107.5 ;
      RECT  9507.5 65972.5 9572.5 66107.5 ;
      RECT  9317.5 65132.5 9382.5 65267.5 ;
      RECT  9507.5 65132.5 9572.5 65267.5 ;
      RECT  9507.5 65132.5 9572.5 65267.5 ;
      RECT  9317.5 65132.5 9382.5 65267.5 ;
      RECT  9507.5 65132.5 9572.5 65267.5 ;
      RECT  9697.5 65132.5 9762.5 65267.5 ;
      RECT  9697.5 65132.5 9762.5 65267.5 ;
      RECT  9507.5 65132.5 9572.5 65267.5 ;
      RECT  9867.5 66062.5 9932.5 66197.5 ;
      RECT  9867.5 65087.5 9932.5 65222.5 ;
      RECT  9702.5 65362.5 9567.5 65427.5 ;
      RECT  9445.0 65577.5 9310.0 65642.5 ;
      RECT  9507.5 65972.5 9572.5 66107.5 ;
      RECT  9697.5 65132.5 9762.5 65267.5 ;
      RECT  9797.5 65577.5 9662.5 65642.5 ;
      RECT  9310.0 65577.5 9445.0 65642.5 ;
      RECT  9567.5 65362.5 9702.5 65427.5 ;
      RECT  9662.5 65577.5 9797.5 65642.5 ;
      RECT  9250.0 66282.5 10170.0 66347.5 ;
      RECT  9250.0 64937.5 10170.0 65002.5 ;
      RECT  10597.5 66130.0 10662.5 66315.0 ;
      RECT  10597.5 64970.0 10662.5 65155.0 ;
      RECT  10237.5 65087.5 10302.5 64937.5 ;
      RECT  10237.5 65972.5 10302.5 66347.5 ;
      RECT  10427.5 65087.5 10492.5 65972.5 ;
      RECT  10237.5 65972.5 10302.5 66107.5 ;
      RECT  10427.5 65972.5 10492.5 66107.5 ;
      RECT  10427.5 65972.5 10492.5 66107.5 ;
      RECT  10237.5 65972.5 10302.5 66107.5 ;
      RECT  10237.5 65087.5 10302.5 65222.5 ;
      RECT  10427.5 65087.5 10492.5 65222.5 ;
      RECT  10427.5 65087.5 10492.5 65222.5 ;
      RECT  10237.5 65087.5 10302.5 65222.5 ;
      RECT  10597.5 66062.5 10662.5 66197.5 ;
      RECT  10597.5 65087.5 10662.5 65222.5 ;
      RECT  10295.0 65530.0 10360.0 65665.0 ;
      RECT  10295.0 65530.0 10360.0 65665.0 ;
      RECT  10460.0 65565.0 10525.0 65630.0 ;
      RECT  10170.0 66282.5 10730.0 66347.5 ;
      RECT  10170.0 64937.5 10730.0 65002.5 ;
      RECT  8432.5 65530.0 8497.5 65665.0 ;
      RECT  8572.5 65257.5 8637.5 65392.5 ;
      RECT  9567.5 65362.5 9432.5 65427.5 ;
      RECT  9117.5 66500.0 9182.5 66315.0 ;
      RECT  9117.5 67660.0 9182.5 67475.0 ;
      RECT  8757.5 67542.5 8822.5 67692.5 ;
      RECT  8757.5 66657.5 8822.5 66282.5 ;
      RECT  8947.5 67542.5 9012.5 66657.5 ;
      RECT  8757.5 66657.5 8822.5 66522.5 ;
      RECT  8947.5 66657.5 9012.5 66522.5 ;
      RECT  8947.5 66657.5 9012.5 66522.5 ;
      RECT  8757.5 66657.5 8822.5 66522.5 ;
      RECT  8757.5 67542.5 8822.5 67407.5 ;
      RECT  8947.5 67542.5 9012.5 67407.5 ;
      RECT  8947.5 67542.5 9012.5 67407.5 ;
      RECT  8757.5 67542.5 8822.5 67407.5 ;
      RECT  9117.5 66567.5 9182.5 66432.5 ;
      RECT  9117.5 67542.5 9182.5 67407.5 ;
      RECT  8815.0 67100.0 8880.0 66965.0 ;
      RECT  8815.0 67100.0 8880.0 66965.0 ;
      RECT  8980.0 67065.0 9045.0 67000.0 ;
      RECT  8690.0 66347.5 9250.0 66282.5 ;
      RECT  8690.0 67692.5 9250.0 67627.5 ;
      RECT  9317.5 67497.5 9382.5 67692.5 ;
      RECT  9317.5 66657.5 9382.5 66282.5 ;
      RECT  9697.5 66657.5 9762.5 66282.5 ;
      RECT  9867.5 66500.0 9932.5 66315.0 ;
      RECT  9867.5 67660.0 9932.5 67475.0 ;
      RECT  9317.5 66657.5 9382.5 66522.5 ;
      RECT  9507.5 66657.5 9572.5 66522.5 ;
      RECT  9507.5 66657.5 9572.5 66522.5 ;
      RECT  9317.5 66657.5 9382.5 66522.5 ;
      RECT  9507.5 66657.5 9572.5 66522.5 ;
      RECT  9697.5 66657.5 9762.5 66522.5 ;
      RECT  9697.5 66657.5 9762.5 66522.5 ;
      RECT  9507.5 66657.5 9572.5 66522.5 ;
      RECT  9317.5 67497.5 9382.5 67362.5 ;
      RECT  9507.5 67497.5 9572.5 67362.5 ;
      RECT  9507.5 67497.5 9572.5 67362.5 ;
      RECT  9317.5 67497.5 9382.5 67362.5 ;
      RECT  9507.5 67497.5 9572.5 67362.5 ;
      RECT  9697.5 67497.5 9762.5 67362.5 ;
      RECT  9697.5 67497.5 9762.5 67362.5 ;
      RECT  9507.5 67497.5 9572.5 67362.5 ;
      RECT  9867.5 66567.5 9932.5 66432.5 ;
      RECT  9867.5 67542.5 9932.5 67407.5 ;
      RECT  9702.5 67267.5 9567.5 67202.5 ;
      RECT  9445.0 67052.5 9310.0 66987.5 ;
      RECT  9507.5 66657.5 9572.5 66522.5 ;
      RECT  9697.5 67497.5 9762.5 67362.5 ;
      RECT  9797.5 67052.5 9662.5 66987.5 ;
      RECT  9310.0 67052.5 9445.0 66987.5 ;
      RECT  9567.5 67267.5 9702.5 67202.5 ;
      RECT  9662.5 67052.5 9797.5 66987.5 ;
      RECT  9250.0 66347.5 10170.0 66282.5 ;
      RECT  9250.0 67692.5 10170.0 67627.5 ;
      RECT  10597.5 66500.0 10662.5 66315.0 ;
      RECT  10597.5 67660.0 10662.5 67475.0 ;
      RECT  10237.5 67542.5 10302.5 67692.5 ;
      RECT  10237.5 66657.5 10302.5 66282.5 ;
      RECT  10427.5 67542.5 10492.5 66657.5 ;
      RECT  10237.5 66657.5 10302.5 66522.5 ;
      RECT  10427.5 66657.5 10492.5 66522.5 ;
      RECT  10427.5 66657.5 10492.5 66522.5 ;
      RECT  10237.5 66657.5 10302.5 66522.5 ;
      RECT  10237.5 67542.5 10302.5 67407.5 ;
      RECT  10427.5 67542.5 10492.5 67407.5 ;
      RECT  10427.5 67542.5 10492.5 67407.5 ;
      RECT  10237.5 67542.5 10302.5 67407.5 ;
      RECT  10597.5 66567.5 10662.5 66432.5 ;
      RECT  10597.5 67542.5 10662.5 67407.5 ;
      RECT  10295.0 67100.0 10360.0 66965.0 ;
      RECT  10295.0 67100.0 10360.0 66965.0 ;
      RECT  10460.0 67065.0 10525.0 67000.0 ;
      RECT  10170.0 66347.5 10730.0 66282.5 ;
      RECT  10170.0 67692.5 10730.0 67627.5 ;
      RECT  8432.5 66965.0 8497.5 67100.0 ;
      RECT  8572.5 67237.5 8637.5 67372.5 ;
      RECT  9567.5 67202.5 9432.5 67267.5 ;
      RECT  9117.5 68820.0 9182.5 69005.0 ;
      RECT  9117.5 67660.0 9182.5 67845.0 ;
      RECT  8757.5 67777.5 8822.5 67627.5 ;
      RECT  8757.5 68662.5 8822.5 69037.5 ;
      RECT  8947.5 67777.5 9012.5 68662.5 ;
      RECT  8757.5 68662.5 8822.5 68797.5 ;
      RECT  8947.5 68662.5 9012.5 68797.5 ;
      RECT  8947.5 68662.5 9012.5 68797.5 ;
      RECT  8757.5 68662.5 8822.5 68797.5 ;
      RECT  8757.5 67777.5 8822.5 67912.5 ;
      RECT  8947.5 67777.5 9012.5 67912.5 ;
      RECT  8947.5 67777.5 9012.5 67912.5 ;
      RECT  8757.5 67777.5 8822.5 67912.5 ;
      RECT  9117.5 68752.5 9182.5 68887.5 ;
      RECT  9117.5 67777.5 9182.5 67912.5 ;
      RECT  8815.0 68220.0 8880.0 68355.0 ;
      RECT  8815.0 68220.0 8880.0 68355.0 ;
      RECT  8980.0 68255.0 9045.0 68320.0 ;
      RECT  8690.0 68972.5 9250.0 69037.5 ;
      RECT  8690.0 67627.5 9250.0 67692.5 ;
      RECT  9317.5 67822.5 9382.5 67627.5 ;
      RECT  9317.5 68662.5 9382.5 69037.5 ;
      RECT  9697.5 68662.5 9762.5 69037.5 ;
      RECT  9867.5 68820.0 9932.5 69005.0 ;
      RECT  9867.5 67660.0 9932.5 67845.0 ;
      RECT  9317.5 68662.5 9382.5 68797.5 ;
      RECT  9507.5 68662.5 9572.5 68797.5 ;
      RECT  9507.5 68662.5 9572.5 68797.5 ;
      RECT  9317.5 68662.5 9382.5 68797.5 ;
      RECT  9507.5 68662.5 9572.5 68797.5 ;
      RECT  9697.5 68662.5 9762.5 68797.5 ;
      RECT  9697.5 68662.5 9762.5 68797.5 ;
      RECT  9507.5 68662.5 9572.5 68797.5 ;
      RECT  9317.5 67822.5 9382.5 67957.5 ;
      RECT  9507.5 67822.5 9572.5 67957.5 ;
      RECT  9507.5 67822.5 9572.5 67957.5 ;
      RECT  9317.5 67822.5 9382.5 67957.5 ;
      RECT  9507.5 67822.5 9572.5 67957.5 ;
      RECT  9697.5 67822.5 9762.5 67957.5 ;
      RECT  9697.5 67822.5 9762.5 67957.5 ;
      RECT  9507.5 67822.5 9572.5 67957.5 ;
      RECT  9867.5 68752.5 9932.5 68887.5 ;
      RECT  9867.5 67777.5 9932.5 67912.5 ;
      RECT  9702.5 68052.5 9567.5 68117.5 ;
      RECT  9445.0 68267.5 9310.0 68332.5 ;
      RECT  9507.5 68662.5 9572.5 68797.5 ;
      RECT  9697.5 67822.5 9762.5 67957.5 ;
      RECT  9797.5 68267.5 9662.5 68332.5 ;
      RECT  9310.0 68267.5 9445.0 68332.5 ;
      RECT  9567.5 68052.5 9702.5 68117.5 ;
      RECT  9662.5 68267.5 9797.5 68332.5 ;
      RECT  9250.0 68972.5 10170.0 69037.5 ;
      RECT  9250.0 67627.5 10170.0 67692.5 ;
      RECT  10597.5 68820.0 10662.5 69005.0 ;
      RECT  10597.5 67660.0 10662.5 67845.0 ;
      RECT  10237.5 67777.5 10302.5 67627.5 ;
      RECT  10237.5 68662.5 10302.5 69037.5 ;
      RECT  10427.5 67777.5 10492.5 68662.5 ;
      RECT  10237.5 68662.5 10302.5 68797.5 ;
      RECT  10427.5 68662.5 10492.5 68797.5 ;
      RECT  10427.5 68662.5 10492.5 68797.5 ;
      RECT  10237.5 68662.5 10302.5 68797.5 ;
      RECT  10237.5 67777.5 10302.5 67912.5 ;
      RECT  10427.5 67777.5 10492.5 67912.5 ;
      RECT  10427.5 67777.5 10492.5 67912.5 ;
      RECT  10237.5 67777.5 10302.5 67912.5 ;
      RECT  10597.5 68752.5 10662.5 68887.5 ;
      RECT  10597.5 67777.5 10662.5 67912.5 ;
      RECT  10295.0 68220.0 10360.0 68355.0 ;
      RECT  10295.0 68220.0 10360.0 68355.0 ;
      RECT  10460.0 68255.0 10525.0 68320.0 ;
      RECT  10170.0 68972.5 10730.0 69037.5 ;
      RECT  10170.0 67627.5 10730.0 67692.5 ;
      RECT  8432.5 68220.0 8497.5 68355.0 ;
      RECT  8572.5 67947.5 8637.5 68082.5 ;
      RECT  9567.5 68052.5 9432.5 68117.5 ;
      RECT  9117.5 69190.0 9182.5 69005.0 ;
      RECT  9117.5 70350.0 9182.5 70165.0 ;
      RECT  8757.5 70232.5 8822.5 70382.5 ;
      RECT  8757.5 69347.5 8822.5 68972.5 ;
      RECT  8947.5 70232.5 9012.5 69347.5 ;
      RECT  8757.5 69347.5 8822.5 69212.5 ;
      RECT  8947.5 69347.5 9012.5 69212.5 ;
      RECT  8947.5 69347.5 9012.5 69212.5 ;
      RECT  8757.5 69347.5 8822.5 69212.5 ;
      RECT  8757.5 70232.5 8822.5 70097.5 ;
      RECT  8947.5 70232.5 9012.5 70097.5 ;
      RECT  8947.5 70232.5 9012.5 70097.5 ;
      RECT  8757.5 70232.5 8822.5 70097.5 ;
      RECT  9117.5 69257.5 9182.5 69122.5 ;
      RECT  9117.5 70232.5 9182.5 70097.5 ;
      RECT  8815.0 69790.0 8880.0 69655.0 ;
      RECT  8815.0 69790.0 8880.0 69655.0 ;
      RECT  8980.0 69755.0 9045.0 69690.0 ;
      RECT  8690.0 69037.5 9250.0 68972.5 ;
      RECT  8690.0 70382.5 9250.0 70317.5 ;
      RECT  9317.5 70187.5 9382.5 70382.5 ;
      RECT  9317.5 69347.5 9382.5 68972.5 ;
      RECT  9697.5 69347.5 9762.5 68972.5 ;
      RECT  9867.5 69190.0 9932.5 69005.0 ;
      RECT  9867.5 70350.0 9932.5 70165.0 ;
      RECT  9317.5 69347.5 9382.5 69212.5 ;
      RECT  9507.5 69347.5 9572.5 69212.5 ;
      RECT  9507.5 69347.5 9572.5 69212.5 ;
      RECT  9317.5 69347.5 9382.5 69212.5 ;
      RECT  9507.5 69347.5 9572.5 69212.5 ;
      RECT  9697.5 69347.5 9762.5 69212.5 ;
      RECT  9697.5 69347.5 9762.5 69212.5 ;
      RECT  9507.5 69347.5 9572.5 69212.5 ;
      RECT  9317.5 70187.5 9382.5 70052.5 ;
      RECT  9507.5 70187.5 9572.5 70052.5 ;
      RECT  9507.5 70187.5 9572.5 70052.5 ;
      RECT  9317.5 70187.5 9382.5 70052.5 ;
      RECT  9507.5 70187.5 9572.5 70052.5 ;
      RECT  9697.5 70187.5 9762.5 70052.5 ;
      RECT  9697.5 70187.5 9762.5 70052.5 ;
      RECT  9507.5 70187.5 9572.5 70052.5 ;
      RECT  9867.5 69257.5 9932.5 69122.5 ;
      RECT  9867.5 70232.5 9932.5 70097.5 ;
      RECT  9702.5 69957.5 9567.5 69892.5 ;
      RECT  9445.0 69742.5 9310.0 69677.5 ;
      RECT  9507.5 69347.5 9572.5 69212.5 ;
      RECT  9697.5 70187.5 9762.5 70052.5 ;
      RECT  9797.5 69742.5 9662.5 69677.5 ;
      RECT  9310.0 69742.5 9445.0 69677.5 ;
      RECT  9567.5 69957.5 9702.5 69892.5 ;
      RECT  9662.5 69742.5 9797.5 69677.5 ;
      RECT  9250.0 69037.5 10170.0 68972.5 ;
      RECT  9250.0 70382.5 10170.0 70317.5 ;
      RECT  10597.5 69190.0 10662.5 69005.0 ;
      RECT  10597.5 70350.0 10662.5 70165.0 ;
      RECT  10237.5 70232.5 10302.5 70382.5 ;
      RECT  10237.5 69347.5 10302.5 68972.5 ;
      RECT  10427.5 70232.5 10492.5 69347.5 ;
      RECT  10237.5 69347.5 10302.5 69212.5 ;
      RECT  10427.5 69347.5 10492.5 69212.5 ;
      RECT  10427.5 69347.5 10492.5 69212.5 ;
      RECT  10237.5 69347.5 10302.5 69212.5 ;
      RECT  10237.5 70232.5 10302.5 70097.5 ;
      RECT  10427.5 70232.5 10492.5 70097.5 ;
      RECT  10427.5 70232.5 10492.5 70097.5 ;
      RECT  10237.5 70232.5 10302.5 70097.5 ;
      RECT  10597.5 69257.5 10662.5 69122.5 ;
      RECT  10597.5 70232.5 10662.5 70097.5 ;
      RECT  10295.0 69790.0 10360.0 69655.0 ;
      RECT  10295.0 69790.0 10360.0 69655.0 ;
      RECT  10460.0 69755.0 10525.0 69690.0 ;
      RECT  10170.0 69037.5 10730.0 68972.5 ;
      RECT  10170.0 70382.5 10730.0 70317.5 ;
      RECT  8432.5 69655.0 8497.5 69790.0 ;
      RECT  8572.5 69927.5 8637.5 70062.5 ;
      RECT  9567.5 69892.5 9432.5 69957.5 ;
      RECT  8235.0 27632.5 8605.0 27697.5 ;
      RECT  8235.0 29612.5 8605.0 29677.5 ;
      RECT  8235.0 30322.5 8605.0 30387.5 ;
      RECT  8235.0 32302.5 8605.0 32367.5 ;
      RECT  8235.0 33012.5 8605.0 33077.5 ;
      RECT  8235.0 34992.5 8605.0 35057.5 ;
      RECT  8235.0 35702.5 8605.0 35767.5 ;
      RECT  8235.0 37682.5 8605.0 37747.5 ;
      RECT  8235.0 38392.5 8605.0 38457.5 ;
      RECT  8235.0 40372.5 8605.0 40437.5 ;
      RECT  8235.0 41082.5 8605.0 41147.5 ;
      RECT  8235.0 43062.5 8605.0 43127.5 ;
      RECT  8235.0 43772.5 8605.0 43837.5 ;
      RECT  8235.0 45752.5 8605.0 45817.5 ;
      RECT  8235.0 46462.5 8605.0 46527.5 ;
      RECT  8235.0 48442.5 8605.0 48507.5 ;
      RECT  8235.0 49152.5 8605.0 49217.5 ;
      RECT  8235.0 51132.5 8605.0 51197.5 ;
      RECT  8235.0 51842.5 8605.0 51907.5 ;
      RECT  8235.0 53822.5 8605.0 53887.5 ;
      RECT  8235.0 54532.5 8605.0 54597.5 ;
      RECT  8235.0 56512.5 8605.0 56577.5 ;
      RECT  8235.0 57222.5 8605.0 57287.5 ;
      RECT  8235.0 59202.5 8605.0 59267.5 ;
      RECT  8235.0 59912.5 8605.0 59977.5 ;
      RECT  8235.0 61892.5 8605.0 61957.5 ;
      RECT  8235.0 62602.5 8605.0 62667.5 ;
      RECT  8235.0 64582.5 8605.0 64647.5 ;
      RECT  8235.0 65292.5 8605.0 65357.5 ;
      RECT  8235.0 67272.5 8605.0 67337.5 ;
      RECT  8235.0 67982.5 8605.0 68047.5 ;
      RECT  8235.0 69962.5 8605.0 70027.5 ;
      RECT  10460.0 27905.0 10525.0 27970.0 ;
      RECT  10460.0 29340.0 10525.0 29405.0 ;
      RECT  10460.0 30595.0 10525.0 30660.0 ;
      RECT  10460.0 32030.0 10525.0 32095.0 ;
      RECT  10460.0 33285.0 10525.0 33350.0 ;
      RECT  10460.0 34720.0 10525.0 34785.0 ;
      RECT  10460.0 35975.0 10525.0 36040.0 ;
      RECT  10460.0 37410.0 10525.0 37475.0 ;
      RECT  10460.0 38665.0 10525.0 38730.0 ;
      RECT  10460.0 40100.0 10525.0 40165.0 ;
      RECT  10460.0 41355.0 10525.0 41420.0 ;
      RECT  10460.0 42790.0 10525.0 42855.0 ;
      RECT  10460.0 44045.0 10525.0 44110.0 ;
      RECT  10460.0 45480.0 10525.0 45545.0 ;
      RECT  10460.0 46735.0 10525.0 46800.0 ;
      RECT  10460.0 48170.0 10525.0 48235.0 ;
      RECT  10460.0 49425.0 10525.0 49490.0 ;
      RECT  10460.0 50860.0 10525.0 50925.0 ;
      RECT  10460.0 52115.0 10525.0 52180.0 ;
      RECT  10460.0 53550.0 10525.0 53615.0 ;
      RECT  10460.0 54805.0 10525.0 54870.0 ;
      RECT  10460.0 56240.0 10525.0 56305.0 ;
      RECT  10460.0 57495.0 10525.0 57560.0 ;
      RECT  10460.0 58930.0 10525.0 58995.0 ;
      RECT  10460.0 60185.0 10525.0 60250.0 ;
      RECT  10460.0 61620.0 10525.0 61685.0 ;
      RECT  10460.0 62875.0 10525.0 62940.0 ;
      RECT  10460.0 64310.0 10525.0 64375.0 ;
      RECT  10460.0 65565.0 10525.0 65630.0 ;
      RECT  10460.0 67000.0 10525.0 67065.0 ;
      RECT  10460.0 68255.0 10525.0 68320.0 ;
      RECT  10460.0 69690.0 10525.0 69755.0 ;
      RECT  8235.0 28622.5 8690.0 28687.5 ;
      RECT  8235.0 31312.5 8690.0 31377.5 ;
      RECT  8235.0 34002.5 8690.0 34067.5 ;
      RECT  8235.0 36692.5 8690.0 36757.5 ;
      RECT  8235.0 39382.5 8690.0 39447.5 ;
      RECT  8235.0 42072.5 8690.0 42137.5 ;
      RECT  8235.0 44762.5 8690.0 44827.5 ;
      RECT  8235.0 47452.5 8690.0 47517.5 ;
      RECT  8235.0 50142.5 8690.0 50207.5 ;
      RECT  8235.0 52832.5 8690.0 52897.5 ;
      RECT  8235.0 55522.5 8690.0 55587.5 ;
      RECT  8235.0 58212.5 8690.0 58277.5 ;
      RECT  8235.0 60902.5 8690.0 60967.5 ;
      RECT  8235.0 63592.5 8690.0 63657.5 ;
      RECT  8235.0 66282.5 8690.0 66347.5 ;
      RECT  8235.0 68972.5 8690.0 69037.5 ;
      RECT  8235.0 27277.5 8690.0 27342.5 ;
      RECT  8235.0 29967.5 8690.0 30032.5 ;
      RECT  8235.0 32657.5 8690.0 32722.5 ;
      RECT  8235.0 35347.5 8690.0 35412.5 ;
      RECT  8235.0 38037.5 8690.0 38102.5 ;
      RECT  8235.0 40727.5 8690.0 40792.5 ;
      RECT  8235.0 43417.5 8690.0 43482.5 ;
      RECT  8235.0 46107.5 8690.0 46172.5 ;
      RECT  8235.0 48797.5 8690.0 48862.5 ;
      RECT  8235.0 51487.5 8690.0 51552.5 ;
      RECT  8235.0 54177.5 8690.0 54242.5 ;
      RECT  8235.0 56867.5 8690.0 56932.5 ;
      RECT  8235.0 59557.5 8690.0 59622.5 ;
      RECT  8235.0 62247.5 8690.0 62312.5 ;
      RECT  8235.0 64937.5 8690.0 65002.5 ;
      RECT  8235.0 67627.5 8690.0 67692.5 ;
      RECT  8235.0 70317.5 8690.0 70382.5 ;
      RECT  4655.0 10760.0 11095.0 10055.0 ;
      RECT  4655.0 9350.0 11095.0 10055.0 ;
      RECT  4655.0 9350.0 11095.0 8645.0 ;
      RECT  4655.0 7940.0 11095.0 8645.0 ;
      RECT  4655.0 7940.0 11095.0 7235.0 ;
      RECT  4655.0 6530.0 11095.0 7235.0 ;
      RECT  4655.0 6530.0 11095.0 5825.0 ;
      RECT  4860.0 10760.0 4925.0 5825.0 ;
      RECT  7865.0 10760.0 7930.0 5825.0 ;
      RECT  10825.0 10760.0 10890.0 5825.0 ;
      RECT  5875.0 10760.0 5940.0 5825.0 ;
      RECT  8835.0 10760.0 8900.0 5825.0 ;
      RECT  5020.0 10760.0 5085.0 5825.0 ;
      RECT  13992.5 27342.5 14127.5 27277.5 ;
      RECT  13992.5 30032.5 14127.5 29967.5 ;
      RECT  13992.5 32722.5 14127.5 32657.5 ;
      RECT  13992.5 35412.5 14127.5 35347.5 ;
      RECT  13992.5 38102.5 14127.5 38037.5 ;
      RECT  13992.5 40792.5 14127.5 40727.5 ;
      RECT  13992.5 43482.5 14127.5 43417.5 ;
      RECT  13992.5 46172.5 14127.5 46107.5 ;
      RECT  13992.5 48862.5 14127.5 48797.5 ;
      RECT  13992.5 51552.5 14127.5 51487.5 ;
      RECT  13992.5 54242.5 14127.5 54177.5 ;
      RECT  13992.5 56932.5 14127.5 56867.5 ;
      RECT  13992.5 59622.5 14127.5 59557.5 ;
      RECT  13992.5 62312.5 14127.5 62247.5 ;
      RECT  13992.5 65002.5 14127.5 64937.5 ;
      RECT  13992.5 67692.5 14127.5 67627.5 ;
      RECT  13992.5 70382.5 14127.5 70317.5 ;
      RECT  10720.0 11342.5 10585.0 11407.5 ;
      RECT  12045.0 11342.5 11910.0 11407.5 ;
      RECT  10445.0 12687.5 10310.0 12752.5 ;
      RECT  12250.0 12687.5 12115.0 12752.5 ;
      RECT  11635.0 16722.5 11500.0 16787.5 ;
      RECT  12455.0 16722.5 12320.0 16787.5 ;
      RECT  11360.0 18067.5 11225.0 18132.5 ;
      RECT  12660.0 18067.5 12525.0 18132.5 ;
      RECT  11085.0 19412.5 10950.0 19477.5 ;
      RECT  12865.0 19412.5 12730.0 19477.5 ;
      RECT  11840.0 11137.5 11705.0 11202.5 ;
      RECT  11840.0 13827.5 11705.0 13892.5 ;
      RECT  11840.0 16517.5 11705.0 16582.5 ;
      RECT  11840.0 19207.5 11705.0 19272.5 ;
      RECT  11840.0 21897.5 11705.0 21962.5 ;
      RECT  11840.0 24587.5 11705.0 24652.5 ;
      RECT  13070.0 25307.5 12935.0 25372.5 ;
      RECT  13275.0 25167.5 13140.0 25232.5 ;
      RECT  13480.0 25027.5 13345.0 25092.5 ;
      RECT  13685.0 24887.5 13550.0 24952.5 ;
      RECT  13070.0 630.0 12935.0 695.0 ;
      RECT  13275.0 2065.0 13140.0 2130.0 ;
      RECT  13480.0 3320.0 13345.0 3385.0 ;
      RECT  13685.0 4755.0 13550.0 4820.0 ;
      RECT  13992.5 67.5 14127.5 2.5 ;
      RECT  13992.5 2757.5 14127.5 2692.5 ;
      RECT  13992.5 5447.5 14127.5 5382.5 ;
      RECT  11162.5 10375.0 11027.5 10440.0 ;
      RECT  12045.0 10375.0 11910.0 10440.0 ;
      RECT  11162.5 9670.0 11027.5 9735.0 ;
      RECT  12250.0 9670.0 12115.0 9735.0 ;
      RECT  11162.5 8965.0 11027.5 9030.0 ;
      RECT  12455.0 8965.0 12320.0 9030.0 ;
      RECT  11162.5 8260.0 11027.5 8325.0 ;
      RECT  12660.0 8260.0 12525.0 8325.0 ;
      RECT  11162.5 7555.0 11027.5 7620.0 ;
      RECT  12865.0 7555.0 12730.0 7620.0 ;
      RECT  11230.0 10727.5 11095.0 10792.5 ;
      RECT  14127.5 10727.5 13992.5 10792.5 ;
      RECT  11230.0 10022.5 11095.0 10087.5 ;
      RECT  14127.5 10022.5 13992.5 10087.5 ;
      RECT  11230.0 9317.5 11095.0 9382.5 ;
      RECT  14127.5 9317.5 13992.5 9382.5 ;
      RECT  11230.0 8612.5 11095.0 8677.5 ;
      RECT  14127.5 8612.5 13992.5 8677.5 ;
      RECT  11230.0 7907.5 11095.0 7972.5 ;
      RECT  14127.5 7907.5 13992.5 7972.5 ;
      RECT  11230.0 7202.5 11095.0 7267.5 ;
      RECT  14127.5 7202.5 13992.5 7267.5 ;
      RECT  11230.0 6497.5 11095.0 6562.5 ;
      RECT  14127.5 6497.5 13992.5 6562.5 ;
      RECT  11230.0 5792.5 11095.0 5857.5 ;
      RECT  14127.5 5792.5 13992.5 5857.5 ;
      RECT  15265.0 9170.0 15130.0 9235.0 ;
      RECT  14855.0 6985.0 14720.0 7050.0 ;
      RECT  15060.0 8532.5 14925.0 8597.5 ;
      RECT  15265.0 71327.5 15130.0 71392.5 ;
      RECT  15470.0 15672.5 15335.0 15737.5 ;
      RECT  15675.0 19697.5 15540.0 19762.5 ;
      RECT  14650.0 10932.5 14515.0 10997.5 ;
      RECT  8532.5 70522.5 8397.5 70587.5 ;
      RECT  14650.0 70522.5 14515.0 70587.5 ;
      RECT  14342.5 8402.5 14207.5 8467.5 ;
      RECT  14342.5 19827.5 14207.5 19892.5 ;
      RECT  14342.5 9330.0 14207.5 9395.0 ;
      RECT  14342.5 16605.0 14207.5 16670.0 ;
      RECT  21920.0 35.0 22270.0 72077.5 ;
      RECT  4175.0 35.0 4525.0 72077.5 ;
      RECT  3455.0 27740.0 3390.0 27805.0 ;
      RECT  3422.5 27740.0 3407.5 27805.0 ;
      RECT  3455.0 27772.5 3390.0 28357.5 ;
      RECT  3455.0 28902.5 3390.0 29297.5 ;
      RECT  3455.0 30222.5 3390.0 30807.5 ;
      RECT  2657.5 30660.0 2280.0 30725.0 ;
      RECT  2657.5 33620.0 2280.0 33685.0 ;
      RECT  2657.5 28670.0 2280.0 28735.0 ;
      RECT  2657.5 31630.0 2280.0 31695.0 ;
      RECT  3440.0 27740.0 3375.0 27805.0 ;
      RECT  3455.0 28870.0 3390.0 28935.0 ;
      RECT  2005.0 39555.0 1940.0 40320.0 ;
      RECT  3455.0 32905.0 3390.0 34335.0 ;
      RECT  2485.0 27655.0 2280.0 27720.0 ;
      RECT  1962.5 34335.0 1897.5 36272.5 ;
      RECT  1747.5 34745.0 1682.5 36530.0 ;
      RECT  3380.0 35770.0 3315.0 36340.0 ;
      RECT  3520.0 35565.0 3455.0 36530.0 ;
      RECT  3660.0 34950.0 3595.0 36720.0 ;
      RECT  3380.0 37280.0 3315.0 37345.0 ;
      RECT  3380.0 36815.0 3315.0 37312.5 ;
      RECT  3407.5 37280.0 3347.5 37345.0 ;
      RECT  3475.0 37445.0 3410.0 37510.0 ;
      RECT  3442.5 37445.0 3407.5 37510.0 ;
      RECT  3475.0 37477.5 3410.0 41017.5 ;
      RECT  690.0 35770.0 625.0 36900.0 ;
      RECT  830.0 34950.0 765.0 37090.0 ;
      RECT  970.0 35155.0 905.0 37280.0 ;
      RECT  690.0 37840.0 625.0 37905.0 ;
      RECT  690.0 37375.0 625.0 37872.5 ;
      RECT  717.5 37840.0 657.5 37905.0 ;
      RECT  750.0 38037.5 685.0 38432.5 ;
      RECT  750.0 38597.5 685.0 38992.5 ;
      RECT  2005.0 39522.5 1940.0 39587.5 ;
      RECT  1972.5 39522.5 1940.0 39587.5 ;
      RECT  2005.0 39430.0 1940.0 39555.0 ;
      RECT  2005.0 38837.5 1940.0 39232.5 ;
      RECT  1962.5 36695.0 1897.5 37065.0 ;
      RECT  2017.5 37770.0 1952.5 38210.0 ;
      RECT  750.0 39157.5 685.0 39395.0 ;
      RECT  2005.0 38435.0 1940.0 38672.5 ;
      RECT  4067.5 27450.0 4002.5 39555.0 ;
      RECT  4067.5 34540.0 4002.5 36145.0 ;
      RECT  2722.5 27450.0 2657.5 39555.0 ;
      RECT  2722.5 35360.0 2657.5 36145.0 ;
      RECT  1377.5 36145.0 1312.5 39555.0 ;
      RECT  1377.5 34540.0 1312.5 36145.0 ;
      RECT  32.5 36145.0 -32.5 39555.0 ;
      RECT  32.5 35360.0 -32.5 36145.0 ;
      RECT  32.5 39522.5 -32.5 39587.5 ;
      RECT  32.5 39350.0 -32.5 39555.0 ;
      RECT  8.881784197e-13 39522.5 -45.0 39587.5 ;
      RECT  165.0 27450.0 870.0 33890.0 ;
      RECT  1575.0 27450.0 870.0 33890.0 ;
      RECT  1575.0 27450.0 2280.0 33890.0 ;
      RECT  165.0 27655.0 2280.0 27720.0 ;
      RECT  165.0 30660.0 2280.0 30725.0 ;
      RECT  165.0 33620.0 2280.0 33685.0 ;
      RECT  165.0 28670.0 2280.0 28735.0 ;
      RECT  165.0 31630.0 2280.0 31695.0 ;
      RECT  165.0 27815.0 2280.0 27880.0 ;
      RECT  2875.0 28067.5 2690.0 28132.5 ;
      RECT  4035.0 28067.5 3850.0 28132.5 ;
      RECT  2832.5 27517.5 2657.5 27962.5 ;
      RECT  3917.5 27707.5 3032.5 27772.5 ;
      RECT  2965.0 27517.5 2800.0 27582.5 ;
      RECT  2965.0 27897.5 2800.0 27962.5 ;
      RECT  3032.5 27517.5 2897.5 27582.5 ;
      RECT  3032.5 27897.5 2897.5 27962.5 ;
      RECT  3032.5 27707.5 2897.5 27772.5 ;
      RECT  3032.5 27707.5 2897.5 27772.5 ;
      RECT  2832.5 27517.5 2767.5 27962.5 ;
      RECT  4015.0 27517.5 3850.0 27582.5 ;
      RECT  4015.0 27897.5 3850.0 27962.5 ;
      RECT  3917.5 27517.5 3782.5 27582.5 ;
      RECT  3917.5 27897.5 3782.5 27962.5 ;
      RECT  3917.5 27707.5 3782.5 27772.5 ;
      RECT  3917.5 27707.5 3782.5 27772.5 ;
      RECT  4047.5 27517.5 3982.5 27962.5 ;
      RECT  2942.5 28067.5 2807.5 28132.5 ;
      RECT  3917.5 28067.5 3782.5 28132.5 ;
      RECT  3475.0 27575.0 3340.0 27640.0 ;
      RECT  3475.0 27575.0 3340.0 27640.0 ;
      RECT  3440.0 27740.0 3375.0 27805.0 ;
      RECT  2722.5 27450.0 2657.5 28200.0 ;
      RECT  4067.5 27450.0 4002.5 28200.0 ;
      RECT  2875.0 29007.5 2690.0 29072.5 ;
      RECT  4035.0 29007.5 3850.0 29072.5 ;
      RECT  2877.5 28267.5 2657.5 28712.5 ;
      RECT  3702.5 28837.5 3207.5 28902.5 ;
      RECT  3010.0 28267.5 2845.0 28332.5 ;
      RECT  3010.0 28647.5 2845.0 28712.5 ;
      RECT  3175.0 28457.5 3010.0 28522.5 ;
      RECT  3175.0 28837.5 3010.0 28902.5 ;
      RECT  3077.5 28267.5 2942.5 28332.5 ;
      RECT  3077.5 28647.5 2942.5 28712.5 ;
      RECT  3077.5 28457.5 2942.5 28522.5 ;
      RECT  3077.5 28837.5 2942.5 28902.5 ;
      RECT  3207.5 28457.5 3142.5 28902.5 ;
      RECT  2877.5 28267.5 2812.5 28712.5 ;
      RECT  4000.0 28267.5 3835.0 28332.5 ;
      RECT  4000.0 28647.5 3835.0 28712.5 ;
      RECT  3835.0 28457.5 3670.0 28522.5 ;
      RECT  3835.0 28837.5 3670.0 28902.5 ;
      RECT  3902.5 28267.5 3767.5 28332.5 ;
      RECT  3902.5 28647.5 3767.5 28712.5 ;
      RECT  3902.5 28457.5 3767.5 28522.5 ;
      RECT  3902.5 28837.5 3767.5 28902.5 ;
      RECT  3702.5 28457.5 3637.5 28902.5 ;
      RECT  4032.5 28267.5 3967.5 28712.5 ;
      RECT  2942.5 29007.5 2807.5 29072.5 ;
      RECT  3917.5 29007.5 3782.5 29072.5 ;
      RECT  3490.0 28325.0 3355.0 28390.0 ;
      RECT  3490.0 28325.0 3355.0 28390.0 ;
      RECT  3455.0 28870.0 3390.0 28935.0 ;
      RECT  2722.5 28200.0 2657.5 29140.0 ;
      RECT  4067.5 28200.0 4002.5 29140.0 ;
      RECT  2875.0 30517.5 2690.0 30582.5 ;
      RECT  4035.0 30517.5 3850.0 30582.5 ;
      RECT  2877.5 29207.5 2657.5 30412.5 ;
      RECT  3702.5 30157.5 3207.5 30222.5 ;
      RECT  3010.0 29207.5 2845.0 29272.5 ;
      RECT  3010.0 29587.5 2845.0 29652.5 ;
      RECT  3010.0 29967.5 2845.0 30032.5 ;
      RECT  3010.0 30347.5 2845.0 30412.5 ;
      RECT  3175.0 29397.5 3010.0 29462.5 ;
      RECT  3175.0 29777.5 3010.0 29842.5 ;
      RECT  3175.0 30157.5 3010.0 30222.5 ;
      RECT  3077.5 29207.5 2942.5 29272.5 ;
      RECT  3077.5 29587.5 2942.5 29652.5 ;
      RECT  3077.5 29967.5 2942.5 30032.5 ;
      RECT  3077.5 30347.5 2942.5 30412.5 ;
      RECT  3077.5 29397.5 2942.5 29462.5 ;
      RECT  3077.5 29777.5 2942.5 29842.5 ;
      RECT  3077.5 30157.5 2942.5 30222.5 ;
      RECT  3207.5 29397.5 3142.5 30222.5 ;
      RECT  2877.5 29207.5 2812.5 30412.5 ;
      RECT  4000.0 29207.5 3835.0 29272.5 ;
      RECT  4000.0 29587.5 3835.0 29652.5 ;
      RECT  4000.0 29967.5 3835.0 30032.5 ;
      RECT  4000.0 30347.5 3835.0 30412.5 ;
      RECT  3835.0 29397.5 3670.0 29462.5 ;
      RECT  3835.0 29777.5 3670.0 29842.5 ;
      RECT  3835.0 30157.5 3670.0 30222.5 ;
      RECT  3902.5 29207.5 3767.5 29272.5 ;
      RECT  3902.5 29587.5 3767.5 29652.5 ;
      RECT  3902.5 29967.5 3767.5 30032.5 ;
      RECT  3902.5 30347.5 3767.5 30412.5 ;
      RECT  3902.5 29397.5 3767.5 29462.5 ;
      RECT  3902.5 29777.5 3767.5 29842.5 ;
      RECT  3902.5 30157.5 3767.5 30222.5 ;
      RECT  3702.5 29397.5 3637.5 30222.5 ;
      RECT  4032.5 29207.5 3967.5 30412.5 ;
      RECT  2942.5 30517.5 2807.5 30582.5 ;
      RECT  3917.5 30517.5 3782.5 30582.5 ;
      RECT  3490.0 29265.0 3355.0 29330.0 ;
      RECT  3490.0 29265.0 3355.0 29330.0 ;
      RECT  3455.0 30190.0 3390.0 30255.0 ;
      RECT  2722.5 29140.0 2657.5 30650.0 ;
      RECT  4067.5 29140.0 4002.5 30650.0 ;
      RECT  2875.0 33167.5 2690.0 33232.5 ;
      RECT  4035.0 33167.5 3850.0 33232.5 ;
      RECT  2877.5 30717.5 2657.5 33062.5 ;
      RECT  3702.5 32807.5 3207.5 32872.5 ;
      RECT  3010.0 30717.5 2845.0 30782.5 ;
      RECT  3010.0 31097.5 2845.0 31162.5 ;
      RECT  3010.0 31477.5 2845.0 31542.5 ;
      RECT  3010.0 31857.5 2845.0 31922.5 ;
      RECT  3010.0 32237.5 2845.0 32302.5 ;
      RECT  3010.0 32617.5 2845.0 32682.5 ;
      RECT  3010.0 32997.5 2845.0 33062.5 ;
      RECT  3175.0 30907.5 3010.0 30972.5 ;
      RECT  3175.0 31287.5 3010.0 31352.5 ;
      RECT  3175.0 31667.5 3010.0 31732.5 ;
      RECT  3175.0 32047.5 3010.0 32112.5 ;
      RECT  3175.0 32427.5 3010.0 32492.5 ;
      RECT  3175.0 32807.5 3010.0 32872.5 ;
      RECT  3077.5 30717.5 2942.5 30782.5 ;
      RECT  3077.5 31097.5 2942.5 31162.5 ;
      RECT  3077.5 31477.5 2942.5 31542.5 ;
      RECT  3077.5 31857.5 2942.5 31922.5 ;
      RECT  3077.5 32237.5 2942.5 32302.5 ;
      RECT  3077.5 32617.5 2942.5 32682.5 ;
      RECT  3077.5 32997.5 2942.5 33062.5 ;
      RECT  3077.5 30907.5 2942.5 30972.5 ;
      RECT  3077.5 31287.5 2942.5 31352.5 ;
      RECT  3077.5 31667.5 2942.5 31732.5 ;
      RECT  3077.5 32047.5 2942.5 32112.5 ;
      RECT  3077.5 32427.5 2942.5 32492.5 ;
      RECT  3077.5 32807.5 2942.5 32872.5 ;
      RECT  3207.5 30907.5 3142.5 32872.5 ;
      RECT  2877.5 30717.5 2812.5 33062.5 ;
      RECT  4000.0 30717.5 3835.0 30782.5 ;
      RECT  4000.0 31097.5 3835.0 31162.5 ;
      RECT  4000.0 31477.5 3835.0 31542.5 ;
      RECT  4000.0 31857.5 3835.0 31922.5 ;
      RECT  4000.0 32237.5 3835.0 32302.5 ;
      RECT  4000.0 32617.5 3835.0 32682.5 ;
      RECT  4000.0 32997.5 3835.0 33062.5 ;
      RECT  3835.0 30907.5 3670.0 30972.5 ;
      RECT  3835.0 31287.5 3670.0 31352.5 ;
      RECT  3835.0 31667.5 3670.0 31732.5 ;
      RECT  3835.0 32047.5 3670.0 32112.5 ;
      RECT  3835.0 32427.5 3670.0 32492.5 ;
      RECT  3835.0 32807.5 3670.0 32872.5 ;
      RECT  3902.5 30717.5 3767.5 30782.5 ;
      RECT  3902.5 31097.5 3767.5 31162.5 ;
      RECT  3902.5 31477.5 3767.5 31542.5 ;
      RECT  3902.5 31857.5 3767.5 31922.5 ;
      RECT  3902.5 32237.5 3767.5 32302.5 ;
      RECT  3902.5 32617.5 3767.5 32682.5 ;
      RECT  3902.5 32997.5 3767.5 33062.5 ;
      RECT  3902.5 30907.5 3767.5 30972.5 ;
      RECT  3902.5 31287.5 3767.5 31352.5 ;
      RECT  3902.5 31667.5 3767.5 31732.5 ;
      RECT  3902.5 32047.5 3767.5 32112.5 ;
      RECT  3902.5 32427.5 3767.5 32492.5 ;
      RECT  3902.5 32807.5 3767.5 32872.5 ;
      RECT  3702.5 30907.5 3637.5 32872.5 ;
      RECT  4032.5 30717.5 3967.5 33062.5 ;
      RECT  2942.5 33167.5 2807.5 33232.5 ;
      RECT  3917.5 33167.5 3782.5 33232.5 ;
      RECT  3490.0 30775.0 3355.0 30840.0 ;
      RECT  3490.0 30775.0 3355.0 30840.0 ;
      RECT  3455.0 32840.0 3390.0 32905.0 ;
      RECT  2722.5 30650.0 2657.5 33300.0 ;
      RECT  4067.5 30650.0 4002.5 33300.0 ;
      RECT  3872.5 36212.5 4067.5 36277.5 ;
      RECT  3032.5 36212.5 2657.5 36277.5 ;
      RECT  3032.5 36592.5 2657.5 36657.5 ;
      RECT  2875.0 36952.5 2690.0 37017.5 ;
      RECT  4035.0 36952.5 3850.0 37017.5 ;
      RECT  3032.5 36212.5 2897.5 36277.5 ;
      RECT  3032.5 36402.5 2897.5 36467.5 ;
      RECT  3032.5 36402.5 2897.5 36467.5 ;
      RECT  3032.5 36212.5 2897.5 36277.5 ;
      RECT  3032.5 36402.5 2897.5 36467.5 ;
      RECT  3032.5 36592.5 2897.5 36657.5 ;
      RECT  3032.5 36592.5 2897.5 36657.5 ;
      RECT  3032.5 36402.5 2897.5 36467.5 ;
      RECT  3032.5 36592.5 2897.5 36657.5 ;
      RECT  3032.5 36782.5 2897.5 36847.5 ;
      RECT  3032.5 36782.5 2897.5 36847.5 ;
      RECT  3032.5 36592.5 2897.5 36657.5 ;
      RECT  3872.5 36212.5 3737.5 36277.5 ;
      RECT  3872.5 36402.5 3737.5 36467.5 ;
      RECT  3872.5 36402.5 3737.5 36467.5 ;
      RECT  3872.5 36212.5 3737.5 36277.5 ;
      RECT  3872.5 36402.5 3737.5 36467.5 ;
      RECT  3872.5 36592.5 3737.5 36657.5 ;
      RECT  3872.5 36592.5 3737.5 36657.5 ;
      RECT  3872.5 36402.5 3737.5 36467.5 ;
      RECT  3872.5 36592.5 3737.5 36657.5 ;
      RECT  3872.5 36782.5 3737.5 36847.5 ;
      RECT  3872.5 36782.5 3737.5 36847.5 ;
      RECT  3872.5 36592.5 3737.5 36657.5 ;
      RECT  2942.5 36952.5 2807.5 37017.5 ;
      RECT  3917.5 36952.5 3782.5 37017.5 ;
      RECT  3660.0 36787.5 3595.0 36652.5 ;
      RECT  3520.0 36597.5 3455.0 36462.5 ;
      RECT  3380.0 36407.5 3315.0 36272.5 ;
      RECT  3032.5 36402.5 2897.5 36467.5 ;
      RECT  3032.5 36782.5 2897.5 36847.5 ;
      RECT  3872.5 36782.5 3737.5 36847.5 ;
      RECT  3415.0 36782.5 3280.0 36847.5 ;
      RECT  3380.0 36272.5 3315.0 36407.5 ;
      RECT  3520.0 36462.5 3455.0 36597.5 ;
      RECT  3660.0 36652.5 3595.0 36787.5 ;
      RECT  3415.0 36782.5 3280.0 36847.5 ;
      RECT  2722.5 36145.0 2657.5 37155.0 ;
      RECT  4067.5 36145.0 4002.5 37155.0 ;
      RECT  2875.0 37582.5 2690.0 37647.5 ;
      RECT  4035.0 37582.5 3850.0 37647.5 ;
      RECT  3917.5 37222.5 4067.5 37287.5 ;
      RECT  3032.5 37222.5 2657.5 37287.5 ;
      RECT  3917.5 37412.5 3032.5 37477.5 ;
      RECT  3032.5 37222.5 2897.5 37287.5 ;
      RECT  3032.5 37412.5 2897.5 37477.5 ;
      RECT  3032.5 37412.5 2897.5 37477.5 ;
      RECT  3032.5 37222.5 2897.5 37287.5 ;
      RECT  3917.5 37222.5 3782.5 37287.5 ;
      RECT  3917.5 37412.5 3782.5 37477.5 ;
      RECT  3917.5 37412.5 3782.5 37477.5 ;
      RECT  3917.5 37222.5 3782.5 37287.5 ;
      RECT  2942.5 37582.5 2807.5 37647.5 ;
      RECT  3917.5 37582.5 3782.5 37647.5 ;
      RECT  3475.0 37280.0 3340.0 37345.0 ;
      RECT  3475.0 37280.0 3340.0 37345.0 ;
      RECT  3440.0 37445.0 3375.0 37510.0 ;
      RECT  2722.5 37155.0 2657.5 37715.0 ;
      RECT  4067.5 37155.0 4002.5 37715.0 ;
      RECT  1462.5 36212.5 1312.5 36277.5 ;
      RECT  1462.5 36592.5 1312.5 36657.5 ;
      RECT  2280.0 36212.5 2722.5 36277.5 ;
      RECT  2505.0 36762.5 2690.0 36827.5 ;
      RECT  1345.0 36762.5 1530.0 36827.5 ;
      RECT  2280.0 36212.5 2415.0 36277.5 ;
      RECT  2280.0 36402.5 2415.0 36467.5 ;
      RECT  2280.0 36402.5 2415.0 36467.5 ;
      RECT  2280.0 36212.5 2415.0 36277.5 ;
      RECT  2280.0 36402.5 2415.0 36467.5 ;
      RECT  2280.0 36592.5 2415.0 36657.5 ;
      RECT  2280.0 36592.5 2415.0 36657.5 ;
      RECT  2280.0 36402.5 2415.0 36467.5 ;
      RECT  1462.5 36212.5 1597.5 36277.5 ;
      RECT  1462.5 36402.5 1597.5 36467.5 ;
      RECT  1462.5 36402.5 1597.5 36467.5 ;
      RECT  1462.5 36212.5 1597.5 36277.5 ;
      RECT  1462.5 36402.5 1597.5 36467.5 ;
      RECT  1462.5 36592.5 1597.5 36657.5 ;
      RECT  1462.5 36592.5 1597.5 36657.5 ;
      RECT  1462.5 36402.5 1597.5 36467.5 ;
      RECT  2437.5 36762.5 2572.5 36827.5 ;
      RECT  1462.5 36762.5 1597.5 36827.5 ;
      RECT  1682.5 36597.5 1747.5 36462.5 ;
      RECT  1897.5 36340.0 1962.5 36205.0 ;
      RECT  2280.0 36592.5 2415.0 36657.5 ;
      RECT  1497.5 36502.5 1562.5 36367.5 ;
      RECT  1897.5 36762.5 1962.5 36627.5 ;
      RECT  1897.5 36205.0 1962.5 36340.0 ;
      RECT  1682.5 36462.5 1747.5 36597.5 ;
      RECT  1897.5 36627.5 1962.5 36762.5 ;
      RECT  2657.5 36145.0 2722.5 37065.0 ;
      RECT  1312.5 36145.0 1377.5 37065.0 ;
      RECT  1507.5 37357.5 1312.5 37422.5 ;
      RECT  2347.5 37357.5 2722.5 37422.5 ;
      RECT  2347.5 37737.5 2722.5 37802.5 ;
      RECT  2505.0 37907.5 2690.0 37972.5 ;
      RECT  1345.0 37907.5 1530.0 37972.5 ;
      RECT  2347.5 37357.5 2482.5 37422.5 ;
      RECT  2347.5 37547.5 2482.5 37612.5 ;
      RECT  2347.5 37547.5 2482.5 37612.5 ;
      RECT  2347.5 37357.5 2482.5 37422.5 ;
      RECT  2347.5 37547.5 2482.5 37612.5 ;
      RECT  2347.5 37737.5 2482.5 37802.5 ;
      RECT  2347.5 37737.5 2482.5 37802.5 ;
      RECT  2347.5 37547.5 2482.5 37612.5 ;
      RECT  1507.5 37357.5 1642.5 37422.5 ;
      RECT  1507.5 37547.5 1642.5 37612.5 ;
      RECT  1507.5 37547.5 1642.5 37612.5 ;
      RECT  1507.5 37357.5 1642.5 37422.5 ;
      RECT  1507.5 37547.5 1642.5 37612.5 ;
      RECT  1507.5 37737.5 1642.5 37802.5 ;
      RECT  1507.5 37737.5 1642.5 37802.5 ;
      RECT  1507.5 37547.5 1642.5 37612.5 ;
      RECT  2437.5 37907.5 2572.5 37972.5 ;
      RECT  1462.5 37907.5 1597.5 37972.5 ;
      RECT  1737.5 37742.5 1802.5 37607.5 ;
      RECT  1952.5 37485.0 2017.5 37350.0 ;
      RECT  2347.5 37547.5 2482.5 37612.5 ;
      RECT  1507.5 37737.5 1642.5 37802.5 ;
      RECT  1952.5 37837.5 2017.5 37702.5 ;
      RECT  1952.5 37350.0 2017.5 37485.0 ;
      RECT  1737.5 37607.5 1802.5 37742.5 ;
      RECT  1952.5 37702.5 2017.5 37837.5 ;
      RECT  2657.5 37290.0 2722.5 38210.0 ;
      RECT  1312.5 37290.0 1377.5 38210.0 ;
      RECT  2505.0 38567.5 2690.0 38502.5 ;
      RECT  1345.0 38567.5 1530.0 38502.5 ;
      RECT  1462.5 38927.5 1312.5 38862.5 ;
      RECT  2347.5 38927.5 2722.5 38862.5 ;
      RECT  1462.5 38737.5 2347.5 38672.5 ;
      RECT  2347.5 38927.5 2482.5 38862.5 ;
      RECT  2347.5 38737.5 2482.5 38672.5 ;
      RECT  2347.5 38737.5 2482.5 38672.5 ;
      RECT  2347.5 38927.5 2482.5 38862.5 ;
      RECT  1462.5 38927.5 1597.5 38862.5 ;
      RECT  1462.5 38737.5 1597.5 38672.5 ;
      RECT  1462.5 38737.5 1597.5 38672.5 ;
      RECT  1462.5 38927.5 1597.5 38862.5 ;
      RECT  2437.5 38567.5 2572.5 38502.5 ;
      RECT  1462.5 38567.5 1597.5 38502.5 ;
      RECT  1905.0 38870.0 2040.0 38805.0 ;
      RECT  1905.0 38870.0 2040.0 38805.0 ;
      RECT  1940.0 38705.0 2005.0 38640.0 ;
      RECT  2657.5 38995.0 2722.5 38435.0 ;
      RECT  1312.5 38995.0 1377.5 38435.0 ;
      RECT  2505.0 39127.5 2690.0 39062.5 ;
      RECT  1345.0 39127.5 1530.0 39062.5 ;
      RECT  1462.5 39487.5 1312.5 39422.5 ;
      RECT  2347.5 39487.5 2722.5 39422.5 ;
      RECT  1462.5 39297.5 2347.5 39232.5 ;
      RECT  2347.5 39487.5 2482.5 39422.5 ;
      RECT  2347.5 39297.5 2482.5 39232.5 ;
      RECT  2347.5 39297.5 2482.5 39232.5 ;
      RECT  2347.5 39487.5 2482.5 39422.5 ;
      RECT  1462.5 39487.5 1597.5 39422.5 ;
      RECT  1462.5 39297.5 1597.5 39232.5 ;
      RECT  1462.5 39297.5 1597.5 39232.5 ;
      RECT  1462.5 39487.5 1597.5 39422.5 ;
      RECT  2437.5 39127.5 2572.5 39062.5 ;
      RECT  1462.5 39127.5 1597.5 39062.5 ;
      RECT  1905.0 39430.0 2040.0 39365.0 ;
      RECT  1905.0 39430.0 2040.0 39365.0 ;
      RECT  1940.0 39265.0 2005.0 39200.0 ;
      RECT  2657.5 39555.0 2722.5 38995.0 ;
      RECT  1312.5 39555.0 1377.5 38995.0 ;
      RECT  1182.5 36772.5 1377.5 36837.5 ;
      RECT  342.5 36772.5 -32.5 36837.5 ;
      RECT  342.5 37152.5 -32.5 37217.5 ;
      RECT  185.0 37512.5 8.881784197e-13 37577.5 ;
      RECT  1345.0 37512.5 1160.0 37577.5 ;
      RECT  342.5 36772.5 207.5 36837.5 ;
      RECT  342.5 36962.5 207.5 37027.5 ;
      RECT  342.5 36962.5 207.5 37027.5 ;
      RECT  342.5 36772.5 207.5 36837.5 ;
      RECT  342.5 36962.5 207.5 37027.5 ;
      RECT  342.5 37152.5 207.5 37217.5 ;
      RECT  342.5 37152.5 207.5 37217.5 ;
      RECT  342.5 36962.5 207.5 37027.5 ;
      RECT  342.5 37152.5 207.5 37217.5 ;
      RECT  342.5 37342.5 207.5 37407.5 ;
      RECT  342.5 37342.5 207.5 37407.5 ;
      RECT  342.5 37152.5 207.5 37217.5 ;
      RECT  1182.5 36772.5 1047.5 36837.5 ;
      RECT  1182.5 36962.5 1047.5 37027.5 ;
      RECT  1182.5 36962.5 1047.5 37027.5 ;
      RECT  1182.5 36772.5 1047.5 36837.5 ;
      RECT  1182.5 36962.5 1047.5 37027.5 ;
      RECT  1182.5 37152.5 1047.5 37217.5 ;
      RECT  1182.5 37152.5 1047.5 37217.5 ;
      RECT  1182.5 36962.5 1047.5 37027.5 ;
      RECT  1182.5 37152.5 1047.5 37217.5 ;
      RECT  1182.5 37342.5 1047.5 37407.5 ;
      RECT  1182.5 37342.5 1047.5 37407.5 ;
      RECT  1182.5 37152.5 1047.5 37217.5 ;
      RECT  252.5 37512.5 117.5 37577.5 ;
      RECT  1227.5 37512.5 1092.5 37577.5 ;
      RECT  970.0 37347.5 905.0 37212.5 ;
      RECT  830.0 37157.5 765.0 37022.5 ;
      RECT  690.0 36967.5 625.0 36832.5 ;
      RECT  342.5 36962.5 207.5 37027.5 ;
      RECT  342.5 37342.5 207.5 37407.5 ;
      RECT  1182.5 37342.5 1047.5 37407.5 ;
      RECT  725.0 37342.5 590.0 37407.5 ;
      RECT  690.0 36832.5 625.0 36967.5 ;
      RECT  830.0 37022.5 765.0 37157.5 ;
      RECT  970.0 37212.5 905.0 37347.5 ;
      RECT  725.0 37342.5 590.0 37407.5 ;
      RECT  32.5 36705.0 -32.5 37715.0 ;
      RECT  1377.5 36705.0 1312.5 37715.0 ;
      RECT  185.0 38142.5 8.881784197e-13 38207.5 ;
      RECT  1345.0 38142.5 1160.0 38207.5 ;
      RECT  1227.5 37782.5 1377.5 37847.5 ;
      RECT  342.5 37782.5 -32.5 37847.5 ;
      RECT  1227.5 37972.5 342.5 38037.5 ;
      RECT  342.5 37782.5 207.5 37847.5 ;
      RECT  342.5 37972.5 207.5 38037.5 ;
      RECT  342.5 37972.5 207.5 38037.5 ;
      RECT  342.5 37782.5 207.5 37847.5 ;
      RECT  1227.5 37782.5 1092.5 37847.5 ;
      RECT  1227.5 37972.5 1092.5 38037.5 ;
      RECT  1227.5 37972.5 1092.5 38037.5 ;
      RECT  1227.5 37782.5 1092.5 37847.5 ;
      RECT  252.5 38142.5 117.5 38207.5 ;
      RECT  1227.5 38142.5 1092.5 38207.5 ;
      RECT  785.0 37840.0 650.0 37905.0 ;
      RECT  785.0 37840.0 650.0 37905.0 ;
      RECT  750.0 38005.0 685.0 38070.0 ;
      RECT  32.5 37715.0 -32.5 38275.0 ;
      RECT  1377.5 37715.0 1312.5 38275.0 ;
      RECT  185.0 38702.5 8.881784197e-13 38767.5 ;
      RECT  1345.0 38702.5 1160.0 38767.5 ;
      RECT  1227.5 38342.5 1377.5 38407.5 ;
      RECT  342.5 38342.5 -32.5 38407.5 ;
      RECT  1227.5 38532.5 342.5 38597.5 ;
      RECT  342.5 38342.5 207.5 38407.5 ;
      RECT  342.5 38532.5 207.5 38597.5 ;
      RECT  342.5 38532.5 207.5 38597.5 ;
      RECT  342.5 38342.5 207.5 38407.5 ;
      RECT  1227.5 38342.5 1092.5 38407.5 ;
      RECT  1227.5 38532.5 1092.5 38597.5 ;
      RECT  1227.5 38532.5 1092.5 38597.5 ;
      RECT  1227.5 38342.5 1092.5 38407.5 ;
      RECT  252.5 38702.5 117.5 38767.5 ;
      RECT  1227.5 38702.5 1092.5 38767.5 ;
      RECT  785.0 38400.0 650.0 38465.0 ;
      RECT  785.0 38400.0 650.0 38465.0 ;
      RECT  750.0 38565.0 685.0 38630.0 ;
      RECT  32.5 38275.0 -32.5 38835.0 ;
      RECT  1377.5 38275.0 1312.5 38835.0 ;
      RECT  185.0 39262.5 8.881784197e-13 39327.5 ;
      RECT  1345.0 39262.5 1160.0 39327.5 ;
      RECT  1227.5 38902.5 1377.5 38967.5 ;
      RECT  342.5 38902.5 -32.5 38967.5 ;
      RECT  1227.5 39092.5 342.5 39157.5 ;
      RECT  342.5 38902.5 207.5 38967.5 ;
      RECT  342.5 39092.5 207.5 39157.5 ;
      RECT  342.5 39092.5 207.5 39157.5 ;
      RECT  342.5 38902.5 207.5 38967.5 ;
      RECT  1227.5 38902.5 1092.5 38967.5 ;
      RECT  1227.5 39092.5 1092.5 39157.5 ;
      RECT  1227.5 39092.5 1092.5 39157.5 ;
      RECT  1227.5 38902.5 1092.5 38967.5 ;
      RECT  252.5 39262.5 117.5 39327.5 ;
      RECT  1227.5 39262.5 1092.5 39327.5 ;
      RECT  785.0 38960.0 650.0 39025.0 ;
      RECT  785.0 38960.0 650.0 39025.0 ;
      RECT  750.0 39125.0 685.0 39190.0 ;
      RECT  32.5 38835.0 -32.5 39395.0 ;
      RECT  1377.5 38835.0 1312.5 39395.0 ;
      RECT  1377.5 52037.5 1312.5 47865.0 ;
      RECT  1312.5 42127.5 1025.0 42192.5 ;
      RECT  1312.5 44537.5 1025.0 44602.5 ;
      RECT  1312.5 44817.5 1025.0 44882.5 ;
      RECT  1312.5 47227.5 1025.0 47292.5 ;
      RECT  1377.5 40082.5 935.0 40147.5 ;
      RECT  935.0 40082.5 230.0 40147.5 ;
      RECT  20.0 43332.5 935.0 43397.5 ;
      RECT  20.0 46022.5 935.0 46087.5 ;
      RECT  20.0 40642.5 935.0 40707.5 ;
      RECT  2005.0 41655.0 1940.0 42355.0 ;
      RECT  2005.0 41847.5 1940.0 41912.5 ;
      RECT  2005.0 41655.0 1940.0 41880.0 ;
      RECT  1972.5 41847.5 1025.0 41912.5 ;
      RECT  2690.0 41717.5 2465.0 41782.5 ;
      RECT  2430.0 40847.5 2365.0 40912.5 ;
      RECT  2005.0 40847.5 1940.0 40912.5 ;
      RECT  2430.0 40880.0 2365.0 41527.5 ;
      RECT  2397.5 40847.5 1972.5 40912.5 ;
      RECT  2005.0 40550.0 1940.0 40880.0 ;
      RECT  1972.5 40847.5 1172.5 40912.5 ;
      RECT  1172.5 40250.0 750.0 40315.0 ;
      RECT  2040.0 40485.0 1905.0 40550.0 ;
      RECT  2005.0 42355.0 1940.0 42560.0 ;
      RECT  2505.0 40247.5 2690.0 40182.5 ;
      RECT  1345.0 40247.5 1530.0 40182.5 ;
      RECT  1462.5 40607.5 1312.5 40542.5 ;
      RECT  2347.5 40607.5 2722.5 40542.5 ;
      RECT  1462.5 40417.5 2347.5 40352.5 ;
      RECT  2347.5 40607.5 2482.5 40542.5 ;
      RECT  2347.5 40417.5 2482.5 40352.5 ;
      RECT  2347.5 40417.5 2482.5 40352.5 ;
      RECT  2347.5 40607.5 2482.5 40542.5 ;
      RECT  1462.5 40607.5 1597.5 40542.5 ;
      RECT  1462.5 40417.5 1597.5 40352.5 ;
      RECT  1462.5 40417.5 1597.5 40352.5 ;
      RECT  1462.5 40607.5 1597.5 40542.5 ;
      RECT  2437.5 40247.5 2572.5 40182.5 ;
      RECT  1462.5 40247.5 1597.5 40182.5 ;
      RECT  1905.0 40550.0 2040.0 40485.0 ;
      RECT  1905.0 40550.0 2040.0 40485.0 ;
      RECT  1940.0 40385.0 2005.0 40320.0 ;
      RECT  2657.5 40675.0 2722.5 40115.0 ;
      RECT  1312.5 40675.0 1377.5 40115.0 ;
      RECT  2330.0 41527.5 2465.0 41592.5 ;
      RECT  2330.0 41717.5 2465.0 41782.5 ;
      RECT  2330.0 41717.5 2465.0 41782.5 ;
      RECT  2330.0 41527.5 2465.0 41592.5 ;
      RECT  1312.5 51972.5 1377.5 52037.5 ;
      RECT  4002.5 51972.5 4067.5 52037.5 ;
      RECT  1312.5 51875.0 1377.5 52005.0 ;
      RECT  1345.0 51972.5 4035.0 52037.5 ;
      RECT  4002.5 51875.0 4067.5 52005.0 ;
      RECT  2875.0 42782.5 2690.0 42847.5 ;
      RECT  4035.0 42782.5 3850.0 42847.5 ;
      RECT  3917.5 42422.5 4067.5 42487.5 ;
      RECT  3032.5 42422.5 2657.5 42487.5 ;
      RECT  3917.5 42612.5 3032.5 42677.5 ;
      RECT  3032.5 42422.5 2897.5 42487.5 ;
      RECT  3032.5 42612.5 2897.5 42677.5 ;
      RECT  3032.5 42612.5 2897.5 42677.5 ;
      RECT  3032.5 42422.5 2897.5 42487.5 ;
      RECT  3917.5 42422.5 3782.5 42487.5 ;
      RECT  3917.5 42612.5 3782.5 42677.5 ;
      RECT  3917.5 42612.5 3782.5 42677.5 ;
      RECT  3917.5 42422.5 3782.5 42487.5 ;
      RECT  2942.5 42782.5 2807.5 42847.5 ;
      RECT  3917.5 42782.5 3782.5 42847.5 ;
      RECT  3475.0 42480.0 3340.0 42545.0 ;
      RECT  3475.0 42480.0 3340.0 42545.0 ;
      RECT  3440.0 42645.0 3375.0 42710.0 ;
      RECT  2722.5 42355.0 2657.5 42915.0 ;
      RECT  4067.5 42355.0 4002.5 42915.0 ;
      RECT  2875.0 43342.5 2690.0 43407.5 ;
      RECT  4035.0 43342.5 3850.0 43407.5 ;
      RECT  3917.5 42982.5 4067.5 43047.5 ;
      RECT  3032.5 42982.5 2657.5 43047.5 ;
      RECT  3917.5 43172.5 3032.5 43237.5 ;
      RECT  3032.5 42982.5 2897.5 43047.5 ;
      RECT  3032.5 43172.5 2897.5 43237.5 ;
      RECT  3032.5 43172.5 2897.5 43237.5 ;
      RECT  3032.5 42982.5 2897.5 43047.5 ;
      RECT  3917.5 42982.5 3782.5 43047.5 ;
      RECT  3917.5 43172.5 3782.5 43237.5 ;
      RECT  3917.5 43172.5 3782.5 43237.5 ;
      RECT  3917.5 42982.5 3782.5 43047.5 ;
      RECT  2942.5 43342.5 2807.5 43407.5 ;
      RECT  3917.5 43342.5 3782.5 43407.5 ;
      RECT  3475.0 43040.0 3340.0 43105.0 ;
      RECT  3475.0 43040.0 3340.0 43105.0 ;
      RECT  3440.0 43205.0 3375.0 43270.0 ;
      RECT  2722.5 42915.0 2657.5 43475.0 ;
      RECT  4067.5 42915.0 4002.5 43475.0 ;
      RECT  3340.0 43040.0 3475.0 43105.0 ;
      RECT  2875.0 43902.5 2690.0 43967.5 ;
      RECT  4035.0 43902.5 3850.0 43967.5 ;
      RECT  3917.5 43542.5 4067.5 43607.5 ;
      RECT  3032.5 43542.5 2657.5 43607.5 ;
      RECT  3917.5 43732.5 3032.5 43797.5 ;
      RECT  3032.5 43542.5 2897.5 43607.5 ;
      RECT  3032.5 43732.5 2897.5 43797.5 ;
      RECT  3032.5 43732.5 2897.5 43797.5 ;
      RECT  3032.5 43542.5 2897.5 43607.5 ;
      RECT  3917.5 43542.5 3782.5 43607.5 ;
      RECT  3917.5 43732.5 3782.5 43797.5 ;
      RECT  3917.5 43732.5 3782.5 43797.5 ;
      RECT  3917.5 43542.5 3782.5 43607.5 ;
      RECT  2942.5 43902.5 2807.5 43967.5 ;
      RECT  3917.5 43902.5 3782.5 43967.5 ;
      RECT  3475.0 43600.0 3340.0 43665.0 ;
      RECT  3475.0 43600.0 3340.0 43665.0 ;
      RECT  3440.0 43765.0 3375.0 43830.0 ;
      RECT  2722.5 43475.0 2657.5 44035.0 ;
      RECT  4067.5 43475.0 4002.5 44035.0 ;
      RECT  3340.0 43600.0 3475.0 43665.0 ;
      RECT  2875.0 44462.5 2690.0 44527.5 ;
      RECT  4035.0 44462.5 3850.0 44527.5 ;
      RECT  3917.5 44102.5 4067.5 44167.5 ;
      RECT  3032.5 44102.5 2657.5 44167.5 ;
      RECT  3917.5 44292.5 3032.5 44357.5 ;
      RECT  3032.5 44102.5 2897.5 44167.5 ;
      RECT  3032.5 44292.5 2897.5 44357.5 ;
      RECT  3032.5 44292.5 2897.5 44357.5 ;
      RECT  3032.5 44102.5 2897.5 44167.5 ;
      RECT  3917.5 44102.5 3782.5 44167.5 ;
      RECT  3917.5 44292.5 3782.5 44357.5 ;
      RECT  3917.5 44292.5 3782.5 44357.5 ;
      RECT  3917.5 44102.5 3782.5 44167.5 ;
      RECT  2942.5 44462.5 2807.5 44527.5 ;
      RECT  3917.5 44462.5 3782.5 44527.5 ;
      RECT  3475.0 44160.0 3340.0 44225.0 ;
      RECT  3475.0 44160.0 3340.0 44225.0 ;
      RECT  3440.0 44325.0 3375.0 44390.0 ;
      RECT  2722.5 44035.0 2657.5 44595.0 ;
      RECT  4067.5 44035.0 4002.5 44595.0 ;
      RECT  3340.0 44160.0 3475.0 44225.0 ;
      RECT  2875.0 45022.5 2690.0 45087.5 ;
      RECT  4035.0 45022.5 3850.0 45087.5 ;
      RECT  3917.5 44662.5 4067.5 44727.5 ;
      RECT  3032.5 44662.5 2657.5 44727.5 ;
      RECT  3917.5 44852.5 3032.5 44917.5 ;
      RECT  3032.5 44662.5 2897.5 44727.5 ;
      RECT  3032.5 44852.5 2897.5 44917.5 ;
      RECT  3032.5 44852.5 2897.5 44917.5 ;
      RECT  3032.5 44662.5 2897.5 44727.5 ;
      RECT  3917.5 44662.5 3782.5 44727.5 ;
      RECT  3917.5 44852.5 3782.5 44917.5 ;
      RECT  3917.5 44852.5 3782.5 44917.5 ;
      RECT  3917.5 44662.5 3782.5 44727.5 ;
      RECT  2942.5 45022.5 2807.5 45087.5 ;
      RECT  3917.5 45022.5 3782.5 45087.5 ;
      RECT  3475.0 44720.0 3340.0 44785.0 ;
      RECT  3475.0 44720.0 3340.0 44785.0 ;
      RECT  3440.0 44885.0 3375.0 44950.0 ;
      RECT  2722.5 44595.0 2657.5 45155.0 ;
      RECT  4067.5 44595.0 4002.5 45155.0 ;
      RECT  3340.0 44720.0 3475.0 44785.0 ;
      RECT  2875.0 45582.5 2690.0 45647.5 ;
      RECT  4035.0 45582.5 3850.0 45647.5 ;
      RECT  3917.5 45222.5 4067.5 45287.5 ;
      RECT  3032.5 45222.5 2657.5 45287.5 ;
      RECT  3917.5 45412.5 3032.5 45477.5 ;
      RECT  3032.5 45222.5 2897.5 45287.5 ;
      RECT  3032.5 45412.5 2897.5 45477.5 ;
      RECT  3032.5 45412.5 2897.5 45477.5 ;
      RECT  3032.5 45222.5 2897.5 45287.5 ;
      RECT  3917.5 45222.5 3782.5 45287.5 ;
      RECT  3917.5 45412.5 3782.5 45477.5 ;
      RECT  3917.5 45412.5 3782.5 45477.5 ;
      RECT  3917.5 45222.5 3782.5 45287.5 ;
      RECT  2942.5 45582.5 2807.5 45647.5 ;
      RECT  3917.5 45582.5 3782.5 45647.5 ;
      RECT  3475.0 45280.0 3340.0 45345.0 ;
      RECT  3475.0 45280.0 3340.0 45345.0 ;
      RECT  3440.0 45445.0 3375.0 45510.0 ;
      RECT  2722.5 45155.0 2657.5 45715.0 ;
      RECT  4067.5 45155.0 4002.5 45715.0 ;
      RECT  3340.0 45280.0 3475.0 45345.0 ;
      RECT  2875.0 46142.5 2690.0 46207.5 ;
      RECT  4035.0 46142.5 3850.0 46207.5 ;
      RECT  3917.5 45782.5 4067.5 45847.5 ;
      RECT  3032.5 45782.5 2657.5 45847.5 ;
      RECT  3917.5 45972.5 3032.5 46037.5 ;
      RECT  3032.5 45782.5 2897.5 45847.5 ;
      RECT  3032.5 45972.5 2897.5 46037.5 ;
      RECT  3032.5 45972.5 2897.5 46037.5 ;
      RECT  3032.5 45782.5 2897.5 45847.5 ;
      RECT  3917.5 45782.5 3782.5 45847.5 ;
      RECT  3917.5 45972.5 3782.5 46037.5 ;
      RECT  3917.5 45972.5 3782.5 46037.5 ;
      RECT  3917.5 45782.5 3782.5 45847.5 ;
      RECT  2942.5 46142.5 2807.5 46207.5 ;
      RECT  3917.5 46142.5 3782.5 46207.5 ;
      RECT  3475.0 45840.0 3340.0 45905.0 ;
      RECT  3475.0 45840.0 3340.0 45905.0 ;
      RECT  3440.0 46005.0 3375.0 46070.0 ;
      RECT  2722.5 45715.0 2657.5 46275.0 ;
      RECT  4067.5 45715.0 4002.5 46275.0 ;
      RECT  3340.0 45840.0 3475.0 45905.0 ;
      RECT  2875.0 46702.5 2690.0 46767.5 ;
      RECT  4035.0 46702.5 3850.0 46767.5 ;
      RECT  3917.5 46342.5 4067.5 46407.5 ;
      RECT  3032.5 46342.5 2657.5 46407.5 ;
      RECT  3917.5 46532.5 3032.5 46597.5 ;
      RECT  3032.5 46342.5 2897.5 46407.5 ;
      RECT  3032.5 46532.5 2897.5 46597.5 ;
      RECT  3032.5 46532.5 2897.5 46597.5 ;
      RECT  3032.5 46342.5 2897.5 46407.5 ;
      RECT  3917.5 46342.5 3782.5 46407.5 ;
      RECT  3917.5 46532.5 3782.5 46597.5 ;
      RECT  3917.5 46532.5 3782.5 46597.5 ;
      RECT  3917.5 46342.5 3782.5 46407.5 ;
      RECT  2942.5 46702.5 2807.5 46767.5 ;
      RECT  3917.5 46702.5 3782.5 46767.5 ;
      RECT  3475.0 46400.0 3340.0 46465.0 ;
      RECT  3475.0 46400.0 3340.0 46465.0 ;
      RECT  3440.0 46565.0 3375.0 46630.0 ;
      RECT  2722.5 46275.0 2657.5 46835.0 ;
      RECT  4067.5 46275.0 4002.5 46835.0 ;
      RECT  3340.0 46400.0 3475.0 46465.0 ;
      RECT  2875.0 47262.5 2690.0 47327.5 ;
      RECT  4035.0 47262.5 3850.0 47327.5 ;
      RECT  3917.5 46902.5 4067.5 46967.5 ;
      RECT  3032.5 46902.5 2657.5 46967.5 ;
      RECT  3917.5 47092.5 3032.5 47157.5 ;
      RECT  3032.5 46902.5 2897.5 46967.5 ;
      RECT  3032.5 47092.5 2897.5 47157.5 ;
      RECT  3032.5 47092.5 2897.5 47157.5 ;
      RECT  3032.5 46902.5 2897.5 46967.5 ;
      RECT  3917.5 46902.5 3782.5 46967.5 ;
      RECT  3917.5 47092.5 3782.5 47157.5 ;
      RECT  3917.5 47092.5 3782.5 47157.5 ;
      RECT  3917.5 46902.5 3782.5 46967.5 ;
      RECT  2942.5 47262.5 2807.5 47327.5 ;
      RECT  3917.5 47262.5 3782.5 47327.5 ;
      RECT  3475.0 46960.0 3340.0 47025.0 ;
      RECT  3475.0 46960.0 3340.0 47025.0 ;
      RECT  3440.0 47125.0 3375.0 47190.0 ;
      RECT  2722.5 46835.0 2657.5 47395.0 ;
      RECT  4067.5 46835.0 4002.5 47395.0 ;
      RECT  3340.0 46960.0 3475.0 47025.0 ;
      RECT  2875.0 47822.5 2690.0 47887.5 ;
      RECT  4035.0 47822.5 3850.0 47887.5 ;
      RECT  3917.5 47462.5 4067.5 47527.5 ;
      RECT  3032.5 47462.5 2657.5 47527.5 ;
      RECT  3917.5 47652.5 3032.5 47717.5 ;
      RECT  3032.5 47462.5 2897.5 47527.5 ;
      RECT  3032.5 47652.5 2897.5 47717.5 ;
      RECT  3032.5 47652.5 2897.5 47717.5 ;
      RECT  3032.5 47462.5 2897.5 47527.5 ;
      RECT  3917.5 47462.5 3782.5 47527.5 ;
      RECT  3917.5 47652.5 3782.5 47717.5 ;
      RECT  3917.5 47652.5 3782.5 47717.5 ;
      RECT  3917.5 47462.5 3782.5 47527.5 ;
      RECT  2942.5 47822.5 2807.5 47887.5 ;
      RECT  3917.5 47822.5 3782.5 47887.5 ;
      RECT  3475.0 47520.0 3340.0 47585.0 ;
      RECT  3475.0 47520.0 3340.0 47585.0 ;
      RECT  3440.0 47685.0 3375.0 47750.0 ;
      RECT  2722.5 47395.0 2657.5 47955.0 ;
      RECT  4067.5 47395.0 4002.5 47955.0 ;
      RECT  3340.0 47520.0 3475.0 47585.0 ;
      RECT  2875.0 48382.5 2690.0 48447.5 ;
      RECT  4035.0 48382.5 3850.0 48447.5 ;
      RECT  3917.5 48022.5 4067.5 48087.5 ;
      RECT  3032.5 48022.5 2657.5 48087.5 ;
      RECT  3917.5 48212.5 3032.5 48277.5 ;
      RECT  3032.5 48022.5 2897.5 48087.5 ;
      RECT  3032.5 48212.5 2897.5 48277.5 ;
      RECT  3032.5 48212.5 2897.5 48277.5 ;
      RECT  3032.5 48022.5 2897.5 48087.5 ;
      RECT  3917.5 48022.5 3782.5 48087.5 ;
      RECT  3917.5 48212.5 3782.5 48277.5 ;
      RECT  3917.5 48212.5 3782.5 48277.5 ;
      RECT  3917.5 48022.5 3782.5 48087.5 ;
      RECT  2942.5 48382.5 2807.5 48447.5 ;
      RECT  3917.5 48382.5 3782.5 48447.5 ;
      RECT  3475.0 48080.0 3340.0 48145.0 ;
      RECT  3475.0 48080.0 3340.0 48145.0 ;
      RECT  3440.0 48245.0 3375.0 48310.0 ;
      RECT  2722.5 47955.0 2657.5 48515.0 ;
      RECT  4067.5 47955.0 4002.5 48515.0 ;
      RECT  3340.0 48080.0 3475.0 48145.0 ;
      RECT  2875.0 48942.5 2690.0 49007.5 ;
      RECT  4035.0 48942.5 3850.0 49007.5 ;
      RECT  3917.5 48582.5 4067.5 48647.5 ;
      RECT  3032.5 48582.5 2657.5 48647.5 ;
      RECT  3917.5 48772.5 3032.5 48837.5 ;
      RECT  3032.5 48582.5 2897.5 48647.5 ;
      RECT  3032.5 48772.5 2897.5 48837.5 ;
      RECT  3032.5 48772.5 2897.5 48837.5 ;
      RECT  3032.5 48582.5 2897.5 48647.5 ;
      RECT  3917.5 48582.5 3782.5 48647.5 ;
      RECT  3917.5 48772.5 3782.5 48837.5 ;
      RECT  3917.5 48772.5 3782.5 48837.5 ;
      RECT  3917.5 48582.5 3782.5 48647.5 ;
      RECT  2942.5 48942.5 2807.5 49007.5 ;
      RECT  3917.5 48942.5 3782.5 49007.5 ;
      RECT  3475.0 48640.0 3340.0 48705.0 ;
      RECT  3475.0 48640.0 3340.0 48705.0 ;
      RECT  3440.0 48805.0 3375.0 48870.0 ;
      RECT  2722.5 48515.0 2657.5 49075.0 ;
      RECT  4067.5 48515.0 4002.5 49075.0 ;
      RECT  3340.0 48640.0 3475.0 48705.0 ;
      RECT  2875.0 49502.5 2690.0 49567.5 ;
      RECT  4035.0 49502.5 3850.0 49567.5 ;
      RECT  3917.5 49142.5 4067.5 49207.5 ;
      RECT  3032.5 49142.5 2657.5 49207.5 ;
      RECT  3917.5 49332.5 3032.5 49397.5 ;
      RECT  3032.5 49142.5 2897.5 49207.5 ;
      RECT  3032.5 49332.5 2897.5 49397.5 ;
      RECT  3032.5 49332.5 2897.5 49397.5 ;
      RECT  3032.5 49142.5 2897.5 49207.5 ;
      RECT  3917.5 49142.5 3782.5 49207.5 ;
      RECT  3917.5 49332.5 3782.5 49397.5 ;
      RECT  3917.5 49332.5 3782.5 49397.5 ;
      RECT  3917.5 49142.5 3782.5 49207.5 ;
      RECT  2942.5 49502.5 2807.5 49567.5 ;
      RECT  3917.5 49502.5 3782.5 49567.5 ;
      RECT  3475.0 49200.0 3340.0 49265.0 ;
      RECT  3475.0 49200.0 3340.0 49265.0 ;
      RECT  3440.0 49365.0 3375.0 49430.0 ;
      RECT  2722.5 49075.0 2657.5 49635.0 ;
      RECT  4067.5 49075.0 4002.5 49635.0 ;
      RECT  3340.0 49200.0 3475.0 49265.0 ;
      RECT  2875.0 50062.5 2690.0 50127.5 ;
      RECT  4035.0 50062.5 3850.0 50127.5 ;
      RECT  3917.5 49702.5 4067.5 49767.5 ;
      RECT  3032.5 49702.5 2657.5 49767.5 ;
      RECT  3917.5 49892.5 3032.5 49957.5 ;
      RECT  3032.5 49702.5 2897.5 49767.5 ;
      RECT  3032.5 49892.5 2897.5 49957.5 ;
      RECT  3032.5 49892.5 2897.5 49957.5 ;
      RECT  3032.5 49702.5 2897.5 49767.5 ;
      RECT  3917.5 49702.5 3782.5 49767.5 ;
      RECT  3917.5 49892.5 3782.5 49957.5 ;
      RECT  3917.5 49892.5 3782.5 49957.5 ;
      RECT  3917.5 49702.5 3782.5 49767.5 ;
      RECT  2942.5 50062.5 2807.5 50127.5 ;
      RECT  3917.5 50062.5 3782.5 50127.5 ;
      RECT  3475.0 49760.0 3340.0 49825.0 ;
      RECT  3475.0 49760.0 3340.0 49825.0 ;
      RECT  3440.0 49925.0 3375.0 49990.0 ;
      RECT  2722.5 49635.0 2657.5 50195.0 ;
      RECT  4067.5 49635.0 4002.5 50195.0 ;
      RECT  3340.0 49760.0 3475.0 49825.0 ;
      RECT  2875.0 50622.5 2690.0 50687.5 ;
      RECT  4035.0 50622.5 3850.0 50687.5 ;
      RECT  3917.5 50262.5 4067.5 50327.5 ;
      RECT  3032.5 50262.5 2657.5 50327.5 ;
      RECT  3917.5 50452.5 3032.5 50517.5 ;
      RECT  3032.5 50262.5 2897.5 50327.5 ;
      RECT  3032.5 50452.5 2897.5 50517.5 ;
      RECT  3032.5 50452.5 2897.5 50517.5 ;
      RECT  3032.5 50262.5 2897.5 50327.5 ;
      RECT  3917.5 50262.5 3782.5 50327.5 ;
      RECT  3917.5 50452.5 3782.5 50517.5 ;
      RECT  3917.5 50452.5 3782.5 50517.5 ;
      RECT  3917.5 50262.5 3782.5 50327.5 ;
      RECT  2942.5 50622.5 2807.5 50687.5 ;
      RECT  3917.5 50622.5 3782.5 50687.5 ;
      RECT  3475.0 50320.0 3340.0 50385.0 ;
      RECT  3475.0 50320.0 3340.0 50385.0 ;
      RECT  3440.0 50485.0 3375.0 50550.0 ;
      RECT  2722.5 50195.0 2657.5 50755.0 ;
      RECT  4067.5 50195.0 4002.5 50755.0 ;
      RECT  3340.0 50320.0 3475.0 50385.0 ;
      RECT  2875.0 51182.5 2690.0 51247.5 ;
      RECT  4035.0 51182.5 3850.0 51247.5 ;
      RECT  3917.5 50822.5 4067.5 50887.5 ;
      RECT  3032.5 50822.5 2657.5 50887.5 ;
      RECT  3917.5 51012.5 3032.5 51077.5 ;
      RECT  3032.5 50822.5 2897.5 50887.5 ;
      RECT  3032.5 51012.5 2897.5 51077.5 ;
      RECT  3032.5 51012.5 2897.5 51077.5 ;
      RECT  3032.5 50822.5 2897.5 50887.5 ;
      RECT  3917.5 50822.5 3782.5 50887.5 ;
      RECT  3917.5 51012.5 3782.5 51077.5 ;
      RECT  3917.5 51012.5 3782.5 51077.5 ;
      RECT  3917.5 50822.5 3782.5 50887.5 ;
      RECT  2942.5 51182.5 2807.5 51247.5 ;
      RECT  3917.5 51182.5 3782.5 51247.5 ;
      RECT  3475.0 50880.0 3340.0 50945.0 ;
      RECT  3475.0 50880.0 3340.0 50945.0 ;
      RECT  3440.0 51045.0 3375.0 51110.0 ;
      RECT  2722.5 50755.0 2657.5 51315.0 ;
      RECT  4067.5 50755.0 4002.5 51315.0 ;
      RECT  3340.0 50880.0 3475.0 50945.0 ;
      RECT  2875.0 51742.5 2690.0 51807.5 ;
      RECT  4035.0 51742.5 3850.0 51807.5 ;
      RECT  3917.5 51382.5 4067.5 51447.5 ;
      RECT  3032.5 51382.5 2657.5 51447.5 ;
      RECT  3917.5 51572.5 3032.5 51637.5 ;
      RECT  3032.5 51382.5 2897.5 51447.5 ;
      RECT  3032.5 51572.5 2897.5 51637.5 ;
      RECT  3032.5 51572.5 2897.5 51637.5 ;
      RECT  3032.5 51382.5 2897.5 51447.5 ;
      RECT  3917.5 51382.5 3782.5 51447.5 ;
      RECT  3917.5 51572.5 3782.5 51637.5 ;
      RECT  3917.5 51572.5 3782.5 51637.5 ;
      RECT  3917.5 51382.5 3782.5 51447.5 ;
      RECT  2942.5 51742.5 2807.5 51807.5 ;
      RECT  3917.5 51742.5 3782.5 51807.5 ;
      RECT  3475.0 51440.0 3340.0 51505.0 ;
      RECT  3475.0 51440.0 3340.0 51505.0 ;
      RECT  3440.0 51605.0 3375.0 51670.0 ;
      RECT  2722.5 51315.0 2657.5 51875.0 ;
      RECT  4067.5 51315.0 4002.5 51875.0 ;
      RECT  3340.0 51440.0 3475.0 51505.0 ;
      RECT  2505.0 50887.5 2690.0 50822.5 ;
      RECT  1345.0 50887.5 1530.0 50822.5 ;
      RECT  1462.5 51247.5 1312.5 51182.5 ;
      RECT  2347.5 51247.5 2722.5 51182.5 ;
      RECT  1462.5 51057.5 2347.5 50992.5 ;
      RECT  2347.5 51247.5 2482.5 51182.5 ;
      RECT  2347.5 51057.5 2482.5 50992.5 ;
      RECT  2347.5 51057.5 2482.5 50992.5 ;
      RECT  2347.5 51247.5 2482.5 51182.5 ;
      RECT  1462.5 51247.5 1597.5 51182.5 ;
      RECT  1462.5 51057.5 1597.5 50992.5 ;
      RECT  1462.5 51057.5 1597.5 50992.5 ;
      RECT  1462.5 51247.5 1597.5 51182.5 ;
      RECT  2437.5 50887.5 2572.5 50822.5 ;
      RECT  1462.5 50887.5 1597.5 50822.5 ;
      RECT  1905.0 51190.0 2040.0 51125.0 ;
      RECT  1905.0 51190.0 2040.0 51125.0 ;
      RECT  1940.0 51025.0 2005.0 50960.0 ;
      RECT  2657.5 51315.0 2722.5 50755.0 ;
      RECT  1312.5 51315.0 1377.5 50755.0 ;
      RECT  1905.0 51125.0 2040.0 51190.0 ;
      RECT  2505.0 50327.5 2690.0 50262.5 ;
      RECT  1345.0 50327.5 1530.0 50262.5 ;
      RECT  1462.5 50687.5 1312.5 50622.5 ;
      RECT  2347.5 50687.5 2722.5 50622.5 ;
      RECT  1462.5 50497.5 2347.5 50432.5 ;
      RECT  2347.5 50687.5 2482.5 50622.5 ;
      RECT  2347.5 50497.5 2482.5 50432.5 ;
      RECT  2347.5 50497.5 2482.5 50432.5 ;
      RECT  2347.5 50687.5 2482.5 50622.5 ;
      RECT  1462.5 50687.5 1597.5 50622.5 ;
      RECT  1462.5 50497.5 1597.5 50432.5 ;
      RECT  1462.5 50497.5 1597.5 50432.5 ;
      RECT  1462.5 50687.5 1597.5 50622.5 ;
      RECT  2437.5 50327.5 2572.5 50262.5 ;
      RECT  1462.5 50327.5 1597.5 50262.5 ;
      RECT  1905.0 50630.0 2040.0 50565.0 ;
      RECT  1905.0 50630.0 2040.0 50565.0 ;
      RECT  1940.0 50465.0 2005.0 50400.0 ;
      RECT  2657.5 50755.0 2722.5 50195.0 ;
      RECT  1312.5 50755.0 1377.5 50195.0 ;
      RECT  1905.0 50565.0 2040.0 50630.0 ;
      RECT  2505.0 49767.5 2690.0 49702.5 ;
      RECT  1345.0 49767.5 1530.0 49702.5 ;
      RECT  1462.5 50127.5 1312.5 50062.5 ;
      RECT  2347.5 50127.5 2722.5 50062.5 ;
      RECT  1462.5 49937.5 2347.5 49872.5 ;
      RECT  2347.5 50127.5 2482.5 50062.5 ;
      RECT  2347.5 49937.5 2482.5 49872.5 ;
      RECT  2347.5 49937.5 2482.5 49872.5 ;
      RECT  2347.5 50127.5 2482.5 50062.5 ;
      RECT  1462.5 50127.5 1597.5 50062.5 ;
      RECT  1462.5 49937.5 1597.5 49872.5 ;
      RECT  1462.5 49937.5 1597.5 49872.5 ;
      RECT  1462.5 50127.5 1597.5 50062.5 ;
      RECT  2437.5 49767.5 2572.5 49702.5 ;
      RECT  1462.5 49767.5 1597.5 49702.5 ;
      RECT  1905.0 50070.0 2040.0 50005.0 ;
      RECT  1905.0 50070.0 2040.0 50005.0 ;
      RECT  1940.0 49905.0 2005.0 49840.0 ;
      RECT  2657.5 50195.0 2722.5 49635.0 ;
      RECT  1312.5 50195.0 1377.5 49635.0 ;
      RECT  1905.0 50005.0 2040.0 50070.0 ;
      RECT  2505.0 49207.5 2690.0 49142.5 ;
      RECT  1345.0 49207.5 1530.0 49142.5 ;
      RECT  1462.5 49567.5 1312.5 49502.5 ;
      RECT  2347.5 49567.5 2722.5 49502.5 ;
      RECT  1462.5 49377.5 2347.5 49312.5 ;
      RECT  2347.5 49567.5 2482.5 49502.5 ;
      RECT  2347.5 49377.5 2482.5 49312.5 ;
      RECT  2347.5 49377.5 2482.5 49312.5 ;
      RECT  2347.5 49567.5 2482.5 49502.5 ;
      RECT  1462.5 49567.5 1597.5 49502.5 ;
      RECT  1462.5 49377.5 1597.5 49312.5 ;
      RECT  1462.5 49377.5 1597.5 49312.5 ;
      RECT  1462.5 49567.5 1597.5 49502.5 ;
      RECT  2437.5 49207.5 2572.5 49142.5 ;
      RECT  1462.5 49207.5 1597.5 49142.5 ;
      RECT  1905.0 49510.0 2040.0 49445.0 ;
      RECT  1905.0 49510.0 2040.0 49445.0 ;
      RECT  1940.0 49345.0 2005.0 49280.0 ;
      RECT  2657.5 49635.0 2722.5 49075.0 ;
      RECT  1312.5 49635.0 1377.5 49075.0 ;
      RECT  1905.0 49445.0 2040.0 49510.0 ;
      RECT  2505.0 48647.5 2690.0 48582.5 ;
      RECT  1345.0 48647.5 1530.0 48582.5 ;
      RECT  1462.5 49007.5 1312.5 48942.5 ;
      RECT  2347.5 49007.5 2722.5 48942.5 ;
      RECT  1462.5 48817.5 2347.5 48752.5 ;
      RECT  2347.5 49007.5 2482.5 48942.5 ;
      RECT  2347.5 48817.5 2482.5 48752.5 ;
      RECT  2347.5 48817.5 2482.5 48752.5 ;
      RECT  2347.5 49007.5 2482.5 48942.5 ;
      RECT  1462.5 49007.5 1597.5 48942.5 ;
      RECT  1462.5 48817.5 1597.5 48752.5 ;
      RECT  1462.5 48817.5 1597.5 48752.5 ;
      RECT  1462.5 49007.5 1597.5 48942.5 ;
      RECT  2437.5 48647.5 2572.5 48582.5 ;
      RECT  1462.5 48647.5 1597.5 48582.5 ;
      RECT  1905.0 48950.0 2040.0 48885.0 ;
      RECT  1905.0 48950.0 2040.0 48885.0 ;
      RECT  1940.0 48785.0 2005.0 48720.0 ;
      RECT  2657.5 49075.0 2722.5 48515.0 ;
      RECT  1312.5 49075.0 1377.5 48515.0 ;
      RECT  1905.0 48885.0 2040.0 48950.0 ;
      RECT  2505.0 48087.5 2690.0 48022.5 ;
      RECT  1345.0 48087.5 1530.0 48022.5 ;
      RECT  1462.5 48447.5 1312.5 48382.5 ;
      RECT  2347.5 48447.5 2722.5 48382.5 ;
      RECT  1462.5 48257.5 2347.5 48192.5 ;
      RECT  2347.5 48447.5 2482.5 48382.5 ;
      RECT  2347.5 48257.5 2482.5 48192.5 ;
      RECT  2347.5 48257.5 2482.5 48192.5 ;
      RECT  2347.5 48447.5 2482.5 48382.5 ;
      RECT  1462.5 48447.5 1597.5 48382.5 ;
      RECT  1462.5 48257.5 1597.5 48192.5 ;
      RECT  1462.5 48257.5 1597.5 48192.5 ;
      RECT  1462.5 48447.5 1597.5 48382.5 ;
      RECT  2437.5 48087.5 2572.5 48022.5 ;
      RECT  1462.5 48087.5 1597.5 48022.5 ;
      RECT  1905.0 48390.0 2040.0 48325.0 ;
      RECT  1905.0 48390.0 2040.0 48325.0 ;
      RECT  1940.0 48225.0 2005.0 48160.0 ;
      RECT  2657.5 48515.0 2722.5 47955.0 ;
      RECT  1312.5 48515.0 1377.5 47955.0 ;
      RECT  1905.0 48325.0 2040.0 48390.0 ;
      RECT  2505.0 47527.5 2690.0 47462.5 ;
      RECT  1345.0 47527.5 1530.0 47462.5 ;
      RECT  1462.5 47887.5 1312.5 47822.5 ;
      RECT  2347.5 47887.5 2722.5 47822.5 ;
      RECT  1462.5 47697.5 2347.5 47632.5 ;
      RECT  2347.5 47887.5 2482.5 47822.5 ;
      RECT  2347.5 47697.5 2482.5 47632.5 ;
      RECT  2347.5 47697.5 2482.5 47632.5 ;
      RECT  2347.5 47887.5 2482.5 47822.5 ;
      RECT  1462.5 47887.5 1597.5 47822.5 ;
      RECT  1462.5 47697.5 1597.5 47632.5 ;
      RECT  1462.5 47697.5 1597.5 47632.5 ;
      RECT  1462.5 47887.5 1597.5 47822.5 ;
      RECT  2437.5 47527.5 2572.5 47462.5 ;
      RECT  1462.5 47527.5 1597.5 47462.5 ;
      RECT  1905.0 47830.0 2040.0 47765.0 ;
      RECT  1905.0 47830.0 2040.0 47765.0 ;
      RECT  1940.0 47665.0 2005.0 47600.0 ;
      RECT  2657.5 47955.0 2722.5 47395.0 ;
      RECT  1312.5 47955.0 1377.5 47395.0 ;
      RECT  1905.0 47765.0 2040.0 47830.0 ;
      RECT  2505.0 46967.5 2690.0 46902.5 ;
      RECT  1345.0 46967.5 1530.0 46902.5 ;
      RECT  1462.5 47327.5 1312.5 47262.5 ;
      RECT  2347.5 47327.5 2722.5 47262.5 ;
      RECT  1462.5 47137.5 2347.5 47072.5 ;
      RECT  2347.5 47327.5 2482.5 47262.5 ;
      RECT  2347.5 47137.5 2482.5 47072.5 ;
      RECT  2347.5 47137.5 2482.5 47072.5 ;
      RECT  2347.5 47327.5 2482.5 47262.5 ;
      RECT  1462.5 47327.5 1597.5 47262.5 ;
      RECT  1462.5 47137.5 1597.5 47072.5 ;
      RECT  1462.5 47137.5 1597.5 47072.5 ;
      RECT  1462.5 47327.5 1597.5 47262.5 ;
      RECT  2437.5 46967.5 2572.5 46902.5 ;
      RECT  1462.5 46967.5 1597.5 46902.5 ;
      RECT  1905.0 47270.0 2040.0 47205.0 ;
      RECT  1905.0 47270.0 2040.0 47205.0 ;
      RECT  1940.0 47105.0 2005.0 47040.0 ;
      RECT  2657.5 47395.0 2722.5 46835.0 ;
      RECT  1312.5 47395.0 1377.5 46835.0 ;
      RECT  1905.0 47205.0 2040.0 47270.0 ;
      RECT  2505.0 46407.5 2690.0 46342.5 ;
      RECT  1345.0 46407.5 1530.0 46342.5 ;
      RECT  1462.5 46767.5 1312.5 46702.5 ;
      RECT  2347.5 46767.5 2722.5 46702.5 ;
      RECT  1462.5 46577.5 2347.5 46512.5 ;
      RECT  2347.5 46767.5 2482.5 46702.5 ;
      RECT  2347.5 46577.5 2482.5 46512.5 ;
      RECT  2347.5 46577.5 2482.5 46512.5 ;
      RECT  2347.5 46767.5 2482.5 46702.5 ;
      RECT  1462.5 46767.5 1597.5 46702.5 ;
      RECT  1462.5 46577.5 1597.5 46512.5 ;
      RECT  1462.5 46577.5 1597.5 46512.5 ;
      RECT  1462.5 46767.5 1597.5 46702.5 ;
      RECT  2437.5 46407.5 2572.5 46342.5 ;
      RECT  1462.5 46407.5 1597.5 46342.5 ;
      RECT  1905.0 46710.0 2040.0 46645.0 ;
      RECT  1905.0 46710.0 2040.0 46645.0 ;
      RECT  1940.0 46545.0 2005.0 46480.0 ;
      RECT  2657.5 46835.0 2722.5 46275.0 ;
      RECT  1312.5 46835.0 1377.5 46275.0 ;
      RECT  1905.0 46645.0 2040.0 46710.0 ;
      RECT  2505.0 45847.5 2690.0 45782.5 ;
      RECT  1345.0 45847.5 1530.0 45782.5 ;
      RECT  1462.5 46207.5 1312.5 46142.5 ;
      RECT  2347.5 46207.5 2722.5 46142.5 ;
      RECT  1462.5 46017.5 2347.5 45952.5 ;
      RECT  2347.5 46207.5 2482.5 46142.5 ;
      RECT  2347.5 46017.5 2482.5 45952.5 ;
      RECT  2347.5 46017.5 2482.5 45952.5 ;
      RECT  2347.5 46207.5 2482.5 46142.5 ;
      RECT  1462.5 46207.5 1597.5 46142.5 ;
      RECT  1462.5 46017.5 1597.5 45952.5 ;
      RECT  1462.5 46017.5 1597.5 45952.5 ;
      RECT  1462.5 46207.5 1597.5 46142.5 ;
      RECT  2437.5 45847.5 2572.5 45782.5 ;
      RECT  1462.5 45847.5 1597.5 45782.5 ;
      RECT  1905.0 46150.0 2040.0 46085.0 ;
      RECT  1905.0 46150.0 2040.0 46085.0 ;
      RECT  1940.0 45985.0 2005.0 45920.0 ;
      RECT  2657.5 46275.0 2722.5 45715.0 ;
      RECT  1312.5 46275.0 1377.5 45715.0 ;
      RECT  1905.0 46085.0 2040.0 46150.0 ;
      RECT  2505.0 45287.5 2690.0 45222.5 ;
      RECT  1345.0 45287.5 1530.0 45222.5 ;
      RECT  1462.5 45647.5 1312.5 45582.5 ;
      RECT  2347.5 45647.5 2722.5 45582.5 ;
      RECT  1462.5 45457.5 2347.5 45392.5 ;
      RECT  2347.5 45647.5 2482.5 45582.5 ;
      RECT  2347.5 45457.5 2482.5 45392.5 ;
      RECT  2347.5 45457.5 2482.5 45392.5 ;
      RECT  2347.5 45647.5 2482.5 45582.5 ;
      RECT  1462.5 45647.5 1597.5 45582.5 ;
      RECT  1462.5 45457.5 1597.5 45392.5 ;
      RECT  1462.5 45457.5 1597.5 45392.5 ;
      RECT  1462.5 45647.5 1597.5 45582.5 ;
      RECT  2437.5 45287.5 2572.5 45222.5 ;
      RECT  1462.5 45287.5 1597.5 45222.5 ;
      RECT  1905.0 45590.0 2040.0 45525.0 ;
      RECT  1905.0 45590.0 2040.0 45525.0 ;
      RECT  1940.0 45425.0 2005.0 45360.0 ;
      RECT  2657.5 45715.0 2722.5 45155.0 ;
      RECT  1312.5 45715.0 1377.5 45155.0 ;
      RECT  1905.0 45525.0 2040.0 45590.0 ;
      RECT  2505.0 44727.5 2690.0 44662.5 ;
      RECT  1345.0 44727.5 1530.0 44662.5 ;
      RECT  1462.5 45087.5 1312.5 45022.5 ;
      RECT  2347.5 45087.5 2722.5 45022.5 ;
      RECT  1462.5 44897.5 2347.5 44832.5 ;
      RECT  2347.5 45087.5 2482.5 45022.5 ;
      RECT  2347.5 44897.5 2482.5 44832.5 ;
      RECT  2347.5 44897.5 2482.5 44832.5 ;
      RECT  2347.5 45087.5 2482.5 45022.5 ;
      RECT  1462.5 45087.5 1597.5 45022.5 ;
      RECT  1462.5 44897.5 1597.5 44832.5 ;
      RECT  1462.5 44897.5 1597.5 44832.5 ;
      RECT  1462.5 45087.5 1597.5 45022.5 ;
      RECT  2437.5 44727.5 2572.5 44662.5 ;
      RECT  1462.5 44727.5 1597.5 44662.5 ;
      RECT  1905.0 45030.0 2040.0 44965.0 ;
      RECT  1905.0 45030.0 2040.0 44965.0 ;
      RECT  1940.0 44865.0 2005.0 44800.0 ;
      RECT  2657.5 45155.0 2722.5 44595.0 ;
      RECT  1312.5 45155.0 1377.5 44595.0 ;
      RECT  1905.0 44965.0 2040.0 45030.0 ;
      RECT  2505.0 44167.5 2690.0 44102.5 ;
      RECT  1345.0 44167.5 1530.0 44102.5 ;
      RECT  1462.5 44527.5 1312.5 44462.5 ;
      RECT  2347.5 44527.5 2722.5 44462.5 ;
      RECT  1462.5 44337.5 2347.5 44272.5 ;
      RECT  2347.5 44527.5 2482.5 44462.5 ;
      RECT  2347.5 44337.5 2482.5 44272.5 ;
      RECT  2347.5 44337.5 2482.5 44272.5 ;
      RECT  2347.5 44527.5 2482.5 44462.5 ;
      RECT  1462.5 44527.5 1597.5 44462.5 ;
      RECT  1462.5 44337.5 1597.5 44272.5 ;
      RECT  1462.5 44337.5 1597.5 44272.5 ;
      RECT  1462.5 44527.5 1597.5 44462.5 ;
      RECT  2437.5 44167.5 2572.5 44102.5 ;
      RECT  1462.5 44167.5 1597.5 44102.5 ;
      RECT  1905.0 44470.0 2040.0 44405.0 ;
      RECT  1905.0 44470.0 2040.0 44405.0 ;
      RECT  1940.0 44305.0 2005.0 44240.0 ;
      RECT  2657.5 44595.0 2722.5 44035.0 ;
      RECT  1312.5 44595.0 1377.5 44035.0 ;
      RECT  1905.0 44405.0 2040.0 44470.0 ;
      RECT  2505.0 43607.5 2690.0 43542.5 ;
      RECT  1345.0 43607.5 1530.0 43542.5 ;
      RECT  1462.5 43967.5 1312.5 43902.5 ;
      RECT  2347.5 43967.5 2722.5 43902.5 ;
      RECT  1462.5 43777.5 2347.5 43712.5 ;
      RECT  2347.5 43967.5 2482.5 43902.5 ;
      RECT  2347.5 43777.5 2482.5 43712.5 ;
      RECT  2347.5 43777.5 2482.5 43712.5 ;
      RECT  2347.5 43967.5 2482.5 43902.5 ;
      RECT  1462.5 43967.5 1597.5 43902.5 ;
      RECT  1462.5 43777.5 1597.5 43712.5 ;
      RECT  1462.5 43777.5 1597.5 43712.5 ;
      RECT  1462.5 43967.5 1597.5 43902.5 ;
      RECT  2437.5 43607.5 2572.5 43542.5 ;
      RECT  1462.5 43607.5 1597.5 43542.5 ;
      RECT  1905.0 43910.0 2040.0 43845.0 ;
      RECT  1905.0 43910.0 2040.0 43845.0 ;
      RECT  1940.0 43745.0 2005.0 43680.0 ;
      RECT  2657.5 44035.0 2722.5 43475.0 ;
      RECT  1312.5 44035.0 1377.5 43475.0 ;
      RECT  1905.0 43845.0 2040.0 43910.0 ;
      RECT  2505.0 43047.5 2690.0 42982.5 ;
      RECT  1345.0 43047.5 1530.0 42982.5 ;
      RECT  1462.5 43407.5 1312.5 43342.5 ;
      RECT  2347.5 43407.5 2722.5 43342.5 ;
      RECT  1462.5 43217.5 2347.5 43152.5 ;
      RECT  2347.5 43407.5 2482.5 43342.5 ;
      RECT  2347.5 43217.5 2482.5 43152.5 ;
      RECT  2347.5 43217.5 2482.5 43152.5 ;
      RECT  2347.5 43407.5 2482.5 43342.5 ;
      RECT  1462.5 43407.5 1597.5 43342.5 ;
      RECT  1462.5 43217.5 1597.5 43152.5 ;
      RECT  1462.5 43217.5 1597.5 43152.5 ;
      RECT  1462.5 43407.5 1597.5 43342.5 ;
      RECT  2437.5 43047.5 2572.5 42982.5 ;
      RECT  1462.5 43047.5 1597.5 42982.5 ;
      RECT  1905.0 43350.0 2040.0 43285.0 ;
      RECT  1905.0 43350.0 2040.0 43285.0 ;
      RECT  1940.0 43185.0 2005.0 43120.0 ;
      RECT  2657.5 43475.0 2722.5 42915.0 ;
      RECT  1312.5 43475.0 1377.5 42915.0 ;
      RECT  1905.0 43285.0 2040.0 43350.0 ;
      RECT  2505.0 42487.5 2690.0 42422.5 ;
      RECT  1345.0 42487.5 1530.0 42422.5 ;
      RECT  1462.5 42847.5 1312.5 42782.5 ;
      RECT  2347.5 42847.5 2722.5 42782.5 ;
      RECT  1462.5 42657.5 2347.5 42592.5 ;
      RECT  2347.5 42847.5 2482.5 42782.5 ;
      RECT  2347.5 42657.5 2482.5 42592.5 ;
      RECT  2347.5 42657.5 2482.5 42592.5 ;
      RECT  2347.5 42847.5 2482.5 42782.5 ;
      RECT  1462.5 42847.5 1597.5 42782.5 ;
      RECT  1462.5 42657.5 1597.5 42592.5 ;
      RECT  1462.5 42657.5 1597.5 42592.5 ;
      RECT  1462.5 42847.5 1597.5 42782.5 ;
      RECT  2437.5 42487.5 2572.5 42422.5 ;
      RECT  1462.5 42487.5 1597.5 42422.5 ;
      RECT  1905.0 42790.0 2040.0 42725.0 ;
      RECT  1905.0 42790.0 2040.0 42725.0 ;
      RECT  1940.0 42625.0 2005.0 42560.0 ;
      RECT  2657.5 42915.0 2722.5 42355.0 ;
      RECT  1312.5 42915.0 1377.5 42355.0 ;
      RECT  1905.0 42725.0 2040.0 42790.0 ;
      RECT  3340.0 42645.0 3475.0 42710.0 ;
      RECT  3340.0 44885.0 3475.0 44950.0 ;
      RECT  3340.0 47125.0 3475.0 47190.0 ;
      RECT  3340.0 49365.0 3475.0 49430.0 ;
      RECT  3340.0 51605.0 3475.0 51670.0 ;
      RECT  1905.0 49280.0 2040.0 49345.0 ;
      RECT  1905.0 47040.0 2040.0 47105.0 ;
      RECT  1905.0 44800.0 2040.0 44865.0 ;
      RECT  3340.0 42480.0 3475.0 42545.0 ;
      RECT  1940.0 42355.0 2005.0 42560.0 ;
      RECT  2657.5 42355.0 2722.5 51875.0 ;
      RECT  1312.5 42355.0 1377.5 51875.0 ;
      RECT  4002.5 42355.0 4067.5 51875.0 ;
      RECT  935.0 42020.0 225.0 40675.0 ;
      RECT  935.0 42020.0 230.0 43365.0 ;
      RECT  935.0 44710.0 230.0 43365.0 ;
      RECT  935.0 44710.0 230.0 46055.0 ;
      RECT  935.0 47400.0 230.0 46055.0 ;
      RECT  1025.0 42127.5 140.0 42192.5 ;
      RECT  1025.0 44537.5 140.0 44602.5 ;
      RECT  1025.0 44817.5 140.0 44882.5 ;
      RECT  1025.0 47227.5 140.0 47292.5 ;
      RECT  1025.0 43332.5 140.0 43397.5 ;
      RECT  1025.0 46022.5 140.0 46087.5 ;
      RECT  1025.0 41987.5 140.0 42052.5 ;
      RECT  1025.0 44677.5 140.0 44742.5 ;
      RECT  1025.0 47367.5 140.0 47432.5 ;
      RECT  1345.0 42092.5 1280.0 42227.5 ;
      RECT  1345.0 44502.5 1280.0 44637.5 ;
      RECT  1345.0 44782.5 1280.0 44917.5 ;
      RECT  1345.0 47192.5 1280.0 47327.5 ;
      RECT  1342.5 42355.0 1277.5 42490.0 ;
      RECT  1377.5 39980.0 1312.5 40115.0 ;
      RECT  867.5 40082.5 1002.5 40147.5 ;
      RECT  162.5 40082.5 297.5 40147.5 ;
      RECT  2005.0 41587.5 1940.0 41722.5 ;
      RECT  1105.0 40847.5 1240.0 40912.5 ;
      RECT  1105.0 40250.0 1240.0 40315.0 ;
      RECT  682.5 40250.0 817.5 40315.0 ;
      RECT  3475.0 39555.0 3410.0 42480.0 ;
      RECT  2005.0 39555.0 1940.0 40320.0 ;
      RECT  20.0 39555.0 -45.0 47487.5 ;
      RECT  2722.5 39555.0 2657.5 42355.0 ;
      RECT  1377.5 39555.0 1312.5 40115.0 ;
      RECT  4067.5 39555.0 4002.5 42355.0 ;
      RECT  3455.0 34402.5 3390.0 34267.5 ;
      RECT  3455.0 30322.5 3390.0 30187.5 ;
      RECT  2517.5 27755.0 2452.5 27620.0 ;
      RECT  1962.5 34402.5 1897.5 34267.5 ;
      RECT  1747.5 34812.5 1682.5 34677.5 ;
      RECT  2017.5 37350.0 1952.5 37215.0 ;
      RECT  1802.5 37607.5 1737.5 37472.5 ;
      RECT  3380.0 35837.5 3315.0 35702.5 ;
      RECT  3520.0 35632.5 3455.0 35497.5 ;
      RECT  3660.0 35017.5 3595.0 34882.5 ;
      RECT  690.0 35837.5 625.0 35702.5 ;
      RECT  830.0 35017.5 765.0 34882.5 ;
      RECT  970.0 35222.5 905.0 35087.5 ;
      RECT  1997.5 37032.5 1862.5 37097.5 ;
      RECT  2052.5 38177.5 1917.5 38242.5 ;
      RECT  785.0 39362.5 650.0 39427.5 ;
      RECT  2040.0 38402.5 1905.0 38467.5 ;
      RECT  4067.5 34607.5 4002.5 34472.5 ;
      RECT  2722.5 35427.5 2657.5 35292.5 ;
      RECT  1377.5 34607.5 1312.5 34472.5 ;
      RECT  32.5 35427.5 -32.5 35292.5 ;
      RECT  3475.0 27450.0 3340.0 27640.0 ;
      RECT  2722.5 27450.0 2657.5 27515.0 ;
      RECT  4067.5 27450.0 4002.5 27515.0 ;
      RECT  4417.5 35327.5 4282.5 35392.5 ;
   LAYER  metal2 ;
      RECT  15572.5 38230.0 15642.5 38435.0 ;
      RECT  15367.5 39190.0 15437.5 39395.0 ;
      RECT  14957.5 36860.0 15027.5 37065.0 ;
      RECT  14752.5 38005.0 14822.5 38210.0 ;
      RECT  15162.5 35565.0 15232.5 35770.0 ;
      RECT  14547.5 34130.0 14617.5 34335.0 ;
      RECT  4035.0 35325.0 4350.0 35395.0 ;
      RECT  14132.5 34335.0 14202.5 34540.0 ;
      RECT  14547.5 35.0 14617.5 72077.5 ;
      RECT  14752.5 35.0 14822.5 72077.5 ;
      RECT  14957.5 35.0 15027.5 72077.5 ;
      RECT  15162.5 35.0 15232.5 72077.5 ;
      RECT  15367.5 35.0 15437.5 72077.5 ;
      RECT  15572.5 35.0 15642.5 72077.5 ;
      RECT  11942.5 35.0 12012.5 27310.0 ;
      RECT  12147.5 35.0 12217.5 27310.0 ;
      RECT  12352.5 35.0 12422.5 27310.0 ;
      RECT  12557.5 35.0 12627.5 27310.0 ;
      RECT  12762.5 35.0 12832.5 27310.0 ;
      RECT  12967.5 35.0 13037.5 27310.0 ;
      RECT  13172.5 35.0 13242.5 27310.0 ;
      RECT  13377.5 35.0 13447.5 27310.0 ;
      RECT  13582.5 35.0 13652.5 27310.0 ;
      RECT  16235.0 70505.0 16305.0 70910.0 ;
      RECT  16570.0 70505.0 16640.0 70910.0 ;
      RECT  16940.0 70505.0 17010.0 70910.0 ;
      RECT  17275.0 70505.0 17345.0 70910.0 ;
      RECT  17645.0 70505.0 17715.0 70910.0 ;
      RECT  17980.0 70505.0 18050.0 70910.0 ;
      RECT  18350.0 70505.0 18420.0 70910.0 ;
      RECT  18685.0 70505.0 18755.0 70910.0 ;
      RECT  19055.0 70505.0 19125.0 70910.0 ;
      RECT  19390.0 70505.0 19460.0 70910.0 ;
      RECT  19760.0 70505.0 19830.0 70910.0 ;
      RECT  20095.0 70505.0 20165.0 70910.0 ;
      RECT  20465.0 70505.0 20535.0 70910.0 ;
      RECT  20800.0 70505.0 20870.0 70910.0 ;
      RECT  21170.0 70505.0 21240.0 70910.0 ;
      RECT  21505.0 70505.0 21575.0 70910.0 ;
      RECT  16402.5 5815.0 16472.5 5885.0 ;
      RECT  16227.5 5815.0 16437.5 5885.0 ;
      RECT  16402.5 5850.0 16472.5 5990.0 ;
      RECT  19222.5 5815.0 19292.5 5885.0 ;
      RECT  19047.5 5815.0 19257.5 5885.0 ;
      RECT  19222.5 5850.0 19292.5 5990.0 ;
      RECT  8430.0 70350.0 8500.0 70555.0 ;
      RECT  16085.0 27310.0 16790.0 28655.0 ;
      RECT  16085.0 30000.0 16790.0 28655.0 ;
      RECT  16085.0 30000.0 16790.0 31345.0 ;
      RECT  16085.0 32690.0 16790.0 31345.0 ;
      RECT  16085.0 32690.0 16790.0 34035.0 ;
      RECT  16085.0 35380.0 16790.0 34035.0 ;
      RECT  16085.0 35380.0 16790.0 36725.0 ;
      RECT  16085.0 38070.0 16790.0 36725.0 ;
      RECT  16085.0 38070.0 16790.0 39415.0 ;
      RECT  16085.0 40760.0 16790.0 39415.0 ;
      RECT  16085.0 40760.0 16790.0 42105.0 ;
      RECT  16085.0 43450.0 16790.0 42105.0 ;
      RECT  16085.0 43450.0 16790.0 44795.0 ;
      RECT  16085.0 46140.0 16790.0 44795.0 ;
      RECT  16085.0 46140.0 16790.0 47485.0 ;
      RECT  16085.0 48830.0 16790.0 47485.0 ;
      RECT  16085.0 48830.0 16790.0 50175.0 ;
      RECT  16085.0 51520.0 16790.0 50175.0 ;
      RECT  16085.0 51520.0 16790.0 52865.0 ;
      RECT  16085.0 54210.0 16790.0 52865.0 ;
      RECT  16085.0 54210.0 16790.0 55555.0 ;
      RECT  16085.0 56900.0 16790.0 55555.0 ;
      RECT  16085.0 56900.0 16790.0 58245.0 ;
      RECT  16085.0 59590.0 16790.0 58245.0 ;
      RECT  16085.0 59590.0 16790.0 60935.0 ;
      RECT  16085.0 62280.0 16790.0 60935.0 ;
      RECT  16085.0 62280.0 16790.0 63625.0 ;
      RECT  16085.0 64970.0 16790.0 63625.0 ;
      RECT  16085.0 64970.0 16790.0 66315.0 ;
      RECT  16085.0 67660.0 16790.0 66315.0 ;
      RECT  16085.0 67660.0 16790.0 69005.0 ;
      RECT  16085.0 70350.0 16790.0 69005.0 ;
      RECT  16790.0 27310.0 17495.0 28655.0 ;
      RECT  16790.0 30000.0 17495.0 28655.0 ;
      RECT  16790.0 30000.0 17495.0 31345.0 ;
      RECT  16790.0 32690.0 17495.0 31345.0 ;
      RECT  16790.0 32690.0 17495.0 34035.0 ;
      RECT  16790.0 35380.0 17495.0 34035.0 ;
      RECT  16790.0 35380.0 17495.0 36725.0 ;
      RECT  16790.0 38070.0 17495.0 36725.0 ;
      RECT  16790.0 38070.0 17495.0 39415.0 ;
      RECT  16790.0 40760.0 17495.0 39415.0 ;
      RECT  16790.0 40760.0 17495.0 42105.0 ;
      RECT  16790.0 43450.0 17495.0 42105.0 ;
      RECT  16790.0 43450.0 17495.0 44795.0 ;
      RECT  16790.0 46140.0 17495.0 44795.0 ;
      RECT  16790.0 46140.0 17495.0 47485.0 ;
      RECT  16790.0 48830.0 17495.0 47485.0 ;
      RECT  16790.0 48830.0 17495.0 50175.0 ;
      RECT  16790.0 51520.0 17495.0 50175.0 ;
      RECT  16790.0 51520.0 17495.0 52865.0 ;
      RECT  16790.0 54210.0 17495.0 52865.0 ;
      RECT  16790.0 54210.0 17495.0 55555.0 ;
      RECT  16790.0 56900.0 17495.0 55555.0 ;
      RECT  16790.0 56900.0 17495.0 58245.0 ;
      RECT  16790.0 59590.0 17495.0 58245.0 ;
      RECT  16790.0 59590.0 17495.0 60935.0 ;
      RECT  16790.0 62280.0 17495.0 60935.0 ;
      RECT  16790.0 62280.0 17495.0 63625.0 ;
      RECT  16790.0 64970.0 17495.0 63625.0 ;
      RECT  16790.0 64970.0 17495.0 66315.0 ;
      RECT  16790.0 67660.0 17495.0 66315.0 ;
      RECT  16790.0 67660.0 17495.0 69005.0 ;
      RECT  16790.0 70350.0 17495.0 69005.0 ;
      RECT  17495.0 27310.0 18200.0 28655.0 ;
      RECT  17495.0 30000.0 18200.0 28655.0 ;
      RECT  17495.0 30000.0 18200.0 31345.0 ;
      RECT  17495.0 32690.0 18200.0 31345.0 ;
      RECT  17495.0 32690.0 18200.0 34035.0 ;
      RECT  17495.0 35380.0 18200.0 34035.0 ;
      RECT  17495.0 35380.0 18200.0 36725.0 ;
      RECT  17495.0 38070.0 18200.0 36725.0 ;
      RECT  17495.0 38070.0 18200.0 39415.0 ;
      RECT  17495.0 40760.0 18200.0 39415.0 ;
      RECT  17495.0 40760.0 18200.0 42105.0 ;
      RECT  17495.0 43450.0 18200.0 42105.0 ;
      RECT  17495.0 43450.0 18200.0 44795.0 ;
      RECT  17495.0 46140.0 18200.0 44795.0 ;
      RECT  17495.0 46140.0 18200.0 47485.0 ;
      RECT  17495.0 48830.0 18200.0 47485.0 ;
      RECT  17495.0 48830.0 18200.0 50175.0 ;
      RECT  17495.0 51520.0 18200.0 50175.0 ;
      RECT  17495.0 51520.0 18200.0 52865.0 ;
      RECT  17495.0 54210.0 18200.0 52865.0 ;
      RECT  17495.0 54210.0 18200.0 55555.0 ;
      RECT  17495.0 56900.0 18200.0 55555.0 ;
      RECT  17495.0 56900.0 18200.0 58245.0 ;
      RECT  17495.0 59590.0 18200.0 58245.0 ;
      RECT  17495.0 59590.0 18200.0 60935.0 ;
      RECT  17495.0 62280.0 18200.0 60935.0 ;
      RECT  17495.0 62280.0 18200.0 63625.0 ;
      RECT  17495.0 64970.0 18200.0 63625.0 ;
      RECT  17495.0 64970.0 18200.0 66315.0 ;
      RECT  17495.0 67660.0 18200.0 66315.0 ;
      RECT  17495.0 67660.0 18200.0 69005.0 ;
      RECT  17495.0 70350.0 18200.0 69005.0 ;
      RECT  18200.0 27310.0 18905.0 28655.0 ;
      RECT  18200.0 30000.0 18905.0 28655.0 ;
      RECT  18200.0 30000.0 18905.0 31345.0 ;
      RECT  18200.0 32690.0 18905.0 31345.0 ;
      RECT  18200.0 32690.0 18905.0 34035.0 ;
      RECT  18200.0 35380.0 18905.0 34035.0 ;
      RECT  18200.0 35380.0 18905.0 36725.0 ;
      RECT  18200.0 38070.0 18905.0 36725.0 ;
      RECT  18200.0 38070.0 18905.0 39415.0 ;
      RECT  18200.0 40760.0 18905.0 39415.0 ;
      RECT  18200.0 40760.0 18905.0 42105.0 ;
      RECT  18200.0 43450.0 18905.0 42105.0 ;
      RECT  18200.0 43450.0 18905.0 44795.0 ;
      RECT  18200.0 46140.0 18905.0 44795.0 ;
      RECT  18200.0 46140.0 18905.0 47485.0 ;
      RECT  18200.0 48830.0 18905.0 47485.0 ;
      RECT  18200.0 48830.0 18905.0 50175.0 ;
      RECT  18200.0 51520.0 18905.0 50175.0 ;
      RECT  18200.0 51520.0 18905.0 52865.0 ;
      RECT  18200.0 54210.0 18905.0 52865.0 ;
      RECT  18200.0 54210.0 18905.0 55555.0 ;
      RECT  18200.0 56900.0 18905.0 55555.0 ;
      RECT  18200.0 56900.0 18905.0 58245.0 ;
      RECT  18200.0 59590.0 18905.0 58245.0 ;
      RECT  18200.0 59590.0 18905.0 60935.0 ;
      RECT  18200.0 62280.0 18905.0 60935.0 ;
      RECT  18200.0 62280.0 18905.0 63625.0 ;
      RECT  18200.0 64970.0 18905.0 63625.0 ;
      RECT  18200.0 64970.0 18905.0 66315.0 ;
      RECT  18200.0 67660.0 18905.0 66315.0 ;
      RECT  18200.0 67660.0 18905.0 69005.0 ;
      RECT  18200.0 70350.0 18905.0 69005.0 ;
      RECT  18905.0 27310.0 19610.0 28655.0 ;
      RECT  18905.0 30000.0 19610.0 28655.0 ;
      RECT  18905.0 30000.0 19610.0 31345.0 ;
      RECT  18905.0 32690.0 19610.0 31345.0 ;
      RECT  18905.0 32690.0 19610.0 34035.0 ;
      RECT  18905.0 35380.0 19610.0 34035.0 ;
      RECT  18905.0 35380.0 19610.0 36725.0 ;
      RECT  18905.0 38070.0 19610.0 36725.0 ;
      RECT  18905.0 38070.0 19610.0 39415.0 ;
      RECT  18905.0 40760.0 19610.0 39415.0 ;
      RECT  18905.0 40760.0 19610.0 42105.0 ;
      RECT  18905.0 43450.0 19610.0 42105.0 ;
      RECT  18905.0 43450.0 19610.0 44795.0 ;
      RECT  18905.0 46140.0 19610.0 44795.0 ;
      RECT  18905.0 46140.0 19610.0 47485.0 ;
      RECT  18905.0 48830.0 19610.0 47485.0 ;
      RECT  18905.0 48830.0 19610.0 50175.0 ;
      RECT  18905.0 51520.0 19610.0 50175.0 ;
      RECT  18905.0 51520.0 19610.0 52865.0 ;
      RECT  18905.0 54210.0 19610.0 52865.0 ;
      RECT  18905.0 54210.0 19610.0 55555.0 ;
      RECT  18905.0 56900.0 19610.0 55555.0 ;
      RECT  18905.0 56900.0 19610.0 58245.0 ;
      RECT  18905.0 59590.0 19610.0 58245.0 ;
      RECT  18905.0 59590.0 19610.0 60935.0 ;
      RECT  18905.0 62280.0 19610.0 60935.0 ;
      RECT  18905.0 62280.0 19610.0 63625.0 ;
      RECT  18905.0 64970.0 19610.0 63625.0 ;
      RECT  18905.0 64970.0 19610.0 66315.0 ;
      RECT  18905.0 67660.0 19610.0 66315.0 ;
      RECT  18905.0 67660.0 19610.0 69005.0 ;
      RECT  18905.0 70350.0 19610.0 69005.0 ;
      RECT  19610.0 27310.0 20315.0 28655.0 ;
      RECT  19610.0 30000.0 20315.0 28655.0 ;
      RECT  19610.0 30000.0 20315.0 31345.0 ;
      RECT  19610.0 32690.0 20315.0 31345.0 ;
      RECT  19610.0 32690.0 20315.0 34035.0 ;
      RECT  19610.0 35380.0 20315.0 34035.0 ;
      RECT  19610.0 35380.0 20315.0 36725.0 ;
      RECT  19610.0 38070.0 20315.0 36725.0 ;
      RECT  19610.0 38070.0 20315.0 39415.0 ;
      RECT  19610.0 40760.0 20315.0 39415.0 ;
      RECT  19610.0 40760.0 20315.0 42105.0 ;
      RECT  19610.0 43450.0 20315.0 42105.0 ;
      RECT  19610.0 43450.0 20315.0 44795.0 ;
      RECT  19610.0 46140.0 20315.0 44795.0 ;
      RECT  19610.0 46140.0 20315.0 47485.0 ;
      RECT  19610.0 48830.0 20315.0 47485.0 ;
      RECT  19610.0 48830.0 20315.0 50175.0 ;
      RECT  19610.0 51520.0 20315.0 50175.0 ;
      RECT  19610.0 51520.0 20315.0 52865.0 ;
      RECT  19610.0 54210.0 20315.0 52865.0 ;
      RECT  19610.0 54210.0 20315.0 55555.0 ;
      RECT  19610.0 56900.0 20315.0 55555.0 ;
      RECT  19610.0 56900.0 20315.0 58245.0 ;
      RECT  19610.0 59590.0 20315.0 58245.0 ;
      RECT  19610.0 59590.0 20315.0 60935.0 ;
      RECT  19610.0 62280.0 20315.0 60935.0 ;
      RECT  19610.0 62280.0 20315.0 63625.0 ;
      RECT  19610.0 64970.0 20315.0 63625.0 ;
      RECT  19610.0 64970.0 20315.0 66315.0 ;
      RECT  19610.0 67660.0 20315.0 66315.0 ;
      RECT  19610.0 67660.0 20315.0 69005.0 ;
      RECT  19610.0 70350.0 20315.0 69005.0 ;
      RECT  20315.0 27310.0 21020.0 28655.0 ;
      RECT  20315.0 30000.0 21020.0 28655.0 ;
      RECT  20315.0 30000.0 21020.0 31345.0 ;
      RECT  20315.0 32690.0 21020.0 31345.0 ;
      RECT  20315.0 32690.0 21020.0 34035.0 ;
      RECT  20315.0 35380.0 21020.0 34035.0 ;
      RECT  20315.0 35380.0 21020.0 36725.0 ;
      RECT  20315.0 38070.0 21020.0 36725.0 ;
      RECT  20315.0 38070.0 21020.0 39415.0 ;
      RECT  20315.0 40760.0 21020.0 39415.0 ;
      RECT  20315.0 40760.0 21020.0 42105.0 ;
      RECT  20315.0 43450.0 21020.0 42105.0 ;
      RECT  20315.0 43450.0 21020.0 44795.0 ;
      RECT  20315.0 46140.0 21020.0 44795.0 ;
      RECT  20315.0 46140.0 21020.0 47485.0 ;
      RECT  20315.0 48830.0 21020.0 47485.0 ;
      RECT  20315.0 48830.0 21020.0 50175.0 ;
      RECT  20315.0 51520.0 21020.0 50175.0 ;
      RECT  20315.0 51520.0 21020.0 52865.0 ;
      RECT  20315.0 54210.0 21020.0 52865.0 ;
      RECT  20315.0 54210.0 21020.0 55555.0 ;
      RECT  20315.0 56900.0 21020.0 55555.0 ;
      RECT  20315.0 56900.0 21020.0 58245.0 ;
      RECT  20315.0 59590.0 21020.0 58245.0 ;
      RECT  20315.0 59590.0 21020.0 60935.0 ;
      RECT  20315.0 62280.0 21020.0 60935.0 ;
      RECT  20315.0 62280.0 21020.0 63625.0 ;
      RECT  20315.0 64970.0 21020.0 63625.0 ;
      RECT  20315.0 64970.0 21020.0 66315.0 ;
      RECT  20315.0 67660.0 21020.0 66315.0 ;
      RECT  20315.0 67660.0 21020.0 69005.0 ;
      RECT  20315.0 70350.0 21020.0 69005.0 ;
      RECT  21020.0 27310.0 21725.0 28655.0 ;
      RECT  21020.0 30000.0 21725.0 28655.0 ;
      RECT  21020.0 30000.0 21725.0 31345.0 ;
      RECT  21020.0 32690.0 21725.0 31345.0 ;
      RECT  21020.0 32690.0 21725.0 34035.0 ;
      RECT  21020.0 35380.0 21725.0 34035.0 ;
      RECT  21020.0 35380.0 21725.0 36725.0 ;
      RECT  21020.0 38070.0 21725.0 36725.0 ;
      RECT  21020.0 38070.0 21725.0 39415.0 ;
      RECT  21020.0 40760.0 21725.0 39415.0 ;
      RECT  21020.0 40760.0 21725.0 42105.0 ;
      RECT  21020.0 43450.0 21725.0 42105.0 ;
      RECT  21020.0 43450.0 21725.0 44795.0 ;
      RECT  21020.0 46140.0 21725.0 44795.0 ;
      RECT  21020.0 46140.0 21725.0 47485.0 ;
      RECT  21020.0 48830.0 21725.0 47485.0 ;
      RECT  21020.0 48830.0 21725.0 50175.0 ;
      RECT  21020.0 51520.0 21725.0 50175.0 ;
      RECT  21020.0 51520.0 21725.0 52865.0 ;
      RECT  21020.0 54210.0 21725.0 52865.0 ;
      RECT  21020.0 54210.0 21725.0 55555.0 ;
      RECT  21020.0 56900.0 21725.0 55555.0 ;
      RECT  21020.0 56900.0 21725.0 58245.0 ;
      RECT  21020.0 59590.0 21725.0 58245.0 ;
      RECT  21020.0 59590.0 21725.0 60935.0 ;
      RECT  21020.0 62280.0 21725.0 60935.0 ;
      RECT  21020.0 62280.0 21725.0 63625.0 ;
      RECT  21020.0 64970.0 21725.0 63625.0 ;
      RECT  21020.0 64970.0 21725.0 66315.0 ;
      RECT  21020.0 67660.0 21725.0 66315.0 ;
      RECT  21020.0 67660.0 21725.0 69005.0 ;
      RECT  21020.0 70350.0 21725.0 69005.0 ;
      RECT  16235.0 27210.0 16305.0 70505.0 ;
      RECT  16570.0 27210.0 16640.0 70505.0 ;
      RECT  16940.0 27210.0 17010.0 70505.0 ;
      RECT  17275.0 27210.0 17345.0 70505.0 ;
      RECT  17645.0 27210.0 17715.0 70505.0 ;
      RECT  17980.0 27210.0 18050.0 70505.0 ;
      RECT  18350.0 27210.0 18420.0 70505.0 ;
      RECT  18685.0 27210.0 18755.0 70505.0 ;
      RECT  19055.0 27210.0 19125.0 70505.0 ;
      RECT  19390.0 27210.0 19460.0 70505.0 ;
      RECT  19760.0 27210.0 19830.0 70505.0 ;
      RECT  20095.0 27210.0 20165.0 70505.0 ;
      RECT  20465.0 27210.0 20535.0 70505.0 ;
      RECT  20800.0 27210.0 20870.0 70505.0 ;
      RECT  21170.0 27210.0 21240.0 70505.0 ;
      RECT  21505.0 27210.0 21575.0 70505.0 ;
      RECT  16050.0 27210.0 16120.0 70505.0 ;
      RECT  16755.0 27210.0 16825.0 70505.0 ;
      RECT  17460.0 27210.0 17530.0 70505.0 ;
      RECT  18165.0 27210.0 18235.0 70505.0 ;
      RECT  18870.0 27210.0 18940.0 70505.0 ;
      RECT  19575.0 27210.0 19645.0 70505.0 ;
      RECT  20280.0 27210.0 20350.0 70505.0 ;
      RECT  20985.0 27210.0 21055.0 70505.0 ;
      RECT  21690.0 27210.0 21760.0 70505.0 ;
      RECT  16235.0 71032.5 16312.5 71167.5 ;
      RECT  16437.5 71032.5 16640.0 71167.5 ;
      RECT  16235.0 71562.5 16312.5 71697.5 ;
      RECT  16570.0 71562.5 16692.5 71697.5 ;
      RECT  16245.0 71032.5 16315.0 71167.5 ;
      RECT  16435.0 71032.5 16505.0 71167.5 ;
      RECT  16245.0 71562.5 16315.0 71697.5 ;
      RECT  16625.0 71562.5 16695.0 71697.5 ;
      RECT  16235.0 70910.0 16305.0 72077.5 ;
      RECT  16570.0 70910.0 16640.0 72077.5 ;
      RECT  16940.0 71032.5 17017.5 71167.5 ;
      RECT  17142.5 71032.5 17345.0 71167.5 ;
      RECT  16940.0 71562.5 17017.5 71697.5 ;
      RECT  17275.0 71562.5 17397.5 71697.5 ;
      RECT  16950.0 71032.5 17020.0 71167.5 ;
      RECT  17140.0 71032.5 17210.0 71167.5 ;
      RECT  16950.0 71562.5 17020.0 71697.5 ;
      RECT  17330.0 71562.5 17400.0 71697.5 ;
      RECT  16940.0 70910.0 17010.0 72077.5 ;
      RECT  17275.0 70910.0 17345.0 72077.5 ;
      RECT  17645.0 71032.5 17722.5 71167.5 ;
      RECT  17847.5 71032.5 18050.0 71167.5 ;
      RECT  17645.0 71562.5 17722.5 71697.5 ;
      RECT  17980.0 71562.5 18102.5 71697.5 ;
      RECT  17655.0 71032.5 17725.0 71167.5 ;
      RECT  17845.0 71032.5 17915.0 71167.5 ;
      RECT  17655.0 71562.5 17725.0 71697.5 ;
      RECT  18035.0 71562.5 18105.0 71697.5 ;
      RECT  17645.0 70910.0 17715.0 72077.5 ;
      RECT  17980.0 70910.0 18050.0 72077.5 ;
      RECT  18350.0 71032.5 18427.5 71167.5 ;
      RECT  18552.5 71032.5 18755.0 71167.5 ;
      RECT  18350.0 71562.5 18427.5 71697.5 ;
      RECT  18685.0 71562.5 18807.5 71697.5 ;
      RECT  18360.0 71032.5 18430.0 71167.5 ;
      RECT  18550.0 71032.5 18620.0 71167.5 ;
      RECT  18360.0 71562.5 18430.0 71697.5 ;
      RECT  18740.0 71562.5 18810.0 71697.5 ;
      RECT  18350.0 70910.0 18420.0 72077.5 ;
      RECT  18685.0 70910.0 18755.0 72077.5 ;
      RECT  19055.0 71032.5 19132.5 71167.5 ;
      RECT  19257.5 71032.5 19460.0 71167.5 ;
      RECT  19055.0 71562.5 19132.5 71697.5 ;
      RECT  19390.0 71562.5 19512.5 71697.5 ;
      RECT  19065.0 71032.5 19135.0 71167.5 ;
      RECT  19255.0 71032.5 19325.0 71167.5 ;
      RECT  19065.0 71562.5 19135.0 71697.5 ;
      RECT  19445.0 71562.5 19515.0 71697.5 ;
      RECT  19055.0 70910.0 19125.0 72077.5 ;
      RECT  19390.0 70910.0 19460.0 72077.5 ;
      RECT  19760.0 71032.5 19837.5 71167.5 ;
      RECT  19962.5 71032.5 20165.0 71167.5 ;
      RECT  19760.0 71562.5 19837.5 71697.5 ;
      RECT  20095.0 71562.5 20217.5 71697.5 ;
      RECT  19770.0 71032.5 19840.0 71167.5 ;
      RECT  19960.0 71032.5 20030.0 71167.5 ;
      RECT  19770.0 71562.5 19840.0 71697.5 ;
      RECT  20150.0 71562.5 20220.0 71697.5 ;
      RECT  19760.0 70910.0 19830.0 72077.5 ;
      RECT  20095.0 70910.0 20165.0 72077.5 ;
      RECT  20465.0 71032.5 20542.5 71167.5 ;
      RECT  20667.5 71032.5 20870.0 71167.5 ;
      RECT  20465.0 71562.5 20542.5 71697.5 ;
      RECT  20800.0 71562.5 20922.5 71697.5 ;
      RECT  20475.0 71032.5 20545.0 71167.5 ;
      RECT  20665.0 71032.5 20735.0 71167.5 ;
      RECT  20475.0 71562.5 20545.0 71697.5 ;
      RECT  20855.0 71562.5 20925.0 71697.5 ;
      RECT  20465.0 70910.0 20535.0 72077.5 ;
      RECT  20800.0 70910.0 20870.0 72077.5 ;
      RECT  21170.0 71032.5 21247.5 71167.5 ;
      RECT  21372.5 71032.5 21575.0 71167.5 ;
      RECT  21170.0 71562.5 21247.5 71697.5 ;
      RECT  21505.0 71562.5 21627.5 71697.5 ;
      RECT  21180.0 71032.5 21250.0 71167.5 ;
      RECT  21370.0 71032.5 21440.0 71167.5 ;
      RECT  21180.0 71562.5 21250.0 71697.5 ;
      RECT  21560.0 71562.5 21630.0 71697.5 ;
      RECT  21170.0 70910.0 21240.0 72077.5 ;
      RECT  21505.0 70910.0 21575.0 72077.5 ;
      RECT  16235.0 70910.0 16305.0 72077.5 ;
      RECT  16570.0 70910.0 16640.0 72077.5 ;
      RECT  16940.0 70910.0 17010.0 72077.5 ;
      RECT  17275.0 70910.0 17345.0 72077.5 ;
      RECT  17645.0 70910.0 17715.0 72077.5 ;
      RECT  17980.0 70910.0 18050.0 72077.5 ;
      RECT  18350.0 70910.0 18420.0 72077.5 ;
      RECT  18685.0 70910.0 18755.0 72077.5 ;
      RECT  19055.0 70910.0 19125.0 72077.5 ;
      RECT  19390.0 70910.0 19460.0 72077.5 ;
      RECT  19760.0 70910.0 19830.0 72077.5 ;
      RECT  20095.0 70910.0 20165.0 72077.5 ;
      RECT  20465.0 70910.0 20535.0 72077.5 ;
      RECT  20800.0 70910.0 20870.0 72077.5 ;
      RECT  21170.0 70910.0 21240.0 72077.5 ;
      RECT  21505.0 70910.0 21575.0 72077.5 ;
      RECT  16940.0 24745.0 17010.0 25445.0 ;
      RECT  17275.0 24605.0 17345.0 25445.0 ;
      RECT  17645.0 24745.0 17715.0 25445.0 ;
      RECT  17980.0 24605.0 18050.0 25445.0 ;
      RECT  18350.0 24745.0 18420.0 25445.0 ;
      RECT  18685.0 24605.0 18755.0 25445.0 ;
      RECT  19760.0 24745.0 19830.0 25445.0 ;
      RECT  20095.0 24605.0 20165.0 25445.0 ;
      RECT  20465.0 24745.0 20535.0 25445.0 ;
      RECT  20800.0 24605.0 20870.0 25445.0 ;
      RECT  21170.0 24745.0 21240.0 25445.0 ;
      RECT  21505.0 24605.0 21575.0 25445.0 ;
      RECT  16235.0 26085.0 16305.0 26155.0 ;
      RECT  16307.5 26085.0 16377.5 26155.0 ;
      RECT  16235.0 25585.0 16305.0 26120.0 ;
      RECT  16270.0 26085.0 16342.5 26155.0 ;
      RECT  16307.5 26120.0 16377.5 26652.5 ;
      RECT  16570.0 26497.5 16640.0 26567.5 ;
      RECT  16497.5 26497.5 16567.5 26567.5 ;
      RECT  16570.0 26532.5 16640.0 27135.0 ;
      RECT  16532.5 26497.5 16605.0 26567.5 ;
      RECT  16497.5 25927.5 16567.5 26532.5 ;
      RECT  16235.0 27067.5 16305.0 27202.5 ;
      RECT  16570.0 25517.5 16640.0 25652.5 ;
      RECT  16307.5 26652.5 16377.5 26787.5 ;
      RECT  16497.5 25792.5 16567.5 25927.5 ;
      RECT  16755.0 25692.5 16825.0 25827.5 ;
      RECT  16235.0 27135.0 16305.0 27275.0 ;
      RECT  16570.0 27135.0 16640.0 27275.0 ;
      RECT  16235.0 25445.0 16305.0 25585.0 ;
      RECT  16570.0 25445.0 16640.0 25585.0 ;
      RECT  16050.0 25445.0 16120.0 27275.0 ;
      RECT  16755.0 25445.0 16825.0 27275.0 ;
      RECT  16940.0 26085.0 17010.0 26155.0 ;
      RECT  17012.5 26085.0 17082.5 26155.0 ;
      RECT  16940.0 25585.0 17010.0 26120.0 ;
      RECT  16975.0 26085.0 17047.5 26155.0 ;
      RECT  17012.5 26120.0 17082.5 26652.5 ;
      RECT  17275.0 26497.5 17345.0 26567.5 ;
      RECT  17202.5 26497.5 17272.5 26567.5 ;
      RECT  17275.0 26532.5 17345.0 27135.0 ;
      RECT  17237.5 26497.5 17310.0 26567.5 ;
      RECT  17202.5 25927.5 17272.5 26532.5 ;
      RECT  16940.0 27067.5 17010.0 27202.5 ;
      RECT  17275.0 25517.5 17345.0 25652.5 ;
      RECT  17012.5 26652.5 17082.5 26787.5 ;
      RECT  17202.5 25792.5 17272.5 25927.5 ;
      RECT  17460.0 25692.5 17530.0 25827.5 ;
      RECT  16940.0 27135.0 17010.0 27275.0 ;
      RECT  17275.0 27135.0 17345.0 27275.0 ;
      RECT  16940.0 25445.0 17010.0 25585.0 ;
      RECT  17275.0 25445.0 17345.0 25585.0 ;
      RECT  16755.0 25445.0 16825.0 27275.0 ;
      RECT  17460.0 25445.0 17530.0 27275.0 ;
      RECT  17645.0 26085.0 17715.0 26155.0 ;
      RECT  17717.5 26085.0 17787.5 26155.0 ;
      RECT  17645.0 25585.0 17715.0 26120.0 ;
      RECT  17680.0 26085.0 17752.5 26155.0 ;
      RECT  17717.5 26120.0 17787.5 26652.5 ;
      RECT  17980.0 26497.5 18050.0 26567.5 ;
      RECT  17907.5 26497.5 17977.5 26567.5 ;
      RECT  17980.0 26532.5 18050.0 27135.0 ;
      RECT  17942.5 26497.5 18015.0 26567.5 ;
      RECT  17907.5 25927.5 17977.5 26532.5 ;
      RECT  17645.0 27067.5 17715.0 27202.5 ;
      RECT  17980.0 25517.5 18050.0 25652.5 ;
      RECT  17717.5 26652.5 17787.5 26787.5 ;
      RECT  17907.5 25792.5 17977.5 25927.5 ;
      RECT  18165.0 25692.5 18235.0 25827.5 ;
      RECT  17645.0 27135.0 17715.0 27275.0 ;
      RECT  17980.0 27135.0 18050.0 27275.0 ;
      RECT  17645.0 25445.0 17715.0 25585.0 ;
      RECT  17980.0 25445.0 18050.0 25585.0 ;
      RECT  17460.0 25445.0 17530.0 27275.0 ;
      RECT  18165.0 25445.0 18235.0 27275.0 ;
      RECT  18350.0 26085.0 18420.0 26155.0 ;
      RECT  18422.5 26085.0 18492.5 26155.0 ;
      RECT  18350.0 25585.0 18420.0 26120.0 ;
      RECT  18385.0 26085.0 18457.5 26155.0 ;
      RECT  18422.5 26120.0 18492.5 26652.5 ;
      RECT  18685.0 26497.5 18755.0 26567.5 ;
      RECT  18612.5 26497.5 18682.5 26567.5 ;
      RECT  18685.0 26532.5 18755.0 27135.0 ;
      RECT  18647.5 26497.5 18720.0 26567.5 ;
      RECT  18612.5 25927.5 18682.5 26532.5 ;
      RECT  18350.0 27067.5 18420.0 27202.5 ;
      RECT  18685.0 25517.5 18755.0 25652.5 ;
      RECT  18422.5 26652.5 18492.5 26787.5 ;
      RECT  18612.5 25792.5 18682.5 25927.5 ;
      RECT  18870.0 25692.5 18940.0 25827.5 ;
      RECT  18350.0 27135.0 18420.0 27275.0 ;
      RECT  18685.0 27135.0 18755.0 27275.0 ;
      RECT  18350.0 25445.0 18420.0 25585.0 ;
      RECT  18685.0 25445.0 18755.0 25585.0 ;
      RECT  18165.0 25445.0 18235.0 27275.0 ;
      RECT  18870.0 25445.0 18940.0 27275.0 ;
      RECT  19055.0 26085.0 19125.0 26155.0 ;
      RECT  19127.5 26085.0 19197.5 26155.0 ;
      RECT  19055.0 25585.0 19125.0 26120.0 ;
      RECT  19090.0 26085.0 19162.5 26155.0 ;
      RECT  19127.5 26120.0 19197.5 26652.5 ;
      RECT  19390.0 26497.5 19460.0 26567.5 ;
      RECT  19317.5 26497.5 19387.5 26567.5 ;
      RECT  19390.0 26532.5 19460.0 27135.0 ;
      RECT  19352.5 26497.5 19425.0 26567.5 ;
      RECT  19317.5 25927.5 19387.5 26532.5 ;
      RECT  19055.0 27067.5 19125.0 27202.5 ;
      RECT  19390.0 25517.5 19460.0 25652.5 ;
      RECT  19127.5 26652.5 19197.5 26787.5 ;
      RECT  19317.5 25792.5 19387.5 25927.5 ;
      RECT  19575.0 25692.5 19645.0 25827.5 ;
      RECT  19055.0 27135.0 19125.0 27275.0 ;
      RECT  19390.0 27135.0 19460.0 27275.0 ;
      RECT  19055.0 25445.0 19125.0 25585.0 ;
      RECT  19390.0 25445.0 19460.0 25585.0 ;
      RECT  18870.0 25445.0 18940.0 27275.0 ;
      RECT  19575.0 25445.0 19645.0 27275.0 ;
      RECT  19760.0 26085.0 19830.0 26155.0 ;
      RECT  19832.5 26085.0 19902.5 26155.0 ;
      RECT  19760.0 25585.0 19830.0 26120.0 ;
      RECT  19795.0 26085.0 19867.5 26155.0 ;
      RECT  19832.5 26120.0 19902.5 26652.5 ;
      RECT  20095.0 26497.5 20165.0 26567.5 ;
      RECT  20022.5 26497.5 20092.5 26567.5 ;
      RECT  20095.0 26532.5 20165.0 27135.0 ;
      RECT  20057.5 26497.5 20130.0 26567.5 ;
      RECT  20022.5 25927.5 20092.5 26532.5 ;
      RECT  19760.0 27067.5 19830.0 27202.5 ;
      RECT  20095.0 25517.5 20165.0 25652.5 ;
      RECT  19832.5 26652.5 19902.5 26787.5 ;
      RECT  20022.5 25792.5 20092.5 25927.5 ;
      RECT  20280.0 25692.5 20350.0 25827.5 ;
      RECT  19760.0 27135.0 19830.0 27275.0 ;
      RECT  20095.0 27135.0 20165.0 27275.0 ;
      RECT  19760.0 25445.0 19830.0 25585.0 ;
      RECT  20095.0 25445.0 20165.0 25585.0 ;
      RECT  19575.0 25445.0 19645.0 27275.0 ;
      RECT  20280.0 25445.0 20350.0 27275.0 ;
      RECT  20465.0 26085.0 20535.0 26155.0 ;
      RECT  20537.5 26085.0 20607.5 26155.0 ;
      RECT  20465.0 25585.0 20535.0 26120.0 ;
      RECT  20500.0 26085.0 20572.5 26155.0 ;
      RECT  20537.5 26120.0 20607.5 26652.5 ;
      RECT  20800.0 26497.5 20870.0 26567.5 ;
      RECT  20727.5 26497.5 20797.5 26567.5 ;
      RECT  20800.0 26532.5 20870.0 27135.0 ;
      RECT  20762.5 26497.5 20835.0 26567.5 ;
      RECT  20727.5 25927.5 20797.5 26532.5 ;
      RECT  20465.0 27067.5 20535.0 27202.5 ;
      RECT  20800.0 25517.5 20870.0 25652.5 ;
      RECT  20537.5 26652.5 20607.5 26787.5 ;
      RECT  20727.5 25792.5 20797.5 25927.5 ;
      RECT  20985.0 25692.5 21055.0 25827.5 ;
      RECT  20465.0 27135.0 20535.0 27275.0 ;
      RECT  20800.0 27135.0 20870.0 27275.0 ;
      RECT  20465.0 25445.0 20535.0 25585.0 ;
      RECT  20800.0 25445.0 20870.0 25585.0 ;
      RECT  20280.0 25445.0 20350.0 27275.0 ;
      RECT  20985.0 25445.0 21055.0 27275.0 ;
      RECT  21170.0 26085.0 21240.0 26155.0 ;
      RECT  21242.5 26085.0 21312.5 26155.0 ;
      RECT  21170.0 25585.0 21240.0 26120.0 ;
      RECT  21205.0 26085.0 21277.5 26155.0 ;
      RECT  21242.5 26120.0 21312.5 26652.5 ;
      RECT  21505.0 26497.5 21575.0 26567.5 ;
      RECT  21432.5 26497.5 21502.5 26567.5 ;
      RECT  21505.0 26532.5 21575.0 27135.0 ;
      RECT  21467.5 26497.5 21540.0 26567.5 ;
      RECT  21432.5 25927.5 21502.5 26532.5 ;
      RECT  21170.0 27067.5 21240.0 27202.5 ;
      RECT  21505.0 25517.5 21575.0 25652.5 ;
      RECT  21242.5 26652.5 21312.5 26787.5 ;
      RECT  21432.5 25792.5 21502.5 25927.5 ;
      RECT  21690.0 25692.5 21760.0 25827.5 ;
      RECT  21170.0 27135.0 21240.0 27275.0 ;
      RECT  21505.0 27135.0 21575.0 27275.0 ;
      RECT  21170.0 25445.0 21240.0 25585.0 ;
      RECT  21505.0 25445.0 21575.0 25585.0 ;
      RECT  20985.0 25445.0 21055.0 27275.0 ;
      RECT  21690.0 25445.0 21760.0 27275.0 ;
      RECT  16370.0 24745.0 16235.0 24815.0 ;
      RECT  16570.0 24605.0 16435.0 24675.0 ;
      RECT  17075.0 24745.0 16940.0 24815.0 ;
      RECT  17275.0 24605.0 17140.0 24675.0 ;
      RECT  17780.0 24745.0 17645.0 24815.0 ;
      RECT  17980.0 24605.0 17845.0 24675.0 ;
      RECT  18485.0 24745.0 18350.0 24815.0 ;
      RECT  18685.0 24605.0 18550.0 24675.0 ;
      RECT  19190.0 24745.0 19055.0 24815.0 ;
      RECT  19390.0 24605.0 19255.0 24675.0 ;
      RECT  19895.0 24745.0 19760.0 24815.0 ;
      RECT  20095.0 24605.0 19960.0 24675.0 ;
      RECT  20600.0 24745.0 20465.0 24815.0 ;
      RECT  20800.0 24605.0 20665.0 24675.0 ;
      RECT  21305.0 24745.0 21170.0 24815.0 ;
      RECT  21505.0 24605.0 21370.0 24675.0 ;
      RECT  16235.0 27135.0 16305.0 27275.0 ;
      RECT  16570.0 27135.0 16640.0 27275.0 ;
      RECT  16940.0 27135.0 17010.0 27275.0 ;
      RECT  17275.0 27135.0 17345.0 27275.0 ;
      RECT  17645.0 27135.0 17715.0 27275.0 ;
      RECT  17980.0 27135.0 18050.0 27275.0 ;
      RECT  18350.0 27135.0 18420.0 27275.0 ;
      RECT  18685.0 27135.0 18755.0 27275.0 ;
      RECT  19055.0 27135.0 19125.0 27275.0 ;
      RECT  19390.0 27135.0 19460.0 27275.0 ;
      RECT  19760.0 27135.0 19830.0 27275.0 ;
      RECT  20095.0 27135.0 20165.0 27275.0 ;
      RECT  20465.0 27135.0 20535.0 27275.0 ;
      RECT  20800.0 27135.0 20870.0 27275.0 ;
      RECT  21170.0 27135.0 21240.0 27275.0 ;
      RECT  21505.0 27135.0 21575.0 27275.0 ;
      RECT  16235.0 24465.0 16305.0 25445.0 ;
      RECT  16570.0 24465.0 16640.0 25445.0 ;
      RECT  19055.0 24465.0 19125.0 25445.0 ;
      RECT  19390.0 24465.0 19460.0 25445.0 ;
      RECT  16050.0 24465.0 16120.0 27275.0 ;
      RECT  16755.0 24465.0 16825.0 27275.0 ;
      RECT  17460.0 24465.0 17530.0 27275.0 ;
      RECT  18165.0 24465.0 18235.0 27275.0 ;
      RECT  18870.0 24465.0 18940.0 27275.0 ;
      RECT  19575.0 24465.0 19645.0 27275.0 ;
      RECT  20280.0 24465.0 20350.0 27275.0 ;
      RECT  20985.0 24465.0 21055.0 27275.0 ;
      RECT  9195.0 35.0 9265.0 5275.0 ;
      RECT  9470.0 35.0 9540.0 5275.0 ;
      RECT  8645.0 35.0 8715.0 5275.0 ;
      RECT  8920.0 35.0 8990.0 5275.0 ;
      RECT  10000.0 640.0 10070.0 710.0 ;
      RECT  10190.0 640.0 10260.0 710.0 ;
      RECT  10000.0 675.0 10070.0 1037.5 ;
      RECT  10035.0 640.0 10225.0 710.0 ;
      RECT  10190.0 332.5 10260.0 675.0 ;
      RECT  10000.0 1037.5 10070.0 1172.5 ;
      RECT  10190.0 197.5 10260.0 332.5 ;
      RECT  10292.5 640.0 10157.5 710.0 ;
      RECT  10000.0 2120.0 10070.0 2050.0 ;
      RECT  10190.0 2120.0 10260.0 2050.0 ;
      RECT  10000.0 2085.0 10070.0 1722.5 ;
      RECT  10035.0 2120.0 10225.0 2050.0 ;
      RECT  10190.0 2427.5 10260.0 2085.0 ;
      RECT  10000.0 1722.5 10070.0 1587.5 ;
      RECT  10190.0 2562.5 10260.0 2427.5 ;
      RECT  10292.5 2120.0 10157.5 2050.0 ;
      RECT  10000.0 3330.0 10070.0 3400.0 ;
      RECT  10190.0 3330.0 10260.0 3400.0 ;
      RECT  10000.0 3365.0 10070.0 3727.5 ;
      RECT  10035.0 3330.0 10225.0 3400.0 ;
      RECT  10190.0 3022.5 10260.0 3365.0 ;
      RECT  10000.0 3727.5 10070.0 3862.5 ;
      RECT  10190.0 2887.5 10260.0 3022.5 ;
      RECT  10292.5 3330.0 10157.5 3400.0 ;
      RECT  10000.0 4810.0 10070.0 4740.0 ;
      RECT  10190.0 4810.0 10260.0 4740.0 ;
      RECT  10000.0 4775.0 10070.0 4412.5 ;
      RECT  10035.0 4810.0 10225.0 4740.0 ;
      RECT  10190.0 5117.5 10260.0 4775.0 ;
      RECT  10000.0 4412.5 10070.0 4277.5 ;
      RECT  10190.0 5252.5 10260.0 5117.5 ;
      RECT  10292.5 4810.0 10157.5 4740.0 ;
      RECT  8747.5 1150.0 8612.5 1220.0 ;
      RECT  7362.5 627.5 7227.5 697.5 ;
      RECT  9022.5 2495.0 8887.5 2565.0 ;
      RECT  7637.5 2062.5 7502.5 2132.5 ;
      RECT  7362.5 2825.0 7227.5 2895.0 ;
      RECT  9297.5 2825.0 9162.5 2895.0 ;
      RECT  7637.5 4170.0 7502.5 4240.0 ;
      RECT  9572.5 4170.0 9437.5 4240.0 ;
      RECT  8747.5 640.0 8612.5 710.0 ;
      RECT  9022.5 425.0 8887.5 495.0 ;
      RECT  9297.5 2050.0 9162.5 2120.0 ;
      RECT  9022.5 2265.0 8887.5 2335.0 ;
      RECT  8747.5 3330.0 8612.5 3400.0 ;
      RECT  9572.5 3115.0 9437.5 3185.0 ;
      RECT  9297.5 4740.0 9162.5 4810.0 ;
      RECT  9572.5 4955.0 9437.5 5025.0 ;
      RECT  7260.0 35.0 7330.0 5275.0 ;
      RECT  7535.0 35.0 7605.0 5275.0 ;
      RECT  16085.0 19580.0 16790.0 24465.0 ;
      RECT  18905.0 19580.0 19610.0 24465.0 ;
      RECT  16235.0 19580.0 16305.0 24465.0 ;
      RECT  16570.0 19580.0 16640.0 23665.0 ;
      RECT  19055.0 19580.0 19125.0 24465.0 ;
      RECT  19390.0 19580.0 19460.0 23665.0 ;
      RECT  16085.0 15405.0 16790.0 19580.0 ;
      RECT  18905.0 15405.0 19610.0 19580.0 ;
      RECT  16402.5 15405.0 16472.5 15545.0 ;
      RECT  19222.5 15405.0 19292.5 15545.0 ;
      RECT  16235.0 19280.0 16305.0 19580.0 ;
      RECT  16570.0 17140.0 16640.0 19580.0 ;
      RECT  19055.0 19280.0 19125.0 19580.0 ;
      RECT  19390.0 17140.0 19460.0 19580.0 ;
      RECT  16085.0 8965.0 16790.0 15405.0 ;
      RECT  18905.0 8965.0 19610.0 15405.0 ;
      RECT  16402.5 8965.0 16472.5 9110.0 ;
      RECT  19222.5 8965.0 19292.5 9110.0 ;
      RECT  16402.5 15135.0 16472.5 15405.0 ;
      RECT  16247.5 14717.5 16317.5 15405.0 ;
      RECT  19222.5 15135.0 19292.5 15405.0 ;
      RECT  19067.5 14717.5 19137.5 15405.0 ;
      RECT  16050.0 8965.0 16120.0 15405.0 ;
      RECT  16755.0 8965.0 16825.0 15405.0 ;
      RECT  18870.0 8965.0 18940.0 15405.0 ;
      RECT  19575.0 8965.0 19645.0 15405.0 ;
      RECT  16085.0 8965.0 16790.0 5990.0 ;
      RECT  18905.0 8965.0 19610.0 5990.0 ;
      RECT  16402.5 6230.0 16472.5 5990.0 ;
      RECT  19222.5 6230.0 19292.5 5990.0 ;
      RECT  16402.5 8965.0 16472.5 8615.0 ;
      RECT  19222.5 8965.0 19292.5 8615.0 ;
      RECT  4655.0 11170.0 4725.0 70350.0 ;
      RECT  4830.0 11170.0 4900.0 70350.0 ;
      RECT  5005.0 11170.0 5075.0 70350.0 ;
      RECT  5180.0 11170.0 5250.0 70350.0 ;
      RECT  5355.0 11170.0 5425.0 70350.0 ;
      RECT  5530.0 11170.0 5600.0 70350.0 ;
      RECT  5705.0 11170.0 5775.0 70350.0 ;
      RECT  5880.0 11170.0 5950.0 70350.0 ;
      RECT  6055.0 11170.0 6125.0 70350.0 ;
      RECT  6230.0 11170.0 6300.0 70350.0 ;
      RECT  6405.0 11170.0 6475.0 70350.0 ;
      RECT  6580.0 11170.0 6650.0 70350.0 ;
      RECT  8785.0 11170.0 8715.0 16410.0 ;
      RECT  8510.0 11170.0 8440.0 16410.0 ;
      RECT  9335.0 11170.0 9265.0 16410.0 ;
      RECT  9060.0 11170.0 8990.0 16410.0 ;
      RECT  7980.0 11775.0 7910.0 11845.0 ;
      RECT  7790.0 11775.0 7720.0 11845.0 ;
      RECT  7980.0 11810.0 7910.0 12172.5 ;
      RECT  7945.0 11775.0 7755.0 11845.0 ;
      RECT  7790.0 11467.5 7720.0 11810.0 ;
      RECT  7980.0 12172.5 7910.0 12307.5 ;
      RECT  7790.0 11332.5 7720.0 11467.5 ;
      RECT  7687.5 11775.0 7822.5 11845.0 ;
      RECT  7980.0 13255.0 7910.0 13185.0 ;
      RECT  7790.0 13255.0 7720.0 13185.0 ;
      RECT  7980.0 13220.0 7910.0 12857.5 ;
      RECT  7945.0 13255.0 7755.0 13185.0 ;
      RECT  7790.0 13562.5 7720.0 13220.0 ;
      RECT  7980.0 12857.5 7910.0 12722.5 ;
      RECT  7790.0 13697.5 7720.0 13562.5 ;
      RECT  7687.5 13255.0 7822.5 13185.0 ;
      RECT  7980.0 14465.0 7910.0 14535.0 ;
      RECT  7790.0 14465.0 7720.0 14535.0 ;
      RECT  7980.0 14500.0 7910.0 14862.5 ;
      RECT  7945.0 14465.0 7755.0 14535.0 ;
      RECT  7790.0 14157.5 7720.0 14500.0 ;
      RECT  7980.0 14862.5 7910.0 14997.5 ;
      RECT  7790.0 14022.5 7720.0 14157.5 ;
      RECT  7687.5 14465.0 7822.5 14535.0 ;
      RECT  7980.0 15945.0 7910.0 15875.0 ;
      RECT  7790.0 15945.0 7720.0 15875.0 ;
      RECT  7980.0 15910.0 7910.0 15547.5 ;
      RECT  7945.0 15945.0 7755.0 15875.0 ;
      RECT  7790.0 16252.5 7720.0 15910.0 ;
      RECT  7980.0 15547.5 7910.0 15412.5 ;
      RECT  7790.0 16387.5 7720.0 16252.5 ;
      RECT  7687.5 15945.0 7822.5 15875.0 ;
      RECT  9232.5 12285.0 9367.5 12355.0 ;
      RECT  10617.5 11762.5 10752.5 11832.5 ;
      RECT  8957.5 13630.0 9092.5 13700.0 ;
      RECT  10342.5 13197.5 10477.5 13267.5 ;
      RECT  10617.5 13960.0 10752.5 14030.0 ;
      RECT  8682.5 13960.0 8817.5 14030.0 ;
      RECT  10342.5 15305.0 10477.5 15375.0 ;
      RECT  8407.5 15305.0 8542.5 15375.0 ;
      RECT  9232.5 11775.0 9367.5 11845.0 ;
      RECT  8957.5 11560.0 9092.5 11630.0 ;
      RECT  8682.5 13185.0 8817.5 13255.0 ;
      RECT  8957.5 13400.0 9092.5 13470.0 ;
      RECT  9232.5 14465.0 9367.5 14535.0 ;
      RECT  8407.5 14250.0 8542.5 14320.0 ;
      RECT  8682.5 15875.0 8817.5 15945.0 ;
      RECT  8407.5 16090.0 8542.5 16160.0 ;
      RECT  10720.0 11170.0 10650.0 16410.0 ;
      RECT  10445.0 11170.0 10375.0 16410.0 ;
      RECT  9425.0 16550.0 9355.0 27170.0 ;
      RECT  9150.0 16550.0 9080.0 27170.0 ;
      RECT  8875.0 16550.0 8805.0 27170.0 ;
      RECT  9975.0 16550.0 9905.0 27170.0 ;
      RECT  9700.0 16550.0 9630.0 27170.0 ;
      RECT  8600.0 16550.0 8530.0 27170.0 ;
      RECT  7690.0 16847.5 7620.0 17552.5 ;
      RECT  8070.0 17202.5 8000.0 17272.5 ;
      RECT  7690.0 17202.5 7620.0 17272.5 ;
      RECT  8070.0 17237.5 8000.0 17552.5 ;
      RECT  8035.0 17202.5 7655.0 17272.5 ;
      RECT  7690.0 16847.5 7620.0 17237.5 ;
      RECT  8070.0 17552.5 8000.0 17687.5 ;
      RECT  7690.0 17552.5 7620.0 17687.5 ;
      RECT  7690.0 16712.5 7620.0 16847.5 ;
      RECT  7690.0 17170.0 7620.0 17305.0 ;
      RECT  7690.0 18942.5 7620.0 18237.5 ;
      RECT  8070.0 18587.5 8000.0 18517.5 ;
      RECT  7690.0 18587.5 7620.0 18517.5 ;
      RECT  8070.0 18552.5 8000.0 18237.5 ;
      RECT  8035.0 18587.5 7655.0 18517.5 ;
      RECT  7690.0 18942.5 7620.0 18552.5 ;
      RECT  8070.0 18237.5 8000.0 18102.5 ;
      RECT  7690.0 18237.5 7620.0 18102.5 ;
      RECT  7690.0 19077.5 7620.0 18942.5 ;
      RECT  7690.0 18620.0 7620.0 18485.0 ;
      RECT  7690.0 19537.5 7620.0 20242.5 ;
      RECT  8070.0 19892.5 8000.0 19962.5 ;
      RECT  7690.0 19892.5 7620.0 19962.5 ;
      RECT  8070.0 19927.5 8000.0 20242.5 ;
      RECT  8035.0 19892.5 7655.0 19962.5 ;
      RECT  7690.0 19537.5 7620.0 19927.5 ;
      RECT  8070.0 20242.5 8000.0 20377.5 ;
      RECT  7690.0 20242.5 7620.0 20377.5 ;
      RECT  7690.0 19402.5 7620.0 19537.5 ;
      RECT  7690.0 19860.0 7620.0 19995.0 ;
      RECT  7690.0 21632.5 7620.0 20927.5 ;
      RECT  8070.0 21277.5 8000.0 21207.5 ;
      RECT  7690.0 21277.5 7620.0 21207.5 ;
      RECT  8070.0 21242.5 8000.0 20927.5 ;
      RECT  8035.0 21277.5 7655.0 21207.5 ;
      RECT  7690.0 21632.5 7620.0 21242.5 ;
      RECT  8070.0 20927.5 8000.0 20792.5 ;
      RECT  7690.0 20927.5 7620.0 20792.5 ;
      RECT  7690.0 21767.5 7620.0 21632.5 ;
      RECT  7690.0 21310.0 7620.0 21175.0 ;
      RECT  7690.0 22227.5 7620.0 22932.5 ;
      RECT  8070.0 22582.5 8000.0 22652.5 ;
      RECT  7690.0 22582.5 7620.0 22652.5 ;
      RECT  8070.0 22617.5 8000.0 22932.5 ;
      RECT  8035.0 22582.5 7655.0 22652.5 ;
      RECT  7690.0 22227.5 7620.0 22617.5 ;
      RECT  8070.0 22932.5 8000.0 23067.5 ;
      RECT  7690.0 22932.5 7620.0 23067.5 ;
      RECT  7690.0 22092.5 7620.0 22227.5 ;
      RECT  7690.0 22550.0 7620.0 22685.0 ;
      RECT  7690.0 24322.5 7620.0 23617.5 ;
      RECT  8070.0 23967.5 8000.0 23897.5 ;
      RECT  7690.0 23967.5 7620.0 23897.5 ;
      RECT  8070.0 23932.5 8000.0 23617.5 ;
      RECT  8035.0 23967.5 7655.0 23897.5 ;
      RECT  7690.0 24322.5 7620.0 23932.5 ;
      RECT  8070.0 23617.5 8000.0 23482.5 ;
      RECT  7690.0 23617.5 7620.0 23482.5 ;
      RECT  7690.0 24457.5 7620.0 24322.5 ;
      RECT  7690.0 24000.0 7620.0 23865.0 ;
      RECT  7690.0 24917.5 7620.0 25622.5 ;
      RECT  8070.0 25272.5 8000.0 25342.5 ;
      RECT  7690.0 25272.5 7620.0 25342.5 ;
      RECT  8070.0 25307.5 8000.0 25622.5 ;
      RECT  8035.0 25272.5 7655.0 25342.5 ;
      RECT  7690.0 24917.5 7620.0 25307.5 ;
      RECT  8070.0 25622.5 8000.0 25757.5 ;
      RECT  7690.0 25622.5 7620.0 25757.5 ;
      RECT  7690.0 24782.5 7620.0 24917.5 ;
      RECT  7690.0 25240.0 7620.0 25375.0 ;
      RECT  7690.0 27012.5 7620.0 26307.5 ;
      RECT  8070.0 26657.5 8000.0 26587.5 ;
      RECT  7690.0 26657.5 7620.0 26587.5 ;
      RECT  8070.0 26622.5 8000.0 26307.5 ;
      RECT  8035.0 26657.5 7655.0 26587.5 ;
      RECT  7690.0 27012.5 7620.0 26622.5 ;
      RECT  8070.0 26307.5 8000.0 26172.5 ;
      RECT  7690.0 26307.5 7620.0 26172.5 ;
      RECT  7690.0 27147.5 7620.0 27012.5 ;
      RECT  7690.0 26690.0 7620.0 26555.0 ;
      RECT  9872.5 17665.0 10007.5 17735.0 ;
      RECT  11532.5 17142.5 11667.5 17212.5 ;
      RECT  9597.5 19010.0 9732.5 19080.0 ;
      RECT  11257.5 18577.5 11392.5 18647.5 ;
      RECT  9322.5 20355.0 9457.5 20425.0 ;
      RECT  10982.5 19832.5 11117.5 19902.5 ;
      RECT  11532.5 20685.0 11667.5 20755.0 ;
      RECT  9047.5 20685.0 9182.5 20755.0 ;
      RECT  11257.5 22030.0 11392.5 22100.0 ;
      RECT  8772.5 22030.0 8907.5 22100.0 ;
      RECT  10982.5 23375.0 11117.5 23445.0 ;
      RECT  8497.5 23375.0 8632.5 23445.0 ;
      RECT  9872.5 17202.5 10007.5 17272.5 ;
      RECT  9597.5 17062.5 9732.5 17132.5 ;
      RECT  9322.5 16922.5 9457.5 16992.5 ;
      RECT  9047.5 18517.5 9182.5 18587.5 ;
      RECT  9597.5 18657.5 9732.5 18727.5 ;
      RECT  9322.5 18797.5 9457.5 18867.5 ;
      RECT  9872.5 19892.5 10007.5 19962.5 ;
      RECT  8772.5 19752.5 8907.5 19822.5 ;
      RECT  9322.5 19612.5 9457.5 19682.5 ;
      RECT  9047.5 21207.5 9182.5 21277.5 ;
      RECT  8772.5 21347.5 8907.5 21417.5 ;
      RECT  9322.5 21487.5 9457.5 21557.5 ;
      RECT  9872.5 22582.5 10007.5 22652.5 ;
      RECT  9597.5 22442.5 9732.5 22512.5 ;
      RECT  8497.5 22302.5 8632.5 22372.5 ;
      RECT  9047.5 23897.5 9182.5 23967.5 ;
      RECT  9597.5 24037.5 9732.5 24107.5 ;
      RECT  8497.5 24177.5 8632.5 24247.5 ;
      RECT  9872.5 25272.5 10007.5 25342.5 ;
      RECT  8772.5 25132.5 8907.5 25202.5 ;
      RECT  8497.5 24992.5 8632.5 25062.5 ;
      RECT  9047.5 26587.5 9182.5 26657.5 ;
      RECT  8772.5 26727.5 8907.5 26797.5 ;
      RECT  8497.5 26867.5 8632.5 26937.5 ;
      RECT  11635.0 16550.0 11565.0 27170.0 ;
      RECT  11360.0 16550.0 11290.0 27170.0 ;
      RECT  11085.0 16550.0 11015.0 27170.0 ;
      RECT  7010.0 27915.0 7080.0 27985.0 ;
      RECT  7200.0 27915.0 7270.0 27985.0 ;
      RECT  7010.0 27950.0 7080.0 28312.5 ;
      RECT  7045.0 27915.0 7235.0 27985.0 ;
      RECT  7200.0 27607.5 7270.0 27950.0 ;
      RECT  7010.0 28312.5 7080.0 28447.5 ;
      RECT  7200.0 27472.5 7270.0 27607.5 ;
      RECT  7302.5 27915.0 7167.5 27985.0 ;
      RECT  7010.0 29395.0 7080.0 29325.0 ;
      RECT  7200.0 29395.0 7270.0 29325.0 ;
      RECT  7010.0 29360.0 7080.0 28997.5 ;
      RECT  7045.0 29395.0 7235.0 29325.0 ;
      RECT  7200.0 29702.5 7270.0 29360.0 ;
      RECT  7010.0 28997.5 7080.0 28862.5 ;
      RECT  7200.0 29837.5 7270.0 29702.5 ;
      RECT  7302.5 29395.0 7167.5 29325.0 ;
      RECT  7010.0 30605.0 7080.0 30675.0 ;
      RECT  7200.0 30605.0 7270.0 30675.0 ;
      RECT  7010.0 30640.0 7080.0 31002.5 ;
      RECT  7045.0 30605.0 7235.0 30675.0 ;
      RECT  7200.0 30297.5 7270.0 30640.0 ;
      RECT  7010.0 31002.5 7080.0 31137.5 ;
      RECT  7200.0 30162.5 7270.0 30297.5 ;
      RECT  7302.5 30605.0 7167.5 30675.0 ;
      RECT  7010.0 32085.0 7080.0 32015.0 ;
      RECT  7200.0 32085.0 7270.0 32015.0 ;
      RECT  7010.0 32050.0 7080.0 31687.5 ;
      RECT  7045.0 32085.0 7235.0 32015.0 ;
      RECT  7200.0 32392.5 7270.0 32050.0 ;
      RECT  7010.0 31687.5 7080.0 31552.5 ;
      RECT  7200.0 32527.5 7270.0 32392.5 ;
      RECT  7302.5 32085.0 7167.5 32015.0 ;
      RECT  7010.0 33295.0 7080.0 33365.0 ;
      RECT  7200.0 33295.0 7270.0 33365.0 ;
      RECT  7010.0 33330.0 7080.0 33692.5 ;
      RECT  7045.0 33295.0 7235.0 33365.0 ;
      RECT  7200.0 32987.5 7270.0 33330.0 ;
      RECT  7010.0 33692.5 7080.0 33827.5 ;
      RECT  7200.0 32852.5 7270.0 32987.5 ;
      RECT  7302.5 33295.0 7167.5 33365.0 ;
      RECT  7010.0 34775.0 7080.0 34705.0 ;
      RECT  7200.0 34775.0 7270.0 34705.0 ;
      RECT  7010.0 34740.0 7080.0 34377.5 ;
      RECT  7045.0 34775.0 7235.0 34705.0 ;
      RECT  7200.0 35082.5 7270.0 34740.0 ;
      RECT  7010.0 34377.5 7080.0 34242.5 ;
      RECT  7200.0 35217.5 7270.0 35082.5 ;
      RECT  7302.5 34775.0 7167.5 34705.0 ;
      RECT  7010.0 35985.0 7080.0 36055.0 ;
      RECT  7200.0 35985.0 7270.0 36055.0 ;
      RECT  7010.0 36020.0 7080.0 36382.5 ;
      RECT  7045.0 35985.0 7235.0 36055.0 ;
      RECT  7200.0 35677.5 7270.0 36020.0 ;
      RECT  7010.0 36382.5 7080.0 36517.5 ;
      RECT  7200.0 35542.5 7270.0 35677.5 ;
      RECT  7302.5 35985.0 7167.5 36055.0 ;
      RECT  7010.0 37465.0 7080.0 37395.0 ;
      RECT  7200.0 37465.0 7270.0 37395.0 ;
      RECT  7010.0 37430.0 7080.0 37067.5 ;
      RECT  7045.0 37465.0 7235.0 37395.0 ;
      RECT  7200.0 37772.5 7270.0 37430.0 ;
      RECT  7010.0 37067.5 7080.0 36932.5 ;
      RECT  7200.0 37907.5 7270.0 37772.5 ;
      RECT  7302.5 37465.0 7167.5 37395.0 ;
      RECT  7010.0 38675.0 7080.0 38745.0 ;
      RECT  7200.0 38675.0 7270.0 38745.0 ;
      RECT  7010.0 38710.0 7080.0 39072.5 ;
      RECT  7045.0 38675.0 7235.0 38745.0 ;
      RECT  7200.0 38367.5 7270.0 38710.0 ;
      RECT  7010.0 39072.5 7080.0 39207.5 ;
      RECT  7200.0 38232.5 7270.0 38367.5 ;
      RECT  7302.5 38675.0 7167.5 38745.0 ;
      RECT  7010.0 40155.0 7080.0 40085.0 ;
      RECT  7200.0 40155.0 7270.0 40085.0 ;
      RECT  7010.0 40120.0 7080.0 39757.5 ;
      RECT  7045.0 40155.0 7235.0 40085.0 ;
      RECT  7200.0 40462.5 7270.0 40120.0 ;
      RECT  7010.0 39757.5 7080.0 39622.5 ;
      RECT  7200.0 40597.5 7270.0 40462.5 ;
      RECT  7302.5 40155.0 7167.5 40085.0 ;
      RECT  7010.0 41365.0 7080.0 41435.0 ;
      RECT  7200.0 41365.0 7270.0 41435.0 ;
      RECT  7010.0 41400.0 7080.0 41762.5 ;
      RECT  7045.0 41365.0 7235.0 41435.0 ;
      RECT  7200.0 41057.5 7270.0 41400.0 ;
      RECT  7010.0 41762.5 7080.0 41897.5 ;
      RECT  7200.0 40922.5 7270.0 41057.5 ;
      RECT  7302.5 41365.0 7167.5 41435.0 ;
      RECT  7010.0 42845.0 7080.0 42775.0 ;
      RECT  7200.0 42845.0 7270.0 42775.0 ;
      RECT  7010.0 42810.0 7080.0 42447.5 ;
      RECT  7045.0 42845.0 7235.0 42775.0 ;
      RECT  7200.0 43152.5 7270.0 42810.0 ;
      RECT  7010.0 42447.5 7080.0 42312.5 ;
      RECT  7200.0 43287.5 7270.0 43152.5 ;
      RECT  7302.5 42845.0 7167.5 42775.0 ;
      RECT  7010.0 44055.0 7080.0 44125.0 ;
      RECT  7200.0 44055.0 7270.0 44125.0 ;
      RECT  7010.0 44090.0 7080.0 44452.5 ;
      RECT  7045.0 44055.0 7235.0 44125.0 ;
      RECT  7200.0 43747.5 7270.0 44090.0 ;
      RECT  7010.0 44452.5 7080.0 44587.5 ;
      RECT  7200.0 43612.5 7270.0 43747.5 ;
      RECT  7302.5 44055.0 7167.5 44125.0 ;
      RECT  7010.0 45535.0 7080.0 45465.0 ;
      RECT  7200.0 45535.0 7270.0 45465.0 ;
      RECT  7010.0 45500.0 7080.0 45137.5 ;
      RECT  7045.0 45535.0 7235.0 45465.0 ;
      RECT  7200.0 45842.5 7270.0 45500.0 ;
      RECT  7010.0 45137.5 7080.0 45002.5 ;
      RECT  7200.0 45977.5 7270.0 45842.5 ;
      RECT  7302.5 45535.0 7167.5 45465.0 ;
      RECT  7010.0 46745.0 7080.0 46815.0 ;
      RECT  7200.0 46745.0 7270.0 46815.0 ;
      RECT  7010.0 46780.0 7080.0 47142.5 ;
      RECT  7045.0 46745.0 7235.0 46815.0 ;
      RECT  7200.0 46437.5 7270.0 46780.0 ;
      RECT  7010.0 47142.5 7080.0 47277.5 ;
      RECT  7200.0 46302.5 7270.0 46437.5 ;
      RECT  7302.5 46745.0 7167.5 46815.0 ;
      RECT  7010.0 48225.0 7080.0 48155.0 ;
      RECT  7200.0 48225.0 7270.0 48155.0 ;
      RECT  7010.0 48190.0 7080.0 47827.5 ;
      RECT  7045.0 48225.0 7235.0 48155.0 ;
      RECT  7200.0 48532.5 7270.0 48190.0 ;
      RECT  7010.0 47827.5 7080.0 47692.5 ;
      RECT  7200.0 48667.5 7270.0 48532.5 ;
      RECT  7302.5 48225.0 7167.5 48155.0 ;
      RECT  7010.0 49435.0 7080.0 49505.0 ;
      RECT  7200.0 49435.0 7270.0 49505.0 ;
      RECT  7010.0 49470.0 7080.0 49832.5 ;
      RECT  7045.0 49435.0 7235.0 49505.0 ;
      RECT  7200.0 49127.5 7270.0 49470.0 ;
      RECT  7010.0 49832.5 7080.0 49967.5 ;
      RECT  7200.0 48992.5 7270.0 49127.5 ;
      RECT  7302.5 49435.0 7167.5 49505.0 ;
      RECT  7010.0 50915.0 7080.0 50845.0 ;
      RECT  7200.0 50915.0 7270.0 50845.0 ;
      RECT  7010.0 50880.0 7080.0 50517.5 ;
      RECT  7045.0 50915.0 7235.0 50845.0 ;
      RECT  7200.0 51222.5 7270.0 50880.0 ;
      RECT  7010.0 50517.5 7080.0 50382.5 ;
      RECT  7200.0 51357.5 7270.0 51222.5 ;
      RECT  7302.5 50915.0 7167.5 50845.0 ;
      RECT  7010.0 52125.0 7080.0 52195.0 ;
      RECT  7200.0 52125.0 7270.0 52195.0 ;
      RECT  7010.0 52160.0 7080.0 52522.5 ;
      RECT  7045.0 52125.0 7235.0 52195.0 ;
      RECT  7200.0 51817.5 7270.0 52160.0 ;
      RECT  7010.0 52522.5 7080.0 52657.5 ;
      RECT  7200.0 51682.5 7270.0 51817.5 ;
      RECT  7302.5 52125.0 7167.5 52195.0 ;
      RECT  7010.0 53605.0 7080.0 53535.0 ;
      RECT  7200.0 53605.0 7270.0 53535.0 ;
      RECT  7010.0 53570.0 7080.0 53207.5 ;
      RECT  7045.0 53605.0 7235.0 53535.0 ;
      RECT  7200.0 53912.5 7270.0 53570.0 ;
      RECT  7010.0 53207.5 7080.0 53072.5 ;
      RECT  7200.0 54047.5 7270.0 53912.5 ;
      RECT  7302.5 53605.0 7167.5 53535.0 ;
      RECT  7010.0 54815.0 7080.0 54885.0 ;
      RECT  7200.0 54815.0 7270.0 54885.0 ;
      RECT  7010.0 54850.0 7080.0 55212.5 ;
      RECT  7045.0 54815.0 7235.0 54885.0 ;
      RECT  7200.0 54507.5 7270.0 54850.0 ;
      RECT  7010.0 55212.5 7080.0 55347.5 ;
      RECT  7200.0 54372.5 7270.0 54507.5 ;
      RECT  7302.5 54815.0 7167.5 54885.0 ;
      RECT  7010.0 56295.0 7080.0 56225.0 ;
      RECT  7200.0 56295.0 7270.0 56225.0 ;
      RECT  7010.0 56260.0 7080.0 55897.5 ;
      RECT  7045.0 56295.0 7235.0 56225.0 ;
      RECT  7200.0 56602.5 7270.0 56260.0 ;
      RECT  7010.0 55897.5 7080.0 55762.5 ;
      RECT  7200.0 56737.5 7270.0 56602.5 ;
      RECT  7302.5 56295.0 7167.5 56225.0 ;
      RECT  7010.0 57505.0 7080.0 57575.0 ;
      RECT  7200.0 57505.0 7270.0 57575.0 ;
      RECT  7010.0 57540.0 7080.0 57902.5 ;
      RECT  7045.0 57505.0 7235.0 57575.0 ;
      RECT  7200.0 57197.5 7270.0 57540.0 ;
      RECT  7010.0 57902.5 7080.0 58037.5 ;
      RECT  7200.0 57062.5 7270.0 57197.5 ;
      RECT  7302.5 57505.0 7167.5 57575.0 ;
      RECT  7010.0 58985.0 7080.0 58915.0 ;
      RECT  7200.0 58985.0 7270.0 58915.0 ;
      RECT  7010.0 58950.0 7080.0 58587.5 ;
      RECT  7045.0 58985.0 7235.0 58915.0 ;
      RECT  7200.0 59292.5 7270.0 58950.0 ;
      RECT  7010.0 58587.5 7080.0 58452.5 ;
      RECT  7200.0 59427.5 7270.0 59292.5 ;
      RECT  7302.5 58985.0 7167.5 58915.0 ;
      RECT  7010.0 60195.0 7080.0 60265.0 ;
      RECT  7200.0 60195.0 7270.0 60265.0 ;
      RECT  7010.0 60230.0 7080.0 60592.5 ;
      RECT  7045.0 60195.0 7235.0 60265.0 ;
      RECT  7200.0 59887.5 7270.0 60230.0 ;
      RECT  7010.0 60592.5 7080.0 60727.5 ;
      RECT  7200.0 59752.5 7270.0 59887.5 ;
      RECT  7302.5 60195.0 7167.5 60265.0 ;
      RECT  7010.0 61675.0 7080.0 61605.0 ;
      RECT  7200.0 61675.0 7270.0 61605.0 ;
      RECT  7010.0 61640.0 7080.0 61277.5 ;
      RECT  7045.0 61675.0 7235.0 61605.0 ;
      RECT  7200.0 61982.5 7270.0 61640.0 ;
      RECT  7010.0 61277.5 7080.0 61142.5 ;
      RECT  7200.0 62117.5 7270.0 61982.5 ;
      RECT  7302.5 61675.0 7167.5 61605.0 ;
      RECT  7010.0 62885.0 7080.0 62955.0 ;
      RECT  7200.0 62885.0 7270.0 62955.0 ;
      RECT  7010.0 62920.0 7080.0 63282.5 ;
      RECT  7045.0 62885.0 7235.0 62955.0 ;
      RECT  7200.0 62577.5 7270.0 62920.0 ;
      RECT  7010.0 63282.5 7080.0 63417.5 ;
      RECT  7200.0 62442.5 7270.0 62577.5 ;
      RECT  7302.5 62885.0 7167.5 62955.0 ;
      RECT  7010.0 64365.0 7080.0 64295.0 ;
      RECT  7200.0 64365.0 7270.0 64295.0 ;
      RECT  7010.0 64330.0 7080.0 63967.5 ;
      RECT  7045.0 64365.0 7235.0 64295.0 ;
      RECT  7200.0 64672.5 7270.0 64330.0 ;
      RECT  7010.0 63967.5 7080.0 63832.5 ;
      RECT  7200.0 64807.5 7270.0 64672.5 ;
      RECT  7302.5 64365.0 7167.5 64295.0 ;
      RECT  7010.0 65575.0 7080.0 65645.0 ;
      RECT  7200.0 65575.0 7270.0 65645.0 ;
      RECT  7010.0 65610.0 7080.0 65972.5 ;
      RECT  7045.0 65575.0 7235.0 65645.0 ;
      RECT  7200.0 65267.5 7270.0 65610.0 ;
      RECT  7010.0 65972.5 7080.0 66107.5 ;
      RECT  7200.0 65132.5 7270.0 65267.5 ;
      RECT  7302.5 65575.0 7167.5 65645.0 ;
      RECT  7010.0 67055.0 7080.0 66985.0 ;
      RECT  7200.0 67055.0 7270.0 66985.0 ;
      RECT  7010.0 67020.0 7080.0 66657.5 ;
      RECT  7045.0 67055.0 7235.0 66985.0 ;
      RECT  7200.0 67362.5 7270.0 67020.0 ;
      RECT  7010.0 66657.5 7080.0 66522.5 ;
      RECT  7200.0 67497.5 7270.0 67362.5 ;
      RECT  7302.5 67055.0 7167.5 66985.0 ;
      RECT  7010.0 68265.0 7080.0 68335.0 ;
      RECT  7200.0 68265.0 7270.0 68335.0 ;
      RECT  7010.0 68300.0 7080.0 68662.5 ;
      RECT  7045.0 68265.0 7235.0 68335.0 ;
      RECT  7200.0 67957.5 7270.0 68300.0 ;
      RECT  7010.0 68662.5 7080.0 68797.5 ;
      RECT  7200.0 67822.5 7270.0 67957.5 ;
      RECT  7302.5 68265.0 7167.5 68335.0 ;
      RECT  7010.0 69745.0 7080.0 69675.0 ;
      RECT  7200.0 69745.0 7270.0 69675.0 ;
      RECT  7010.0 69710.0 7080.0 69347.5 ;
      RECT  7045.0 69745.0 7235.0 69675.0 ;
      RECT  7200.0 70052.5 7270.0 69710.0 ;
      RECT  7010.0 69347.5 7080.0 69212.5 ;
      RECT  7200.0 70187.5 7270.0 70052.5 ;
      RECT  7302.5 69745.0 7167.5 69675.0 ;
      RECT  4757.5 11762.5 4622.5 11832.5 ;
      RECT  4932.5 13197.5 4797.5 13267.5 ;
      RECT  5107.5 14452.5 4972.5 14522.5 ;
      RECT  5282.5 15887.5 5147.5 15957.5 ;
      RECT  5457.5 17142.5 5322.5 17212.5 ;
      RECT  5632.5 18577.5 5497.5 18647.5 ;
      RECT  5807.5 19832.5 5672.5 19902.5 ;
      RECT  5982.5 21267.5 5847.5 21337.5 ;
      RECT  6157.5 22522.5 6022.5 22592.5 ;
      RECT  6332.5 23957.5 6197.5 24027.5 ;
      RECT  6507.5 25212.5 6372.5 25282.5 ;
      RECT  6682.5 26647.5 6547.5 26717.5 ;
      RECT  4757.5 27915.0 4622.5 27985.0 ;
      RECT  5457.5 27700.0 5322.5 27770.0 ;
      RECT  4757.5 29325.0 4622.5 29395.0 ;
      RECT  5632.5 29540.0 5497.5 29610.0 ;
      RECT  4757.5 30605.0 4622.5 30675.0 ;
      RECT  5807.5 30390.0 5672.5 30460.0 ;
      RECT  4757.5 32015.0 4622.5 32085.0 ;
      RECT  5982.5 32230.0 5847.5 32300.0 ;
      RECT  4757.5 33295.0 4622.5 33365.0 ;
      RECT  6157.5 33080.0 6022.5 33150.0 ;
      RECT  4757.5 34705.0 4622.5 34775.0 ;
      RECT  6332.5 34920.0 6197.5 34990.0 ;
      RECT  4757.5 35985.0 4622.5 36055.0 ;
      RECT  6507.5 35770.0 6372.5 35840.0 ;
      RECT  4757.5 37395.0 4622.5 37465.0 ;
      RECT  6682.5 37610.0 6547.5 37680.0 ;
      RECT  4932.5 38675.0 4797.5 38745.0 ;
      RECT  5457.5 38460.0 5322.5 38530.0 ;
      RECT  4932.5 40085.0 4797.5 40155.0 ;
      RECT  5632.5 40300.0 5497.5 40370.0 ;
      RECT  4932.5 41365.0 4797.5 41435.0 ;
      RECT  5807.5 41150.0 5672.5 41220.0 ;
      RECT  4932.5 42775.0 4797.5 42845.0 ;
      RECT  5982.5 42990.0 5847.5 43060.0 ;
      RECT  4932.5 44055.0 4797.5 44125.0 ;
      RECT  6157.5 43840.0 6022.5 43910.0 ;
      RECT  4932.5 45465.0 4797.5 45535.0 ;
      RECT  6332.5 45680.0 6197.5 45750.0 ;
      RECT  4932.5 46745.0 4797.5 46815.0 ;
      RECT  6507.5 46530.0 6372.5 46600.0 ;
      RECT  4932.5 48155.0 4797.5 48225.0 ;
      RECT  6682.5 48370.0 6547.5 48440.0 ;
      RECT  5107.5 49435.0 4972.5 49505.0 ;
      RECT  5457.5 49220.0 5322.5 49290.0 ;
      RECT  5107.5 50845.0 4972.5 50915.0 ;
      RECT  5632.5 51060.0 5497.5 51130.0 ;
      RECT  5107.5 52125.0 4972.5 52195.0 ;
      RECT  5807.5 51910.0 5672.5 51980.0 ;
      RECT  5107.5 53535.0 4972.5 53605.0 ;
      RECT  5982.5 53750.0 5847.5 53820.0 ;
      RECT  5107.5 54815.0 4972.5 54885.0 ;
      RECT  6157.5 54600.0 6022.5 54670.0 ;
      RECT  5107.5 56225.0 4972.5 56295.0 ;
      RECT  6332.5 56440.0 6197.5 56510.0 ;
      RECT  5107.5 57505.0 4972.5 57575.0 ;
      RECT  6507.5 57290.0 6372.5 57360.0 ;
      RECT  5107.5 58915.0 4972.5 58985.0 ;
      RECT  6682.5 59130.0 6547.5 59200.0 ;
      RECT  5282.5 60195.0 5147.5 60265.0 ;
      RECT  5457.5 59980.0 5322.5 60050.0 ;
      RECT  5282.5 61605.0 5147.5 61675.0 ;
      RECT  5632.5 61820.0 5497.5 61890.0 ;
      RECT  5282.5 62885.0 5147.5 62955.0 ;
      RECT  5807.5 62670.0 5672.5 62740.0 ;
      RECT  5282.5 64295.0 5147.5 64365.0 ;
      RECT  5982.5 64510.0 5847.5 64580.0 ;
      RECT  5282.5 65575.0 5147.5 65645.0 ;
      RECT  6157.5 65360.0 6022.5 65430.0 ;
      RECT  5282.5 66985.0 5147.5 67055.0 ;
      RECT  6332.5 67200.0 6197.5 67270.0 ;
      RECT  5282.5 68265.0 5147.5 68335.0 ;
      RECT  6507.5 68050.0 6372.5 68120.0 ;
      RECT  5282.5 69675.0 5147.5 69745.0 ;
      RECT  6682.5 69890.0 6547.5 69960.0 ;
      RECT  10650.0 11170.0 10720.0 16410.0 ;
      RECT  10375.0 11170.0 10445.0 16410.0 ;
      RECT  11565.0 16550.0 11635.0 27170.0 ;
      RECT  11290.0 16550.0 11360.0 27170.0 ;
      RECT  11015.0 16550.0 11085.0 27170.0 ;
      RECT  8570.0 27700.0 8640.0 27770.0 ;
      RECT  8570.0 27665.0 8640.0 27735.0 ;
      RECT  8605.0 27700.0 9567.5 27770.0 ;
      RECT  8570.0 29540.0 8640.0 29610.0 ;
      RECT  8570.0 29575.0 8640.0 29645.0 ;
      RECT  8605.0 29540.0 9567.5 29610.0 ;
      RECT  8570.0 30390.0 8640.0 30460.0 ;
      RECT  8570.0 30355.0 8640.0 30425.0 ;
      RECT  8605.0 30390.0 9567.5 30460.0 ;
      RECT  8570.0 32230.0 8640.0 32300.0 ;
      RECT  8570.0 32265.0 8640.0 32335.0 ;
      RECT  8605.0 32230.0 9567.5 32300.0 ;
      RECT  8570.0 33080.0 8640.0 33150.0 ;
      RECT  8570.0 33045.0 8640.0 33115.0 ;
      RECT  8605.0 33080.0 9567.5 33150.0 ;
      RECT  8570.0 34920.0 8640.0 34990.0 ;
      RECT  8570.0 34955.0 8640.0 35025.0 ;
      RECT  8605.0 34920.0 9567.5 34990.0 ;
      RECT  8570.0 35770.0 8640.0 35840.0 ;
      RECT  8570.0 35735.0 8640.0 35805.0 ;
      RECT  8605.0 35770.0 9567.5 35840.0 ;
      RECT  8570.0 37610.0 8640.0 37680.0 ;
      RECT  8570.0 37645.0 8640.0 37715.0 ;
      RECT  8605.0 37610.0 9567.5 37680.0 ;
      RECT  8570.0 38460.0 8640.0 38530.0 ;
      RECT  8570.0 38425.0 8640.0 38495.0 ;
      RECT  8605.0 38460.0 9567.5 38530.0 ;
      RECT  8570.0 40300.0 8640.0 40370.0 ;
      RECT  8570.0 40335.0 8640.0 40405.0 ;
      RECT  8605.0 40300.0 9567.5 40370.0 ;
      RECT  8570.0 41150.0 8640.0 41220.0 ;
      RECT  8570.0 41115.0 8640.0 41185.0 ;
      RECT  8605.0 41150.0 9567.5 41220.0 ;
      RECT  8570.0 42990.0 8640.0 43060.0 ;
      RECT  8570.0 43025.0 8640.0 43095.0 ;
      RECT  8605.0 42990.0 9567.5 43060.0 ;
      RECT  8570.0 43840.0 8640.0 43910.0 ;
      RECT  8570.0 43805.0 8640.0 43875.0 ;
      RECT  8605.0 43840.0 9567.5 43910.0 ;
      RECT  8570.0 45680.0 8640.0 45750.0 ;
      RECT  8570.0 45715.0 8640.0 45785.0 ;
      RECT  8605.0 45680.0 9567.5 45750.0 ;
      RECT  8570.0 46530.0 8640.0 46600.0 ;
      RECT  8570.0 46495.0 8640.0 46565.0 ;
      RECT  8605.0 46530.0 9567.5 46600.0 ;
      RECT  8570.0 48370.0 8640.0 48440.0 ;
      RECT  8570.0 48405.0 8640.0 48475.0 ;
      RECT  8605.0 48370.0 9567.5 48440.0 ;
      RECT  8570.0 49220.0 8640.0 49290.0 ;
      RECT  8570.0 49185.0 8640.0 49255.0 ;
      RECT  8605.0 49220.0 9567.5 49290.0 ;
      RECT  8570.0 51060.0 8640.0 51130.0 ;
      RECT  8570.0 51095.0 8640.0 51165.0 ;
      RECT  8605.0 51060.0 9567.5 51130.0 ;
      RECT  8570.0 51910.0 8640.0 51980.0 ;
      RECT  8570.0 51875.0 8640.0 51945.0 ;
      RECT  8605.0 51910.0 9567.5 51980.0 ;
      RECT  8570.0 53750.0 8640.0 53820.0 ;
      RECT  8570.0 53785.0 8640.0 53855.0 ;
      RECT  8605.0 53750.0 9567.5 53820.0 ;
      RECT  8570.0 54600.0 8640.0 54670.0 ;
      RECT  8570.0 54565.0 8640.0 54635.0 ;
      RECT  8605.0 54600.0 9567.5 54670.0 ;
      RECT  8570.0 56440.0 8640.0 56510.0 ;
      RECT  8570.0 56475.0 8640.0 56545.0 ;
      RECT  8605.0 56440.0 9567.5 56510.0 ;
      RECT  8570.0 57290.0 8640.0 57360.0 ;
      RECT  8570.0 57255.0 8640.0 57325.0 ;
      RECT  8605.0 57290.0 9567.5 57360.0 ;
      RECT  8570.0 59130.0 8640.0 59200.0 ;
      RECT  8570.0 59165.0 8640.0 59235.0 ;
      RECT  8605.0 59130.0 9567.5 59200.0 ;
      RECT  8570.0 59980.0 8640.0 60050.0 ;
      RECT  8570.0 59945.0 8640.0 60015.0 ;
      RECT  8605.0 59980.0 9567.5 60050.0 ;
      RECT  8570.0 61820.0 8640.0 61890.0 ;
      RECT  8570.0 61855.0 8640.0 61925.0 ;
      RECT  8605.0 61820.0 9567.5 61890.0 ;
      RECT  8570.0 62670.0 8640.0 62740.0 ;
      RECT  8570.0 62635.0 8640.0 62705.0 ;
      RECT  8605.0 62670.0 9567.5 62740.0 ;
      RECT  8570.0 64510.0 8640.0 64580.0 ;
      RECT  8570.0 64545.0 8640.0 64615.0 ;
      RECT  8605.0 64510.0 9567.5 64580.0 ;
      RECT  8570.0 65360.0 8640.0 65430.0 ;
      RECT  8570.0 65325.0 8640.0 65395.0 ;
      RECT  8605.0 65360.0 9567.5 65430.0 ;
      RECT  8570.0 67200.0 8640.0 67270.0 ;
      RECT  8570.0 67235.0 8640.0 67305.0 ;
      RECT  8605.0 67200.0 9567.5 67270.0 ;
      RECT  8570.0 68050.0 8640.0 68120.0 ;
      RECT  8570.0 68015.0 8640.0 68085.0 ;
      RECT  8605.0 68050.0 9567.5 68120.0 ;
      RECT  8570.0 69890.0 8640.0 69960.0 ;
      RECT  8570.0 69925.0 8640.0 69995.0 ;
      RECT  8605.0 69890.0 9567.5 69960.0 ;
      RECT  9505.0 27915.0 9575.0 27985.0 ;
      RECT  9695.0 27915.0 9765.0 27985.0 ;
      RECT  9505.0 27950.0 9575.0 28312.5 ;
      RECT  9540.0 27915.0 9730.0 27985.0 ;
      RECT  9695.0 27607.5 9765.0 27950.0 ;
      RECT  9505.0 28312.5 9575.0 28447.5 ;
      RECT  9695.0 27472.5 9765.0 27607.5 ;
      RECT  9797.5 27915.0 9662.5 27985.0 ;
      RECT  8430.0 27870.0 8500.0 28005.0 ;
      RECT  8570.0 27597.5 8640.0 27732.5 ;
      RECT  9567.5 27700.0 9432.5 27770.0 ;
      RECT  9505.0 29395.0 9575.0 29325.0 ;
      RECT  9695.0 29395.0 9765.0 29325.0 ;
      RECT  9505.0 29360.0 9575.0 28997.5 ;
      RECT  9540.0 29395.0 9730.0 29325.0 ;
      RECT  9695.0 29702.5 9765.0 29360.0 ;
      RECT  9505.0 28997.5 9575.0 28862.5 ;
      RECT  9695.0 29837.5 9765.0 29702.5 ;
      RECT  9797.5 29395.0 9662.5 29325.0 ;
      RECT  8430.0 29305.0 8500.0 29440.0 ;
      RECT  8570.0 29577.5 8640.0 29712.5 ;
      RECT  9567.5 29540.0 9432.5 29610.0 ;
      RECT  9505.0 30605.0 9575.0 30675.0 ;
      RECT  9695.0 30605.0 9765.0 30675.0 ;
      RECT  9505.0 30640.0 9575.0 31002.5 ;
      RECT  9540.0 30605.0 9730.0 30675.0 ;
      RECT  9695.0 30297.5 9765.0 30640.0 ;
      RECT  9505.0 31002.5 9575.0 31137.5 ;
      RECT  9695.0 30162.5 9765.0 30297.5 ;
      RECT  9797.5 30605.0 9662.5 30675.0 ;
      RECT  8430.0 30560.0 8500.0 30695.0 ;
      RECT  8570.0 30287.5 8640.0 30422.5 ;
      RECT  9567.5 30390.0 9432.5 30460.0 ;
      RECT  9505.0 32085.0 9575.0 32015.0 ;
      RECT  9695.0 32085.0 9765.0 32015.0 ;
      RECT  9505.0 32050.0 9575.0 31687.5 ;
      RECT  9540.0 32085.0 9730.0 32015.0 ;
      RECT  9695.0 32392.5 9765.0 32050.0 ;
      RECT  9505.0 31687.5 9575.0 31552.5 ;
      RECT  9695.0 32527.5 9765.0 32392.5 ;
      RECT  9797.5 32085.0 9662.5 32015.0 ;
      RECT  8430.0 31995.0 8500.0 32130.0 ;
      RECT  8570.0 32267.5 8640.0 32402.5 ;
      RECT  9567.5 32230.0 9432.5 32300.0 ;
      RECT  9505.0 33295.0 9575.0 33365.0 ;
      RECT  9695.0 33295.0 9765.0 33365.0 ;
      RECT  9505.0 33330.0 9575.0 33692.5 ;
      RECT  9540.0 33295.0 9730.0 33365.0 ;
      RECT  9695.0 32987.5 9765.0 33330.0 ;
      RECT  9505.0 33692.5 9575.0 33827.5 ;
      RECT  9695.0 32852.5 9765.0 32987.5 ;
      RECT  9797.5 33295.0 9662.5 33365.0 ;
      RECT  8430.0 33250.0 8500.0 33385.0 ;
      RECT  8570.0 32977.5 8640.0 33112.5 ;
      RECT  9567.5 33080.0 9432.5 33150.0 ;
      RECT  9505.0 34775.0 9575.0 34705.0 ;
      RECT  9695.0 34775.0 9765.0 34705.0 ;
      RECT  9505.0 34740.0 9575.0 34377.5 ;
      RECT  9540.0 34775.0 9730.0 34705.0 ;
      RECT  9695.0 35082.5 9765.0 34740.0 ;
      RECT  9505.0 34377.5 9575.0 34242.5 ;
      RECT  9695.0 35217.5 9765.0 35082.5 ;
      RECT  9797.5 34775.0 9662.5 34705.0 ;
      RECT  8430.0 34685.0 8500.0 34820.0 ;
      RECT  8570.0 34957.5 8640.0 35092.5 ;
      RECT  9567.5 34920.0 9432.5 34990.0 ;
      RECT  9505.0 35985.0 9575.0 36055.0 ;
      RECT  9695.0 35985.0 9765.0 36055.0 ;
      RECT  9505.0 36020.0 9575.0 36382.5 ;
      RECT  9540.0 35985.0 9730.0 36055.0 ;
      RECT  9695.0 35677.5 9765.0 36020.0 ;
      RECT  9505.0 36382.5 9575.0 36517.5 ;
      RECT  9695.0 35542.5 9765.0 35677.5 ;
      RECT  9797.5 35985.0 9662.5 36055.0 ;
      RECT  8430.0 35940.0 8500.0 36075.0 ;
      RECT  8570.0 35667.5 8640.0 35802.5 ;
      RECT  9567.5 35770.0 9432.5 35840.0 ;
      RECT  9505.0 37465.0 9575.0 37395.0 ;
      RECT  9695.0 37465.0 9765.0 37395.0 ;
      RECT  9505.0 37430.0 9575.0 37067.5 ;
      RECT  9540.0 37465.0 9730.0 37395.0 ;
      RECT  9695.0 37772.5 9765.0 37430.0 ;
      RECT  9505.0 37067.5 9575.0 36932.5 ;
      RECT  9695.0 37907.5 9765.0 37772.5 ;
      RECT  9797.5 37465.0 9662.5 37395.0 ;
      RECT  8430.0 37375.0 8500.0 37510.0 ;
      RECT  8570.0 37647.5 8640.0 37782.5 ;
      RECT  9567.5 37610.0 9432.5 37680.0 ;
      RECT  9505.0 38675.0 9575.0 38745.0 ;
      RECT  9695.0 38675.0 9765.0 38745.0 ;
      RECT  9505.0 38710.0 9575.0 39072.5 ;
      RECT  9540.0 38675.0 9730.0 38745.0 ;
      RECT  9695.0 38367.5 9765.0 38710.0 ;
      RECT  9505.0 39072.5 9575.0 39207.5 ;
      RECT  9695.0 38232.5 9765.0 38367.5 ;
      RECT  9797.5 38675.0 9662.5 38745.0 ;
      RECT  8430.0 38630.0 8500.0 38765.0 ;
      RECT  8570.0 38357.5 8640.0 38492.5 ;
      RECT  9567.5 38460.0 9432.5 38530.0 ;
      RECT  9505.0 40155.0 9575.0 40085.0 ;
      RECT  9695.0 40155.0 9765.0 40085.0 ;
      RECT  9505.0 40120.0 9575.0 39757.5 ;
      RECT  9540.0 40155.0 9730.0 40085.0 ;
      RECT  9695.0 40462.5 9765.0 40120.0 ;
      RECT  9505.0 39757.5 9575.0 39622.5 ;
      RECT  9695.0 40597.5 9765.0 40462.5 ;
      RECT  9797.5 40155.0 9662.5 40085.0 ;
      RECT  8430.0 40065.0 8500.0 40200.0 ;
      RECT  8570.0 40337.5 8640.0 40472.5 ;
      RECT  9567.5 40300.0 9432.5 40370.0 ;
      RECT  9505.0 41365.0 9575.0 41435.0 ;
      RECT  9695.0 41365.0 9765.0 41435.0 ;
      RECT  9505.0 41400.0 9575.0 41762.5 ;
      RECT  9540.0 41365.0 9730.0 41435.0 ;
      RECT  9695.0 41057.5 9765.0 41400.0 ;
      RECT  9505.0 41762.5 9575.0 41897.5 ;
      RECT  9695.0 40922.5 9765.0 41057.5 ;
      RECT  9797.5 41365.0 9662.5 41435.0 ;
      RECT  8430.0 41320.0 8500.0 41455.0 ;
      RECT  8570.0 41047.5 8640.0 41182.5 ;
      RECT  9567.5 41150.0 9432.5 41220.0 ;
      RECT  9505.0 42845.0 9575.0 42775.0 ;
      RECT  9695.0 42845.0 9765.0 42775.0 ;
      RECT  9505.0 42810.0 9575.0 42447.5 ;
      RECT  9540.0 42845.0 9730.0 42775.0 ;
      RECT  9695.0 43152.5 9765.0 42810.0 ;
      RECT  9505.0 42447.5 9575.0 42312.5 ;
      RECT  9695.0 43287.5 9765.0 43152.5 ;
      RECT  9797.5 42845.0 9662.5 42775.0 ;
      RECT  8430.0 42755.0 8500.0 42890.0 ;
      RECT  8570.0 43027.5 8640.0 43162.5 ;
      RECT  9567.5 42990.0 9432.5 43060.0 ;
      RECT  9505.0 44055.0 9575.0 44125.0 ;
      RECT  9695.0 44055.0 9765.0 44125.0 ;
      RECT  9505.0 44090.0 9575.0 44452.5 ;
      RECT  9540.0 44055.0 9730.0 44125.0 ;
      RECT  9695.0 43747.5 9765.0 44090.0 ;
      RECT  9505.0 44452.5 9575.0 44587.5 ;
      RECT  9695.0 43612.5 9765.0 43747.5 ;
      RECT  9797.5 44055.0 9662.5 44125.0 ;
      RECT  8430.0 44010.0 8500.0 44145.0 ;
      RECT  8570.0 43737.5 8640.0 43872.5 ;
      RECT  9567.5 43840.0 9432.5 43910.0 ;
      RECT  9505.0 45535.0 9575.0 45465.0 ;
      RECT  9695.0 45535.0 9765.0 45465.0 ;
      RECT  9505.0 45500.0 9575.0 45137.5 ;
      RECT  9540.0 45535.0 9730.0 45465.0 ;
      RECT  9695.0 45842.5 9765.0 45500.0 ;
      RECT  9505.0 45137.5 9575.0 45002.5 ;
      RECT  9695.0 45977.5 9765.0 45842.5 ;
      RECT  9797.5 45535.0 9662.5 45465.0 ;
      RECT  8430.0 45445.0 8500.0 45580.0 ;
      RECT  8570.0 45717.5 8640.0 45852.5 ;
      RECT  9567.5 45680.0 9432.5 45750.0 ;
      RECT  9505.0 46745.0 9575.0 46815.0 ;
      RECT  9695.0 46745.0 9765.0 46815.0 ;
      RECT  9505.0 46780.0 9575.0 47142.5 ;
      RECT  9540.0 46745.0 9730.0 46815.0 ;
      RECT  9695.0 46437.5 9765.0 46780.0 ;
      RECT  9505.0 47142.5 9575.0 47277.5 ;
      RECT  9695.0 46302.5 9765.0 46437.5 ;
      RECT  9797.5 46745.0 9662.5 46815.0 ;
      RECT  8430.0 46700.0 8500.0 46835.0 ;
      RECT  8570.0 46427.5 8640.0 46562.5 ;
      RECT  9567.5 46530.0 9432.5 46600.0 ;
      RECT  9505.0 48225.0 9575.0 48155.0 ;
      RECT  9695.0 48225.0 9765.0 48155.0 ;
      RECT  9505.0 48190.0 9575.0 47827.5 ;
      RECT  9540.0 48225.0 9730.0 48155.0 ;
      RECT  9695.0 48532.5 9765.0 48190.0 ;
      RECT  9505.0 47827.5 9575.0 47692.5 ;
      RECT  9695.0 48667.5 9765.0 48532.5 ;
      RECT  9797.5 48225.0 9662.5 48155.0 ;
      RECT  8430.0 48135.0 8500.0 48270.0 ;
      RECT  8570.0 48407.5 8640.0 48542.5 ;
      RECT  9567.5 48370.0 9432.5 48440.0 ;
      RECT  9505.0 49435.0 9575.0 49505.0 ;
      RECT  9695.0 49435.0 9765.0 49505.0 ;
      RECT  9505.0 49470.0 9575.0 49832.5 ;
      RECT  9540.0 49435.0 9730.0 49505.0 ;
      RECT  9695.0 49127.5 9765.0 49470.0 ;
      RECT  9505.0 49832.5 9575.0 49967.5 ;
      RECT  9695.0 48992.5 9765.0 49127.5 ;
      RECT  9797.5 49435.0 9662.5 49505.0 ;
      RECT  8430.0 49390.0 8500.0 49525.0 ;
      RECT  8570.0 49117.5 8640.0 49252.5 ;
      RECT  9567.5 49220.0 9432.5 49290.0 ;
      RECT  9505.0 50915.0 9575.0 50845.0 ;
      RECT  9695.0 50915.0 9765.0 50845.0 ;
      RECT  9505.0 50880.0 9575.0 50517.5 ;
      RECT  9540.0 50915.0 9730.0 50845.0 ;
      RECT  9695.0 51222.5 9765.0 50880.0 ;
      RECT  9505.0 50517.5 9575.0 50382.5 ;
      RECT  9695.0 51357.5 9765.0 51222.5 ;
      RECT  9797.5 50915.0 9662.5 50845.0 ;
      RECT  8430.0 50825.0 8500.0 50960.0 ;
      RECT  8570.0 51097.5 8640.0 51232.5 ;
      RECT  9567.5 51060.0 9432.5 51130.0 ;
      RECT  9505.0 52125.0 9575.0 52195.0 ;
      RECT  9695.0 52125.0 9765.0 52195.0 ;
      RECT  9505.0 52160.0 9575.0 52522.5 ;
      RECT  9540.0 52125.0 9730.0 52195.0 ;
      RECT  9695.0 51817.5 9765.0 52160.0 ;
      RECT  9505.0 52522.5 9575.0 52657.5 ;
      RECT  9695.0 51682.5 9765.0 51817.5 ;
      RECT  9797.5 52125.0 9662.5 52195.0 ;
      RECT  8430.0 52080.0 8500.0 52215.0 ;
      RECT  8570.0 51807.5 8640.0 51942.5 ;
      RECT  9567.5 51910.0 9432.5 51980.0 ;
      RECT  9505.0 53605.0 9575.0 53535.0 ;
      RECT  9695.0 53605.0 9765.0 53535.0 ;
      RECT  9505.0 53570.0 9575.0 53207.5 ;
      RECT  9540.0 53605.0 9730.0 53535.0 ;
      RECT  9695.0 53912.5 9765.0 53570.0 ;
      RECT  9505.0 53207.5 9575.0 53072.5 ;
      RECT  9695.0 54047.5 9765.0 53912.5 ;
      RECT  9797.5 53605.0 9662.5 53535.0 ;
      RECT  8430.0 53515.0 8500.0 53650.0 ;
      RECT  8570.0 53787.5 8640.0 53922.5 ;
      RECT  9567.5 53750.0 9432.5 53820.0 ;
      RECT  9505.0 54815.0 9575.0 54885.0 ;
      RECT  9695.0 54815.0 9765.0 54885.0 ;
      RECT  9505.0 54850.0 9575.0 55212.5 ;
      RECT  9540.0 54815.0 9730.0 54885.0 ;
      RECT  9695.0 54507.5 9765.0 54850.0 ;
      RECT  9505.0 55212.5 9575.0 55347.5 ;
      RECT  9695.0 54372.5 9765.0 54507.5 ;
      RECT  9797.5 54815.0 9662.5 54885.0 ;
      RECT  8430.0 54770.0 8500.0 54905.0 ;
      RECT  8570.0 54497.5 8640.0 54632.5 ;
      RECT  9567.5 54600.0 9432.5 54670.0 ;
      RECT  9505.0 56295.0 9575.0 56225.0 ;
      RECT  9695.0 56295.0 9765.0 56225.0 ;
      RECT  9505.0 56260.0 9575.0 55897.5 ;
      RECT  9540.0 56295.0 9730.0 56225.0 ;
      RECT  9695.0 56602.5 9765.0 56260.0 ;
      RECT  9505.0 55897.5 9575.0 55762.5 ;
      RECT  9695.0 56737.5 9765.0 56602.5 ;
      RECT  9797.5 56295.0 9662.5 56225.0 ;
      RECT  8430.0 56205.0 8500.0 56340.0 ;
      RECT  8570.0 56477.5 8640.0 56612.5 ;
      RECT  9567.5 56440.0 9432.5 56510.0 ;
      RECT  9505.0 57505.0 9575.0 57575.0 ;
      RECT  9695.0 57505.0 9765.0 57575.0 ;
      RECT  9505.0 57540.0 9575.0 57902.5 ;
      RECT  9540.0 57505.0 9730.0 57575.0 ;
      RECT  9695.0 57197.5 9765.0 57540.0 ;
      RECT  9505.0 57902.5 9575.0 58037.5 ;
      RECT  9695.0 57062.5 9765.0 57197.5 ;
      RECT  9797.5 57505.0 9662.5 57575.0 ;
      RECT  8430.0 57460.0 8500.0 57595.0 ;
      RECT  8570.0 57187.5 8640.0 57322.5 ;
      RECT  9567.5 57290.0 9432.5 57360.0 ;
      RECT  9505.0 58985.0 9575.0 58915.0 ;
      RECT  9695.0 58985.0 9765.0 58915.0 ;
      RECT  9505.0 58950.0 9575.0 58587.5 ;
      RECT  9540.0 58985.0 9730.0 58915.0 ;
      RECT  9695.0 59292.5 9765.0 58950.0 ;
      RECT  9505.0 58587.5 9575.0 58452.5 ;
      RECT  9695.0 59427.5 9765.0 59292.5 ;
      RECT  9797.5 58985.0 9662.5 58915.0 ;
      RECT  8430.0 58895.0 8500.0 59030.0 ;
      RECT  8570.0 59167.5 8640.0 59302.5 ;
      RECT  9567.5 59130.0 9432.5 59200.0 ;
      RECT  9505.0 60195.0 9575.0 60265.0 ;
      RECT  9695.0 60195.0 9765.0 60265.0 ;
      RECT  9505.0 60230.0 9575.0 60592.5 ;
      RECT  9540.0 60195.0 9730.0 60265.0 ;
      RECT  9695.0 59887.5 9765.0 60230.0 ;
      RECT  9505.0 60592.5 9575.0 60727.5 ;
      RECT  9695.0 59752.5 9765.0 59887.5 ;
      RECT  9797.5 60195.0 9662.5 60265.0 ;
      RECT  8430.0 60150.0 8500.0 60285.0 ;
      RECT  8570.0 59877.5 8640.0 60012.5 ;
      RECT  9567.5 59980.0 9432.5 60050.0 ;
      RECT  9505.0 61675.0 9575.0 61605.0 ;
      RECT  9695.0 61675.0 9765.0 61605.0 ;
      RECT  9505.0 61640.0 9575.0 61277.5 ;
      RECT  9540.0 61675.0 9730.0 61605.0 ;
      RECT  9695.0 61982.5 9765.0 61640.0 ;
      RECT  9505.0 61277.5 9575.0 61142.5 ;
      RECT  9695.0 62117.5 9765.0 61982.5 ;
      RECT  9797.5 61675.0 9662.5 61605.0 ;
      RECT  8430.0 61585.0 8500.0 61720.0 ;
      RECT  8570.0 61857.5 8640.0 61992.5 ;
      RECT  9567.5 61820.0 9432.5 61890.0 ;
      RECT  9505.0 62885.0 9575.0 62955.0 ;
      RECT  9695.0 62885.0 9765.0 62955.0 ;
      RECT  9505.0 62920.0 9575.0 63282.5 ;
      RECT  9540.0 62885.0 9730.0 62955.0 ;
      RECT  9695.0 62577.5 9765.0 62920.0 ;
      RECT  9505.0 63282.5 9575.0 63417.5 ;
      RECT  9695.0 62442.5 9765.0 62577.5 ;
      RECT  9797.5 62885.0 9662.5 62955.0 ;
      RECT  8430.0 62840.0 8500.0 62975.0 ;
      RECT  8570.0 62567.5 8640.0 62702.5 ;
      RECT  9567.5 62670.0 9432.5 62740.0 ;
      RECT  9505.0 64365.0 9575.0 64295.0 ;
      RECT  9695.0 64365.0 9765.0 64295.0 ;
      RECT  9505.0 64330.0 9575.0 63967.5 ;
      RECT  9540.0 64365.0 9730.0 64295.0 ;
      RECT  9695.0 64672.5 9765.0 64330.0 ;
      RECT  9505.0 63967.5 9575.0 63832.5 ;
      RECT  9695.0 64807.5 9765.0 64672.5 ;
      RECT  9797.5 64365.0 9662.5 64295.0 ;
      RECT  8430.0 64275.0 8500.0 64410.0 ;
      RECT  8570.0 64547.5 8640.0 64682.5 ;
      RECT  9567.5 64510.0 9432.5 64580.0 ;
      RECT  9505.0 65575.0 9575.0 65645.0 ;
      RECT  9695.0 65575.0 9765.0 65645.0 ;
      RECT  9505.0 65610.0 9575.0 65972.5 ;
      RECT  9540.0 65575.0 9730.0 65645.0 ;
      RECT  9695.0 65267.5 9765.0 65610.0 ;
      RECT  9505.0 65972.5 9575.0 66107.5 ;
      RECT  9695.0 65132.5 9765.0 65267.5 ;
      RECT  9797.5 65575.0 9662.5 65645.0 ;
      RECT  8430.0 65530.0 8500.0 65665.0 ;
      RECT  8570.0 65257.5 8640.0 65392.5 ;
      RECT  9567.5 65360.0 9432.5 65430.0 ;
      RECT  9505.0 67055.0 9575.0 66985.0 ;
      RECT  9695.0 67055.0 9765.0 66985.0 ;
      RECT  9505.0 67020.0 9575.0 66657.5 ;
      RECT  9540.0 67055.0 9730.0 66985.0 ;
      RECT  9695.0 67362.5 9765.0 67020.0 ;
      RECT  9505.0 66657.5 9575.0 66522.5 ;
      RECT  9695.0 67497.5 9765.0 67362.5 ;
      RECT  9797.5 67055.0 9662.5 66985.0 ;
      RECT  8430.0 66965.0 8500.0 67100.0 ;
      RECT  8570.0 67237.5 8640.0 67372.5 ;
      RECT  9567.5 67200.0 9432.5 67270.0 ;
      RECT  9505.0 68265.0 9575.0 68335.0 ;
      RECT  9695.0 68265.0 9765.0 68335.0 ;
      RECT  9505.0 68300.0 9575.0 68662.5 ;
      RECT  9540.0 68265.0 9730.0 68335.0 ;
      RECT  9695.0 67957.5 9765.0 68300.0 ;
      RECT  9505.0 68662.5 9575.0 68797.5 ;
      RECT  9695.0 67822.5 9765.0 67957.5 ;
      RECT  9797.5 68265.0 9662.5 68335.0 ;
      RECT  8430.0 68220.0 8500.0 68355.0 ;
      RECT  8570.0 67947.5 8640.0 68082.5 ;
      RECT  9567.5 68050.0 9432.5 68120.0 ;
      RECT  9505.0 69745.0 9575.0 69675.0 ;
      RECT  9695.0 69745.0 9765.0 69675.0 ;
      RECT  9505.0 69710.0 9575.0 69347.5 ;
      RECT  9540.0 69745.0 9730.0 69675.0 ;
      RECT  9695.0 70052.5 9765.0 69710.0 ;
      RECT  9505.0 69347.5 9575.0 69212.5 ;
      RECT  9695.0 70187.5 9765.0 70052.5 ;
      RECT  9797.5 69745.0 9662.5 69675.0 ;
      RECT  8430.0 69655.0 8500.0 69790.0 ;
      RECT  8570.0 69927.5 8640.0 70062.5 ;
      RECT  9567.5 69890.0 9432.5 69960.0 ;
      RECT  8430.0 27310.0 8500.0 70350.0 ;
      RECT  4655.0 10760.0 11095.0 10055.0 ;
      RECT  4655.0 9350.0 11095.0 10055.0 ;
      RECT  4655.0 9350.0 11095.0 8645.0 ;
      RECT  4655.0 7940.0 11095.0 8645.0 ;
      RECT  4655.0 7940.0 11095.0 7235.0 ;
      RECT  4655.0 6530.0 11095.0 7235.0 ;
      RECT  4655.0 6530.0 11095.0 5825.0 ;
      RECT  4655.0 10442.5 4800.0 10372.5 ;
      RECT  4655.0 9737.5 4800.0 9667.5 ;
      RECT  4655.0 9032.5 4800.0 8962.5 ;
      RECT  4655.0 8327.5 4800.0 8257.5 ;
      RECT  4655.0 7622.5 4800.0 7552.5 ;
      RECT  4655.0 6917.5 4800.0 6847.5 ;
      RECT  4655.0 6212.5 4800.0 6142.5 ;
      RECT  10825.0 10442.5 11095.0 10372.5 ;
      RECT  10407.5 10597.5 11095.0 10527.5 ;
      RECT  10825.0 9737.5 11095.0 9667.5 ;
      RECT  10407.5 9582.5 11095.0 9512.5 ;
      RECT  10825.0 9032.5 11095.0 8962.5 ;
      RECT  10407.5 9187.5 11095.0 9117.5 ;
      RECT  10825.0 8327.5 11095.0 8257.5 ;
      RECT  10407.5 8172.5 11095.0 8102.5 ;
      RECT  10825.0 7622.5 11095.0 7552.5 ;
      RECT  10407.5 7777.5 11095.0 7707.5 ;
      RECT  10825.0 6917.5 11095.0 6847.5 ;
      RECT  10407.5 6762.5 11095.0 6692.5 ;
      RECT  10825.0 6212.5 11095.0 6142.5 ;
      RECT  10407.5 6367.5 11095.0 6297.5 ;
      RECT  4655.0 10795.0 11095.0 10725.0 ;
      RECT  4655.0 10090.0 11095.0 10020.0 ;
      RECT  4655.0 9385.0 11095.0 9315.0 ;
      RECT  4655.0 8680.0 11095.0 8610.0 ;
      RECT  4655.0 7975.0 11095.0 7905.0 ;
      RECT  4655.0 7270.0 11095.0 7200.0 ;
      RECT  4655.0 6565.0 11095.0 6495.0 ;
      RECT  4655.0 5860.0 11095.0 5790.0 ;
      RECT  16192.5 5815.0 16262.5 5950.0 ;
      RECT  19012.5 5815.0 19082.5 5950.0 ;
      RECT  16402.5 35.0 16472.5 170.0 ;
      RECT  19222.5 35.0 19292.5 170.0 ;
      RECT  13992.5 27345.0 14127.5 27275.0 ;
      RECT  13992.5 30035.0 14127.5 29965.0 ;
      RECT  13992.5 32725.0 14127.5 32655.0 ;
      RECT  13992.5 35415.0 14127.5 35345.0 ;
      RECT  13992.5 38105.0 14127.5 38035.0 ;
      RECT  13992.5 40795.0 14127.5 40725.0 ;
      RECT  13992.5 43485.0 14127.5 43415.0 ;
      RECT  13992.5 46175.0 14127.5 46105.0 ;
      RECT  13992.5 48865.0 14127.5 48795.0 ;
      RECT  13992.5 51555.0 14127.5 51485.0 ;
      RECT  13992.5 54245.0 14127.5 54175.0 ;
      RECT  13992.5 56935.0 14127.5 56865.0 ;
      RECT  13992.5 59625.0 14127.5 59555.0 ;
      RECT  13992.5 62315.0 14127.5 62245.0 ;
      RECT  13992.5 65005.0 14127.5 64935.0 ;
      RECT  13992.5 67695.0 14127.5 67625.0 ;
      RECT  13992.5 70385.0 14127.5 70315.0 ;
      RECT  10720.0 11340.0 10585.0 11410.0 ;
      RECT  12045.0 11340.0 11910.0 11410.0 ;
      RECT  10445.0 12685.0 10310.0 12755.0 ;
      RECT  12250.0 12685.0 12115.0 12755.0 ;
      RECT  11635.0 16720.0 11500.0 16790.0 ;
      RECT  12455.0 16720.0 12320.0 16790.0 ;
      RECT  11360.0 18065.0 11225.0 18135.0 ;
      RECT  12660.0 18065.0 12525.0 18135.0 ;
      RECT  11085.0 19410.0 10950.0 19480.0 ;
      RECT  12865.0 19410.0 12730.0 19480.0 ;
      RECT  11840.0 11135.0 11705.0 11205.0 ;
      RECT  11840.0 11135.0 11705.0 11205.0 ;
      RECT  13925.0 11205.0 14060.0 11135.0 ;
      RECT  11840.0 13825.0 11705.0 13895.0 ;
      RECT  11840.0 13825.0 11705.0 13895.0 ;
      RECT  13925.0 13895.0 14060.0 13825.0 ;
      RECT  11840.0 16515.0 11705.0 16585.0 ;
      RECT  11840.0 16515.0 11705.0 16585.0 ;
      RECT  13925.0 16585.0 14060.0 16515.0 ;
      RECT  11840.0 19205.0 11705.0 19275.0 ;
      RECT  11840.0 19205.0 11705.0 19275.0 ;
      RECT  13925.0 19275.0 14060.0 19205.0 ;
      RECT  11840.0 21895.0 11705.0 21965.0 ;
      RECT  11840.0 21895.0 11705.0 21965.0 ;
      RECT  13925.0 21965.0 14060.0 21895.0 ;
      RECT  11840.0 24585.0 11705.0 24655.0 ;
      RECT  11840.0 24585.0 11705.0 24655.0 ;
      RECT  13925.0 24655.0 14060.0 24585.0 ;
      RECT  13070.0 25305.0 12935.0 25375.0 ;
      RECT  13275.0 25165.0 13140.0 25235.0 ;
      RECT  13480.0 25025.0 13345.0 25095.0 ;
      RECT  13685.0 24885.0 13550.0 24955.0 ;
      RECT  13070.0 627.5 12935.0 697.5 ;
      RECT  13275.0 2062.5 13140.0 2132.5 ;
      RECT  13480.0 3317.5 13345.0 3387.5 ;
      RECT  13685.0 4752.5 13550.0 4822.5 ;
      RECT  13992.5 70.0 14127.5 2.49800180541e-13 ;
      RECT  13992.5 2760.0 14127.5 2690.0 ;
      RECT  13992.5 5450.0 14127.5 5380.0 ;
      RECT  11162.5 6847.5 11027.5 6917.5 ;
      RECT  7260.0 5207.5 7330.0 5342.5 ;
      RECT  11162.5 6142.5 11027.5 6212.5 ;
      RECT  7535.0 5207.5 7605.0 5342.5 ;
      RECT  11162.5 10372.5 11027.5 10442.5 ;
      RECT  12045.0 10372.5 11910.0 10442.5 ;
      RECT  11162.5 9667.5 11027.5 9737.5 ;
      RECT  12250.0 9667.5 12115.0 9737.5 ;
      RECT  11162.5 8962.5 11027.5 9032.5 ;
      RECT  12455.0 8962.5 12320.0 9032.5 ;
      RECT  11162.5 8257.5 11027.5 8327.5 ;
      RECT  12660.0 8257.5 12525.0 8327.5 ;
      RECT  11162.5 7552.5 11027.5 7622.5 ;
      RECT  12865.0 7552.5 12730.0 7622.5 ;
      RECT  11230.0 10725.0 11095.0 10795.0 ;
      RECT  14127.5 10725.0 13992.5 10795.0 ;
      RECT  11230.0 10020.0 11095.0 10090.0 ;
      RECT  14127.5 10020.0 13992.5 10090.0 ;
      RECT  11230.0 9315.0 11095.0 9385.0 ;
      RECT  14127.5 9315.0 13992.5 9385.0 ;
      RECT  11230.0 8610.0 11095.0 8680.0 ;
      RECT  14127.5 8610.0 13992.5 8680.0 ;
      RECT  11230.0 7905.0 11095.0 7975.0 ;
      RECT  14127.5 7905.0 13992.5 7975.0 ;
      RECT  11230.0 7200.0 11095.0 7270.0 ;
      RECT  14127.5 7200.0 13992.5 7270.0 ;
      RECT  11230.0 6495.0 11095.0 6565.0 ;
      RECT  14127.5 6495.0 13992.5 6565.0 ;
      RECT  11230.0 5790.0 11095.0 5860.0 ;
      RECT  14127.5 5790.0 13992.5 5860.0 ;
      RECT  15265.0 9167.5 15130.0 9237.5 ;
      RECT  14855.0 6982.5 14720.0 7052.5 ;
      RECT  15060.0 8530.0 14925.0 8600.0 ;
      RECT  15265.0 71325.0 15130.0 71395.0 ;
      RECT  15470.0 15670.0 15335.0 15740.0 ;
      RECT  15675.0 19695.0 15540.0 19765.0 ;
      RECT  14650.0 10930.0 14515.0 11000.0 ;
      RECT  8532.5 70520.0 8397.5 70590.0 ;
      RECT  14650.0 70520.0 14515.0 70590.0 ;
      RECT  14342.5 8400.0 14207.5 8470.0 ;
      RECT  14342.5 19825.0 14207.5 19895.0 ;
      RECT  14342.5 9327.5 14207.5 9397.5 ;
      RECT  14342.5 16602.5 14207.5 16672.5 ;
      RECT  16402.5 35.0 16472.5 175.0 ;
      RECT  19222.5 35.0 19292.5 175.0 ;
      RECT  15572.5 35.0 15642.5 72077.5 ;
      RECT  15367.5 35.0 15437.5 72077.5 ;
      RECT  14752.5 35.0 14822.5 72077.5 ;
      RECT  14957.5 35.0 15027.5 72077.5 ;
      RECT  15162.5 35.0 15232.5 72077.5 ;
      RECT  14547.5 35.0 14617.5 72077.5 ;
      RECT  13992.5 35.0 14342.5 72077.5 ;
      RECT  4035.0 34710.0 8.881784197e-13 34780.0 ;
      RECT  4035.0 34915.0 8.881784197e-13 34985.0 ;
      RECT  4035.0 35120.0 8.881784197e-13 35190.0 ;
      RECT  4035.0 35530.0 8.881784197e-13 35600.0 ;
      RECT  3422.5 30220.0 2690.0 30290.0 ;
      RECT  2520.0 27687.5 2450.0 34335.0 ;
      RECT  4035.0 34505.0 3830.0 34575.0 ;
      RECT  2895.0 35325.0 2690.0 35395.0 ;
      RECT  1550.0 34505.0 1345.0 34575.0 ;
      RECT  205.0 35325.0 8.881784197e-13 35395.0 ;
      RECT  165.0 27450.0 870.0 33890.0 ;
      RECT  1575.0 27450.0 870.0 33890.0 ;
      RECT  1575.0 27450.0 2280.0 33890.0 ;
      RECT  482.5 27450.0 552.5 27595.0 ;
      RECT  1187.5 27450.0 1257.5 27595.0 ;
      RECT  1892.5 27450.0 1962.5 27595.0 ;
      RECT  482.5 33620.0 552.5 33890.0 ;
      RECT  327.5 33202.5 397.5 33890.0 ;
      RECT  1187.5 33620.0 1257.5 33890.0 ;
      RECT  1342.5 33202.5 1412.5 33890.0 ;
      RECT  1892.5 33620.0 1962.5 33890.0 ;
      RECT  1737.5 33202.5 1807.5 33890.0 ;
      RECT  130.0 27450.0 200.0 33890.0 ;
      RECT  835.0 27450.0 905.0 33890.0 ;
      RECT  1540.0 27450.0 1610.0 33890.0 ;
      RECT  2245.0 27450.0 2315.0 33890.0 ;
      RECT  3737.5 36780.0 3032.5 36850.0 ;
      RECT  3382.5 36400.0 3312.5 36470.0 ;
      RECT  3382.5 36780.0 3312.5 36850.0 ;
      RECT  3347.5 36400.0 3032.5 36470.0 ;
      RECT  3382.5 36435.0 3312.5 36815.0 ;
      RECT  3737.5 36780.0 3347.5 36850.0 ;
      RECT  3032.5 36400.0 2897.5 36470.0 ;
      RECT  3032.5 36780.0 2897.5 36850.0 ;
      RECT  3872.5 36780.0 3737.5 36850.0 ;
      RECT  3415.0 36780.0 3280.0 36850.0 ;
      RECT  1895.0 36590.0 1965.0 36660.0 ;
      RECT  1930.0 36590.0 2280.0 36660.0 ;
      RECT  1895.0 36625.0 1965.0 36695.0 ;
      RECT  1495.0 36590.0 1565.0 36660.0 ;
      RECT  1495.0 36467.5 1565.0 36625.0 ;
      RECT  1530.0 36590.0 1930.0 36660.0 ;
      RECT  2280.0 36590.0 2415.0 36660.0 ;
      RECT  1495.0 36502.5 1565.0 36367.5 ;
      RECT  1895.0 36762.5 1965.0 36627.5 ;
      RECT  1950.0 37545.0 2020.0 37615.0 ;
      RECT  1950.0 37735.0 2020.0 37805.0 ;
      RECT  1985.0 37545.0 2347.5 37615.0 ;
      RECT  1950.0 37580.0 2020.0 37770.0 ;
      RECT  1642.5 37735.0 1985.0 37805.0 ;
      RECT  2347.5 37545.0 2482.5 37615.0 ;
      RECT  1507.5 37735.0 1642.5 37805.0 ;
      RECT  1950.0 37837.5 2020.0 37702.5 ;
      RECT  1047.5 37340.0 342.5 37410.0 ;
      RECT  692.5 36960.0 622.5 37030.0 ;
      RECT  692.5 37340.0 622.5 37410.0 ;
      RECT  657.5 36960.0 342.5 37030.0 ;
      RECT  692.5 36995.0 622.5 37375.0 ;
      RECT  1047.5 37340.0 657.5 37410.0 ;
      RECT  342.5 36960.0 207.5 37030.0 ;
      RECT  342.5 37340.0 207.5 37410.0 ;
      RECT  1182.5 37340.0 1047.5 37410.0 ;
      RECT  725.0 37340.0 590.0 37410.0 ;
      RECT  397.5 33957.5 327.5 33822.5 ;
      RECT  397.5 35632.5 327.5 35497.5 ;
      RECT  552.5 33957.5 482.5 33822.5 ;
      RECT  552.5 34812.5 482.5 34677.5 ;
      RECT  1412.5 33957.5 1342.5 33822.5 ;
      RECT  1412.5 35017.5 1342.5 34882.5 ;
      RECT  1807.5 33957.5 1737.5 33822.5 ;
      RECT  1807.5 35222.5 1737.5 35087.5 ;
      RECT  200.0 33957.5 130.0 33822.5 ;
      RECT  200.0 34607.5 130.0 34472.5 ;
      RECT  905.0 33957.5 835.0 33822.5 ;
      RECT  905.0 34607.5 835.0 34472.5 ;
      RECT  1610.0 33957.5 1540.0 33822.5 ;
      RECT  1610.0 34607.5 1540.0 34472.5 ;
      RECT  2315.0 33957.5 2245.0 33822.5 ;
      RECT  2315.0 34607.5 2245.0 34472.5 ;
      RECT  1380.0 40115.0 1310.0 47865.0 ;
      RECT  970.0 40115.0 900.0 47555.0 ;
      RECT  265.0 40115.0 195.0 47555.0 ;
      RECT  1207.5 40282.5 1137.5 40880.0 ;
      RECT  785.0 40282.5 715.0 40562.5 ;
      RECT  3372.5 42677.5 3442.5 43072.5 ;
      RECT  3372.5 43072.5 3442.5 43632.5 ;
      RECT  3372.5 43632.5 3442.5 44192.5 ;
      RECT  3372.5 44192.5 3442.5 44752.5 ;
      RECT  3372.5 44917.5 3442.5 45312.5 ;
      RECT  3372.5 45312.5 3442.5 45872.5 ;
      RECT  3372.5 45872.5 3442.5 46432.5 ;
      RECT  3372.5 46432.5 3442.5 46992.5 ;
      RECT  3372.5 47157.5 3442.5 47552.5 ;
      RECT  3372.5 47552.5 3442.5 48112.5 ;
      RECT  3372.5 48112.5 3442.5 48672.5 ;
      RECT  3372.5 48672.5 3442.5 49232.5 ;
      RECT  3372.5 49397.5 3442.5 49792.5 ;
      RECT  3372.5 49792.5 3442.5 50352.5 ;
      RECT  3372.5 50352.5 3442.5 50912.5 ;
      RECT  3372.5 50912.5 3442.5 51472.5 ;
      RECT  2655.0 51602.5 2725.0 51672.5 ;
      RECT  2655.0 51122.5 2725.0 51192.5 ;
      RECT  2690.0 51602.5 3407.5 51672.5 ;
      RECT  2655.0 51157.5 2725.0 51637.5 ;
      RECT  1972.5 51122.5 2690.0 51192.5 ;
      RECT  1937.5 50597.5 2007.5 51157.5 ;
      RECT  1937.5 50037.5 2007.5 50597.5 ;
      RECT  1937.5 49477.5 2007.5 50037.5 ;
      RECT  1937.5 48917.5 2007.5 49312.5 ;
      RECT  1937.5 48357.5 2007.5 48917.5 ;
      RECT  1937.5 47797.5 2007.5 48357.5 ;
      RECT  1937.5 47237.5 2007.5 47797.5 ;
      RECT  1937.5 46677.5 2007.5 47072.5 ;
      RECT  1937.5 46117.5 2007.5 46677.5 ;
      RECT  1937.5 45557.5 2007.5 46117.5 ;
      RECT  1937.5 44997.5 2007.5 45557.5 ;
      RECT  1937.5 44437.5 2007.5 44832.5 ;
      RECT  1937.5 43877.5 2007.5 44437.5 ;
      RECT  1937.5 43317.5 2007.5 43877.5 ;
      RECT  1937.5 42757.5 2007.5 43317.5 ;
      RECT  3340.0 43037.5 3475.0 43107.5 ;
      RECT  3340.0 43597.5 3475.0 43667.5 ;
      RECT  3340.0 44157.5 3475.0 44227.5 ;
      RECT  3340.0 44717.5 3475.0 44787.5 ;
      RECT  3340.0 45277.5 3475.0 45347.5 ;
      RECT  3340.0 45837.5 3475.0 45907.5 ;
      RECT  3340.0 46397.5 3475.0 46467.5 ;
      RECT  3340.0 46957.5 3475.0 47027.5 ;
      RECT  3340.0 47517.5 3475.0 47587.5 ;
      RECT  3340.0 48077.5 3475.0 48147.5 ;
      RECT  3340.0 48637.5 3475.0 48707.5 ;
      RECT  3340.0 49197.5 3475.0 49267.5 ;
      RECT  3340.0 49757.5 3475.0 49827.5 ;
      RECT  3340.0 50317.5 3475.0 50387.5 ;
      RECT  3340.0 50877.5 3475.0 50947.5 ;
      RECT  3340.0 51437.5 3475.0 51507.5 ;
      RECT  1905.0 51122.5 2040.0 51192.5 ;
      RECT  1905.0 50562.5 2040.0 50632.5 ;
      RECT  1905.0 50002.5 2040.0 50072.5 ;
      RECT  1905.0 49442.5 2040.0 49512.5 ;
      RECT  1905.0 48882.5 2040.0 48952.5 ;
      RECT  1905.0 48322.5 2040.0 48392.5 ;
      RECT  1905.0 47762.5 2040.0 47832.5 ;
      RECT  1905.0 47202.5 2040.0 47272.5 ;
      RECT  1905.0 46642.5 2040.0 46712.5 ;
      RECT  1905.0 46082.5 2040.0 46152.5 ;
      RECT  1905.0 45522.5 2040.0 45592.5 ;
      RECT  1905.0 44962.5 2040.0 45032.5 ;
      RECT  1905.0 44402.5 2040.0 44472.5 ;
      RECT  1905.0 43842.5 2040.0 43912.5 ;
      RECT  1905.0 43282.5 2040.0 43352.5 ;
      RECT  1905.0 42722.5 2040.0 42792.5 ;
      RECT  3340.0 42642.5 3475.0 42712.5 ;
      RECT  3340.0 44882.5 3475.0 44952.5 ;
      RECT  3340.0 47122.5 3475.0 47192.5 ;
      RECT  3340.0 49362.5 3475.0 49432.5 ;
      RECT  3340.0 51602.5 3475.0 51672.5 ;
      RECT  1905.0 49277.5 2040.0 49347.5 ;
      RECT  1905.0 47037.5 2040.0 47107.5 ;
      RECT  1905.0 44797.5 2040.0 44867.5 ;
      RECT  935.0 42020.0 225.0 40675.0 ;
      RECT  935.0 42020.0 230.0 43365.0 ;
      RECT  935.0 44710.0 230.0 43365.0 ;
      RECT  935.0 44710.0 230.0 46055.0 ;
      RECT  935.0 47400.0 230.0 46055.0 ;
      RECT  785.0 41920.0 715.0 47555.0 ;
      RECT  450.0 41920.0 380.0 47555.0 ;
      RECT  970.0 41920.0 900.0 47555.0 ;
      RECT  265.0 41920.0 195.0 47555.0 ;
      RECT  1347.5 42092.5 1277.5 42227.5 ;
      RECT  1347.5 44502.5 1277.5 44637.5 ;
      RECT  1347.5 44782.5 1277.5 44917.5 ;
      RECT  1347.5 47192.5 1277.5 47327.5 ;
      RECT  1345.0 42355.0 1275.0 42490.0 ;
      RECT  1380.0 39980.0 1310.0 40115.0 ;
      RECT  867.5 40080.0 1002.5 40150.0 ;
      RECT  162.5 40080.0 297.5 40150.0 ;
      RECT  1105.0 40845.0 1240.0 40915.0 ;
      RECT  1105.0 40247.5 1240.0 40317.5 ;
      RECT  682.5 40247.5 817.5 40317.5 ;
      RECT  3457.5 34402.5 3387.5 34267.5 ;
      RECT  3457.5 30322.5 3387.5 30187.5 ;
      RECT  2725.0 30322.5 2655.0 30187.5 ;
      RECT  2725.0 35837.5 2655.0 35702.5 ;
      RECT  2520.0 27755.0 2450.0 27620.0 ;
      RECT  1965.0 34402.5 1895.0 34267.5 ;
      RECT  1750.0 34812.5 1680.0 34677.5 ;
      RECT  2020.0 37350.0 1950.0 37215.0 ;
      RECT  2020.0 37350.0 1950.0 37215.0 ;
      RECT  2020.0 35837.5 1950.0 35702.5 ;
      RECT  1805.0 37607.5 1735.0 37472.5 ;
      RECT  1805.0 37607.5 1735.0 37472.5 ;
      RECT  1805.0 35632.5 1735.0 35497.5 ;
      RECT  3382.5 35837.5 3312.5 35702.5 ;
      RECT  3522.5 35632.5 3452.5 35497.5 ;
      RECT  3662.5 35017.5 3592.5 34882.5 ;
      RECT  692.5 35837.5 622.5 35702.5 ;
      RECT  832.5 35017.5 762.5 34882.5 ;
      RECT  972.5 35222.5 902.5 35087.5 ;
      RECT  1997.5 37030.0 1862.5 37100.0 ;
      RECT  2052.5 38175.0 1917.5 38245.0 ;
      RECT  785.0 39360.0 650.0 39430.0 ;
      RECT  2040.0 38400.0 1905.0 38470.0 ;
      RECT  4070.0 34607.5 4000.0 34472.5 ;
      RECT  2725.0 35427.5 2655.0 35292.5 ;
      RECT  1380.0 34607.5 1310.0 34472.5 ;
      RECT  35.0 35427.5 -35.0 35292.5 ;
      RECT  4035.0 38400.0 1972.5 38470.0 ;
      RECT  4035.0 39360.0 717.5 39430.0 ;
      RECT  4035.0 37030.0 1930.0 37100.0 ;
      RECT  4035.0 38175.0 1985.0 38245.0 ;
      RECT  4035.0 35735.0 8.881784197e-13 35805.0 ;
      RECT  4035.0 34300.0 0.0 34370.0 ;
      RECT  4035.0 35325.0 8.881784197e-13 35395.0 ;
      RECT  4035.0 34505.0 0.0 34575.0 ;
      RECT  15675.0 38400.0 15540.0 38470.0 ;
      RECT  4035.0 38400.0 3900.0 38470.0 ;
      RECT  15470.0 39360.0 15335.0 39430.0 ;
      RECT  4035.0 39360.0 3900.0 39430.0 ;
      RECT  15060.0 37030.0 14925.0 37100.0 ;
      RECT  4035.0 37030.0 3900.0 37100.0 ;
      RECT  14855.0 38175.0 14720.0 38245.0 ;
      RECT  4035.0 38175.0 3900.0 38245.0 ;
      RECT  15265.0 35735.0 15130.0 35805.0 ;
      RECT  4035.0 35735.0 3900.0 35805.0 ;
      RECT  14650.0 34300.0 14515.0 34370.0 ;
      RECT  4035.0 34300.0 3900.0 34370.0 ;
      RECT  4417.5 35325.0 4282.5 35395.0 ;
      RECT  14235.0 34505.0 14100.0 34575.0 ;
      RECT  4035.0 34505.0 3900.0 34575.0 ;
   LAYER  metal3 ;
      RECT  4035.0 38400.0 15607.5 38470.0 ;
      RECT  4035.0 39360.0 15402.5 39430.0 ;
      RECT  4035.0 37030.0 14992.5 37100.0 ;
      RECT  4035.0 38175.0 14787.5 38245.0 ;
      RECT  4035.0 35735.0 15197.5 35805.0 ;
      RECT  4035.0 34300.0 14582.5 34370.0 ;
      RECT  4035.0 34505.0 14167.5 34575.0 ;
      RECT  16192.5 24360.0 16262.5 24430.0 ;
      RECT  16192.5 5850.0 16262.5 24395.0 ;
      RECT  16227.5 24360.0 16397.5 24430.0 ;
      RECT  19012.5 24360.0 19082.5 24430.0 ;
      RECT  19012.5 5850.0 19082.5 24395.0 ;
      RECT  19047.5 24360.0 19217.5 24430.0 ;
      RECT  16402.5 35.0 16472.5 8965.0 ;
      RECT  19222.5 35.0 19292.5 8965.0 ;
      RECT  11772.5 11135.0 13992.5 11205.0 ;
      RECT  11772.5 13825.0 13992.5 13895.0 ;
      RECT  11772.5 16515.0 13992.5 16585.0 ;
      RECT  11772.5 19205.0 13992.5 19275.0 ;
      RECT  11772.5 21895.0 13992.5 21965.0 ;
      RECT  11772.5 24585.0 13992.5 24655.0 ;
      RECT  7260.0 6847.5 7330.0 6917.5 ;
      RECT  7295.0 6847.5 11095.0 6917.5 ;
      RECT  7260.0 5275.0 7330.0 6882.5 ;
      RECT  7535.0 6142.5 7605.0 6212.5 ;
      RECT  7570.0 6142.5 11095.0 6212.5 ;
      RECT  7535.0 5275.0 7605.0 6177.5 ;
      RECT  16397.5 24325.0 16467.5 24465.0 ;
      RECT  19217.5 24325.0 19287.5 24465.0 ;
      RECT  16402.5 8965.0 16472.5 9105.0 ;
      RECT  19222.5 8965.0 19292.5 9105.0 ;
      RECT  4655.0 10442.5 4795.0 10372.5 ;
      RECT  4655.0 9737.5 4795.0 9667.5 ;
      RECT  4655.0 9032.5 4795.0 8962.5 ;
      RECT  4655.0 8327.5 4795.0 8257.5 ;
      RECT  4655.0 7622.5 4795.0 7552.5 ;
      RECT  4655.0 6917.5 4795.0 6847.5 ;
      RECT  4655.0 6212.5 4795.0 6142.5 ;
      RECT  16192.5 5815.0 16262.5 5950.0 ;
      RECT  19012.5 5815.0 19082.5 5950.0 ;
      RECT  16402.5 35.0 16472.5 170.0 ;
      RECT  19222.5 35.0 19292.5 170.0 ;
      RECT  11840.0 11135.0 11705.0 11205.0 ;
      RECT  13925.0 11205.0 14060.0 11135.0 ;
      RECT  11840.0 13825.0 11705.0 13895.0 ;
      RECT  13925.0 13895.0 14060.0 13825.0 ;
      RECT  11840.0 16515.0 11705.0 16585.0 ;
      RECT  13925.0 16585.0 14060.0 16515.0 ;
      RECT  11840.0 19205.0 11705.0 19275.0 ;
      RECT  13925.0 19275.0 14060.0 19205.0 ;
      RECT  11840.0 21895.0 11705.0 21965.0 ;
      RECT  13925.0 21965.0 14060.0 21895.0 ;
      RECT  11840.0 24585.0 11705.0 24655.0 ;
      RECT  13925.0 24655.0 14060.0 24585.0 ;
      RECT  11162.5 6847.5 11027.5 6917.5 ;
      RECT  7260.0 5207.5 7330.0 5342.5 ;
      RECT  11162.5 6142.5 11027.5 6212.5 ;
      RECT  7535.0 5207.5 7605.0 5342.5 ;
      RECT  4175.0 10372.5 4655.0 10442.5 ;
      RECT  4175.0 9667.5 4655.0 9737.5 ;
      RECT  4175.0 8962.5 4655.0 9032.5 ;
      RECT  4175.0 8257.5 4655.0 8327.5 ;
      RECT  4175.0 7552.5 4655.0 7622.5 ;
      RECT  4175.0 6847.5 4655.0 6917.5 ;
      RECT  4175.0 6142.5 4655.0 6212.5 ;
      RECT  397.5 33890.0 327.5 35565.0 ;
      RECT  552.5 33890.0 482.5 34745.0 ;
      RECT  1412.5 33890.0 1342.5 34950.0 ;
      RECT  1807.5 33890.0 1737.5 35155.0 ;
      RECT  200.0 33890.0 130.0 34540.0 ;
      RECT  905.0 33890.0 835.0 34540.0 ;
      RECT  1610.0 33890.0 1540.0 34540.0 ;
      RECT  2315.0 33890.0 2245.0 34540.0 ;
      RECT  2725.0 30255.0 2655.0 35770.0 ;
      RECT  2020.0 35770.0 1950.0 37282.5 ;
      RECT  1805.0 35565.0 1735.0 37540.0 ;
      RECT  482.5 27450.0 552.5 27590.0 ;
      RECT  1187.5 27450.0 1257.5 27590.0 ;
      RECT  1892.5 27450.0 1962.5 27590.0 ;
      RECT  397.5 33957.5 327.5 33822.5 ;
      RECT  397.5 35632.5 327.5 35497.5 ;
      RECT  552.5 33957.5 482.5 33822.5 ;
      RECT  552.5 34812.5 482.5 34677.5 ;
      RECT  1412.5 33957.5 1342.5 33822.5 ;
      RECT  1412.5 35017.5 1342.5 34882.5 ;
      RECT  1807.5 33957.5 1737.5 33822.5 ;
      RECT  1807.5 35222.5 1737.5 35087.5 ;
      RECT  200.0 33957.5 130.0 33822.5 ;
      RECT  200.0 34607.5 130.0 34472.5 ;
      RECT  905.0 33957.5 835.0 33822.5 ;
      RECT  905.0 34607.5 835.0 34472.5 ;
      RECT  1610.0 33957.5 1540.0 33822.5 ;
      RECT  1610.0 34607.5 1540.0 34472.5 ;
      RECT  2315.0 33957.5 2245.0 33822.5 ;
      RECT  2315.0 34607.5 2245.0 34472.5 ;
      RECT  2725.0 30322.5 2655.0 30187.5 ;
      RECT  2725.0 35837.5 2655.0 35702.5 ;
      RECT  2020.0 37350.0 1950.0 37215.0 ;
      RECT  2020.0 35837.5 1950.0 35702.5 ;
      RECT  1805.0 37607.5 1735.0 37472.5 ;
      RECT  1805.0 35632.5 1735.0 35497.5 ;
      RECT  1257.5 27450.0 1187.5 27590.0 ;
      RECT  1962.5 27450.0 1892.5 27590.0 ;
      RECT  552.5 27450.0 482.5 27590.0 ;
      RECT  15675.0 38400.0 15540.0 38470.0 ;
      RECT  4035.0 38400.0 3900.0 38470.0 ;
      RECT  15470.0 39360.0 15335.0 39430.0 ;
      RECT  4035.0 39360.0 3900.0 39430.0 ;
      RECT  15060.0 37030.0 14925.0 37100.0 ;
      RECT  4035.0 37030.0 3900.0 37100.0 ;
      RECT  14855.0 38175.0 14720.0 38245.0 ;
      RECT  4035.0 38175.0 3900.0 38245.0 ;
      RECT  15265.0 35735.0 15130.0 35805.0 ;
      RECT  4035.0 35735.0 3900.0 35805.0 ;
      RECT  14650.0 34300.0 14515.0 34370.0 ;
      RECT  4035.0 34300.0 3900.0 34370.0 ;
      RECT  14235.0 34505.0 14100.0 34575.0 ;
      RECT  4035.0 34505.0 3900.0 34575.0 ;
   END
   END    sram_2_16_1_freepdk45
END    LIBRARY
