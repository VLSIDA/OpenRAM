magic
tech sky130A
magscale 1 2
timestamp 1595931502
<< checkpaint >>
rect -1296 -1309 3136 11397
<< metal1 >>
rect 624 10054 688 10106
rect 1360 10054 1424 10106
rect 49 9456 113 9508
rect 164 9456 228 9508
rect 417 9456 481 9508
rect 785 9456 849 9508
rect 1153 9456 1217 9508
rect 1521 9456 1585 9508
rect 624 8934 688 8986
rect 1360 8934 1424 8986
rect 49 8412 113 8464
rect 164 8412 228 8464
rect 417 8412 481 8464
rect 785 8412 849 8464
rect 1153 8412 1217 8464
rect 1521 8412 1585 8464
rect 624 7814 688 7866
rect 1360 7814 1424 7866
rect 49 7216 113 7268
rect 164 7216 228 7268
rect 417 7216 481 7268
rect 785 7216 849 7268
rect 1153 7216 1217 7268
rect 1521 7216 1585 7268
rect 624 6694 688 6746
rect 1360 6694 1424 6746
rect 49 6172 113 6224
rect 164 6172 228 6224
rect 417 6172 481 6224
rect 785 6172 849 6224
rect 1153 6172 1217 6224
rect 1521 6172 1585 6224
rect 624 5574 688 5626
rect 1360 5574 1424 5626
rect 49 4976 113 5028
rect 164 4976 228 5028
rect 417 4976 481 5028
rect 785 4976 849 5028
rect 1153 4976 1217 5028
rect 1521 4976 1585 5028
rect 624 4454 688 4506
rect 1360 4454 1424 4506
rect 49 3932 113 3984
rect 164 3932 228 3984
rect 417 3932 481 3984
rect 785 3932 849 3984
rect 1153 3932 1217 3984
rect 1521 3932 1585 3984
rect 624 3334 688 3386
rect 1360 3334 1424 3386
rect 49 2736 113 2788
rect 164 2736 228 2788
rect 417 2736 481 2788
rect 785 2736 849 2788
rect 1153 2736 1217 2788
rect 1521 2736 1585 2788
rect 624 2214 688 2266
rect 1360 2214 1424 2266
rect 49 1692 113 1744
rect 164 1692 228 1744
rect 417 1692 481 1744
rect 785 1692 849 1744
rect 1153 1692 1217 1744
rect 1521 1692 1585 1744
rect 624 1094 688 1146
rect 1360 1094 1424 1146
rect 49 496 113 548
rect 164 496 228 548
rect 417 496 481 548
rect 785 496 849 548
rect 1153 496 1217 548
rect 1521 496 1585 548
rect 624 -26 688 26
rect 1360 -26 1424 26
<< metal2 >>
rect 628 10056 684 10104
rect 1364 10056 1420 10104
rect 67 8974 95 9482
rect 168 9458 224 9506
rect 421 9458 477 9506
rect 789 9458 845 9506
rect 1157 9458 1213 9506
rect 1525 9496 1581 9506
rect 1525 9468 1651 9496
rect 1525 9458 1581 9468
rect 67 8946 210 8974
rect 182 8462 210 8946
rect 628 8936 684 8984
rect 1364 8936 1420 8984
rect 67 7854 95 8438
rect 168 8414 224 8462
rect 421 8414 477 8462
rect 789 8414 845 8462
rect 1157 8414 1213 8462
rect 1525 8414 1581 8462
rect 67 7826 210 7854
rect 182 7266 210 7826
rect 628 7816 684 7864
rect 1364 7816 1420 7864
rect 67 6734 95 7242
rect 168 7218 224 7266
rect 421 7218 477 7266
rect 789 7218 845 7266
rect 1157 7218 1213 7266
rect 1525 7218 1581 7266
rect 67 6706 210 6734
rect 182 6222 210 6706
rect 628 6696 684 6744
rect 1364 6696 1420 6744
rect 67 5614 95 6198
rect 168 6174 224 6222
rect 421 6174 477 6222
rect 789 6174 845 6222
rect 1157 6174 1213 6222
rect 1525 6174 1581 6222
rect 67 5586 210 5614
rect 182 5026 210 5586
rect 628 5576 684 5624
rect 1364 5576 1420 5624
rect 67 4494 95 5002
rect 168 4978 224 5026
rect 421 4978 477 5026
rect 789 4978 845 5026
rect 1157 4978 1213 5026
rect 1525 4978 1581 5026
rect 67 4466 210 4494
rect 182 3982 210 4466
rect 628 4456 684 4504
rect 1364 4456 1420 4504
rect 67 3374 95 3958
rect 168 3934 224 3982
rect 421 3934 477 3982
rect 789 3934 845 3982
rect 1157 3934 1213 3982
rect 1525 3934 1581 3982
rect 67 3346 210 3374
rect 182 2786 210 3346
rect 628 3336 684 3384
rect 1364 3336 1420 3384
rect 67 2254 95 2762
rect 168 2738 224 2786
rect 421 2738 477 2786
rect 789 2738 845 2786
rect 1157 2738 1213 2786
rect 1525 2738 1581 2786
rect 67 2226 210 2254
rect 182 1742 210 2226
rect 628 2216 684 2264
rect 1364 2216 1420 2264
rect 67 1134 95 1718
rect 168 1694 224 1742
rect 421 1694 477 1742
rect 789 1694 845 1742
rect 1157 1694 1213 1742
rect 1525 1694 1581 1742
rect 67 1106 210 1134
rect 182 546 210 1106
rect 628 1096 684 1144
rect 1364 1096 1420 1144
rect 64 0 92 522
rect 168 498 224 546
rect 421 498 477 546
rect 789 498 845 546
rect 1157 498 1213 546
rect 1525 498 1581 546
rect 628 -24 684 24
rect 1364 -24 1420 24
rect 1623 0 1651 9468
<< metal3 >>
rect 607 10031 705 10129
rect 1343 10031 1441 10129
rect 196 9452 1553 9512
rect 607 8911 705 9009
rect 1343 8911 1441 9009
rect 196 8408 1553 8468
rect 607 7791 705 7889
rect 1343 7791 1441 7889
rect 196 7212 1553 7272
rect 607 6671 705 6769
rect 1343 6671 1441 6769
rect 196 6168 1553 6228
rect 607 5551 705 5649
rect 1343 5551 1441 5649
rect 196 4972 1553 5032
rect 607 4431 705 4529
rect 1343 4431 1441 4529
rect 196 3928 1553 3988
rect 607 3311 705 3409
rect 1343 3311 1441 3409
rect 196 2732 1553 2792
rect 607 2191 705 2289
rect 1343 2191 1441 2289
rect 196 1688 1553 1748
rect 607 1071 705 1169
rect 1343 1071 1441 1169
rect 196 492 1553 552
rect 607 -49 705 49
rect 1343 -49 1441 49
use contact_9  contact_9_80
timestamp 1595931502
transform 1 0 416 0 1 485
box 0 0 66 74
use contact_9  contact_9_79
timestamp 1595931502
transform 1 0 784 0 1 485
box 0 0 66 74
use contact_9  contact_9_78
timestamp 1595931502
transform 1 0 1152 0 1 485
box 0 0 66 74
use contact_9  contact_9_77
timestamp 1595931502
transform 1 0 1520 0 1 485
box 0 0 66 74
use contact_9  contact_9_76
timestamp 1595931502
transform 1 0 163 0 1 485
box 0 0 66 74
use contact_9  contact_9_75
timestamp 1595931502
transform 1 0 416 0 1 1681
box 0 0 66 74
use contact_9  contact_9_74
timestamp 1595931502
transform 1 0 784 0 1 1681
box 0 0 66 74
use contact_9  contact_9_73
timestamp 1595931502
transform 1 0 1152 0 1 1681
box 0 0 66 74
use contact_9  contact_9_72
timestamp 1595931502
transform 1 0 1520 0 1 1681
box 0 0 66 74
use contact_9  contact_9_71
timestamp 1595931502
transform 1 0 163 0 1 1681
box 0 0 66 74
use contact_9  contact_9_70
timestamp 1595931502
transform 1 0 416 0 1 2725
box 0 0 66 74
use contact_9  contact_9_69
timestamp 1595931502
transform 1 0 784 0 1 2725
box 0 0 66 74
use contact_9  contact_9_68
timestamp 1595931502
transform 1 0 1152 0 1 2725
box 0 0 66 74
use contact_9  contact_9_67
timestamp 1595931502
transform 1 0 1520 0 1 2725
box 0 0 66 74
use contact_9  contact_9_66
timestamp 1595931502
transform 1 0 163 0 1 2725
box 0 0 66 74
use contact_9  contact_9_65
timestamp 1595931502
transform 1 0 416 0 1 3921
box 0 0 66 74
use contact_9  contact_9_64
timestamp 1595931502
transform 1 0 784 0 1 3921
box 0 0 66 74
use contact_9  contact_9_63
timestamp 1595931502
transform 1 0 1152 0 1 3921
box 0 0 66 74
use contact_9  contact_9_62
timestamp 1595931502
transform 1 0 1520 0 1 3921
box 0 0 66 74
use contact_9  contact_9_61
timestamp 1595931502
transform 1 0 163 0 1 3921
box 0 0 66 74
use contact_9  contact_9_60
timestamp 1595931502
transform 1 0 416 0 1 4965
box 0 0 66 74
use contact_9  contact_9_59
timestamp 1595931502
transform 1 0 784 0 1 4965
box 0 0 66 74
use contact_9  contact_9_58
timestamp 1595931502
transform 1 0 1152 0 1 4965
box 0 0 66 74
use contact_9  contact_9_57
timestamp 1595931502
transform 1 0 1520 0 1 4965
box 0 0 66 74
use contact_9  contact_9_56
timestamp 1595931502
transform 1 0 163 0 1 4965
box 0 0 66 74
use contact_9  contact_9_55
timestamp 1595931502
transform 1 0 416 0 1 6161
box 0 0 66 74
use contact_9  contact_9_54
timestamp 1595931502
transform 1 0 784 0 1 6161
box 0 0 66 74
use contact_9  contact_9_53
timestamp 1595931502
transform 1 0 1152 0 1 6161
box 0 0 66 74
use contact_9  contact_9_52
timestamp 1595931502
transform 1 0 1520 0 1 6161
box 0 0 66 74
use contact_9  contact_9_51
timestamp 1595931502
transform 1 0 163 0 1 6161
box 0 0 66 74
use contact_9  contact_9_50
timestamp 1595931502
transform 1 0 416 0 1 7205
box 0 0 66 74
use contact_9  contact_9_49
timestamp 1595931502
transform 1 0 784 0 1 7205
box 0 0 66 74
use contact_9  contact_9_48
timestamp 1595931502
transform 1 0 1152 0 1 7205
box 0 0 66 74
use contact_9  contact_9_47
timestamp 1595931502
transform 1 0 1520 0 1 7205
box 0 0 66 74
use contact_9  contact_9_46
timestamp 1595931502
transform 1 0 163 0 1 7205
box 0 0 66 74
use contact_9  contact_9_45
timestamp 1595931502
transform 1 0 416 0 1 8401
box 0 0 66 74
use contact_9  contact_9_44
timestamp 1595931502
transform 1 0 784 0 1 8401
box 0 0 66 74
use contact_9  contact_9_43
timestamp 1595931502
transform 1 0 1152 0 1 8401
box 0 0 66 74
use contact_9  contact_9_42
timestamp 1595931502
transform 1 0 1520 0 1 8401
box 0 0 66 74
use contact_9  contact_9_41
timestamp 1595931502
transform 1 0 163 0 1 8401
box 0 0 66 74
use contact_9  contact_9_40
timestamp 1595931502
transform 1 0 416 0 1 9445
box 0 0 66 74
use contact_9  contact_9_39
timestamp 1595931502
transform 1 0 784 0 1 9445
box 0 0 66 74
use contact_9  contact_9_38
timestamp 1595931502
transform 1 0 1152 0 1 9445
box 0 0 66 74
use contact_9  contact_9_37
timestamp 1595931502
transform 1 0 1520 0 1 9445
box 0 0 66 74
use contact_9  contact_9_36
timestamp 1595931502
transform 1 0 163 0 1 9445
box 0 0 66 74
use contact_9  contact_9_35
timestamp 1595931502
transform 1 0 623 0 1 1083
box 0 0 66 74
use contact_9  contact_9_34
timestamp 1595931502
transform 1 0 1359 0 1 1083
box 0 0 66 74
use contact_9  contact_9_33
timestamp 1595931502
transform 1 0 623 0 1 -37
box 0 0 66 74
use contact_9  contact_9_32
timestamp 1595931502
transform 1 0 1359 0 1 -37
box 0 0 66 74
use contact_9  contact_9_31
timestamp 1595931502
transform 1 0 623 0 1 1083
box 0 0 66 74
use contact_9  contact_9_30
timestamp 1595931502
transform 1 0 1359 0 1 1083
box 0 0 66 74
use contact_9  contact_9_29
timestamp 1595931502
transform 1 0 623 0 1 2203
box 0 0 66 74
use contact_9  contact_9_28
timestamp 1595931502
transform 1 0 1359 0 1 2203
box 0 0 66 74
use contact_9  contact_9_27
timestamp 1595931502
transform 1 0 623 0 1 3323
box 0 0 66 74
use contact_9  contact_9_26
timestamp 1595931502
transform 1 0 1359 0 1 3323
box 0 0 66 74
use contact_9  contact_9_25
timestamp 1595931502
transform 1 0 623 0 1 2203
box 0 0 66 74
use contact_9  contact_9_24
timestamp 1595931502
transform 1 0 1359 0 1 2203
box 0 0 66 74
use contact_9  contact_9_23
timestamp 1595931502
transform 1 0 623 0 1 3323
box 0 0 66 74
use contact_9  contact_9_22
timestamp 1595931502
transform 1 0 1359 0 1 3323
box 0 0 66 74
use contact_9  contact_9_21
timestamp 1595931502
transform 1 0 623 0 1 4443
box 0 0 66 74
use contact_9  contact_9_20
timestamp 1595931502
transform 1 0 1359 0 1 4443
box 0 0 66 74
use contact_9  contact_9_19
timestamp 1595931502
transform 1 0 623 0 1 5563
box 0 0 66 74
use contact_9  contact_9_18
timestamp 1595931502
transform 1 0 1359 0 1 5563
box 0 0 66 74
use contact_9  contact_9_17
timestamp 1595931502
transform 1 0 623 0 1 4443
box 0 0 66 74
use contact_9  contact_9_16
timestamp 1595931502
transform 1 0 1359 0 1 4443
box 0 0 66 74
use contact_9  contact_9_15
timestamp 1595931502
transform 1 0 623 0 1 5563
box 0 0 66 74
use contact_9  contact_9_14
timestamp 1595931502
transform 1 0 1359 0 1 5563
box 0 0 66 74
use contact_9  contact_9_13
timestamp 1595931502
transform 1 0 623 0 1 6683
box 0 0 66 74
use contact_9  contact_9_12
timestamp 1595931502
transform 1 0 1359 0 1 6683
box 0 0 66 74
use contact_9  contact_9_11
timestamp 1595931502
transform 1 0 623 0 1 7803
box 0 0 66 74
use contact_9  contact_9_10
timestamp 1595931502
transform 1 0 1359 0 1 7803
box 0 0 66 74
use contact_9  contact_9_9
timestamp 1595931502
transform 1 0 623 0 1 6683
box 0 0 66 74
use contact_9  contact_9_8
timestamp 1595931502
transform 1 0 1359 0 1 6683
box 0 0 66 74
use contact_9  contact_9_7
timestamp 1595931502
transform 1 0 623 0 1 7803
box 0 0 66 74
use contact_9  contact_9_6
timestamp 1595931502
transform 1 0 1359 0 1 7803
box 0 0 66 74
use contact_9  contact_9_5
timestamp 1595931502
transform 1 0 623 0 1 8923
box 0 0 66 74
use contact_9  contact_9_4
timestamp 1595931502
transform 1 0 1359 0 1 8923
box 0 0 66 74
use contact_9  contact_9_3
timestamp 1595931502
transform 1 0 623 0 1 10043
box 0 0 66 74
use contact_9  contact_9_2
timestamp 1595931502
transform 1 0 1359 0 1 10043
box 0 0 66 74
use contact_9  contact_9_1
timestamp 1595931502
transform 1 0 623 0 1 8923
box 0 0 66 74
use contact_9  contact_9_0
timestamp 1595931502
transform 1 0 1359 0 1 8923
box 0 0 66 74
use pinv_10  pinv_10_44
timestamp 1595931502
transform 1 0 0 0 1 0
box -36 -17 404 1177
use pinv_10  pinv_10_43
timestamp 1595931502
transform 1 0 368 0 1 0
box -36 -17 404 1177
use pinv_10  pinv_10_42
timestamp 1595931502
transform 1 0 736 0 1 0
box -36 -17 404 1177
use pinv_10  pinv_10_41
timestamp 1595931502
transform 1 0 1104 0 1 0
box -36 -17 404 1177
use pinv_10  pinv_10_40
timestamp 1595931502
transform 1 0 1472 0 1 0
box -36 -17 404 1177
use pinv_10  pinv_10_39
timestamp 1595931502
transform 1 0 0 0 -1 2240
box -36 -17 404 1177
use pinv_10  pinv_10_38
timestamp 1595931502
transform 1 0 368 0 -1 2240
box -36 -17 404 1177
use pinv_10  pinv_10_37
timestamp 1595931502
transform 1 0 736 0 -1 2240
box -36 -17 404 1177
use pinv_10  pinv_10_36
timestamp 1595931502
transform 1 0 1104 0 -1 2240
box -36 -17 404 1177
use pinv_10  pinv_10_35
timestamp 1595931502
transform 1 0 1472 0 -1 2240
box -36 -17 404 1177
use pinv_10  pinv_10_34
timestamp 1595931502
transform 1 0 0 0 1 2240
box -36 -17 404 1177
use pinv_10  pinv_10_33
timestamp 1595931502
transform 1 0 368 0 1 2240
box -36 -17 404 1177
use pinv_10  pinv_10_32
timestamp 1595931502
transform 1 0 736 0 1 2240
box -36 -17 404 1177
use pinv_10  pinv_10_31
timestamp 1595931502
transform 1 0 1104 0 1 2240
box -36 -17 404 1177
use pinv_10  pinv_10_30
timestamp 1595931502
transform 1 0 1472 0 1 2240
box -36 -17 404 1177
use pinv_10  pinv_10_29
timestamp 1595931502
transform 1 0 0 0 -1 4480
box -36 -17 404 1177
use pinv_10  pinv_10_28
timestamp 1595931502
transform 1 0 368 0 -1 4480
box -36 -17 404 1177
use pinv_10  pinv_10_27
timestamp 1595931502
transform 1 0 736 0 -1 4480
box -36 -17 404 1177
use pinv_10  pinv_10_26
timestamp 1595931502
transform 1 0 1104 0 -1 4480
box -36 -17 404 1177
use pinv_10  pinv_10_25
timestamp 1595931502
transform 1 0 1472 0 -1 4480
box -36 -17 404 1177
use pinv_10  pinv_10_24
timestamp 1595931502
transform 1 0 0 0 1 4480
box -36 -17 404 1177
use pinv_10  pinv_10_23
timestamp 1595931502
transform 1 0 368 0 1 4480
box -36 -17 404 1177
use pinv_10  pinv_10_22
timestamp 1595931502
transform 1 0 736 0 1 4480
box -36 -17 404 1177
use pinv_10  pinv_10_21
timestamp 1595931502
transform 1 0 1104 0 1 4480
box -36 -17 404 1177
use pinv_10  pinv_10_20
timestamp 1595931502
transform 1 0 1472 0 1 4480
box -36 -17 404 1177
use pinv_10  pinv_10_19
timestamp 1595931502
transform 1 0 0 0 -1 6720
box -36 -17 404 1177
use pinv_10  pinv_10_18
timestamp 1595931502
transform 1 0 368 0 -1 6720
box -36 -17 404 1177
use pinv_10  pinv_10_17
timestamp 1595931502
transform 1 0 736 0 -1 6720
box -36 -17 404 1177
use pinv_10  pinv_10_16
timestamp 1595931502
transform 1 0 1104 0 -1 6720
box -36 -17 404 1177
use pinv_10  pinv_10_15
timestamp 1595931502
transform 1 0 1472 0 -1 6720
box -36 -17 404 1177
use pinv_10  pinv_10_14
timestamp 1595931502
transform 1 0 0 0 1 6720
box -36 -17 404 1177
use pinv_10  pinv_10_13
timestamp 1595931502
transform 1 0 368 0 1 6720
box -36 -17 404 1177
use pinv_10  pinv_10_12
timestamp 1595931502
transform 1 0 736 0 1 6720
box -36 -17 404 1177
use pinv_10  pinv_10_11
timestamp 1595931502
transform 1 0 1104 0 1 6720
box -36 -17 404 1177
use pinv_10  pinv_10_10
timestamp 1595931502
transform 1 0 1472 0 1 6720
box -36 -17 404 1177
use pinv_10  pinv_10_9
timestamp 1595931502
transform 1 0 0 0 -1 8960
box -36 -17 404 1177
use pinv_10  pinv_10_8
timestamp 1595931502
transform 1 0 368 0 -1 8960
box -36 -17 404 1177
use pinv_10  pinv_10_7
timestamp 1595931502
transform 1 0 736 0 -1 8960
box -36 -17 404 1177
use pinv_10  pinv_10_6
timestamp 1595931502
transform 1 0 1104 0 -1 8960
box -36 -17 404 1177
use pinv_10  pinv_10_5
timestamp 1595931502
transform 1 0 1472 0 -1 8960
box -36 -17 404 1177
use pinv_10  pinv_10_4
timestamp 1595931502
transform 1 0 0 0 1 8960
box -36 -17 404 1177
use pinv_10  pinv_10_3
timestamp 1595931502
transform 1 0 368 0 1 8960
box -36 -17 404 1177
use pinv_10  pinv_10_2
timestamp 1595931502
transform 1 0 736 0 1 8960
box -36 -17 404 1177
use pinv_10  pinv_10_1
timestamp 1595931502
transform 1 0 1104 0 1 8960
box -36 -17 404 1177
use pinv_10  pinv_10_0
timestamp 1595931502
transform 1 0 1472 0 1 8960
box -36 -17 404 1177
use contact_8  contact_8_91
timestamp 1595931502
transform 1 0 417 0 1 490
box 0 0 64 64
use contact_8  contact_8_90
timestamp 1595931502
transform 1 0 785 0 1 490
box 0 0 64 64
use contact_8  contact_8_89
timestamp 1595931502
transform 1 0 1153 0 1 490
box 0 0 64 64
use contact_8  contact_8_88
timestamp 1595931502
transform 1 0 1521 0 1 490
box 0 0 64 64
use contact_8  contact_8_87
timestamp 1595931502
transform 1 0 49 0 1 490
box 0 0 64 64
use contact_8  contact_8_86
timestamp 1595931502
transform 1 0 164 0 1 490
box 0 0 64 64
use contact_8  contact_8_85
timestamp 1595931502
transform 1 0 417 0 1 1686
box 0 0 64 64
use contact_8  contact_8_84
timestamp 1595931502
transform 1 0 785 0 1 1686
box 0 0 64 64
use contact_8  contact_8_83
timestamp 1595931502
transform 1 0 1153 0 1 1686
box 0 0 64 64
use contact_8  contact_8_82
timestamp 1595931502
transform 1 0 1521 0 1 1686
box 0 0 64 64
use contact_8  contact_8_81
timestamp 1595931502
transform 1 0 49 0 1 1686
box 0 0 64 64
use contact_8  contact_8_80
timestamp 1595931502
transform 1 0 164 0 1 1686
box 0 0 64 64
use contact_8  contact_8_79
timestamp 1595931502
transform 1 0 417 0 1 2730
box 0 0 64 64
use contact_8  contact_8_78
timestamp 1595931502
transform 1 0 785 0 1 2730
box 0 0 64 64
use contact_8  contact_8_77
timestamp 1595931502
transform 1 0 1153 0 1 2730
box 0 0 64 64
use contact_8  contact_8_76
timestamp 1595931502
transform 1 0 1521 0 1 2730
box 0 0 64 64
use contact_8  contact_8_75
timestamp 1595931502
transform 1 0 49 0 1 2730
box 0 0 64 64
use contact_8  contact_8_74
timestamp 1595931502
transform 1 0 164 0 1 2730
box 0 0 64 64
use contact_8  contact_8_73
timestamp 1595931502
transform 1 0 417 0 1 3926
box 0 0 64 64
use contact_8  contact_8_72
timestamp 1595931502
transform 1 0 785 0 1 3926
box 0 0 64 64
use contact_8  contact_8_71
timestamp 1595931502
transform 1 0 1153 0 1 3926
box 0 0 64 64
use contact_8  contact_8_70
timestamp 1595931502
transform 1 0 1521 0 1 3926
box 0 0 64 64
use contact_8  contact_8_69
timestamp 1595931502
transform 1 0 49 0 1 3926
box 0 0 64 64
use contact_8  contact_8_68
timestamp 1595931502
transform 1 0 164 0 1 3926
box 0 0 64 64
use contact_8  contact_8_67
timestamp 1595931502
transform 1 0 417 0 1 4970
box 0 0 64 64
use contact_8  contact_8_66
timestamp 1595931502
transform 1 0 785 0 1 4970
box 0 0 64 64
use contact_8  contact_8_65
timestamp 1595931502
transform 1 0 1153 0 1 4970
box 0 0 64 64
use contact_8  contact_8_64
timestamp 1595931502
transform 1 0 1521 0 1 4970
box 0 0 64 64
use contact_8  contact_8_63
timestamp 1595931502
transform 1 0 49 0 1 4970
box 0 0 64 64
use contact_8  contact_8_62
timestamp 1595931502
transform 1 0 164 0 1 4970
box 0 0 64 64
use contact_8  contact_8_61
timestamp 1595931502
transform 1 0 417 0 1 6166
box 0 0 64 64
use contact_8  contact_8_60
timestamp 1595931502
transform 1 0 785 0 1 6166
box 0 0 64 64
use contact_8  contact_8_59
timestamp 1595931502
transform 1 0 1153 0 1 6166
box 0 0 64 64
use contact_8  contact_8_58
timestamp 1595931502
transform 1 0 1521 0 1 6166
box 0 0 64 64
use contact_8  contact_8_57
timestamp 1595931502
transform 1 0 49 0 1 6166
box 0 0 64 64
use contact_8  contact_8_56
timestamp 1595931502
transform 1 0 164 0 1 6166
box 0 0 64 64
use contact_8  contact_8_55
timestamp 1595931502
transform 1 0 417 0 1 7210
box 0 0 64 64
use contact_8  contact_8_54
timestamp 1595931502
transform 1 0 785 0 1 7210
box 0 0 64 64
use contact_8  contact_8_53
timestamp 1595931502
transform 1 0 1153 0 1 7210
box 0 0 64 64
use contact_8  contact_8_52
timestamp 1595931502
transform 1 0 1521 0 1 7210
box 0 0 64 64
use contact_8  contact_8_51
timestamp 1595931502
transform 1 0 49 0 1 7210
box 0 0 64 64
use contact_8  contact_8_50
timestamp 1595931502
transform 1 0 164 0 1 7210
box 0 0 64 64
use contact_8  contact_8_49
timestamp 1595931502
transform 1 0 417 0 1 8406
box 0 0 64 64
use contact_8  contact_8_48
timestamp 1595931502
transform 1 0 785 0 1 8406
box 0 0 64 64
use contact_8  contact_8_47
timestamp 1595931502
transform 1 0 1153 0 1 8406
box 0 0 64 64
use contact_8  contact_8_46
timestamp 1595931502
transform 1 0 1521 0 1 8406
box 0 0 64 64
use contact_8  contact_8_45
timestamp 1595931502
transform 1 0 49 0 1 8406
box 0 0 64 64
use contact_8  contact_8_44
timestamp 1595931502
transform 1 0 164 0 1 8406
box 0 0 64 64
use contact_8  contact_8_43
timestamp 1595931502
transform 1 0 417 0 1 9450
box 0 0 64 64
use contact_8  contact_8_42
timestamp 1595931502
transform 1 0 785 0 1 9450
box 0 0 64 64
use contact_8  contact_8_41
timestamp 1595931502
transform 1 0 1153 0 1 9450
box 0 0 64 64
use contact_8  contact_8_40
timestamp 1595931502
transform 1 0 1521 0 1 9450
box 0 0 64 64
use contact_8  contact_8_39
timestamp 1595931502
transform 1 0 49 0 1 9450
box 0 0 64 64
use contact_8  contact_8_38
timestamp 1595931502
transform 1 0 164 0 1 9450
box 0 0 64 64
use contact_8  contact_8_37
timestamp 1595931502
transform 1 0 624 0 1 1088
box 0 0 64 64
use contact_8  contact_8_36
timestamp 1595931502
transform 1 0 1360 0 1 1088
box 0 0 64 64
use contact_8  contact_8_35
timestamp 1595931502
transform 1 0 624 0 1 -32
box 0 0 64 64
use contact_8  contact_8_34
timestamp 1595931502
transform 1 0 1360 0 1 -32
box 0 0 64 64
use contact_8  contact_8_33
timestamp 1595931502
transform 1 0 624 0 1 1088
box 0 0 64 64
use contact_8  contact_8_32
timestamp 1595931502
transform 1 0 1360 0 1 1088
box 0 0 64 64
use contact_8  contact_8_31
timestamp 1595931502
transform 1 0 624 0 1 2208
box 0 0 64 64
use contact_8  contact_8_30
timestamp 1595931502
transform 1 0 1360 0 1 2208
box 0 0 64 64
use contact_8  contact_8_29
timestamp 1595931502
transform 1 0 624 0 1 3328
box 0 0 64 64
use contact_8  contact_8_28
timestamp 1595931502
transform 1 0 1360 0 1 3328
box 0 0 64 64
use contact_8  contact_8_27
timestamp 1595931502
transform 1 0 624 0 1 2208
box 0 0 64 64
use contact_8  contact_8_26
timestamp 1595931502
transform 1 0 1360 0 1 2208
box 0 0 64 64
use contact_8  contact_8_25
timestamp 1595931502
transform 1 0 624 0 1 3328
box 0 0 64 64
use contact_8  contact_8_24
timestamp 1595931502
transform 1 0 1360 0 1 3328
box 0 0 64 64
use contact_8  contact_8_23
timestamp 1595931502
transform 1 0 624 0 1 4448
box 0 0 64 64
use contact_8  contact_8_22
timestamp 1595931502
transform 1 0 1360 0 1 4448
box 0 0 64 64
use contact_8  contact_8_21
timestamp 1595931502
transform 1 0 624 0 1 5568
box 0 0 64 64
use contact_8  contact_8_20
timestamp 1595931502
transform 1 0 1360 0 1 5568
box 0 0 64 64
use contact_8  contact_8_19
timestamp 1595931502
transform 1 0 624 0 1 4448
box 0 0 64 64
use contact_8  contact_8_18
timestamp 1595931502
transform 1 0 1360 0 1 4448
box 0 0 64 64
use contact_8  contact_8_17
timestamp 1595931502
transform 1 0 624 0 1 5568
box 0 0 64 64
use contact_8  contact_8_16
timestamp 1595931502
transform 1 0 1360 0 1 5568
box 0 0 64 64
use contact_8  contact_8_15
timestamp 1595931502
transform 1 0 624 0 1 6688
box 0 0 64 64
use contact_8  contact_8_14
timestamp 1595931502
transform 1 0 1360 0 1 6688
box 0 0 64 64
use contact_8  contact_8_13
timestamp 1595931502
transform 1 0 624 0 1 7808
box 0 0 64 64
use contact_8  contact_8_12
timestamp 1595931502
transform 1 0 1360 0 1 7808
box 0 0 64 64
use contact_8  contact_8_11
timestamp 1595931502
transform 1 0 624 0 1 6688
box 0 0 64 64
use contact_8  contact_8_10
timestamp 1595931502
transform 1 0 1360 0 1 6688
box 0 0 64 64
use contact_8  contact_8_9
timestamp 1595931502
transform 1 0 624 0 1 7808
box 0 0 64 64
use contact_8  contact_8_8
timestamp 1595931502
transform 1 0 1360 0 1 7808
box 0 0 64 64
use contact_8  contact_8_7
timestamp 1595931502
transform 1 0 624 0 1 8928
box 0 0 64 64
use contact_8  contact_8_6
timestamp 1595931502
transform 1 0 1360 0 1 8928
box 0 0 64 64
use contact_8  contact_8_5
timestamp 1595931502
transform 1 0 624 0 1 10048
box 0 0 64 64
use contact_8  contact_8_4
timestamp 1595931502
transform 1 0 1360 0 1 10048
box 0 0 64 64
use contact_8  contact_8_3
timestamp 1595931502
transform 1 0 624 0 1 8928
box 0 0 64 64
use contact_8  contact_8_2
timestamp 1595931502
transform 1 0 1360 0 1 8928
box 0 0 64 64
use contact_8  contact_8_1
timestamp 1595931502
transform 1 0 49 0 1 490
box 0 0 64 64
use contact_8  contact_8_0
timestamp 1595931502
transform 1 0 1521 0 1 9450
box 0 0 64 64
use contact_7  contact_7_91
timestamp 1595931502
transform 1 0 420 0 1 489
box 0 0 58 66
use contact_7  contact_7_90
timestamp 1595931502
transform 1 0 788 0 1 489
box 0 0 58 66
use contact_7  contact_7_89
timestamp 1595931502
transform 1 0 1156 0 1 489
box 0 0 58 66
use contact_7  contact_7_88
timestamp 1595931502
transform 1 0 1524 0 1 489
box 0 0 58 66
use contact_7  contact_7_87
timestamp 1595931502
transform 1 0 52 0 1 489
box 0 0 58 66
use contact_7  contact_7_86
timestamp 1595931502
transform 1 0 167 0 1 489
box 0 0 58 66
use contact_7  contact_7_85
timestamp 1595931502
transform 1 0 420 0 1 1685
box 0 0 58 66
use contact_7  contact_7_84
timestamp 1595931502
transform 1 0 788 0 1 1685
box 0 0 58 66
use contact_7  contact_7_83
timestamp 1595931502
transform 1 0 1156 0 1 1685
box 0 0 58 66
use contact_7  contact_7_82
timestamp 1595931502
transform 1 0 1524 0 1 1685
box 0 0 58 66
use contact_7  contact_7_81
timestamp 1595931502
transform 1 0 52 0 1 1685
box 0 0 58 66
use contact_7  contact_7_80
timestamp 1595931502
transform 1 0 167 0 1 1685
box 0 0 58 66
use contact_7  contact_7_79
timestamp 1595931502
transform 1 0 420 0 1 2729
box 0 0 58 66
use contact_7  contact_7_78
timestamp 1595931502
transform 1 0 788 0 1 2729
box 0 0 58 66
use contact_7  contact_7_77
timestamp 1595931502
transform 1 0 1156 0 1 2729
box 0 0 58 66
use contact_7  contact_7_76
timestamp 1595931502
transform 1 0 1524 0 1 2729
box 0 0 58 66
use contact_7  contact_7_75
timestamp 1595931502
transform 1 0 52 0 1 2729
box 0 0 58 66
use contact_7  contact_7_74
timestamp 1595931502
transform 1 0 167 0 1 2729
box 0 0 58 66
use contact_7  contact_7_73
timestamp 1595931502
transform 1 0 420 0 1 3925
box 0 0 58 66
use contact_7  contact_7_72
timestamp 1595931502
transform 1 0 788 0 1 3925
box 0 0 58 66
use contact_7  contact_7_71
timestamp 1595931502
transform 1 0 1156 0 1 3925
box 0 0 58 66
use contact_7  contact_7_70
timestamp 1595931502
transform 1 0 1524 0 1 3925
box 0 0 58 66
use contact_7  contact_7_69
timestamp 1595931502
transform 1 0 52 0 1 3925
box 0 0 58 66
use contact_7  contact_7_68
timestamp 1595931502
transform 1 0 167 0 1 3925
box 0 0 58 66
use contact_7  contact_7_67
timestamp 1595931502
transform 1 0 420 0 1 4969
box 0 0 58 66
use contact_7  contact_7_66
timestamp 1595931502
transform 1 0 788 0 1 4969
box 0 0 58 66
use contact_7  contact_7_65
timestamp 1595931502
transform 1 0 1156 0 1 4969
box 0 0 58 66
use contact_7  contact_7_64
timestamp 1595931502
transform 1 0 1524 0 1 4969
box 0 0 58 66
use contact_7  contact_7_63
timestamp 1595931502
transform 1 0 52 0 1 4969
box 0 0 58 66
use contact_7  contact_7_62
timestamp 1595931502
transform 1 0 167 0 1 4969
box 0 0 58 66
use contact_7  contact_7_61
timestamp 1595931502
transform 1 0 420 0 1 6165
box 0 0 58 66
use contact_7  contact_7_60
timestamp 1595931502
transform 1 0 788 0 1 6165
box 0 0 58 66
use contact_7  contact_7_59
timestamp 1595931502
transform 1 0 1156 0 1 6165
box 0 0 58 66
use contact_7  contact_7_58
timestamp 1595931502
transform 1 0 1524 0 1 6165
box 0 0 58 66
use contact_7  contact_7_57
timestamp 1595931502
transform 1 0 52 0 1 6165
box 0 0 58 66
use contact_7  contact_7_56
timestamp 1595931502
transform 1 0 167 0 1 6165
box 0 0 58 66
use contact_7  contact_7_55
timestamp 1595931502
transform 1 0 420 0 1 7209
box 0 0 58 66
use contact_7  contact_7_54
timestamp 1595931502
transform 1 0 788 0 1 7209
box 0 0 58 66
use contact_7  contact_7_53
timestamp 1595931502
transform 1 0 1156 0 1 7209
box 0 0 58 66
use contact_7  contact_7_52
timestamp 1595931502
transform 1 0 1524 0 1 7209
box 0 0 58 66
use contact_7  contact_7_51
timestamp 1595931502
transform 1 0 52 0 1 7209
box 0 0 58 66
use contact_7  contact_7_50
timestamp 1595931502
transform 1 0 167 0 1 7209
box 0 0 58 66
use contact_7  contact_7_49
timestamp 1595931502
transform 1 0 420 0 1 8405
box 0 0 58 66
use contact_7  contact_7_48
timestamp 1595931502
transform 1 0 788 0 1 8405
box 0 0 58 66
use contact_7  contact_7_47
timestamp 1595931502
transform 1 0 1156 0 1 8405
box 0 0 58 66
use contact_7  contact_7_46
timestamp 1595931502
transform 1 0 1524 0 1 8405
box 0 0 58 66
use contact_7  contact_7_45
timestamp 1595931502
transform 1 0 52 0 1 8405
box 0 0 58 66
use contact_7  contact_7_44
timestamp 1595931502
transform 1 0 167 0 1 8405
box 0 0 58 66
use contact_7  contact_7_43
timestamp 1595931502
transform 1 0 420 0 1 9449
box 0 0 58 66
use contact_7  contact_7_42
timestamp 1595931502
transform 1 0 788 0 1 9449
box 0 0 58 66
use contact_7  contact_7_41
timestamp 1595931502
transform 1 0 1156 0 1 9449
box 0 0 58 66
use contact_7  contact_7_40
timestamp 1595931502
transform 1 0 1524 0 1 9449
box 0 0 58 66
use contact_7  contact_7_39
timestamp 1595931502
transform 1 0 52 0 1 9449
box 0 0 58 66
use contact_7  contact_7_38
timestamp 1595931502
transform 1 0 167 0 1 9449
box 0 0 58 66
use contact_7  contact_7_37
timestamp 1595931502
transform 1 0 627 0 1 1087
box 0 0 58 66
use contact_7  contact_7_36
timestamp 1595931502
transform 1 0 1363 0 1 1087
box 0 0 58 66
use contact_7  contact_7_35
timestamp 1595931502
transform 1 0 627 0 1 -33
box 0 0 58 66
use contact_7  contact_7_34
timestamp 1595931502
transform 1 0 1363 0 1 -33
box 0 0 58 66
use contact_7  contact_7_33
timestamp 1595931502
transform 1 0 627 0 1 1087
box 0 0 58 66
use contact_7  contact_7_32
timestamp 1595931502
transform 1 0 1363 0 1 1087
box 0 0 58 66
use contact_7  contact_7_31
timestamp 1595931502
transform 1 0 627 0 1 2207
box 0 0 58 66
use contact_7  contact_7_30
timestamp 1595931502
transform 1 0 1363 0 1 2207
box 0 0 58 66
use contact_7  contact_7_29
timestamp 1595931502
transform 1 0 627 0 1 3327
box 0 0 58 66
use contact_7  contact_7_28
timestamp 1595931502
transform 1 0 1363 0 1 3327
box 0 0 58 66
use contact_7  contact_7_27
timestamp 1595931502
transform 1 0 627 0 1 2207
box 0 0 58 66
use contact_7  contact_7_26
timestamp 1595931502
transform 1 0 1363 0 1 2207
box 0 0 58 66
use contact_7  contact_7_25
timestamp 1595931502
transform 1 0 627 0 1 3327
box 0 0 58 66
use contact_7  contact_7_24
timestamp 1595931502
transform 1 0 1363 0 1 3327
box 0 0 58 66
use contact_7  contact_7_23
timestamp 1595931502
transform 1 0 627 0 1 4447
box 0 0 58 66
use contact_7  contact_7_22
timestamp 1595931502
transform 1 0 1363 0 1 4447
box 0 0 58 66
use contact_7  contact_7_21
timestamp 1595931502
transform 1 0 627 0 1 5567
box 0 0 58 66
use contact_7  contact_7_20
timestamp 1595931502
transform 1 0 1363 0 1 5567
box 0 0 58 66
use contact_7  contact_7_19
timestamp 1595931502
transform 1 0 627 0 1 4447
box 0 0 58 66
use contact_7  contact_7_18
timestamp 1595931502
transform 1 0 1363 0 1 4447
box 0 0 58 66
use contact_7  contact_7_17
timestamp 1595931502
transform 1 0 627 0 1 5567
box 0 0 58 66
use contact_7  contact_7_16
timestamp 1595931502
transform 1 0 1363 0 1 5567
box 0 0 58 66
use contact_7  contact_7_15
timestamp 1595931502
transform 1 0 627 0 1 6687
box 0 0 58 66
use contact_7  contact_7_14
timestamp 1595931502
transform 1 0 1363 0 1 6687
box 0 0 58 66
use contact_7  contact_7_13
timestamp 1595931502
transform 1 0 627 0 1 7807
box 0 0 58 66
use contact_7  contact_7_12
timestamp 1595931502
transform 1 0 1363 0 1 7807
box 0 0 58 66
use contact_7  contact_7_11
timestamp 1595931502
transform 1 0 627 0 1 6687
box 0 0 58 66
use contact_7  contact_7_10
timestamp 1595931502
transform 1 0 1363 0 1 6687
box 0 0 58 66
use contact_7  contact_7_9
timestamp 1595931502
transform 1 0 627 0 1 7807
box 0 0 58 66
use contact_7  contact_7_8
timestamp 1595931502
transform 1 0 1363 0 1 7807
box 0 0 58 66
use contact_7  contact_7_7
timestamp 1595931502
transform 1 0 627 0 1 8927
box 0 0 58 66
use contact_7  contact_7_6
timestamp 1595931502
transform 1 0 1363 0 1 8927
box 0 0 58 66
use contact_7  contact_7_5
timestamp 1595931502
transform 1 0 627 0 1 10047
box 0 0 58 66
use contact_7  contact_7_4
timestamp 1595931502
transform 1 0 1363 0 1 10047
box 0 0 58 66
use contact_7  contact_7_3
timestamp 1595931502
transform 1 0 627 0 1 8927
box 0 0 58 66
use contact_7  contact_7_2
timestamp 1595931502
transform 1 0 1363 0 1 8927
box 0 0 58 66
use contact_7  contact_7_1
timestamp 1595931502
transform 1 0 52 0 1 489
box 0 0 58 66
use contact_7  contact_7_0
timestamp 1595931502
transform 1 0 1524 0 1 9449
box 0 0 58 66
<< labels >>
rlabel metal3 s 1392 4480 1392 4480 4 gnd
rlabel metal3 s 1392 6720 1392 6720 4 gnd
rlabel metal3 s 1392 2240 1392 2240 4 gnd
rlabel metal3 s 1392 8960 1392 8960 4 gnd
rlabel metal3 s 656 6720 656 6720 4 gnd
rlabel metal3 s 656 2240 656 2240 4 gnd
rlabel metal3 s 656 4480 656 4480 4 gnd
rlabel metal3 s 656 0 656 0 4 gnd
rlabel metal3 s 656 8960 656 8960 4 gnd
rlabel metal3 s 1392 0 1392 0 4 gnd
rlabel metal2 s 78 261 78 261 4 in
rlabel metal2 s 1637 4741 1637 4741 4 out
rlabel metal3 s 1392 3360 1392 3360 4 vdd
rlabel metal3 s 1392 3360 1392 3360 4 vdd
rlabel metal3 s 656 7840 656 7840 4 vdd
rlabel metal3 s 1392 10080 1392 10080 4 vdd
rlabel metal3 s 1392 1120 1392 1120 4 vdd
rlabel metal3 s 1392 1120 1392 1120 4 vdd
rlabel metal3 s 1392 5600 1392 5600 4 vdd
rlabel metal3 s 656 1120 656 1120 4 vdd
rlabel metal3 s 656 10080 656 10080 4 vdd
rlabel metal3 s 1392 7840 1392 7840 4 vdd
rlabel metal3 s 656 5600 656 5600 4 vdd
rlabel metal3 s 656 3360 656 3360 4 vdd
rlabel metal3 s 656 3360 656 3360 4 vdd
rlabel metal3 s 656 1120 656 1120 4 vdd
<< properties >>
string FIXED_BBOX 0 0 1840 10080
<< end >>
