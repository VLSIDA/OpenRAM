VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 1000 ;
END UNITS
SITE  MacroSite
   CLASS Core ;
   SIZE 324000.0 by 421500.0 ;
END  MacroSite
MACRO sram1
   CLASS BLOCK ;
   SIZE 324000.0 BY 421500.0 ;
   SYMMETRY X Y R90 ;
   SITE MacroSite ;
   PIN DIN[0]
      DIRECTION INPUT ;
      PORT
