VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 1000 ;
END UNITS
SITE  MacroSite
   CLASS Core ;
   SIZE 2250.0 by 1200.0 ;
END  MacroSite
MACRO sram_2_16_1_scn3me_subm
   CLASS BLOCK ;
   SIZE 2250.0 BY 1200.0 ;
   SYMMETRY X Y R90 ;
   SITE MacroSite ;
   PIN DATA[0]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  180000.0 0.0 180900.0 1800.0 ;
      END
   END DATA[0]
   PIN DATA[1]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  190200.0 0.0 191100.0 1800.0 ;
      END
   END DATA[1]
   PIN ADDR[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  52800.0 77400.0 60000.0 78900.0 ;
      END
   END ADDR[0]
   PIN ADDR[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  52800.0 67200.0 60000.0 68700.0 ;
      END
   END ADDR[1]
   PIN ADDR[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  52800.0 57000.0 60000.0 58500.0 ;
      END
   END ADDR[2]
   PIN ADDR[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  52800.0 46800.0 60000.0 48300.0 ;
      END
   END ADDR[3]
   PIN CSb
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  14400.0 203100.0 16200.0 204900.0 ;
      END
   END CSb
   PIN WEb
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  24600.0 203100.0 26400.0 204900.0 ;
      END
   END WEb
   PIN OEb
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  4200.0 203100.0 6000.0 204900.0 ;
      END
   END OEb
   PIN clk
      DIRECTION INPUT ;
      PORT
         LAYER metal1 ;
         RECT  42600.0 202200.0 43800.0 205800.0 ;
      END
   END clk
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal1 ;
         RECT  198600.0 0.0 203100.0 436800.0 ;
         LAYER metal1 ;
         RECT  52800.0 0.0 57300.0 436800.0 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal2 ;
         RECT  148050.0 0.0 152550.0 436800.0 ;
      END
   END gnd
   OBS
   LAYER  metal1 ;
      RECT  54600.0 295650.0 55500.0 298350.0 ;
      RECT  97500.0 205350.0 98400.0 206250.0 ;
      RECT  97500.0 202950.0 98400.0 203850.0 ;
      RECT  96150.0 205350.0 97950.0 206250.0 ;
      RECT  97500.0 203400.0 98400.0 205800.0 ;
      RECT  97950.0 202950.0 99900.0 203850.0 ;
      RECT  154950.0 205350.0 155850.0 206250.0 ;
      RECT  154950.0 200850.0 155850.0 201750.0 ;
      RECT  136050.0 205350.0 155400.0 206250.0 ;
      RECT  154950.0 201300.0 155850.0 205800.0 ;
      RECT  155400.0 200850.0 174900.0 201750.0 ;
      RECT  97500.0 219750.0 98400.0 220650.0 ;
      RECT  97500.0 222150.0 98400.0 223050.0 ;
      RECT  96150.0 219750.0 97950.0 220650.0 ;
      RECT  97500.0 220200.0 98400.0 222600.0 ;
      RECT  97950.0 222150.0 99900.0 223050.0 ;
      RECT  154950.0 219750.0 155850.0 220650.0 ;
      RECT  154950.0 224250.0 155850.0 225150.0 ;
      RECT  136050.0 219750.0 155400.0 220650.0 ;
      RECT  154950.0 220200.0 155850.0 224700.0 ;
      RECT  155400.0 224250.0 174900.0 225150.0 ;
      RECT  97500.0 232950.0 98400.0 233850.0 ;
      RECT  97500.0 230550.0 98400.0 231450.0 ;
      RECT  96150.0 232950.0 97950.0 233850.0 ;
      RECT  97500.0 231000.0 98400.0 233400.0 ;
      RECT  97950.0 230550.0 99900.0 231450.0 ;
      RECT  154950.0 232950.0 155850.0 233850.0 ;
      RECT  154950.0 228450.0 155850.0 229350.0 ;
      RECT  136050.0 232950.0 155400.0 233850.0 ;
      RECT  154950.0 228900.0 155850.0 233400.0 ;
      RECT  155400.0 228450.0 174900.0 229350.0 ;
      RECT  97500.0 247350.0 98400.0 248250.0 ;
      RECT  97500.0 249750.0 98400.0 250650.0 ;
      RECT  96150.0 247350.0 97950.0 248250.0 ;
      RECT  97500.0 247800.0 98400.0 250200.0 ;
      RECT  97950.0 249750.0 99900.0 250650.0 ;
      RECT  154950.0 247350.0 155850.0 248250.0 ;
      RECT  154950.0 251850.0 155850.0 252750.0 ;
      RECT  136050.0 247350.0 155400.0 248250.0 ;
      RECT  154950.0 247800.0 155850.0 252300.0 ;
      RECT  155400.0 251850.0 174900.0 252750.0 ;
      RECT  97500.0 260550.0 98400.0 261450.0 ;
      RECT  97500.0 258150.0 98400.0 259050.0 ;
      RECT  96150.0 260550.0 97950.0 261450.0 ;
      RECT  97500.0 258600.0 98400.0 261000.0 ;
      RECT  97950.0 258150.0 99900.0 259050.0 ;
      RECT  154950.0 260550.0 155850.0 261450.0 ;
      RECT  154950.0 256050.0 155850.0 256950.0 ;
      RECT  136050.0 260550.0 155400.0 261450.0 ;
      RECT  154950.0 256500.0 155850.0 261000.0 ;
      RECT  155400.0 256050.0 174900.0 256950.0 ;
      RECT  97500.0 274950.0 98400.0 275850.0 ;
      RECT  97500.0 277350.0 98400.0 278250.0 ;
      RECT  96150.0 274950.0 97950.0 275850.0 ;
      RECT  97500.0 275400.0 98400.0 277800.0 ;
      RECT  97950.0 277350.0 99900.0 278250.0 ;
      RECT  154950.0 274950.0 155850.0 275850.0 ;
      RECT  154950.0 279450.0 155850.0 280350.0 ;
      RECT  136050.0 274950.0 155400.0 275850.0 ;
      RECT  154950.0 275400.0 155850.0 279900.0 ;
      RECT  155400.0 279450.0 174900.0 280350.0 ;
      RECT  97500.0 288150.0 98400.0 289050.0 ;
      RECT  97500.0 285750.0 98400.0 286650.0 ;
      RECT  96150.0 288150.0 97950.0 289050.0 ;
      RECT  97500.0 286200.0 98400.0 288600.0 ;
      RECT  97950.0 285750.0 99900.0 286650.0 ;
      RECT  154950.0 288150.0 155850.0 289050.0 ;
      RECT  154950.0 283650.0 155850.0 284550.0 ;
      RECT  136050.0 288150.0 155400.0 289050.0 ;
      RECT  154950.0 284100.0 155850.0 288600.0 ;
      RECT  155400.0 283650.0 174900.0 284550.0 ;
      RECT  97500.0 302550.0 98400.0 303450.0 ;
      RECT  97500.0 304950.0 98400.0 305850.0 ;
      RECT  96150.0 302550.0 97950.0 303450.0 ;
      RECT  97500.0 303000.0 98400.0 305400.0 ;
      RECT  97950.0 304950.0 99900.0 305850.0 ;
      RECT  154950.0 302550.0 155850.0 303450.0 ;
      RECT  154950.0 307050.0 155850.0 307950.0 ;
      RECT  136050.0 302550.0 155400.0 303450.0 ;
      RECT  154950.0 303000.0 155850.0 307500.0 ;
      RECT  155400.0 307050.0 174900.0 307950.0 ;
      RECT  97500.0 315750.0 98400.0 316650.0 ;
      RECT  97500.0 313350.0 98400.0 314250.0 ;
      RECT  96150.0 315750.0 97950.0 316650.0 ;
      RECT  97500.0 313800.0 98400.0 316200.0 ;
      RECT  97950.0 313350.0 99900.0 314250.0 ;
      RECT  154950.0 315750.0 155850.0 316650.0 ;
      RECT  154950.0 311250.0 155850.0 312150.0 ;
      RECT  136050.0 315750.0 155400.0 316650.0 ;
      RECT  154950.0 311700.0 155850.0 316200.0 ;
      RECT  155400.0 311250.0 174900.0 312150.0 ;
      RECT  97500.0 330150.0 98400.0 331050.0 ;
      RECT  97500.0 332550.0 98400.0 333450.0 ;
      RECT  96150.0 330150.0 97950.0 331050.0 ;
      RECT  97500.0 330600.0 98400.0 333000.0 ;
      RECT  97950.0 332550.0 99900.0 333450.0 ;
      RECT  154950.0 330150.0 155850.0 331050.0 ;
      RECT  154950.0 334650.0 155850.0 335550.0 ;
      RECT  136050.0 330150.0 155400.0 331050.0 ;
      RECT  154950.0 330600.0 155850.0 335100.0 ;
      RECT  155400.0 334650.0 174900.0 335550.0 ;
      RECT  97500.0 343350.0 98400.0 344250.0 ;
      RECT  97500.0 340950.0 98400.0 341850.0 ;
      RECT  96150.0 343350.0 97950.0 344250.0 ;
      RECT  97500.0 341400.0 98400.0 343800.0 ;
      RECT  97950.0 340950.0 99900.0 341850.0 ;
      RECT  154950.0 343350.0 155850.0 344250.0 ;
      RECT  154950.0 338850.0 155850.0 339750.0 ;
      RECT  136050.0 343350.0 155400.0 344250.0 ;
      RECT  154950.0 339300.0 155850.0 343800.0 ;
      RECT  155400.0 338850.0 174900.0 339750.0 ;
      RECT  97500.0 357750.0 98400.0 358650.0 ;
      RECT  97500.0 360150.0 98400.0 361050.0 ;
      RECT  96150.0 357750.0 97950.0 358650.0 ;
      RECT  97500.0 358200.0 98400.0 360600.0 ;
      RECT  97950.0 360150.0 99900.0 361050.0 ;
      RECT  154950.0 357750.0 155850.0 358650.0 ;
      RECT  154950.0 362250.0 155850.0 363150.0 ;
      RECT  136050.0 357750.0 155400.0 358650.0 ;
      RECT  154950.0 358200.0 155850.0 362700.0 ;
      RECT  155400.0 362250.0 174900.0 363150.0 ;
      RECT  97500.0 370950.0 98400.0 371850.0 ;
      RECT  97500.0 368550.0 98400.0 369450.0 ;
      RECT  96150.0 370950.0 97950.0 371850.0 ;
      RECT  97500.0 369000.0 98400.0 371400.0 ;
      RECT  97950.0 368550.0 99900.0 369450.0 ;
      RECT  154950.0 370950.0 155850.0 371850.0 ;
      RECT  154950.0 366450.0 155850.0 367350.0 ;
      RECT  136050.0 370950.0 155400.0 371850.0 ;
      RECT  154950.0 366900.0 155850.0 371400.0 ;
      RECT  155400.0 366450.0 174900.0 367350.0 ;
      RECT  97500.0 385350.0 98400.0 386250.0 ;
      RECT  97500.0 387750.0 98400.0 388650.0 ;
      RECT  96150.0 385350.0 97950.0 386250.0 ;
      RECT  97500.0 385800.0 98400.0 388200.0 ;
      RECT  97950.0 387750.0 99900.0 388650.0 ;
      RECT  154950.0 385350.0 155850.0 386250.0 ;
      RECT  154950.0 389850.0 155850.0 390750.0 ;
      RECT  136050.0 385350.0 155400.0 386250.0 ;
      RECT  154950.0 385800.0 155850.0 390300.0 ;
      RECT  155400.0 389850.0 174900.0 390750.0 ;
      RECT  97500.0 398550.0 98400.0 399450.0 ;
      RECT  97500.0 396150.0 98400.0 397050.0 ;
      RECT  96150.0 398550.0 97950.0 399450.0 ;
      RECT  97500.0 396600.0 98400.0 399000.0 ;
      RECT  97950.0 396150.0 99900.0 397050.0 ;
      RECT  154950.0 398550.0 155850.0 399450.0 ;
      RECT  154950.0 394050.0 155850.0 394950.0 ;
      RECT  136050.0 398550.0 155400.0 399450.0 ;
      RECT  154950.0 394500.0 155850.0 399000.0 ;
      RECT  155400.0 394050.0 174900.0 394950.0 ;
      RECT  97500.0 412950.0 98400.0 413850.0 ;
      RECT  97500.0 415350.0 98400.0 416250.0 ;
      RECT  96150.0 412950.0 97950.0 413850.0 ;
      RECT  97500.0 413400.0 98400.0 415800.0 ;
      RECT  97950.0 415350.0 99900.0 416250.0 ;
      RECT  154950.0 412950.0 155850.0 413850.0 ;
      RECT  154950.0 417450.0 155850.0 418350.0 ;
      RECT  136050.0 412950.0 155400.0 413850.0 ;
      RECT  154950.0 413400.0 155850.0 417900.0 ;
      RECT  155400.0 417450.0 174900.0 418350.0 ;
      RECT  106200.0 198750.0 175500.0 199650.0 ;
      RECT  106200.0 226350.0 175500.0 227250.0 ;
      RECT  106200.0 253950.0 175500.0 254850.0 ;
      RECT  106200.0 281550.0 175500.0 282450.0 ;
      RECT  106200.0 309150.0 175500.0 310050.0 ;
      RECT  106200.0 336750.0 175500.0 337650.0 ;
      RECT  106200.0 364350.0 175500.0 365250.0 ;
      RECT  106200.0 391950.0 175500.0 392850.0 ;
      RECT  106200.0 419550.0 175500.0 420450.0 ;
      RECT  52800.0 212550.0 203100.0 213450.0 ;
      RECT  52800.0 240150.0 203100.0 241050.0 ;
      RECT  52800.0 267750.0 203100.0 268650.0 ;
      RECT  52800.0 295350.0 203100.0 296250.0 ;
      RECT  52800.0 322950.0 203100.0 323850.0 ;
      RECT  52800.0 350550.0 203100.0 351450.0 ;
      RECT  52800.0 378150.0 203100.0 379050.0 ;
      RECT  52800.0 405750.0 203100.0 406650.0 ;
      RECT  130500.0 91050.0 135000.0 91950.0 ;
      RECT  127500.0 104850.0 137700.0 105750.0 ;
      RECT  130500.0 146250.0 140400.0 147150.0 ;
      RECT  127500.0 160050.0 143100.0 160950.0 ;
      RECT  130500.0 88350.0 132000.0 89250.0 ;
      RECT  130500.0 115950.0 132000.0 116850.0 ;
      RECT  130500.0 143550.0 132000.0 144450.0 ;
      RECT  130500.0 171150.0 132000.0 172050.0 ;
      RECT  52800.0 102150.0 130500.0 103050.0 ;
      RECT  52800.0 129750.0 130500.0 130650.0 ;
      RECT  52800.0 157350.0 130500.0 158250.0 ;
      RECT  52800.0 184950.0 130500.0 185850.0 ;
      RECT  117900.0 77100.0 135000.0 78000.0 ;
      RECT  117900.0 68400.0 137700.0 69300.0 ;
      RECT  117900.0 56700.0 140400.0 57600.0 ;
      RECT  117900.0 48000.0 143100.0 48900.0 ;
      RECT  119100.0 72750.0 149250.0 73650.0 ;
      RECT  119100.0 52350.0 149250.0 53250.0 ;
      RECT  115500.0 40050.0 116400.0 40950.0 ;
      RECT  115500.0 40500.0 116400.0 42600.0 ;
      RECT  52800.0 40050.0 115950.0 40950.0 ;
      RECT  163800.0 32400.0 175500.0 33300.0 ;
      RECT  158400.0 27900.0 175500.0 28800.0 ;
      RECT  161100.0 25500.0 175500.0 26400.0 ;
      RECT  163800.0 424800.0 175500.0 425700.0 ;
      RECT  166500.0 96900.0 175500.0 97800.0 ;
      RECT  169200.0 195000.0 175500.0 195900.0 ;
      RECT  61500.0 85050.0 62400.0 85950.0 ;
      RECT  61500.0 83400.0 62400.0 85500.0 ;
      RECT  61950.0 85050.0 155700.0 85950.0 ;
      RECT  103050.0 421650.0 156600.0 422550.0 ;
      RECT  175500.0 435900.0 198600.0 436800.0 ;
      RECT  175500.0 167700.0 198600.0 168600.0 ;
      RECT  175500.0 99000.0 198600.0 99900.0 ;
      RECT  175500.0 86400.0 198600.0 87300.0 ;
      RECT  175500.0 9600.0 198600.0 10500.0 ;
      RECT  152550.0 23400.0 175500.0 24300.0 ;
      RECT  152550.0 192900.0 175500.0 193800.0 ;
      RECT  152550.0 94800.0 175500.0 95700.0 ;
      RECT  175500.0 199200.0 185700.0 213000.0 ;
      RECT  175500.0 226800.0 185700.0 213000.0 ;
      RECT  175500.0 226800.0 185700.0 240600.0 ;
      RECT  175500.0 254400.0 185700.0 240600.0 ;
      RECT  175500.0 254400.0 185700.0 268200.0 ;
      RECT  175500.0 282000.0 185700.0 268200.0 ;
      RECT  175500.0 282000.0 185700.0 295800.0 ;
      RECT  175500.0 309600.0 185700.0 295800.0 ;
      RECT  175500.0 309600.0 185700.0 323400.0 ;
      RECT  175500.0 337200.0 185700.0 323400.0 ;
      RECT  175500.0 337200.0 185700.0 351000.0 ;
      RECT  175500.0 364800.0 185700.0 351000.0 ;
      RECT  175500.0 364800.0 185700.0 378600.0 ;
      RECT  175500.0 392400.0 185700.0 378600.0 ;
      RECT  175500.0 392400.0 185700.0 406200.0 ;
      RECT  175500.0 420000.0 185700.0 406200.0 ;
      RECT  185700.0 199200.0 195900.0 213000.0 ;
      RECT  185700.0 226800.0 195900.0 213000.0 ;
      RECT  185700.0 226800.0 195900.0 240600.0 ;
      RECT  185700.0 254400.0 195900.0 240600.0 ;
      RECT  185700.0 254400.0 195900.0 268200.0 ;
      RECT  185700.0 282000.0 195900.0 268200.0 ;
      RECT  185700.0 282000.0 195900.0 295800.0 ;
      RECT  185700.0 309600.0 195900.0 295800.0 ;
      RECT  185700.0 309600.0 195900.0 323400.0 ;
      RECT  185700.0 337200.0 195900.0 323400.0 ;
      RECT  185700.0 337200.0 195900.0 351000.0 ;
      RECT  185700.0 364800.0 195900.0 351000.0 ;
      RECT  185700.0 364800.0 195900.0 378600.0 ;
      RECT  185700.0 392400.0 195900.0 378600.0 ;
      RECT  185700.0 392400.0 195900.0 406200.0 ;
      RECT  185700.0 420000.0 195900.0 406200.0 ;
      RECT  174900.0 200700.0 196500.0 201900.0 ;
      RECT  174900.0 224100.0 196500.0 225300.0 ;
      RECT  174900.0 228300.0 196500.0 229500.0 ;
      RECT  174900.0 251700.0 196500.0 252900.0 ;
      RECT  174900.0 255900.0 196500.0 257100.0 ;
      RECT  174900.0 279300.0 196500.0 280500.0 ;
      RECT  174900.0 283500.0 196500.0 284700.0 ;
      RECT  174900.0 306900.0 196500.0 308100.0 ;
      RECT  174900.0 311100.0 196500.0 312300.0 ;
      RECT  174900.0 334500.0 196500.0 335700.0 ;
      RECT  174900.0 338700.0 196500.0 339900.0 ;
      RECT  174900.0 362100.0 196500.0 363300.0 ;
      RECT  174900.0 366300.0 196500.0 367500.0 ;
      RECT  174900.0 389700.0 196500.0 390900.0 ;
      RECT  174900.0 393900.0 196500.0 395100.0 ;
      RECT  174900.0 417300.0 196500.0 418500.0 ;
      RECT  174900.0 212400.0 196500.0 213300.0 ;
      RECT  174900.0 240000.0 196500.0 240900.0 ;
      RECT  174900.0 267600.0 196500.0 268500.0 ;
      RECT  174900.0 295200.0 196500.0 296100.0 ;
      RECT  174900.0 322800.0 196500.0 323700.0 ;
      RECT  174900.0 350400.0 196500.0 351300.0 ;
      RECT  174900.0 378000.0 196500.0 378900.0 ;
      RECT  174900.0 405600.0 196500.0 406500.0 ;
      RECT  180900.0 429600.0 182100.0 436800.0 ;
      RECT  178500.0 422400.0 179700.0 423600.0 ;
      RECT  180900.0 422400.0 182100.0 423600.0 ;
      RECT  180900.0 422400.0 182100.0 423600.0 ;
      RECT  178500.0 422400.0 179700.0 423600.0 ;
      RECT  178500.0 429600.0 179700.0 430800.0 ;
      RECT  180900.0 429600.0 182100.0 430800.0 ;
      RECT  180900.0 429600.0 182100.0 430800.0 ;
      RECT  178500.0 429600.0 179700.0 430800.0 ;
      RECT  180900.0 429600.0 182100.0 430800.0 ;
      RECT  183300.0 429600.0 184500.0 430800.0 ;
      RECT  183300.0 429600.0 184500.0 430800.0 ;
      RECT  180900.0 429600.0 182100.0 430800.0 ;
      RECT  180600.0 424650.0 179400.0 425850.0 ;
      RECT  180900.0 435000.0 182100.0 436200.0 ;
      RECT  178500.0 422400.0 179700.0 423600.0 ;
      RECT  180900.0 422400.0 182100.0 423600.0 ;
      RECT  178500.0 429600.0 179700.0 430800.0 ;
      RECT  183300.0 429600.0 184500.0 430800.0 ;
      RECT  175500.0 424800.0 185700.0 425700.0 ;
      RECT  175500.0 435900.0 185700.0 436800.0 ;
      RECT  191100.0 429600.0 192300.0 436800.0 ;
      RECT  188700.0 422400.0 189900.0 423600.0 ;
      RECT  191100.0 422400.0 192300.0 423600.0 ;
      RECT  191100.0 422400.0 192300.0 423600.0 ;
      RECT  188700.0 422400.0 189900.0 423600.0 ;
      RECT  188700.0 429600.0 189900.0 430800.0 ;
      RECT  191100.0 429600.0 192300.0 430800.0 ;
      RECT  191100.0 429600.0 192300.0 430800.0 ;
      RECT  188700.0 429600.0 189900.0 430800.0 ;
      RECT  191100.0 429600.0 192300.0 430800.0 ;
      RECT  193500.0 429600.0 194700.0 430800.0 ;
      RECT  193500.0 429600.0 194700.0 430800.0 ;
      RECT  191100.0 429600.0 192300.0 430800.0 ;
      RECT  190800.0 424650.0 189600.0 425850.0 ;
      RECT  191100.0 435000.0 192300.0 436200.0 ;
      RECT  188700.0 422400.0 189900.0 423600.0 ;
      RECT  191100.0 422400.0 192300.0 423600.0 ;
      RECT  188700.0 429600.0 189900.0 430800.0 ;
      RECT  193500.0 429600.0 194700.0 430800.0 ;
      RECT  185700.0 424800.0 195900.0 425700.0 ;
      RECT  185700.0 435900.0 195900.0 436800.0 ;
      RECT  175500.0 424800.0 195900.0 425700.0 ;
      RECT  175500.0 435900.0 195900.0 436800.0 ;
      RECT  175500.0 150300.0 185700.0 199200.0 ;
      RECT  185700.0 150300.0 195900.0 199200.0 ;
      RECT  175500.0 195000.0 195900.0 195900.0 ;
      RECT  175500.0 167700.0 195900.0 168600.0 ;
      RECT  175500.0 192900.0 195900.0 193800.0 ;
      RECT  175500.0 90000.0 185700.0 150300.0 ;
      RECT  185700.0 90000.0 195900.0 150300.0 ;
      RECT  175500.0 96900.0 195900.0 97800.0 ;
      RECT  175500.0 99000.0 195900.0 99900.0 ;
      RECT  175500.0 94800.0 195900.0 95700.0 ;
      RECT  175500.0 30000.0 185700.0 90000.0 ;
      RECT  195900.0 30000.0 185700.0 90000.0 ;
      RECT  175500.0 32400.0 195900.0 33300.0 ;
      RECT  175500.0 86400.0 195900.0 87300.0 ;
      RECT  175500.0 30000.0 185700.0 8100.0 ;
      RECT  185700.0 30000.0 195900.0 8100.0 ;
      RECT  175500.0 26400.0 195900.0 25500.0 ;
      RECT  175500.0 28800.0 195900.0 27900.0 ;
      RECT  175500.0 10500.0 195900.0 9600.0 ;
      RECT  175500.0 24300.0 195900.0 23400.0 ;
      RECT  87750.0 206550.0 88650.0 207450.0 ;
      RECT  87750.0 205350.0 88650.0 206250.0 ;
      RECT  83700.0 206550.0 88200.0 207450.0 ;
      RECT  87750.0 205800.0 88650.0 207000.0 ;
      RECT  88200.0 205350.0 92700.0 206250.0 ;
      RECT  87750.0 218550.0 88650.0 219450.0 ;
      RECT  87750.0 219750.0 88650.0 220650.0 ;
      RECT  83700.0 218550.0 88200.0 219450.0 ;
      RECT  87750.0 219000.0 88650.0 220200.0 ;
      RECT  88200.0 219750.0 92700.0 220650.0 ;
      RECT  87750.0 234150.0 88650.0 235050.0 ;
      RECT  87750.0 232950.0 88650.0 233850.0 ;
      RECT  83700.0 234150.0 88200.0 235050.0 ;
      RECT  87750.0 233400.0 88650.0 234600.0 ;
      RECT  88200.0 232950.0 92700.0 233850.0 ;
      RECT  87750.0 246150.0 88650.0 247050.0 ;
      RECT  87750.0 247350.0 88650.0 248250.0 ;
      RECT  83700.0 246150.0 88200.0 247050.0 ;
      RECT  87750.0 246600.0 88650.0 247800.0 ;
      RECT  88200.0 247350.0 92700.0 248250.0 ;
      RECT  87750.0 261750.0 88650.0 262650.0 ;
      RECT  87750.0 260550.0 88650.0 261450.0 ;
      RECT  83700.0 261750.0 88200.0 262650.0 ;
      RECT  87750.0 261000.0 88650.0 262200.0 ;
      RECT  88200.0 260550.0 92700.0 261450.0 ;
      RECT  87750.0 273750.0 88650.0 274650.0 ;
      RECT  87750.0 274950.0 88650.0 275850.0 ;
      RECT  83700.0 273750.0 88200.0 274650.0 ;
      RECT  87750.0 274200.0 88650.0 275400.0 ;
      RECT  88200.0 274950.0 92700.0 275850.0 ;
      RECT  87750.0 289350.0 88650.0 290250.0 ;
      RECT  87750.0 288150.0 88650.0 289050.0 ;
      RECT  83700.0 289350.0 88200.0 290250.0 ;
      RECT  87750.0 288600.0 88650.0 289800.0 ;
      RECT  88200.0 288150.0 92700.0 289050.0 ;
      RECT  87750.0 301350.0 88650.0 302250.0 ;
      RECT  87750.0 302550.0 88650.0 303450.0 ;
      RECT  83700.0 301350.0 88200.0 302250.0 ;
      RECT  87750.0 301800.0 88650.0 303000.0 ;
      RECT  88200.0 302550.0 92700.0 303450.0 ;
      RECT  87750.0 316950.0 88650.0 317850.0 ;
      RECT  87750.0 315750.0 88650.0 316650.0 ;
      RECT  83700.0 316950.0 88200.0 317850.0 ;
      RECT  87750.0 316200.0 88650.0 317400.0 ;
      RECT  88200.0 315750.0 92700.0 316650.0 ;
      RECT  87750.0 328950.0 88650.0 329850.0 ;
      RECT  87750.0 330150.0 88650.0 331050.0 ;
      RECT  83700.0 328950.0 88200.0 329850.0 ;
      RECT  87750.0 329400.0 88650.0 330600.0 ;
      RECT  88200.0 330150.0 92700.0 331050.0 ;
      RECT  87750.0 344550.0 88650.0 345450.0 ;
      RECT  87750.0 343350.0 88650.0 344250.0 ;
      RECT  83700.0 344550.0 88200.0 345450.0 ;
      RECT  87750.0 343800.0 88650.0 345000.0 ;
      RECT  88200.0 343350.0 92700.0 344250.0 ;
      RECT  87750.0 356550.0 88650.0 357450.0 ;
      RECT  87750.0 357750.0 88650.0 358650.0 ;
      RECT  83700.0 356550.0 88200.0 357450.0 ;
      RECT  87750.0 357000.0 88650.0 358200.0 ;
      RECT  88200.0 357750.0 92700.0 358650.0 ;
      RECT  87750.0 372150.0 88650.0 373050.0 ;
      RECT  87750.0 370950.0 88650.0 371850.0 ;
      RECT  83700.0 372150.0 88200.0 373050.0 ;
      RECT  87750.0 371400.0 88650.0 372600.0 ;
      RECT  88200.0 370950.0 92700.0 371850.0 ;
      RECT  87750.0 384150.0 88650.0 385050.0 ;
      RECT  87750.0 385350.0 88650.0 386250.0 ;
      RECT  83700.0 384150.0 88200.0 385050.0 ;
      RECT  87750.0 384600.0 88650.0 385800.0 ;
      RECT  88200.0 385350.0 92700.0 386250.0 ;
      RECT  87750.0 399750.0 88650.0 400650.0 ;
      RECT  87750.0 398550.0 88650.0 399450.0 ;
      RECT  83700.0 399750.0 88200.0 400650.0 ;
      RECT  87750.0 399000.0 88650.0 400200.0 ;
      RECT  88200.0 398550.0 92700.0 399450.0 ;
      RECT  87750.0 411750.0 88650.0 412650.0 ;
      RECT  87750.0 412950.0 88650.0 413850.0 ;
      RECT  83700.0 411750.0 88200.0 412650.0 ;
      RECT  87750.0 412200.0 88650.0 413400.0 ;
      RECT  88200.0 412950.0 92700.0 413850.0 ;
      RECT  59550.0 94950.0 75900.0 95850.0 ;
      RECT  61650.0 109350.0 75900.0 110250.0 ;
      RECT  63750.0 122550.0 75900.0 123450.0 ;
      RECT  65850.0 136950.0 75900.0 137850.0 ;
      RECT  67950.0 150150.0 75900.0 151050.0 ;
      RECT  70050.0 164550.0 75900.0 165450.0 ;
      RECT  72150.0 177750.0 75900.0 178650.0 ;
      RECT  74250.0 192150.0 75900.0 193050.0 ;
      RECT  59550.0 206550.0 78300.0 207450.0 ;
      RECT  67950.0 203850.0 81300.0 204750.0 ;
      RECT  59550.0 218550.0 78300.0 219450.0 ;
      RECT  70050.0 221250.0 81300.0 222150.0 ;
      RECT  59550.0 234150.0 78300.0 235050.0 ;
      RECT  72150.0 231450.0 81300.0 232350.0 ;
      RECT  59550.0 246150.0 78300.0 247050.0 ;
      RECT  74250.0 248850.0 81300.0 249750.0 ;
      RECT  61650.0 261750.0 78300.0 262650.0 ;
      RECT  67950.0 259050.0 81300.0 259950.0 ;
      RECT  61650.0 273750.0 78300.0 274650.0 ;
      RECT  70050.0 276450.0 81300.0 277350.0 ;
      RECT  61650.0 289350.0 78300.0 290250.0 ;
      RECT  72150.0 286650.0 81300.0 287550.0 ;
      RECT  61650.0 301350.0 78300.0 302250.0 ;
      RECT  74250.0 304050.0 81300.0 304950.0 ;
      RECT  63750.0 316950.0 78300.0 317850.0 ;
      RECT  67950.0 314250.0 81300.0 315150.0 ;
      RECT  63750.0 328950.0 78300.0 329850.0 ;
      RECT  70050.0 331650.0 81300.0 332550.0 ;
      RECT  63750.0 344550.0 78300.0 345450.0 ;
      RECT  72150.0 341850.0 81300.0 342750.0 ;
      RECT  63750.0 356550.0 78300.0 357450.0 ;
      RECT  74250.0 359250.0 81300.0 360150.0 ;
      RECT  65850.0 372150.0 78300.0 373050.0 ;
      RECT  67950.0 369450.0 81300.0 370350.0 ;
      RECT  65850.0 384150.0 78300.0 385050.0 ;
      RECT  70050.0 386850.0 81300.0 387750.0 ;
      RECT  65850.0 399750.0 78300.0 400650.0 ;
      RECT  72150.0 397050.0 81300.0 397950.0 ;
      RECT  65850.0 411750.0 78300.0 412650.0 ;
      RECT  74250.0 414450.0 81300.0 415350.0 ;
      RECT  114450.0 94950.0 113550.0 95850.0 ;
      RECT  114450.0 99450.0 113550.0 100350.0 ;
      RECT  118650.0 94950.0 114000.0 95850.0 ;
      RECT  114450.0 95400.0 113550.0 99900.0 ;
      RECT  114000.0 99450.0 111450.0 100350.0 ;
      RECT  130050.0 94950.0 122100.0 95850.0 ;
      RECT  114450.0 109350.0 113550.0 110250.0 ;
      RECT  114450.0 113250.0 113550.0 114150.0 ;
      RECT  118650.0 109350.0 114000.0 110250.0 ;
      RECT  114450.0 109800.0 113550.0 113700.0 ;
      RECT  114000.0 113250.0 108450.0 114150.0 ;
      RECT  127050.0 109350.0 122100.0 110250.0 ;
      RECT  130050.0 118050.0 105450.0 118950.0 ;
      RECT  127050.0 131850.0 102450.0 132750.0 ;
      RECT  111450.0 93450.0 94500.0 94350.0 ;
      RECT  108450.0 96150.0 97500.0 97050.0 ;
      RECT  105450.0 110850.0 94500.0 111750.0 ;
      RECT  108450.0 108150.0 97500.0 109050.0 ;
      RECT  111450.0 121050.0 94500.0 121950.0 ;
      RECT  102450.0 123750.0 97500.0 124650.0 ;
      RECT  105450.0 138450.0 94500.0 139350.0 ;
      RECT  102450.0 135750.0 97500.0 136650.0 ;
      RECT  88050.0 96150.0 87150.0 97050.0 ;
      RECT  88050.0 94950.0 87150.0 95850.0 ;
      RECT  92100.0 96150.0 87600.0 97050.0 ;
      RECT  88050.0 95400.0 87150.0 96600.0 ;
      RECT  87600.0 94950.0 83100.0 95850.0 ;
      RECT  88050.0 108150.0 87150.0 109050.0 ;
      RECT  88050.0 109350.0 87150.0 110250.0 ;
      RECT  92100.0 108150.0 87600.0 109050.0 ;
      RECT  88050.0 108600.0 87150.0 109800.0 ;
      RECT  87600.0 109350.0 83100.0 110250.0 ;
      RECT  88050.0 123750.0 87150.0 124650.0 ;
      RECT  88050.0 122550.0 87150.0 123450.0 ;
      RECT  92100.0 123750.0 87600.0 124650.0 ;
      RECT  88050.0 123000.0 87150.0 124200.0 ;
      RECT  87600.0 122550.0 83100.0 123450.0 ;
      RECT  88050.0 135750.0 87150.0 136650.0 ;
      RECT  88050.0 136950.0 87150.0 137850.0 ;
      RECT  92100.0 135750.0 87600.0 136650.0 ;
      RECT  88050.0 136200.0 87150.0 137400.0 ;
      RECT  87600.0 136950.0 83100.0 137850.0 ;
      RECT  117900.0 100650.0 116700.0 102600.0 ;
      RECT  117900.0 88800.0 116700.0 90750.0 ;
      RECT  122700.0 90150.0 121500.0 88350.0 ;
      RECT  122700.0 99450.0 121500.0 103050.0 ;
      RECT  120000.0 90150.0 119100.0 99450.0 ;
      RECT  122700.0 99450.0 121500.0 100650.0 ;
      RECT  120300.0 99450.0 119100.0 100650.0 ;
      RECT  120300.0 99450.0 119100.0 100650.0 ;
      RECT  122700.0 99450.0 121500.0 100650.0 ;
      RECT  122700.0 90150.0 121500.0 91350.0 ;
      RECT  120300.0 90150.0 119100.0 91350.0 ;
      RECT  120300.0 90150.0 119100.0 91350.0 ;
      RECT  122700.0 90150.0 121500.0 91350.0 ;
      RECT  117900.0 100050.0 116700.0 101250.0 ;
      RECT  117900.0 90150.0 116700.0 91350.0 ;
      RECT  122100.0 94800.0 120900.0 96000.0 ;
      RECT  122100.0 94800.0 120900.0 96000.0 ;
      RECT  119550.0 94950.0 118650.0 95850.0 ;
      RECT  124500.0 102150.0 114900.0 103050.0 ;
      RECT  124500.0 88350.0 114900.0 89250.0 ;
      RECT  117900.0 104550.0 116700.0 102600.0 ;
      RECT  117900.0 116400.0 116700.0 114450.0 ;
      RECT  122700.0 115050.0 121500.0 116850.0 ;
      RECT  122700.0 105750.0 121500.0 102150.0 ;
      RECT  120000.0 115050.0 119100.0 105750.0 ;
      RECT  122700.0 105750.0 121500.0 104550.0 ;
      RECT  120300.0 105750.0 119100.0 104550.0 ;
      RECT  120300.0 105750.0 119100.0 104550.0 ;
      RECT  122700.0 105750.0 121500.0 104550.0 ;
      RECT  122700.0 115050.0 121500.0 113850.0 ;
      RECT  120300.0 115050.0 119100.0 113850.0 ;
      RECT  120300.0 115050.0 119100.0 113850.0 ;
      RECT  122700.0 115050.0 121500.0 113850.0 ;
      RECT  117900.0 105150.0 116700.0 103950.0 ;
      RECT  117900.0 115050.0 116700.0 113850.0 ;
      RECT  122100.0 110400.0 120900.0 109200.0 ;
      RECT  122100.0 110400.0 120900.0 109200.0 ;
      RECT  119550.0 110250.0 118650.0 109350.0 ;
      RECT  124500.0 103050.0 114900.0 102150.0 ;
      RECT  124500.0 116850.0 114900.0 115950.0 ;
      RECT  78900.0 100650.0 77700.0 102600.0 ;
      RECT  78900.0 88800.0 77700.0 90750.0 ;
      RECT  83700.0 90150.0 82500.0 88350.0 ;
      RECT  83700.0 99450.0 82500.0 103050.0 ;
      RECT  81000.0 90150.0 80100.0 99450.0 ;
      RECT  83700.0 99450.0 82500.0 100650.0 ;
      RECT  81300.0 99450.0 80100.0 100650.0 ;
      RECT  81300.0 99450.0 80100.0 100650.0 ;
      RECT  83700.0 99450.0 82500.0 100650.0 ;
      RECT  83700.0 90150.0 82500.0 91350.0 ;
      RECT  81300.0 90150.0 80100.0 91350.0 ;
      RECT  81300.0 90150.0 80100.0 91350.0 ;
      RECT  83700.0 90150.0 82500.0 91350.0 ;
      RECT  78900.0 100050.0 77700.0 101250.0 ;
      RECT  78900.0 90150.0 77700.0 91350.0 ;
      RECT  83100.0 94800.0 81900.0 96000.0 ;
      RECT  83100.0 94800.0 81900.0 96000.0 ;
      RECT  80550.0 94950.0 79650.0 95850.0 ;
      RECT  85500.0 102150.0 75900.0 103050.0 ;
      RECT  85500.0 88350.0 75900.0 89250.0 ;
      RECT  78900.0 104550.0 77700.0 102600.0 ;
      RECT  78900.0 116400.0 77700.0 114450.0 ;
      RECT  83700.0 115050.0 82500.0 116850.0 ;
      RECT  83700.0 105750.0 82500.0 102150.0 ;
      RECT  81000.0 115050.0 80100.0 105750.0 ;
      RECT  83700.0 105750.0 82500.0 104550.0 ;
      RECT  81300.0 105750.0 80100.0 104550.0 ;
      RECT  81300.0 105750.0 80100.0 104550.0 ;
      RECT  83700.0 105750.0 82500.0 104550.0 ;
      RECT  83700.0 115050.0 82500.0 113850.0 ;
      RECT  81300.0 115050.0 80100.0 113850.0 ;
      RECT  81300.0 115050.0 80100.0 113850.0 ;
      RECT  83700.0 115050.0 82500.0 113850.0 ;
      RECT  78900.0 105150.0 77700.0 103950.0 ;
      RECT  78900.0 115050.0 77700.0 113850.0 ;
      RECT  83100.0 110400.0 81900.0 109200.0 ;
      RECT  83100.0 110400.0 81900.0 109200.0 ;
      RECT  80550.0 110250.0 79650.0 109350.0 ;
      RECT  85500.0 103050.0 75900.0 102150.0 ;
      RECT  85500.0 116850.0 75900.0 115950.0 ;
      RECT  78900.0 128250.0 77700.0 130200.0 ;
      RECT  78900.0 116400.0 77700.0 118350.0 ;
      RECT  83700.0 117750.0 82500.0 115950.0 ;
      RECT  83700.0 127050.0 82500.0 130650.0 ;
      RECT  81000.0 117750.0 80100.0 127050.0 ;
      RECT  83700.0 127050.0 82500.0 128250.0 ;
      RECT  81300.0 127050.0 80100.0 128250.0 ;
      RECT  81300.0 127050.0 80100.0 128250.0 ;
      RECT  83700.0 127050.0 82500.0 128250.0 ;
      RECT  83700.0 117750.0 82500.0 118950.0 ;
      RECT  81300.0 117750.0 80100.0 118950.0 ;
      RECT  81300.0 117750.0 80100.0 118950.0 ;
      RECT  83700.0 117750.0 82500.0 118950.0 ;
      RECT  78900.0 127650.0 77700.0 128850.0 ;
      RECT  78900.0 117750.0 77700.0 118950.0 ;
      RECT  83100.0 122400.0 81900.0 123600.0 ;
      RECT  83100.0 122400.0 81900.0 123600.0 ;
      RECT  80550.0 122550.0 79650.0 123450.0 ;
      RECT  85500.0 129750.0 75900.0 130650.0 ;
      RECT  85500.0 115950.0 75900.0 116850.0 ;
      RECT  78900.0 132150.0 77700.0 130200.0 ;
      RECT  78900.0 144000.0 77700.0 142050.0 ;
      RECT  83700.0 142650.0 82500.0 144450.0 ;
      RECT  83700.0 133350.0 82500.0 129750.0 ;
      RECT  81000.0 142650.0 80100.0 133350.0 ;
      RECT  83700.0 133350.0 82500.0 132150.0 ;
      RECT  81300.0 133350.0 80100.0 132150.0 ;
      RECT  81300.0 133350.0 80100.0 132150.0 ;
      RECT  83700.0 133350.0 82500.0 132150.0 ;
      RECT  83700.0 142650.0 82500.0 141450.0 ;
      RECT  81300.0 142650.0 80100.0 141450.0 ;
      RECT  81300.0 142650.0 80100.0 141450.0 ;
      RECT  83700.0 142650.0 82500.0 141450.0 ;
      RECT  78900.0 132750.0 77700.0 131550.0 ;
      RECT  78900.0 142650.0 77700.0 141450.0 ;
      RECT  83100.0 138000.0 81900.0 136800.0 ;
      RECT  83100.0 138000.0 81900.0 136800.0 ;
      RECT  80550.0 137850.0 79650.0 136950.0 ;
      RECT  85500.0 130650.0 75900.0 129750.0 ;
      RECT  85500.0 144450.0 75900.0 143550.0 ;
      RECT  98100.0 90750.0 96900.0 88350.0 ;
      RECT  98100.0 99450.0 96900.0 103050.0 ;
      RECT  93300.0 99450.0 92100.0 103050.0 ;
      RECT  90900.0 100650.0 89700.0 102600.0 ;
      RECT  90900.0 88800.0 89700.0 90750.0 ;
      RECT  98100.0 99450.0 96900.0 100650.0 ;
      RECT  95700.0 99450.0 94500.0 100650.0 ;
      RECT  95700.0 99450.0 94500.0 100650.0 ;
      RECT  98100.0 99450.0 96900.0 100650.0 ;
      RECT  95700.0 99450.0 94500.0 100650.0 ;
      RECT  93300.0 99450.0 92100.0 100650.0 ;
      RECT  93300.0 99450.0 92100.0 100650.0 ;
      RECT  95700.0 99450.0 94500.0 100650.0 ;
      RECT  98100.0 90750.0 96900.0 91950.0 ;
      RECT  95700.0 90750.0 94500.0 91950.0 ;
      RECT  95700.0 90750.0 94500.0 91950.0 ;
      RECT  98100.0 90750.0 96900.0 91950.0 ;
      RECT  95700.0 90750.0 94500.0 91950.0 ;
      RECT  93300.0 90750.0 92100.0 91950.0 ;
      RECT  93300.0 90750.0 92100.0 91950.0 ;
      RECT  95700.0 90750.0 94500.0 91950.0 ;
      RECT  90900.0 100050.0 89700.0 101250.0 ;
      RECT  90900.0 90150.0 89700.0 91350.0 ;
      RECT  93300.0 93300.0 94500.0 94500.0 ;
      RECT  96300.0 96000.0 97500.0 97200.0 ;
      RECT  95700.0 99450.0 94500.0 100650.0 ;
      RECT  93300.0 90750.0 92100.0 91950.0 ;
      RECT  92100.0 96000.0 93300.0 97200.0 ;
      RECT  97500.0 96000.0 96300.0 97200.0 ;
      RECT  94500.0 93300.0 93300.0 94500.0 ;
      RECT  93300.0 96000.0 92100.0 97200.0 ;
      RECT  99900.0 102150.0 85500.0 103050.0 ;
      RECT  99900.0 88350.0 85500.0 89250.0 ;
      RECT  98100.0 114450.0 96900.0 116850.0 ;
      RECT  98100.0 105750.0 96900.0 102150.0 ;
      RECT  93300.0 105750.0 92100.0 102150.0 ;
      RECT  90900.0 104550.0 89700.0 102600.0 ;
      RECT  90900.0 116400.0 89700.0 114450.0 ;
      RECT  98100.0 105750.0 96900.0 104550.0 ;
      RECT  95700.0 105750.0 94500.0 104550.0 ;
      RECT  95700.0 105750.0 94500.0 104550.0 ;
      RECT  98100.0 105750.0 96900.0 104550.0 ;
      RECT  95700.0 105750.0 94500.0 104550.0 ;
      RECT  93300.0 105750.0 92100.0 104550.0 ;
      RECT  93300.0 105750.0 92100.0 104550.0 ;
      RECT  95700.0 105750.0 94500.0 104550.0 ;
      RECT  98100.0 114450.0 96900.0 113250.0 ;
      RECT  95700.0 114450.0 94500.0 113250.0 ;
      RECT  95700.0 114450.0 94500.0 113250.0 ;
      RECT  98100.0 114450.0 96900.0 113250.0 ;
      RECT  95700.0 114450.0 94500.0 113250.0 ;
      RECT  93300.0 114450.0 92100.0 113250.0 ;
      RECT  93300.0 114450.0 92100.0 113250.0 ;
      RECT  95700.0 114450.0 94500.0 113250.0 ;
      RECT  90900.0 105150.0 89700.0 103950.0 ;
      RECT  90900.0 115050.0 89700.0 113850.0 ;
      RECT  93300.0 111900.0 94500.0 110700.0 ;
      RECT  96300.0 109200.0 97500.0 108000.0 ;
      RECT  95700.0 105750.0 94500.0 104550.0 ;
      RECT  93300.0 114450.0 92100.0 113250.0 ;
      RECT  92100.0 109200.0 93300.0 108000.0 ;
      RECT  97500.0 109200.0 96300.0 108000.0 ;
      RECT  94500.0 111900.0 93300.0 110700.0 ;
      RECT  93300.0 109200.0 92100.0 108000.0 ;
      RECT  99900.0 103050.0 85500.0 102150.0 ;
      RECT  99900.0 116850.0 85500.0 115950.0 ;
      RECT  98100.0 118350.0 96900.0 115950.0 ;
      RECT  98100.0 127050.0 96900.0 130650.0 ;
      RECT  93300.0 127050.0 92100.0 130650.0 ;
      RECT  90900.0 128250.0 89700.0 130200.0 ;
      RECT  90900.0 116400.0 89700.0 118350.0 ;
      RECT  98100.0 127050.0 96900.0 128250.0 ;
      RECT  95700.0 127050.0 94500.0 128250.0 ;
      RECT  95700.0 127050.0 94500.0 128250.0 ;
      RECT  98100.0 127050.0 96900.0 128250.0 ;
      RECT  95700.0 127050.0 94500.0 128250.0 ;
      RECT  93300.0 127050.0 92100.0 128250.0 ;
      RECT  93300.0 127050.0 92100.0 128250.0 ;
      RECT  95700.0 127050.0 94500.0 128250.0 ;
      RECT  98100.0 118350.0 96900.0 119550.0 ;
      RECT  95700.0 118350.0 94500.0 119550.0 ;
      RECT  95700.0 118350.0 94500.0 119550.0 ;
      RECT  98100.0 118350.0 96900.0 119550.0 ;
      RECT  95700.0 118350.0 94500.0 119550.0 ;
      RECT  93300.0 118350.0 92100.0 119550.0 ;
      RECT  93300.0 118350.0 92100.0 119550.0 ;
      RECT  95700.0 118350.0 94500.0 119550.0 ;
      RECT  90900.0 127650.0 89700.0 128850.0 ;
      RECT  90900.0 117750.0 89700.0 118950.0 ;
      RECT  93300.0 120900.0 94500.0 122100.0 ;
      RECT  96300.0 123600.0 97500.0 124800.0 ;
      RECT  95700.0 127050.0 94500.0 128250.0 ;
      RECT  93300.0 118350.0 92100.0 119550.0 ;
      RECT  92100.0 123600.0 93300.0 124800.0 ;
      RECT  97500.0 123600.0 96300.0 124800.0 ;
      RECT  94500.0 120900.0 93300.0 122100.0 ;
      RECT  93300.0 123600.0 92100.0 124800.0 ;
      RECT  99900.0 129750.0 85500.0 130650.0 ;
      RECT  99900.0 115950.0 85500.0 116850.0 ;
      RECT  98100.0 142050.0 96900.0 144450.0 ;
      RECT  98100.0 133350.0 96900.0 129750.0 ;
      RECT  93300.0 133350.0 92100.0 129750.0 ;
      RECT  90900.0 132150.0 89700.0 130200.0 ;
      RECT  90900.0 144000.0 89700.0 142050.0 ;
      RECT  98100.0 133350.0 96900.0 132150.0 ;
      RECT  95700.0 133350.0 94500.0 132150.0 ;
      RECT  95700.0 133350.0 94500.0 132150.0 ;
      RECT  98100.0 133350.0 96900.0 132150.0 ;
      RECT  95700.0 133350.0 94500.0 132150.0 ;
      RECT  93300.0 133350.0 92100.0 132150.0 ;
      RECT  93300.0 133350.0 92100.0 132150.0 ;
      RECT  95700.0 133350.0 94500.0 132150.0 ;
      RECT  98100.0 142050.0 96900.0 140850.0 ;
      RECT  95700.0 142050.0 94500.0 140850.0 ;
      RECT  95700.0 142050.0 94500.0 140850.0 ;
      RECT  98100.0 142050.0 96900.0 140850.0 ;
      RECT  95700.0 142050.0 94500.0 140850.0 ;
      RECT  93300.0 142050.0 92100.0 140850.0 ;
      RECT  93300.0 142050.0 92100.0 140850.0 ;
      RECT  95700.0 142050.0 94500.0 140850.0 ;
      RECT  90900.0 132750.0 89700.0 131550.0 ;
      RECT  90900.0 142650.0 89700.0 141450.0 ;
      RECT  93300.0 139500.0 94500.0 138300.0 ;
      RECT  96300.0 136800.0 97500.0 135600.0 ;
      RECT  95700.0 133350.0 94500.0 132150.0 ;
      RECT  93300.0 142050.0 92100.0 140850.0 ;
      RECT  92100.0 136800.0 93300.0 135600.0 ;
      RECT  97500.0 136800.0 96300.0 135600.0 ;
      RECT  94500.0 139500.0 93300.0 138300.0 ;
      RECT  93300.0 136800.0 92100.0 135600.0 ;
      RECT  99900.0 130650.0 85500.0 129750.0 ;
      RECT  99900.0 144450.0 85500.0 143550.0 ;
      RECT  110850.0 99300.0 112050.0 100500.0 ;
      RECT  129450.0 94800.0 130650.0 96000.0 ;
      RECT  107850.0 113100.0 109050.0 114300.0 ;
      RECT  126450.0 109200.0 127650.0 110400.0 ;
      RECT  129450.0 117900.0 130650.0 119100.0 ;
      RECT  104850.0 117900.0 106050.0 119100.0 ;
      RECT  126450.0 131700.0 127650.0 132900.0 ;
      RECT  101850.0 131700.0 103050.0 132900.0 ;
      RECT  110850.0 93300.0 112050.0 94500.0 ;
      RECT  107850.0 96000.0 109050.0 97200.0 ;
      RECT  104850.0 110700.0 106050.0 111900.0 ;
      RECT  107850.0 108000.0 109050.0 109200.0 ;
      RECT  110850.0 120900.0 112050.0 122100.0 ;
      RECT  101850.0 123600.0 103050.0 124800.0 ;
      RECT  104850.0 138300.0 106050.0 139500.0 ;
      RECT  101850.0 135600.0 103050.0 136800.0 ;
      RECT  79650.0 94950.0 75900.0 95850.0 ;
      RECT  79650.0 109350.0 75900.0 110250.0 ;
      RECT  79650.0 122550.0 75900.0 123450.0 ;
      RECT  79650.0 136950.0 75900.0 137850.0 ;
      RECT  130500.0 102150.0 75900.0 103050.0 ;
      RECT  130500.0 129750.0 75900.0 130650.0 ;
      RECT  130500.0 88350.0 75900.0 89250.0 ;
      RECT  130500.0 115950.0 75900.0 116850.0 ;
      RECT  130500.0 143550.0 75900.0 144450.0 ;
      RECT  114450.0 150150.0 113550.0 151050.0 ;
      RECT  114450.0 154650.0 113550.0 155550.0 ;
      RECT  118650.0 150150.0 114000.0 151050.0 ;
      RECT  114450.0 150600.0 113550.0 155100.0 ;
      RECT  114000.0 154650.0 111450.0 155550.0 ;
      RECT  130050.0 150150.0 122100.0 151050.0 ;
      RECT  114450.0 164550.0 113550.0 165450.0 ;
      RECT  114450.0 168450.0 113550.0 169350.0 ;
      RECT  118650.0 164550.0 114000.0 165450.0 ;
      RECT  114450.0 165000.0 113550.0 168900.0 ;
      RECT  114000.0 168450.0 108450.0 169350.0 ;
      RECT  127050.0 164550.0 122100.0 165450.0 ;
      RECT  130050.0 173250.0 105450.0 174150.0 ;
      RECT  127050.0 187050.0 102450.0 187950.0 ;
      RECT  111450.0 148650.0 94500.0 149550.0 ;
      RECT  108450.0 151350.0 97500.0 152250.0 ;
      RECT  105450.0 166050.0 94500.0 166950.0 ;
      RECT  108450.0 163350.0 97500.0 164250.0 ;
      RECT  111450.0 176250.0 94500.0 177150.0 ;
      RECT  102450.0 178950.0 97500.0 179850.0 ;
      RECT  105450.0 193650.0 94500.0 194550.0 ;
      RECT  102450.0 190950.0 97500.0 191850.0 ;
      RECT  88050.0 151350.0 87150.0 152250.0 ;
      RECT  88050.0 150150.0 87150.0 151050.0 ;
      RECT  92100.0 151350.0 87600.0 152250.0 ;
      RECT  88050.0 150600.0 87150.0 151800.0 ;
      RECT  87600.0 150150.0 83100.0 151050.0 ;
      RECT  88050.0 163350.0 87150.0 164250.0 ;
      RECT  88050.0 164550.0 87150.0 165450.0 ;
      RECT  92100.0 163350.0 87600.0 164250.0 ;
      RECT  88050.0 163800.0 87150.0 165000.0 ;
      RECT  87600.0 164550.0 83100.0 165450.0 ;
      RECT  88050.0 178950.0 87150.0 179850.0 ;
      RECT  88050.0 177750.0 87150.0 178650.0 ;
      RECT  92100.0 178950.0 87600.0 179850.0 ;
      RECT  88050.0 178200.0 87150.0 179400.0 ;
      RECT  87600.0 177750.0 83100.0 178650.0 ;
      RECT  88050.0 190950.0 87150.0 191850.0 ;
      RECT  88050.0 192150.0 87150.0 193050.0 ;
      RECT  92100.0 190950.0 87600.0 191850.0 ;
      RECT  88050.0 191400.0 87150.0 192600.0 ;
      RECT  87600.0 192150.0 83100.0 193050.0 ;
      RECT  117900.0 155850.0 116700.0 157800.0 ;
      RECT  117900.0 144000.0 116700.0 145950.0 ;
      RECT  122700.0 145350.0 121500.0 143550.0 ;
      RECT  122700.0 154650.0 121500.0 158250.0 ;
      RECT  120000.0 145350.0 119100.0 154650.0 ;
      RECT  122700.0 154650.0 121500.0 155850.0 ;
      RECT  120300.0 154650.0 119100.0 155850.0 ;
      RECT  120300.0 154650.0 119100.0 155850.0 ;
      RECT  122700.0 154650.0 121500.0 155850.0 ;
      RECT  122700.0 145350.0 121500.0 146550.0 ;
      RECT  120300.0 145350.0 119100.0 146550.0 ;
      RECT  120300.0 145350.0 119100.0 146550.0 ;
      RECT  122700.0 145350.0 121500.0 146550.0 ;
      RECT  117900.0 155250.0 116700.0 156450.0 ;
      RECT  117900.0 145350.0 116700.0 146550.0 ;
      RECT  122100.0 150000.0 120900.0 151200.0 ;
      RECT  122100.0 150000.0 120900.0 151200.0 ;
      RECT  119550.0 150150.0 118650.0 151050.0 ;
      RECT  124500.0 157350.0 114900.0 158250.0 ;
      RECT  124500.0 143550.0 114900.0 144450.0 ;
      RECT  117900.0 159750.0 116700.0 157800.0 ;
      RECT  117900.0 171600.0 116700.0 169650.0 ;
      RECT  122700.0 170250.0 121500.0 172050.0 ;
      RECT  122700.0 160950.0 121500.0 157350.0 ;
      RECT  120000.0 170250.0 119100.0 160950.0 ;
      RECT  122700.0 160950.0 121500.0 159750.0 ;
      RECT  120300.0 160950.0 119100.0 159750.0 ;
      RECT  120300.0 160950.0 119100.0 159750.0 ;
      RECT  122700.0 160950.0 121500.0 159750.0 ;
      RECT  122700.0 170250.0 121500.0 169050.0 ;
      RECT  120300.0 170250.0 119100.0 169050.0 ;
      RECT  120300.0 170250.0 119100.0 169050.0 ;
      RECT  122700.0 170250.0 121500.0 169050.0 ;
      RECT  117900.0 160350.0 116700.0 159150.0 ;
      RECT  117900.0 170250.0 116700.0 169050.0 ;
      RECT  122100.0 165600.0 120900.0 164400.0 ;
      RECT  122100.0 165600.0 120900.0 164400.0 ;
      RECT  119550.0 165450.0 118650.0 164550.0 ;
      RECT  124500.0 158250.0 114900.0 157350.0 ;
      RECT  124500.0 172050.0 114900.0 171150.0 ;
      RECT  78900.0 155850.0 77700.0 157800.0 ;
      RECT  78900.0 144000.0 77700.0 145950.0 ;
      RECT  83700.0 145350.0 82500.0 143550.0 ;
      RECT  83700.0 154650.0 82500.0 158250.0 ;
      RECT  81000.0 145350.0 80100.0 154650.0 ;
      RECT  83700.0 154650.0 82500.0 155850.0 ;
      RECT  81300.0 154650.0 80100.0 155850.0 ;
      RECT  81300.0 154650.0 80100.0 155850.0 ;
      RECT  83700.0 154650.0 82500.0 155850.0 ;
      RECT  83700.0 145350.0 82500.0 146550.0 ;
      RECT  81300.0 145350.0 80100.0 146550.0 ;
      RECT  81300.0 145350.0 80100.0 146550.0 ;
      RECT  83700.0 145350.0 82500.0 146550.0 ;
      RECT  78900.0 155250.0 77700.0 156450.0 ;
      RECT  78900.0 145350.0 77700.0 146550.0 ;
      RECT  83100.0 150000.0 81900.0 151200.0 ;
      RECT  83100.0 150000.0 81900.0 151200.0 ;
      RECT  80550.0 150150.0 79650.0 151050.0 ;
      RECT  85500.0 157350.0 75900.0 158250.0 ;
      RECT  85500.0 143550.0 75900.0 144450.0 ;
      RECT  78900.0 159750.0 77700.0 157800.0 ;
      RECT  78900.0 171600.0 77700.0 169650.0 ;
      RECT  83700.0 170250.0 82500.0 172050.0 ;
      RECT  83700.0 160950.0 82500.0 157350.0 ;
      RECT  81000.0 170250.0 80100.0 160950.0 ;
      RECT  83700.0 160950.0 82500.0 159750.0 ;
      RECT  81300.0 160950.0 80100.0 159750.0 ;
      RECT  81300.0 160950.0 80100.0 159750.0 ;
      RECT  83700.0 160950.0 82500.0 159750.0 ;
      RECT  83700.0 170250.0 82500.0 169050.0 ;
      RECT  81300.0 170250.0 80100.0 169050.0 ;
      RECT  81300.0 170250.0 80100.0 169050.0 ;
      RECT  83700.0 170250.0 82500.0 169050.0 ;
      RECT  78900.0 160350.0 77700.0 159150.0 ;
      RECT  78900.0 170250.0 77700.0 169050.0 ;
      RECT  83100.0 165600.0 81900.0 164400.0 ;
      RECT  83100.0 165600.0 81900.0 164400.0 ;
      RECT  80550.0 165450.0 79650.0 164550.0 ;
      RECT  85500.0 158250.0 75900.0 157350.0 ;
      RECT  85500.0 172050.0 75900.0 171150.0 ;
      RECT  78900.0 183450.0 77700.0 185400.0 ;
      RECT  78900.0 171600.0 77700.0 173550.0 ;
      RECT  83700.0 172950.0 82500.0 171150.0 ;
      RECT  83700.0 182250.0 82500.0 185850.0 ;
      RECT  81000.0 172950.0 80100.0 182250.0 ;
      RECT  83700.0 182250.0 82500.0 183450.0 ;
      RECT  81300.0 182250.0 80100.0 183450.0 ;
      RECT  81300.0 182250.0 80100.0 183450.0 ;
      RECT  83700.0 182250.0 82500.0 183450.0 ;
      RECT  83700.0 172950.0 82500.0 174150.0 ;
      RECT  81300.0 172950.0 80100.0 174150.0 ;
      RECT  81300.0 172950.0 80100.0 174150.0 ;
      RECT  83700.0 172950.0 82500.0 174150.0 ;
      RECT  78900.0 182850.0 77700.0 184050.0 ;
      RECT  78900.0 172950.0 77700.0 174150.0 ;
      RECT  83100.0 177600.0 81900.0 178800.0 ;
      RECT  83100.0 177600.0 81900.0 178800.0 ;
      RECT  80550.0 177750.0 79650.0 178650.0 ;
      RECT  85500.0 184950.0 75900.0 185850.0 ;
      RECT  85500.0 171150.0 75900.0 172050.0 ;
      RECT  78900.0 187350.0 77700.0 185400.0 ;
      RECT  78900.0 199200.0 77700.0 197250.0 ;
      RECT  83700.0 197850.0 82500.0 199650.0 ;
      RECT  83700.0 188550.0 82500.0 184950.0 ;
      RECT  81000.0 197850.0 80100.0 188550.0 ;
      RECT  83700.0 188550.0 82500.0 187350.0 ;
      RECT  81300.0 188550.0 80100.0 187350.0 ;
      RECT  81300.0 188550.0 80100.0 187350.0 ;
      RECT  83700.0 188550.0 82500.0 187350.0 ;
      RECT  83700.0 197850.0 82500.0 196650.0 ;
      RECT  81300.0 197850.0 80100.0 196650.0 ;
      RECT  81300.0 197850.0 80100.0 196650.0 ;
      RECT  83700.0 197850.0 82500.0 196650.0 ;
      RECT  78900.0 187950.0 77700.0 186750.0 ;
      RECT  78900.0 197850.0 77700.0 196650.0 ;
      RECT  83100.0 193200.0 81900.0 192000.0 ;
      RECT  83100.0 193200.0 81900.0 192000.0 ;
      RECT  80550.0 193050.0 79650.0 192150.0 ;
      RECT  85500.0 185850.0 75900.0 184950.0 ;
      RECT  85500.0 199650.0 75900.0 198750.0 ;
      RECT  98100.0 145950.0 96900.0 143550.0 ;
      RECT  98100.0 154650.0 96900.0 158250.0 ;
      RECT  93300.0 154650.0 92100.0 158250.0 ;
      RECT  90900.0 155850.0 89700.0 157800.0 ;
      RECT  90900.0 144000.0 89700.0 145950.0 ;
      RECT  98100.0 154650.0 96900.0 155850.0 ;
      RECT  95700.0 154650.0 94500.0 155850.0 ;
      RECT  95700.0 154650.0 94500.0 155850.0 ;
      RECT  98100.0 154650.0 96900.0 155850.0 ;
      RECT  95700.0 154650.0 94500.0 155850.0 ;
      RECT  93300.0 154650.0 92100.0 155850.0 ;
      RECT  93300.0 154650.0 92100.0 155850.0 ;
      RECT  95700.0 154650.0 94500.0 155850.0 ;
      RECT  98100.0 145950.0 96900.0 147150.0 ;
      RECT  95700.0 145950.0 94500.0 147150.0 ;
      RECT  95700.0 145950.0 94500.0 147150.0 ;
      RECT  98100.0 145950.0 96900.0 147150.0 ;
      RECT  95700.0 145950.0 94500.0 147150.0 ;
      RECT  93300.0 145950.0 92100.0 147150.0 ;
      RECT  93300.0 145950.0 92100.0 147150.0 ;
      RECT  95700.0 145950.0 94500.0 147150.0 ;
      RECT  90900.0 155250.0 89700.0 156450.0 ;
      RECT  90900.0 145350.0 89700.0 146550.0 ;
      RECT  93300.0 148500.0 94500.0 149700.0 ;
      RECT  96300.0 151200.0 97500.0 152400.0 ;
      RECT  95700.0 154650.0 94500.0 155850.0 ;
      RECT  93300.0 145950.0 92100.0 147150.0 ;
      RECT  92100.0 151200.0 93300.0 152400.0 ;
      RECT  97500.0 151200.0 96300.0 152400.0 ;
      RECT  94500.0 148500.0 93300.0 149700.0 ;
      RECT  93300.0 151200.0 92100.0 152400.0 ;
      RECT  99900.0 157350.0 85500.0 158250.0 ;
      RECT  99900.0 143550.0 85500.0 144450.0 ;
      RECT  98100.0 169650.0 96900.0 172050.0 ;
      RECT  98100.0 160950.0 96900.0 157350.0 ;
      RECT  93300.0 160950.0 92100.0 157350.0 ;
      RECT  90900.0 159750.0 89700.0 157800.0 ;
      RECT  90900.0 171600.0 89700.0 169650.0 ;
      RECT  98100.0 160950.0 96900.0 159750.0 ;
      RECT  95700.0 160950.0 94500.0 159750.0 ;
      RECT  95700.0 160950.0 94500.0 159750.0 ;
      RECT  98100.0 160950.0 96900.0 159750.0 ;
      RECT  95700.0 160950.0 94500.0 159750.0 ;
      RECT  93300.0 160950.0 92100.0 159750.0 ;
      RECT  93300.0 160950.0 92100.0 159750.0 ;
      RECT  95700.0 160950.0 94500.0 159750.0 ;
      RECT  98100.0 169650.0 96900.0 168450.0 ;
      RECT  95700.0 169650.0 94500.0 168450.0 ;
      RECT  95700.0 169650.0 94500.0 168450.0 ;
      RECT  98100.0 169650.0 96900.0 168450.0 ;
      RECT  95700.0 169650.0 94500.0 168450.0 ;
      RECT  93300.0 169650.0 92100.0 168450.0 ;
      RECT  93300.0 169650.0 92100.0 168450.0 ;
      RECT  95700.0 169650.0 94500.0 168450.0 ;
      RECT  90900.0 160350.0 89700.0 159150.0 ;
      RECT  90900.0 170250.0 89700.0 169050.0 ;
      RECT  93300.0 167100.0 94500.0 165900.0 ;
      RECT  96300.0 164400.0 97500.0 163200.0 ;
      RECT  95700.0 160950.0 94500.0 159750.0 ;
      RECT  93300.0 169650.0 92100.0 168450.0 ;
      RECT  92100.0 164400.0 93300.0 163200.0 ;
      RECT  97500.0 164400.0 96300.0 163200.0 ;
      RECT  94500.0 167100.0 93300.0 165900.0 ;
      RECT  93300.0 164400.0 92100.0 163200.0 ;
      RECT  99900.0 158250.0 85500.0 157350.0 ;
      RECT  99900.0 172050.0 85500.0 171150.0 ;
      RECT  98100.0 173550.0 96900.0 171150.0 ;
      RECT  98100.0 182250.0 96900.0 185850.0 ;
      RECT  93300.0 182250.0 92100.0 185850.0 ;
      RECT  90900.0 183450.0 89700.0 185400.0 ;
      RECT  90900.0 171600.0 89700.0 173550.0 ;
      RECT  98100.0 182250.0 96900.0 183450.0 ;
      RECT  95700.0 182250.0 94500.0 183450.0 ;
      RECT  95700.0 182250.0 94500.0 183450.0 ;
      RECT  98100.0 182250.0 96900.0 183450.0 ;
      RECT  95700.0 182250.0 94500.0 183450.0 ;
      RECT  93300.0 182250.0 92100.0 183450.0 ;
      RECT  93300.0 182250.0 92100.0 183450.0 ;
      RECT  95700.0 182250.0 94500.0 183450.0 ;
      RECT  98100.0 173550.0 96900.0 174750.0 ;
      RECT  95700.0 173550.0 94500.0 174750.0 ;
      RECT  95700.0 173550.0 94500.0 174750.0 ;
      RECT  98100.0 173550.0 96900.0 174750.0 ;
      RECT  95700.0 173550.0 94500.0 174750.0 ;
      RECT  93300.0 173550.0 92100.0 174750.0 ;
      RECT  93300.0 173550.0 92100.0 174750.0 ;
      RECT  95700.0 173550.0 94500.0 174750.0 ;
      RECT  90900.0 182850.0 89700.0 184050.0 ;
      RECT  90900.0 172950.0 89700.0 174150.0 ;
      RECT  93300.0 176100.0 94500.0 177300.0 ;
      RECT  96300.0 178800.0 97500.0 180000.0 ;
      RECT  95700.0 182250.0 94500.0 183450.0 ;
      RECT  93300.0 173550.0 92100.0 174750.0 ;
      RECT  92100.0 178800.0 93300.0 180000.0 ;
      RECT  97500.0 178800.0 96300.0 180000.0 ;
      RECT  94500.0 176100.0 93300.0 177300.0 ;
      RECT  93300.0 178800.0 92100.0 180000.0 ;
      RECT  99900.0 184950.0 85500.0 185850.0 ;
      RECT  99900.0 171150.0 85500.0 172050.0 ;
      RECT  98100.0 197250.0 96900.0 199650.0 ;
      RECT  98100.0 188550.0 96900.0 184950.0 ;
      RECT  93300.0 188550.0 92100.0 184950.0 ;
      RECT  90900.0 187350.0 89700.0 185400.0 ;
      RECT  90900.0 199200.0 89700.0 197250.0 ;
      RECT  98100.0 188550.0 96900.0 187350.0 ;
      RECT  95700.0 188550.0 94500.0 187350.0 ;
      RECT  95700.0 188550.0 94500.0 187350.0 ;
      RECT  98100.0 188550.0 96900.0 187350.0 ;
      RECT  95700.0 188550.0 94500.0 187350.0 ;
      RECT  93300.0 188550.0 92100.0 187350.0 ;
      RECT  93300.0 188550.0 92100.0 187350.0 ;
      RECT  95700.0 188550.0 94500.0 187350.0 ;
      RECT  98100.0 197250.0 96900.0 196050.0 ;
      RECT  95700.0 197250.0 94500.0 196050.0 ;
      RECT  95700.0 197250.0 94500.0 196050.0 ;
      RECT  98100.0 197250.0 96900.0 196050.0 ;
      RECT  95700.0 197250.0 94500.0 196050.0 ;
      RECT  93300.0 197250.0 92100.0 196050.0 ;
      RECT  93300.0 197250.0 92100.0 196050.0 ;
      RECT  95700.0 197250.0 94500.0 196050.0 ;
      RECT  90900.0 187950.0 89700.0 186750.0 ;
      RECT  90900.0 197850.0 89700.0 196650.0 ;
      RECT  93300.0 194700.0 94500.0 193500.0 ;
      RECT  96300.0 192000.0 97500.0 190800.0 ;
      RECT  95700.0 188550.0 94500.0 187350.0 ;
      RECT  93300.0 197250.0 92100.0 196050.0 ;
      RECT  92100.0 192000.0 93300.0 190800.0 ;
      RECT  97500.0 192000.0 96300.0 190800.0 ;
      RECT  94500.0 194700.0 93300.0 193500.0 ;
      RECT  93300.0 192000.0 92100.0 190800.0 ;
      RECT  99900.0 185850.0 85500.0 184950.0 ;
      RECT  99900.0 199650.0 85500.0 198750.0 ;
      RECT  110850.0 154500.0 112050.0 155700.0 ;
      RECT  129450.0 150000.0 130650.0 151200.0 ;
      RECT  107850.0 168300.0 109050.0 169500.0 ;
      RECT  126450.0 164400.0 127650.0 165600.0 ;
      RECT  129450.0 173100.0 130650.0 174300.0 ;
      RECT  104850.0 173100.0 106050.0 174300.0 ;
      RECT  126450.0 186900.0 127650.0 188100.0 ;
      RECT  101850.0 186900.0 103050.0 188100.0 ;
      RECT  110850.0 148500.0 112050.0 149700.0 ;
      RECT  107850.0 151200.0 109050.0 152400.0 ;
      RECT  104850.0 165900.0 106050.0 167100.0 ;
      RECT  107850.0 163200.0 109050.0 164400.0 ;
      RECT  110850.0 176100.0 112050.0 177300.0 ;
      RECT  101850.0 178800.0 103050.0 180000.0 ;
      RECT  104850.0 193500.0 106050.0 194700.0 ;
      RECT  101850.0 190800.0 103050.0 192000.0 ;
      RECT  79650.0 150150.0 75900.0 151050.0 ;
      RECT  79650.0 164550.0 75900.0 165450.0 ;
      RECT  79650.0 177750.0 75900.0 178650.0 ;
      RECT  79650.0 192150.0 75900.0 193050.0 ;
      RECT  130500.0 157350.0 75900.0 158250.0 ;
      RECT  130500.0 184950.0 75900.0 185850.0 ;
      RECT  130500.0 143550.0 75900.0 144450.0 ;
      RECT  130500.0 171150.0 75900.0 172050.0 ;
      RECT  130500.0 198750.0 75900.0 199650.0 ;
      RECT  77700.0 201150.0 78900.0 198750.0 ;
      RECT  77700.0 209850.0 78900.0 213450.0 ;
      RECT  82500.0 209850.0 83700.0 213450.0 ;
      RECT  84900.0 211050.0 86100.0 213000.0 ;
      RECT  84900.0 199200.0 86100.0 201150.0 ;
      RECT  77700.0 209850.0 78900.0 211050.0 ;
      RECT  80100.0 209850.0 81300.0 211050.0 ;
      RECT  80100.0 209850.0 81300.0 211050.0 ;
      RECT  77700.0 209850.0 78900.0 211050.0 ;
      RECT  80100.0 209850.0 81300.0 211050.0 ;
      RECT  82500.0 209850.0 83700.0 211050.0 ;
      RECT  82500.0 209850.0 83700.0 211050.0 ;
      RECT  80100.0 209850.0 81300.0 211050.0 ;
      RECT  77700.0 201150.0 78900.0 202350.0 ;
      RECT  80100.0 201150.0 81300.0 202350.0 ;
      RECT  80100.0 201150.0 81300.0 202350.0 ;
      RECT  77700.0 201150.0 78900.0 202350.0 ;
      RECT  80100.0 201150.0 81300.0 202350.0 ;
      RECT  82500.0 201150.0 83700.0 202350.0 ;
      RECT  82500.0 201150.0 83700.0 202350.0 ;
      RECT  80100.0 201150.0 81300.0 202350.0 ;
      RECT  84900.0 210450.0 86100.0 211650.0 ;
      RECT  84900.0 200550.0 86100.0 201750.0 ;
      RECT  82500.0 203700.0 81300.0 204900.0 ;
      RECT  79500.0 206400.0 78300.0 207600.0 ;
      RECT  80100.0 209850.0 81300.0 211050.0 ;
      RECT  82500.0 201150.0 83700.0 202350.0 ;
      RECT  83700.0 206400.0 82500.0 207600.0 ;
      RECT  78300.0 206400.0 79500.0 207600.0 ;
      RECT  81300.0 203700.0 82500.0 204900.0 ;
      RECT  82500.0 206400.0 83700.0 207600.0 ;
      RECT  75900.0 212550.0 90300.0 213450.0 ;
      RECT  75900.0 198750.0 90300.0 199650.0 ;
      RECT  77700.0 224850.0 78900.0 227250.0 ;
      RECT  77700.0 216150.0 78900.0 212550.0 ;
      RECT  82500.0 216150.0 83700.0 212550.0 ;
      RECT  84900.0 214950.0 86100.0 213000.0 ;
      RECT  84900.0 226800.0 86100.0 224850.0 ;
      RECT  77700.0 216150.0 78900.0 214950.0 ;
      RECT  80100.0 216150.0 81300.0 214950.0 ;
      RECT  80100.0 216150.0 81300.0 214950.0 ;
      RECT  77700.0 216150.0 78900.0 214950.0 ;
      RECT  80100.0 216150.0 81300.0 214950.0 ;
      RECT  82500.0 216150.0 83700.0 214950.0 ;
      RECT  82500.0 216150.0 83700.0 214950.0 ;
      RECT  80100.0 216150.0 81300.0 214950.0 ;
      RECT  77700.0 224850.0 78900.0 223650.0 ;
      RECT  80100.0 224850.0 81300.0 223650.0 ;
      RECT  80100.0 224850.0 81300.0 223650.0 ;
      RECT  77700.0 224850.0 78900.0 223650.0 ;
      RECT  80100.0 224850.0 81300.0 223650.0 ;
      RECT  82500.0 224850.0 83700.0 223650.0 ;
      RECT  82500.0 224850.0 83700.0 223650.0 ;
      RECT  80100.0 224850.0 81300.0 223650.0 ;
      RECT  84900.0 215550.0 86100.0 214350.0 ;
      RECT  84900.0 225450.0 86100.0 224250.0 ;
      RECT  82500.0 222300.0 81300.0 221100.0 ;
      RECT  79500.0 219600.0 78300.0 218400.0 ;
      RECT  80100.0 216150.0 81300.0 214950.0 ;
      RECT  82500.0 224850.0 83700.0 223650.0 ;
      RECT  83700.0 219600.0 82500.0 218400.0 ;
      RECT  78300.0 219600.0 79500.0 218400.0 ;
      RECT  81300.0 222300.0 82500.0 221100.0 ;
      RECT  82500.0 219600.0 83700.0 218400.0 ;
      RECT  75900.0 213450.0 90300.0 212550.0 ;
      RECT  75900.0 227250.0 90300.0 226350.0 ;
      RECT  77700.0 228750.0 78900.0 226350.0 ;
      RECT  77700.0 237450.0 78900.0 241050.0 ;
      RECT  82500.0 237450.0 83700.0 241050.0 ;
      RECT  84900.0 238650.0 86100.0 240600.0 ;
      RECT  84900.0 226800.0 86100.0 228750.0 ;
      RECT  77700.0 237450.0 78900.0 238650.0 ;
      RECT  80100.0 237450.0 81300.0 238650.0 ;
      RECT  80100.0 237450.0 81300.0 238650.0 ;
      RECT  77700.0 237450.0 78900.0 238650.0 ;
      RECT  80100.0 237450.0 81300.0 238650.0 ;
      RECT  82500.0 237450.0 83700.0 238650.0 ;
      RECT  82500.0 237450.0 83700.0 238650.0 ;
      RECT  80100.0 237450.0 81300.0 238650.0 ;
      RECT  77700.0 228750.0 78900.0 229950.0 ;
      RECT  80100.0 228750.0 81300.0 229950.0 ;
      RECT  80100.0 228750.0 81300.0 229950.0 ;
      RECT  77700.0 228750.0 78900.0 229950.0 ;
      RECT  80100.0 228750.0 81300.0 229950.0 ;
      RECT  82500.0 228750.0 83700.0 229950.0 ;
      RECT  82500.0 228750.0 83700.0 229950.0 ;
      RECT  80100.0 228750.0 81300.0 229950.0 ;
      RECT  84900.0 238050.0 86100.0 239250.0 ;
      RECT  84900.0 228150.0 86100.0 229350.0 ;
      RECT  82500.0 231300.0 81300.0 232500.0 ;
      RECT  79500.0 234000.0 78300.0 235200.0 ;
      RECT  80100.0 237450.0 81300.0 238650.0 ;
      RECT  82500.0 228750.0 83700.0 229950.0 ;
      RECT  83700.0 234000.0 82500.0 235200.0 ;
      RECT  78300.0 234000.0 79500.0 235200.0 ;
      RECT  81300.0 231300.0 82500.0 232500.0 ;
      RECT  82500.0 234000.0 83700.0 235200.0 ;
      RECT  75900.0 240150.0 90300.0 241050.0 ;
      RECT  75900.0 226350.0 90300.0 227250.0 ;
      RECT  77700.0 252450.0 78900.0 254850.0 ;
      RECT  77700.0 243750.0 78900.0 240150.0 ;
      RECT  82500.0 243750.0 83700.0 240150.0 ;
      RECT  84900.0 242550.0 86100.0 240600.0 ;
      RECT  84900.0 254400.0 86100.0 252450.0 ;
      RECT  77700.0 243750.0 78900.0 242550.0 ;
      RECT  80100.0 243750.0 81300.0 242550.0 ;
      RECT  80100.0 243750.0 81300.0 242550.0 ;
      RECT  77700.0 243750.0 78900.0 242550.0 ;
      RECT  80100.0 243750.0 81300.0 242550.0 ;
      RECT  82500.0 243750.0 83700.0 242550.0 ;
      RECT  82500.0 243750.0 83700.0 242550.0 ;
      RECT  80100.0 243750.0 81300.0 242550.0 ;
      RECT  77700.0 252450.0 78900.0 251250.0 ;
      RECT  80100.0 252450.0 81300.0 251250.0 ;
      RECT  80100.0 252450.0 81300.0 251250.0 ;
      RECT  77700.0 252450.0 78900.0 251250.0 ;
      RECT  80100.0 252450.0 81300.0 251250.0 ;
      RECT  82500.0 252450.0 83700.0 251250.0 ;
      RECT  82500.0 252450.0 83700.0 251250.0 ;
      RECT  80100.0 252450.0 81300.0 251250.0 ;
      RECT  84900.0 243150.0 86100.0 241950.0 ;
      RECT  84900.0 253050.0 86100.0 251850.0 ;
      RECT  82500.0 249900.0 81300.0 248700.0 ;
      RECT  79500.0 247200.0 78300.0 246000.0 ;
      RECT  80100.0 243750.0 81300.0 242550.0 ;
      RECT  82500.0 252450.0 83700.0 251250.0 ;
      RECT  83700.0 247200.0 82500.0 246000.0 ;
      RECT  78300.0 247200.0 79500.0 246000.0 ;
      RECT  81300.0 249900.0 82500.0 248700.0 ;
      RECT  82500.0 247200.0 83700.0 246000.0 ;
      RECT  75900.0 241050.0 90300.0 240150.0 ;
      RECT  75900.0 254850.0 90300.0 253950.0 ;
      RECT  77700.0 256350.0 78900.0 253950.0 ;
      RECT  77700.0 265050.0 78900.0 268650.0 ;
      RECT  82500.0 265050.0 83700.0 268650.0 ;
      RECT  84900.0 266250.0 86100.0 268200.0 ;
      RECT  84900.0 254400.0 86100.0 256350.0 ;
      RECT  77700.0 265050.0 78900.0 266250.0 ;
      RECT  80100.0 265050.0 81300.0 266250.0 ;
      RECT  80100.0 265050.0 81300.0 266250.0 ;
      RECT  77700.0 265050.0 78900.0 266250.0 ;
      RECT  80100.0 265050.0 81300.0 266250.0 ;
      RECT  82500.0 265050.0 83700.0 266250.0 ;
      RECT  82500.0 265050.0 83700.0 266250.0 ;
      RECT  80100.0 265050.0 81300.0 266250.0 ;
      RECT  77700.0 256350.0 78900.0 257550.0 ;
      RECT  80100.0 256350.0 81300.0 257550.0 ;
      RECT  80100.0 256350.0 81300.0 257550.0 ;
      RECT  77700.0 256350.0 78900.0 257550.0 ;
      RECT  80100.0 256350.0 81300.0 257550.0 ;
      RECT  82500.0 256350.0 83700.0 257550.0 ;
      RECT  82500.0 256350.0 83700.0 257550.0 ;
      RECT  80100.0 256350.0 81300.0 257550.0 ;
      RECT  84900.0 265650.0 86100.0 266850.0 ;
      RECT  84900.0 255750.0 86100.0 256950.0 ;
      RECT  82500.0 258900.0 81300.0 260100.0 ;
      RECT  79500.0 261600.0 78300.0 262800.0 ;
      RECT  80100.0 265050.0 81300.0 266250.0 ;
      RECT  82500.0 256350.0 83700.0 257550.0 ;
      RECT  83700.0 261600.0 82500.0 262800.0 ;
      RECT  78300.0 261600.0 79500.0 262800.0 ;
      RECT  81300.0 258900.0 82500.0 260100.0 ;
      RECT  82500.0 261600.0 83700.0 262800.0 ;
      RECT  75900.0 267750.0 90300.0 268650.0 ;
      RECT  75900.0 253950.0 90300.0 254850.0 ;
      RECT  77700.0 280050.0 78900.0 282450.0 ;
      RECT  77700.0 271350.0 78900.0 267750.0 ;
      RECT  82500.0 271350.0 83700.0 267750.0 ;
      RECT  84900.0 270150.0 86100.0 268200.0 ;
      RECT  84900.0 282000.0 86100.0 280050.0 ;
      RECT  77700.0 271350.0 78900.0 270150.0 ;
      RECT  80100.0 271350.0 81300.0 270150.0 ;
      RECT  80100.0 271350.0 81300.0 270150.0 ;
      RECT  77700.0 271350.0 78900.0 270150.0 ;
      RECT  80100.0 271350.0 81300.0 270150.0 ;
      RECT  82500.0 271350.0 83700.0 270150.0 ;
      RECT  82500.0 271350.0 83700.0 270150.0 ;
      RECT  80100.0 271350.0 81300.0 270150.0 ;
      RECT  77700.0 280050.0 78900.0 278850.0 ;
      RECT  80100.0 280050.0 81300.0 278850.0 ;
      RECT  80100.0 280050.0 81300.0 278850.0 ;
      RECT  77700.0 280050.0 78900.0 278850.0 ;
      RECT  80100.0 280050.0 81300.0 278850.0 ;
      RECT  82500.0 280050.0 83700.0 278850.0 ;
      RECT  82500.0 280050.0 83700.0 278850.0 ;
      RECT  80100.0 280050.0 81300.0 278850.0 ;
      RECT  84900.0 270750.0 86100.0 269550.0 ;
      RECT  84900.0 280650.0 86100.0 279450.0 ;
      RECT  82500.0 277500.0 81300.0 276300.0 ;
      RECT  79500.0 274800.0 78300.0 273600.0 ;
      RECT  80100.0 271350.0 81300.0 270150.0 ;
      RECT  82500.0 280050.0 83700.0 278850.0 ;
      RECT  83700.0 274800.0 82500.0 273600.0 ;
      RECT  78300.0 274800.0 79500.0 273600.0 ;
      RECT  81300.0 277500.0 82500.0 276300.0 ;
      RECT  82500.0 274800.0 83700.0 273600.0 ;
      RECT  75900.0 268650.0 90300.0 267750.0 ;
      RECT  75900.0 282450.0 90300.0 281550.0 ;
      RECT  77700.0 283950.0 78900.0 281550.0 ;
      RECT  77700.0 292650.0 78900.0 296250.0 ;
      RECT  82500.0 292650.0 83700.0 296250.0 ;
      RECT  84900.0 293850.0 86100.0 295800.0 ;
      RECT  84900.0 282000.0 86100.0 283950.0 ;
      RECT  77700.0 292650.0 78900.0 293850.0 ;
      RECT  80100.0 292650.0 81300.0 293850.0 ;
      RECT  80100.0 292650.0 81300.0 293850.0 ;
      RECT  77700.0 292650.0 78900.0 293850.0 ;
      RECT  80100.0 292650.0 81300.0 293850.0 ;
      RECT  82500.0 292650.0 83700.0 293850.0 ;
      RECT  82500.0 292650.0 83700.0 293850.0 ;
      RECT  80100.0 292650.0 81300.0 293850.0 ;
      RECT  77700.0 283950.0 78900.0 285150.0 ;
      RECT  80100.0 283950.0 81300.0 285150.0 ;
      RECT  80100.0 283950.0 81300.0 285150.0 ;
      RECT  77700.0 283950.0 78900.0 285150.0 ;
      RECT  80100.0 283950.0 81300.0 285150.0 ;
      RECT  82500.0 283950.0 83700.0 285150.0 ;
      RECT  82500.0 283950.0 83700.0 285150.0 ;
      RECT  80100.0 283950.0 81300.0 285150.0 ;
      RECT  84900.0 293250.0 86100.0 294450.0 ;
      RECT  84900.0 283350.0 86100.0 284550.0 ;
      RECT  82500.0 286500.0 81300.0 287700.0 ;
      RECT  79500.0 289200.0 78300.0 290400.0 ;
      RECT  80100.0 292650.0 81300.0 293850.0 ;
      RECT  82500.0 283950.0 83700.0 285150.0 ;
      RECT  83700.0 289200.0 82500.0 290400.0 ;
      RECT  78300.0 289200.0 79500.0 290400.0 ;
      RECT  81300.0 286500.0 82500.0 287700.0 ;
      RECT  82500.0 289200.0 83700.0 290400.0 ;
      RECT  75900.0 295350.0 90300.0 296250.0 ;
      RECT  75900.0 281550.0 90300.0 282450.0 ;
      RECT  77700.0 307650.0 78900.0 310050.0 ;
      RECT  77700.0 298950.0 78900.0 295350.0 ;
      RECT  82500.0 298950.0 83700.0 295350.0 ;
      RECT  84900.0 297750.0 86100.0 295800.0 ;
      RECT  84900.0 309600.0 86100.0 307650.0 ;
      RECT  77700.0 298950.0 78900.0 297750.0 ;
      RECT  80100.0 298950.0 81300.0 297750.0 ;
      RECT  80100.0 298950.0 81300.0 297750.0 ;
      RECT  77700.0 298950.0 78900.0 297750.0 ;
      RECT  80100.0 298950.0 81300.0 297750.0 ;
      RECT  82500.0 298950.0 83700.0 297750.0 ;
      RECT  82500.0 298950.0 83700.0 297750.0 ;
      RECT  80100.0 298950.0 81300.0 297750.0 ;
      RECT  77700.0 307650.0 78900.0 306450.0 ;
      RECT  80100.0 307650.0 81300.0 306450.0 ;
      RECT  80100.0 307650.0 81300.0 306450.0 ;
      RECT  77700.0 307650.0 78900.0 306450.0 ;
      RECT  80100.0 307650.0 81300.0 306450.0 ;
      RECT  82500.0 307650.0 83700.0 306450.0 ;
      RECT  82500.0 307650.0 83700.0 306450.0 ;
      RECT  80100.0 307650.0 81300.0 306450.0 ;
      RECT  84900.0 298350.0 86100.0 297150.0 ;
      RECT  84900.0 308250.0 86100.0 307050.0 ;
      RECT  82500.0 305100.0 81300.0 303900.0 ;
      RECT  79500.0 302400.0 78300.0 301200.0 ;
      RECT  80100.0 298950.0 81300.0 297750.0 ;
      RECT  82500.0 307650.0 83700.0 306450.0 ;
      RECT  83700.0 302400.0 82500.0 301200.0 ;
      RECT  78300.0 302400.0 79500.0 301200.0 ;
      RECT  81300.0 305100.0 82500.0 303900.0 ;
      RECT  82500.0 302400.0 83700.0 301200.0 ;
      RECT  75900.0 296250.0 90300.0 295350.0 ;
      RECT  75900.0 310050.0 90300.0 309150.0 ;
      RECT  77700.0 311550.0 78900.0 309150.0 ;
      RECT  77700.0 320250.0 78900.0 323850.0 ;
      RECT  82500.0 320250.0 83700.0 323850.0 ;
      RECT  84900.0 321450.0 86100.0 323400.0 ;
      RECT  84900.0 309600.0 86100.0 311550.0 ;
      RECT  77700.0 320250.0 78900.0 321450.0 ;
      RECT  80100.0 320250.0 81300.0 321450.0 ;
      RECT  80100.0 320250.0 81300.0 321450.0 ;
      RECT  77700.0 320250.0 78900.0 321450.0 ;
      RECT  80100.0 320250.0 81300.0 321450.0 ;
      RECT  82500.0 320250.0 83700.0 321450.0 ;
      RECT  82500.0 320250.0 83700.0 321450.0 ;
      RECT  80100.0 320250.0 81300.0 321450.0 ;
      RECT  77700.0 311550.0 78900.0 312750.0 ;
      RECT  80100.0 311550.0 81300.0 312750.0 ;
      RECT  80100.0 311550.0 81300.0 312750.0 ;
      RECT  77700.0 311550.0 78900.0 312750.0 ;
      RECT  80100.0 311550.0 81300.0 312750.0 ;
      RECT  82500.0 311550.0 83700.0 312750.0 ;
      RECT  82500.0 311550.0 83700.0 312750.0 ;
      RECT  80100.0 311550.0 81300.0 312750.0 ;
      RECT  84900.0 320850.0 86100.0 322050.0 ;
      RECT  84900.0 310950.0 86100.0 312150.0 ;
      RECT  82500.0 314100.0 81300.0 315300.0 ;
      RECT  79500.0 316800.0 78300.0 318000.0 ;
      RECT  80100.0 320250.0 81300.0 321450.0 ;
      RECT  82500.0 311550.0 83700.0 312750.0 ;
      RECT  83700.0 316800.0 82500.0 318000.0 ;
      RECT  78300.0 316800.0 79500.0 318000.0 ;
      RECT  81300.0 314100.0 82500.0 315300.0 ;
      RECT  82500.0 316800.0 83700.0 318000.0 ;
      RECT  75900.0 322950.0 90300.0 323850.0 ;
      RECT  75900.0 309150.0 90300.0 310050.0 ;
      RECT  77700.0 335250.0 78900.0 337650.0 ;
      RECT  77700.0 326550.0 78900.0 322950.0 ;
      RECT  82500.0 326550.0 83700.0 322950.0 ;
      RECT  84900.0 325350.0 86100.0 323400.0 ;
      RECT  84900.0 337200.0 86100.0 335250.0 ;
      RECT  77700.0 326550.0 78900.0 325350.0 ;
      RECT  80100.0 326550.0 81300.0 325350.0 ;
      RECT  80100.0 326550.0 81300.0 325350.0 ;
      RECT  77700.0 326550.0 78900.0 325350.0 ;
      RECT  80100.0 326550.0 81300.0 325350.0 ;
      RECT  82500.0 326550.0 83700.0 325350.0 ;
      RECT  82500.0 326550.0 83700.0 325350.0 ;
      RECT  80100.0 326550.0 81300.0 325350.0 ;
      RECT  77700.0 335250.0 78900.0 334050.0 ;
      RECT  80100.0 335250.0 81300.0 334050.0 ;
      RECT  80100.0 335250.0 81300.0 334050.0 ;
      RECT  77700.0 335250.0 78900.0 334050.0 ;
      RECT  80100.0 335250.0 81300.0 334050.0 ;
      RECT  82500.0 335250.0 83700.0 334050.0 ;
      RECT  82500.0 335250.0 83700.0 334050.0 ;
      RECT  80100.0 335250.0 81300.0 334050.0 ;
      RECT  84900.0 325950.0 86100.0 324750.0 ;
      RECT  84900.0 335850.0 86100.0 334650.0 ;
      RECT  82500.0 332700.0 81300.0 331500.0 ;
      RECT  79500.0 330000.0 78300.0 328800.0 ;
      RECT  80100.0 326550.0 81300.0 325350.0 ;
      RECT  82500.0 335250.0 83700.0 334050.0 ;
      RECT  83700.0 330000.0 82500.0 328800.0 ;
      RECT  78300.0 330000.0 79500.0 328800.0 ;
      RECT  81300.0 332700.0 82500.0 331500.0 ;
      RECT  82500.0 330000.0 83700.0 328800.0 ;
      RECT  75900.0 323850.0 90300.0 322950.0 ;
      RECT  75900.0 337650.0 90300.0 336750.0 ;
      RECT  77700.0 339150.0 78900.0 336750.0 ;
      RECT  77700.0 347850.0 78900.0 351450.0 ;
      RECT  82500.0 347850.0 83700.0 351450.0 ;
      RECT  84900.0 349050.0 86100.0 351000.0 ;
      RECT  84900.0 337200.0 86100.0 339150.0 ;
      RECT  77700.0 347850.0 78900.0 349050.0 ;
      RECT  80100.0 347850.0 81300.0 349050.0 ;
      RECT  80100.0 347850.0 81300.0 349050.0 ;
      RECT  77700.0 347850.0 78900.0 349050.0 ;
      RECT  80100.0 347850.0 81300.0 349050.0 ;
      RECT  82500.0 347850.0 83700.0 349050.0 ;
      RECT  82500.0 347850.0 83700.0 349050.0 ;
      RECT  80100.0 347850.0 81300.0 349050.0 ;
      RECT  77700.0 339150.0 78900.0 340350.0 ;
      RECT  80100.0 339150.0 81300.0 340350.0 ;
      RECT  80100.0 339150.0 81300.0 340350.0 ;
      RECT  77700.0 339150.0 78900.0 340350.0 ;
      RECT  80100.0 339150.0 81300.0 340350.0 ;
      RECT  82500.0 339150.0 83700.0 340350.0 ;
      RECT  82500.0 339150.0 83700.0 340350.0 ;
      RECT  80100.0 339150.0 81300.0 340350.0 ;
      RECT  84900.0 348450.0 86100.0 349650.0 ;
      RECT  84900.0 338550.0 86100.0 339750.0 ;
      RECT  82500.0 341700.0 81300.0 342900.0 ;
      RECT  79500.0 344400.0 78300.0 345600.0 ;
      RECT  80100.0 347850.0 81300.0 349050.0 ;
      RECT  82500.0 339150.0 83700.0 340350.0 ;
      RECT  83700.0 344400.0 82500.0 345600.0 ;
      RECT  78300.0 344400.0 79500.0 345600.0 ;
      RECT  81300.0 341700.0 82500.0 342900.0 ;
      RECT  82500.0 344400.0 83700.0 345600.0 ;
      RECT  75900.0 350550.0 90300.0 351450.0 ;
      RECT  75900.0 336750.0 90300.0 337650.0 ;
      RECT  77700.0 362850.0 78900.0 365250.0 ;
      RECT  77700.0 354150.0 78900.0 350550.0 ;
      RECT  82500.0 354150.0 83700.0 350550.0 ;
      RECT  84900.0 352950.0 86100.0 351000.0 ;
      RECT  84900.0 364800.0 86100.0 362850.0 ;
      RECT  77700.0 354150.0 78900.0 352950.0 ;
      RECT  80100.0 354150.0 81300.0 352950.0 ;
      RECT  80100.0 354150.0 81300.0 352950.0 ;
      RECT  77700.0 354150.0 78900.0 352950.0 ;
      RECT  80100.0 354150.0 81300.0 352950.0 ;
      RECT  82500.0 354150.0 83700.0 352950.0 ;
      RECT  82500.0 354150.0 83700.0 352950.0 ;
      RECT  80100.0 354150.0 81300.0 352950.0 ;
      RECT  77700.0 362850.0 78900.0 361650.0 ;
      RECT  80100.0 362850.0 81300.0 361650.0 ;
      RECT  80100.0 362850.0 81300.0 361650.0 ;
      RECT  77700.0 362850.0 78900.0 361650.0 ;
      RECT  80100.0 362850.0 81300.0 361650.0 ;
      RECT  82500.0 362850.0 83700.0 361650.0 ;
      RECT  82500.0 362850.0 83700.0 361650.0 ;
      RECT  80100.0 362850.0 81300.0 361650.0 ;
      RECT  84900.0 353550.0 86100.0 352350.0 ;
      RECT  84900.0 363450.0 86100.0 362250.0 ;
      RECT  82500.0 360300.0 81300.0 359100.0 ;
      RECT  79500.0 357600.0 78300.0 356400.0 ;
      RECT  80100.0 354150.0 81300.0 352950.0 ;
      RECT  82500.0 362850.0 83700.0 361650.0 ;
      RECT  83700.0 357600.0 82500.0 356400.0 ;
      RECT  78300.0 357600.0 79500.0 356400.0 ;
      RECT  81300.0 360300.0 82500.0 359100.0 ;
      RECT  82500.0 357600.0 83700.0 356400.0 ;
      RECT  75900.0 351450.0 90300.0 350550.0 ;
      RECT  75900.0 365250.0 90300.0 364350.0 ;
      RECT  77700.0 366750.0 78900.0 364350.0 ;
      RECT  77700.0 375450.0 78900.0 379050.0 ;
      RECT  82500.0 375450.0 83700.0 379050.0 ;
      RECT  84900.0 376650.0 86100.0 378600.0 ;
      RECT  84900.0 364800.0 86100.0 366750.0 ;
      RECT  77700.0 375450.0 78900.0 376650.0 ;
      RECT  80100.0 375450.0 81300.0 376650.0 ;
      RECT  80100.0 375450.0 81300.0 376650.0 ;
      RECT  77700.0 375450.0 78900.0 376650.0 ;
      RECT  80100.0 375450.0 81300.0 376650.0 ;
      RECT  82500.0 375450.0 83700.0 376650.0 ;
      RECT  82500.0 375450.0 83700.0 376650.0 ;
      RECT  80100.0 375450.0 81300.0 376650.0 ;
      RECT  77700.0 366750.0 78900.0 367950.0 ;
      RECT  80100.0 366750.0 81300.0 367950.0 ;
      RECT  80100.0 366750.0 81300.0 367950.0 ;
      RECT  77700.0 366750.0 78900.0 367950.0 ;
      RECT  80100.0 366750.0 81300.0 367950.0 ;
      RECT  82500.0 366750.0 83700.0 367950.0 ;
      RECT  82500.0 366750.0 83700.0 367950.0 ;
      RECT  80100.0 366750.0 81300.0 367950.0 ;
      RECT  84900.0 376050.0 86100.0 377250.0 ;
      RECT  84900.0 366150.0 86100.0 367350.0 ;
      RECT  82500.0 369300.0 81300.0 370500.0 ;
      RECT  79500.0 372000.0 78300.0 373200.0 ;
      RECT  80100.0 375450.0 81300.0 376650.0 ;
      RECT  82500.0 366750.0 83700.0 367950.0 ;
      RECT  83700.0 372000.0 82500.0 373200.0 ;
      RECT  78300.0 372000.0 79500.0 373200.0 ;
      RECT  81300.0 369300.0 82500.0 370500.0 ;
      RECT  82500.0 372000.0 83700.0 373200.0 ;
      RECT  75900.0 378150.0 90300.0 379050.0 ;
      RECT  75900.0 364350.0 90300.0 365250.0 ;
      RECT  77700.0 390450.0 78900.0 392850.0 ;
      RECT  77700.0 381750.0 78900.0 378150.0 ;
      RECT  82500.0 381750.0 83700.0 378150.0 ;
      RECT  84900.0 380550.0 86100.0 378600.0 ;
      RECT  84900.0 392400.0 86100.0 390450.0 ;
      RECT  77700.0 381750.0 78900.0 380550.0 ;
      RECT  80100.0 381750.0 81300.0 380550.0 ;
      RECT  80100.0 381750.0 81300.0 380550.0 ;
      RECT  77700.0 381750.0 78900.0 380550.0 ;
      RECT  80100.0 381750.0 81300.0 380550.0 ;
      RECT  82500.0 381750.0 83700.0 380550.0 ;
      RECT  82500.0 381750.0 83700.0 380550.0 ;
      RECT  80100.0 381750.0 81300.0 380550.0 ;
      RECT  77700.0 390450.0 78900.0 389250.0 ;
      RECT  80100.0 390450.0 81300.0 389250.0 ;
      RECT  80100.0 390450.0 81300.0 389250.0 ;
      RECT  77700.0 390450.0 78900.0 389250.0 ;
      RECT  80100.0 390450.0 81300.0 389250.0 ;
      RECT  82500.0 390450.0 83700.0 389250.0 ;
      RECT  82500.0 390450.0 83700.0 389250.0 ;
      RECT  80100.0 390450.0 81300.0 389250.0 ;
      RECT  84900.0 381150.0 86100.0 379950.0 ;
      RECT  84900.0 391050.0 86100.0 389850.0 ;
      RECT  82500.0 387900.0 81300.0 386700.0 ;
      RECT  79500.0 385200.0 78300.0 384000.0 ;
      RECT  80100.0 381750.0 81300.0 380550.0 ;
      RECT  82500.0 390450.0 83700.0 389250.0 ;
      RECT  83700.0 385200.0 82500.0 384000.0 ;
      RECT  78300.0 385200.0 79500.0 384000.0 ;
      RECT  81300.0 387900.0 82500.0 386700.0 ;
      RECT  82500.0 385200.0 83700.0 384000.0 ;
      RECT  75900.0 379050.0 90300.0 378150.0 ;
      RECT  75900.0 392850.0 90300.0 391950.0 ;
      RECT  77700.0 394350.0 78900.0 391950.0 ;
      RECT  77700.0 403050.0 78900.0 406650.0 ;
      RECT  82500.0 403050.0 83700.0 406650.0 ;
      RECT  84900.0 404250.0 86100.0 406200.0 ;
      RECT  84900.0 392400.0 86100.0 394350.0 ;
      RECT  77700.0 403050.0 78900.0 404250.0 ;
      RECT  80100.0 403050.0 81300.0 404250.0 ;
      RECT  80100.0 403050.0 81300.0 404250.0 ;
      RECT  77700.0 403050.0 78900.0 404250.0 ;
      RECT  80100.0 403050.0 81300.0 404250.0 ;
      RECT  82500.0 403050.0 83700.0 404250.0 ;
      RECT  82500.0 403050.0 83700.0 404250.0 ;
      RECT  80100.0 403050.0 81300.0 404250.0 ;
      RECT  77700.0 394350.0 78900.0 395550.0 ;
      RECT  80100.0 394350.0 81300.0 395550.0 ;
      RECT  80100.0 394350.0 81300.0 395550.0 ;
      RECT  77700.0 394350.0 78900.0 395550.0 ;
      RECT  80100.0 394350.0 81300.0 395550.0 ;
      RECT  82500.0 394350.0 83700.0 395550.0 ;
      RECT  82500.0 394350.0 83700.0 395550.0 ;
      RECT  80100.0 394350.0 81300.0 395550.0 ;
      RECT  84900.0 403650.0 86100.0 404850.0 ;
      RECT  84900.0 393750.0 86100.0 394950.0 ;
      RECT  82500.0 396900.0 81300.0 398100.0 ;
      RECT  79500.0 399600.0 78300.0 400800.0 ;
      RECT  80100.0 403050.0 81300.0 404250.0 ;
      RECT  82500.0 394350.0 83700.0 395550.0 ;
      RECT  83700.0 399600.0 82500.0 400800.0 ;
      RECT  78300.0 399600.0 79500.0 400800.0 ;
      RECT  81300.0 396900.0 82500.0 398100.0 ;
      RECT  82500.0 399600.0 83700.0 400800.0 ;
      RECT  75900.0 405750.0 90300.0 406650.0 ;
      RECT  75900.0 391950.0 90300.0 392850.0 ;
      RECT  77700.0 418050.0 78900.0 420450.0 ;
      RECT  77700.0 409350.0 78900.0 405750.0 ;
      RECT  82500.0 409350.0 83700.0 405750.0 ;
      RECT  84900.0 408150.0 86100.0 406200.0 ;
      RECT  84900.0 420000.0 86100.0 418050.0 ;
      RECT  77700.0 409350.0 78900.0 408150.0 ;
      RECT  80100.0 409350.0 81300.0 408150.0 ;
      RECT  80100.0 409350.0 81300.0 408150.0 ;
      RECT  77700.0 409350.0 78900.0 408150.0 ;
      RECT  80100.0 409350.0 81300.0 408150.0 ;
      RECT  82500.0 409350.0 83700.0 408150.0 ;
      RECT  82500.0 409350.0 83700.0 408150.0 ;
      RECT  80100.0 409350.0 81300.0 408150.0 ;
      RECT  77700.0 418050.0 78900.0 416850.0 ;
      RECT  80100.0 418050.0 81300.0 416850.0 ;
      RECT  80100.0 418050.0 81300.0 416850.0 ;
      RECT  77700.0 418050.0 78900.0 416850.0 ;
      RECT  80100.0 418050.0 81300.0 416850.0 ;
      RECT  82500.0 418050.0 83700.0 416850.0 ;
      RECT  82500.0 418050.0 83700.0 416850.0 ;
      RECT  80100.0 418050.0 81300.0 416850.0 ;
      RECT  84900.0 408750.0 86100.0 407550.0 ;
      RECT  84900.0 418650.0 86100.0 417450.0 ;
      RECT  82500.0 415500.0 81300.0 414300.0 ;
      RECT  79500.0 412800.0 78300.0 411600.0 ;
      RECT  80100.0 409350.0 81300.0 408150.0 ;
      RECT  82500.0 418050.0 83700.0 416850.0 ;
      RECT  83700.0 412800.0 82500.0 411600.0 ;
      RECT  78300.0 412800.0 79500.0 411600.0 ;
      RECT  81300.0 415500.0 82500.0 414300.0 ;
      RECT  82500.0 412800.0 83700.0 411600.0 ;
      RECT  75900.0 406650.0 90300.0 405750.0 ;
      RECT  75900.0 420450.0 90300.0 419550.0 ;
      RECT  96900.0 211050.0 98100.0 213000.0 ;
      RECT  96900.0 199200.0 98100.0 201150.0 ;
      RECT  92100.0 200550.0 93300.0 198750.0 ;
      RECT  92100.0 209850.0 93300.0 213450.0 ;
      RECT  94800.0 200550.0 95700.0 209850.0 ;
      RECT  92100.0 209850.0 93300.0 211050.0 ;
      RECT  94500.0 209850.0 95700.0 211050.0 ;
      RECT  94500.0 209850.0 95700.0 211050.0 ;
      RECT  92100.0 209850.0 93300.0 211050.0 ;
      RECT  92100.0 200550.0 93300.0 201750.0 ;
      RECT  94500.0 200550.0 95700.0 201750.0 ;
      RECT  94500.0 200550.0 95700.0 201750.0 ;
      RECT  92100.0 200550.0 93300.0 201750.0 ;
      RECT  96900.0 210450.0 98100.0 211650.0 ;
      RECT  96900.0 200550.0 98100.0 201750.0 ;
      RECT  92700.0 205200.0 93900.0 206400.0 ;
      RECT  92700.0 205200.0 93900.0 206400.0 ;
      RECT  95250.0 205350.0 96150.0 206250.0 ;
      RECT  90300.0 212550.0 99900.0 213450.0 ;
      RECT  90300.0 198750.0 99900.0 199650.0 ;
      RECT  96900.0 214950.0 98100.0 213000.0 ;
      RECT  96900.0 226800.0 98100.0 224850.0 ;
      RECT  92100.0 225450.0 93300.0 227250.0 ;
      RECT  92100.0 216150.0 93300.0 212550.0 ;
      RECT  94800.0 225450.0 95700.0 216150.0 ;
      RECT  92100.0 216150.0 93300.0 214950.0 ;
      RECT  94500.0 216150.0 95700.0 214950.0 ;
      RECT  94500.0 216150.0 95700.0 214950.0 ;
      RECT  92100.0 216150.0 93300.0 214950.0 ;
      RECT  92100.0 225450.0 93300.0 224250.0 ;
      RECT  94500.0 225450.0 95700.0 224250.0 ;
      RECT  94500.0 225450.0 95700.0 224250.0 ;
      RECT  92100.0 225450.0 93300.0 224250.0 ;
      RECT  96900.0 215550.0 98100.0 214350.0 ;
      RECT  96900.0 225450.0 98100.0 224250.0 ;
      RECT  92700.0 220800.0 93900.0 219600.0 ;
      RECT  92700.0 220800.0 93900.0 219600.0 ;
      RECT  95250.0 220650.0 96150.0 219750.0 ;
      RECT  90300.0 213450.0 99900.0 212550.0 ;
      RECT  90300.0 227250.0 99900.0 226350.0 ;
      RECT  96900.0 238650.0 98100.0 240600.0 ;
      RECT  96900.0 226800.0 98100.0 228750.0 ;
      RECT  92100.0 228150.0 93300.0 226350.0 ;
      RECT  92100.0 237450.0 93300.0 241050.0 ;
      RECT  94800.0 228150.0 95700.0 237450.0 ;
      RECT  92100.0 237450.0 93300.0 238650.0 ;
      RECT  94500.0 237450.0 95700.0 238650.0 ;
      RECT  94500.0 237450.0 95700.0 238650.0 ;
      RECT  92100.0 237450.0 93300.0 238650.0 ;
      RECT  92100.0 228150.0 93300.0 229350.0 ;
      RECT  94500.0 228150.0 95700.0 229350.0 ;
      RECT  94500.0 228150.0 95700.0 229350.0 ;
      RECT  92100.0 228150.0 93300.0 229350.0 ;
      RECT  96900.0 238050.0 98100.0 239250.0 ;
      RECT  96900.0 228150.0 98100.0 229350.0 ;
      RECT  92700.0 232800.0 93900.0 234000.0 ;
      RECT  92700.0 232800.0 93900.0 234000.0 ;
      RECT  95250.0 232950.0 96150.0 233850.0 ;
      RECT  90300.0 240150.0 99900.0 241050.0 ;
      RECT  90300.0 226350.0 99900.0 227250.0 ;
      RECT  96900.0 242550.0 98100.0 240600.0 ;
      RECT  96900.0 254400.0 98100.0 252450.0 ;
      RECT  92100.0 253050.0 93300.0 254850.0 ;
      RECT  92100.0 243750.0 93300.0 240150.0 ;
      RECT  94800.0 253050.0 95700.0 243750.0 ;
      RECT  92100.0 243750.0 93300.0 242550.0 ;
      RECT  94500.0 243750.0 95700.0 242550.0 ;
      RECT  94500.0 243750.0 95700.0 242550.0 ;
      RECT  92100.0 243750.0 93300.0 242550.0 ;
      RECT  92100.0 253050.0 93300.0 251850.0 ;
      RECT  94500.0 253050.0 95700.0 251850.0 ;
      RECT  94500.0 253050.0 95700.0 251850.0 ;
      RECT  92100.0 253050.0 93300.0 251850.0 ;
      RECT  96900.0 243150.0 98100.0 241950.0 ;
      RECT  96900.0 253050.0 98100.0 251850.0 ;
      RECT  92700.0 248400.0 93900.0 247200.0 ;
      RECT  92700.0 248400.0 93900.0 247200.0 ;
      RECT  95250.0 248250.0 96150.0 247350.0 ;
      RECT  90300.0 241050.0 99900.0 240150.0 ;
      RECT  90300.0 254850.0 99900.0 253950.0 ;
      RECT  96900.0 266250.0 98100.0 268200.0 ;
      RECT  96900.0 254400.0 98100.0 256350.0 ;
      RECT  92100.0 255750.0 93300.0 253950.0 ;
      RECT  92100.0 265050.0 93300.0 268650.0 ;
      RECT  94800.0 255750.0 95700.0 265050.0 ;
      RECT  92100.0 265050.0 93300.0 266250.0 ;
      RECT  94500.0 265050.0 95700.0 266250.0 ;
      RECT  94500.0 265050.0 95700.0 266250.0 ;
      RECT  92100.0 265050.0 93300.0 266250.0 ;
      RECT  92100.0 255750.0 93300.0 256950.0 ;
      RECT  94500.0 255750.0 95700.0 256950.0 ;
      RECT  94500.0 255750.0 95700.0 256950.0 ;
      RECT  92100.0 255750.0 93300.0 256950.0 ;
      RECT  96900.0 265650.0 98100.0 266850.0 ;
      RECT  96900.0 255750.0 98100.0 256950.0 ;
      RECT  92700.0 260400.0 93900.0 261600.0 ;
      RECT  92700.0 260400.0 93900.0 261600.0 ;
      RECT  95250.0 260550.0 96150.0 261450.0 ;
      RECT  90300.0 267750.0 99900.0 268650.0 ;
      RECT  90300.0 253950.0 99900.0 254850.0 ;
      RECT  96900.0 270150.0 98100.0 268200.0 ;
      RECT  96900.0 282000.0 98100.0 280050.0 ;
      RECT  92100.0 280650.0 93300.0 282450.0 ;
      RECT  92100.0 271350.0 93300.0 267750.0 ;
      RECT  94800.0 280650.0 95700.0 271350.0 ;
      RECT  92100.0 271350.0 93300.0 270150.0 ;
      RECT  94500.0 271350.0 95700.0 270150.0 ;
      RECT  94500.0 271350.0 95700.0 270150.0 ;
      RECT  92100.0 271350.0 93300.0 270150.0 ;
      RECT  92100.0 280650.0 93300.0 279450.0 ;
      RECT  94500.0 280650.0 95700.0 279450.0 ;
      RECT  94500.0 280650.0 95700.0 279450.0 ;
      RECT  92100.0 280650.0 93300.0 279450.0 ;
      RECT  96900.0 270750.0 98100.0 269550.0 ;
      RECT  96900.0 280650.0 98100.0 279450.0 ;
      RECT  92700.0 276000.0 93900.0 274800.0 ;
      RECT  92700.0 276000.0 93900.0 274800.0 ;
      RECT  95250.0 275850.0 96150.0 274950.0 ;
      RECT  90300.0 268650.0 99900.0 267750.0 ;
      RECT  90300.0 282450.0 99900.0 281550.0 ;
      RECT  96900.0 293850.0 98100.0 295800.0 ;
      RECT  96900.0 282000.0 98100.0 283950.0 ;
      RECT  92100.0 283350.0 93300.0 281550.0 ;
      RECT  92100.0 292650.0 93300.0 296250.0 ;
      RECT  94800.0 283350.0 95700.0 292650.0 ;
      RECT  92100.0 292650.0 93300.0 293850.0 ;
      RECT  94500.0 292650.0 95700.0 293850.0 ;
      RECT  94500.0 292650.0 95700.0 293850.0 ;
      RECT  92100.0 292650.0 93300.0 293850.0 ;
      RECT  92100.0 283350.0 93300.0 284550.0 ;
      RECT  94500.0 283350.0 95700.0 284550.0 ;
      RECT  94500.0 283350.0 95700.0 284550.0 ;
      RECT  92100.0 283350.0 93300.0 284550.0 ;
      RECT  96900.0 293250.0 98100.0 294450.0 ;
      RECT  96900.0 283350.0 98100.0 284550.0 ;
      RECT  92700.0 288000.0 93900.0 289200.0 ;
      RECT  92700.0 288000.0 93900.0 289200.0 ;
      RECT  95250.0 288150.0 96150.0 289050.0 ;
      RECT  90300.0 295350.0 99900.0 296250.0 ;
      RECT  90300.0 281550.0 99900.0 282450.0 ;
      RECT  96900.0 297750.0 98100.0 295800.0 ;
      RECT  96900.0 309600.0 98100.0 307650.0 ;
      RECT  92100.0 308250.0 93300.0 310050.0 ;
      RECT  92100.0 298950.0 93300.0 295350.0 ;
      RECT  94800.0 308250.0 95700.0 298950.0 ;
      RECT  92100.0 298950.0 93300.0 297750.0 ;
      RECT  94500.0 298950.0 95700.0 297750.0 ;
      RECT  94500.0 298950.0 95700.0 297750.0 ;
      RECT  92100.0 298950.0 93300.0 297750.0 ;
      RECT  92100.0 308250.0 93300.0 307050.0 ;
      RECT  94500.0 308250.0 95700.0 307050.0 ;
      RECT  94500.0 308250.0 95700.0 307050.0 ;
      RECT  92100.0 308250.0 93300.0 307050.0 ;
      RECT  96900.0 298350.0 98100.0 297150.0 ;
      RECT  96900.0 308250.0 98100.0 307050.0 ;
      RECT  92700.0 303600.0 93900.0 302400.0 ;
      RECT  92700.0 303600.0 93900.0 302400.0 ;
      RECT  95250.0 303450.0 96150.0 302550.0 ;
      RECT  90300.0 296250.0 99900.0 295350.0 ;
      RECT  90300.0 310050.0 99900.0 309150.0 ;
      RECT  96900.0 321450.0 98100.0 323400.0 ;
      RECT  96900.0 309600.0 98100.0 311550.0 ;
      RECT  92100.0 310950.0 93300.0 309150.0 ;
      RECT  92100.0 320250.0 93300.0 323850.0 ;
      RECT  94800.0 310950.0 95700.0 320250.0 ;
      RECT  92100.0 320250.0 93300.0 321450.0 ;
      RECT  94500.0 320250.0 95700.0 321450.0 ;
      RECT  94500.0 320250.0 95700.0 321450.0 ;
      RECT  92100.0 320250.0 93300.0 321450.0 ;
      RECT  92100.0 310950.0 93300.0 312150.0 ;
      RECT  94500.0 310950.0 95700.0 312150.0 ;
      RECT  94500.0 310950.0 95700.0 312150.0 ;
      RECT  92100.0 310950.0 93300.0 312150.0 ;
      RECT  96900.0 320850.0 98100.0 322050.0 ;
      RECT  96900.0 310950.0 98100.0 312150.0 ;
      RECT  92700.0 315600.0 93900.0 316800.0 ;
      RECT  92700.0 315600.0 93900.0 316800.0 ;
      RECT  95250.0 315750.0 96150.0 316650.0 ;
      RECT  90300.0 322950.0 99900.0 323850.0 ;
      RECT  90300.0 309150.0 99900.0 310050.0 ;
      RECT  96900.0 325350.0 98100.0 323400.0 ;
      RECT  96900.0 337200.0 98100.0 335250.0 ;
      RECT  92100.0 335850.0 93300.0 337650.0 ;
      RECT  92100.0 326550.0 93300.0 322950.0 ;
      RECT  94800.0 335850.0 95700.0 326550.0 ;
      RECT  92100.0 326550.0 93300.0 325350.0 ;
      RECT  94500.0 326550.0 95700.0 325350.0 ;
      RECT  94500.0 326550.0 95700.0 325350.0 ;
      RECT  92100.0 326550.0 93300.0 325350.0 ;
      RECT  92100.0 335850.0 93300.0 334650.0 ;
      RECT  94500.0 335850.0 95700.0 334650.0 ;
      RECT  94500.0 335850.0 95700.0 334650.0 ;
      RECT  92100.0 335850.0 93300.0 334650.0 ;
      RECT  96900.0 325950.0 98100.0 324750.0 ;
      RECT  96900.0 335850.0 98100.0 334650.0 ;
      RECT  92700.0 331200.0 93900.0 330000.0 ;
      RECT  92700.0 331200.0 93900.0 330000.0 ;
      RECT  95250.0 331050.0 96150.0 330150.0 ;
      RECT  90300.0 323850.0 99900.0 322950.0 ;
      RECT  90300.0 337650.0 99900.0 336750.0 ;
      RECT  96900.0 349050.0 98100.0 351000.0 ;
      RECT  96900.0 337200.0 98100.0 339150.0 ;
      RECT  92100.0 338550.0 93300.0 336750.0 ;
      RECT  92100.0 347850.0 93300.0 351450.0 ;
      RECT  94800.0 338550.0 95700.0 347850.0 ;
      RECT  92100.0 347850.0 93300.0 349050.0 ;
      RECT  94500.0 347850.0 95700.0 349050.0 ;
      RECT  94500.0 347850.0 95700.0 349050.0 ;
      RECT  92100.0 347850.0 93300.0 349050.0 ;
      RECT  92100.0 338550.0 93300.0 339750.0 ;
      RECT  94500.0 338550.0 95700.0 339750.0 ;
      RECT  94500.0 338550.0 95700.0 339750.0 ;
      RECT  92100.0 338550.0 93300.0 339750.0 ;
      RECT  96900.0 348450.0 98100.0 349650.0 ;
      RECT  96900.0 338550.0 98100.0 339750.0 ;
      RECT  92700.0 343200.0 93900.0 344400.0 ;
      RECT  92700.0 343200.0 93900.0 344400.0 ;
      RECT  95250.0 343350.0 96150.0 344250.0 ;
      RECT  90300.0 350550.0 99900.0 351450.0 ;
      RECT  90300.0 336750.0 99900.0 337650.0 ;
      RECT  96900.0 352950.0 98100.0 351000.0 ;
      RECT  96900.0 364800.0 98100.0 362850.0 ;
      RECT  92100.0 363450.0 93300.0 365250.0 ;
      RECT  92100.0 354150.0 93300.0 350550.0 ;
      RECT  94800.0 363450.0 95700.0 354150.0 ;
      RECT  92100.0 354150.0 93300.0 352950.0 ;
      RECT  94500.0 354150.0 95700.0 352950.0 ;
      RECT  94500.0 354150.0 95700.0 352950.0 ;
      RECT  92100.0 354150.0 93300.0 352950.0 ;
      RECT  92100.0 363450.0 93300.0 362250.0 ;
      RECT  94500.0 363450.0 95700.0 362250.0 ;
      RECT  94500.0 363450.0 95700.0 362250.0 ;
      RECT  92100.0 363450.0 93300.0 362250.0 ;
      RECT  96900.0 353550.0 98100.0 352350.0 ;
      RECT  96900.0 363450.0 98100.0 362250.0 ;
      RECT  92700.0 358800.0 93900.0 357600.0 ;
      RECT  92700.0 358800.0 93900.0 357600.0 ;
      RECT  95250.0 358650.0 96150.0 357750.0 ;
      RECT  90300.0 351450.0 99900.0 350550.0 ;
      RECT  90300.0 365250.0 99900.0 364350.0 ;
      RECT  96900.0 376650.0 98100.0 378600.0 ;
      RECT  96900.0 364800.0 98100.0 366750.0 ;
      RECT  92100.0 366150.0 93300.0 364350.0 ;
      RECT  92100.0 375450.0 93300.0 379050.0 ;
      RECT  94800.0 366150.0 95700.0 375450.0 ;
      RECT  92100.0 375450.0 93300.0 376650.0 ;
      RECT  94500.0 375450.0 95700.0 376650.0 ;
      RECT  94500.0 375450.0 95700.0 376650.0 ;
      RECT  92100.0 375450.0 93300.0 376650.0 ;
      RECT  92100.0 366150.0 93300.0 367350.0 ;
      RECT  94500.0 366150.0 95700.0 367350.0 ;
      RECT  94500.0 366150.0 95700.0 367350.0 ;
      RECT  92100.0 366150.0 93300.0 367350.0 ;
      RECT  96900.0 376050.0 98100.0 377250.0 ;
      RECT  96900.0 366150.0 98100.0 367350.0 ;
      RECT  92700.0 370800.0 93900.0 372000.0 ;
      RECT  92700.0 370800.0 93900.0 372000.0 ;
      RECT  95250.0 370950.0 96150.0 371850.0 ;
      RECT  90300.0 378150.0 99900.0 379050.0 ;
      RECT  90300.0 364350.0 99900.0 365250.0 ;
      RECT  96900.0 380550.0 98100.0 378600.0 ;
      RECT  96900.0 392400.0 98100.0 390450.0 ;
      RECT  92100.0 391050.0 93300.0 392850.0 ;
      RECT  92100.0 381750.0 93300.0 378150.0 ;
      RECT  94800.0 391050.0 95700.0 381750.0 ;
      RECT  92100.0 381750.0 93300.0 380550.0 ;
      RECT  94500.0 381750.0 95700.0 380550.0 ;
      RECT  94500.0 381750.0 95700.0 380550.0 ;
      RECT  92100.0 381750.0 93300.0 380550.0 ;
      RECT  92100.0 391050.0 93300.0 389850.0 ;
      RECT  94500.0 391050.0 95700.0 389850.0 ;
      RECT  94500.0 391050.0 95700.0 389850.0 ;
      RECT  92100.0 391050.0 93300.0 389850.0 ;
      RECT  96900.0 381150.0 98100.0 379950.0 ;
      RECT  96900.0 391050.0 98100.0 389850.0 ;
      RECT  92700.0 386400.0 93900.0 385200.0 ;
      RECT  92700.0 386400.0 93900.0 385200.0 ;
      RECT  95250.0 386250.0 96150.0 385350.0 ;
      RECT  90300.0 379050.0 99900.0 378150.0 ;
      RECT  90300.0 392850.0 99900.0 391950.0 ;
      RECT  96900.0 404250.0 98100.0 406200.0 ;
      RECT  96900.0 392400.0 98100.0 394350.0 ;
      RECT  92100.0 393750.0 93300.0 391950.0 ;
      RECT  92100.0 403050.0 93300.0 406650.0 ;
      RECT  94800.0 393750.0 95700.0 403050.0 ;
      RECT  92100.0 403050.0 93300.0 404250.0 ;
      RECT  94500.0 403050.0 95700.0 404250.0 ;
      RECT  94500.0 403050.0 95700.0 404250.0 ;
      RECT  92100.0 403050.0 93300.0 404250.0 ;
      RECT  92100.0 393750.0 93300.0 394950.0 ;
      RECT  94500.0 393750.0 95700.0 394950.0 ;
      RECT  94500.0 393750.0 95700.0 394950.0 ;
      RECT  92100.0 393750.0 93300.0 394950.0 ;
      RECT  96900.0 403650.0 98100.0 404850.0 ;
      RECT  96900.0 393750.0 98100.0 394950.0 ;
      RECT  92700.0 398400.0 93900.0 399600.0 ;
      RECT  92700.0 398400.0 93900.0 399600.0 ;
      RECT  95250.0 398550.0 96150.0 399450.0 ;
      RECT  90300.0 405750.0 99900.0 406650.0 ;
      RECT  90300.0 391950.0 99900.0 392850.0 ;
      RECT  96900.0 408150.0 98100.0 406200.0 ;
      RECT  96900.0 420000.0 98100.0 418050.0 ;
      RECT  92100.0 418650.0 93300.0 420450.0 ;
      RECT  92100.0 409350.0 93300.0 405750.0 ;
      RECT  94800.0 418650.0 95700.0 409350.0 ;
      RECT  92100.0 409350.0 93300.0 408150.0 ;
      RECT  94500.0 409350.0 95700.0 408150.0 ;
      RECT  94500.0 409350.0 95700.0 408150.0 ;
      RECT  92100.0 409350.0 93300.0 408150.0 ;
      RECT  92100.0 418650.0 93300.0 417450.0 ;
      RECT  94500.0 418650.0 95700.0 417450.0 ;
      RECT  94500.0 418650.0 95700.0 417450.0 ;
      RECT  92100.0 418650.0 93300.0 417450.0 ;
      RECT  96900.0 408750.0 98100.0 407550.0 ;
      RECT  96900.0 418650.0 98100.0 417450.0 ;
      RECT  92700.0 414000.0 93900.0 412800.0 ;
      RECT  92700.0 414000.0 93900.0 412800.0 ;
      RECT  95250.0 413850.0 96150.0 412950.0 ;
      RECT  90300.0 406650.0 99900.0 405750.0 ;
      RECT  90300.0 420450.0 99900.0 419550.0 ;
      RECT  60150.0 94800.0 58950.0 96000.0 ;
      RECT  62250.0 109200.0 61050.0 110400.0 ;
      RECT  64350.0 122400.0 63150.0 123600.0 ;
      RECT  66450.0 136800.0 65250.0 138000.0 ;
      RECT  68550.0 150000.0 67350.0 151200.0 ;
      RECT  70650.0 164400.0 69450.0 165600.0 ;
      RECT  72750.0 177600.0 71550.0 178800.0 ;
      RECT  74850.0 192000.0 73650.0 193200.0 ;
      RECT  60150.0 206400.0 58950.0 207600.0 ;
      RECT  68550.0 203700.0 67350.0 204900.0 ;
      RECT  60150.0 218400.0 58950.0 219600.0 ;
      RECT  70650.0 221100.0 69450.0 222300.0 ;
      RECT  60150.0 234000.0 58950.0 235200.0 ;
      RECT  72750.0 231300.0 71550.0 232500.0 ;
      RECT  60150.0 246000.0 58950.0 247200.0 ;
      RECT  74850.0 248700.0 73650.0 249900.0 ;
      RECT  62250.0 261600.0 61050.0 262800.0 ;
      RECT  68550.0 258900.0 67350.0 260100.0 ;
      RECT  62250.0 273600.0 61050.0 274800.0 ;
      RECT  70650.0 276300.0 69450.0 277500.0 ;
      RECT  62250.0 289200.0 61050.0 290400.0 ;
      RECT  72750.0 286500.0 71550.0 287700.0 ;
      RECT  62250.0 301200.0 61050.0 302400.0 ;
      RECT  74850.0 303900.0 73650.0 305100.0 ;
      RECT  64350.0 316800.0 63150.0 318000.0 ;
      RECT  68550.0 314100.0 67350.0 315300.0 ;
      RECT  64350.0 328800.0 63150.0 330000.0 ;
      RECT  70650.0 331500.0 69450.0 332700.0 ;
      RECT  64350.0 344400.0 63150.0 345600.0 ;
      RECT  72750.0 341700.0 71550.0 342900.0 ;
      RECT  64350.0 356400.0 63150.0 357600.0 ;
      RECT  74850.0 359100.0 73650.0 360300.0 ;
      RECT  66450.0 372000.0 65250.0 373200.0 ;
      RECT  68550.0 369300.0 67350.0 370500.0 ;
      RECT  66450.0 384000.0 65250.0 385200.0 ;
      RECT  70650.0 386700.0 69450.0 387900.0 ;
      RECT  66450.0 399600.0 65250.0 400800.0 ;
      RECT  72750.0 396900.0 71550.0 398100.0 ;
      RECT  66450.0 411600.0 65250.0 412800.0 ;
      RECT  74850.0 414300.0 73650.0 415500.0 ;
      RECT  95250.0 205350.0 96150.0 206250.0 ;
      RECT  95250.0 219750.0 96150.0 220650.0 ;
      RECT  95250.0 232950.0 96150.0 233850.0 ;
      RECT  95250.0 247350.0 96150.0 248250.0 ;
      RECT  95250.0 260550.0 96150.0 261450.0 ;
      RECT  95250.0 274950.0 96150.0 275850.0 ;
      RECT  95250.0 288150.0 96150.0 289050.0 ;
      RECT  95250.0 302550.0 96150.0 303450.0 ;
      RECT  95250.0 315750.0 96150.0 316650.0 ;
      RECT  95250.0 330150.0 96150.0 331050.0 ;
      RECT  95250.0 343350.0 96150.0 344250.0 ;
      RECT  95250.0 357750.0 96150.0 358650.0 ;
      RECT  95250.0 370950.0 96150.0 371850.0 ;
      RECT  95250.0 385350.0 96150.0 386250.0 ;
      RECT  95250.0 398550.0 96150.0 399450.0 ;
      RECT  95250.0 412950.0 96150.0 413850.0 ;
      RECT  59100.0 102150.0 130500.0 103050.0 ;
      RECT  59100.0 129750.0 130500.0 130650.0 ;
      RECT  59100.0 157350.0 130500.0 158250.0 ;
      RECT  59100.0 184950.0 130500.0 185850.0 ;
      RECT  59100.0 212550.0 130500.0 213450.0 ;
      RECT  59100.0 240150.0 130500.0 241050.0 ;
      RECT  59100.0 267750.0 130500.0 268650.0 ;
      RECT  59100.0 295350.0 130500.0 296250.0 ;
      RECT  59100.0 322950.0 130500.0 323850.0 ;
      RECT  59100.0 350550.0 130500.0 351450.0 ;
      RECT  59100.0 378150.0 130500.0 379050.0 ;
      RECT  59100.0 405750.0 130500.0 406650.0 ;
      RECT  59100.0 88350.0 130500.0 89250.0 ;
      RECT  59100.0 115950.0 130500.0 116850.0 ;
      RECT  59100.0 143550.0 130500.0 144450.0 ;
      RECT  59100.0 171150.0 130500.0 172050.0 ;
      RECT  59100.0 198750.0 130500.0 199650.0 ;
      RECT  59100.0 226350.0 130500.0 227250.0 ;
      RECT  59100.0 253950.0 130500.0 254850.0 ;
      RECT  59100.0 281550.0 130500.0 282450.0 ;
      RECT  59100.0 309150.0 130500.0 310050.0 ;
      RECT  59100.0 336750.0 130500.0 337650.0 ;
      RECT  59100.0 364350.0 130500.0 365250.0 ;
      RECT  59100.0 391950.0 130500.0 392850.0 ;
      RECT  59100.0 419550.0 130500.0 420450.0 ;
      RECT  103050.0 205350.0 108600.0 206250.0 ;
      RECT  111150.0 206550.0 112050.0 207450.0 ;
      RECT  111150.0 205350.0 112050.0 206250.0 ;
      RECT  111150.0 206250.0 112050.0 207000.0 ;
      RECT  111600.0 206550.0 118200.0 207450.0 ;
      RECT  118200.0 206550.0 119400.0 207450.0 ;
      RECT  127650.0 206550.0 128550.0 207450.0 ;
      RECT  127650.0 205350.0 128550.0 206250.0 ;
      RECT  123600.0 206550.0 128100.0 207450.0 ;
      RECT  127650.0 205800.0 128550.0 207000.0 ;
      RECT  128100.0 205350.0 132600.0 206250.0 ;
      RECT  103050.0 219750.0 108600.0 220650.0 ;
      RECT  111150.0 218550.0 112050.0 219450.0 ;
      RECT  111150.0 219750.0 112050.0 220650.0 ;
      RECT  111150.0 219000.0 112050.0 220650.0 ;
      RECT  111600.0 218550.0 118200.0 219450.0 ;
      RECT  118200.0 218550.0 119400.0 219450.0 ;
      RECT  127650.0 218550.0 128550.0 219450.0 ;
      RECT  127650.0 219750.0 128550.0 220650.0 ;
      RECT  123600.0 218550.0 128100.0 219450.0 ;
      RECT  127650.0 219000.0 128550.0 220200.0 ;
      RECT  128100.0 219750.0 132600.0 220650.0 ;
      RECT  103050.0 232950.0 108600.0 233850.0 ;
      RECT  111150.0 234150.0 112050.0 235050.0 ;
      RECT  111150.0 232950.0 112050.0 233850.0 ;
      RECT  111150.0 233850.0 112050.0 234600.0 ;
      RECT  111600.0 234150.0 118200.0 235050.0 ;
      RECT  118200.0 234150.0 119400.0 235050.0 ;
      RECT  127650.0 234150.0 128550.0 235050.0 ;
      RECT  127650.0 232950.0 128550.0 233850.0 ;
      RECT  123600.0 234150.0 128100.0 235050.0 ;
      RECT  127650.0 233400.0 128550.0 234600.0 ;
      RECT  128100.0 232950.0 132600.0 233850.0 ;
      RECT  103050.0 247350.0 108600.0 248250.0 ;
      RECT  111150.0 246150.0 112050.0 247050.0 ;
      RECT  111150.0 247350.0 112050.0 248250.0 ;
      RECT  111150.0 246600.0 112050.0 248250.0 ;
      RECT  111600.0 246150.0 118200.0 247050.0 ;
      RECT  118200.0 246150.0 119400.0 247050.0 ;
      RECT  127650.0 246150.0 128550.0 247050.0 ;
      RECT  127650.0 247350.0 128550.0 248250.0 ;
      RECT  123600.0 246150.0 128100.0 247050.0 ;
      RECT  127650.0 246600.0 128550.0 247800.0 ;
      RECT  128100.0 247350.0 132600.0 248250.0 ;
      RECT  103050.0 260550.0 108600.0 261450.0 ;
      RECT  111150.0 261750.0 112050.0 262650.0 ;
      RECT  111150.0 260550.0 112050.0 261450.0 ;
      RECT  111150.0 261450.0 112050.0 262200.0 ;
      RECT  111600.0 261750.0 118200.0 262650.0 ;
      RECT  118200.0 261750.0 119400.0 262650.0 ;
      RECT  127650.0 261750.0 128550.0 262650.0 ;
      RECT  127650.0 260550.0 128550.0 261450.0 ;
      RECT  123600.0 261750.0 128100.0 262650.0 ;
      RECT  127650.0 261000.0 128550.0 262200.0 ;
      RECT  128100.0 260550.0 132600.0 261450.0 ;
      RECT  103050.0 274950.0 108600.0 275850.0 ;
      RECT  111150.0 273750.0 112050.0 274650.0 ;
      RECT  111150.0 274950.0 112050.0 275850.0 ;
      RECT  111150.0 274200.0 112050.0 275850.0 ;
      RECT  111600.0 273750.0 118200.0 274650.0 ;
      RECT  118200.0 273750.0 119400.0 274650.0 ;
      RECT  127650.0 273750.0 128550.0 274650.0 ;
      RECT  127650.0 274950.0 128550.0 275850.0 ;
      RECT  123600.0 273750.0 128100.0 274650.0 ;
      RECT  127650.0 274200.0 128550.0 275400.0 ;
      RECT  128100.0 274950.0 132600.0 275850.0 ;
      RECT  103050.0 288150.0 108600.0 289050.0 ;
      RECT  111150.0 289350.0 112050.0 290250.0 ;
      RECT  111150.0 288150.0 112050.0 289050.0 ;
      RECT  111150.0 289050.0 112050.0 289800.0 ;
      RECT  111600.0 289350.0 118200.0 290250.0 ;
      RECT  118200.0 289350.0 119400.0 290250.0 ;
      RECT  127650.0 289350.0 128550.0 290250.0 ;
      RECT  127650.0 288150.0 128550.0 289050.0 ;
      RECT  123600.0 289350.0 128100.0 290250.0 ;
      RECT  127650.0 288600.0 128550.0 289800.0 ;
      RECT  128100.0 288150.0 132600.0 289050.0 ;
      RECT  103050.0 302550.0 108600.0 303450.0 ;
      RECT  111150.0 301350.0 112050.0 302250.0 ;
      RECT  111150.0 302550.0 112050.0 303450.0 ;
      RECT  111150.0 301800.0 112050.0 303450.0 ;
      RECT  111600.0 301350.0 118200.0 302250.0 ;
      RECT  118200.0 301350.0 119400.0 302250.0 ;
      RECT  127650.0 301350.0 128550.0 302250.0 ;
      RECT  127650.0 302550.0 128550.0 303450.0 ;
      RECT  123600.0 301350.0 128100.0 302250.0 ;
      RECT  127650.0 301800.0 128550.0 303000.0 ;
      RECT  128100.0 302550.0 132600.0 303450.0 ;
      RECT  103050.0 315750.0 108600.0 316650.0 ;
      RECT  111150.0 316950.0 112050.0 317850.0 ;
      RECT  111150.0 315750.0 112050.0 316650.0 ;
      RECT  111150.0 316650.0 112050.0 317400.0 ;
      RECT  111600.0 316950.0 118200.0 317850.0 ;
      RECT  118200.0 316950.0 119400.0 317850.0 ;
      RECT  127650.0 316950.0 128550.0 317850.0 ;
      RECT  127650.0 315750.0 128550.0 316650.0 ;
      RECT  123600.0 316950.0 128100.0 317850.0 ;
      RECT  127650.0 316200.0 128550.0 317400.0 ;
      RECT  128100.0 315750.0 132600.0 316650.0 ;
      RECT  103050.0 330150.0 108600.0 331050.0 ;
      RECT  111150.0 328950.0 112050.0 329850.0 ;
      RECT  111150.0 330150.0 112050.0 331050.0 ;
      RECT  111150.0 329400.0 112050.0 331050.0 ;
      RECT  111600.0 328950.0 118200.0 329850.0 ;
      RECT  118200.0 328950.0 119400.0 329850.0 ;
      RECT  127650.0 328950.0 128550.0 329850.0 ;
      RECT  127650.0 330150.0 128550.0 331050.0 ;
      RECT  123600.0 328950.0 128100.0 329850.0 ;
      RECT  127650.0 329400.0 128550.0 330600.0 ;
      RECT  128100.0 330150.0 132600.0 331050.0 ;
      RECT  103050.0 343350.0 108600.0 344250.0 ;
      RECT  111150.0 344550.0 112050.0 345450.0 ;
      RECT  111150.0 343350.0 112050.0 344250.0 ;
      RECT  111150.0 344250.0 112050.0 345000.0 ;
      RECT  111600.0 344550.0 118200.0 345450.0 ;
      RECT  118200.0 344550.0 119400.0 345450.0 ;
      RECT  127650.0 344550.0 128550.0 345450.0 ;
      RECT  127650.0 343350.0 128550.0 344250.0 ;
      RECT  123600.0 344550.0 128100.0 345450.0 ;
      RECT  127650.0 343800.0 128550.0 345000.0 ;
      RECT  128100.0 343350.0 132600.0 344250.0 ;
      RECT  103050.0 357750.0 108600.0 358650.0 ;
      RECT  111150.0 356550.0 112050.0 357450.0 ;
      RECT  111150.0 357750.0 112050.0 358650.0 ;
      RECT  111150.0 357000.0 112050.0 358650.0 ;
      RECT  111600.0 356550.0 118200.0 357450.0 ;
      RECT  118200.0 356550.0 119400.0 357450.0 ;
      RECT  127650.0 356550.0 128550.0 357450.0 ;
      RECT  127650.0 357750.0 128550.0 358650.0 ;
      RECT  123600.0 356550.0 128100.0 357450.0 ;
      RECT  127650.0 357000.0 128550.0 358200.0 ;
      RECT  128100.0 357750.0 132600.0 358650.0 ;
      RECT  103050.0 370950.0 108600.0 371850.0 ;
      RECT  111150.0 372150.0 112050.0 373050.0 ;
      RECT  111150.0 370950.0 112050.0 371850.0 ;
      RECT  111150.0 371850.0 112050.0 372600.0 ;
      RECT  111600.0 372150.0 118200.0 373050.0 ;
      RECT  118200.0 372150.0 119400.0 373050.0 ;
      RECT  127650.0 372150.0 128550.0 373050.0 ;
      RECT  127650.0 370950.0 128550.0 371850.0 ;
      RECT  123600.0 372150.0 128100.0 373050.0 ;
      RECT  127650.0 371400.0 128550.0 372600.0 ;
      RECT  128100.0 370950.0 132600.0 371850.0 ;
      RECT  103050.0 385350.0 108600.0 386250.0 ;
      RECT  111150.0 384150.0 112050.0 385050.0 ;
      RECT  111150.0 385350.0 112050.0 386250.0 ;
      RECT  111150.0 384600.0 112050.0 386250.0 ;
      RECT  111600.0 384150.0 118200.0 385050.0 ;
      RECT  118200.0 384150.0 119400.0 385050.0 ;
      RECT  127650.0 384150.0 128550.0 385050.0 ;
      RECT  127650.0 385350.0 128550.0 386250.0 ;
      RECT  123600.0 384150.0 128100.0 385050.0 ;
      RECT  127650.0 384600.0 128550.0 385800.0 ;
      RECT  128100.0 385350.0 132600.0 386250.0 ;
      RECT  103050.0 398550.0 108600.0 399450.0 ;
      RECT  111150.0 399750.0 112050.0 400650.0 ;
      RECT  111150.0 398550.0 112050.0 399450.0 ;
      RECT  111150.0 399450.0 112050.0 400200.0 ;
      RECT  111600.0 399750.0 118200.0 400650.0 ;
      RECT  118200.0 399750.0 119400.0 400650.0 ;
      RECT  127650.0 399750.0 128550.0 400650.0 ;
      RECT  127650.0 398550.0 128550.0 399450.0 ;
      RECT  123600.0 399750.0 128100.0 400650.0 ;
      RECT  127650.0 399000.0 128550.0 400200.0 ;
      RECT  128100.0 398550.0 132600.0 399450.0 ;
      RECT  103050.0 412950.0 108600.0 413850.0 ;
      RECT  111150.0 411750.0 112050.0 412650.0 ;
      RECT  111150.0 412950.0 112050.0 413850.0 ;
      RECT  111150.0 412200.0 112050.0 413850.0 ;
      RECT  111600.0 411750.0 118200.0 412650.0 ;
      RECT  118200.0 411750.0 119400.0 412650.0 ;
      RECT  127650.0 411750.0 128550.0 412650.0 ;
      RECT  127650.0 412950.0 128550.0 413850.0 ;
      RECT  123600.0 411750.0 128100.0 412650.0 ;
      RECT  127650.0 412200.0 128550.0 413400.0 ;
      RECT  128100.0 412950.0 132600.0 413850.0 ;
      RECT  112800.0 211050.0 114000.0 213000.0 ;
      RECT  112800.0 199200.0 114000.0 201150.0 ;
      RECT  108000.0 200550.0 109200.0 198750.0 ;
      RECT  108000.0 209850.0 109200.0 213450.0 ;
      RECT  110700.0 200550.0 111600.0 209850.0 ;
      RECT  108000.0 209850.0 109200.0 211050.0 ;
      RECT  110400.0 209850.0 111600.0 211050.0 ;
      RECT  110400.0 209850.0 111600.0 211050.0 ;
      RECT  108000.0 209850.0 109200.0 211050.0 ;
      RECT  108000.0 200550.0 109200.0 201750.0 ;
      RECT  110400.0 200550.0 111600.0 201750.0 ;
      RECT  110400.0 200550.0 111600.0 201750.0 ;
      RECT  108000.0 200550.0 109200.0 201750.0 ;
      RECT  112800.0 210450.0 114000.0 211650.0 ;
      RECT  112800.0 200550.0 114000.0 201750.0 ;
      RECT  108600.0 205200.0 109800.0 206400.0 ;
      RECT  108600.0 205200.0 109800.0 206400.0 ;
      RECT  111150.0 205350.0 112050.0 206250.0 ;
      RECT  106200.0 212550.0 115800.0 213450.0 ;
      RECT  106200.0 198750.0 115800.0 199650.0 ;
      RECT  117600.0 201150.0 118800.0 198750.0 ;
      RECT  117600.0 209850.0 118800.0 213450.0 ;
      RECT  122400.0 209850.0 123600.0 213450.0 ;
      RECT  124800.0 211050.0 126000.0 213000.0 ;
      RECT  124800.0 199200.0 126000.0 201150.0 ;
      RECT  117600.0 209850.0 118800.0 211050.0 ;
      RECT  120000.0 209850.0 121200.0 211050.0 ;
      RECT  120000.0 209850.0 121200.0 211050.0 ;
      RECT  117600.0 209850.0 118800.0 211050.0 ;
      RECT  120000.0 209850.0 121200.0 211050.0 ;
      RECT  122400.0 209850.0 123600.0 211050.0 ;
      RECT  122400.0 209850.0 123600.0 211050.0 ;
      RECT  120000.0 209850.0 121200.0 211050.0 ;
      RECT  117600.0 201150.0 118800.0 202350.0 ;
      RECT  120000.0 201150.0 121200.0 202350.0 ;
      RECT  120000.0 201150.0 121200.0 202350.0 ;
      RECT  117600.0 201150.0 118800.0 202350.0 ;
      RECT  120000.0 201150.0 121200.0 202350.0 ;
      RECT  122400.0 201150.0 123600.0 202350.0 ;
      RECT  122400.0 201150.0 123600.0 202350.0 ;
      RECT  120000.0 201150.0 121200.0 202350.0 ;
      RECT  124800.0 210450.0 126000.0 211650.0 ;
      RECT  124800.0 200550.0 126000.0 201750.0 ;
      RECT  122400.0 203700.0 121200.0 204900.0 ;
      RECT  119400.0 206400.0 118200.0 207600.0 ;
      RECT  120000.0 209850.0 121200.0 211050.0 ;
      RECT  122400.0 201150.0 123600.0 202350.0 ;
      RECT  123600.0 206400.0 122400.0 207600.0 ;
      RECT  118200.0 206400.0 119400.0 207600.0 ;
      RECT  121200.0 203700.0 122400.0 204900.0 ;
      RECT  122400.0 206400.0 123600.0 207600.0 ;
      RECT  115800.0 212550.0 130200.0 213450.0 ;
      RECT  115800.0 198750.0 130200.0 199650.0 ;
      RECT  136800.0 211050.0 138000.0 213000.0 ;
      RECT  136800.0 199200.0 138000.0 201150.0 ;
      RECT  132000.0 200550.0 133200.0 198750.0 ;
      RECT  132000.0 209850.0 133200.0 213450.0 ;
      RECT  134700.0 200550.0 135600.0 209850.0 ;
      RECT  132000.0 209850.0 133200.0 211050.0 ;
      RECT  134400.0 209850.0 135600.0 211050.0 ;
      RECT  134400.0 209850.0 135600.0 211050.0 ;
      RECT  132000.0 209850.0 133200.0 211050.0 ;
      RECT  132000.0 200550.0 133200.0 201750.0 ;
      RECT  134400.0 200550.0 135600.0 201750.0 ;
      RECT  134400.0 200550.0 135600.0 201750.0 ;
      RECT  132000.0 200550.0 133200.0 201750.0 ;
      RECT  136800.0 210450.0 138000.0 211650.0 ;
      RECT  136800.0 200550.0 138000.0 201750.0 ;
      RECT  132600.0 205200.0 133800.0 206400.0 ;
      RECT  132600.0 205200.0 133800.0 206400.0 ;
      RECT  135150.0 205350.0 136050.0 206250.0 ;
      RECT  130200.0 212550.0 139800.0 213450.0 ;
      RECT  130200.0 198750.0 139800.0 199650.0 ;
      RECT  102450.0 205200.0 103650.0 206400.0 ;
      RECT  104400.0 202800.0 105600.0 204000.0 ;
      RECT  121200.0 203700.0 120000.0 204900.0 ;
      RECT  112800.0 214950.0 114000.0 213000.0 ;
      RECT  112800.0 226800.0 114000.0 224850.0 ;
      RECT  108000.0 225450.0 109200.0 227250.0 ;
      RECT  108000.0 216150.0 109200.0 212550.0 ;
      RECT  110700.0 225450.0 111600.0 216150.0 ;
      RECT  108000.0 216150.0 109200.0 214950.0 ;
      RECT  110400.0 216150.0 111600.0 214950.0 ;
      RECT  110400.0 216150.0 111600.0 214950.0 ;
      RECT  108000.0 216150.0 109200.0 214950.0 ;
      RECT  108000.0 225450.0 109200.0 224250.0 ;
      RECT  110400.0 225450.0 111600.0 224250.0 ;
      RECT  110400.0 225450.0 111600.0 224250.0 ;
      RECT  108000.0 225450.0 109200.0 224250.0 ;
      RECT  112800.0 215550.0 114000.0 214350.0 ;
      RECT  112800.0 225450.0 114000.0 224250.0 ;
      RECT  108600.0 220800.0 109800.0 219600.0 ;
      RECT  108600.0 220800.0 109800.0 219600.0 ;
      RECT  111150.0 220650.0 112050.0 219750.0 ;
      RECT  106200.0 213450.0 115800.0 212550.0 ;
      RECT  106200.0 227250.0 115800.0 226350.0 ;
      RECT  117600.0 224850.0 118800.0 227250.0 ;
      RECT  117600.0 216150.0 118800.0 212550.0 ;
      RECT  122400.0 216150.0 123600.0 212550.0 ;
      RECT  124800.0 214950.0 126000.0 213000.0 ;
      RECT  124800.0 226800.0 126000.0 224850.0 ;
      RECT  117600.0 216150.0 118800.0 214950.0 ;
      RECT  120000.0 216150.0 121200.0 214950.0 ;
      RECT  120000.0 216150.0 121200.0 214950.0 ;
      RECT  117600.0 216150.0 118800.0 214950.0 ;
      RECT  120000.0 216150.0 121200.0 214950.0 ;
      RECT  122400.0 216150.0 123600.0 214950.0 ;
      RECT  122400.0 216150.0 123600.0 214950.0 ;
      RECT  120000.0 216150.0 121200.0 214950.0 ;
      RECT  117600.0 224850.0 118800.0 223650.0 ;
      RECT  120000.0 224850.0 121200.0 223650.0 ;
      RECT  120000.0 224850.0 121200.0 223650.0 ;
      RECT  117600.0 224850.0 118800.0 223650.0 ;
      RECT  120000.0 224850.0 121200.0 223650.0 ;
      RECT  122400.0 224850.0 123600.0 223650.0 ;
      RECT  122400.0 224850.0 123600.0 223650.0 ;
      RECT  120000.0 224850.0 121200.0 223650.0 ;
      RECT  124800.0 215550.0 126000.0 214350.0 ;
      RECT  124800.0 225450.0 126000.0 224250.0 ;
      RECT  122400.0 222300.0 121200.0 221100.0 ;
      RECT  119400.0 219600.0 118200.0 218400.0 ;
      RECT  120000.0 216150.0 121200.0 214950.0 ;
      RECT  122400.0 224850.0 123600.0 223650.0 ;
      RECT  123600.0 219600.0 122400.0 218400.0 ;
      RECT  118200.0 219600.0 119400.0 218400.0 ;
      RECT  121200.0 222300.0 122400.0 221100.0 ;
      RECT  122400.0 219600.0 123600.0 218400.0 ;
      RECT  115800.0 213450.0 130200.0 212550.0 ;
      RECT  115800.0 227250.0 130200.0 226350.0 ;
      RECT  136800.0 214950.0 138000.0 213000.0 ;
      RECT  136800.0 226800.0 138000.0 224850.0 ;
      RECT  132000.0 225450.0 133200.0 227250.0 ;
      RECT  132000.0 216150.0 133200.0 212550.0 ;
      RECT  134700.0 225450.0 135600.0 216150.0 ;
      RECT  132000.0 216150.0 133200.0 214950.0 ;
      RECT  134400.0 216150.0 135600.0 214950.0 ;
      RECT  134400.0 216150.0 135600.0 214950.0 ;
      RECT  132000.0 216150.0 133200.0 214950.0 ;
      RECT  132000.0 225450.0 133200.0 224250.0 ;
      RECT  134400.0 225450.0 135600.0 224250.0 ;
      RECT  134400.0 225450.0 135600.0 224250.0 ;
      RECT  132000.0 225450.0 133200.0 224250.0 ;
      RECT  136800.0 215550.0 138000.0 214350.0 ;
      RECT  136800.0 225450.0 138000.0 224250.0 ;
      RECT  132600.0 220800.0 133800.0 219600.0 ;
      RECT  132600.0 220800.0 133800.0 219600.0 ;
      RECT  135150.0 220650.0 136050.0 219750.0 ;
      RECT  130200.0 213450.0 139800.0 212550.0 ;
      RECT  130200.0 227250.0 139800.0 226350.0 ;
      RECT  102450.0 219600.0 103650.0 220800.0 ;
      RECT  104400.0 222000.0 105600.0 223200.0 ;
      RECT  121200.0 221100.0 120000.0 222300.0 ;
      RECT  112800.0 238650.0 114000.0 240600.0 ;
      RECT  112800.0 226800.0 114000.0 228750.0 ;
      RECT  108000.0 228150.0 109200.0 226350.0 ;
      RECT  108000.0 237450.0 109200.0 241050.0 ;
      RECT  110700.0 228150.0 111600.0 237450.0 ;
      RECT  108000.0 237450.0 109200.0 238650.0 ;
      RECT  110400.0 237450.0 111600.0 238650.0 ;
      RECT  110400.0 237450.0 111600.0 238650.0 ;
      RECT  108000.0 237450.0 109200.0 238650.0 ;
      RECT  108000.0 228150.0 109200.0 229350.0 ;
      RECT  110400.0 228150.0 111600.0 229350.0 ;
      RECT  110400.0 228150.0 111600.0 229350.0 ;
      RECT  108000.0 228150.0 109200.0 229350.0 ;
      RECT  112800.0 238050.0 114000.0 239250.0 ;
      RECT  112800.0 228150.0 114000.0 229350.0 ;
      RECT  108600.0 232800.0 109800.0 234000.0 ;
      RECT  108600.0 232800.0 109800.0 234000.0 ;
      RECT  111150.0 232950.0 112050.0 233850.0 ;
      RECT  106200.0 240150.0 115800.0 241050.0 ;
      RECT  106200.0 226350.0 115800.0 227250.0 ;
      RECT  117600.0 228750.0 118800.0 226350.0 ;
      RECT  117600.0 237450.0 118800.0 241050.0 ;
      RECT  122400.0 237450.0 123600.0 241050.0 ;
      RECT  124800.0 238650.0 126000.0 240600.0 ;
      RECT  124800.0 226800.0 126000.0 228750.0 ;
      RECT  117600.0 237450.0 118800.0 238650.0 ;
      RECT  120000.0 237450.0 121200.0 238650.0 ;
      RECT  120000.0 237450.0 121200.0 238650.0 ;
      RECT  117600.0 237450.0 118800.0 238650.0 ;
      RECT  120000.0 237450.0 121200.0 238650.0 ;
      RECT  122400.0 237450.0 123600.0 238650.0 ;
      RECT  122400.0 237450.0 123600.0 238650.0 ;
      RECT  120000.0 237450.0 121200.0 238650.0 ;
      RECT  117600.0 228750.0 118800.0 229950.0 ;
      RECT  120000.0 228750.0 121200.0 229950.0 ;
      RECT  120000.0 228750.0 121200.0 229950.0 ;
      RECT  117600.0 228750.0 118800.0 229950.0 ;
      RECT  120000.0 228750.0 121200.0 229950.0 ;
      RECT  122400.0 228750.0 123600.0 229950.0 ;
      RECT  122400.0 228750.0 123600.0 229950.0 ;
      RECT  120000.0 228750.0 121200.0 229950.0 ;
      RECT  124800.0 238050.0 126000.0 239250.0 ;
      RECT  124800.0 228150.0 126000.0 229350.0 ;
      RECT  122400.0 231300.0 121200.0 232500.0 ;
      RECT  119400.0 234000.0 118200.0 235200.0 ;
      RECT  120000.0 237450.0 121200.0 238650.0 ;
      RECT  122400.0 228750.0 123600.0 229950.0 ;
      RECT  123600.0 234000.0 122400.0 235200.0 ;
      RECT  118200.0 234000.0 119400.0 235200.0 ;
      RECT  121200.0 231300.0 122400.0 232500.0 ;
      RECT  122400.0 234000.0 123600.0 235200.0 ;
      RECT  115800.0 240150.0 130200.0 241050.0 ;
      RECT  115800.0 226350.0 130200.0 227250.0 ;
      RECT  136800.0 238650.0 138000.0 240600.0 ;
      RECT  136800.0 226800.0 138000.0 228750.0 ;
      RECT  132000.0 228150.0 133200.0 226350.0 ;
      RECT  132000.0 237450.0 133200.0 241050.0 ;
      RECT  134700.0 228150.0 135600.0 237450.0 ;
      RECT  132000.0 237450.0 133200.0 238650.0 ;
      RECT  134400.0 237450.0 135600.0 238650.0 ;
      RECT  134400.0 237450.0 135600.0 238650.0 ;
      RECT  132000.0 237450.0 133200.0 238650.0 ;
      RECT  132000.0 228150.0 133200.0 229350.0 ;
      RECT  134400.0 228150.0 135600.0 229350.0 ;
      RECT  134400.0 228150.0 135600.0 229350.0 ;
      RECT  132000.0 228150.0 133200.0 229350.0 ;
      RECT  136800.0 238050.0 138000.0 239250.0 ;
      RECT  136800.0 228150.0 138000.0 229350.0 ;
      RECT  132600.0 232800.0 133800.0 234000.0 ;
      RECT  132600.0 232800.0 133800.0 234000.0 ;
      RECT  135150.0 232950.0 136050.0 233850.0 ;
      RECT  130200.0 240150.0 139800.0 241050.0 ;
      RECT  130200.0 226350.0 139800.0 227250.0 ;
      RECT  102450.0 232800.0 103650.0 234000.0 ;
      RECT  104400.0 230400.0 105600.0 231600.0 ;
      RECT  121200.0 231300.0 120000.0 232500.0 ;
      RECT  112800.0 242550.0 114000.0 240600.0 ;
      RECT  112800.0 254400.0 114000.0 252450.0 ;
      RECT  108000.0 253050.0 109200.0 254850.0 ;
      RECT  108000.0 243750.0 109200.0 240150.0 ;
      RECT  110700.0 253050.0 111600.0 243750.0 ;
      RECT  108000.0 243750.0 109200.0 242550.0 ;
      RECT  110400.0 243750.0 111600.0 242550.0 ;
      RECT  110400.0 243750.0 111600.0 242550.0 ;
      RECT  108000.0 243750.0 109200.0 242550.0 ;
      RECT  108000.0 253050.0 109200.0 251850.0 ;
      RECT  110400.0 253050.0 111600.0 251850.0 ;
      RECT  110400.0 253050.0 111600.0 251850.0 ;
      RECT  108000.0 253050.0 109200.0 251850.0 ;
      RECT  112800.0 243150.0 114000.0 241950.0 ;
      RECT  112800.0 253050.0 114000.0 251850.0 ;
      RECT  108600.0 248400.0 109800.0 247200.0 ;
      RECT  108600.0 248400.0 109800.0 247200.0 ;
      RECT  111150.0 248250.0 112050.0 247350.0 ;
      RECT  106200.0 241050.0 115800.0 240150.0 ;
      RECT  106200.0 254850.0 115800.0 253950.0 ;
      RECT  117600.0 252450.0 118800.0 254850.0 ;
      RECT  117600.0 243750.0 118800.0 240150.0 ;
      RECT  122400.0 243750.0 123600.0 240150.0 ;
      RECT  124800.0 242550.0 126000.0 240600.0 ;
      RECT  124800.0 254400.0 126000.0 252450.0 ;
      RECT  117600.0 243750.0 118800.0 242550.0 ;
      RECT  120000.0 243750.0 121200.0 242550.0 ;
      RECT  120000.0 243750.0 121200.0 242550.0 ;
      RECT  117600.0 243750.0 118800.0 242550.0 ;
      RECT  120000.0 243750.0 121200.0 242550.0 ;
      RECT  122400.0 243750.0 123600.0 242550.0 ;
      RECT  122400.0 243750.0 123600.0 242550.0 ;
      RECT  120000.0 243750.0 121200.0 242550.0 ;
      RECT  117600.0 252450.0 118800.0 251250.0 ;
      RECT  120000.0 252450.0 121200.0 251250.0 ;
      RECT  120000.0 252450.0 121200.0 251250.0 ;
      RECT  117600.0 252450.0 118800.0 251250.0 ;
      RECT  120000.0 252450.0 121200.0 251250.0 ;
      RECT  122400.0 252450.0 123600.0 251250.0 ;
      RECT  122400.0 252450.0 123600.0 251250.0 ;
      RECT  120000.0 252450.0 121200.0 251250.0 ;
      RECT  124800.0 243150.0 126000.0 241950.0 ;
      RECT  124800.0 253050.0 126000.0 251850.0 ;
      RECT  122400.0 249900.0 121200.0 248700.0 ;
      RECT  119400.0 247200.0 118200.0 246000.0 ;
      RECT  120000.0 243750.0 121200.0 242550.0 ;
      RECT  122400.0 252450.0 123600.0 251250.0 ;
      RECT  123600.0 247200.0 122400.0 246000.0 ;
      RECT  118200.0 247200.0 119400.0 246000.0 ;
      RECT  121200.0 249900.0 122400.0 248700.0 ;
      RECT  122400.0 247200.0 123600.0 246000.0 ;
      RECT  115800.0 241050.0 130200.0 240150.0 ;
      RECT  115800.0 254850.0 130200.0 253950.0 ;
      RECT  136800.0 242550.0 138000.0 240600.0 ;
      RECT  136800.0 254400.0 138000.0 252450.0 ;
      RECT  132000.0 253050.0 133200.0 254850.0 ;
      RECT  132000.0 243750.0 133200.0 240150.0 ;
      RECT  134700.0 253050.0 135600.0 243750.0 ;
      RECT  132000.0 243750.0 133200.0 242550.0 ;
      RECT  134400.0 243750.0 135600.0 242550.0 ;
      RECT  134400.0 243750.0 135600.0 242550.0 ;
      RECT  132000.0 243750.0 133200.0 242550.0 ;
      RECT  132000.0 253050.0 133200.0 251850.0 ;
      RECT  134400.0 253050.0 135600.0 251850.0 ;
      RECT  134400.0 253050.0 135600.0 251850.0 ;
      RECT  132000.0 253050.0 133200.0 251850.0 ;
      RECT  136800.0 243150.0 138000.0 241950.0 ;
      RECT  136800.0 253050.0 138000.0 251850.0 ;
      RECT  132600.0 248400.0 133800.0 247200.0 ;
      RECT  132600.0 248400.0 133800.0 247200.0 ;
      RECT  135150.0 248250.0 136050.0 247350.0 ;
      RECT  130200.0 241050.0 139800.0 240150.0 ;
      RECT  130200.0 254850.0 139800.0 253950.0 ;
      RECT  102450.0 247200.0 103650.0 248400.0 ;
      RECT  104400.0 249600.0 105600.0 250800.0 ;
      RECT  121200.0 248700.0 120000.0 249900.0 ;
      RECT  112800.0 266250.0 114000.0 268200.0 ;
      RECT  112800.0 254400.0 114000.0 256350.0 ;
      RECT  108000.0 255750.0 109200.0 253950.0 ;
      RECT  108000.0 265050.0 109200.0 268650.0 ;
      RECT  110700.0 255750.0 111600.0 265050.0 ;
      RECT  108000.0 265050.0 109200.0 266250.0 ;
      RECT  110400.0 265050.0 111600.0 266250.0 ;
      RECT  110400.0 265050.0 111600.0 266250.0 ;
      RECT  108000.0 265050.0 109200.0 266250.0 ;
      RECT  108000.0 255750.0 109200.0 256950.0 ;
      RECT  110400.0 255750.0 111600.0 256950.0 ;
      RECT  110400.0 255750.0 111600.0 256950.0 ;
      RECT  108000.0 255750.0 109200.0 256950.0 ;
      RECT  112800.0 265650.0 114000.0 266850.0 ;
      RECT  112800.0 255750.0 114000.0 256950.0 ;
      RECT  108600.0 260400.0 109800.0 261600.0 ;
      RECT  108600.0 260400.0 109800.0 261600.0 ;
      RECT  111150.0 260550.0 112050.0 261450.0 ;
      RECT  106200.0 267750.0 115800.0 268650.0 ;
      RECT  106200.0 253950.0 115800.0 254850.0 ;
      RECT  117600.0 256350.0 118800.0 253950.0 ;
      RECT  117600.0 265050.0 118800.0 268650.0 ;
      RECT  122400.0 265050.0 123600.0 268650.0 ;
      RECT  124800.0 266250.0 126000.0 268200.0 ;
      RECT  124800.0 254400.0 126000.0 256350.0 ;
      RECT  117600.0 265050.0 118800.0 266250.0 ;
      RECT  120000.0 265050.0 121200.0 266250.0 ;
      RECT  120000.0 265050.0 121200.0 266250.0 ;
      RECT  117600.0 265050.0 118800.0 266250.0 ;
      RECT  120000.0 265050.0 121200.0 266250.0 ;
      RECT  122400.0 265050.0 123600.0 266250.0 ;
      RECT  122400.0 265050.0 123600.0 266250.0 ;
      RECT  120000.0 265050.0 121200.0 266250.0 ;
      RECT  117600.0 256350.0 118800.0 257550.0 ;
      RECT  120000.0 256350.0 121200.0 257550.0 ;
      RECT  120000.0 256350.0 121200.0 257550.0 ;
      RECT  117600.0 256350.0 118800.0 257550.0 ;
      RECT  120000.0 256350.0 121200.0 257550.0 ;
      RECT  122400.0 256350.0 123600.0 257550.0 ;
      RECT  122400.0 256350.0 123600.0 257550.0 ;
      RECT  120000.0 256350.0 121200.0 257550.0 ;
      RECT  124800.0 265650.0 126000.0 266850.0 ;
      RECT  124800.0 255750.0 126000.0 256950.0 ;
      RECT  122400.0 258900.0 121200.0 260100.0 ;
      RECT  119400.0 261600.0 118200.0 262800.0 ;
      RECT  120000.0 265050.0 121200.0 266250.0 ;
      RECT  122400.0 256350.0 123600.0 257550.0 ;
      RECT  123600.0 261600.0 122400.0 262800.0 ;
      RECT  118200.0 261600.0 119400.0 262800.0 ;
      RECT  121200.0 258900.0 122400.0 260100.0 ;
      RECT  122400.0 261600.0 123600.0 262800.0 ;
      RECT  115800.0 267750.0 130200.0 268650.0 ;
      RECT  115800.0 253950.0 130200.0 254850.0 ;
      RECT  136800.0 266250.0 138000.0 268200.0 ;
      RECT  136800.0 254400.0 138000.0 256350.0 ;
      RECT  132000.0 255750.0 133200.0 253950.0 ;
      RECT  132000.0 265050.0 133200.0 268650.0 ;
      RECT  134700.0 255750.0 135600.0 265050.0 ;
      RECT  132000.0 265050.0 133200.0 266250.0 ;
      RECT  134400.0 265050.0 135600.0 266250.0 ;
      RECT  134400.0 265050.0 135600.0 266250.0 ;
      RECT  132000.0 265050.0 133200.0 266250.0 ;
      RECT  132000.0 255750.0 133200.0 256950.0 ;
      RECT  134400.0 255750.0 135600.0 256950.0 ;
      RECT  134400.0 255750.0 135600.0 256950.0 ;
      RECT  132000.0 255750.0 133200.0 256950.0 ;
      RECT  136800.0 265650.0 138000.0 266850.0 ;
      RECT  136800.0 255750.0 138000.0 256950.0 ;
      RECT  132600.0 260400.0 133800.0 261600.0 ;
      RECT  132600.0 260400.0 133800.0 261600.0 ;
      RECT  135150.0 260550.0 136050.0 261450.0 ;
      RECT  130200.0 267750.0 139800.0 268650.0 ;
      RECT  130200.0 253950.0 139800.0 254850.0 ;
      RECT  102450.0 260400.0 103650.0 261600.0 ;
      RECT  104400.0 258000.0 105600.0 259200.0 ;
      RECT  121200.0 258900.0 120000.0 260100.0 ;
      RECT  112800.0 270150.0 114000.0 268200.0 ;
      RECT  112800.0 282000.0 114000.0 280050.0 ;
      RECT  108000.0 280650.0 109200.0 282450.0 ;
      RECT  108000.0 271350.0 109200.0 267750.0 ;
      RECT  110700.0 280650.0 111600.0 271350.0 ;
      RECT  108000.0 271350.0 109200.0 270150.0 ;
      RECT  110400.0 271350.0 111600.0 270150.0 ;
      RECT  110400.0 271350.0 111600.0 270150.0 ;
      RECT  108000.0 271350.0 109200.0 270150.0 ;
      RECT  108000.0 280650.0 109200.0 279450.0 ;
      RECT  110400.0 280650.0 111600.0 279450.0 ;
      RECT  110400.0 280650.0 111600.0 279450.0 ;
      RECT  108000.0 280650.0 109200.0 279450.0 ;
      RECT  112800.0 270750.0 114000.0 269550.0 ;
      RECT  112800.0 280650.0 114000.0 279450.0 ;
      RECT  108600.0 276000.0 109800.0 274800.0 ;
      RECT  108600.0 276000.0 109800.0 274800.0 ;
      RECT  111150.0 275850.0 112050.0 274950.0 ;
      RECT  106200.0 268650.0 115800.0 267750.0 ;
      RECT  106200.0 282450.0 115800.0 281550.0 ;
      RECT  117600.0 280050.0 118800.0 282450.0 ;
      RECT  117600.0 271350.0 118800.0 267750.0 ;
      RECT  122400.0 271350.0 123600.0 267750.0 ;
      RECT  124800.0 270150.0 126000.0 268200.0 ;
      RECT  124800.0 282000.0 126000.0 280050.0 ;
      RECT  117600.0 271350.0 118800.0 270150.0 ;
      RECT  120000.0 271350.0 121200.0 270150.0 ;
      RECT  120000.0 271350.0 121200.0 270150.0 ;
      RECT  117600.0 271350.0 118800.0 270150.0 ;
      RECT  120000.0 271350.0 121200.0 270150.0 ;
      RECT  122400.0 271350.0 123600.0 270150.0 ;
      RECT  122400.0 271350.0 123600.0 270150.0 ;
      RECT  120000.0 271350.0 121200.0 270150.0 ;
      RECT  117600.0 280050.0 118800.0 278850.0 ;
      RECT  120000.0 280050.0 121200.0 278850.0 ;
      RECT  120000.0 280050.0 121200.0 278850.0 ;
      RECT  117600.0 280050.0 118800.0 278850.0 ;
      RECT  120000.0 280050.0 121200.0 278850.0 ;
      RECT  122400.0 280050.0 123600.0 278850.0 ;
      RECT  122400.0 280050.0 123600.0 278850.0 ;
      RECT  120000.0 280050.0 121200.0 278850.0 ;
      RECT  124800.0 270750.0 126000.0 269550.0 ;
      RECT  124800.0 280650.0 126000.0 279450.0 ;
      RECT  122400.0 277500.0 121200.0 276300.0 ;
      RECT  119400.0 274800.0 118200.0 273600.0 ;
      RECT  120000.0 271350.0 121200.0 270150.0 ;
      RECT  122400.0 280050.0 123600.0 278850.0 ;
      RECT  123600.0 274800.0 122400.0 273600.0 ;
      RECT  118200.0 274800.0 119400.0 273600.0 ;
      RECT  121200.0 277500.0 122400.0 276300.0 ;
      RECT  122400.0 274800.0 123600.0 273600.0 ;
      RECT  115800.0 268650.0 130200.0 267750.0 ;
      RECT  115800.0 282450.0 130200.0 281550.0 ;
      RECT  136800.0 270150.0 138000.0 268200.0 ;
      RECT  136800.0 282000.0 138000.0 280050.0 ;
      RECT  132000.0 280650.0 133200.0 282450.0 ;
      RECT  132000.0 271350.0 133200.0 267750.0 ;
      RECT  134700.0 280650.0 135600.0 271350.0 ;
      RECT  132000.0 271350.0 133200.0 270150.0 ;
      RECT  134400.0 271350.0 135600.0 270150.0 ;
      RECT  134400.0 271350.0 135600.0 270150.0 ;
      RECT  132000.0 271350.0 133200.0 270150.0 ;
      RECT  132000.0 280650.0 133200.0 279450.0 ;
      RECT  134400.0 280650.0 135600.0 279450.0 ;
      RECT  134400.0 280650.0 135600.0 279450.0 ;
      RECT  132000.0 280650.0 133200.0 279450.0 ;
      RECT  136800.0 270750.0 138000.0 269550.0 ;
      RECT  136800.0 280650.0 138000.0 279450.0 ;
      RECT  132600.0 276000.0 133800.0 274800.0 ;
      RECT  132600.0 276000.0 133800.0 274800.0 ;
      RECT  135150.0 275850.0 136050.0 274950.0 ;
      RECT  130200.0 268650.0 139800.0 267750.0 ;
      RECT  130200.0 282450.0 139800.0 281550.0 ;
      RECT  102450.0 274800.0 103650.0 276000.0 ;
      RECT  104400.0 277200.0 105600.0 278400.0 ;
      RECT  121200.0 276300.0 120000.0 277500.0 ;
      RECT  112800.0 293850.0 114000.0 295800.0 ;
      RECT  112800.0 282000.0 114000.0 283950.0 ;
      RECT  108000.0 283350.0 109200.0 281550.0 ;
      RECT  108000.0 292650.0 109200.0 296250.0 ;
      RECT  110700.0 283350.0 111600.0 292650.0 ;
      RECT  108000.0 292650.0 109200.0 293850.0 ;
      RECT  110400.0 292650.0 111600.0 293850.0 ;
      RECT  110400.0 292650.0 111600.0 293850.0 ;
      RECT  108000.0 292650.0 109200.0 293850.0 ;
      RECT  108000.0 283350.0 109200.0 284550.0 ;
      RECT  110400.0 283350.0 111600.0 284550.0 ;
      RECT  110400.0 283350.0 111600.0 284550.0 ;
      RECT  108000.0 283350.0 109200.0 284550.0 ;
      RECT  112800.0 293250.0 114000.0 294450.0 ;
      RECT  112800.0 283350.0 114000.0 284550.0 ;
      RECT  108600.0 288000.0 109800.0 289200.0 ;
      RECT  108600.0 288000.0 109800.0 289200.0 ;
      RECT  111150.0 288150.0 112050.0 289050.0 ;
      RECT  106200.0 295350.0 115800.0 296250.0 ;
      RECT  106200.0 281550.0 115800.0 282450.0 ;
      RECT  117600.0 283950.0 118800.0 281550.0 ;
      RECT  117600.0 292650.0 118800.0 296250.0 ;
      RECT  122400.0 292650.0 123600.0 296250.0 ;
      RECT  124800.0 293850.0 126000.0 295800.0 ;
      RECT  124800.0 282000.0 126000.0 283950.0 ;
      RECT  117600.0 292650.0 118800.0 293850.0 ;
      RECT  120000.0 292650.0 121200.0 293850.0 ;
      RECT  120000.0 292650.0 121200.0 293850.0 ;
      RECT  117600.0 292650.0 118800.0 293850.0 ;
      RECT  120000.0 292650.0 121200.0 293850.0 ;
      RECT  122400.0 292650.0 123600.0 293850.0 ;
      RECT  122400.0 292650.0 123600.0 293850.0 ;
      RECT  120000.0 292650.0 121200.0 293850.0 ;
      RECT  117600.0 283950.0 118800.0 285150.0 ;
      RECT  120000.0 283950.0 121200.0 285150.0 ;
      RECT  120000.0 283950.0 121200.0 285150.0 ;
      RECT  117600.0 283950.0 118800.0 285150.0 ;
      RECT  120000.0 283950.0 121200.0 285150.0 ;
      RECT  122400.0 283950.0 123600.0 285150.0 ;
      RECT  122400.0 283950.0 123600.0 285150.0 ;
      RECT  120000.0 283950.0 121200.0 285150.0 ;
      RECT  124800.0 293250.0 126000.0 294450.0 ;
      RECT  124800.0 283350.0 126000.0 284550.0 ;
      RECT  122400.0 286500.0 121200.0 287700.0 ;
      RECT  119400.0 289200.0 118200.0 290400.0 ;
      RECT  120000.0 292650.0 121200.0 293850.0 ;
      RECT  122400.0 283950.0 123600.0 285150.0 ;
      RECT  123600.0 289200.0 122400.0 290400.0 ;
      RECT  118200.0 289200.0 119400.0 290400.0 ;
      RECT  121200.0 286500.0 122400.0 287700.0 ;
      RECT  122400.0 289200.0 123600.0 290400.0 ;
      RECT  115800.0 295350.0 130200.0 296250.0 ;
      RECT  115800.0 281550.0 130200.0 282450.0 ;
      RECT  136800.0 293850.0 138000.0 295800.0 ;
      RECT  136800.0 282000.0 138000.0 283950.0 ;
      RECT  132000.0 283350.0 133200.0 281550.0 ;
      RECT  132000.0 292650.0 133200.0 296250.0 ;
      RECT  134700.0 283350.0 135600.0 292650.0 ;
      RECT  132000.0 292650.0 133200.0 293850.0 ;
      RECT  134400.0 292650.0 135600.0 293850.0 ;
      RECT  134400.0 292650.0 135600.0 293850.0 ;
      RECT  132000.0 292650.0 133200.0 293850.0 ;
      RECT  132000.0 283350.0 133200.0 284550.0 ;
      RECT  134400.0 283350.0 135600.0 284550.0 ;
      RECT  134400.0 283350.0 135600.0 284550.0 ;
      RECT  132000.0 283350.0 133200.0 284550.0 ;
      RECT  136800.0 293250.0 138000.0 294450.0 ;
      RECT  136800.0 283350.0 138000.0 284550.0 ;
      RECT  132600.0 288000.0 133800.0 289200.0 ;
      RECT  132600.0 288000.0 133800.0 289200.0 ;
      RECT  135150.0 288150.0 136050.0 289050.0 ;
      RECT  130200.0 295350.0 139800.0 296250.0 ;
      RECT  130200.0 281550.0 139800.0 282450.0 ;
      RECT  102450.0 288000.0 103650.0 289200.0 ;
      RECT  104400.0 285600.0 105600.0 286800.0 ;
      RECT  121200.0 286500.0 120000.0 287700.0 ;
      RECT  112800.0 297750.0 114000.0 295800.0 ;
      RECT  112800.0 309600.0 114000.0 307650.0 ;
      RECT  108000.0 308250.0 109200.0 310050.0 ;
      RECT  108000.0 298950.0 109200.0 295350.0 ;
      RECT  110700.0 308250.0 111600.0 298950.0 ;
      RECT  108000.0 298950.0 109200.0 297750.0 ;
      RECT  110400.0 298950.0 111600.0 297750.0 ;
      RECT  110400.0 298950.0 111600.0 297750.0 ;
      RECT  108000.0 298950.0 109200.0 297750.0 ;
      RECT  108000.0 308250.0 109200.0 307050.0 ;
      RECT  110400.0 308250.0 111600.0 307050.0 ;
      RECT  110400.0 308250.0 111600.0 307050.0 ;
      RECT  108000.0 308250.0 109200.0 307050.0 ;
      RECT  112800.0 298350.0 114000.0 297150.0 ;
      RECT  112800.0 308250.0 114000.0 307050.0 ;
      RECT  108600.0 303600.0 109800.0 302400.0 ;
      RECT  108600.0 303600.0 109800.0 302400.0 ;
      RECT  111150.0 303450.0 112050.0 302550.0 ;
      RECT  106200.0 296250.0 115800.0 295350.0 ;
      RECT  106200.0 310050.0 115800.0 309150.0 ;
      RECT  117600.0 307650.0 118800.0 310050.0 ;
      RECT  117600.0 298950.0 118800.0 295350.0 ;
      RECT  122400.0 298950.0 123600.0 295350.0 ;
      RECT  124800.0 297750.0 126000.0 295800.0 ;
      RECT  124800.0 309600.0 126000.0 307650.0 ;
      RECT  117600.0 298950.0 118800.0 297750.0 ;
      RECT  120000.0 298950.0 121200.0 297750.0 ;
      RECT  120000.0 298950.0 121200.0 297750.0 ;
      RECT  117600.0 298950.0 118800.0 297750.0 ;
      RECT  120000.0 298950.0 121200.0 297750.0 ;
      RECT  122400.0 298950.0 123600.0 297750.0 ;
      RECT  122400.0 298950.0 123600.0 297750.0 ;
      RECT  120000.0 298950.0 121200.0 297750.0 ;
      RECT  117600.0 307650.0 118800.0 306450.0 ;
      RECT  120000.0 307650.0 121200.0 306450.0 ;
      RECT  120000.0 307650.0 121200.0 306450.0 ;
      RECT  117600.0 307650.0 118800.0 306450.0 ;
      RECT  120000.0 307650.0 121200.0 306450.0 ;
      RECT  122400.0 307650.0 123600.0 306450.0 ;
      RECT  122400.0 307650.0 123600.0 306450.0 ;
      RECT  120000.0 307650.0 121200.0 306450.0 ;
      RECT  124800.0 298350.0 126000.0 297150.0 ;
      RECT  124800.0 308250.0 126000.0 307050.0 ;
      RECT  122400.0 305100.0 121200.0 303900.0 ;
      RECT  119400.0 302400.0 118200.0 301200.0 ;
      RECT  120000.0 298950.0 121200.0 297750.0 ;
      RECT  122400.0 307650.0 123600.0 306450.0 ;
      RECT  123600.0 302400.0 122400.0 301200.0 ;
      RECT  118200.0 302400.0 119400.0 301200.0 ;
      RECT  121200.0 305100.0 122400.0 303900.0 ;
      RECT  122400.0 302400.0 123600.0 301200.0 ;
      RECT  115800.0 296250.0 130200.0 295350.0 ;
      RECT  115800.0 310050.0 130200.0 309150.0 ;
      RECT  136800.0 297750.0 138000.0 295800.0 ;
      RECT  136800.0 309600.0 138000.0 307650.0 ;
      RECT  132000.0 308250.0 133200.0 310050.0 ;
      RECT  132000.0 298950.0 133200.0 295350.0 ;
      RECT  134700.0 308250.0 135600.0 298950.0 ;
      RECT  132000.0 298950.0 133200.0 297750.0 ;
      RECT  134400.0 298950.0 135600.0 297750.0 ;
      RECT  134400.0 298950.0 135600.0 297750.0 ;
      RECT  132000.0 298950.0 133200.0 297750.0 ;
      RECT  132000.0 308250.0 133200.0 307050.0 ;
      RECT  134400.0 308250.0 135600.0 307050.0 ;
      RECT  134400.0 308250.0 135600.0 307050.0 ;
      RECT  132000.0 308250.0 133200.0 307050.0 ;
      RECT  136800.0 298350.0 138000.0 297150.0 ;
      RECT  136800.0 308250.0 138000.0 307050.0 ;
      RECT  132600.0 303600.0 133800.0 302400.0 ;
      RECT  132600.0 303600.0 133800.0 302400.0 ;
      RECT  135150.0 303450.0 136050.0 302550.0 ;
      RECT  130200.0 296250.0 139800.0 295350.0 ;
      RECT  130200.0 310050.0 139800.0 309150.0 ;
      RECT  102450.0 302400.0 103650.0 303600.0 ;
      RECT  104400.0 304800.0 105600.0 306000.0 ;
      RECT  121200.0 303900.0 120000.0 305100.0 ;
      RECT  112800.0 321450.0 114000.0 323400.0 ;
      RECT  112800.0 309600.0 114000.0 311550.0 ;
      RECT  108000.0 310950.0 109200.0 309150.0 ;
      RECT  108000.0 320250.0 109200.0 323850.0 ;
      RECT  110700.0 310950.0 111600.0 320250.0 ;
      RECT  108000.0 320250.0 109200.0 321450.0 ;
      RECT  110400.0 320250.0 111600.0 321450.0 ;
      RECT  110400.0 320250.0 111600.0 321450.0 ;
      RECT  108000.0 320250.0 109200.0 321450.0 ;
      RECT  108000.0 310950.0 109200.0 312150.0 ;
      RECT  110400.0 310950.0 111600.0 312150.0 ;
      RECT  110400.0 310950.0 111600.0 312150.0 ;
      RECT  108000.0 310950.0 109200.0 312150.0 ;
      RECT  112800.0 320850.0 114000.0 322050.0 ;
      RECT  112800.0 310950.0 114000.0 312150.0 ;
      RECT  108600.0 315600.0 109800.0 316800.0 ;
      RECT  108600.0 315600.0 109800.0 316800.0 ;
      RECT  111150.0 315750.0 112050.0 316650.0 ;
      RECT  106200.0 322950.0 115800.0 323850.0 ;
      RECT  106200.0 309150.0 115800.0 310050.0 ;
      RECT  117600.0 311550.0 118800.0 309150.0 ;
      RECT  117600.0 320250.0 118800.0 323850.0 ;
      RECT  122400.0 320250.0 123600.0 323850.0 ;
      RECT  124800.0 321450.0 126000.0 323400.0 ;
      RECT  124800.0 309600.0 126000.0 311550.0 ;
      RECT  117600.0 320250.0 118800.0 321450.0 ;
      RECT  120000.0 320250.0 121200.0 321450.0 ;
      RECT  120000.0 320250.0 121200.0 321450.0 ;
      RECT  117600.0 320250.0 118800.0 321450.0 ;
      RECT  120000.0 320250.0 121200.0 321450.0 ;
      RECT  122400.0 320250.0 123600.0 321450.0 ;
      RECT  122400.0 320250.0 123600.0 321450.0 ;
      RECT  120000.0 320250.0 121200.0 321450.0 ;
      RECT  117600.0 311550.0 118800.0 312750.0 ;
      RECT  120000.0 311550.0 121200.0 312750.0 ;
      RECT  120000.0 311550.0 121200.0 312750.0 ;
      RECT  117600.0 311550.0 118800.0 312750.0 ;
      RECT  120000.0 311550.0 121200.0 312750.0 ;
      RECT  122400.0 311550.0 123600.0 312750.0 ;
      RECT  122400.0 311550.0 123600.0 312750.0 ;
      RECT  120000.0 311550.0 121200.0 312750.0 ;
      RECT  124800.0 320850.0 126000.0 322050.0 ;
      RECT  124800.0 310950.0 126000.0 312150.0 ;
      RECT  122400.0 314100.0 121200.0 315300.0 ;
      RECT  119400.0 316800.0 118200.0 318000.0 ;
      RECT  120000.0 320250.0 121200.0 321450.0 ;
      RECT  122400.0 311550.0 123600.0 312750.0 ;
      RECT  123600.0 316800.0 122400.0 318000.0 ;
      RECT  118200.0 316800.0 119400.0 318000.0 ;
      RECT  121200.0 314100.0 122400.0 315300.0 ;
      RECT  122400.0 316800.0 123600.0 318000.0 ;
      RECT  115800.0 322950.0 130200.0 323850.0 ;
      RECT  115800.0 309150.0 130200.0 310050.0 ;
      RECT  136800.0 321450.0 138000.0 323400.0 ;
      RECT  136800.0 309600.0 138000.0 311550.0 ;
      RECT  132000.0 310950.0 133200.0 309150.0 ;
      RECT  132000.0 320250.0 133200.0 323850.0 ;
      RECT  134700.0 310950.0 135600.0 320250.0 ;
      RECT  132000.0 320250.0 133200.0 321450.0 ;
      RECT  134400.0 320250.0 135600.0 321450.0 ;
      RECT  134400.0 320250.0 135600.0 321450.0 ;
      RECT  132000.0 320250.0 133200.0 321450.0 ;
      RECT  132000.0 310950.0 133200.0 312150.0 ;
      RECT  134400.0 310950.0 135600.0 312150.0 ;
      RECT  134400.0 310950.0 135600.0 312150.0 ;
      RECT  132000.0 310950.0 133200.0 312150.0 ;
      RECT  136800.0 320850.0 138000.0 322050.0 ;
      RECT  136800.0 310950.0 138000.0 312150.0 ;
      RECT  132600.0 315600.0 133800.0 316800.0 ;
      RECT  132600.0 315600.0 133800.0 316800.0 ;
      RECT  135150.0 315750.0 136050.0 316650.0 ;
      RECT  130200.0 322950.0 139800.0 323850.0 ;
      RECT  130200.0 309150.0 139800.0 310050.0 ;
      RECT  102450.0 315600.0 103650.0 316800.0 ;
      RECT  104400.0 313200.0 105600.0 314400.0 ;
      RECT  121200.0 314100.0 120000.0 315300.0 ;
      RECT  112800.0 325350.0 114000.0 323400.0 ;
      RECT  112800.0 337200.0 114000.0 335250.0 ;
      RECT  108000.0 335850.0 109200.0 337650.0 ;
      RECT  108000.0 326550.0 109200.0 322950.0 ;
      RECT  110700.0 335850.0 111600.0 326550.0 ;
      RECT  108000.0 326550.0 109200.0 325350.0 ;
      RECT  110400.0 326550.0 111600.0 325350.0 ;
      RECT  110400.0 326550.0 111600.0 325350.0 ;
      RECT  108000.0 326550.0 109200.0 325350.0 ;
      RECT  108000.0 335850.0 109200.0 334650.0 ;
      RECT  110400.0 335850.0 111600.0 334650.0 ;
      RECT  110400.0 335850.0 111600.0 334650.0 ;
      RECT  108000.0 335850.0 109200.0 334650.0 ;
      RECT  112800.0 325950.0 114000.0 324750.0 ;
      RECT  112800.0 335850.0 114000.0 334650.0 ;
      RECT  108600.0 331200.0 109800.0 330000.0 ;
      RECT  108600.0 331200.0 109800.0 330000.0 ;
      RECT  111150.0 331050.0 112050.0 330150.0 ;
      RECT  106200.0 323850.0 115800.0 322950.0 ;
      RECT  106200.0 337650.0 115800.0 336750.0 ;
      RECT  117600.0 335250.0 118800.0 337650.0 ;
      RECT  117600.0 326550.0 118800.0 322950.0 ;
      RECT  122400.0 326550.0 123600.0 322950.0 ;
      RECT  124800.0 325350.0 126000.0 323400.0 ;
      RECT  124800.0 337200.0 126000.0 335250.0 ;
      RECT  117600.0 326550.0 118800.0 325350.0 ;
      RECT  120000.0 326550.0 121200.0 325350.0 ;
      RECT  120000.0 326550.0 121200.0 325350.0 ;
      RECT  117600.0 326550.0 118800.0 325350.0 ;
      RECT  120000.0 326550.0 121200.0 325350.0 ;
      RECT  122400.0 326550.0 123600.0 325350.0 ;
      RECT  122400.0 326550.0 123600.0 325350.0 ;
      RECT  120000.0 326550.0 121200.0 325350.0 ;
      RECT  117600.0 335250.0 118800.0 334050.0 ;
      RECT  120000.0 335250.0 121200.0 334050.0 ;
      RECT  120000.0 335250.0 121200.0 334050.0 ;
      RECT  117600.0 335250.0 118800.0 334050.0 ;
      RECT  120000.0 335250.0 121200.0 334050.0 ;
      RECT  122400.0 335250.0 123600.0 334050.0 ;
      RECT  122400.0 335250.0 123600.0 334050.0 ;
      RECT  120000.0 335250.0 121200.0 334050.0 ;
      RECT  124800.0 325950.0 126000.0 324750.0 ;
      RECT  124800.0 335850.0 126000.0 334650.0 ;
      RECT  122400.0 332700.0 121200.0 331500.0 ;
      RECT  119400.0 330000.0 118200.0 328800.0 ;
      RECT  120000.0 326550.0 121200.0 325350.0 ;
      RECT  122400.0 335250.0 123600.0 334050.0 ;
      RECT  123600.0 330000.0 122400.0 328800.0 ;
      RECT  118200.0 330000.0 119400.0 328800.0 ;
      RECT  121200.0 332700.0 122400.0 331500.0 ;
      RECT  122400.0 330000.0 123600.0 328800.0 ;
      RECT  115800.0 323850.0 130200.0 322950.0 ;
      RECT  115800.0 337650.0 130200.0 336750.0 ;
      RECT  136800.0 325350.0 138000.0 323400.0 ;
      RECT  136800.0 337200.0 138000.0 335250.0 ;
      RECT  132000.0 335850.0 133200.0 337650.0 ;
      RECT  132000.0 326550.0 133200.0 322950.0 ;
      RECT  134700.0 335850.0 135600.0 326550.0 ;
      RECT  132000.0 326550.0 133200.0 325350.0 ;
      RECT  134400.0 326550.0 135600.0 325350.0 ;
      RECT  134400.0 326550.0 135600.0 325350.0 ;
      RECT  132000.0 326550.0 133200.0 325350.0 ;
      RECT  132000.0 335850.0 133200.0 334650.0 ;
      RECT  134400.0 335850.0 135600.0 334650.0 ;
      RECT  134400.0 335850.0 135600.0 334650.0 ;
      RECT  132000.0 335850.0 133200.0 334650.0 ;
      RECT  136800.0 325950.0 138000.0 324750.0 ;
      RECT  136800.0 335850.0 138000.0 334650.0 ;
      RECT  132600.0 331200.0 133800.0 330000.0 ;
      RECT  132600.0 331200.0 133800.0 330000.0 ;
      RECT  135150.0 331050.0 136050.0 330150.0 ;
      RECT  130200.0 323850.0 139800.0 322950.0 ;
      RECT  130200.0 337650.0 139800.0 336750.0 ;
      RECT  102450.0 330000.0 103650.0 331200.0 ;
      RECT  104400.0 332400.0 105600.0 333600.0 ;
      RECT  121200.0 331500.0 120000.0 332700.0 ;
      RECT  112800.0 349050.0 114000.0 351000.0 ;
      RECT  112800.0 337200.0 114000.0 339150.0 ;
      RECT  108000.0 338550.0 109200.0 336750.0 ;
      RECT  108000.0 347850.0 109200.0 351450.0 ;
      RECT  110700.0 338550.0 111600.0 347850.0 ;
      RECT  108000.0 347850.0 109200.0 349050.0 ;
      RECT  110400.0 347850.0 111600.0 349050.0 ;
      RECT  110400.0 347850.0 111600.0 349050.0 ;
      RECT  108000.0 347850.0 109200.0 349050.0 ;
      RECT  108000.0 338550.0 109200.0 339750.0 ;
      RECT  110400.0 338550.0 111600.0 339750.0 ;
      RECT  110400.0 338550.0 111600.0 339750.0 ;
      RECT  108000.0 338550.0 109200.0 339750.0 ;
      RECT  112800.0 348450.0 114000.0 349650.0 ;
      RECT  112800.0 338550.0 114000.0 339750.0 ;
      RECT  108600.0 343200.0 109800.0 344400.0 ;
      RECT  108600.0 343200.0 109800.0 344400.0 ;
      RECT  111150.0 343350.0 112050.0 344250.0 ;
      RECT  106200.0 350550.0 115800.0 351450.0 ;
      RECT  106200.0 336750.0 115800.0 337650.0 ;
      RECT  117600.0 339150.0 118800.0 336750.0 ;
      RECT  117600.0 347850.0 118800.0 351450.0 ;
      RECT  122400.0 347850.0 123600.0 351450.0 ;
      RECT  124800.0 349050.0 126000.0 351000.0 ;
      RECT  124800.0 337200.0 126000.0 339150.0 ;
      RECT  117600.0 347850.0 118800.0 349050.0 ;
      RECT  120000.0 347850.0 121200.0 349050.0 ;
      RECT  120000.0 347850.0 121200.0 349050.0 ;
      RECT  117600.0 347850.0 118800.0 349050.0 ;
      RECT  120000.0 347850.0 121200.0 349050.0 ;
      RECT  122400.0 347850.0 123600.0 349050.0 ;
      RECT  122400.0 347850.0 123600.0 349050.0 ;
      RECT  120000.0 347850.0 121200.0 349050.0 ;
      RECT  117600.0 339150.0 118800.0 340350.0 ;
      RECT  120000.0 339150.0 121200.0 340350.0 ;
      RECT  120000.0 339150.0 121200.0 340350.0 ;
      RECT  117600.0 339150.0 118800.0 340350.0 ;
      RECT  120000.0 339150.0 121200.0 340350.0 ;
      RECT  122400.0 339150.0 123600.0 340350.0 ;
      RECT  122400.0 339150.0 123600.0 340350.0 ;
      RECT  120000.0 339150.0 121200.0 340350.0 ;
      RECT  124800.0 348450.0 126000.0 349650.0 ;
      RECT  124800.0 338550.0 126000.0 339750.0 ;
      RECT  122400.0 341700.0 121200.0 342900.0 ;
      RECT  119400.0 344400.0 118200.0 345600.0 ;
      RECT  120000.0 347850.0 121200.0 349050.0 ;
      RECT  122400.0 339150.0 123600.0 340350.0 ;
      RECT  123600.0 344400.0 122400.0 345600.0 ;
      RECT  118200.0 344400.0 119400.0 345600.0 ;
      RECT  121200.0 341700.0 122400.0 342900.0 ;
      RECT  122400.0 344400.0 123600.0 345600.0 ;
      RECT  115800.0 350550.0 130200.0 351450.0 ;
      RECT  115800.0 336750.0 130200.0 337650.0 ;
      RECT  136800.0 349050.0 138000.0 351000.0 ;
      RECT  136800.0 337200.0 138000.0 339150.0 ;
      RECT  132000.0 338550.0 133200.0 336750.0 ;
      RECT  132000.0 347850.0 133200.0 351450.0 ;
      RECT  134700.0 338550.0 135600.0 347850.0 ;
      RECT  132000.0 347850.0 133200.0 349050.0 ;
      RECT  134400.0 347850.0 135600.0 349050.0 ;
      RECT  134400.0 347850.0 135600.0 349050.0 ;
      RECT  132000.0 347850.0 133200.0 349050.0 ;
      RECT  132000.0 338550.0 133200.0 339750.0 ;
      RECT  134400.0 338550.0 135600.0 339750.0 ;
      RECT  134400.0 338550.0 135600.0 339750.0 ;
      RECT  132000.0 338550.0 133200.0 339750.0 ;
      RECT  136800.0 348450.0 138000.0 349650.0 ;
      RECT  136800.0 338550.0 138000.0 339750.0 ;
      RECT  132600.0 343200.0 133800.0 344400.0 ;
      RECT  132600.0 343200.0 133800.0 344400.0 ;
      RECT  135150.0 343350.0 136050.0 344250.0 ;
      RECT  130200.0 350550.0 139800.0 351450.0 ;
      RECT  130200.0 336750.0 139800.0 337650.0 ;
      RECT  102450.0 343200.0 103650.0 344400.0 ;
      RECT  104400.0 340800.0 105600.0 342000.0 ;
      RECT  121200.0 341700.0 120000.0 342900.0 ;
      RECT  112800.0 352950.0 114000.0 351000.0 ;
      RECT  112800.0 364800.0 114000.0 362850.0 ;
      RECT  108000.0 363450.0 109200.0 365250.0 ;
      RECT  108000.0 354150.0 109200.0 350550.0 ;
      RECT  110700.0 363450.0 111600.0 354150.0 ;
      RECT  108000.0 354150.0 109200.0 352950.0 ;
      RECT  110400.0 354150.0 111600.0 352950.0 ;
      RECT  110400.0 354150.0 111600.0 352950.0 ;
      RECT  108000.0 354150.0 109200.0 352950.0 ;
      RECT  108000.0 363450.0 109200.0 362250.0 ;
      RECT  110400.0 363450.0 111600.0 362250.0 ;
      RECT  110400.0 363450.0 111600.0 362250.0 ;
      RECT  108000.0 363450.0 109200.0 362250.0 ;
      RECT  112800.0 353550.0 114000.0 352350.0 ;
      RECT  112800.0 363450.0 114000.0 362250.0 ;
      RECT  108600.0 358800.0 109800.0 357600.0 ;
      RECT  108600.0 358800.0 109800.0 357600.0 ;
      RECT  111150.0 358650.0 112050.0 357750.0 ;
      RECT  106200.0 351450.0 115800.0 350550.0 ;
      RECT  106200.0 365250.0 115800.0 364350.0 ;
      RECT  117600.0 362850.0 118800.0 365250.0 ;
      RECT  117600.0 354150.0 118800.0 350550.0 ;
      RECT  122400.0 354150.0 123600.0 350550.0 ;
      RECT  124800.0 352950.0 126000.0 351000.0 ;
      RECT  124800.0 364800.0 126000.0 362850.0 ;
      RECT  117600.0 354150.0 118800.0 352950.0 ;
      RECT  120000.0 354150.0 121200.0 352950.0 ;
      RECT  120000.0 354150.0 121200.0 352950.0 ;
      RECT  117600.0 354150.0 118800.0 352950.0 ;
      RECT  120000.0 354150.0 121200.0 352950.0 ;
      RECT  122400.0 354150.0 123600.0 352950.0 ;
      RECT  122400.0 354150.0 123600.0 352950.0 ;
      RECT  120000.0 354150.0 121200.0 352950.0 ;
      RECT  117600.0 362850.0 118800.0 361650.0 ;
      RECT  120000.0 362850.0 121200.0 361650.0 ;
      RECT  120000.0 362850.0 121200.0 361650.0 ;
      RECT  117600.0 362850.0 118800.0 361650.0 ;
      RECT  120000.0 362850.0 121200.0 361650.0 ;
      RECT  122400.0 362850.0 123600.0 361650.0 ;
      RECT  122400.0 362850.0 123600.0 361650.0 ;
      RECT  120000.0 362850.0 121200.0 361650.0 ;
      RECT  124800.0 353550.0 126000.0 352350.0 ;
      RECT  124800.0 363450.0 126000.0 362250.0 ;
      RECT  122400.0 360300.0 121200.0 359100.0 ;
      RECT  119400.0 357600.0 118200.0 356400.0 ;
      RECT  120000.0 354150.0 121200.0 352950.0 ;
      RECT  122400.0 362850.0 123600.0 361650.0 ;
      RECT  123600.0 357600.0 122400.0 356400.0 ;
      RECT  118200.0 357600.0 119400.0 356400.0 ;
      RECT  121200.0 360300.0 122400.0 359100.0 ;
      RECT  122400.0 357600.0 123600.0 356400.0 ;
      RECT  115800.0 351450.0 130200.0 350550.0 ;
      RECT  115800.0 365250.0 130200.0 364350.0 ;
      RECT  136800.0 352950.0 138000.0 351000.0 ;
      RECT  136800.0 364800.0 138000.0 362850.0 ;
      RECT  132000.0 363450.0 133200.0 365250.0 ;
      RECT  132000.0 354150.0 133200.0 350550.0 ;
      RECT  134700.0 363450.0 135600.0 354150.0 ;
      RECT  132000.0 354150.0 133200.0 352950.0 ;
      RECT  134400.0 354150.0 135600.0 352950.0 ;
      RECT  134400.0 354150.0 135600.0 352950.0 ;
      RECT  132000.0 354150.0 133200.0 352950.0 ;
      RECT  132000.0 363450.0 133200.0 362250.0 ;
      RECT  134400.0 363450.0 135600.0 362250.0 ;
      RECT  134400.0 363450.0 135600.0 362250.0 ;
      RECT  132000.0 363450.0 133200.0 362250.0 ;
      RECT  136800.0 353550.0 138000.0 352350.0 ;
      RECT  136800.0 363450.0 138000.0 362250.0 ;
      RECT  132600.0 358800.0 133800.0 357600.0 ;
      RECT  132600.0 358800.0 133800.0 357600.0 ;
      RECT  135150.0 358650.0 136050.0 357750.0 ;
      RECT  130200.0 351450.0 139800.0 350550.0 ;
      RECT  130200.0 365250.0 139800.0 364350.0 ;
      RECT  102450.0 357600.0 103650.0 358800.0 ;
      RECT  104400.0 360000.0 105600.0 361200.0 ;
      RECT  121200.0 359100.0 120000.0 360300.0 ;
      RECT  112800.0 376650.0 114000.0 378600.0 ;
      RECT  112800.0 364800.0 114000.0 366750.0 ;
      RECT  108000.0 366150.0 109200.0 364350.0 ;
      RECT  108000.0 375450.0 109200.0 379050.0 ;
      RECT  110700.0 366150.0 111600.0 375450.0 ;
      RECT  108000.0 375450.0 109200.0 376650.0 ;
      RECT  110400.0 375450.0 111600.0 376650.0 ;
      RECT  110400.0 375450.0 111600.0 376650.0 ;
      RECT  108000.0 375450.0 109200.0 376650.0 ;
      RECT  108000.0 366150.0 109200.0 367350.0 ;
      RECT  110400.0 366150.0 111600.0 367350.0 ;
      RECT  110400.0 366150.0 111600.0 367350.0 ;
      RECT  108000.0 366150.0 109200.0 367350.0 ;
      RECT  112800.0 376050.0 114000.0 377250.0 ;
      RECT  112800.0 366150.0 114000.0 367350.0 ;
      RECT  108600.0 370800.0 109800.0 372000.0 ;
      RECT  108600.0 370800.0 109800.0 372000.0 ;
      RECT  111150.0 370950.0 112050.0 371850.0 ;
      RECT  106200.0 378150.0 115800.0 379050.0 ;
      RECT  106200.0 364350.0 115800.0 365250.0 ;
      RECT  117600.0 366750.0 118800.0 364350.0 ;
      RECT  117600.0 375450.0 118800.0 379050.0 ;
      RECT  122400.0 375450.0 123600.0 379050.0 ;
      RECT  124800.0 376650.0 126000.0 378600.0 ;
      RECT  124800.0 364800.0 126000.0 366750.0 ;
      RECT  117600.0 375450.0 118800.0 376650.0 ;
      RECT  120000.0 375450.0 121200.0 376650.0 ;
      RECT  120000.0 375450.0 121200.0 376650.0 ;
      RECT  117600.0 375450.0 118800.0 376650.0 ;
      RECT  120000.0 375450.0 121200.0 376650.0 ;
      RECT  122400.0 375450.0 123600.0 376650.0 ;
      RECT  122400.0 375450.0 123600.0 376650.0 ;
      RECT  120000.0 375450.0 121200.0 376650.0 ;
      RECT  117600.0 366750.0 118800.0 367950.0 ;
      RECT  120000.0 366750.0 121200.0 367950.0 ;
      RECT  120000.0 366750.0 121200.0 367950.0 ;
      RECT  117600.0 366750.0 118800.0 367950.0 ;
      RECT  120000.0 366750.0 121200.0 367950.0 ;
      RECT  122400.0 366750.0 123600.0 367950.0 ;
      RECT  122400.0 366750.0 123600.0 367950.0 ;
      RECT  120000.0 366750.0 121200.0 367950.0 ;
      RECT  124800.0 376050.0 126000.0 377250.0 ;
      RECT  124800.0 366150.0 126000.0 367350.0 ;
      RECT  122400.0 369300.0 121200.0 370500.0 ;
      RECT  119400.0 372000.0 118200.0 373200.0 ;
      RECT  120000.0 375450.0 121200.0 376650.0 ;
      RECT  122400.0 366750.0 123600.0 367950.0 ;
      RECT  123600.0 372000.0 122400.0 373200.0 ;
      RECT  118200.0 372000.0 119400.0 373200.0 ;
      RECT  121200.0 369300.0 122400.0 370500.0 ;
      RECT  122400.0 372000.0 123600.0 373200.0 ;
      RECT  115800.0 378150.0 130200.0 379050.0 ;
      RECT  115800.0 364350.0 130200.0 365250.0 ;
      RECT  136800.0 376650.0 138000.0 378600.0 ;
      RECT  136800.0 364800.0 138000.0 366750.0 ;
      RECT  132000.0 366150.0 133200.0 364350.0 ;
      RECT  132000.0 375450.0 133200.0 379050.0 ;
      RECT  134700.0 366150.0 135600.0 375450.0 ;
      RECT  132000.0 375450.0 133200.0 376650.0 ;
      RECT  134400.0 375450.0 135600.0 376650.0 ;
      RECT  134400.0 375450.0 135600.0 376650.0 ;
      RECT  132000.0 375450.0 133200.0 376650.0 ;
      RECT  132000.0 366150.0 133200.0 367350.0 ;
      RECT  134400.0 366150.0 135600.0 367350.0 ;
      RECT  134400.0 366150.0 135600.0 367350.0 ;
      RECT  132000.0 366150.0 133200.0 367350.0 ;
      RECT  136800.0 376050.0 138000.0 377250.0 ;
      RECT  136800.0 366150.0 138000.0 367350.0 ;
      RECT  132600.0 370800.0 133800.0 372000.0 ;
      RECT  132600.0 370800.0 133800.0 372000.0 ;
      RECT  135150.0 370950.0 136050.0 371850.0 ;
      RECT  130200.0 378150.0 139800.0 379050.0 ;
      RECT  130200.0 364350.0 139800.0 365250.0 ;
      RECT  102450.0 370800.0 103650.0 372000.0 ;
      RECT  104400.0 368400.0 105600.0 369600.0 ;
      RECT  121200.0 369300.0 120000.0 370500.0 ;
      RECT  112800.0 380550.0 114000.0 378600.0 ;
      RECT  112800.0 392400.0 114000.0 390450.0 ;
      RECT  108000.0 391050.0 109200.0 392850.0 ;
      RECT  108000.0 381750.0 109200.0 378150.0 ;
      RECT  110700.0 391050.0 111600.0 381750.0 ;
      RECT  108000.0 381750.0 109200.0 380550.0 ;
      RECT  110400.0 381750.0 111600.0 380550.0 ;
      RECT  110400.0 381750.0 111600.0 380550.0 ;
      RECT  108000.0 381750.0 109200.0 380550.0 ;
      RECT  108000.0 391050.0 109200.0 389850.0 ;
      RECT  110400.0 391050.0 111600.0 389850.0 ;
      RECT  110400.0 391050.0 111600.0 389850.0 ;
      RECT  108000.0 391050.0 109200.0 389850.0 ;
      RECT  112800.0 381150.0 114000.0 379950.0 ;
      RECT  112800.0 391050.0 114000.0 389850.0 ;
      RECT  108600.0 386400.0 109800.0 385200.0 ;
      RECT  108600.0 386400.0 109800.0 385200.0 ;
      RECT  111150.0 386250.0 112050.0 385350.0 ;
      RECT  106200.0 379050.0 115800.0 378150.0 ;
      RECT  106200.0 392850.0 115800.0 391950.0 ;
      RECT  117600.0 390450.0 118800.0 392850.0 ;
      RECT  117600.0 381750.0 118800.0 378150.0 ;
      RECT  122400.0 381750.0 123600.0 378150.0 ;
      RECT  124800.0 380550.0 126000.0 378600.0 ;
      RECT  124800.0 392400.0 126000.0 390450.0 ;
      RECT  117600.0 381750.0 118800.0 380550.0 ;
      RECT  120000.0 381750.0 121200.0 380550.0 ;
      RECT  120000.0 381750.0 121200.0 380550.0 ;
      RECT  117600.0 381750.0 118800.0 380550.0 ;
      RECT  120000.0 381750.0 121200.0 380550.0 ;
      RECT  122400.0 381750.0 123600.0 380550.0 ;
      RECT  122400.0 381750.0 123600.0 380550.0 ;
      RECT  120000.0 381750.0 121200.0 380550.0 ;
      RECT  117600.0 390450.0 118800.0 389250.0 ;
      RECT  120000.0 390450.0 121200.0 389250.0 ;
      RECT  120000.0 390450.0 121200.0 389250.0 ;
      RECT  117600.0 390450.0 118800.0 389250.0 ;
      RECT  120000.0 390450.0 121200.0 389250.0 ;
      RECT  122400.0 390450.0 123600.0 389250.0 ;
      RECT  122400.0 390450.0 123600.0 389250.0 ;
      RECT  120000.0 390450.0 121200.0 389250.0 ;
      RECT  124800.0 381150.0 126000.0 379950.0 ;
      RECT  124800.0 391050.0 126000.0 389850.0 ;
      RECT  122400.0 387900.0 121200.0 386700.0 ;
      RECT  119400.0 385200.0 118200.0 384000.0 ;
      RECT  120000.0 381750.0 121200.0 380550.0 ;
      RECT  122400.0 390450.0 123600.0 389250.0 ;
      RECT  123600.0 385200.0 122400.0 384000.0 ;
      RECT  118200.0 385200.0 119400.0 384000.0 ;
      RECT  121200.0 387900.0 122400.0 386700.0 ;
      RECT  122400.0 385200.0 123600.0 384000.0 ;
      RECT  115800.0 379050.0 130200.0 378150.0 ;
      RECT  115800.0 392850.0 130200.0 391950.0 ;
      RECT  136800.0 380550.0 138000.0 378600.0 ;
      RECT  136800.0 392400.0 138000.0 390450.0 ;
      RECT  132000.0 391050.0 133200.0 392850.0 ;
      RECT  132000.0 381750.0 133200.0 378150.0 ;
      RECT  134700.0 391050.0 135600.0 381750.0 ;
      RECT  132000.0 381750.0 133200.0 380550.0 ;
      RECT  134400.0 381750.0 135600.0 380550.0 ;
      RECT  134400.0 381750.0 135600.0 380550.0 ;
      RECT  132000.0 381750.0 133200.0 380550.0 ;
      RECT  132000.0 391050.0 133200.0 389850.0 ;
      RECT  134400.0 391050.0 135600.0 389850.0 ;
      RECT  134400.0 391050.0 135600.0 389850.0 ;
      RECT  132000.0 391050.0 133200.0 389850.0 ;
      RECT  136800.0 381150.0 138000.0 379950.0 ;
      RECT  136800.0 391050.0 138000.0 389850.0 ;
      RECT  132600.0 386400.0 133800.0 385200.0 ;
      RECT  132600.0 386400.0 133800.0 385200.0 ;
      RECT  135150.0 386250.0 136050.0 385350.0 ;
      RECT  130200.0 379050.0 139800.0 378150.0 ;
      RECT  130200.0 392850.0 139800.0 391950.0 ;
      RECT  102450.0 385200.0 103650.0 386400.0 ;
      RECT  104400.0 387600.0 105600.0 388800.0 ;
      RECT  121200.0 386700.0 120000.0 387900.0 ;
      RECT  112800.0 404250.0 114000.0 406200.0 ;
      RECT  112800.0 392400.0 114000.0 394350.0 ;
      RECT  108000.0 393750.0 109200.0 391950.0 ;
      RECT  108000.0 403050.0 109200.0 406650.0 ;
      RECT  110700.0 393750.0 111600.0 403050.0 ;
      RECT  108000.0 403050.0 109200.0 404250.0 ;
      RECT  110400.0 403050.0 111600.0 404250.0 ;
      RECT  110400.0 403050.0 111600.0 404250.0 ;
      RECT  108000.0 403050.0 109200.0 404250.0 ;
      RECT  108000.0 393750.0 109200.0 394950.0 ;
      RECT  110400.0 393750.0 111600.0 394950.0 ;
      RECT  110400.0 393750.0 111600.0 394950.0 ;
      RECT  108000.0 393750.0 109200.0 394950.0 ;
      RECT  112800.0 403650.0 114000.0 404850.0 ;
      RECT  112800.0 393750.0 114000.0 394950.0 ;
      RECT  108600.0 398400.0 109800.0 399600.0 ;
      RECT  108600.0 398400.0 109800.0 399600.0 ;
      RECT  111150.0 398550.0 112050.0 399450.0 ;
      RECT  106200.0 405750.0 115800.0 406650.0 ;
      RECT  106200.0 391950.0 115800.0 392850.0 ;
      RECT  117600.0 394350.0 118800.0 391950.0 ;
      RECT  117600.0 403050.0 118800.0 406650.0 ;
      RECT  122400.0 403050.0 123600.0 406650.0 ;
      RECT  124800.0 404250.0 126000.0 406200.0 ;
      RECT  124800.0 392400.0 126000.0 394350.0 ;
      RECT  117600.0 403050.0 118800.0 404250.0 ;
      RECT  120000.0 403050.0 121200.0 404250.0 ;
      RECT  120000.0 403050.0 121200.0 404250.0 ;
      RECT  117600.0 403050.0 118800.0 404250.0 ;
      RECT  120000.0 403050.0 121200.0 404250.0 ;
      RECT  122400.0 403050.0 123600.0 404250.0 ;
      RECT  122400.0 403050.0 123600.0 404250.0 ;
      RECT  120000.0 403050.0 121200.0 404250.0 ;
      RECT  117600.0 394350.0 118800.0 395550.0 ;
      RECT  120000.0 394350.0 121200.0 395550.0 ;
      RECT  120000.0 394350.0 121200.0 395550.0 ;
      RECT  117600.0 394350.0 118800.0 395550.0 ;
      RECT  120000.0 394350.0 121200.0 395550.0 ;
      RECT  122400.0 394350.0 123600.0 395550.0 ;
      RECT  122400.0 394350.0 123600.0 395550.0 ;
      RECT  120000.0 394350.0 121200.0 395550.0 ;
      RECT  124800.0 403650.0 126000.0 404850.0 ;
      RECT  124800.0 393750.0 126000.0 394950.0 ;
      RECT  122400.0 396900.0 121200.0 398100.0 ;
      RECT  119400.0 399600.0 118200.0 400800.0 ;
      RECT  120000.0 403050.0 121200.0 404250.0 ;
      RECT  122400.0 394350.0 123600.0 395550.0 ;
      RECT  123600.0 399600.0 122400.0 400800.0 ;
      RECT  118200.0 399600.0 119400.0 400800.0 ;
      RECT  121200.0 396900.0 122400.0 398100.0 ;
      RECT  122400.0 399600.0 123600.0 400800.0 ;
      RECT  115800.0 405750.0 130200.0 406650.0 ;
      RECT  115800.0 391950.0 130200.0 392850.0 ;
      RECT  136800.0 404250.0 138000.0 406200.0 ;
      RECT  136800.0 392400.0 138000.0 394350.0 ;
      RECT  132000.0 393750.0 133200.0 391950.0 ;
      RECT  132000.0 403050.0 133200.0 406650.0 ;
      RECT  134700.0 393750.0 135600.0 403050.0 ;
      RECT  132000.0 403050.0 133200.0 404250.0 ;
      RECT  134400.0 403050.0 135600.0 404250.0 ;
      RECT  134400.0 403050.0 135600.0 404250.0 ;
      RECT  132000.0 403050.0 133200.0 404250.0 ;
      RECT  132000.0 393750.0 133200.0 394950.0 ;
      RECT  134400.0 393750.0 135600.0 394950.0 ;
      RECT  134400.0 393750.0 135600.0 394950.0 ;
      RECT  132000.0 393750.0 133200.0 394950.0 ;
      RECT  136800.0 403650.0 138000.0 404850.0 ;
      RECT  136800.0 393750.0 138000.0 394950.0 ;
      RECT  132600.0 398400.0 133800.0 399600.0 ;
      RECT  132600.0 398400.0 133800.0 399600.0 ;
      RECT  135150.0 398550.0 136050.0 399450.0 ;
      RECT  130200.0 405750.0 139800.0 406650.0 ;
      RECT  130200.0 391950.0 139800.0 392850.0 ;
      RECT  102450.0 398400.0 103650.0 399600.0 ;
      RECT  104400.0 396000.0 105600.0 397200.0 ;
      RECT  121200.0 396900.0 120000.0 398100.0 ;
      RECT  112800.0 408150.0 114000.0 406200.0 ;
      RECT  112800.0 420000.0 114000.0 418050.0 ;
      RECT  108000.0 418650.0 109200.0 420450.0 ;
      RECT  108000.0 409350.0 109200.0 405750.0 ;
      RECT  110700.0 418650.0 111600.0 409350.0 ;
      RECT  108000.0 409350.0 109200.0 408150.0 ;
      RECT  110400.0 409350.0 111600.0 408150.0 ;
      RECT  110400.0 409350.0 111600.0 408150.0 ;
      RECT  108000.0 409350.0 109200.0 408150.0 ;
      RECT  108000.0 418650.0 109200.0 417450.0 ;
      RECT  110400.0 418650.0 111600.0 417450.0 ;
      RECT  110400.0 418650.0 111600.0 417450.0 ;
      RECT  108000.0 418650.0 109200.0 417450.0 ;
      RECT  112800.0 408750.0 114000.0 407550.0 ;
      RECT  112800.0 418650.0 114000.0 417450.0 ;
      RECT  108600.0 414000.0 109800.0 412800.0 ;
      RECT  108600.0 414000.0 109800.0 412800.0 ;
      RECT  111150.0 413850.0 112050.0 412950.0 ;
      RECT  106200.0 406650.0 115800.0 405750.0 ;
      RECT  106200.0 420450.0 115800.0 419550.0 ;
      RECT  117600.0 418050.0 118800.0 420450.0 ;
      RECT  117600.0 409350.0 118800.0 405750.0 ;
      RECT  122400.0 409350.0 123600.0 405750.0 ;
      RECT  124800.0 408150.0 126000.0 406200.0 ;
      RECT  124800.0 420000.0 126000.0 418050.0 ;
      RECT  117600.0 409350.0 118800.0 408150.0 ;
      RECT  120000.0 409350.0 121200.0 408150.0 ;
      RECT  120000.0 409350.0 121200.0 408150.0 ;
      RECT  117600.0 409350.0 118800.0 408150.0 ;
      RECT  120000.0 409350.0 121200.0 408150.0 ;
      RECT  122400.0 409350.0 123600.0 408150.0 ;
      RECT  122400.0 409350.0 123600.0 408150.0 ;
      RECT  120000.0 409350.0 121200.0 408150.0 ;
      RECT  117600.0 418050.0 118800.0 416850.0 ;
      RECT  120000.0 418050.0 121200.0 416850.0 ;
      RECT  120000.0 418050.0 121200.0 416850.0 ;
      RECT  117600.0 418050.0 118800.0 416850.0 ;
      RECT  120000.0 418050.0 121200.0 416850.0 ;
      RECT  122400.0 418050.0 123600.0 416850.0 ;
      RECT  122400.0 418050.0 123600.0 416850.0 ;
      RECT  120000.0 418050.0 121200.0 416850.0 ;
      RECT  124800.0 408750.0 126000.0 407550.0 ;
      RECT  124800.0 418650.0 126000.0 417450.0 ;
      RECT  122400.0 415500.0 121200.0 414300.0 ;
      RECT  119400.0 412800.0 118200.0 411600.0 ;
      RECT  120000.0 409350.0 121200.0 408150.0 ;
      RECT  122400.0 418050.0 123600.0 416850.0 ;
      RECT  123600.0 412800.0 122400.0 411600.0 ;
      RECT  118200.0 412800.0 119400.0 411600.0 ;
      RECT  121200.0 415500.0 122400.0 414300.0 ;
      RECT  122400.0 412800.0 123600.0 411600.0 ;
      RECT  115800.0 406650.0 130200.0 405750.0 ;
      RECT  115800.0 420450.0 130200.0 419550.0 ;
      RECT  136800.0 408150.0 138000.0 406200.0 ;
      RECT  136800.0 420000.0 138000.0 418050.0 ;
      RECT  132000.0 418650.0 133200.0 420450.0 ;
      RECT  132000.0 409350.0 133200.0 405750.0 ;
      RECT  134700.0 418650.0 135600.0 409350.0 ;
      RECT  132000.0 409350.0 133200.0 408150.0 ;
      RECT  134400.0 409350.0 135600.0 408150.0 ;
      RECT  134400.0 409350.0 135600.0 408150.0 ;
      RECT  132000.0 409350.0 133200.0 408150.0 ;
      RECT  132000.0 418650.0 133200.0 417450.0 ;
      RECT  134400.0 418650.0 135600.0 417450.0 ;
      RECT  134400.0 418650.0 135600.0 417450.0 ;
      RECT  132000.0 418650.0 133200.0 417450.0 ;
      RECT  136800.0 408750.0 138000.0 407550.0 ;
      RECT  136800.0 418650.0 138000.0 417450.0 ;
      RECT  132600.0 414000.0 133800.0 412800.0 ;
      RECT  132600.0 414000.0 133800.0 412800.0 ;
      RECT  135150.0 413850.0 136050.0 412950.0 ;
      RECT  130200.0 406650.0 139800.0 405750.0 ;
      RECT  130200.0 420450.0 139800.0 419550.0 ;
      RECT  102450.0 412800.0 103650.0 414000.0 ;
      RECT  104400.0 415200.0 105600.0 416400.0 ;
      RECT  121200.0 414300.0 120000.0 415500.0 ;
      RECT  99900.0 202950.0 105000.0 203850.0 ;
      RECT  99900.0 222150.0 105000.0 223050.0 ;
      RECT  99900.0 230550.0 105000.0 231450.0 ;
      RECT  99900.0 249750.0 105000.0 250650.0 ;
      RECT  99900.0 258150.0 105000.0 259050.0 ;
      RECT  99900.0 277350.0 105000.0 278250.0 ;
      RECT  99900.0 285750.0 105000.0 286650.0 ;
      RECT  99900.0 304950.0 105000.0 305850.0 ;
      RECT  99900.0 313350.0 105000.0 314250.0 ;
      RECT  99900.0 332550.0 105000.0 333450.0 ;
      RECT  99900.0 340950.0 105000.0 341850.0 ;
      RECT  99900.0 360150.0 105000.0 361050.0 ;
      RECT  99900.0 368550.0 105000.0 369450.0 ;
      RECT  99900.0 387750.0 105000.0 388650.0 ;
      RECT  99900.0 396150.0 105000.0 397050.0 ;
      RECT  99900.0 415350.0 105000.0 416250.0 ;
      RECT  135150.0 205350.0 136050.0 206250.0 ;
      RECT  135150.0 219750.0 136050.0 220650.0 ;
      RECT  135150.0 232950.0 136050.0 233850.0 ;
      RECT  135150.0 247350.0 136050.0 248250.0 ;
      RECT  135150.0 260550.0 136050.0 261450.0 ;
      RECT  135150.0 274950.0 136050.0 275850.0 ;
      RECT  135150.0 288150.0 136050.0 289050.0 ;
      RECT  135150.0 302550.0 136050.0 303450.0 ;
      RECT  135150.0 315750.0 136050.0 316650.0 ;
      RECT  135150.0 330150.0 136050.0 331050.0 ;
      RECT  135150.0 343350.0 136050.0 344250.0 ;
      RECT  135150.0 357750.0 136050.0 358650.0 ;
      RECT  135150.0 370950.0 136050.0 371850.0 ;
      RECT  135150.0 385350.0 136050.0 386250.0 ;
      RECT  135150.0 398550.0 136050.0 399450.0 ;
      RECT  135150.0 412950.0 136050.0 413850.0 ;
      RECT  99900.0 212550.0 106200.0 213450.0 ;
      RECT  99900.0 240150.0 106200.0 241050.0 ;
      RECT  99900.0 267750.0 106200.0 268650.0 ;
      RECT  99900.0 295350.0 106200.0 296250.0 ;
      RECT  99900.0 322950.0 106200.0 323850.0 ;
      RECT  99900.0 350550.0 106200.0 351450.0 ;
      RECT  99900.0 378150.0 106200.0 379050.0 ;
      RECT  99900.0 405750.0 106200.0 406650.0 ;
      RECT  99900.0 198750.0 106200.0 199650.0 ;
      RECT  99900.0 226350.0 106200.0 227250.0 ;
      RECT  99900.0 253950.0 106200.0 254850.0 ;
      RECT  99900.0 281550.0 106200.0 282450.0 ;
      RECT  99900.0 309150.0 106200.0 310050.0 ;
      RECT  99900.0 336750.0 106200.0 337650.0 ;
      RECT  99900.0 364350.0 106200.0 365250.0 ;
      RECT  99900.0 391950.0 106200.0 392850.0 ;
      RECT  99900.0 419550.0 106200.0 420450.0 ;
      RECT  59100.0 83400.0 119100.0 73200.0 ;
      RECT  59100.0 63000.0 119100.0 73200.0 ;
      RECT  59100.0 63000.0 119100.0 52800.0 ;
      RECT  59100.0 42600.0 119100.0 52800.0 ;
      RECT  61500.0 83400.0 62400.0 42600.0 ;
      RECT  115500.0 83400.0 116400.0 42600.0 ;
      RECT  148050.0 199800.0 149250.0 198600.0 ;
      RECT  148050.0 227400.0 149250.0 226200.0 ;
      RECT  148050.0 255000.0 149250.0 253800.0 ;
      RECT  148050.0 282600.0 149250.0 281400.0 ;
      RECT  148050.0 310200.0 149250.0 309000.0 ;
      RECT  148050.0 337800.0 149250.0 336600.0 ;
      RECT  148050.0 365400.0 149250.0 364200.0 ;
      RECT  148050.0 393000.0 149250.0 391800.0 ;
      RECT  148050.0 420600.0 149250.0 419400.0 ;
      RECT  130500.0 91050.0 129300.0 92250.0 ;
      RECT  135600.0 90900.0 134400.0 92100.0 ;
      RECT  127500.0 104850.0 126300.0 106050.0 ;
      RECT  138300.0 104700.0 137100.0 105900.0 ;
      RECT  130500.0 146250.0 129300.0 147450.0 ;
      RECT  141000.0 146100.0 139800.0 147300.0 ;
      RECT  127500.0 160050.0 126300.0 161250.0 ;
      RECT  143700.0 159900.0 142500.0 161100.0 ;
      RECT  132600.0 88200.0 131400.0 89400.0 ;
      RECT  132600.0 115800.0 131400.0 117000.0 ;
      RECT  132600.0 143400.0 131400.0 144600.0 ;
      RECT  132600.0 171000.0 131400.0 172200.0 ;
      RECT  118500.0 76950.0 117300.0 78150.0 ;
      RECT  135600.0 76950.0 134400.0 78150.0 ;
      RECT  118500.0 68250.0 117300.0 69450.0 ;
      RECT  138300.0 68250.0 137100.0 69450.0 ;
      RECT  118500.0 56550.0 117300.0 57750.0 ;
      RECT  141000.0 56550.0 139800.0 57750.0 ;
      RECT  118500.0 47850.0 117300.0 49050.0 ;
      RECT  143700.0 47850.0 142500.0 49050.0 ;
      RECT  120300.0 72600.0 119100.0 73800.0 ;
      RECT  149250.0 72750.0 148050.0 73950.0 ;
      RECT  120300.0 52200.0 119100.0 53400.0 ;
      RECT  149250.0 52350.0 148050.0 53550.0 ;
      RECT  164400.0 32250.0 163200.0 33450.0 ;
      RECT  159000.0 27750.0 157800.0 28950.0 ;
      RECT  161700.0 25350.0 160500.0 26550.0 ;
      RECT  164400.0 424650.0 163200.0 425850.0 ;
      RECT  167100.0 96750.0 165900.0 97950.0 ;
      RECT  169800.0 194850.0 168600.0 196050.0 ;
      RECT  156300.0 84900.0 155100.0 86100.0 ;
      RECT  103650.0 421500.0 102450.0 422700.0 ;
      RECT  156300.0 421500.0 155100.0 422700.0 ;
      RECT  152550.0 23400.0 151350.0 24600.0 ;
      RECT  152550.0 192900.0 151350.0 194100.0 ;
      RECT  152550.0 94800.0 151350.0 96000.0 ;
      RECT  198600.0 0.0 203100.0 436800.0 ;
      RECT  52800.0 0.0 57300.0 436800.0 ;
      RECT  43650.0 207600.0 42750.0 217200.0 ;
      RECT  43800.0 223800.0 42900.0 224700.0 ;
      RECT  43350.0 223800.0 43200.0 224700.0 ;
      RECT  43800.0 224250.0 42900.0 231600.0 ;
      RECT  43800.0 243450.0 42900.0 250800.0 ;
      RECT  35550.0 258600.0 30600.0 259500.0 ;
      RECT  43650.0 207150.0 42750.0 208050.0 ;
      RECT  43650.0 223800.0 42750.0 224700.0 ;
      RECT  29250.0 362100.0 28350.0 375450.0 ;
      RECT  43800.0 272700.0 42900.0 284850.0 ;
      RECT  33300.0 204600.0 30600.0 205500.0 ;
      RECT  29700.0 284850.0 28800.0 311700.0 ;
      RECT  27000.0 290250.0 26100.0 314700.0 ;
      RECT  41700.0 303750.0 40800.0 312300.0 ;
      RECT  43650.0 301050.0 42750.0 314700.0 ;
      RECT  45600.0 292950.0 44700.0 317100.0 ;
      RECT  41700.0 326850.0 40800.0 327750.0 ;
      RECT  41700.0 318300.0 40800.0 327300.0 ;
      RECT  43200.0 326850.0 41250.0 327750.0 ;
      RECT  43800.0 329250.0 42900.0 330150.0 ;
      RECT  43350.0 329250.0 43200.0 330150.0 ;
      RECT  43800.0 329700.0 42900.0 387300.0 ;
      RECT  14100.0 303750.0 13200.0 321900.0 ;
      RECT  16050.0 292950.0 15150.0 324300.0 ;
      RECT  18000.0 295650.0 17100.0 326700.0 ;
      RECT  14100.0 336450.0 13200.0 337350.0 ;
      RECT  14100.0 327900.0 13200.0 336900.0 ;
      RECT  15600.0 336450.0 13650.0 337350.0 ;
      RECT  16050.0 339300.0 15150.0 346500.0 ;
      RECT  16050.0 348900.0 15150.0 356100.0 ;
      RECT  29250.0 361650.0 28350.0 362550.0 ;
      RECT  28800.0 361650.0 28350.0 362550.0 ;
      RECT  29250.0 359700.0 28350.0 362100.0 ;
      RECT  29250.0 349500.0 28350.0 356700.0 ;
      RECT  29700.0 316800.0 28800.0 323100.0 ;
      RECT  30450.0 333000.0 29550.0 340200.0 ;
      RECT  16050.0 358500.0 15150.0 362700.0 ;
      RECT  29250.0 342900.0 28350.0 347100.0 ;
      RECT  50250.0 202200.0 49350.0 362100.0 ;
      RECT  50250.0 287550.0 49350.0 308700.0 ;
      RECT  36450.0 202200.0 35550.0 362100.0 ;
      RECT  36450.0 298350.0 35550.0 308700.0 ;
      RECT  22650.0 308700.0 21750.0 362100.0 ;
      RECT  22650.0 287550.0 21750.0 308700.0 ;
      RECT  8850.0 308700.0 7950.0 362100.0 ;
      RECT  8850.0 298350.0 7950.0 308700.0 ;
      RECT  8850.0 361650.0 7950.0 362550.0 ;
      RECT  8850.0 360000.0 7950.0 362100.0 ;
      RECT  8400.0 361650.0 3600.0 362550.0 ;
      RECT  7.1054273576e-12 202200.0 10200.0 262200.0 ;
      RECT  20400.0 202200.0 10200.0 262200.0 ;
      RECT  20400.0 202200.0 30600.0 262200.0 ;
      RECT  7.1054273576e-12 204600.0 30600.0 205500.0 ;
      RECT  1.42108547152e-11 258600.0 30600.0 259500.0 ;
      RECT  37950.0 211200.0 36000.0 212400.0 ;
      RECT  49800.0 211200.0 47850.0 212400.0 ;
      RECT  48450.0 206700.0 39150.0 207600.0 ;
      RECT  38550.0 204150.0 36600.0 205050.0 ;
      RECT  38550.0 208950.0 36600.0 209850.0 ;
      RECT  39150.0 204000.0 37950.0 205200.0 ;
      RECT  39150.0 208800.0 37950.0 210000.0 ;
      RECT  39150.0 206400.0 37950.0 207600.0 ;
      RECT  39150.0 206400.0 37950.0 207600.0 ;
      RECT  37050.0 204150.0 36150.0 209850.0 ;
      RECT  49800.0 204150.0 47850.0 205050.0 ;
      RECT  49800.0 208950.0 47850.0 209850.0 ;
      RECT  48450.0 204000.0 47250.0 205200.0 ;
      RECT  48450.0 208800.0 47250.0 210000.0 ;
      RECT  48450.0 206400.0 47250.0 207600.0 ;
      RECT  48450.0 206400.0 47250.0 207600.0 ;
      RECT  50250.0 204150.0 49350.0 209850.0 ;
      RECT  38550.0 211200.0 37350.0 212400.0 ;
      RECT  48450.0 211200.0 47250.0 212400.0 ;
      RECT  43800.0 204600.0 42600.0 205800.0 ;
      RECT  43800.0 204600.0 42600.0 205800.0 ;
      RECT  43650.0 207150.0 42750.0 208050.0 ;
      RECT  36450.0 202200.0 35550.0 214200.0 ;
      RECT  50250.0 202200.0 49350.0 214200.0 ;
      RECT  37950.0 225600.0 36000.0 226800.0 ;
      RECT  49800.0 225600.0 47850.0 226800.0 ;
      RECT  37350.0 216150.0 35550.0 221850.0 ;
      RECT  46050.0 223350.0 41250.0 224250.0 ;
      RECT  38850.0 216150.0 36900.0 217050.0 ;
      RECT  38850.0 220950.0 36900.0 221850.0 ;
      RECT  40800.0 218550.0 38850.0 219450.0 ;
      RECT  40800.0 223350.0 38850.0 224250.0 ;
      RECT  39450.0 216000.0 38250.0 217200.0 ;
      RECT  39450.0 220800.0 38250.0 222000.0 ;
      RECT  39450.0 218400.0 38250.0 219600.0 ;
      RECT  39450.0 223200.0 38250.0 224400.0 ;
      RECT  41250.0 218550.0 40350.0 224250.0 ;
      RECT  37350.0 216150.0 36450.0 221850.0 ;
      RECT  49500.0 216150.0 47550.0 217050.0 ;
      RECT  49500.0 220950.0 47550.0 221850.0 ;
      RECT  47550.0 218550.0 45600.0 219450.0 ;
      RECT  47550.0 223350.0 45600.0 224250.0 ;
      RECT  48150.0 216000.0 46950.0 217200.0 ;
      RECT  48150.0 220800.0 46950.0 222000.0 ;
      RECT  48150.0 218400.0 46950.0 219600.0 ;
      RECT  48150.0 223200.0 46950.0 224400.0 ;
      RECT  46050.0 218550.0 45150.0 224250.0 ;
      RECT  49950.0 216150.0 49050.0 221850.0 ;
      RECT  38550.0 225600.0 37350.0 226800.0 ;
      RECT  48450.0 225600.0 47250.0 226800.0 ;
      RECT  43800.0 216600.0 42600.0 217800.0 ;
      RECT  43800.0 216600.0 42600.0 217800.0 ;
      RECT  43650.0 223800.0 42750.0 224700.0 ;
      RECT  36450.0 214200.0 35550.0 228600.0 ;
      RECT  50250.0 214200.0 49350.0 228600.0 ;
      RECT  37950.0 244800.0 36000.0 246000.0 ;
      RECT  49800.0 244800.0 47850.0 246000.0 ;
      RECT  37800.0 230550.0 35550.0 241050.0 ;
      RECT  45900.0 242550.0 41700.0 243450.0 ;
      RECT  39300.0 230550.0 37350.0 231450.0 ;
      RECT  39300.0 235350.0 37350.0 236250.0 ;
      RECT  39300.0 240150.0 37350.0 241050.0 ;
      RECT  41250.0 232950.0 39300.0 233850.0 ;
      RECT  41250.0 237750.0 39300.0 238650.0 ;
      RECT  41250.0 242550.0 39300.0 243450.0 ;
      RECT  39900.0 230400.0 38700.0 231600.0 ;
      RECT  39900.0 235200.0 38700.0 236400.0 ;
      RECT  39900.0 240000.0 38700.0 241200.0 ;
      RECT  39900.0 232800.0 38700.0 234000.0 ;
      RECT  39900.0 237600.0 38700.0 238800.0 ;
      RECT  39900.0 242400.0 38700.0 243600.0 ;
      RECT  41700.0 232950.0 40800.0 243450.0 ;
      RECT  37800.0 230550.0 36900.0 241050.0 ;
      RECT  49350.0 230550.0 47400.0 231450.0 ;
      RECT  49350.0 235350.0 47400.0 236250.0 ;
      RECT  49350.0 240150.0 47400.0 241050.0 ;
      RECT  47400.0 232950.0 45450.0 233850.0 ;
      RECT  47400.0 237750.0 45450.0 238650.0 ;
      RECT  47400.0 242550.0 45450.0 243450.0 ;
      RECT  48000.0 230400.0 46800.0 231600.0 ;
      RECT  48000.0 235200.0 46800.0 236400.0 ;
      RECT  48000.0 240000.0 46800.0 241200.0 ;
      RECT  48000.0 232800.0 46800.0 234000.0 ;
      RECT  48000.0 237600.0 46800.0 238800.0 ;
      RECT  48000.0 242400.0 46800.0 243600.0 ;
      RECT  45900.0 232950.0 45000.0 243450.0 ;
      RECT  49800.0 230550.0 48900.0 241050.0 ;
      RECT  38550.0 244800.0 37350.0 246000.0 ;
      RECT  48450.0 244800.0 47250.0 246000.0 ;
      RECT  43950.0 231000.0 42750.0 232200.0 ;
      RECT  43950.0 231000.0 42750.0 232200.0 ;
      RECT  43800.0 243000.0 42900.0 243900.0 ;
      RECT  36450.0 228600.0 35550.0 247800.0 ;
      RECT  50250.0 228600.0 49350.0 247800.0 ;
      RECT  37950.0 276000.0 36000.0 277200.0 ;
      RECT  49800.0 276000.0 47850.0 277200.0 ;
      RECT  37800.0 249750.0 35550.0 274650.0 ;
      RECT  45900.0 271350.0 41700.0 272250.0 ;
      RECT  39300.0 249750.0 37350.0 250650.0 ;
      RECT  39300.0 254550.0 37350.0 255450.0 ;
      RECT  39300.0 259350.0 37350.0 260250.0 ;
      RECT  39300.0 264150.0 37350.0 265050.0 ;
      RECT  39300.0 268950.0 37350.0 269850.0 ;
      RECT  39300.0 273750.0 37350.0 274650.0 ;
      RECT  41250.0 252150.0 39300.0 253050.0 ;
      RECT  41250.0 256950.0 39300.0 257850.0 ;
      RECT  41250.0 261750.0 39300.0 262650.0 ;
      RECT  41250.0 266550.0 39300.0 267450.0 ;
      RECT  41250.0 271350.0 39300.0 272250.0 ;
      RECT  39900.0 249600.0 38700.0 250800.0 ;
      RECT  39900.0 254400.0 38700.0 255600.0 ;
      RECT  39900.0 259200.0 38700.0 260400.0 ;
      RECT  39900.0 264000.0 38700.0 265200.0 ;
      RECT  39900.0 268800.0 38700.0 270000.0 ;
      RECT  39900.0 273600.0 38700.0 274800.0 ;
      RECT  39900.0 252000.0 38700.0 253200.0 ;
      RECT  39900.0 256800.0 38700.0 258000.0 ;
      RECT  39900.0 261600.0 38700.0 262800.0 ;
      RECT  39900.0 266400.0 38700.0 267600.0 ;
      RECT  39900.0 271200.0 38700.0 272400.0 ;
      RECT  41700.0 252150.0 40800.0 272250.0 ;
      RECT  37800.0 249750.0 36900.0 274650.0 ;
      RECT  49350.0 249750.0 47400.0 250650.0 ;
      RECT  49350.0 254550.0 47400.0 255450.0 ;
      RECT  49350.0 259350.0 47400.0 260250.0 ;
      RECT  49350.0 264150.0 47400.0 265050.0 ;
      RECT  49350.0 268950.0 47400.0 269850.0 ;
      RECT  49350.0 273750.0 47400.0 274650.0 ;
      RECT  47400.0 252150.0 45450.0 253050.0 ;
      RECT  47400.0 256950.0 45450.0 257850.0 ;
      RECT  47400.0 261750.0 45450.0 262650.0 ;
      RECT  47400.0 266550.0 45450.0 267450.0 ;
      RECT  47400.0 271350.0 45450.0 272250.0 ;
      RECT  48000.0 249600.0 46800.0 250800.0 ;
      RECT  48000.0 254400.0 46800.0 255600.0 ;
      RECT  48000.0 259200.0 46800.0 260400.0 ;
      RECT  48000.0 264000.0 46800.0 265200.0 ;
      RECT  48000.0 268800.0 46800.0 270000.0 ;
      RECT  48000.0 273600.0 46800.0 274800.0 ;
      RECT  48000.0 252000.0 46800.0 253200.0 ;
      RECT  48000.0 256800.0 46800.0 258000.0 ;
      RECT  48000.0 261600.0 46800.0 262800.0 ;
      RECT  48000.0 266400.0 46800.0 267600.0 ;
      RECT  48000.0 271200.0 46800.0 272400.0 ;
      RECT  45900.0 252150.0 45000.0 272250.0 ;
      RECT  49800.0 249750.0 48900.0 274650.0 ;
      RECT  38550.0 276000.0 37350.0 277200.0 ;
      RECT  48450.0 276000.0 47250.0 277200.0 ;
      RECT  43950.0 250200.0 42750.0 251400.0 ;
      RECT  43950.0 250200.0 42750.0 251400.0 ;
      RECT  43800.0 271800.0 42900.0 272700.0 ;
      RECT  36450.0 247800.0 35550.0 279000.0 ;
      RECT  50250.0 247800.0 49350.0 279000.0 ;
      RECT  47850.0 310500.0 50250.0 311700.0 ;
      RECT  39150.0 310500.0 35550.0 311700.0 ;
      RECT  39150.0 315300.0 35550.0 316500.0 ;
      RECT  37950.0 320100.0 36000.0 321300.0 ;
      RECT  49800.0 320100.0 47850.0 321300.0 ;
      RECT  39150.0 310500.0 37950.0 311700.0 ;
      RECT  39150.0 312900.0 37950.0 314100.0 ;
      RECT  39150.0 312900.0 37950.0 314100.0 ;
      RECT  39150.0 310500.0 37950.0 311700.0 ;
      RECT  39150.0 312900.0 37950.0 314100.0 ;
      RECT  39150.0 315300.0 37950.0 316500.0 ;
      RECT  39150.0 315300.0 37950.0 316500.0 ;
      RECT  39150.0 312900.0 37950.0 314100.0 ;
      RECT  39150.0 315300.0 37950.0 316500.0 ;
      RECT  39150.0 317700.0 37950.0 318900.0 ;
      RECT  39150.0 317700.0 37950.0 318900.0 ;
      RECT  39150.0 315300.0 37950.0 316500.0 ;
      RECT  47850.0 310500.0 46650.0 311700.0 ;
      RECT  47850.0 312900.0 46650.0 314100.0 ;
      RECT  47850.0 312900.0 46650.0 314100.0 ;
      RECT  47850.0 310500.0 46650.0 311700.0 ;
      RECT  47850.0 312900.0 46650.0 314100.0 ;
      RECT  47850.0 315300.0 46650.0 316500.0 ;
      RECT  47850.0 315300.0 46650.0 316500.0 ;
      RECT  47850.0 312900.0 46650.0 314100.0 ;
      RECT  47850.0 315300.0 46650.0 316500.0 ;
      RECT  47850.0 317700.0 46650.0 318900.0 ;
      RECT  47850.0 317700.0 46650.0 318900.0 ;
      RECT  47850.0 315300.0 46650.0 316500.0 ;
      RECT  38550.0 320100.0 37350.0 321300.0 ;
      RECT  48450.0 320100.0 47250.0 321300.0 ;
      RECT  45750.0 317700.0 44550.0 316500.0 ;
      RECT  43800.0 315300.0 42600.0 314100.0 ;
      RECT  41850.0 312900.0 40650.0 311700.0 ;
      RECT  39150.0 312900.0 37950.0 314100.0 ;
      RECT  39150.0 317700.0 37950.0 318900.0 ;
      RECT  47850.0 317700.0 46650.0 318900.0 ;
      RECT  41850.0 317700.0 40650.0 318900.0 ;
      RECT  41850.0 311700.0 40650.0 312900.0 ;
      RECT  43800.0 314100.0 42600.0 315300.0 ;
      RECT  45750.0 316500.0 44550.0 317700.0 ;
      RECT  41850.0 317700.0 40650.0 318900.0 ;
      RECT  36450.0 308700.0 35550.0 324300.0 ;
      RECT  50250.0 308700.0 49350.0 324300.0 ;
      RECT  37950.0 330900.0 36000.0 332100.0 ;
      RECT  49800.0 330900.0 47850.0 332100.0 ;
      RECT  48450.0 326100.0 50250.0 327300.0 ;
      RECT  39150.0 326100.0 35550.0 327300.0 ;
      RECT  48450.0 328800.0 39150.0 329700.0 ;
      RECT  39150.0 326100.0 37950.0 327300.0 ;
      RECT  39150.0 328500.0 37950.0 329700.0 ;
      RECT  39150.0 328500.0 37950.0 329700.0 ;
      RECT  39150.0 326100.0 37950.0 327300.0 ;
      RECT  48450.0 326100.0 47250.0 327300.0 ;
      RECT  48450.0 328500.0 47250.0 329700.0 ;
      RECT  48450.0 328500.0 47250.0 329700.0 ;
      RECT  48450.0 326100.0 47250.0 327300.0 ;
      RECT  38550.0 330900.0 37350.0 332100.0 ;
      RECT  48450.0 330900.0 47250.0 332100.0 ;
      RECT  43800.0 326700.0 42600.0 327900.0 ;
      RECT  43800.0 326700.0 42600.0 327900.0 ;
      RECT  43650.0 329250.0 42750.0 330150.0 ;
      RECT  36450.0 324300.0 35550.0 333900.0 ;
      RECT  50250.0 324300.0 49350.0 333900.0 ;
      RECT  23550.0 310500.0 21750.0 311700.0 ;
      RECT  23550.0 315300.0 21750.0 316500.0 ;
      RECT  32250.0 310500.0 36450.0 311700.0 ;
      RECT  34050.0 317700.0 36000.0 318900.0 ;
      RECT  22200.0 317700.0 24150.0 318900.0 ;
      RECT  32250.0 310500.0 33450.0 311700.0 ;
      RECT  32250.0 312900.0 33450.0 314100.0 ;
      RECT  32250.0 312900.0 33450.0 314100.0 ;
      RECT  32250.0 310500.0 33450.0 311700.0 ;
      RECT  32250.0 312900.0 33450.0 314100.0 ;
      RECT  32250.0 315300.0 33450.0 316500.0 ;
      RECT  32250.0 315300.0 33450.0 316500.0 ;
      RECT  32250.0 312900.0 33450.0 314100.0 ;
      RECT  23550.0 310500.0 24750.0 311700.0 ;
      RECT  23550.0 312900.0 24750.0 314100.0 ;
      RECT  23550.0 312900.0 24750.0 314100.0 ;
      RECT  23550.0 310500.0 24750.0 311700.0 ;
      RECT  23550.0 312900.0 24750.0 314100.0 ;
      RECT  23550.0 315300.0 24750.0 316500.0 ;
      RECT  23550.0 315300.0 24750.0 316500.0 ;
      RECT  23550.0 312900.0 24750.0 314100.0 ;
      RECT  33450.0 317700.0 34650.0 318900.0 ;
      RECT  23550.0 317700.0 24750.0 318900.0 ;
      RECT  25950.0 315300.0 27150.0 314100.0 ;
      RECT  28650.0 312300.0 29850.0 311100.0 ;
      RECT  32250.0 315300.0 33450.0 316500.0 ;
      RECT  23550.0 314100.0 24750.0 312900.0 ;
      RECT  28650.0 317400.0 29850.0 316200.0 ;
      RECT  28650.0 311100.0 29850.0 312300.0 ;
      RECT  25950.0 314100.0 27150.0 315300.0 ;
      RECT  28650.0 316200.0 29850.0 317400.0 ;
      RECT  35550.0 308700.0 36450.0 323100.0 ;
      RECT  21750.0 308700.0 22650.0 323100.0 ;
      RECT  24150.0 327600.0 21750.0 328800.0 ;
      RECT  32850.0 327600.0 36450.0 328800.0 ;
      RECT  32850.0 332400.0 36450.0 333600.0 ;
      RECT  34050.0 334800.0 36000.0 336000.0 ;
      RECT  22200.0 334800.0 24150.0 336000.0 ;
      RECT  32850.0 327600.0 34050.0 328800.0 ;
      RECT  32850.0 330000.0 34050.0 331200.0 ;
      RECT  32850.0 330000.0 34050.0 331200.0 ;
      RECT  32850.0 327600.0 34050.0 328800.0 ;
      RECT  32850.0 330000.0 34050.0 331200.0 ;
      RECT  32850.0 332400.0 34050.0 333600.0 ;
      RECT  32850.0 332400.0 34050.0 333600.0 ;
      RECT  32850.0 330000.0 34050.0 331200.0 ;
      RECT  24150.0 327600.0 25350.0 328800.0 ;
      RECT  24150.0 330000.0 25350.0 331200.0 ;
      RECT  24150.0 330000.0 25350.0 331200.0 ;
      RECT  24150.0 327600.0 25350.0 328800.0 ;
      RECT  24150.0 330000.0 25350.0 331200.0 ;
      RECT  24150.0 332400.0 25350.0 333600.0 ;
      RECT  24150.0 332400.0 25350.0 333600.0 ;
      RECT  24150.0 330000.0 25350.0 331200.0 ;
      RECT  33450.0 334800.0 34650.0 336000.0 ;
      RECT  23550.0 334800.0 24750.0 336000.0 ;
      RECT  26700.0 332400.0 27900.0 331200.0 ;
      RECT  29400.0 329400.0 30600.0 328200.0 ;
      RECT  32850.0 330000.0 34050.0 331200.0 ;
      RECT  24150.0 332400.0 25350.0 333600.0 ;
      RECT  29400.0 333600.0 30600.0 332400.0 ;
      RECT  29400.0 328200.0 30600.0 329400.0 ;
      RECT  26700.0 331200.0 27900.0 332400.0 ;
      RECT  29400.0 332400.0 30600.0 333600.0 ;
      RECT  35550.0 325800.0 36450.0 340200.0 ;
      RECT  21750.0 325800.0 22650.0 340200.0 ;
      RECT  34050.0 345900.0 36000.0 344700.0 ;
      RECT  22200.0 345900.0 24150.0 344700.0 ;
      RECT  23550.0 350700.0 21750.0 349500.0 ;
      RECT  32850.0 350700.0 36450.0 349500.0 ;
      RECT  23550.0 348000.0 32850.0 347100.0 ;
      RECT  32850.0 350700.0 34050.0 349500.0 ;
      RECT  32850.0 348300.0 34050.0 347100.0 ;
      RECT  32850.0 348300.0 34050.0 347100.0 ;
      RECT  32850.0 350700.0 34050.0 349500.0 ;
      RECT  23550.0 350700.0 24750.0 349500.0 ;
      RECT  23550.0 348300.0 24750.0 347100.0 ;
      RECT  23550.0 348300.0 24750.0 347100.0 ;
      RECT  23550.0 350700.0 24750.0 349500.0 ;
      RECT  33450.0 345900.0 34650.0 344700.0 ;
      RECT  23550.0 345900.0 24750.0 344700.0 ;
      RECT  28200.0 350100.0 29400.0 348900.0 ;
      RECT  28200.0 350100.0 29400.0 348900.0 ;
      RECT  28350.0 347550.0 29250.0 346650.0 ;
      RECT  35550.0 352500.0 36450.0 342900.0 ;
      RECT  21750.0 352500.0 22650.0 342900.0 ;
      RECT  34050.0 355500.0 36000.0 354300.0 ;
      RECT  22200.0 355500.0 24150.0 354300.0 ;
      RECT  23550.0 360300.0 21750.0 359100.0 ;
      RECT  32850.0 360300.0 36450.0 359100.0 ;
      RECT  23550.0 357600.0 32850.0 356700.0 ;
      RECT  32850.0 360300.0 34050.0 359100.0 ;
      RECT  32850.0 357900.0 34050.0 356700.0 ;
      RECT  32850.0 357900.0 34050.0 356700.0 ;
      RECT  32850.0 360300.0 34050.0 359100.0 ;
      RECT  23550.0 360300.0 24750.0 359100.0 ;
      RECT  23550.0 357900.0 24750.0 356700.0 ;
      RECT  23550.0 357900.0 24750.0 356700.0 ;
      RECT  23550.0 360300.0 24750.0 359100.0 ;
      RECT  33450.0 355500.0 34650.0 354300.0 ;
      RECT  23550.0 355500.0 24750.0 354300.0 ;
      RECT  28200.0 359700.0 29400.0 358500.0 ;
      RECT  28200.0 359700.0 29400.0 358500.0 ;
      RECT  28350.0 357150.0 29250.0 356250.0 ;
      RECT  35550.0 362100.0 36450.0 352500.0 ;
      RECT  21750.0 362100.0 22650.0 352500.0 ;
      RECT  20250.0 320100.0 22650.0 321300.0 ;
      RECT  11550.0 320100.0 7950.0 321300.0 ;
      RECT  11550.0 324900.0 7950.0 326100.0 ;
      RECT  10350.0 329700.0 8400.0 330900.0 ;
      RECT  22200.0 329700.0 20250.0 330900.0 ;
      RECT  11550.0 320100.0 10350.0 321300.0 ;
      RECT  11550.0 322500.0 10350.0 323700.0 ;
      RECT  11550.0 322500.0 10350.0 323700.0 ;
      RECT  11550.0 320100.0 10350.0 321300.0 ;
      RECT  11550.0 322500.0 10350.0 323700.0 ;
      RECT  11550.0 324900.0 10350.0 326100.0 ;
      RECT  11550.0 324900.0 10350.0 326100.0 ;
      RECT  11550.0 322500.0 10350.0 323700.0 ;
      RECT  11550.0 324900.0 10350.0 326100.0 ;
      RECT  11550.0 327300.0 10350.0 328500.0 ;
      RECT  11550.0 327300.0 10350.0 328500.0 ;
      RECT  11550.0 324900.0 10350.0 326100.0 ;
      RECT  20250.0 320100.0 19050.0 321300.0 ;
      RECT  20250.0 322500.0 19050.0 323700.0 ;
      RECT  20250.0 322500.0 19050.0 323700.0 ;
      RECT  20250.0 320100.0 19050.0 321300.0 ;
      RECT  20250.0 322500.0 19050.0 323700.0 ;
      RECT  20250.0 324900.0 19050.0 326100.0 ;
      RECT  20250.0 324900.0 19050.0 326100.0 ;
      RECT  20250.0 322500.0 19050.0 323700.0 ;
      RECT  20250.0 324900.0 19050.0 326100.0 ;
      RECT  20250.0 327300.0 19050.0 328500.0 ;
      RECT  20250.0 327300.0 19050.0 328500.0 ;
      RECT  20250.0 324900.0 19050.0 326100.0 ;
      RECT  10950.0 329700.0 9750.0 330900.0 ;
      RECT  20850.0 329700.0 19650.0 330900.0 ;
      RECT  18150.0 327300.0 16950.0 326100.0 ;
      RECT  16200.0 324900.0 15000.0 323700.0 ;
      RECT  14250.0 322500.0 13050.0 321300.0 ;
      RECT  11550.0 322500.0 10350.0 323700.0 ;
      RECT  11550.0 327300.0 10350.0 328500.0 ;
      RECT  20250.0 327300.0 19050.0 328500.0 ;
      RECT  14250.0 327300.0 13050.0 328500.0 ;
      RECT  14250.0 321300.0 13050.0 322500.0 ;
      RECT  16200.0 323700.0 15000.0 324900.0 ;
      RECT  18150.0 326100.0 16950.0 327300.0 ;
      RECT  14250.0 327300.0 13050.0 328500.0 ;
      RECT  8850.0 318300.0 7950.0 333900.0 ;
      RECT  22650.0 318300.0 21750.0 333900.0 ;
      RECT  10350.0 340500.0 8400.0 341700.0 ;
      RECT  22200.0 340500.0 20250.0 341700.0 ;
      RECT  20850.0 335700.0 22650.0 336900.0 ;
      RECT  11550.0 335700.0 7950.0 336900.0 ;
      RECT  20850.0 338400.0 11550.0 339300.0 ;
      RECT  11550.0 335700.0 10350.0 336900.0 ;
      RECT  11550.0 338100.0 10350.0 339300.0 ;
      RECT  11550.0 338100.0 10350.0 339300.0 ;
      RECT  11550.0 335700.0 10350.0 336900.0 ;
      RECT  20850.0 335700.0 19650.0 336900.0 ;
      RECT  20850.0 338100.0 19650.0 339300.0 ;
      RECT  20850.0 338100.0 19650.0 339300.0 ;
      RECT  20850.0 335700.0 19650.0 336900.0 ;
      RECT  10950.0 340500.0 9750.0 341700.0 ;
      RECT  20850.0 340500.0 19650.0 341700.0 ;
      RECT  16200.0 336300.0 15000.0 337500.0 ;
      RECT  16200.0 336300.0 15000.0 337500.0 ;
      RECT  16050.0 338850.0 15150.0 339750.0 ;
      RECT  8850.0 333900.0 7950.0 343500.0 ;
      RECT  22650.0 333900.0 21750.0 343500.0 ;
      RECT  10350.0 350100.0 8400.0 351300.0 ;
      RECT  22200.0 350100.0 20250.0 351300.0 ;
      RECT  20850.0 345300.0 22650.0 346500.0 ;
      RECT  11550.0 345300.0 7950.0 346500.0 ;
      RECT  20850.0 348000.0 11550.0 348900.0 ;
      RECT  11550.0 345300.0 10350.0 346500.0 ;
      RECT  11550.0 347700.0 10350.0 348900.0 ;
      RECT  11550.0 347700.0 10350.0 348900.0 ;
      RECT  11550.0 345300.0 10350.0 346500.0 ;
      RECT  20850.0 345300.0 19650.0 346500.0 ;
      RECT  20850.0 347700.0 19650.0 348900.0 ;
      RECT  20850.0 347700.0 19650.0 348900.0 ;
      RECT  20850.0 345300.0 19650.0 346500.0 ;
      RECT  10950.0 350100.0 9750.0 351300.0 ;
      RECT  20850.0 350100.0 19650.0 351300.0 ;
      RECT  16200.0 345900.0 15000.0 347100.0 ;
      RECT  16200.0 345900.0 15000.0 347100.0 ;
      RECT  16050.0 348450.0 15150.0 349350.0 ;
      RECT  8850.0 343500.0 7950.0 353100.0 ;
      RECT  22650.0 343500.0 21750.0 353100.0 ;
      RECT  10350.0 359700.0 8400.0 360900.0 ;
      RECT  22200.0 359700.0 20250.0 360900.0 ;
      RECT  20850.0 354900.0 22650.0 356100.0 ;
      RECT  11550.0 354900.0 7950.0 356100.0 ;
      RECT  20850.0 357600.0 11550.0 358500.0 ;
      RECT  11550.0 354900.0 10350.0 356100.0 ;
      RECT  11550.0 357300.0 10350.0 358500.0 ;
      RECT  11550.0 357300.0 10350.0 358500.0 ;
      RECT  11550.0 354900.0 10350.0 356100.0 ;
      RECT  20850.0 354900.0 19650.0 356100.0 ;
      RECT  20850.0 357300.0 19650.0 358500.0 ;
      RECT  20850.0 357300.0 19650.0 358500.0 ;
      RECT  20850.0 354900.0 19650.0 356100.0 ;
      RECT  10950.0 359700.0 9750.0 360900.0 ;
      RECT  20850.0 359700.0 19650.0 360900.0 ;
      RECT  16200.0 355500.0 15000.0 356700.0 ;
      RECT  16200.0 355500.0 15000.0 356700.0 ;
      RECT  16050.0 358050.0 15150.0 358950.0 ;
      RECT  8850.0 353100.0 7950.0 362700.0 ;
      RECT  22650.0 353100.0 21750.0 362700.0 ;
      RECT  22650.0 396600.0 16800.0 397500.0 ;
      RECT  22650.0 420000.0 16800.0 420900.0 ;
      RECT  22200.0 425550.0 16800.0 426450.0 ;
      RECT  4500.0 408300.0 16800.0 409200.0 ;
      RECT  4500.0 380700.0 16800.0 381600.0 ;
      RECT  29250.0 397500.0 28350.0 410100.0 ;
      RECT  29250.0 392550.0 28350.0 393450.0 ;
      RECT  29250.0 393000.0 28350.0 397500.0 ;
      RECT  28800.0 392550.0 17400.0 393450.0 ;
      RECT  36000.0 398250.0 33750.0 399150.0 ;
      RECT  33600.0 383550.0 32700.0 384450.0 ;
      RECT  29250.0 383550.0 28350.0 384450.0 ;
      RECT  33600.0 384000.0 32700.0 395700.0 ;
      RECT  33150.0 383550.0 28800.0 384450.0 ;
      RECT  29250.0 378900.0 28350.0 384000.0 ;
      RECT  28800.0 383550.0 19950.0 384450.0 ;
      RECT  19950.0 375450.0 13200.0 376350.0 ;
      RECT  29400.0 377700.0 28200.0 378900.0 ;
      RECT  29250.0 410100.0 28350.0 413850.0 ;
      RECT  34050.0 374700.0 36000.0 373500.0 ;
      RECT  22200.0 374700.0 24150.0 373500.0 ;
      RECT  23550.0 379500.0 21750.0 378300.0 ;
      RECT  32850.0 379500.0 36450.0 378300.0 ;
      RECT  23550.0 376800.0 32850.0 375900.0 ;
      RECT  32850.0 379500.0 34050.0 378300.0 ;
      RECT  32850.0 377100.0 34050.0 375900.0 ;
      RECT  32850.0 377100.0 34050.0 375900.0 ;
      RECT  32850.0 379500.0 34050.0 378300.0 ;
      RECT  23550.0 379500.0 24750.0 378300.0 ;
      RECT  23550.0 377100.0 24750.0 375900.0 ;
      RECT  23550.0 377100.0 24750.0 375900.0 ;
      RECT  23550.0 379500.0 24750.0 378300.0 ;
      RECT  33450.0 374700.0 34650.0 373500.0 ;
      RECT  23550.0 374700.0 24750.0 373500.0 ;
      RECT  28200.0 378900.0 29400.0 377700.0 ;
      RECT  28200.0 378900.0 29400.0 377700.0 ;
      RECT  28350.0 376350.0 29250.0 375450.0 ;
      RECT  35550.0 381300.0 36450.0 371700.0 ;
      RECT  21750.0 381300.0 22650.0 371700.0 ;
      RECT  32550.0 395700.0 33750.0 396900.0 ;
      RECT  32550.0 398100.0 33750.0 399300.0 ;
      RECT  32550.0 398100.0 33750.0 399300.0 ;
      RECT  32550.0 395700.0 33750.0 396900.0 ;
      RECT  21750.0 430650.0 22650.0 431550.0 ;
      RECT  49350.0 430650.0 50250.0 431550.0 ;
      RECT  21750.0 429300.0 22650.0 431100.0 ;
      RECT  22200.0 430650.0 49800.0 431550.0 ;
      RECT  49350.0 429300.0 50250.0 431100.0 ;
      RECT  37950.0 416700.0 36000.0 417900.0 ;
      RECT  49800.0 416700.0 47850.0 417900.0 ;
      RECT  48450.0 411900.0 50250.0 413100.0 ;
      RECT  39150.0 411900.0 35550.0 413100.0 ;
      RECT  48450.0 414600.0 39150.0 415500.0 ;
      RECT  39150.0 411900.0 37950.0 413100.0 ;
      RECT  39150.0 414300.0 37950.0 415500.0 ;
      RECT  39150.0 414300.0 37950.0 415500.0 ;
      RECT  39150.0 411900.0 37950.0 413100.0 ;
      RECT  48450.0 411900.0 47250.0 413100.0 ;
      RECT  48450.0 414300.0 47250.0 415500.0 ;
      RECT  48450.0 414300.0 47250.0 415500.0 ;
      RECT  48450.0 411900.0 47250.0 413100.0 ;
      RECT  38550.0 416700.0 37350.0 417900.0 ;
      RECT  48450.0 416700.0 47250.0 417900.0 ;
      RECT  43800.0 412500.0 42600.0 413700.0 ;
      RECT  43800.0 412500.0 42600.0 413700.0 ;
      RECT  43650.0 415050.0 42750.0 415950.0 ;
      RECT  36450.0 410100.0 35550.0 419700.0 ;
      RECT  50250.0 410100.0 49350.0 419700.0 ;
      RECT  37950.0 426300.0 36000.0 427500.0 ;
      RECT  49800.0 426300.0 47850.0 427500.0 ;
      RECT  48450.0 421500.0 50250.0 422700.0 ;
      RECT  39150.0 421500.0 35550.0 422700.0 ;
      RECT  48450.0 424200.0 39150.0 425100.0 ;
      RECT  39150.0 421500.0 37950.0 422700.0 ;
      RECT  39150.0 423900.0 37950.0 425100.0 ;
      RECT  39150.0 423900.0 37950.0 425100.0 ;
      RECT  39150.0 421500.0 37950.0 422700.0 ;
      RECT  48450.0 421500.0 47250.0 422700.0 ;
      RECT  48450.0 423900.0 47250.0 425100.0 ;
      RECT  48450.0 423900.0 47250.0 425100.0 ;
      RECT  48450.0 421500.0 47250.0 422700.0 ;
      RECT  38550.0 426300.0 37350.0 427500.0 ;
      RECT  48450.0 426300.0 47250.0 427500.0 ;
      RECT  43800.0 422100.0 42600.0 423300.0 ;
      RECT  43800.0 422100.0 42600.0 423300.0 ;
      RECT  43650.0 424650.0 42750.0 425550.0 ;
      RECT  36450.0 419700.0 35550.0 429300.0 ;
      RECT  50250.0 419700.0 49350.0 429300.0 ;
      RECT  42600.0 422100.0 43800.0 423300.0 ;
      RECT  34050.0 422700.0 36000.0 421500.0 ;
      RECT  22200.0 422700.0 24150.0 421500.0 ;
      RECT  23550.0 427500.0 21750.0 426300.0 ;
      RECT  32850.0 427500.0 36450.0 426300.0 ;
      RECT  23550.0 424800.0 32850.0 423900.0 ;
      RECT  32850.0 427500.0 34050.0 426300.0 ;
      RECT  32850.0 425100.0 34050.0 423900.0 ;
      RECT  32850.0 425100.0 34050.0 423900.0 ;
      RECT  32850.0 427500.0 34050.0 426300.0 ;
      RECT  23550.0 427500.0 24750.0 426300.0 ;
      RECT  23550.0 425100.0 24750.0 423900.0 ;
      RECT  23550.0 425100.0 24750.0 423900.0 ;
      RECT  23550.0 427500.0 24750.0 426300.0 ;
      RECT  33450.0 422700.0 34650.0 421500.0 ;
      RECT  23550.0 422700.0 24750.0 421500.0 ;
      RECT  28200.0 426900.0 29400.0 425700.0 ;
      RECT  28200.0 426900.0 29400.0 425700.0 ;
      RECT  28350.0 424350.0 29250.0 423450.0 ;
      RECT  35550.0 429300.0 36450.0 419700.0 ;
      RECT  21750.0 429300.0 22650.0 419700.0 ;
      RECT  28200.0 425700.0 29400.0 426900.0 ;
      RECT  34050.0 413100.0 36000.0 411900.0 ;
      RECT  22200.0 413100.0 24150.0 411900.0 ;
      RECT  23550.0 417900.0 21750.0 416700.0 ;
      RECT  32850.0 417900.0 36450.0 416700.0 ;
      RECT  23550.0 415200.0 32850.0 414300.0 ;
      RECT  32850.0 417900.0 34050.0 416700.0 ;
      RECT  32850.0 415500.0 34050.0 414300.0 ;
      RECT  32850.0 415500.0 34050.0 414300.0 ;
      RECT  32850.0 417900.0 34050.0 416700.0 ;
      RECT  23550.0 417900.0 24750.0 416700.0 ;
      RECT  23550.0 415500.0 24750.0 414300.0 ;
      RECT  23550.0 415500.0 24750.0 414300.0 ;
      RECT  23550.0 417900.0 24750.0 416700.0 ;
      RECT  33450.0 413100.0 34650.0 411900.0 ;
      RECT  23550.0 413100.0 24750.0 411900.0 ;
      RECT  28200.0 417300.0 29400.0 416100.0 ;
      RECT  28200.0 417300.0 29400.0 416100.0 ;
      RECT  28350.0 414750.0 29250.0 413850.0 ;
      RECT  35550.0 419700.0 36450.0 410100.0 ;
      RECT  21750.0 419700.0 22650.0 410100.0 ;
      RECT  28200.0 416100.0 29400.0 417300.0 ;
      RECT  42600.0 414900.0 43800.0 416100.0 ;
      RECT  42600.0 424500.0 43800.0 425700.0 ;
      RECT  28200.0 423300.0 29400.0 424500.0 ;
      RECT  42600.0 412500.0 43800.0 413700.0 ;
      RECT  28350.0 410100.0 29250.0 413850.0 ;
      RECT  35550.0 410100.0 36450.0 429300.0 ;
      RECT  21750.0 410100.0 22650.0 429300.0 ;
      RECT  49350.0 410100.0 50250.0 429300.0 ;
      RECT  16800.0 395100.0 6600.0 381300.0 ;
      RECT  16800.0 395100.0 6600.0 408900.0 ;
      RECT  16800.0 422700.0 6600.0 408900.0 ;
      RECT  17400.0 396600.0 6000.0 397800.0 ;
      RECT  17400.0 420000.0 6000.0 421200.0 ;
      RECT  17400.0 408300.0 6000.0 409200.0 ;
      RECT  22650.0 396600.0 21450.0 397800.0 ;
      RECT  22650.0 420000.0 21450.0 421200.0 ;
      RECT  22650.0 410100.0 21450.0 411300.0 ;
      RECT  22650.0 370500.0 21450.0 371700.0 ;
      RECT  21600.0 425400.0 22800.0 426600.0 ;
      RECT  16200.0 425400.0 17400.0 426600.0 ;
      RECT  29400.0 396900.0 28200.0 398100.0 ;
      RECT  19350.0 383400.0 20550.0 384600.0 ;
      RECT  19350.0 375300.0 20550.0 376500.0 ;
      RECT  12600.0 375300.0 13800.0 376500.0 ;
      RECT  43800.0 362100.0 42900.0 412500.0 ;
      RECT  29250.0 362100.0 28350.0 375450.0 ;
      RECT  4500.0 362100.0 3600.0 423150.0 ;
      RECT  36450.0 362100.0 35550.0 410100.0 ;
      RECT  22650.0 362100.0 21750.0 381300.0 ;
      RECT  50250.0 362100.0 49350.0 410100.0 ;
      RECT  43950.0 285450.0 42750.0 284250.0 ;
      RECT  43950.0 244500.0 42750.0 243300.0 ;
      RECT  33900.0 205650.0 32700.0 204450.0 ;
      RECT  29850.0 285450.0 28650.0 284250.0 ;
      RECT  27150.0 290850.0 25950.0 289650.0 ;
      RECT  30600.0 328200.0 29400.0 327000.0 ;
      RECT  27900.0 331200.0 26700.0 330000.0 ;
      RECT  41850.0 304350.0 40650.0 303150.0 ;
      RECT  43800.0 301650.0 42600.0 300450.0 ;
      RECT  45750.0 293550.0 44550.0 292350.0 ;
      RECT  14250.0 304350.0 13050.0 303150.0 ;
      RECT  16200.0 293550.0 15000.0 292350.0 ;
      RECT  18150.0 296250.0 16950.0 295050.0 ;
      RECT  29850.0 322500.0 28650.0 323700.0 ;
      RECT  30600.0 339600.0 29400.0 340800.0 ;
      RECT  16200.0 362100.0 15000.0 363300.0 ;
      RECT  29400.0 342300.0 28200.0 343500.0 ;
      RECT  50400.0 288150.0 49200.0 286950.0 ;
      RECT  36600.0 298950.0 35400.0 297750.0 ;
      RECT  22800.0 288150.0 21600.0 286950.0 ;
      RECT  9000.0 298950.0 7800.0 297750.0 ;
      RECT  43800.0 202200.0 42600.0 205800.0 ;
      RECT  36450.0 202200.0 35550.0 203100.0 ;
      RECT  50250.0 202200.0 49350.0 203100.0 ;
      RECT  55650.0 297750.0 54450.0 298950.0 ;
   LAYER  metal2 ;
      RECT  168750.0 340200.0 169650.0 342900.0 ;
      RECT  166050.0 360000.0 166950.0 362700.0 ;
      RECT  160650.0 320400.0 161550.0 323100.0 ;
      RECT  157950.0 337500.0 158850.0 340200.0 ;
      RECT  163350.0 301050.0 164250.0 303750.0 ;
      RECT  155250.0 282150.0 156150.0 284850.0 ;
      RECT  49800.0 297900.0 55050.0 298800.0 ;
      RECT  149850.0 284850.0 150750.0 287550.0 ;
      RECT  155250.0 0.0 156150.0 436800.0 ;
      RECT  157950.0 0.0 158850.0 436800.0 ;
      RECT  160650.0 0.0 161550.0 436800.0 ;
      RECT  163350.0 0.0 164250.0 436800.0 ;
      RECT  166050.0 0.0 166950.0 436800.0 ;
      RECT  168750.0 0.0 169650.0 436800.0 ;
      RECT  134550.0 37200.0 135450.0 199200.0 ;
      RECT  137250.0 37200.0 138150.0 199200.0 ;
      RECT  139950.0 37200.0 140850.0 199200.0 ;
      RECT  142650.0 37200.0 143550.0 199200.0 ;
      RECT  178650.0 420000.0 179550.0 421800.0 ;
      RECT  181650.0 420000.0 182550.0 420600.0 ;
      RECT  188850.0 420000.0 189750.0 421800.0 ;
      RECT  191850.0 420000.0 192750.0 420600.0 ;
      RECT  180150.0 5850.0 181050.0 6750.0 ;
      RECT  177000.0 5850.0 180600.0 6750.0 ;
      RECT  180150.0 6300.0 181050.0 8100.0 ;
      RECT  190350.0 5850.0 191250.0 6750.0 ;
      RECT  187200.0 5850.0 190800.0 6750.0 ;
      RECT  190350.0 6300.0 191250.0 8100.0 ;
      RECT  102600.0 420000.0 103500.0 422100.0 ;
      RECT  175500.0 199200.0 185700.0 213000.0 ;
      RECT  175500.0 226800.0 185700.0 213000.0 ;
      RECT  175500.0 226800.0 185700.0 240600.0 ;
      RECT  175500.0 254400.0 185700.0 240600.0 ;
      RECT  175500.0 254400.0 185700.0 268200.0 ;
      RECT  175500.0 282000.0 185700.0 268200.0 ;
      RECT  175500.0 282000.0 185700.0 295800.0 ;
      RECT  175500.0 309600.0 185700.0 295800.0 ;
      RECT  175500.0 309600.0 185700.0 323400.0 ;
      RECT  175500.0 337200.0 185700.0 323400.0 ;
      RECT  175500.0 337200.0 185700.0 351000.0 ;
      RECT  175500.0 364800.0 185700.0 351000.0 ;
      RECT  175500.0 364800.0 185700.0 378600.0 ;
      RECT  175500.0 392400.0 185700.0 378600.0 ;
      RECT  175500.0 392400.0 185700.0 406200.0 ;
      RECT  175500.0 420000.0 185700.0 406200.0 ;
      RECT  185700.0 199200.0 195900.0 213000.0 ;
      RECT  185700.0 226800.0 195900.0 213000.0 ;
      RECT  185700.0 226800.0 195900.0 240600.0 ;
      RECT  185700.0 254400.0 195900.0 240600.0 ;
      RECT  185700.0 254400.0 195900.0 268200.0 ;
      RECT  185700.0 282000.0 195900.0 268200.0 ;
      RECT  185700.0 282000.0 195900.0 295800.0 ;
      RECT  185700.0 309600.0 195900.0 295800.0 ;
      RECT  185700.0 309600.0 195900.0 323400.0 ;
      RECT  185700.0 337200.0 195900.0 323400.0 ;
      RECT  185700.0 337200.0 195900.0 351000.0 ;
      RECT  185700.0 364800.0 195900.0 351000.0 ;
      RECT  185700.0 364800.0 195900.0 378600.0 ;
      RECT  185700.0 392400.0 195900.0 378600.0 ;
      RECT  185700.0 392400.0 195900.0 406200.0 ;
      RECT  185700.0 420000.0 195900.0 406200.0 ;
      RECT  178500.0 199800.0 179700.0 421800.0 ;
      RECT  181500.0 198600.0 182700.0 420600.0 ;
      RECT  188700.0 199800.0 189900.0 421800.0 ;
      RECT  191700.0 198600.0 192900.0 420600.0 ;
      RECT  174900.0 198600.0 176100.0 420600.0 ;
      RECT  185100.0 198600.0 186300.0 420600.0 ;
      RECT  195300.0 198600.0 196500.0 420600.0 ;
      RECT  178500.0 422400.0 179700.0 423600.0 ;
      RECT  180900.0 422400.0 182550.0 423600.0 ;
      RECT  178500.0 429600.0 179700.0 430800.0 ;
      RECT  181650.0 429600.0 184500.0 430800.0 ;
      RECT  178500.0 422400.0 179700.0 423600.0 ;
      RECT  180900.0 422400.0 182100.0 423600.0 ;
      RECT  178500.0 429600.0 179700.0 430800.0 ;
      RECT  183300.0 429600.0 184500.0 430800.0 ;
      RECT  178650.0 420000.0 179550.0 436800.0 ;
      RECT  181650.0 420000.0 182550.0 436800.0 ;
      RECT  188700.0 422400.0 189900.0 423600.0 ;
      RECT  191100.0 422400.0 192750.0 423600.0 ;
      RECT  188700.0 429600.0 189900.0 430800.0 ;
      RECT  191850.0 429600.0 194700.0 430800.0 ;
      RECT  188700.0 422400.0 189900.0 423600.0 ;
      RECT  191100.0 422400.0 192300.0 423600.0 ;
      RECT  188700.0 429600.0 189900.0 430800.0 ;
      RECT  193500.0 429600.0 194700.0 430800.0 ;
      RECT  188850.0 420000.0 189750.0 436800.0 ;
      RECT  191850.0 420000.0 192750.0 436800.0 ;
      RECT  178650.0 420000.0 179550.0 436800.0 ;
      RECT  181650.0 420000.0 182550.0 436800.0 ;
      RECT  188850.0 420000.0 189750.0 436800.0 ;
      RECT  191850.0 420000.0 192750.0 436800.0 ;
      RECT  175500.0 150300.0 185700.0 199200.0 ;
      RECT  185700.0 150300.0 195900.0 199200.0 ;
      RECT  178500.0 150300.0 179700.0 163500.0 ;
      RECT  181500.0 150300.0 182700.0 163500.0 ;
      RECT  188700.0 150300.0 189900.0 163500.0 ;
      RECT  191700.0 150300.0 192900.0 163500.0 ;
      RECT  175500.0 90000.0 185700.0 150300.0 ;
      RECT  185700.0 90000.0 195900.0 150300.0 ;
      RECT  180000.0 90000.0 181200.0 92700.0 ;
      RECT  190200.0 90000.0 191400.0 92700.0 ;
      RECT  178500.0 148200.0 179700.0 150300.0 ;
      RECT  181500.0 142800.0 182700.0 150300.0 ;
      RECT  188700.0 148200.0 189900.0 150300.0 ;
      RECT  191700.0 142800.0 192900.0 150300.0 ;
      RECT  175500.0 30000.0 185700.0 90000.0 ;
      RECT  195900.0 30000.0 185700.0 90000.0 ;
      RECT  180000.0 87600.0 182700.0 88800.0 ;
      RECT  177300.0 85500.0 178500.0 90000.0 ;
      RECT  188700.0 87600.0 191400.0 88800.0 ;
      RECT  192900.0 85500.0 194100.0 90000.0 ;
      RECT  185100.0 30000.0 186300.0 90000.0 ;
      RECT  175500.0 30000.0 185700.0 8100.0 ;
      RECT  185700.0 30000.0 195900.0 8100.0 ;
      RECT  180000.0 15000.0 181200.0 8100.0 ;
      RECT  190200.0 15000.0 191400.0 8100.0 ;
      RECT  180000.0 30000.0 181200.0 28500.0 ;
      RECT  190200.0 30000.0 191400.0 28500.0 ;
      RECT  59100.0 88800.0 60000.0 420000.0 ;
      RECT  61200.0 88800.0 62100.0 420000.0 ;
      RECT  63300.0 88800.0 64200.0 420000.0 ;
      RECT  65400.0 88800.0 66300.0 420000.0 ;
      RECT  67500.0 88800.0 68400.0 420000.0 ;
      RECT  69600.0 88800.0 70500.0 420000.0 ;
      RECT  71700.0 88800.0 72600.0 420000.0 ;
      RECT  73800.0 88800.0 74700.0 420000.0 ;
      RECT  105900.0 88800.0 105000.0 142200.0 ;
      RECT  102900.0 88800.0 102000.0 142200.0 ;
      RECT  111900.0 88800.0 111000.0 142200.0 ;
      RECT  108900.0 88800.0 108000.0 142200.0 ;
      RECT  95550.0 96150.0 94650.0 97050.0 ;
      RECT  93150.0 96150.0 92250.0 97050.0 ;
      RECT  95550.0 96600.0 94650.0 99450.0 ;
      RECT  95100.0 96150.0 92700.0 97050.0 ;
      RECT  93150.0 91950.0 92250.0 96600.0 ;
      RECT  95700.0 99450.0 94500.0 100650.0 ;
      RECT  93300.0 90750.0 92100.0 91950.0 ;
      RECT  92100.0 96000.0 93300.0 97200.0 ;
      RECT  95550.0 109050.0 94650.0 108150.0 ;
      RECT  93150.0 109050.0 92250.0 108150.0 ;
      RECT  95550.0 108600.0 94650.0 105750.0 ;
      RECT  95100.0 109050.0 92700.0 108150.0 ;
      RECT  93150.0 113250.0 92250.0 108600.0 ;
      RECT  95700.0 105750.0 94500.0 104550.0 ;
      RECT  93300.0 114450.0 92100.0 113250.0 ;
      RECT  92100.0 109200.0 93300.0 108000.0 ;
      RECT  95550.0 123750.0 94650.0 124650.0 ;
      RECT  93150.0 123750.0 92250.0 124650.0 ;
      RECT  95550.0 124200.0 94650.0 127050.0 ;
      RECT  95100.0 123750.0 92700.0 124650.0 ;
      RECT  93150.0 119550.0 92250.0 124200.0 ;
      RECT  95700.0 127050.0 94500.0 128250.0 ;
      RECT  93300.0 118350.0 92100.0 119550.0 ;
      RECT  92100.0 123600.0 93300.0 124800.0 ;
      RECT  95550.0 136650.0 94650.0 135750.0 ;
      RECT  93150.0 136650.0 92250.0 135750.0 ;
      RECT  95550.0 136200.0 94650.0 133350.0 ;
      RECT  95100.0 136650.0 92700.0 135750.0 ;
      RECT  93150.0 140850.0 92250.0 136200.0 ;
      RECT  95700.0 133350.0 94500.0 132150.0 ;
      RECT  93300.0 142050.0 92100.0 140850.0 ;
      RECT  92100.0 136800.0 93300.0 135600.0 ;
      RECT  110850.0 99300.0 112050.0 100500.0 ;
      RECT  129450.0 94800.0 130650.0 96000.0 ;
      RECT  107850.0 113100.0 109050.0 114300.0 ;
      RECT  126450.0 109200.0 127650.0 110400.0 ;
      RECT  129450.0 117900.0 130650.0 119100.0 ;
      RECT  104850.0 117900.0 106050.0 119100.0 ;
      RECT  126450.0 131700.0 127650.0 132900.0 ;
      RECT  101850.0 131700.0 103050.0 132900.0 ;
      RECT  110850.0 93300.0 112050.0 94500.0 ;
      RECT  107850.0 96000.0 109050.0 97200.0 ;
      RECT  104850.0 110700.0 106050.0 111900.0 ;
      RECT  107850.0 108000.0 109050.0 109200.0 ;
      RECT  110850.0 120900.0 112050.0 122100.0 ;
      RECT  101850.0 123600.0 103050.0 124800.0 ;
      RECT  104850.0 138300.0 106050.0 139500.0 ;
      RECT  101850.0 135600.0 103050.0 136800.0 ;
      RECT  130500.0 88800.0 129600.0 142200.0 ;
      RECT  127500.0 88800.0 126600.0 142200.0 ;
      RECT  105900.0 144000.0 105000.0 197400.0 ;
      RECT  102900.0 144000.0 102000.0 197400.0 ;
      RECT  111900.0 144000.0 111000.0 197400.0 ;
      RECT  108900.0 144000.0 108000.0 197400.0 ;
      RECT  95550.0 151350.0 94650.0 152250.0 ;
      RECT  93150.0 151350.0 92250.0 152250.0 ;
      RECT  95550.0 151800.0 94650.0 154650.0 ;
      RECT  95100.0 151350.0 92700.0 152250.0 ;
      RECT  93150.0 147150.0 92250.0 151800.0 ;
      RECT  95700.0 154650.0 94500.0 155850.0 ;
      RECT  93300.0 145950.0 92100.0 147150.0 ;
      RECT  92100.0 151200.0 93300.0 152400.0 ;
      RECT  95550.0 164250.0 94650.0 163350.0 ;
      RECT  93150.0 164250.0 92250.0 163350.0 ;
      RECT  95550.0 163800.0 94650.0 160950.0 ;
      RECT  95100.0 164250.0 92700.0 163350.0 ;
      RECT  93150.0 168450.0 92250.0 163800.0 ;
      RECT  95700.0 160950.0 94500.0 159750.0 ;
      RECT  93300.0 169650.0 92100.0 168450.0 ;
      RECT  92100.0 164400.0 93300.0 163200.0 ;
      RECT  95550.0 178950.0 94650.0 179850.0 ;
      RECT  93150.0 178950.0 92250.0 179850.0 ;
      RECT  95550.0 179400.0 94650.0 182250.0 ;
      RECT  95100.0 178950.0 92700.0 179850.0 ;
      RECT  93150.0 174750.0 92250.0 179400.0 ;
      RECT  95700.0 182250.0 94500.0 183450.0 ;
      RECT  93300.0 173550.0 92100.0 174750.0 ;
      RECT  92100.0 178800.0 93300.0 180000.0 ;
      RECT  95550.0 191850.0 94650.0 190950.0 ;
      RECT  93150.0 191850.0 92250.0 190950.0 ;
      RECT  95550.0 191400.0 94650.0 188550.0 ;
      RECT  95100.0 191850.0 92700.0 190950.0 ;
      RECT  93150.0 196050.0 92250.0 191400.0 ;
      RECT  95700.0 188550.0 94500.0 187350.0 ;
      RECT  93300.0 197250.0 92100.0 196050.0 ;
      RECT  92100.0 192000.0 93300.0 190800.0 ;
      RECT  110850.0 154500.0 112050.0 155700.0 ;
      RECT  129450.0 150000.0 130650.0 151200.0 ;
      RECT  107850.0 168300.0 109050.0 169500.0 ;
      RECT  126450.0 164400.0 127650.0 165600.0 ;
      RECT  129450.0 173100.0 130650.0 174300.0 ;
      RECT  104850.0 173100.0 106050.0 174300.0 ;
      RECT  126450.0 186900.0 127650.0 188100.0 ;
      RECT  101850.0 186900.0 103050.0 188100.0 ;
      RECT  110850.0 148500.0 112050.0 149700.0 ;
      RECT  107850.0 151200.0 109050.0 152400.0 ;
      RECT  104850.0 165900.0 106050.0 167100.0 ;
      RECT  107850.0 163200.0 109050.0 164400.0 ;
      RECT  110850.0 176100.0 112050.0 177300.0 ;
      RECT  101850.0 178800.0 103050.0 180000.0 ;
      RECT  104850.0 193500.0 106050.0 194700.0 ;
      RECT  101850.0 190800.0 103050.0 192000.0 ;
      RECT  130500.0 144000.0 129600.0 197400.0 ;
      RECT  127500.0 144000.0 126600.0 197400.0 ;
      RECT  80250.0 206550.0 81150.0 207450.0 ;
      RECT  82650.0 206550.0 83550.0 207450.0 ;
      RECT  80250.0 207000.0 81150.0 209850.0 ;
      RECT  80700.0 206550.0 83100.0 207450.0 ;
      RECT  82650.0 202350.0 83550.0 207000.0 ;
      RECT  80100.0 209850.0 81300.0 211050.0 ;
      RECT  82500.0 201150.0 83700.0 202350.0 ;
      RECT  83700.0 206400.0 82500.0 207600.0 ;
      RECT  80250.0 219450.0 81150.0 218550.0 ;
      RECT  82650.0 219450.0 83550.0 218550.0 ;
      RECT  80250.0 219000.0 81150.0 216150.0 ;
      RECT  80700.0 219450.0 83100.0 218550.0 ;
      RECT  82650.0 223650.0 83550.0 219000.0 ;
      RECT  80100.0 216150.0 81300.0 214950.0 ;
      RECT  82500.0 224850.0 83700.0 223650.0 ;
      RECT  83700.0 219600.0 82500.0 218400.0 ;
      RECT  80250.0 234150.0 81150.0 235050.0 ;
      RECT  82650.0 234150.0 83550.0 235050.0 ;
      RECT  80250.0 234600.0 81150.0 237450.0 ;
      RECT  80700.0 234150.0 83100.0 235050.0 ;
      RECT  82650.0 229950.0 83550.0 234600.0 ;
      RECT  80100.0 237450.0 81300.0 238650.0 ;
      RECT  82500.0 228750.0 83700.0 229950.0 ;
      RECT  83700.0 234000.0 82500.0 235200.0 ;
      RECT  80250.0 247050.0 81150.0 246150.0 ;
      RECT  82650.0 247050.0 83550.0 246150.0 ;
      RECT  80250.0 246600.0 81150.0 243750.0 ;
      RECT  80700.0 247050.0 83100.0 246150.0 ;
      RECT  82650.0 251250.0 83550.0 246600.0 ;
      RECT  80100.0 243750.0 81300.0 242550.0 ;
      RECT  82500.0 252450.0 83700.0 251250.0 ;
      RECT  83700.0 247200.0 82500.0 246000.0 ;
      RECT  80250.0 261750.0 81150.0 262650.0 ;
      RECT  82650.0 261750.0 83550.0 262650.0 ;
      RECT  80250.0 262200.0 81150.0 265050.0 ;
      RECT  80700.0 261750.0 83100.0 262650.0 ;
      RECT  82650.0 257550.0 83550.0 262200.0 ;
      RECT  80100.0 265050.0 81300.0 266250.0 ;
      RECT  82500.0 256350.0 83700.0 257550.0 ;
      RECT  83700.0 261600.0 82500.0 262800.0 ;
      RECT  80250.0 274650.0 81150.0 273750.0 ;
      RECT  82650.0 274650.0 83550.0 273750.0 ;
      RECT  80250.0 274200.0 81150.0 271350.0 ;
      RECT  80700.0 274650.0 83100.0 273750.0 ;
      RECT  82650.0 278850.0 83550.0 274200.0 ;
      RECT  80100.0 271350.0 81300.0 270150.0 ;
      RECT  82500.0 280050.0 83700.0 278850.0 ;
      RECT  83700.0 274800.0 82500.0 273600.0 ;
      RECT  80250.0 289350.0 81150.0 290250.0 ;
      RECT  82650.0 289350.0 83550.0 290250.0 ;
      RECT  80250.0 289800.0 81150.0 292650.0 ;
      RECT  80700.0 289350.0 83100.0 290250.0 ;
      RECT  82650.0 285150.0 83550.0 289800.0 ;
      RECT  80100.0 292650.0 81300.0 293850.0 ;
      RECT  82500.0 283950.0 83700.0 285150.0 ;
      RECT  83700.0 289200.0 82500.0 290400.0 ;
      RECT  80250.0 302250.0 81150.0 301350.0 ;
      RECT  82650.0 302250.0 83550.0 301350.0 ;
      RECT  80250.0 301800.0 81150.0 298950.0 ;
      RECT  80700.0 302250.0 83100.0 301350.0 ;
      RECT  82650.0 306450.0 83550.0 301800.0 ;
      RECT  80100.0 298950.0 81300.0 297750.0 ;
      RECT  82500.0 307650.0 83700.0 306450.0 ;
      RECT  83700.0 302400.0 82500.0 301200.0 ;
      RECT  80250.0 316950.0 81150.0 317850.0 ;
      RECT  82650.0 316950.0 83550.0 317850.0 ;
      RECT  80250.0 317400.0 81150.0 320250.0 ;
      RECT  80700.0 316950.0 83100.0 317850.0 ;
      RECT  82650.0 312750.0 83550.0 317400.0 ;
      RECT  80100.0 320250.0 81300.0 321450.0 ;
      RECT  82500.0 311550.0 83700.0 312750.0 ;
      RECT  83700.0 316800.0 82500.0 318000.0 ;
      RECT  80250.0 329850.0 81150.0 328950.0 ;
      RECT  82650.0 329850.0 83550.0 328950.0 ;
      RECT  80250.0 329400.0 81150.0 326550.0 ;
      RECT  80700.0 329850.0 83100.0 328950.0 ;
      RECT  82650.0 334050.0 83550.0 329400.0 ;
      RECT  80100.0 326550.0 81300.0 325350.0 ;
      RECT  82500.0 335250.0 83700.0 334050.0 ;
      RECT  83700.0 330000.0 82500.0 328800.0 ;
      RECT  80250.0 344550.0 81150.0 345450.0 ;
      RECT  82650.0 344550.0 83550.0 345450.0 ;
      RECT  80250.0 345000.0 81150.0 347850.0 ;
      RECT  80700.0 344550.0 83100.0 345450.0 ;
      RECT  82650.0 340350.0 83550.0 345000.0 ;
      RECT  80100.0 347850.0 81300.0 349050.0 ;
      RECT  82500.0 339150.0 83700.0 340350.0 ;
      RECT  83700.0 344400.0 82500.0 345600.0 ;
      RECT  80250.0 357450.0 81150.0 356550.0 ;
      RECT  82650.0 357450.0 83550.0 356550.0 ;
      RECT  80250.0 357000.0 81150.0 354150.0 ;
      RECT  80700.0 357450.0 83100.0 356550.0 ;
      RECT  82650.0 361650.0 83550.0 357000.0 ;
      RECT  80100.0 354150.0 81300.0 352950.0 ;
      RECT  82500.0 362850.0 83700.0 361650.0 ;
      RECT  83700.0 357600.0 82500.0 356400.0 ;
      RECT  80250.0 372150.0 81150.0 373050.0 ;
      RECT  82650.0 372150.0 83550.0 373050.0 ;
      RECT  80250.0 372600.0 81150.0 375450.0 ;
      RECT  80700.0 372150.0 83100.0 373050.0 ;
      RECT  82650.0 367950.0 83550.0 372600.0 ;
      RECT  80100.0 375450.0 81300.0 376650.0 ;
      RECT  82500.0 366750.0 83700.0 367950.0 ;
      RECT  83700.0 372000.0 82500.0 373200.0 ;
      RECT  80250.0 385050.0 81150.0 384150.0 ;
      RECT  82650.0 385050.0 83550.0 384150.0 ;
      RECT  80250.0 384600.0 81150.0 381750.0 ;
      RECT  80700.0 385050.0 83100.0 384150.0 ;
      RECT  82650.0 389250.0 83550.0 384600.0 ;
      RECT  80100.0 381750.0 81300.0 380550.0 ;
      RECT  82500.0 390450.0 83700.0 389250.0 ;
      RECT  83700.0 385200.0 82500.0 384000.0 ;
      RECT  80250.0 399750.0 81150.0 400650.0 ;
      RECT  82650.0 399750.0 83550.0 400650.0 ;
      RECT  80250.0 400200.0 81150.0 403050.0 ;
      RECT  80700.0 399750.0 83100.0 400650.0 ;
      RECT  82650.0 395550.0 83550.0 400200.0 ;
      RECT  80100.0 403050.0 81300.0 404250.0 ;
      RECT  82500.0 394350.0 83700.0 395550.0 ;
      RECT  83700.0 399600.0 82500.0 400800.0 ;
      RECT  80250.0 412650.0 81150.0 411750.0 ;
      RECT  82650.0 412650.0 83550.0 411750.0 ;
      RECT  80250.0 412200.0 81150.0 409350.0 ;
      RECT  80700.0 412650.0 83100.0 411750.0 ;
      RECT  82650.0 416850.0 83550.0 412200.0 ;
      RECT  80100.0 409350.0 81300.0 408150.0 ;
      RECT  82500.0 418050.0 83700.0 416850.0 ;
      RECT  83700.0 412800.0 82500.0 411600.0 ;
      RECT  60150.0 94800.0 58950.0 96000.0 ;
      RECT  62250.0 109200.0 61050.0 110400.0 ;
      RECT  64350.0 122400.0 63150.0 123600.0 ;
      RECT  66450.0 136800.0 65250.0 138000.0 ;
      RECT  68550.0 150000.0 67350.0 151200.0 ;
      RECT  70650.0 164400.0 69450.0 165600.0 ;
      RECT  72750.0 177600.0 71550.0 178800.0 ;
      RECT  74850.0 192000.0 73650.0 193200.0 ;
      RECT  60150.0 206400.0 58950.0 207600.0 ;
      RECT  68550.0 203700.0 67350.0 204900.0 ;
      RECT  60150.0 218400.0 58950.0 219600.0 ;
      RECT  70650.0 221100.0 69450.0 222300.0 ;
      RECT  60150.0 234000.0 58950.0 235200.0 ;
      RECT  72750.0 231300.0 71550.0 232500.0 ;
      RECT  60150.0 246000.0 58950.0 247200.0 ;
      RECT  74850.0 248700.0 73650.0 249900.0 ;
      RECT  62250.0 261600.0 61050.0 262800.0 ;
      RECT  68550.0 258900.0 67350.0 260100.0 ;
      RECT  62250.0 273600.0 61050.0 274800.0 ;
      RECT  70650.0 276300.0 69450.0 277500.0 ;
      RECT  62250.0 289200.0 61050.0 290400.0 ;
      RECT  72750.0 286500.0 71550.0 287700.0 ;
      RECT  62250.0 301200.0 61050.0 302400.0 ;
      RECT  74850.0 303900.0 73650.0 305100.0 ;
      RECT  64350.0 316800.0 63150.0 318000.0 ;
      RECT  68550.0 314100.0 67350.0 315300.0 ;
      RECT  64350.0 328800.0 63150.0 330000.0 ;
      RECT  70650.0 331500.0 69450.0 332700.0 ;
      RECT  64350.0 344400.0 63150.0 345600.0 ;
      RECT  72750.0 341700.0 71550.0 342900.0 ;
      RECT  64350.0 356400.0 63150.0 357600.0 ;
      RECT  74850.0 359100.0 73650.0 360300.0 ;
      RECT  66450.0 372000.0 65250.0 373200.0 ;
      RECT  68550.0 369300.0 67350.0 370500.0 ;
      RECT  66450.0 384000.0 65250.0 385200.0 ;
      RECT  70650.0 386700.0 69450.0 387900.0 ;
      RECT  66450.0 399600.0 65250.0 400800.0 ;
      RECT  72750.0 396900.0 71550.0 398100.0 ;
      RECT  66450.0 411600.0 65250.0 412800.0 ;
      RECT  74850.0 414300.0 73650.0 415500.0 ;
      RECT  129600.0 88800.0 130500.0 142200.0 ;
      RECT  126600.0 88800.0 127500.0 142200.0 ;
      RECT  129600.0 144000.0 130500.0 197400.0 ;
      RECT  126600.0 144000.0 127500.0 197400.0 ;
      RECT  104550.0 203850.0 105450.0 204750.0 ;
      RECT  104550.0 203400.0 105450.0 204300.0 ;
      RECT  105000.0 203850.0 121200.0 204750.0 ;
      RECT  104550.0 221250.0 105450.0 222150.0 ;
      RECT  104550.0 221700.0 105450.0 222600.0 ;
      RECT  105000.0 221250.0 121200.0 222150.0 ;
      RECT  104550.0 231450.0 105450.0 232350.0 ;
      RECT  104550.0 231000.0 105450.0 231900.0 ;
      RECT  105000.0 231450.0 121200.0 232350.0 ;
      RECT  104550.0 248850.0 105450.0 249750.0 ;
      RECT  104550.0 249300.0 105450.0 250200.0 ;
      RECT  105000.0 248850.0 121200.0 249750.0 ;
      RECT  104550.0 259050.0 105450.0 259950.0 ;
      RECT  104550.0 258600.0 105450.0 259500.0 ;
      RECT  105000.0 259050.0 121200.0 259950.0 ;
      RECT  104550.0 276450.0 105450.0 277350.0 ;
      RECT  104550.0 276900.0 105450.0 277800.0 ;
      RECT  105000.0 276450.0 121200.0 277350.0 ;
      RECT  104550.0 286650.0 105450.0 287550.0 ;
      RECT  104550.0 286200.0 105450.0 287100.0 ;
      RECT  105000.0 286650.0 121200.0 287550.0 ;
      RECT  104550.0 304050.0 105450.0 304950.0 ;
      RECT  104550.0 304500.0 105450.0 305400.0 ;
      RECT  105000.0 304050.0 121200.0 304950.0 ;
      RECT  104550.0 314250.0 105450.0 315150.0 ;
      RECT  104550.0 313800.0 105450.0 314700.0 ;
      RECT  105000.0 314250.0 121200.0 315150.0 ;
      RECT  104550.0 331650.0 105450.0 332550.0 ;
      RECT  104550.0 332100.0 105450.0 333000.0 ;
      RECT  105000.0 331650.0 121200.0 332550.0 ;
      RECT  104550.0 341850.0 105450.0 342750.0 ;
      RECT  104550.0 341400.0 105450.0 342300.0 ;
      RECT  105000.0 341850.0 121200.0 342750.0 ;
      RECT  104550.0 359250.0 105450.0 360150.0 ;
      RECT  104550.0 359700.0 105450.0 360600.0 ;
      RECT  105000.0 359250.0 121200.0 360150.0 ;
      RECT  104550.0 369450.0 105450.0 370350.0 ;
      RECT  104550.0 369000.0 105450.0 369900.0 ;
      RECT  105000.0 369450.0 121200.0 370350.0 ;
      RECT  104550.0 386850.0 105450.0 387750.0 ;
      RECT  104550.0 387300.0 105450.0 388200.0 ;
      RECT  105000.0 386850.0 121200.0 387750.0 ;
      RECT  104550.0 397050.0 105450.0 397950.0 ;
      RECT  104550.0 396600.0 105450.0 397500.0 ;
      RECT  105000.0 397050.0 121200.0 397950.0 ;
      RECT  104550.0 414450.0 105450.0 415350.0 ;
      RECT  104550.0 414900.0 105450.0 415800.0 ;
      RECT  105000.0 414450.0 121200.0 415350.0 ;
      RECT  120150.0 206550.0 121050.0 207450.0 ;
      RECT  122550.0 206550.0 123450.0 207450.0 ;
      RECT  120150.0 207000.0 121050.0 209850.0 ;
      RECT  120600.0 206550.0 123000.0 207450.0 ;
      RECT  122550.0 202350.0 123450.0 207000.0 ;
      RECT  120000.0 209850.0 121200.0 211050.0 ;
      RECT  122400.0 201150.0 123600.0 202350.0 ;
      RECT  123600.0 206400.0 122400.0 207600.0 ;
      RECT  102450.0 205200.0 103650.0 206400.0 ;
      RECT  104400.0 202800.0 105600.0 204000.0 ;
      RECT  121200.0 203700.0 120000.0 204900.0 ;
      RECT  120150.0 219450.0 121050.0 218550.0 ;
      RECT  122550.0 219450.0 123450.0 218550.0 ;
      RECT  120150.0 219000.0 121050.0 216150.0 ;
      RECT  120600.0 219450.0 123000.0 218550.0 ;
      RECT  122550.0 223650.0 123450.0 219000.0 ;
      RECT  120000.0 216150.0 121200.0 214950.0 ;
      RECT  122400.0 224850.0 123600.0 223650.0 ;
      RECT  123600.0 219600.0 122400.0 218400.0 ;
      RECT  102450.0 219600.0 103650.0 220800.0 ;
      RECT  104400.0 222000.0 105600.0 223200.0 ;
      RECT  121200.0 221100.0 120000.0 222300.0 ;
      RECT  120150.0 234150.0 121050.0 235050.0 ;
      RECT  122550.0 234150.0 123450.0 235050.0 ;
      RECT  120150.0 234600.0 121050.0 237450.0 ;
      RECT  120600.0 234150.0 123000.0 235050.0 ;
      RECT  122550.0 229950.0 123450.0 234600.0 ;
      RECT  120000.0 237450.0 121200.0 238650.0 ;
      RECT  122400.0 228750.0 123600.0 229950.0 ;
      RECT  123600.0 234000.0 122400.0 235200.0 ;
      RECT  102450.0 232800.0 103650.0 234000.0 ;
      RECT  104400.0 230400.0 105600.0 231600.0 ;
      RECT  121200.0 231300.0 120000.0 232500.0 ;
      RECT  120150.0 247050.0 121050.0 246150.0 ;
      RECT  122550.0 247050.0 123450.0 246150.0 ;
      RECT  120150.0 246600.0 121050.0 243750.0 ;
      RECT  120600.0 247050.0 123000.0 246150.0 ;
      RECT  122550.0 251250.0 123450.0 246600.0 ;
      RECT  120000.0 243750.0 121200.0 242550.0 ;
      RECT  122400.0 252450.0 123600.0 251250.0 ;
      RECT  123600.0 247200.0 122400.0 246000.0 ;
      RECT  102450.0 247200.0 103650.0 248400.0 ;
      RECT  104400.0 249600.0 105600.0 250800.0 ;
      RECT  121200.0 248700.0 120000.0 249900.0 ;
      RECT  120150.0 261750.0 121050.0 262650.0 ;
      RECT  122550.0 261750.0 123450.0 262650.0 ;
      RECT  120150.0 262200.0 121050.0 265050.0 ;
      RECT  120600.0 261750.0 123000.0 262650.0 ;
      RECT  122550.0 257550.0 123450.0 262200.0 ;
      RECT  120000.0 265050.0 121200.0 266250.0 ;
      RECT  122400.0 256350.0 123600.0 257550.0 ;
      RECT  123600.0 261600.0 122400.0 262800.0 ;
      RECT  102450.0 260400.0 103650.0 261600.0 ;
      RECT  104400.0 258000.0 105600.0 259200.0 ;
      RECT  121200.0 258900.0 120000.0 260100.0 ;
      RECT  120150.0 274650.0 121050.0 273750.0 ;
      RECT  122550.0 274650.0 123450.0 273750.0 ;
      RECT  120150.0 274200.0 121050.0 271350.0 ;
      RECT  120600.0 274650.0 123000.0 273750.0 ;
      RECT  122550.0 278850.0 123450.0 274200.0 ;
      RECT  120000.0 271350.0 121200.0 270150.0 ;
      RECT  122400.0 280050.0 123600.0 278850.0 ;
      RECT  123600.0 274800.0 122400.0 273600.0 ;
      RECT  102450.0 274800.0 103650.0 276000.0 ;
      RECT  104400.0 277200.0 105600.0 278400.0 ;
      RECT  121200.0 276300.0 120000.0 277500.0 ;
      RECT  120150.0 289350.0 121050.0 290250.0 ;
      RECT  122550.0 289350.0 123450.0 290250.0 ;
      RECT  120150.0 289800.0 121050.0 292650.0 ;
      RECT  120600.0 289350.0 123000.0 290250.0 ;
      RECT  122550.0 285150.0 123450.0 289800.0 ;
      RECT  120000.0 292650.0 121200.0 293850.0 ;
      RECT  122400.0 283950.0 123600.0 285150.0 ;
      RECT  123600.0 289200.0 122400.0 290400.0 ;
      RECT  102450.0 288000.0 103650.0 289200.0 ;
      RECT  104400.0 285600.0 105600.0 286800.0 ;
      RECT  121200.0 286500.0 120000.0 287700.0 ;
      RECT  120150.0 302250.0 121050.0 301350.0 ;
      RECT  122550.0 302250.0 123450.0 301350.0 ;
      RECT  120150.0 301800.0 121050.0 298950.0 ;
      RECT  120600.0 302250.0 123000.0 301350.0 ;
      RECT  122550.0 306450.0 123450.0 301800.0 ;
      RECT  120000.0 298950.0 121200.0 297750.0 ;
      RECT  122400.0 307650.0 123600.0 306450.0 ;
      RECT  123600.0 302400.0 122400.0 301200.0 ;
      RECT  102450.0 302400.0 103650.0 303600.0 ;
      RECT  104400.0 304800.0 105600.0 306000.0 ;
      RECT  121200.0 303900.0 120000.0 305100.0 ;
      RECT  120150.0 316950.0 121050.0 317850.0 ;
      RECT  122550.0 316950.0 123450.0 317850.0 ;
      RECT  120150.0 317400.0 121050.0 320250.0 ;
      RECT  120600.0 316950.0 123000.0 317850.0 ;
      RECT  122550.0 312750.0 123450.0 317400.0 ;
      RECT  120000.0 320250.0 121200.0 321450.0 ;
      RECT  122400.0 311550.0 123600.0 312750.0 ;
      RECT  123600.0 316800.0 122400.0 318000.0 ;
      RECT  102450.0 315600.0 103650.0 316800.0 ;
      RECT  104400.0 313200.0 105600.0 314400.0 ;
      RECT  121200.0 314100.0 120000.0 315300.0 ;
      RECT  120150.0 329850.0 121050.0 328950.0 ;
      RECT  122550.0 329850.0 123450.0 328950.0 ;
      RECT  120150.0 329400.0 121050.0 326550.0 ;
      RECT  120600.0 329850.0 123000.0 328950.0 ;
      RECT  122550.0 334050.0 123450.0 329400.0 ;
      RECT  120000.0 326550.0 121200.0 325350.0 ;
      RECT  122400.0 335250.0 123600.0 334050.0 ;
      RECT  123600.0 330000.0 122400.0 328800.0 ;
      RECT  102450.0 330000.0 103650.0 331200.0 ;
      RECT  104400.0 332400.0 105600.0 333600.0 ;
      RECT  121200.0 331500.0 120000.0 332700.0 ;
      RECT  120150.0 344550.0 121050.0 345450.0 ;
      RECT  122550.0 344550.0 123450.0 345450.0 ;
      RECT  120150.0 345000.0 121050.0 347850.0 ;
      RECT  120600.0 344550.0 123000.0 345450.0 ;
      RECT  122550.0 340350.0 123450.0 345000.0 ;
      RECT  120000.0 347850.0 121200.0 349050.0 ;
      RECT  122400.0 339150.0 123600.0 340350.0 ;
      RECT  123600.0 344400.0 122400.0 345600.0 ;
      RECT  102450.0 343200.0 103650.0 344400.0 ;
      RECT  104400.0 340800.0 105600.0 342000.0 ;
      RECT  121200.0 341700.0 120000.0 342900.0 ;
      RECT  120150.0 357450.0 121050.0 356550.0 ;
      RECT  122550.0 357450.0 123450.0 356550.0 ;
      RECT  120150.0 357000.0 121050.0 354150.0 ;
      RECT  120600.0 357450.0 123000.0 356550.0 ;
      RECT  122550.0 361650.0 123450.0 357000.0 ;
      RECT  120000.0 354150.0 121200.0 352950.0 ;
      RECT  122400.0 362850.0 123600.0 361650.0 ;
      RECT  123600.0 357600.0 122400.0 356400.0 ;
      RECT  102450.0 357600.0 103650.0 358800.0 ;
      RECT  104400.0 360000.0 105600.0 361200.0 ;
      RECT  121200.0 359100.0 120000.0 360300.0 ;
      RECT  120150.0 372150.0 121050.0 373050.0 ;
      RECT  122550.0 372150.0 123450.0 373050.0 ;
      RECT  120150.0 372600.0 121050.0 375450.0 ;
      RECT  120600.0 372150.0 123000.0 373050.0 ;
      RECT  122550.0 367950.0 123450.0 372600.0 ;
      RECT  120000.0 375450.0 121200.0 376650.0 ;
      RECT  122400.0 366750.0 123600.0 367950.0 ;
      RECT  123600.0 372000.0 122400.0 373200.0 ;
      RECT  102450.0 370800.0 103650.0 372000.0 ;
      RECT  104400.0 368400.0 105600.0 369600.0 ;
      RECT  121200.0 369300.0 120000.0 370500.0 ;
      RECT  120150.0 385050.0 121050.0 384150.0 ;
      RECT  122550.0 385050.0 123450.0 384150.0 ;
      RECT  120150.0 384600.0 121050.0 381750.0 ;
      RECT  120600.0 385050.0 123000.0 384150.0 ;
      RECT  122550.0 389250.0 123450.0 384600.0 ;
      RECT  120000.0 381750.0 121200.0 380550.0 ;
      RECT  122400.0 390450.0 123600.0 389250.0 ;
      RECT  123600.0 385200.0 122400.0 384000.0 ;
      RECT  102450.0 385200.0 103650.0 386400.0 ;
      RECT  104400.0 387600.0 105600.0 388800.0 ;
      RECT  121200.0 386700.0 120000.0 387900.0 ;
      RECT  120150.0 399750.0 121050.0 400650.0 ;
      RECT  122550.0 399750.0 123450.0 400650.0 ;
      RECT  120150.0 400200.0 121050.0 403050.0 ;
      RECT  120600.0 399750.0 123000.0 400650.0 ;
      RECT  122550.0 395550.0 123450.0 400200.0 ;
      RECT  120000.0 403050.0 121200.0 404250.0 ;
      RECT  122400.0 394350.0 123600.0 395550.0 ;
      RECT  123600.0 399600.0 122400.0 400800.0 ;
      RECT  102450.0 398400.0 103650.0 399600.0 ;
      RECT  104400.0 396000.0 105600.0 397200.0 ;
      RECT  121200.0 396900.0 120000.0 398100.0 ;
      RECT  120150.0 412650.0 121050.0 411750.0 ;
      RECT  122550.0 412650.0 123450.0 411750.0 ;
      RECT  120150.0 412200.0 121050.0 409350.0 ;
      RECT  120600.0 412650.0 123000.0 411750.0 ;
      RECT  122550.0 416850.0 123450.0 412200.0 ;
      RECT  120000.0 409350.0 121200.0 408150.0 ;
      RECT  122400.0 418050.0 123600.0 416850.0 ;
      RECT  123600.0 412800.0 122400.0 411600.0 ;
      RECT  102450.0 412800.0 103650.0 414000.0 ;
      RECT  104400.0 415200.0 105600.0 416400.0 ;
      RECT  121200.0 414300.0 120000.0 415500.0 ;
      RECT  102600.0 199200.0 103500.0 420000.0 ;
      RECT  59100.0 83400.0 119100.0 73200.0 ;
      RECT  59100.0 63000.0 119100.0 73200.0 ;
      RECT  59100.0 63000.0 119100.0 52800.0 ;
      RECT  59100.0 42600.0 119100.0 52800.0 ;
      RECT  116700.0 78900.0 117900.0 76200.0 ;
      RECT  114600.0 81600.0 119100.0 80400.0 ;
      RECT  116700.0 70200.0 117900.0 67500.0 ;
      RECT  114600.0 66000.0 119100.0 64800.0 ;
      RECT  116700.0 58500.0 117900.0 55800.0 ;
      RECT  114600.0 61200.0 119100.0 60000.0 ;
      RECT  116700.0 49800.0 117900.0 47100.0 ;
      RECT  114600.0 45600.0 119100.0 44400.0 ;
      RECT  59100.0 73800.0 119100.0 72600.0 ;
      RECT  59100.0 53400.0 119100.0 52200.0 ;
      RECT  176550.0 5850.0 177750.0 7050.0 ;
      RECT  186750.0 5850.0 187950.0 7050.0 ;
      RECT  180300.0 300.0 181500.0 1500.0 ;
      RECT  190500.0 300.0 191700.0 1500.0 ;
      RECT  148050.0 199800.0 149250.0 198600.0 ;
      RECT  148050.0 227400.0 149250.0 226200.0 ;
      RECT  148050.0 255000.0 149250.0 253800.0 ;
      RECT  148050.0 282600.0 149250.0 281400.0 ;
      RECT  148050.0 310200.0 149250.0 309000.0 ;
      RECT  148050.0 337800.0 149250.0 336600.0 ;
      RECT  148050.0 365400.0 149250.0 364200.0 ;
      RECT  148050.0 393000.0 149250.0 391800.0 ;
      RECT  148050.0 420600.0 149250.0 419400.0 ;
      RECT  130500.0 91050.0 129300.0 92250.0 ;
      RECT  135600.0 90900.0 134400.0 92100.0 ;
      RECT  127500.0 104850.0 126300.0 106050.0 ;
      RECT  138300.0 104700.0 137100.0 105900.0 ;
      RECT  130500.0 146250.0 129300.0 147450.0 ;
      RECT  141000.0 146100.0 139800.0 147300.0 ;
      RECT  127500.0 160050.0 126300.0 161250.0 ;
      RECT  143700.0 159900.0 142500.0 161100.0 ;
      RECT  132600.0 88200.0 131400.0 89400.0 ;
      RECT  132600.0 88200.0 131400.0 89400.0 ;
      RECT  147450.0 89400.0 148650.0 88200.0 ;
      RECT  132600.0 115800.0 131400.0 117000.0 ;
      RECT  132600.0 115800.0 131400.0 117000.0 ;
      RECT  147450.0 117000.0 148650.0 115800.0 ;
      RECT  132600.0 143400.0 131400.0 144600.0 ;
      RECT  132600.0 143400.0 131400.0 144600.0 ;
      RECT  147450.0 144600.0 148650.0 143400.0 ;
      RECT  132600.0 171000.0 131400.0 172200.0 ;
      RECT  132600.0 171000.0 131400.0 172200.0 ;
      RECT  147450.0 172200.0 148650.0 171000.0 ;
      RECT  118500.0 76950.0 117300.0 78150.0 ;
      RECT  135600.0 76950.0 134400.0 78150.0 ;
      RECT  118500.0 68250.0 117300.0 69450.0 ;
      RECT  138300.0 68250.0 137100.0 69450.0 ;
      RECT  118500.0 56550.0 117300.0 57750.0 ;
      RECT  141000.0 56550.0 139800.0 57750.0 ;
      RECT  118500.0 47850.0 117300.0 49050.0 ;
      RECT  143700.0 47850.0 142500.0 49050.0 ;
      RECT  120300.0 72600.0 119100.0 73800.0 ;
      RECT  149250.0 72750.0 148050.0 73950.0 ;
      RECT  120300.0 52200.0 119100.0 53400.0 ;
      RECT  149250.0 52350.0 148050.0 53550.0 ;
      RECT  164400.0 32250.0 163200.0 33450.0 ;
      RECT  159000.0 27750.0 157800.0 28950.0 ;
      RECT  161700.0 25350.0 160500.0 26550.0 ;
      RECT  164400.0 424650.0 163200.0 425850.0 ;
      RECT  167100.0 96750.0 165900.0 97950.0 ;
      RECT  169800.0 194850.0 168600.0 196050.0 ;
      RECT  156300.0 84900.0 155100.0 86100.0 ;
      RECT  103650.0 421500.0 102450.0 422700.0 ;
      RECT  156300.0 421500.0 155100.0 422700.0 ;
      RECT  152550.0 23400.0 151350.0 24600.0 ;
      RECT  152550.0 192900.0 151350.0 194100.0 ;
      RECT  152550.0 94800.0 151350.0 96000.0 ;
      RECT  180000.0 0.0 180900.0 1800.0 ;
      RECT  190200.0 0.0 191100.0 1800.0 ;
      RECT  168750.0 0.0 169650.0 436800.0 ;
      RECT  166050.0 0.0 166950.0 436800.0 ;
      RECT  157950.0 0.0 158850.0 436800.0 ;
      RECT  160650.0 0.0 161550.0 436800.0 ;
      RECT  163350.0 0.0 164250.0 436800.0 ;
      RECT  155250.0 0.0 156150.0 436800.0 ;
      RECT  148050.0 0.0 152550.0 436800.0 ;
      RECT  49800.0 289800.0 1.42108547152e-11 290700.0 ;
      RECT  49800.0 292500.0 1.42108547152e-11 293400.0 ;
      RECT  49800.0 295200.0 1.42108547152e-11 296100.0 ;
      RECT  49800.0 300600.0 1.42108547152e-11 301500.0 ;
      RECT  33750.0 205050.0 32850.0 284850.0 ;
      RECT  49800.0 287100.0 47100.0 288000.0 ;
      RECT  38700.0 297900.0 36000.0 298800.0 ;
      RECT  24900.0 287100.0 22200.0 288000.0 ;
      RECT  11100.0 297900.0 8400.0 298800.0 ;
      RECT  7.1054273576e-12 202200.0 10200.0 262200.0 ;
      RECT  20400.0 202200.0 10200.0 262200.0 ;
      RECT  20400.0 202200.0 30600.0 262200.0 ;
      RECT  4500.0 259800.0 7200.0 261000.0 ;
      RECT  1800.0 257700.0 3000.0 262200.0 ;
      RECT  13200.0 259800.0 15900.0 261000.0 ;
      RECT  17400.0 257700.0 18600.0 262200.0 ;
      RECT  24900.0 259800.0 27600.0 261000.0 ;
      RECT  22200.0 257700.0 23400.0 262200.0 ;
      RECT  9600.0 202200.0 10800.0 262200.0 ;
      RECT  30000.0 202200.0 31200.0 262200.0 ;
      RECT  46650.0 317850.0 39150.0 318750.0 ;
      RECT  41700.0 313050.0 40800.0 313950.0 ;
      RECT  41700.0 317850.0 40800.0 318750.0 ;
      RECT  41250.0 313050.0 39150.0 313950.0 ;
      RECT  41700.0 313500.0 40800.0 318300.0 ;
      RECT  46650.0 317850.0 41250.0 318750.0 ;
      RECT  39150.0 312900.0 37950.0 314100.0 ;
      RECT  39150.0 317700.0 37950.0 318900.0 ;
      RECT  47850.0 317700.0 46650.0 318900.0 ;
      RECT  41850.0 317700.0 40650.0 318900.0 ;
      RECT  28800.0 315450.0 29700.0 316350.0 ;
      RECT  29250.0 315450.0 32250.0 316350.0 ;
      RECT  28800.0 315900.0 29700.0 316800.0 ;
      RECT  23700.0 315450.0 24600.0 316350.0 ;
      RECT  23700.0 314100.0 24600.0 315900.0 ;
      RECT  24150.0 315450.0 29250.0 316350.0 ;
      RECT  32250.0 315300.0 33450.0 316500.0 ;
      RECT  23550.0 314100.0 24750.0 312900.0 ;
      RECT  28650.0 317400.0 29850.0 316200.0 ;
      RECT  29550.0 330150.0 30450.0 331050.0 ;
      RECT  29550.0 332550.0 30450.0 333450.0 ;
      RECT  30000.0 330150.0 32850.0 331050.0 ;
      RECT  29550.0 330600.0 30450.0 333000.0 ;
      RECT  25350.0 332550.0 30000.0 333450.0 ;
      RECT  32850.0 330000.0 34050.0 331200.0 ;
      RECT  24150.0 332400.0 25350.0 333600.0 ;
      RECT  29400.0 333600.0 30600.0 332400.0 ;
      RECT  19050.0 327450.0 11550.0 328350.0 ;
      RECT  14100.0 322650.0 13200.0 323550.0 ;
      RECT  14100.0 327450.0 13200.0 328350.0 ;
      RECT  13650.0 322650.0 11550.0 323550.0 ;
      RECT  14100.0 323100.0 13200.0 327900.0 ;
      RECT  19050.0 327450.0 13650.0 328350.0 ;
      RECT  11550.0 322500.0 10350.0 323700.0 ;
      RECT  11550.0 327300.0 10350.0 328500.0 ;
      RECT  20250.0 327300.0 19050.0 328500.0 ;
      RECT  14250.0 327300.0 13050.0 328500.0 ;
      RECT  3000.0 262800.0 1800.0 261600.0 ;
      RECT  3000.0 301650.0 1800.0 300450.0 ;
      RECT  6450.0 261600.0 5250.0 260400.0 ;
      RECT  6450.0 290850.0 5250.0 289650.0 ;
      RECT  18600.0 262800.0 17400.0 261600.0 ;
      RECT  18600.0 293550.0 17400.0 292350.0 ;
      RECT  23400.0 262800.0 22200.0 261600.0 ;
      RECT  23400.0 296250.0 22200.0 295050.0 ;
      RECT  10800.0 262800.0 9600.0 261600.0 ;
      RECT  10800.0 288150.0 9600.0 286950.0 ;
      RECT  31200.0 262800.0 30000.0 261600.0 ;
      RECT  31200.0 288150.0 30000.0 286950.0 ;
      RECT  22650.0 371700.0 21750.0 425400.0 ;
      RECT  22650.0 381300.0 21750.0 384000.0 ;
      RECT  22650.0 384000.0 21750.0 426000.0 ;
      RECT  17250.0 423300.0 16350.0 426000.0 ;
      RECT  20400.0 375900.0 19500.0 384000.0 ;
      RECT  13650.0 375900.0 12750.0 380700.0 ;
      RECT  42750.0 415500.0 43650.0 422700.0 ;
      RECT  35550.0 424650.0 36450.0 425550.0 ;
      RECT  35550.0 425850.0 36450.0 426750.0 ;
      RECT  36000.0 424650.0 43200.0 425550.0 ;
      RECT  35550.0 425100.0 36450.0 426300.0 ;
      RECT  28800.0 425850.0 36000.0 426750.0 ;
      RECT  28350.0 416700.0 29250.0 423900.0 ;
      RECT  42600.0 422100.0 43800.0 423300.0 ;
      RECT  28200.0 425700.0 29400.0 426900.0 ;
      RECT  28200.0 416100.0 29400.0 417300.0 ;
      RECT  42600.0 414900.0 43800.0 416100.0 ;
      RECT  42600.0 424500.0 43800.0 425700.0 ;
      RECT  28200.0 423300.0 29400.0 424500.0 ;
      RECT  16800.0 395100.0 6600.0 381300.0 ;
      RECT  16800.0 395100.0 6600.0 408900.0 ;
      RECT  16800.0 422700.0 6600.0 408900.0 ;
      RECT  13800.0 395700.0 12600.0 424500.0 ;
      RECT  10800.0 394500.0 9600.0 423300.0 ;
      RECT  17400.0 394500.0 16200.0 423300.0 ;
      RECT  7200.0 394500.0 6000.0 423300.0 ;
      RECT  22650.0 396600.0 21450.0 397800.0 ;
      RECT  22650.0 420000.0 21450.0 421200.0 ;
      RECT  22650.0 410100.0 21450.0 411300.0 ;
      RECT  22650.0 370500.0 21450.0 371700.0 ;
      RECT  21600.0 425400.0 22800.0 426600.0 ;
      RECT  16200.0 425400.0 17400.0 426600.0 ;
      RECT  19350.0 383400.0 20550.0 384600.0 ;
      RECT  19350.0 375300.0 20550.0 376500.0 ;
      RECT  12600.0 375300.0 13800.0 376500.0 ;
      RECT  43950.0 285450.0 42750.0 284250.0 ;
      RECT  43950.0 244500.0 42750.0 243300.0 ;
      RECT  43950.0 304350.0 42750.0 303150.0 ;
      RECT  43950.0 244500.0 42750.0 243300.0 ;
      RECT  33900.0 205650.0 32700.0 204450.0 ;
      RECT  29850.0 285450.0 28650.0 284250.0 ;
      RECT  27150.0 290850.0 25950.0 289650.0 ;
      RECT  30600.0 328200.0 29400.0 327000.0 ;
      RECT  30600.0 328200.0 29400.0 327000.0 ;
      RECT  30600.0 304350.0 29400.0 303150.0 ;
      RECT  27900.0 331200.0 26700.0 330000.0 ;
      RECT  27900.0 331200.0 26700.0 330000.0 ;
      RECT  27900.0 301650.0 26700.0 300450.0 ;
      RECT  41850.0 304350.0 40650.0 303150.0 ;
      RECT  43800.0 301650.0 42600.0 300450.0 ;
      RECT  45750.0 293550.0 44550.0 292350.0 ;
      RECT  14250.0 304350.0 13050.0 303150.0 ;
      RECT  16200.0 293550.0 15000.0 292350.0 ;
      RECT  18150.0 296250.0 16950.0 295050.0 ;
      RECT  29850.0 322500.0 28650.0 323700.0 ;
      RECT  30600.0 339600.0 29400.0 340800.0 ;
      RECT  16200.0 362100.0 15000.0 363300.0 ;
      RECT  29400.0 342300.0 28200.0 343500.0 ;
      RECT  50400.0 288150.0 49200.0 286950.0 ;
      RECT  36600.0 298950.0 35400.0 297750.0 ;
      RECT  22800.0 288150.0 21600.0 286950.0 ;
      RECT  9000.0 298950.0 7800.0 297750.0 ;
      RECT  49800.0 342450.0 28800.0 343350.0 ;
      RECT  49800.0 362250.0 15600.0 363150.0 ;
      RECT  49800.0 322650.0 29250.0 323550.0 ;
      RECT  49800.0 339750.0 30000.0 340650.0 ;
      RECT  49800.0 303300.0 1.42108547152e-11 304200.0 ;
      RECT  49800.0 284400.0 1.42108547152e-11 285300.0 ;
      RECT  49800.0 297900.0 1.42108547152e-11 298800.0 ;
      RECT  49800.0 287100.0 1.42108547152e-11 288000.0 ;
      RECT  169800.0 342300.0 168600.0 343500.0 ;
      RECT  49500.0 342450.0 48300.0 343650.0 ;
      RECT  167100.0 362100.0 165900.0 363300.0 ;
      RECT  49500.0 362250.0 48300.0 363450.0 ;
      RECT  161700.0 322500.0 160500.0 323700.0 ;
      RECT  49500.0 322650.0 48300.0 323850.0 ;
      RECT  159000.0 339600.0 157800.0 340800.0 ;
      RECT  49500.0 339750.0 48300.0 340950.0 ;
      RECT  164400.0 303150.0 163200.0 304350.0 ;
      RECT  49500.0 303300.0 48300.0 304500.0 ;
      RECT  156300.0 284250.0 155100.0 285450.0 ;
      RECT  49500.0 284400.0 48300.0 285600.0 ;
      RECT  55650.0 297750.0 54450.0 298950.0 ;
      RECT  150900.0 286950.0 149700.0 288150.0 ;
      RECT  49500.0 287100.0 48300.0 288300.0 ;
   LAYER  metal3 ;
      RECT  49800.0 342150.0 169200.0 343650.0 ;
      RECT  49800.0 361950.0 166500.0 363450.0 ;
      RECT  49800.0 322350.0 161100.0 323850.0 ;
      RECT  49800.0 339450.0 158400.0 340950.0 ;
      RECT  49800.0 303000.0 163800.0 304500.0 ;
      RECT  49800.0 284100.0 155700.0 285600.0 ;
      RECT  49800.0 286800.0 150300.0 288300.0 ;
      RECT  176250.0 6300.0 177750.0 151200.0 ;
      RECT  186450.0 6300.0 187950.0 151200.0 ;
      RECT  180000.0 0.0 181500.0 30000.0 ;
      RECT  190200.0 0.0 191700.0 30000.0 ;
      RECT  132000.0 88050.0 148050.0 89550.0 ;
      RECT  132000.0 115650.0 148050.0 117150.0 ;
      RECT  132000.0 143250.0 148050.0 144750.0 ;
      RECT  132000.0 170850.0 148050.0 172350.0 ;
      RECT  176100.0 151200.0 177900.0 153000.0 ;
      RECT  186300.0 151200.0 188100.0 153000.0 ;
      RECT  179700.0 30900.0 181500.0 32700.0 ;
      RECT  189900.0 30900.0 191700.0 32700.0 ;
      RECT  60000.0 79200.0 61800.0 77400.0 ;
      RECT  60000.0 69000.0 61800.0 67200.0 ;
      RECT  60000.0 58800.0 61800.0 57000.0 ;
      RECT  60000.0 48600.0 61800.0 46800.0 ;
      RECT  176250.0 5550.0 178050.0 7350.0 ;
      RECT  186450.0 5550.0 188250.0 7350.0 ;
      RECT  180000.0 0.0 181800.0 1800.0 ;
      RECT  190200.0 0.0 192000.0 1800.0 ;
      RECT  132900.0 87900.0 131100.0 89700.0 ;
      RECT  147150.0 89700.0 148950.0 87900.0 ;
      RECT  132900.0 115500.0 131100.0 117300.0 ;
      RECT  147150.0 117300.0 148950.0 115500.0 ;
      RECT  132900.0 143100.0 131100.0 144900.0 ;
      RECT  147150.0 144900.0 148950.0 143100.0 ;
      RECT  132900.0 170700.0 131100.0 172500.0 ;
      RECT  147150.0 172500.0 148950.0 170700.0 ;
      RECT  52800.0 77400.0 60000.0 78900.0 ;
      RECT  52800.0 67200.0 60000.0 68700.0 ;
      RECT  52800.0 57000.0 60000.0 58500.0 ;
      RECT  52800.0 46800.0 60000.0 48300.0 ;
      RECT  3150.0 262200.0 1650.0 301050.0 ;
      RECT  6600.0 261000.0 5100.0 290250.0 ;
      RECT  18750.0 262200.0 17250.0 292950.0 ;
      RECT  23550.0 262200.0 22050.0 295650.0 ;
      RECT  10950.0 262200.0 9450.0 287550.0 ;
      RECT  31350.0 262200.0 29850.0 287550.0 ;
      RECT  44100.0 243900.0 42600.0 303750.0 ;
      RECT  30750.0 303750.0 29250.0 327600.0 ;
      RECT  28050.0 301050.0 26550.0 330600.0 ;
      RECT  4200.0 203100.0 6000.0 204900.0 ;
      RECT  14400.0 203100.0 16200.0 204900.0 ;
      RECT  24600.0 203100.0 26400.0 204900.0 ;
      RECT  3300.0 263100.0 1500.0 261300.0 ;
      RECT  3300.0 301950.0 1500.0 300150.0 ;
      RECT  6750.0 261900.0 4950.0 260100.0 ;
      RECT  6750.0 291150.0 4950.0 289350.0 ;
      RECT  18900.0 263100.0 17100.0 261300.0 ;
      RECT  18900.0 293850.0 17100.0 292050.0 ;
      RECT  23700.0 263100.0 21900.0 261300.0 ;
      RECT  23700.0 296550.0 21900.0 294750.0 ;
      RECT  11100.0 263100.0 9300.0 261300.0 ;
      RECT  11100.0 288450.0 9300.0 286650.0 ;
      RECT  31500.0 263100.0 29700.0 261300.0 ;
      RECT  31500.0 288450.0 29700.0 286650.0 ;
      RECT  44250.0 244800.0 42450.0 243000.0 ;
      RECT  44250.0 304650.0 42450.0 302850.0 ;
      RECT  30900.0 328500.0 29100.0 326700.0 ;
      RECT  30900.0 304650.0 29100.0 302850.0 ;
      RECT  28200.0 331500.0 26400.0 329700.0 ;
      RECT  28200.0 301950.0 26400.0 300150.0 ;
      RECT  16200.0 203100.0 14400.0 204900.0 ;
      RECT  26400.0 203100.0 24600.0 204900.0 ;
      RECT  6000.0 203100.0 4200.0 204900.0 ;
      RECT  170100.0 342000.0 168300.0 343800.0 ;
      RECT  49800.0 342150.0 48000.0 343950.0 ;
      RECT  167400.0 361800.0 165600.0 363600.0 ;
      RECT  49800.0 361950.0 48000.0 363750.0 ;
      RECT  162000.0 322200.0 160200.0 324000.0 ;
      RECT  49800.0 322350.0 48000.0 324150.0 ;
      RECT  159300.0 339300.0 157500.0 341100.0 ;
      RECT  49800.0 339450.0 48000.0 341250.0 ;
      RECT  164700.0 302850.0 162900.0 304650.0 ;
      RECT  49800.0 303000.0 48000.0 304800.0 ;
      RECT  156600.0 283950.0 154800.0 285750.0 ;
      RECT  49800.0 284100.0 48000.0 285900.0 ;
      RECT  151200.0 286650.0 149400.0 288450.0 ;
      RECT  49800.0 286800.0 48000.0 288600.0 ;
   END
   END    sram_2_16_1_scn3me_subm
END    LIBRARY
