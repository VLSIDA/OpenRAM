magic
tech sky130A
magscale 1 2
timestamp 1595931502
<< checkpaint >>
rect -1302 -1364 2550 7684
<< ndiffc >>
rect 42 6256 76 6258
rect 1172 6256 1206 6258
rect 42 6224 76 6226
rect 1172 6224 1206 6226
rect 14 6067 17 6099
rect 463 6067 466 6099
rect 596 6067 599 6099
rect 649 6067 652 6099
rect 782 6067 785 6099
rect 1231 6067 1234 6099
rect 42 5908 76 5942
rect 404 5908 438 5942
rect 810 5908 844 5942
rect 1172 5908 1206 5942
rect 14 5751 17 5783
rect 463 5751 466 5783
rect 596 5751 599 5783
rect 649 5751 652 5783
rect 782 5751 785 5783
rect 1231 5751 1234 5783
rect 42 5624 76 5626
rect 1172 5624 1206 5626
rect 42 5592 76 5594
rect 1172 5592 1206 5594
rect 42 5466 76 5468
rect 1172 5466 1206 5468
rect 42 5434 76 5436
rect 1172 5434 1206 5436
rect 14 5277 17 5309
rect 463 5277 466 5309
rect 596 5277 599 5309
rect 649 5277 652 5309
rect 782 5277 785 5309
rect 1231 5277 1234 5309
rect 42 5118 76 5152
rect 404 5118 438 5152
rect 810 5118 844 5152
rect 1172 5118 1206 5152
rect 14 4961 17 4993
rect 463 4961 466 4993
rect 596 4961 599 4993
rect 649 4961 652 4993
rect 782 4961 785 4993
rect 1231 4961 1234 4993
rect 42 4834 76 4836
rect 1172 4834 1206 4836
rect 42 4802 76 4804
rect 1172 4802 1206 4804
rect 42 4676 76 4678
rect 1172 4676 1206 4678
rect 42 4644 76 4646
rect 1172 4644 1206 4646
rect 14 4487 17 4519
rect 463 4487 466 4519
rect 596 4487 599 4519
rect 649 4487 652 4519
rect 782 4487 785 4519
rect 1231 4487 1234 4519
rect 42 4328 76 4362
rect 404 4328 438 4362
rect 810 4328 844 4362
rect 1172 4328 1206 4362
rect 14 4171 17 4203
rect 463 4171 466 4203
rect 596 4171 599 4203
rect 649 4171 652 4203
rect 782 4171 785 4203
rect 1231 4171 1234 4203
rect 42 4044 76 4046
rect 1172 4044 1206 4046
rect 42 4012 76 4014
rect 1172 4012 1206 4014
rect 42 3886 76 3888
rect 1172 3886 1206 3888
rect 42 3854 76 3856
rect 1172 3854 1206 3856
rect 14 3697 17 3729
rect 463 3697 466 3729
rect 596 3697 599 3729
rect 649 3697 652 3729
rect 782 3697 785 3729
rect 1231 3697 1234 3729
rect 42 3538 76 3572
rect 404 3538 438 3572
rect 810 3538 844 3572
rect 1172 3538 1206 3572
rect 14 3381 17 3413
rect 463 3381 466 3413
rect 596 3381 599 3413
rect 649 3381 652 3413
rect 782 3381 785 3413
rect 1231 3381 1234 3413
rect 42 3254 76 3256
rect 1172 3254 1206 3256
rect 42 3222 76 3224
rect 1172 3222 1206 3224
rect 42 3096 76 3098
rect 1172 3096 1206 3098
rect 42 3064 76 3066
rect 1172 3064 1206 3066
rect 14 2907 17 2939
rect 463 2907 466 2939
rect 596 2907 599 2939
rect 649 2907 652 2939
rect 782 2907 785 2939
rect 1231 2907 1234 2939
rect 42 2748 76 2782
rect 404 2748 438 2782
rect 810 2748 844 2782
rect 1172 2748 1206 2782
rect 14 2591 17 2623
rect 463 2591 466 2623
rect 596 2591 599 2623
rect 649 2591 652 2623
rect 782 2591 785 2623
rect 1231 2591 1234 2623
rect 42 2464 76 2466
rect 1172 2464 1206 2466
rect 42 2432 76 2434
rect 1172 2432 1206 2434
rect 42 2306 76 2308
rect 1172 2306 1206 2308
rect 42 2274 76 2276
rect 1172 2274 1206 2276
rect 14 2117 17 2149
rect 463 2117 466 2149
rect 596 2117 599 2149
rect 649 2117 652 2149
rect 782 2117 785 2149
rect 1231 2117 1234 2149
rect 42 1958 76 1992
rect 404 1958 438 1992
rect 810 1958 844 1992
rect 1172 1958 1206 1992
rect 14 1801 17 1833
rect 463 1801 466 1833
rect 596 1801 599 1833
rect 649 1801 652 1833
rect 782 1801 785 1833
rect 1231 1801 1234 1833
rect 42 1674 76 1676
rect 1172 1674 1206 1676
rect 42 1642 76 1644
rect 1172 1642 1206 1644
rect 42 1516 76 1518
rect 1172 1516 1206 1518
rect 42 1484 76 1486
rect 1172 1484 1206 1486
rect 14 1327 17 1359
rect 463 1327 466 1359
rect 596 1327 599 1359
rect 649 1327 652 1359
rect 782 1327 785 1359
rect 1231 1327 1234 1359
rect 42 1168 76 1202
rect 404 1168 438 1202
rect 810 1168 844 1202
rect 1172 1168 1206 1202
rect 14 1011 17 1043
rect 463 1011 466 1043
rect 596 1011 599 1043
rect 649 1011 652 1043
rect 782 1011 785 1043
rect 1231 1011 1234 1043
rect 42 884 76 886
rect 1172 884 1206 886
rect 42 852 76 854
rect 1172 852 1206 854
rect 42 726 76 728
rect 1172 726 1206 728
rect 42 694 76 696
rect 1172 694 1206 696
rect 14 537 17 569
rect 463 537 466 569
rect 596 537 599 569
rect 649 537 652 569
rect 782 537 785 569
rect 1231 537 1234 569
rect 42 378 76 412
rect 404 378 438 412
rect 810 378 844 412
rect 1172 378 1206 412
rect 14 221 17 253
rect 463 221 466 253
rect 596 221 599 253
rect 649 221 652 253
rect 782 221 785 253
rect 1231 221 1234 253
rect 42 94 76 96
rect 1172 94 1206 96
rect 42 62 76 64
rect 1172 62 1206 64
<< locali >>
rect 193 6147 196 6181
rect 224 6147 227 6181
rect 1021 6147 1024 6181
rect 1052 6147 1055 6181
rect -14 6099 14 6100
rect -14 6067 0 6099
rect 107 6079 109 6107
rect 139 6079 141 6113
rect -14 6066 14 6067
rect 193 6066 196 6100
rect 224 6066 227 6100
rect 466 6099 497 6100
rect 565 6099 596 6100
rect 652 6099 683 6100
rect 751 6099 782 6100
rect 271 6062 278 6096
rect 339 6053 341 6087
rect 371 6059 373 6087
rect 466 6066 497 6067
rect 565 6066 596 6067
rect 652 6066 683 6067
rect 751 6066 782 6067
rect 875 6059 877 6087
rect 907 6053 909 6087
rect 970 6062 977 6096
rect 1021 6066 1024 6100
rect 1052 6066 1055 6100
rect 1107 6079 1109 6113
rect 1139 6079 1141 6107
rect 1234 6099 1262 6100
rect 1248 6067 1262 6099
rect 1234 6066 1262 6067
rect 193 5985 196 6019
rect 224 5985 227 6019
rect 1021 5985 1024 6019
rect 1052 5985 1055 6019
rect 193 5831 196 5865
rect 224 5831 227 5865
rect 1021 5831 1024 5865
rect 1052 5831 1055 5865
rect -14 5783 14 5784
rect -14 5751 0 5783
rect -14 5750 14 5751
rect 107 5743 109 5771
rect 139 5737 141 5771
rect 193 5750 196 5784
rect 224 5750 227 5784
rect 271 5754 278 5788
rect 339 5763 341 5797
rect 371 5763 373 5791
rect 466 5783 497 5784
rect 565 5783 596 5784
rect 652 5783 683 5784
rect 751 5783 782 5784
rect 875 5763 877 5791
rect 907 5763 909 5797
rect 970 5754 977 5788
rect 466 5750 497 5751
rect 565 5750 596 5751
rect 652 5750 683 5751
rect 751 5750 782 5751
rect 1021 5750 1024 5784
rect 1052 5750 1055 5784
rect 1234 5783 1262 5784
rect 1107 5737 1109 5771
rect 1139 5743 1141 5771
rect 1248 5751 1262 5783
rect 1234 5750 1262 5751
rect 193 5669 196 5703
rect 224 5669 227 5703
rect 1021 5669 1024 5703
rect 1052 5669 1055 5703
rect 193 5357 196 5391
rect 224 5357 227 5391
rect 1021 5357 1024 5391
rect 1052 5357 1055 5391
rect -14 5309 14 5310
rect -14 5277 0 5309
rect 107 5289 109 5317
rect 139 5289 141 5323
rect -14 5276 14 5277
rect 193 5276 196 5310
rect 224 5276 227 5310
rect 466 5309 497 5310
rect 565 5309 596 5310
rect 652 5309 683 5310
rect 751 5309 782 5310
rect 271 5272 278 5306
rect 339 5263 341 5297
rect 371 5269 373 5297
rect 466 5276 497 5277
rect 565 5276 596 5277
rect 652 5276 683 5277
rect 751 5276 782 5277
rect 875 5269 877 5297
rect 907 5263 909 5297
rect 970 5272 977 5306
rect 1021 5276 1024 5310
rect 1052 5276 1055 5310
rect 1107 5289 1109 5323
rect 1139 5289 1141 5317
rect 1234 5309 1262 5310
rect 1248 5277 1262 5309
rect 1234 5276 1262 5277
rect 193 5195 196 5229
rect 224 5195 227 5229
rect 1021 5195 1024 5229
rect 1052 5195 1055 5229
rect 193 5041 196 5075
rect 224 5041 227 5075
rect 1021 5041 1024 5075
rect 1052 5041 1055 5075
rect -14 4993 14 4994
rect -14 4961 0 4993
rect -14 4960 14 4961
rect 107 4953 109 4981
rect 139 4947 141 4981
rect 193 4960 196 4994
rect 224 4960 227 4994
rect 271 4964 278 4998
rect 339 4973 341 5007
rect 371 4973 373 5001
rect 466 4993 497 4994
rect 565 4993 596 4994
rect 652 4993 683 4994
rect 751 4993 782 4994
rect 875 4973 877 5001
rect 907 4973 909 5007
rect 970 4964 977 4998
rect 466 4960 497 4961
rect 565 4960 596 4961
rect 652 4960 683 4961
rect 751 4960 782 4961
rect 1021 4960 1024 4994
rect 1052 4960 1055 4994
rect 1234 4993 1262 4994
rect 1107 4947 1109 4981
rect 1139 4953 1141 4981
rect 1248 4961 1262 4993
rect 1234 4960 1262 4961
rect 193 4879 196 4913
rect 224 4879 227 4913
rect 1021 4879 1024 4913
rect 1052 4879 1055 4913
rect 193 4567 196 4601
rect 224 4567 227 4601
rect 1021 4567 1024 4601
rect 1052 4567 1055 4601
rect -14 4519 14 4520
rect -14 4487 0 4519
rect 107 4499 109 4527
rect 139 4499 141 4533
rect -14 4486 14 4487
rect 193 4486 196 4520
rect 224 4486 227 4520
rect 466 4519 497 4520
rect 565 4519 596 4520
rect 652 4519 683 4520
rect 751 4519 782 4520
rect 271 4482 278 4516
rect 339 4473 341 4507
rect 371 4479 373 4507
rect 466 4486 497 4487
rect 565 4486 596 4487
rect 652 4486 683 4487
rect 751 4486 782 4487
rect 875 4479 877 4507
rect 907 4473 909 4507
rect 970 4482 977 4516
rect 1021 4486 1024 4520
rect 1052 4486 1055 4520
rect 1107 4499 1109 4533
rect 1139 4499 1141 4527
rect 1234 4519 1262 4520
rect 1248 4487 1262 4519
rect 1234 4486 1262 4487
rect 193 4405 196 4439
rect 224 4405 227 4439
rect 1021 4405 1024 4439
rect 1052 4405 1055 4439
rect 193 4251 196 4285
rect 224 4251 227 4285
rect 1021 4251 1024 4285
rect 1052 4251 1055 4285
rect -14 4203 14 4204
rect -14 4171 0 4203
rect -14 4170 14 4171
rect 107 4163 109 4191
rect 139 4157 141 4191
rect 193 4170 196 4204
rect 224 4170 227 4204
rect 271 4174 278 4208
rect 339 4183 341 4217
rect 371 4183 373 4211
rect 466 4203 497 4204
rect 565 4203 596 4204
rect 652 4203 683 4204
rect 751 4203 782 4204
rect 875 4183 877 4211
rect 907 4183 909 4217
rect 970 4174 977 4208
rect 466 4170 497 4171
rect 565 4170 596 4171
rect 652 4170 683 4171
rect 751 4170 782 4171
rect 1021 4170 1024 4204
rect 1052 4170 1055 4204
rect 1234 4203 1262 4204
rect 1107 4157 1109 4191
rect 1139 4163 1141 4191
rect 1248 4171 1262 4203
rect 1234 4170 1262 4171
rect 193 4089 196 4123
rect 224 4089 227 4123
rect 1021 4089 1024 4123
rect 1052 4089 1055 4123
rect 193 3777 196 3811
rect 224 3777 227 3811
rect 1021 3777 1024 3811
rect 1052 3777 1055 3811
rect -14 3729 14 3730
rect -14 3697 0 3729
rect 107 3709 109 3737
rect 139 3709 141 3743
rect -14 3696 14 3697
rect 193 3696 196 3730
rect 224 3696 227 3730
rect 466 3729 497 3730
rect 565 3729 596 3730
rect 652 3729 683 3730
rect 751 3729 782 3730
rect 271 3692 278 3726
rect 339 3683 341 3717
rect 371 3689 373 3717
rect 466 3696 497 3697
rect 565 3696 596 3697
rect 652 3696 683 3697
rect 751 3696 782 3697
rect 875 3689 877 3717
rect 907 3683 909 3717
rect 970 3692 977 3726
rect 1021 3696 1024 3730
rect 1052 3696 1055 3730
rect 1107 3709 1109 3743
rect 1139 3709 1141 3737
rect 1234 3729 1262 3730
rect 1248 3697 1262 3729
rect 1234 3696 1262 3697
rect 193 3615 196 3649
rect 224 3615 227 3649
rect 1021 3615 1024 3649
rect 1052 3615 1055 3649
rect 193 3461 196 3495
rect 224 3461 227 3495
rect 1021 3461 1024 3495
rect 1052 3461 1055 3495
rect -14 3413 14 3414
rect -14 3381 0 3413
rect -14 3380 14 3381
rect 107 3373 109 3401
rect 139 3367 141 3401
rect 193 3380 196 3414
rect 224 3380 227 3414
rect 271 3384 278 3418
rect 339 3393 341 3427
rect 371 3393 373 3421
rect 466 3413 497 3414
rect 565 3413 596 3414
rect 652 3413 683 3414
rect 751 3413 782 3414
rect 875 3393 877 3421
rect 907 3393 909 3427
rect 970 3384 977 3418
rect 466 3380 497 3381
rect 565 3380 596 3381
rect 652 3380 683 3381
rect 751 3380 782 3381
rect 1021 3380 1024 3414
rect 1052 3380 1055 3414
rect 1234 3413 1262 3414
rect 1107 3367 1109 3401
rect 1139 3373 1141 3401
rect 1248 3381 1262 3413
rect 1234 3380 1262 3381
rect 193 3299 196 3333
rect 224 3299 227 3333
rect 1021 3299 1024 3333
rect 1052 3299 1055 3333
rect 193 2987 196 3021
rect 224 2987 227 3021
rect 1021 2987 1024 3021
rect 1052 2987 1055 3021
rect -14 2939 14 2940
rect -14 2907 0 2939
rect 107 2919 109 2947
rect 139 2919 141 2953
rect -14 2906 14 2907
rect 193 2906 196 2940
rect 224 2906 227 2940
rect 466 2939 497 2940
rect 565 2939 596 2940
rect 652 2939 683 2940
rect 751 2939 782 2940
rect 271 2902 278 2936
rect 339 2893 341 2927
rect 371 2899 373 2927
rect 466 2906 497 2907
rect 565 2906 596 2907
rect 652 2906 683 2907
rect 751 2906 782 2907
rect 875 2899 877 2927
rect 907 2893 909 2927
rect 970 2902 977 2936
rect 1021 2906 1024 2940
rect 1052 2906 1055 2940
rect 1107 2919 1109 2953
rect 1139 2919 1141 2947
rect 1234 2939 1262 2940
rect 1248 2907 1262 2939
rect 1234 2906 1262 2907
rect 193 2825 196 2859
rect 224 2825 227 2859
rect 1021 2825 1024 2859
rect 1052 2825 1055 2859
rect 193 2671 196 2705
rect 224 2671 227 2705
rect 1021 2671 1024 2705
rect 1052 2671 1055 2705
rect -14 2623 14 2624
rect -14 2591 0 2623
rect -14 2590 14 2591
rect 107 2583 109 2611
rect 139 2577 141 2611
rect 193 2590 196 2624
rect 224 2590 227 2624
rect 271 2594 278 2628
rect 339 2603 341 2637
rect 371 2603 373 2631
rect 466 2623 497 2624
rect 565 2623 596 2624
rect 652 2623 683 2624
rect 751 2623 782 2624
rect 875 2603 877 2631
rect 907 2603 909 2637
rect 970 2594 977 2628
rect 466 2590 497 2591
rect 565 2590 596 2591
rect 652 2590 683 2591
rect 751 2590 782 2591
rect 1021 2590 1024 2624
rect 1052 2590 1055 2624
rect 1234 2623 1262 2624
rect 1107 2577 1109 2611
rect 1139 2583 1141 2611
rect 1248 2591 1262 2623
rect 1234 2590 1262 2591
rect 193 2509 196 2543
rect 224 2509 227 2543
rect 1021 2509 1024 2543
rect 1052 2509 1055 2543
rect 193 2197 196 2231
rect 224 2197 227 2231
rect 1021 2197 1024 2231
rect 1052 2197 1055 2231
rect -14 2149 14 2150
rect -14 2117 0 2149
rect 107 2129 109 2157
rect 139 2129 141 2163
rect -14 2116 14 2117
rect 193 2116 196 2150
rect 224 2116 227 2150
rect 466 2149 497 2150
rect 565 2149 596 2150
rect 652 2149 683 2150
rect 751 2149 782 2150
rect 271 2112 278 2146
rect 339 2103 341 2137
rect 371 2109 373 2137
rect 466 2116 497 2117
rect 565 2116 596 2117
rect 652 2116 683 2117
rect 751 2116 782 2117
rect 875 2109 877 2137
rect 907 2103 909 2137
rect 970 2112 977 2146
rect 1021 2116 1024 2150
rect 1052 2116 1055 2150
rect 1107 2129 1109 2163
rect 1139 2129 1141 2157
rect 1234 2149 1262 2150
rect 1248 2117 1262 2149
rect 1234 2116 1262 2117
rect 193 2035 196 2069
rect 224 2035 227 2069
rect 1021 2035 1024 2069
rect 1052 2035 1055 2069
rect 193 1881 196 1915
rect 224 1881 227 1915
rect 1021 1881 1024 1915
rect 1052 1881 1055 1915
rect -14 1833 14 1834
rect -14 1801 0 1833
rect -14 1800 14 1801
rect 107 1793 109 1821
rect 139 1787 141 1821
rect 193 1800 196 1834
rect 224 1800 227 1834
rect 271 1804 278 1838
rect 339 1813 341 1847
rect 371 1813 373 1841
rect 466 1833 497 1834
rect 565 1833 596 1834
rect 652 1833 683 1834
rect 751 1833 782 1834
rect 875 1813 877 1841
rect 907 1813 909 1847
rect 970 1804 977 1838
rect 466 1800 497 1801
rect 565 1800 596 1801
rect 652 1800 683 1801
rect 751 1800 782 1801
rect 1021 1800 1024 1834
rect 1052 1800 1055 1834
rect 1234 1833 1262 1834
rect 1107 1787 1109 1821
rect 1139 1793 1141 1821
rect 1248 1801 1262 1833
rect 1234 1800 1262 1801
rect 193 1719 196 1753
rect 224 1719 227 1753
rect 1021 1719 1024 1753
rect 1052 1719 1055 1753
rect 193 1407 196 1441
rect 224 1407 227 1441
rect 1021 1407 1024 1441
rect 1052 1407 1055 1441
rect -14 1359 14 1360
rect -14 1327 0 1359
rect 107 1339 109 1367
rect 139 1339 141 1373
rect -14 1326 14 1327
rect 193 1326 196 1360
rect 224 1326 227 1360
rect 466 1359 497 1360
rect 565 1359 596 1360
rect 652 1359 683 1360
rect 751 1359 782 1360
rect 271 1322 278 1356
rect 339 1313 341 1347
rect 371 1319 373 1347
rect 466 1326 497 1327
rect 565 1326 596 1327
rect 652 1326 683 1327
rect 751 1326 782 1327
rect 875 1319 877 1347
rect 907 1313 909 1347
rect 970 1322 977 1356
rect 1021 1326 1024 1360
rect 1052 1326 1055 1360
rect 1107 1339 1109 1373
rect 1139 1339 1141 1367
rect 1234 1359 1262 1360
rect 1248 1327 1262 1359
rect 1234 1326 1262 1327
rect 193 1245 196 1279
rect 224 1245 227 1279
rect 1021 1245 1024 1279
rect 1052 1245 1055 1279
rect 193 1091 196 1125
rect 224 1091 227 1125
rect 1021 1091 1024 1125
rect 1052 1091 1055 1125
rect -14 1043 14 1044
rect -14 1011 0 1043
rect -14 1010 14 1011
rect 107 1003 109 1031
rect 139 997 141 1031
rect 193 1010 196 1044
rect 224 1010 227 1044
rect 271 1014 278 1048
rect 339 1023 341 1057
rect 371 1023 373 1051
rect 466 1043 497 1044
rect 565 1043 596 1044
rect 652 1043 683 1044
rect 751 1043 782 1044
rect 875 1023 877 1051
rect 907 1023 909 1057
rect 970 1014 977 1048
rect 466 1010 497 1011
rect 565 1010 596 1011
rect 652 1010 683 1011
rect 751 1010 782 1011
rect 1021 1010 1024 1044
rect 1052 1010 1055 1044
rect 1234 1043 1262 1044
rect 1107 997 1109 1031
rect 1139 1003 1141 1031
rect 1248 1011 1262 1043
rect 1234 1010 1262 1011
rect 193 929 196 963
rect 224 929 227 963
rect 1021 929 1024 963
rect 1052 929 1055 963
rect 193 617 196 651
rect 224 617 227 651
rect 1021 617 1024 651
rect 1052 617 1055 651
rect -14 569 14 570
rect -14 537 0 569
rect 107 549 109 577
rect 139 549 141 583
rect -14 536 14 537
rect 193 536 196 570
rect 224 536 227 570
rect 466 569 497 570
rect 565 569 596 570
rect 652 569 683 570
rect 751 569 782 570
rect 271 532 278 566
rect 339 523 341 557
rect 371 529 373 557
rect 466 536 497 537
rect 565 536 596 537
rect 652 536 683 537
rect 751 536 782 537
rect 875 529 877 557
rect 907 523 909 557
rect 970 532 977 566
rect 1021 536 1024 570
rect 1052 536 1055 570
rect 1107 549 1109 583
rect 1139 549 1141 577
rect 1234 569 1262 570
rect 1248 537 1262 569
rect 1234 536 1262 537
rect 193 455 196 489
rect 224 455 227 489
rect 1021 455 1024 489
rect 1052 455 1055 489
rect 193 301 196 335
rect 224 301 227 335
rect 1021 301 1024 335
rect 1052 301 1055 335
rect -14 253 14 254
rect -14 221 0 253
rect -14 220 14 221
rect 107 213 109 241
rect 139 207 141 241
rect 193 220 196 254
rect 224 220 227 254
rect 271 224 278 258
rect 339 233 341 267
rect 371 233 373 261
rect 466 253 497 254
rect 565 253 596 254
rect 652 253 683 254
rect 751 253 782 254
rect 875 233 877 261
rect 907 233 909 267
rect 970 224 977 258
rect 466 220 497 221
rect 565 220 596 221
rect 652 220 683 221
rect 751 220 782 221
rect 1021 220 1024 254
rect 1052 220 1055 254
rect 1234 253 1262 254
rect 1107 207 1109 241
rect 1139 213 1141 241
rect 1248 221 1262 253
rect 1234 220 1262 221
rect 193 139 196 173
rect 224 139 227 173
rect 1021 139 1024 173
rect 1052 139 1055 173
<< metal1 >>
rect 78 0 114 6320
rect 150 0 186 6320
rect 222 5609 258 6241
rect 222 4819 258 5451
rect 222 4029 258 4661
rect 222 3239 258 3871
rect 222 2449 258 3081
rect 222 1659 258 2291
rect 222 869 258 1501
rect 222 79 258 711
rect 294 0 330 6320
rect 366 0 402 6320
rect 846 0 882 6320
rect 918 0 954 6320
rect 990 5609 1026 6241
rect 990 4819 1026 5451
rect 990 4029 1026 4661
rect 990 3239 1026 3871
rect 990 2449 1026 3081
rect 990 1659 1026 2291
rect 990 869 1026 1501
rect 990 79 1026 711
rect 1062 0 1098 6320
rect 1134 0 1170 6320
<< metal2 >>
rect 186 6265 294 6375
rect 954 6265 1062 6375
rect 0 6169 1248 6217
rect 186 6045 294 6121
rect 954 6045 1062 6121
rect 0 5949 1248 5997
rect 0 5853 1248 5901
rect 186 5729 294 5805
rect 954 5729 1062 5805
rect 0 5633 1248 5681
rect 186 5475 294 5585
rect 954 5475 1062 5585
rect 0 5379 1248 5427
rect 186 5255 294 5331
rect 954 5255 1062 5331
rect 0 5159 1248 5207
rect 0 5063 1248 5111
rect 186 4939 294 5015
rect 954 4939 1062 5015
rect 0 4843 1248 4891
rect 186 4685 294 4795
rect 954 4685 1062 4795
rect 0 4589 1248 4637
rect 186 4465 294 4541
rect 954 4465 1062 4541
rect 0 4369 1248 4417
rect 0 4273 1248 4321
rect 186 4149 294 4225
rect 954 4149 1062 4225
rect 0 4053 1248 4101
rect 186 3895 294 4005
rect 954 3895 1062 4005
rect 0 3799 1248 3847
rect 186 3675 294 3751
rect 954 3675 1062 3751
rect 0 3579 1248 3627
rect 0 3483 1248 3531
rect 186 3359 294 3435
rect 954 3359 1062 3435
rect 0 3263 1248 3311
rect 186 3105 294 3215
rect 954 3105 1062 3215
rect 0 3009 1248 3057
rect 186 2885 294 2961
rect 954 2885 1062 2961
rect 0 2789 1248 2837
rect 0 2693 1248 2741
rect 186 2569 294 2645
rect 954 2569 1062 2645
rect 0 2473 1248 2521
rect 186 2315 294 2425
rect 954 2315 1062 2425
rect 0 2219 1248 2267
rect 186 2095 294 2171
rect 954 2095 1062 2171
rect 0 1999 1248 2047
rect 0 1903 1248 1951
rect 186 1779 294 1855
rect 954 1779 1062 1855
rect 0 1683 1248 1731
rect 186 1525 294 1635
rect 954 1525 1062 1635
rect 0 1429 1248 1477
rect 186 1305 294 1381
rect 954 1305 1062 1381
rect 0 1209 1248 1257
rect 0 1113 1248 1161
rect 186 989 294 1065
rect 954 989 1062 1065
rect 0 893 1248 941
rect 186 735 294 845
rect 954 735 1062 845
rect 0 639 1248 687
rect 186 515 294 591
rect 954 515 1062 591
rect 0 419 1248 467
rect 0 323 1248 371
rect 186 199 294 275
rect 954 199 1062 275
rect 0 103 1248 151
rect 186 -55 294 55
rect 954 -55 1062 55
use cell_1rw_1r  cell_1rw_1r_0
timestamp 1595931502
transform -1 0 1248 0 -1 6320
box -42 -104 624 420
use cell_1rw_1r  cell_1rw_1r_1
timestamp 1595931502
transform -1 0 1248 0 1 5530
box -42 -104 624 420
use cell_1rw_1r  cell_1rw_1r_2
timestamp 1595931502
transform -1 0 1248 0 -1 5530
box -42 -104 624 420
use cell_1rw_1r  cell_1rw_1r_3
timestamp 1595931502
transform -1 0 1248 0 1 4740
box -42 -104 624 420
use cell_1rw_1r  cell_1rw_1r_4
timestamp 1595931502
transform -1 0 1248 0 -1 4740
box -42 -104 624 420
use cell_1rw_1r  cell_1rw_1r_5
timestamp 1595931502
transform -1 0 1248 0 1 3950
box -42 -104 624 420
use cell_1rw_1r  cell_1rw_1r_6
timestamp 1595931502
transform -1 0 1248 0 -1 3950
box -42 -104 624 420
use cell_1rw_1r  cell_1rw_1r_7
timestamp 1595931502
transform -1 0 1248 0 1 3160
box -42 -104 624 420
use cell_1rw_1r  cell_1rw_1r_8
timestamp 1595931502
transform -1 0 1248 0 -1 3160
box -42 -104 624 420
use cell_1rw_1r  cell_1rw_1r_9
timestamp 1595931502
transform -1 0 1248 0 1 2370
box -42 -104 624 420
use cell_1rw_1r  cell_1rw_1r_10
timestamp 1595931502
transform -1 0 1248 0 -1 2370
box -42 -104 624 420
use cell_1rw_1r  cell_1rw_1r_11
timestamp 1595931502
transform -1 0 1248 0 1 1580
box -42 -104 624 420
use cell_1rw_1r  cell_1rw_1r_12
timestamp 1595931502
transform -1 0 1248 0 -1 1580
box -42 -104 624 420
use cell_1rw_1r  cell_1rw_1r_13
timestamp 1595931502
transform -1 0 1248 0 1 790
box -42 -104 624 420
use cell_1rw_1r  cell_1rw_1r_14
timestamp 1595931502
transform -1 0 1248 0 -1 790
box -42 -104 624 420
use cell_1rw_1r  cell_1rw_1r_15
timestamp 1595931502
transform -1 0 1248 0 1 0
box -42 -104 624 420
use cell_1rw_1r  cell_1rw_1r_16
timestamp 1595931502
transform 1 0 0 0 -1 6320
box -42 -104 624 420
use cell_1rw_1r  cell_1rw_1r_17
timestamp 1595931502
transform 1 0 0 0 1 5530
box -42 -104 624 420
use cell_1rw_1r  cell_1rw_1r_18
timestamp 1595931502
transform 1 0 0 0 -1 5530
box -42 -104 624 420
use cell_1rw_1r  cell_1rw_1r_19
timestamp 1595931502
transform 1 0 0 0 1 4740
box -42 -104 624 420
use cell_1rw_1r  cell_1rw_1r_20
timestamp 1595931502
transform 1 0 0 0 -1 4740
box -42 -104 624 420
use cell_1rw_1r  cell_1rw_1r_21
timestamp 1595931502
transform 1 0 0 0 1 3950
box -42 -104 624 420
use cell_1rw_1r  cell_1rw_1r_22
timestamp 1595931502
transform 1 0 0 0 -1 3950
box -42 -104 624 420
use cell_1rw_1r  cell_1rw_1r_23
timestamp 1595931502
transform 1 0 0 0 1 3160
box -42 -104 624 420
use cell_1rw_1r  cell_1rw_1r_24
timestamp 1595931502
transform 1 0 0 0 -1 3160
box -42 -104 624 420
use cell_1rw_1r  cell_1rw_1r_25
timestamp 1595931502
transform 1 0 0 0 1 2370
box -42 -104 624 420
use cell_1rw_1r  cell_1rw_1r_26
timestamp 1595931502
transform 1 0 0 0 -1 2370
box -42 -104 624 420
use cell_1rw_1r  cell_1rw_1r_27
timestamp 1595931502
transform 1 0 0 0 1 1580
box -42 -104 624 420
use cell_1rw_1r  cell_1rw_1r_28
timestamp 1595931502
transform 1 0 0 0 -1 1580
box -42 -104 624 420
use cell_1rw_1r  cell_1rw_1r_29
timestamp 1595931502
transform 1 0 0 0 1 790
box -42 -104 624 420
use cell_1rw_1r  cell_1rw_1r_30
timestamp 1595931502
transform 1 0 0 0 -1 790
box -42 -104 624 420
use cell_1rw_1r  cell_1rw_1r_31
timestamp 1595931502
transform 1 0 0 0 1 0
box -42 -104 624 420
<< labels >>
rlabel metal1 s 168 3160 168 3160 4 br0_0
rlabel metal2 s 624 4613 624 4613 4 wl1_11
rlabel metal1 s 1080 3160 1080 3160 4 br0_1
rlabel metal1 s 384 3160 384 3160 4 br1_0
rlabel metal2 s 624 917 624 917 4 wl1_2
rlabel metal2 s 624 5403 624 5403 4 wl1_13
rlabel metal1 s 936 3160 936 3160 4 bl1_1
rlabel metal2 s 624 1927 624 1927 4 wl0_4
rlabel metal2 s 624 3823 624 3823 4 wl1_9
rlabel metal2 s 624 347 624 347 4 wl0_0
rlabel metal2 s 624 1137 624 1137 4 wl0_2
rlabel metal2 s 624 3033 624 3033 4 wl1_7
rlabel metal2 s 624 663 624 663 4 wl1_1
rlabel metal2 s 624 5657 624 5657 4 wl1_14
rlabel metal2 s 624 4393 624 4393 4 wl0_11
rlabel metal1 s 864 3160 864 3160 4 br1_1
rlabel metal2 s 624 6193 624 6193 4 wl1_15
rlabel metal2 s 624 4077 624 4077 4 wl1_10
rlabel metal2 s 624 1707 624 1707 4 wl1_4
rlabel metal2 s 624 1233 624 1233 4 wl0_3
rlabel metal2 s 1008 6083 1008 6083 4 gnd
rlabel metal2 s 240 3397 240 3397 4 gnd
rlabel metal2 s 240 1027 240 1027 4 gnd
rlabel metal2 s 240 237 240 237 4 gnd
rlabel metal2 s 240 3713 240 3713 4 gnd
rlabel metal2 s 240 553 240 553 4 gnd
rlabel metal2 s 1008 5767 1008 5767 4 gnd
rlabel metal2 s 240 3160 240 3160 4 gnd
rlabel metal2 s 1008 4740 1008 4740 4 gnd
rlabel metal2 s 1008 5530 1008 5530 4 gnd
rlabel metal2 s 1008 1027 1008 1027 4 gnd
rlabel metal2 s 240 2923 240 2923 4 gnd
rlabel metal2 s 240 0 240 0 4 gnd
rlabel metal2 s 1008 3950 1008 3950 4 gnd
rlabel metal2 s 240 4187 240 4187 4 gnd
rlabel metal2 s 240 4740 240 4740 4 gnd
rlabel metal2 s 240 5767 240 5767 4 gnd
rlabel metal2 s 240 1343 240 1343 4 gnd
rlabel metal2 s 1008 1580 1008 1580 4 gnd
rlabel metal2 s 240 2133 240 2133 4 gnd
rlabel metal2 s 1008 237 1008 237 4 gnd
rlabel metal2 s 1008 1817 1008 1817 4 gnd
rlabel metal2 s 1008 3397 1008 3397 4 gnd
rlabel metal2 s 240 6320 240 6320 4 gnd
rlabel metal2 s 1008 1343 1008 1343 4 gnd
rlabel metal2 s 240 2370 240 2370 4 gnd
rlabel metal2 s 240 4977 240 4977 4 gnd
rlabel metal2 s 1008 6320 1008 6320 4 gnd
rlabel metal2 s 1008 2923 1008 2923 4 gnd
rlabel metal2 s 240 3950 240 3950 4 gnd
rlabel metal2 s 1008 0 1008 0 4 gnd
rlabel metal2 s 240 2607 240 2607 4 gnd
rlabel metal2 s 1008 5293 1008 5293 4 gnd
rlabel metal2 s 240 5530 240 5530 4 gnd
rlabel metal2 s 240 790 240 790 4 gnd
rlabel metal2 s 240 6083 240 6083 4 gnd
rlabel metal2 s 1008 4977 1008 4977 4 gnd
rlabel metal2 s 1008 2370 1008 2370 4 gnd
rlabel metal2 s 1008 3160 1008 3160 4 gnd
rlabel metal2 s 1008 4503 1008 4503 4 gnd
rlabel metal2 s 240 1580 240 1580 4 gnd
rlabel metal2 s 1008 553 1008 553 4 gnd
rlabel metal2 s 240 5293 240 5293 4 gnd
rlabel metal2 s 240 1817 240 1817 4 gnd
rlabel metal2 s 1008 2133 1008 2133 4 gnd
rlabel metal2 s 1008 790 1008 790 4 gnd
rlabel metal2 s 1008 2607 1008 2607 4 gnd
rlabel metal2 s 1008 4187 1008 4187 4 gnd
rlabel metal2 s 240 4503 240 4503 4 gnd
rlabel metal2 s 1008 3713 1008 3713 4 gnd
rlabel metal2 s 624 3507 624 3507 4 wl0_8
rlabel metal2 s 624 2497 624 2497 4 wl1_6
rlabel metal2 s 624 2717 624 2717 4 wl0_6
rlabel metal2 s 624 127 624 127 4 wl1_0
rlabel metal2 s 624 2813 624 2813 4 wl0_7
rlabel metal1 s 1008 2120 1008 2120 4 vdd
rlabel metal1 s 1008 3409 1008 3409 4 vdd
rlabel metal1 s 240 4199 240 4199 4 vdd
rlabel metal1 s 240 1829 240 1829 4 vdd
rlabel metal1 s 1008 4989 1008 4989 4 vdd
rlabel metal1 s 1008 5280 1008 5280 4 vdd
rlabel metal1 s 1008 249 1008 249 4 vdd
rlabel metal1 s 1008 1039 1008 1039 4 vdd
rlabel metal1 s 240 1039 240 1039 4 vdd
rlabel metal1 s 240 2120 240 2120 4 vdd
rlabel metal1 s 240 4989 240 4989 4 vdd
rlabel metal1 s 1008 5779 1008 5779 4 vdd
rlabel metal1 s 240 3409 240 3409 4 vdd
rlabel metal1 s 1008 3700 1008 3700 4 vdd
rlabel metal1 s 240 6070 240 6070 4 vdd
rlabel metal1 s 240 4490 240 4490 4 vdd
rlabel metal1 s 1008 1330 1008 1330 4 vdd
rlabel metal1 s 1008 2910 1008 2910 4 vdd
rlabel metal1 s 240 2619 240 2619 4 vdd
rlabel metal1 s 1008 2619 1008 2619 4 vdd
rlabel metal1 s 240 249 240 249 4 vdd
rlabel metal1 s 240 2910 240 2910 4 vdd
rlabel metal1 s 240 5280 240 5280 4 vdd
rlabel metal1 s 240 3700 240 3700 4 vdd
rlabel metal1 s 240 540 240 540 4 vdd
rlabel metal1 s 1008 1829 1008 1829 4 vdd
rlabel metal1 s 1008 6070 1008 6070 4 vdd
rlabel metal1 s 240 1330 240 1330 4 vdd
rlabel metal1 s 240 5779 240 5779 4 vdd
rlabel metal1 s 1008 540 1008 540 4 vdd
rlabel metal1 s 1008 4490 1008 4490 4 vdd
rlabel metal1 s 1008 4199 1008 4199 4 vdd
rlabel metal2 s 624 5973 624 5973 4 wl0_15
rlabel metal2 s 624 3287 624 3287 4 wl1_8
rlabel metal2 s 624 5087 624 5087 4 wl0_12
rlabel metal2 s 624 4867 624 4867 4 wl1_12
rlabel metal2 s 624 5877 624 5877 4 wl0_14
rlabel metal2 s 624 3603 624 3603 4 wl0_9
rlabel metal2 s 624 2243 624 2243 4 wl1_5
rlabel metal1 s 96 3160 96 3160 4 bl0_0
rlabel metal2 s 624 2023 624 2023 4 wl0_5
rlabel metal2 s 624 5183 624 5183 4 wl0_13
rlabel metal2 s 624 443 624 443 4 wl0_1
rlabel metal2 s 624 1453 624 1453 4 wl1_3
rlabel metal1 s 1152 3160 1152 3160 4 bl0_1
rlabel metal2 s 624 4297 624 4297 4 wl0_10
rlabel metal1 s 312 3160 312 3160 4 bl1_0
<< properties >>
string FIXED_BBOX 0 0 1248 6320
<< end >>
