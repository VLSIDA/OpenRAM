VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 1000 ;
END UNITS
SITE  MacroSite
   CLASS Core ;
   SIZE 277800.0 by 440700.0 ;
END  MacroSite
MACRO sram_2_16_1_scn3me_subm
   CLASS BLOCK ;
   SIZE 277800.0 BY 440700.0 ;
   SYMMETRY X Y R90 ;
   SITE MacroSite ;
   PIN DATA[0]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  180000.0 0.0 180900.0 1800.0 ;
      END
   END DATA[0]
   PIN DATA[1]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  190200.0 0.0 191100.0 1800.0 ;
      END
   END DATA[1]
   PIN ADDR[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  52800.0 77700.0 60000.0 79200.0 ;
      END
   END ADDR[0]
   PIN ADDR[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  52800.0 67500.0 60000.0 69000.0 ;
      END
   END ADDR[1]
   PIN ADDR[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  52800.0 57300.0 60000.0 58800.0 ;
      END
   END ADDR[2]
   PIN ADDR[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  52800.0 47100.0 60000.0 48600.0 ;
      END
   END ADDR[3]
   PIN CSb
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  14400.0 203400.0 16200.0 205200.0 ;
      END
   END CSb
   PIN WEb
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  24600.0 203400.0 26400.0 205200.0 ;
      END
   END WEb
   PIN OEb
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  4200.0 203400.0 6000.0 205200.0 ;
      END
   END OEb
   PIN clk
      DIRECTION INPUT ;
      PORT
         LAYER metal1 ;
         RECT  42600.0 202500.0 43800.0 206100.0 ;
      END
   END clk
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal1 ;
         RECT  198600.0 0.0 203100.0 440700.0 ;
         LAYER metal1 ;
         RECT  52800.0 0.0 57300.0 440700.0 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal2 ;
         RECT  148050.0 0.0 152550.0 440700.0 ;
      END
   END gnd
   OBS
   LAYER  metal1 ;
      RECT  54600.0 295950.0 55500.0 298650.0 ;
      RECT  97500.0 205650.0 98400.0 206550.0 ;
      RECT  97500.0 203250.0 98400.0 204150.0 ;
      RECT  96150.0 205650.0 97950.0 206550.0 ;
      RECT  97500.0 203700.0 98400.0 206100.0 ;
      RECT  97950.0 203250.0 99900.0 204150.0 ;
      RECT  154950.0 205650.0 155850.0 206550.0 ;
      RECT  154950.0 201150.0 155850.0 202050.0 ;
      RECT  136050.0 205650.0 155400.0 206550.0 ;
      RECT  154950.0 201600.0 155850.0 206100.0 ;
      RECT  155400.0 201150.0 174900.0 202050.0 ;
      RECT  97500.0 220050.0 98400.0 220950.0 ;
      RECT  97500.0 222450.0 98400.0 223350.0 ;
      RECT  96150.0 220050.0 97950.0 220950.0 ;
      RECT  97500.0 220500.0 98400.0 222900.0 ;
      RECT  97950.0 222450.0 99900.0 223350.0 ;
      RECT  154950.0 220050.0 155850.0 220950.0 ;
      RECT  154950.0 224550.0 155850.0 225450.0 ;
      RECT  136050.0 220050.0 155400.0 220950.0 ;
      RECT  154950.0 220500.0 155850.0 225000.0 ;
      RECT  155400.0 224550.0 174900.0 225450.0 ;
      RECT  97500.0 233250.0 98400.0 234150.0 ;
      RECT  97500.0 230850.0 98400.0 231750.0 ;
      RECT  96150.0 233250.0 97950.0 234150.0 ;
      RECT  97500.0 231300.0 98400.0 233700.0 ;
      RECT  97950.0 230850.0 99900.0 231750.0 ;
      RECT  154950.0 233250.0 155850.0 234150.0 ;
      RECT  154950.0 228750.0 155850.0 229650.0 ;
      RECT  136050.0 233250.0 155400.0 234150.0 ;
      RECT  154950.0 229200.0 155850.0 233700.0 ;
      RECT  155400.0 228750.0 174900.0 229650.0 ;
      RECT  97500.0 247650.0 98400.0 248550.0 ;
      RECT  97500.0 250050.0 98400.0 250950.0 ;
      RECT  96150.0 247650.0 97950.0 248550.0 ;
      RECT  97500.0 248100.0 98400.0 250500.0 ;
      RECT  97950.0 250050.0 99900.0 250950.0 ;
      RECT  154950.0 247650.0 155850.0 248550.0 ;
      RECT  154950.0 252150.0 155850.0 253050.0 ;
      RECT  136050.0 247650.0 155400.0 248550.0 ;
      RECT  154950.0 248100.0 155850.0 252600.0 ;
      RECT  155400.0 252150.0 174900.0 253050.0 ;
      RECT  97500.0 260850.0 98400.0 261750.0 ;
      RECT  97500.0 258450.0 98400.0 259350.0 ;
      RECT  96150.0 260850.0 97950.0 261750.0 ;
      RECT  97500.0 258900.0 98400.0 261300.0 ;
      RECT  97950.0 258450.0 99900.0 259350.0 ;
      RECT  154950.0 260850.0 155850.0 261750.0 ;
      RECT  154950.0 256350.0 155850.0 257250.0 ;
      RECT  136050.0 260850.0 155400.0 261750.0 ;
      RECT  154950.0 256800.0 155850.0 261300.0 ;
      RECT  155400.0 256350.0 174900.0 257250.0 ;
      RECT  97500.0 275250.0 98400.0 276150.0 ;
      RECT  97500.0 277650.0 98400.0 278550.0 ;
      RECT  96150.0 275250.0 97950.0 276150.0 ;
      RECT  97500.0 275700.0 98400.0 278100.0 ;
      RECT  97950.0 277650.0 99900.0 278550.0 ;
      RECT  154950.0 275250.0 155850.0 276150.0 ;
      RECT  154950.0 279750.0 155850.0 280650.0 ;
      RECT  136050.0 275250.0 155400.0 276150.0 ;
      RECT  154950.0 275700.0 155850.0 280200.0 ;
      RECT  155400.0 279750.0 174900.0 280650.0 ;
      RECT  97500.0 288450.0 98400.0 289350.0 ;
      RECT  97500.0 286050.0 98400.0 286950.0 ;
      RECT  96150.0 288450.0 97950.0 289350.0 ;
      RECT  97500.0 286500.0 98400.0 288900.0 ;
      RECT  97950.0 286050.0 99900.0 286950.0 ;
      RECT  154950.0 288450.0 155850.0 289350.0 ;
      RECT  154950.0 283950.0 155850.0 284850.0 ;
      RECT  136050.0 288450.0 155400.0 289350.0 ;
      RECT  154950.0 284400.0 155850.0 288900.0 ;
      RECT  155400.0 283950.0 174900.0 284850.0 ;
      RECT  97500.0 302850.0 98400.0 303750.0 ;
      RECT  97500.0 305250.0 98400.0 306150.0 ;
      RECT  96150.0 302850.0 97950.0 303750.0 ;
      RECT  97500.0 303300.0 98400.0 305700.0 ;
      RECT  97950.0 305250.0 99900.0 306150.0 ;
      RECT  154950.0 302850.0 155850.0 303750.0 ;
      RECT  154950.0 307350.0 155850.0 308250.0 ;
      RECT  136050.0 302850.0 155400.0 303750.0 ;
      RECT  154950.0 303300.0 155850.0 307800.0 ;
      RECT  155400.0 307350.0 174900.0 308250.0 ;
      RECT  97500.0 316050.0 98400.0 316950.0 ;
      RECT  97500.0 313650.0 98400.0 314550.0 ;
      RECT  96150.0 316050.0 97950.0 316950.0 ;
      RECT  97500.0 314100.0 98400.0 316500.0 ;
      RECT  97950.0 313650.0 99900.0 314550.0 ;
      RECT  154950.0 316050.0 155850.0 316950.0 ;
      RECT  154950.0 311550.0 155850.0 312450.0 ;
      RECT  136050.0 316050.0 155400.0 316950.0 ;
      RECT  154950.0 312000.0 155850.0 316500.0 ;
      RECT  155400.0 311550.0 174900.0 312450.0 ;
      RECT  97500.0 330450.0 98400.0 331350.0 ;
      RECT  97500.0 332850.0 98400.0 333750.0 ;
      RECT  96150.0 330450.0 97950.0 331350.0 ;
      RECT  97500.0 330900.0 98400.0 333300.0 ;
      RECT  97950.0 332850.0 99900.0 333750.0 ;
      RECT  154950.0 330450.0 155850.0 331350.0 ;
      RECT  154950.0 334950.0 155850.0 335850.0 ;
      RECT  136050.0 330450.0 155400.0 331350.0 ;
      RECT  154950.0 330900.0 155850.0 335400.0 ;
      RECT  155400.0 334950.0 174900.0 335850.0 ;
      RECT  97500.0 343650.0 98400.0 344550.0 ;
      RECT  97500.0 341250.0 98400.0 342150.0 ;
      RECT  96150.0 343650.0 97950.0 344550.0 ;
      RECT  97500.0 341700.0 98400.0 344100.0 ;
      RECT  97950.0 341250.0 99900.0 342150.0 ;
      RECT  154950.0 343650.0 155850.0 344550.0 ;
      RECT  154950.0 339150.0 155850.0 340050.0 ;
      RECT  136050.0 343650.0 155400.0 344550.0 ;
      RECT  154950.0 339600.0 155850.0 344100.0 ;
      RECT  155400.0 339150.0 174900.0 340050.0 ;
      RECT  97500.0 358050.0 98400.0 358950.0 ;
      RECT  97500.0 360450.0 98400.0 361350.0 ;
      RECT  96150.0 358050.0 97950.0 358950.0 ;
      RECT  97500.0 358500.0 98400.0 360900.0 ;
      RECT  97950.0 360450.0 99900.0 361350.0 ;
      RECT  154950.0 358050.0 155850.0 358950.0 ;
      RECT  154950.0 362550.0 155850.0 363450.0 ;
      RECT  136050.0 358050.0 155400.0 358950.0 ;
      RECT  154950.0 358500.0 155850.0 363000.0 ;
      RECT  155400.0 362550.0 174900.0 363450.0 ;
      RECT  97500.0 371250.0 98400.0 372150.0 ;
      RECT  97500.0 368850.0 98400.0 369750.0 ;
      RECT  96150.0 371250.0 97950.0 372150.0 ;
      RECT  97500.0 369300.0 98400.0 371700.0 ;
      RECT  97950.0 368850.0 99900.0 369750.0 ;
      RECT  154950.0 371250.0 155850.0 372150.0 ;
      RECT  154950.0 366750.0 155850.0 367650.0 ;
      RECT  136050.0 371250.0 155400.0 372150.0 ;
      RECT  154950.0 367200.0 155850.0 371700.0 ;
      RECT  155400.0 366750.0 174900.0 367650.0 ;
      RECT  97500.0 385650.0 98400.0 386550.0 ;
      RECT  97500.0 388050.0 98400.0 388950.0 ;
      RECT  96150.0 385650.0 97950.0 386550.0 ;
      RECT  97500.0 386100.0 98400.0 388500.0 ;
      RECT  97950.0 388050.0 99900.0 388950.0 ;
      RECT  154950.0 385650.0 155850.0 386550.0 ;
      RECT  154950.0 390150.0 155850.0 391050.0 ;
      RECT  136050.0 385650.0 155400.0 386550.0 ;
      RECT  154950.0 386100.0 155850.0 390600.0 ;
      RECT  155400.0 390150.0 174900.0 391050.0 ;
      RECT  97500.0 398850.0 98400.0 399750.0 ;
      RECT  97500.0 396450.0 98400.0 397350.0 ;
      RECT  96150.0 398850.0 97950.0 399750.0 ;
      RECT  97500.0 396900.0 98400.0 399300.0 ;
      RECT  97950.0 396450.0 99900.0 397350.0 ;
      RECT  154950.0 398850.0 155850.0 399750.0 ;
      RECT  154950.0 394350.0 155850.0 395250.0 ;
      RECT  136050.0 398850.0 155400.0 399750.0 ;
      RECT  154950.0 394800.0 155850.0 399300.0 ;
      RECT  155400.0 394350.0 174900.0 395250.0 ;
      RECT  97500.0 413250.0 98400.0 414150.0 ;
      RECT  97500.0 415650.0 98400.0 416550.0 ;
      RECT  96150.0 413250.0 97950.0 414150.0 ;
      RECT  97500.0 413700.0 98400.0 416100.0 ;
      RECT  97950.0 415650.0 99900.0 416550.0 ;
      RECT  154950.0 413250.0 155850.0 414150.0 ;
      RECT  154950.0 417750.0 155850.0 418650.0 ;
      RECT  136050.0 413250.0 155400.0 414150.0 ;
      RECT  154950.0 413700.0 155850.0 418200.0 ;
      RECT  155400.0 417750.0 174900.0 418650.0 ;
      RECT  106200.0 199050.0 175500.0 199950.0 ;
      RECT  106200.0 226650.0 175500.0 227550.0 ;
      RECT  106200.0 254250.0 175500.0 255150.0 ;
      RECT  106200.0 281850.0 175500.0 282750.0 ;
      RECT  106200.0 309450.0 175500.0 310350.0 ;
      RECT  106200.0 337050.0 175500.0 337950.0 ;
      RECT  106200.0 364650.0 175500.0 365550.0 ;
      RECT  106200.0 392250.0 175500.0 393150.0 ;
      RECT  106200.0 419850.0 175500.0 420750.0 ;
      RECT  52800.0 212850.0 203100.0 213750.0 ;
      RECT  52800.0 240450.0 203100.0 241350.0 ;
      RECT  52800.0 268050.0 203100.0 268950.0 ;
      RECT  52800.0 295650.0 203100.0 296550.0 ;
      RECT  52800.0 323250.0 203100.0 324150.0 ;
      RECT  52800.0 350850.0 203100.0 351750.0 ;
      RECT  52800.0 378450.0 203100.0 379350.0 ;
      RECT  52800.0 406050.0 203100.0 406950.0 ;
      RECT  130500.0 91350.0 135000.0 92250.0 ;
      RECT  127500.0 105150.0 137700.0 106050.0 ;
      RECT  130500.0 146550.0 140400.0 147450.0 ;
      RECT  127500.0 160350.0 143100.0 161250.0 ;
      RECT  130500.0 88650.0 132000.0 89550.0 ;
      RECT  130500.0 116250.0 132000.0 117150.0 ;
      RECT  130500.0 143850.0 132000.0 144750.0 ;
      RECT  130500.0 171450.0 132000.0 172350.0 ;
      RECT  52800.0 102450.0 130500.0 103350.0 ;
      RECT  52800.0 130050.0 130500.0 130950.0 ;
      RECT  52800.0 157650.0 130500.0 158550.0 ;
      RECT  52800.0 185250.0 130500.0 186150.0 ;
      RECT  117900.0 77400.0 135000.0 78300.0 ;
      RECT  117900.0 68700.0 137700.0 69600.0 ;
      RECT  117900.0 57000.0 140400.0 57900.0 ;
      RECT  117900.0 48300.0 143100.0 49200.0 ;
      RECT  119100.0 73050.0 149250.0 73950.0 ;
      RECT  119100.0 52650.0 149250.0 53550.0 ;
      RECT  115500.0 40350.0 116400.0 41250.0 ;
      RECT  115500.0 40800.0 116400.0 42900.0 ;
      RECT  52800.0 40350.0 115950.0 41250.0 ;
      RECT  163800.0 32400.0 175500.0 33300.0 ;
      RECT  158400.0 27900.0 175500.0 28800.0 ;
      RECT  161100.0 25500.0 175500.0 26400.0 ;
      RECT  163800.0 428700.0 175500.0 429600.0 ;
      RECT  166500.0 97200.0 175500.0 98100.0 ;
      RECT  169200.0 195300.0 175500.0 196200.0 ;
      RECT  61500.0 85350.0 62400.0 86250.0 ;
      RECT  61500.0 83700.0 62400.0 85800.0 ;
      RECT  61950.0 85350.0 155700.0 86250.0 ;
      RECT  103050.0 421950.0 156600.0 422850.0 ;
      RECT  175500.0 439800.0 198600.0 440700.0 ;
      RECT  175500.0 168000.0 198600.0 168900.0 ;
      RECT  175500.0 99300.0 198600.0 100200.0 ;
      RECT  175500.0 86400.0 198600.0 87300.0 ;
      RECT  175500.0 9600.0 198600.0 10500.0 ;
      RECT  152550.0 23400.0 175500.0 24300.0 ;
      RECT  152550.0 193200.0 175500.0 194100.0 ;
      RECT  152550.0 95100.0 175500.0 96000.0 ;
      RECT  175500.0 199500.0 185700.0 213300.0 ;
      RECT  175500.0 227100.0 185700.0 213300.0 ;
      RECT  175500.0 227100.0 185700.0 240900.0 ;
      RECT  175500.0 254700.0 185700.0 240900.0 ;
      RECT  175500.0 254700.0 185700.0 268500.0 ;
      RECT  175500.0 282300.0 185700.0 268500.0 ;
      RECT  175500.0 282300.0 185700.0 296100.0 ;
      RECT  175500.0 309900.0 185700.0 296100.0 ;
      RECT  175500.0 309900.0 185700.0 323700.0 ;
      RECT  175500.0 337500.0 185700.0 323700.0 ;
      RECT  175500.0 337500.0 185700.0 351300.0 ;
      RECT  175500.0 365100.0 185700.0 351300.0 ;
      RECT  175500.0 365100.0 185700.0 378900.0 ;
      RECT  175500.0 392700.0 185700.0 378900.0 ;
      RECT  175500.0 392700.0 185700.0 406500.0 ;
      RECT  175500.0 420300.0 185700.0 406500.0 ;
      RECT  185700.0 199500.0 195900.0 213300.0 ;
      RECT  185700.0 227100.0 195900.0 213300.0 ;
      RECT  185700.0 227100.0 195900.0 240900.0 ;
      RECT  185700.0 254700.0 195900.0 240900.0 ;
      RECT  185700.0 254700.0 195900.0 268500.0 ;
      RECT  185700.0 282300.0 195900.0 268500.0 ;
      RECT  185700.0 282300.0 195900.0 296100.0 ;
      RECT  185700.0 309900.0 195900.0 296100.0 ;
      RECT  185700.0 309900.0 195900.0 323700.0 ;
      RECT  185700.0 337500.0 195900.0 323700.0 ;
      RECT  185700.0 337500.0 195900.0 351300.0 ;
      RECT  185700.0 365100.0 195900.0 351300.0 ;
      RECT  185700.0 365100.0 195900.0 378900.0 ;
      RECT  185700.0 392700.0 195900.0 378900.0 ;
      RECT  185700.0 392700.0 195900.0 406500.0 ;
      RECT  185700.0 420300.0 195900.0 406500.0 ;
      RECT  174900.0 201000.0 196500.0 202200.0 ;
      RECT  174900.0 224400.0 196500.0 225600.0 ;
      RECT  174900.0 228600.0 196500.0 229800.0 ;
      RECT  174900.0 252000.0 196500.0 253200.0 ;
      RECT  174900.0 256200.0 196500.0 257400.0 ;
      RECT  174900.0 279600.0 196500.0 280800.0 ;
      RECT  174900.0 283800.0 196500.0 285000.0 ;
      RECT  174900.0 307200.0 196500.0 308400.0 ;
      RECT  174900.0 311400.0 196500.0 312600.0 ;
      RECT  174900.0 334800.0 196500.0 336000.0 ;
      RECT  174900.0 339000.0 196500.0 340200.0 ;
      RECT  174900.0 362400.0 196500.0 363600.0 ;
      RECT  174900.0 366600.0 196500.0 367800.0 ;
      RECT  174900.0 390000.0 196500.0 391200.0 ;
      RECT  174900.0 394200.0 196500.0 395400.0 ;
      RECT  174900.0 417600.0 196500.0 418800.0 ;
      RECT  174900.0 212700.0 196500.0 213600.0 ;
      RECT  174900.0 240300.0 196500.0 241200.0 ;
      RECT  174900.0 267900.0 196500.0 268800.0 ;
      RECT  174900.0 295500.0 196500.0 296400.0 ;
      RECT  174900.0 323100.0 196500.0 324000.0 ;
      RECT  174900.0 350700.0 196500.0 351600.0 ;
      RECT  174900.0 378300.0 196500.0 379200.0 ;
      RECT  174900.0 405900.0 196500.0 406800.0 ;
      RECT  180900.0 433500.0 182100.0 440700.0 ;
      RECT  178500.0 426300.0 179700.0 427500.0 ;
      RECT  180900.0 426300.0 182100.0 427500.0 ;
      RECT  180900.0 426300.0 182100.0 427500.0 ;
      RECT  178500.0 426300.0 179700.0 427500.0 ;
      RECT  178500.0 433500.0 179700.0 434700.0 ;
      RECT  180900.0 433500.0 182100.0 434700.0 ;
      RECT  180900.0 433500.0 182100.0 434700.0 ;
      RECT  178500.0 433500.0 179700.0 434700.0 ;
      RECT  180900.0 433500.0 182100.0 434700.0 ;
      RECT  183300.0 433500.0 184500.0 434700.0 ;
      RECT  183300.0 433500.0 184500.0 434700.0 ;
      RECT  180900.0 433500.0 182100.0 434700.0 ;
      RECT  180600.0 428550.0 179400.0 429750.0 ;
      RECT  180900.0 438900.0 182100.0 440100.0 ;
      RECT  178500.0 426300.0 179700.0 427500.0 ;
      RECT  180900.0 426300.0 182100.0 427500.0 ;
      RECT  178500.0 433500.0 179700.0 434700.0 ;
      RECT  183300.0 433500.0 184500.0 434700.0 ;
      RECT  175500.0 428700.0 185700.0 429600.0 ;
      RECT  175500.0 439800.0 185700.0 440700.0 ;
      RECT  191100.0 433500.0 192300.0 440700.0 ;
      RECT  188700.0 426300.0 189900.0 427500.0 ;
      RECT  191100.0 426300.0 192300.0 427500.0 ;
      RECT  191100.0 426300.0 192300.0 427500.0 ;
      RECT  188700.0 426300.0 189900.0 427500.0 ;
      RECT  188700.0 433500.0 189900.0 434700.0 ;
      RECT  191100.0 433500.0 192300.0 434700.0 ;
      RECT  191100.0 433500.0 192300.0 434700.0 ;
      RECT  188700.0 433500.0 189900.0 434700.0 ;
      RECT  191100.0 433500.0 192300.0 434700.0 ;
      RECT  193500.0 433500.0 194700.0 434700.0 ;
      RECT  193500.0 433500.0 194700.0 434700.0 ;
      RECT  191100.0 433500.0 192300.0 434700.0 ;
      RECT  190800.0 428550.0 189600.0 429750.0 ;
      RECT  191100.0 438900.0 192300.0 440100.0 ;
      RECT  188700.0 426300.0 189900.0 427500.0 ;
      RECT  191100.0 426300.0 192300.0 427500.0 ;
      RECT  188700.0 433500.0 189900.0 434700.0 ;
      RECT  193500.0 433500.0 194700.0 434700.0 ;
      RECT  185700.0 428700.0 195900.0 429600.0 ;
      RECT  185700.0 439800.0 195900.0 440700.0 ;
      RECT  175500.0 428700.0 195900.0 429600.0 ;
      RECT  175500.0 439800.0 195900.0 440700.0 ;
      RECT  175500.0 150600.0 185700.0 199500.0 ;
      RECT  185700.0 150600.0 195900.0 199500.0 ;
      RECT  175500.0 195300.0 195900.0 196200.0 ;
      RECT  175500.0 168000.0 195900.0 168900.0 ;
      RECT  175500.0 193200.0 195900.0 194100.0 ;
      RECT  175500.0 90000.0 185700.0 150600.0 ;
      RECT  185700.0 90000.0 195900.0 150600.0 ;
      RECT  175500.0 97200.0 195900.0 98100.0 ;
      RECT  175500.0 99300.0 195900.0 100200.0 ;
      RECT  175500.0 95100.0 195900.0 96000.0 ;
      RECT  175500.0 30000.0 185700.0 90000.0 ;
      RECT  195900.0 30000.0 185700.0 90000.0 ;
      RECT  175500.0 32400.0 195900.0 33300.0 ;
      RECT  175500.0 86400.0 195900.0 87300.0 ;
      RECT  175500.0 30000.0 185700.0 8100.0 ;
      RECT  185700.0 30000.0 195900.0 8100.0 ;
      RECT  175500.0 26400.0 195900.0 25500.0 ;
      RECT  175500.0 28800.0 195900.0 27900.0 ;
      RECT  175500.0 10500.0 195900.0 9600.0 ;
      RECT  175500.0 24300.0 195900.0 23400.0 ;
      RECT  87750.0 206850.0 88650.0 207750.0 ;
      RECT  87750.0 205650.0 88650.0 206550.0 ;
      RECT  83700.0 206850.0 88200.0 207750.0 ;
      RECT  87750.0 206100.0 88650.0 207300.0 ;
      RECT  88200.0 205650.0 92700.0 206550.0 ;
      RECT  87750.0 218850.0 88650.0 219750.0 ;
      RECT  87750.0 220050.0 88650.0 220950.0 ;
      RECT  83700.0 218850.0 88200.0 219750.0 ;
      RECT  87750.0 219300.0 88650.0 220500.0 ;
      RECT  88200.0 220050.0 92700.0 220950.0 ;
      RECT  87750.0 234450.0 88650.0 235350.0 ;
      RECT  87750.0 233250.0 88650.0 234150.0 ;
      RECT  83700.0 234450.0 88200.0 235350.0 ;
      RECT  87750.0 233700.0 88650.0 234900.0 ;
      RECT  88200.0 233250.0 92700.0 234150.0 ;
      RECT  87750.0 246450.0 88650.0 247350.0 ;
      RECT  87750.0 247650.0 88650.0 248550.0 ;
      RECT  83700.0 246450.0 88200.0 247350.0 ;
      RECT  87750.0 246900.0 88650.0 248100.0 ;
      RECT  88200.0 247650.0 92700.0 248550.0 ;
      RECT  87750.0 262050.0 88650.0 262950.0 ;
      RECT  87750.0 260850.0 88650.0 261750.0 ;
      RECT  83700.0 262050.0 88200.0 262950.0 ;
      RECT  87750.0 261300.0 88650.0 262500.0 ;
      RECT  88200.0 260850.0 92700.0 261750.0 ;
      RECT  87750.0 274050.0 88650.0 274950.0 ;
      RECT  87750.0 275250.0 88650.0 276150.0 ;
      RECT  83700.0 274050.0 88200.0 274950.0 ;
      RECT  87750.0 274500.0 88650.0 275700.0 ;
      RECT  88200.0 275250.0 92700.0 276150.0 ;
      RECT  87750.0 289650.0 88650.0 290550.0 ;
      RECT  87750.0 288450.0 88650.0 289350.0 ;
      RECT  83700.0 289650.0 88200.0 290550.0 ;
      RECT  87750.0 288900.0 88650.0 290100.0 ;
      RECT  88200.0 288450.0 92700.0 289350.0 ;
      RECT  87750.0 301650.0 88650.0 302550.0 ;
      RECT  87750.0 302850.0 88650.0 303750.0 ;
      RECT  83700.0 301650.0 88200.0 302550.0 ;
      RECT  87750.0 302100.0 88650.0 303300.0 ;
      RECT  88200.0 302850.0 92700.0 303750.0 ;
      RECT  87750.0 317250.0 88650.0 318150.0 ;
      RECT  87750.0 316050.0 88650.0 316950.0 ;
      RECT  83700.0 317250.0 88200.0 318150.0 ;
      RECT  87750.0 316500.0 88650.0 317700.0 ;
      RECT  88200.0 316050.0 92700.0 316950.0 ;
      RECT  87750.0 329250.0 88650.0 330150.0 ;
      RECT  87750.0 330450.0 88650.0 331350.0 ;
      RECT  83700.0 329250.0 88200.0 330150.0 ;
      RECT  87750.0 329700.0 88650.0 330900.0 ;
      RECT  88200.0 330450.0 92700.0 331350.0 ;
      RECT  87750.0 344850.0 88650.0 345750.0 ;
      RECT  87750.0 343650.0 88650.0 344550.0 ;
      RECT  83700.0 344850.0 88200.0 345750.0 ;
      RECT  87750.0 344100.0 88650.0 345300.0 ;
      RECT  88200.0 343650.0 92700.0 344550.0 ;
      RECT  87750.0 356850.0 88650.0 357750.0 ;
      RECT  87750.0 358050.0 88650.0 358950.0 ;
      RECT  83700.0 356850.0 88200.0 357750.0 ;
      RECT  87750.0 357300.0 88650.0 358500.0 ;
      RECT  88200.0 358050.0 92700.0 358950.0 ;
      RECT  87750.0 372450.0 88650.0 373350.0 ;
      RECT  87750.0 371250.0 88650.0 372150.0 ;
      RECT  83700.0 372450.0 88200.0 373350.0 ;
      RECT  87750.0 371700.0 88650.0 372900.0 ;
      RECT  88200.0 371250.0 92700.0 372150.0 ;
      RECT  87750.0 384450.0 88650.0 385350.0 ;
      RECT  87750.0 385650.0 88650.0 386550.0 ;
      RECT  83700.0 384450.0 88200.0 385350.0 ;
      RECT  87750.0 384900.0 88650.0 386100.0 ;
      RECT  88200.0 385650.0 92700.0 386550.0 ;
      RECT  87750.0 400050.0 88650.0 400950.0 ;
      RECT  87750.0 398850.0 88650.0 399750.0 ;
      RECT  83700.0 400050.0 88200.0 400950.0 ;
      RECT  87750.0 399300.0 88650.0 400500.0 ;
      RECT  88200.0 398850.0 92700.0 399750.0 ;
      RECT  87750.0 412050.0 88650.0 412950.0 ;
      RECT  87750.0 413250.0 88650.0 414150.0 ;
      RECT  83700.0 412050.0 88200.0 412950.0 ;
      RECT  87750.0 412500.0 88650.0 413700.0 ;
      RECT  88200.0 413250.0 92700.0 414150.0 ;
      RECT  59550.0 95250.0 75900.0 96150.0 ;
      RECT  61650.0 109650.0 75900.0 110550.0 ;
      RECT  63750.0 122850.0 75900.0 123750.0 ;
      RECT  65850.0 137250.0 75900.0 138150.0 ;
      RECT  67950.0 150450.0 75900.0 151350.0 ;
      RECT  70050.0 164850.0 75900.0 165750.0 ;
      RECT  72150.0 178050.0 75900.0 178950.0 ;
      RECT  74250.0 192450.0 75900.0 193350.0 ;
      RECT  59550.0 206850.0 78300.0 207750.0 ;
      RECT  67950.0 204150.0 81300.0 205050.0 ;
      RECT  59550.0 218850.0 78300.0 219750.0 ;
      RECT  70050.0 221550.0 81300.0 222450.0 ;
      RECT  59550.0 234450.0 78300.0 235350.0 ;
      RECT  72150.0 231750.0 81300.0 232650.0 ;
      RECT  59550.0 246450.0 78300.0 247350.0 ;
      RECT  74250.0 249150.0 81300.0 250050.0 ;
      RECT  61650.0 262050.0 78300.0 262950.0 ;
      RECT  67950.0 259350.0 81300.0 260250.0 ;
      RECT  61650.0 274050.0 78300.0 274950.0 ;
      RECT  70050.0 276750.0 81300.0 277650.0 ;
      RECT  61650.0 289650.0 78300.0 290550.0 ;
      RECT  72150.0 286950.0 81300.0 287850.0 ;
      RECT  61650.0 301650.0 78300.0 302550.0 ;
      RECT  74250.0 304350.0 81300.0 305250.0 ;
      RECT  63750.0 317250.0 78300.0 318150.0 ;
      RECT  67950.0 314550.0 81300.0 315450.0 ;
      RECT  63750.0 329250.0 78300.0 330150.0 ;
      RECT  70050.0 331950.0 81300.0 332850.0 ;
      RECT  63750.0 344850.0 78300.0 345750.0 ;
      RECT  72150.0 342150.0 81300.0 343050.0 ;
      RECT  63750.0 356850.0 78300.0 357750.0 ;
      RECT  74250.0 359550.0 81300.0 360450.0 ;
      RECT  65850.0 372450.0 78300.0 373350.0 ;
      RECT  67950.0 369750.0 81300.0 370650.0 ;
      RECT  65850.0 384450.0 78300.0 385350.0 ;
      RECT  70050.0 387150.0 81300.0 388050.0 ;
      RECT  65850.0 400050.0 78300.0 400950.0 ;
      RECT  72150.0 397350.0 81300.0 398250.0 ;
      RECT  65850.0 412050.0 78300.0 412950.0 ;
      RECT  74250.0 414750.0 81300.0 415650.0 ;
      RECT  114450.0 95250.0 113550.0 96150.0 ;
      RECT  114450.0 99750.0 113550.0 100650.0 ;
      RECT  118650.0 95250.0 114000.0 96150.0 ;
      RECT  114450.0 95700.0 113550.0 100200.0 ;
      RECT  114000.0 99750.0 111450.0 100650.0 ;
      RECT  130050.0 95250.0 122100.0 96150.0 ;
      RECT  114450.0 109650.0 113550.0 110550.0 ;
      RECT  114450.0 113550.0 113550.0 114450.0 ;
      RECT  118650.0 109650.0 114000.0 110550.0 ;
      RECT  114450.0 110100.0 113550.0 114000.0 ;
      RECT  114000.0 113550.0 108450.0 114450.0 ;
      RECT  127050.0 109650.0 122100.0 110550.0 ;
      RECT  130050.0 118350.0 105450.0 119250.0 ;
      RECT  127050.0 132150.0 102450.0 133050.0 ;
      RECT  111450.0 96450.0 97500.0 97350.0 ;
      RECT  108450.0 93750.0 94500.0 94650.0 ;
      RECT  105450.0 108450.0 97500.0 109350.0 ;
      RECT  108450.0 111150.0 94500.0 112050.0 ;
      RECT  111450.0 124050.0 97500.0 124950.0 ;
      RECT  102450.0 121350.0 94500.0 122250.0 ;
      RECT  105450.0 136050.0 97500.0 136950.0 ;
      RECT  102450.0 138750.0 94500.0 139650.0 ;
      RECT  88050.0 96450.0 87150.0 97350.0 ;
      RECT  88050.0 95250.0 87150.0 96150.0 ;
      RECT  92100.0 96450.0 87600.0 97350.0 ;
      RECT  88050.0 95700.0 87150.0 96900.0 ;
      RECT  87600.0 95250.0 83100.0 96150.0 ;
      RECT  88050.0 108450.0 87150.0 109350.0 ;
      RECT  88050.0 109650.0 87150.0 110550.0 ;
      RECT  92100.0 108450.0 87600.0 109350.0 ;
      RECT  88050.0 108900.0 87150.0 110100.0 ;
      RECT  87600.0 109650.0 83100.0 110550.0 ;
      RECT  88050.0 124050.0 87150.0 124950.0 ;
      RECT  88050.0 122850.0 87150.0 123750.0 ;
      RECT  92100.0 124050.0 87600.0 124950.0 ;
      RECT  88050.0 123300.0 87150.0 124500.0 ;
      RECT  87600.0 122850.0 83100.0 123750.0 ;
      RECT  88050.0 136050.0 87150.0 136950.0 ;
      RECT  88050.0 137250.0 87150.0 138150.0 ;
      RECT  92100.0 136050.0 87600.0 136950.0 ;
      RECT  88050.0 136500.0 87150.0 137700.0 ;
      RECT  87600.0 137250.0 83100.0 138150.0 ;
      RECT  117900.0 100950.0 116700.0 102900.0 ;
      RECT  117900.0 89100.0 116700.0 91050.0 ;
      RECT  122700.0 90450.0 121500.0 88650.0 ;
      RECT  122700.0 99750.0 121500.0 103350.0 ;
      RECT  120000.0 90450.0 119100.0 99750.0 ;
      RECT  122700.0 99750.0 121500.0 100950.0 ;
      RECT  120300.0 99750.0 119100.0 100950.0 ;
      RECT  120300.0 99750.0 119100.0 100950.0 ;
      RECT  122700.0 99750.0 121500.0 100950.0 ;
      RECT  122700.0 90450.0 121500.0 91650.0 ;
      RECT  120300.0 90450.0 119100.0 91650.0 ;
      RECT  120300.0 90450.0 119100.0 91650.0 ;
      RECT  122700.0 90450.0 121500.0 91650.0 ;
      RECT  117900.0 100350.0 116700.0 101550.0 ;
      RECT  117900.0 90450.0 116700.0 91650.0 ;
      RECT  122100.0 95100.0 120900.0 96300.0 ;
      RECT  122100.0 95100.0 120900.0 96300.0 ;
      RECT  119550.0 95250.0 118650.0 96150.0 ;
      RECT  124500.0 102450.0 114900.0 103350.0 ;
      RECT  124500.0 88650.0 114900.0 89550.0 ;
      RECT  117900.0 104850.0 116700.0 102900.0 ;
      RECT  117900.0 116700.0 116700.0 114750.0 ;
      RECT  122700.0 115350.0 121500.0 117150.0 ;
      RECT  122700.0 106050.0 121500.0 102450.0 ;
      RECT  120000.0 115350.0 119100.0 106050.0 ;
      RECT  122700.0 106050.0 121500.0 104850.0 ;
      RECT  120300.0 106050.0 119100.0 104850.0 ;
      RECT  120300.0 106050.0 119100.0 104850.0 ;
      RECT  122700.0 106050.0 121500.0 104850.0 ;
      RECT  122700.0 115350.0 121500.0 114150.0 ;
      RECT  120300.0 115350.0 119100.0 114150.0 ;
      RECT  120300.0 115350.0 119100.0 114150.0 ;
      RECT  122700.0 115350.0 121500.0 114150.0 ;
      RECT  117900.0 105450.0 116700.0 104250.0 ;
      RECT  117900.0 115350.0 116700.0 114150.0 ;
      RECT  122100.0 110700.0 120900.0 109500.0 ;
      RECT  122100.0 110700.0 120900.0 109500.0 ;
      RECT  119550.0 110550.0 118650.0 109650.0 ;
      RECT  124500.0 103350.0 114900.0 102450.0 ;
      RECT  124500.0 117150.0 114900.0 116250.0 ;
      RECT  78900.0 100950.0 77700.0 102900.0 ;
      RECT  78900.0 89100.0 77700.0 91050.0 ;
      RECT  83700.0 90450.0 82500.0 88650.0 ;
      RECT  83700.0 99750.0 82500.0 103350.0 ;
      RECT  81000.0 90450.0 80100.0 99750.0 ;
      RECT  83700.0 99750.0 82500.0 100950.0 ;
      RECT  81300.0 99750.0 80100.0 100950.0 ;
      RECT  81300.0 99750.0 80100.0 100950.0 ;
      RECT  83700.0 99750.0 82500.0 100950.0 ;
      RECT  83700.0 90450.0 82500.0 91650.0 ;
      RECT  81300.0 90450.0 80100.0 91650.0 ;
      RECT  81300.0 90450.0 80100.0 91650.0 ;
      RECT  83700.0 90450.0 82500.0 91650.0 ;
      RECT  78900.0 100350.0 77700.0 101550.0 ;
      RECT  78900.0 90450.0 77700.0 91650.0 ;
      RECT  83100.0 95100.0 81900.0 96300.0 ;
      RECT  83100.0 95100.0 81900.0 96300.0 ;
      RECT  80550.0 95250.0 79650.0 96150.0 ;
      RECT  85500.0 102450.0 75900.0 103350.0 ;
      RECT  85500.0 88650.0 75900.0 89550.0 ;
      RECT  78900.0 104850.0 77700.0 102900.0 ;
      RECT  78900.0 116700.0 77700.0 114750.0 ;
      RECT  83700.0 115350.0 82500.0 117150.0 ;
      RECT  83700.0 106050.0 82500.0 102450.0 ;
      RECT  81000.0 115350.0 80100.0 106050.0 ;
      RECT  83700.0 106050.0 82500.0 104850.0 ;
      RECT  81300.0 106050.0 80100.0 104850.0 ;
      RECT  81300.0 106050.0 80100.0 104850.0 ;
      RECT  83700.0 106050.0 82500.0 104850.0 ;
      RECT  83700.0 115350.0 82500.0 114150.0 ;
      RECT  81300.0 115350.0 80100.0 114150.0 ;
      RECT  81300.0 115350.0 80100.0 114150.0 ;
      RECT  83700.0 115350.0 82500.0 114150.0 ;
      RECT  78900.0 105450.0 77700.0 104250.0 ;
      RECT  78900.0 115350.0 77700.0 114150.0 ;
      RECT  83100.0 110700.0 81900.0 109500.0 ;
      RECT  83100.0 110700.0 81900.0 109500.0 ;
      RECT  80550.0 110550.0 79650.0 109650.0 ;
      RECT  85500.0 103350.0 75900.0 102450.0 ;
      RECT  85500.0 117150.0 75900.0 116250.0 ;
      RECT  78900.0 128550.0 77700.0 130500.0 ;
      RECT  78900.0 116700.0 77700.0 118650.0 ;
      RECT  83700.0 118050.0 82500.0 116250.0 ;
      RECT  83700.0 127350.0 82500.0 130950.0 ;
      RECT  81000.0 118050.0 80100.0 127350.0 ;
      RECT  83700.0 127350.0 82500.0 128550.0 ;
      RECT  81300.0 127350.0 80100.0 128550.0 ;
      RECT  81300.0 127350.0 80100.0 128550.0 ;
      RECT  83700.0 127350.0 82500.0 128550.0 ;
      RECT  83700.0 118050.0 82500.0 119250.0 ;
      RECT  81300.0 118050.0 80100.0 119250.0 ;
      RECT  81300.0 118050.0 80100.0 119250.0 ;
      RECT  83700.0 118050.0 82500.0 119250.0 ;
      RECT  78900.0 127950.0 77700.0 129150.0 ;
      RECT  78900.0 118050.0 77700.0 119250.0 ;
      RECT  83100.0 122700.0 81900.0 123900.0 ;
      RECT  83100.0 122700.0 81900.0 123900.0 ;
      RECT  80550.0 122850.0 79650.0 123750.0 ;
      RECT  85500.0 130050.0 75900.0 130950.0 ;
      RECT  85500.0 116250.0 75900.0 117150.0 ;
      RECT  78900.0 132450.0 77700.0 130500.0 ;
      RECT  78900.0 144300.0 77700.0 142350.0 ;
      RECT  83700.0 142950.0 82500.0 144750.0 ;
      RECT  83700.0 133650.0 82500.0 130050.0 ;
      RECT  81000.0 142950.0 80100.0 133650.0 ;
      RECT  83700.0 133650.0 82500.0 132450.0 ;
      RECT  81300.0 133650.0 80100.0 132450.0 ;
      RECT  81300.0 133650.0 80100.0 132450.0 ;
      RECT  83700.0 133650.0 82500.0 132450.0 ;
      RECT  83700.0 142950.0 82500.0 141750.0 ;
      RECT  81300.0 142950.0 80100.0 141750.0 ;
      RECT  81300.0 142950.0 80100.0 141750.0 ;
      RECT  83700.0 142950.0 82500.0 141750.0 ;
      RECT  78900.0 133050.0 77700.0 131850.0 ;
      RECT  78900.0 142950.0 77700.0 141750.0 ;
      RECT  83100.0 138300.0 81900.0 137100.0 ;
      RECT  83100.0 138300.0 81900.0 137100.0 ;
      RECT  80550.0 138150.0 79650.0 137250.0 ;
      RECT  85500.0 130950.0 75900.0 130050.0 ;
      RECT  85500.0 144750.0 75900.0 143850.0 ;
      RECT  98100.0 91050.0 96900.0 88650.0 ;
      RECT  98100.0 99750.0 96900.0 103350.0 ;
      RECT  93300.0 99750.0 92100.0 103350.0 ;
      RECT  90900.0 100950.0 89700.0 102900.0 ;
      RECT  90900.0 89100.0 89700.0 91050.0 ;
      RECT  98100.0 99750.0 96900.0 100950.0 ;
      RECT  95700.0 99750.0 94500.0 100950.0 ;
      RECT  95700.0 99750.0 94500.0 100950.0 ;
      RECT  98100.0 99750.0 96900.0 100950.0 ;
      RECT  95700.0 99750.0 94500.0 100950.0 ;
      RECT  93300.0 99750.0 92100.0 100950.0 ;
      RECT  93300.0 99750.0 92100.0 100950.0 ;
      RECT  95700.0 99750.0 94500.0 100950.0 ;
      RECT  98100.0 91050.0 96900.0 92250.0 ;
      RECT  95700.0 91050.0 94500.0 92250.0 ;
      RECT  95700.0 91050.0 94500.0 92250.0 ;
      RECT  98100.0 91050.0 96900.0 92250.0 ;
      RECT  95700.0 91050.0 94500.0 92250.0 ;
      RECT  93300.0 91050.0 92100.0 92250.0 ;
      RECT  93300.0 91050.0 92100.0 92250.0 ;
      RECT  95700.0 91050.0 94500.0 92250.0 ;
      RECT  90900.0 100350.0 89700.0 101550.0 ;
      RECT  90900.0 90450.0 89700.0 91650.0 ;
      RECT  93300.0 93600.0 94500.0 94800.0 ;
      RECT  96300.0 96300.0 97500.0 97500.0 ;
      RECT  95700.0 99750.0 94500.0 100950.0 ;
      RECT  93300.0 91050.0 92100.0 92250.0 ;
      RECT  92100.0 96300.0 93300.0 97500.0 ;
      RECT  97500.0 96300.0 96300.0 97500.0 ;
      RECT  94500.0 93600.0 93300.0 94800.0 ;
      RECT  93300.0 96300.0 92100.0 97500.0 ;
      RECT  99900.0 102450.0 85500.0 103350.0 ;
      RECT  99900.0 88650.0 85500.0 89550.0 ;
      RECT  98100.0 114750.0 96900.0 117150.0 ;
      RECT  98100.0 106050.0 96900.0 102450.0 ;
      RECT  93300.0 106050.0 92100.0 102450.0 ;
      RECT  90900.0 104850.0 89700.0 102900.0 ;
      RECT  90900.0 116700.0 89700.0 114750.0 ;
      RECT  98100.0 106050.0 96900.0 104850.0 ;
      RECT  95700.0 106050.0 94500.0 104850.0 ;
      RECT  95700.0 106050.0 94500.0 104850.0 ;
      RECT  98100.0 106050.0 96900.0 104850.0 ;
      RECT  95700.0 106050.0 94500.0 104850.0 ;
      RECT  93300.0 106050.0 92100.0 104850.0 ;
      RECT  93300.0 106050.0 92100.0 104850.0 ;
      RECT  95700.0 106050.0 94500.0 104850.0 ;
      RECT  98100.0 114750.0 96900.0 113550.0 ;
      RECT  95700.0 114750.0 94500.0 113550.0 ;
      RECT  95700.0 114750.0 94500.0 113550.0 ;
      RECT  98100.0 114750.0 96900.0 113550.0 ;
      RECT  95700.0 114750.0 94500.0 113550.0 ;
      RECT  93300.0 114750.0 92100.0 113550.0 ;
      RECT  93300.0 114750.0 92100.0 113550.0 ;
      RECT  95700.0 114750.0 94500.0 113550.0 ;
      RECT  90900.0 105450.0 89700.0 104250.0 ;
      RECT  90900.0 115350.0 89700.0 114150.0 ;
      RECT  93300.0 112200.0 94500.0 111000.0 ;
      RECT  96300.0 109500.0 97500.0 108300.0 ;
      RECT  95700.0 106050.0 94500.0 104850.0 ;
      RECT  93300.0 114750.0 92100.0 113550.0 ;
      RECT  92100.0 109500.0 93300.0 108300.0 ;
      RECT  97500.0 109500.0 96300.0 108300.0 ;
      RECT  94500.0 112200.0 93300.0 111000.0 ;
      RECT  93300.0 109500.0 92100.0 108300.0 ;
      RECT  99900.0 103350.0 85500.0 102450.0 ;
      RECT  99900.0 117150.0 85500.0 116250.0 ;
      RECT  98100.0 118650.0 96900.0 116250.0 ;
      RECT  98100.0 127350.0 96900.0 130950.0 ;
      RECT  93300.0 127350.0 92100.0 130950.0 ;
      RECT  90900.0 128550.0 89700.0 130500.0 ;
      RECT  90900.0 116700.0 89700.0 118650.0 ;
      RECT  98100.0 127350.0 96900.0 128550.0 ;
      RECT  95700.0 127350.0 94500.0 128550.0 ;
      RECT  95700.0 127350.0 94500.0 128550.0 ;
      RECT  98100.0 127350.0 96900.0 128550.0 ;
      RECT  95700.0 127350.0 94500.0 128550.0 ;
      RECT  93300.0 127350.0 92100.0 128550.0 ;
      RECT  93300.0 127350.0 92100.0 128550.0 ;
      RECT  95700.0 127350.0 94500.0 128550.0 ;
      RECT  98100.0 118650.0 96900.0 119850.0 ;
      RECT  95700.0 118650.0 94500.0 119850.0 ;
      RECT  95700.0 118650.0 94500.0 119850.0 ;
      RECT  98100.0 118650.0 96900.0 119850.0 ;
      RECT  95700.0 118650.0 94500.0 119850.0 ;
      RECT  93300.0 118650.0 92100.0 119850.0 ;
      RECT  93300.0 118650.0 92100.0 119850.0 ;
      RECT  95700.0 118650.0 94500.0 119850.0 ;
      RECT  90900.0 127950.0 89700.0 129150.0 ;
      RECT  90900.0 118050.0 89700.0 119250.0 ;
      RECT  93300.0 121200.0 94500.0 122400.0 ;
      RECT  96300.0 123900.0 97500.0 125100.0 ;
      RECT  95700.0 127350.0 94500.0 128550.0 ;
      RECT  93300.0 118650.0 92100.0 119850.0 ;
      RECT  92100.0 123900.0 93300.0 125100.0 ;
      RECT  97500.0 123900.0 96300.0 125100.0 ;
      RECT  94500.0 121200.0 93300.0 122400.0 ;
      RECT  93300.0 123900.0 92100.0 125100.0 ;
      RECT  99900.0 130050.0 85500.0 130950.0 ;
      RECT  99900.0 116250.0 85500.0 117150.0 ;
      RECT  98100.0 142350.0 96900.0 144750.0 ;
      RECT  98100.0 133650.0 96900.0 130050.0 ;
      RECT  93300.0 133650.0 92100.0 130050.0 ;
      RECT  90900.0 132450.0 89700.0 130500.0 ;
      RECT  90900.0 144300.0 89700.0 142350.0 ;
      RECT  98100.0 133650.0 96900.0 132450.0 ;
      RECT  95700.0 133650.0 94500.0 132450.0 ;
      RECT  95700.0 133650.0 94500.0 132450.0 ;
      RECT  98100.0 133650.0 96900.0 132450.0 ;
      RECT  95700.0 133650.0 94500.0 132450.0 ;
      RECT  93300.0 133650.0 92100.0 132450.0 ;
      RECT  93300.0 133650.0 92100.0 132450.0 ;
      RECT  95700.0 133650.0 94500.0 132450.0 ;
      RECT  98100.0 142350.0 96900.0 141150.0 ;
      RECT  95700.0 142350.0 94500.0 141150.0 ;
      RECT  95700.0 142350.0 94500.0 141150.0 ;
      RECT  98100.0 142350.0 96900.0 141150.0 ;
      RECT  95700.0 142350.0 94500.0 141150.0 ;
      RECT  93300.0 142350.0 92100.0 141150.0 ;
      RECT  93300.0 142350.0 92100.0 141150.0 ;
      RECT  95700.0 142350.0 94500.0 141150.0 ;
      RECT  90900.0 133050.0 89700.0 131850.0 ;
      RECT  90900.0 142950.0 89700.0 141750.0 ;
      RECT  93300.0 139800.0 94500.0 138600.0 ;
      RECT  96300.0 137100.0 97500.0 135900.0 ;
      RECT  95700.0 133650.0 94500.0 132450.0 ;
      RECT  93300.0 142350.0 92100.0 141150.0 ;
      RECT  92100.0 137100.0 93300.0 135900.0 ;
      RECT  97500.0 137100.0 96300.0 135900.0 ;
      RECT  94500.0 139800.0 93300.0 138600.0 ;
      RECT  93300.0 137100.0 92100.0 135900.0 ;
      RECT  99900.0 130950.0 85500.0 130050.0 ;
      RECT  99900.0 144750.0 85500.0 143850.0 ;
      RECT  110850.0 99600.0 112050.0 100800.0 ;
      RECT  129450.0 95100.0 130650.0 96300.0 ;
      RECT  107850.0 113400.0 109050.0 114600.0 ;
      RECT  126450.0 109500.0 127650.0 110700.0 ;
      RECT  129450.0 118200.0 130650.0 119400.0 ;
      RECT  104850.0 118200.0 106050.0 119400.0 ;
      RECT  126450.0 132000.0 127650.0 133200.0 ;
      RECT  101850.0 132000.0 103050.0 133200.0 ;
      RECT  110850.0 96300.0 112050.0 97500.0 ;
      RECT  107850.0 93600.0 109050.0 94800.0 ;
      RECT  104850.0 108300.0 106050.0 109500.0 ;
      RECT  107850.0 111000.0 109050.0 112200.0 ;
      RECT  110850.0 123900.0 112050.0 125100.0 ;
      RECT  101850.0 121200.0 103050.0 122400.0 ;
      RECT  104850.0 135900.0 106050.0 137100.0 ;
      RECT  101850.0 138600.0 103050.0 139800.0 ;
      RECT  79650.0 95250.0 75900.0 96150.0 ;
      RECT  79650.0 109650.0 75900.0 110550.0 ;
      RECT  79650.0 122850.0 75900.0 123750.0 ;
      RECT  79650.0 137250.0 75900.0 138150.0 ;
      RECT  130500.0 102450.0 75900.0 103350.0 ;
      RECT  130500.0 130050.0 75900.0 130950.0 ;
      RECT  130500.0 88650.0 75900.0 89550.0 ;
      RECT  130500.0 116250.0 75900.0 117150.0 ;
      RECT  130500.0 143850.0 75900.0 144750.0 ;
      RECT  114450.0 150450.0 113550.0 151350.0 ;
      RECT  114450.0 154950.0 113550.0 155850.0 ;
      RECT  118650.0 150450.0 114000.0 151350.0 ;
      RECT  114450.0 150900.0 113550.0 155400.0 ;
      RECT  114000.0 154950.0 111450.0 155850.0 ;
      RECT  130050.0 150450.0 122100.0 151350.0 ;
      RECT  114450.0 164850.0 113550.0 165750.0 ;
      RECT  114450.0 168750.0 113550.0 169650.0 ;
      RECT  118650.0 164850.0 114000.0 165750.0 ;
      RECT  114450.0 165300.0 113550.0 169200.0 ;
      RECT  114000.0 168750.0 108450.0 169650.0 ;
      RECT  127050.0 164850.0 122100.0 165750.0 ;
      RECT  130050.0 173550.0 105450.0 174450.0 ;
      RECT  127050.0 187350.0 102450.0 188250.0 ;
      RECT  111450.0 151650.0 97500.0 152550.0 ;
      RECT  108450.0 148950.0 94500.0 149850.0 ;
      RECT  105450.0 163650.0 97500.0 164550.0 ;
      RECT  108450.0 166350.0 94500.0 167250.0 ;
      RECT  111450.0 179250.0 97500.0 180150.0 ;
      RECT  102450.0 176550.0 94500.0 177450.0 ;
      RECT  105450.0 191250.0 97500.0 192150.0 ;
      RECT  102450.0 193950.0 94500.0 194850.0 ;
      RECT  88050.0 151650.0 87150.0 152550.0 ;
      RECT  88050.0 150450.0 87150.0 151350.0 ;
      RECT  92100.0 151650.0 87600.0 152550.0 ;
      RECT  88050.0 150900.0 87150.0 152100.0 ;
      RECT  87600.0 150450.0 83100.0 151350.0 ;
      RECT  88050.0 163650.0 87150.0 164550.0 ;
      RECT  88050.0 164850.0 87150.0 165750.0 ;
      RECT  92100.0 163650.0 87600.0 164550.0 ;
      RECT  88050.0 164100.0 87150.0 165300.0 ;
      RECT  87600.0 164850.0 83100.0 165750.0 ;
      RECT  88050.0 179250.0 87150.0 180150.0 ;
      RECT  88050.0 178050.0 87150.0 178950.0 ;
      RECT  92100.0 179250.0 87600.0 180150.0 ;
      RECT  88050.0 178500.0 87150.0 179700.0 ;
      RECT  87600.0 178050.0 83100.0 178950.0 ;
      RECT  88050.0 191250.0 87150.0 192150.0 ;
      RECT  88050.0 192450.0 87150.0 193350.0 ;
      RECT  92100.0 191250.0 87600.0 192150.0 ;
      RECT  88050.0 191700.0 87150.0 192900.0 ;
      RECT  87600.0 192450.0 83100.0 193350.0 ;
      RECT  117900.0 156150.0 116700.0 158100.0 ;
      RECT  117900.0 144300.0 116700.0 146250.0 ;
      RECT  122700.0 145650.0 121500.0 143850.0 ;
      RECT  122700.0 154950.0 121500.0 158550.0 ;
      RECT  120000.0 145650.0 119100.0 154950.0 ;
      RECT  122700.0 154950.0 121500.0 156150.0 ;
      RECT  120300.0 154950.0 119100.0 156150.0 ;
      RECT  120300.0 154950.0 119100.0 156150.0 ;
      RECT  122700.0 154950.0 121500.0 156150.0 ;
      RECT  122700.0 145650.0 121500.0 146850.0 ;
      RECT  120300.0 145650.0 119100.0 146850.0 ;
      RECT  120300.0 145650.0 119100.0 146850.0 ;
      RECT  122700.0 145650.0 121500.0 146850.0 ;
      RECT  117900.0 155550.0 116700.0 156750.0 ;
      RECT  117900.0 145650.0 116700.0 146850.0 ;
      RECT  122100.0 150300.0 120900.0 151500.0 ;
      RECT  122100.0 150300.0 120900.0 151500.0 ;
      RECT  119550.0 150450.0 118650.0 151350.0 ;
      RECT  124500.0 157650.0 114900.0 158550.0 ;
      RECT  124500.0 143850.0 114900.0 144750.0 ;
      RECT  117900.0 160050.0 116700.0 158100.0 ;
      RECT  117900.0 171900.0 116700.0 169950.0 ;
      RECT  122700.0 170550.0 121500.0 172350.0 ;
      RECT  122700.0 161250.0 121500.0 157650.0 ;
      RECT  120000.0 170550.0 119100.0 161250.0 ;
      RECT  122700.0 161250.0 121500.0 160050.0 ;
      RECT  120300.0 161250.0 119100.0 160050.0 ;
      RECT  120300.0 161250.0 119100.0 160050.0 ;
      RECT  122700.0 161250.0 121500.0 160050.0 ;
      RECT  122700.0 170550.0 121500.0 169350.0 ;
      RECT  120300.0 170550.0 119100.0 169350.0 ;
      RECT  120300.0 170550.0 119100.0 169350.0 ;
      RECT  122700.0 170550.0 121500.0 169350.0 ;
      RECT  117900.0 160650.0 116700.0 159450.0 ;
      RECT  117900.0 170550.0 116700.0 169350.0 ;
      RECT  122100.0 165900.0 120900.0 164700.0 ;
      RECT  122100.0 165900.0 120900.0 164700.0 ;
      RECT  119550.0 165750.0 118650.0 164850.0 ;
      RECT  124500.0 158550.0 114900.0 157650.0 ;
      RECT  124500.0 172350.0 114900.0 171450.0 ;
      RECT  78900.0 156150.0 77700.0 158100.0 ;
      RECT  78900.0 144300.0 77700.0 146250.0 ;
      RECT  83700.0 145650.0 82500.0 143850.0 ;
      RECT  83700.0 154950.0 82500.0 158550.0 ;
      RECT  81000.0 145650.0 80100.0 154950.0 ;
      RECT  83700.0 154950.0 82500.0 156150.0 ;
      RECT  81300.0 154950.0 80100.0 156150.0 ;
      RECT  81300.0 154950.0 80100.0 156150.0 ;
      RECT  83700.0 154950.0 82500.0 156150.0 ;
      RECT  83700.0 145650.0 82500.0 146850.0 ;
      RECT  81300.0 145650.0 80100.0 146850.0 ;
      RECT  81300.0 145650.0 80100.0 146850.0 ;
      RECT  83700.0 145650.0 82500.0 146850.0 ;
      RECT  78900.0 155550.0 77700.0 156750.0 ;
      RECT  78900.0 145650.0 77700.0 146850.0 ;
      RECT  83100.0 150300.0 81900.0 151500.0 ;
      RECT  83100.0 150300.0 81900.0 151500.0 ;
      RECT  80550.0 150450.0 79650.0 151350.0 ;
      RECT  85500.0 157650.0 75900.0 158550.0 ;
      RECT  85500.0 143850.0 75900.0 144750.0 ;
      RECT  78900.0 160050.0 77700.0 158100.0 ;
      RECT  78900.0 171900.0 77700.0 169950.0 ;
      RECT  83700.0 170550.0 82500.0 172350.0 ;
      RECT  83700.0 161250.0 82500.0 157650.0 ;
      RECT  81000.0 170550.0 80100.0 161250.0 ;
      RECT  83700.0 161250.0 82500.0 160050.0 ;
      RECT  81300.0 161250.0 80100.0 160050.0 ;
      RECT  81300.0 161250.0 80100.0 160050.0 ;
      RECT  83700.0 161250.0 82500.0 160050.0 ;
      RECT  83700.0 170550.0 82500.0 169350.0 ;
      RECT  81300.0 170550.0 80100.0 169350.0 ;
      RECT  81300.0 170550.0 80100.0 169350.0 ;
      RECT  83700.0 170550.0 82500.0 169350.0 ;
      RECT  78900.0 160650.0 77700.0 159450.0 ;
      RECT  78900.0 170550.0 77700.0 169350.0 ;
      RECT  83100.0 165900.0 81900.0 164700.0 ;
      RECT  83100.0 165900.0 81900.0 164700.0 ;
      RECT  80550.0 165750.0 79650.0 164850.0 ;
      RECT  85500.0 158550.0 75900.0 157650.0 ;
      RECT  85500.0 172350.0 75900.0 171450.0 ;
      RECT  78900.0 183750.0 77700.0 185700.0 ;
      RECT  78900.0 171900.0 77700.0 173850.0 ;
      RECT  83700.0 173250.0 82500.0 171450.0 ;
      RECT  83700.0 182550.0 82500.0 186150.0 ;
      RECT  81000.0 173250.0 80100.0 182550.0 ;
      RECT  83700.0 182550.0 82500.0 183750.0 ;
      RECT  81300.0 182550.0 80100.0 183750.0 ;
      RECT  81300.0 182550.0 80100.0 183750.0 ;
      RECT  83700.0 182550.0 82500.0 183750.0 ;
      RECT  83700.0 173250.0 82500.0 174450.0 ;
      RECT  81300.0 173250.0 80100.0 174450.0 ;
      RECT  81300.0 173250.0 80100.0 174450.0 ;
      RECT  83700.0 173250.0 82500.0 174450.0 ;
      RECT  78900.0 183150.0 77700.0 184350.0 ;
      RECT  78900.0 173250.0 77700.0 174450.0 ;
      RECT  83100.0 177900.0 81900.0 179100.0 ;
      RECT  83100.0 177900.0 81900.0 179100.0 ;
      RECT  80550.0 178050.0 79650.0 178950.0 ;
      RECT  85500.0 185250.0 75900.0 186150.0 ;
      RECT  85500.0 171450.0 75900.0 172350.0 ;
      RECT  78900.0 187650.0 77700.0 185700.0 ;
      RECT  78900.0 199500.0 77700.0 197550.0 ;
      RECT  83700.0 198150.0 82500.0 199950.0 ;
      RECT  83700.0 188850.0 82500.0 185250.0 ;
      RECT  81000.0 198150.0 80100.0 188850.0 ;
      RECT  83700.0 188850.0 82500.0 187650.0 ;
      RECT  81300.0 188850.0 80100.0 187650.0 ;
      RECT  81300.0 188850.0 80100.0 187650.0 ;
      RECT  83700.0 188850.0 82500.0 187650.0 ;
      RECT  83700.0 198150.0 82500.0 196950.0 ;
      RECT  81300.0 198150.0 80100.0 196950.0 ;
      RECT  81300.0 198150.0 80100.0 196950.0 ;
      RECT  83700.0 198150.0 82500.0 196950.0 ;
      RECT  78900.0 188250.0 77700.0 187050.0 ;
      RECT  78900.0 198150.0 77700.0 196950.0 ;
      RECT  83100.0 193500.0 81900.0 192300.0 ;
      RECT  83100.0 193500.0 81900.0 192300.0 ;
      RECT  80550.0 193350.0 79650.0 192450.0 ;
      RECT  85500.0 186150.0 75900.0 185250.0 ;
      RECT  85500.0 199950.0 75900.0 199050.0 ;
      RECT  98100.0 146250.0 96900.0 143850.0 ;
      RECT  98100.0 154950.0 96900.0 158550.0 ;
      RECT  93300.0 154950.0 92100.0 158550.0 ;
      RECT  90900.0 156150.0 89700.0 158100.0 ;
      RECT  90900.0 144300.0 89700.0 146250.0 ;
      RECT  98100.0 154950.0 96900.0 156150.0 ;
      RECT  95700.0 154950.0 94500.0 156150.0 ;
      RECT  95700.0 154950.0 94500.0 156150.0 ;
      RECT  98100.0 154950.0 96900.0 156150.0 ;
      RECT  95700.0 154950.0 94500.0 156150.0 ;
      RECT  93300.0 154950.0 92100.0 156150.0 ;
      RECT  93300.0 154950.0 92100.0 156150.0 ;
      RECT  95700.0 154950.0 94500.0 156150.0 ;
      RECT  98100.0 146250.0 96900.0 147450.0 ;
      RECT  95700.0 146250.0 94500.0 147450.0 ;
      RECT  95700.0 146250.0 94500.0 147450.0 ;
      RECT  98100.0 146250.0 96900.0 147450.0 ;
      RECT  95700.0 146250.0 94500.0 147450.0 ;
      RECT  93300.0 146250.0 92100.0 147450.0 ;
      RECT  93300.0 146250.0 92100.0 147450.0 ;
      RECT  95700.0 146250.0 94500.0 147450.0 ;
      RECT  90900.0 155550.0 89700.0 156750.0 ;
      RECT  90900.0 145650.0 89700.0 146850.0 ;
      RECT  93300.0 148800.0 94500.0 150000.0 ;
      RECT  96300.0 151500.0 97500.0 152700.0 ;
      RECT  95700.0 154950.0 94500.0 156150.0 ;
      RECT  93300.0 146250.0 92100.0 147450.0 ;
      RECT  92100.0 151500.0 93300.0 152700.0 ;
      RECT  97500.0 151500.0 96300.0 152700.0 ;
      RECT  94500.0 148800.0 93300.0 150000.0 ;
      RECT  93300.0 151500.0 92100.0 152700.0 ;
      RECT  99900.0 157650.0 85500.0 158550.0 ;
      RECT  99900.0 143850.0 85500.0 144750.0 ;
      RECT  98100.0 169950.0 96900.0 172350.0 ;
      RECT  98100.0 161250.0 96900.0 157650.0 ;
      RECT  93300.0 161250.0 92100.0 157650.0 ;
      RECT  90900.0 160050.0 89700.0 158100.0 ;
      RECT  90900.0 171900.0 89700.0 169950.0 ;
      RECT  98100.0 161250.0 96900.0 160050.0 ;
      RECT  95700.0 161250.0 94500.0 160050.0 ;
      RECT  95700.0 161250.0 94500.0 160050.0 ;
      RECT  98100.0 161250.0 96900.0 160050.0 ;
      RECT  95700.0 161250.0 94500.0 160050.0 ;
      RECT  93300.0 161250.0 92100.0 160050.0 ;
      RECT  93300.0 161250.0 92100.0 160050.0 ;
      RECT  95700.0 161250.0 94500.0 160050.0 ;
      RECT  98100.0 169950.0 96900.0 168750.0 ;
      RECT  95700.0 169950.0 94500.0 168750.0 ;
      RECT  95700.0 169950.0 94500.0 168750.0 ;
      RECT  98100.0 169950.0 96900.0 168750.0 ;
      RECT  95700.0 169950.0 94500.0 168750.0 ;
      RECT  93300.0 169950.0 92100.0 168750.0 ;
      RECT  93300.0 169950.0 92100.0 168750.0 ;
      RECT  95700.0 169950.0 94500.0 168750.0 ;
      RECT  90900.0 160650.0 89700.0 159450.0 ;
      RECT  90900.0 170550.0 89700.0 169350.0 ;
      RECT  93300.0 167400.0 94500.0 166200.0 ;
      RECT  96300.0 164700.0 97500.0 163500.0 ;
      RECT  95700.0 161250.0 94500.0 160050.0 ;
      RECT  93300.0 169950.0 92100.0 168750.0 ;
      RECT  92100.0 164700.0 93300.0 163500.0 ;
      RECT  97500.0 164700.0 96300.0 163500.0 ;
      RECT  94500.0 167400.0 93300.0 166200.0 ;
      RECT  93300.0 164700.0 92100.0 163500.0 ;
      RECT  99900.0 158550.0 85500.0 157650.0 ;
      RECT  99900.0 172350.0 85500.0 171450.0 ;
      RECT  98100.0 173850.0 96900.0 171450.0 ;
      RECT  98100.0 182550.0 96900.0 186150.0 ;
      RECT  93300.0 182550.0 92100.0 186150.0 ;
      RECT  90900.0 183750.0 89700.0 185700.0 ;
      RECT  90900.0 171900.0 89700.0 173850.0 ;
      RECT  98100.0 182550.0 96900.0 183750.0 ;
      RECT  95700.0 182550.0 94500.0 183750.0 ;
      RECT  95700.0 182550.0 94500.0 183750.0 ;
      RECT  98100.0 182550.0 96900.0 183750.0 ;
      RECT  95700.0 182550.0 94500.0 183750.0 ;
      RECT  93300.0 182550.0 92100.0 183750.0 ;
      RECT  93300.0 182550.0 92100.0 183750.0 ;
      RECT  95700.0 182550.0 94500.0 183750.0 ;
      RECT  98100.0 173850.0 96900.0 175050.0 ;
      RECT  95700.0 173850.0 94500.0 175050.0 ;
      RECT  95700.0 173850.0 94500.0 175050.0 ;
      RECT  98100.0 173850.0 96900.0 175050.0 ;
      RECT  95700.0 173850.0 94500.0 175050.0 ;
      RECT  93300.0 173850.0 92100.0 175050.0 ;
      RECT  93300.0 173850.0 92100.0 175050.0 ;
      RECT  95700.0 173850.0 94500.0 175050.0 ;
      RECT  90900.0 183150.0 89700.0 184350.0 ;
      RECT  90900.0 173250.0 89700.0 174450.0 ;
      RECT  93300.0 176400.0 94500.0 177600.0 ;
      RECT  96300.0 179100.0 97500.0 180300.0 ;
      RECT  95700.0 182550.0 94500.0 183750.0 ;
      RECT  93300.0 173850.0 92100.0 175050.0 ;
      RECT  92100.0 179100.0 93300.0 180300.0 ;
      RECT  97500.0 179100.0 96300.0 180300.0 ;
      RECT  94500.0 176400.0 93300.0 177600.0 ;
      RECT  93300.0 179100.0 92100.0 180300.0 ;
      RECT  99900.0 185250.0 85500.0 186150.0 ;
      RECT  99900.0 171450.0 85500.0 172350.0 ;
      RECT  98100.0 197550.0 96900.0 199950.0 ;
      RECT  98100.0 188850.0 96900.0 185250.0 ;
      RECT  93300.0 188850.0 92100.0 185250.0 ;
      RECT  90900.0 187650.0 89700.0 185700.0 ;
      RECT  90900.0 199500.0 89700.0 197550.0 ;
      RECT  98100.0 188850.0 96900.0 187650.0 ;
      RECT  95700.0 188850.0 94500.0 187650.0 ;
      RECT  95700.0 188850.0 94500.0 187650.0 ;
      RECT  98100.0 188850.0 96900.0 187650.0 ;
      RECT  95700.0 188850.0 94500.0 187650.0 ;
      RECT  93300.0 188850.0 92100.0 187650.0 ;
      RECT  93300.0 188850.0 92100.0 187650.0 ;
      RECT  95700.0 188850.0 94500.0 187650.0 ;
      RECT  98100.0 197550.0 96900.0 196350.0 ;
      RECT  95700.0 197550.0 94500.0 196350.0 ;
      RECT  95700.0 197550.0 94500.0 196350.0 ;
      RECT  98100.0 197550.0 96900.0 196350.0 ;
      RECT  95700.0 197550.0 94500.0 196350.0 ;
      RECT  93300.0 197550.0 92100.0 196350.0 ;
      RECT  93300.0 197550.0 92100.0 196350.0 ;
      RECT  95700.0 197550.0 94500.0 196350.0 ;
      RECT  90900.0 188250.0 89700.0 187050.0 ;
      RECT  90900.0 198150.0 89700.0 196950.0 ;
      RECT  93300.0 195000.0 94500.0 193800.0 ;
      RECT  96300.0 192300.0 97500.0 191100.0 ;
      RECT  95700.0 188850.0 94500.0 187650.0 ;
      RECT  93300.0 197550.0 92100.0 196350.0 ;
      RECT  92100.0 192300.0 93300.0 191100.0 ;
      RECT  97500.0 192300.0 96300.0 191100.0 ;
      RECT  94500.0 195000.0 93300.0 193800.0 ;
      RECT  93300.0 192300.0 92100.0 191100.0 ;
      RECT  99900.0 186150.0 85500.0 185250.0 ;
      RECT  99900.0 199950.0 85500.0 199050.0 ;
      RECT  110850.0 154800.0 112050.0 156000.0 ;
      RECT  129450.0 150300.0 130650.0 151500.0 ;
      RECT  107850.0 168600.0 109050.0 169800.0 ;
      RECT  126450.0 164700.0 127650.0 165900.0 ;
      RECT  129450.0 173400.0 130650.0 174600.0 ;
      RECT  104850.0 173400.0 106050.0 174600.0 ;
      RECT  126450.0 187200.0 127650.0 188400.0 ;
      RECT  101850.0 187200.0 103050.0 188400.0 ;
      RECT  110850.0 151500.0 112050.0 152700.0 ;
      RECT  107850.0 148800.0 109050.0 150000.0 ;
      RECT  104850.0 163500.0 106050.0 164700.0 ;
      RECT  107850.0 166200.0 109050.0 167400.0 ;
      RECT  110850.0 179100.0 112050.0 180300.0 ;
      RECT  101850.0 176400.0 103050.0 177600.0 ;
      RECT  104850.0 191100.0 106050.0 192300.0 ;
      RECT  101850.0 193800.0 103050.0 195000.0 ;
      RECT  79650.0 150450.0 75900.0 151350.0 ;
      RECT  79650.0 164850.0 75900.0 165750.0 ;
      RECT  79650.0 178050.0 75900.0 178950.0 ;
      RECT  79650.0 192450.0 75900.0 193350.0 ;
      RECT  130500.0 157650.0 75900.0 158550.0 ;
      RECT  130500.0 185250.0 75900.0 186150.0 ;
      RECT  130500.0 143850.0 75900.0 144750.0 ;
      RECT  130500.0 171450.0 75900.0 172350.0 ;
      RECT  130500.0 199050.0 75900.0 199950.0 ;
      RECT  77700.0 201450.0 78900.0 199050.0 ;
      RECT  77700.0 210150.0 78900.0 213750.0 ;
      RECT  82500.0 210150.0 83700.0 213750.0 ;
      RECT  84900.0 211350.0 86100.0 213300.0 ;
      RECT  84900.0 199500.0 86100.0 201450.0 ;
      RECT  77700.0 210150.0 78900.0 211350.0 ;
      RECT  80100.0 210150.0 81300.0 211350.0 ;
      RECT  80100.0 210150.0 81300.0 211350.0 ;
      RECT  77700.0 210150.0 78900.0 211350.0 ;
      RECT  80100.0 210150.0 81300.0 211350.0 ;
      RECT  82500.0 210150.0 83700.0 211350.0 ;
      RECT  82500.0 210150.0 83700.0 211350.0 ;
      RECT  80100.0 210150.0 81300.0 211350.0 ;
      RECT  77700.0 201450.0 78900.0 202650.0 ;
      RECT  80100.0 201450.0 81300.0 202650.0 ;
      RECT  80100.0 201450.0 81300.0 202650.0 ;
      RECT  77700.0 201450.0 78900.0 202650.0 ;
      RECT  80100.0 201450.0 81300.0 202650.0 ;
      RECT  82500.0 201450.0 83700.0 202650.0 ;
      RECT  82500.0 201450.0 83700.0 202650.0 ;
      RECT  80100.0 201450.0 81300.0 202650.0 ;
      RECT  84900.0 210750.0 86100.0 211950.0 ;
      RECT  84900.0 200850.0 86100.0 202050.0 ;
      RECT  82500.0 204000.0 81300.0 205200.0 ;
      RECT  79500.0 206700.0 78300.0 207900.0 ;
      RECT  80100.0 210150.0 81300.0 211350.0 ;
      RECT  82500.0 201450.0 83700.0 202650.0 ;
      RECT  83700.0 206700.0 82500.0 207900.0 ;
      RECT  78300.0 206700.0 79500.0 207900.0 ;
      RECT  81300.0 204000.0 82500.0 205200.0 ;
      RECT  82500.0 206700.0 83700.0 207900.0 ;
      RECT  75900.0 212850.0 90300.0 213750.0 ;
      RECT  75900.0 199050.0 90300.0 199950.0 ;
      RECT  77700.0 225150.0 78900.0 227550.0 ;
      RECT  77700.0 216450.0 78900.0 212850.0 ;
      RECT  82500.0 216450.0 83700.0 212850.0 ;
      RECT  84900.0 215250.0 86100.0 213300.0 ;
      RECT  84900.0 227100.0 86100.0 225150.0 ;
      RECT  77700.0 216450.0 78900.0 215250.0 ;
      RECT  80100.0 216450.0 81300.0 215250.0 ;
      RECT  80100.0 216450.0 81300.0 215250.0 ;
      RECT  77700.0 216450.0 78900.0 215250.0 ;
      RECT  80100.0 216450.0 81300.0 215250.0 ;
      RECT  82500.0 216450.0 83700.0 215250.0 ;
      RECT  82500.0 216450.0 83700.0 215250.0 ;
      RECT  80100.0 216450.0 81300.0 215250.0 ;
      RECT  77700.0 225150.0 78900.0 223950.0 ;
      RECT  80100.0 225150.0 81300.0 223950.0 ;
      RECT  80100.0 225150.0 81300.0 223950.0 ;
      RECT  77700.0 225150.0 78900.0 223950.0 ;
      RECT  80100.0 225150.0 81300.0 223950.0 ;
      RECT  82500.0 225150.0 83700.0 223950.0 ;
      RECT  82500.0 225150.0 83700.0 223950.0 ;
      RECT  80100.0 225150.0 81300.0 223950.0 ;
      RECT  84900.0 215850.0 86100.0 214650.0 ;
      RECT  84900.0 225750.0 86100.0 224550.0 ;
      RECT  82500.0 222600.0 81300.0 221400.0 ;
      RECT  79500.0 219900.0 78300.0 218700.0 ;
      RECT  80100.0 216450.0 81300.0 215250.0 ;
      RECT  82500.0 225150.0 83700.0 223950.0 ;
      RECT  83700.0 219900.0 82500.0 218700.0 ;
      RECT  78300.0 219900.0 79500.0 218700.0 ;
      RECT  81300.0 222600.0 82500.0 221400.0 ;
      RECT  82500.0 219900.0 83700.0 218700.0 ;
      RECT  75900.0 213750.0 90300.0 212850.0 ;
      RECT  75900.0 227550.0 90300.0 226650.0 ;
      RECT  77700.0 229050.0 78900.0 226650.0 ;
      RECT  77700.0 237750.0 78900.0 241350.0 ;
      RECT  82500.0 237750.0 83700.0 241350.0 ;
      RECT  84900.0 238950.0 86100.0 240900.0 ;
      RECT  84900.0 227100.0 86100.0 229050.0 ;
      RECT  77700.0 237750.0 78900.0 238950.0 ;
      RECT  80100.0 237750.0 81300.0 238950.0 ;
      RECT  80100.0 237750.0 81300.0 238950.0 ;
      RECT  77700.0 237750.0 78900.0 238950.0 ;
      RECT  80100.0 237750.0 81300.0 238950.0 ;
      RECT  82500.0 237750.0 83700.0 238950.0 ;
      RECT  82500.0 237750.0 83700.0 238950.0 ;
      RECT  80100.0 237750.0 81300.0 238950.0 ;
      RECT  77700.0 229050.0 78900.0 230250.0 ;
      RECT  80100.0 229050.0 81300.0 230250.0 ;
      RECT  80100.0 229050.0 81300.0 230250.0 ;
      RECT  77700.0 229050.0 78900.0 230250.0 ;
      RECT  80100.0 229050.0 81300.0 230250.0 ;
      RECT  82500.0 229050.0 83700.0 230250.0 ;
      RECT  82500.0 229050.0 83700.0 230250.0 ;
      RECT  80100.0 229050.0 81300.0 230250.0 ;
      RECT  84900.0 238350.0 86100.0 239550.0 ;
      RECT  84900.0 228450.0 86100.0 229650.0 ;
      RECT  82500.0 231600.0 81300.0 232800.0 ;
      RECT  79500.0 234300.0 78300.0 235500.0 ;
      RECT  80100.0 237750.0 81300.0 238950.0 ;
      RECT  82500.0 229050.0 83700.0 230250.0 ;
      RECT  83700.0 234300.0 82500.0 235500.0 ;
      RECT  78300.0 234300.0 79500.0 235500.0 ;
      RECT  81300.0 231600.0 82500.0 232800.0 ;
      RECT  82500.0 234300.0 83700.0 235500.0 ;
      RECT  75900.0 240450.0 90300.0 241350.0 ;
      RECT  75900.0 226650.0 90300.0 227550.0 ;
      RECT  77700.0 252750.0 78900.0 255150.0 ;
      RECT  77700.0 244050.0 78900.0 240450.0 ;
      RECT  82500.0 244050.0 83700.0 240450.0 ;
      RECT  84900.0 242850.0 86100.0 240900.0 ;
      RECT  84900.0 254700.0 86100.0 252750.0 ;
      RECT  77700.0 244050.0 78900.0 242850.0 ;
      RECT  80100.0 244050.0 81300.0 242850.0 ;
      RECT  80100.0 244050.0 81300.0 242850.0 ;
      RECT  77700.0 244050.0 78900.0 242850.0 ;
      RECT  80100.0 244050.0 81300.0 242850.0 ;
      RECT  82500.0 244050.0 83700.0 242850.0 ;
      RECT  82500.0 244050.0 83700.0 242850.0 ;
      RECT  80100.0 244050.0 81300.0 242850.0 ;
      RECT  77700.0 252750.0 78900.0 251550.0 ;
      RECT  80100.0 252750.0 81300.0 251550.0 ;
      RECT  80100.0 252750.0 81300.0 251550.0 ;
      RECT  77700.0 252750.0 78900.0 251550.0 ;
      RECT  80100.0 252750.0 81300.0 251550.0 ;
      RECT  82500.0 252750.0 83700.0 251550.0 ;
      RECT  82500.0 252750.0 83700.0 251550.0 ;
      RECT  80100.0 252750.0 81300.0 251550.0 ;
      RECT  84900.0 243450.0 86100.0 242250.0 ;
      RECT  84900.0 253350.0 86100.0 252150.0 ;
      RECT  82500.0 250200.0 81300.0 249000.0 ;
      RECT  79500.0 247500.0 78300.0 246300.0 ;
      RECT  80100.0 244050.0 81300.0 242850.0 ;
      RECT  82500.0 252750.0 83700.0 251550.0 ;
      RECT  83700.0 247500.0 82500.0 246300.0 ;
      RECT  78300.0 247500.0 79500.0 246300.0 ;
      RECT  81300.0 250200.0 82500.0 249000.0 ;
      RECT  82500.0 247500.0 83700.0 246300.0 ;
      RECT  75900.0 241350.0 90300.0 240450.0 ;
      RECT  75900.0 255150.0 90300.0 254250.0 ;
      RECT  77700.0 256650.0 78900.0 254250.0 ;
      RECT  77700.0 265350.0 78900.0 268950.0 ;
      RECT  82500.0 265350.0 83700.0 268950.0 ;
      RECT  84900.0 266550.0 86100.0 268500.0 ;
      RECT  84900.0 254700.0 86100.0 256650.0 ;
      RECT  77700.0 265350.0 78900.0 266550.0 ;
      RECT  80100.0 265350.0 81300.0 266550.0 ;
      RECT  80100.0 265350.0 81300.0 266550.0 ;
      RECT  77700.0 265350.0 78900.0 266550.0 ;
      RECT  80100.0 265350.0 81300.0 266550.0 ;
      RECT  82500.0 265350.0 83700.0 266550.0 ;
      RECT  82500.0 265350.0 83700.0 266550.0 ;
      RECT  80100.0 265350.0 81300.0 266550.0 ;
      RECT  77700.0 256650.0 78900.0 257850.0 ;
      RECT  80100.0 256650.0 81300.0 257850.0 ;
      RECT  80100.0 256650.0 81300.0 257850.0 ;
      RECT  77700.0 256650.0 78900.0 257850.0 ;
      RECT  80100.0 256650.0 81300.0 257850.0 ;
      RECT  82500.0 256650.0 83700.0 257850.0 ;
      RECT  82500.0 256650.0 83700.0 257850.0 ;
      RECT  80100.0 256650.0 81300.0 257850.0 ;
      RECT  84900.0 265950.0 86100.0 267150.0 ;
      RECT  84900.0 256050.0 86100.0 257250.0 ;
      RECT  82500.0 259200.0 81300.0 260400.0 ;
      RECT  79500.0 261900.0 78300.0 263100.0 ;
      RECT  80100.0 265350.0 81300.0 266550.0 ;
      RECT  82500.0 256650.0 83700.0 257850.0 ;
      RECT  83700.0 261900.0 82500.0 263100.0 ;
      RECT  78300.0 261900.0 79500.0 263100.0 ;
      RECT  81300.0 259200.0 82500.0 260400.0 ;
      RECT  82500.0 261900.0 83700.0 263100.0 ;
      RECT  75900.0 268050.0 90300.0 268950.0 ;
      RECT  75900.0 254250.0 90300.0 255150.0 ;
      RECT  77700.0 280350.0 78900.0 282750.0 ;
      RECT  77700.0 271650.0 78900.0 268050.0 ;
      RECT  82500.0 271650.0 83700.0 268050.0 ;
      RECT  84900.0 270450.0 86100.0 268500.0 ;
      RECT  84900.0 282300.0 86100.0 280350.0 ;
      RECT  77700.0 271650.0 78900.0 270450.0 ;
      RECT  80100.0 271650.0 81300.0 270450.0 ;
      RECT  80100.0 271650.0 81300.0 270450.0 ;
      RECT  77700.0 271650.0 78900.0 270450.0 ;
      RECT  80100.0 271650.0 81300.0 270450.0 ;
      RECT  82500.0 271650.0 83700.0 270450.0 ;
      RECT  82500.0 271650.0 83700.0 270450.0 ;
      RECT  80100.0 271650.0 81300.0 270450.0 ;
      RECT  77700.0 280350.0 78900.0 279150.0 ;
      RECT  80100.0 280350.0 81300.0 279150.0 ;
      RECT  80100.0 280350.0 81300.0 279150.0 ;
      RECT  77700.0 280350.0 78900.0 279150.0 ;
      RECT  80100.0 280350.0 81300.0 279150.0 ;
      RECT  82500.0 280350.0 83700.0 279150.0 ;
      RECT  82500.0 280350.0 83700.0 279150.0 ;
      RECT  80100.0 280350.0 81300.0 279150.0 ;
      RECT  84900.0 271050.0 86100.0 269850.0 ;
      RECT  84900.0 280950.0 86100.0 279750.0 ;
      RECT  82500.0 277800.0 81300.0 276600.0 ;
      RECT  79500.0 275100.0 78300.0 273900.0 ;
      RECT  80100.0 271650.0 81300.0 270450.0 ;
      RECT  82500.0 280350.0 83700.0 279150.0 ;
      RECT  83700.0 275100.0 82500.0 273900.0 ;
      RECT  78300.0 275100.0 79500.0 273900.0 ;
      RECT  81300.0 277800.0 82500.0 276600.0 ;
      RECT  82500.0 275100.0 83700.0 273900.0 ;
      RECT  75900.0 268950.0 90300.0 268050.0 ;
      RECT  75900.0 282750.0 90300.0 281850.0 ;
      RECT  77700.0 284250.0 78900.0 281850.0 ;
      RECT  77700.0 292950.0 78900.0 296550.0 ;
      RECT  82500.0 292950.0 83700.0 296550.0 ;
      RECT  84900.0 294150.0 86100.0 296100.0 ;
      RECT  84900.0 282300.0 86100.0 284250.0 ;
      RECT  77700.0 292950.0 78900.0 294150.0 ;
      RECT  80100.0 292950.0 81300.0 294150.0 ;
      RECT  80100.0 292950.0 81300.0 294150.0 ;
      RECT  77700.0 292950.0 78900.0 294150.0 ;
      RECT  80100.0 292950.0 81300.0 294150.0 ;
      RECT  82500.0 292950.0 83700.0 294150.0 ;
      RECT  82500.0 292950.0 83700.0 294150.0 ;
      RECT  80100.0 292950.0 81300.0 294150.0 ;
      RECT  77700.0 284250.0 78900.0 285450.0 ;
      RECT  80100.0 284250.0 81300.0 285450.0 ;
      RECT  80100.0 284250.0 81300.0 285450.0 ;
      RECT  77700.0 284250.0 78900.0 285450.0 ;
      RECT  80100.0 284250.0 81300.0 285450.0 ;
      RECT  82500.0 284250.0 83700.0 285450.0 ;
      RECT  82500.0 284250.0 83700.0 285450.0 ;
      RECT  80100.0 284250.0 81300.0 285450.0 ;
      RECT  84900.0 293550.0 86100.0 294750.0 ;
      RECT  84900.0 283650.0 86100.0 284850.0 ;
      RECT  82500.0 286800.0 81300.0 288000.0 ;
      RECT  79500.0 289500.0 78300.0 290700.0 ;
      RECT  80100.0 292950.0 81300.0 294150.0 ;
      RECT  82500.0 284250.0 83700.0 285450.0 ;
      RECT  83700.0 289500.0 82500.0 290700.0 ;
      RECT  78300.0 289500.0 79500.0 290700.0 ;
      RECT  81300.0 286800.0 82500.0 288000.0 ;
      RECT  82500.0 289500.0 83700.0 290700.0 ;
      RECT  75900.0 295650.0 90300.0 296550.0 ;
      RECT  75900.0 281850.0 90300.0 282750.0 ;
      RECT  77700.0 307950.0 78900.0 310350.0 ;
      RECT  77700.0 299250.0 78900.0 295650.0 ;
      RECT  82500.0 299250.0 83700.0 295650.0 ;
      RECT  84900.0 298050.0 86100.0 296100.0 ;
      RECT  84900.0 309900.0 86100.0 307950.0 ;
      RECT  77700.0 299250.0 78900.0 298050.0 ;
      RECT  80100.0 299250.0 81300.0 298050.0 ;
      RECT  80100.0 299250.0 81300.0 298050.0 ;
      RECT  77700.0 299250.0 78900.0 298050.0 ;
      RECT  80100.0 299250.0 81300.0 298050.0 ;
      RECT  82500.0 299250.0 83700.0 298050.0 ;
      RECT  82500.0 299250.0 83700.0 298050.0 ;
      RECT  80100.0 299250.0 81300.0 298050.0 ;
      RECT  77700.0 307950.0 78900.0 306750.0 ;
      RECT  80100.0 307950.0 81300.0 306750.0 ;
      RECT  80100.0 307950.0 81300.0 306750.0 ;
      RECT  77700.0 307950.0 78900.0 306750.0 ;
      RECT  80100.0 307950.0 81300.0 306750.0 ;
      RECT  82500.0 307950.0 83700.0 306750.0 ;
      RECT  82500.0 307950.0 83700.0 306750.0 ;
      RECT  80100.0 307950.0 81300.0 306750.0 ;
      RECT  84900.0 298650.0 86100.0 297450.0 ;
      RECT  84900.0 308550.0 86100.0 307350.0 ;
      RECT  82500.0 305400.0 81300.0 304200.0 ;
      RECT  79500.0 302700.0 78300.0 301500.0 ;
      RECT  80100.0 299250.0 81300.0 298050.0 ;
      RECT  82500.0 307950.0 83700.0 306750.0 ;
      RECT  83700.0 302700.0 82500.0 301500.0 ;
      RECT  78300.0 302700.0 79500.0 301500.0 ;
      RECT  81300.0 305400.0 82500.0 304200.0 ;
      RECT  82500.0 302700.0 83700.0 301500.0 ;
      RECT  75900.0 296550.0 90300.0 295650.0 ;
      RECT  75900.0 310350.0 90300.0 309450.0 ;
      RECT  77700.0 311850.0 78900.0 309450.0 ;
      RECT  77700.0 320550.0 78900.0 324150.0 ;
      RECT  82500.0 320550.0 83700.0 324150.0 ;
      RECT  84900.0 321750.0 86100.0 323700.0 ;
      RECT  84900.0 309900.0 86100.0 311850.0 ;
      RECT  77700.0 320550.0 78900.0 321750.0 ;
      RECT  80100.0 320550.0 81300.0 321750.0 ;
      RECT  80100.0 320550.0 81300.0 321750.0 ;
      RECT  77700.0 320550.0 78900.0 321750.0 ;
      RECT  80100.0 320550.0 81300.0 321750.0 ;
      RECT  82500.0 320550.0 83700.0 321750.0 ;
      RECT  82500.0 320550.0 83700.0 321750.0 ;
      RECT  80100.0 320550.0 81300.0 321750.0 ;
      RECT  77700.0 311850.0 78900.0 313050.0 ;
      RECT  80100.0 311850.0 81300.0 313050.0 ;
      RECT  80100.0 311850.0 81300.0 313050.0 ;
      RECT  77700.0 311850.0 78900.0 313050.0 ;
      RECT  80100.0 311850.0 81300.0 313050.0 ;
      RECT  82500.0 311850.0 83700.0 313050.0 ;
      RECT  82500.0 311850.0 83700.0 313050.0 ;
      RECT  80100.0 311850.0 81300.0 313050.0 ;
      RECT  84900.0 321150.0 86100.0 322350.0 ;
      RECT  84900.0 311250.0 86100.0 312450.0 ;
      RECT  82500.0 314400.0 81300.0 315600.0 ;
      RECT  79500.0 317100.0 78300.0 318300.0 ;
      RECT  80100.0 320550.0 81300.0 321750.0 ;
      RECT  82500.0 311850.0 83700.0 313050.0 ;
      RECT  83700.0 317100.0 82500.0 318300.0 ;
      RECT  78300.0 317100.0 79500.0 318300.0 ;
      RECT  81300.0 314400.0 82500.0 315600.0 ;
      RECT  82500.0 317100.0 83700.0 318300.0 ;
      RECT  75900.0 323250.0 90300.0 324150.0 ;
      RECT  75900.0 309450.0 90300.0 310350.0 ;
      RECT  77700.0 335550.0 78900.0 337950.0 ;
      RECT  77700.0 326850.0 78900.0 323250.0 ;
      RECT  82500.0 326850.0 83700.0 323250.0 ;
      RECT  84900.0 325650.0 86100.0 323700.0 ;
      RECT  84900.0 337500.0 86100.0 335550.0 ;
      RECT  77700.0 326850.0 78900.0 325650.0 ;
      RECT  80100.0 326850.0 81300.0 325650.0 ;
      RECT  80100.0 326850.0 81300.0 325650.0 ;
      RECT  77700.0 326850.0 78900.0 325650.0 ;
      RECT  80100.0 326850.0 81300.0 325650.0 ;
      RECT  82500.0 326850.0 83700.0 325650.0 ;
      RECT  82500.0 326850.0 83700.0 325650.0 ;
      RECT  80100.0 326850.0 81300.0 325650.0 ;
      RECT  77700.0 335550.0 78900.0 334350.0 ;
      RECT  80100.0 335550.0 81300.0 334350.0 ;
      RECT  80100.0 335550.0 81300.0 334350.0 ;
      RECT  77700.0 335550.0 78900.0 334350.0 ;
      RECT  80100.0 335550.0 81300.0 334350.0 ;
      RECT  82500.0 335550.0 83700.0 334350.0 ;
      RECT  82500.0 335550.0 83700.0 334350.0 ;
      RECT  80100.0 335550.0 81300.0 334350.0 ;
      RECT  84900.0 326250.0 86100.0 325050.0 ;
      RECT  84900.0 336150.0 86100.0 334950.0 ;
      RECT  82500.0 333000.0 81300.0 331800.0 ;
      RECT  79500.0 330300.0 78300.0 329100.0 ;
      RECT  80100.0 326850.0 81300.0 325650.0 ;
      RECT  82500.0 335550.0 83700.0 334350.0 ;
      RECT  83700.0 330300.0 82500.0 329100.0 ;
      RECT  78300.0 330300.0 79500.0 329100.0 ;
      RECT  81300.0 333000.0 82500.0 331800.0 ;
      RECT  82500.0 330300.0 83700.0 329100.0 ;
      RECT  75900.0 324150.0 90300.0 323250.0 ;
      RECT  75900.0 337950.0 90300.0 337050.0 ;
      RECT  77700.0 339450.0 78900.0 337050.0 ;
      RECT  77700.0 348150.0 78900.0 351750.0 ;
      RECT  82500.0 348150.0 83700.0 351750.0 ;
      RECT  84900.0 349350.0 86100.0 351300.0 ;
      RECT  84900.0 337500.0 86100.0 339450.0 ;
      RECT  77700.0 348150.0 78900.0 349350.0 ;
      RECT  80100.0 348150.0 81300.0 349350.0 ;
      RECT  80100.0 348150.0 81300.0 349350.0 ;
      RECT  77700.0 348150.0 78900.0 349350.0 ;
      RECT  80100.0 348150.0 81300.0 349350.0 ;
      RECT  82500.0 348150.0 83700.0 349350.0 ;
      RECT  82500.0 348150.0 83700.0 349350.0 ;
      RECT  80100.0 348150.0 81300.0 349350.0 ;
      RECT  77700.0 339450.0 78900.0 340650.0 ;
      RECT  80100.0 339450.0 81300.0 340650.0 ;
      RECT  80100.0 339450.0 81300.0 340650.0 ;
      RECT  77700.0 339450.0 78900.0 340650.0 ;
      RECT  80100.0 339450.0 81300.0 340650.0 ;
      RECT  82500.0 339450.0 83700.0 340650.0 ;
      RECT  82500.0 339450.0 83700.0 340650.0 ;
      RECT  80100.0 339450.0 81300.0 340650.0 ;
      RECT  84900.0 348750.0 86100.0 349950.0 ;
      RECT  84900.0 338850.0 86100.0 340050.0 ;
      RECT  82500.0 342000.0 81300.0 343200.0 ;
      RECT  79500.0 344700.0 78300.0 345900.0 ;
      RECT  80100.0 348150.0 81300.0 349350.0 ;
      RECT  82500.0 339450.0 83700.0 340650.0 ;
      RECT  83700.0 344700.0 82500.0 345900.0 ;
      RECT  78300.0 344700.0 79500.0 345900.0 ;
      RECT  81300.0 342000.0 82500.0 343200.0 ;
      RECT  82500.0 344700.0 83700.0 345900.0 ;
      RECT  75900.0 350850.0 90300.0 351750.0 ;
      RECT  75900.0 337050.0 90300.0 337950.0 ;
      RECT  77700.0 363150.0 78900.0 365550.0 ;
      RECT  77700.0 354450.0 78900.0 350850.0 ;
      RECT  82500.0 354450.0 83700.0 350850.0 ;
      RECT  84900.0 353250.0 86100.0 351300.0 ;
      RECT  84900.0 365100.0 86100.0 363150.0 ;
      RECT  77700.0 354450.0 78900.0 353250.0 ;
      RECT  80100.0 354450.0 81300.0 353250.0 ;
      RECT  80100.0 354450.0 81300.0 353250.0 ;
      RECT  77700.0 354450.0 78900.0 353250.0 ;
      RECT  80100.0 354450.0 81300.0 353250.0 ;
      RECT  82500.0 354450.0 83700.0 353250.0 ;
      RECT  82500.0 354450.0 83700.0 353250.0 ;
      RECT  80100.0 354450.0 81300.0 353250.0 ;
      RECT  77700.0 363150.0 78900.0 361950.0 ;
      RECT  80100.0 363150.0 81300.0 361950.0 ;
      RECT  80100.0 363150.0 81300.0 361950.0 ;
      RECT  77700.0 363150.0 78900.0 361950.0 ;
      RECT  80100.0 363150.0 81300.0 361950.0 ;
      RECT  82500.0 363150.0 83700.0 361950.0 ;
      RECT  82500.0 363150.0 83700.0 361950.0 ;
      RECT  80100.0 363150.0 81300.0 361950.0 ;
      RECT  84900.0 353850.0 86100.0 352650.0 ;
      RECT  84900.0 363750.0 86100.0 362550.0 ;
      RECT  82500.0 360600.0 81300.0 359400.0 ;
      RECT  79500.0 357900.0 78300.0 356700.0 ;
      RECT  80100.0 354450.0 81300.0 353250.0 ;
      RECT  82500.0 363150.0 83700.0 361950.0 ;
      RECT  83700.0 357900.0 82500.0 356700.0 ;
      RECT  78300.0 357900.0 79500.0 356700.0 ;
      RECT  81300.0 360600.0 82500.0 359400.0 ;
      RECT  82500.0 357900.0 83700.0 356700.0 ;
      RECT  75900.0 351750.0 90300.0 350850.0 ;
      RECT  75900.0 365550.0 90300.0 364650.0 ;
      RECT  77700.0 367050.0 78900.0 364650.0 ;
      RECT  77700.0 375750.0 78900.0 379350.0 ;
      RECT  82500.0 375750.0 83700.0 379350.0 ;
      RECT  84900.0 376950.0 86100.0 378900.0 ;
      RECT  84900.0 365100.0 86100.0 367050.0 ;
      RECT  77700.0 375750.0 78900.0 376950.0 ;
      RECT  80100.0 375750.0 81300.0 376950.0 ;
      RECT  80100.0 375750.0 81300.0 376950.0 ;
      RECT  77700.0 375750.0 78900.0 376950.0 ;
      RECT  80100.0 375750.0 81300.0 376950.0 ;
      RECT  82500.0 375750.0 83700.0 376950.0 ;
      RECT  82500.0 375750.0 83700.0 376950.0 ;
      RECT  80100.0 375750.0 81300.0 376950.0 ;
      RECT  77700.0 367050.0 78900.0 368250.0 ;
      RECT  80100.0 367050.0 81300.0 368250.0 ;
      RECT  80100.0 367050.0 81300.0 368250.0 ;
      RECT  77700.0 367050.0 78900.0 368250.0 ;
      RECT  80100.0 367050.0 81300.0 368250.0 ;
      RECT  82500.0 367050.0 83700.0 368250.0 ;
      RECT  82500.0 367050.0 83700.0 368250.0 ;
      RECT  80100.0 367050.0 81300.0 368250.0 ;
      RECT  84900.0 376350.0 86100.0 377550.0 ;
      RECT  84900.0 366450.0 86100.0 367650.0 ;
      RECT  82500.0 369600.0 81300.0 370800.0 ;
      RECT  79500.0 372300.0 78300.0 373500.0 ;
      RECT  80100.0 375750.0 81300.0 376950.0 ;
      RECT  82500.0 367050.0 83700.0 368250.0 ;
      RECT  83700.0 372300.0 82500.0 373500.0 ;
      RECT  78300.0 372300.0 79500.0 373500.0 ;
      RECT  81300.0 369600.0 82500.0 370800.0 ;
      RECT  82500.0 372300.0 83700.0 373500.0 ;
      RECT  75900.0 378450.0 90300.0 379350.0 ;
      RECT  75900.0 364650.0 90300.0 365550.0 ;
      RECT  77700.0 390750.0 78900.0 393150.0 ;
      RECT  77700.0 382050.0 78900.0 378450.0 ;
      RECT  82500.0 382050.0 83700.0 378450.0 ;
      RECT  84900.0 380850.0 86100.0 378900.0 ;
      RECT  84900.0 392700.0 86100.0 390750.0 ;
      RECT  77700.0 382050.0 78900.0 380850.0 ;
      RECT  80100.0 382050.0 81300.0 380850.0 ;
      RECT  80100.0 382050.0 81300.0 380850.0 ;
      RECT  77700.0 382050.0 78900.0 380850.0 ;
      RECT  80100.0 382050.0 81300.0 380850.0 ;
      RECT  82500.0 382050.0 83700.0 380850.0 ;
      RECT  82500.0 382050.0 83700.0 380850.0 ;
      RECT  80100.0 382050.0 81300.0 380850.0 ;
      RECT  77700.0 390750.0 78900.0 389550.0 ;
      RECT  80100.0 390750.0 81300.0 389550.0 ;
      RECT  80100.0 390750.0 81300.0 389550.0 ;
      RECT  77700.0 390750.0 78900.0 389550.0 ;
      RECT  80100.0 390750.0 81300.0 389550.0 ;
      RECT  82500.0 390750.0 83700.0 389550.0 ;
      RECT  82500.0 390750.0 83700.0 389550.0 ;
      RECT  80100.0 390750.0 81300.0 389550.0 ;
      RECT  84900.0 381450.0 86100.0 380250.0 ;
      RECT  84900.0 391350.0 86100.0 390150.0 ;
      RECT  82500.0 388200.0 81300.0 387000.0 ;
      RECT  79500.0 385500.0 78300.0 384300.0 ;
      RECT  80100.0 382050.0 81300.0 380850.0 ;
      RECT  82500.0 390750.0 83700.0 389550.0 ;
      RECT  83700.0 385500.0 82500.0 384300.0 ;
      RECT  78300.0 385500.0 79500.0 384300.0 ;
      RECT  81300.0 388200.0 82500.0 387000.0 ;
      RECT  82500.0 385500.0 83700.0 384300.0 ;
      RECT  75900.0 379350.0 90300.0 378450.0 ;
      RECT  75900.0 393150.0 90300.0 392250.0 ;
      RECT  77700.0 394650.0 78900.0 392250.0 ;
      RECT  77700.0 403350.0 78900.0 406950.0 ;
      RECT  82500.0 403350.0 83700.0 406950.0 ;
      RECT  84900.0 404550.0 86100.0 406500.0 ;
      RECT  84900.0 392700.0 86100.0 394650.0 ;
      RECT  77700.0 403350.0 78900.0 404550.0 ;
      RECT  80100.0 403350.0 81300.0 404550.0 ;
      RECT  80100.0 403350.0 81300.0 404550.0 ;
      RECT  77700.0 403350.0 78900.0 404550.0 ;
      RECT  80100.0 403350.0 81300.0 404550.0 ;
      RECT  82500.0 403350.0 83700.0 404550.0 ;
      RECT  82500.0 403350.0 83700.0 404550.0 ;
      RECT  80100.0 403350.0 81300.0 404550.0 ;
      RECT  77700.0 394650.0 78900.0 395850.0 ;
      RECT  80100.0 394650.0 81300.0 395850.0 ;
      RECT  80100.0 394650.0 81300.0 395850.0 ;
      RECT  77700.0 394650.0 78900.0 395850.0 ;
      RECT  80100.0 394650.0 81300.0 395850.0 ;
      RECT  82500.0 394650.0 83700.0 395850.0 ;
      RECT  82500.0 394650.0 83700.0 395850.0 ;
      RECT  80100.0 394650.0 81300.0 395850.0 ;
      RECT  84900.0 403950.0 86100.0 405150.0 ;
      RECT  84900.0 394050.0 86100.0 395250.0 ;
      RECT  82500.0 397200.0 81300.0 398400.0 ;
      RECT  79500.0 399900.0 78300.0 401100.0 ;
      RECT  80100.0 403350.0 81300.0 404550.0 ;
      RECT  82500.0 394650.0 83700.0 395850.0 ;
      RECT  83700.0 399900.0 82500.0 401100.0 ;
      RECT  78300.0 399900.0 79500.0 401100.0 ;
      RECT  81300.0 397200.0 82500.0 398400.0 ;
      RECT  82500.0 399900.0 83700.0 401100.0 ;
      RECT  75900.0 406050.0 90300.0 406950.0 ;
      RECT  75900.0 392250.0 90300.0 393150.0 ;
      RECT  77700.0 418350.0 78900.0 420750.0 ;
      RECT  77700.0 409650.0 78900.0 406050.0 ;
      RECT  82500.0 409650.0 83700.0 406050.0 ;
      RECT  84900.0 408450.0 86100.0 406500.0 ;
      RECT  84900.0 420300.0 86100.0 418350.0 ;
      RECT  77700.0 409650.0 78900.0 408450.0 ;
      RECT  80100.0 409650.0 81300.0 408450.0 ;
      RECT  80100.0 409650.0 81300.0 408450.0 ;
      RECT  77700.0 409650.0 78900.0 408450.0 ;
      RECT  80100.0 409650.0 81300.0 408450.0 ;
      RECT  82500.0 409650.0 83700.0 408450.0 ;
      RECT  82500.0 409650.0 83700.0 408450.0 ;
      RECT  80100.0 409650.0 81300.0 408450.0 ;
      RECT  77700.0 418350.0 78900.0 417150.0 ;
      RECT  80100.0 418350.0 81300.0 417150.0 ;
      RECT  80100.0 418350.0 81300.0 417150.0 ;
      RECT  77700.0 418350.0 78900.0 417150.0 ;
      RECT  80100.0 418350.0 81300.0 417150.0 ;
      RECT  82500.0 418350.0 83700.0 417150.0 ;
      RECT  82500.0 418350.0 83700.0 417150.0 ;
      RECT  80100.0 418350.0 81300.0 417150.0 ;
      RECT  84900.0 409050.0 86100.0 407850.0 ;
      RECT  84900.0 418950.0 86100.0 417750.0 ;
      RECT  82500.0 415800.0 81300.0 414600.0 ;
      RECT  79500.0 413100.0 78300.0 411900.0 ;
      RECT  80100.0 409650.0 81300.0 408450.0 ;
      RECT  82500.0 418350.0 83700.0 417150.0 ;
      RECT  83700.0 413100.0 82500.0 411900.0 ;
      RECT  78300.0 413100.0 79500.0 411900.0 ;
      RECT  81300.0 415800.0 82500.0 414600.0 ;
      RECT  82500.0 413100.0 83700.0 411900.0 ;
      RECT  75900.0 406950.0 90300.0 406050.0 ;
      RECT  75900.0 420750.0 90300.0 419850.0 ;
      RECT  96900.0 211350.0 98100.0 213300.0 ;
      RECT  96900.0 199500.0 98100.0 201450.0 ;
      RECT  92100.0 200850.0 93300.0 199050.0 ;
      RECT  92100.0 210150.0 93300.0 213750.0 ;
      RECT  94800.0 200850.0 95700.0 210150.0 ;
      RECT  92100.0 210150.0 93300.0 211350.0 ;
      RECT  94500.0 210150.0 95700.0 211350.0 ;
      RECT  94500.0 210150.0 95700.0 211350.0 ;
      RECT  92100.0 210150.0 93300.0 211350.0 ;
      RECT  92100.0 200850.0 93300.0 202050.0 ;
      RECT  94500.0 200850.0 95700.0 202050.0 ;
      RECT  94500.0 200850.0 95700.0 202050.0 ;
      RECT  92100.0 200850.0 93300.0 202050.0 ;
      RECT  96900.0 210750.0 98100.0 211950.0 ;
      RECT  96900.0 200850.0 98100.0 202050.0 ;
      RECT  92700.0 205500.0 93900.0 206700.0 ;
      RECT  92700.0 205500.0 93900.0 206700.0 ;
      RECT  95250.0 205650.0 96150.0 206550.0 ;
      RECT  90300.0 212850.0 99900.0 213750.0 ;
      RECT  90300.0 199050.0 99900.0 199950.0 ;
      RECT  96900.0 215250.0 98100.0 213300.0 ;
      RECT  96900.0 227100.0 98100.0 225150.0 ;
      RECT  92100.0 225750.0 93300.0 227550.0 ;
      RECT  92100.0 216450.0 93300.0 212850.0 ;
      RECT  94800.0 225750.0 95700.0 216450.0 ;
      RECT  92100.0 216450.0 93300.0 215250.0 ;
      RECT  94500.0 216450.0 95700.0 215250.0 ;
      RECT  94500.0 216450.0 95700.0 215250.0 ;
      RECT  92100.0 216450.0 93300.0 215250.0 ;
      RECT  92100.0 225750.0 93300.0 224550.0 ;
      RECT  94500.0 225750.0 95700.0 224550.0 ;
      RECT  94500.0 225750.0 95700.0 224550.0 ;
      RECT  92100.0 225750.0 93300.0 224550.0 ;
      RECT  96900.0 215850.0 98100.0 214650.0 ;
      RECT  96900.0 225750.0 98100.0 224550.0 ;
      RECT  92700.0 221100.0 93900.0 219900.0 ;
      RECT  92700.0 221100.0 93900.0 219900.0 ;
      RECT  95250.0 220950.0 96150.0 220050.0 ;
      RECT  90300.0 213750.0 99900.0 212850.0 ;
      RECT  90300.0 227550.0 99900.0 226650.0 ;
      RECT  96900.0 238950.0 98100.0 240900.0 ;
      RECT  96900.0 227100.0 98100.0 229050.0 ;
      RECT  92100.0 228450.0 93300.0 226650.0 ;
      RECT  92100.0 237750.0 93300.0 241350.0 ;
      RECT  94800.0 228450.0 95700.0 237750.0 ;
      RECT  92100.0 237750.0 93300.0 238950.0 ;
      RECT  94500.0 237750.0 95700.0 238950.0 ;
      RECT  94500.0 237750.0 95700.0 238950.0 ;
      RECT  92100.0 237750.0 93300.0 238950.0 ;
      RECT  92100.0 228450.0 93300.0 229650.0 ;
      RECT  94500.0 228450.0 95700.0 229650.0 ;
      RECT  94500.0 228450.0 95700.0 229650.0 ;
      RECT  92100.0 228450.0 93300.0 229650.0 ;
      RECT  96900.0 238350.0 98100.0 239550.0 ;
      RECT  96900.0 228450.0 98100.0 229650.0 ;
      RECT  92700.0 233100.0 93900.0 234300.0 ;
      RECT  92700.0 233100.0 93900.0 234300.0 ;
      RECT  95250.0 233250.0 96150.0 234150.0 ;
      RECT  90300.0 240450.0 99900.0 241350.0 ;
      RECT  90300.0 226650.0 99900.0 227550.0 ;
      RECT  96900.0 242850.0 98100.0 240900.0 ;
      RECT  96900.0 254700.0 98100.0 252750.0 ;
      RECT  92100.0 253350.0 93300.0 255150.0 ;
      RECT  92100.0 244050.0 93300.0 240450.0 ;
      RECT  94800.0 253350.0 95700.0 244050.0 ;
      RECT  92100.0 244050.0 93300.0 242850.0 ;
      RECT  94500.0 244050.0 95700.0 242850.0 ;
      RECT  94500.0 244050.0 95700.0 242850.0 ;
      RECT  92100.0 244050.0 93300.0 242850.0 ;
      RECT  92100.0 253350.0 93300.0 252150.0 ;
      RECT  94500.0 253350.0 95700.0 252150.0 ;
      RECT  94500.0 253350.0 95700.0 252150.0 ;
      RECT  92100.0 253350.0 93300.0 252150.0 ;
      RECT  96900.0 243450.0 98100.0 242250.0 ;
      RECT  96900.0 253350.0 98100.0 252150.0 ;
      RECT  92700.0 248700.0 93900.0 247500.0 ;
      RECT  92700.0 248700.0 93900.0 247500.0 ;
      RECT  95250.0 248550.0 96150.0 247650.0 ;
      RECT  90300.0 241350.0 99900.0 240450.0 ;
      RECT  90300.0 255150.0 99900.0 254250.0 ;
      RECT  96900.0 266550.0 98100.0 268500.0 ;
      RECT  96900.0 254700.0 98100.0 256650.0 ;
      RECT  92100.0 256050.0 93300.0 254250.0 ;
      RECT  92100.0 265350.0 93300.0 268950.0 ;
      RECT  94800.0 256050.0 95700.0 265350.0 ;
      RECT  92100.0 265350.0 93300.0 266550.0 ;
      RECT  94500.0 265350.0 95700.0 266550.0 ;
      RECT  94500.0 265350.0 95700.0 266550.0 ;
      RECT  92100.0 265350.0 93300.0 266550.0 ;
      RECT  92100.0 256050.0 93300.0 257250.0 ;
      RECT  94500.0 256050.0 95700.0 257250.0 ;
      RECT  94500.0 256050.0 95700.0 257250.0 ;
      RECT  92100.0 256050.0 93300.0 257250.0 ;
      RECT  96900.0 265950.0 98100.0 267150.0 ;
      RECT  96900.0 256050.0 98100.0 257250.0 ;
      RECT  92700.0 260700.0 93900.0 261900.0 ;
      RECT  92700.0 260700.0 93900.0 261900.0 ;
      RECT  95250.0 260850.0 96150.0 261750.0 ;
      RECT  90300.0 268050.0 99900.0 268950.0 ;
      RECT  90300.0 254250.0 99900.0 255150.0 ;
      RECT  96900.0 270450.0 98100.0 268500.0 ;
      RECT  96900.0 282300.0 98100.0 280350.0 ;
      RECT  92100.0 280950.0 93300.0 282750.0 ;
      RECT  92100.0 271650.0 93300.0 268050.0 ;
      RECT  94800.0 280950.0 95700.0 271650.0 ;
      RECT  92100.0 271650.0 93300.0 270450.0 ;
      RECT  94500.0 271650.0 95700.0 270450.0 ;
      RECT  94500.0 271650.0 95700.0 270450.0 ;
      RECT  92100.0 271650.0 93300.0 270450.0 ;
      RECT  92100.0 280950.0 93300.0 279750.0 ;
      RECT  94500.0 280950.0 95700.0 279750.0 ;
      RECT  94500.0 280950.0 95700.0 279750.0 ;
      RECT  92100.0 280950.0 93300.0 279750.0 ;
      RECT  96900.0 271050.0 98100.0 269850.0 ;
      RECT  96900.0 280950.0 98100.0 279750.0 ;
      RECT  92700.0 276300.0 93900.0 275100.0 ;
      RECT  92700.0 276300.0 93900.0 275100.0 ;
      RECT  95250.0 276150.0 96150.0 275250.0 ;
      RECT  90300.0 268950.0 99900.0 268050.0 ;
      RECT  90300.0 282750.0 99900.0 281850.0 ;
      RECT  96900.0 294150.0 98100.0 296100.0 ;
      RECT  96900.0 282300.0 98100.0 284250.0 ;
      RECT  92100.0 283650.0 93300.0 281850.0 ;
      RECT  92100.0 292950.0 93300.0 296550.0 ;
      RECT  94800.0 283650.0 95700.0 292950.0 ;
      RECT  92100.0 292950.0 93300.0 294150.0 ;
      RECT  94500.0 292950.0 95700.0 294150.0 ;
      RECT  94500.0 292950.0 95700.0 294150.0 ;
      RECT  92100.0 292950.0 93300.0 294150.0 ;
      RECT  92100.0 283650.0 93300.0 284850.0 ;
      RECT  94500.0 283650.0 95700.0 284850.0 ;
      RECT  94500.0 283650.0 95700.0 284850.0 ;
      RECT  92100.0 283650.0 93300.0 284850.0 ;
      RECT  96900.0 293550.0 98100.0 294750.0 ;
      RECT  96900.0 283650.0 98100.0 284850.0 ;
      RECT  92700.0 288300.0 93900.0 289500.0 ;
      RECT  92700.0 288300.0 93900.0 289500.0 ;
      RECT  95250.0 288450.0 96150.0 289350.0 ;
      RECT  90300.0 295650.0 99900.0 296550.0 ;
      RECT  90300.0 281850.0 99900.0 282750.0 ;
      RECT  96900.0 298050.0 98100.0 296100.0 ;
      RECT  96900.0 309900.0 98100.0 307950.0 ;
      RECT  92100.0 308550.0 93300.0 310350.0 ;
      RECT  92100.0 299250.0 93300.0 295650.0 ;
      RECT  94800.0 308550.0 95700.0 299250.0 ;
      RECT  92100.0 299250.0 93300.0 298050.0 ;
      RECT  94500.0 299250.0 95700.0 298050.0 ;
      RECT  94500.0 299250.0 95700.0 298050.0 ;
      RECT  92100.0 299250.0 93300.0 298050.0 ;
      RECT  92100.0 308550.0 93300.0 307350.0 ;
      RECT  94500.0 308550.0 95700.0 307350.0 ;
      RECT  94500.0 308550.0 95700.0 307350.0 ;
      RECT  92100.0 308550.0 93300.0 307350.0 ;
      RECT  96900.0 298650.0 98100.0 297450.0 ;
      RECT  96900.0 308550.0 98100.0 307350.0 ;
      RECT  92700.0 303900.0 93900.0 302700.0 ;
      RECT  92700.0 303900.0 93900.0 302700.0 ;
      RECT  95250.0 303750.0 96150.0 302850.0 ;
      RECT  90300.0 296550.0 99900.0 295650.0 ;
      RECT  90300.0 310350.0 99900.0 309450.0 ;
      RECT  96900.0 321750.0 98100.0 323700.0 ;
      RECT  96900.0 309900.0 98100.0 311850.0 ;
      RECT  92100.0 311250.0 93300.0 309450.0 ;
      RECT  92100.0 320550.0 93300.0 324150.0 ;
      RECT  94800.0 311250.0 95700.0 320550.0 ;
      RECT  92100.0 320550.0 93300.0 321750.0 ;
      RECT  94500.0 320550.0 95700.0 321750.0 ;
      RECT  94500.0 320550.0 95700.0 321750.0 ;
      RECT  92100.0 320550.0 93300.0 321750.0 ;
      RECT  92100.0 311250.0 93300.0 312450.0 ;
      RECT  94500.0 311250.0 95700.0 312450.0 ;
      RECT  94500.0 311250.0 95700.0 312450.0 ;
      RECT  92100.0 311250.0 93300.0 312450.0 ;
      RECT  96900.0 321150.0 98100.0 322350.0 ;
      RECT  96900.0 311250.0 98100.0 312450.0 ;
      RECT  92700.0 315900.0 93900.0 317100.0 ;
      RECT  92700.0 315900.0 93900.0 317100.0 ;
      RECT  95250.0 316050.0 96150.0 316950.0 ;
      RECT  90300.0 323250.0 99900.0 324150.0 ;
      RECT  90300.0 309450.0 99900.0 310350.0 ;
      RECT  96900.0 325650.0 98100.0 323700.0 ;
      RECT  96900.0 337500.0 98100.0 335550.0 ;
      RECT  92100.0 336150.0 93300.0 337950.0 ;
      RECT  92100.0 326850.0 93300.0 323250.0 ;
      RECT  94800.0 336150.0 95700.0 326850.0 ;
      RECT  92100.0 326850.0 93300.0 325650.0 ;
      RECT  94500.0 326850.0 95700.0 325650.0 ;
      RECT  94500.0 326850.0 95700.0 325650.0 ;
      RECT  92100.0 326850.0 93300.0 325650.0 ;
      RECT  92100.0 336150.0 93300.0 334950.0 ;
      RECT  94500.0 336150.0 95700.0 334950.0 ;
      RECT  94500.0 336150.0 95700.0 334950.0 ;
      RECT  92100.0 336150.0 93300.0 334950.0 ;
      RECT  96900.0 326250.0 98100.0 325050.0 ;
      RECT  96900.0 336150.0 98100.0 334950.0 ;
      RECT  92700.0 331500.0 93900.0 330300.0 ;
      RECT  92700.0 331500.0 93900.0 330300.0 ;
      RECT  95250.0 331350.0 96150.0 330450.0 ;
      RECT  90300.0 324150.0 99900.0 323250.0 ;
      RECT  90300.0 337950.0 99900.0 337050.0 ;
      RECT  96900.0 349350.0 98100.0 351300.0 ;
      RECT  96900.0 337500.0 98100.0 339450.0 ;
      RECT  92100.0 338850.0 93300.0 337050.0 ;
      RECT  92100.0 348150.0 93300.0 351750.0 ;
      RECT  94800.0 338850.0 95700.0 348150.0 ;
      RECT  92100.0 348150.0 93300.0 349350.0 ;
      RECT  94500.0 348150.0 95700.0 349350.0 ;
      RECT  94500.0 348150.0 95700.0 349350.0 ;
      RECT  92100.0 348150.0 93300.0 349350.0 ;
      RECT  92100.0 338850.0 93300.0 340050.0 ;
      RECT  94500.0 338850.0 95700.0 340050.0 ;
      RECT  94500.0 338850.0 95700.0 340050.0 ;
      RECT  92100.0 338850.0 93300.0 340050.0 ;
      RECT  96900.0 348750.0 98100.0 349950.0 ;
      RECT  96900.0 338850.0 98100.0 340050.0 ;
      RECT  92700.0 343500.0 93900.0 344700.0 ;
      RECT  92700.0 343500.0 93900.0 344700.0 ;
      RECT  95250.0 343650.0 96150.0 344550.0 ;
      RECT  90300.0 350850.0 99900.0 351750.0 ;
      RECT  90300.0 337050.0 99900.0 337950.0 ;
      RECT  96900.0 353250.0 98100.0 351300.0 ;
      RECT  96900.0 365100.0 98100.0 363150.0 ;
      RECT  92100.0 363750.0 93300.0 365550.0 ;
      RECT  92100.0 354450.0 93300.0 350850.0 ;
      RECT  94800.0 363750.0 95700.0 354450.0 ;
      RECT  92100.0 354450.0 93300.0 353250.0 ;
      RECT  94500.0 354450.0 95700.0 353250.0 ;
      RECT  94500.0 354450.0 95700.0 353250.0 ;
      RECT  92100.0 354450.0 93300.0 353250.0 ;
      RECT  92100.0 363750.0 93300.0 362550.0 ;
      RECT  94500.0 363750.0 95700.0 362550.0 ;
      RECT  94500.0 363750.0 95700.0 362550.0 ;
      RECT  92100.0 363750.0 93300.0 362550.0 ;
      RECT  96900.0 353850.0 98100.0 352650.0 ;
      RECT  96900.0 363750.0 98100.0 362550.0 ;
      RECT  92700.0 359100.0 93900.0 357900.0 ;
      RECT  92700.0 359100.0 93900.0 357900.0 ;
      RECT  95250.0 358950.0 96150.0 358050.0 ;
      RECT  90300.0 351750.0 99900.0 350850.0 ;
      RECT  90300.0 365550.0 99900.0 364650.0 ;
      RECT  96900.0 376950.0 98100.0 378900.0 ;
      RECT  96900.0 365100.0 98100.0 367050.0 ;
      RECT  92100.0 366450.0 93300.0 364650.0 ;
      RECT  92100.0 375750.0 93300.0 379350.0 ;
      RECT  94800.0 366450.0 95700.0 375750.0 ;
      RECT  92100.0 375750.0 93300.0 376950.0 ;
      RECT  94500.0 375750.0 95700.0 376950.0 ;
      RECT  94500.0 375750.0 95700.0 376950.0 ;
      RECT  92100.0 375750.0 93300.0 376950.0 ;
      RECT  92100.0 366450.0 93300.0 367650.0 ;
      RECT  94500.0 366450.0 95700.0 367650.0 ;
      RECT  94500.0 366450.0 95700.0 367650.0 ;
      RECT  92100.0 366450.0 93300.0 367650.0 ;
      RECT  96900.0 376350.0 98100.0 377550.0 ;
      RECT  96900.0 366450.0 98100.0 367650.0 ;
      RECT  92700.0 371100.0 93900.0 372300.0 ;
      RECT  92700.0 371100.0 93900.0 372300.0 ;
      RECT  95250.0 371250.0 96150.0 372150.0 ;
      RECT  90300.0 378450.0 99900.0 379350.0 ;
      RECT  90300.0 364650.0 99900.0 365550.0 ;
      RECT  96900.0 380850.0 98100.0 378900.0 ;
      RECT  96900.0 392700.0 98100.0 390750.0 ;
      RECT  92100.0 391350.0 93300.0 393150.0 ;
      RECT  92100.0 382050.0 93300.0 378450.0 ;
      RECT  94800.0 391350.0 95700.0 382050.0 ;
      RECT  92100.0 382050.0 93300.0 380850.0 ;
      RECT  94500.0 382050.0 95700.0 380850.0 ;
      RECT  94500.0 382050.0 95700.0 380850.0 ;
      RECT  92100.0 382050.0 93300.0 380850.0 ;
      RECT  92100.0 391350.0 93300.0 390150.0 ;
      RECT  94500.0 391350.0 95700.0 390150.0 ;
      RECT  94500.0 391350.0 95700.0 390150.0 ;
      RECT  92100.0 391350.0 93300.0 390150.0 ;
      RECT  96900.0 381450.0 98100.0 380250.0 ;
      RECT  96900.0 391350.0 98100.0 390150.0 ;
      RECT  92700.0 386700.0 93900.0 385500.0 ;
      RECT  92700.0 386700.0 93900.0 385500.0 ;
      RECT  95250.0 386550.0 96150.0 385650.0 ;
      RECT  90300.0 379350.0 99900.0 378450.0 ;
      RECT  90300.0 393150.0 99900.0 392250.0 ;
      RECT  96900.0 404550.0 98100.0 406500.0 ;
      RECT  96900.0 392700.0 98100.0 394650.0 ;
      RECT  92100.0 394050.0 93300.0 392250.0 ;
      RECT  92100.0 403350.0 93300.0 406950.0 ;
      RECT  94800.0 394050.0 95700.0 403350.0 ;
      RECT  92100.0 403350.0 93300.0 404550.0 ;
      RECT  94500.0 403350.0 95700.0 404550.0 ;
      RECT  94500.0 403350.0 95700.0 404550.0 ;
      RECT  92100.0 403350.0 93300.0 404550.0 ;
      RECT  92100.0 394050.0 93300.0 395250.0 ;
      RECT  94500.0 394050.0 95700.0 395250.0 ;
      RECT  94500.0 394050.0 95700.0 395250.0 ;
      RECT  92100.0 394050.0 93300.0 395250.0 ;
      RECT  96900.0 403950.0 98100.0 405150.0 ;
      RECT  96900.0 394050.0 98100.0 395250.0 ;
      RECT  92700.0 398700.0 93900.0 399900.0 ;
      RECT  92700.0 398700.0 93900.0 399900.0 ;
      RECT  95250.0 398850.0 96150.0 399750.0 ;
      RECT  90300.0 406050.0 99900.0 406950.0 ;
      RECT  90300.0 392250.0 99900.0 393150.0 ;
      RECT  96900.0 408450.0 98100.0 406500.0 ;
      RECT  96900.0 420300.0 98100.0 418350.0 ;
      RECT  92100.0 418950.0 93300.0 420750.0 ;
      RECT  92100.0 409650.0 93300.0 406050.0 ;
      RECT  94800.0 418950.0 95700.0 409650.0 ;
      RECT  92100.0 409650.0 93300.0 408450.0 ;
      RECT  94500.0 409650.0 95700.0 408450.0 ;
      RECT  94500.0 409650.0 95700.0 408450.0 ;
      RECT  92100.0 409650.0 93300.0 408450.0 ;
      RECT  92100.0 418950.0 93300.0 417750.0 ;
      RECT  94500.0 418950.0 95700.0 417750.0 ;
      RECT  94500.0 418950.0 95700.0 417750.0 ;
      RECT  92100.0 418950.0 93300.0 417750.0 ;
      RECT  96900.0 409050.0 98100.0 407850.0 ;
      RECT  96900.0 418950.0 98100.0 417750.0 ;
      RECT  92700.0 414300.0 93900.0 413100.0 ;
      RECT  92700.0 414300.0 93900.0 413100.0 ;
      RECT  95250.0 414150.0 96150.0 413250.0 ;
      RECT  90300.0 406950.0 99900.0 406050.0 ;
      RECT  90300.0 420750.0 99900.0 419850.0 ;
      RECT  60150.0 95100.0 58950.0 96300.0 ;
      RECT  62250.0 109500.0 61050.0 110700.0 ;
      RECT  64350.0 122700.0 63150.0 123900.0 ;
      RECT  66450.0 137100.0 65250.0 138300.0 ;
      RECT  68550.0 150300.0 67350.0 151500.0 ;
      RECT  70650.0 164700.0 69450.0 165900.0 ;
      RECT  72750.0 177900.0 71550.0 179100.0 ;
      RECT  74850.0 192300.0 73650.0 193500.0 ;
      RECT  60150.0 206700.0 58950.0 207900.0 ;
      RECT  68550.0 204000.0 67350.0 205200.0 ;
      RECT  60150.0 218700.0 58950.0 219900.0 ;
      RECT  70650.0 221400.0 69450.0 222600.0 ;
      RECT  60150.0 234300.0 58950.0 235500.0 ;
      RECT  72750.0 231600.0 71550.0 232800.0 ;
      RECT  60150.0 246300.0 58950.0 247500.0 ;
      RECT  74850.0 249000.0 73650.0 250200.0 ;
      RECT  62250.0 261900.0 61050.0 263100.0 ;
      RECT  68550.0 259200.0 67350.0 260400.0 ;
      RECT  62250.0 273900.0 61050.0 275100.0 ;
      RECT  70650.0 276600.0 69450.0 277800.0 ;
      RECT  62250.0 289500.0 61050.0 290700.0 ;
      RECT  72750.0 286800.0 71550.0 288000.0 ;
      RECT  62250.0 301500.0 61050.0 302700.0 ;
      RECT  74850.0 304200.0 73650.0 305400.0 ;
      RECT  64350.0 317100.0 63150.0 318300.0 ;
      RECT  68550.0 314400.0 67350.0 315600.0 ;
      RECT  64350.0 329100.0 63150.0 330300.0 ;
      RECT  70650.0 331800.0 69450.0 333000.0 ;
      RECT  64350.0 344700.0 63150.0 345900.0 ;
      RECT  72750.0 342000.0 71550.0 343200.0 ;
      RECT  64350.0 356700.0 63150.0 357900.0 ;
      RECT  74850.0 359400.0 73650.0 360600.0 ;
      RECT  66450.0 372300.0 65250.0 373500.0 ;
      RECT  68550.0 369600.0 67350.0 370800.0 ;
      RECT  66450.0 384300.0 65250.0 385500.0 ;
      RECT  70650.0 387000.0 69450.0 388200.0 ;
      RECT  66450.0 399900.0 65250.0 401100.0 ;
      RECT  72750.0 397200.0 71550.0 398400.0 ;
      RECT  66450.0 411900.0 65250.0 413100.0 ;
      RECT  74850.0 414600.0 73650.0 415800.0 ;
      RECT  95250.0 205650.0 96150.0 206550.0 ;
      RECT  95250.0 220050.0 96150.0 220950.0 ;
      RECT  95250.0 233250.0 96150.0 234150.0 ;
      RECT  95250.0 247650.0 96150.0 248550.0 ;
      RECT  95250.0 260850.0 96150.0 261750.0 ;
      RECT  95250.0 275250.0 96150.0 276150.0 ;
      RECT  95250.0 288450.0 96150.0 289350.0 ;
      RECT  95250.0 302850.0 96150.0 303750.0 ;
      RECT  95250.0 316050.0 96150.0 316950.0 ;
      RECT  95250.0 330450.0 96150.0 331350.0 ;
      RECT  95250.0 343650.0 96150.0 344550.0 ;
      RECT  95250.0 358050.0 96150.0 358950.0 ;
      RECT  95250.0 371250.0 96150.0 372150.0 ;
      RECT  95250.0 385650.0 96150.0 386550.0 ;
      RECT  95250.0 398850.0 96150.0 399750.0 ;
      RECT  95250.0 413250.0 96150.0 414150.0 ;
      RECT  59100.0 102450.0 130500.0 103350.0 ;
      RECT  59100.0 130050.0 130500.0 130950.0 ;
      RECT  59100.0 157650.0 130500.0 158550.0 ;
      RECT  59100.0 185250.0 130500.0 186150.0 ;
      RECT  59100.0 212850.0 130500.0 213750.0 ;
      RECT  59100.0 240450.0 130500.0 241350.0 ;
      RECT  59100.0 268050.0 130500.0 268950.0 ;
      RECT  59100.0 295650.0 130500.0 296550.0 ;
      RECT  59100.0 323250.0 130500.0 324150.0 ;
      RECT  59100.0 350850.0 130500.0 351750.0 ;
      RECT  59100.0 378450.0 130500.0 379350.0 ;
      RECT  59100.0 406050.0 130500.0 406950.0 ;
      RECT  59100.0 88650.0 130500.0 89550.0 ;
      RECT  59100.0 116250.0 130500.0 117150.0 ;
      RECT  59100.0 143850.0 130500.0 144750.0 ;
      RECT  59100.0 171450.0 130500.0 172350.0 ;
      RECT  59100.0 199050.0 130500.0 199950.0 ;
      RECT  59100.0 226650.0 130500.0 227550.0 ;
      RECT  59100.0 254250.0 130500.0 255150.0 ;
      RECT  59100.0 281850.0 130500.0 282750.0 ;
      RECT  59100.0 309450.0 130500.0 310350.0 ;
      RECT  59100.0 337050.0 130500.0 337950.0 ;
      RECT  59100.0 364650.0 130500.0 365550.0 ;
      RECT  59100.0 392250.0 130500.0 393150.0 ;
      RECT  59100.0 419850.0 130500.0 420750.0 ;
      RECT  103050.0 205650.0 108600.0 206550.0 ;
      RECT  111150.0 206850.0 112050.0 207750.0 ;
      RECT  111150.0 205650.0 112050.0 206550.0 ;
      RECT  111150.0 206550.0 112050.0 207300.0 ;
      RECT  111600.0 206850.0 118200.0 207750.0 ;
      RECT  118200.0 206850.0 119400.0 207750.0 ;
      RECT  127650.0 206850.0 128550.0 207750.0 ;
      RECT  127650.0 205650.0 128550.0 206550.0 ;
      RECT  123600.0 206850.0 128100.0 207750.0 ;
      RECT  127650.0 206100.0 128550.0 207300.0 ;
      RECT  128100.0 205650.0 132600.0 206550.0 ;
      RECT  103050.0 220050.0 108600.0 220950.0 ;
      RECT  111150.0 218850.0 112050.0 219750.0 ;
      RECT  111150.0 220050.0 112050.0 220950.0 ;
      RECT  111150.0 219300.0 112050.0 220950.0 ;
      RECT  111600.0 218850.0 118200.0 219750.0 ;
      RECT  118200.0 218850.0 119400.0 219750.0 ;
      RECT  127650.0 218850.0 128550.0 219750.0 ;
      RECT  127650.0 220050.0 128550.0 220950.0 ;
      RECT  123600.0 218850.0 128100.0 219750.0 ;
      RECT  127650.0 219300.0 128550.0 220500.0 ;
      RECT  128100.0 220050.0 132600.0 220950.0 ;
      RECT  103050.0 233250.0 108600.0 234150.0 ;
      RECT  111150.0 234450.0 112050.0 235350.0 ;
      RECT  111150.0 233250.0 112050.0 234150.0 ;
      RECT  111150.0 234150.0 112050.0 234900.0 ;
      RECT  111600.0 234450.0 118200.0 235350.0 ;
      RECT  118200.0 234450.0 119400.0 235350.0 ;
      RECT  127650.0 234450.0 128550.0 235350.0 ;
      RECT  127650.0 233250.0 128550.0 234150.0 ;
      RECT  123600.0 234450.0 128100.0 235350.0 ;
      RECT  127650.0 233700.0 128550.0 234900.0 ;
      RECT  128100.0 233250.0 132600.0 234150.0 ;
      RECT  103050.0 247650.0 108600.0 248550.0 ;
      RECT  111150.0 246450.0 112050.0 247350.0 ;
      RECT  111150.0 247650.0 112050.0 248550.0 ;
      RECT  111150.0 246900.0 112050.0 248550.0 ;
      RECT  111600.0 246450.0 118200.0 247350.0 ;
      RECT  118200.0 246450.0 119400.0 247350.0 ;
      RECT  127650.0 246450.0 128550.0 247350.0 ;
      RECT  127650.0 247650.0 128550.0 248550.0 ;
      RECT  123600.0 246450.0 128100.0 247350.0 ;
      RECT  127650.0 246900.0 128550.0 248100.0 ;
      RECT  128100.0 247650.0 132600.0 248550.0 ;
      RECT  103050.0 260850.0 108600.0 261750.0 ;
      RECT  111150.0 262050.0 112050.0 262950.0 ;
      RECT  111150.0 260850.0 112050.0 261750.0 ;
      RECT  111150.0 261750.0 112050.0 262500.0 ;
      RECT  111600.0 262050.0 118200.0 262950.0 ;
      RECT  118200.0 262050.0 119400.0 262950.0 ;
      RECT  127650.0 262050.0 128550.0 262950.0 ;
      RECT  127650.0 260850.0 128550.0 261750.0 ;
      RECT  123600.0 262050.0 128100.0 262950.0 ;
      RECT  127650.0 261300.0 128550.0 262500.0 ;
      RECT  128100.0 260850.0 132600.0 261750.0 ;
      RECT  103050.0 275250.0 108600.0 276150.0 ;
      RECT  111150.0 274050.0 112050.0 274950.0 ;
      RECT  111150.0 275250.0 112050.0 276150.0 ;
      RECT  111150.0 274500.0 112050.0 276150.0 ;
      RECT  111600.0 274050.0 118200.0 274950.0 ;
      RECT  118200.0 274050.0 119400.0 274950.0 ;
      RECT  127650.0 274050.0 128550.0 274950.0 ;
      RECT  127650.0 275250.0 128550.0 276150.0 ;
      RECT  123600.0 274050.0 128100.0 274950.0 ;
      RECT  127650.0 274500.0 128550.0 275700.0 ;
      RECT  128100.0 275250.0 132600.0 276150.0 ;
      RECT  103050.0 288450.0 108600.0 289350.0 ;
      RECT  111150.0 289650.0 112050.0 290550.0 ;
      RECT  111150.0 288450.0 112050.0 289350.0 ;
      RECT  111150.0 289350.0 112050.0 290100.0 ;
      RECT  111600.0 289650.0 118200.0 290550.0 ;
      RECT  118200.0 289650.0 119400.0 290550.0 ;
      RECT  127650.0 289650.0 128550.0 290550.0 ;
      RECT  127650.0 288450.0 128550.0 289350.0 ;
      RECT  123600.0 289650.0 128100.0 290550.0 ;
      RECT  127650.0 288900.0 128550.0 290100.0 ;
      RECT  128100.0 288450.0 132600.0 289350.0 ;
      RECT  103050.0 302850.0 108600.0 303750.0 ;
      RECT  111150.0 301650.0 112050.0 302550.0 ;
      RECT  111150.0 302850.0 112050.0 303750.0 ;
      RECT  111150.0 302100.0 112050.0 303750.0 ;
      RECT  111600.0 301650.0 118200.0 302550.0 ;
      RECT  118200.0 301650.0 119400.0 302550.0 ;
      RECT  127650.0 301650.0 128550.0 302550.0 ;
      RECT  127650.0 302850.0 128550.0 303750.0 ;
      RECT  123600.0 301650.0 128100.0 302550.0 ;
      RECT  127650.0 302100.0 128550.0 303300.0 ;
      RECT  128100.0 302850.0 132600.0 303750.0 ;
      RECT  103050.0 316050.0 108600.0 316950.0 ;
      RECT  111150.0 317250.0 112050.0 318150.0 ;
      RECT  111150.0 316050.0 112050.0 316950.0 ;
      RECT  111150.0 316950.0 112050.0 317700.0 ;
      RECT  111600.0 317250.0 118200.0 318150.0 ;
      RECT  118200.0 317250.0 119400.0 318150.0 ;
      RECT  127650.0 317250.0 128550.0 318150.0 ;
      RECT  127650.0 316050.0 128550.0 316950.0 ;
      RECT  123600.0 317250.0 128100.0 318150.0 ;
      RECT  127650.0 316500.0 128550.0 317700.0 ;
      RECT  128100.0 316050.0 132600.0 316950.0 ;
      RECT  103050.0 330450.0 108600.0 331350.0 ;
      RECT  111150.0 329250.0 112050.0 330150.0 ;
      RECT  111150.0 330450.0 112050.0 331350.0 ;
      RECT  111150.0 329700.0 112050.0 331350.0 ;
      RECT  111600.0 329250.0 118200.0 330150.0 ;
      RECT  118200.0 329250.0 119400.0 330150.0 ;
      RECT  127650.0 329250.0 128550.0 330150.0 ;
      RECT  127650.0 330450.0 128550.0 331350.0 ;
      RECT  123600.0 329250.0 128100.0 330150.0 ;
      RECT  127650.0 329700.0 128550.0 330900.0 ;
      RECT  128100.0 330450.0 132600.0 331350.0 ;
      RECT  103050.0 343650.0 108600.0 344550.0 ;
      RECT  111150.0 344850.0 112050.0 345750.0 ;
      RECT  111150.0 343650.0 112050.0 344550.0 ;
      RECT  111150.0 344550.0 112050.0 345300.0 ;
      RECT  111600.0 344850.0 118200.0 345750.0 ;
      RECT  118200.0 344850.0 119400.0 345750.0 ;
      RECT  127650.0 344850.0 128550.0 345750.0 ;
      RECT  127650.0 343650.0 128550.0 344550.0 ;
      RECT  123600.0 344850.0 128100.0 345750.0 ;
      RECT  127650.0 344100.0 128550.0 345300.0 ;
      RECT  128100.0 343650.0 132600.0 344550.0 ;
      RECT  103050.0 358050.0 108600.0 358950.0 ;
      RECT  111150.0 356850.0 112050.0 357750.0 ;
      RECT  111150.0 358050.0 112050.0 358950.0 ;
      RECT  111150.0 357300.0 112050.0 358950.0 ;
      RECT  111600.0 356850.0 118200.0 357750.0 ;
      RECT  118200.0 356850.0 119400.0 357750.0 ;
      RECT  127650.0 356850.0 128550.0 357750.0 ;
      RECT  127650.0 358050.0 128550.0 358950.0 ;
      RECT  123600.0 356850.0 128100.0 357750.0 ;
      RECT  127650.0 357300.0 128550.0 358500.0 ;
      RECT  128100.0 358050.0 132600.0 358950.0 ;
      RECT  103050.0 371250.0 108600.0 372150.0 ;
      RECT  111150.0 372450.0 112050.0 373350.0 ;
      RECT  111150.0 371250.0 112050.0 372150.0 ;
      RECT  111150.0 372150.0 112050.0 372900.0 ;
      RECT  111600.0 372450.0 118200.0 373350.0 ;
      RECT  118200.0 372450.0 119400.0 373350.0 ;
      RECT  127650.0 372450.0 128550.0 373350.0 ;
      RECT  127650.0 371250.0 128550.0 372150.0 ;
      RECT  123600.0 372450.0 128100.0 373350.0 ;
      RECT  127650.0 371700.0 128550.0 372900.0 ;
      RECT  128100.0 371250.0 132600.0 372150.0 ;
      RECT  103050.0 385650.0 108600.0 386550.0 ;
      RECT  111150.0 384450.0 112050.0 385350.0 ;
      RECT  111150.0 385650.0 112050.0 386550.0 ;
      RECT  111150.0 384900.0 112050.0 386550.0 ;
      RECT  111600.0 384450.0 118200.0 385350.0 ;
      RECT  118200.0 384450.0 119400.0 385350.0 ;
      RECT  127650.0 384450.0 128550.0 385350.0 ;
      RECT  127650.0 385650.0 128550.0 386550.0 ;
      RECT  123600.0 384450.0 128100.0 385350.0 ;
      RECT  127650.0 384900.0 128550.0 386100.0 ;
      RECT  128100.0 385650.0 132600.0 386550.0 ;
      RECT  103050.0 398850.0 108600.0 399750.0 ;
      RECT  111150.0 400050.0 112050.0 400950.0 ;
      RECT  111150.0 398850.0 112050.0 399750.0 ;
      RECT  111150.0 399750.0 112050.0 400500.0 ;
      RECT  111600.0 400050.0 118200.0 400950.0 ;
      RECT  118200.0 400050.0 119400.0 400950.0 ;
      RECT  127650.0 400050.0 128550.0 400950.0 ;
      RECT  127650.0 398850.0 128550.0 399750.0 ;
      RECT  123600.0 400050.0 128100.0 400950.0 ;
      RECT  127650.0 399300.0 128550.0 400500.0 ;
      RECT  128100.0 398850.0 132600.0 399750.0 ;
      RECT  103050.0 413250.0 108600.0 414150.0 ;
      RECT  111150.0 412050.0 112050.0 412950.0 ;
      RECT  111150.0 413250.0 112050.0 414150.0 ;
      RECT  111150.0 412500.0 112050.0 414150.0 ;
      RECT  111600.0 412050.0 118200.0 412950.0 ;
      RECT  118200.0 412050.0 119400.0 412950.0 ;
      RECT  127650.0 412050.0 128550.0 412950.0 ;
      RECT  127650.0 413250.0 128550.0 414150.0 ;
      RECT  123600.0 412050.0 128100.0 412950.0 ;
      RECT  127650.0 412500.0 128550.0 413700.0 ;
      RECT  128100.0 413250.0 132600.0 414150.0 ;
      RECT  112800.0 211350.0 114000.0 213300.0 ;
      RECT  112800.0 199500.0 114000.0 201450.0 ;
      RECT  108000.0 200850.0 109200.0 199050.0 ;
      RECT  108000.0 210150.0 109200.0 213750.0 ;
      RECT  110700.0 200850.0 111600.0 210150.0 ;
      RECT  108000.0 210150.0 109200.0 211350.0 ;
      RECT  110400.0 210150.0 111600.0 211350.0 ;
      RECT  110400.0 210150.0 111600.0 211350.0 ;
      RECT  108000.0 210150.0 109200.0 211350.0 ;
      RECT  108000.0 200850.0 109200.0 202050.0 ;
      RECT  110400.0 200850.0 111600.0 202050.0 ;
      RECT  110400.0 200850.0 111600.0 202050.0 ;
      RECT  108000.0 200850.0 109200.0 202050.0 ;
      RECT  112800.0 210750.0 114000.0 211950.0 ;
      RECT  112800.0 200850.0 114000.0 202050.0 ;
      RECT  108600.0 205500.0 109800.0 206700.0 ;
      RECT  108600.0 205500.0 109800.0 206700.0 ;
      RECT  111150.0 205650.0 112050.0 206550.0 ;
      RECT  106200.0 212850.0 115800.0 213750.0 ;
      RECT  106200.0 199050.0 115800.0 199950.0 ;
      RECT  117600.0 201450.0 118800.0 199050.0 ;
      RECT  117600.0 210150.0 118800.0 213750.0 ;
      RECT  122400.0 210150.0 123600.0 213750.0 ;
      RECT  124800.0 211350.0 126000.0 213300.0 ;
      RECT  124800.0 199500.0 126000.0 201450.0 ;
      RECT  117600.0 210150.0 118800.0 211350.0 ;
      RECT  120000.0 210150.0 121200.0 211350.0 ;
      RECT  120000.0 210150.0 121200.0 211350.0 ;
      RECT  117600.0 210150.0 118800.0 211350.0 ;
      RECT  120000.0 210150.0 121200.0 211350.0 ;
      RECT  122400.0 210150.0 123600.0 211350.0 ;
      RECT  122400.0 210150.0 123600.0 211350.0 ;
      RECT  120000.0 210150.0 121200.0 211350.0 ;
      RECT  117600.0 201450.0 118800.0 202650.0 ;
      RECT  120000.0 201450.0 121200.0 202650.0 ;
      RECT  120000.0 201450.0 121200.0 202650.0 ;
      RECT  117600.0 201450.0 118800.0 202650.0 ;
      RECT  120000.0 201450.0 121200.0 202650.0 ;
      RECT  122400.0 201450.0 123600.0 202650.0 ;
      RECT  122400.0 201450.0 123600.0 202650.0 ;
      RECT  120000.0 201450.0 121200.0 202650.0 ;
      RECT  124800.0 210750.0 126000.0 211950.0 ;
      RECT  124800.0 200850.0 126000.0 202050.0 ;
      RECT  122400.0 204000.0 121200.0 205200.0 ;
      RECT  119400.0 206700.0 118200.0 207900.0 ;
      RECT  120000.0 210150.0 121200.0 211350.0 ;
      RECT  122400.0 201450.0 123600.0 202650.0 ;
      RECT  123600.0 206700.0 122400.0 207900.0 ;
      RECT  118200.0 206700.0 119400.0 207900.0 ;
      RECT  121200.0 204000.0 122400.0 205200.0 ;
      RECT  122400.0 206700.0 123600.0 207900.0 ;
      RECT  115800.0 212850.0 130200.0 213750.0 ;
      RECT  115800.0 199050.0 130200.0 199950.0 ;
      RECT  136800.0 211350.0 138000.0 213300.0 ;
      RECT  136800.0 199500.0 138000.0 201450.0 ;
      RECT  132000.0 200850.0 133200.0 199050.0 ;
      RECT  132000.0 210150.0 133200.0 213750.0 ;
      RECT  134700.0 200850.0 135600.0 210150.0 ;
      RECT  132000.0 210150.0 133200.0 211350.0 ;
      RECT  134400.0 210150.0 135600.0 211350.0 ;
      RECT  134400.0 210150.0 135600.0 211350.0 ;
      RECT  132000.0 210150.0 133200.0 211350.0 ;
      RECT  132000.0 200850.0 133200.0 202050.0 ;
      RECT  134400.0 200850.0 135600.0 202050.0 ;
      RECT  134400.0 200850.0 135600.0 202050.0 ;
      RECT  132000.0 200850.0 133200.0 202050.0 ;
      RECT  136800.0 210750.0 138000.0 211950.0 ;
      RECT  136800.0 200850.0 138000.0 202050.0 ;
      RECT  132600.0 205500.0 133800.0 206700.0 ;
      RECT  132600.0 205500.0 133800.0 206700.0 ;
      RECT  135150.0 205650.0 136050.0 206550.0 ;
      RECT  130200.0 212850.0 139800.0 213750.0 ;
      RECT  130200.0 199050.0 139800.0 199950.0 ;
      RECT  102450.0 205500.0 103650.0 206700.0 ;
      RECT  104400.0 203100.0 105600.0 204300.0 ;
      RECT  121200.0 204000.0 120000.0 205200.0 ;
      RECT  112800.0 215250.0 114000.0 213300.0 ;
      RECT  112800.0 227100.0 114000.0 225150.0 ;
      RECT  108000.0 225750.0 109200.0 227550.0 ;
      RECT  108000.0 216450.0 109200.0 212850.0 ;
      RECT  110700.0 225750.0 111600.0 216450.0 ;
      RECT  108000.0 216450.0 109200.0 215250.0 ;
      RECT  110400.0 216450.0 111600.0 215250.0 ;
      RECT  110400.0 216450.0 111600.0 215250.0 ;
      RECT  108000.0 216450.0 109200.0 215250.0 ;
      RECT  108000.0 225750.0 109200.0 224550.0 ;
      RECT  110400.0 225750.0 111600.0 224550.0 ;
      RECT  110400.0 225750.0 111600.0 224550.0 ;
      RECT  108000.0 225750.0 109200.0 224550.0 ;
      RECT  112800.0 215850.0 114000.0 214650.0 ;
      RECT  112800.0 225750.0 114000.0 224550.0 ;
      RECT  108600.0 221100.0 109800.0 219900.0 ;
      RECT  108600.0 221100.0 109800.0 219900.0 ;
      RECT  111150.0 220950.0 112050.0 220050.0 ;
      RECT  106200.0 213750.0 115800.0 212850.0 ;
      RECT  106200.0 227550.0 115800.0 226650.0 ;
      RECT  117600.0 225150.0 118800.0 227550.0 ;
      RECT  117600.0 216450.0 118800.0 212850.0 ;
      RECT  122400.0 216450.0 123600.0 212850.0 ;
      RECT  124800.0 215250.0 126000.0 213300.0 ;
      RECT  124800.0 227100.0 126000.0 225150.0 ;
      RECT  117600.0 216450.0 118800.0 215250.0 ;
      RECT  120000.0 216450.0 121200.0 215250.0 ;
      RECT  120000.0 216450.0 121200.0 215250.0 ;
      RECT  117600.0 216450.0 118800.0 215250.0 ;
      RECT  120000.0 216450.0 121200.0 215250.0 ;
      RECT  122400.0 216450.0 123600.0 215250.0 ;
      RECT  122400.0 216450.0 123600.0 215250.0 ;
      RECT  120000.0 216450.0 121200.0 215250.0 ;
      RECT  117600.0 225150.0 118800.0 223950.0 ;
      RECT  120000.0 225150.0 121200.0 223950.0 ;
      RECT  120000.0 225150.0 121200.0 223950.0 ;
      RECT  117600.0 225150.0 118800.0 223950.0 ;
      RECT  120000.0 225150.0 121200.0 223950.0 ;
      RECT  122400.0 225150.0 123600.0 223950.0 ;
      RECT  122400.0 225150.0 123600.0 223950.0 ;
      RECT  120000.0 225150.0 121200.0 223950.0 ;
      RECT  124800.0 215850.0 126000.0 214650.0 ;
      RECT  124800.0 225750.0 126000.0 224550.0 ;
      RECT  122400.0 222600.0 121200.0 221400.0 ;
      RECT  119400.0 219900.0 118200.0 218700.0 ;
      RECT  120000.0 216450.0 121200.0 215250.0 ;
      RECT  122400.0 225150.0 123600.0 223950.0 ;
      RECT  123600.0 219900.0 122400.0 218700.0 ;
      RECT  118200.0 219900.0 119400.0 218700.0 ;
      RECT  121200.0 222600.0 122400.0 221400.0 ;
      RECT  122400.0 219900.0 123600.0 218700.0 ;
      RECT  115800.0 213750.0 130200.0 212850.0 ;
      RECT  115800.0 227550.0 130200.0 226650.0 ;
      RECT  136800.0 215250.0 138000.0 213300.0 ;
      RECT  136800.0 227100.0 138000.0 225150.0 ;
      RECT  132000.0 225750.0 133200.0 227550.0 ;
      RECT  132000.0 216450.0 133200.0 212850.0 ;
      RECT  134700.0 225750.0 135600.0 216450.0 ;
      RECT  132000.0 216450.0 133200.0 215250.0 ;
      RECT  134400.0 216450.0 135600.0 215250.0 ;
      RECT  134400.0 216450.0 135600.0 215250.0 ;
      RECT  132000.0 216450.0 133200.0 215250.0 ;
      RECT  132000.0 225750.0 133200.0 224550.0 ;
      RECT  134400.0 225750.0 135600.0 224550.0 ;
      RECT  134400.0 225750.0 135600.0 224550.0 ;
      RECT  132000.0 225750.0 133200.0 224550.0 ;
      RECT  136800.0 215850.0 138000.0 214650.0 ;
      RECT  136800.0 225750.0 138000.0 224550.0 ;
      RECT  132600.0 221100.0 133800.0 219900.0 ;
      RECT  132600.0 221100.0 133800.0 219900.0 ;
      RECT  135150.0 220950.0 136050.0 220050.0 ;
      RECT  130200.0 213750.0 139800.0 212850.0 ;
      RECT  130200.0 227550.0 139800.0 226650.0 ;
      RECT  102450.0 219900.0 103650.0 221100.0 ;
      RECT  104400.0 222300.0 105600.0 223500.0 ;
      RECT  121200.0 221400.0 120000.0 222600.0 ;
      RECT  112800.0 238950.0 114000.0 240900.0 ;
      RECT  112800.0 227100.0 114000.0 229050.0 ;
      RECT  108000.0 228450.0 109200.0 226650.0 ;
      RECT  108000.0 237750.0 109200.0 241350.0 ;
      RECT  110700.0 228450.0 111600.0 237750.0 ;
      RECT  108000.0 237750.0 109200.0 238950.0 ;
      RECT  110400.0 237750.0 111600.0 238950.0 ;
      RECT  110400.0 237750.0 111600.0 238950.0 ;
      RECT  108000.0 237750.0 109200.0 238950.0 ;
      RECT  108000.0 228450.0 109200.0 229650.0 ;
      RECT  110400.0 228450.0 111600.0 229650.0 ;
      RECT  110400.0 228450.0 111600.0 229650.0 ;
      RECT  108000.0 228450.0 109200.0 229650.0 ;
      RECT  112800.0 238350.0 114000.0 239550.0 ;
      RECT  112800.0 228450.0 114000.0 229650.0 ;
      RECT  108600.0 233100.0 109800.0 234300.0 ;
      RECT  108600.0 233100.0 109800.0 234300.0 ;
      RECT  111150.0 233250.0 112050.0 234150.0 ;
      RECT  106200.0 240450.0 115800.0 241350.0 ;
      RECT  106200.0 226650.0 115800.0 227550.0 ;
      RECT  117600.0 229050.0 118800.0 226650.0 ;
      RECT  117600.0 237750.0 118800.0 241350.0 ;
      RECT  122400.0 237750.0 123600.0 241350.0 ;
      RECT  124800.0 238950.0 126000.0 240900.0 ;
      RECT  124800.0 227100.0 126000.0 229050.0 ;
      RECT  117600.0 237750.0 118800.0 238950.0 ;
      RECT  120000.0 237750.0 121200.0 238950.0 ;
      RECT  120000.0 237750.0 121200.0 238950.0 ;
      RECT  117600.0 237750.0 118800.0 238950.0 ;
      RECT  120000.0 237750.0 121200.0 238950.0 ;
      RECT  122400.0 237750.0 123600.0 238950.0 ;
      RECT  122400.0 237750.0 123600.0 238950.0 ;
      RECT  120000.0 237750.0 121200.0 238950.0 ;
      RECT  117600.0 229050.0 118800.0 230250.0 ;
      RECT  120000.0 229050.0 121200.0 230250.0 ;
      RECT  120000.0 229050.0 121200.0 230250.0 ;
      RECT  117600.0 229050.0 118800.0 230250.0 ;
      RECT  120000.0 229050.0 121200.0 230250.0 ;
      RECT  122400.0 229050.0 123600.0 230250.0 ;
      RECT  122400.0 229050.0 123600.0 230250.0 ;
      RECT  120000.0 229050.0 121200.0 230250.0 ;
      RECT  124800.0 238350.0 126000.0 239550.0 ;
      RECT  124800.0 228450.0 126000.0 229650.0 ;
      RECT  122400.0 231600.0 121200.0 232800.0 ;
      RECT  119400.0 234300.0 118200.0 235500.0 ;
      RECT  120000.0 237750.0 121200.0 238950.0 ;
      RECT  122400.0 229050.0 123600.0 230250.0 ;
      RECT  123600.0 234300.0 122400.0 235500.0 ;
      RECT  118200.0 234300.0 119400.0 235500.0 ;
      RECT  121200.0 231600.0 122400.0 232800.0 ;
      RECT  122400.0 234300.0 123600.0 235500.0 ;
      RECT  115800.0 240450.0 130200.0 241350.0 ;
      RECT  115800.0 226650.0 130200.0 227550.0 ;
      RECT  136800.0 238950.0 138000.0 240900.0 ;
      RECT  136800.0 227100.0 138000.0 229050.0 ;
      RECT  132000.0 228450.0 133200.0 226650.0 ;
      RECT  132000.0 237750.0 133200.0 241350.0 ;
      RECT  134700.0 228450.0 135600.0 237750.0 ;
      RECT  132000.0 237750.0 133200.0 238950.0 ;
      RECT  134400.0 237750.0 135600.0 238950.0 ;
      RECT  134400.0 237750.0 135600.0 238950.0 ;
      RECT  132000.0 237750.0 133200.0 238950.0 ;
      RECT  132000.0 228450.0 133200.0 229650.0 ;
      RECT  134400.0 228450.0 135600.0 229650.0 ;
      RECT  134400.0 228450.0 135600.0 229650.0 ;
      RECT  132000.0 228450.0 133200.0 229650.0 ;
      RECT  136800.0 238350.0 138000.0 239550.0 ;
      RECT  136800.0 228450.0 138000.0 229650.0 ;
      RECT  132600.0 233100.0 133800.0 234300.0 ;
      RECT  132600.0 233100.0 133800.0 234300.0 ;
      RECT  135150.0 233250.0 136050.0 234150.0 ;
      RECT  130200.0 240450.0 139800.0 241350.0 ;
      RECT  130200.0 226650.0 139800.0 227550.0 ;
      RECT  102450.0 233100.0 103650.0 234300.0 ;
      RECT  104400.0 230700.0 105600.0 231900.0 ;
      RECT  121200.0 231600.0 120000.0 232800.0 ;
      RECT  112800.0 242850.0 114000.0 240900.0 ;
      RECT  112800.0 254700.0 114000.0 252750.0 ;
      RECT  108000.0 253350.0 109200.0 255150.0 ;
      RECT  108000.0 244050.0 109200.0 240450.0 ;
      RECT  110700.0 253350.0 111600.0 244050.0 ;
      RECT  108000.0 244050.0 109200.0 242850.0 ;
      RECT  110400.0 244050.0 111600.0 242850.0 ;
      RECT  110400.0 244050.0 111600.0 242850.0 ;
      RECT  108000.0 244050.0 109200.0 242850.0 ;
      RECT  108000.0 253350.0 109200.0 252150.0 ;
      RECT  110400.0 253350.0 111600.0 252150.0 ;
      RECT  110400.0 253350.0 111600.0 252150.0 ;
      RECT  108000.0 253350.0 109200.0 252150.0 ;
      RECT  112800.0 243450.0 114000.0 242250.0 ;
      RECT  112800.0 253350.0 114000.0 252150.0 ;
      RECT  108600.0 248700.0 109800.0 247500.0 ;
      RECT  108600.0 248700.0 109800.0 247500.0 ;
      RECT  111150.0 248550.0 112050.0 247650.0 ;
      RECT  106200.0 241350.0 115800.0 240450.0 ;
      RECT  106200.0 255150.0 115800.0 254250.0 ;
      RECT  117600.0 252750.0 118800.0 255150.0 ;
      RECT  117600.0 244050.0 118800.0 240450.0 ;
      RECT  122400.0 244050.0 123600.0 240450.0 ;
      RECT  124800.0 242850.0 126000.0 240900.0 ;
      RECT  124800.0 254700.0 126000.0 252750.0 ;
      RECT  117600.0 244050.0 118800.0 242850.0 ;
      RECT  120000.0 244050.0 121200.0 242850.0 ;
      RECT  120000.0 244050.0 121200.0 242850.0 ;
      RECT  117600.0 244050.0 118800.0 242850.0 ;
      RECT  120000.0 244050.0 121200.0 242850.0 ;
      RECT  122400.0 244050.0 123600.0 242850.0 ;
      RECT  122400.0 244050.0 123600.0 242850.0 ;
      RECT  120000.0 244050.0 121200.0 242850.0 ;
      RECT  117600.0 252750.0 118800.0 251550.0 ;
      RECT  120000.0 252750.0 121200.0 251550.0 ;
      RECT  120000.0 252750.0 121200.0 251550.0 ;
      RECT  117600.0 252750.0 118800.0 251550.0 ;
      RECT  120000.0 252750.0 121200.0 251550.0 ;
      RECT  122400.0 252750.0 123600.0 251550.0 ;
      RECT  122400.0 252750.0 123600.0 251550.0 ;
      RECT  120000.0 252750.0 121200.0 251550.0 ;
      RECT  124800.0 243450.0 126000.0 242250.0 ;
      RECT  124800.0 253350.0 126000.0 252150.0 ;
      RECT  122400.0 250200.0 121200.0 249000.0 ;
      RECT  119400.0 247500.0 118200.0 246300.0 ;
      RECT  120000.0 244050.0 121200.0 242850.0 ;
      RECT  122400.0 252750.0 123600.0 251550.0 ;
      RECT  123600.0 247500.0 122400.0 246300.0 ;
      RECT  118200.0 247500.0 119400.0 246300.0 ;
      RECT  121200.0 250200.0 122400.0 249000.0 ;
      RECT  122400.0 247500.0 123600.0 246300.0 ;
      RECT  115800.0 241350.0 130200.0 240450.0 ;
      RECT  115800.0 255150.0 130200.0 254250.0 ;
      RECT  136800.0 242850.0 138000.0 240900.0 ;
      RECT  136800.0 254700.0 138000.0 252750.0 ;
      RECT  132000.0 253350.0 133200.0 255150.0 ;
      RECT  132000.0 244050.0 133200.0 240450.0 ;
      RECT  134700.0 253350.0 135600.0 244050.0 ;
      RECT  132000.0 244050.0 133200.0 242850.0 ;
      RECT  134400.0 244050.0 135600.0 242850.0 ;
      RECT  134400.0 244050.0 135600.0 242850.0 ;
      RECT  132000.0 244050.0 133200.0 242850.0 ;
      RECT  132000.0 253350.0 133200.0 252150.0 ;
      RECT  134400.0 253350.0 135600.0 252150.0 ;
      RECT  134400.0 253350.0 135600.0 252150.0 ;
      RECT  132000.0 253350.0 133200.0 252150.0 ;
      RECT  136800.0 243450.0 138000.0 242250.0 ;
      RECT  136800.0 253350.0 138000.0 252150.0 ;
      RECT  132600.0 248700.0 133800.0 247500.0 ;
      RECT  132600.0 248700.0 133800.0 247500.0 ;
      RECT  135150.0 248550.0 136050.0 247650.0 ;
      RECT  130200.0 241350.0 139800.0 240450.0 ;
      RECT  130200.0 255150.0 139800.0 254250.0 ;
      RECT  102450.0 247500.0 103650.0 248700.0 ;
      RECT  104400.0 249900.0 105600.0 251100.0 ;
      RECT  121200.0 249000.0 120000.0 250200.0 ;
      RECT  112800.0 266550.0 114000.0 268500.0 ;
      RECT  112800.0 254700.0 114000.0 256650.0 ;
      RECT  108000.0 256050.0 109200.0 254250.0 ;
      RECT  108000.0 265350.0 109200.0 268950.0 ;
      RECT  110700.0 256050.0 111600.0 265350.0 ;
      RECT  108000.0 265350.0 109200.0 266550.0 ;
      RECT  110400.0 265350.0 111600.0 266550.0 ;
      RECT  110400.0 265350.0 111600.0 266550.0 ;
      RECT  108000.0 265350.0 109200.0 266550.0 ;
      RECT  108000.0 256050.0 109200.0 257250.0 ;
      RECT  110400.0 256050.0 111600.0 257250.0 ;
      RECT  110400.0 256050.0 111600.0 257250.0 ;
      RECT  108000.0 256050.0 109200.0 257250.0 ;
      RECT  112800.0 265950.0 114000.0 267150.0 ;
      RECT  112800.0 256050.0 114000.0 257250.0 ;
      RECT  108600.0 260700.0 109800.0 261900.0 ;
      RECT  108600.0 260700.0 109800.0 261900.0 ;
      RECT  111150.0 260850.0 112050.0 261750.0 ;
      RECT  106200.0 268050.0 115800.0 268950.0 ;
      RECT  106200.0 254250.0 115800.0 255150.0 ;
      RECT  117600.0 256650.0 118800.0 254250.0 ;
      RECT  117600.0 265350.0 118800.0 268950.0 ;
      RECT  122400.0 265350.0 123600.0 268950.0 ;
      RECT  124800.0 266550.0 126000.0 268500.0 ;
      RECT  124800.0 254700.0 126000.0 256650.0 ;
      RECT  117600.0 265350.0 118800.0 266550.0 ;
      RECT  120000.0 265350.0 121200.0 266550.0 ;
      RECT  120000.0 265350.0 121200.0 266550.0 ;
      RECT  117600.0 265350.0 118800.0 266550.0 ;
      RECT  120000.0 265350.0 121200.0 266550.0 ;
      RECT  122400.0 265350.0 123600.0 266550.0 ;
      RECT  122400.0 265350.0 123600.0 266550.0 ;
      RECT  120000.0 265350.0 121200.0 266550.0 ;
      RECT  117600.0 256650.0 118800.0 257850.0 ;
      RECT  120000.0 256650.0 121200.0 257850.0 ;
      RECT  120000.0 256650.0 121200.0 257850.0 ;
      RECT  117600.0 256650.0 118800.0 257850.0 ;
      RECT  120000.0 256650.0 121200.0 257850.0 ;
      RECT  122400.0 256650.0 123600.0 257850.0 ;
      RECT  122400.0 256650.0 123600.0 257850.0 ;
      RECT  120000.0 256650.0 121200.0 257850.0 ;
      RECT  124800.0 265950.0 126000.0 267150.0 ;
      RECT  124800.0 256050.0 126000.0 257250.0 ;
      RECT  122400.0 259200.0 121200.0 260400.0 ;
      RECT  119400.0 261900.0 118200.0 263100.0 ;
      RECT  120000.0 265350.0 121200.0 266550.0 ;
      RECT  122400.0 256650.0 123600.0 257850.0 ;
      RECT  123600.0 261900.0 122400.0 263100.0 ;
      RECT  118200.0 261900.0 119400.0 263100.0 ;
      RECT  121200.0 259200.0 122400.0 260400.0 ;
      RECT  122400.0 261900.0 123600.0 263100.0 ;
      RECT  115800.0 268050.0 130200.0 268950.0 ;
      RECT  115800.0 254250.0 130200.0 255150.0 ;
      RECT  136800.0 266550.0 138000.0 268500.0 ;
      RECT  136800.0 254700.0 138000.0 256650.0 ;
      RECT  132000.0 256050.0 133200.0 254250.0 ;
      RECT  132000.0 265350.0 133200.0 268950.0 ;
      RECT  134700.0 256050.0 135600.0 265350.0 ;
      RECT  132000.0 265350.0 133200.0 266550.0 ;
      RECT  134400.0 265350.0 135600.0 266550.0 ;
      RECT  134400.0 265350.0 135600.0 266550.0 ;
      RECT  132000.0 265350.0 133200.0 266550.0 ;
      RECT  132000.0 256050.0 133200.0 257250.0 ;
      RECT  134400.0 256050.0 135600.0 257250.0 ;
      RECT  134400.0 256050.0 135600.0 257250.0 ;
      RECT  132000.0 256050.0 133200.0 257250.0 ;
      RECT  136800.0 265950.0 138000.0 267150.0 ;
      RECT  136800.0 256050.0 138000.0 257250.0 ;
      RECT  132600.0 260700.0 133800.0 261900.0 ;
      RECT  132600.0 260700.0 133800.0 261900.0 ;
      RECT  135150.0 260850.0 136050.0 261750.0 ;
      RECT  130200.0 268050.0 139800.0 268950.0 ;
      RECT  130200.0 254250.0 139800.0 255150.0 ;
      RECT  102450.0 260700.0 103650.0 261900.0 ;
      RECT  104400.0 258300.0 105600.0 259500.0 ;
      RECT  121200.0 259200.0 120000.0 260400.0 ;
      RECT  112800.0 270450.0 114000.0 268500.0 ;
      RECT  112800.0 282300.0 114000.0 280350.0 ;
      RECT  108000.0 280950.0 109200.0 282750.0 ;
      RECT  108000.0 271650.0 109200.0 268050.0 ;
      RECT  110700.0 280950.0 111600.0 271650.0 ;
      RECT  108000.0 271650.0 109200.0 270450.0 ;
      RECT  110400.0 271650.0 111600.0 270450.0 ;
      RECT  110400.0 271650.0 111600.0 270450.0 ;
      RECT  108000.0 271650.0 109200.0 270450.0 ;
      RECT  108000.0 280950.0 109200.0 279750.0 ;
      RECT  110400.0 280950.0 111600.0 279750.0 ;
      RECT  110400.0 280950.0 111600.0 279750.0 ;
      RECT  108000.0 280950.0 109200.0 279750.0 ;
      RECT  112800.0 271050.0 114000.0 269850.0 ;
      RECT  112800.0 280950.0 114000.0 279750.0 ;
      RECT  108600.0 276300.0 109800.0 275100.0 ;
      RECT  108600.0 276300.0 109800.0 275100.0 ;
      RECT  111150.0 276150.0 112050.0 275250.0 ;
      RECT  106200.0 268950.0 115800.0 268050.0 ;
      RECT  106200.0 282750.0 115800.0 281850.0 ;
      RECT  117600.0 280350.0 118800.0 282750.0 ;
      RECT  117600.0 271650.0 118800.0 268050.0 ;
      RECT  122400.0 271650.0 123600.0 268050.0 ;
      RECT  124800.0 270450.0 126000.0 268500.0 ;
      RECT  124800.0 282300.0 126000.0 280350.0 ;
      RECT  117600.0 271650.0 118800.0 270450.0 ;
      RECT  120000.0 271650.0 121200.0 270450.0 ;
      RECT  120000.0 271650.0 121200.0 270450.0 ;
      RECT  117600.0 271650.0 118800.0 270450.0 ;
      RECT  120000.0 271650.0 121200.0 270450.0 ;
      RECT  122400.0 271650.0 123600.0 270450.0 ;
      RECT  122400.0 271650.0 123600.0 270450.0 ;
      RECT  120000.0 271650.0 121200.0 270450.0 ;
      RECT  117600.0 280350.0 118800.0 279150.0 ;
      RECT  120000.0 280350.0 121200.0 279150.0 ;
      RECT  120000.0 280350.0 121200.0 279150.0 ;
      RECT  117600.0 280350.0 118800.0 279150.0 ;
      RECT  120000.0 280350.0 121200.0 279150.0 ;
      RECT  122400.0 280350.0 123600.0 279150.0 ;
      RECT  122400.0 280350.0 123600.0 279150.0 ;
      RECT  120000.0 280350.0 121200.0 279150.0 ;
      RECT  124800.0 271050.0 126000.0 269850.0 ;
      RECT  124800.0 280950.0 126000.0 279750.0 ;
      RECT  122400.0 277800.0 121200.0 276600.0 ;
      RECT  119400.0 275100.0 118200.0 273900.0 ;
      RECT  120000.0 271650.0 121200.0 270450.0 ;
      RECT  122400.0 280350.0 123600.0 279150.0 ;
      RECT  123600.0 275100.0 122400.0 273900.0 ;
      RECT  118200.0 275100.0 119400.0 273900.0 ;
      RECT  121200.0 277800.0 122400.0 276600.0 ;
      RECT  122400.0 275100.0 123600.0 273900.0 ;
      RECT  115800.0 268950.0 130200.0 268050.0 ;
      RECT  115800.0 282750.0 130200.0 281850.0 ;
      RECT  136800.0 270450.0 138000.0 268500.0 ;
      RECT  136800.0 282300.0 138000.0 280350.0 ;
      RECT  132000.0 280950.0 133200.0 282750.0 ;
      RECT  132000.0 271650.0 133200.0 268050.0 ;
      RECT  134700.0 280950.0 135600.0 271650.0 ;
      RECT  132000.0 271650.0 133200.0 270450.0 ;
      RECT  134400.0 271650.0 135600.0 270450.0 ;
      RECT  134400.0 271650.0 135600.0 270450.0 ;
      RECT  132000.0 271650.0 133200.0 270450.0 ;
      RECT  132000.0 280950.0 133200.0 279750.0 ;
      RECT  134400.0 280950.0 135600.0 279750.0 ;
      RECT  134400.0 280950.0 135600.0 279750.0 ;
      RECT  132000.0 280950.0 133200.0 279750.0 ;
      RECT  136800.0 271050.0 138000.0 269850.0 ;
      RECT  136800.0 280950.0 138000.0 279750.0 ;
      RECT  132600.0 276300.0 133800.0 275100.0 ;
      RECT  132600.0 276300.0 133800.0 275100.0 ;
      RECT  135150.0 276150.0 136050.0 275250.0 ;
      RECT  130200.0 268950.0 139800.0 268050.0 ;
      RECT  130200.0 282750.0 139800.0 281850.0 ;
      RECT  102450.0 275100.0 103650.0 276300.0 ;
      RECT  104400.0 277500.0 105600.0 278700.0 ;
      RECT  121200.0 276600.0 120000.0 277800.0 ;
      RECT  112800.0 294150.0 114000.0 296100.0 ;
      RECT  112800.0 282300.0 114000.0 284250.0 ;
      RECT  108000.0 283650.0 109200.0 281850.0 ;
      RECT  108000.0 292950.0 109200.0 296550.0 ;
      RECT  110700.0 283650.0 111600.0 292950.0 ;
      RECT  108000.0 292950.0 109200.0 294150.0 ;
      RECT  110400.0 292950.0 111600.0 294150.0 ;
      RECT  110400.0 292950.0 111600.0 294150.0 ;
      RECT  108000.0 292950.0 109200.0 294150.0 ;
      RECT  108000.0 283650.0 109200.0 284850.0 ;
      RECT  110400.0 283650.0 111600.0 284850.0 ;
      RECT  110400.0 283650.0 111600.0 284850.0 ;
      RECT  108000.0 283650.0 109200.0 284850.0 ;
      RECT  112800.0 293550.0 114000.0 294750.0 ;
      RECT  112800.0 283650.0 114000.0 284850.0 ;
      RECT  108600.0 288300.0 109800.0 289500.0 ;
      RECT  108600.0 288300.0 109800.0 289500.0 ;
      RECT  111150.0 288450.0 112050.0 289350.0 ;
      RECT  106200.0 295650.0 115800.0 296550.0 ;
      RECT  106200.0 281850.0 115800.0 282750.0 ;
      RECT  117600.0 284250.0 118800.0 281850.0 ;
      RECT  117600.0 292950.0 118800.0 296550.0 ;
      RECT  122400.0 292950.0 123600.0 296550.0 ;
      RECT  124800.0 294150.0 126000.0 296100.0 ;
      RECT  124800.0 282300.0 126000.0 284250.0 ;
      RECT  117600.0 292950.0 118800.0 294150.0 ;
      RECT  120000.0 292950.0 121200.0 294150.0 ;
      RECT  120000.0 292950.0 121200.0 294150.0 ;
      RECT  117600.0 292950.0 118800.0 294150.0 ;
      RECT  120000.0 292950.0 121200.0 294150.0 ;
      RECT  122400.0 292950.0 123600.0 294150.0 ;
      RECT  122400.0 292950.0 123600.0 294150.0 ;
      RECT  120000.0 292950.0 121200.0 294150.0 ;
      RECT  117600.0 284250.0 118800.0 285450.0 ;
      RECT  120000.0 284250.0 121200.0 285450.0 ;
      RECT  120000.0 284250.0 121200.0 285450.0 ;
      RECT  117600.0 284250.0 118800.0 285450.0 ;
      RECT  120000.0 284250.0 121200.0 285450.0 ;
      RECT  122400.0 284250.0 123600.0 285450.0 ;
      RECT  122400.0 284250.0 123600.0 285450.0 ;
      RECT  120000.0 284250.0 121200.0 285450.0 ;
      RECT  124800.0 293550.0 126000.0 294750.0 ;
      RECT  124800.0 283650.0 126000.0 284850.0 ;
      RECT  122400.0 286800.0 121200.0 288000.0 ;
      RECT  119400.0 289500.0 118200.0 290700.0 ;
      RECT  120000.0 292950.0 121200.0 294150.0 ;
      RECT  122400.0 284250.0 123600.0 285450.0 ;
      RECT  123600.0 289500.0 122400.0 290700.0 ;
      RECT  118200.0 289500.0 119400.0 290700.0 ;
      RECT  121200.0 286800.0 122400.0 288000.0 ;
      RECT  122400.0 289500.0 123600.0 290700.0 ;
      RECT  115800.0 295650.0 130200.0 296550.0 ;
      RECT  115800.0 281850.0 130200.0 282750.0 ;
      RECT  136800.0 294150.0 138000.0 296100.0 ;
      RECT  136800.0 282300.0 138000.0 284250.0 ;
      RECT  132000.0 283650.0 133200.0 281850.0 ;
      RECT  132000.0 292950.0 133200.0 296550.0 ;
      RECT  134700.0 283650.0 135600.0 292950.0 ;
      RECT  132000.0 292950.0 133200.0 294150.0 ;
      RECT  134400.0 292950.0 135600.0 294150.0 ;
      RECT  134400.0 292950.0 135600.0 294150.0 ;
      RECT  132000.0 292950.0 133200.0 294150.0 ;
      RECT  132000.0 283650.0 133200.0 284850.0 ;
      RECT  134400.0 283650.0 135600.0 284850.0 ;
      RECT  134400.0 283650.0 135600.0 284850.0 ;
      RECT  132000.0 283650.0 133200.0 284850.0 ;
      RECT  136800.0 293550.0 138000.0 294750.0 ;
      RECT  136800.0 283650.0 138000.0 284850.0 ;
      RECT  132600.0 288300.0 133800.0 289500.0 ;
      RECT  132600.0 288300.0 133800.0 289500.0 ;
      RECT  135150.0 288450.0 136050.0 289350.0 ;
      RECT  130200.0 295650.0 139800.0 296550.0 ;
      RECT  130200.0 281850.0 139800.0 282750.0 ;
      RECT  102450.0 288300.0 103650.0 289500.0 ;
      RECT  104400.0 285900.0 105600.0 287100.0 ;
      RECT  121200.0 286800.0 120000.0 288000.0 ;
      RECT  112800.0 298050.0 114000.0 296100.0 ;
      RECT  112800.0 309900.0 114000.0 307950.0 ;
      RECT  108000.0 308550.0 109200.0 310350.0 ;
      RECT  108000.0 299250.0 109200.0 295650.0 ;
      RECT  110700.0 308550.0 111600.0 299250.0 ;
      RECT  108000.0 299250.0 109200.0 298050.0 ;
      RECT  110400.0 299250.0 111600.0 298050.0 ;
      RECT  110400.0 299250.0 111600.0 298050.0 ;
      RECT  108000.0 299250.0 109200.0 298050.0 ;
      RECT  108000.0 308550.0 109200.0 307350.0 ;
      RECT  110400.0 308550.0 111600.0 307350.0 ;
      RECT  110400.0 308550.0 111600.0 307350.0 ;
      RECT  108000.0 308550.0 109200.0 307350.0 ;
      RECT  112800.0 298650.0 114000.0 297450.0 ;
      RECT  112800.0 308550.0 114000.0 307350.0 ;
      RECT  108600.0 303900.0 109800.0 302700.0 ;
      RECT  108600.0 303900.0 109800.0 302700.0 ;
      RECT  111150.0 303750.0 112050.0 302850.0 ;
      RECT  106200.0 296550.0 115800.0 295650.0 ;
      RECT  106200.0 310350.0 115800.0 309450.0 ;
      RECT  117600.0 307950.0 118800.0 310350.0 ;
      RECT  117600.0 299250.0 118800.0 295650.0 ;
      RECT  122400.0 299250.0 123600.0 295650.0 ;
      RECT  124800.0 298050.0 126000.0 296100.0 ;
      RECT  124800.0 309900.0 126000.0 307950.0 ;
      RECT  117600.0 299250.0 118800.0 298050.0 ;
      RECT  120000.0 299250.0 121200.0 298050.0 ;
      RECT  120000.0 299250.0 121200.0 298050.0 ;
      RECT  117600.0 299250.0 118800.0 298050.0 ;
      RECT  120000.0 299250.0 121200.0 298050.0 ;
      RECT  122400.0 299250.0 123600.0 298050.0 ;
      RECT  122400.0 299250.0 123600.0 298050.0 ;
      RECT  120000.0 299250.0 121200.0 298050.0 ;
      RECT  117600.0 307950.0 118800.0 306750.0 ;
      RECT  120000.0 307950.0 121200.0 306750.0 ;
      RECT  120000.0 307950.0 121200.0 306750.0 ;
      RECT  117600.0 307950.0 118800.0 306750.0 ;
      RECT  120000.0 307950.0 121200.0 306750.0 ;
      RECT  122400.0 307950.0 123600.0 306750.0 ;
      RECT  122400.0 307950.0 123600.0 306750.0 ;
      RECT  120000.0 307950.0 121200.0 306750.0 ;
      RECT  124800.0 298650.0 126000.0 297450.0 ;
      RECT  124800.0 308550.0 126000.0 307350.0 ;
      RECT  122400.0 305400.0 121200.0 304200.0 ;
      RECT  119400.0 302700.0 118200.0 301500.0 ;
      RECT  120000.0 299250.0 121200.0 298050.0 ;
      RECT  122400.0 307950.0 123600.0 306750.0 ;
      RECT  123600.0 302700.0 122400.0 301500.0 ;
      RECT  118200.0 302700.0 119400.0 301500.0 ;
      RECT  121200.0 305400.0 122400.0 304200.0 ;
      RECT  122400.0 302700.0 123600.0 301500.0 ;
      RECT  115800.0 296550.0 130200.0 295650.0 ;
      RECT  115800.0 310350.0 130200.0 309450.0 ;
      RECT  136800.0 298050.0 138000.0 296100.0 ;
      RECT  136800.0 309900.0 138000.0 307950.0 ;
      RECT  132000.0 308550.0 133200.0 310350.0 ;
      RECT  132000.0 299250.0 133200.0 295650.0 ;
      RECT  134700.0 308550.0 135600.0 299250.0 ;
      RECT  132000.0 299250.0 133200.0 298050.0 ;
      RECT  134400.0 299250.0 135600.0 298050.0 ;
      RECT  134400.0 299250.0 135600.0 298050.0 ;
      RECT  132000.0 299250.0 133200.0 298050.0 ;
      RECT  132000.0 308550.0 133200.0 307350.0 ;
      RECT  134400.0 308550.0 135600.0 307350.0 ;
      RECT  134400.0 308550.0 135600.0 307350.0 ;
      RECT  132000.0 308550.0 133200.0 307350.0 ;
      RECT  136800.0 298650.0 138000.0 297450.0 ;
      RECT  136800.0 308550.0 138000.0 307350.0 ;
      RECT  132600.0 303900.0 133800.0 302700.0 ;
      RECT  132600.0 303900.0 133800.0 302700.0 ;
      RECT  135150.0 303750.0 136050.0 302850.0 ;
      RECT  130200.0 296550.0 139800.0 295650.0 ;
      RECT  130200.0 310350.0 139800.0 309450.0 ;
      RECT  102450.0 302700.0 103650.0 303900.0 ;
      RECT  104400.0 305100.0 105600.0 306300.0 ;
      RECT  121200.0 304200.0 120000.0 305400.0 ;
      RECT  112800.0 321750.0 114000.0 323700.0 ;
      RECT  112800.0 309900.0 114000.0 311850.0 ;
      RECT  108000.0 311250.0 109200.0 309450.0 ;
      RECT  108000.0 320550.0 109200.0 324150.0 ;
      RECT  110700.0 311250.0 111600.0 320550.0 ;
      RECT  108000.0 320550.0 109200.0 321750.0 ;
      RECT  110400.0 320550.0 111600.0 321750.0 ;
      RECT  110400.0 320550.0 111600.0 321750.0 ;
      RECT  108000.0 320550.0 109200.0 321750.0 ;
      RECT  108000.0 311250.0 109200.0 312450.0 ;
      RECT  110400.0 311250.0 111600.0 312450.0 ;
      RECT  110400.0 311250.0 111600.0 312450.0 ;
      RECT  108000.0 311250.0 109200.0 312450.0 ;
      RECT  112800.0 321150.0 114000.0 322350.0 ;
      RECT  112800.0 311250.0 114000.0 312450.0 ;
      RECT  108600.0 315900.0 109800.0 317100.0 ;
      RECT  108600.0 315900.0 109800.0 317100.0 ;
      RECT  111150.0 316050.0 112050.0 316950.0 ;
      RECT  106200.0 323250.0 115800.0 324150.0 ;
      RECT  106200.0 309450.0 115800.0 310350.0 ;
      RECT  117600.0 311850.0 118800.0 309450.0 ;
      RECT  117600.0 320550.0 118800.0 324150.0 ;
      RECT  122400.0 320550.0 123600.0 324150.0 ;
      RECT  124800.0 321750.0 126000.0 323700.0 ;
      RECT  124800.0 309900.0 126000.0 311850.0 ;
      RECT  117600.0 320550.0 118800.0 321750.0 ;
      RECT  120000.0 320550.0 121200.0 321750.0 ;
      RECT  120000.0 320550.0 121200.0 321750.0 ;
      RECT  117600.0 320550.0 118800.0 321750.0 ;
      RECT  120000.0 320550.0 121200.0 321750.0 ;
      RECT  122400.0 320550.0 123600.0 321750.0 ;
      RECT  122400.0 320550.0 123600.0 321750.0 ;
      RECT  120000.0 320550.0 121200.0 321750.0 ;
      RECT  117600.0 311850.0 118800.0 313050.0 ;
      RECT  120000.0 311850.0 121200.0 313050.0 ;
      RECT  120000.0 311850.0 121200.0 313050.0 ;
      RECT  117600.0 311850.0 118800.0 313050.0 ;
      RECT  120000.0 311850.0 121200.0 313050.0 ;
      RECT  122400.0 311850.0 123600.0 313050.0 ;
      RECT  122400.0 311850.0 123600.0 313050.0 ;
      RECT  120000.0 311850.0 121200.0 313050.0 ;
      RECT  124800.0 321150.0 126000.0 322350.0 ;
      RECT  124800.0 311250.0 126000.0 312450.0 ;
      RECT  122400.0 314400.0 121200.0 315600.0 ;
      RECT  119400.0 317100.0 118200.0 318300.0 ;
      RECT  120000.0 320550.0 121200.0 321750.0 ;
      RECT  122400.0 311850.0 123600.0 313050.0 ;
      RECT  123600.0 317100.0 122400.0 318300.0 ;
      RECT  118200.0 317100.0 119400.0 318300.0 ;
      RECT  121200.0 314400.0 122400.0 315600.0 ;
      RECT  122400.0 317100.0 123600.0 318300.0 ;
      RECT  115800.0 323250.0 130200.0 324150.0 ;
      RECT  115800.0 309450.0 130200.0 310350.0 ;
      RECT  136800.0 321750.0 138000.0 323700.0 ;
      RECT  136800.0 309900.0 138000.0 311850.0 ;
      RECT  132000.0 311250.0 133200.0 309450.0 ;
      RECT  132000.0 320550.0 133200.0 324150.0 ;
      RECT  134700.0 311250.0 135600.0 320550.0 ;
      RECT  132000.0 320550.0 133200.0 321750.0 ;
      RECT  134400.0 320550.0 135600.0 321750.0 ;
      RECT  134400.0 320550.0 135600.0 321750.0 ;
      RECT  132000.0 320550.0 133200.0 321750.0 ;
      RECT  132000.0 311250.0 133200.0 312450.0 ;
      RECT  134400.0 311250.0 135600.0 312450.0 ;
      RECT  134400.0 311250.0 135600.0 312450.0 ;
      RECT  132000.0 311250.0 133200.0 312450.0 ;
      RECT  136800.0 321150.0 138000.0 322350.0 ;
      RECT  136800.0 311250.0 138000.0 312450.0 ;
      RECT  132600.0 315900.0 133800.0 317100.0 ;
      RECT  132600.0 315900.0 133800.0 317100.0 ;
      RECT  135150.0 316050.0 136050.0 316950.0 ;
      RECT  130200.0 323250.0 139800.0 324150.0 ;
      RECT  130200.0 309450.0 139800.0 310350.0 ;
      RECT  102450.0 315900.0 103650.0 317100.0 ;
      RECT  104400.0 313500.0 105600.0 314700.0 ;
      RECT  121200.0 314400.0 120000.0 315600.0 ;
      RECT  112800.0 325650.0 114000.0 323700.0 ;
      RECT  112800.0 337500.0 114000.0 335550.0 ;
      RECT  108000.0 336150.0 109200.0 337950.0 ;
      RECT  108000.0 326850.0 109200.0 323250.0 ;
      RECT  110700.0 336150.0 111600.0 326850.0 ;
      RECT  108000.0 326850.0 109200.0 325650.0 ;
      RECT  110400.0 326850.0 111600.0 325650.0 ;
      RECT  110400.0 326850.0 111600.0 325650.0 ;
      RECT  108000.0 326850.0 109200.0 325650.0 ;
      RECT  108000.0 336150.0 109200.0 334950.0 ;
      RECT  110400.0 336150.0 111600.0 334950.0 ;
      RECT  110400.0 336150.0 111600.0 334950.0 ;
      RECT  108000.0 336150.0 109200.0 334950.0 ;
      RECT  112800.0 326250.0 114000.0 325050.0 ;
      RECT  112800.0 336150.0 114000.0 334950.0 ;
      RECT  108600.0 331500.0 109800.0 330300.0 ;
      RECT  108600.0 331500.0 109800.0 330300.0 ;
      RECT  111150.0 331350.0 112050.0 330450.0 ;
      RECT  106200.0 324150.0 115800.0 323250.0 ;
      RECT  106200.0 337950.0 115800.0 337050.0 ;
      RECT  117600.0 335550.0 118800.0 337950.0 ;
      RECT  117600.0 326850.0 118800.0 323250.0 ;
      RECT  122400.0 326850.0 123600.0 323250.0 ;
      RECT  124800.0 325650.0 126000.0 323700.0 ;
      RECT  124800.0 337500.0 126000.0 335550.0 ;
      RECT  117600.0 326850.0 118800.0 325650.0 ;
      RECT  120000.0 326850.0 121200.0 325650.0 ;
      RECT  120000.0 326850.0 121200.0 325650.0 ;
      RECT  117600.0 326850.0 118800.0 325650.0 ;
      RECT  120000.0 326850.0 121200.0 325650.0 ;
      RECT  122400.0 326850.0 123600.0 325650.0 ;
      RECT  122400.0 326850.0 123600.0 325650.0 ;
      RECT  120000.0 326850.0 121200.0 325650.0 ;
      RECT  117600.0 335550.0 118800.0 334350.0 ;
      RECT  120000.0 335550.0 121200.0 334350.0 ;
      RECT  120000.0 335550.0 121200.0 334350.0 ;
      RECT  117600.0 335550.0 118800.0 334350.0 ;
      RECT  120000.0 335550.0 121200.0 334350.0 ;
      RECT  122400.0 335550.0 123600.0 334350.0 ;
      RECT  122400.0 335550.0 123600.0 334350.0 ;
      RECT  120000.0 335550.0 121200.0 334350.0 ;
      RECT  124800.0 326250.0 126000.0 325050.0 ;
      RECT  124800.0 336150.0 126000.0 334950.0 ;
      RECT  122400.0 333000.0 121200.0 331800.0 ;
      RECT  119400.0 330300.0 118200.0 329100.0 ;
      RECT  120000.0 326850.0 121200.0 325650.0 ;
      RECT  122400.0 335550.0 123600.0 334350.0 ;
      RECT  123600.0 330300.0 122400.0 329100.0 ;
      RECT  118200.0 330300.0 119400.0 329100.0 ;
      RECT  121200.0 333000.0 122400.0 331800.0 ;
      RECT  122400.0 330300.0 123600.0 329100.0 ;
      RECT  115800.0 324150.0 130200.0 323250.0 ;
      RECT  115800.0 337950.0 130200.0 337050.0 ;
      RECT  136800.0 325650.0 138000.0 323700.0 ;
      RECT  136800.0 337500.0 138000.0 335550.0 ;
      RECT  132000.0 336150.0 133200.0 337950.0 ;
      RECT  132000.0 326850.0 133200.0 323250.0 ;
      RECT  134700.0 336150.0 135600.0 326850.0 ;
      RECT  132000.0 326850.0 133200.0 325650.0 ;
      RECT  134400.0 326850.0 135600.0 325650.0 ;
      RECT  134400.0 326850.0 135600.0 325650.0 ;
      RECT  132000.0 326850.0 133200.0 325650.0 ;
      RECT  132000.0 336150.0 133200.0 334950.0 ;
      RECT  134400.0 336150.0 135600.0 334950.0 ;
      RECT  134400.0 336150.0 135600.0 334950.0 ;
      RECT  132000.0 336150.0 133200.0 334950.0 ;
      RECT  136800.0 326250.0 138000.0 325050.0 ;
      RECT  136800.0 336150.0 138000.0 334950.0 ;
      RECT  132600.0 331500.0 133800.0 330300.0 ;
      RECT  132600.0 331500.0 133800.0 330300.0 ;
      RECT  135150.0 331350.0 136050.0 330450.0 ;
      RECT  130200.0 324150.0 139800.0 323250.0 ;
      RECT  130200.0 337950.0 139800.0 337050.0 ;
      RECT  102450.0 330300.0 103650.0 331500.0 ;
      RECT  104400.0 332700.0 105600.0 333900.0 ;
      RECT  121200.0 331800.0 120000.0 333000.0 ;
      RECT  112800.0 349350.0 114000.0 351300.0 ;
      RECT  112800.0 337500.0 114000.0 339450.0 ;
      RECT  108000.0 338850.0 109200.0 337050.0 ;
      RECT  108000.0 348150.0 109200.0 351750.0 ;
      RECT  110700.0 338850.0 111600.0 348150.0 ;
      RECT  108000.0 348150.0 109200.0 349350.0 ;
      RECT  110400.0 348150.0 111600.0 349350.0 ;
      RECT  110400.0 348150.0 111600.0 349350.0 ;
      RECT  108000.0 348150.0 109200.0 349350.0 ;
      RECT  108000.0 338850.0 109200.0 340050.0 ;
      RECT  110400.0 338850.0 111600.0 340050.0 ;
      RECT  110400.0 338850.0 111600.0 340050.0 ;
      RECT  108000.0 338850.0 109200.0 340050.0 ;
      RECT  112800.0 348750.0 114000.0 349950.0 ;
      RECT  112800.0 338850.0 114000.0 340050.0 ;
      RECT  108600.0 343500.0 109800.0 344700.0 ;
      RECT  108600.0 343500.0 109800.0 344700.0 ;
      RECT  111150.0 343650.0 112050.0 344550.0 ;
      RECT  106200.0 350850.0 115800.0 351750.0 ;
      RECT  106200.0 337050.0 115800.0 337950.0 ;
      RECT  117600.0 339450.0 118800.0 337050.0 ;
      RECT  117600.0 348150.0 118800.0 351750.0 ;
      RECT  122400.0 348150.0 123600.0 351750.0 ;
      RECT  124800.0 349350.0 126000.0 351300.0 ;
      RECT  124800.0 337500.0 126000.0 339450.0 ;
      RECT  117600.0 348150.0 118800.0 349350.0 ;
      RECT  120000.0 348150.0 121200.0 349350.0 ;
      RECT  120000.0 348150.0 121200.0 349350.0 ;
      RECT  117600.0 348150.0 118800.0 349350.0 ;
      RECT  120000.0 348150.0 121200.0 349350.0 ;
      RECT  122400.0 348150.0 123600.0 349350.0 ;
      RECT  122400.0 348150.0 123600.0 349350.0 ;
      RECT  120000.0 348150.0 121200.0 349350.0 ;
      RECT  117600.0 339450.0 118800.0 340650.0 ;
      RECT  120000.0 339450.0 121200.0 340650.0 ;
      RECT  120000.0 339450.0 121200.0 340650.0 ;
      RECT  117600.0 339450.0 118800.0 340650.0 ;
      RECT  120000.0 339450.0 121200.0 340650.0 ;
      RECT  122400.0 339450.0 123600.0 340650.0 ;
      RECT  122400.0 339450.0 123600.0 340650.0 ;
      RECT  120000.0 339450.0 121200.0 340650.0 ;
      RECT  124800.0 348750.0 126000.0 349950.0 ;
      RECT  124800.0 338850.0 126000.0 340050.0 ;
      RECT  122400.0 342000.0 121200.0 343200.0 ;
      RECT  119400.0 344700.0 118200.0 345900.0 ;
      RECT  120000.0 348150.0 121200.0 349350.0 ;
      RECT  122400.0 339450.0 123600.0 340650.0 ;
      RECT  123600.0 344700.0 122400.0 345900.0 ;
      RECT  118200.0 344700.0 119400.0 345900.0 ;
      RECT  121200.0 342000.0 122400.0 343200.0 ;
      RECT  122400.0 344700.0 123600.0 345900.0 ;
      RECT  115800.0 350850.0 130200.0 351750.0 ;
      RECT  115800.0 337050.0 130200.0 337950.0 ;
      RECT  136800.0 349350.0 138000.0 351300.0 ;
      RECT  136800.0 337500.0 138000.0 339450.0 ;
      RECT  132000.0 338850.0 133200.0 337050.0 ;
      RECT  132000.0 348150.0 133200.0 351750.0 ;
      RECT  134700.0 338850.0 135600.0 348150.0 ;
      RECT  132000.0 348150.0 133200.0 349350.0 ;
      RECT  134400.0 348150.0 135600.0 349350.0 ;
      RECT  134400.0 348150.0 135600.0 349350.0 ;
      RECT  132000.0 348150.0 133200.0 349350.0 ;
      RECT  132000.0 338850.0 133200.0 340050.0 ;
      RECT  134400.0 338850.0 135600.0 340050.0 ;
      RECT  134400.0 338850.0 135600.0 340050.0 ;
      RECT  132000.0 338850.0 133200.0 340050.0 ;
      RECT  136800.0 348750.0 138000.0 349950.0 ;
      RECT  136800.0 338850.0 138000.0 340050.0 ;
      RECT  132600.0 343500.0 133800.0 344700.0 ;
      RECT  132600.0 343500.0 133800.0 344700.0 ;
      RECT  135150.0 343650.0 136050.0 344550.0 ;
      RECT  130200.0 350850.0 139800.0 351750.0 ;
      RECT  130200.0 337050.0 139800.0 337950.0 ;
      RECT  102450.0 343500.0 103650.0 344700.0 ;
      RECT  104400.0 341100.0 105600.0 342300.0 ;
      RECT  121200.0 342000.0 120000.0 343200.0 ;
      RECT  112800.0 353250.0 114000.0 351300.0 ;
      RECT  112800.0 365100.0 114000.0 363150.0 ;
      RECT  108000.0 363750.0 109200.0 365550.0 ;
      RECT  108000.0 354450.0 109200.0 350850.0 ;
      RECT  110700.0 363750.0 111600.0 354450.0 ;
      RECT  108000.0 354450.0 109200.0 353250.0 ;
      RECT  110400.0 354450.0 111600.0 353250.0 ;
      RECT  110400.0 354450.0 111600.0 353250.0 ;
      RECT  108000.0 354450.0 109200.0 353250.0 ;
      RECT  108000.0 363750.0 109200.0 362550.0 ;
      RECT  110400.0 363750.0 111600.0 362550.0 ;
      RECT  110400.0 363750.0 111600.0 362550.0 ;
      RECT  108000.0 363750.0 109200.0 362550.0 ;
      RECT  112800.0 353850.0 114000.0 352650.0 ;
      RECT  112800.0 363750.0 114000.0 362550.0 ;
      RECT  108600.0 359100.0 109800.0 357900.0 ;
      RECT  108600.0 359100.0 109800.0 357900.0 ;
      RECT  111150.0 358950.0 112050.0 358050.0 ;
      RECT  106200.0 351750.0 115800.0 350850.0 ;
      RECT  106200.0 365550.0 115800.0 364650.0 ;
      RECT  117600.0 363150.0 118800.0 365550.0 ;
      RECT  117600.0 354450.0 118800.0 350850.0 ;
      RECT  122400.0 354450.0 123600.0 350850.0 ;
      RECT  124800.0 353250.0 126000.0 351300.0 ;
      RECT  124800.0 365100.0 126000.0 363150.0 ;
      RECT  117600.0 354450.0 118800.0 353250.0 ;
      RECT  120000.0 354450.0 121200.0 353250.0 ;
      RECT  120000.0 354450.0 121200.0 353250.0 ;
      RECT  117600.0 354450.0 118800.0 353250.0 ;
      RECT  120000.0 354450.0 121200.0 353250.0 ;
      RECT  122400.0 354450.0 123600.0 353250.0 ;
      RECT  122400.0 354450.0 123600.0 353250.0 ;
      RECT  120000.0 354450.0 121200.0 353250.0 ;
      RECT  117600.0 363150.0 118800.0 361950.0 ;
      RECT  120000.0 363150.0 121200.0 361950.0 ;
      RECT  120000.0 363150.0 121200.0 361950.0 ;
      RECT  117600.0 363150.0 118800.0 361950.0 ;
      RECT  120000.0 363150.0 121200.0 361950.0 ;
      RECT  122400.0 363150.0 123600.0 361950.0 ;
      RECT  122400.0 363150.0 123600.0 361950.0 ;
      RECT  120000.0 363150.0 121200.0 361950.0 ;
      RECT  124800.0 353850.0 126000.0 352650.0 ;
      RECT  124800.0 363750.0 126000.0 362550.0 ;
      RECT  122400.0 360600.0 121200.0 359400.0 ;
      RECT  119400.0 357900.0 118200.0 356700.0 ;
      RECT  120000.0 354450.0 121200.0 353250.0 ;
      RECT  122400.0 363150.0 123600.0 361950.0 ;
      RECT  123600.0 357900.0 122400.0 356700.0 ;
      RECT  118200.0 357900.0 119400.0 356700.0 ;
      RECT  121200.0 360600.0 122400.0 359400.0 ;
      RECT  122400.0 357900.0 123600.0 356700.0 ;
      RECT  115800.0 351750.0 130200.0 350850.0 ;
      RECT  115800.0 365550.0 130200.0 364650.0 ;
      RECT  136800.0 353250.0 138000.0 351300.0 ;
      RECT  136800.0 365100.0 138000.0 363150.0 ;
      RECT  132000.0 363750.0 133200.0 365550.0 ;
      RECT  132000.0 354450.0 133200.0 350850.0 ;
      RECT  134700.0 363750.0 135600.0 354450.0 ;
      RECT  132000.0 354450.0 133200.0 353250.0 ;
      RECT  134400.0 354450.0 135600.0 353250.0 ;
      RECT  134400.0 354450.0 135600.0 353250.0 ;
      RECT  132000.0 354450.0 133200.0 353250.0 ;
      RECT  132000.0 363750.0 133200.0 362550.0 ;
      RECT  134400.0 363750.0 135600.0 362550.0 ;
      RECT  134400.0 363750.0 135600.0 362550.0 ;
      RECT  132000.0 363750.0 133200.0 362550.0 ;
      RECT  136800.0 353850.0 138000.0 352650.0 ;
      RECT  136800.0 363750.0 138000.0 362550.0 ;
      RECT  132600.0 359100.0 133800.0 357900.0 ;
      RECT  132600.0 359100.0 133800.0 357900.0 ;
      RECT  135150.0 358950.0 136050.0 358050.0 ;
      RECT  130200.0 351750.0 139800.0 350850.0 ;
      RECT  130200.0 365550.0 139800.0 364650.0 ;
      RECT  102450.0 357900.0 103650.0 359100.0 ;
      RECT  104400.0 360300.0 105600.0 361500.0 ;
      RECT  121200.0 359400.0 120000.0 360600.0 ;
      RECT  112800.0 376950.0 114000.0 378900.0 ;
      RECT  112800.0 365100.0 114000.0 367050.0 ;
      RECT  108000.0 366450.0 109200.0 364650.0 ;
      RECT  108000.0 375750.0 109200.0 379350.0 ;
      RECT  110700.0 366450.0 111600.0 375750.0 ;
      RECT  108000.0 375750.0 109200.0 376950.0 ;
      RECT  110400.0 375750.0 111600.0 376950.0 ;
      RECT  110400.0 375750.0 111600.0 376950.0 ;
      RECT  108000.0 375750.0 109200.0 376950.0 ;
      RECT  108000.0 366450.0 109200.0 367650.0 ;
      RECT  110400.0 366450.0 111600.0 367650.0 ;
      RECT  110400.0 366450.0 111600.0 367650.0 ;
      RECT  108000.0 366450.0 109200.0 367650.0 ;
      RECT  112800.0 376350.0 114000.0 377550.0 ;
      RECT  112800.0 366450.0 114000.0 367650.0 ;
      RECT  108600.0 371100.0 109800.0 372300.0 ;
      RECT  108600.0 371100.0 109800.0 372300.0 ;
      RECT  111150.0 371250.0 112050.0 372150.0 ;
      RECT  106200.0 378450.0 115800.0 379350.0 ;
      RECT  106200.0 364650.0 115800.0 365550.0 ;
      RECT  117600.0 367050.0 118800.0 364650.0 ;
      RECT  117600.0 375750.0 118800.0 379350.0 ;
      RECT  122400.0 375750.0 123600.0 379350.0 ;
      RECT  124800.0 376950.0 126000.0 378900.0 ;
      RECT  124800.0 365100.0 126000.0 367050.0 ;
      RECT  117600.0 375750.0 118800.0 376950.0 ;
      RECT  120000.0 375750.0 121200.0 376950.0 ;
      RECT  120000.0 375750.0 121200.0 376950.0 ;
      RECT  117600.0 375750.0 118800.0 376950.0 ;
      RECT  120000.0 375750.0 121200.0 376950.0 ;
      RECT  122400.0 375750.0 123600.0 376950.0 ;
      RECT  122400.0 375750.0 123600.0 376950.0 ;
      RECT  120000.0 375750.0 121200.0 376950.0 ;
      RECT  117600.0 367050.0 118800.0 368250.0 ;
      RECT  120000.0 367050.0 121200.0 368250.0 ;
      RECT  120000.0 367050.0 121200.0 368250.0 ;
      RECT  117600.0 367050.0 118800.0 368250.0 ;
      RECT  120000.0 367050.0 121200.0 368250.0 ;
      RECT  122400.0 367050.0 123600.0 368250.0 ;
      RECT  122400.0 367050.0 123600.0 368250.0 ;
      RECT  120000.0 367050.0 121200.0 368250.0 ;
      RECT  124800.0 376350.0 126000.0 377550.0 ;
      RECT  124800.0 366450.0 126000.0 367650.0 ;
      RECT  122400.0 369600.0 121200.0 370800.0 ;
      RECT  119400.0 372300.0 118200.0 373500.0 ;
      RECT  120000.0 375750.0 121200.0 376950.0 ;
      RECT  122400.0 367050.0 123600.0 368250.0 ;
      RECT  123600.0 372300.0 122400.0 373500.0 ;
      RECT  118200.0 372300.0 119400.0 373500.0 ;
      RECT  121200.0 369600.0 122400.0 370800.0 ;
      RECT  122400.0 372300.0 123600.0 373500.0 ;
      RECT  115800.0 378450.0 130200.0 379350.0 ;
      RECT  115800.0 364650.0 130200.0 365550.0 ;
      RECT  136800.0 376950.0 138000.0 378900.0 ;
      RECT  136800.0 365100.0 138000.0 367050.0 ;
      RECT  132000.0 366450.0 133200.0 364650.0 ;
      RECT  132000.0 375750.0 133200.0 379350.0 ;
      RECT  134700.0 366450.0 135600.0 375750.0 ;
      RECT  132000.0 375750.0 133200.0 376950.0 ;
      RECT  134400.0 375750.0 135600.0 376950.0 ;
      RECT  134400.0 375750.0 135600.0 376950.0 ;
      RECT  132000.0 375750.0 133200.0 376950.0 ;
      RECT  132000.0 366450.0 133200.0 367650.0 ;
      RECT  134400.0 366450.0 135600.0 367650.0 ;
      RECT  134400.0 366450.0 135600.0 367650.0 ;
      RECT  132000.0 366450.0 133200.0 367650.0 ;
      RECT  136800.0 376350.0 138000.0 377550.0 ;
      RECT  136800.0 366450.0 138000.0 367650.0 ;
      RECT  132600.0 371100.0 133800.0 372300.0 ;
      RECT  132600.0 371100.0 133800.0 372300.0 ;
      RECT  135150.0 371250.0 136050.0 372150.0 ;
      RECT  130200.0 378450.0 139800.0 379350.0 ;
      RECT  130200.0 364650.0 139800.0 365550.0 ;
      RECT  102450.0 371100.0 103650.0 372300.0 ;
      RECT  104400.0 368700.0 105600.0 369900.0 ;
      RECT  121200.0 369600.0 120000.0 370800.0 ;
      RECT  112800.0 380850.0 114000.0 378900.0 ;
      RECT  112800.0 392700.0 114000.0 390750.0 ;
      RECT  108000.0 391350.0 109200.0 393150.0 ;
      RECT  108000.0 382050.0 109200.0 378450.0 ;
      RECT  110700.0 391350.0 111600.0 382050.0 ;
      RECT  108000.0 382050.0 109200.0 380850.0 ;
      RECT  110400.0 382050.0 111600.0 380850.0 ;
      RECT  110400.0 382050.0 111600.0 380850.0 ;
      RECT  108000.0 382050.0 109200.0 380850.0 ;
      RECT  108000.0 391350.0 109200.0 390150.0 ;
      RECT  110400.0 391350.0 111600.0 390150.0 ;
      RECT  110400.0 391350.0 111600.0 390150.0 ;
      RECT  108000.0 391350.0 109200.0 390150.0 ;
      RECT  112800.0 381450.0 114000.0 380250.0 ;
      RECT  112800.0 391350.0 114000.0 390150.0 ;
      RECT  108600.0 386700.0 109800.0 385500.0 ;
      RECT  108600.0 386700.0 109800.0 385500.0 ;
      RECT  111150.0 386550.0 112050.0 385650.0 ;
      RECT  106200.0 379350.0 115800.0 378450.0 ;
      RECT  106200.0 393150.0 115800.0 392250.0 ;
      RECT  117600.0 390750.0 118800.0 393150.0 ;
      RECT  117600.0 382050.0 118800.0 378450.0 ;
      RECT  122400.0 382050.0 123600.0 378450.0 ;
      RECT  124800.0 380850.0 126000.0 378900.0 ;
      RECT  124800.0 392700.0 126000.0 390750.0 ;
      RECT  117600.0 382050.0 118800.0 380850.0 ;
      RECT  120000.0 382050.0 121200.0 380850.0 ;
      RECT  120000.0 382050.0 121200.0 380850.0 ;
      RECT  117600.0 382050.0 118800.0 380850.0 ;
      RECT  120000.0 382050.0 121200.0 380850.0 ;
      RECT  122400.0 382050.0 123600.0 380850.0 ;
      RECT  122400.0 382050.0 123600.0 380850.0 ;
      RECT  120000.0 382050.0 121200.0 380850.0 ;
      RECT  117600.0 390750.0 118800.0 389550.0 ;
      RECT  120000.0 390750.0 121200.0 389550.0 ;
      RECT  120000.0 390750.0 121200.0 389550.0 ;
      RECT  117600.0 390750.0 118800.0 389550.0 ;
      RECT  120000.0 390750.0 121200.0 389550.0 ;
      RECT  122400.0 390750.0 123600.0 389550.0 ;
      RECT  122400.0 390750.0 123600.0 389550.0 ;
      RECT  120000.0 390750.0 121200.0 389550.0 ;
      RECT  124800.0 381450.0 126000.0 380250.0 ;
      RECT  124800.0 391350.0 126000.0 390150.0 ;
      RECT  122400.0 388200.0 121200.0 387000.0 ;
      RECT  119400.0 385500.0 118200.0 384300.0 ;
      RECT  120000.0 382050.0 121200.0 380850.0 ;
      RECT  122400.0 390750.0 123600.0 389550.0 ;
      RECT  123600.0 385500.0 122400.0 384300.0 ;
      RECT  118200.0 385500.0 119400.0 384300.0 ;
      RECT  121200.0 388200.0 122400.0 387000.0 ;
      RECT  122400.0 385500.0 123600.0 384300.0 ;
      RECT  115800.0 379350.0 130200.0 378450.0 ;
      RECT  115800.0 393150.0 130200.0 392250.0 ;
      RECT  136800.0 380850.0 138000.0 378900.0 ;
      RECT  136800.0 392700.0 138000.0 390750.0 ;
      RECT  132000.0 391350.0 133200.0 393150.0 ;
      RECT  132000.0 382050.0 133200.0 378450.0 ;
      RECT  134700.0 391350.0 135600.0 382050.0 ;
      RECT  132000.0 382050.0 133200.0 380850.0 ;
      RECT  134400.0 382050.0 135600.0 380850.0 ;
      RECT  134400.0 382050.0 135600.0 380850.0 ;
      RECT  132000.0 382050.0 133200.0 380850.0 ;
      RECT  132000.0 391350.0 133200.0 390150.0 ;
      RECT  134400.0 391350.0 135600.0 390150.0 ;
      RECT  134400.0 391350.0 135600.0 390150.0 ;
      RECT  132000.0 391350.0 133200.0 390150.0 ;
      RECT  136800.0 381450.0 138000.0 380250.0 ;
      RECT  136800.0 391350.0 138000.0 390150.0 ;
      RECT  132600.0 386700.0 133800.0 385500.0 ;
      RECT  132600.0 386700.0 133800.0 385500.0 ;
      RECT  135150.0 386550.0 136050.0 385650.0 ;
      RECT  130200.0 379350.0 139800.0 378450.0 ;
      RECT  130200.0 393150.0 139800.0 392250.0 ;
      RECT  102450.0 385500.0 103650.0 386700.0 ;
      RECT  104400.0 387900.0 105600.0 389100.0 ;
      RECT  121200.0 387000.0 120000.0 388200.0 ;
      RECT  112800.0 404550.0 114000.0 406500.0 ;
      RECT  112800.0 392700.0 114000.0 394650.0 ;
      RECT  108000.0 394050.0 109200.0 392250.0 ;
      RECT  108000.0 403350.0 109200.0 406950.0 ;
      RECT  110700.0 394050.0 111600.0 403350.0 ;
      RECT  108000.0 403350.0 109200.0 404550.0 ;
      RECT  110400.0 403350.0 111600.0 404550.0 ;
      RECT  110400.0 403350.0 111600.0 404550.0 ;
      RECT  108000.0 403350.0 109200.0 404550.0 ;
      RECT  108000.0 394050.0 109200.0 395250.0 ;
      RECT  110400.0 394050.0 111600.0 395250.0 ;
      RECT  110400.0 394050.0 111600.0 395250.0 ;
      RECT  108000.0 394050.0 109200.0 395250.0 ;
      RECT  112800.0 403950.0 114000.0 405150.0 ;
      RECT  112800.0 394050.0 114000.0 395250.0 ;
      RECT  108600.0 398700.0 109800.0 399900.0 ;
      RECT  108600.0 398700.0 109800.0 399900.0 ;
      RECT  111150.0 398850.0 112050.0 399750.0 ;
      RECT  106200.0 406050.0 115800.0 406950.0 ;
      RECT  106200.0 392250.0 115800.0 393150.0 ;
      RECT  117600.0 394650.0 118800.0 392250.0 ;
      RECT  117600.0 403350.0 118800.0 406950.0 ;
      RECT  122400.0 403350.0 123600.0 406950.0 ;
      RECT  124800.0 404550.0 126000.0 406500.0 ;
      RECT  124800.0 392700.0 126000.0 394650.0 ;
      RECT  117600.0 403350.0 118800.0 404550.0 ;
      RECT  120000.0 403350.0 121200.0 404550.0 ;
      RECT  120000.0 403350.0 121200.0 404550.0 ;
      RECT  117600.0 403350.0 118800.0 404550.0 ;
      RECT  120000.0 403350.0 121200.0 404550.0 ;
      RECT  122400.0 403350.0 123600.0 404550.0 ;
      RECT  122400.0 403350.0 123600.0 404550.0 ;
      RECT  120000.0 403350.0 121200.0 404550.0 ;
      RECT  117600.0 394650.0 118800.0 395850.0 ;
      RECT  120000.0 394650.0 121200.0 395850.0 ;
      RECT  120000.0 394650.0 121200.0 395850.0 ;
      RECT  117600.0 394650.0 118800.0 395850.0 ;
      RECT  120000.0 394650.0 121200.0 395850.0 ;
      RECT  122400.0 394650.0 123600.0 395850.0 ;
      RECT  122400.0 394650.0 123600.0 395850.0 ;
      RECT  120000.0 394650.0 121200.0 395850.0 ;
      RECT  124800.0 403950.0 126000.0 405150.0 ;
      RECT  124800.0 394050.0 126000.0 395250.0 ;
      RECT  122400.0 397200.0 121200.0 398400.0 ;
      RECT  119400.0 399900.0 118200.0 401100.0 ;
      RECT  120000.0 403350.0 121200.0 404550.0 ;
      RECT  122400.0 394650.0 123600.0 395850.0 ;
      RECT  123600.0 399900.0 122400.0 401100.0 ;
      RECT  118200.0 399900.0 119400.0 401100.0 ;
      RECT  121200.0 397200.0 122400.0 398400.0 ;
      RECT  122400.0 399900.0 123600.0 401100.0 ;
      RECT  115800.0 406050.0 130200.0 406950.0 ;
      RECT  115800.0 392250.0 130200.0 393150.0 ;
      RECT  136800.0 404550.0 138000.0 406500.0 ;
      RECT  136800.0 392700.0 138000.0 394650.0 ;
      RECT  132000.0 394050.0 133200.0 392250.0 ;
      RECT  132000.0 403350.0 133200.0 406950.0 ;
      RECT  134700.0 394050.0 135600.0 403350.0 ;
      RECT  132000.0 403350.0 133200.0 404550.0 ;
      RECT  134400.0 403350.0 135600.0 404550.0 ;
      RECT  134400.0 403350.0 135600.0 404550.0 ;
      RECT  132000.0 403350.0 133200.0 404550.0 ;
      RECT  132000.0 394050.0 133200.0 395250.0 ;
      RECT  134400.0 394050.0 135600.0 395250.0 ;
      RECT  134400.0 394050.0 135600.0 395250.0 ;
      RECT  132000.0 394050.0 133200.0 395250.0 ;
      RECT  136800.0 403950.0 138000.0 405150.0 ;
      RECT  136800.0 394050.0 138000.0 395250.0 ;
      RECT  132600.0 398700.0 133800.0 399900.0 ;
      RECT  132600.0 398700.0 133800.0 399900.0 ;
      RECT  135150.0 398850.0 136050.0 399750.0 ;
      RECT  130200.0 406050.0 139800.0 406950.0 ;
      RECT  130200.0 392250.0 139800.0 393150.0 ;
      RECT  102450.0 398700.0 103650.0 399900.0 ;
      RECT  104400.0 396300.0 105600.0 397500.0 ;
      RECT  121200.0 397200.0 120000.0 398400.0 ;
      RECT  112800.0 408450.0 114000.0 406500.0 ;
      RECT  112800.0 420300.0 114000.0 418350.0 ;
      RECT  108000.0 418950.0 109200.0 420750.0 ;
      RECT  108000.0 409650.0 109200.0 406050.0 ;
      RECT  110700.0 418950.0 111600.0 409650.0 ;
      RECT  108000.0 409650.0 109200.0 408450.0 ;
      RECT  110400.0 409650.0 111600.0 408450.0 ;
      RECT  110400.0 409650.0 111600.0 408450.0 ;
      RECT  108000.0 409650.0 109200.0 408450.0 ;
      RECT  108000.0 418950.0 109200.0 417750.0 ;
      RECT  110400.0 418950.0 111600.0 417750.0 ;
      RECT  110400.0 418950.0 111600.0 417750.0 ;
      RECT  108000.0 418950.0 109200.0 417750.0 ;
      RECT  112800.0 409050.0 114000.0 407850.0 ;
      RECT  112800.0 418950.0 114000.0 417750.0 ;
      RECT  108600.0 414300.0 109800.0 413100.0 ;
      RECT  108600.0 414300.0 109800.0 413100.0 ;
      RECT  111150.0 414150.0 112050.0 413250.0 ;
      RECT  106200.0 406950.0 115800.0 406050.0 ;
      RECT  106200.0 420750.0 115800.0 419850.0 ;
      RECT  117600.0 418350.0 118800.0 420750.0 ;
      RECT  117600.0 409650.0 118800.0 406050.0 ;
      RECT  122400.0 409650.0 123600.0 406050.0 ;
      RECT  124800.0 408450.0 126000.0 406500.0 ;
      RECT  124800.0 420300.0 126000.0 418350.0 ;
      RECT  117600.0 409650.0 118800.0 408450.0 ;
      RECT  120000.0 409650.0 121200.0 408450.0 ;
      RECT  120000.0 409650.0 121200.0 408450.0 ;
      RECT  117600.0 409650.0 118800.0 408450.0 ;
      RECT  120000.0 409650.0 121200.0 408450.0 ;
      RECT  122400.0 409650.0 123600.0 408450.0 ;
      RECT  122400.0 409650.0 123600.0 408450.0 ;
      RECT  120000.0 409650.0 121200.0 408450.0 ;
      RECT  117600.0 418350.0 118800.0 417150.0 ;
      RECT  120000.0 418350.0 121200.0 417150.0 ;
      RECT  120000.0 418350.0 121200.0 417150.0 ;
      RECT  117600.0 418350.0 118800.0 417150.0 ;
      RECT  120000.0 418350.0 121200.0 417150.0 ;
      RECT  122400.0 418350.0 123600.0 417150.0 ;
      RECT  122400.0 418350.0 123600.0 417150.0 ;
      RECT  120000.0 418350.0 121200.0 417150.0 ;
      RECT  124800.0 409050.0 126000.0 407850.0 ;
      RECT  124800.0 418950.0 126000.0 417750.0 ;
      RECT  122400.0 415800.0 121200.0 414600.0 ;
      RECT  119400.0 413100.0 118200.0 411900.0 ;
      RECT  120000.0 409650.0 121200.0 408450.0 ;
      RECT  122400.0 418350.0 123600.0 417150.0 ;
      RECT  123600.0 413100.0 122400.0 411900.0 ;
      RECT  118200.0 413100.0 119400.0 411900.0 ;
      RECT  121200.0 415800.0 122400.0 414600.0 ;
      RECT  122400.0 413100.0 123600.0 411900.0 ;
      RECT  115800.0 406950.0 130200.0 406050.0 ;
      RECT  115800.0 420750.0 130200.0 419850.0 ;
      RECT  136800.0 408450.0 138000.0 406500.0 ;
      RECT  136800.0 420300.0 138000.0 418350.0 ;
      RECT  132000.0 418950.0 133200.0 420750.0 ;
      RECT  132000.0 409650.0 133200.0 406050.0 ;
      RECT  134700.0 418950.0 135600.0 409650.0 ;
      RECT  132000.0 409650.0 133200.0 408450.0 ;
      RECT  134400.0 409650.0 135600.0 408450.0 ;
      RECT  134400.0 409650.0 135600.0 408450.0 ;
      RECT  132000.0 409650.0 133200.0 408450.0 ;
      RECT  132000.0 418950.0 133200.0 417750.0 ;
      RECT  134400.0 418950.0 135600.0 417750.0 ;
      RECT  134400.0 418950.0 135600.0 417750.0 ;
      RECT  132000.0 418950.0 133200.0 417750.0 ;
      RECT  136800.0 409050.0 138000.0 407850.0 ;
      RECT  136800.0 418950.0 138000.0 417750.0 ;
      RECT  132600.0 414300.0 133800.0 413100.0 ;
      RECT  132600.0 414300.0 133800.0 413100.0 ;
      RECT  135150.0 414150.0 136050.0 413250.0 ;
      RECT  130200.0 406950.0 139800.0 406050.0 ;
      RECT  130200.0 420750.0 139800.0 419850.0 ;
      RECT  102450.0 413100.0 103650.0 414300.0 ;
      RECT  104400.0 415500.0 105600.0 416700.0 ;
      RECT  121200.0 414600.0 120000.0 415800.0 ;
      RECT  99900.0 203250.0 105000.0 204150.0 ;
      RECT  99900.0 222450.0 105000.0 223350.0 ;
      RECT  99900.0 230850.0 105000.0 231750.0 ;
      RECT  99900.0 250050.0 105000.0 250950.0 ;
      RECT  99900.0 258450.0 105000.0 259350.0 ;
      RECT  99900.0 277650.0 105000.0 278550.0 ;
      RECT  99900.0 286050.0 105000.0 286950.0 ;
      RECT  99900.0 305250.0 105000.0 306150.0 ;
      RECT  99900.0 313650.0 105000.0 314550.0 ;
      RECT  99900.0 332850.0 105000.0 333750.0 ;
      RECT  99900.0 341250.0 105000.0 342150.0 ;
      RECT  99900.0 360450.0 105000.0 361350.0 ;
      RECT  99900.0 368850.0 105000.0 369750.0 ;
      RECT  99900.0 388050.0 105000.0 388950.0 ;
      RECT  99900.0 396450.0 105000.0 397350.0 ;
      RECT  99900.0 415650.0 105000.0 416550.0 ;
      RECT  135150.0 205650.0 136050.0 206550.0 ;
      RECT  135150.0 220050.0 136050.0 220950.0 ;
      RECT  135150.0 233250.0 136050.0 234150.0 ;
      RECT  135150.0 247650.0 136050.0 248550.0 ;
      RECT  135150.0 260850.0 136050.0 261750.0 ;
      RECT  135150.0 275250.0 136050.0 276150.0 ;
      RECT  135150.0 288450.0 136050.0 289350.0 ;
      RECT  135150.0 302850.0 136050.0 303750.0 ;
      RECT  135150.0 316050.0 136050.0 316950.0 ;
      RECT  135150.0 330450.0 136050.0 331350.0 ;
      RECT  135150.0 343650.0 136050.0 344550.0 ;
      RECT  135150.0 358050.0 136050.0 358950.0 ;
      RECT  135150.0 371250.0 136050.0 372150.0 ;
      RECT  135150.0 385650.0 136050.0 386550.0 ;
      RECT  135150.0 398850.0 136050.0 399750.0 ;
      RECT  135150.0 413250.0 136050.0 414150.0 ;
      RECT  99900.0 212850.0 106200.0 213750.0 ;
      RECT  99900.0 240450.0 106200.0 241350.0 ;
      RECT  99900.0 268050.0 106200.0 268950.0 ;
      RECT  99900.0 295650.0 106200.0 296550.0 ;
      RECT  99900.0 323250.0 106200.0 324150.0 ;
      RECT  99900.0 350850.0 106200.0 351750.0 ;
      RECT  99900.0 378450.0 106200.0 379350.0 ;
      RECT  99900.0 406050.0 106200.0 406950.0 ;
      RECT  99900.0 199050.0 106200.0 199950.0 ;
      RECT  99900.0 226650.0 106200.0 227550.0 ;
      RECT  99900.0 254250.0 106200.0 255150.0 ;
      RECT  99900.0 281850.0 106200.0 282750.0 ;
      RECT  99900.0 309450.0 106200.0 310350.0 ;
      RECT  99900.0 337050.0 106200.0 337950.0 ;
      RECT  99900.0 364650.0 106200.0 365550.0 ;
      RECT  99900.0 392250.0 106200.0 393150.0 ;
      RECT  99900.0 419850.0 106200.0 420750.0 ;
      RECT  59100.0 83700.0 119100.0 73500.0 ;
      RECT  59100.0 63300.0 119100.0 73500.0 ;
      RECT  59100.0 63300.0 119100.0 53100.0 ;
      RECT  59100.0 42900.0 119100.0 53100.0 ;
      RECT  61500.0 83700.0 62400.0 42900.0 ;
      RECT  115500.0 83700.0 116400.0 42900.0 ;
      RECT  148050.0 200100.0 149250.0 198900.0 ;
      RECT  148050.0 227700.0 149250.0 226500.0 ;
      RECT  148050.0 255300.0 149250.0 254100.0 ;
      RECT  148050.0 282900.0 149250.0 281700.0 ;
      RECT  148050.0 310500.0 149250.0 309300.0 ;
      RECT  148050.0 338100.0 149250.0 336900.0 ;
      RECT  148050.0 365700.0 149250.0 364500.0 ;
      RECT  148050.0 393300.0 149250.0 392100.0 ;
      RECT  148050.0 420900.0 149250.0 419700.0 ;
      RECT  130500.0 91350.0 129300.0 92550.0 ;
      RECT  135600.0 91200.0 134400.0 92400.0 ;
      RECT  127500.0 105150.0 126300.0 106350.0 ;
      RECT  138300.0 105000.0 137100.0 106200.0 ;
      RECT  130500.0 146550.0 129300.0 147750.0 ;
      RECT  141000.0 146400.0 139800.0 147600.0 ;
      RECT  127500.0 160350.0 126300.0 161550.0 ;
      RECT  143700.0 160200.0 142500.0 161400.0 ;
      RECT  132600.0 88500.0 131400.0 89700.0 ;
      RECT  132600.0 116100.0 131400.0 117300.0 ;
      RECT  132600.0 143700.0 131400.0 144900.0 ;
      RECT  132600.0 171300.0 131400.0 172500.0 ;
      RECT  118500.0 77250.0 117300.0 78450.0 ;
      RECT  135600.0 77250.0 134400.0 78450.0 ;
      RECT  118500.0 68550.0 117300.0 69750.0 ;
      RECT  138300.0 68550.0 137100.0 69750.0 ;
      RECT  118500.0 56850.0 117300.0 58050.0 ;
      RECT  141000.0 56850.0 139800.0 58050.0 ;
      RECT  118500.0 48150.0 117300.0 49350.0 ;
      RECT  143700.0 48150.0 142500.0 49350.0 ;
      RECT  120300.0 72900.0 119100.0 74100.0 ;
      RECT  149250.0 73050.0 148050.0 74250.0 ;
      RECT  120300.0 52500.0 119100.0 53700.0 ;
      RECT  149250.0 52650.0 148050.0 53850.0 ;
      RECT  164400.0 32250.0 163200.0 33450.0 ;
      RECT  159000.0 27750.0 157800.0 28950.0 ;
      RECT  161700.0 25350.0 160500.0 26550.0 ;
      RECT  164400.0 428550.0 163200.0 429750.0 ;
      RECT  167100.0 97050.0 165900.0 98250.0 ;
      RECT  169800.0 195150.0 168600.0 196350.0 ;
      RECT  156300.0 85200.0 155100.0 86400.0 ;
      RECT  103650.0 421800.0 102450.0 423000.0 ;
      RECT  156300.0 421800.0 155100.0 423000.0 ;
      RECT  152550.0 23400.0 151350.0 24600.0 ;
      RECT  152550.0 193200.0 151350.0 194400.0 ;
      RECT  152550.0 95100.0 151350.0 96300.0 ;
      RECT  198600.0 0.0 203100.0 440700.0 ;
      RECT  52800.0 0.0 57300.0 440700.0 ;
      RECT  43650.0 207900.0 42750.0 217500.0 ;
      RECT  43800.0 224100.0 42900.0 225000.0 ;
      RECT  43350.0 224100.0 43200.0 225000.0 ;
      RECT  43800.0 224550.0 42900.0 231900.0 ;
      RECT  43800.0 243750.0 42900.0 251100.0 ;
      RECT  35550.0 258900.0 30600.0 259800.0 ;
      RECT  43650.0 207450.0 42750.0 208350.0 ;
      RECT  43650.0 224100.0 42750.0 225000.0 ;
      RECT  29250.0 362400.0 28350.0 375750.0 ;
      RECT  43800.0 273000.0 42900.0 285150.0 ;
      RECT  33300.0 204900.0 30600.0 205800.0 ;
      RECT  29700.0 285150.0 28800.0 312000.0 ;
      RECT  27000.0 290550.0 26100.0 315000.0 ;
      RECT  41700.0 304050.0 40800.0 312600.0 ;
      RECT  43650.0 301350.0 42750.0 315000.0 ;
      RECT  45600.0 293250.0 44700.0 317400.0 ;
      RECT  41700.0 327150.0 40800.0 328050.0 ;
      RECT  41700.0 318600.0 40800.0 327600.0 ;
      RECT  43200.0 327150.0 41250.0 328050.0 ;
      RECT  43800.0 329550.0 42900.0 330450.0 ;
      RECT  43350.0 329550.0 43200.0 330450.0 ;
      RECT  43800.0 330000.0 42900.0 387600.0 ;
      RECT  14100.0 304050.0 13200.0 322200.0 ;
      RECT  16050.0 293250.0 15150.0 324600.0 ;
      RECT  18000.0 295950.0 17100.0 327000.0 ;
      RECT  14100.0 336750.0 13200.0 337650.0 ;
      RECT  14100.0 328200.0 13200.0 337200.0 ;
      RECT  15600.0 336750.0 13650.0 337650.0 ;
      RECT  16050.0 339600.0 15150.0 346800.0 ;
      RECT  16050.0 349200.0 15150.0 356400.0 ;
      RECT  29250.0 361950.0 28350.0 362850.0 ;
      RECT  28800.0 361950.0 28350.0 362850.0 ;
      RECT  29250.0 360000.0 28350.0 362400.0 ;
      RECT  29250.0 349800.0 28350.0 357000.0 ;
      RECT  29700.0 317100.0 28800.0 323400.0 ;
      RECT  30450.0 333300.0 29550.0 340500.0 ;
      RECT  16050.0 358800.0 15150.0 363000.0 ;
      RECT  29250.0 343200.0 28350.0 347400.0 ;
      RECT  50250.0 202500.0 49350.0 362400.0 ;
      RECT  50250.0 287850.0 49350.0 309000.0 ;
      RECT  36450.0 202500.0 35550.0 362400.0 ;
      RECT  36450.0 298650.0 35550.0 309000.0 ;
      RECT  22650.0 309000.0 21750.0 362400.0 ;
      RECT  22650.0 287850.0 21750.0 309000.0 ;
      RECT  8850.0 309000.0 7950.0 362400.0 ;
      RECT  8850.0 298650.0 7950.0 309000.0 ;
      RECT  8850.0 361950.0 7950.0 362850.0 ;
      RECT  8850.0 360300.0 7950.0 362400.0 ;
      RECT  8400.0 361950.0 3600.0 362850.0 ;
      RECT  7.1054273576e-12 202500.0 10200.0 262500.0 ;
      RECT  20400.0 202500.0 10200.0 262500.0 ;
      RECT  20400.0 202500.0 30600.0 262500.0 ;
      RECT  7.1054273576e-12 204900.0 30600.0 205800.0 ;
      RECT  1.42108547152e-11 258900.0 30600.0 259800.0 ;
      RECT  37950.0 211500.0 36000.0 212700.0 ;
      RECT  49800.0 211500.0 47850.0 212700.0 ;
      RECT  48450.0 207000.0 39150.0 207900.0 ;
      RECT  38550.0 204450.0 36600.0 205350.0 ;
      RECT  38550.0 209250.0 36600.0 210150.0 ;
      RECT  39150.0 204300.0 37950.0 205500.0 ;
      RECT  39150.0 209100.0 37950.0 210300.0 ;
      RECT  39150.0 206700.0 37950.0 207900.0 ;
      RECT  39150.0 206700.0 37950.0 207900.0 ;
      RECT  37050.0 204450.0 36150.0 210150.0 ;
      RECT  49800.0 204450.0 47850.0 205350.0 ;
      RECT  49800.0 209250.0 47850.0 210150.0 ;
      RECT  48450.0 204300.0 47250.0 205500.0 ;
      RECT  48450.0 209100.0 47250.0 210300.0 ;
      RECT  48450.0 206700.0 47250.0 207900.0 ;
      RECT  48450.0 206700.0 47250.0 207900.0 ;
      RECT  50250.0 204450.0 49350.0 210150.0 ;
      RECT  38550.0 211500.0 37350.0 212700.0 ;
      RECT  48450.0 211500.0 47250.0 212700.0 ;
      RECT  43800.0 204900.0 42600.0 206100.0 ;
      RECT  43800.0 204900.0 42600.0 206100.0 ;
      RECT  43650.0 207450.0 42750.0 208350.0 ;
      RECT  36450.0 202500.0 35550.0 214500.0 ;
      RECT  50250.0 202500.0 49350.0 214500.0 ;
      RECT  37950.0 225900.0 36000.0 227100.0 ;
      RECT  49800.0 225900.0 47850.0 227100.0 ;
      RECT  37350.0 216450.0 35550.0 222150.0 ;
      RECT  46050.0 223650.0 41250.0 224550.0 ;
      RECT  38850.0 216450.0 36900.0 217350.0 ;
      RECT  38850.0 221250.0 36900.0 222150.0 ;
      RECT  40800.0 218850.0 38850.0 219750.0 ;
      RECT  40800.0 223650.0 38850.0 224550.0 ;
      RECT  39450.0 216300.0 38250.0 217500.0 ;
      RECT  39450.0 221100.0 38250.0 222300.0 ;
      RECT  39450.0 218700.0 38250.0 219900.0 ;
      RECT  39450.0 223500.0 38250.0 224700.0 ;
      RECT  41250.0 218850.0 40350.0 224550.0 ;
      RECT  37350.0 216450.0 36450.0 222150.0 ;
      RECT  49500.0 216450.0 47550.0 217350.0 ;
      RECT  49500.0 221250.0 47550.0 222150.0 ;
      RECT  47550.0 218850.0 45600.0 219750.0 ;
      RECT  47550.0 223650.0 45600.0 224550.0 ;
      RECT  48150.0 216300.0 46950.0 217500.0 ;
      RECT  48150.0 221100.0 46950.0 222300.0 ;
      RECT  48150.0 218700.0 46950.0 219900.0 ;
      RECT  48150.0 223500.0 46950.0 224700.0 ;
      RECT  46050.0 218850.0 45150.0 224550.0 ;
      RECT  49950.0 216450.0 49050.0 222150.0 ;
      RECT  38550.0 225900.0 37350.0 227100.0 ;
      RECT  48450.0 225900.0 47250.0 227100.0 ;
      RECT  43800.0 216900.0 42600.0 218100.0 ;
      RECT  43800.0 216900.0 42600.0 218100.0 ;
      RECT  43650.0 224100.0 42750.0 225000.0 ;
      RECT  36450.0 214500.0 35550.0 228900.0 ;
      RECT  50250.0 214500.0 49350.0 228900.0 ;
      RECT  37950.0 245100.0 36000.0 246300.0 ;
      RECT  49800.0 245100.0 47850.0 246300.0 ;
      RECT  37800.0 230850.0 35550.0 241350.0 ;
      RECT  45900.0 242850.0 41700.0 243750.0 ;
      RECT  39300.0 230850.0 37350.0 231750.0 ;
      RECT  39300.0 235650.0 37350.0 236550.0 ;
      RECT  39300.0 240450.0 37350.0 241350.0 ;
      RECT  41250.0 233250.0 39300.0 234150.0 ;
      RECT  41250.0 238050.0 39300.0 238950.0 ;
      RECT  41250.0 242850.0 39300.0 243750.0 ;
      RECT  39900.0 230700.0 38700.0 231900.0 ;
      RECT  39900.0 235500.0 38700.0 236700.0 ;
      RECT  39900.0 240300.0 38700.0 241500.0 ;
      RECT  39900.0 233100.0 38700.0 234300.0 ;
      RECT  39900.0 237900.0 38700.0 239100.0 ;
      RECT  39900.0 242700.0 38700.0 243900.0 ;
      RECT  41700.0 233250.0 40800.0 243750.0 ;
      RECT  37800.0 230850.0 36900.0 241350.0 ;
      RECT  49350.0 230850.0 47400.0 231750.0 ;
      RECT  49350.0 235650.0 47400.0 236550.0 ;
      RECT  49350.0 240450.0 47400.0 241350.0 ;
      RECT  47400.0 233250.0 45450.0 234150.0 ;
      RECT  47400.0 238050.0 45450.0 238950.0 ;
      RECT  47400.0 242850.0 45450.0 243750.0 ;
      RECT  48000.0 230700.0 46800.0 231900.0 ;
      RECT  48000.0 235500.0 46800.0 236700.0 ;
      RECT  48000.0 240300.0 46800.0 241500.0 ;
      RECT  48000.0 233100.0 46800.0 234300.0 ;
      RECT  48000.0 237900.0 46800.0 239100.0 ;
      RECT  48000.0 242700.0 46800.0 243900.0 ;
      RECT  45900.0 233250.0 45000.0 243750.0 ;
      RECT  49800.0 230850.0 48900.0 241350.0 ;
      RECT  38550.0 245100.0 37350.0 246300.0 ;
      RECT  48450.0 245100.0 47250.0 246300.0 ;
      RECT  43950.0 231300.0 42750.0 232500.0 ;
      RECT  43950.0 231300.0 42750.0 232500.0 ;
      RECT  43800.0 243300.0 42900.0 244200.0 ;
      RECT  36450.0 228900.0 35550.0 248100.0 ;
      RECT  50250.0 228900.0 49350.0 248100.0 ;
      RECT  37950.0 276300.0 36000.0 277500.0 ;
      RECT  49800.0 276300.0 47850.0 277500.0 ;
      RECT  37800.0 250050.0 35550.0 274950.0 ;
      RECT  45900.0 271650.0 41700.0 272550.0 ;
      RECT  39300.0 250050.0 37350.0 250950.0 ;
      RECT  39300.0 254850.0 37350.0 255750.0 ;
      RECT  39300.0 259650.0 37350.0 260550.0 ;
      RECT  39300.0 264450.0 37350.0 265350.0 ;
      RECT  39300.0 269250.0 37350.0 270150.0 ;
      RECT  39300.0 274050.0 37350.0 274950.0 ;
      RECT  41250.0 252450.0 39300.0 253350.0 ;
      RECT  41250.0 257250.0 39300.0 258150.0 ;
      RECT  41250.0 262050.0 39300.0 262950.0 ;
      RECT  41250.0 266850.0 39300.0 267750.0 ;
      RECT  41250.0 271650.0 39300.0 272550.0 ;
      RECT  39900.0 249900.0 38700.0 251100.0 ;
      RECT  39900.0 254700.0 38700.0 255900.0 ;
      RECT  39900.0 259500.0 38700.0 260700.0 ;
      RECT  39900.0 264300.0 38700.0 265500.0 ;
      RECT  39900.0 269100.0 38700.0 270300.0 ;
      RECT  39900.0 273900.0 38700.0 275100.0 ;
      RECT  39900.0 252300.0 38700.0 253500.0 ;
      RECT  39900.0 257100.0 38700.0 258300.0 ;
      RECT  39900.0 261900.0 38700.0 263100.0 ;
      RECT  39900.0 266700.0 38700.0 267900.0 ;
      RECT  39900.0 271500.0 38700.0 272700.0 ;
      RECT  41700.0 252450.0 40800.0 272550.0 ;
      RECT  37800.0 250050.0 36900.0 274950.0 ;
      RECT  49350.0 250050.0 47400.0 250950.0 ;
      RECT  49350.0 254850.0 47400.0 255750.0 ;
      RECT  49350.0 259650.0 47400.0 260550.0 ;
      RECT  49350.0 264450.0 47400.0 265350.0 ;
      RECT  49350.0 269250.0 47400.0 270150.0 ;
      RECT  49350.0 274050.0 47400.0 274950.0 ;
      RECT  47400.0 252450.0 45450.0 253350.0 ;
      RECT  47400.0 257250.0 45450.0 258150.0 ;
      RECT  47400.0 262050.0 45450.0 262950.0 ;
      RECT  47400.0 266850.0 45450.0 267750.0 ;
      RECT  47400.0 271650.0 45450.0 272550.0 ;
      RECT  48000.0 249900.0 46800.0 251100.0 ;
      RECT  48000.0 254700.0 46800.0 255900.0 ;
      RECT  48000.0 259500.0 46800.0 260700.0 ;
      RECT  48000.0 264300.0 46800.0 265500.0 ;
      RECT  48000.0 269100.0 46800.0 270300.0 ;
      RECT  48000.0 273900.0 46800.0 275100.0 ;
      RECT  48000.0 252300.0 46800.0 253500.0 ;
      RECT  48000.0 257100.0 46800.0 258300.0 ;
      RECT  48000.0 261900.0 46800.0 263100.0 ;
      RECT  48000.0 266700.0 46800.0 267900.0 ;
      RECT  48000.0 271500.0 46800.0 272700.0 ;
      RECT  45900.0 252450.0 45000.0 272550.0 ;
      RECT  49800.0 250050.0 48900.0 274950.0 ;
      RECT  38550.0 276300.0 37350.0 277500.0 ;
      RECT  48450.0 276300.0 47250.0 277500.0 ;
      RECT  43950.0 250500.0 42750.0 251700.0 ;
      RECT  43950.0 250500.0 42750.0 251700.0 ;
      RECT  43800.0 272100.0 42900.0 273000.0 ;
      RECT  36450.0 248100.0 35550.0 279300.0 ;
      RECT  50250.0 248100.0 49350.0 279300.0 ;
      RECT  47850.0 310800.0 50250.0 312000.0 ;
      RECT  39150.0 310800.0 35550.0 312000.0 ;
      RECT  39150.0 315600.0 35550.0 316800.0 ;
      RECT  37950.0 320400.0 36000.0 321600.0 ;
      RECT  49800.0 320400.0 47850.0 321600.0 ;
      RECT  39150.0 310800.0 37950.0 312000.0 ;
      RECT  39150.0 313200.0 37950.0 314400.0 ;
      RECT  39150.0 313200.0 37950.0 314400.0 ;
      RECT  39150.0 310800.0 37950.0 312000.0 ;
      RECT  39150.0 313200.0 37950.0 314400.0 ;
      RECT  39150.0 315600.0 37950.0 316800.0 ;
      RECT  39150.0 315600.0 37950.0 316800.0 ;
      RECT  39150.0 313200.0 37950.0 314400.0 ;
      RECT  39150.0 315600.0 37950.0 316800.0 ;
      RECT  39150.0 318000.0 37950.0 319200.0 ;
      RECT  39150.0 318000.0 37950.0 319200.0 ;
      RECT  39150.0 315600.0 37950.0 316800.0 ;
      RECT  47850.0 310800.0 46650.0 312000.0 ;
      RECT  47850.0 313200.0 46650.0 314400.0 ;
      RECT  47850.0 313200.0 46650.0 314400.0 ;
      RECT  47850.0 310800.0 46650.0 312000.0 ;
      RECT  47850.0 313200.0 46650.0 314400.0 ;
      RECT  47850.0 315600.0 46650.0 316800.0 ;
      RECT  47850.0 315600.0 46650.0 316800.0 ;
      RECT  47850.0 313200.0 46650.0 314400.0 ;
      RECT  47850.0 315600.0 46650.0 316800.0 ;
      RECT  47850.0 318000.0 46650.0 319200.0 ;
      RECT  47850.0 318000.0 46650.0 319200.0 ;
      RECT  47850.0 315600.0 46650.0 316800.0 ;
      RECT  38550.0 320400.0 37350.0 321600.0 ;
      RECT  48450.0 320400.0 47250.0 321600.0 ;
      RECT  45750.0 318000.0 44550.0 316800.0 ;
      RECT  43800.0 315600.0 42600.0 314400.0 ;
      RECT  41850.0 313200.0 40650.0 312000.0 ;
      RECT  39150.0 313200.0 37950.0 314400.0 ;
      RECT  39150.0 318000.0 37950.0 319200.0 ;
      RECT  47850.0 318000.0 46650.0 319200.0 ;
      RECT  41850.0 318000.0 40650.0 319200.0 ;
      RECT  41850.0 312000.0 40650.0 313200.0 ;
      RECT  43800.0 314400.0 42600.0 315600.0 ;
      RECT  45750.0 316800.0 44550.0 318000.0 ;
      RECT  41850.0 318000.0 40650.0 319200.0 ;
      RECT  36450.0 309000.0 35550.0 324600.0 ;
      RECT  50250.0 309000.0 49350.0 324600.0 ;
      RECT  37950.0 331200.0 36000.0 332400.0 ;
      RECT  49800.0 331200.0 47850.0 332400.0 ;
      RECT  48450.0 326400.0 50250.0 327600.0 ;
      RECT  39150.0 326400.0 35550.0 327600.0 ;
      RECT  48450.0 329100.0 39150.0 330000.0 ;
      RECT  39150.0 326400.0 37950.0 327600.0 ;
      RECT  39150.0 328800.0 37950.0 330000.0 ;
      RECT  39150.0 328800.0 37950.0 330000.0 ;
      RECT  39150.0 326400.0 37950.0 327600.0 ;
      RECT  48450.0 326400.0 47250.0 327600.0 ;
      RECT  48450.0 328800.0 47250.0 330000.0 ;
      RECT  48450.0 328800.0 47250.0 330000.0 ;
      RECT  48450.0 326400.0 47250.0 327600.0 ;
      RECT  38550.0 331200.0 37350.0 332400.0 ;
      RECT  48450.0 331200.0 47250.0 332400.0 ;
      RECT  43800.0 327000.0 42600.0 328200.0 ;
      RECT  43800.0 327000.0 42600.0 328200.0 ;
      RECT  43650.0 329550.0 42750.0 330450.0 ;
      RECT  36450.0 324600.0 35550.0 334200.0 ;
      RECT  50250.0 324600.0 49350.0 334200.0 ;
      RECT  23550.0 310800.0 21750.0 312000.0 ;
      RECT  23550.0 315600.0 21750.0 316800.0 ;
      RECT  32250.0 310800.0 36450.0 312000.0 ;
      RECT  34050.0 318000.0 36000.0 319200.0 ;
      RECT  22200.0 318000.0 24150.0 319200.0 ;
      RECT  32250.0 310800.0 33450.0 312000.0 ;
      RECT  32250.0 313200.0 33450.0 314400.0 ;
      RECT  32250.0 313200.0 33450.0 314400.0 ;
      RECT  32250.0 310800.0 33450.0 312000.0 ;
      RECT  32250.0 313200.0 33450.0 314400.0 ;
      RECT  32250.0 315600.0 33450.0 316800.0 ;
      RECT  32250.0 315600.0 33450.0 316800.0 ;
      RECT  32250.0 313200.0 33450.0 314400.0 ;
      RECT  23550.0 310800.0 24750.0 312000.0 ;
      RECT  23550.0 313200.0 24750.0 314400.0 ;
      RECT  23550.0 313200.0 24750.0 314400.0 ;
      RECT  23550.0 310800.0 24750.0 312000.0 ;
      RECT  23550.0 313200.0 24750.0 314400.0 ;
      RECT  23550.0 315600.0 24750.0 316800.0 ;
      RECT  23550.0 315600.0 24750.0 316800.0 ;
      RECT  23550.0 313200.0 24750.0 314400.0 ;
      RECT  33450.0 318000.0 34650.0 319200.0 ;
      RECT  23550.0 318000.0 24750.0 319200.0 ;
      RECT  25950.0 315600.0 27150.0 314400.0 ;
      RECT  28650.0 312600.0 29850.0 311400.0 ;
      RECT  32250.0 315600.0 33450.0 316800.0 ;
      RECT  23550.0 314400.0 24750.0 313200.0 ;
      RECT  28650.0 317700.0 29850.0 316500.0 ;
      RECT  28650.0 311400.0 29850.0 312600.0 ;
      RECT  25950.0 314400.0 27150.0 315600.0 ;
      RECT  28650.0 316500.0 29850.0 317700.0 ;
      RECT  35550.0 309000.0 36450.0 323400.0 ;
      RECT  21750.0 309000.0 22650.0 323400.0 ;
      RECT  24150.0 327900.0 21750.0 329100.0 ;
      RECT  32850.0 327900.0 36450.0 329100.0 ;
      RECT  32850.0 332700.0 36450.0 333900.0 ;
      RECT  34050.0 335100.0 36000.0 336300.0 ;
      RECT  22200.0 335100.0 24150.0 336300.0 ;
      RECT  32850.0 327900.0 34050.0 329100.0 ;
      RECT  32850.0 330300.0 34050.0 331500.0 ;
      RECT  32850.0 330300.0 34050.0 331500.0 ;
      RECT  32850.0 327900.0 34050.0 329100.0 ;
      RECT  32850.0 330300.0 34050.0 331500.0 ;
      RECT  32850.0 332700.0 34050.0 333900.0 ;
      RECT  32850.0 332700.0 34050.0 333900.0 ;
      RECT  32850.0 330300.0 34050.0 331500.0 ;
      RECT  24150.0 327900.0 25350.0 329100.0 ;
      RECT  24150.0 330300.0 25350.0 331500.0 ;
      RECT  24150.0 330300.0 25350.0 331500.0 ;
      RECT  24150.0 327900.0 25350.0 329100.0 ;
      RECT  24150.0 330300.0 25350.0 331500.0 ;
      RECT  24150.0 332700.0 25350.0 333900.0 ;
      RECT  24150.0 332700.0 25350.0 333900.0 ;
      RECT  24150.0 330300.0 25350.0 331500.0 ;
      RECT  33450.0 335100.0 34650.0 336300.0 ;
      RECT  23550.0 335100.0 24750.0 336300.0 ;
      RECT  26700.0 332700.0 27900.0 331500.0 ;
      RECT  29400.0 329700.0 30600.0 328500.0 ;
      RECT  32850.0 330300.0 34050.0 331500.0 ;
      RECT  24150.0 332700.0 25350.0 333900.0 ;
      RECT  29400.0 333900.0 30600.0 332700.0 ;
      RECT  29400.0 328500.0 30600.0 329700.0 ;
      RECT  26700.0 331500.0 27900.0 332700.0 ;
      RECT  29400.0 332700.0 30600.0 333900.0 ;
      RECT  35550.0 326100.0 36450.0 340500.0 ;
      RECT  21750.0 326100.0 22650.0 340500.0 ;
      RECT  34050.0 346200.0 36000.0 345000.0 ;
      RECT  22200.0 346200.0 24150.0 345000.0 ;
      RECT  23550.0 351000.0 21750.0 349800.0 ;
      RECT  32850.0 351000.0 36450.0 349800.0 ;
      RECT  23550.0 348300.0 32850.0 347400.0 ;
      RECT  32850.0 351000.0 34050.0 349800.0 ;
      RECT  32850.0 348600.0 34050.0 347400.0 ;
      RECT  32850.0 348600.0 34050.0 347400.0 ;
      RECT  32850.0 351000.0 34050.0 349800.0 ;
      RECT  23550.0 351000.0 24750.0 349800.0 ;
      RECT  23550.0 348600.0 24750.0 347400.0 ;
      RECT  23550.0 348600.0 24750.0 347400.0 ;
      RECT  23550.0 351000.0 24750.0 349800.0 ;
      RECT  33450.0 346200.0 34650.0 345000.0 ;
      RECT  23550.0 346200.0 24750.0 345000.0 ;
      RECT  28200.0 350400.0 29400.0 349200.0 ;
      RECT  28200.0 350400.0 29400.0 349200.0 ;
      RECT  28350.0 347850.0 29250.0 346950.0 ;
      RECT  35550.0 352800.0 36450.0 343200.0 ;
      RECT  21750.0 352800.0 22650.0 343200.0 ;
      RECT  34050.0 355800.0 36000.0 354600.0 ;
      RECT  22200.0 355800.0 24150.0 354600.0 ;
      RECT  23550.0 360600.0 21750.0 359400.0 ;
      RECT  32850.0 360600.0 36450.0 359400.0 ;
      RECT  23550.0 357900.0 32850.0 357000.0 ;
      RECT  32850.0 360600.0 34050.0 359400.0 ;
      RECT  32850.0 358200.0 34050.0 357000.0 ;
      RECT  32850.0 358200.0 34050.0 357000.0 ;
      RECT  32850.0 360600.0 34050.0 359400.0 ;
      RECT  23550.0 360600.0 24750.0 359400.0 ;
      RECT  23550.0 358200.0 24750.0 357000.0 ;
      RECT  23550.0 358200.0 24750.0 357000.0 ;
      RECT  23550.0 360600.0 24750.0 359400.0 ;
      RECT  33450.0 355800.0 34650.0 354600.0 ;
      RECT  23550.0 355800.0 24750.0 354600.0 ;
      RECT  28200.0 360000.0 29400.0 358800.0 ;
      RECT  28200.0 360000.0 29400.0 358800.0 ;
      RECT  28350.0 357450.0 29250.0 356550.0 ;
      RECT  35550.0 362400.0 36450.0 352800.0 ;
      RECT  21750.0 362400.0 22650.0 352800.0 ;
      RECT  20250.0 320400.0 22650.0 321600.0 ;
      RECT  11550.0 320400.0 7950.0 321600.0 ;
      RECT  11550.0 325200.0 7950.0 326400.0 ;
      RECT  10350.0 330000.0 8400.0 331200.0 ;
      RECT  22200.0 330000.0 20250.0 331200.0 ;
      RECT  11550.0 320400.0 10350.0 321600.0 ;
      RECT  11550.0 322800.0 10350.0 324000.0 ;
      RECT  11550.0 322800.0 10350.0 324000.0 ;
      RECT  11550.0 320400.0 10350.0 321600.0 ;
      RECT  11550.0 322800.0 10350.0 324000.0 ;
      RECT  11550.0 325200.0 10350.0 326400.0 ;
      RECT  11550.0 325200.0 10350.0 326400.0 ;
      RECT  11550.0 322800.0 10350.0 324000.0 ;
      RECT  11550.0 325200.0 10350.0 326400.0 ;
      RECT  11550.0 327600.0 10350.0 328800.0 ;
      RECT  11550.0 327600.0 10350.0 328800.0 ;
      RECT  11550.0 325200.0 10350.0 326400.0 ;
      RECT  20250.0 320400.0 19050.0 321600.0 ;
      RECT  20250.0 322800.0 19050.0 324000.0 ;
      RECT  20250.0 322800.0 19050.0 324000.0 ;
      RECT  20250.0 320400.0 19050.0 321600.0 ;
      RECT  20250.0 322800.0 19050.0 324000.0 ;
      RECT  20250.0 325200.0 19050.0 326400.0 ;
      RECT  20250.0 325200.0 19050.0 326400.0 ;
      RECT  20250.0 322800.0 19050.0 324000.0 ;
      RECT  20250.0 325200.0 19050.0 326400.0 ;
      RECT  20250.0 327600.0 19050.0 328800.0 ;
      RECT  20250.0 327600.0 19050.0 328800.0 ;
      RECT  20250.0 325200.0 19050.0 326400.0 ;
      RECT  10950.0 330000.0 9750.0 331200.0 ;
      RECT  20850.0 330000.0 19650.0 331200.0 ;
      RECT  18150.0 327600.0 16950.0 326400.0 ;
      RECT  16200.0 325200.0 15000.0 324000.0 ;
      RECT  14250.0 322800.0 13050.0 321600.0 ;
      RECT  11550.0 322800.0 10350.0 324000.0 ;
      RECT  11550.0 327600.0 10350.0 328800.0 ;
      RECT  20250.0 327600.0 19050.0 328800.0 ;
      RECT  14250.0 327600.0 13050.0 328800.0 ;
      RECT  14250.0 321600.0 13050.0 322800.0 ;
      RECT  16200.0 324000.0 15000.0 325200.0 ;
      RECT  18150.0 326400.0 16950.0 327600.0 ;
      RECT  14250.0 327600.0 13050.0 328800.0 ;
      RECT  8850.0 318600.0 7950.0 334200.0 ;
      RECT  22650.0 318600.0 21750.0 334200.0 ;
      RECT  10350.0 340800.0 8400.0 342000.0 ;
      RECT  22200.0 340800.0 20250.0 342000.0 ;
      RECT  20850.0 336000.0 22650.0 337200.0 ;
      RECT  11550.0 336000.0 7950.0 337200.0 ;
      RECT  20850.0 338700.0 11550.0 339600.0 ;
      RECT  11550.0 336000.0 10350.0 337200.0 ;
      RECT  11550.0 338400.0 10350.0 339600.0 ;
      RECT  11550.0 338400.0 10350.0 339600.0 ;
      RECT  11550.0 336000.0 10350.0 337200.0 ;
      RECT  20850.0 336000.0 19650.0 337200.0 ;
      RECT  20850.0 338400.0 19650.0 339600.0 ;
      RECT  20850.0 338400.0 19650.0 339600.0 ;
      RECT  20850.0 336000.0 19650.0 337200.0 ;
      RECT  10950.0 340800.0 9750.0 342000.0 ;
      RECT  20850.0 340800.0 19650.0 342000.0 ;
      RECT  16200.0 336600.0 15000.0 337800.0 ;
      RECT  16200.0 336600.0 15000.0 337800.0 ;
      RECT  16050.0 339150.0 15150.0 340050.0 ;
      RECT  8850.0 334200.0 7950.0 343800.0 ;
      RECT  22650.0 334200.0 21750.0 343800.0 ;
      RECT  10350.0 350400.0 8400.0 351600.0 ;
      RECT  22200.0 350400.0 20250.0 351600.0 ;
      RECT  20850.0 345600.0 22650.0 346800.0 ;
      RECT  11550.0 345600.0 7950.0 346800.0 ;
      RECT  20850.0 348300.0 11550.0 349200.0 ;
      RECT  11550.0 345600.0 10350.0 346800.0 ;
      RECT  11550.0 348000.0 10350.0 349200.0 ;
      RECT  11550.0 348000.0 10350.0 349200.0 ;
      RECT  11550.0 345600.0 10350.0 346800.0 ;
      RECT  20850.0 345600.0 19650.0 346800.0 ;
      RECT  20850.0 348000.0 19650.0 349200.0 ;
      RECT  20850.0 348000.0 19650.0 349200.0 ;
      RECT  20850.0 345600.0 19650.0 346800.0 ;
      RECT  10950.0 350400.0 9750.0 351600.0 ;
      RECT  20850.0 350400.0 19650.0 351600.0 ;
      RECT  16200.0 346200.0 15000.0 347400.0 ;
      RECT  16200.0 346200.0 15000.0 347400.0 ;
      RECT  16050.0 348750.0 15150.0 349650.0 ;
      RECT  8850.0 343800.0 7950.0 353400.0 ;
      RECT  22650.0 343800.0 21750.0 353400.0 ;
      RECT  10350.0 360000.0 8400.0 361200.0 ;
      RECT  22200.0 360000.0 20250.0 361200.0 ;
      RECT  20850.0 355200.0 22650.0 356400.0 ;
      RECT  11550.0 355200.0 7950.0 356400.0 ;
      RECT  20850.0 357900.0 11550.0 358800.0 ;
      RECT  11550.0 355200.0 10350.0 356400.0 ;
      RECT  11550.0 357600.0 10350.0 358800.0 ;
      RECT  11550.0 357600.0 10350.0 358800.0 ;
      RECT  11550.0 355200.0 10350.0 356400.0 ;
      RECT  20850.0 355200.0 19650.0 356400.0 ;
      RECT  20850.0 357600.0 19650.0 358800.0 ;
      RECT  20850.0 357600.0 19650.0 358800.0 ;
      RECT  20850.0 355200.0 19650.0 356400.0 ;
      RECT  10950.0 360000.0 9750.0 361200.0 ;
      RECT  20850.0 360000.0 19650.0 361200.0 ;
      RECT  16200.0 355800.0 15000.0 357000.0 ;
      RECT  16200.0 355800.0 15000.0 357000.0 ;
      RECT  16050.0 358350.0 15150.0 359250.0 ;
      RECT  8850.0 353400.0 7950.0 363000.0 ;
      RECT  22650.0 353400.0 21750.0 363000.0 ;
      RECT  22650.0 499050.0 21750.0 430200.0 ;
      RECT  21750.0 397050.0 17400.0 397950.0 ;
      RECT  21750.0 420450.0 17400.0 421350.0 ;
      RECT  22650.0 371550.0 16800.0 372450.0 ;
      RECT  16800.0 371550.0 6600.0 372450.0 ;
      RECT  4500.0 408600.0 16800.0 409500.0 ;
      RECT  4500.0 381000.0 16800.0 381900.0 ;
      RECT  29250.0 397800.0 28350.0 410400.0 ;
      RECT  29250.0 392850.0 28350.0 393750.0 ;
      RECT  29250.0 393300.0 28350.0 397800.0 ;
      RECT  28800.0 392850.0 17400.0 393750.0 ;
      RECT  36000.0 398550.0 33750.0 399450.0 ;
      RECT  33600.0 383850.0 32700.0 384750.0 ;
      RECT  29250.0 383850.0 28350.0 384750.0 ;
      RECT  33600.0 384300.0 32700.0 396000.0 ;
      RECT  33150.0 383850.0 28800.0 384750.0 ;
      RECT  29250.0 379200.0 28350.0 384300.0 ;
      RECT  28800.0 383850.0 19950.0 384750.0 ;
      RECT  19950.0 375750.0 13200.0 376650.0 ;
      RECT  29400.0 378000.0 28200.0 379200.0 ;
      RECT  29250.0 410400.0 28350.0 414150.0 ;
      RECT  34050.0 375000.0 36000.0 373800.0 ;
      RECT  22200.0 375000.0 24150.0 373800.0 ;
      RECT  23550.0 379800.0 21750.0 378600.0 ;
      RECT  32850.0 379800.0 36450.0 378600.0 ;
      RECT  23550.0 377100.0 32850.0 376200.0 ;
      RECT  32850.0 379800.0 34050.0 378600.0 ;
      RECT  32850.0 377400.0 34050.0 376200.0 ;
      RECT  32850.0 377400.0 34050.0 376200.0 ;
      RECT  32850.0 379800.0 34050.0 378600.0 ;
      RECT  23550.0 379800.0 24750.0 378600.0 ;
      RECT  23550.0 377400.0 24750.0 376200.0 ;
      RECT  23550.0 377400.0 24750.0 376200.0 ;
      RECT  23550.0 379800.0 24750.0 378600.0 ;
      RECT  33450.0 375000.0 34650.0 373800.0 ;
      RECT  23550.0 375000.0 24750.0 373800.0 ;
      RECT  28200.0 379200.0 29400.0 378000.0 ;
      RECT  28200.0 379200.0 29400.0 378000.0 ;
      RECT  28350.0 376650.0 29250.0 375750.0 ;
      RECT  35550.0 381600.0 36450.0 372000.0 ;
      RECT  21750.0 381600.0 22650.0 372000.0 ;
      RECT  32550.0 396000.0 33750.0 397200.0 ;
      RECT  32550.0 398400.0 33750.0 399600.0 ;
      RECT  32550.0 398400.0 33750.0 399600.0 ;
      RECT  32550.0 396000.0 33750.0 397200.0 ;
      RECT  21750.0 498150.0 22650.0 499050.0 ;
      RECT  49350.0 498150.0 50250.0 499050.0 ;
      RECT  21750.0 496800.0 22650.0 498600.0 ;
      RECT  22200.0 498150.0 49800.0 499050.0 ;
      RECT  49350.0 496800.0 50250.0 498600.0 ;
      RECT  37950.0 417000.0 36000.0 418200.0 ;
      RECT  49800.0 417000.0 47850.0 418200.0 ;
      RECT  48450.0 412200.0 50250.0 413400.0 ;
      RECT  39150.0 412200.0 35550.0 413400.0 ;
      RECT  48450.0 414900.0 39150.0 415800.0 ;
      RECT  39150.0 412200.0 37950.0 413400.0 ;
      RECT  39150.0 414600.0 37950.0 415800.0 ;
      RECT  39150.0 414600.0 37950.0 415800.0 ;
      RECT  39150.0 412200.0 37950.0 413400.0 ;
      RECT  48450.0 412200.0 47250.0 413400.0 ;
      RECT  48450.0 414600.0 47250.0 415800.0 ;
      RECT  48450.0 414600.0 47250.0 415800.0 ;
      RECT  48450.0 412200.0 47250.0 413400.0 ;
      RECT  38550.0 417000.0 37350.0 418200.0 ;
      RECT  48450.0 417000.0 47250.0 418200.0 ;
      RECT  43800.0 412800.0 42600.0 414000.0 ;
      RECT  43800.0 412800.0 42600.0 414000.0 ;
      RECT  43650.0 415350.0 42750.0 416250.0 ;
      RECT  36450.0 410400.0 35550.0 420000.0 ;
      RECT  50250.0 410400.0 49350.0 420000.0 ;
      RECT  37950.0 426600.0 36000.0 427800.0 ;
      RECT  49800.0 426600.0 47850.0 427800.0 ;
      RECT  48450.0 421800.0 50250.0 423000.0 ;
      RECT  39150.0 421800.0 35550.0 423000.0 ;
      RECT  48450.0 424500.0 39150.0 425400.0 ;
      RECT  39150.0 421800.0 37950.0 423000.0 ;
      RECT  39150.0 424200.0 37950.0 425400.0 ;
      RECT  39150.0 424200.0 37950.0 425400.0 ;
      RECT  39150.0 421800.0 37950.0 423000.0 ;
      RECT  48450.0 421800.0 47250.0 423000.0 ;
      RECT  48450.0 424200.0 47250.0 425400.0 ;
      RECT  48450.0 424200.0 47250.0 425400.0 ;
      RECT  48450.0 421800.0 47250.0 423000.0 ;
      RECT  38550.0 426600.0 37350.0 427800.0 ;
      RECT  48450.0 426600.0 47250.0 427800.0 ;
      RECT  43800.0 422400.0 42600.0 423600.0 ;
      RECT  43800.0 422400.0 42600.0 423600.0 ;
      RECT  43650.0 424950.0 42750.0 425850.0 ;
      RECT  36450.0 420000.0 35550.0 429600.0 ;
      RECT  50250.0 420000.0 49350.0 429600.0 ;
      RECT  42600.0 422400.0 43800.0 423600.0 ;
      RECT  37950.0 436200.0 36000.0 437400.0 ;
      RECT  49800.0 436200.0 47850.0 437400.0 ;
      RECT  48450.0 431400.0 50250.0 432600.0 ;
      RECT  39150.0 431400.0 35550.0 432600.0 ;
      RECT  48450.0 434100.0 39150.0 435000.0 ;
      RECT  39150.0 431400.0 37950.0 432600.0 ;
      RECT  39150.0 433800.0 37950.0 435000.0 ;
      RECT  39150.0 433800.0 37950.0 435000.0 ;
      RECT  39150.0 431400.0 37950.0 432600.0 ;
      RECT  48450.0 431400.0 47250.0 432600.0 ;
      RECT  48450.0 433800.0 47250.0 435000.0 ;
      RECT  48450.0 433800.0 47250.0 435000.0 ;
      RECT  48450.0 431400.0 47250.0 432600.0 ;
      RECT  38550.0 436200.0 37350.0 437400.0 ;
      RECT  48450.0 436200.0 47250.0 437400.0 ;
      RECT  43800.0 432000.0 42600.0 433200.0 ;
      RECT  43800.0 432000.0 42600.0 433200.0 ;
      RECT  43650.0 434550.0 42750.0 435450.0 ;
      RECT  36450.0 429600.0 35550.0 439200.0 ;
      RECT  50250.0 429600.0 49350.0 439200.0 ;
      RECT  42600.0 432000.0 43800.0 433200.0 ;
      RECT  37950.0 445800.0 36000.0 447000.0 ;
      RECT  49800.0 445800.0 47850.0 447000.0 ;
      RECT  48450.0 441000.0 50250.0 442200.0 ;
      RECT  39150.0 441000.0 35550.0 442200.0 ;
      RECT  48450.0 443700.0 39150.0 444600.0 ;
      RECT  39150.0 441000.0 37950.0 442200.0 ;
      RECT  39150.0 443400.0 37950.0 444600.0 ;
      RECT  39150.0 443400.0 37950.0 444600.0 ;
      RECT  39150.0 441000.0 37950.0 442200.0 ;
      RECT  48450.0 441000.0 47250.0 442200.0 ;
      RECT  48450.0 443400.0 47250.0 444600.0 ;
      RECT  48450.0 443400.0 47250.0 444600.0 ;
      RECT  48450.0 441000.0 47250.0 442200.0 ;
      RECT  38550.0 445800.0 37350.0 447000.0 ;
      RECT  48450.0 445800.0 47250.0 447000.0 ;
      RECT  43800.0 441600.0 42600.0 442800.0 ;
      RECT  43800.0 441600.0 42600.0 442800.0 ;
      RECT  43650.0 444150.0 42750.0 445050.0 ;
      RECT  36450.0 439200.0 35550.0 448800.0 ;
      RECT  50250.0 439200.0 49350.0 448800.0 ;
      RECT  42600.0 441600.0 43800.0 442800.0 ;
      RECT  37950.0 455400.0 36000.0 456600.0 ;
      RECT  49800.0 455400.0 47850.0 456600.0 ;
      RECT  48450.0 450600.0 50250.0 451800.0 ;
      RECT  39150.0 450600.0 35550.0 451800.0 ;
      RECT  48450.0 453300.0 39150.0 454200.0 ;
      RECT  39150.0 450600.0 37950.0 451800.0 ;
      RECT  39150.0 453000.0 37950.0 454200.0 ;
      RECT  39150.0 453000.0 37950.0 454200.0 ;
      RECT  39150.0 450600.0 37950.0 451800.0 ;
      RECT  48450.0 450600.0 47250.0 451800.0 ;
      RECT  48450.0 453000.0 47250.0 454200.0 ;
      RECT  48450.0 453000.0 47250.0 454200.0 ;
      RECT  48450.0 450600.0 47250.0 451800.0 ;
      RECT  38550.0 455400.0 37350.0 456600.0 ;
      RECT  48450.0 455400.0 47250.0 456600.0 ;
      RECT  43800.0 451200.0 42600.0 452400.0 ;
      RECT  43800.0 451200.0 42600.0 452400.0 ;
      RECT  43650.0 453750.0 42750.0 454650.0 ;
      RECT  36450.0 448800.0 35550.0 458400.0 ;
      RECT  50250.0 448800.0 49350.0 458400.0 ;
      RECT  42600.0 451200.0 43800.0 452400.0 ;
      RECT  37950.0 465000.0 36000.0 466200.0 ;
      RECT  49800.0 465000.0 47850.0 466200.0 ;
      RECT  48450.0 460200.0 50250.0 461400.0 ;
      RECT  39150.0 460200.0 35550.0 461400.0 ;
      RECT  48450.0 462900.0 39150.0 463800.0 ;
      RECT  39150.0 460200.0 37950.0 461400.0 ;
      RECT  39150.0 462600.0 37950.0 463800.0 ;
      RECT  39150.0 462600.0 37950.0 463800.0 ;
      RECT  39150.0 460200.0 37950.0 461400.0 ;
      RECT  48450.0 460200.0 47250.0 461400.0 ;
      RECT  48450.0 462600.0 47250.0 463800.0 ;
      RECT  48450.0 462600.0 47250.0 463800.0 ;
      RECT  48450.0 460200.0 47250.0 461400.0 ;
      RECT  38550.0 465000.0 37350.0 466200.0 ;
      RECT  48450.0 465000.0 47250.0 466200.0 ;
      RECT  43800.0 460800.0 42600.0 462000.0 ;
      RECT  43800.0 460800.0 42600.0 462000.0 ;
      RECT  43650.0 463350.0 42750.0 464250.0 ;
      RECT  36450.0 458400.0 35550.0 468000.0 ;
      RECT  50250.0 458400.0 49350.0 468000.0 ;
      RECT  42600.0 460800.0 43800.0 462000.0 ;
      RECT  37950.0 474600.0 36000.0 475800.0 ;
      RECT  49800.0 474600.0 47850.0 475800.0 ;
      RECT  48450.0 469800.0 50250.0 471000.0 ;
      RECT  39150.0 469800.0 35550.0 471000.0 ;
      RECT  48450.0 472500.0 39150.0 473400.0 ;
      RECT  39150.0 469800.0 37950.0 471000.0 ;
      RECT  39150.0 472200.0 37950.0 473400.0 ;
      RECT  39150.0 472200.0 37950.0 473400.0 ;
      RECT  39150.0 469800.0 37950.0 471000.0 ;
      RECT  48450.0 469800.0 47250.0 471000.0 ;
      RECT  48450.0 472200.0 47250.0 473400.0 ;
      RECT  48450.0 472200.0 47250.0 473400.0 ;
      RECT  48450.0 469800.0 47250.0 471000.0 ;
      RECT  38550.0 474600.0 37350.0 475800.0 ;
      RECT  48450.0 474600.0 47250.0 475800.0 ;
      RECT  43800.0 470400.0 42600.0 471600.0 ;
      RECT  43800.0 470400.0 42600.0 471600.0 ;
      RECT  43650.0 472950.0 42750.0 473850.0 ;
      RECT  36450.0 468000.0 35550.0 477600.0 ;
      RECT  50250.0 468000.0 49350.0 477600.0 ;
      RECT  42600.0 470400.0 43800.0 471600.0 ;
      RECT  37950.0 484200.0 36000.0 485400.0 ;
      RECT  49800.0 484200.0 47850.0 485400.0 ;
      RECT  48450.0 479400.0 50250.0 480600.0 ;
      RECT  39150.0 479400.0 35550.0 480600.0 ;
      RECT  48450.0 482100.0 39150.0 483000.0 ;
      RECT  39150.0 479400.0 37950.0 480600.0 ;
      RECT  39150.0 481800.0 37950.0 483000.0 ;
      RECT  39150.0 481800.0 37950.0 483000.0 ;
      RECT  39150.0 479400.0 37950.0 480600.0 ;
      RECT  48450.0 479400.0 47250.0 480600.0 ;
      RECT  48450.0 481800.0 47250.0 483000.0 ;
      RECT  48450.0 481800.0 47250.0 483000.0 ;
      RECT  48450.0 479400.0 47250.0 480600.0 ;
      RECT  38550.0 484200.0 37350.0 485400.0 ;
      RECT  48450.0 484200.0 47250.0 485400.0 ;
      RECT  43800.0 480000.0 42600.0 481200.0 ;
      RECT  43800.0 480000.0 42600.0 481200.0 ;
      RECT  43650.0 482550.0 42750.0 483450.0 ;
      RECT  36450.0 477600.0 35550.0 487200.0 ;
      RECT  50250.0 477600.0 49350.0 487200.0 ;
      RECT  42600.0 480000.0 43800.0 481200.0 ;
      RECT  37950.0 493800.0 36000.0 495000.0 ;
      RECT  49800.0 493800.0 47850.0 495000.0 ;
      RECT  48450.0 489000.0 50250.0 490200.0 ;
      RECT  39150.0 489000.0 35550.0 490200.0 ;
      RECT  48450.0 491700.0 39150.0 492600.0 ;
      RECT  39150.0 489000.0 37950.0 490200.0 ;
      RECT  39150.0 491400.0 37950.0 492600.0 ;
      RECT  39150.0 491400.0 37950.0 492600.0 ;
      RECT  39150.0 489000.0 37950.0 490200.0 ;
      RECT  48450.0 489000.0 47250.0 490200.0 ;
      RECT  48450.0 491400.0 47250.0 492600.0 ;
      RECT  48450.0 491400.0 47250.0 492600.0 ;
      RECT  48450.0 489000.0 47250.0 490200.0 ;
      RECT  38550.0 493800.0 37350.0 495000.0 ;
      RECT  48450.0 493800.0 47250.0 495000.0 ;
      RECT  43800.0 489600.0 42600.0 490800.0 ;
      RECT  43800.0 489600.0 42600.0 490800.0 ;
      RECT  43650.0 492150.0 42750.0 493050.0 ;
      RECT  36450.0 487200.0 35550.0 496800.0 ;
      RECT  50250.0 487200.0 49350.0 496800.0 ;
      RECT  42600.0 489600.0 43800.0 490800.0 ;
      RECT  34050.0 480600.0 36000.0 479400.0 ;
      RECT  22200.0 480600.0 24150.0 479400.0 ;
      RECT  23550.0 485400.0 21750.0 484200.0 ;
      RECT  32850.0 485400.0 36450.0 484200.0 ;
      RECT  23550.0 482700.0 32850.0 481800.0 ;
      RECT  32850.0 485400.0 34050.0 484200.0 ;
      RECT  32850.0 483000.0 34050.0 481800.0 ;
      RECT  32850.0 483000.0 34050.0 481800.0 ;
      RECT  32850.0 485400.0 34050.0 484200.0 ;
      RECT  23550.0 485400.0 24750.0 484200.0 ;
      RECT  23550.0 483000.0 24750.0 481800.0 ;
      RECT  23550.0 483000.0 24750.0 481800.0 ;
      RECT  23550.0 485400.0 24750.0 484200.0 ;
      RECT  33450.0 480600.0 34650.0 479400.0 ;
      RECT  23550.0 480600.0 24750.0 479400.0 ;
      RECT  28200.0 484800.0 29400.0 483600.0 ;
      RECT  28200.0 484800.0 29400.0 483600.0 ;
      RECT  28350.0 482250.0 29250.0 481350.0 ;
      RECT  35550.0 487200.0 36450.0 477600.0 ;
      RECT  21750.0 487200.0 22650.0 477600.0 ;
      RECT  28200.0 483600.0 29400.0 484800.0 ;
      RECT  34050.0 471000.0 36000.0 469800.0 ;
      RECT  22200.0 471000.0 24150.0 469800.0 ;
      RECT  23550.0 475800.0 21750.0 474600.0 ;
      RECT  32850.0 475800.0 36450.0 474600.0 ;
      RECT  23550.0 473100.0 32850.0 472200.0 ;
      RECT  32850.0 475800.0 34050.0 474600.0 ;
      RECT  32850.0 473400.0 34050.0 472200.0 ;
      RECT  32850.0 473400.0 34050.0 472200.0 ;
      RECT  32850.0 475800.0 34050.0 474600.0 ;
      RECT  23550.0 475800.0 24750.0 474600.0 ;
      RECT  23550.0 473400.0 24750.0 472200.0 ;
      RECT  23550.0 473400.0 24750.0 472200.0 ;
      RECT  23550.0 475800.0 24750.0 474600.0 ;
      RECT  33450.0 471000.0 34650.0 469800.0 ;
      RECT  23550.0 471000.0 24750.0 469800.0 ;
      RECT  28200.0 475200.0 29400.0 474000.0 ;
      RECT  28200.0 475200.0 29400.0 474000.0 ;
      RECT  28350.0 472650.0 29250.0 471750.0 ;
      RECT  35550.0 477600.0 36450.0 468000.0 ;
      RECT  21750.0 477600.0 22650.0 468000.0 ;
      RECT  28200.0 474000.0 29400.0 475200.0 ;
      RECT  34050.0 461400.0 36000.0 460200.0 ;
      RECT  22200.0 461400.0 24150.0 460200.0 ;
      RECT  23550.0 466200.0 21750.0 465000.0 ;
      RECT  32850.0 466200.0 36450.0 465000.0 ;
      RECT  23550.0 463500.0 32850.0 462600.0 ;
      RECT  32850.0 466200.0 34050.0 465000.0 ;
      RECT  32850.0 463800.0 34050.0 462600.0 ;
      RECT  32850.0 463800.0 34050.0 462600.0 ;
      RECT  32850.0 466200.0 34050.0 465000.0 ;
      RECT  23550.0 466200.0 24750.0 465000.0 ;
      RECT  23550.0 463800.0 24750.0 462600.0 ;
      RECT  23550.0 463800.0 24750.0 462600.0 ;
      RECT  23550.0 466200.0 24750.0 465000.0 ;
      RECT  33450.0 461400.0 34650.0 460200.0 ;
      RECT  23550.0 461400.0 24750.0 460200.0 ;
      RECT  28200.0 465600.0 29400.0 464400.0 ;
      RECT  28200.0 465600.0 29400.0 464400.0 ;
      RECT  28350.0 463050.0 29250.0 462150.0 ;
      RECT  35550.0 468000.0 36450.0 458400.0 ;
      RECT  21750.0 468000.0 22650.0 458400.0 ;
      RECT  28200.0 464400.0 29400.0 465600.0 ;
      RECT  34050.0 451800.0 36000.0 450600.0 ;
      RECT  22200.0 451800.0 24150.0 450600.0 ;
      RECT  23550.0 456600.0 21750.0 455400.0 ;
      RECT  32850.0 456600.0 36450.0 455400.0 ;
      RECT  23550.0 453900.0 32850.0 453000.0 ;
      RECT  32850.0 456600.0 34050.0 455400.0 ;
      RECT  32850.0 454200.0 34050.0 453000.0 ;
      RECT  32850.0 454200.0 34050.0 453000.0 ;
      RECT  32850.0 456600.0 34050.0 455400.0 ;
      RECT  23550.0 456600.0 24750.0 455400.0 ;
      RECT  23550.0 454200.0 24750.0 453000.0 ;
      RECT  23550.0 454200.0 24750.0 453000.0 ;
      RECT  23550.0 456600.0 24750.0 455400.0 ;
      RECT  33450.0 451800.0 34650.0 450600.0 ;
      RECT  23550.0 451800.0 24750.0 450600.0 ;
      RECT  28200.0 456000.0 29400.0 454800.0 ;
      RECT  28200.0 456000.0 29400.0 454800.0 ;
      RECT  28350.0 453450.0 29250.0 452550.0 ;
      RECT  35550.0 458400.0 36450.0 448800.0 ;
      RECT  21750.0 458400.0 22650.0 448800.0 ;
      RECT  28200.0 454800.0 29400.0 456000.0 ;
      RECT  34050.0 442200.0 36000.0 441000.0 ;
      RECT  22200.0 442200.0 24150.0 441000.0 ;
      RECT  23550.0 447000.0 21750.0 445800.0 ;
      RECT  32850.0 447000.0 36450.0 445800.0 ;
      RECT  23550.0 444300.0 32850.0 443400.0 ;
      RECT  32850.0 447000.0 34050.0 445800.0 ;
      RECT  32850.0 444600.0 34050.0 443400.0 ;
      RECT  32850.0 444600.0 34050.0 443400.0 ;
      RECT  32850.0 447000.0 34050.0 445800.0 ;
      RECT  23550.0 447000.0 24750.0 445800.0 ;
      RECT  23550.0 444600.0 24750.0 443400.0 ;
      RECT  23550.0 444600.0 24750.0 443400.0 ;
      RECT  23550.0 447000.0 24750.0 445800.0 ;
      RECT  33450.0 442200.0 34650.0 441000.0 ;
      RECT  23550.0 442200.0 24750.0 441000.0 ;
      RECT  28200.0 446400.0 29400.0 445200.0 ;
      RECT  28200.0 446400.0 29400.0 445200.0 ;
      RECT  28350.0 443850.0 29250.0 442950.0 ;
      RECT  35550.0 448800.0 36450.0 439200.0 ;
      RECT  21750.0 448800.0 22650.0 439200.0 ;
      RECT  28200.0 445200.0 29400.0 446400.0 ;
      RECT  34050.0 432600.0 36000.0 431400.0 ;
      RECT  22200.0 432600.0 24150.0 431400.0 ;
      RECT  23550.0 437400.0 21750.0 436200.0 ;
      RECT  32850.0 437400.0 36450.0 436200.0 ;
      RECT  23550.0 434700.0 32850.0 433800.0 ;
      RECT  32850.0 437400.0 34050.0 436200.0 ;
      RECT  32850.0 435000.0 34050.0 433800.0 ;
      RECT  32850.0 435000.0 34050.0 433800.0 ;
      RECT  32850.0 437400.0 34050.0 436200.0 ;
      RECT  23550.0 437400.0 24750.0 436200.0 ;
      RECT  23550.0 435000.0 24750.0 433800.0 ;
      RECT  23550.0 435000.0 24750.0 433800.0 ;
      RECT  23550.0 437400.0 24750.0 436200.0 ;
      RECT  33450.0 432600.0 34650.0 431400.0 ;
      RECT  23550.0 432600.0 24750.0 431400.0 ;
      RECT  28200.0 436800.0 29400.0 435600.0 ;
      RECT  28200.0 436800.0 29400.0 435600.0 ;
      RECT  28350.0 434250.0 29250.0 433350.0 ;
      RECT  35550.0 439200.0 36450.0 429600.0 ;
      RECT  21750.0 439200.0 22650.0 429600.0 ;
      RECT  28200.0 435600.0 29400.0 436800.0 ;
      RECT  34050.0 423000.0 36000.0 421800.0 ;
      RECT  22200.0 423000.0 24150.0 421800.0 ;
      RECT  23550.0 427800.0 21750.0 426600.0 ;
      RECT  32850.0 427800.0 36450.0 426600.0 ;
      RECT  23550.0 425100.0 32850.0 424200.0 ;
      RECT  32850.0 427800.0 34050.0 426600.0 ;
      RECT  32850.0 425400.0 34050.0 424200.0 ;
      RECT  32850.0 425400.0 34050.0 424200.0 ;
      RECT  32850.0 427800.0 34050.0 426600.0 ;
      RECT  23550.0 427800.0 24750.0 426600.0 ;
      RECT  23550.0 425400.0 24750.0 424200.0 ;
      RECT  23550.0 425400.0 24750.0 424200.0 ;
      RECT  23550.0 427800.0 24750.0 426600.0 ;
      RECT  33450.0 423000.0 34650.0 421800.0 ;
      RECT  23550.0 423000.0 24750.0 421800.0 ;
      RECT  28200.0 427200.0 29400.0 426000.0 ;
      RECT  28200.0 427200.0 29400.0 426000.0 ;
      RECT  28350.0 424650.0 29250.0 423750.0 ;
      RECT  35550.0 429600.0 36450.0 420000.0 ;
      RECT  21750.0 429600.0 22650.0 420000.0 ;
      RECT  28200.0 426000.0 29400.0 427200.0 ;
      RECT  34050.0 413400.0 36000.0 412200.0 ;
      RECT  22200.0 413400.0 24150.0 412200.0 ;
      RECT  23550.0 418200.0 21750.0 417000.0 ;
      RECT  32850.0 418200.0 36450.0 417000.0 ;
      RECT  23550.0 415500.0 32850.0 414600.0 ;
      RECT  32850.0 418200.0 34050.0 417000.0 ;
      RECT  32850.0 415800.0 34050.0 414600.0 ;
      RECT  32850.0 415800.0 34050.0 414600.0 ;
      RECT  32850.0 418200.0 34050.0 417000.0 ;
      RECT  23550.0 418200.0 24750.0 417000.0 ;
      RECT  23550.0 415800.0 24750.0 414600.0 ;
      RECT  23550.0 415800.0 24750.0 414600.0 ;
      RECT  23550.0 418200.0 24750.0 417000.0 ;
      RECT  33450.0 413400.0 34650.0 412200.0 ;
      RECT  23550.0 413400.0 24750.0 412200.0 ;
      RECT  28200.0 417600.0 29400.0 416400.0 ;
      RECT  28200.0 417600.0 29400.0 416400.0 ;
      RECT  28350.0 415050.0 29250.0 414150.0 ;
      RECT  35550.0 420000.0 36450.0 410400.0 ;
      RECT  21750.0 420000.0 22650.0 410400.0 ;
      RECT  28200.0 416400.0 29400.0 417600.0 ;
      RECT  42600.0 415200.0 43800.0 416400.0 ;
      RECT  42600.0 453600.0 43800.0 454800.0 ;
      RECT  42600.0 492000.0 43800.0 493200.0 ;
      RECT  28200.0 452400.0 29400.0 453600.0 ;
      RECT  42600.0 412800.0 43800.0 414000.0 ;
      RECT  28350.0 410400.0 29250.0 414150.0 ;
      RECT  35550.0 410400.0 36450.0 496800.0 ;
      RECT  21750.0 410400.0 22650.0 496800.0 ;
      RECT  49350.0 410400.0 50250.0 496800.0 ;
      RECT  16800.0 395400.0 6600.0 381600.0 ;
      RECT  16800.0 395400.0 6600.0 409200.0 ;
      RECT  16800.0 423000.0 6600.0 409200.0 ;
      RECT  17400.0 396900.0 6000.0 398100.0 ;
      RECT  17400.0 420300.0 6000.0 421500.0 ;
      RECT  17400.0 408600.0 6000.0 409500.0 ;
      RECT  22350.0 396900.0 21150.0 398100.0 ;
      RECT  22350.0 420300.0 21150.0 421500.0 ;
      RECT  22200.0 410400.0 21000.0 411600.0 ;
      RECT  22800.0 370800.0 21600.0 372000.0 ;
      RECT  16200.0 371400.0 17400.0 372600.0 ;
      RECT  6000.0 371400.0 7200.0 372600.0 ;
      RECT  29400.0 397200.0 28200.0 398400.0 ;
      RECT  19350.0 383700.0 20550.0 384900.0 ;
      RECT  19350.0 375600.0 20550.0 376800.0 ;
      RECT  12600.0 375600.0 13800.0 376800.0 ;
      RECT  43800.0 362400.0 42900.0 412800.0 ;
      RECT  29250.0 362400.0 28350.0 375750.0 ;
      RECT  4500.0 362400.0 3600.0 425250.0 ;
      RECT  36450.0 362400.0 35550.0 410400.0 ;
      RECT  22650.0 362400.0 21750.0 372000.0 ;
      RECT  50250.0 362400.0 49350.0 410400.0 ;
      RECT  43950.0 285750.0 42750.0 284550.0 ;
      RECT  43950.0 244800.0 42750.0 243600.0 ;
      RECT  33900.0 205950.0 32700.0 204750.0 ;
      RECT  29850.0 285750.0 28650.0 284550.0 ;
      RECT  27150.0 291150.0 25950.0 289950.0 ;
      RECT  30600.0 328500.0 29400.0 327300.0 ;
      RECT  27900.0 331500.0 26700.0 330300.0 ;
      RECT  41850.0 304650.0 40650.0 303450.0 ;
      RECT  43800.0 301950.0 42600.0 300750.0 ;
      RECT  45750.0 293850.0 44550.0 292650.0 ;
      RECT  14250.0 304650.0 13050.0 303450.0 ;
      RECT  16200.0 293850.0 15000.0 292650.0 ;
      RECT  18150.0 296550.0 16950.0 295350.0 ;
      RECT  29850.0 322800.0 28650.0 324000.0 ;
      RECT  30600.0 339900.0 29400.0 341100.0 ;
      RECT  16200.0 362400.0 15000.0 363600.0 ;
      RECT  29400.0 342600.0 28200.0 343800.0 ;
      RECT  50400.0 288450.0 49200.0 287250.0 ;
      RECT  36600.0 299250.0 35400.0 298050.0 ;
      RECT  22800.0 288450.0 21600.0 287250.0 ;
      RECT  9000.0 299250.0 7800.0 298050.0 ;
      RECT  43800.0 202500.0 42600.0 206100.0 ;
      RECT  36450.0 202500.0 35550.0 203400.0 ;
      RECT  50250.0 202500.0 49350.0 203400.0 ;
      RECT  55650.0 298050.0 54450.0 299250.0 ;
   LAYER  metal2 ;
      RECT  168750.0 340500.0 169650.0 343200.0 ;
      RECT  166050.0 360300.0 166950.0 363000.0 ;
      RECT  160650.0 320700.0 161550.0 323400.0 ;
      RECT  157950.0 337800.0 158850.0 340500.0 ;
      RECT  163350.0 301350.0 164250.0 304050.0 ;
      RECT  155250.0 282450.0 156150.0 285150.0 ;
      RECT  49800.0 298200.0 55050.0 299100.0 ;
      RECT  149850.0 285150.0 150750.0 287850.0 ;
      RECT  155250.0 0.0 156150.0 440700.0 ;
      RECT  157950.0 0.0 158850.0 440700.0 ;
      RECT  160650.0 0.0 161550.0 440700.0 ;
      RECT  163350.0 0.0 164250.0 440700.0 ;
      RECT  166050.0 0.0 166950.0 440700.0 ;
      RECT  168750.0 0.0 169650.0 440700.0 ;
      RECT  134550.0 37500.0 135450.0 199500.0 ;
      RECT  137250.0 37500.0 138150.0 199500.0 ;
      RECT  139950.0 37500.0 140850.0 199500.0 ;
      RECT  142650.0 37500.0 143550.0 199500.0 ;
      RECT  181650.0 422700.0 182550.0 423900.0 ;
      RECT  191850.0 422700.0 192750.0 423900.0 ;
      RECT  180150.0 5850.0 181050.0 6750.0 ;
      RECT  177000.0 5850.0 180600.0 6750.0 ;
      RECT  180150.0 6300.0 181050.0 8100.0 ;
      RECT  190350.0 5850.0 191250.0 6750.0 ;
      RECT  187200.0 5850.0 190800.0 6750.0 ;
      RECT  190350.0 6300.0 191250.0 8100.0 ;
      RECT  102600.0 420300.0 103500.0 422400.0 ;
      RECT  175500.0 199500.0 185700.0 213300.0 ;
      RECT  175500.0 227100.0 185700.0 213300.0 ;
      RECT  175500.0 227100.0 185700.0 240900.0 ;
      RECT  175500.0 254700.0 185700.0 240900.0 ;
      RECT  175500.0 254700.0 185700.0 268500.0 ;
      RECT  175500.0 282300.0 185700.0 268500.0 ;
      RECT  175500.0 282300.0 185700.0 296100.0 ;
      RECT  175500.0 309900.0 185700.0 296100.0 ;
      RECT  175500.0 309900.0 185700.0 323700.0 ;
      RECT  175500.0 337500.0 185700.0 323700.0 ;
      RECT  175500.0 337500.0 185700.0 351300.0 ;
      RECT  175500.0 365100.0 185700.0 351300.0 ;
      RECT  175500.0 365100.0 185700.0 378900.0 ;
      RECT  175500.0 392700.0 185700.0 378900.0 ;
      RECT  175500.0 392700.0 185700.0 406500.0 ;
      RECT  175500.0 420300.0 185700.0 406500.0 ;
      RECT  185700.0 199500.0 195900.0 213300.0 ;
      RECT  185700.0 227100.0 195900.0 213300.0 ;
      RECT  185700.0 227100.0 195900.0 240900.0 ;
      RECT  185700.0 254700.0 195900.0 240900.0 ;
      RECT  185700.0 254700.0 195900.0 268500.0 ;
      RECT  185700.0 282300.0 195900.0 268500.0 ;
      RECT  185700.0 282300.0 195900.0 296100.0 ;
      RECT  185700.0 309900.0 195900.0 296100.0 ;
      RECT  185700.0 309900.0 195900.0 323700.0 ;
      RECT  185700.0 337500.0 195900.0 323700.0 ;
      RECT  185700.0 337500.0 195900.0 351300.0 ;
      RECT  185700.0 365100.0 195900.0 351300.0 ;
      RECT  185700.0 365100.0 195900.0 378900.0 ;
      RECT  185700.0 392700.0 195900.0 378900.0 ;
      RECT  185700.0 392700.0 195900.0 406500.0 ;
      RECT  185700.0 420300.0 195900.0 406500.0 ;
      RECT  178500.0 200100.0 179700.0 423900.0 ;
      RECT  181500.0 198900.0 182700.0 422700.0 ;
      RECT  188700.0 200100.0 189900.0 423900.0 ;
      RECT  191700.0 198900.0 192900.0 422700.0 ;
      RECT  174900.0 198900.0 176100.0 422700.0 ;
      RECT  185100.0 198900.0 186300.0 422700.0 ;
      RECT  195300.0 198900.0 196500.0 422700.0 ;
      RECT  178500.0 426300.0 179700.0 427500.0 ;
      RECT  180900.0 426300.0 182550.0 427500.0 ;
      RECT  178500.0 433500.0 179700.0 434700.0 ;
      RECT  181650.0 433500.0 184500.0 434700.0 ;
      RECT  178500.0 426300.0 179700.0 427500.0 ;
      RECT  180900.0 426300.0 182100.0 427500.0 ;
      RECT  178500.0 433500.0 179700.0 434700.0 ;
      RECT  183300.0 433500.0 184500.0 434700.0 ;
      RECT  178650.0 423900.0 179550.0 440700.0 ;
      RECT  181650.0 423900.0 182550.0 440700.0 ;
      RECT  188700.0 426300.0 189900.0 427500.0 ;
      RECT  191100.0 426300.0 192750.0 427500.0 ;
      RECT  188700.0 433500.0 189900.0 434700.0 ;
      RECT  191850.0 433500.0 194700.0 434700.0 ;
      RECT  188700.0 426300.0 189900.0 427500.0 ;
      RECT  191100.0 426300.0 192300.0 427500.0 ;
      RECT  188700.0 433500.0 189900.0 434700.0 ;
      RECT  193500.0 433500.0 194700.0 434700.0 ;
      RECT  188850.0 423900.0 189750.0 440700.0 ;
      RECT  191850.0 423900.0 192750.0 440700.0 ;
      RECT  178650.0 423900.0 179550.0 440700.0 ;
      RECT  181650.0 423900.0 182550.0 440700.0 ;
      RECT  188850.0 423900.0 189750.0 440700.0 ;
      RECT  191850.0 423900.0 192750.0 440700.0 ;
      RECT  175500.0 150600.0 185700.0 199500.0 ;
      RECT  185700.0 150600.0 195900.0 199500.0 ;
      RECT  178500.0 150600.0 179700.0 163800.0 ;
      RECT  181500.0 150600.0 182700.0 163800.0 ;
      RECT  188700.0 150600.0 189900.0 163800.0 ;
      RECT  191700.0 150600.0 192900.0 163800.0 ;
      RECT  175500.0 90000.0 185700.0 150600.0 ;
      RECT  185700.0 90000.0 195900.0 150600.0 ;
      RECT  180000.0 90000.0 181200.0 93000.0 ;
      RECT  190200.0 90000.0 191400.0 93000.0 ;
      RECT  178500.0 148500.0 179700.0 150600.0 ;
      RECT  181500.0 143100.0 182700.0 150600.0 ;
      RECT  188700.0 148500.0 189900.0 150600.0 ;
      RECT  191700.0 143100.0 192900.0 150600.0 ;
      RECT  175500.0 30000.0 185700.0 90000.0 ;
      RECT  195900.0 30000.0 185700.0 90000.0 ;
      RECT  180000.0 87600.0 182700.0 88800.0 ;
      RECT  177300.0 85500.0 178500.0 90000.0 ;
      RECT  188700.0 87600.0 191400.0 88800.0 ;
      RECT  192900.0 85500.0 194100.0 90000.0 ;
      RECT  185100.0 30000.0 186300.0 90000.0 ;
      RECT  175500.0 30000.0 185700.0 8100.0 ;
      RECT  185700.0 30000.0 195900.0 8100.0 ;
      RECT  180000.0 15000.0 181200.0 8100.0 ;
      RECT  190200.0 15000.0 191400.0 8100.0 ;
      RECT  180000.0 30000.0 181200.0 28500.0 ;
      RECT  190200.0 30000.0 191400.0 28500.0 ;
      RECT  59100.0 89100.0 60000.0 420300.0 ;
      RECT  61200.0 89100.0 62100.0 420300.0 ;
      RECT  63300.0 89100.0 64200.0 420300.0 ;
      RECT  65400.0 89100.0 66300.0 420300.0 ;
      RECT  67500.0 89100.0 68400.0 420300.0 ;
      RECT  69600.0 89100.0 70500.0 420300.0 ;
      RECT  71700.0 89100.0 72600.0 420300.0 ;
      RECT  73800.0 89100.0 74700.0 420300.0 ;
      RECT  105900.0 89100.0 105000.0 142500.0 ;
      RECT  102900.0 89100.0 102000.0 142500.0 ;
      RECT  111900.0 89100.0 111000.0 142500.0 ;
      RECT  108900.0 89100.0 108000.0 142500.0 ;
      RECT  95550.0 96450.0 94650.0 97350.0 ;
      RECT  93150.0 96450.0 92250.0 97350.0 ;
      RECT  95550.0 96900.0 94650.0 99750.0 ;
      RECT  95100.0 96450.0 92700.0 97350.0 ;
      RECT  93150.0 92250.0 92250.0 96900.0 ;
      RECT  95700.0 99750.0 94500.0 100950.0 ;
      RECT  93300.0 91050.0 92100.0 92250.0 ;
      RECT  92100.0 96300.0 93300.0 97500.0 ;
      RECT  95550.0 109350.0 94650.0 108450.0 ;
      RECT  93150.0 109350.0 92250.0 108450.0 ;
      RECT  95550.0 108900.0 94650.0 106050.0 ;
      RECT  95100.0 109350.0 92700.0 108450.0 ;
      RECT  93150.0 113550.0 92250.0 108900.0 ;
      RECT  95700.0 106050.0 94500.0 104850.0 ;
      RECT  93300.0 114750.0 92100.0 113550.0 ;
      RECT  92100.0 109500.0 93300.0 108300.0 ;
      RECT  95550.0 124050.0 94650.0 124950.0 ;
      RECT  93150.0 124050.0 92250.0 124950.0 ;
      RECT  95550.0 124500.0 94650.0 127350.0 ;
      RECT  95100.0 124050.0 92700.0 124950.0 ;
      RECT  93150.0 119850.0 92250.0 124500.0 ;
      RECT  95700.0 127350.0 94500.0 128550.0 ;
      RECT  93300.0 118650.0 92100.0 119850.0 ;
      RECT  92100.0 123900.0 93300.0 125100.0 ;
      RECT  95550.0 136950.0 94650.0 136050.0 ;
      RECT  93150.0 136950.0 92250.0 136050.0 ;
      RECT  95550.0 136500.0 94650.0 133650.0 ;
      RECT  95100.0 136950.0 92700.0 136050.0 ;
      RECT  93150.0 141150.0 92250.0 136500.0 ;
      RECT  95700.0 133650.0 94500.0 132450.0 ;
      RECT  93300.0 142350.0 92100.0 141150.0 ;
      RECT  92100.0 137100.0 93300.0 135900.0 ;
      RECT  110850.0 99600.0 112050.0 100800.0 ;
      RECT  129450.0 95100.0 130650.0 96300.0 ;
      RECT  107850.0 113400.0 109050.0 114600.0 ;
      RECT  126450.0 109500.0 127650.0 110700.0 ;
      RECT  129450.0 118200.0 130650.0 119400.0 ;
      RECT  104850.0 118200.0 106050.0 119400.0 ;
      RECT  126450.0 132000.0 127650.0 133200.0 ;
      RECT  101850.0 132000.0 103050.0 133200.0 ;
      RECT  110850.0 96300.0 112050.0 97500.0 ;
      RECT  107850.0 93600.0 109050.0 94800.0 ;
      RECT  104850.0 108300.0 106050.0 109500.0 ;
      RECT  107850.0 111000.0 109050.0 112200.0 ;
      RECT  110850.0 123900.0 112050.0 125100.0 ;
      RECT  101850.0 121200.0 103050.0 122400.0 ;
      RECT  104850.0 135900.0 106050.0 137100.0 ;
      RECT  101850.0 138600.0 103050.0 139800.0 ;
      RECT  130500.0 89100.0 129600.0 142500.0 ;
      RECT  127500.0 89100.0 126600.0 142500.0 ;
      RECT  105900.0 144300.0 105000.0 197700.0 ;
      RECT  102900.0 144300.0 102000.0 197700.0 ;
      RECT  111900.0 144300.0 111000.0 197700.0 ;
      RECT  108900.0 144300.0 108000.0 197700.0 ;
      RECT  95550.0 151650.0 94650.0 152550.0 ;
      RECT  93150.0 151650.0 92250.0 152550.0 ;
      RECT  95550.0 152100.0 94650.0 154950.0 ;
      RECT  95100.0 151650.0 92700.0 152550.0 ;
      RECT  93150.0 147450.0 92250.0 152100.0 ;
      RECT  95700.0 154950.0 94500.0 156150.0 ;
      RECT  93300.0 146250.0 92100.0 147450.0 ;
      RECT  92100.0 151500.0 93300.0 152700.0 ;
      RECT  95550.0 164550.0 94650.0 163650.0 ;
      RECT  93150.0 164550.0 92250.0 163650.0 ;
      RECT  95550.0 164100.0 94650.0 161250.0 ;
      RECT  95100.0 164550.0 92700.0 163650.0 ;
      RECT  93150.0 168750.0 92250.0 164100.0 ;
      RECT  95700.0 161250.0 94500.0 160050.0 ;
      RECT  93300.0 169950.0 92100.0 168750.0 ;
      RECT  92100.0 164700.0 93300.0 163500.0 ;
      RECT  95550.0 179250.0 94650.0 180150.0 ;
      RECT  93150.0 179250.0 92250.0 180150.0 ;
      RECT  95550.0 179700.0 94650.0 182550.0 ;
      RECT  95100.0 179250.0 92700.0 180150.0 ;
      RECT  93150.0 175050.0 92250.0 179700.0 ;
      RECT  95700.0 182550.0 94500.0 183750.0 ;
      RECT  93300.0 173850.0 92100.0 175050.0 ;
      RECT  92100.0 179100.0 93300.0 180300.0 ;
      RECT  95550.0 192150.0 94650.0 191250.0 ;
      RECT  93150.0 192150.0 92250.0 191250.0 ;
      RECT  95550.0 191700.0 94650.0 188850.0 ;
      RECT  95100.0 192150.0 92700.0 191250.0 ;
      RECT  93150.0 196350.0 92250.0 191700.0 ;
      RECT  95700.0 188850.0 94500.0 187650.0 ;
      RECT  93300.0 197550.0 92100.0 196350.0 ;
      RECT  92100.0 192300.0 93300.0 191100.0 ;
      RECT  110850.0 154800.0 112050.0 156000.0 ;
      RECT  129450.0 150300.0 130650.0 151500.0 ;
      RECT  107850.0 168600.0 109050.0 169800.0 ;
      RECT  126450.0 164700.0 127650.0 165900.0 ;
      RECT  129450.0 173400.0 130650.0 174600.0 ;
      RECT  104850.0 173400.0 106050.0 174600.0 ;
      RECT  126450.0 187200.0 127650.0 188400.0 ;
      RECT  101850.0 187200.0 103050.0 188400.0 ;
      RECT  110850.0 151500.0 112050.0 152700.0 ;
      RECT  107850.0 148800.0 109050.0 150000.0 ;
      RECT  104850.0 163500.0 106050.0 164700.0 ;
      RECT  107850.0 166200.0 109050.0 167400.0 ;
      RECT  110850.0 179100.0 112050.0 180300.0 ;
      RECT  101850.0 176400.0 103050.0 177600.0 ;
      RECT  104850.0 191100.0 106050.0 192300.0 ;
      RECT  101850.0 193800.0 103050.0 195000.0 ;
      RECT  130500.0 144300.0 129600.0 197700.0 ;
      RECT  127500.0 144300.0 126600.0 197700.0 ;
      RECT  80250.0 206850.0 81150.0 207750.0 ;
      RECT  82650.0 206850.0 83550.0 207750.0 ;
      RECT  80250.0 207300.0 81150.0 210150.0 ;
      RECT  80700.0 206850.0 83100.0 207750.0 ;
      RECT  82650.0 202650.0 83550.0 207300.0 ;
      RECT  80100.0 210150.0 81300.0 211350.0 ;
      RECT  82500.0 201450.0 83700.0 202650.0 ;
      RECT  83700.0 206700.0 82500.0 207900.0 ;
      RECT  80250.0 219750.0 81150.0 218850.0 ;
      RECT  82650.0 219750.0 83550.0 218850.0 ;
      RECT  80250.0 219300.0 81150.0 216450.0 ;
      RECT  80700.0 219750.0 83100.0 218850.0 ;
      RECT  82650.0 223950.0 83550.0 219300.0 ;
      RECT  80100.0 216450.0 81300.0 215250.0 ;
      RECT  82500.0 225150.0 83700.0 223950.0 ;
      RECT  83700.0 219900.0 82500.0 218700.0 ;
      RECT  80250.0 234450.0 81150.0 235350.0 ;
      RECT  82650.0 234450.0 83550.0 235350.0 ;
      RECT  80250.0 234900.0 81150.0 237750.0 ;
      RECT  80700.0 234450.0 83100.0 235350.0 ;
      RECT  82650.0 230250.0 83550.0 234900.0 ;
      RECT  80100.0 237750.0 81300.0 238950.0 ;
      RECT  82500.0 229050.0 83700.0 230250.0 ;
      RECT  83700.0 234300.0 82500.0 235500.0 ;
      RECT  80250.0 247350.0 81150.0 246450.0 ;
      RECT  82650.0 247350.0 83550.0 246450.0 ;
      RECT  80250.0 246900.0 81150.0 244050.0 ;
      RECT  80700.0 247350.0 83100.0 246450.0 ;
      RECT  82650.0 251550.0 83550.0 246900.0 ;
      RECT  80100.0 244050.0 81300.0 242850.0 ;
      RECT  82500.0 252750.0 83700.0 251550.0 ;
      RECT  83700.0 247500.0 82500.0 246300.0 ;
      RECT  80250.0 262050.0 81150.0 262950.0 ;
      RECT  82650.0 262050.0 83550.0 262950.0 ;
      RECT  80250.0 262500.0 81150.0 265350.0 ;
      RECT  80700.0 262050.0 83100.0 262950.0 ;
      RECT  82650.0 257850.0 83550.0 262500.0 ;
      RECT  80100.0 265350.0 81300.0 266550.0 ;
      RECT  82500.0 256650.0 83700.0 257850.0 ;
      RECT  83700.0 261900.0 82500.0 263100.0 ;
      RECT  80250.0 274950.0 81150.0 274050.0 ;
      RECT  82650.0 274950.0 83550.0 274050.0 ;
      RECT  80250.0 274500.0 81150.0 271650.0 ;
      RECT  80700.0 274950.0 83100.0 274050.0 ;
      RECT  82650.0 279150.0 83550.0 274500.0 ;
      RECT  80100.0 271650.0 81300.0 270450.0 ;
      RECT  82500.0 280350.0 83700.0 279150.0 ;
      RECT  83700.0 275100.0 82500.0 273900.0 ;
      RECT  80250.0 289650.0 81150.0 290550.0 ;
      RECT  82650.0 289650.0 83550.0 290550.0 ;
      RECT  80250.0 290100.0 81150.0 292950.0 ;
      RECT  80700.0 289650.0 83100.0 290550.0 ;
      RECT  82650.0 285450.0 83550.0 290100.0 ;
      RECT  80100.0 292950.0 81300.0 294150.0 ;
      RECT  82500.0 284250.0 83700.0 285450.0 ;
      RECT  83700.0 289500.0 82500.0 290700.0 ;
      RECT  80250.0 302550.0 81150.0 301650.0 ;
      RECT  82650.0 302550.0 83550.0 301650.0 ;
      RECT  80250.0 302100.0 81150.0 299250.0 ;
      RECT  80700.0 302550.0 83100.0 301650.0 ;
      RECT  82650.0 306750.0 83550.0 302100.0 ;
      RECT  80100.0 299250.0 81300.0 298050.0 ;
      RECT  82500.0 307950.0 83700.0 306750.0 ;
      RECT  83700.0 302700.0 82500.0 301500.0 ;
      RECT  80250.0 317250.0 81150.0 318150.0 ;
      RECT  82650.0 317250.0 83550.0 318150.0 ;
      RECT  80250.0 317700.0 81150.0 320550.0 ;
      RECT  80700.0 317250.0 83100.0 318150.0 ;
      RECT  82650.0 313050.0 83550.0 317700.0 ;
      RECT  80100.0 320550.0 81300.0 321750.0 ;
      RECT  82500.0 311850.0 83700.0 313050.0 ;
      RECT  83700.0 317100.0 82500.0 318300.0 ;
      RECT  80250.0 330150.0 81150.0 329250.0 ;
      RECT  82650.0 330150.0 83550.0 329250.0 ;
      RECT  80250.0 329700.0 81150.0 326850.0 ;
      RECT  80700.0 330150.0 83100.0 329250.0 ;
      RECT  82650.0 334350.0 83550.0 329700.0 ;
      RECT  80100.0 326850.0 81300.0 325650.0 ;
      RECT  82500.0 335550.0 83700.0 334350.0 ;
      RECT  83700.0 330300.0 82500.0 329100.0 ;
      RECT  80250.0 344850.0 81150.0 345750.0 ;
      RECT  82650.0 344850.0 83550.0 345750.0 ;
      RECT  80250.0 345300.0 81150.0 348150.0 ;
      RECT  80700.0 344850.0 83100.0 345750.0 ;
      RECT  82650.0 340650.0 83550.0 345300.0 ;
      RECT  80100.0 348150.0 81300.0 349350.0 ;
      RECT  82500.0 339450.0 83700.0 340650.0 ;
      RECT  83700.0 344700.0 82500.0 345900.0 ;
      RECT  80250.0 357750.0 81150.0 356850.0 ;
      RECT  82650.0 357750.0 83550.0 356850.0 ;
      RECT  80250.0 357300.0 81150.0 354450.0 ;
      RECT  80700.0 357750.0 83100.0 356850.0 ;
      RECT  82650.0 361950.0 83550.0 357300.0 ;
      RECT  80100.0 354450.0 81300.0 353250.0 ;
      RECT  82500.0 363150.0 83700.0 361950.0 ;
      RECT  83700.0 357900.0 82500.0 356700.0 ;
      RECT  80250.0 372450.0 81150.0 373350.0 ;
      RECT  82650.0 372450.0 83550.0 373350.0 ;
      RECT  80250.0 372900.0 81150.0 375750.0 ;
      RECT  80700.0 372450.0 83100.0 373350.0 ;
      RECT  82650.0 368250.0 83550.0 372900.0 ;
      RECT  80100.0 375750.0 81300.0 376950.0 ;
      RECT  82500.0 367050.0 83700.0 368250.0 ;
      RECT  83700.0 372300.0 82500.0 373500.0 ;
      RECT  80250.0 385350.0 81150.0 384450.0 ;
      RECT  82650.0 385350.0 83550.0 384450.0 ;
      RECT  80250.0 384900.0 81150.0 382050.0 ;
      RECT  80700.0 385350.0 83100.0 384450.0 ;
      RECT  82650.0 389550.0 83550.0 384900.0 ;
      RECT  80100.0 382050.0 81300.0 380850.0 ;
      RECT  82500.0 390750.0 83700.0 389550.0 ;
      RECT  83700.0 385500.0 82500.0 384300.0 ;
      RECT  80250.0 400050.0 81150.0 400950.0 ;
      RECT  82650.0 400050.0 83550.0 400950.0 ;
      RECT  80250.0 400500.0 81150.0 403350.0 ;
      RECT  80700.0 400050.0 83100.0 400950.0 ;
      RECT  82650.0 395850.0 83550.0 400500.0 ;
      RECT  80100.0 403350.0 81300.0 404550.0 ;
      RECT  82500.0 394650.0 83700.0 395850.0 ;
      RECT  83700.0 399900.0 82500.0 401100.0 ;
      RECT  80250.0 412950.0 81150.0 412050.0 ;
      RECT  82650.0 412950.0 83550.0 412050.0 ;
      RECT  80250.0 412500.0 81150.0 409650.0 ;
      RECT  80700.0 412950.0 83100.0 412050.0 ;
      RECT  82650.0 417150.0 83550.0 412500.0 ;
      RECT  80100.0 409650.0 81300.0 408450.0 ;
      RECT  82500.0 418350.0 83700.0 417150.0 ;
      RECT  83700.0 413100.0 82500.0 411900.0 ;
      RECT  60150.0 95100.0 58950.0 96300.0 ;
      RECT  62250.0 109500.0 61050.0 110700.0 ;
      RECT  64350.0 122700.0 63150.0 123900.0 ;
      RECT  66450.0 137100.0 65250.0 138300.0 ;
      RECT  68550.0 150300.0 67350.0 151500.0 ;
      RECT  70650.0 164700.0 69450.0 165900.0 ;
      RECT  72750.0 177900.0 71550.0 179100.0 ;
      RECT  74850.0 192300.0 73650.0 193500.0 ;
      RECT  60150.0 206700.0 58950.0 207900.0 ;
      RECT  68550.0 204000.0 67350.0 205200.0 ;
      RECT  60150.0 218700.0 58950.0 219900.0 ;
      RECT  70650.0 221400.0 69450.0 222600.0 ;
      RECT  60150.0 234300.0 58950.0 235500.0 ;
      RECT  72750.0 231600.0 71550.0 232800.0 ;
      RECT  60150.0 246300.0 58950.0 247500.0 ;
      RECT  74850.0 249000.0 73650.0 250200.0 ;
      RECT  62250.0 261900.0 61050.0 263100.0 ;
      RECT  68550.0 259200.0 67350.0 260400.0 ;
      RECT  62250.0 273900.0 61050.0 275100.0 ;
      RECT  70650.0 276600.0 69450.0 277800.0 ;
      RECT  62250.0 289500.0 61050.0 290700.0 ;
      RECT  72750.0 286800.0 71550.0 288000.0 ;
      RECT  62250.0 301500.0 61050.0 302700.0 ;
      RECT  74850.0 304200.0 73650.0 305400.0 ;
      RECT  64350.0 317100.0 63150.0 318300.0 ;
      RECT  68550.0 314400.0 67350.0 315600.0 ;
      RECT  64350.0 329100.0 63150.0 330300.0 ;
      RECT  70650.0 331800.0 69450.0 333000.0 ;
      RECT  64350.0 344700.0 63150.0 345900.0 ;
      RECT  72750.0 342000.0 71550.0 343200.0 ;
      RECT  64350.0 356700.0 63150.0 357900.0 ;
      RECT  74850.0 359400.0 73650.0 360600.0 ;
      RECT  66450.0 372300.0 65250.0 373500.0 ;
      RECT  68550.0 369600.0 67350.0 370800.0 ;
      RECT  66450.0 384300.0 65250.0 385500.0 ;
      RECT  70650.0 387000.0 69450.0 388200.0 ;
      RECT  66450.0 399900.0 65250.0 401100.0 ;
      RECT  72750.0 397200.0 71550.0 398400.0 ;
      RECT  66450.0 411900.0 65250.0 413100.0 ;
      RECT  74850.0 414600.0 73650.0 415800.0 ;
      RECT  129600.0 89100.0 130500.0 142500.0 ;
      RECT  126600.0 89100.0 127500.0 142500.0 ;
      RECT  129600.0 144300.0 130500.0 197700.0 ;
      RECT  126600.0 144300.0 127500.0 197700.0 ;
      RECT  104550.0 204150.0 105450.0 205050.0 ;
      RECT  104550.0 203700.0 105450.0 204600.0 ;
      RECT  105000.0 204150.0 121200.0 205050.0 ;
      RECT  104550.0 221550.0 105450.0 222450.0 ;
      RECT  104550.0 222000.0 105450.0 222900.0 ;
      RECT  105000.0 221550.0 121200.0 222450.0 ;
      RECT  104550.0 231750.0 105450.0 232650.0 ;
      RECT  104550.0 231300.0 105450.0 232200.0 ;
      RECT  105000.0 231750.0 121200.0 232650.0 ;
      RECT  104550.0 249150.0 105450.0 250050.0 ;
      RECT  104550.0 249600.0 105450.0 250500.0 ;
      RECT  105000.0 249150.0 121200.0 250050.0 ;
      RECT  104550.0 259350.0 105450.0 260250.0 ;
      RECT  104550.0 258900.0 105450.0 259800.0 ;
      RECT  105000.0 259350.0 121200.0 260250.0 ;
      RECT  104550.0 276750.0 105450.0 277650.0 ;
      RECT  104550.0 277200.0 105450.0 278100.0 ;
      RECT  105000.0 276750.0 121200.0 277650.0 ;
      RECT  104550.0 286950.0 105450.0 287850.0 ;
      RECT  104550.0 286500.0 105450.0 287400.0 ;
      RECT  105000.0 286950.0 121200.0 287850.0 ;
      RECT  104550.0 304350.0 105450.0 305250.0 ;
      RECT  104550.0 304800.0 105450.0 305700.0 ;
      RECT  105000.0 304350.0 121200.0 305250.0 ;
      RECT  104550.0 314550.0 105450.0 315450.0 ;
      RECT  104550.0 314100.0 105450.0 315000.0 ;
      RECT  105000.0 314550.0 121200.0 315450.0 ;
      RECT  104550.0 331950.0 105450.0 332850.0 ;
      RECT  104550.0 332400.0 105450.0 333300.0 ;
      RECT  105000.0 331950.0 121200.0 332850.0 ;
      RECT  104550.0 342150.0 105450.0 343050.0 ;
      RECT  104550.0 341700.0 105450.0 342600.0 ;
      RECT  105000.0 342150.0 121200.0 343050.0 ;
      RECT  104550.0 359550.0 105450.0 360450.0 ;
      RECT  104550.0 360000.0 105450.0 360900.0 ;
      RECT  105000.0 359550.0 121200.0 360450.0 ;
      RECT  104550.0 369750.0 105450.0 370650.0 ;
      RECT  104550.0 369300.0 105450.0 370200.0 ;
      RECT  105000.0 369750.0 121200.0 370650.0 ;
      RECT  104550.0 387150.0 105450.0 388050.0 ;
      RECT  104550.0 387600.0 105450.0 388500.0 ;
      RECT  105000.0 387150.0 121200.0 388050.0 ;
      RECT  104550.0 397350.0 105450.0 398250.0 ;
      RECT  104550.0 396900.0 105450.0 397800.0 ;
      RECT  105000.0 397350.0 121200.0 398250.0 ;
      RECT  104550.0 414750.0 105450.0 415650.0 ;
      RECT  104550.0 415200.0 105450.0 416100.0 ;
      RECT  105000.0 414750.0 121200.0 415650.0 ;
      RECT  120150.0 206850.0 121050.0 207750.0 ;
      RECT  122550.0 206850.0 123450.0 207750.0 ;
      RECT  120150.0 207300.0 121050.0 210150.0 ;
      RECT  120600.0 206850.0 123000.0 207750.0 ;
      RECT  122550.0 202650.0 123450.0 207300.0 ;
      RECT  120000.0 210150.0 121200.0 211350.0 ;
      RECT  122400.0 201450.0 123600.0 202650.0 ;
      RECT  123600.0 206700.0 122400.0 207900.0 ;
      RECT  102450.0 205500.0 103650.0 206700.0 ;
      RECT  104400.0 203100.0 105600.0 204300.0 ;
      RECT  121200.0 204000.0 120000.0 205200.0 ;
      RECT  120150.0 219750.0 121050.0 218850.0 ;
      RECT  122550.0 219750.0 123450.0 218850.0 ;
      RECT  120150.0 219300.0 121050.0 216450.0 ;
      RECT  120600.0 219750.0 123000.0 218850.0 ;
      RECT  122550.0 223950.0 123450.0 219300.0 ;
      RECT  120000.0 216450.0 121200.0 215250.0 ;
      RECT  122400.0 225150.0 123600.0 223950.0 ;
      RECT  123600.0 219900.0 122400.0 218700.0 ;
      RECT  102450.0 219900.0 103650.0 221100.0 ;
      RECT  104400.0 222300.0 105600.0 223500.0 ;
      RECT  121200.0 221400.0 120000.0 222600.0 ;
      RECT  120150.0 234450.0 121050.0 235350.0 ;
      RECT  122550.0 234450.0 123450.0 235350.0 ;
      RECT  120150.0 234900.0 121050.0 237750.0 ;
      RECT  120600.0 234450.0 123000.0 235350.0 ;
      RECT  122550.0 230250.0 123450.0 234900.0 ;
      RECT  120000.0 237750.0 121200.0 238950.0 ;
      RECT  122400.0 229050.0 123600.0 230250.0 ;
      RECT  123600.0 234300.0 122400.0 235500.0 ;
      RECT  102450.0 233100.0 103650.0 234300.0 ;
      RECT  104400.0 230700.0 105600.0 231900.0 ;
      RECT  121200.0 231600.0 120000.0 232800.0 ;
      RECT  120150.0 247350.0 121050.0 246450.0 ;
      RECT  122550.0 247350.0 123450.0 246450.0 ;
      RECT  120150.0 246900.0 121050.0 244050.0 ;
      RECT  120600.0 247350.0 123000.0 246450.0 ;
      RECT  122550.0 251550.0 123450.0 246900.0 ;
      RECT  120000.0 244050.0 121200.0 242850.0 ;
      RECT  122400.0 252750.0 123600.0 251550.0 ;
      RECT  123600.0 247500.0 122400.0 246300.0 ;
      RECT  102450.0 247500.0 103650.0 248700.0 ;
      RECT  104400.0 249900.0 105600.0 251100.0 ;
      RECT  121200.0 249000.0 120000.0 250200.0 ;
      RECT  120150.0 262050.0 121050.0 262950.0 ;
      RECT  122550.0 262050.0 123450.0 262950.0 ;
      RECT  120150.0 262500.0 121050.0 265350.0 ;
      RECT  120600.0 262050.0 123000.0 262950.0 ;
      RECT  122550.0 257850.0 123450.0 262500.0 ;
      RECT  120000.0 265350.0 121200.0 266550.0 ;
      RECT  122400.0 256650.0 123600.0 257850.0 ;
      RECT  123600.0 261900.0 122400.0 263100.0 ;
      RECT  102450.0 260700.0 103650.0 261900.0 ;
      RECT  104400.0 258300.0 105600.0 259500.0 ;
      RECT  121200.0 259200.0 120000.0 260400.0 ;
      RECT  120150.0 274950.0 121050.0 274050.0 ;
      RECT  122550.0 274950.0 123450.0 274050.0 ;
      RECT  120150.0 274500.0 121050.0 271650.0 ;
      RECT  120600.0 274950.0 123000.0 274050.0 ;
      RECT  122550.0 279150.0 123450.0 274500.0 ;
      RECT  120000.0 271650.0 121200.0 270450.0 ;
      RECT  122400.0 280350.0 123600.0 279150.0 ;
      RECT  123600.0 275100.0 122400.0 273900.0 ;
      RECT  102450.0 275100.0 103650.0 276300.0 ;
      RECT  104400.0 277500.0 105600.0 278700.0 ;
      RECT  121200.0 276600.0 120000.0 277800.0 ;
      RECT  120150.0 289650.0 121050.0 290550.0 ;
      RECT  122550.0 289650.0 123450.0 290550.0 ;
      RECT  120150.0 290100.0 121050.0 292950.0 ;
      RECT  120600.0 289650.0 123000.0 290550.0 ;
      RECT  122550.0 285450.0 123450.0 290100.0 ;
      RECT  120000.0 292950.0 121200.0 294150.0 ;
      RECT  122400.0 284250.0 123600.0 285450.0 ;
      RECT  123600.0 289500.0 122400.0 290700.0 ;
      RECT  102450.0 288300.0 103650.0 289500.0 ;
      RECT  104400.0 285900.0 105600.0 287100.0 ;
      RECT  121200.0 286800.0 120000.0 288000.0 ;
      RECT  120150.0 302550.0 121050.0 301650.0 ;
      RECT  122550.0 302550.0 123450.0 301650.0 ;
      RECT  120150.0 302100.0 121050.0 299250.0 ;
      RECT  120600.0 302550.0 123000.0 301650.0 ;
      RECT  122550.0 306750.0 123450.0 302100.0 ;
      RECT  120000.0 299250.0 121200.0 298050.0 ;
      RECT  122400.0 307950.0 123600.0 306750.0 ;
      RECT  123600.0 302700.0 122400.0 301500.0 ;
      RECT  102450.0 302700.0 103650.0 303900.0 ;
      RECT  104400.0 305100.0 105600.0 306300.0 ;
      RECT  121200.0 304200.0 120000.0 305400.0 ;
      RECT  120150.0 317250.0 121050.0 318150.0 ;
      RECT  122550.0 317250.0 123450.0 318150.0 ;
      RECT  120150.0 317700.0 121050.0 320550.0 ;
      RECT  120600.0 317250.0 123000.0 318150.0 ;
      RECT  122550.0 313050.0 123450.0 317700.0 ;
      RECT  120000.0 320550.0 121200.0 321750.0 ;
      RECT  122400.0 311850.0 123600.0 313050.0 ;
      RECT  123600.0 317100.0 122400.0 318300.0 ;
      RECT  102450.0 315900.0 103650.0 317100.0 ;
      RECT  104400.0 313500.0 105600.0 314700.0 ;
      RECT  121200.0 314400.0 120000.0 315600.0 ;
      RECT  120150.0 330150.0 121050.0 329250.0 ;
      RECT  122550.0 330150.0 123450.0 329250.0 ;
      RECT  120150.0 329700.0 121050.0 326850.0 ;
      RECT  120600.0 330150.0 123000.0 329250.0 ;
      RECT  122550.0 334350.0 123450.0 329700.0 ;
      RECT  120000.0 326850.0 121200.0 325650.0 ;
      RECT  122400.0 335550.0 123600.0 334350.0 ;
      RECT  123600.0 330300.0 122400.0 329100.0 ;
      RECT  102450.0 330300.0 103650.0 331500.0 ;
      RECT  104400.0 332700.0 105600.0 333900.0 ;
      RECT  121200.0 331800.0 120000.0 333000.0 ;
      RECT  120150.0 344850.0 121050.0 345750.0 ;
      RECT  122550.0 344850.0 123450.0 345750.0 ;
      RECT  120150.0 345300.0 121050.0 348150.0 ;
      RECT  120600.0 344850.0 123000.0 345750.0 ;
      RECT  122550.0 340650.0 123450.0 345300.0 ;
      RECT  120000.0 348150.0 121200.0 349350.0 ;
      RECT  122400.0 339450.0 123600.0 340650.0 ;
      RECT  123600.0 344700.0 122400.0 345900.0 ;
      RECT  102450.0 343500.0 103650.0 344700.0 ;
      RECT  104400.0 341100.0 105600.0 342300.0 ;
      RECT  121200.0 342000.0 120000.0 343200.0 ;
      RECT  120150.0 357750.0 121050.0 356850.0 ;
      RECT  122550.0 357750.0 123450.0 356850.0 ;
      RECT  120150.0 357300.0 121050.0 354450.0 ;
      RECT  120600.0 357750.0 123000.0 356850.0 ;
      RECT  122550.0 361950.0 123450.0 357300.0 ;
      RECT  120000.0 354450.0 121200.0 353250.0 ;
      RECT  122400.0 363150.0 123600.0 361950.0 ;
      RECT  123600.0 357900.0 122400.0 356700.0 ;
      RECT  102450.0 357900.0 103650.0 359100.0 ;
      RECT  104400.0 360300.0 105600.0 361500.0 ;
      RECT  121200.0 359400.0 120000.0 360600.0 ;
      RECT  120150.0 372450.0 121050.0 373350.0 ;
      RECT  122550.0 372450.0 123450.0 373350.0 ;
      RECT  120150.0 372900.0 121050.0 375750.0 ;
      RECT  120600.0 372450.0 123000.0 373350.0 ;
      RECT  122550.0 368250.0 123450.0 372900.0 ;
      RECT  120000.0 375750.0 121200.0 376950.0 ;
      RECT  122400.0 367050.0 123600.0 368250.0 ;
      RECT  123600.0 372300.0 122400.0 373500.0 ;
      RECT  102450.0 371100.0 103650.0 372300.0 ;
      RECT  104400.0 368700.0 105600.0 369900.0 ;
      RECT  121200.0 369600.0 120000.0 370800.0 ;
      RECT  120150.0 385350.0 121050.0 384450.0 ;
      RECT  122550.0 385350.0 123450.0 384450.0 ;
      RECT  120150.0 384900.0 121050.0 382050.0 ;
      RECT  120600.0 385350.0 123000.0 384450.0 ;
      RECT  122550.0 389550.0 123450.0 384900.0 ;
      RECT  120000.0 382050.0 121200.0 380850.0 ;
      RECT  122400.0 390750.0 123600.0 389550.0 ;
      RECT  123600.0 385500.0 122400.0 384300.0 ;
      RECT  102450.0 385500.0 103650.0 386700.0 ;
      RECT  104400.0 387900.0 105600.0 389100.0 ;
      RECT  121200.0 387000.0 120000.0 388200.0 ;
      RECT  120150.0 400050.0 121050.0 400950.0 ;
      RECT  122550.0 400050.0 123450.0 400950.0 ;
      RECT  120150.0 400500.0 121050.0 403350.0 ;
      RECT  120600.0 400050.0 123000.0 400950.0 ;
      RECT  122550.0 395850.0 123450.0 400500.0 ;
      RECT  120000.0 403350.0 121200.0 404550.0 ;
      RECT  122400.0 394650.0 123600.0 395850.0 ;
      RECT  123600.0 399900.0 122400.0 401100.0 ;
      RECT  102450.0 398700.0 103650.0 399900.0 ;
      RECT  104400.0 396300.0 105600.0 397500.0 ;
      RECT  121200.0 397200.0 120000.0 398400.0 ;
      RECT  120150.0 412950.0 121050.0 412050.0 ;
      RECT  122550.0 412950.0 123450.0 412050.0 ;
      RECT  120150.0 412500.0 121050.0 409650.0 ;
      RECT  120600.0 412950.0 123000.0 412050.0 ;
      RECT  122550.0 417150.0 123450.0 412500.0 ;
      RECT  120000.0 409650.0 121200.0 408450.0 ;
      RECT  122400.0 418350.0 123600.0 417150.0 ;
      RECT  123600.0 413100.0 122400.0 411900.0 ;
      RECT  102450.0 413100.0 103650.0 414300.0 ;
      RECT  104400.0 415500.0 105600.0 416700.0 ;
      RECT  121200.0 414600.0 120000.0 415800.0 ;
      RECT  102600.0 199500.0 103500.0 420300.0 ;
      RECT  59100.0 83700.0 119100.0 73500.0 ;
      RECT  59100.0 63300.0 119100.0 73500.0 ;
      RECT  59100.0 63300.0 119100.0 53100.0 ;
      RECT  59100.0 42900.0 119100.0 53100.0 ;
      RECT  116700.0 79200.0 117900.0 76500.0 ;
      RECT  114600.0 81900.0 119100.0 80700.0 ;
      RECT  116700.0 70500.0 117900.0 67800.0 ;
      RECT  114600.0 66300.0 119100.0 65100.0 ;
      RECT  116700.0 58800.0 117900.0 56100.0 ;
      RECT  114600.0 61500.0 119100.0 60300.0 ;
      RECT  116700.0 50100.0 117900.0 47400.0 ;
      RECT  114600.0 45900.0 119100.0 44700.0 ;
      RECT  59100.0 74100.0 119100.0 72900.0 ;
      RECT  59100.0 53700.0 119100.0 52500.0 ;
      RECT  176550.0 5850.0 177750.0 7050.0 ;
      RECT  186750.0 5850.0 187950.0 7050.0 ;
      RECT  180300.0 300.0 181500.0 1500.0 ;
      RECT  190500.0 300.0 191700.0 1500.0 ;
      RECT  148050.0 200100.0 149250.0 198900.0 ;
      RECT  148050.0 227700.0 149250.0 226500.0 ;
      RECT  148050.0 255300.0 149250.0 254100.0 ;
      RECT  148050.0 282900.0 149250.0 281700.0 ;
      RECT  148050.0 310500.0 149250.0 309300.0 ;
      RECT  148050.0 338100.0 149250.0 336900.0 ;
      RECT  148050.0 365700.0 149250.0 364500.0 ;
      RECT  148050.0 393300.0 149250.0 392100.0 ;
      RECT  148050.0 420900.0 149250.0 419700.0 ;
      RECT  130500.0 91350.0 129300.0 92550.0 ;
      RECT  135600.0 91200.0 134400.0 92400.0 ;
      RECT  127500.0 105150.0 126300.0 106350.0 ;
      RECT  138300.0 105000.0 137100.0 106200.0 ;
      RECT  130500.0 146550.0 129300.0 147750.0 ;
      RECT  141000.0 146400.0 139800.0 147600.0 ;
      RECT  127500.0 160350.0 126300.0 161550.0 ;
      RECT  143700.0 160200.0 142500.0 161400.0 ;
      RECT  132600.0 88500.0 131400.0 89700.0 ;
      RECT  132600.0 88500.0 131400.0 89700.0 ;
      RECT  147450.0 89700.0 148650.0 88500.0 ;
      RECT  132600.0 116100.0 131400.0 117300.0 ;
      RECT  132600.0 116100.0 131400.0 117300.0 ;
      RECT  147450.0 117300.0 148650.0 116100.0 ;
      RECT  132600.0 143700.0 131400.0 144900.0 ;
      RECT  132600.0 143700.0 131400.0 144900.0 ;
      RECT  147450.0 144900.0 148650.0 143700.0 ;
      RECT  132600.0 171300.0 131400.0 172500.0 ;
      RECT  132600.0 171300.0 131400.0 172500.0 ;
      RECT  147450.0 172500.0 148650.0 171300.0 ;
      RECT  118500.0 77250.0 117300.0 78450.0 ;
      RECT  135600.0 77250.0 134400.0 78450.0 ;
      RECT  118500.0 68550.0 117300.0 69750.0 ;
      RECT  138300.0 68550.0 137100.0 69750.0 ;
      RECT  118500.0 56850.0 117300.0 58050.0 ;
      RECT  141000.0 56850.0 139800.0 58050.0 ;
      RECT  118500.0 48150.0 117300.0 49350.0 ;
      RECT  143700.0 48150.0 142500.0 49350.0 ;
      RECT  120300.0 72900.0 119100.0 74100.0 ;
      RECT  149250.0 73050.0 148050.0 74250.0 ;
      RECT  120300.0 52500.0 119100.0 53700.0 ;
      RECT  149250.0 52650.0 148050.0 53850.0 ;
      RECT  164400.0 32250.0 163200.0 33450.0 ;
      RECT  159000.0 27750.0 157800.0 28950.0 ;
      RECT  161700.0 25350.0 160500.0 26550.0 ;
      RECT  164400.0 428550.0 163200.0 429750.0 ;
      RECT  167100.0 97050.0 165900.0 98250.0 ;
      RECT  169800.0 195150.0 168600.0 196350.0 ;
      RECT  156300.0 85200.0 155100.0 86400.0 ;
      RECT  103650.0 421800.0 102450.0 423000.0 ;
      RECT  156300.0 421800.0 155100.0 423000.0 ;
      RECT  152550.0 23400.0 151350.0 24600.0 ;
      RECT  152550.0 193200.0 151350.0 194400.0 ;
      RECT  152550.0 95100.0 151350.0 96300.0 ;
      RECT  180000.0 0.0 180900.0 1800.0 ;
      RECT  190200.0 0.0 191100.0 1800.0 ;
      RECT  168750.0 0.0 169650.0 440700.0 ;
      RECT  166050.0 0.0 166950.0 440700.0 ;
      RECT  157950.0 0.0 158850.0 440700.0 ;
      RECT  160650.0 0.0 161550.0 440700.0 ;
      RECT  163350.0 0.0 164250.0 440700.0 ;
      RECT  155250.0 0.0 156150.0 440700.0 ;
      RECT  148050.0 0.0 152550.0 440700.0 ;
      RECT  49800.0 290100.0 1.42108547152e-11 291000.0 ;
      RECT  49800.0 292800.0 1.42108547152e-11 293700.0 ;
      RECT  49800.0 295500.0 1.42108547152e-11 296400.0 ;
      RECT  49800.0 300900.0 1.42108547152e-11 301800.0 ;
      RECT  43350.0 243750.0 36000.0 244650.0 ;
      RECT  33750.0 205350.0 32850.0 285150.0 ;
      RECT  49800.0 287400.0 47100.0 288300.0 ;
      RECT  38700.0 298200.0 36000.0 299100.0 ;
      RECT  24900.0 287400.0 22200.0 288300.0 ;
      RECT  11100.0 298200.0 8400.0 299100.0 ;
      RECT  7.1054273576e-12 202500.0 10200.0 262500.0 ;
      RECT  20400.0 202500.0 10200.0 262500.0 ;
      RECT  20400.0 202500.0 30600.0 262500.0 ;
      RECT  4500.0 260100.0 7200.0 261300.0 ;
      RECT  1800.0 258000.0 3000.0 262500.0 ;
      RECT  13200.0 260100.0 15900.0 261300.0 ;
      RECT  17400.0 258000.0 18600.0 262500.0 ;
      RECT  24900.0 260100.0 27600.0 261300.0 ;
      RECT  22200.0 258000.0 23400.0 262500.0 ;
      RECT  9600.0 202500.0 10800.0 262500.0 ;
      RECT  30000.0 202500.0 31200.0 262500.0 ;
      RECT  46650.0 318150.0 39150.0 319050.0 ;
      RECT  41700.0 313350.0 40800.0 314250.0 ;
      RECT  41700.0 318150.0 40800.0 319050.0 ;
      RECT  41250.0 313350.0 39150.0 314250.0 ;
      RECT  41700.0 313800.0 40800.0 318600.0 ;
      RECT  46650.0 318150.0 41250.0 319050.0 ;
      RECT  39150.0 313200.0 37950.0 314400.0 ;
      RECT  39150.0 318000.0 37950.0 319200.0 ;
      RECT  47850.0 318000.0 46650.0 319200.0 ;
      RECT  41850.0 318000.0 40650.0 319200.0 ;
      RECT  28800.0 315750.0 29700.0 316650.0 ;
      RECT  29250.0 315750.0 32250.0 316650.0 ;
      RECT  28800.0 316200.0 29700.0 317100.0 ;
      RECT  23700.0 315750.0 24600.0 316650.0 ;
      RECT  23700.0 314400.0 24600.0 316200.0 ;
      RECT  24150.0 315750.0 29250.0 316650.0 ;
      RECT  32250.0 315600.0 33450.0 316800.0 ;
      RECT  23550.0 314400.0 24750.0 313200.0 ;
      RECT  28650.0 317700.0 29850.0 316500.0 ;
      RECT  29550.0 330450.0 30450.0 331350.0 ;
      RECT  29550.0 332850.0 30450.0 333750.0 ;
      RECT  30000.0 330450.0 32850.0 331350.0 ;
      RECT  29550.0 330900.0 30450.0 333300.0 ;
      RECT  25350.0 332850.0 30000.0 333750.0 ;
      RECT  32850.0 330300.0 34050.0 331500.0 ;
      RECT  24150.0 332700.0 25350.0 333900.0 ;
      RECT  29400.0 333900.0 30600.0 332700.0 ;
      RECT  19050.0 327750.0 11550.0 328650.0 ;
      RECT  14100.0 322950.0 13200.0 323850.0 ;
      RECT  14100.0 327750.0 13200.0 328650.0 ;
      RECT  13650.0 322950.0 11550.0 323850.0 ;
      RECT  14100.0 323400.0 13200.0 328200.0 ;
      RECT  19050.0 327750.0 13650.0 328650.0 ;
      RECT  11550.0 322800.0 10350.0 324000.0 ;
      RECT  11550.0 327600.0 10350.0 328800.0 ;
      RECT  20250.0 327600.0 19050.0 328800.0 ;
      RECT  14250.0 327600.0 13050.0 328800.0 ;
      RECT  3000.0 263100.0 1800.0 261900.0 ;
      RECT  3000.0 301950.0 1800.0 300750.0 ;
      RECT  6450.0 261900.0 5250.0 260700.0 ;
      RECT  6450.0 291150.0 5250.0 289950.0 ;
      RECT  18600.0 263100.0 17400.0 261900.0 ;
      RECT  18600.0 293850.0 17400.0 292650.0 ;
      RECT  23400.0 263100.0 22200.0 261900.0 ;
      RECT  23400.0 296550.0 22200.0 295350.0 ;
      RECT  10800.0 263100.0 9600.0 261900.0 ;
      RECT  10800.0 288450.0 9600.0 287250.0 ;
      RECT  31200.0 263100.0 30000.0 261900.0 ;
      RECT  31200.0 288450.0 30000.0 287250.0 ;
      RECT  22650.0 372000.0 21750.0 430200.0 ;
      RECT  17250.0 372000.0 16350.0 425400.0 ;
      RECT  7050.0 372000.0 6150.0 425400.0 ;
      RECT  20400.0 376200.0 19500.0 384300.0 ;
      RECT  13650.0 376200.0 12750.0 381000.0 ;
      RECT  42750.0 415800.0 43650.0 423000.0 ;
      RECT  42750.0 423000.0 43650.0 432600.0 ;
      RECT  42750.0 432600.0 43650.0 442200.0 ;
      RECT  42750.0 442200.0 43650.0 451800.0 ;
      RECT  42750.0 454200.0 43650.0 461400.0 ;
      RECT  42750.0 461400.0 43650.0 471000.0 ;
      RECT  42750.0 471000.0 43650.0 480600.0 ;
      RECT  42750.0 480600.0 43650.0 490200.0 ;
      RECT  35550.0 492150.0 36450.0 493050.0 ;
      RECT  35550.0 483750.0 36450.0 484650.0 ;
      RECT  36000.0 492150.0 43200.0 493050.0 ;
      RECT  35550.0 484200.0 36450.0 492600.0 ;
      RECT  28800.0 483750.0 36000.0 484650.0 ;
      RECT  28350.0 474600.0 29250.0 484200.0 ;
      RECT  28350.0 465000.0 29250.0 474600.0 ;
      RECT  28350.0 455400.0 29250.0 465000.0 ;
      RECT  28350.0 445800.0 29250.0 453000.0 ;
      RECT  28350.0 436200.0 29250.0 445800.0 ;
      RECT  28350.0 426600.0 29250.0 436200.0 ;
      RECT  28350.0 417000.0 29250.0 426600.0 ;
      RECT  42600.0 422400.0 43800.0 423600.0 ;
      RECT  42600.0 432000.0 43800.0 433200.0 ;
      RECT  42600.0 441600.0 43800.0 442800.0 ;
      RECT  42600.0 451200.0 43800.0 452400.0 ;
      RECT  42600.0 460800.0 43800.0 462000.0 ;
      RECT  42600.0 470400.0 43800.0 471600.0 ;
      RECT  42600.0 480000.0 43800.0 481200.0 ;
      RECT  42600.0 489600.0 43800.0 490800.0 ;
      RECT  28200.0 483600.0 29400.0 484800.0 ;
      RECT  28200.0 474000.0 29400.0 475200.0 ;
      RECT  28200.0 464400.0 29400.0 465600.0 ;
      RECT  28200.0 454800.0 29400.0 456000.0 ;
      RECT  28200.0 445200.0 29400.0 446400.0 ;
      RECT  28200.0 435600.0 29400.0 436800.0 ;
      RECT  28200.0 426000.0 29400.0 427200.0 ;
      RECT  28200.0 416400.0 29400.0 417600.0 ;
      RECT  42600.0 415200.0 43800.0 416400.0 ;
      RECT  42600.0 453600.0 43800.0 454800.0 ;
      RECT  42600.0 492000.0 43800.0 493200.0 ;
      RECT  28200.0 452400.0 29400.0 453600.0 ;
      RECT  16800.0 395400.0 6600.0 381600.0 ;
      RECT  16800.0 395400.0 6600.0 409200.0 ;
      RECT  16800.0 423000.0 6600.0 409200.0 ;
      RECT  13800.0 396000.0 12600.0 426600.0 ;
      RECT  10800.0 394800.0 9600.0 425400.0 ;
      RECT  17400.0 394800.0 16200.0 425400.0 ;
      RECT  7200.0 394800.0 6000.0 425400.0 ;
      RECT  22350.0 396900.0 21150.0 398100.0 ;
      RECT  22350.0 420300.0 21150.0 421500.0 ;
      RECT  22200.0 410400.0 21000.0 411600.0 ;
      RECT  22800.0 370800.0 21600.0 372000.0 ;
      RECT  16200.0 371400.0 17400.0 372600.0 ;
      RECT  6000.0 371400.0 7200.0 372600.0 ;
      RECT  19350.0 383700.0 20550.0 384900.0 ;
      RECT  19350.0 375600.0 20550.0 376800.0 ;
      RECT  12600.0 375600.0 13800.0 376800.0 ;
      RECT  43950.0 285750.0 42750.0 284550.0 ;
      RECT  43950.0 244800.0 42750.0 243600.0 ;
      RECT  36600.0 244800.0 35400.0 243600.0 ;
      RECT  36600.0 304650.0 35400.0 303450.0 ;
      RECT  33900.0 205950.0 32700.0 204750.0 ;
      RECT  29850.0 285750.0 28650.0 284550.0 ;
      RECT  27150.0 291150.0 25950.0 289950.0 ;
      RECT  30600.0 328500.0 29400.0 327300.0 ;
      RECT  30600.0 328500.0 29400.0 327300.0 ;
      RECT  30600.0 304650.0 29400.0 303450.0 ;
      RECT  27900.0 331500.0 26700.0 330300.0 ;
      RECT  27900.0 331500.0 26700.0 330300.0 ;
      RECT  27900.0 301950.0 26700.0 300750.0 ;
      RECT  41850.0 304650.0 40650.0 303450.0 ;
      RECT  43800.0 301950.0 42600.0 300750.0 ;
      RECT  45750.0 293850.0 44550.0 292650.0 ;
      RECT  14250.0 304650.0 13050.0 303450.0 ;
      RECT  16200.0 293850.0 15000.0 292650.0 ;
      RECT  18150.0 296550.0 16950.0 295350.0 ;
      RECT  29850.0 322800.0 28650.0 324000.0 ;
      RECT  30600.0 339900.0 29400.0 341100.0 ;
      RECT  16200.0 362400.0 15000.0 363600.0 ;
      RECT  29400.0 342600.0 28200.0 343800.0 ;
      RECT  50400.0 288450.0 49200.0 287250.0 ;
      RECT  36600.0 299250.0 35400.0 298050.0 ;
      RECT  22800.0 288450.0 21600.0 287250.0 ;
      RECT  9000.0 299250.0 7800.0 298050.0 ;
      RECT  49800.0 342750.0 28800.0 343650.0 ;
      RECT  49800.0 362550.0 15600.0 363450.0 ;
      RECT  49800.0 322950.0 29250.0 323850.0 ;
      RECT  49800.0 340050.0 30000.0 340950.0 ;
      RECT  49800.0 303600.0 1.42108547152e-11 304500.0 ;
      RECT  49800.0 284700.0 1.42108547152e-11 285600.0 ;
      RECT  49800.0 298200.0 1.42108547152e-11 299100.0 ;
      RECT  49800.0 287400.0 1.42108547152e-11 288300.0 ;
      RECT  169800.0 342600.0 168600.0 343800.0 ;
      RECT  49500.0 342750.0 48300.0 343950.0 ;
      RECT  167100.0 362400.0 165900.0 363600.0 ;
      RECT  49500.0 362550.0 48300.0 363750.0 ;
      RECT  161700.0 322800.0 160500.0 324000.0 ;
      RECT  49500.0 322950.0 48300.0 324150.0 ;
      RECT  159000.0 339900.0 157800.0 341100.0 ;
      RECT  49500.0 340050.0 48300.0 341250.0 ;
      RECT  164400.0 303450.0 163200.0 304650.0 ;
      RECT  49500.0 303600.0 48300.0 304800.0 ;
      RECT  156300.0 284550.0 155100.0 285750.0 ;
      RECT  49500.0 284700.0 48300.0 285900.0 ;
      RECT  55650.0 298050.0 54450.0 299250.0 ;
      RECT  150900.0 287250.0 149700.0 288450.0 ;
      RECT  49500.0 287400.0 48300.0 288600.0 ;
   LAYER  metal3 ;
      RECT  49800.0 342450.0 169200.0 343950.0 ;
      RECT  49800.0 362250.0 166500.0 363750.0 ;
      RECT  49800.0 322650.0 161100.0 324150.0 ;
      RECT  49800.0 339750.0 158400.0 341250.0 ;
      RECT  49800.0 303300.0 163800.0 304800.0 ;
      RECT  49800.0 284400.0 155700.0 285900.0 ;
      RECT  49800.0 287100.0 150300.0 288600.0 ;
      RECT  176250.0 6300.0 177750.0 151500.0 ;
      RECT  186450.0 6300.0 187950.0 151500.0 ;
      RECT  180000.0 0.0 181500.0 30000.0 ;
      RECT  190200.0 0.0 191700.0 30000.0 ;
      RECT  132000.0 88350.0 148050.0 89850.0 ;
      RECT  132000.0 115950.0 148050.0 117450.0 ;
      RECT  132000.0 143550.0 148050.0 145050.0 ;
      RECT  132000.0 171150.0 148050.0 172650.0 ;
      RECT  176100.0 151500.0 177900.0 153300.0 ;
      RECT  186300.0 151500.0 188100.0 153300.0 ;
      RECT  179700.0 30900.0 181500.0 32700.0 ;
      RECT  189900.0 30900.0 191700.0 32700.0 ;
      RECT  60000.0 79500.0 61800.0 77700.0 ;
      RECT  60000.0 69300.0 61800.0 67500.0 ;
      RECT  60000.0 59100.0 61800.0 57300.0 ;
      RECT  60000.0 48900.0 61800.0 47100.0 ;
      RECT  176250.0 5550.0 178050.0 7350.0 ;
      RECT  186450.0 5550.0 188250.0 7350.0 ;
      RECT  180000.0 0.0 181800.0 1800.0 ;
      RECT  190200.0 0.0 192000.0 1800.0 ;
      RECT  132900.0 88200.0 131100.0 90000.0 ;
      RECT  147150.0 90000.0 148950.0 88200.0 ;
      RECT  132900.0 115800.0 131100.0 117600.0 ;
      RECT  147150.0 117600.0 148950.0 115800.0 ;
      RECT  132900.0 143400.0 131100.0 145200.0 ;
      RECT  147150.0 145200.0 148950.0 143400.0 ;
      RECT  132900.0 171000.0 131100.0 172800.0 ;
      RECT  147150.0 172800.0 148950.0 171000.0 ;
      RECT  52800.0 77700.0 60000.0 79200.0 ;
      RECT  52800.0 67500.0 60000.0 69000.0 ;
      RECT  52800.0 57300.0 60000.0 58800.0 ;
      RECT  52800.0 47100.0 60000.0 48600.0 ;
      RECT  3150.0 262500.0 1650.0 301350.0 ;
      RECT  6600.0 261300.0 5100.0 290550.0 ;
      RECT  18750.0 262500.0 17250.0 293250.0 ;
      RECT  23550.0 262500.0 22050.0 295950.0 ;
      RECT  10950.0 262500.0 9450.0 287850.0 ;
      RECT  31350.0 262500.0 29850.0 287850.0 ;
      RECT  36750.0 244200.0 35250.0 304050.0 ;
      RECT  30750.0 304050.0 29250.0 327900.0 ;
      RECT  28050.0 301350.0 26550.0 330900.0 ;
      RECT  4200.0 203400.0 6000.0 205200.0 ;
      RECT  14400.0 203400.0 16200.0 205200.0 ;
      RECT  24600.0 203400.0 26400.0 205200.0 ;
      RECT  3300.0 263400.0 1500.0 261600.0 ;
      RECT  3300.0 302250.0 1500.0 300450.0 ;
      RECT  6750.0 262200.0 4950.0 260400.0 ;
      RECT  6750.0 291450.0 4950.0 289650.0 ;
      RECT  18900.0 263400.0 17100.0 261600.0 ;
      RECT  18900.0 294150.0 17100.0 292350.0 ;
      RECT  23700.0 263400.0 21900.0 261600.0 ;
      RECT  23700.0 296850.0 21900.0 295050.0 ;
      RECT  11100.0 263400.0 9300.0 261600.0 ;
      RECT  11100.0 288750.0 9300.0 286950.0 ;
      RECT  31500.0 263400.0 29700.0 261600.0 ;
      RECT  31500.0 288750.0 29700.0 286950.0 ;
      RECT  36900.0 245100.0 35100.0 243300.0 ;
      RECT  36900.0 304950.0 35100.0 303150.0 ;
      RECT  30900.0 328800.0 29100.0 327000.0 ;
      RECT  30900.0 304950.0 29100.0 303150.0 ;
      RECT  28200.0 331800.0 26400.0 330000.0 ;
      RECT  28200.0 302250.0 26400.0 300450.0 ;
      RECT  16200.0 203400.0 14400.0 205200.0 ;
      RECT  26400.0 203400.0 24600.0 205200.0 ;
      RECT  6000.0 203400.0 4200.0 205200.0 ;
      RECT  170100.0 342300.0 168300.0 344100.0 ;
      RECT  49800.0 342450.0 48000.0 344250.0 ;
      RECT  167400.0 362100.0 165600.0 363900.0 ;
      RECT  49800.0 362250.0 48000.0 364050.0 ;
      RECT  162000.0 322500.0 160200.0 324300.0 ;
      RECT  49800.0 322650.0 48000.0 324450.0 ;
      RECT  159300.0 339600.0 157500.0 341400.0 ;
      RECT  49800.0 339750.0 48000.0 341550.0 ;
      RECT  164700.0 303150.0 162900.0 304950.0 ;
      RECT  49800.0 303300.0 48000.0 305100.0 ;
      RECT  156600.0 284250.0 154800.0 286050.0 ;
      RECT  49800.0 284400.0 48000.0 286200.0 ;
      RECT  151200.0 286950.0 149400.0 288750.0 ;
      RECT  49800.0 287100.0 48000.0 288900.0 ;
   END
   END    sram_2_16_1_scn3me_subm
END    LIBRARY
