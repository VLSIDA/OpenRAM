VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO sram_16_16_sky130_0.05
   CLASS BLOCK ;
   SIZE 240.74 BY 171.035 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  58.355 3.03 58.685 3.29 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  64.195 3.03 64.525 3.29 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  70.035 3.03 70.365 3.29 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  75.875 3.03 76.205 3.29 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  81.715 3.03 82.045 3.29 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  87.555 3.03 87.885 3.29 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  93.395 3.03 93.725 3.29 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  99.235 3.03 99.565 3.29 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  105.075 3.03 105.405 3.29 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  110.915 3.03 111.245 3.29 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  116.755 3.03 117.085 3.29 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  122.595 3.03 122.925 3.29 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  128.435 3.03 128.765 3.29 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  134.275 3.03 134.605 3.29 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  140.115 3.03 140.445 3.29 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  145.955 3.03 146.285 3.29 ;
      END
   END din0[15]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  34.995 142.185 35.325 142.445 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  34.995 150.685 35.325 150.945 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  34.995 156.325 35.325 156.585 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  34.995 164.825 35.325 165.085 ;
      END
   END addr0[3]
   PIN addr1[0]
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  207.535 73.645 207.865 73.905 ;
      END
   END addr1[0]
   PIN addr1[1]
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  207.535 65.145 207.865 65.405 ;
      END
   END addr1[1]
   PIN addr1[2]
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  207.535 59.505 207.865 59.765 ;
      END
   END addr1[2]
   PIN addr1[3]
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  207.535 51.005 207.865 51.265 ;
      END
   END addr1[3]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  1.305 33.625 1.635 33.885 ;
      END
   END csb0
   PIN csb1
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  239.725 168.065 240.055 168.325 ;
      END
   END csb1
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  1.305 42.125 1.635 42.385 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  16.055 34.21 16.195 34.35 ;
      END
   END clk0
   PIN clk1
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  225.585 167.6 225.725 167.74 ;
      END
   END clk1
   PIN wmask0[0]
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  46.675 3.03 47.005 3.29 ;
      END
   END wmask0[0]
   PIN wmask0[1]
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  52.515 3.03 52.845 3.29 ;
      END
   END wmask0[1]
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER m1 ;
         RECT  96.78 70.725 97.01 71.995 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER m1 ;
         RECT  101.13 70.725 101.36 71.995 ;
      END
   END dout0[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER m1 ;
         RECT  103.02 70.725 103.25 71.995 ;
      END
   END dout0[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER m1 ;
         RECT  107.37 70.725 107.6 71.995 ;
      END
   END dout0[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER m1 ;
         RECT  109.26 70.725 109.49 71.995 ;
      END
   END dout0[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER m1 ;
         RECT  113.61 70.725 113.84 71.995 ;
      END
   END dout0[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER m1 ;
         RECT  115.5 70.725 115.73 71.995 ;
      END
   END dout0[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER m1 ;
         RECT  119.85 70.725 120.08 71.995 ;
      END
   END dout0[7]
   PIN dout0[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER m1 ;
         RECT  121.74 70.725 121.97 71.995 ;
      END
   END dout0[8]
   PIN dout0[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER m1 ;
         RECT  126.09 70.725 126.32 71.995 ;
      END
   END dout0[9]
   PIN dout0[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER m1 ;
         RECT  127.98 70.725 128.21 71.995 ;
      END
   END dout0[10]
   PIN dout0[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER m1 ;
         RECT  132.33 70.725 132.56 71.995 ;
      END
   END dout0[11]
   PIN dout0[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER m1 ;
         RECT  134.22 70.725 134.45 71.995 ;
      END
   END dout0[12]
   PIN dout0[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER m1 ;
         RECT  138.57 70.725 138.8 71.995 ;
      END
   END dout0[13]
   PIN dout0[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER m1 ;
         RECT  140.46 70.725 140.69 71.995 ;
      END
   END dout0[14]
   PIN dout0[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER m1 ;
         RECT  144.81 70.725 145.04 71.995 ;
      END
   END dout0[15]
   PIN dout1[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER m1 ;
         RECT  96.78 144.095 97.01 145.365 ;
      END
   END dout1[0]
   PIN dout1[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER m1 ;
         RECT  101.13 144.095 101.36 145.365 ;
      END
   END dout1[1]
   PIN dout1[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER m1 ;
         RECT  103.02 144.095 103.25 145.365 ;
      END
   END dout1[2]
   PIN dout1[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER m1 ;
         RECT  107.37 144.095 107.6 145.365 ;
      END
   END dout1[3]
   PIN dout1[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER m1 ;
         RECT  109.26 144.095 109.49 145.365 ;
      END
   END dout1[4]
   PIN dout1[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER m1 ;
         RECT  113.61 144.095 113.84 145.365 ;
      END
   END dout1[5]
   PIN dout1[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER m1 ;
         RECT  115.5 144.095 115.73 145.365 ;
      END
   END dout1[6]
   PIN dout1[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER m1 ;
         RECT  119.85 144.095 120.08 145.365 ;
      END
   END dout1[7]
   PIN dout1[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER m1 ;
         RECT  121.74 144.095 121.97 145.365 ;
      END
   END dout1[8]
   PIN dout1[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER m1 ;
         RECT  126.09 144.095 126.32 145.365 ;
      END
   END dout1[9]
   PIN dout1[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER m1 ;
         RECT  127.98 144.095 128.21 145.365 ;
      END
   END dout1[10]
   PIN dout1[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER m1 ;
         RECT  132.33 144.095 132.56 145.365 ;
      END
   END dout1[11]
   PIN dout1[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER m1 ;
         RECT  134.22 144.095 134.45 145.365 ;
      END
   END dout1[12]
   PIN dout1[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER m1 ;
         RECT  138.57 144.095 138.8 145.365 ;
      END
   END dout1[13]
   PIN dout1[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER m1 ;
         RECT  140.46 144.095 140.69 145.365 ;
      END
   END dout1[14]
   PIN dout1[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER m1 ;
         RECT  144.81 144.095 145.04 145.365 ;
      END
   END dout1[15]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER m3 ;
         RECT  67.465 100.045 67.955 100.535 ;
         LAYER m4 ;
         RECT  46.92 0.0 47.3 171.06 ;
         LAYER m3 ;
         RECT  97.67 89.29 97.97 89.59 ;
         LAYER m3 ;
         RECT  2.615 116.05 3.105 116.54 ;
         LAYER m4 ;
         RECT  143.48 0.0 143.86 7.86 ;
         LAYER m3 ;
         RECT  147.495 89.195 147.985 89.685 ;
         LAYER m3 ;
         RECT  38.08 153.0 220.02 153.38 ;
         LAYER m3 ;
         RECT  104.16 142.97 104.65 143.46 ;
         LAYER m3 ;
         RECT  174.485 109.92 174.975 110.41 ;
         LAYER m4 ;
         RECT  6.12 0.0 6.5 171.06 ;
         LAYER m3 ;
         RECT  121.94 129.36 122.43 129.85 ;
         LAYER m3 ;
         RECT  137.17 142.97 137.66 143.46 ;
         LAYER m3 ;
         RECT  134.835 60.12 135.325 60.61 ;
         LAYER m3 ;
         RECT  92.48 101.32 149.98 101.7 ;
         LAYER m3 ;
         RECT  0.0 55.08 38.46 55.46 ;
         LAYER m3 ;
         RECT  68.0 116.28 89.46 116.66 ;
         LAYER m3 ;
         RECT  107.53 129.36 108.02 129.85 ;
         LAYER m3 ;
         RECT  177.74 113.905 178.23 114.395 ;
         LAYER m3 ;
         RECT  0.0 22.44 240.42 22.82 ;
         LAYER m4 ;
         RECT  79.56 0.0 79.94 171.06 ;
         LAYER m4 ;
         RECT  128.52 61.2 128.9 171.06 ;
         LAYER m4 ;
         RECT  49.64 0.0 50.02 171.06 ;
         LAYER m3 ;
         RECT  155.72 133.96 240.42 134.34 ;
         LAYER m3 ;
         RECT  207.4 48.28 240.42 48.66 ;
         LAYER m3 ;
         RECT  40.8 72.76 199.62 73.14 ;
         LAYER m4 ;
         RECT  131.24 61.2 131.62 171.06 ;
         LAYER m3 ;
         RECT  0.0 51.0 198.94 51.38 ;
         LAYER m3 ;
         RECT  0.0 150.28 38.46 150.66 ;
         LAYER m4 ;
         RECT  89.08 0.0 89.46 171.06 ;
         LAYER m4 ;
         RECT  76.84 0.0 77.22 171.06 ;
         LAYER m3 ;
         RECT  0.0 26.52 240.42 26.9 ;
         LAYER m3 ;
         RECT  92.48 108.12 149.98 108.5 ;
         LAYER m3 ;
         RECT  92.48 97.24 149.98 97.62 ;
         LAYER m4 ;
         RECT  161.16 0.0 161.54 171.06 ;
         LAYER m4 ;
         RECT  238.68 0.0 239.06 171.06 ;
         LAYER m4 ;
         RECT  42.84 0.0 43.22 171.06 ;
         LAYER m3 ;
         RECT  95.05 86.24 95.54 86.73 ;
         LAYER m3 ;
         RECT  112.835 64.87 113.325 65.36 ;
         LAYER m3 ;
         RECT  141.6 142.97 142.09 143.46 ;
         LAYER m3 ;
         RECT  0.0 56.44 240.42 56.82 ;
         LAYER m3 ;
         RECT  43.52 163.88 240.42 164.26 ;
         LAYER m4 ;
         RECT  19.72 0.0 20.1 171.06 ;
         LAYER m3 ;
         RECT  40.8 87.72 240.42 88.1 ;
         LAYER m4 ;
         RECT  8.84 0.0 9.22 171.06 ;
         LAYER m3 ;
         RECT  174.485 117.82 174.975 118.31 ;
         LAYER m3 ;
         RECT  42.16 140.76 240.42 141.14 ;
         LAYER m3 ;
         RECT  0.0 161.16 240.42 161.54 ;
         LAYER m4 ;
         RECT  240.04 0.0 240.42 171.06 ;
         LAYER m4 ;
         RECT  133.96 0.0 134.34 171.06 ;
         LAYER m3 ;
         RECT  92.48 93.16 149.98 93.54 ;
         LAYER m4 ;
         RECT  67.32 0.0 67.7 171.06 ;
         LAYER m3 ;
         RECT  109.775 64.87 110.265 65.36 ;
         LAYER m4 ;
         RECT  223.72 0.0 224.1 171.06 ;
         LAYER m3 ;
         RECT  0.0 49.64 240.42 50.02 ;
         LAYER m3 ;
         RECT  204.68 142.12 240.42 142.5 ;
         LAYER m3 ;
         RECT  101.225 7.165 101.715 7.655 ;
         LAYER m3 ;
         RECT  143.47 76.82 143.96 77.31 ;
         LAYER m3 ;
         RECT  106.595 64.87 107.085 65.36 ;
         LAYER m3 ;
         RECT  174.485 103.995 174.975 104.485 ;
         LAYER m3 ;
         RECT  15.64 34.68 240.42 35.06 ;
         LAYER m3 ;
         RECT  106.03 76.82 106.52 77.31 ;
         LAYER m3 ;
         RECT  67.465 117.82 67.955 118.31 ;
         LAYER m4 ;
         RECT  153.0 0.0 153.38 171.06 ;
         LAYER m3 ;
         RECT  207.4 76.84 240.42 77.22 ;
         LAYER m4 ;
         RECT  91.8 16.32 92.18 171.06 ;
         LAYER m4 ;
         RECT  31.96 0.0 32.34 171.06 ;
         LAYER m3 ;
         RECT  0.0 27.88 240.42 28.26 ;
         LAYER m3 ;
         RECT  42.84 142.12 201.66 142.5 ;
         LAYER m4 ;
         RECT  144.84 8.84 145.22 171.06 ;
         LAYER m3 ;
         RECT  0.0 78.2 240.42 78.58 ;
         LAYER m3 ;
         RECT  153.0 114.92 240.42 115.3 ;
         LAYER m3 ;
         RECT  0.0 71.4 96.26 71.78 ;
         LAYER m4 ;
         RECT  108.12 0.0 108.5 171.06 ;
         LAYER m3 ;
         RECT  68.0 98.6 89.46 98.98 ;
         LAYER m3 ;
         RECT  0.0 67.32 96.26 67.7 ;
         LAYER m3 ;
         RECT  141.6 72.63 142.09 73.12 ;
         LAYER m3 ;
         RECT  174.485 119.795 174.975 120.285 ;
         LAYER m4 ;
         RECT  78.2 0.0 78.58 171.06 ;
         LAYER m4 ;
         RECT  138.04 61.2 138.42 171.06 ;
         LAYER m3 ;
         RECT  122.88 72.63 123.37 73.12 ;
         LAYER m3 ;
         RECT  92.48 105.4 149.98 105.78 ;
         LAYER m3 ;
         RECT  67.465 96.095 67.955 96.585 ;
         LAYER m3 ;
         RECT  147.56 83.64 240.42 84.02 ;
         LAYER m3 ;
         RECT  0.0 6.12 240.42 6.5 ;
         LAYER m3 ;
         RECT  92.48 94.52 149.98 94.9 ;
         LAYER m3 ;
         RECT  229.16 170.68 239.06 171.06 ;
         LAYER m3 ;
         RECT  0.0 4.76 240.42 5.14 ;
         LAYER m4 ;
         RECT  123.08 61.2 123.46 171.06 ;
         LAYER m4 ;
         RECT  234.6 0.0 234.98 171.06 ;
         LAYER m3 ;
         RECT  135.36 142.97 135.85 143.46 ;
         LAYER m3 ;
         RECT  174.485 107.945 174.975 108.435 ;
         LAYER m3 ;
         RECT  103.635 60.12 104.125 60.61 ;
         LAYER m3 ;
         RECT  174.485 111.895 174.975 112.385 ;
         LAYER m3 ;
         RECT  0.0 104.04 60.9 104.42 ;
         LAYER m4 ;
         RECT  75.48 0.0 75.86 171.06 ;
         LAYER m4 ;
         RECT  123.08 0.0 123.46 9.22 ;
         LAYER m3 ;
         RECT  43.52 157.08 201.66 157.46 ;
         LAYER m3 ;
         RECT  9.52 135.32 96.94 135.7 ;
         LAYER m3 ;
         RECT  177.74 94.155 178.23 94.645 ;
         LAYER m3 ;
         RECT  0.0 48.28 11.94 48.66 ;
         LAYER m3 ;
         RECT  153.0 105.4 174.46 105.78 ;
         LAYER m4 ;
         RECT  15.64 0.0 16.02 171.06 ;
         LAYER m3 ;
         RECT  145.52 59.16 198.94 59.54 ;
         LAYER m3 ;
         RECT  0.0 19.72 240.42 20.1 ;
         LAYER m3 ;
         RECT  0.0 70.04 38.46 70.42 ;
         LAYER m3 ;
         RECT  0.0 136.68 240.42 137.06 ;
         LAYER m3 ;
         RECT  119.075 64.87 119.565 65.36 ;
         LAYER m3 ;
         RECT  140.66 129.36 141.15 129.85 ;
         LAYER m3 ;
         RECT  21.08 48.28 204.38 48.66 ;
         LAYER m3 ;
         RECT  125.12 52.36 240.42 52.74 ;
         LAYER m3 ;
         RECT  40.8 30.6 240.42 30.98 ;
         LAYER m3 ;
         RECT  118.45 142.97 118.94 143.46 ;
         LAYER m3 ;
         RECT  97.86 138.78 98.35 139.27 ;
         LAYER m3 ;
         RECT  0.0 155.72 240.42 156.1 ;
         LAYER m3 ;
         RECT  0.0 154.36 240.42 154.74 ;
         LAYER m4 ;
         RECT  197.88 0.0 198.26 171.06 ;
         LAYER m4 ;
         RECT  219.64 0.0 220.02 171.06 ;
         LAYER m3 ;
         RECT  234.575 88.35 235.065 88.84 ;
         LAYER m4 ;
         RECT  154.36 0.0 154.74 171.06 ;
         LAYER m3 ;
         RECT  130.93 142.97 131.42 143.46 ;
         LAYER m3 ;
         RECT  238.255 99.55 238.745 100.04 ;
         LAYER m3 ;
         RECT  177.74 100.205 178.23 100.695 ;
         LAYER m3 ;
         RECT  141.35 89.29 141.65 89.59 ;
         LAYER m3 ;
         RECT  0.0 153.0 35.74 153.38 ;
         LAYER m4 ;
         RECT  157.08 0.0 157.46 171.06 ;
         LAYER m4 ;
         RECT  99.96 61.2 100.34 171.06 ;
         LAYER m3 ;
         RECT  0.0 158.44 240.42 158.82 ;
         LAYER m3 ;
         RECT  7.48 121.72 60.9 122.1 ;
         LAYER m3 ;
         RECT  53.14 98.105 53.63 98.595 ;
         LAYER m4 ;
         RECT  56.44 0.0 56.82 171.06 ;
         LAYER m4 ;
         RECT  192.44 0.0 192.82 171.06 ;
         LAYER m3 ;
         RECT  2.615 127.25 3.105 127.74 ;
         LAYER m3 ;
         RECT  34.68 31.96 240.42 32.34 ;
         LAYER m4 ;
         RECT  116.28 61.2 116.66 171.06 ;
         LAYER m3 ;
         RECT  181.56 112.2 240.42 112.58 ;
         LAYER m3 ;
         RECT  106.495 60.12 106.985 60.61 ;
         LAYER m3 ;
         RECT  122.82 76.82 123.31 77.31 ;
         LAYER m3 ;
         RECT  89.76 70.04 240.42 70.42 ;
         LAYER m3 ;
         RECT  195.425 94.12 195.915 94.61 ;
         LAYER m3 ;
         RECT  112.27 76.82 112.76 77.31 ;
         LAYER m3 ;
         RECT  92.48 123.08 149.98 123.46 ;
         LAYER m4 ;
         RECT  200.6 0.0 200.98 171.06 ;
         LAYER m3 ;
         RECT  112.735 60.12 113.225 60.61 ;
         LAYER m3 ;
         RECT  101.29 86.24 101.78 86.73 ;
         LAYER m4 ;
         RECT  139.4 8.84 139.78 171.06 ;
         LAYER m3 ;
         RECT  107.03 89.29 107.33 89.59 ;
         LAYER m3 ;
         RECT  204.68 65.96 240.42 66.34 ;
         LAYER m3 ;
         RECT  137.695 60.12 138.185 60.61 ;
         LAYER m3 ;
         RECT  100.355 64.87 100.845 65.36 ;
         LAYER m3 ;
         RECT  0.0 131.24 240.42 131.62 ;
         LAYER m3 ;
         RECT  177.74 117.855 178.23 118.345 ;
         LAYER m3 ;
         RECT  144.47 126.5 144.77 126.8 ;
         LAYER m4 ;
         RECT  61.88 0.0 62.26 171.06 ;
         LAYER m3 ;
         RECT  210.12 75.48 240.42 75.86 ;
         LAYER m3 ;
         RECT  94.455 89.195 94.945 89.685 ;
         LAYER m3 ;
         RECT  0.0 127.16 232.94 127.54 ;
         LAYER m3 ;
         RECT  0.0 37.4 240.42 37.78 ;
         LAYER m4 ;
         RECT  222.36 0.0 222.74 171.06 ;
         LAYER m3 ;
         RECT  110.15 126.5 110.45 126.8 ;
         LAYER m3 ;
         RECT  0.0 91.8 89.46 92.18 ;
         LAYER m3 ;
         RECT  146.2 7.48 240.42 7.86 ;
         LAYER m3 ;
         RECT  64.21 100.205 64.7 100.695 ;
         LAYER m3 ;
         RECT  153.0 99.96 174.46 100.34 ;
         LAYER m3 ;
         RECT  143.41 72.63 143.9 73.12 ;
         LAYER m3 ;
         RECT  64.21 102.055 64.7 102.545 ;
         LAYER m3 ;
         RECT  56.395 109.92 56.885 110.41 ;
         LAYER m3 ;
         RECT  0.0 117.64 60.9 118.02 ;
         LAYER m3 ;
         RECT  0.0 82.28 7.86 82.66 ;
         LAYER m3 ;
         RECT  92.48 91.8 149.98 92.18 ;
         LAYER m4 ;
         RECT  204.68 0.0 205.06 171.06 ;
         LAYER m3 ;
         RECT  120.01 86.24 120.5 86.73 ;
         LAYER m4 ;
         RECT  22.44 0.0 22.82 171.06 ;
         LAYER m3 ;
         RECT  92.48 110.84 149.98 111.22 ;
         LAYER m3 ;
         RECT  153.0 116.28 174.46 116.66 ;
         LAYER m3 ;
         RECT  144.84 135.32 240.42 135.7 ;
         LAYER m4 ;
         RECT  136.68 0.0 137.06 171.06 ;
         LAYER m3 ;
         RECT  138.23 89.29 138.53 89.59 ;
         LAYER m3 ;
         RECT  153.0 119.0 230.9 119.38 ;
         LAYER m4 ;
         RECT  162.52 0.0 162.9 171.06 ;
         LAYER m3 ;
         RECT  152.32 3.4 240.42 3.78 ;
         LAYER m4 ;
         RECT  97.24 61.2 97.62 171.06 ;
         LAYER m3 ;
         RECT  181.56 117.64 240.42 118.02 ;
         LAYER m4 ;
         RECT  193.8 0.0 194.18 171.06 ;
         LAYER m3 ;
         RECT  157.295 107.8 157.785 108.29 ;
         LAYER m3 ;
         RECT  97.395 60.12 97.885 60.61 ;
         LAYER m3 ;
         RECT  238.255 77.15 238.745 77.64 ;
         LAYER m3 ;
         RECT  77.865 7.165 78.355 7.655 ;
         LAYER m3 ;
         RECT  97.24 82.28 232.94 82.66 ;
         LAYER m4 ;
         RECT  30.6 0.0 30.98 171.06 ;
         LAYER m3 ;
         RECT  64.21 108.105 64.7 108.595 ;
         LAYER m3 ;
         RECT  112.905 7.165 113.395 7.655 ;
         LAYER m3 ;
         RECT  177.74 98.105 178.23 98.595 ;
         LAYER m3 ;
         RECT  99.79 76.82 100.28 77.31 ;
         LAYER m4 ;
         RECT  221.0 0.0 221.38 171.06 ;
         LAYER m3 ;
         RECT  155.04 132.6 172.42 132.98 ;
         LAYER m3 ;
         RECT  185.555 105.97 186.045 106.46 ;
         LAYER m3 ;
         RECT  92.48 98.6 149.98 98.98 ;
         LAYER m3 ;
         RECT  188.81 98.105 189.3 98.595 ;
         LAYER m4 ;
         RECT  203.32 0.0 203.7 171.06 ;
         LAYER m3 ;
         RECT  144.035 64.87 144.525 65.36 ;
         LAYER m3 ;
         RECT  100.255 60.12 100.745 60.61 ;
         LAYER m3 ;
         RECT  0.0 10.2 67.7 10.58 ;
         LAYER m3 ;
         RECT  6.295 127.25 6.785 127.74 ;
         LAYER m4 ;
         RECT  106.76 61.2 107.14 171.06 ;
         LAYER m3 ;
         RECT  0.0 63.24 96.26 63.62 ;
         LAYER m4 ;
         RECT  37.4 0.0 37.78 171.06 ;
         LAYER m3 ;
         RECT  125.75 89.29 126.05 89.59 ;
         LAYER m3 ;
         RECT  92.48 104.04 149.98 104.42 ;
         LAYER m3 ;
         RECT  202.885 135.42 203.375 135.91 ;
         LAYER m4 ;
         RECT  34.68 0.0 35.06 171.06 ;
         LAYER m4 ;
         RECT  104.04 61.2 104.42 171.06 ;
         LAYER m4 ;
         RECT  173.4 0.0 173.78 171.06 ;
         LAYER m3 ;
         RECT  71.82 107.72 72.31 108.21 ;
         LAYER m3 ;
         RECT  36.985 146.32 37.475 146.81 ;
         LAYER m4 ;
         RECT  155.72 0.0 156.1 171.06 ;
         LAYER m3 ;
         RECT  135.11 89.29 135.41 89.59 ;
         LAYER m3 ;
         RECT  137.23 138.78 137.72 139.27 ;
         LAYER m4 ;
         RECT  174.76 0.0 175.14 171.06 ;
         LAYER m4 ;
         RECT  7.48 0.0 7.86 171.06 ;
         LAYER m3 ;
         RECT  103.22 86.24 103.71 86.73 ;
         LAYER m3 ;
         RECT  116.58 138.78 117.07 139.27 ;
         LAYER m3 ;
         RECT  92.48 124.44 149.98 124.82 ;
         LAYER m3 ;
         RECT  133.28 8.84 142.5 9.22 ;
         LAYER m3 ;
         RECT  0.0 38.76 11.26 39.14 ;
         LAYER m3 ;
         RECT  198.56 106.76 240.42 107.14 ;
         LAYER m3 ;
         RECT  131.99 126.5 132.29 126.8 ;
         LAYER m3 ;
         RECT  153.0 113.56 174.46 113.94 ;
         LAYER m3 ;
         RECT  153.0 106.76 174.46 107.14 ;
         LAYER m3 ;
         RECT  9.52 119.0 89.46 119.38 ;
         LAYER m3 ;
         RECT  146.9 129.36 147.39 129.85 ;
         LAYER m3 ;
         RECT  68.0 117.64 89.46 118.02 ;
         LAYER m3 ;
         RECT  134.42 129.36 134.91 129.85 ;
         LAYER m3 ;
         RECT  204.0 146.2 240.42 146.58 ;
         LAYER m3 ;
         RECT  144.47 89.29 144.77 89.59 ;
         LAYER m4 ;
         RECT  112.2 0.0 112.58 13.98 ;
         LAYER m3 ;
         RECT  128.495 64.87 128.985 65.36 ;
         LAYER m3 ;
         RECT  111.52 14.28 240.42 14.66 ;
         LAYER m4 ;
         RECT  195.16 0.0 195.54 171.06 ;
         LAYER m3 ;
         RECT  116.39 126.5 116.69 126.8 ;
         LAYER m3 ;
         RECT  113.77 129.36 114.26 129.85 ;
         LAYER m3 ;
         RECT  103.22 129.36 103.71 129.85 ;
         LAYER m3 ;
         RECT  60.345 7.165 60.835 7.655 ;
         LAYER m3 ;
         RECT  140.66 86.24 141.15 86.73 ;
         LAYER m3 ;
         RECT  238.255 110.75 238.745 111.24 ;
         LAYER m3 ;
         RECT  105.4 11.56 114.62 11.94 ;
         LAYER m3 ;
         RECT  0.0 80.92 85.38 81.3 ;
         LAYER m3 ;
         RECT  104.1 138.78 104.59 139.27 ;
         LAYER m4 ;
         RECT  97.24 0.0 97.62 16.7 ;
         LAYER m4 ;
         RECT  57.8 10.2 58.18 171.06 ;
         LAYER m3 ;
         RECT  138.73 86.24 139.22 86.73 ;
         LAYER m3 ;
         RECT  38.08 167.96 225.46 168.34 ;
         LAYER m3 ;
         RECT  67.465 111.895 67.955 112.385 ;
         LAYER m3 ;
         RECT  110.4 72.63 110.89 73.12 ;
         LAYER m3 ;
         RECT  131.555 64.87 132.045 65.36 ;
         LAYER m4 ;
         RECT  158.44 0.0 158.82 171.06 ;
         LAYER m3 ;
         RECT  2.615 93.65 3.105 94.14 ;
         LAYER m3 ;
         RECT  118.51 138.78 119.0 139.27 ;
         LAYER m3 ;
         RECT  153.0 109.48 174.46 109.86 ;
         LAYER m3 ;
         RECT  7.48 132.6 94.9 132.98 ;
         LAYER m4 ;
         RECT  201.96 0.0 202.34 171.06 ;
         LAYER m4 ;
         RECT  191.08 0.0 191.46 171.06 ;
         LAYER m3 ;
         RECT  128.595 60.12 129.085 60.61 ;
         LAYER m3 ;
         RECT  92.48 116.28 149.98 116.66 ;
         LAYER m3 ;
         RECT  7.48 110.84 89.46 111.22 ;
         LAYER m3 ;
         RECT  0.0 142.12 38.46 142.5 ;
         LAYER m3 ;
         RECT  153.0 91.8 230.9 92.18 ;
         LAYER m3 ;
         RECT  174.485 98.07 174.975 98.56 ;
         LAYER m3 ;
         RECT  204.0 139.4 240.42 139.78 ;
         LAYER m4 ;
         RECT  53.72 0.0 54.1 171.06 ;
         LAYER m4 ;
         RECT  48.28 0.0 48.66 171.06 ;
         LAYER m3 ;
         RECT  97.92 72.63 98.41 73.12 ;
         LAYER m3 ;
         RECT  132.49 129.36 132.98 129.85 ;
         LAYER m3 ;
         RECT  53.14 94.155 53.63 94.645 ;
         LAYER m3 ;
         RECT  134.42 86.24 134.91 86.73 ;
         LAYER m3 ;
         RECT  181.56 95.88 240.42 96.26 ;
         LAYER m4 ;
         RECT  163.88 0.0 164.26 171.06 ;
         LAYER m3 ;
         RECT  54.505 7.165 54.995 7.655 ;
         LAYER m3 ;
         RECT  122.82 138.78 123.31 139.27 ;
         LAYER m4 ;
         RECT  176.12 0.0 176.5 171.06 ;
         LAYER m3 ;
         RECT  84.655 107.8 85.145 108.29 ;
         LAYER m3 ;
         RECT  153.0 110.84 240.42 111.22 ;
         LAYER m4 ;
         RECT  150.28 10.2 150.66 171.06 ;
         LAYER m3 ;
         RECT  64.21 109.955 64.7 110.445 ;
         LAYER m3 ;
         RECT  141.35 126.5 141.65 126.8 ;
         LAYER m3 ;
         RECT  40.8 45.56 240.42 45.94 ;
         LAYER m3 ;
         RECT  153.0 123.08 240.42 123.46 ;
         LAYER m3 ;
         RECT  143.935 60.12 144.425 60.61 ;
         LAYER m3 ;
         RECT  100.79 89.29 101.09 89.59 ;
         LAYER m3 ;
         RECT  0.0 21.08 240.42 21.46 ;
         LAYER m4 ;
         RECT  86.36 14.96 86.74 171.06 ;
         LAYER m4 ;
         RECT  18.36 0.0 18.74 171.06 ;
         LAYER m4 ;
         RECT  227.8 0.0 228.18 171.06 ;
         LAYER m3 ;
         RECT  7.48 87.72 38.46 88.1 ;
         LAYER m3 ;
         RECT  64.21 119.955 64.7 120.445 ;
         LAYER m3 ;
         RECT  137.23 76.82 137.72 77.31 ;
         LAYER m3 ;
         RECT  130.99 76.82 131.48 77.31 ;
         LAYER m3 ;
         RECT  64.21 112.055 64.7 112.545 ;
         LAYER m3 ;
         RECT  97.67 126.5 97.97 126.8 ;
         LAYER m3 ;
         RECT  112.21 72.63 112.7 73.12 ;
         LAYER m3 ;
         RECT  78.88 108.12 89.46 108.5 ;
         LAYER m3 ;
         RECT  0.0 17.0 96.94 17.38 ;
         LAYER m3 ;
         RECT  67.465 109.92 67.955 110.41 ;
         LAYER m3 ;
         RECT  112.27 138.78 112.76 139.27 ;
         LAYER m3 ;
         RECT  119.51 89.29 119.81 89.59 ;
         LAYER m3 ;
         RECT  1.36 45.56 38.46 45.94 ;
         LAYER m3 ;
         RECT  145.52 61.88 204.38 62.26 ;
         LAYER m3 ;
         RECT  177.74 121.805 178.23 122.295 ;
         LAYER m3 ;
         RECT  0.0 0.68 47.3 1.06 ;
         LAYER m4 ;
         RECT  26.52 0.0 26.9 171.06 ;
         LAYER m3 ;
         RECT  64.21 104.155 64.7 104.645 ;
         LAYER m3 ;
         RECT  0.0 112.2 60.9 112.58 ;
         LAYER m3 ;
         RECT  130.99 138.78 131.48 139.27 ;
         LAYER m3 ;
         RECT  0.0 165.24 240.42 165.62 ;
         LAYER m3 ;
         RECT  68.0 99.96 89.46 100.34 ;
         LAYER m4 ;
         RECT  40.12 0.0 40.5 171.06 ;
         LAYER m3 ;
         RECT  108.12 12.92 240.42 13.3 ;
         LAYER m3 ;
         RECT  0.0 144.84 96.26 145.22 ;
         LAYER m3 ;
         RECT  152.32 8.84 240.42 9.22 ;
         LAYER m3 ;
         RECT  7.48 99.96 60.9 100.34 ;
         LAYER m4 ;
         RECT  25.16 0.0 25.54 171.06 ;
         LAYER m3 ;
         RECT  116.64 72.63 117.13 73.12 ;
         LAYER m3 ;
         RECT  0.0 94.52 43.9 94.9 ;
         LAYER m3 ;
         RECT  188.81 106.005 189.3 106.495 ;
         LAYER m3 ;
         RECT  68.0 106.76 89.46 107.14 ;
         LAYER m3 ;
         RECT  95.385 7.165 95.875 7.655 ;
         LAYER m3 ;
         RECT  234.575 99.55 235.065 100.04 ;
         LAYER m3 ;
         RECT  67.465 103.995 67.955 104.485 ;
         LAYER m3 ;
         RECT  130.93 72.63 131.42 73.12 ;
         LAYER m3 ;
         RECT  138.73 129.36 139.22 129.85 ;
         LAYER m3 ;
         RECT  67.465 94.12 67.955 94.61 ;
         LAYER m3 ;
         RECT  135.3 76.82 135.79 77.31 ;
         LAYER m3 ;
         RECT  177.74 106.005 178.23 106.495 ;
         LAYER m3 ;
         RECT  0.0 31.96 13.3 32.34 ;
         LAYER m4 ;
         RECT  21.08 0.0 21.46 171.06 ;
         LAYER m4 ;
         RECT  159.8 0.0 160.18 171.06 ;
         LAYER m4 ;
         RECT  151.64 0.0 152.02 171.06 ;
         LAYER m3 ;
         RECT  0.0 166.6 225.46 166.98 ;
         LAYER m3 ;
         RECT  92.48 114.92 149.98 115.3 ;
         LAYER m3 ;
         RECT  0.0 151.64 240.42 152.02 ;
         LAYER m3 ;
         RECT  181.56 104.04 240.42 104.42 ;
         LAYER m3 ;
         RECT  124.75 76.82 125.24 77.31 ;
         LAYER m3 ;
         RECT  0.0 106.76 43.9 107.14 ;
         LAYER m3 ;
         RECT  0.0 86.36 240.42 86.74 ;
         LAYER m4 ;
         RECT  199.24 0.0 199.62 171.06 ;
         LAYER m3 ;
         RECT  96.98 129.36 97.47 129.85 ;
         LAYER m3 ;
         RECT  56.395 94.12 56.885 94.61 ;
         LAYER m3 ;
         RECT  147.495 126.405 147.985 126.895 ;
         LAYER m4 ;
         RECT  41.48 0.0 41.86 171.06 ;
         LAYER m3 ;
         RECT  0.0 75.48 200.98 75.86 ;
         LAYER m4 ;
         RECT  52.36 0.0 52.74 171.06 ;
         LAYER m3 ;
         RECT  123.11 57.905 123.6 58.395 ;
         LAYER m3 ;
         RECT  115.7 129.36 116.19 129.85 ;
         LAYER m3 ;
         RECT  46.525 105.97 47.015 106.46 ;
         LAYER m3 ;
         RECT  153.0 117.64 174.46 118.02 ;
         LAYER m4 ;
         RECT  74.12 12.92 74.5 171.06 ;
         LAYER m3 ;
         RECT  153.0 94.52 174.46 94.9 ;
         LAYER m3 ;
         RECT  147.56 80.92 240.42 81.3 ;
         LAYER m3 ;
         RECT  109.875 60.12 110.365 60.61 ;
         LAYER m3 ;
         RECT  145.52 63.24 240.42 63.62 ;
         LAYER m3 ;
         RECT  170.13 107.72 170.62 108.21 ;
         LAYER m4 ;
         RECT  207.4 0.0 207.78 171.06 ;
         LAYER m4 ;
         RECT  117.64 0.0 118.02 171.06 ;
         LAYER m3 ;
         RECT  92.48 90.44 149.98 90.82 ;
         LAYER m3 ;
         RECT  64.21 121.805 64.7 122.295 ;
         LAYER m4 ;
         RECT  110.84 0.0 111.22 171.06 ;
         LAYER m3 ;
         RECT  141.54 138.78 142.03 139.27 ;
         LAYER m3 ;
         RECT  177.74 116.005 178.23 116.495 ;
         LAYER m3 ;
         RECT  97.92 142.97 98.41 143.46 ;
         LAYER m3 ;
         RECT  68.0 112.2 89.46 112.58 ;
         LAYER m3 ;
         RECT  0.0 36.04 240.42 36.42 ;
         LAYER m4 ;
         RECT  59.16 0.0 59.54 171.06 ;
         LAYER m4 ;
         RECT  114.92 0.0 115.3 171.06 ;
         LAYER m4 ;
         RECT  112.2 61.2 112.58 171.06 ;
         LAYER m4 ;
         RECT  68.68 11.56 69.06 171.06 ;
         LAYER m3 ;
         RECT  153.0 97.24 230.9 97.62 ;
         LAYER m3 ;
         RECT  0.0 128.52 201.66 128.9 ;
         LAYER m4 ;
         RECT  226.44 0.0 226.82 171.06 ;
         LAYER m3 ;
         RECT  0.0 65.96 199.62 66.34 ;
         LAYER m4 ;
         RECT  14.28 0.0 14.66 171.06 ;
         LAYER m3 ;
         RECT  152.32 2.04 240.42 2.42 ;
         LAYER m3 ;
         RECT  0.0 18.36 61.58 18.74 ;
         LAYER m3 ;
         RECT  6.295 93.65 6.785 94.14 ;
         LAYER m3 ;
         RECT  175.44 132.6 230.22 132.98 ;
         LAYER m3 ;
         RECT  204.68 72.76 240.42 73.14 ;
         LAYER m3 ;
         RECT  192.44 98.6 240.42 98.98 ;
         LAYER m3 ;
         RECT  64.21 113.905 64.7 114.395 ;
         LAYER m3 ;
         RECT  118.745 7.165 119.235 7.655 ;
         LAYER m3 ;
         RECT  0.0 85.0 230.9 85.38 ;
         LAYER m3 ;
         RECT  116.015 64.87 116.505 65.36 ;
         LAYER m3 ;
         RECT  177.74 119.955 178.23 120.445 ;
         LAYER m3 ;
         RECT  23.12 38.76 240.42 39.14 ;
         LAYER m3 ;
         RECT  153.0 90.44 240.42 90.82 ;
         LAYER m3 ;
         RECT  0.0 143.48 240.42 143.86 ;
         LAYER m3 ;
         RECT  116.64 142.97 117.13 143.46 ;
         LAYER m3 ;
         RECT  39.485 80.18 39.975 80.67 ;
         LAYER m3 ;
         RECT  92.48 106.76 149.98 107.14 ;
         LAYER m3 ;
         RECT  135.11 126.5 135.41 126.8 ;
         LAYER m3 ;
         RECT  177.74 96.255 178.23 96.745 ;
         LAYER m3 ;
         RECT  135.36 72.63 135.85 73.12 ;
         LAYER m3 ;
         RECT  0.0 95.88 60.9 96.26 ;
         LAYER m3 ;
         RECT  0.375 37.76 0.865 38.25 ;
         LAYER m3 ;
         RECT  89.545 7.165 90.035 7.655 ;
         LAYER m3 ;
         RECT  9.52 113.56 60.9 113.94 ;
         LAYER m4 ;
         RECT  0.68 0.0 1.06 171.06 ;
         LAYER m3 ;
         RECT  9.52 124.44 89.46 124.82 ;
         LAYER m4 ;
         RECT  147.56 0.0 147.94 171.06 ;
         LAYER m3 ;
         RECT  92.48 102.68 149.98 103.06 ;
         LAYER m3 ;
         RECT  185.555 98.07 186.045 98.56 ;
         LAYER m4 ;
         RECT  120.36 0.0 120.74 171.06 ;
         LAYER m3 ;
         RECT  116.115 60.12 116.605 60.61 ;
         LAYER m3 ;
         RECT  153.0 112.2 174.46 112.58 ;
         LAYER m3 ;
         RECT  0.0 140.76 33.02 141.14 ;
         LAYER m4 ;
         RECT  214.2 0.0 214.58 171.06 ;
         LAYER m3 ;
         RECT  174.485 96.095 174.975 96.585 ;
         LAYER m3 ;
         RECT  104.1 76.82 104.59 77.31 ;
         LAYER m4 ;
         RECT  125.8 0.0 126.18 10.58 ;
         LAYER m3 ;
         RECT  177.74 109.955 178.23 110.445 ;
         LAYER m3 ;
         RECT  0.0 33.32 240.42 33.7 ;
         LAYER m3 ;
         RECT  0.0 148.92 240.42 149.3 ;
         LAYER m3 ;
         RECT  198.56 94.52 232.94 94.9 ;
         LAYER m3 ;
         RECT  92.48 95.88 149.98 96.26 ;
         LAYER m3 ;
         RECT  0.0 11.56 73.14 11.94 ;
         LAYER m3 ;
         RECT  131.455 60.12 131.945 60.61 ;
         LAYER m4 ;
         RECT  27.88 0.0 28.26 171.06 ;
         LAYER m4 ;
         RECT  182.92 0.0 183.3 171.06 ;
         LAYER m3 ;
         RECT  0.0 15.64 90.82 16.02 ;
         LAYER m3 ;
         RECT  174.485 105.97 174.975 106.46 ;
         LAYER m4 ;
         RECT  188.36 0.0 188.74 171.06 ;
         LAYER m4 ;
         RECT  218.28 0.0 218.66 171.06 ;
         LAYER m3 ;
         RECT  106.03 138.78 106.52 139.27 ;
         LAYER m4 ;
         RECT  63.24 19.04 63.62 171.06 ;
         LAYER m4 ;
         RECT  132.6 8.84 132.98 171.06 ;
         LAYER m3 ;
         RECT  67.465 119.795 67.955 120.285 ;
         LAYER m3 ;
         RECT  0.0 25.16 240.42 25.54 ;
         LAYER m3 ;
         RECT  0.0 53.72 94.9 54.1 ;
         LAYER m3 ;
         RECT  120.01 129.36 120.5 129.85 ;
         LAYER m3 ;
         RECT  64.21 94.155 64.7 94.645 ;
         LAYER m3 ;
         RECT  0.0 72.76 38.46 73.14 ;
         LAYER m4 ;
         RECT  4.76 0.0 5.14 171.06 ;
         LAYER m4 ;
         RECT  82.28 0.0 82.66 171.06 ;
         LAYER m3 ;
         RECT  116.58 76.82 117.07 77.31 ;
         LAYER m3 ;
         RECT  147.945 7.165 148.435 7.655 ;
         LAYER m3 ;
         RECT  9.52 97.24 89.46 97.62 ;
         LAYER m4 ;
         RECT  230.52 0.0 230.9 171.06 ;
         LAYER m3 ;
         RECT  0.0 64.6 240.42 64.98 ;
         LAYER m3 ;
         RECT  0.0 29.24 240.42 29.62 ;
         LAYER m3 ;
         RECT  0.0 167.96 35.74 168.34 ;
         LAYER m4 ;
         RECT  85.0 0.0 85.38 171.06 ;
         LAYER m3 ;
         RECT  67.465 121.77 67.955 122.26 ;
         LAYER m4 ;
         RECT  212.84 0.0 213.22 171.06 ;
         LAYER m3 ;
         RECT  92.48 99.96 149.98 100.34 ;
         LAYER m3 ;
         RECT  0.0 12.92 79.26 13.3 ;
         LAYER m3 ;
         RECT  0.0 105.4 43.9 105.78 ;
         LAYER m3 ;
         RECT  114.24 15.64 240.42 16.02 ;
         LAYER m3 ;
         RECT  118.975 60.12 119.465 60.61 ;
         LAYER m4 ;
         RECT  177.48 0.0 177.86 171.06 ;
         LAYER m3 ;
         RECT  0.0 109.48 50.02 109.86 ;
         LAYER m4 ;
         RECT  102.68 0.0 103.06 171.06 ;
         LAYER m3 ;
         RECT  129.12 142.97 129.61 143.46 ;
         LAYER m3 ;
         RECT  105.97 142.97 106.46 143.46 ;
         LAYER m4 ;
         RECT  235.96 0.0 236.34 171.06 ;
         LAYER m3 ;
         RECT  109.46 129.36 109.95 129.85 ;
         LAYER m4 ;
         RECT  38.76 0.0 39.14 171.06 ;
         LAYER m4 ;
         RECT  36.04 0.0 36.42 171.06 ;
         LAYER m3 ;
         RECT  64.21 116.005 64.7 116.495 ;
         LAYER m3 ;
         RECT  131.99 89.29 132.29 89.59 ;
         LAYER m3 ;
         RECT  0.0 146.2 151.34 146.58 ;
         LAYER m3 ;
         RECT  0.0 8.84 56.14 9.22 ;
         LAYER m3 ;
         RECT  68.0 102.68 89.46 103.06 ;
         LAYER m3 ;
         RECT  144.97 129.36 145.46 129.85 ;
         LAYER m4 ;
         RECT  45.56 0.0 45.94 171.06 ;
         LAYER m3 ;
         RECT  6.295 116.05 6.785 116.54 ;
         LAYER m4 ;
         RECT  208.76 0.0 209.14 171.06 ;
         LAYER m3 ;
         RECT  119.51 126.5 119.81 126.8 ;
         LAYER m4 ;
         RECT  172.04 0.0 172.42 171.06 ;
         LAYER m4 ;
         RECT  211.48 0.0 211.86 171.06 ;
         LAYER m3 ;
         RECT  0.0 83.64 38.46 84.02 ;
         LAYER m3 ;
         RECT  48.665 7.165 49.155 7.655 ;
         LAYER m3 ;
         RECT  129.06 138.78 129.55 139.27 ;
         LAYER m4 ;
         RECT  95.88 55.08 96.26 171.06 ;
         LAYER m3 ;
         RECT  174.485 100.045 174.975 100.535 ;
         LAYER m3 ;
         RECT  68.0 113.56 89.46 113.94 ;
         LAYER m4 ;
         RECT  196.52 0.0 196.9 171.06 ;
         LAYER m3 ;
         RECT  72.025 7.165 72.515 7.655 ;
         LAYER m4 ;
         RECT  44.2 0.0 44.58 171.06 ;
         LAYER m3 ;
         RECT  96.98 86.24 97.47 86.73 ;
         LAYER m3 ;
         RECT  92.48 113.56 149.98 113.94 ;
         LAYER m3 ;
         RECT  134.735 64.87 135.225 65.36 ;
         LAYER m4 ;
         RECT  121.72 8.84 122.1 171.06 ;
         LAYER m3 ;
         RECT  128.87 126.5 129.17 126.8 ;
         LAYER m3 ;
         RECT  98.15 57.905 98.64 58.395 ;
         LAYER m4 ;
         RECT  23.8 0.0 24.18 171.06 ;
         LAYER m4 ;
         RECT  119.0 61.2 119.38 171.06 ;
         LAYER m3 ;
         RECT  129.06 76.82 129.55 77.31 ;
         LAYER m3 ;
         RECT  68.0 121.72 174.46 122.1 ;
         LAYER m3 ;
         RECT  238.255 88.35 238.745 88.84 ;
         LAYER m3 ;
         RECT  38.08 139.4 152.02 139.78 ;
         LAYER m4 ;
         RECT  105.4 0.0 105.78 171.06 ;
         LAYER m3 ;
         RECT  0.0 147.56 240.42 147.94 ;
         LAYER m4 ;
         RECT  210.12 0.0 210.5 171.06 ;
         LAYER m3 ;
         RECT  2.615 104.85 3.105 105.34 ;
         LAYER m3 ;
         RECT  107.065 7.165 107.555 7.655 ;
         LAYER m3 ;
         RECT  188.81 94.155 189.3 94.645 ;
         LAYER m3 ;
         RECT  153.0 120.36 174.46 120.74 ;
         LAYER m3 ;
         RECT  153.0 108.12 163.58 108.5 ;
         LAYER m3 ;
         RECT  122.63 89.29 122.93 89.59 ;
         LAYER m3 ;
         RECT  39.485 37.76 39.975 38.25 ;
         LAYER m3 ;
         RECT  174.485 115.845 174.975 116.335 ;
         LAYER m3 ;
         RECT  0.0 61.88 96.26 62.26 ;
         LAYER m3 ;
         RECT  181.56 116.28 232.94 116.66 ;
         LAYER m3 ;
         RECT  36.985 160.46 37.475 160.95 ;
         LAYER m4 ;
         RECT  98.6 17.68 98.98 171.06 ;
         LAYER m3 ;
         RECT  83.705 7.165 84.195 7.655 ;
         LAYER m4 ;
         RECT  12.92 0.0 13.3 171.06 ;
         LAYER m3 ;
         RECT  234.575 77.15 235.065 77.64 ;
         LAYER m3 ;
         RECT  68.0 104.04 89.46 104.42 ;
         LAYER m4 ;
         RECT  169.32 0.0 169.7 171.06 ;
         LAYER m3 ;
         RECT  125.75 126.5 126.05 126.8 ;
         LAYER m3 ;
         RECT  174.485 102.02 174.975 102.51 ;
         LAYER m3 ;
         RECT  68.0 95.88 89.46 96.26 ;
         LAYER m3 ;
         RECT  67.465 115.845 67.955 116.335 ;
         LAYER m3 ;
         RECT  99.73 142.97 100.22 143.46 ;
         LAYER m4 ;
         RECT  124.44 0.0 124.82 171.06 ;
         LAYER m3 ;
         RECT  9.52 129.88 240.42 130.26 ;
         LAYER m3 ;
         RECT  92.48 117.64 149.98 118.02 ;
         LAYER m3 ;
         RECT  113.27 126.5 113.57 126.8 ;
         LAYER m3 ;
         RECT  0.0 138.04 240.42 138.42 ;
         LAYER m3 ;
         RECT  40.8 59.16 96.26 59.54 ;
         LAYER m4 ;
         RECT  166.6 0.0 166.98 171.06 ;
         LAYER m3 ;
         RECT  153.0 104.04 174.46 104.42 ;
         LAYER m3 ;
         RECT  0.0 120.36 60.9 120.74 ;
         LAYER m3 ;
         RECT  127.16 11.56 240.42 11.94 ;
         LAYER m4 ;
         RECT  127.16 10.2 127.54 171.06 ;
         LAYER m4 ;
         RECT  148.92 0.0 149.3 171.06 ;
         LAYER m3 ;
         RECT  202.885 163.7 203.375 164.19 ;
         LAYER m3 ;
         RECT  204.68 59.16 240.42 59.54 ;
         LAYER m3 ;
         RECT  185.555 109.92 186.045 110.41 ;
         LAYER m3 ;
         RECT  2.615 138.45 3.105 138.94 ;
         LAYER m3 ;
         RECT  6.295 104.85 6.785 105.34 ;
         LAYER m3 ;
         RECT  68.0 94.52 89.46 94.9 ;
         LAYER m3 ;
         RECT  64.21 106.005 64.7 106.495 ;
         LAYER m3 ;
         RECT  130.425 7.165 130.915 7.655 ;
         LAYER m3 ;
         RECT  125.315 64.87 125.805 65.36 ;
         LAYER m3 ;
         RECT  1.36 44.2 38.46 44.58 ;
         LAYER m3 ;
         RECT  185.555 94.12 186.045 94.61 ;
         LAYER m3 ;
         RECT  53.14 109.955 53.63 110.445 ;
         LAYER m3 ;
         RECT  118.45 72.63 118.94 73.12 ;
         LAYER m4 ;
         RECT  231.88 0.0 232.26 171.06 ;
         LAYER m3 ;
         RECT  97.86 76.82 98.35 77.31 ;
         LAYER m3 ;
         RECT  153.0 98.6 174.46 98.98 ;
         LAYER m3 ;
         RECT  99.73 72.63 100.22 73.12 ;
         LAYER m3 ;
         RECT  234.575 121.95 235.065 122.44 ;
         LAYER m3 ;
         RECT  0.0 2.04 39.14 2.42 ;
         LAYER m3 ;
         RECT  122.355 60.12 122.845 60.61 ;
         LAYER m3 ;
         RECT  177.74 112.055 178.23 112.545 ;
         LAYER m3 ;
         RECT  122.63 126.5 122.93 126.8 ;
         LAYER m3 ;
         RECT  192.44 109.48 240.42 109.86 ;
         LAYER m3 ;
         RECT  147.56 55.08 240.42 55.46 ;
         LAYER m3 ;
         RECT  124.44 10.2 240.42 10.58 ;
         LAYER m3 ;
         RECT  177.74 102.055 178.23 102.545 ;
         LAYER m3 ;
         RECT  153.0 101.32 240.42 101.7 ;
         LAYER m3 ;
         RECT  135.3 138.78 135.79 139.27 ;
         LAYER m3 ;
         RECT  137.17 72.63 137.66 73.12 ;
         LAYER m3 ;
         RECT  136.265 7.165 136.755 7.655 ;
         LAYER m3 ;
         RECT  107.03 126.5 107.33 126.8 ;
         LAYER m3 ;
         RECT  0.0 46.92 240.42 47.3 ;
         LAYER m3 ;
         RECT  143.47 138.78 143.96 139.27 ;
         LAYER m3 ;
         RECT  0.0 116.28 60.9 116.66 ;
         LAYER m4 ;
         RECT  11.56 0.0 11.94 171.06 ;
         LAYER m3 ;
         RECT  181.56 121.72 240.42 122.1 ;
         LAYER m3 ;
         RECT  67.465 113.87 67.955 114.36 ;
         LAYER m3 ;
         RECT  104.16 72.63 104.65 73.12 ;
         LAYER m3 ;
         RECT  229.84 162.52 240.42 162.9 ;
         LAYER m3 ;
         RECT  0.0 79.56 230.9 79.94 ;
         LAYER m3 ;
         RECT  174.485 113.87 174.975 114.36 ;
         LAYER m3 ;
         RECT  9.52 101.32 89.46 101.7 ;
         LAYER m3 ;
         RECT  177.74 108.105 178.23 108.595 ;
         LAYER m3 ;
         RECT  125.215 60.12 125.705 60.61 ;
         LAYER m3 ;
         RECT  0.0 159.8 221.38 160.18 ;
         LAYER m3 ;
         RECT  105.97 72.63 106.46 73.12 ;
         LAYER m4 ;
         RECT  87.72 0.0 88.1 171.06 ;
         LAYER m3 ;
         RECT  67.465 107.945 67.955 108.435 ;
         LAYER m3 ;
         RECT  0.0 76.84 204.38 77.22 ;
         LAYER m3 ;
         RECT  97.92 53.72 119.38 54.1 ;
         LAYER m4 ;
         RECT  70.04 0.0 70.42 171.06 ;
         LAYER m4 ;
         RECT  229.16 0.0 229.54 171.06 ;
         LAYER m3 ;
         RECT  0.0 125.8 240.42 126.18 ;
         LAYER m4 ;
         RECT  131.24 0.0 131.62 7.86 ;
         LAYER m4 ;
         RECT  233.24 0.0 233.62 171.06 ;
         LAYER m3 ;
         RECT  107.53 86.24 108.02 86.73 ;
         LAYER m3 ;
         RECT  112.21 142.97 112.7 143.46 ;
         LAYER m4 ;
         RECT  225.08 0.0 225.46 171.06 ;
         LAYER m3 ;
         RECT  103.91 126.5 104.21 126.8 ;
         LAYER m3 ;
         RECT  0.0 3.4 50.02 3.78 ;
         LAYER m3 ;
         RECT  153.0 102.68 174.46 103.06 ;
         LAYER m3 ;
         RECT  153.0 93.16 240.42 93.54 ;
         LAYER m3 ;
         RECT  234.575 110.75 235.065 111.24 ;
         LAYER m3 ;
         RECT  92.48 109.48 149.98 109.86 ;
         LAYER m4 ;
         RECT  167.96 0.0 168.34 171.06 ;
         LAYER m3 ;
         RECT  231.88 167.96 240.42 168.34 ;
         LAYER m4 ;
         RECT  237.32 0.0 237.7 171.06 ;
         LAYER m3 ;
         RECT  14.28 40.12 240.42 40.5 ;
         LAYER m4 ;
         RECT  143.48 61.2 143.86 171.06 ;
         LAYER m3 ;
         RECT  0.0 169.32 240.42 169.7 ;
         LAYER m3 ;
         RECT  174.485 121.77 174.975 122.26 ;
         LAYER m3 ;
         RECT  113.27 89.29 113.57 89.59 ;
         LAYER m3 ;
         RECT  53.14 106.005 53.63 106.495 ;
         LAYER m3 ;
         RECT  92.48 120.36 149.98 120.74 ;
         LAYER m3 ;
         RECT  0.0 133.96 94.9 134.34 ;
         LAYER m3 ;
         RECT  141.075 60.12 141.565 60.61 ;
         LAYER m4 ;
         RECT  101.32 0.0 101.7 171.06 ;
         LAYER m3 ;
         RECT  124.69 72.63 125.18 73.12 ;
         LAYER m3 ;
         RECT  140.975 64.87 141.465 65.36 ;
         LAYER m3 ;
         RECT  99.79 138.78 100.28 139.27 ;
         LAYER m3 ;
         RECT  6.295 138.45 6.785 138.94 ;
         LAYER m4 ;
         RECT  3.4 0.0 3.78 171.06 ;
         LAYER m4 ;
         RECT  17.0 0.0 17.38 171.06 ;
         LAYER m4 ;
         RECT  165.24 0.0 165.62 171.06 ;
         LAYER m3 ;
         RECT  204.68 157.08 240.42 157.46 ;
         LAYER m3 ;
         RECT  195.425 105.97 195.915 106.46 ;
         LAYER m4 ;
         RECT  93.16 0.0 93.54 171.06 ;
         LAYER m4 ;
         RECT  170.68 0.0 171.06 171.06 ;
         LAYER m3 ;
         RECT  229.84 153.0 240.42 153.38 ;
         LAYER m3 ;
         RECT  64.21 98.105 64.7 98.595 ;
         LAYER m3 ;
         RECT  42.84 150.28 240.42 150.66 ;
         LAYER m4 ;
         RECT  216.92 0.0 217.3 171.06 ;
         LAYER m3 ;
         RECT  0.0 41.48 240.42 41.86 ;
         LAYER m3 ;
         RECT  204.68 128.52 240.42 128.9 ;
         LAYER m3 ;
         RECT  64.21 96.255 64.7 96.745 ;
         LAYER m3 ;
         RECT  101.29 129.36 101.78 129.85 ;
         LAYER m3 ;
         RECT  0.0 89.08 240.42 89.46 ;
         LAYER m3 ;
         RECT  0.0 42.84 9.9 43.22 ;
         LAYER m3 ;
         RECT  0.0 7.48 50.02 7.86 ;
         LAYER m3 ;
         RECT  188.81 109.955 189.3 110.445 ;
         LAYER m3 ;
         RECT  128.18 129.36 128.67 129.85 ;
         LAYER m4 ;
         RECT  187.0 0.0 187.38 171.06 ;
         LAYER m4 ;
         RECT  65.96 0.0 66.34 171.06 ;
         LAYER m3 ;
         RECT  92.48 112.2 149.98 112.58 ;
         LAYER m3 ;
         RECT  142.105 7.165 142.595 7.655 ;
         LAYER m4 ;
         RECT  181.56 0.0 181.94 171.06 ;
         LAYER m3 ;
         RECT  0.0 57.8 240.42 58.18 ;
         LAYER m3 ;
         RECT  1.36 30.6 38.46 30.98 ;
         LAYER m4 ;
         RECT  72.76 0.0 73.14 171.06 ;
         LAYER m4 ;
         RECT  109.48 61.2 109.86 171.06 ;
         LAYER m3 ;
         RECT  204.68 51.0 240.42 51.38 ;
         LAYER m4 ;
         RECT  55.08 0.0 55.46 171.06 ;
         LAYER m4 ;
         RECT  99.96 0.0 100.34 9.22 ;
         LAYER m3 ;
         RECT  238.255 121.95 238.745 122.44 ;
         LAYER m3 ;
         RECT  0.0 68.68 240.42 69.06 ;
         LAYER m3 ;
         RECT  228.48 159.8 240.42 160.18 ;
         LAYER m3 ;
         RECT  0.0 52.36 96.94 52.74 ;
         LAYER m3 ;
         RECT  0.0 74.12 10.58 74.5 ;
         LAYER m3 ;
         RECT  109.46 86.24 109.95 86.73 ;
         LAYER m3 ;
         RECT  0.0 60.52 240.42 60.9 ;
         LAYER m3 ;
         RECT  145.52 67.32 240.42 67.7 ;
         LAYER m4 ;
         RECT  60.52 0.0 60.9 171.06 ;
         LAYER m3 ;
         RECT  124.69 142.97 125.18 143.46 ;
         LAYER m3 ;
         RECT  110.4 142.97 110.89 143.46 ;
         LAYER m4 ;
         RECT  113.56 0.0 113.94 171.06 ;
         LAYER m3 ;
         RECT  0.0 14.28 85.38 14.66 ;
         LAYER m4 ;
         RECT  189.72 0.0 190.1 171.06 ;
         LAYER m4 ;
         RECT  180.2 0.0 180.58 171.06 ;
         LAYER m3 ;
         RECT  68.0 105.4 89.46 105.78 ;
         LAYER m3 ;
         RECT  240.495 163.7 240.985 164.19 ;
         LAYER m3 ;
         RECT  39.485 51.9 39.975 52.39 ;
         LAYER m3 ;
         RECT  0.0 59.16 38.46 59.54 ;
         LAYER m3 ;
         RECT  132.49 86.24 132.98 86.73 ;
         LAYER m3 ;
         RECT  205.385 55.14 205.875 55.63 ;
         LAYER m3 ;
         RECT  68.0 120.36 89.46 120.74 ;
         LAYER m3 ;
         RECT  115.7 86.24 116.19 86.73 ;
         LAYER m3 ;
         RECT  56.395 105.97 56.885 106.46 ;
         LAYER m3 ;
         RECT  39.485 66.04 39.975 66.53 ;
         LAYER m4 ;
         RECT  51.0 8.84 51.38 171.06 ;
         LAYER m4 ;
         RECT  71.4 0.0 71.78 171.06 ;
         LAYER m3 ;
         RECT  153.0 124.44 230.9 124.82 ;
         LAYER m4 ;
         RECT  146.2 0.0 146.58 171.06 ;
         LAYER m3 ;
         RECT  137.795 64.87 138.285 65.36 ;
         LAYER m4 ;
         RECT  129.88 0.0 130.26 171.06 ;
         LAYER m4 ;
         RECT  90.44 0.0 90.82 171.06 ;
         LAYER m4 ;
         RECT  106.76 0.0 107.14 11.94 ;
         LAYER m3 ;
         RECT  181.56 99.96 240.42 100.34 ;
         LAYER m3 ;
         RECT  94.455 126.405 94.945 126.895 ;
         LAYER m3 ;
         RECT  99.96 52.36 122.1 52.74 ;
         LAYER m3 ;
         RECT  103.91 89.29 104.21 89.59 ;
         LAYER m3 ;
         RECT  0.0 163.88 38.46 164.26 ;
         LAYER m3 ;
         RECT  143.41 142.97 143.9 143.46 ;
         LAYER m3 ;
         RECT  113.77 86.24 114.26 86.73 ;
         LAYER m3 ;
         RECT  181.56 120.36 240.42 120.74 ;
         LAYER m4 ;
         RECT  29.24 0.0 29.62 171.06 ;
         LAYER m3 ;
         RECT  174.485 94.12 174.975 94.61 ;
         LAYER m3 ;
         RECT  110.15 89.29 110.45 89.59 ;
         LAYER m3 ;
         RECT  126.25 129.36 126.74 129.85 ;
         LAYER m3 ;
         RECT  153.0 95.88 174.46 96.26 ;
         LAYER m4 ;
         RECT  140.76 61.2 141.14 171.06 ;
         LAYER m3 ;
         RECT  141.54 76.82 142.03 77.31 ;
         LAYER m3 ;
         RECT  122.88 142.97 123.37 143.46 ;
         LAYER m3 ;
         RECT  100.79 126.5 101.09 126.8 ;
         LAYER m4 ;
         RECT  178.84 0.0 179.22 171.06 ;
         LAYER m3 ;
         RECT  123.08 53.72 240.42 54.1 ;
         LAYER m4 ;
         RECT  185.64 0.0 186.02 171.06 ;
         LAYER m3 ;
         RECT  144.97 86.24 145.46 86.73 ;
         LAYER m3 ;
         RECT  116.39 89.29 116.69 89.59 ;
         LAYER m3 ;
         RECT  198.56 105.4 232.94 105.78 ;
         LAYER m3 ;
         RECT  68.0 109.48 89.46 109.86 ;
         LAYER m3 ;
         RECT  177.74 104.155 178.23 104.645 ;
         LAYER m3 ;
         RECT  121.94 86.24 122.43 86.73 ;
         LAYER m3 ;
         RECT  181.56 102.68 230.9 103.06 ;
         LAYER m3 ;
         RECT  110.34 76.82 110.83 77.31 ;
         LAYER m3 ;
         RECT  0.0 139.4 35.74 139.78 ;
         LAYER m4 ;
         RECT  94.52 0.0 94.9 171.06 ;
         LAYER m3 ;
         RECT  149.6 0.68 240.42 1.06 ;
         LAYER m4 ;
         RECT  83.64 0.0 84.02 171.06 ;
         LAYER m3 ;
         RECT  0.0 123.08 89.46 123.46 ;
         LAYER m4 ;
         RECT  125.8 61.2 126.18 171.06 ;
         LAYER m3 ;
         RECT  0.0 93.16 89.46 93.54 ;
         LAYER m3 ;
         RECT  46.525 94.12 47.015 94.61 ;
         LAYER m3 ;
         RECT  117.64 17.0 240.42 17.38 ;
         LAYER m3 ;
         RECT  103.535 64.87 104.025 65.36 ;
         LAYER m3 ;
         RECT  67.465 102.02 67.955 102.51 ;
         LAYER m3 ;
         RECT  181.56 113.56 230.9 113.94 ;
         LAYER m3 ;
         RECT  19.72 42.84 240.42 43.22 ;
         LAYER m3 ;
         RECT  9.52 108.12 60.9 108.5 ;
         LAYER m3 ;
         RECT  64.21 117.855 64.7 118.345 ;
         LAYER m3 ;
         RECT  110.34 138.78 110.83 139.27 ;
         LAYER m3 ;
         RECT  97.295 64.87 97.785 65.36 ;
         LAYER m4 ;
         RECT  215.56 0.0 215.94 171.06 ;
         LAYER m3 ;
         RECT  40.8 44.2 240.42 44.58 ;
         LAYER m4 ;
         RECT  142.12 0.0 142.5 171.06 ;
         LAYER m4 ;
         RECT  33.32 0.0 33.7 171.06 ;
         LAYER m3 ;
         RECT  67.465 105.97 67.955 106.46 ;
         LAYER m3 ;
         RECT  124.585 7.165 125.075 7.655 ;
         LAYER m3 ;
         RECT  128.87 89.29 129.17 89.59 ;
         LAYER m3 ;
         RECT  124.75 138.78 125.24 139.27 ;
         LAYER m3 ;
         RECT  66.185 7.165 66.675 7.655 ;
         LAYER m3 ;
         RECT  9.52 90.44 89.46 90.82 ;
         LAYER m3 ;
         RECT  0.0 170.68 201.66 171.06 ;
         LAYER m3 ;
         RECT  126.25 86.24 126.74 86.73 ;
         LAYER m3 ;
         RECT  205.385 69.28 205.875 69.77 ;
         LAYER m3 ;
         RECT  7.48 98.6 50.02 98.98 ;
         LAYER m3 ;
         RECT  202.885 149.56 203.375 150.05 ;
         LAYER m4 ;
         RECT  80.92 13.6 81.3 171.06 ;
         LAYER m3 ;
         RECT  0.0 23.8 240.42 24.18 ;
         LAYER m3 ;
         RECT  207.4 61.88 240.42 62.26 ;
         LAYER m4 ;
         RECT  116.28 0.0 116.66 15.34 ;
         LAYER m3 ;
         RECT  17.68 74.12 240.42 74.5 ;
         LAYER m3 ;
         RECT  128.18 86.24 128.67 86.73 ;
         LAYER m4 ;
         RECT  184.28 0.0 184.66 171.06 ;
         LAYER m3 ;
         RECT  67.465 98.07 67.955 98.56 ;
         LAYER m3 ;
         RECT  145.52 144.84 240.42 145.22 ;
         LAYER m3 ;
         RECT  118.51 76.82 119.0 77.31 ;
         LAYER m3 ;
         RECT  181.56 108.12 230.9 108.5 ;
         LAYER m3 ;
         RECT  138.23 126.5 138.53 126.8 ;
         LAYER m3 ;
         RECT  129.12 72.63 129.61 73.12 ;
         LAYER m3 ;
         RECT  0.0 157.08 38.46 157.46 ;
         LAYER m4 ;
         RECT  206.04 0.0 206.42 171.06 ;
         LAYER m4 ;
         RECT  135.32 61.2 135.7 171.06 ;
         LAYER m3 ;
         RECT  145.52 71.4 240.42 71.78 ;
         LAYER m3 ;
         RECT  122.255 64.87 122.745 65.36 ;
         LAYER m3 ;
         RECT  0.0 102.68 60.9 103.06 ;
         LAYER m3 ;
         RECT  0.0 114.92 89.46 115.3 ;
         LAYER m4 ;
         RECT  2.04 0.0 2.42 171.06 ;
         LAYER m3 ;
         RECT  99.28 18.36 240.42 18.74 ;
         LAYER m4 ;
         RECT  10.2 0.0 10.58 171.06 ;
         LAYER m3 ;
         RECT  0.0 162.52 217.98 162.9 ;
         LAYER m3 ;
         RECT  92.48 119.0 149.98 119.38 ;
         LAYER m4 ;
         RECT  64.6 0.0 64.98 171.06 ;
         LAYER m3 ;
         RECT  56.395 98.07 56.885 98.56 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER m3 ;
         RECT  205.385 62.21 205.875 62.7 ;
         LAYER m3 ;
         RECT  0.0 17.68 61.58 18.06 ;
         LAYER m3 ;
         RECT  0.0 167.28 240.42 167.66 ;
         LAYER m3 ;
         RECT  179.865 112.045 180.355 112.535 ;
         LAYER m4 ;
         RECT  182.24 0.0 182.62 171.06 ;
         LAYER m3 ;
         RECT  2.615 121.65 3.105 122.14 ;
         LAYER m4 ;
         RECT  225.76 0.0 226.14 171.06 ;
         LAYER m3 ;
         RECT  7.48 138.72 96.26 139.1 ;
         LAYER m4 ;
         RECT  54.4 0.0 54.78 171.06 ;
         LAYER m3 ;
         RECT  55.035 105.97 55.525 106.46 ;
         LAYER m4 ;
         RECT  24.48 0.0 24.86 171.06 ;
         LAYER m4 ;
         RECT  212.16 0.0 212.54 171.06 ;
         LAYER m3 ;
         RECT  0.0 161.84 240.42 162.22 ;
         LAYER m3 ;
         RECT  124.585 0.095 125.075 0.585 ;
         LAYER m4 ;
         RECT  29.92 0.0 30.3 171.06 ;
         LAYER m4 ;
         RECT  160.48 0.0 160.86 171.06 ;
         LAYER m3 ;
         RECT  23.12 38.08 38.46 38.46 ;
         LAYER m3 ;
         RECT  77.035 107.8 77.525 108.29 ;
         LAYER m3 ;
         RECT  179.52 119.68 240.42 120.06 ;
         LAYER m3 ;
         RECT  6.295 121.65 6.785 122.14 ;
         LAYER m3 ;
         RECT  69.36 100.64 173.1 101.02 ;
         LAYER m3 ;
         RECT  98.15 52.305 98.64 52.795 ;
         LAYER m3 ;
         RECT  118.45 144.58 118.94 145.07 ;
         LAYER m3 ;
         RECT  118.1 134.91 118.59 135.4 ;
         LAYER m4 ;
         RECT  95.2 0.0 95.58 171.06 ;
         LAYER m3 ;
         RECT  0.375 44.84 0.865 45.33 ;
         LAYER m3 ;
         RECT  0.0 134.64 94.9 135.02 ;
         LAYER m4 ;
         RECT  76.16 0.0 76.54 171.06 ;
         LAYER m4 ;
         RECT  146.88 0.0 147.26 171.06 ;
         LAYER m3 ;
         RECT  62.085 117.855 62.575 118.345 ;
         LAYER m3 ;
         RECT  116.07 67.055 116.56 67.545 ;
         LAYER m3 ;
         RECT  197.2 106.08 240.42 106.46 ;
         LAYER m3 ;
         RECT  0.0 84.32 38.46 84.7 ;
         LAYER m3 ;
         RECT  0.0 73.44 10.58 73.82 ;
         LAYER m3 ;
         RECT  62.085 100.195 62.575 100.685 ;
         LAYER m3 ;
         RECT  0.0 25.84 240.42 26.22 ;
         LAYER m3 ;
         RECT  91.07 90.91 91.37 91.21 ;
         LAYER m3 ;
         RECT  17.68 73.44 199.62 73.82 ;
         LAYER m3 ;
         RECT  97.325 62.2 97.815 62.69 ;
         LAYER m3 ;
         RECT  238.255 127.55 238.745 128.04 ;
         LAYER m3 ;
         RECT  147.56 54.4 240.42 54.78 ;
         LAYER m4 ;
         RECT  20.4 0.0 20.78 171.06 ;
         LAYER m3 ;
         RECT  0.0 72.08 96.26 72.46 ;
         LAYER m3 ;
         RECT  149.6 126.48 240.42 126.86 ;
         LAYER m3 ;
         RECT  91.07 116.98 91.37 117.28 ;
         LAYER m3 ;
         RECT  0.0 165.92 240.42 166.3 ;
         LAYER m3 ;
         RECT  147.56 81.6 240.42 81.98 ;
         LAYER m3 ;
         RECT  62.085 108.095 62.575 108.585 ;
         LAYER m3 ;
         RECT  2.615 132.85 3.105 133.34 ;
         LAYER m3 ;
         RECT  51.015 109.955 51.505 110.445 ;
         LAYER m3 ;
         RECT  210.12 74.8 240.42 75.18 ;
         LAYER m3 ;
         RECT  97.92 144.58 98.41 145.07 ;
         LAYER m3 ;
         RECT  145.52 77.52 232.94 77.9 ;
         LAYER m3 ;
         RECT  0.0 85.68 93.54 86.06 ;
         LAYER m3 ;
         RECT  86.36 107.44 156.1 107.82 ;
         LAYER m3 ;
         RECT  0.0 31.28 13.3 31.66 ;
         LAYER m3 ;
         RECT  118.45 71.02 118.94 71.51 ;
         LAYER m3 ;
         RECT  2.615 99.25 3.105 99.74 ;
         LAYER m4 ;
         RECT  221.68 0.0 222.06 171.06 ;
         LAYER m3 ;
         RECT  124.69 144.58 125.18 145.07 ;
         LAYER m3 ;
         RECT  69.36 93.84 173.1 94.22 ;
         LAYER m3 ;
         RECT  186.915 94.12 187.405 94.61 ;
         LAYER m4 ;
         RECT  106.08 0.0 106.46 11.94 ;
         LAYER m3 ;
         RECT  9.52 102.0 62.94 102.38 ;
         LAYER m3 ;
         RECT  0.0 43.52 240.42 43.9 ;
         LAYER m3 ;
         RECT  119.045 62.2 119.535 62.69 ;
         LAYER m3 ;
         RECT  91.07 115.795 91.37 116.095 ;
         LAYER m3 ;
         RECT  91.07 96.045 91.37 96.345 ;
         LAYER m3 ;
         RECT  104.16 144.58 104.65 145.07 ;
         LAYER m3 ;
         RECT  125.26 67.055 125.75 67.545 ;
         LAYER m3 ;
         RECT  196.785 94.12 197.275 94.61 ;
         LAYER m3 ;
         RECT  62.085 106.005 62.575 106.495 ;
         LAYER m3 ;
         RECT  127.16 12.24 240.42 12.62 ;
         LAYER m4 ;
         RECT  148.24 0.0 148.62 171.06 ;
         LAYER m3 ;
         RECT  148.92 129.2 240.42 129.58 ;
         LAYER m3 ;
         RECT  172.255 107.725 172.745 108.215 ;
         LAYER m3 ;
         RECT  151.07 116.98 151.37 117.28 ;
         LAYER m3 ;
         RECT  62.085 115.995 62.575 116.485 ;
         LAYER m3 ;
         RECT  116.64 144.58 117.13 145.07 ;
         LAYER m3 ;
         RECT  9.52 136.0 201.66 136.38 ;
         LAYER m4 ;
         RECT  161.84 0.0 162.22 171.06 ;
         LAYER m3 ;
         RECT  145.52 65.28 199.62 65.66 ;
         LAYER m3 ;
         RECT  122.31 67.055 122.8 67.545 ;
         LAYER m3 ;
         RECT  0.0 108.8 62.94 109.18 ;
         LAYER m3 ;
         RECT  175.845 121.77 176.335 122.26 ;
         LAYER m3 ;
         RECT  106.565 62.2 107.055 62.69 ;
         LAYER m3 ;
         RECT  60.345 0.095 60.835 0.585 ;
         LAYER m4 ;
         RECT  36.72 0.0 37.1 171.06 ;
         LAYER m3 ;
         RECT  0.0 82.96 7.86 83.34 ;
         LAYER m3 ;
         RECT  91.07 113.03 91.37 113.33 ;
         LAYER m3 ;
         RECT  134.79 67.055 135.28 67.545 ;
         LAYER m3 ;
         RECT  147.56 82.96 240.42 83.34 ;
         LAYER m3 ;
         RECT  62.085 94.155 62.575 94.645 ;
         LAYER m3 ;
         RECT  131.5 67.055 131.99 67.545 ;
         LAYER m3 ;
         RECT  0.0 103.36 66.34 103.74 ;
         LAYER m3 ;
         RECT  0.0 24.48 240.42 24.86 ;
         LAYER m3 ;
         RECT  118.745 0.095 119.235 0.585 ;
         LAYER m3 ;
         RECT  147.945 0.095 148.435 0.585 ;
         LAYER m4 ;
         RECT  191.76 0.0 192.14 171.06 ;
         LAYER m4 ;
         RECT  150.96 10.2 151.34 171.06 ;
         LAYER m3 ;
         RECT  112.805 62.2 113.295 62.69 ;
         LAYER m3 ;
         RECT  176.12 103.36 240.42 103.74 ;
         LAYER m4 ;
         RECT  112.88 61.2 113.26 171.06 ;
         LAYER m3 ;
         RECT  38.08 146.88 240.42 147.26 ;
         LAYER m3 ;
         RECT  141.6 71.02 142.09 71.51 ;
         LAYER m4 ;
         RECT  174.08 0.0 174.46 171.06 ;
         LAYER m4 ;
         RECT  10.88 0.0 11.26 171.06 ;
         LAYER m3 ;
         RECT  164.915 107.8 165.405 108.29 ;
         LAYER m3 ;
         RECT  118.47 63.21 118.96 63.7 ;
         LAYER m3 ;
         RECT  202.885 156.63 203.375 157.12 ;
         LAYER m3 ;
         RECT  205.385 48.07 205.875 48.56 ;
         LAYER m3 ;
         RECT  69.36 111.52 173.1 111.9 ;
         LAYER m3 ;
         RECT  116.64 71.02 117.13 71.51 ;
         LAYER m3 ;
         RECT  105.62 134.91 106.11 135.4 ;
         LAYER m3 ;
         RECT  0.0 76.16 96.26 76.54 ;
         LAYER m3 ;
         RECT  99.73 144.58 100.22 145.07 ;
         LAYER m3 ;
         RECT  0.0 12.24 73.14 12.62 ;
         LAYER m4 ;
         RECT  127.84 10.2 128.22 171.06 ;
         LAYER m3 ;
         RECT  151.07 114.61 151.37 114.91 ;
         LAYER m3 ;
         RECT  159.12 107.44 169.02 107.82 ;
         LAYER m4 ;
         RECT  210.8 0.0 211.18 171.06 ;
         LAYER m4 ;
         RECT  167.28 0.0 167.66 171.06 ;
         LAYER m3 ;
         RECT  234.575 105.15 235.065 105.64 ;
         LAYER m3 ;
         RECT  179.865 121.805 180.355 122.295 ;
         LAYER m3 ;
         RECT  89.08 62.56 240.42 62.94 ;
         LAYER m3 ;
         RECT  204.0 145.52 240.42 145.9 ;
         LAYER m3 ;
         RECT  91.07 99.995 91.37 100.295 ;
         LAYER m3 ;
         RECT  190.4 110.16 232.94 110.54 ;
         LAYER m4 ;
         RECT  28.56 0.0 28.94 171.06 ;
         LAYER m3 ;
         RECT  229.16 170.0 240.42 170.38 ;
         LAYER m4 ;
         RECT  131.92 61.2 132.3 171.06 ;
         LAYER m3 ;
         RECT  0.0 51.68 38.46 52.06 ;
         LAYER m3 ;
         RECT  110.38 63.21 110.87 63.7 ;
         LAYER m3 ;
         RECT  124.44 10.88 240.42 11.26 ;
         LAYER m4 ;
         RECT  13.6 0.0 13.98 171.06 ;
         LAYER m3 ;
         RECT  137.765 62.2 138.255 62.69 ;
         LAYER m4 ;
         RECT  194.48 0.0 194.86 171.06 ;
         LAYER m3 ;
         RECT  69.36 102.0 173.1 102.38 ;
         LAYER m4 ;
         RECT  63.92 0.0 64.3 171.06 ;
         LAYER m3 ;
         RECT  105.99 63.21 106.48 63.7 ;
         LAYER m3 ;
         RECT  69.36 115.6 173.1 115.98 ;
         LAYER m3 ;
         RECT  143.41 71.02 143.9 71.51 ;
         LAYER m3 ;
         RECT  104.14 63.21 104.63 63.7 ;
         LAYER m3 ;
         RECT  151.07 96.045 151.37 96.345 ;
         LAYER m4 ;
         RECT  141.44 61.2 141.82 171.06 ;
         LAYER m4 ;
         RECT  231.2 0.0 231.58 171.06 ;
         LAYER m3 ;
         RECT  112.23 63.21 112.72 63.7 ;
         LAYER m3 ;
         RECT  97.9 63.21 98.39 63.7 ;
         LAYER m3 ;
         RECT  179.865 102.055 180.355 102.545 ;
         LAYER m3 ;
         RECT  0.0 106.08 45.26 106.46 ;
         LAYER m3 ;
         RECT  0.0 47.6 240.42 47.98 ;
         LAYER m3 ;
         RECT  196.785 105.97 197.275 106.46 ;
         LAYER m3 ;
         RECT  0.0 42.16 9.9 42.54 ;
         LAYER m3 ;
         RECT  0.0 118.32 62.94 118.7 ;
         LAYER m3 ;
         RECT  0.0 141.44 33.02 141.82 ;
         LAYER m3 ;
         RECT  151.07 111.845 151.37 112.145 ;
         LAYER m3 ;
         RECT  0.0 155.04 240.42 155.42 ;
         LAYER m3 ;
         RECT  123.11 52.305 123.6 52.795 ;
         LAYER m3 ;
         RECT  0.0 21.76 240.42 22.14 ;
         LAYER m3 ;
         RECT  111.52 13.6 240.42 13.98 ;
         LAYER m3 ;
         RECT  151.07 94.86 151.37 95.16 ;
         LAYER m4 ;
         RECT  8.16 0.0 8.54 171.06 ;
         LAYER m4 ;
         RECT  180.88 0.0 181.26 171.06 ;
         LAYER m4 ;
         RECT  223.04 0.0 223.42 171.06 ;
         LAYER m3 ;
         RECT  0.0 100.64 62.94 101.02 ;
         LAYER m4 ;
         RECT  179.52 0.0 179.9 171.06 ;
         LAYER m3 ;
         RECT  135.71 134.91 136.2 135.4 ;
         LAYER m3 ;
         RECT  151.07 124.88 151.37 125.18 ;
         LAYER m3 ;
         RECT  0.0 140.08 240.42 140.46 ;
         LAYER m3 ;
         RECT  202.885 128.35 203.375 128.84 ;
         LAYER m3 ;
         RECT  204.0 131.92 240.42 132.3 ;
         LAYER m3 ;
         RECT  0.0 53.04 94.9 53.42 ;
         LAYER m3 ;
         RECT  179.52 122.4 232.94 122.78 ;
         LAYER m4 ;
         RECT  137.36 61.2 137.74 171.06 ;
         LAYER m3 ;
         RECT  91.07 102.76 91.37 103.06 ;
         LAYER m4 ;
         RECT  119.68 0.0 120.06 171.06 ;
         LAYER m4 ;
         RECT  23.12 0.0 23.5 171.06 ;
         LAYER m3 ;
         RECT  229.84 153.68 240.42 154.06 ;
         LAYER m3 ;
         RECT  0.0 157.76 240.42 158.14 ;
         LAYER m4 ;
         RECT  145.52 0.0 145.9 171.06 ;
         LAYER m4 ;
         RECT  122.4 0.0 122.78 9.22 ;
         LAYER m4 ;
         RECT  220.32 0.0 220.7 171.06 ;
         LAYER m3 ;
         RECT  204.68 58.48 240.42 58.86 ;
         LAYER m3 ;
         RECT  190.935 106.005 191.425 106.495 ;
         LAYER m3 ;
         RECT  39.485 58.97 39.975 59.46 ;
         LAYER m3 ;
         RECT  122.88 71.02 123.37 71.51 ;
         LAYER m3 ;
         RECT  238.255 116.35 238.745 116.84 ;
         LAYER m3 ;
         RECT  9.52 91.12 230.9 91.5 ;
         LAYER m4 ;
         RECT  27.2 0.0 27.58 171.06 ;
         LAYER m3 ;
         RECT  238.255 105.15 238.745 105.64 ;
         LAYER m4 ;
         RECT  44.88 0.0 45.26 171.06 ;
         LAYER m3 ;
         RECT  83.705 0.095 84.195 0.585 ;
         LAYER m3 ;
         RECT  62.085 121.805 62.575 122.295 ;
         LAYER m3 ;
         RECT  69.36 110.16 173.1 110.54 ;
         LAYER m3 ;
         RECT  0.0 88.4 232.94 88.78 ;
         LAYER m3 ;
         RECT  0.0 16.32 96.94 16.7 ;
         LAYER m3 ;
         RECT  149.6 6.8 240.42 7.18 ;
         LAYER m3 ;
         RECT  112.21 71.02 112.7 71.51 ;
         LAYER m3 ;
         RECT  130.425 0.095 130.915 0.585 ;
         LAYER m4 ;
         RECT  235.28 0.0 235.66 171.06 ;
         LAYER m3 ;
         RECT  136.82 134.91 137.31 135.4 ;
         LAYER m4 ;
         RECT  89.76 0.0 90.14 171.06 ;
         LAYER m4 ;
         RECT  57.12 10.2 57.5 171.06 ;
         LAYER m3 ;
         RECT  179.865 119.945 180.355 120.435 ;
         LAYER m4 ;
         RECT  193.12 0.0 193.5 171.06 ;
         LAYER m3 ;
         RECT  99.75 63.21 100.24 63.7 ;
         LAYER m3 ;
         RECT  6.295 88.05 6.785 88.54 ;
         LAYER m3 ;
         RECT  117.64 16.32 240.42 16.7 ;
         LAYER m4 ;
         RECT  171.36 0.0 171.74 171.06 ;
         LAYER m4 ;
         RECT  201.28 0.0 201.66 171.06 ;
         LAYER m3 ;
         RECT  43.52 156.4 240.42 156.78 ;
         LAYER m3 ;
         RECT  0.0 1.36 39.14 1.74 ;
         LAYER m3 ;
         RECT  0.0 68.0 240.42 68.38 ;
         LAYER m4 ;
         RECT  40.8 0.0 41.18 171.06 ;
         LAYER m3 ;
         RECT  0.0 28.56 240.42 28.94 ;
         LAYER m3 ;
         RECT  0.0 59.84 96.26 60.22 ;
         LAYER m4 ;
         RECT  93.84 0.0 94.22 171.06 ;
         LAYER m3 ;
         RECT  0.0 32.64 240.42 33.02 ;
         LAYER m4 ;
         RECT  2.72 0.0 3.1 171.06 ;
         LAYER m4 ;
         RECT  178.16 0.0 178.54 171.06 ;
         LAYER m4 ;
         RECT  123.76 0.0 124.14 171.06 ;
         LAYER m3 ;
         RECT  0.0 92.48 240.42 92.86 ;
         LAYER m3 ;
         RECT  100.3 67.055 100.79 67.545 ;
         LAYER m3 ;
         RECT  175.845 96.095 176.335 96.585 ;
         LAYER m4 ;
         RECT  134.64 61.2 135.02 171.06 ;
         LAYER m4 ;
         RECT  144.16 61.2 144.54 171.06 ;
         LAYER m3 ;
         RECT  99.96 58.48 122.1 58.86 ;
         LAYER m3 ;
         RECT  112.78 67.055 113.27 67.545 ;
         LAYER m3 ;
         RECT  151.07 110.66 151.37 110.96 ;
         LAYER m3 ;
         RECT  204.68 73.44 240.42 73.82 ;
         LAYER m4 ;
         RECT  133.28 8.84 133.66 171.06 ;
         LAYER m3 ;
         RECT  179.52 107.44 230.9 107.82 ;
         LAYER m4 ;
         RECT  238.0 0.0 238.38 171.06 ;
         LAYER m3 ;
         RECT  179.865 113.905 180.355 114.395 ;
         LAYER m3 ;
         RECT  39.485 73.11 39.975 73.6 ;
         LAYER m3 ;
         RECT  9.52 112.88 240.42 113.26 ;
         LAYER m3 ;
         RECT  0.0 133.28 145.22 133.66 ;
         LAYER m3 ;
         RECT  66.105 119.795 66.595 120.285 ;
         LAYER m3 ;
         RECT  234.575 93.95 235.065 94.44 ;
         LAYER m3 ;
         RECT  152.32 4.08 240.42 4.46 ;
         LAYER m4 ;
         RECT  164.56 0.0 164.94 171.06 ;
         LAYER m3 ;
         RECT  190.935 109.955 191.425 110.445 ;
         LAYER m4 ;
         RECT  100.64 0.0 101.02 9.22 ;
         LAYER m3 ;
         RECT  129.12 71.02 129.61 71.51 ;
         LAYER m3 ;
         RECT  144.005 62.2 144.495 62.69 ;
         LAYER m3 ;
         RECT  0.0 70.72 240.42 71.1 ;
         LAYER m3 ;
         RECT  103.59 67.055 104.08 67.545 ;
         LAYER m4 ;
         RECT  172.72 0.0 173.1 171.06 ;
         LAYER m3 ;
         RECT  130.58 134.91 131.07 135.4 ;
         LAYER m3 ;
         RECT  0.0 4.08 50.02 4.46 ;
         LAYER m4 ;
         RECT  21.76 0.0 22.14 171.06 ;
         LAYER m4 ;
         RECT  184.96 0.0 185.34 171.06 ;
         LAYER m3 ;
         RECT  179.52 114.24 230.9 114.62 ;
         LAYER m3 ;
         RECT  91.07 122.51 91.37 122.81 ;
         LAYER m3 ;
         RECT  151.07 103.945 151.37 104.245 ;
         LAYER m4 ;
         RECT  4.08 0.0 4.46 171.06 ;
         LAYER m3 ;
         RECT  0.0 61.2 240.42 61.58 ;
         LAYER m3 ;
         RECT  141.58 63.21 142.07 63.7 ;
         LAYER m3 ;
         RECT  69.36 119.68 173.1 120.06 ;
         LAYER m4 ;
         RECT  72.08 0.0 72.46 171.06 ;
         LAYER m3 ;
         RECT  151.07 113.03 151.37 113.33 ;
         LAYER m3 ;
         RECT  6.295 99.25 6.785 99.74 ;
         LAYER m3 ;
         RECT  0.0 14.96 90.82 15.34 ;
         LAYER m4 ;
         RECT  214.88 0.0 215.26 171.06 ;
         LAYER m3 ;
         RECT  151.07 106.71 151.37 107.01 ;
         LAYER m4 ;
         RECT  84.32 0.0 84.7 171.06 ;
         LAYER m3 ;
         RECT  175.845 107.945 176.335 108.435 ;
         LAYER m3 ;
         RECT  145.52 76.16 240.42 76.54 ;
         LAYER m3 ;
         RECT  62.085 113.905 62.575 114.395 ;
         LAYER m3 ;
         RECT  152.32 9.52 240.42 9.9 ;
         LAYER m3 ;
         RECT  179.865 115.995 180.355 116.485 ;
         LAYER m4 ;
         RECT  224.4 0.0 224.78 171.06 ;
         LAYER m4 ;
         RECT  70.72 0.0 71.1 171.06 ;
         LAYER m3 ;
         RECT  66.105 109.92 66.595 110.41 ;
         LAYER m3 ;
         RECT  175.845 103.995 176.335 104.485 ;
         LAYER m3 ;
         RECT  9.52 107.44 62.94 107.82 ;
         LAYER m3 ;
         RECT  0.0 29.92 240.42 30.3 ;
         LAYER m3 ;
         RECT  141.95 80.69 142.44 81.18 ;
         LAYER m4 ;
         RECT  53.04 0.0 53.42 171.06 ;
         LAYER m3 ;
         RECT  105.4 12.24 114.62 12.62 ;
         LAYER m3 ;
         RECT  62.085 96.245 62.575 96.735 ;
         LAYER m3 ;
         RECT  0.0 9.52 56.14 9.9 ;
         LAYER m3 ;
         RECT  145.52 72.08 240.42 72.46 ;
         LAYER m3 ;
         RECT  151.07 119.745 151.37 120.045 ;
         LAYER m3 ;
         RECT  179.52 100.64 240.42 101.02 ;
         LAYER m3 ;
         RECT  175.845 113.87 176.335 114.36 ;
         LAYER m3 ;
         RECT  0.0 111.52 62.94 111.9 ;
         LAYER m3 ;
         RECT  66.105 115.845 66.595 116.335 ;
         LAYER m3 ;
         RECT  114.24 14.96 240.42 15.34 ;
         LAYER m4 ;
         RECT  55.76 0.0 56.14 171.06 ;
         LAYER m3 ;
         RECT  0.0 110.16 52.06 110.54 ;
         LAYER m3 ;
         RECT  0.0 63.92 240.42 64.3 ;
         LAYER m3 ;
         RECT  137.17 71.02 137.66 71.51 ;
         LAYER m3 ;
         RECT  66.105 105.97 66.595 106.46 ;
         LAYER m4 ;
         RECT  125.12 61.2 125.5 171.06 ;
         LAYER m3 ;
         RECT  91.07 103.945 91.37 104.245 ;
         LAYER m3 ;
         RECT  0.0 13.6 85.38 13.98 ;
         LAYER m3 ;
         RECT  151.07 105.13 151.37 105.43 ;
         LAYER m3 ;
         RECT  69.36 114.24 173.1 114.62 ;
         LAYER m3 ;
         RECT  0.0 146.88 35.74 147.26 ;
         LAYER m3 ;
         RECT  116.62 63.21 117.11 63.7 ;
         LAYER m4 ;
         RECT  104.72 0.0 105.1 171.06 ;
         LAYER m3 ;
         RECT  179.52 104.72 240.42 105.1 ;
         LAYER m3 ;
         RECT  0.0 131.92 94.9 132.3 ;
         LAYER m3 ;
         RECT  151.07 120.93 151.37 121.23 ;
         LAYER m3 ;
         RECT  151.07 123.695 151.37 123.995 ;
         LAYER m3 ;
         RECT  91.07 109.08 91.37 109.38 ;
         LAYER m4 ;
         RECT  183.6 0.0 183.98 171.06 ;
         LAYER m3 ;
         RECT  0.0 163.2 201.66 163.58 ;
         LAYER m3 ;
         RECT  0.0 126.48 92.86 126.86 ;
         LAYER m3 ;
         RECT  45.165 94.12 45.655 94.61 ;
         LAYER m3 ;
         RECT  2.615 110.45 3.105 110.94 ;
         LAYER m3 ;
         RECT  142.105 0.095 142.595 0.585 ;
         LAYER m4 ;
         RECT  129.2 61.2 129.58 171.06 ;
         LAYER m4 ;
         RECT  39.44 0.0 39.82 171.06 ;
         LAYER m4 ;
         RECT  208.08 0.0 208.46 171.06 ;
         LAYER m3 ;
         RECT  36.985 167.53 37.475 168.02 ;
         LAYER m3 ;
         RECT  0.0 159.12 221.38 159.5 ;
         LAYER m4 ;
         RECT  186.32 0.0 186.7 171.06 ;
         LAYER m3 ;
         RECT  205.385 76.35 205.875 76.84 ;
         LAYER m3 ;
         RECT  103.565 62.2 104.055 62.69 ;
         LAYER m3 ;
         RECT  62.085 102.055 62.575 102.545 ;
         LAYER m3 ;
         RECT  0.0 89.76 92.86 90.14 ;
         LAYER m3 ;
         RECT  0.0 46.24 240.42 46.62 ;
         LAYER m3 ;
         RECT  48.665 0.095 49.155 0.585 ;
         LAYER m4 ;
         RECT  199.92 0.0 200.3 171.06 ;
         LAYER m4 ;
         RECT  25.84 0.0 26.22 171.06 ;
         LAYER m3 ;
         RECT  151.07 90.91 151.37 91.21 ;
         LAYER m3 ;
         RECT  97.92 71.02 98.41 71.51 ;
         LAYER m3 ;
         RECT  179.865 94.155 180.355 94.645 ;
         LAYER m3 ;
         RECT  91.07 106.71 91.37 107.01 ;
         LAYER m4 ;
         RECT  165.92 0.0 166.3 171.06 ;
         LAYER m3 ;
         RECT  0.0 10.88 67.7 11.26 ;
         LAYER m3 ;
         RECT  0.0 50.32 240.42 50.7 ;
         LAYER m3 ;
         RECT  69.36 96.56 173.1 96.94 ;
         LAYER m3 ;
         RECT  91.07 119.745 91.37 120.045 ;
         LAYER m3 ;
         RECT  0.0 87.04 240.42 87.42 ;
         LAYER m3 ;
         RECT  69.36 106.08 173.1 106.46 ;
         LAYER m4 ;
         RECT  190.4 0.0 190.78 171.06 ;
         LAYER m4 ;
         RECT  97.92 61.2 98.3 171.06 ;
         LAYER m3 ;
         RECT  0.0 57.12 240.42 57.5 ;
         LAYER m3 ;
         RECT  66.105 100.045 66.595 100.535 ;
         LAYER m3 ;
         RECT  119.02 67.055 119.51 67.545 ;
         LAYER m4 ;
         RECT  175.44 0.0 175.82 171.06 ;
         LAYER m3 ;
         RECT  0.0 168.64 225.46 169.02 ;
         LAYER m3 ;
         RECT  62.085 112.045 62.575 112.535 ;
         LAYER m3 ;
         RECT  69.36 104.72 173.1 105.1 ;
         LAYER m3 ;
         RECT  91.07 123.695 91.37 123.995 ;
         LAYER m4 ;
         RECT  159.12 0.0 159.5 171.06 ;
         LAYER m3 ;
         RECT  91.07 105.13 91.37 105.43 ;
         LAYER m3 ;
         RECT  0.0 99.28 232.94 99.66 ;
         LAYER m4 ;
         RECT  176.8 0.0 177.18 171.06 ;
         LAYER m3 ;
         RECT  107.065 0.095 107.555 0.585 ;
         LAYER m3 ;
         RECT  151.07 118.56 151.37 118.86 ;
         LAYER m3 ;
         RECT  231.88 168.64 240.42 169.02 ;
         LAYER m4 ;
         RECT  114.24 0.0 114.62 171.06 ;
         LAYER m3 ;
         RECT  175.845 105.97 176.335 106.46 ;
         LAYER m3 ;
         RECT  7.48 127.84 240.42 128.22 ;
         LAYER m4 ;
         RECT  168.64 0.0 169.02 171.06 ;
         LAYER m3 ;
         RECT  141.6 144.58 142.09 145.07 ;
         LAYER m3 ;
         RECT  0.0 145.52 151.34 145.9 ;
         LAYER m3 ;
         RECT  123.23 80.69 123.72 81.18 ;
         LAYER m4 ;
         RECT  17.68 0.0 18.06 171.06 ;
         LAYER m3 ;
         RECT  0.0 149.6 201.66 149.98 ;
         LAYER m4 ;
         RECT  87.04 14.96 87.42 171.06 ;
         LAYER m3 ;
         RECT  19.72 42.16 240.42 42.54 ;
         LAYER m4 ;
         RECT  34.0 0.0 34.38 171.06 ;
         LAYER m3 ;
         RECT  0.0 170.0 207.1 170.38 ;
         LAYER m4 ;
         RECT  66.64 0.0 67.02 171.06 ;
         LAYER m4 ;
         RECT  65.28 0.0 65.66 171.06 ;
         LAYER m3 ;
         RECT  179.52 111.52 232.94 111.9 ;
         LAYER m3 ;
         RECT  0.0 80.24 38.46 80.62 ;
         LAYER m4 ;
         RECT  102.0 0.0 102.38 171.06 ;
         LAYER m4 ;
         RECT  126.48 0.0 126.86 171.06 ;
         LAYER m3 ;
         RECT  0.0 122.4 62.94 122.78 ;
         LAYER m3 ;
         RECT  179.52 118.32 240.42 118.7 ;
         LAYER m3 ;
         RECT  40.8 51.68 198.94 52.06 ;
         LAYER m3 ;
         RECT  175.845 119.795 176.335 120.285 ;
         LAYER m3 ;
         RECT  204.68 163.2 217.98 163.58 ;
         LAYER m4 ;
         RECT  155.04 0.0 155.42 171.06 ;
         LAYER m4 ;
         RECT  218.96 0.0 219.34 171.06 ;
         LAYER m3 ;
         RECT  0.0 65.28 96.26 65.66 ;
         LAYER m4 ;
         RECT  136.0 0.0 136.38 171.06 ;
         LAYER m4 ;
         RECT  131.92 0.0 132.3 7.86 ;
         LAYER m3 ;
         RECT  0.0 62.56 38.46 62.94 ;
         LAYER m3 ;
         RECT  43.52 164.56 240.42 164.94 ;
         LAYER m3 ;
         RECT  146.2 8.16 240.42 8.54 ;
         LAYER m3 ;
         RECT  54.505 0.095 54.995 0.585 ;
         LAYER m3 ;
         RECT  179.865 104.145 180.355 104.635 ;
         LAYER m3 ;
         RECT  91.07 92.095 91.37 92.395 ;
         LAYER m3 ;
         RECT  130.95 63.21 131.44 63.7 ;
         LAYER m3 ;
         RECT  97.35 67.055 97.84 67.545 ;
         LAYER m3 ;
         RECT  135.71 80.69 136.2 81.18 ;
         LAYER m3 ;
         RECT  101.225 0.095 101.715 0.585 ;
         LAYER m3 ;
         RECT  62.085 109.955 62.575 110.445 ;
         LAYER m3 ;
         RECT  207.4 55.76 240.42 56.14 ;
         LAYER m4 ;
         RECT  48.96 0.0 49.34 171.06 ;
         LAYER m4 ;
         RECT  96.56 55.08 96.94 171.06 ;
         LAYER m4 ;
         RECT  206.72 0.0 207.1 171.06 ;
         LAYER m3 ;
         RECT  99.73 71.02 100.22 71.51 ;
         LAYER m4 ;
         RECT  50.32 0.0 50.7 171.06 ;
         LAYER m3 ;
         RECT  179.865 98.105 180.355 98.595 ;
         LAYER m3 ;
         RECT  204.68 51.68 240.42 52.06 ;
         LAYER m3 ;
         RECT  77.865 0.095 78.355 0.585 ;
         LAYER m3 ;
         RECT  175.845 109.92 176.335 110.41 ;
         LAYER m3 ;
         RECT  21.08 48.96 240.42 49.34 ;
         LAYER m3 ;
         RECT  135.34 63.21 135.83 63.7 ;
         LAYER m3 ;
         RECT  143.41 144.58 143.9 145.07 ;
         LAYER m3 ;
         RECT  0.0 19.04 240.42 19.42 ;
         LAYER m3 ;
         RECT  15.64 35.36 240.42 35.74 ;
         LAYER m4 ;
         RECT  157.76 0.0 158.14 171.06 ;
         LAYER m3 ;
         RECT  91.07 124.88 91.37 125.18 ;
         LAYER m3 ;
         RECT  116.99 80.69 117.48 81.18 ;
         LAYER m4 ;
         RECT  88.4 0.0 88.78 171.06 ;
         LAYER m3 ;
         RECT  130.93 144.58 131.42 145.07 ;
         LAYER m3 ;
         RECT  95.385 0.095 95.875 0.585 ;
         LAYER m3 ;
         RECT  141.005 62.2 141.495 62.69 ;
         LAYER m4 ;
         RECT  138.72 8.84 139.1 171.06 ;
         LAYER m3 ;
         RECT  0.0 39.44 240.42 39.82 ;
         LAYER m3 ;
         RECT  0.0 114.24 62.94 114.62 ;
         LAYER m3 ;
         RECT  105.97 144.58 106.46 145.07 ;
         LAYER m4 ;
         RECT  78.88 0.0 79.26 171.06 ;
         LAYER m3 ;
         RECT  0.0 8.16 50.02 8.54 ;
         LAYER m4 ;
         RECT  31.28 0.0 31.66 171.06 ;
         LAYER m3 ;
         RECT  66.105 121.77 66.595 122.26 ;
         LAYER m3 ;
         RECT  0.0 54.4 86.06 54.78 ;
         LAYER m3 ;
         RECT  204.68 136.0 240.42 136.38 ;
         LAYER m3 ;
         RECT  186.915 109.92 187.405 110.41 ;
         LAYER m3 ;
         RECT  91.07 118.56 91.37 118.86 ;
         LAYER m3 ;
         RECT  0.0 95.2 240.42 95.58 ;
         LAYER m3 ;
         RECT  0.0 77.52 96.26 77.9 ;
         LAYER m4 ;
         RECT  110.16 61.2 110.54 171.06 ;
         LAYER m3 ;
         RECT  0.0 23.12 240.42 23.5 ;
         LAYER m3 ;
         RECT  130.93 71.02 131.42 71.51 ;
         LAYER m4 ;
         RECT  236.64 0.0 237.02 171.06 ;
         LAYER m3 ;
         RECT  137.19 63.21 137.68 63.7 ;
         LAYER m3 ;
         RECT  112.905 0.095 113.395 0.585 ;
         LAYER m3 ;
         RECT  91.07 111.845 91.37 112.145 ;
         LAYER m3 ;
         RECT  66.105 107.945 66.595 108.435 ;
         LAYER m4 ;
         RECT  107.44 0.0 107.82 171.06 ;
         LAYER m3 ;
         RECT  89.76 69.36 204.38 69.74 ;
         LAYER m3 ;
         RECT  0.0 97.92 52.06 98.3 ;
         LAYER m3 ;
         RECT  62.085 119.945 62.575 120.435 ;
         LAYER m3 ;
         RECT  91.07 93.28 91.37 93.58 ;
         LAYER m3 ;
         RECT  6.295 132.85 6.785 133.34 ;
         LAYER m4 ;
         RECT  125.12 0.0 125.5 10.58 ;
         LAYER m3 ;
         RECT  112.21 144.58 112.7 145.07 ;
         LAYER m3 ;
         RECT  66.105 96.095 66.595 96.585 ;
         LAYER m3 ;
         RECT  66.105 102.02 66.595 102.51 ;
         LAYER m3 ;
         RECT  69.36 118.32 173.1 118.7 ;
         LAYER m3 ;
         RECT  55.035 98.07 55.525 98.56 ;
         LAYER m4 ;
         RECT  19.04 0.0 19.42 171.06 ;
         LAYER m3 ;
         RECT  0.0 78.88 240.42 79.26 ;
         LAYER m3 ;
         RECT  151.07 99.995 151.37 100.295 ;
         LAYER m3 ;
         RECT  7.48 104.72 62.94 105.1 ;
         LAYER m4 ;
         RECT  12.24 0.0 12.62 171.06 ;
         LAYER m3 ;
         RECT  234.575 116.35 235.065 116.84 ;
         LAYER m3 ;
         RECT  179.865 117.855 180.355 118.345 ;
         LAYER m4 ;
         RECT  202.64 0.0 203.02 171.06 ;
         LAYER m3 ;
         RECT  151.07 109.08 151.37 109.38 ;
         LAYER m3 ;
         RECT  124.69 71.02 125.18 71.51 ;
         LAYER m3 ;
         RECT  146.88 85.68 230.9 86.06 ;
         LAYER m3 ;
         RECT  66.105 113.87 66.595 114.36 ;
         LAYER m3 ;
         RECT  179.865 96.245 180.355 96.735 ;
         LAYER m4 ;
         RECT  111.52 0.0 111.9 171.06 ;
         LAYER m4 ;
         RECT  140.08 0.0 140.46 171.06 ;
         LAYER m3 ;
         RECT  110.4 71.02 110.89 71.51 ;
         LAYER m3 ;
         RECT  136.265 0.095 136.755 0.585 ;
         LAYER m3 ;
         RECT  204.68 149.6 240.42 149.98 ;
         LAYER m3 ;
         RECT  69.36 103.36 173.1 103.74 ;
         LAYER m3 ;
         RECT  104.51 80.69 105.0 81.18 ;
         LAYER m4 ;
         RECT  82.96 0.0 83.34 171.06 ;
         LAYER m3 ;
         RECT  0.0 150.96 240.42 151.34 ;
         LAYER m4 ;
         RECT  163.2 0.0 163.58 171.06 ;
         LAYER m3 ;
         RECT  118.1 80.69 118.59 81.18 ;
         LAYER m3 ;
         RECT  122.285 62.2 122.775 62.69 ;
         LAYER m3 ;
         RECT  98.27 134.91 98.76 135.4 ;
         LAYER m3 ;
         RECT  136.82 80.69 137.31 81.18 ;
         LAYER m3 ;
         RECT  110.75 80.69 111.24 81.18 ;
         LAYER m4 ;
         RECT  233.92 0.0 234.3 171.06 ;
         LAYER m3 ;
         RECT  99.38 80.69 99.87 81.18 ;
         LAYER m3 ;
         RECT  91.07 110.66 91.37 110.96 ;
         LAYER m3 ;
         RECT  129.12 144.58 129.61 145.07 ;
         LAYER m3 ;
         RECT  91.07 120.93 91.37 121.23 ;
         LAYER m4 ;
         RECT  0.0 0.0 0.38 171.06 ;
         LAYER m4 ;
         RECT  108.8 0.0 109.18 171.06 ;
         LAYER m4 ;
         RECT  116.96 0.0 117.34 171.06 ;
         LAYER m3 ;
         RECT  42.84 142.8 96.26 143.18 ;
         LAYER m3 ;
         RECT  155.72 134.64 240.42 135.02 ;
         LAYER m3 ;
         RECT  175.845 98.07 176.335 98.56 ;
         LAYER m4 ;
         RECT  106.08 61.2 106.46 171.06 ;
         LAYER m3 ;
         RECT  122.88 144.58 123.37 145.07 ;
         LAYER m3 ;
         RECT  9.52 130.56 240.42 130.94 ;
         LAYER m3 ;
         RECT  105.62 80.69 106.11 81.18 ;
         LAYER m3 ;
         RECT  0.0 164.56 38.46 164.94 ;
         LAYER m3 ;
         RECT  0.0 74.8 200.98 75.18 ;
         LAYER m4 ;
         RECT  9.52 0.0 9.9 171.06 ;
         LAYER m3 ;
         RECT  109.83 67.055 110.32 67.545 ;
         LAYER m3 ;
         RECT  0.0 55.76 38.46 56.14 ;
         LAYER m3 ;
         RECT  91.07 107.895 91.37 108.195 ;
         LAYER m3 ;
         RECT  97.92 53.04 119.38 53.42 ;
         LAYER m3 ;
         RECT  40.8 66.64 240.42 67.02 ;
         LAYER m4 ;
         RECT  46.24 0.0 46.62 171.06 ;
         LAYER m3 ;
         RECT  143.98 67.055 144.47 67.545 ;
         LAYER m4 ;
         RECT  130.56 0.0 130.94 171.06 ;
         LAYER m3 ;
         RECT  66.105 94.12 66.595 94.61 ;
         LAYER m3 ;
         RECT  62.085 98.105 62.575 98.595 ;
         LAYER m3 ;
         RECT  110.4 144.58 110.89 145.07 ;
         LAYER m3 ;
         RECT  40.8 80.24 230.9 80.62 ;
         LAYER m3 ;
         RECT  186.915 105.97 187.405 106.46 ;
         LAYER m3 ;
         RECT  0.375 30.68 0.865 31.17 ;
         LAYER m3 ;
         RECT  204.68 65.28 240.42 65.66 ;
         LAYER m4 ;
         RECT  156.4 0.0 156.78 171.06 ;
         LAYER m3 ;
         RECT  186.915 98.07 187.405 98.56 ;
         LAYER m3 ;
         RECT  98.27 80.69 98.76 81.18 ;
         LAYER m3 ;
         RECT  111.86 80.69 112.35 81.18 ;
         LAYER m3 ;
         RECT  151.07 97.23 151.37 97.53 ;
         LAYER m3 ;
         RECT  0.0 48.96 11.94 49.34 ;
         LAYER m4 ;
         RECT  227.12 0.0 227.5 171.06 ;
         LAYER m3 ;
         RECT  204.0 138.72 240.42 139.1 ;
         LAYER m3 ;
         RECT  0.0 66.64 38.46 67.02 ;
         LAYER m3 ;
         RECT  240.495 170.78 240.985 171.27 ;
         LAYER m4 ;
         RECT  42.16 0.0 42.54 171.06 ;
         LAYER m3 ;
         RECT  179.52 96.56 230.9 96.94 ;
         LAYER m3 ;
         RECT  9.52 123.76 240.42 124.14 ;
         LAYER m3 ;
         RECT  45.165 105.97 45.655 106.46 ;
         LAYER m3 ;
         RECT  137.17 144.58 137.66 145.07 ;
         LAYER m3 ;
         RECT  66.185 0.095 66.675 0.585 ;
         LAYER m4 ;
         RECT  43.52 0.0 43.9 171.06 ;
         LAYER m3 ;
         RECT  129.1 63.21 129.59 63.7 ;
         LAYER m3 ;
         RECT  66.105 98.07 66.595 98.56 ;
         LAYER m3 ;
         RECT  125.12 58.48 198.94 58.86 ;
         LAYER m3 ;
         RECT  202.885 170.77 203.375 171.26 ;
         LAYER m3 ;
         RECT  6.295 110.45 6.785 110.94 ;
         LAYER m4 ;
         RECT  1.36 0.0 1.74 171.06 ;
         LAYER m3 ;
         RECT  40.8 38.08 240.42 38.46 ;
         LAYER m3 ;
         RECT  179.865 108.095 180.355 108.585 ;
         LAYER m4 ;
         RECT  228.48 0.0 228.86 171.06 ;
         LAYER m4 ;
         RECT  74.8 12.92 75.18 171.06 ;
         LAYER m3 ;
         RECT  55.035 94.12 55.525 94.61 ;
         LAYER m4 ;
         RECT  47.6 0.0 47.98 171.06 ;
         LAYER m3 ;
         RECT  0.0 144.16 240.42 144.54 ;
         LAYER m3 ;
         RECT  141.03 67.055 141.52 67.545 ;
         LAYER m3 ;
         RECT  0.0 0.0 240.42 0.38 ;
         LAYER m3 ;
         RECT  175.845 117.82 176.335 118.31 ;
         LAYER m3 ;
         RECT  90.44 55.76 204.38 56.14 ;
         LAYER m3 ;
         RECT  190.935 98.105 191.425 98.595 ;
         LAYER m4 ;
         RECT  217.6 0.0 217.98 171.06 ;
         LAYER m3 ;
         RECT  145.52 142.8 240.42 143.18 ;
         LAYER m3 ;
         RECT  100.325 62.2 100.815 62.69 ;
         LAYER m4 ;
         RECT  81.6 0.0 81.98 171.06 ;
         LAYER m4 ;
         RECT  152.32 0.0 152.7 171.06 ;
         LAYER m3 ;
         RECT  91.07 94.86 91.37 95.16 ;
         LAYER m4 ;
         RECT  197.2 0.0 197.58 171.06 ;
         LAYER m3 ;
         RECT  39.485 44.83 39.975 45.32 ;
         LAYER m3 ;
         RECT  151.07 122.51 151.37 122.81 ;
         LAYER m3 ;
         RECT  39.485 30.69 39.975 31.18 ;
         LAYER m3 ;
         RECT  179.865 109.955 180.355 110.445 ;
         LAYER m3 ;
         RECT  149.6 89.76 240.42 90.14 ;
         LAYER m3 ;
         RECT  88.4 84.32 240.42 84.7 ;
         LAYER m4 ;
         RECT  16.32 0.0 16.7 171.06 ;
         LAYER m3 ;
         RECT  0.0 44.88 240.42 45.26 ;
         LAYER m4 ;
         RECT  38.08 0.0 38.46 171.06 ;
         LAYER m4 ;
         RECT  58.48 0.0 58.86 171.06 ;
         LAYER m3 ;
         RECT  7.48 115.6 62.94 115.98 ;
         LAYER m3 ;
         RECT  9.52 119.68 62.94 120.06 ;
         LAYER m3 ;
         RECT  69.36 122.4 173.1 122.78 ;
         LAYER m3 ;
         RECT  91.07 101.18 91.37 101.48 ;
         LAYER m3 ;
         RECT  0.0 152.32 240.42 152.7 ;
         LAYER m3 ;
         RECT  0.0 20.4 240.42 20.78 ;
         LAYER m3 ;
         RECT  130.58 80.69 131.07 81.18 ;
         LAYER m4 ;
         RECT  73.44 0.0 73.82 171.06 ;
         LAYER m3 ;
         RECT  116.99 134.91 117.48 135.4 ;
         LAYER m3 ;
         RECT  106.54 67.055 107.03 67.545 ;
         LAYER m4 ;
         RECT  144.16 0.0 144.54 7.86 ;
         LAYER m4 ;
         RECT  68.0 0.0 68.38 171.06 ;
         LAYER m3 ;
         RECT  238.255 93.95 238.745 94.44 ;
         LAYER m3 ;
         RECT  0.0 153.68 220.02 154.06 ;
         LAYER m4 ;
         RECT  100.64 61.2 101.02 171.06 ;
         LAYER m4 ;
         RECT  204.0 0.0 204.38 171.06 ;
         LAYER m4 ;
         RECT  59.84 0.0 60.22 171.06 ;
         LAYER m3 ;
         RECT  128.525 62.2 129.015 62.69 ;
         LAYER m4 ;
         RECT  232.56 0.0 232.94 171.06 ;
         LAYER m3 ;
         RECT  124.34 134.91 124.83 135.4 ;
         LAYER m3 ;
         RECT  134.765 62.2 135.255 62.69 ;
         LAYER m3 ;
         RECT  0.0 125.12 230.9 125.5 ;
         LAYER m3 ;
         RECT  0.0 156.4 38.46 156.78 ;
         LAYER m4 ;
         RECT  195.84 0.0 196.22 171.06 ;
         LAYER m3 ;
         RECT  202.885 142.49 203.375 142.98 ;
         LAYER m3 ;
         RECT  66.105 103.995 66.595 104.485 ;
         LAYER m3 ;
         RECT  55.035 109.92 55.525 110.41 ;
         LAYER m3 ;
         RECT  0.0 5.44 240.42 5.82 ;
         LAYER m3 ;
         RECT  14.28 40.8 240.42 41.18 ;
         LAYER m3 ;
         RECT  65.96 108.8 176.5 109.18 ;
         LAYER m3 ;
         RECT  0.0 160.48 35.74 160.86 ;
         LAYER m3 ;
         RECT  0.0 34.0 240.42 34.38 ;
         LAYER m3 ;
         RECT  124.71 63.21 125.2 63.7 ;
         LAYER m4 ;
         RECT  118.32 0.0 118.7 171.06 ;
         LAYER m3 ;
         RECT  152.32 1.36 240.42 1.74 ;
         LAYER m3 ;
         RECT  175.845 94.12 176.335 94.61 ;
         LAYER m4 ;
         RECT  122.4 61.2 122.78 171.06 ;
         LAYER m4 ;
         RECT  112.88 0.0 113.26 13.98 ;
         LAYER m3 ;
         RECT  69.695 107.725 70.185 108.215 ;
         LAYER m3 ;
         RECT  207.4 69.36 240.42 69.74 ;
         LAYER m3 ;
         RECT  133.28 9.52 142.5 9.9 ;
         LAYER m3 ;
         RECT  38.08 160.48 240.42 160.86 ;
         LAYER m4 ;
         RECT  189.04 0.0 189.42 171.06 ;
         LAYER m3 ;
         RECT  2.615 88.05 3.105 88.54 ;
         LAYER m3 ;
         RECT  122.86 63.21 123.35 63.7 ;
         LAYER m3 ;
         RECT  124.34 80.69 124.83 81.18 ;
         LAYER m3 ;
         RECT  51.015 98.105 51.505 98.595 ;
         LAYER m3 ;
         RECT  145.52 59.84 240.42 60.22 ;
         LAYER m3 ;
         RECT  228.48 159.12 240.42 159.5 ;
         LAYER m3 ;
         RECT  175.845 102.02 176.335 102.51 ;
         LAYER m4 ;
         RECT  187.68 0.0 188.06 171.06 ;
         LAYER m3 ;
         RECT  141.95 134.91 142.44 135.4 ;
         LAYER m4 ;
         RECT  229.84 0.0 230.22 171.06 ;
         LAYER m3 ;
         RECT  151.07 93.28 151.37 93.58 ;
         LAYER m3 ;
         RECT  1.36 38.08 11.26 38.46 ;
         LAYER m3 ;
         RECT  125.285 62.2 125.775 62.69 ;
         LAYER m3 ;
         RECT  116.045 62.2 116.535 62.69 ;
         LAYER m4 ;
         RECT  14.96 0.0 15.34 171.06 ;
         LAYER m3 ;
         RECT  0.0 6.8 47.3 7.18 ;
         LAYER m4 ;
         RECT  85.68 0.0 86.06 171.06 ;
         LAYER m4 ;
         RECT  209.44 0.0 209.82 171.06 ;
         LAYER m4 ;
         RECT  51.68 8.84 52.06 171.06 ;
         LAYER m3 ;
         RECT  105.97 71.02 106.46 71.51 ;
         LAYER m3 ;
         RECT  179.52 115.6 240.42 115.98 ;
         LAYER m4 ;
         RECT  153.68 0.0 154.06 171.06 ;
         LAYER m3 ;
         RECT  229.84 163.2 239.06 163.58 ;
         LAYER m3 ;
         RECT  151.07 107.895 151.37 108.195 ;
         LAYER m4 ;
         RECT  213.52 0.0 213.9 171.06 ;
         LAYER m3 ;
         RECT  0.0 2.72 240.42 3.1 ;
         LAYER m4 ;
         RECT  5.44 0.0 5.82 171.06 ;
         LAYER m3 ;
         RECT  51.015 94.155 51.505 94.645 ;
         LAYER m3 ;
         RECT  143.06 80.69 143.55 81.18 ;
         LAYER m3 ;
         RECT  175.845 115.845 176.335 116.335 ;
         LAYER m3 ;
         RECT  66.105 111.895 66.595 112.385 ;
         LAYER m3 ;
         RECT  135.36 144.58 135.85 145.07 ;
         LAYER m4 ;
         RECT  216.24 0.0 216.62 171.06 ;
         LAYER m3 ;
         RECT  42.16 141.44 240.42 141.82 ;
         LAYER m4 ;
         RECT  239.36 0.0 239.74 171.06 ;
         LAYER m3 ;
         RECT  0.0 58.48 96.94 58.86 ;
         LAYER m3 ;
         RECT  175.845 100.045 176.335 100.535 ;
         LAYER m4 ;
         RECT  91.12 0.0 91.5 171.06 ;
         LAYER m4 ;
         RECT  80.24 13.6 80.62 171.06 ;
         LAYER m3 ;
         RECT  72.025 0.095 72.515 0.585 ;
         LAYER m4 ;
         RECT  170.0 0.0 170.38 171.06 ;
         LAYER m3 ;
         RECT  69.36 97.92 173.1 98.3 ;
         LAYER m3 ;
         RECT  91.07 98.81 91.37 99.11 ;
         LAYER m3 ;
         RECT  109.805 62.2 110.295 62.69 ;
         LAYER m4 ;
         RECT  62.56 19.04 62.94 171.06 ;
         LAYER m3 ;
         RECT  137.74 67.055 138.23 67.545 ;
         LAYER m3 ;
         RECT  175.845 111.895 176.335 112.385 ;
         LAYER m3 ;
         RECT  143.43 63.21 143.92 63.7 ;
         LAYER m3 ;
         RECT  151.07 102.76 151.37 103.06 ;
         LAYER m3 ;
         RECT  0.0 142.8 38.46 143.18 ;
         LAYER m3 ;
         RECT  128.55 67.055 129.04 67.545 ;
         LAYER m3 ;
         RECT  0.0 148.24 240.42 148.62 ;
         LAYER m3 ;
         RECT  0.0 27.2 240.42 27.58 ;
         LAYER m3 ;
         RECT  9.52 96.56 62.94 96.94 ;
         LAYER m3 ;
         RECT  91.07 114.61 91.37 114.91 ;
         LAYER m3 ;
         RECT  51.015 106.005 51.505 106.495 ;
         LAYER m4 ;
         RECT  103.36 61.2 103.74 171.06 ;
         LAYER m3 ;
         RECT  151.07 115.795 151.37 116.095 ;
         LAYER m3 ;
         RECT  36.985 139.25 37.475 139.74 ;
         LAYER m3 ;
         RECT  110.75 134.91 111.24 135.4 ;
         LAYER m3 ;
         RECT  0.0 81.6 85.38 81.98 ;
         LAYER m4 ;
         RECT  77.52 0.0 77.9 171.06 ;
         LAYER m3 ;
         RECT  99.28 17.68 240.42 18.06 ;
         LAYER m3 ;
         RECT  66.105 117.82 66.595 118.31 ;
         LAYER m4 ;
         RECT  99.28 0.0 99.66 171.06 ;
         LAYER m3 ;
         RECT  129.47 134.91 129.96 135.4 ;
         LAYER m4 ;
         RECT  142.8 0.0 143.18 171.06 ;
         LAYER m3 ;
         RECT  34.68 31.28 240.42 31.66 ;
         LAYER m4 ;
         RECT  149.6 0.0 149.98 171.06 ;
         LAYER m3 ;
         RECT  135.36 71.02 135.85 71.51 ;
         LAYER m3 ;
         RECT  104.16 71.02 104.65 71.51 ;
         LAYER m4 ;
         RECT  121.04 55.08 121.42 171.06 ;
         LAYER m3 ;
         RECT  89.545 0.095 90.035 0.585 ;
         LAYER m3 ;
         RECT  73.44 107.44 83.34 107.82 ;
         LAYER m3 ;
         RECT  39.485 87.25 39.975 87.74 ;
         LAYER m3 ;
         RECT  179.865 100.195 180.355 100.685 ;
         LAYER m3 ;
         RECT  0.0 69.36 38.46 69.74 ;
         LAYER m3 ;
         RECT  91.07 97.23 91.37 97.53 ;
         LAYER m3 ;
         RECT  0.0 137.36 240.42 137.74 ;
         LAYER m3 ;
         RECT  143.06 134.91 143.55 135.4 ;
         LAYER m3 ;
         RECT  179.865 106.005 180.355 106.495 ;
         LAYER m3 ;
         RECT  123.23 134.91 123.72 135.4 ;
         LAYER m3 ;
         RECT  179.52 102.0 230.9 102.38 ;
         LAYER m4 ;
         RECT  205.36 0.0 205.74 171.06 ;
         LAYER m3 ;
         RECT  131.525 62.2 132.015 62.69 ;
         LAYER m3 ;
         RECT  36.985 153.39 37.475 153.88 ;
         LAYER m3 ;
         RECT  123.08 53.04 240.42 53.42 ;
         LAYER m3 ;
         RECT  197.2 93.84 240.42 94.22 ;
         LAYER m3 ;
         RECT  0.0 36.72 240.42 37.1 ;
         LAYER m3 ;
         RECT  0.0 121.04 240.42 121.42 ;
         LAYER m4 ;
         RECT  32.64 0.0 33.02 171.06 ;
         LAYER m4 ;
         RECT  115.6 61.2 115.98 171.06 ;
         LAYER m4 ;
         RECT  69.36 11.56 69.74 171.06 ;
         LAYER m3 ;
         RECT  62.085 104.145 62.575 104.635 ;
         LAYER m3 ;
         RECT  0.0 116.96 240.42 117.34 ;
         LAYER m3 ;
         RECT  129.47 80.69 129.96 81.18 ;
         LAYER m3 ;
         RECT  151.07 98.81 151.37 99.11 ;
         LAYER m3 ;
         RECT  151.07 101.18 151.37 101.48 ;
         LAYER m3 ;
         RECT  7.48 93.84 45.26 94.22 ;
         LAYER m3 ;
         RECT  104.51 134.91 105.0 135.4 ;
         LAYER m3 ;
         RECT  179.52 108.8 240.42 109.18 ;
         LAYER m4 ;
         RECT  198.56 0.0 198.94 171.06 ;
         LAYER m4 ;
         RECT  6.8 0.0 7.18 171.06 ;
         LAYER m3 ;
         RECT  151.07 92.095 151.37 92.395 ;
         LAYER m3 ;
         RECT  99.38 134.91 99.87 135.4 ;
         LAYER m3 ;
         RECT  0.0 129.2 95.58 129.58 ;
         LAYER m4 ;
         RECT  61.2 0.0 61.58 171.06 ;
         LAYER m4 ;
         RECT  92.48 16.32 92.86 171.06 ;
         LAYER m3 ;
         RECT  234.575 82.75 235.065 83.24 ;
         LAYER m3 ;
         RECT  234.575 127.55 235.065 128.04 ;
         LAYER m3 ;
         RECT  111.86 134.91 112.35 135.4 ;
         LAYER m4 ;
         RECT  35.36 0.0 35.74 171.06 ;
         LAYER m3 ;
         RECT  238.255 82.75 238.745 83.24 ;
         LAYER m3 ;
         RECT  190.4 97.92 240.42 98.3 ;
         LAYER m3 ;
         RECT  190.935 94.155 191.425 94.645 ;
      END
   END gnd
   OBS
   LAYER  m1 ;
      RECT  98.45 92.73 98.66 93.14 ;
      RECT  96.05 91.725 96.26 92.055 ;
      RECT  99.095 92.64 99.17 94.345 ;
      RECT  99.01 93.225 99.095 93.635 ;
      RECT  98.09 91.725 98.27 92.64 ;
      POLYGON  99.095 91.725 99.095 92.055 98.66 92.055 98.66 92.435 99.095 92.435 99.095 92.64 99.17 92.64 99.17 91.725 99.095 91.725 ;
      RECT  99.17 92.64 99.38 94.345 ;
      POLYGON  98.66 92.73 98.66 93.14 98.835 93.14 98.915 93.06 98.915 92.73 98.66 92.73 ;
      RECT  96.05 92.64 96.26 94.345 ;
      RECT  97.73 91.725 97.91 92.64 ;
      RECT  96.65 92.64 96.83 94.345 ;
      RECT  98.45 93.72 98.66 94.13 ;
      RECT  99.17 92.435 99.38 92.64 ;
      RECT  96.26 92.64 96.47 94.345 ;
      RECT  98.45 92.055 98.66 92.435 ;
      RECT  97.01 92.64 97.19 94.345 ;
      RECT  97.73 92.64 97.91 94.345 ;
      RECT  97.01 91.725 97.19 92.64 ;
      RECT  99.17 91.725 99.38 92.055 ;
      RECT  97.37 92.64 97.55 94.345 ;
      RECT  97.37 91.725 97.55 92.64 ;
      RECT  96.05 92.435 96.26 92.64 ;
      RECT  99.17 92.055 99.38 92.435 ;
      RECT  98.09 92.64 98.27 94.345 ;
      RECT  96.26 92.435 96.47 92.64 ;
      RECT  96.05 92.055 96.26 92.435 ;
      POLYGON  98.66 93.72 98.66 94.13 98.915 94.13 98.915 93.8 98.835 93.72 98.66 93.72 ;
      RECT  96.65 91.725 96.83 92.64 ;
      RECT  96.26 91.725 96.47 92.055 ;
      RECT  96.26 92.055 96.47 92.435 ;
      RECT  98.45 95.71 98.66 95.3 ;
      RECT  96.05 96.715 96.26 96.385 ;
      RECT  99.095 95.8 99.17 94.095 ;
      RECT  99.01 95.215 99.095 94.805 ;
      RECT  98.09 96.715 98.27 95.8 ;
      POLYGON  99.095 96.715 99.095 96.385 98.66 96.385 98.66 96.005 99.095 96.005 99.095 95.8 99.17 95.8 99.17 96.715 99.095 96.715 ;
      RECT  99.17 95.8 99.38 94.095 ;
      POLYGON  98.66 95.71 98.66 95.3 98.835 95.3 98.915 95.38 98.915 95.71 98.66 95.71 ;
      RECT  96.05 95.8 96.26 94.095 ;
      RECT  97.73 96.715 97.91 95.8 ;
      RECT  96.65 95.8 96.83 94.095 ;
      RECT  98.45 94.72 98.66 94.31 ;
      RECT  99.17 96.005 99.38 95.8 ;
      RECT  96.26 95.8 96.47 94.095 ;
      RECT  98.45 96.385 98.66 96.005 ;
      RECT  97.01 95.8 97.19 94.095 ;
      RECT  97.73 95.8 97.91 94.095 ;
      RECT  97.01 96.715 97.19 95.8 ;
      RECT  99.17 96.715 99.38 96.385 ;
      RECT  97.37 95.8 97.55 94.095 ;
      RECT  97.37 96.715 97.55 95.8 ;
      RECT  96.05 96.005 96.26 95.8 ;
      RECT  99.17 96.385 99.38 96.005 ;
      RECT  98.09 95.8 98.27 94.095 ;
      RECT  96.26 96.005 96.47 95.8 ;
      RECT  96.05 96.385 96.26 96.005 ;
      POLYGON  98.66 94.72 98.66 94.31 98.915 94.31 98.915 94.64 98.835 94.72 98.66 94.72 ;
      RECT  96.65 96.715 96.83 95.8 ;
      RECT  96.26 96.715 96.47 96.385 ;
      RECT  96.26 96.385 96.47 96.005 ;
      RECT  98.45 96.68 98.66 97.09 ;
      RECT  96.05 95.675 96.26 96.005 ;
      RECT  99.095 96.59 99.17 98.295 ;
      RECT  99.01 97.175 99.095 97.585 ;
      RECT  98.09 95.675 98.27 96.59 ;
      POLYGON  99.095 95.675 99.095 96.005 98.66 96.005 98.66 96.385 99.095 96.385 99.095 96.59 99.17 96.59 99.17 95.675 99.095 95.675 ;
      RECT  99.17 96.59 99.38 98.295 ;
      POLYGON  98.66 96.68 98.66 97.09 98.835 97.09 98.915 97.01 98.915 96.68 98.66 96.68 ;
      RECT  96.05 96.59 96.26 98.295 ;
      RECT  97.73 95.675 97.91 96.59 ;
      RECT  96.65 96.59 96.83 98.295 ;
      RECT  98.45 97.67 98.66 98.08 ;
      RECT  99.17 96.385 99.38 96.59 ;
      RECT  96.26 96.59 96.47 98.295 ;
      RECT  98.45 96.005 98.66 96.385 ;
      RECT  97.01 96.59 97.19 98.295 ;
      RECT  97.73 96.59 97.91 98.295 ;
      RECT  97.01 95.675 97.19 96.59 ;
      RECT  99.17 95.675 99.38 96.005 ;
      RECT  97.37 96.59 97.55 98.295 ;
      RECT  97.37 95.675 97.55 96.59 ;
      RECT  96.05 96.385 96.26 96.59 ;
      RECT  99.17 96.005 99.38 96.385 ;
      RECT  98.09 96.59 98.27 98.295 ;
      RECT  96.26 96.385 96.47 96.59 ;
      RECT  96.05 96.005 96.26 96.385 ;
      POLYGON  98.66 97.67 98.66 98.08 98.915 98.08 98.915 97.75 98.835 97.67 98.66 97.67 ;
      RECT  96.65 95.675 96.83 96.59 ;
      RECT  96.26 95.675 96.47 96.005 ;
      RECT  96.26 96.005 96.47 96.385 ;
      RECT  98.45 99.66 98.66 99.25 ;
      RECT  96.05 100.665 96.26 100.335 ;
      RECT  99.095 99.75 99.17 98.045 ;
      RECT  99.01 99.165 99.095 98.755 ;
      RECT  98.09 100.665 98.27 99.75 ;
      POLYGON  99.095 100.665 99.095 100.335 98.66 100.335 98.66 99.955 99.095 99.955 99.095 99.75 99.17 99.75 99.17 100.665 99.095 100.665 ;
      RECT  99.17 99.75 99.38 98.045 ;
      POLYGON  98.66 99.66 98.66 99.25 98.835 99.25 98.915 99.33 98.915 99.66 98.66 99.66 ;
      RECT  96.05 99.75 96.26 98.045 ;
      RECT  97.73 100.665 97.91 99.75 ;
      RECT  96.65 99.75 96.83 98.045 ;
      RECT  98.45 98.67 98.66 98.26 ;
      RECT  99.17 99.955 99.38 99.75 ;
      RECT  96.26 99.75 96.47 98.045 ;
      RECT  98.45 100.335 98.66 99.955 ;
      RECT  97.01 99.75 97.19 98.045 ;
      RECT  97.73 99.75 97.91 98.045 ;
      RECT  97.01 100.665 97.19 99.75 ;
      RECT  99.17 100.665 99.38 100.335 ;
      RECT  97.37 99.75 97.55 98.045 ;
      RECT  97.37 100.665 97.55 99.75 ;
      RECT  96.05 99.955 96.26 99.75 ;
      RECT  99.17 100.335 99.38 99.955 ;
      RECT  98.09 99.75 98.27 98.045 ;
      RECT  96.26 99.955 96.47 99.75 ;
      RECT  96.05 100.335 96.26 99.955 ;
      POLYGON  98.66 98.67 98.66 98.26 98.915 98.26 98.915 98.59 98.835 98.67 98.66 98.67 ;
      RECT  96.65 100.665 96.83 99.75 ;
      RECT  96.26 100.665 96.47 100.335 ;
      RECT  96.26 100.335 96.47 99.955 ;
      RECT  98.45 100.63 98.66 101.04 ;
      RECT  96.05 99.625 96.26 99.955 ;
      RECT  99.095 100.54 99.17 102.245 ;
      RECT  99.01 101.125 99.095 101.535 ;
      RECT  98.09 99.625 98.27 100.54 ;
      POLYGON  99.095 99.625 99.095 99.955 98.66 99.955 98.66 100.335 99.095 100.335 99.095 100.54 99.17 100.54 99.17 99.625 99.095 99.625 ;
      RECT  99.17 100.54 99.38 102.245 ;
      POLYGON  98.66 100.63 98.66 101.04 98.835 101.04 98.915 100.96 98.915 100.63 98.66 100.63 ;
      RECT  96.05 100.54 96.26 102.245 ;
      RECT  97.73 99.625 97.91 100.54 ;
      RECT  96.65 100.54 96.83 102.245 ;
      RECT  98.45 101.62 98.66 102.03 ;
      RECT  99.17 100.335 99.38 100.54 ;
      RECT  96.26 100.54 96.47 102.245 ;
      RECT  98.45 99.955 98.66 100.335 ;
      RECT  97.01 100.54 97.19 102.245 ;
      RECT  97.73 100.54 97.91 102.245 ;
      RECT  97.01 99.625 97.19 100.54 ;
      RECT  99.17 99.625 99.38 99.955 ;
      RECT  97.37 100.54 97.55 102.245 ;
      RECT  97.37 99.625 97.55 100.54 ;
      RECT  96.05 100.335 96.26 100.54 ;
      RECT  99.17 99.955 99.38 100.335 ;
      RECT  98.09 100.54 98.27 102.245 ;
      RECT  96.26 100.335 96.47 100.54 ;
      RECT  96.05 99.955 96.26 100.335 ;
      POLYGON  98.66 101.62 98.66 102.03 98.915 102.03 98.915 101.7 98.835 101.62 98.66 101.62 ;
      RECT  96.65 99.625 96.83 100.54 ;
      RECT  96.26 99.625 96.47 99.955 ;
      RECT  96.26 99.955 96.47 100.335 ;
      RECT  98.45 103.61 98.66 103.2 ;
      RECT  96.05 104.615 96.26 104.285 ;
      RECT  99.095 103.7 99.17 101.995 ;
      RECT  99.01 103.115 99.095 102.705 ;
      RECT  98.09 104.615 98.27 103.7 ;
      POLYGON  99.095 104.615 99.095 104.285 98.66 104.285 98.66 103.905 99.095 103.905 99.095 103.7 99.17 103.7 99.17 104.615 99.095 104.615 ;
      RECT  99.17 103.7 99.38 101.995 ;
      POLYGON  98.66 103.61 98.66 103.2 98.835 103.2 98.915 103.28 98.915 103.61 98.66 103.61 ;
      RECT  96.05 103.7 96.26 101.995 ;
      RECT  97.73 104.615 97.91 103.7 ;
      RECT  96.65 103.7 96.83 101.995 ;
      RECT  98.45 102.62 98.66 102.21 ;
      RECT  99.17 103.905 99.38 103.7 ;
      RECT  96.26 103.7 96.47 101.995 ;
      RECT  98.45 104.285 98.66 103.905 ;
      RECT  97.01 103.7 97.19 101.995 ;
      RECT  97.73 103.7 97.91 101.995 ;
      RECT  97.01 104.615 97.19 103.7 ;
      RECT  99.17 104.615 99.38 104.285 ;
      RECT  97.37 103.7 97.55 101.995 ;
      RECT  97.37 104.615 97.55 103.7 ;
      RECT  96.05 103.905 96.26 103.7 ;
      RECT  99.17 104.285 99.38 103.905 ;
      RECT  98.09 103.7 98.27 101.995 ;
      RECT  96.26 103.905 96.47 103.7 ;
      RECT  96.05 104.285 96.26 103.905 ;
      POLYGON  98.66 102.62 98.66 102.21 98.915 102.21 98.915 102.54 98.835 102.62 98.66 102.62 ;
      RECT  96.65 104.615 96.83 103.7 ;
      RECT  96.26 104.615 96.47 104.285 ;
      RECT  96.26 104.285 96.47 103.905 ;
      RECT  98.45 104.58 98.66 104.99 ;
      RECT  96.05 103.575 96.26 103.905 ;
      RECT  99.095 104.49 99.17 106.195 ;
      RECT  99.01 105.075 99.095 105.485 ;
      RECT  98.09 103.575 98.27 104.49 ;
      POLYGON  99.095 103.575 99.095 103.905 98.66 103.905 98.66 104.285 99.095 104.285 99.095 104.49 99.17 104.49 99.17 103.575 99.095 103.575 ;
      RECT  99.17 104.49 99.38 106.195 ;
      POLYGON  98.66 104.58 98.66 104.99 98.835 104.99 98.915 104.91 98.915 104.58 98.66 104.58 ;
      RECT  96.05 104.49 96.26 106.195 ;
      RECT  97.73 103.575 97.91 104.49 ;
      RECT  96.65 104.49 96.83 106.195 ;
      RECT  98.45 105.57 98.66 105.98 ;
      RECT  99.17 104.285 99.38 104.49 ;
      RECT  96.26 104.49 96.47 106.195 ;
      RECT  98.45 103.905 98.66 104.285 ;
      RECT  97.01 104.49 97.19 106.195 ;
      RECT  97.73 104.49 97.91 106.195 ;
      RECT  97.01 103.575 97.19 104.49 ;
      RECT  99.17 103.575 99.38 103.905 ;
      RECT  97.37 104.49 97.55 106.195 ;
      RECT  97.37 103.575 97.55 104.49 ;
      RECT  96.05 104.285 96.26 104.49 ;
      RECT  99.17 103.905 99.38 104.285 ;
      RECT  98.09 104.49 98.27 106.195 ;
      RECT  96.26 104.285 96.47 104.49 ;
      RECT  96.05 103.905 96.26 104.285 ;
      POLYGON  98.66 105.57 98.66 105.98 98.915 105.98 98.915 105.65 98.835 105.57 98.66 105.57 ;
      RECT  96.65 103.575 96.83 104.49 ;
      RECT  96.26 103.575 96.47 103.905 ;
      RECT  96.26 103.905 96.47 104.285 ;
      RECT  98.45 107.56 98.66 107.15 ;
      RECT  96.05 108.565 96.26 108.235 ;
      RECT  99.095 107.65 99.17 105.945 ;
      RECT  99.01 107.065 99.095 106.655 ;
      RECT  98.09 108.565 98.27 107.65 ;
      POLYGON  99.095 108.565 99.095 108.235 98.66 108.235 98.66 107.855 99.095 107.855 99.095 107.65 99.17 107.65 99.17 108.565 99.095 108.565 ;
      RECT  99.17 107.65 99.38 105.945 ;
      POLYGON  98.66 107.56 98.66 107.15 98.835 107.15 98.915 107.23 98.915 107.56 98.66 107.56 ;
      RECT  96.05 107.65 96.26 105.945 ;
      RECT  97.73 108.565 97.91 107.65 ;
      RECT  96.65 107.65 96.83 105.945 ;
      RECT  98.45 106.57 98.66 106.16 ;
      RECT  99.17 107.855 99.38 107.65 ;
      RECT  96.26 107.65 96.47 105.945 ;
      RECT  98.45 108.235 98.66 107.855 ;
      RECT  97.01 107.65 97.19 105.945 ;
      RECT  97.73 107.65 97.91 105.945 ;
      RECT  97.01 108.565 97.19 107.65 ;
      RECT  99.17 108.565 99.38 108.235 ;
      RECT  97.37 107.65 97.55 105.945 ;
      RECT  97.37 108.565 97.55 107.65 ;
      RECT  96.05 107.855 96.26 107.65 ;
      RECT  99.17 108.235 99.38 107.855 ;
      RECT  98.09 107.65 98.27 105.945 ;
      RECT  96.26 107.855 96.47 107.65 ;
      RECT  96.05 108.235 96.26 107.855 ;
      POLYGON  98.66 106.57 98.66 106.16 98.915 106.16 98.915 106.49 98.835 106.57 98.66 106.57 ;
      RECT  96.65 108.565 96.83 107.65 ;
      RECT  96.26 108.565 96.47 108.235 ;
      RECT  96.26 108.235 96.47 107.855 ;
      RECT  98.45 108.53 98.66 108.94 ;
      RECT  96.05 107.525 96.26 107.855 ;
      RECT  99.095 108.44 99.17 110.145 ;
      RECT  99.01 109.025 99.095 109.435 ;
      RECT  98.09 107.525 98.27 108.44 ;
      POLYGON  99.095 107.525 99.095 107.855 98.66 107.855 98.66 108.235 99.095 108.235 99.095 108.44 99.17 108.44 99.17 107.525 99.095 107.525 ;
      RECT  99.17 108.44 99.38 110.145 ;
      POLYGON  98.66 108.53 98.66 108.94 98.835 108.94 98.915 108.86 98.915 108.53 98.66 108.53 ;
      RECT  96.05 108.44 96.26 110.145 ;
      RECT  97.73 107.525 97.91 108.44 ;
      RECT  96.65 108.44 96.83 110.145 ;
      RECT  98.45 109.52 98.66 109.93 ;
      RECT  99.17 108.235 99.38 108.44 ;
      RECT  96.26 108.44 96.47 110.145 ;
      RECT  98.45 107.855 98.66 108.235 ;
      RECT  97.01 108.44 97.19 110.145 ;
      RECT  97.73 108.44 97.91 110.145 ;
      RECT  97.01 107.525 97.19 108.44 ;
      RECT  99.17 107.525 99.38 107.855 ;
      RECT  97.37 108.44 97.55 110.145 ;
      RECT  97.37 107.525 97.55 108.44 ;
      RECT  96.05 108.235 96.26 108.44 ;
      RECT  99.17 107.855 99.38 108.235 ;
      RECT  98.09 108.44 98.27 110.145 ;
      RECT  96.26 108.235 96.47 108.44 ;
      RECT  96.05 107.855 96.26 108.235 ;
      POLYGON  98.66 109.52 98.66 109.93 98.915 109.93 98.915 109.6 98.835 109.52 98.66 109.52 ;
      RECT  96.65 107.525 96.83 108.44 ;
      RECT  96.26 107.525 96.47 107.855 ;
      RECT  96.26 107.855 96.47 108.235 ;
      RECT  98.45 111.51 98.66 111.1 ;
      RECT  96.05 112.515 96.26 112.185 ;
      RECT  99.095 111.6 99.17 109.895 ;
      RECT  99.01 111.015 99.095 110.605 ;
      RECT  98.09 112.515 98.27 111.6 ;
      POLYGON  99.095 112.515 99.095 112.185 98.66 112.185 98.66 111.805 99.095 111.805 99.095 111.6 99.17 111.6 99.17 112.515 99.095 112.515 ;
      RECT  99.17 111.6 99.38 109.895 ;
      POLYGON  98.66 111.51 98.66 111.1 98.835 111.1 98.915 111.18 98.915 111.51 98.66 111.51 ;
      RECT  96.05 111.6 96.26 109.895 ;
      RECT  97.73 112.515 97.91 111.6 ;
      RECT  96.65 111.6 96.83 109.895 ;
      RECT  98.45 110.52 98.66 110.11 ;
      RECT  99.17 111.805 99.38 111.6 ;
      RECT  96.26 111.6 96.47 109.895 ;
      RECT  98.45 112.185 98.66 111.805 ;
      RECT  97.01 111.6 97.19 109.895 ;
      RECT  97.73 111.6 97.91 109.895 ;
      RECT  97.01 112.515 97.19 111.6 ;
      RECT  99.17 112.515 99.38 112.185 ;
      RECT  97.37 111.6 97.55 109.895 ;
      RECT  97.37 112.515 97.55 111.6 ;
      RECT  96.05 111.805 96.26 111.6 ;
      RECT  99.17 112.185 99.38 111.805 ;
      RECT  98.09 111.6 98.27 109.895 ;
      RECT  96.26 111.805 96.47 111.6 ;
      RECT  96.05 112.185 96.26 111.805 ;
      POLYGON  98.66 110.52 98.66 110.11 98.915 110.11 98.915 110.44 98.835 110.52 98.66 110.52 ;
      RECT  96.65 112.515 96.83 111.6 ;
      RECT  96.26 112.515 96.47 112.185 ;
      RECT  96.26 112.185 96.47 111.805 ;
      RECT  98.45 112.48 98.66 112.89 ;
      RECT  96.05 111.475 96.26 111.805 ;
      RECT  99.095 112.39 99.17 114.095 ;
      RECT  99.01 112.975 99.095 113.385 ;
      RECT  98.09 111.475 98.27 112.39 ;
      POLYGON  99.095 111.475 99.095 111.805 98.66 111.805 98.66 112.185 99.095 112.185 99.095 112.39 99.17 112.39 99.17 111.475 99.095 111.475 ;
      RECT  99.17 112.39 99.38 114.095 ;
      POLYGON  98.66 112.48 98.66 112.89 98.835 112.89 98.915 112.81 98.915 112.48 98.66 112.48 ;
      RECT  96.05 112.39 96.26 114.095 ;
      RECT  97.73 111.475 97.91 112.39 ;
      RECT  96.65 112.39 96.83 114.095 ;
      RECT  98.45 113.47 98.66 113.88 ;
      RECT  99.17 112.185 99.38 112.39 ;
      RECT  96.26 112.39 96.47 114.095 ;
      RECT  98.45 111.805 98.66 112.185 ;
      RECT  97.01 112.39 97.19 114.095 ;
      RECT  97.73 112.39 97.91 114.095 ;
      RECT  97.01 111.475 97.19 112.39 ;
      RECT  99.17 111.475 99.38 111.805 ;
      RECT  97.37 112.39 97.55 114.095 ;
      RECT  97.37 111.475 97.55 112.39 ;
      RECT  96.05 112.185 96.26 112.39 ;
      RECT  99.17 111.805 99.38 112.185 ;
      RECT  98.09 112.39 98.27 114.095 ;
      RECT  96.26 112.185 96.47 112.39 ;
      RECT  96.05 111.805 96.26 112.185 ;
      POLYGON  98.66 113.47 98.66 113.88 98.915 113.88 98.915 113.55 98.835 113.47 98.66 113.47 ;
      RECT  96.65 111.475 96.83 112.39 ;
      RECT  96.26 111.475 96.47 111.805 ;
      RECT  96.26 111.805 96.47 112.185 ;
      RECT  98.45 115.46 98.66 115.05 ;
      RECT  96.05 116.465 96.26 116.135 ;
      RECT  99.095 115.55 99.17 113.845 ;
      RECT  99.01 114.965 99.095 114.555 ;
      RECT  98.09 116.465 98.27 115.55 ;
      POLYGON  99.095 116.465 99.095 116.135 98.66 116.135 98.66 115.755 99.095 115.755 99.095 115.55 99.17 115.55 99.17 116.465 99.095 116.465 ;
      RECT  99.17 115.55 99.38 113.845 ;
      POLYGON  98.66 115.46 98.66 115.05 98.835 115.05 98.915 115.13 98.915 115.46 98.66 115.46 ;
      RECT  96.05 115.55 96.26 113.845 ;
      RECT  97.73 116.465 97.91 115.55 ;
      RECT  96.65 115.55 96.83 113.845 ;
      RECT  98.45 114.47 98.66 114.06 ;
      RECT  99.17 115.755 99.38 115.55 ;
      RECT  96.26 115.55 96.47 113.845 ;
      RECT  98.45 116.135 98.66 115.755 ;
      RECT  97.01 115.55 97.19 113.845 ;
      RECT  97.73 115.55 97.91 113.845 ;
      RECT  97.01 116.465 97.19 115.55 ;
      RECT  99.17 116.465 99.38 116.135 ;
      RECT  97.37 115.55 97.55 113.845 ;
      RECT  97.37 116.465 97.55 115.55 ;
      RECT  96.05 115.755 96.26 115.55 ;
      RECT  99.17 116.135 99.38 115.755 ;
      RECT  98.09 115.55 98.27 113.845 ;
      RECT  96.26 115.755 96.47 115.55 ;
      RECT  96.05 116.135 96.26 115.755 ;
      POLYGON  98.66 114.47 98.66 114.06 98.915 114.06 98.915 114.39 98.835 114.47 98.66 114.47 ;
      RECT  96.65 116.465 96.83 115.55 ;
      RECT  96.26 116.465 96.47 116.135 ;
      RECT  96.26 116.135 96.47 115.755 ;
      RECT  98.45 116.43 98.66 116.84 ;
      RECT  96.05 115.425 96.26 115.755 ;
      RECT  99.095 116.34 99.17 118.045 ;
      RECT  99.01 116.925 99.095 117.335 ;
      RECT  98.09 115.425 98.27 116.34 ;
      POLYGON  99.095 115.425 99.095 115.755 98.66 115.755 98.66 116.135 99.095 116.135 99.095 116.34 99.17 116.34 99.17 115.425 99.095 115.425 ;
      RECT  99.17 116.34 99.38 118.045 ;
      POLYGON  98.66 116.43 98.66 116.84 98.835 116.84 98.915 116.76 98.915 116.43 98.66 116.43 ;
      RECT  96.05 116.34 96.26 118.045 ;
      RECT  97.73 115.425 97.91 116.34 ;
      RECT  96.65 116.34 96.83 118.045 ;
      RECT  98.45 117.42 98.66 117.83 ;
      RECT  99.17 116.135 99.38 116.34 ;
      RECT  96.26 116.34 96.47 118.045 ;
      RECT  98.45 115.755 98.66 116.135 ;
      RECT  97.01 116.34 97.19 118.045 ;
      RECT  97.73 116.34 97.91 118.045 ;
      RECT  97.01 115.425 97.19 116.34 ;
      RECT  99.17 115.425 99.38 115.755 ;
      RECT  97.37 116.34 97.55 118.045 ;
      RECT  97.37 115.425 97.55 116.34 ;
      RECT  96.05 116.135 96.26 116.34 ;
      RECT  99.17 115.755 99.38 116.135 ;
      RECT  98.09 116.34 98.27 118.045 ;
      RECT  96.26 116.135 96.47 116.34 ;
      RECT  96.05 115.755 96.26 116.135 ;
      POLYGON  98.66 117.42 98.66 117.83 98.915 117.83 98.915 117.5 98.835 117.42 98.66 117.42 ;
      RECT  96.65 115.425 96.83 116.34 ;
      RECT  96.26 115.425 96.47 115.755 ;
      RECT  96.26 115.755 96.47 116.135 ;
      RECT  98.45 119.41 98.66 119.0 ;
      RECT  96.05 120.415 96.26 120.085 ;
      RECT  99.095 119.5 99.17 117.795 ;
      RECT  99.01 118.915 99.095 118.505 ;
      RECT  98.09 120.415 98.27 119.5 ;
      POLYGON  99.095 120.415 99.095 120.085 98.66 120.085 98.66 119.705 99.095 119.705 99.095 119.5 99.17 119.5 99.17 120.415 99.095 120.415 ;
      RECT  99.17 119.5 99.38 117.795 ;
      POLYGON  98.66 119.41 98.66 119.0 98.835 119.0 98.915 119.08 98.915 119.41 98.66 119.41 ;
      RECT  96.05 119.5 96.26 117.795 ;
      RECT  97.73 120.415 97.91 119.5 ;
      RECT  96.65 119.5 96.83 117.795 ;
      RECT  98.45 118.42 98.66 118.01 ;
      RECT  99.17 119.705 99.38 119.5 ;
      RECT  96.26 119.5 96.47 117.795 ;
      RECT  98.45 120.085 98.66 119.705 ;
      RECT  97.01 119.5 97.19 117.795 ;
      RECT  97.73 119.5 97.91 117.795 ;
      RECT  97.01 120.415 97.19 119.5 ;
      RECT  99.17 120.415 99.38 120.085 ;
      RECT  97.37 119.5 97.55 117.795 ;
      RECT  97.37 120.415 97.55 119.5 ;
      RECT  96.05 119.705 96.26 119.5 ;
      RECT  99.17 120.085 99.38 119.705 ;
      RECT  98.09 119.5 98.27 117.795 ;
      RECT  96.26 119.705 96.47 119.5 ;
      RECT  96.05 120.085 96.26 119.705 ;
      POLYGON  98.66 118.42 98.66 118.01 98.915 118.01 98.915 118.34 98.835 118.42 98.66 118.42 ;
      RECT  96.65 120.415 96.83 119.5 ;
      RECT  96.26 120.415 96.47 120.085 ;
      RECT  96.26 120.085 96.47 119.705 ;
      RECT  98.45 120.38 98.66 120.79 ;
      RECT  96.05 119.375 96.26 119.705 ;
      RECT  99.095 120.29 99.17 121.995 ;
      RECT  99.01 120.875 99.095 121.285 ;
      RECT  98.09 119.375 98.27 120.29 ;
      POLYGON  99.095 119.375 99.095 119.705 98.66 119.705 98.66 120.085 99.095 120.085 99.095 120.29 99.17 120.29 99.17 119.375 99.095 119.375 ;
      RECT  99.17 120.29 99.38 121.995 ;
      POLYGON  98.66 120.38 98.66 120.79 98.835 120.79 98.915 120.71 98.915 120.38 98.66 120.38 ;
      RECT  96.05 120.29 96.26 121.995 ;
      RECT  97.73 119.375 97.91 120.29 ;
      RECT  96.65 120.29 96.83 121.995 ;
      RECT  98.45 121.37 98.66 121.78 ;
      RECT  99.17 120.085 99.38 120.29 ;
      RECT  96.26 120.29 96.47 121.995 ;
      RECT  98.45 119.705 98.66 120.085 ;
      RECT  97.01 120.29 97.19 121.995 ;
      RECT  97.73 120.29 97.91 121.995 ;
      RECT  97.01 119.375 97.19 120.29 ;
      RECT  99.17 119.375 99.38 119.705 ;
      RECT  97.37 120.29 97.55 121.995 ;
      RECT  97.37 119.375 97.55 120.29 ;
      RECT  96.05 120.085 96.26 120.29 ;
      RECT  99.17 119.705 99.38 120.085 ;
      RECT  98.09 120.29 98.27 121.995 ;
      RECT  96.26 120.085 96.47 120.29 ;
      RECT  96.05 119.705 96.26 120.085 ;
      POLYGON  98.66 121.37 98.66 121.78 98.915 121.78 98.915 121.45 98.835 121.37 98.66 121.37 ;
      RECT  96.65 119.375 96.83 120.29 ;
      RECT  96.26 119.375 96.47 119.705 ;
      RECT  96.26 119.705 96.47 120.085 ;
      RECT  98.45 123.36 98.66 122.95 ;
      RECT  96.05 124.365 96.26 124.035 ;
      RECT  99.095 123.45 99.17 121.745 ;
      RECT  99.01 122.865 99.095 122.455 ;
      RECT  98.09 124.365 98.27 123.45 ;
      POLYGON  99.095 124.365 99.095 124.035 98.66 124.035 98.66 123.655 99.095 123.655 99.095 123.45 99.17 123.45 99.17 124.365 99.095 124.365 ;
      RECT  99.17 123.45 99.38 121.745 ;
      POLYGON  98.66 123.36 98.66 122.95 98.835 122.95 98.915 123.03 98.915 123.36 98.66 123.36 ;
      RECT  96.05 123.45 96.26 121.745 ;
      RECT  97.73 124.365 97.91 123.45 ;
      RECT  96.65 123.45 96.83 121.745 ;
      RECT  98.45 122.37 98.66 121.96 ;
      RECT  99.17 123.655 99.38 123.45 ;
      RECT  96.26 123.45 96.47 121.745 ;
      RECT  98.45 124.035 98.66 123.655 ;
      RECT  97.01 123.45 97.19 121.745 ;
      RECT  97.73 123.45 97.91 121.745 ;
      RECT  97.01 124.365 97.19 123.45 ;
      RECT  99.17 124.365 99.38 124.035 ;
      RECT  97.37 123.45 97.55 121.745 ;
      RECT  97.37 124.365 97.55 123.45 ;
      RECT  96.05 123.655 96.26 123.45 ;
      RECT  99.17 124.035 99.38 123.655 ;
      RECT  98.09 123.45 98.27 121.745 ;
      RECT  96.26 123.655 96.47 123.45 ;
      RECT  96.05 124.035 96.26 123.655 ;
      POLYGON  98.66 122.37 98.66 121.96 98.915 121.96 98.915 122.29 98.835 122.37 98.66 122.37 ;
      RECT  96.65 124.365 96.83 123.45 ;
      RECT  96.26 124.365 96.47 124.035 ;
      RECT  96.26 124.035 96.47 123.655 ;
      RECT  100.31 92.73 100.1 93.14 ;
      RECT  102.71 91.725 102.5 92.055 ;
      RECT  99.665 92.64 99.59 94.345 ;
      RECT  99.75 93.225 99.665 93.635 ;
      RECT  100.67 91.725 100.49 92.64 ;
      POLYGON  99.665 91.725 99.665 92.055 100.1 92.055 100.1 92.435 99.665 92.435 99.665 92.64 99.59 92.64 99.59 91.725 99.665 91.725 ;
      RECT  99.59 92.64 99.38 94.345 ;
      POLYGON  100.1 92.73 100.1 93.14 99.925 93.14 99.845 93.06 99.845 92.73 100.1 92.73 ;
      RECT  102.71 92.64 102.5 94.345 ;
      RECT  101.03 91.725 100.85 92.64 ;
      RECT  102.11 92.64 101.93 94.345 ;
      RECT  100.31 93.72 100.1 94.13 ;
      RECT  99.59 92.435 99.38 92.64 ;
      RECT  102.5 92.64 102.29 94.345 ;
      RECT  100.31 92.055 100.1 92.435 ;
      RECT  101.75 92.64 101.57 94.345 ;
      RECT  101.03 92.64 100.85 94.345 ;
      RECT  101.75 91.725 101.57 92.64 ;
      RECT  99.59 91.725 99.38 92.055 ;
      RECT  101.39 92.64 101.21 94.345 ;
      RECT  101.39 91.725 101.21 92.64 ;
      RECT  102.71 92.435 102.5 92.64 ;
      RECT  99.59 92.055 99.38 92.435 ;
      RECT  100.67 92.64 100.49 94.345 ;
      RECT  102.5 92.435 102.29 92.64 ;
      RECT  102.71 92.055 102.5 92.435 ;
      POLYGON  100.1 93.72 100.1 94.13 99.845 94.13 99.845 93.8 99.925 93.72 100.1 93.72 ;
      RECT  102.11 91.725 101.93 92.64 ;
      RECT  102.5 91.725 102.29 92.055 ;
      RECT  102.5 92.055 102.29 92.435 ;
      RECT  100.31 95.71 100.1 95.3 ;
      RECT  102.71 96.715 102.5 96.385 ;
      RECT  99.665 95.8 99.59 94.095 ;
      RECT  99.75 95.215 99.665 94.805 ;
      RECT  100.67 96.715 100.49 95.8 ;
      POLYGON  99.665 96.715 99.665 96.385 100.1 96.385 100.1 96.005 99.665 96.005 99.665 95.8 99.59 95.8 99.59 96.715 99.665 96.715 ;
      RECT  99.59 95.8 99.38 94.095 ;
      POLYGON  100.1 95.71 100.1 95.3 99.925 95.3 99.845 95.38 99.845 95.71 100.1 95.71 ;
      RECT  102.71 95.8 102.5 94.095 ;
      RECT  101.03 96.715 100.85 95.8 ;
      RECT  102.11 95.8 101.93 94.095 ;
      RECT  100.31 94.72 100.1 94.31 ;
      RECT  99.59 96.005 99.38 95.8 ;
      RECT  102.5 95.8 102.29 94.095 ;
      RECT  100.31 96.385 100.1 96.005 ;
      RECT  101.75 95.8 101.57 94.095 ;
      RECT  101.03 95.8 100.85 94.095 ;
      RECT  101.75 96.715 101.57 95.8 ;
      RECT  99.59 96.715 99.38 96.385 ;
      RECT  101.39 95.8 101.21 94.095 ;
      RECT  101.39 96.715 101.21 95.8 ;
      RECT  102.71 96.005 102.5 95.8 ;
      RECT  99.59 96.385 99.38 96.005 ;
      RECT  100.67 95.8 100.49 94.095 ;
      RECT  102.5 96.005 102.29 95.8 ;
      RECT  102.71 96.385 102.5 96.005 ;
      POLYGON  100.1 94.72 100.1 94.31 99.845 94.31 99.845 94.64 99.925 94.72 100.1 94.72 ;
      RECT  102.11 96.715 101.93 95.8 ;
      RECT  102.5 96.715 102.29 96.385 ;
      RECT  102.5 96.385 102.29 96.005 ;
      RECT  100.31 96.68 100.1 97.09 ;
      RECT  102.71 95.675 102.5 96.005 ;
      RECT  99.665 96.59 99.59 98.295 ;
      RECT  99.75 97.175 99.665 97.585 ;
      RECT  100.67 95.675 100.49 96.59 ;
      POLYGON  99.665 95.675 99.665 96.005 100.1 96.005 100.1 96.385 99.665 96.385 99.665 96.59 99.59 96.59 99.59 95.675 99.665 95.675 ;
      RECT  99.59 96.59 99.38 98.295 ;
      POLYGON  100.1 96.68 100.1 97.09 99.925 97.09 99.845 97.01 99.845 96.68 100.1 96.68 ;
      RECT  102.71 96.59 102.5 98.295 ;
      RECT  101.03 95.675 100.85 96.59 ;
      RECT  102.11 96.59 101.93 98.295 ;
      RECT  100.31 97.67 100.1 98.08 ;
      RECT  99.59 96.385 99.38 96.59 ;
      RECT  102.5 96.59 102.29 98.295 ;
      RECT  100.31 96.005 100.1 96.385 ;
      RECT  101.75 96.59 101.57 98.295 ;
      RECT  101.03 96.59 100.85 98.295 ;
      RECT  101.75 95.675 101.57 96.59 ;
      RECT  99.59 95.675 99.38 96.005 ;
      RECT  101.39 96.59 101.21 98.295 ;
      RECT  101.39 95.675 101.21 96.59 ;
      RECT  102.71 96.385 102.5 96.59 ;
      RECT  99.59 96.005 99.38 96.385 ;
      RECT  100.67 96.59 100.49 98.295 ;
      RECT  102.5 96.385 102.29 96.59 ;
      RECT  102.71 96.005 102.5 96.385 ;
      POLYGON  100.1 97.67 100.1 98.08 99.845 98.08 99.845 97.75 99.925 97.67 100.1 97.67 ;
      RECT  102.11 95.675 101.93 96.59 ;
      RECT  102.5 95.675 102.29 96.005 ;
      RECT  102.5 96.005 102.29 96.385 ;
      RECT  100.31 99.66 100.1 99.25 ;
      RECT  102.71 100.665 102.5 100.335 ;
      RECT  99.665 99.75 99.59 98.045 ;
      RECT  99.75 99.165 99.665 98.755 ;
      RECT  100.67 100.665 100.49 99.75 ;
      POLYGON  99.665 100.665 99.665 100.335 100.1 100.335 100.1 99.955 99.665 99.955 99.665 99.75 99.59 99.75 99.59 100.665 99.665 100.665 ;
      RECT  99.59 99.75 99.38 98.045 ;
      POLYGON  100.1 99.66 100.1 99.25 99.925 99.25 99.845 99.33 99.845 99.66 100.1 99.66 ;
      RECT  102.71 99.75 102.5 98.045 ;
      RECT  101.03 100.665 100.85 99.75 ;
      RECT  102.11 99.75 101.93 98.045 ;
      RECT  100.31 98.67 100.1 98.26 ;
      RECT  99.59 99.955 99.38 99.75 ;
      RECT  102.5 99.75 102.29 98.045 ;
      RECT  100.31 100.335 100.1 99.955 ;
      RECT  101.75 99.75 101.57 98.045 ;
      RECT  101.03 99.75 100.85 98.045 ;
      RECT  101.75 100.665 101.57 99.75 ;
      RECT  99.59 100.665 99.38 100.335 ;
      RECT  101.39 99.75 101.21 98.045 ;
      RECT  101.39 100.665 101.21 99.75 ;
      RECT  102.71 99.955 102.5 99.75 ;
      RECT  99.59 100.335 99.38 99.955 ;
      RECT  100.67 99.75 100.49 98.045 ;
      RECT  102.5 99.955 102.29 99.75 ;
      RECT  102.71 100.335 102.5 99.955 ;
      POLYGON  100.1 98.67 100.1 98.26 99.845 98.26 99.845 98.59 99.925 98.67 100.1 98.67 ;
      RECT  102.11 100.665 101.93 99.75 ;
      RECT  102.5 100.665 102.29 100.335 ;
      RECT  102.5 100.335 102.29 99.955 ;
      RECT  100.31 100.63 100.1 101.04 ;
      RECT  102.71 99.625 102.5 99.955 ;
      RECT  99.665 100.54 99.59 102.245 ;
      RECT  99.75 101.125 99.665 101.535 ;
      RECT  100.67 99.625 100.49 100.54 ;
      POLYGON  99.665 99.625 99.665 99.955 100.1 99.955 100.1 100.335 99.665 100.335 99.665 100.54 99.59 100.54 99.59 99.625 99.665 99.625 ;
      RECT  99.59 100.54 99.38 102.245 ;
      POLYGON  100.1 100.63 100.1 101.04 99.925 101.04 99.845 100.96 99.845 100.63 100.1 100.63 ;
      RECT  102.71 100.54 102.5 102.245 ;
      RECT  101.03 99.625 100.85 100.54 ;
      RECT  102.11 100.54 101.93 102.245 ;
      RECT  100.31 101.62 100.1 102.03 ;
      RECT  99.59 100.335 99.38 100.54 ;
      RECT  102.5 100.54 102.29 102.245 ;
      RECT  100.31 99.955 100.1 100.335 ;
      RECT  101.75 100.54 101.57 102.245 ;
      RECT  101.03 100.54 100.85 102.245 ;
      RECT  101.75 99.625 101.57 100.54 ;
      RECT  99.59 99.625 99.38 99.955 ;
      RECT  101.39 100.54 101.21 102.245 ;
      RECT  101.39 99.625 101.21 100.54 ;
      RECT  102.71 100.335 102.5 100.54 ;
      RECT  99.59 99.955 99.38 100.335 ;
      RECT  100.67 100.54 100.49 102.245 ;
      RECT  102.5 100.335 102.29 100.54 ;
      RECT  102.71 99.955 102.5 100.335 ;
      POLYGON  100.1 101.62 100.1 102.03 99.845 102.03 99.845 101.7 99.925 101.62 100.1 101.62 ;
      RECT  102.11 99.625 101.93 100.54 ;
      RECT  102.5 99.625 102.29 99.955 ;
      RECT  102.5 99.955 102.29 100.335 ;
      RECT  100.31 103.61 100.1 103.2 ;
      RECT  102.71 104.615 102.5 104.285 ;
      RECT  99.665 103.7 99.59 101.995 ;
      RECT  99.75 103.115 99.665 102.705 ;
      RECT  100.67 104.615 100.49 103.7 ;
      POLYGON  99.665 104.615 99.665 104.285 100.1 104.285 100.1 103.905 99.665 103.905 99.665 103.7 99.59 103.7 99.59 104.615 99.665 104.615 ;
      RECT  99.59 103.7 99.38 101.995 ;
      POLYGON  100.1 103.61 100.1 103.2 99.925 103.2 99.845 103.28 99.845 103.61 100.1 103.61 ;
      RECT  102.71 103.7 102.5 101.995 ;
      RECT  101.03 104.615 100.85 103.7 ;
      RECT  102.11 103.7 101.93 101.995 ;
      RECT  100.31 102.62 100.1 102.21 ;
      RECT  99.59 103.905 99.38 103.7 ;
      RECT  102.5 103.7 102.29 101.995 ;
      RECT  100.31 104.285 100.1 103.905 ;
      RECT  101.75 103.7 101.57 101.995 ;
      RECT  101.03 103.7 100.85 101.995 ;
      RECT  101.75 104.615 101.57 103.7 ;
      RECT  99.59 104.615 99.38 104.285 ;
      RECT  101.39 103.7 101.21 101.995 ;
      RECT  101.39 104.615 101.21 103.7 ;
      RECT  102.71 103.905 102.5 103.7 ;
      RECT  99.59 104.285 99.38 103.905 ;
      RECT  100.67 103.7 100.49 101.995 ;
      RECT  102.5 103.905 102.29 103.7 ;
      RECT  102.71 104.285 102.5 103.905 ;
      POLYGON  100.1 102.62 100.1 102.21 99.845 102.21 99.845 102.54 99.925 102.62 100.1 102.62 ;
      RECT  102.11 104.615 101.93 103.7 ;
      RECT  102.5 104.615 102.29 104.285 ;
      RECT  102.5 104.285 102.29 103.905 ;
      RECT  100.31 104.58 100.1 104.99 ;
      RECT  102.71 103.575 102.5 103.905 ;
      RECT  99.665 104.49 99.59 106.195 ;
      RECT  99.75 105.075 99.665 105.485 ;
      RECT  100.67 103.575 100.49 104.49 ;
      POLYGON  99.665 103.575 99.665 103.905 100.1 103.905 100.1 104.285 99.665 104.285 99.665 104.49 99.59 104.49 99.59 103.575 99.665 103.575 ;
      RECT  99.59 104.49 99.38 106.195 ;
      POLYGON  100.1 104.58 100.1 104.99 99.925 104.99 99.845 104.91 99.845 104.58 100.1 104.58 ;
      RECT  102.71 104.49 102.5 106.195 ;
      RECT  101.03 103.575 100.85 104.49 ;
      RECT  102.11 104.49 101.93 106.195 ;
      RECT  100.31 105.57 100.1 105.98 ;
      RECT  99.59 104.285 99.38 104.49 ;
      RECT  102.5 104.49 102.29 106.195 ;
      RECT  100.31 103.905 100.1 104.285 ;
      RECT  101.75 104.49 101.57 106.195 ;
      RECT  101.03 104.49 100.85 106.195 ;
      RECT  101.75 103.575 101.57 104.49 ;
      RECT  99.59 103.575 99.38 103.905 ;
      RECT  101.39 104.49 101.21 106.195 ;
      RECT  101.39 103.575 101.21 104.49 ;
      RECT  102.71 104.285 102.5 104.49 ;
      RECT  99.59 103.905 99.38 104.285 ;
      RECT  100.67 104.49 100.49 106.195 ;
      RECT  102.5 104.285 102.29 104.49 ;
      RECT  102.71 103.905 102.5 104.285 ;
      POLYGON  100.1 105.57 100.1 105.98 99.845 105.98 99.845 105.65 99.925 105.57 100.1 105.57 ;
      RECT  102.11 103.575 101.93 104.49 ;
      RECT  102.5 103.575 102.29 103.905 ;
      RECT  102.5 103.905 102.29 104.285 ;
      RECT  100.31 107.56 100.1 107.15 ;
      RECT  102.71 108.565 102.5 108.235 ;
      RECT  99.665 107.65 99.59 105.945 ;
      RECT  99.75 107.065 99.665 106.655 ;
      RECT  100.67 108.565 100.49 107.65 ;
      POLYGON  99.665 108.565 99.665 108.235 100.1 108.235 100.1 107.855 99.665 107.855 99.665 107.65 99.59 107.65 99.59 108.565 99.665 108.565 ;
      RECT  99.59 107.65 99.38 105.945 ;
      POLYGON  100.1 107.56 100.1 107.15 99.925 107.15 99.845 107.23 99.845 107.56 100.1 107.56 ;
      RECT  102.71 107.65 102.5 105.945 ;
      RECT  101.03 108.565 100.85 107.65 ;
      RECT  102.11 107.65 101.93 105.945 ;
      RECT  100.31 106.57 100.1 106.16 ;
      RECT  99.59 107.855 99.38 107.65 ;
      RECT  102.5 107.65 102.29 105.945 ;
      RECT  100.31 108.235 100.1 107.855 ;
      RECT  101.75 107.65 101.57 105.945 ;
      RECT  101.03 107.65 100.85 105.945 ;
      RECT  101.75 108.565 101.57 107.65 ;
      RECT  99.59 108.565 99.38 108.235 ;
      RECT  101.39 107.65 101.21 105.945 ;
      RECT  101.39 108.565 101.21 107.65 ;
      RECT  102.71 107.855 102.5 107.65 ;
      RECT  99.59 108.235 99.38 107.855 ;
      RECT  100.67 107.65 100.49 105.945 ;
      RECT  102.5 107.855 102.29 107.65 ;
      RECT  102.71 108.235 102.5 107.855 ;
      POLYGON  100.1 106.57 100.1 106.16 99.845 106.16 99.845 106.49 99.925 106.57 100.1 106.57 ;
      RECT  102.11 108.565 101.93 107.65 ;
      RECT  102.5 108.565 102.29 108.235 ;
      RECT  102.5 108.235 102.29 107.855 ;
      RECT  100.31 108.53 100.1 108.94 ;
      RECT  102.71 107.525 102.5 107.855 ;
      RECT  99.665 108.44 99.59 110.145 ;
      RECT  99.75 109.025 99.665 109.435 ;
      RECT  100.67 107.525 100.49 108.44 ;
      POLYGON  99.665 107.525 99.665 107.855 100.1 107.855 100.1 108.235 99.665 108.235 99.665 108.44 99.59 108.44 99.59 107.525 99.665 107.525 ;
      RECT  99.59 108.44 99.38 110.145 ;
      POLYGON  100.1 108.53 100.1 108.94 99.925 108.94 99.845 108.86 99.845 108.53 100.1 108.53 ;
      RECT  102.71 108.44 102.5 110.145 ;
      RECT  101.03 107.525 100.85 108.44 ;
      RECT  102.11 108.44 101.93 110.145 ;
      RECT  100.31 109.52 100.1 109.93 ;
      RECT  99.59 108.235 99.38 108.44 ;
      RECT  102.5 108.44 102.29 110.145 ;
      RECT  100.31 107.855 100.1 108.235 ;
      RECT  101.75 108.44 101.57 110.145 ;
      RECT  101.03 108.44 100.85 110.145 ;
      RECT  101.75 107.525 101.57 108.44 ;
      RECT  99.59 107.525 99.38 107.855 ;
      RECT  101.39 108.44 101.21 110.145 ;
      RECT  101.39 107.525 101.21 108.44 ;
      RECT  102.71 108.235 102.5 108.44 ;
      RECT  99.59 107.855 99.38 108.235 ;
      RECT  100.67 108.44 100.49 110.145 ;
      RECT  102.5 108.235 102.29 108.44 ;
      RECT  102.71 107.855 102.5 108.235 ;
      POLYGON  100.1 109.52 100.1 109.93 99.845 109.93 99.845 109.6 99.925 109.52 100.1 109.52 ;
      RECT  102.11 107.525 101.93 108.44 ;
      RECT  102.5 107.525 102.29 107.855 ;
      RECT  102.5 107.855 102.29 108.235 ;
      RECT  100.31 111.51 100.1 111.1 ;
      RECT  102.71 112.515 102.5 112.185 ;
      RECT  99.665 111.6 99.59 109.895 ;
      RECT  99.75 111.015 99.665 110.605 ;
      RECT  100.67 112.515 100.49 111.6 ;
      POLYGON  99.665 112.515 99.665 112.185 100.1 112.185 100.1 111.805 99.665 111.805 99.665 111.6 99.59 111.6 99.59 112.515 99.665 112.515 ;
      RECT  99.59 111.6 99.38 109.895 ;
      POLYGON  100.1 111.51 100.1 111.1 99.925 111.1 99.845 111.18 99.845 111.51 100.1 111.51 ;
      RECT  102.71 111.6 102.5 109.895 ;
      RECT  101.03 112.515 100.85 111.6 ;
      RECT  102.11 111.6 101.93 109.895 ;
      RECT  100.31 110.52 100.1 110.11 ;
      RECT  99.59 111.805 99.38 111.6 ;
      RECT  102.5 111.6 102.29 109.895 ;
      RECT  100.31 112.185 100.1 111.805 ;
      RECT  101.75 111.6 101.57 109.895 ;
      RECT  101.03 111.6 100.85 109.895 ;
      RECT  101.75 112.515 101.57 111.6 ;
      RECT  99.59 112.515 99.38 112.185 ;
      RECT  101.39 111.6 101.21 109.895 ;
      RECT  101.39 112.515 101.21 111.6 ;
      RECT  102.71 111.805 102.5 111.6 ;
      RECT  99.59 112.185 99.38 111.805 ;
      RECT  100.67 111.6 100.49 109.895 ;
      RECT  102.5 111.805 102.29 111.6 ;
      RECT  102.71 112.185 102.5 111.805 ;
      POLYGON  100.1 110.52 100.1 110.11 99.845 110.11 99.845 110.44 99.925 110.52 100.1 110.52 ;
      RECT  102.11 112.515 101.93 111.6 ;
      RECT  102.5 112.515 102.29 112.185 ;
      RECT  102.5 112.185 102.29 111.805 ;
      RECT  100.31 112.48 100.1 112.89 ;
      RECT  102.71 111.475 102.5 111.805 ;
      RECT  99.665 112.39 99.59 114.095 ;
      RECT  99.75 112.975 99.665 113.385 ;
      RECT  100.67 111.475 100.49 112.39 ;
      POLYGON  99.665 111.475 99.665 111.805 100.1 111.805 100.1 112.185 99.665 112.185 99.665 112.39 99.59 112.39 99.59 111.475 99.665 111.475 ;
      RECT  99.59 112.39 99.38 114.095 ;
      POLYGON  100.1 112.48 100.1 112.89 99.925 112.89 99.845 112.81 99.845 112.48 100.1 112.48 ;
      RECT  102.71 112.39 102.5 114.095 ;
      RECT  101.03 111.475 100.85 112.39 ;
      RECT  102.11 112.39 101.93 114.095 ;
      RECT  100.31 113.47 100.1 113.88 ;
      RECT  99.59 112.185 99.38 112.39 ;
      RECT  102.5 112.39 102.29 114.095 ;
      RECT  100.31 111.805 100.1 112.185 ;
      RECT  101.75 112.39 101.57 114.095 ;
      RECT  101.03 112.39 100.85 114.095 ;
      RECT  101.75 111.475 101.57 112.39 ;
      RECT  99.59 111.475 99.38 111.805 ;
      RECT  101.39 112.39 101.21 114.095 ;
      RECT  101.39 111.475 101.21 112.39 ;
      RECT  102.71 112.185 102.5 112.39 ;
      RECT  99.59 111.805 99.38 112.185 ;
      RECT  100.67 112.39 100.49 114.095 ;
      RECT  102.5 112.185 102.29 112.39 ;
      RECT  102.71 111.805 102.5 112.185 ;
      POLYGON  100.1 113.47 100.1 113.88 99.845 113.88 99.845 113.55 99.925 113.47 100.1 113.47 ;
      RECT  102.11 111.475 101.93 112.39 ;
      RECT  102.5 111.475 102.29 111.805 ;
      RECT  102.5 111.805 102.29 112.185 ;
      RECT  100.31 115.46 100.1 115.05 ;
      RECT  102.71 116.465 102.5 116.135 ;
      RECT  99.665 115.55 99.59 113.845 ;
      RECT  99.75 114.965 99.665 114.555 ;
      RECT  100.67 116.465 100.49 115.55 ;
      POLYGON  99.665 116.465 99.665 116.135 100.1 116.135 100.1 115.755 99.665 115.755 99.665 115.55 99.59 115.55 99.59 116.465 99.665 116.465 ;
      RECT  99.59 115.55 99.38 113.845 ;
      POLYGON  100.1 115.46 100.1 115.05 99.925 115.05 99.845 115.13 99.845 115.46 100.1 115.46 ;
      RECT  102.71 115.55 102.5 113.845 ;
      RECT  101.03 116.465 100.85 115.55 ;
      RECT  102.11 115.55 101.93 113.845 ;
      RECT  100.31 114.47 100.1 114.06 ;
      RECT  99.59 115.755 99.38 115.55 ;
      RECT  102.5 115.55 102.29 113.845 ;
      RECT  100.31 116.135 100.1 115.755 ;
      RECT  101.75 115.55 101.57 113.845 ;
      RECT  101.03 115.55 100.85 113.845 ;
      RECT  101.75 116.465 101.57 115.55 ;
      RECT  99.59 116.465 99.38 116.135 ;
      RECT  101.39 115.55 101.21 113.845 ;
      RECT  101.39 116.465 101.21 115.55 ;
      RECT  102.71 115.755 102.5 115.55 ;
      RECT  99.59 116.135 99.38 115.755 ;
      RECT  100.67 115.55 100.49 113.845 ;
      RECT  102.5 115.755 102.29 115.55 ;
      RECT  102.71 116.135 102.5 115.755 ;
      POLYGON  100.1 114.47 100.1 114.06 99.845 114.06 99.845 114.39 99.925 114.47 100.1 114.47 ;
      RECT  102.11 116.465 101.93 115.55 ;
      RECT  102.5 116.465 102.29 116.135 ;
      RECT  102.5 116.135 102.29 115.755 ;
      RECT  100.31 116.43 100.1 116.84 ;
      RECT  102.71 115.425 102.5 115.755 ;
      RECT  99.665 116.34 99.59 118.045 ;
      RECT  99.75 116.925 99.665 117.335 ;
      RECT  100.67 115.425 100.49 116.34 ;
      POLYGON  99.665 115.425 99.665 115.755 100.1 115.755 100.1 116.135 99.665 116.135 99.665 116.34 99.59 116.34 99.59 115.425 99.665 115.425 ;
      RECT  99.59 116.34 99.38 118.045 ;
      POLYGON  100.1 116.43 100.1 116.84 99.925 116.84 99.845 116.76 99.845 116.43 100.1 116.43 ;
      RECT  102.71 116.34 102.5 118.045 ;
      RECT  101.03 115.425 100.85 116.34 ;
      RECT  102.11 116.34 101.93 118.045 ;
      RECT  100.31 117.42 100.1 117.83 ;
      RECT  99.59 116.135 99.38 116.34 ;
      RECT  102.5 116.34 102.29 118.045 ;
      RECT  100.31 115.755 100.1 116.135 ;
      RECT  101.75 116.34 101.57 118.045 ;
      RECT  101.03 116.34 100.85 118.045 ;
      RECT  101.75 115.425 101.57 116.34 ;
      RECT  99.59 115.425 99.38 115.755 ;
      RECT  101.39 116.34 101.21 118.045 ;
      RECT  101.39 115.425 101.21 116.34 ;
      RECT  102.71 116.135 102.5 116.34 ;
      RECT  99.59 115.755 99.38 116.135 ;
      RECT  100.67 116.34 100.49 118.045 ;
      RECT  102.5 116.135 102.29 116.34 ;
      RECT  102.71 115.755 102.5 116.135 ;
      POLYGON  100.1 117.42 100.1 117.83 99.845 117.83 99.845 117.5 99.925 117.42 100.1 117.42 ;
      RECT  102.11 115.425 101.93 116.34 ;
      RECT  102.5 115.425 102.29 115.755 ;
      RECT  102.5 115.755 102.29 116.135 ;
      RECT  100.31 119.41 100.1 119.0 ;
      RECT  102.71 120.415 102.5 120.085 ;
      RECT  99.665 119.5 99.59 117.795 ;
      RECT  99.75 118.915 99.665 118.505 ;
      RECT  100.67 120.415 100.49 119.5 ;
      POLYGON  99.665 120.415 99.665 120.085 100.1 120.085 100.1 119.705 99.665 119.705 99.665 119.5 99.59 119.5 99.59 120.415 99.665 120.415 ;
      RECT  99.59 119.5 99.38 117.795 ;
      POLYGON  100.1 119.41 100.1 119.0 99.925 119.0 99.845 119.08 99.845 119.41 100.1 119.41 ;
      RECT  102.71 119.5 102.5 117.795 ;
      RECT  101.03 120.415 100.85 119.5 ;
      RECT  102.11 119.5 101.93 117.795 ;
      RECT  100.31 118.42 100.1 118.01 ;
      RECT  99.59 119.705 99.38 119.5 ;
      RECT  102.5 119.5 102.29 117.795 ;
      RECT  100.31 120.085 100.1 119.705 ;
      RECT  101.75 119.5 101.57 117.795 ;
      RECT  101.03 119.5 100.85 117.795 ;
      RECT  101.75 120.415 101.57 119.5 ;
      RECT  99.59 120.415 99.38 120.085 ;
      RECT  101.39 119.5 101.21 117.795 ;
      RECT  101.39 120.415 101.21 119.5 ;
      RECT  102.71 119.705 102.5 119.5 ;
      RECT  99.59 120.085 99.38 119.705 ;
      RECT  100.67 119.5 100.49 117.795 ;
      RECT  102.5 119.705 102.29 119.5 ;
      RECT  102.71 120.085 102.5 119.705 ;
      POLYGON  100.1 118.42 100.1 118.01 99.845 118.01 99.845 118.34 99.925 118.42 100.1 118.42 ;
      RECT  102.11 120.415 101.93 119.5 ;
      RECT  102.5 120.415 102.29 120.085 ;
      RECT  102.5 120.085 102.29 119.705 ;
      RECT  100.31 120.38 100.1 120.79 ;
      RECT  102.71 119.375 102.5 119.705 ;
      RECT  99.665 120.29 99.59 121.995 ;
      RECT  99.75 120.875 99.665 121.285 ;
      RECT  100.67 119.375 100.49 120.29 ;
      POLYGON  99.665 119.375 99.665 119.705 100.1 119.705 100.1 120.085 99.665 120.085 99.665 120.29 99.59 120.29 99.59 119.375 99.665 119.375 ;
      RECT  99.59 120.29 99.38 121.995 ;
      POLYGON  100.1 120.38 100.1 120.79 99.925 120.79 99.845 120.71 99.845 120.38 100.1 120.38 ;
      RECT  102.71 120.29 102.5 121.995 ;
      RECT  101.03 119.375 100.85 120.29 ;
      RECT  102.11 120.29 101.93 121.995 ;
      RECT  100.31 121.37 100.1 121.78 ;
      RECT  99.59 120.085 99.38 120.29 ;
      RECT  102.5 120.29 102.29 121.995 ;
      RECT  100.31 119.705 100.1 120.085 ;
      RECT  101.75 120.29 101.57 121.995 ;
      RECT  101.03 120.29 100.85 121.995 ;
      RECT  101.75 119.375 101.57 120.29 ;
      RECT  99.59 119.375 99.38 119.705 ;
      RECT  101.39 120.29 101.21 121.995 ;
      RECT  101.39 119.375 101.21 120.29 ;
      RECT  102.71 120.085 102.5 120.29 ;
      RECT  99.59 119.705 99.38 120.085 ;
      RECT  100.67 120.29 100.49 121.995 ;
      RECT  102.5 120.085 102.29 120.29 ;
      RECT  102.71 119.705 102.5 120.085 ;
      POLYGON  100.1 121.37 100.1 121.78 99.845 121.78 99.845 121.45 99.925 121.37 100.1 121.37 ;
      RECT  102.11 119.375 101.93 120.29 ;
      RECT  102.5 119.375 102.29 119.705 ;
      RECT  102.5 119.705 102.29 120.085 ;
      RECT  100.31 123.36 100.1 122.95 ;
      RECT  102.71 124.365 102.5 124.035 ;
      RECT  99.665 123.45 99.59 121.745 ;
      RECT  99.75 122.865 99.665 122.455 ;
      RECT  100.67 124.365 100.49 123.45 ;
      POLYGON  99.665 124.365 99.665 124.035 100.1 124.035 100.1 123.655 99.665 123.655 99.665 123.45 99.59 123.45 99.59 124.365 99.665 124.365 ;
      RECT  99.59 123.45 99.38 121.745 ;
      POLYGON  100.1 123.36 100.1 122.95 99.925 122.95 99.845 123.03 99.845 123.36 100.1 123.36 ;
      RECT  102.71 123.45 102.5 121.745 ;
      RECT  101.03 124.365 100.85 123.45 ;
      RECT  102.11 123.45 101.93 121.745 ;
      RECT  100.31 122.37 100.1 121.96 ;
      RECT  99.59 123.655 99.38 123.45 ;
      RECT  102.5 123.45 102.29 121.745 ;
      RECT  100.31 124.035 100.1 123.655 ;
      RECT  101.75 123.45 101.57 121.745 ;
      RECT  101.03 123.45 100.85 121.745 ;
      RECT  101.75 124.365 101.57 123.45 ;
      RECT  99.59 124.365 99.38 124.035 ;
      RECT  101.39 123.45 101.21 121.745 ;
      RECT  101.39 124.365 101.21 123.45 ;
      RECT  102.71 123.655 102.5 123.45 ;
      RECT  99.59 124.035 99.38 123.655 ;
      RECT  100.67 123.45 100.49 121.745 ;
      RECT  102.5 123.655 102.29 123.45 ;
      RECT  102.71 124.035 102.5 123.655 ;
      POLYGON  100.1 122.37 100.1 121.96 99.845 121.96 99.845 122.29 99.925 122.37 100.1 122.37 ;
      RECT  102.11 124.365 101.93 123.45 ;
      RECT  102.5 124.365 102.29 124.035 ;
      RECT  102.5 124.035 102.29 123.655 ;
      RECT  104.69 92.73 104.9 93.14 ;
      RECT  102.29 91.725 102.5 92.055 ;
      RECT  105.335 92.64 105.41 94.345 ;
      RECT  105.25 93.225 105.335 93.635 ;
      RECT  104.33 91.725 104.51 92.64 ;
      POLYGON  105.335 91.725 105.335 92.055 104.9 92.055 104.9 92.435 105.335 92.435 105.335 92.64 105.41 92.64 105.41 91.725 105.335 91.725 ;
      RECT  105.41 92.64 105.62 94.345 ;
      POLYGON  104.9 92.73 104.9 93.14 105.075 93.14 105.155 93.06 105.155 92.73 104.9 92.73 ;
      RECT  102.29 92.64 102.5 94.345 ;
      RECT  103.97 91.725 104.15 92.64 ;
      RECT  102.89 92.64 103.07 94.345 ;
      RECT  104.69 93.72 104.9 94.13 ;
      RECT  105.41 92.435 105.62 92.64 ;
      RECT  102.5 92.64 102.71 94.345 ;
      RECT  104.69 92.055 104.9 92.435 ;
      RECT  103.25 92.64 103.43 94.345 ;
      RECT  103.97 92.64 104.15 94.345 ;
      RECT  103.25 91.725 103.43 92.64 ;
      RECT  105.41 91.725 105.62 92.055 ;
      RECT  103.61 92.64 103.79 94.345 ;
      RECT  103.61 91.725 103.79 92.64 ;
      RECT  102.29 92.435 102.5 92.64 ;
      RECT  105.41 92.055 105.62 92.435 ;
      RECT  104.33 92.64 104.51 94.345 ;
      RECT  102.5 92.435 102.71 92.64 ;
      RECT  102.29 92.055 102.5 92.435 ;
      POLYGON  104.9 93.72 104.9 94.13 105.155 94.13 105.155 93.8 105.075 93.72 104.9 93.72 ;
      RECT  102.89 91.725 103.07 92.64 ;
      RECT  102.5 91.725 102.71 92.055 ;
      RECT  102.5 92.055 102.71 92.435 ;
      RECT  104.69 95.71 104.9 95.3 ;
      RECT  102.29 96.715 102.5 96.385 ;
      RECT  105.335 95.8 105.41 94.095 ;
      RECT  105.25 95.215 105.335 94.805 ;
      RECT  104.33 96.715 104.51 95.8 ;
      POLYGON  105.335 96.715 105.335 96.385 104.9 96.385 104.9 96.005 105.335 96.005 105.335 95.8 105.41 95.8 105.41 96.715 105.335 96.715 ;
      RECT  105.41 95.8 105.62 94.095 ;
      POLYGON  104.9 95.71 104.9 95.3 105.075 95.3 105.155 95.38 105.155 95.71 104.9 95.71 ;
      RECT  102.29 95.8 102.5 94.095 ;
      RECT  103.97 96.715 104.15 95.8 ;
      RECT  102.89 95.8 103.07 94.095 ;
      RECT  104.69 94.72 104.9 94.31 ;
      RECT  105.41 96.005 105.62 95.8 ;
      RECT  102.5 95.8 102.71 94.095 ;
      RECT  104.69 96.385 104.9 96.005 ;
      RECT  103.25 95.8 103.43 94.095 ;
      RECT  103.97 95.8 104.15 94.095 ;
      RECT  103.25 96.715 103.43 95.8 ;
      RECT  105.41 96.715 105.62 96.385 ;
      RECT  103.61 95.8 103.79 94.095 ;
      RECT  103.61 96.715 103.79 95.8 ;
      RECT  102.29 96.005 102.5 95.8 ;
      RECT  105.41 96.385 105.62 96.005 ;
      RECT  104.33 95.8 104.51 94.095 ;
      RECT  102.5 96.005 102.71 95.8 ;
      RECT  102.29 96.385 102.5 96.005 ;
      POLYGON  104.9 94.72 104.9 94.31 105.155 94.31 105.155 94.64 105.075 94.72 104.9 94.72 ;
      RECT  102.89 96.715 103.07 95.8 ;
      RECT  102.5 96.715 102.71 96.385 ;
      RECT  102.5 96.385 102.71 96.005 ;
      RECT  104.69 96.68 104.9 97.09 ;
      RECT  102.29 95.675 102.5 96.005 ;
      RECT  105.335 96.59 105.41 98.295 ;
      RECT  105.25 97.175 105.335 97.585 ;
      RECT  104.33 95.675 104.51 96.59 ;
      POLYGON  105.335 95.675 105.335 96.005 104.9 96.005 104.9 96.385 105.335 96.385 105.335 96.59 105.41 96.59 105.41 95.675 105.335 95.675 ;
      RECT  105.41 96.59 105.62 98.295 ;
      POLYGON  104.9 96.68 104.9 97.09 105.075 97.09 105.155 97.01 105.155 96.68 104.9 96.68 ;
      RECT  102.29 96.59 102.5 98.295 ;
      RECT  103.97 95.675 104.15 96.59 ;
      RECT  102.89 96.59 103.07 98.295 ;
      RECT  104.69 97.67 104.9 98.08 ;
      RECT  105.41 96.385 105.62 96.59 ;
      RECT  102.5 96.59 102.71 98.295 ;
      RECT  104.69 96.005 104.9 96.385 ;
      RECT  103.25 96.59 103.43 98.295 ;
      RECT  103.97 96.59 104.15 98.295 ;
      RECT  103.25 95.675 103.43 96.59 ;
      RECT  105.41 95.675 105.62 96.005 ;
      RECT  103.61 96.59 103.79 98.295 ;
      RECT  103.61 95.675 103.79 96.59 ;
      RECT  102.29 96.385 102.5 96.59 ;
      RECT  105.41 96.005 105.62 96.385 ;
      RECT  104.33 96.59 104.51 98.295 ;
      RECT  102.5 96.385 102.71 96.59 ;
      RECT  102.29 96.005 102.5 96.385 ;
      POLYGON  104.9 97.67 104.9 98.08 105.155 98.08 105.155 97.75 105.075 97.67 104.9 97.67 ;
      RECT  102.89 95.675 103.07 96.59 ;
      RECT  102.5 95.675 102.71 96.005 ;
      RECT  102.5 96.005 102.71 96.385 ;
      RECT  104.69 99.66 104.9 99.25 ;
      RECT  102.29 100.665 102.5 100.335 ;
      RECT  105.335 99.75 105.41 98.045 ;
      RECT  105.25 99.165 105.335 98.755 ;
      RECT  104.33 100.665 104.51 99.75 ;
      POLYGON  105.335 100.665 105.335 100.335 104.9 100.335 104.9 99.955 105.335 99.955 105.335 99.75 105.41 99.75 105.41 100.665 105.335 100.665 ;
      RECT  105.41 99.75 105.62 98.045 ;
      POLYGON  104.9 99.66 104.9 99.25 105.075 99.25 105.155 99.33 105.155 99.66 104.9 99.66 ;
      RECT  102.29 99.75 102.5 98.045 ;
      RECT  103.97 100.665 104.15 99.75 ;
      RECT  102.89 99.75 103.07 98.045 ;
      RECT  104.69 98.67 104.9 98.26 ;
      RECT  105.41 99.955 105.62 99.75 ;
      RECT  102.5 99.75 102.71 98.045 ;
      RECT  104.69 100.335 104.9 99.955 ;
      RECT  103.25 99.75 103.43 98.045 ;
      RECT  103.97 99.75 104.15 98.045 ;
      RECT  103.25 100.665 103.43 99.75 ;
      RECT  105.41 100.665 105.62 100.335 ;
      RECT  103.61 99.75 103.79 98.045 ;
      RECT  103.61 100.665 103.79 99.75 ;
      RECT  102.29 99.955 102.5 99.75 ;
      RECT  105.41 100.335 105.62 99.955 ;
      RECT  104.33 99.75 104.51 98.045 ;
      RECT  102.5 99.955 102.71 99.75 ;
      RECT  102.29 100.335 102.5 99.955 ;
      POLYGON  104.9 98.67 104.9 98.26 105.155 98.26 105.155 98.59 105.075 98.67 104.9 98.67 ;
      RECT  102.89 100.665 103.07 99.75 ;
      RECT  102.5 100.665 102.71 100.335 ;
      RECT  102.5 100.335 102.71 99.955 ;
      RECT  104.69 100.63 104.9 101.04 ;
      RECT  102.29 99.625 102.5 99.955 ;
      RECT  105.335 100.54 105.41 102.245 ;
      RECT  105.25 101.125 105.335 101.535 ;
      RECT  104.33 99.625 104.51 100.54 ;
      POLYGON  105.335 99.625 105.335 99.955 104.9 99.955 104.9 100.335 105.335 100.335 105.335 100.54 105.41 100.54 105.41 99.625 105.335 99.625 ;
      RECT  105.41 100.54 105.62 102.245 ;
      POLYGON  104.9 100.63 104.9 101.04 105.075 101.04 105.155 100.96 105.155 100.63 104.9 100.63 ;
      RECT  102.29 100.54 102.5 102.245 ;
      RECT  103.97 99.625 104.15 100.54 ;
      RECT  102.89 100.54 103.07 102.245 ;
      RECT  104.69 101.62 104.9 102.03 ;
      RECT  105.41 100.335 105.62 100.54 ;
      RECT  102.5 100.54 102.71 102.245 ;
      RECT  104.69 99.955 104.9 100.335 ;
      RECT  103.25 100.54 103.43 102.245 ;
      RECT  103.97 100.54 104.15 102.245 ;
      RECT  103.25 99.625 103.43 100.54 ;
      RECT  105.41 99.625 105.62 99.955 ;
      RECT  103.61 100.54 103.79 102.245 ;
      RECT  103.61 99.625 103.79 100.54 ;
      RECT  102.29 100.335 102.5 100.54 ;
      RECT  105.41 99.955 105.62 100.335 ;
      RECT  104.33 100.54 104.51 102.245 ;
      RECT  102.5 100.335 102.71 100.54 ;
      RECT  102.29 99.955 102.5 100.335 ;
      POLYGON  104.9 101.62 104.9 102.03 105.155 102.03 105.155 101.7 105.075 101.62 104.9 101.62 ;
      RECT  102.89 99.625 103.07 100.54 ;
      RECT  102.5 99.625 102.71 99.955 ;
      RECT  102.5 99.955 102.71 100.335 ;
      RECT  104.69 103.61 104.9 103.2 ;
      RECT  102.29 104.615 102.5 104.285 ;
      RECT  105.335 103.7 105.41 101.995 ;
      RECT  105.25 103.115 105.335 102.705 ;
      RECT  104.33 104.615 104.51 103.7 ;
      POLYGON  105.335 104.615 105.335 104.285 104.9 104.285 104.9 103.905 105.335 103.905 105.335 103.7 105.41 103.7 105.41 104.615 105.335 104.615 ;
      RECT  105.41 103.7 105.62 101.995 ;
      POLYGON  104.9 103.61 104.9 103.2 105.075 103.2 105.155 103.28 105.155 103.61 104.9 103.61 ;
      RECT  102.29 103.7 102.5 101.995 ;
      RECT  103.97 104.615 104.15 103.7 ;
      RECT  102.89 103.7 103.07 101.995 ;
      RECT  104.69 102.62 104.9 102.21 ;
      RECT  105.41 103.905 105.62 103.7 ;
      RECT  102.5 103.7 102.71 101.995 ;
      RECT  104.69 104.285 104.9 103.905 ;
      RECT  103.25 103.7 103.43 101.995 ;
      RECT  103.97 103.7 104.15 101.995 ;
      RECT  103.25 104.615 103.43 103.7 ;
      RECT  105.41 104.615 105.62 104.285 ;
      RECT  103.61 103.7 103.79 101.995 ;
      RECT  103.61 104.615 103.79 103.7 ;
      RECT  102.29 103.905 102.5 103.7 ;
      RECT  105.41 104.285 105.62 103.905 ;
      RECT  104.33 103.7 104.51 101.995 ;
      RECT  102.5 103.905 102.71 103.7 ;
      RECT  102.29 104.285 102.5 103.905 ;
      POLYGON  104.9 102.62 104.9 102.21 105.155 102.21 105.155 102.54 105.075 102.62 104.9 102.62 ;
      RECT  102.89 104.615 103.07 103.7 ;
      RECT  102.5 104.615 102.71 104.285 ;
      RECT  102.5 104.285 102.71 103.905 ;
      RECT  104.69 104.58 104.9 104.99 ;
      RECT  102.29 103.575 102.5 103.905 ;
      RECT  105.335 104.49 105.41 106.195 ;
      RECT  105.25 105.075 105.335 105.485 ;
      RECT  104.33 103.575 104.51 104.49 ;
      POLYGON  105.335 103.575 105.335 103.905 104.9 103.905 104.9 104.285 105.335 104.285 105.335 104.49 105.41 104.49 105.41 103.575 105.335 103.575 ;
      RECT  105.41 104.49 105.62 106.195 ;
      POLYGON  104.9 104.58 104.9 104.99 105.075 104.99 105.155 104.91 105.155 104.58 104.9 104.58 ;
      RECT  102.29 104.49 102.5 106.195 ;
      RECT  103.97 103.575 104.15 104.49 ;
      RECT  102.89 104.49 103.07 106.195 ;
      RECT  104.69 105.57 104.9 105.98 ;
      RECT  105.41 104.285 105.62 104.49 ;
      RECT  102.5 104.49 102.71 106.195 ;
      RECT  104.69 103.905 104.9 104.285 ;
      RECT  103.25 104.49 103.43 106.195 ;
      RECT  103.97 104.49 104.15 106.195 ;
      RECT  103.25 103.575 103.43 104.49 ;
      RECT  105.41 103.575 105.62 103.905 ;
      RECT  103.61 104.49 103.79 106.195 ;
      RECT  103.61 103.575 103.79 104.49 ;
      RECT  102.29 104.285 102.5 104.49 ;
      RECT  105.41 103.905 105.62 104.285 ;
      RECT  104.33 104.49 104.51 106.195 ;
      RECT  102.5 104.285 102.71 104.49 ;
      RECT  102.29 103.905 102.5 104.285 ;
      POLYGON  104.9 105.57 104.9 105.98 105.155 105.98 105.155 105.65 105.075 105.57 104.9 105.57 ;
      RECT  102.89 103.575 103.07 104.49 ;
      RECT  102.5 103.575 102.71 103.905 ;
      RECT  102.5 103.905 102.71 104.285 ;
      RECT  104.69 107.56 104.9 107.15 ;
      RECT  102.29 108.565 102.5 108.235 ;
      RECT  105.335 107.65 105.41 105.945 ;
      RECT  105.25 107.065 105.335 106.655 ;
      RECT  104.33 108.565 104.51 107.65 ;
      POLYGON  105.335 108.565 105.335 108.235 104.9 108.235 104.9 107.855 105.335 107.855 105.335 107.65 105.41 107.65 105.41 108.565 105.335 108.565 ;
      RECT  105.41 107.65 105.62 105.945 ;
      POLYGON  104.9 107.56 104.9 107.15 105.075 107.15 105.155 107.23 105.155 107.56 104.9 107.56 ;
      RECT  102.29 107.65 102.5 105.945 ;
      RECT  103.97 108.565 104.15 107.65 ;
      RECT  102.89 107.65 103.07 105.945 ;
      RECT  104.69 106.57 104.9 106.16 ;
      RECT  105.41 107.855 105.62 107.65 ;
      RECT  102.5 107.65 102.71 105.945 ;
      RECT  104.69 108.235 104.9 107.855 ;
      RECT  103.25 107.65 103.43 105.945 ;
      RECT  103.97 107.65 104.15 105.945 ;
      RECT  103.25 108.565 103.43 107.65 ;
      RECT  105.41 108.565 105.62 108.235 ;
      RECT  103.61 107.65 103.79 105.945 ;
      RECT  103.61 108.565 103.79 107.65 ;
      RECT  102.29 107.855 102.5 107.65 ;
      RECT  105.41 108.235 105.62 107.855 ;
      RECT  104.33 107.65 104.51 105.945 ;
      RECT  102.5 107.855 102.71 107.65 ;
      RECT  102.29 108.235 102.5 107.855 ;
      POLYGON  104.9 106.57 104.9 106.16 105.155 106.16 105.155 106.49 105.075 106.57 104.9 106.57 ;
      RECT  102.89 108.565 103.07 107.65 ;
      RECT  102.5 108.565 102.71 108.235 ;
      RECT  102.5 108.235 102.71 107.855 ;
      RECT  104.69 108.53 104.9 108.94 ;
      RECT  102.29 107.525 102.5 107.855 ;
      RECT  105.335 108.44 105.41 110.145 ;
      RECT  105.25 109.025 105.335 109.435 ;
      RECT  104.33 107.525 104.51 108.44 ;
      POLYGON  105.335 107.525 105.335 107.855 104.9 107.855 104.9 108.235 105.335 108.235 105.335 108.44 105.41 108.44 105.41 107.525 105.335 107.525 ;
      RECT  105.41 108.44 105.62 110.145 ;
      POLYGON  104.9 108.53 104.9 108.94 105.075 108.94 105.155 108.86 105.155 108.53 104.9 108.53 ;
      RECT  102.29 108.44 102.5 110.145 ;
      RECT  103.97 107.525 104.15 108.44 ;
      RECT  102.89 108.44 103.07 110.145 ;
      RECT  104.69 109.52 104.9 109.93 ;
      RECT  105.41 108.235 105.62 108.44 ;
      RECT  102.5 108.44 102.71 110.145 ;
      RECT  104.69 107.855 104.9 108.235 ;
      RECT  103.25 108.44 103.43 110.145 ;
      RECT  103.97 108.44 104.15 110.145 ;
      RECT  103.25 107.525 103.43 108.44 ;
      RECT  105.41 107.525 105.62 107.855 ;
      RECT  103.61 108.44 103.79 110.145 ;
      RECT  103.61 107.525 103.79 108.44 ;
      RECT  102.29 108.235 102.5 108.44 ;
      RECT  105.41 107.855 105.62 108.235 ;
      RECT  104.33 108.44 104.51 110.145 ;
      RECT  102.5 108.235 102.71 108.44 ;
      RECT  102.29 107.855 102.5 108.235 ;
      POLYGON  104.9 109.52 104.9 109.93 105.155 109.93 105.155 109.6 105.075 109.52 104.9 109.52 ;
      RECT  102.89 107.525 103.07 108.44 ;
      RECT  102.5 107.525 102.71 107.855 ;
      RECT  102.5 107.855 102.71 108.235 ;
      RECT  104.69 111.51 104.9 111.1 ;
      RECT  102.29 112.515 102.5 112.185 ;
      RECT  105.335 111.6 105.41 109.895 ;
      RECT  105.25 111.015 105.335 110.605 ;
      RECT  104.33 112.515 104.51 111.6 ;
      POLYGON  105.335 112.515 105.335 112.185 104.9 112.185 104.9 111.805 105.335 111.805 105.335 111.6 105.41 111.6 105.41 112.515 105.335 112.515 ;
      RECT  105.41 111.6 105.62 109.895 ;
      POLYGON  104.9 111.51 104.9 111.1 105.075 111.1 105.155 111.18 105.155 111.51 104.9 111.51 ;
      RECT  102.29 111.6 102.5 109.895 ;
      RECT  103.97 112.515 104.15 111.6 ;
      RECT  102.89 111.6 103.07 109.895 ;
      RECT  104.69 110.52 104.9 110.11 ;
      RECT  105.41 111.805 105.62 111.6 ;
      RECT  102.5 111.6 102.71 109.895 ;
      RECT  104.69 112.185 104.9 111.805 ;
      RECT  103.25 111.6 103.43 109.895 ;
      RECT  103.97 111.6 104.15 109.895 ;
      RECT  103.25 112.515 103.43 111.6 ;
      RECT  105.41 112.515 105.62 112.185 ;
      RECT  103.61 111.6 103.79 109.895 ;
      RECT  103.61 112.515 103.79 111.6 ;
      RECT  102.29 111.805 102.5 111.6 ;
      RECT  105.41 112.185 105.62 111.805 ;
      RECT  104.33 111.6 104.51 109.895 ;
      RECT  102.5 111.805 102.71 111.6 ;
      RECT  102.29 112.185 102.5 111.805 ;
      POLYGON  104.9 110.52 104.9 110.11 105.155 110.11 105.155 110.44 105.075 110.52 104.9 110.52 ;
      RECT  102.89 112.515 103.07 111.6 ;
      RECT  102.5 112.515 102.71 112.185 ;
      RECT  102.5 112.185 102.71 111.805 ;
      RECT  104.69 112.48 104.9 112.89 ;
      RECT  102.29 111.475 102.5 111.805 ;
      RECT  105.335 112.39 105.41 114.095 ;
      RECT  105.25 112.975 105.335 113.385 ;
      RECT  104.33 111.475 104.51 112.39 ;
      POLYGON  105.335 111.475 105.335 111.805 104.9 111.805 104.9 112.185 105.335 112.185 105.335 112.39 105.41 112.39 105.41 111.475 105.335 111.475 ;
      RECT  105.41 112.39 105.62 114.095 ;
      POLYGON  104.9 112.48 104.9 112.89 105.075 112.89 105.155 112.81 105.155 112.48 104.9 112.48 ;
      RECT  102.29 112.39 102.5 114.095 ;
      RECT  103.97 111.475 104.15 112.39 ;
      RECT  102.89 112.39 103.07 114.095 ;
      RECT  104.69 113.47 104.9 113.88 ;
      RECT  105.41 112.185 105.62 112.39 ;
      RECT  102.5 112.39 102.71 114.095 ;
      RECT  104.69 111.805 104.9 112.185 ;
      RECT  103.25 112.39 103.43 114.095 ;
      RECT  103.97 112.39 104.15 114.095 ;
      RECT  103.25 111.475 103.43 112.39 ;
      RECT  105.41 111.475 105.62 111.805 ;
      RECT  103.61 112.39 103.79 114.095 ;
      RECT  103.61 111.475 103.79 112.39 ;
      RECT  102.29 112.185 102.5 112.39 ;
      RECT  105.41 111.805 105.62 112.185 ;
      RECT  104.33 112.39 104.51 114.095 ;
      RECT  102.5 112.185 102.71 112.39 ;
      RECT  102.29 111.805 102.5 112.185 ;
      POLYGON  104.9 113.47 104.9 113.88 105.155 113.88 105.155 113.55 105.075 113.47 104.9 113.47 ;
      RECT  102.89 111.475 103.07 112.39 ;
      RECT  102.5 111.475 102.71 111.805 ;
      RECT  102.5 111.805 102.71 112.185 ;
      RECT  104.69 115.46 104.9 115.05 ;
      RECT  102.29 116.465 102.5 116.135 ;
      RECT  105.335 115.55 105.41 113.845 ;
      RECT  105.25 114.965 105.335 114.555 ;
      RECT  104.33 116.465 104.51 115.55 ;
      POLYGON  105.335 116.465 105.335 116.135 104.9 116.135 104.9 115.755 105.335 115.755 105.335 115.55 105.41 115.55 105.41 116.465 105.335 116.465 ;
      RECT  105.41 115.55 105.62 113.845 ;
      POLYGON  104.9 115.46 104.9 115.05 105.075 115.05 105.155 115.13 105.155 115.46 104.9 115.46 ;
      RECT  102.29 115.55 102.5 113.845 ;
      RECT  103.97 116.465 104.15 115.55 ;
      RECT  102.89 115.55 103.07 113.845 ;
      RECT  104.69 114.47 104.9 114.06 ;
      RECT  105.41 115.755 105.62 115.55 ;
      RECT  102.5 115.55 102.71 113.845 ;
      RECT  104.69 116.135 104.9 115.755 ;
      RECT  103.25 115.55 103.43 113.845 ;
      RECT  103.97 115.55 104.15 113.845 ;
      RECT  103.25 116.465 103.43 115.55 ;
      RECT  105.41 116.465 105.62 116.135 ;
      RECT  103.61 115.55 103.79 113.845 ;
      RECT  103.61 116.465 103.79 115.55 ;
      RECT  102.29 115.755 102.5 115.55 ;
      RECT  105.41 116.135 105.62 115.755 ;
      RECT  104.33 115.55 104.51 113.845 ;
      RECT  102.5 115.755 102.71 115.55 ;
      RECT  102.29 116.135 102.5 115.755 ;
      POLYGON  104.9 114.47 104.9 114.06 105.155 114.06 105.155 114.39 105.075 114.47 104.9 114.47 ;
      RECT  102.89 116.465 103.07 115.55 ;
      RECT  102.5 116.465 102.71 116.135 ;
      RECT  102.5 116.135 102.71 115.755 ;
      RECT  104.69 116.43 104.9 116.84 ;
      RECT  102.29 115.425 102.5 115.755 ;
      RECT  105.335 116.34 105.41 118.045 ;
      RECT  105.25 116.925 105.335 117.335 ;
      RECT  104.33 115.425 104.51 116.34 ;
      POLYGON  105.335 115.425 105.335 115.755 104.9 115.755 104.9 116.135 105.335 116.135 105.335 116.34 105.41 116.34 105.41 115.425 105.335 115.425 ;
      RECT  105.41 116.34 105.62 118.045 ;
      POLYGON  104.9 116.43 104.9 116.84 105.075 116.84 105.155 116.76 105.155 116.43 104.9 116.43 ;
      RECT  102.29 116.34 102.5 118.045 ;
      RECT  103.97 115.425 104.15 116.34 ;
      RECT  102.89 116.34 103.07 118.045 ;
      RECT  104.69 117.42 104.9 117.83 ;
      RECT  105.41 116.135 105.62 116.34 ;
      RECT  102.5 116.34 102.71 118.045 ;
      RECT  104.69 115.755 104.9 116.135 ;
      RECT  103.25 116.34 103.43 118.045 ;
      RECT  103.97 116.34 104.15 118.045 ;
      RECT  103.25 115.425 103.43 116.34 ;
      RECT  105.41 115.425 105.62 115.755 ;
      RECT  103.61 116.34 103.79 118.045 ;
      RECT  103.61 115.425 103.79 116.34 ;
      RECT  102.29 116.135 102.5 116.34 ;
      RECT  105.41 115.755 105.62 116.135 ;
      RECT  104.33 116.34 104.51 118.045 ;
      RECT  102.5 116.135 102.71 116.34 ;
      RECT  102.29 115.755 102.5 116.135 ;
      POLYGON  104.9 117.42 104.9 117.83 105.155 117.83 105.155 117.5 105.075 117.42 104.9 117.42 ;
      RECT  102.89 115.425 103.07 116.34 ;
      RECT  102.5 115.425 102.71 115.755 ;
      RECT  102.5 115.755 102.71 116.135 ;
      RECT  104.69 119.41 104.9 119.0 ;
      RECT  102.29 120.415 102.5 120.085 ;
      RECT  105.335 119.5 105.41 117.795 ;
      RECT  105.25 118.915 105.335 118.505 ;
      RECT  104.33 120.415 104.51 119.5 ;
      POLYGON  105.335 120.415 105.335 120.085 104.9 120.085 104.9 119.705 105.335 119.705 105.335 119.5 105.41 119.5 105.41 120.415 105.335 120.415 ;
      RECT  105.41 119.5 105.62 117.795 ;
      POLYGON  104.9 119.41 104.9 119.0 105.075 119.0 105.155 119.08 105.155 119.41 104.9 119.41 ;
      RECT  102.29 119.5 102.5 117.795 ;
      RECT  103.97 120.415 104.15 119.5 ;
      RECT  102.89 119.5 103.07 117.795 ;
      RECT  104.69 118.42 104.9 118.01 ;
      RECT  105.41 119.705 105.62 119.5 ;
      RECT  102.5 119.5 102.71 117.795 ;
      RECT  104.69 120.085 104.9 119.705 ;
      RECT  103.25 119.5 103.43 117.795 ;
      RECT  103.97 119.5 104.15 117.795 ;
      RECT  103.25 120.415 103.43 119.5 ;
      RECT  105.41 120.415 105.62 120.085 ;
      RECT  103.61 119.5 103.79 117.795 ;
      RECT  103.61 120.415 103.79 119.5 ;
      RECT  102.29 119.705 102.5 119.5 ;
      RECT  105.41 120.085 105.62 119.705 ;
      RECT  104.33 119.5 104.51 117.795 ;
      RECT  102.5 119.705 102.71 119.5 ;
      RECT  102.29 120.085 102.5 119.705 ;
      POLYGON  104.9 118.42 104.9 118.01 105.155 118.01 105.155 118.34 105.075 118.42 104.9 118.42 ;
      RECT  102.89 120.415 103.07 119.5 ;
      RECT  102.5 120.415 102.71 120.085 ;
      RECT  102.5 120.085 102.71 119.705 ;
      RECT  104.69 120.38 104.9 120.79 ;
      RECT  102.29 119.375 102.5 119.705 ;
      RECT  105.335 120.29 105.41 121.995 ;
      RECT  105.25 120.875 105.335 121.285 ;
      RECT  104.33 119.375 104.51 120.29 ;
      POLYGON  105.335 119.375 105.335 119.705 104.9 119.705 104.9 120.085 105.335 120.085 105.335 120.29 105.41 120.29 105.41 119.375 105.335 119.375 ;
      RECT  105.41 120.29 105.62 121.995 ;
      POLYGON  104.9 120.38 104.9 120.79 105.075 120.79 105.155 120.71 105.155 120.38 104.9 120.38 ;
      RECT  102.29 120.29 102.5 121.995 ;
      RECT  103.97 119.375 104.15 120.29 ;
      RECT  102.89 120.29 103.07 121.995 ;
      RECT  104.69 121.37 104.9 121.78 ;
      RECT  105.41 120.085 105.62 120.29 ;
      RECT  102.5 120.29 102.71 121.995 ;
      RECT  104.69 119.705 104.9 120.085 ;
      RECT  103.25 120.29 103.43 121.995 ;
      RECT  103.97 120.29 104.15 121.995 ;
      RECT  103.25 119.375 103.43 120.29 ;
      RECT  105.41 119.375 105.62 119.705 ;
      RECT  103.61 120.29 103.79 121.995 ;
      RECT  103.61 119.375 103.79 120.29 ;
      RECT  102.29 120.085 102.5 120.29 ;
      RECT  105.41 119.705 105.62 120.085 ;
      RECT  104.33 120.29 104.51 121.995 ;
      RECT  102.5 120.085 102.71 120.29 ;
      RECT  102.29 119.705 102.5 120.085 ;
      POLYGON  104.9 121.37 104.9 121.78 105.155 121.78 105.155 121.45 105.075 121.37 104.9 121.37 ;
      RECT  102.89 119.375 103.07 120.29 ;
      RECT  102.5 119.375 102.71 119.705 ;
      RECT  102.5 119.705 102.71 120.085 ;
      RECT  104.69 123.36 104.9 122.95 ;
      RECT  102.29 124.365 102.5 124.035 ;
      RECT  105.335 123.45 105.41 121.745 ;
      RECT  105.25 122.865 105.335 122.455 ;
      RECT  104.33 124.365 104.51 123.45 ;
      POLYGON  105.335 124.365 105.335 124.035 104.9 124.035 104.9 123.655 105.335 123.655 105.335 123.45 105.41 123.45 105.41 124.365 105.335 124.365 ;
      RECT  105.41 123.45 105.62 121.745 ;
      POLYGON  104.9 123.36 104.9 122.95 105.075 122.95 105.155 123.03 105.155 123.36 104.9 123.36 ;
      RECT  102.29 123.45 102.5 121.745 ;
      RECT  103.97 124.365 104.15 123.45 ;
      RECT  102.89 123.45 103.07 121.745 ;
      RECT  104.69 122.37 104.9 121.96 ;
      RECT  105.41 123.655 105.62 123.45 ;
      RECT  102.5 123.45 102.71 121.745 ;
      RECT  104.69 124.035 104.9 123.655 ;
      RECT  103.25 123.45 103.43 121.745 ;
      RECT  103.97 123.45 104.15 121.745 ;
      RECT  103.25 124.365 103.43 123.45 ;
      RECT  105.41 124.365 105.62 124.035 ;
      RECT  103.61 123.45 103.79 121.745 ;
      RECT  103.61 124.365 103.79 123.45 ;
      RECT  102.29 123.655 102.5 123.45 ;
      RECT  105.41 124.035 105.62 123.655 ;
      RECT  104.33 123.45 104.51 121.745 ;
      RECT  102.5 123.655 102.71 123.45 ;
      RECT  102.29 124.035 102.5 123.655 ;
      POLYGON  104.9 122.37 104.9 121.96 105.155 121.96 105.155 122.29 105.075 122.37 104.9 122.37 ;
      RECT  102.89 124.365 103.07 123.45 ;
      RECT  102.5 124.365 102.71 124.035 ;
      RECT  102.5 124.035 102.71 123.655 ;
      RECT  106.55 92.73 106.34 93.14 ;
      RECT  108.95 91.725 108.74 92.055 ;
      RECT  105.905 92.64 105.83 94.345 ;
      RECT  105.99 93.225 105.905 93.635 ;
      RECT  106.91 91.725 106.73 92.64 ;
      POLYGON  105.905 91.725 105.905 92.055 106.34 92.055 106.34 92.435 105.905 92.435 105.905 92.64 105.83 92.64 105.83 91.725 105.905 91.725 ;
      RECT  105.83 92.64 105.62 94.345 ;
      POLYGON  106.34 92.73 106.34 93.14 106.165 93.14 106.085 93.06 106.085 92.73 106.34 92.73 ;
      RECT  108.95 92.64 108.74 94.345 ;
      RECT  107.27 91.725 107.09 92.64 ;
      RECT  108.35 92.64 108.17 94.345 ;
      RECT  106.55 93.72 106.34 94.13 ;
      RECT  105.83 92.435 105.62 92.64 ;
      RECT  108.74 92.64 108.53 94.345 ;
      RECT  106.55 92.055 106.34 92.435 ;
      RECT  107.99 92.64 107.81 94.345 ;
      RECT  107.27 92.64 107.09 94.345 ;
      RECT  107.99 91.725 107.81 92.64 ;
      RECT  105.83 91.725 105.62 92.055 ;
      RECT  107.63 92.64 107.45 94.345 ;
      RECT  107.63 91.725 107.45 92.64 ;
      RECT  108.95 92.435 108.74 92.64 ;
      RECT  105.83 92.055 105.62 92.435 ;
      RECT  106.91 92.64 106.73 94.345 ;
      RECT  108.74 92.435 108.53 92.64 ;
      RECT  108.95 92.055 108.74 92.435 ;
      POLYGON  106.34 93.72 106.34 94.13 106.085 94.13 106.085 93.8 106.165 93.72 106.34 93.72 ;
      RECT  108.35 91.725 108.17 92.64 ;
      RECT  108.74 91.725 108.53 92.055 ;
      RECT  108.74 92.055 108.53 92.435 ;
      RECT  106.55 95.71 106.34 95.3 ;
      RECT  108.95 96.715 108.74 96.385 ;
      RECT  105.905 95.8 105.83 94.095 ;
      RECT  105.99 95.215 105.905 94.805 ;
      RECT  106.91 96.715 106.73 95.8 ;
      POLYGON  105.905 96.715 105.905 96.385 106.34 96.385 106.34 96.005 105.905 96.005 105.905 95.8 105.83 95.8 105.83 96.715 105.905 96.715 ;
      RECT  105.83 95.8 105.62 94.095 ;
      POLYGON  106.34 95.71 106.34 95.3 106.165 95.3 106.085 95.38 106.085 95.71 106.34 95.71 ;
      RECT  108.95 95.8 108.74 94.095 ;
      RECT  107.27 96.715 107.09 95.8 ;
      RECT  108.35 95.8 108.17 94.095 ;
      RECT  106.55 94.72 106.34 94.31 ;
      RECT  105.83 96.005 105.62 95.8 ;
      RECT  108.74 95.8 108.53 94.095 ;
      RECT  106.55 96.385 106.34 96.005 ;
      RECT  107.99 95.8 107.81 94.095 ;
      RECT  107.27 95.8 107.09 94.095 ;
      RECT  107.99 96.715 107.81 95.8 ;
      RECT  105.83 96.715 105.62 96.385 ;
      RECT  107.63 95.8 107.45 94.095 ;
      RECT  107.63 96.715 107.45 95.8 ;
      RECT  108.95 96.005 108.74 95.8 ;
      RECT  105.83 96.385 105.62 96.005 ;
      RECT  106.91 95.8 106.73 94.095 ;
      RECT  108.74 96.005 108.53 95.8 ;
      RECT  108.95 96.385 108.74 96.005 ;
      POLYGON  106.34 94.72 106.34 94.31 106.085 94.31 106.085 94.64 106.165 94.72 106.34 94.72 ;
      RECT  108.35 96.715 108.17 95.8 ;
      RECT  108.74 96.715 108.53 96.385 ;
      RECT  108.74 96.385 108.53 96.005 ;
      RECT  106.55 96.68 106.34 97.09 ;
      RECT  108.95 95.675 108.74 96.005 ;
      RECT  105.905 96.59 105.83 98.295 ;
      RECT  105.99 97.175 105.905 97.585 ;
      RECT  106.91 95.675 106.73 96.59 ;
      POLYGON  105.905 95.675 105.905 96.005 106.34 96.005 106.34 96.385 105.905 96.385 105.905 96.59 105.83 96.59 105.83 95.675 105.905 95.675 ;
      RECT  105.83 96.59 105.62 98.295 ;
      POLYGON  106.34 96.68 106.34 97.09 106.165 97.09 106.085 97.01 106.085 96.68 106.34 96.68 ;
      RECT  108.95 96.59 108.74 98.295 ;
      RECT  107.27 95.675 107.09 96.59 ;
      RECT  108.35 96.59 108.17 98.295 ;
      RECT  106.55 97.67 106.34 98.08 ;
      RECT  105.83 96.385 105.62 96.59 ;
      RECT  108.74 96.59 108.53 98.295 ;
      RECT  106.55 96.005 106.34 96.385 ;
      RECT  107.99 96.59 107.81 98.295 ;
      RECT  107.27 96.59 107.09 98.295 ;
      RECT  107.99 95.675 107.81 96.59 ;
      RECT  105.83 95.675 105.62 96.005 ;
      RECT  107.63 96.59 107.45 98.295 ;
      RECT  107.63 95.675 107.45 96.59 ;
      RECT  108.95 96.385 108.74 96.59 ;
      RECT  105.83 96.005 105.62 96.385 ;
      RECT  106.91 96.59 106.73 98.295 ;
      RECT  108.74 96.385 108.53 96.59 ;
      RECT  108.95 96.005 108.74 96.385 ;
      POLYGON  106.34 97.67 106.34 98.08 106.085 98.08 106.085 97.75 106.165 97.67 106.34 97.67 ;
      RECT  108.35 95.675 108.17 96.59 ;
      RECT  108.74 95.675 108.53 96.005 ;
      RECT  108.74 96.005 108.53 96.385 ;
      RECT  106.55 99.66 106.34 99.25 ;
      RECT  108.95 100.665 108.74 100.335 ;
      RECT  105.905 99.75 105.83 98.045 ;
      RECT  105.99 99.165 105.905 98.755 ;
      RECT  106.91 100.665 106.73 99.75 ;
      POLYGON  105.905 100.665 105.905 100.335 106.34 100.335 106.34 99.955 105.905 99.955 105.905 99.75 105.83 99.75 105.83 100.665 105.905 100.665 ;
      RECT  105.83 99.75 105.62 98.045 ;
      POLYGON  106.34 99.66 106.34 99.25 106.165 99.25 106.085 99.33 106.085 99.66 106.34 99.66 ;
      RECT  108.95 99.75 108.74 98.045 ;
      RECT  107.27 100.665 107.09 99.75 ;
      RECT  108.35 99.75 108.17 98.045 ;
      RECT  106.55 98.67 106.34 98.26 ;
      RECT  105.83 99.955 105.62 99.75 ;
      RECT  108.74 99.75 108.53 98.045 ;
      RECT  106.55 100.335 106.34 99.955 ;
      RECT  107.99 99.75 107.81 98.045 ;
      RECT  107.27 99.75 107.09 98.045 ;
      RECT  107.99 100.665 107.81 99.75 ;
      RECT  105.83 100.665 105.62 100.335 ;
      RECT  107.63 99.75 107.45 98.045 ;
      RECT  107.63 100.665 107.45 99.75 ;
      RECT  108.95 99.955 108.74 99.75 ;
      RECT  105.83 100.335 105.62 99.955 ;
      RECT  106.91 99.75 106.73 98.045 ;
      RECT  108.74 99.955 108.53 99.75 ;
      RECT  108.95 100.335 108.74 99.955 ;
      POLYGON  106.34 98.67 106.34 98.26 106.085 98.26 106.085 98.59 106.165 98.67 106.34 98.67 ;
      RECT  108.35 100.665 108.17 99.75 ;
      RECT  108.74 100.665 108.53 100.335 ;
      RECT  108.74 100.335 108.53 99.955 ;
      RECT  106.55 100.63 106.34 101.04 ;
      RECT  108.95 99.625 108.74 99.955 ;
      RECT  105.905 100.54 105.83 102.245 ;
      RECT  105.99 101.125 105.905 101.535 ;
      RECT  106.91 99.625 106.73 100.54 ;
      POLYGON  105.905 99.625 105.905 99.955 106.34 99.955 106.34 100.335 105.905 100.335 105.905 100.54 105.83 100.54 105.83 99.625 105.905 99.625 ;
      RECT  105.83 100.54 105.62 102.245 ;
      POLYGON  106.34 100.63 106.34 101.04 106.165 101.04 106.085 100.96 106.085 100.63 106.34 100.63 ;
      RECT  108.95 100.54 108.74 102.245 ;
      RECT  107.27 99.625 107.09 100.54 ;
      RECT  108.35 100.54 108.17 102.245 ;
      RECT  106.55 101.62 106.34 102.03 ;
      RECT  105.83 100.335 105.62 100.54 ;
      RECT  108.74 100.54 108.53 102.245 ;
      RECT  106.55 99.955 106.34 100.335 ;
      RECT  107.99 100.54 107.81 102.245 ;
      RECT  107.27 100.54 107.09 102.245 ;
      RECT  107.99 99.625 107.81 100.54 ;
      RECT  105.83 99.625 105.62 99.955 ;
      RECT  107.63 100.54 107.45 102.245 ;
      RECT  107.63 99.625 107.45 100.54 ;
      RECT  108.95 100.335 108.74 100.54 ;
      RECT  105.83 99.955 105.62 100.335 ;
      RECT  106.91 100.54 106.73 102.245 ;
      RECT  108.74 100.335 108.53 100.54 ;
      RECT  108.95 99.955 108.74 100.335 ;
      POLYGON  106.34 101.62 106.34 102.03 106.085 102.03 106.085 101.7 106.165 101.62 106.34 101.62 ;
      RECT  108.35 99.625 108.17 100.54 ;
      RECT  108.74 99.625 108.53 99.955 ;
      RECT  108.74 99.955 108.53 100.335 ;
      RECT  106.55 103.61 106.34 103.2 ;
      RECT  108.95 104.615 108.74 104.285 ;
      RECT  105.905 103.7 105.83 101.995 ;
      RECT  105.99 103.115 105.905 102.705 ;
      RECT  106.91 104.615 106.73 103.7 ;
      POLYGON  105.905 104.615 105.905 104.285 106.34 104.285 106.34 103.905 105.905 103.905 105.905 103.7 105.83 103.7 105.83 104.615 105.905 104.615 ;
      RECT  105.83 103.7 105.62 101.995 ;
      POLYGON  106.34 103.61 106.34 103.2 106.165 103.2 106.085 103.28 106.085 103.61 106.34 103.61 ;
      RECT  108.95 103.7 108.74 101.995 ;
      RECT  107.27 104.615 107.09 103.7 ;
      RECT  108.35 103.7 108.17 101.995 ;
      RECT  106.55 102.62 106.34 102.21 ;
      RECT  105.83 103.905 105.62 103.7 ;
      RECT  108.74 103.7 108.53 101.995 ;
      RECT  106.55 104.285 106.34 103.905 ;
      RECT  107.99 103.7 107.81 101.995 ;
      RECT  107.27 103.7 107.09 101.995 ;
      RECT  107.99 104.615 107.81 103.7 ;
      RECT  105.83 104.615 105.62 104.285 ;
      RECT  107.63 103.7 107.45 101.995 ;
      RECT  107.63 104.615 107.45 103.7 ;
      RECT  108.95 103.905 108.74 103.7 ;
      RECT  105.83 104.285 105.62 103.905 ;
      RECT  106.91 103.7 106.73 101.995 ;
      RECT  108.74 103.905 108.53 103.7 ;
      RECT  108.95 104.285 108.74 103.905 ;
      POLYGON  106.34 102.62 106.34 102.21 106.085 102.21 106.085 102.54 106.165 102.62 106.34 102.62 ;
      RECT  108.35 104.615 108.17 103.7 ;
      RECT  108.74 104.615 108.53 104.285 ;
      RECT  108.74 104.285 108.53 103.905 ;
      RECT  106.55 104.58 106.34 104.99 ;
      RECT  108.95 103.575 108.74 103.905 ;
      RECT  105.905 104.49 105.83 106.195 ;
      RECT  105.99 105.075 105.905 105.485 ;
      RECT  106.91 103.575 106.73 104.49 ;
      POLYGON  105.905 103.575 105.905 103.905 106.34 103.905 106.34 104.285 105.905 104.285 105.905 104.49 105.83 104.49 105.83 103.575 105.905 103.575 ;
      RECT  105.83 104.49 105.62 106.195 ;
      POLYGON  106.34 104.58 106.34 104.99 106.165 104.99 106.085 104.91 106.085 104.58 106.34 104.58 ;
      RECT  108.95 104.49 108.74 106.195 ;
      RECT  107.27 103.575 107.09 104.49 ;
      RECT  108.35 104.49 108.17 106.195 ;
      RECT  106.55 105.57 106.34 105.98 ;
      RECT  105.83 104.285 105.62 104.49 ;
      RECT  108.74 104.49 108.53 106.195 ;
      RECT  106.55 103.905 106.34 104.285 ;
      RECT  107.99 104.49 107.81 106.195 ;
      RECT  107.27 104.49 107.09 106.195 ;
      RECT  107.99 103.575 107.81 104.49 ;
      RECT  105.83 103.575 105.62 103.905 ;
      RECT  107.63 104.49 107.45 106.195 ;
      RECT  107.63 103.575 107.45 104.49 ;
      RECT  108.95 104.285 108.74 104.49 ;
      RECT  105.83 103.905 105.62 104.285 ;
      RECT  106.91 104.49 106.73 106.195 ;
      RECT  108.74 104.285 108.53 104.49 ;
      RECT  108.95 103.905 108.74 104.285 ;
      POLYGON  106.34 105.57 106.34 105.98 106.085 105.98 106.085 105.65 106.165 105.57 106.34 105.57 ;
      RECT  108.35 103.575 108.17 104.49 ;
      RECT  108.74 103.575 108.53 103.905 ;
      RECT  108.74 103.905 108.53 104.285 ;
      RECT  106.55 107.56 106.34 107.15 ;
      RECT  108.95 108.565 108.74 108.235 ;
      RECT  105.905 107.65 105.83 105.945 ;
      RECT  105.99 107.065 105.905 106.655 ;
      RECT  106.91 108.565 106.73 107.65 ;
      POLYGON  105.905 108.565 105.905 108.235 106.34 108.235 106.34 107.855 105.905 107.855 105.905 107.65 105.83 107.65 105.83 108.565 105.905 108.565 ;
      RECT  105.83 107.65 105.62 105.945 ;
      POLYGON  106.34 107.56 106.34 107.15 106.165 107.15 106.085 107.23 106.085 107.56 106.34 107.56 ;
      RECT  108.95 107.65 108.74 105.945 ;
      RECT  107.27 108.565 107.09 107.65 ;
      RECT  108.35 107.65 108.17 105.945 ;
      RECT  106.55 106.57 106.34 106.16 ;
      RECT  105.83 107.855 105.62 107.65 ;
      RECT  108.74 107.65 108.53 105.945 ;
      RECT  106.55 108.235 106.34 107.855 ;
      RECT  107.99 107.65 107.81 105.945 ;
      RECT  107.27 107.65 107.09 105.945 ;
      RECT  107.99 108.565 107.81 107.65 ;
      RECT  105.83 108.565 105.62 108.235 ;
      RECT  107.63 107.65 107.45 105.945 ;
      RECT  107.63 108.565 107.45 107.65 ;
      RECT  108.95 107.855 108.74 107.65 ;
      RECT  105.83 108.235 105.62 107.855 ;
      RECT  106.91 107.65 106.73 105.945 ;
      RECT  108.74 107.855 108.53 107.65 ;
      RECT  108.95 108.235 108.74 107.855 ;
      POLYGON  106.34 106.57 106.34 106.16 106.085 106.16 106.085 106.49 106.165 106.57 106.34 106.57 ;
      RECT  108.35 108.565 108.17 107.65 ;
      RECT  108.74 108.565 108.53 108.235 ;
      RECT  108.74 108.235 108.53 107.855 ;
      RECT  106.55 108.53 106.34 108.94 ;
      RECT  108.95 107.525 108.74 107.855 ;
      RECT  105.905 108.44 105.83 110.145 ;
      RECT  105.99 109.025 105.905 109.435 ;
      RECT  106.91 107.525 106.73 108.44 ;
      POLYGON  105.905 107.525 105.905 107.855 106.34 107.855 106.34 108.235 105.905 108.235 105.905 108.44 105.83 108.44 105.83 107.525 105.905 107.525 ;
      RECT  105.83 108.44 105.62 110.145 ;
      POLYGON  106.34 108.53 106.34 108.94 106.165 108.94 106.085 108.86 106.085 108.53 106.34 108.53 ;
      RECT  108.95 108.44 108.74 110.145 ;
      RECT  107.27 107.525 107.09 108.44 ;
      RECT  108.35 108.44 108.17 110.145 ;
      RECT  106.55 109.52 106.34 109.93 ;
      RECT  105.83 108.235 105.62 108.44 ;
      RECT  108.74 108.44 108.53 110.145 ;
      RECT  106.55 107.855 106.34 108.235 ;
      RECT  107.99 108.44 107.81 110.145 ;
      RECT  107.27 108.44 107.09 110.145 ;
      RECT  107.99 107.525 107.81 108.44 ;
      RECT  105.83 107.525 105.62 107.855 ;
      RECT  107.63 108.44 107.45 110.145 ;
      RECT  107.63 107.525 107.45 108.44 ;
      RECT  108.95 108.235 108.74 108.44 ;
      RECT  105.83 107.855 105.62 108.235 ;
      RECT  106.91 108.44 106.73 110.145 ;
      RECT  108.74 108.235 108.53 108.44 ;
      RECT  108.95 107.855 108.74 108.235 ;
      POLYGON  106.34 109.52 106.34 109.93 106.085 109.93 106.085 109.6 106.165 109.52 106.34 109.52 ;
      RECT  108.35 107.525 108.17 108.44 ;
      RECT  108.74 107.525 108.53 107.855 ;
      RECT  108.74 107.855 108.53 108.235 ;
      RECT  106.55 111.51 106.34 111.1 ;
      RECT  108.95 112.515 108.74 112.185 ;
      RECT  105.905 111.6 105.83 109.895 ;
      RECT  105.99 111.015 105.905 110.605 ;
      RECT  106.91 112.515 106.73 111.6 ;
      POLYGON  105.905 112.515 105.905 112.185 106.34 112.185 106.34 111.805 105.905 111.805 105.905 111.6 105.83 111.6 105.83 112.515 105.905 112.515 ;
      RECT  105.83 111.6 105.62 109.895 ;
      POLYGON  106.34 111.51 106.34 111.1 106.165 111.1 106.085 111.18 106.085 111.51 106.34 111.51 ;
      RECT  108.95 111.6 108.74 109.895 ;
      RECT  107.27 112.515 107.09 111.6 ;
      RECT  108.35 111.6 108.17 109.895 ;
      RECT  106.55 110.52 106.34 110.11 ;
      RECT  105.83 111.805 105.62 111.6 ;
      RECT  108.74 111.6 108.53 109.895 ;
      RECT  106.55 112.185 106.34 111.805 ;
      RECT  107.99 111.6 107.81 109.895 ;
      RECT  107.27 111.6 107.09 109.895 ;
      RECT  107.99 112.515 107.81 111.6 ;
      RECT  105.83 112.515 105.62 112.185 ;
      RECT  107.63 111.6 107.45 109.895 ;
      RECT  107.63 112.515 107.45 111.6 ;
      RECT  108.95 111.805 108.74 111.6 ;
      RECT  105.83 112.185 105.62 111.805 ;
      RECT  106.91 111.6 106.73 109.895 ;
      RECT  108.74 111.805 108.53 111.6 ;
      RECT  108.95 112.185 108.74 111.805 ;
      POLYGON  106.34 110.52 106.34 110.11 106.085 110.11 106.085 110.44 106.165 110.52 106.34 110.52 ;
      RECT  108.35 112.515 108.17 111.6 ;
      RECT  108.74 112.515 108.53 112.185 ;
      RECT  108.74 112.185 108.53 111.805 ;
      RECT  106.55 112.48 106.34 112.89 ;
      RECT  108.95 111.475 108.74 111.805 ;
      RECT  105.905 112.39 105.83 114.095 ;
      RECT  105.99 112.975 105.905 113.385 ;
      RECT  106.91 111.475 106.73 112.39 ;
      POLYGON  105.905 111.475 105.905 111.805 106.34 111.805 106.34 112.185 105.905 112.185 105.905 112.39 105.83 112.39 105.83 111.475 105.905 111.475 ;
      RECT  105.83 112.39 105.62 114.095 ;
      POLYGON  106.34 112.48 106.34 112.89 106.165 112.89 106.085 112.81 106.085 112.48 106.34 112.48 ;
      RECT  108.95 112.39 108.74 114.095 ;
      RECT  107.27 111.475 107.09 112.39 ;
      RECT  108.35 112.39 108.17 114.095 ;
      RECT  106.55 113.47 106.34 113.88 ;
      RECT  105.83 112.185 105.62 112.39 ;
      RECT  108.74 112.39 108.53 114.095 ;
      RECT  106.55 111.805 106.34 112.185 ;
      RECT  107.99 112.39 107.81 114.095 ;
      RECT  107.27 112.39 107.09 114.095 ;
      RECT  107.99 111.475 107.81 112.39 ;
      RECT  105.83 111.475 105.62 111.805 ;
      RECT  107.63 112.39 107.45 114.095 ;
      RECT  107.63 111.475 107.45 112.39 ;
      RECT  108.95 112.185 108.74 112.39 ;
      RECT  105.83 111.805 105.62 112.185 ;
      RECT  106.91 112.39 106.73 114.095 ;
      RECT  108.74 112.185 108.53 112.39 ;
      RECT  108.95 111.805 108.74 112.185 ;
      POLYGON  106.34 113.47 106.34 113.88 106.085 113.88 106.085 113.55 106.165 113.47 106.34 113.47 ;
      RECT  108.35 111.475 108.17 112.39 ;
      RECT  108.74 111.475 108.53 111.805 ;
      RECT  108.74 111.805 108.53 112.185 ;
      RECT  106.55 115.46 106.34 115.05 ;
      RECT  108.95 116.465 108.74 116.135 ;
      RECT  105.905 115.55 105.83 113.845 ;
      RECT  105.99 114.965 105.905 114.555 ;
      RECT  106.91 116.465 106.73 115.55 ;
      POLYGON  105.905 116.465 105.905 116.135 106.34 116.135 106.34 115.755 105.905 115.755 105.905 115.55 105.83 115.55 105.83 116.465 105.905 116.465 ;
      RECT  105.83 115.55 105.62 113.845 ;
      POLYGON  106.34 115.46 106.34 115.05 106.165 115.05 106.085 115.13 106.085 115.46 106.34 115.46 ;
      RECT  108.95 115.55 108.74 113.845 ;
      RECT  107.27 116.465 107.09 115.55 ;
      RECT  108.35 115.55 108.17 113.845 ;
      RECT  106.55 114.47 106.34 114.06 ;
      RECT  105.83 115.755 105.62 115.55 ;
      RECT  108.74 115.55 108.53 113.845 ;
      RECT  106.55 116.135 106.34 115.755 ;
      RECT  107.99 115.55 107.81 113.845 ;
      RECT  107.27 115.55 107.09 113.845 ;
      RECT  107.99 116.465 107.81 115.55 ;
      RECT  105.83 116.465 105.62 116.135 ;
      RECT  107.63 115.55 107.45 113.845 ;
      RECT  107.63 116.465 107.45 115.55 ;
      RECT  108.95 115.755 108.74 115.55 ;
      RECT  105.83 116.135 105.62 115.755 ;
      RECT  106.91 115.55 106.73 113.845 ;
      RECT  108.74 115.755 108.53 115.55 ;
      RECT  108.95 116.135 108.74 115.755 ;
      POLYGON  106.34 114.47 106.34 114.06 106.085 114.06 106.085 114.39 106.165 114.47 106.34 114.47 ;
      RECT  108.35 116.465 108.17 115.55 ;
      RECT  108.74 116.465 108.53 116.135 ;
      RECT  108.74 116.135 108.53 115.755 ;
      RECT  106.55 116.43 106.34 116.84 ;
      RECT  108.95 115.425 108.74 115.755 ;
      RECT  105.905 116.34 105.83 118.045 ;
      RECT  105.99 116.925 105.905 117.335 ;
      RECT  106.91 115.425 106.73 116.34 ;
      POLYGON  105.905 115.425 105.905 115.755 106.34 115.755 106.34 116.135 105.905 116.135 105.905 116.34 105.83 116.34 105.83 115.425 105.905 115.425 ;
      RECT  105.83 116.34 105.62 118.045 ;
      POLYGON  106.34 116.43 106.34 116.84 106.165 116.84 106.085 116.76 106.085 116.43 106.34 116.43 ;
      RECT  108.95 116.34 108.74 118.045 ;
      RECT  107.27 115.425 107.09 116.34 ;
      RECT  108.35 116.34 108.17 118.045 ;
      RECT  106.55 117.42 106.34 117.83 ;
      RECT  105.83 116.135 105.62 116.34 ;
      RECT  108.74 116.34 108.53 118.045 ;
      RECT  106.55 115.755 106.34 116.135 ;
      RECT  107.99 116.34 107.81 118.045 ;
      RECT  107.27 116.34 107.09 118.045 ;
      RECT  107.99 115.425 107.81 116.34 ;
      RECT  105.83 115.425 105.62 115.755 ;
      RECT  107.63 116.34 107.45 118.045 ;
      RECT  107.63 115.425 107.45 116.34 ;
      RECT  108.95 116.135 108.74 116.34 ;
      RECT  105.83 115.755 105.62 116.135 ;
      RECT  106.91 116.34 106.73 118.045 ;
      RECT  108.74 116.135 108.53 116.34 ;
      RECT  108.95 115.755 108.74 116.135 ;
      POLYGON  106.34 117.42 106.34 117.83 106.085 117.83 106.085 117.5 106.165 117.42 106.34 117.42 ;
      RECT  108.35 115.425 108.17 116.34 ;
      RECT  108.74 115.425 108.53 115.755 ;
      RECT  108.74 115.755 108.53 116.135 ;
      RECT  106.55 119.41 106.34 119.0 ;
      RECT  108.95 120.415 108.74 120.085 ;
      RECT  105.905 119.5 105.83 117.795 ;
      RECT  105.99 118.915 105.905 118.505 ;
      RECT  106.91 120.415 106.73 119.5 ;
      POLYGON  105.905 120.415 105.905 120.085 106.34 120.085 106.34 119.705 105.905 119.705 105.905 119.5 105.83 119.5 105.83 120.415 105.905 120.415 ;
      RECT  105.83 119.5 105.62 117.795 ;
      POLYGON  106.34 119.41 106.34 119.0 106.165 119.0 106.085 119.08 106.085 119.41 106.34 119.41 ;
      RECT  108.95 119.5 108.74 117.795 ;
      RECT  107.27 120.415 107.09 119.5 ;
      RECT  108.35 119.5 108.17 117.795 ;
      RECT  106.55 118.42 106.34 118.01 ;
      RECT  105.83 119.705 105.62 119.5 ;
      RECT  108.74 119.5 108.53 117.795 ;
      RECT  106.55 120.085 106.34 119.705 ;
      RECT  107.99 119.5 107.81 117.795 ;
      RECT  107.27 119.5 107.09 117.795 ;
      RECT  107.99 120.415 107.81 119.5 ;
      RECT  105.83 120.415 105.62 120.085 ;
      RECT  107.63 119.5 107.45 117.795 ;
      RECT  107.63 120.415 107.45 119.5 ;
      RECT  108.95 119.705 108.74 119.5 ;
      RECT  105.83 120.085 105.62 119.705 ;
      RECT  106.91 119.5 106.73 117.795 ;
      RECT  108.74 119.705 108.53 119.5 ;
      RECT  108.95 120.085 108.74 119.705 ;
      POLYGON  106.34 118.42 106.34 118.01 106.085 118.01 106.085 118.34 106.165 118.42 106.34 118.42 ;
      RECT  108.35 120.415 108.17 119.5 ;
      RECT  108.74 120.415 108.53 120.085 ;
      RECT  108.74 120.085 108.53 119.705 ;
      RECT  106.55 120.38 106.34 120.79 ;
      RECT  108.95 119.375 108.74 119.705 ;
      RECT  105.905 120.29 105.83 121.995 ;
      RECT  105.99 120.875 105.905 121.285 ;
      RECT  106.91 119.375 106.73 120.29 ;
      POLYGON  105.905 119.375 105.905 119.705 106.34 119.705 106.34 120.085 105.905 120.085 105.905 120.29 105.83 120.29 105.83 119.375 105.905 119.375 ;
      RECT  105.83 120.29 105.62 121.995 ;
      POLYGON  106.34 120.38 106.34 120.79 106.165 120.79 106.085 120.71 106.085 120.38 106.34 120.38 ;
      RECT  108.95 120.29 108.74 121.995 ;
      RECT  107.27 119.375 107.09 120.29 ;
      RECT  108.35 120.29 108.17 121.995 ;
      RECT  106.55 121.37 106.34 121.78 ;
      RECT  105.83 120.085 105.62 120.29 ;
      RECT  108.74 120.29 108.53 121.995 ;
      RECT  106.55 119.705 106.34 120.085 ;
      RECT  107.99 120.29 107.81 121.995 ;
      RECT  107.27 120.29 107.09 121.995 ;
      RECT  107.99 119.375 107.81 120.29 ;
      RECT  105.83 119.375 105.62 119.705 ;
      RECT  107.63 120.29 107.45 121.995 ;
      RECT  107.63 119.375 107.45 120.29 ;
      RECT  108.95 120.085 108.74 120.29 ;
      RECT  105.83 119.705 105.62 120.085 ;
      RECT  106.91 120.29 106.73 121.995 ;
      RECT  108.74 120.085 108.53 120.29 ;
      RECT  108.95 119.705 108.74 120.085 ;
      POLYGON  106.34 121.37 106.34 121.78 106.085 121.78 106.085 121.45 106.165 121.37 106.34 121.37 ;
      RECT  108.35 119.375 108.17 120.29 ;
      RECT  108.74 119.375 108.53 119.705 ;
      RECT  108.74 119.705 108.53 120.085 ;
      RECT  106.55 123.36 106.34 122.95 ;
      RECT  108.95 124.365 108.74 124.035 ;
      RECT  105.905 123.45 105.83 121.745 ;
      RECT  105.99 122.865 105.905 122.455 ;
      RECT  106.91 124.365 106.73 123.45 ;
      POLYGON  105.905 124.365 105.905 124.035 106.34 124.035 106.34 123.655 105.905 123.655 105.905 123.45 105.83 123.45 105.83 124.365 105.905 124.365 ;
      RECT  105.83 123.45 105.62 121.745 ;
      POLYGON  106.34 123.36 106.34 122.95 106.165 122.95 106.085 123.03 106.085 123.36 106.34 123.36 ;
      RECT  108.95 123.45 108.74 121.745 ;
      RECT  107.27 124.365 107.09 123.45 ;
      RECT  108.35 123.45 108.17 121.745 ;
      RECT  106.55 122.37 106.34 121.96 ;
      RECT  105.83 123.655 105.62 123.45 ;
      RECT  108.74 123.45 108.53 121.745 ;
      RECT  106.55 124.035 106.34 123.655 ;
      RECT  107.99 123.45 107.81 121.745 ;
      RECT  107.27 123.45 107.09 121.745 ;
      RECT  107.99 124.365 107.81 123.45 ;
      RECT  105.83 124.365 105.62 124.035 ;
      RECT  107.63 123.45 107.45 121.745 ;
      RECT  107.63 124.365 107.45 123.45 ;
      RECT  108.95 123.655 108.74 123.45 ;
      RECT  105.83 124.035 105.62 123.655 ;
      RECT  106.91 123.45 106.73 121.745 ;
      RECT  108.74 123.655 108.53 123.45 ;
      RECT  108.95 124.035 108.74 123.655 ;
      POLYGON  106.34 122.37 106.34 121.96 106.085 121.96 106.085 122.29 106.165 122.37 106.34 122.37 ;
      RECT  108.35 124.365 108.17 123.45 ;
      RECT  108.74 124.365 108.53 124.035 ;
      RECT  108.74 124.035 108.53 123.655 ;
      RECT  110.93 92.73 111.14 93.14 ;
      RECT  108.53 91.725 108.74 92.055 ;
      RECT  111.575 92.64 111.65 94.345 ;
      RECT  111.49 93.225 111.575 93.635 ;
      RECT  110.57 91.725 110.75 92.64 ;
      POLYGON  111.575 91.725 111.575 92.055 111.14 92.055 111.14 92.435 111.575 92.435 111.575 92.64 111.65 92.64 111.65 91.725 111.575 91.725 ;
      RECT  111.65 92.64 111.86 94.345 ;
      POLYGON  111.14 92.73 111.14 93.14 111.315 93.14 111.395 93.06 111.395 92.73 111.14 92.73 ;
      RECT  108.53 92.64 108.74 94.345 ;
      RECT  110.21 91.725 110.39 92.64 ;
      RECT  109.13 92.64 109.31 94.345 ;
      RECT  110.93 93.72 111.14 94.13 ;
      RECT  111.65 92.435 111.86 92.64 ;
      RECT  108.74 92.64 108.95 94.345 ;
      RECT  110.93 92.055 111.14 92.435 ;
      RECT  109.49 92.64 109.67 94.345 ;
      RECT  110.21 92.64 110.39 94.345 ;
      RECT  109.49 91.725 109.67 92.64 ;
      RECT  111.65 91.725 111.86 92.055 ;
      RECT  109.85 92.64 110.03 94.345 ;
      RECT  109.85 91.725 110.03 92.64 ;
      RECT  108.53 92.435 108.74 92.64 ;
      RECT  111.65 92.055 111.86 92.435 ;
      RECT  110.57 92.64 110.75 94.345 ;
      RECT  108.74 92.435 108.95 92.64 ;
      RECT  108.53 92.055 108.74 92.435 ;
      POLYGON  111.14 93.72 111.14 94.13 111.395 94.13 111.395 93.8 111.315 93.72 111.14 93.72 ;
      RECT  109.13 91.725 109.31 92.64 ;
      RECT  108.74 91.725 108.95 92.055 ;
      RECT  108.74 92.055 108.95 92.435 ;
      RECT  110.93 95.71 111.14 95.3 ;
      RECT  108.53 96.715 108.74 96.385 ;
      RECT  111.575 95.8 111.65 94.095 ;
      RECT  111.49 95.215 111.575 94.805 ;
      RECT  110.57 96.715 110.75 95.8 ;
      POLYGON  111.575 96.715 111.575 96.385 111.14 96.385 111.14 96.005 111.575 96.005 111.575 95.8 111.65 95.8 111.65 96.715 111.575 96.715 ;
      RECT  111.65 95.8 111.86 94.095 ;
      POLYGON  111.14 95.71 111.14 95.3 111.315 95.3 111.395 95.38 111.395 95.71 111.14 95.71 ;
      RECT  108.53 95.8 108.74 94.095 ;
      RECT  110.21 96.715 110.39 95.8 ;
      RECT  109.13 95.8 109.31 94.095 ;
      RECT  110.93 94.72 111.14 94.31 ;
      RECT  111.65 96.005 111.86 95.8 ;
      RECT  108.74 95.8 108.95 94.095 ;
      RECT  110.93 96.385 111.14 96.005 ;
      RECT  109.49 95.8 109.67 94.095 ;
      RECT  110.21 95.8 110.39 94.095 ;
      RECT  109.49 96.715 109.67 95.8 ;
      RECT  111.65 96.715 111.86 96.385 ;
      RECT  109.85 95.8 110.03 94.095 ;
      RECT  109.85 96.715 110.03 95.8 ;
      RECT  108.53 96.005 108.74 95.8 ;
      RECT  111.65 96.385 111.86 96.005 ;
      RECT  110.57 95.8 110.75 94.095 ;
      RECT  108.74 96.005 108.95 95.8 ;
      RECT  108.53 96.385 108.74 96.005 ;
      POLYGON  111.14 94.72 111.14 94.31 111.395 94.31 111.395 94.64 111.315 94.72 111.14 94.72 ;
      RECT  109.13 96.715 109.31 95.8 ;
      RECT  108.74 96.715 108.95 96.385 ;
      RECT  108.74 96.385 108.95 96.005 ;
      RECT  110.93 96.68 111.14 97.09 ;
      RECT  108.53 95.675 108.74 96.005 ;
      RECT  111.575 96.59 111.65 98.295 ;
      RECT  111.49 97.175 111.575 97.585 ;
      RECT  110.57 95.675 110.75 96.59 ;
      POLYGON  111.575 95.675 111.575 96.005 111.14 96.005 111.14 96.385 111.575 96.385 111.575 96.59 111.65 96.59 111.65 95.675 111.575 95.675 ;
      RECT  111.65 96.59 111.86 98.295 ;
      POLYGON  111.14 96.68 111.14 97.09 111.315 97.09 111.395 97.01 111.395 96.68 111.14 96.68 ;
      RECT  108.53 96.59 108.74 98.295 ;
      RECT  110.21 95.675 110.39 96.59 ;
      RECT  109.13 96.59 109.31 98.295 ;
      RECT  110.93 97.67 111.14 98.08 ;
      RECT  111.65 96.385 111.86 96.59 ;
      RECT  108.74 96.59 108.95 98.295 ;
      RECT  110.93 96.005 111.14 96.385 ;
      RECT  109.49 96.59 109.67 98.295 ;
      RECT  110.21 96.59 110.39 98.295 ;
      RECT  109.49 95.675 109.67 96.59 ;
      RECT  111.65 95.675 111.86 96.005 ;
      RECT  109.85 96.59 110.03 98.295 ;
      RECT  109.85 95.675 110.03 96.59 ;
      RECT  108.53 96.385 108.74 96.59 ;
      RECT  111.65 96.005 111.86 96.385 ;
      RECT  110.57 96.59 110.75 98.295 ;
      RECT  108.74 96.385 108.95 96.59 ;
      RECT  108.53 96.005 108.74 96.385 ;
      POLYGON  111.14 97.67 111.14 98.08 111.395 98.08 111.395 97.75 111.315 97.67 111.14 97.67 ;
      RECT  109.13 95.675 109.31 96.59 ;
      RECT  108.74 95.675 108.95 96.005 ;
      RECT  108.74 96.005 108.95 96.385 ;
      RECT  110.93 99.66 111.14 99.25 ;
      RECT  108.53 100.665 108.74 100.335 ;
      RECT  111.575 99.75 111.65 98.045 ;
      RECT  111.49 99.165 111.575 98.755 ;
      RECT  110.57 100.665 110.75 99.75 ;
      POLYGON  111.575 100.665 111.575 100.335 111.14 100.335 111.14 99.955 111.575 99.955 111.575 99.75 111.65 99.75 111.65 100.665 111.575 100.665 ;
      RECT  111.65 99.75 111.86 98.045 ;
      POLYGON  111.14 99.66 111.14 99.25 111.315 99.25 111.395 99.33 111.395 99.66 111.14 99.66 ;
      RECT  108.53 99.75 108.74 98.045 ;
      RECT  110.21 100.665 110.39 99.75 ;
      RECT  109.13 99.75 109.31 98.045 ;
      RECT  110.93 98.67 111.14 98.26 ;
      RECT  111.65 99.955 111.86 99.75 ;
      RECT  108.74 99.75 108.95 98.045 ;
      RECT  110.93 100.335 111.14 99.955 ;
      RECT  109.49 99.75 109.67 98.045 ;
      RECT  110.21 99.75 110.39 98.045 ;
      RECT  109.49 100.665 109.67 99.75 ;
      RECT  111.65 100.665 111.86 100.335 ;
      RECT  109.85 99.75 110.03 98.045 ;
      RECT  109.85 100.665 110.03 99.75 ;
      RECT  108.53 99.955 108.74 99.75 ;
      RECT  111.65 100.335 111.86 99.955 ;
      RECT  110.57 99.75 110.75 98.045 ;
      RECT  108.74 99.955 108.95 99.75 ;
      RECT  108.53 100.335 108.74 99.955 ;
      POLYGON  111.14 98.67 111.14 98.26 111.395 98.26 111.395 98.59 111.315 98.67 111.14 98.67 ;
      RECT  109.13 100.665 109.31 99.75 ;
      RECT  108.74 100.665 108.95 100.335 ;
      RECT  108.74 100.335 108.95 99.955 ;
      RECT  110.93 100.63 111.14 101.04 ;
      RECT  108.53 99.625 108.74 99.955 ;
      RECT  111.575 100.54 111.65 102.245 ;
      RECT  111.49 101.125 111.575 101.535 ;
      RECT  110.57 99.625 110.75 100.54 ;
      POLYGON  111.575 99.625 111.575 99.955 111.14 99.955 111.14 100.335 111.575 100.335 111.575 100.54 111.65 100.54 111.65 99.625 111.575 99.625 ;
      RECT  111.65 100.54 111.86 102.245 ;
      POLYGON  111.14 100.63 111.14 101.04 111.315 101.04 111.395 100.96 111.395 100.63 111.14 100.63 ;
      RECT  108.53 100.54 108.74 102.245 ;
      RECT  110.21 99.625 110.39 100.54 ;
      RECT  109.13 100.54 109.31 102.245 ;
      RECT  110.93 101.62 111.14 102.03 ;
      RECT  111.65 100.335 111.86 100.54 ;
      RECT  108.74 100.54 108.95 102.245 ;
      RECT  110.93 99.955 111.14 100.335 ;
      RECT  109.49 100.54 109.67 102.245 ;
      RECT  110.21 100.54 110.39 102.245 ;
      RECT  109.49 99.625 109.67 100.54 ;
      RECT  111.65 99.625 111.86 99.955 ;
      RECT  109.85 100.54 110.03 102.245 ;
      RECT  109.85 99.625 110.03 100.54 ;
      RECT  108.53 100.335 108.74 100.54 ;
      RECT  111.65 99.955 111.86 100.335 ;
      RECT  110.57 100.54 110.75 102.245 ;
      RECT  108.74 100.335 108.95 100.54 ;
      RECT  108.53 99.955 108.74 100.335 ;
      POLYGON  111.14 101.62 111.14 102.03 111.395 102.03 111.395 101.7 111.315 101.62 111.14 101.62 ;
      RECT  109.13 99.625 109.31 100.54 ;
      RECT  108.74 99.625 108.95 99.955 ;
      RECT  108.74 99.955 108.95 100.335 ;
      RECT  110.93 103.61 111.14 103.2 ;
      RECT  108.53 104.615 108.74 104.285 ;
      RECT  111.575 103.7 111.65 101.995 ;
      RECT  111.49 103.115 111.575 102.705 ;
      RECT  110.57 104.615 110.75 103.7 ;
      POLYGON  111.575 104.615 111.575 104.285 111.14 104.285 111.14 103.905 111.575 103.905 111.575 103.7 111.65 103.7 111.65 104.615 111.575 104.615 ;
      RECT  111.65 103.7 111.86 101.995 ;
      POLYGON  111.14 103.61 111.14 103.2 111.315 103.2 111.395 103.28 111.395 103.61 111.14 103.61 ;
      RECT  108.53 103.7 108.74 101.995 ;
      RECT  110.21 104.615 110.39 103.7 ;
      RECT  109.13 103.7 109.31 101.995 ;
      RECT  110.93 102.62 111.14 102.21 ;
      RECT  111.65 103.905 111.86 103.7 ;
      RECT  108.74 103.7 108.95 101.995 ;
      RECT  110.93 104.285 111.14 103.905 ;
      RECT  109.49 103.7 109.67 101.995 ;
      RECT  110.21 103.7 110.39 101.995 ;
      RECT  109.49 104.615 109.67 103.7 ;
      RECT  111.65 104.615 111.86 104.285 ;
      RECT  109.85 103.7 110.03 101.995 ;
      RECT  109.85 104.615 110.03 103.7 ;
      RECT  108.53 103.905 108.74 103.7 ;
      RECT  111.65 104.285 111.86 103.905 ;
      RECT  110.57 103.7 110.75 101.995 ;
      RECT  108.74 103.905 108.95 103.7 ;
      RECT  108.53 104.285 108.74 103.905 ;
      POLYGON  111.14 102.62 111.14 102.21 111.395 102.21 111.395 102.54 111.315 102.62 111.14 102.62 ;
      RECT  109.13 104.615 109.31 103.7 ;
      RECT  108.74 104.615 108.95 104.285 ;
      RECT  108.74 104.285 108.95 103.905 ;
      RECT  110.93 104.58 111.14 104.99 ;
      RECT  108.53 103.575 108.74 103.905 ;
      RECT  111.575 104.49 111.65 106.195 ;
      RECT  111.49 105.075 111.575 105.485 ;
      RECT  110.57 103.575 110.75 104.49 ;
      POLYGON  111.575 103.575 111.575 103.905 111.14 103.905 111.14 104.285 111.575 104.285 111.575 104.49 111.65 104.49 111.65 103.575 111.575 103.575 ;
      RECT  111.65 104.49 111.86 106.195 ;
      POLYGON  111.14 104.58 111.14 104.99 111.315 104.99 111.395 104.91 111.395 104.58 111.14 104.58 ;
      RECT  108.53 104.49 108.74 106.195 ;
      RECT  110.21 103.575 110.39 104.49 ;
      RECT  109.13 104.49 109.31 106.195 ;
      RECT  110.93 105.57 111.14 105.98 ;
      RECT  111.65 104.285 111.86 104.49 ;
      RECT  108.74 104.49 108.95 106.195 ;
      RECT  110.93 103.905 111.14 104.285 ;
      RECT  109.49 104.49 109.67 106.195 ;
      RECT  110.21 104.49 110.39 106.195 ;
      RECT  109.49 103.575 109.67 104.49 ;
      RECT  111.65 103.575 111.86 103.905 ;
      RECT  109.85 104.49 110.03 106.195 ;
      RECT  109.85 103.575 110.03 104.49 ;
      RECT  108.53 104.285 108.74 104.49 ;
      RECT  111.65 103.905 111.86 104.285 ;
      RECT  110.57 104.49 110.75 106.195 ;
      RECT  108.74 104.285 108.95 104.49 ;
      RECT  108.53 103.905 108.74 104.285 ;
      POLYGON  111.14 105.57 111.14 105.98 111.395 105.98 111.395 105.65 111.315 105.57 111.14 105.57 ;
      RECT  109.13 103.575 109.31 104.49 ;
      RECT  108.74 103.575 108.95 103.905 ;
      RECT  108.74 103.905 108.95 104.285 ;
      RECT  110.93 107.56 111.14 107.15 ;
      RECT  108.53 108.565 108.74 108.235 ;
      RECT  111.575 107.65 111.65 105.945 ;
      RECT  111.49 107.065 111.575 106.655 ;
      RECT  110.57 108.565 110.75 107.65 ;
      POLYGON  111.575 108.565 111.575 108.235 111.14 108.235 111.14 107.855 111.575 107.855 111.575 107.65 111.65 107.65 111.65 108.565 111.575 108.565 ;
      RECT  111.65 107.65 111.86 105.945 ;
      POLYGON  111.14 107.56 111.14 107.15 111.315 107.15 111.395 107.23 111.395 107.56 111.14 107.56 ;
      RECT  108.53 107.65 108.74 105.945 ;
      RECT  110.21 108.565 110.39 107.65 ;
      RECT  109.13 107.65 109.31 105.945 ;
      RECT  110.93 106.57 111.14 106.16 ;
      RECT  111.65 107.855 111.86 107.65 ;
      RECT  108.74 107.65 108.95 105.945 ;
      RECT  110.93 108.235 111.14 107.855 ;
      RECT  109.49 107.65 109.67 105.945 ;
      RECT  110.21 107.65 110.39 105.945 ;
      RECT  109.49 108.565 109.67 107.65 ;
      RECT  111.65 108.565 111.86 108.235 ;
      RECT  109.85 107.65 110.03 105.945 ;
      RECT  109.85 108.565 110.03 107.65 ;
      RECT  108.53 107.855 108.74 107.65 ;
      RECT  111.65 108.235 111.86 107.855 ;
      RECT  110.57 107.65 110.75 105.945 ;
      RECT  108.74 107.855 108.95 107.65 ;
      RECT  108.53 108.235 108.74 107.855 ;
      POLYGON  111.14 106.57 111.14 106.16 111.395 106.16 111.395 106.49 111.315 106.57 111.14 106.57 ;
      RECT  109.13 108.565 109.31 107.65 ;
      RECT  108.74 108.565 108.95 108.235 ;
      RECT  108.74 108.235 108.95 107.855 ;
      RECT  110.93 108.53 111.14 108.94 ;
      RECT  108.53 107.525 108.74 107.855 ;
      RECT  111.575 108.44 111.65 110.145 ;
      RECT  111.49 109.025 111.575 109.435 ;
      RECT  110.57 107.525 110.75 108.44 ;
      POLYGON  111.575 107.525 111.575 107.855 111.14 107.855 111.14 108.235 111.575 108.235 111.575 108.44 111.65 108.44 111.65 107.525 111.575 107.525 ;
      RECT  111.65 108.44 111.86 110.145 ;
      POLYGON  111.14 108.53 111.14 108.94 111.315 108.94 111.395 108.86 111.395 108.53 111.14 108.53 ;
      RECT  108.53 108.44 108.74 110.145 ;
      RECT  110.21 107.525 110.39 108.44 ;
      RECT  109.13 108.44 109.31 110.145 ;
      RECT  110.93 109.52 111.14 109.93 ;
      RECT  111.65 108.235 111.86 108.44 ;
      RECT  108.74 108.44 108.95 110.145 ;
      RECT  110.93 107.855 111.14 108.235 ;
      RECT  109.49 108.44 109.67 110.145 ;
      RECT  110.21 108.44 110.39 110.145 ;
      RECT  109.49 107.525 109.67 108.44 ;
      RECT  111.65 107.525 111.86 107.855 ;
      RECT  109.85 108.44 110.03 110.145 ;
      RECT  109.85 107.525 110.03 108.44 ;
      RECT  108.53 108.235 108.74 108.44 ;
      RECT  111.65 107.855 111.86 108.235 ;
      RECT  110.57 108.44 110.75 110.145 ;
      RECT  108.74 108.235 108.95 108.44 ;
      RECT  108.53 107.855 108.74 108.235 ;
      POLYGON  111.14 109.52 111.14 109.93 111.395 109.93 111.395 109.6 111.315 109.52 111.14 109.52 ;
      RECT  109.13 107.525 109.31 108.44 ;
      RECT  108.74 107.525 108.95 107.855 ;
      RECT  108.74 107.855 108.95 108.235 ;
      RECT  110.93 111.51 111.14 111.1 ;
      RECT  108.53 112.515 108.74 112.185 ;
      RECT  111.575 111.6 111.65 109.895 ;
      RECT  111.49 111.015 111.575 110.605 ;
      RECT  110.57 112.515 110.75 111.6 ;
      POLYGON  111.575 112.515 111.575 112.185 111.14 112.185 111.14 111.805 111.575 111.805 111.575 111.6 111.65 111.6 111.65 112.515 111.575 112.515 ;
      RECT  111.65 111.6 111.86 109.895 ;
      POLYGON  111.14 111.51 111.14 111.1 111.315 111.1 111.395 111.18 111.395 111.51 111.14 111.51 ;
      RECT  108.53 111.6 108.74 109.895 ;
      RECT  110.21 112.515 110.39 111.6 ;
      RECT  109.13 111.6 109.31 109.895 ;
      RECT  110.93 110.52 111.14 110.11 ;
      RECT  111.65 111.805 111.86 111.6 ;
      RECT  108.74 111.6 108.95 109.895 ;
      RECT  110.93 112.185 111.14 111.805 ;
      RECT  109.49 111.6 109.67 109.895 ;
      RECT  110.21 111.6 110.39 109.895 ;
      RECT  109.49 112.515 109.67 111.6 ;
      RECT  111.65 112.515 111.86 112.185 ;
      RECT  109.85 111.6 110.03 109.895 ;
      RECT  109.85 112.515 110.03 111.6 ;
      RECT  108.53 111.805 108.74 111.6 ;
      RECT  111.65 112.185 111.86 111.805 ;
      RECT  110.57 111.6 110.75 109.895 ;
      RECT  108.74 111.805 108.95 111.6 ;
      RECT  108.53 112.185 108.74 111.805 ;
      POLYGON  111.14 110.52 111.14 110.11 111.395 110.11 111.395 110.44 111.315 110.52 111.14 110.52 ;
      RECT  109.13 112.515 109.31 111.6 ;
      RECT  108.74 112.515 108.95 112.185 ;
      RECT  108.74 112.185 108.95 111.805 ;
      RECT  110.93 112.48 111.14 112.89 ;
      RECT  108.53 111.475 108.74 111.805 ;
      RECT  111.575 112.39 111.65 114.095 ;
      RECT  111.49 112.975 111.575 113.385 ;
      RECT  110.57 111.475 110.75 112.39 ;
      POLYGON  111.575 111.475 111.575 111.805 111.14 111.805 111.14 112.185 111.575 112.185 111.575 112.39 111.65 112.39 111.65 111.475 111.575 111.475 ;
      RECT  111.65 112.39 111.86 114.095 ;
      POLYGON  111.14 112.48 111.14 112.89 111.315 112.89 111.395 112.81 111.395 112.48 111.14 112.48 ;
      RECT  108.53 112.39 108.74 114.095 ;
      RECT  110.21 111.475 110.39 112.39 ;
      RECT  109.13 112.39 109.31 114.095 ;
      RECT  110.93 113.47 111.14 113.88 ;
      RECT  111.65 112.185 111.86 112.39 ;
      RECT  108.74 112.39 108.95 114.095 ;
      RECT  110.93 111.805 111.14 112.185 ;
      RECT  109.49 112.39 109.67 114.095 ;
      RECT  110.21 112.39 110.39 114.095 ;
      RECT  109.49 111.475 109.67 112.39 ;
      RECT  111.65 111.475 111.86 111.805 ;
      RECT  109.85 112.39 110.03 114.095 ;
      RECT  109.85 111.475 110.03 112.39 ;
      RECT  108.53 112.185 108.74 112.39 ;
      RECT  111.65 111.805 111.86 112.185 ;
      RECT  110.57 112.39 110.75 114.095 ;
      RECT  108.74 112.185 108.95 112.39 ;
      RECT  108.53 111.805 108.74 112.185 ;
      POLYGON  111.14 113.47 111.14 113.88 111.395 113.88 111.395 113.55 111.315 113.47 111.14 113.47 ;
      RECT  109.13 111.475 109.31 112.39 ;
      RECT  108.74 111.475 108.95 111.805 ;
      RECT  108.74 111.805 108.95 112.185 ;
      RECT  110.93 115.46 111.14 115.05 ;
      RECT  108.53 116.465 108.74 116.135 ;
      RECT  111.575 115.55 111.65 113.845 ;
      RECT  111.49 114.965 111.575 114.555 ;
      RECT  110.57 116.465 110.75 115.55 ;
      POLYGON  111.575 116.465 111.575 116.135 111.14 116.135 111.14 115.755 111.575 115.755 111.575 115.55 111.65 115.55 111.65 116.465 111.575 116.465 ;
      RECT  111.65 115.55 111.86 113.845 ;
      POLYGON  111.14 115.46 111.14 115.05 111.315 115.05 111.395 115.13 111.395 115.46 111.14 115.46 ;
      RECT  108.53 115.55 108.74 113.845 ;
      RECT  110.21 116.465 110.39 115.55 ;
      RECT  109.13 115.55 109.31 113.845 ;
      RECT  110.93 114.47 111.14 114.06 ;
      RECT  111.65 115.755 111.86 115.55 ;
      RECT  108.74 115.55 108.95 113.845 ;
      RECT  110.93 116.135 111.14 115.755 ;
      RECT  109.49 115.55 109.67 113.845 ;
      RECT  110.21 115.55 110.39 113.845 ;
      RECT  109.49 116.465 109.67 115.55 ;
      RECT  111.65 116.465 111.86 116.135 ;
      RECT  109.85 115.55 110.03 113.845 ;
      RECT  109.85 116.465 110.03 115.55 ;
      RECT  108.53 115.755 108.74 115.55 ;
      RECT  111.65 116.135 111.86 115.755 ;
      RECT  110.57 115.55 110.75 113.845 ;
      RECT  108.74 115.755 108.95 115.55 ;
      RECT  108.53 116.135 108.74 115.755 ;
      POLYGON  111.14 114.47 111.14 114.06 111.395 114.06 111.395 114.39 111.315 114.47 111.14 114.47 ;
      RECT  109.13 116.465 109.31 115.55 ;
      RECT  108.74 116.465 108.95 116.135 ;
      RECT  108.74 116.135 108.95 115.755 ;
      RECT  110.93 116.43 111.14 116.84 ;
      RECT  108.53 115.425 108.74 115.755 ;
      RECT  111.575 116.34 111.65 118.045 ;
      RECT  111.49 116.925 111.575 117.335 ;
      RECT  110.57 115.425 110.75 116.34 ;
      POLYGON  111.575 115.425 111.575 115.755 111.14 115.755 111.14 116.135 111.575 116.135 111.575 116.34 111.65 116.34 111.65 115.425 111.575 115.425 ;
      RECT  111.65 116.34 111.86 118.045 ;
      POLYGON  111.14 116.43 111.14 116.84 111.315 116.84 111.395 116.76 111.395 116.43 111.14 116.43 ;
      RECT  108.53 116.34 108.74 118.045 ;
      RECT  110.21 115.425 110.39 116.34 ;
      RECT  109.13 116.34 109.31 118.045 ;
      RECT  110.93 117.42 111.14 117.83 ;
      RECT  111.65 116.135 111.86 116.34 ;
      RECT  108.74 116.34 108.95 118.045 ;
      RECT  110.93 115.755 111.14 116.135 ;
      RECT  109.49 116.34 109.67 118.045 ;
      RECT  110.21 116.34 110.39 118.045 ;
      RECT  109.49 115.425 109.67 116.34 ;
      RECT  111.65 115.425 111.86 115.755 ;
      RECT  109.85 116.34 110.03 118.045 ;
      RECT  109.85 115.425 110.03 116.34 ;
      RECT  108.53 116.135 108.74 116.34 ;
      RECT  111.65 115.755 111.86 116.135 ;
      RECT  110.57 116.34 110.75 118.045 ;
      RECT  108.74 116.135 108.95 116.34 ;
      RECT  108.53 115.755 108.74 116.135 ;
      POLYGON  111.14 117.42 111.14 117.83 111.395 117.83 111.395 117.5 111.315 117.42 111.14 117.42 ;
      RECT  109.13 115.425 109.31 116.34 ;
      RECT  108.74 115.425 108.95 115.755 ;
      RECT  108.74 115.755 108.95 116.135 ;
      RECT  110.93 119.41 111.14 119.0 ;
      RECT  108.53 120.415 108.74 120.085 ;
      RECT  111.575 119.5 111.65 117.795 ;
      RECT  111.49 118.915 111.575 118.505 ;
      RECT  110.57 120.415 110.75 119.5 ;
      POLYGON  111.575 120.415 111.575 120.085 111.14 120.085 111.14 119.705 111.575 119.705 111.575 119.5 111.65 119.5 111.65 120.415 111.575 120.415 ;
      RECT  111.65 119.5 111.86 117.795 ;
      POLYGON  111.14 119.41 111.14 119.0 111.315 119.0 111.395 119.08 111.395 119.41 111.14 119.41 ;
      RECT  108.53 119.5 108.74 117.795 ;
      RECT  110.21 120.415 110.39 119.5 ;
      RECT  109.13 119.5 109.31 117.795 ;
      RECT  110.93 118.42 111.14 118.01 ;
      RECT  111.65 119.705 111.86 119.5 ;
      RECT  108.74 119.5 108.95 117.795 ;
      RECT  110.93 120.085 111.14 119.705 ;
      RECT  109.49 119.5 109.67 117.795 ;
      RECT  110.21 119.5 110.39 117.795 ;
      RECT  109.49 120.415 109.67 119.5 ;
      RECT  111.65 120.415 111.86 120.085 ;
      RECT  109.85 119.5 110.03 117.795 ;
      RECT  109.85 120.415 110.03 119.5 ;
      RECT  108.53 119.705 108.74 119.5 ;
      RECT  111.65 120.085 111.86 119.705 ;
      RECT  110.57 119.5 110.75 117.795 ;
      RECT  108.74 119.705 108.95 119.5 ;
      RECT  108.53 120.085 108.74 119.705 ;
      POLYGON  111.14 118.42 111.14 118.01 111.395 118.01 111.395 118.34 111.315 118.42 111.14 118.42 ;
      RECT  109.13 120.415 109.31 119.5 ;
      RECT  108.74 120.415 108.95 120.085 ;
      RECT  108.74 120.085 108.95 119.705 ;
      RECT  110.93 120.38 111.14 120.79 ;
      RECT  108.53 119.375 108.74 119.705 ;
      RECT  111.575 120.29 111.65 121.995 ;
      RECT  111.49 120.875 111.575 121.285 ;
      RECT  110.57 119.375 110.75 120.29 ;
      POLYGON  111.575 119.375 111.575 119.705 111.14 119.705 111.14 120.085 111.575 120.085 111.575 120.29 111.65 120.29 111.65 119.375 111.575 119.375 ;
      RECT  111.65 120.29 111.86 121.995 ;
      POLYGON  111.14 120.38 111.14 120.79 111.315 120.79 111.395 120.71 111.395 120.38 111.14 120.38 ;
      RECT  108.53 120.29 108.74 121.995 ;
      RECT  110.21 119.375 110.39 120.29 ;
      RECT  109.13 120.29 109.31 121.995 ;
      RECT  110.93 121.37 111.14 121.78 ;
      RECT  111.65 120.085 111.86 120.29 ;
      RECT  108.74 120.29 108.95 121.995 ;
      RECT  110.93 119.705 111.14 120.085 ;
      RECT  109.49 120.29 109.67 121.995 ;
      RECT  110.21 120.29 110.39 121.995 ;
      RECT  109.49 119.375 109.67 120.29 ;
      RECT  111.65 119.375 111.86 119.705 ;
      RECT  109.85 120.29 110.03 121.995 ;
      RECT  109.85 119.375 110.03 120.29 ;
      RECT  108.53 120.085 108.74 120.29 ;
      RECT  111.65 119.705 111.86 120.085 ;
      RECT  110.57 120.29 110.75 121.995 ;
      RECT  108.74 120.085 108.95 120.29 ;
      RECT  108.53 119.705 108.74 120.085 ;
      POLYGON  111.14 121.37 111.14 121.78 111.395 121.78 111.395 121.45 111.315 121.37 111.14 121.37 ;
      RECT  109.13 119.375 109.31 120.29 ;
      RECT  108.74 119.375 108.95 119.705 ;
      RECT  108.74 119.705 108.95 120.085 ;
      RECT  110.93 123.36 111.14 122.95 ;
      RECT  108.53 124.365 108.74 124.035 ;
      RECT  111.575 123.45 111.65 121.745 ;
      RECT  111.49 122.865 111.575 122.455 ;
      RECT  110.57 124.365 110.75 123.45 ;
      POLYGON  111.575 124.365 111.575 124.035 111.14 124.035 111.14 123.655 111.575 123.655 111.575 123.45 111.65 123.45 111.65 124.365 111.575 124.365 ;
      RECT  111.65 123.45 111.86 121.745 ;
      POLYGON  111.14 123.36 111.14 122.95 111.315 122.95 111.395 123.03 111.395 123.36 111.14 123.36 ;
      RECT  108.53 123.45 108.74 121.745 ;
      RECT  110.21 124.365 110.39 123.45 ;
      RECT  109.13 123.45 109.31 121.745 ;
      RECT  110.93 122.37 111.14 121.96 ;
      RECT  111.65 123.655 111.86 123.45 ;
      RECT  108.74 123.45 108.95 121.745 ;
      RECT  110.93 124.035 111.14 123.655 ;
      RECT  109.49 123.45 109.67 121.745 ;
      RECT  110.21 123.45 110.39 121.745 ;
      RECT  109.49 124.365 109.67 123.45 ;
      RECT  111.65 124.365 111.86 124.035 ;
      RECT  109.85 123.45 110.03 121.745 ;
      RECT  109.85 124.365 110.03 123.45 ;
      RECT  108.53 123.655 108.74 123.45 ;
      RECT  111.65 124.035 111.86 123.655 ;
      RECT  110.57 123.45 110.75 121.745 ;
      RECT  108.74 123.655 108.95 123.45 ;
      RECT  108.53 124.035 108.74 123.655 ;
      POLYGON  111.14 122.37 111.14 121.96 111.395 121.96 111.395 122.29 111.315 122.37 111.14 122.37 ;
      RECT  109.13 124.365 109.31 123.45 ;
      RECT  108.74 124.365 108.95 124.035 ;
      RECT  108.74 124.035 108.95 123.655 ;
      RECT  112.79 92.73 112.58 93.14 ;
      RECT  115.19 91.725 114.98 92.055 ;
      RECT  112.145 92.64 112.07 94.345 ;
      RECT  112.23 93.225 112.145 93.635 ;
      RECT  113.15 91.725 112.97 92.64 ;
      POLYGON  112.145 91.725 112.145 92.055 112.58 92.055 112.58 92.435 112.145 92.435 112.145 92.64 112.07 92.64 112.07 91.725 112.145 91.725 ;
      RECT  112.07 92.64 111.86 94.345 ;
      POLYGON  112.58 92.73 112.58 93.14 112.405 93.14 112.325 93.06 112.325 92.73 112.58 92.73 ;
      RECT  115.19 92.64 114.98 94.345 ;
      RECT  113.51 91.725 113.33 92.64 ;
      RECT  114.59 92.64 114.41 94.345 ;
      RECT  112.79 93.72 112.58 94.13 ;
      RECT  112.07 92.435 111.86 92.64 ;
      RECT  114.98 92.64 114.77 94.345 ;
      RECT  112.79 92.055 112.58 92.435 ;
      RECT  114.23 92.64 114.05 94.345 ;
      RECT  113.51 92.64 113.33 94.345 ;
      RECT  114.23 91.725 114.05 92.64 ;
      RECT  112.07 91.725 111.86 92.055 ;
      RECT  113.87 92.64 113.69 94.345 ;
      RECT  113.87 91.725 113.69 92.64 ;
      RECT  115.19 92.435 114.98 92.64 ;
      RECT  112.07 92.055 111.86 92.435 ;
      RECT  113.15 92.64 112.97 94.345 ;
      RECT  114.98 92.435 114.77 92.64 ;
      RECT  115.19 92.055 114.98 92.435 ;
      POLYGON  112.58 93.72 112.58 94.13 112.325 94.13 112.325 93.8 112.405 93.72 112.58 93.72 ;
      RECT  114.59 91.725 114.41 92.64 ;
      RECT  114.98 91.725 114.77 92.055 ;
      RECT  114.98 92.055 114.77 92.435 ;
      RECT  112.79 95.71 112.58 95.3 ;
      RECT  115.19 96.715 114.98 96.385 ;
      RECT  112.145 95.8 112.07 94.095 ;
      RECT  112.23 95.215 112.145 94.805 ;
      RECT  113.15 96.715 112.97 95.8 ;
      POLYGON  112.145 96.715 112.145 96.385 112.58 96.385 112.58 96.005 112.145 96.005 112.145 95.8 112.07 95.8 112.07 96.715 112.145 96.715 ;
      RECT  112.07 95.8 111.86 94.095 ;
      POLYGON  112.58 95.71 112.58 95.3 112.405 95.3 112.325 95.38 112.325 95.71 112.58 95.71 ;
      RECT  115.19 95.8 114.98 94.095 ;
      RECT  113.51 96.715 113.33 95.8 ;
      RECT  114.59 95.8 114.41 94.095 ;
      RECT  112.79 94.72 112.58 94.31 ;
      RECT  112.07 96.005 111.86 95.8 ;
      RECT  114.98 95.8 114.77 94.095 ;
      RECT  112.79 96.385 112.58 96.005 ;
      RECT  114.23 95.8 114.05 94.095 ;
      RECT  113.51 95.8 113.33 94.095 ;
      RECT  114.23 96.715 114.05 95.8 ;
      RECT  112.07 96.715 111.86 96.385 ;
      RECT  113.87 95.8 113.69 94.095 ;
      RECT  113.87 96.715 113.69 95.8 ;
      RECT  115.19 96.005 114.98 95.8 ;
      RECT  112.07 96.385 111.86 96.005 ;
      RECT  113.15 95.8 112.97 94.095 ;
      RECT  114.98 96.005 114.77 95.8 ;
      RECT  115.19 96.385 114.98 96.005 ;
      POLYGON  112.58 94.72 112.58 94.31 112.325 94.31 112.325 94.64 112.405 94.72 112.58 94.72 ;
      RECT  114.59 96.715 114.41 95.8 ;
      RECT  114.98 96.715 114.77 96.385 ;
      RECT  114.98 96.385 114.77 96.005 ;
      RECT  112.79 96.68 112.58 97.09 ;
      RECT  115.19 95.675 114.98 96.005 ;
      RECT  112.145 96.59 112.07 98.295 ;
      RECT  112.23 97.175 112.145 97.585 ;
      RECT  113.15 95.675 112.97 96.59 ;
      POLYGON  112.145 95.675 112.145 96.005 112.58 96.005 112.58 96.385 112.145 96.385 112.145 96.59 112.07 96.59 112.07 95.675 112.145 95.675 ;
      RECT  112.07 96.59 111.86 98.295 ;
      POLYGON  112.58 96.68 112.58 97.09 112.405 97.09 112.325 97.01 112.325 96.68 112.58 96.68 ;
      RECT  115.19 96.59 114.98 98.295 ;
      RECT  113.51 95.675 113.33 96.59 ;
      RECT  114.59 96.59 114.41 98.295 ;
      RECT  112.79 97.67 112.58 98.08 ;
      RECT  112.07 96.385 111.86 96.59 ;
      RECT  114.98 96.59 114.77 98.295 ;
      RECT  112.79 96.005 112.58 96.385 ;
      RECT  114.23 96.59 114.05 98.295 ;
      RECT  113.51 96.59 113.33 98.295 ;
      RECT  114.23 95.675 114.05 96.59 ;
      RECT  112.07 95.675 111.86 96.005 ;
      RECT  113.87 96.59 113.69 98.295 ;
      RECT  113.87 95.675 113.69 96.59 ;
      RECT  115.19 96.385 114.98 96.59 ;
      RECT  112.07 96.005 111.86 96.385 ;
      RECT  113.15 96.59 112.97 98.295 ;
      RECT  114.98 96.385 114.77 96.59 ;
      RECT  115.19 96.005 114.98 96.385 ;
      POLYGON  112.58 97.67 112.58 98.08 112.325 98.08 112.325 97.75 112.405 97.67 112.58 97.67 ;
      RECT  114.59 95.675 114.41 96.59 ;
      RECT  114.98 95.675 114.77 96.005 ;
      RECT  114.98 96.005 114.77 96.385 ;
      RECT  112.79 99.66 112.58 99.25 ;
      RECT  115.19 100.665 114.98 100.335 ;
      RECT  112.145 99.75 112.07 98.045 ;
      RECT  112.23 99.165 112.145 98.755 ;
      RECT  113.15 100.665 112.97 99.75 ;
      POLYGON  112.145 100.665 112.145 100.335 112.58 100.335 112.58 99.955 112.145 99.955 112.145 99.75 112.07 99.75 112.07 100.665 112.145 100.665 ;
      RECT  112.07 99.75 111.86 98.045 ;
      POLYGON  112.58 99.66 112.58 99.25 112.405 99.25 112.325 99.33 112.325 99.66 112.58 99.66 ;
      RECT  115.19 99.75 114.98 98.045 ;
      RECT  113.51 100.665 113.33 99.75 ;
      RECT  114.59 99.75 114.41 98.045 ;
      RECT  112.79 98.67 112.58 98.26 ;
      RECT  112.07 99.955 111.86 99.75 ;
      RECT  114.98 99.75 114.77 98.045 ;
      RECT  112.79 100.335 112.58 99.955 ;
      RECT  114.23 99.75 114.05 98.045 ;
      RECT  113.51 99.75 113.33 98.045 ;
      RECT  114.23 100.665 114.05 99.75 ;
      RECT  112.07 100.665 111.86 100.335 ;
      RECT  113.87 99.75 113.69 98.045 ;
      RECT  113.87 100.665 113.69 99.75 ;
      RECT  115.19 99.955 114.98 99.75 ;
      RECT  112.07 100.335 111.86 99.955 ;
      RECT  113.15 99.75 112.97 98.045 ;
      RECT  114.98 99.955 114.77 99.75 ;
      RECT  115.19 100.335 114.98 99.955 ;
      POLYGON  112.58 98.67 112.58 98.26 112.325 98.26 112.325 98.59 112.405 98.67 112.58 98.67 ;
      RECT  114.59 100.665 114.41 99.75 ;
      RECT  114.98 100.665 114.77 100.335 ;
      RECT  114.98 100.335 114.77 99.955 ;
      RECT  112.79 100.63 112.58 101.04 ;
      RECT  115.19 99.625 114.98 99.955 ;
      RECT  112.145 100.54 112.07 102.245 ;
      RECT  112.23 101.125 112.145 101.535 ;
      RECT  113.15 99.625 112.97 100.54 ;
      POLYGON  112.145 99.625 112.145 99.955 112.58 99.955 112.58 100.335 112.145 100.335 112.145 100.54 112.07 100.54 112.07 99.625 112.145 99.625 ;
      RECT  112.07 100.54 111.86 102.245 ;
      POLYGON  112.58 100.63 112.58 101.04 112.405 101.04 112.325 100.96 112.325 100.63 112.58 100.63 ;
      RECT  115.19 100.54 114.98 102.245 ;
      RECT  113.51 99.625 113.33 100.54 ;
      RECT  114.59 100.54 114.41 102.245 ;
      RECT  112.79 101.62 112.58 102.03 ;
      RECT  112.07 100.335 111.86 100.54 ;
      RECT  114.98 100.54 114.77 102.245 ;
      RECT  112.79 99.955 112.58 100.335 ;
      RECT  114.23 100.54 114.05 102.245 ;
      RECT  113.51 100.54 113.33 102.245 ;
      RECT  114.23 99.625 114.05 100.54 ;
      RECT  112.07 99.625 111.86 99.955 ;
      RECT  113.87 100.54 113.69 102.245 ;
      RECT  113.87 99.625 113.69 100.54 ;
      RECT  115.19 100.335 114.98 100.54 ;
      RECT  112.07 99.955 111.86 100.335 ;
      RECT  113.15 100.54 112.97 102.245 ;
      RECT  114.98 100.335 114.77 100.54 ;
      RECT  115.19 99.955 114.98 100.335 ;
      POLYGON  112.58 101.62 112.58 102.03 112.325 102.03 112.325 101.7 112.405 101.62 112.58 101.62 ;
      RECT  114.59 99.625 114.41 100.54 ;
      RECT  114.98 99.625 114.77 99.955 ;
      RECT  114.98 99.955 114.77 100.335 ;
      RECT  112.79 103.61 112.58 103.2 ;
      RECT  115.19 104.615 114.98 104.285 ;
      RECT  112.145 103.7 112.07 101.995 ;
      RECT  112.23 103.115 112.145 102.705 ;
      RECT  113.15 104.615 112.97 103.7 ;
      POLYGON  112.145 104.615 112.145 104.285 112.58 104.285 112.58 103.905 112.145 103.905 112.145 103.7 112.07 103.7 112.07 104.615 112.145 104.615 ;
      RECT  112.07 103.7 111.86 101.995 ;
      POLYGON  112.58 103.61 112.58 103.2 112.405 103.2 112.325 103.28 112.325 103.61 112.58 103.61 ;
      RECT  115.19 103.7 114.98 101.995 ;
      RECT  113.51 104.615 113.33 103.7 ;
      RECT  114.59 103.7 114.41 101.995 ;
      RECT  112.79 102.62 112.58 102.21 ;
      RECT  112.07 103.905 111.86 103.7 ;
      RECT  114.98 103.7 114.77 101.995 ;
      RECT  112.79 104.285 112.58 103.905 ;
      RECT  114.23 103.7 114.05 101.995 ;
      RECT  113.51 103.7 113.33 101.995 ;
      RECT  114.23 104.615 114.05 103.7 ;
      RECT  112.07 104.615 111.86 104.285 ;
      RECT  113.87 103.7 113.69 101.995 ;
      RECT  113.87 104.615 113.69 103.7 ;
      RECT  115.19 103.905 114.98 103.7 ;
      RECT  112.07 104.285 111.86 103.905 ;
      RECT  113.15 103.7 112.97 101.995 ;
      RECT  114.98 103.905 114.77 103.7 ;
      RECT  115.19 104.285 114.98 103.905 ;
      POLYGON  112.58 102.62 112.58 102.21 112.325 102.21 112.325 102.54 112.405 102.62 112.58 102.62 ;
      RECT  114.59 104.615 114.41 103.7 ;
      RECT  114.98 104.615 114.77 104.285 ;
      RECT  114.98 104.285 114.77 103.905 ;
      RECT  112.79 104.58 112.58 104.99 ;
      RECT  115.19 103.575 114.98 103.905 ;
      RECT  112.145 104.49 112.07 106.195 ;
      RECT  112.23 105.075 112.145 105.485 ;
      RECT  113.15 103.575 112.97 104.49 ;
      POLYGON  112.145 103.575 112.145 103.905 112.58 103.905 112.58 104.285 112.145 104.285 112.145 104.49 112.07 104.49 112.07 103.575 112.145 103.575 ;
      RECT  112.07 104.49 111.86 106.195 ;
      POLYGON  112.58 104.58 112.58 104.99 112.405 104.99 112.325 104.91 112.325 104.58 112.58 104.58 ;
      RECT  115.19 104.49 114.98 106.195 ;
      RECT  113.51 103.575 113.33 104.49 ;
      RECT  114.59 104.49 114.41 106.195 ;
      RECT  112.79 105.57 112.58 105.98 ;
      RECT  112.07 104.285 111.86 104.49 ;
      RECT  114.98 104.49 114.77 106.195 ;
      RECT  112.79 103.905 112.58 104.285 ;
      RECT  114.23 104.49 114.05 106.195 ;
      RECT  113.51 104.49 113.33 106.195 ;
      RECT  114.23 103.575 114.05 104.49 ;
      RECT  112.07 103.575 111.86 103.905 ;
      RECT  113.87 104.49 113.69 106.195 ;
      RECT  113.87 103.575 113.69 104.49 ;
      RECT  115.19 104.285 114.98 104.49 ;
      RECT  112.07 103.905 111.86 104.285 ;
      RECT  113.15 104.49 112.97 106.195 ;
      RECT  114.98 104.285 114.77 104.49 ;
      RECT  115.19 103.905 114.98 104.285 ;
      POLYGON  112.58 105.57 112.58 105.98 112.325 105.98 112.325 105.65 112.405 105.57 112.58 105.57 ;
      RECT  114.59 103.575 114.41 104.49 ;
      RECT  114.98 103.575 114.77 103.905 ;
      RECT  114.98 103.905 114.77 104.285 ;
      RECT  112.79 107.56 112.58 107.15 ;
      RECT  115.19 108.565 114.98 108.235 ;
      RECT  112.145 107.65 112.07 105.945 ;
      RECT  112.23 107.065 112.145 106.655 ;
      RECT  113.15 108.565 112.97 107.65 ;
      POLYGON  112.145 108.565 112.145 108.235 112.58 108.235 112.58 107.855 112.145 107.855 112.145 107.65 112.07 107.65 112.07 108.565 112.145 108.565 ;
      RECT  112.07 107.65 111.86 105.945 ;
      POLYGON  112.58 107.56 112.58 107.15 112.405 107.15 112.325 107.23 112.325 107.56 112.58 107.56 ;
      RECT  115.19 107.65 114.98 105.945 ;
      RECT  113.51 108.565 113.33 107.65 ;
      RECT  114.59 107.65 114.41 105.945 ;
      RECT  112.79 106.57 112.58 106.16 ;
      RECT  112.07 107.855 111.86 107.65 ;
      RECT  114.98 107.65 114.77 105.945 ;
      RECT  112.79 108.235 112.58 107.855 ;
      RECT  114.23 107.65 114.05 105.945 ;
      RECT  113.51 107.65 113.33 105.945 ;
      RECT  114.23 108.565 114.05 107.65 ;
      RECT  112.07 108.565 111.86 108.235 ;
      RECT  113.87 107.65 113.69 105.945 ;
      RECT  113.87 108.565 113.69 107.65 ;
      RECT  115.19 107.855 114.98 107.65 ;
      RECT  112.07 108.235 111.86 107.855 ;
      RECT  113.15 107.65 112.97 105.945 ;
      RECT  114.98 107.855 114.77 107.65 ;
      RECT  115.19 108.235 114.98 107.855 ;
      POLYGON  112.58 106.57 112.58 106.16 112.325 106.16 112.325 106.49 112.405 106.57 112.58 106.57 ;
      RECT  114.59 108.565 114.41 107.65 ;
      RECT  114.98 108.565 114.77 108.235 ;
      RECT  114.98 108.235 114.77 107.855 ;
      RECT  112.79 108.53 112.58 108.94 ;
      RECT  115.19 107.525 114.98 107.855 ;
      RECT  112.145 108.44 112.07 110.145 ;
      RECT  112.23 109.025 112.145 109.435 ;
      RECT  113.15 107.525 112.97 108.44 ;
      POLYGON  112.145 107.525 112.145 107.855 112.58 107.855 112.58 108.235 112.145 108.235 112.145 108.44 112.07 108.44 112.07 107.525 112.145 107.525 ;
      RECT  112.07 108.44 111.86 110.145 ;
      POLYGON  112.58 108.53 112.58 108.94 112.405 108.94 112.325 108.86 112.325 108.53 112.58 108.53 ;
      RECT  115.19 108.44 114.98 110.145 ;
      RECT  113.51 107.525 113.33 108.44 ;
      RECT  114.59 108.44 114.41 110.145 ;
      RECT  112.79 109.52 112.58 109.93 ;
      RECT  112.07 108.235 111.86 108.44 ;
      RECT  114.98 108.44 114.77 110.145 ;
      RECT  112.79 107.855 112.58 108.235 ;
      RECT  114.23 108.44 114.05 110.145 ;
      RECT  113.51 108.44 113.33 110.145 ;
      RECT  114.23 107.525 114.05 108.44 ;
      RECT  112.07 107.525 111.86 107.855 ;
      RECT  113.87 108.44 113.69 110.145 ;
      RECT  113.87 107.525 113.69 108.44 ;
      RECT  115.19 108.235 114.98 108.44 ;
      RECT  112.07 107.855 111.86 108.235 ;
      RECT  113.15 108.44 112.97 110.145 ;
      RECT  114.98 108.235 114.77 108.44 ;
      RECT  115.19 107.855 114.98 108.235 ;
      POLYGON  112.58 109.52 112.58 109.93 112.325 109.93 112.325 109.6 112.405 109.52 112.58 109.52 ;
      RECT  114.59 107.525 114.41 108.44 ;
      RECT  114.98 107.525 114.77 107.855 ;
      RECT  114.98 107.855 114.77 108.235 ;
      RECT  112.79 111.51 112.58 111.1 ;
      RECT  115.19 112.515 114.98 112.185 ;
      RECT  112.145 111.6 112.07 109.895 ;
      RECT  112.23 111.015 112.145 110.605 ;
      RECT  113.15 112.515 112.97 111.6 ;
      POLYGON  112.145 112.515 112.145 112.185 112.58 112.185 112.58 111.805 112.145 111.805 112.145 111.6 112.07 111.6 112.07 112.515 112.145 112.515 ;
      RECT  112.07 111.6 111.86 109.895 ;
      POLYGON  112.58 111.51 112.58 111.1 112.405 111.1 112.325 111.18 112.325 111.51 112.58 111.51 ;
      RECT  115.19 111.6 114.98 109.895 ;
      RECT  113.51 112.515 113.33 111.6 ;
      RECT  114.59 111.6 114.41 109.895 ;
      RECT  112.79 110.52 112.58 110.11 ;
      RECT  112.07 111.805 111.86 111.6 ;
      RECT  114.98 111.6 114.77 109.895 ;
      RECT  112.79 112.185 112.58 111.805 ;
      RECT  114.23 111.6 114.05 109.895 ;
      RECT  113.51 111.6 113.33 109.895 ;
      RECT  114.23 112.515 114.05 111.6 ;
      RECT  112.07 112.515 111.86 112.185 ;
      RECT  113.87 111.6 113.69 109.895 ;
      RECT  113.87 112.515 113.69 111.6 ;
      RECT  115.19 111.805 114.98 111.6 ;
      RECT  112.07 112.185 111.86 111.805 ;
      RECT  113.15 111.6 112.97 109.895 ;
      RECT  114.98 111.805 114.77 111.6 ;
      RECT  115.19 112.185 114.98 111.805 ;
      POLYGON  112.58 110.52 112.58 110.11 112.325 110.11 112.325 110.44 112.405 110.52 112.58 110.52 ;
      RECT  114.59 112.515 114.41 111.6 ;
      RECT  114.98 112.515 114.77 112.185 ;
      RECT  114.98 112.185 114.77 111.805 ;
      RECT  112.79 112.48 112.58 112.89 ;
      RECT  115.19 111.475 114.98 111.805 ;
      RECT  112.145 112.39 112.07 114.095 ;
      RECT  112.23 112.975 112.145 113.385 ;
      RECT  113.15 111.475 112.97 112.39 ;
      POLYGON  112.145 111.475 112.145 111.805 112.58 111.805 112.58 112.185 112.145 112.185 112.145 112.39 112.07 112.39 112.07 111.475 112.145 111.475 ;
      RECT  112.07 112.39 111.86 114.095 ;
      POLYGON  112.58 112.48 112.58 112.89 112.405 112.89 112.325 112.81 112.325 112.48 112.58 112.48 ;
      RECT  115.19 112.39 114.98 114.095 ;
      RECT  113.51 111.475 113.33 112.39 ;
      RECT  114.59 112.39 114.41 114.095 ;
      RECT  112.79 113.47 112.58 113.88 ;
      RECT  112.07 112.185 111.86 112.39 ;
      RECT  114.98 112.39 114.77 114.095 ;
      RECT  112.79 111.805 112.58 112.185 ;
      RECT  114.23 112.39 114.05 114.095 ;
      RECT  113.51 112.39 113.33 114.095 ;
      RECT  114.23 111.475 114.05 112.39 ;
      RECT  112.07 111.475 111.86 111.805 ;
      RECT  113.87 112.39 113.69 114.095 ;
      RECT  113.87 111.475 113.69 112.39 ;
      RECT  115.19 112.185 114.98 112.39 ;
      RECT  112.07 111.805 111.86 112.185 ;
      RECT  113.15 112.39 112.97 114.095 ;
      RECT  114.98 112.185 114.77 112.39 ;
      RECT  115.19 111.805 114.98 112.185 ;
      POLYGON  112.58 113.47 112.58 113.88 112.325 113.88 112.325 113.55 112.405 113.47 112.58 113.47 ;
      RECT  114.59 111.475 114.41 112.39 ;
      RECT  114.98 111.475 114.77 111.805 ;
      RECT  114.98 111.805 114.77 112.185 ;
      RECT  112.79 115.46 112.58 115.05 ;
      RECT  115.19 116.465 114.98 116.135 ;
      RECT  112.145 115.55 112.07 113.845 ;
      RECT  112.23 114.965 112.145 114.555 ;
      RECT  113.15 116.465 112.97 115.55 ;
      POLYGON  112.145 116.465 112.145 116.135 112.58 116.135 112.58 115.755 112.145 115.755 112.145 115.55 112.07 115.55 112.07 116.465 112.145 116.465 ;
      RECT  112.07 115.55 111.86 113.845 ;
      POLYGON  112.58 115.46 112.58 115.05 112.405 115.05 112.325 115.13 112.325 115.46 112.58 115.46 ;
      RECT  115.19 115.55 114.98 113.845 ;
      RECT  113.51 116.465 113.33 115.55 ;
      RECT  114.59 115.55 114.41 113.845 ;
      RECT  112.79 114.47 112.58 114.06 ;
      RECT  112.07 115.755 111.86 115.55 ;
      RECT  114.98 115.55 114.77 113.845 ;
      RECT  112.79 116.135 112.58 115.755 ;
      RECT  114.23 115.55 114.05 113.845 ;
      RECT  113.51 115.55 113.33 113.845 ;
      RECT  114.23 116.465 114.05 115.55 ;
      RECT  112.07 116.465 111.86 116.135 ;
      RECT  113.87 115.55 113.69 113.845 ;
      RECT  113.87 116.465 113.69 115.55 ;
      RECT  115.19 115.755 114.98 115.55 ;
      RECT  112.07 116.135 111.86 115.755 ;
      RECT  113.15 115.55 112.97 113.845 ;
      RECT  114.98 115.755 114.77 115.55 ;
      RECT  115.19 116.135 114.98 115.755 ;
      POLYGON  112.58 114.47 112.58 114.06 112.325 114.06 112.325 114.39 112.405 114.47 112.58 114.47 ;
      RECT  114.59 116.465 114.41 115.55 ;
      RECT  114.98 116.465 114.77 116.135 ;
      RECT  114.98 116.135 114.77 115.755 ;
      RECT  112.79 116.43 112.58 116.84 ;
      RECT  115.19 115.425 114.98 115.755 ;
      RECT  112.145 116.34 112.07 118.045 ;
      RECT  112.23 116.925 112.145 117.335 ;
      RECT  113.15 115.425 112.97 116.34 ;
      POLYGON  112.145 115.425 112.145 115.755 112.58 115.755 112.58 116.135 112.145 116.135 112.145 116.34 112.07 116.34 112.07 115.425 112.145 115.425 ;
      RECT  112.07 116.34 111.86 118.045 ;
      POLYGON  112.58 116.43 112.58 116.84 112.405 116.84 112.325 116.76 112.325 116.43 112.58 116.43 ;
      RECT  115.19 116.34 114.98 118.045 ;
      RECT  113.51 115.425 113.33 116.34 ;
      RECT  114.59 116.34 114.41 118.045 ;
      RECT  112.79 117.42 112.58 117.83 ;
      RECT  112.07 116.135 111.86 116.34 ;
      RECT  114.98 116.34 114.77 118.045 ;
      RECT  112.79 115.755 112.58 116.135 ;
      RECT  114.23 116.34 114.05 118.045 ;
      RECT  113.51 116.34 113.33 118.045 ;
      RECT  114.23 115.425 114.05 116.34 ;
      RECT  112.07 115.425 111.86 115.755 ;
      RECT  113.87 116.34 113.69 118.045 ;
      RECT  113.87 115.425 113.69 116.34 ;
      RECT  115.19 116.135 114.98 116.34 ;
      RECT  112.07 115.755 111.86 116.135 ;
      RECT  113.15 116.34 112.97 118.045 ;
      RECT  114.98 116.135 114.77 116.34 ;
      RECT  115.19 115.755 114.98 116.135 ;
      POLYGON  112.58 117.42 112.58 117.83 112.325 117.83 112.325 117.5 112.405 117.42 112.58 117.42 ;
      RECT  114.59 115.425 114.41 116.34 ;
      RECT  114.98 115.425 114.77 115.755 ;
      RECT  114.98 115.755 114.77 116.135 ;
      RECT  112.79 119.41 112.58 119.0 ;
      RECT  115.19 120.415 114.98 120.085 ;
      RECT  112.145 119.5 112.07 117.795 ;
      RECT  112.23 118.915 112.145 118.505 ;
      RECT  113.15 120.415 112.97 119.5 ;
      POLYGON  112.145 120.415 112.145 120.085 112.58 120.085 112.58 119.705 112.145 119.705 112.145 119.5 112.07 119.5 112.07 120.415 112.145 120.415 ;
      RECT  112.07 119.5 111.86 117.795 ;
      POLYGON  112.58 119.41 112.58 119.0 112.405 119.0 112.325 119.08 112.325 119.41 112.58 119.41 ;
      RECT  115.19 119.5 114.98 117.795 ;
      RECT  113.51 120.415 113.33 119.5 ;
      RECT  114.59 119.5 114.41 117.795 ;
      RECT  112.79 118.42 112.58 118.01 ;
      RECT  112.07 119.705 111.86 119.5 ;
      RECT  114.98 119.5 114.77 117.795 ;
      RECT  112.79 120.085 112.58 119.705 ;
      RECT  114.23 119.5 114.05 117.795 ;
      RECT  113.51 119.5 113.33 117.795 ;
      RECT  114.23 120.415 114.05 119.5 ;
      RECT  112.07 120.415 111.86 120.085 ;
      RECT  113.87 119.5 113.69 117.795 ;
      RECT  113.87 120.415 113.69 119.5 ;
      RECT  115.19 119.705 114.98 119.5 ;
      RECT  112.07 120.085 111.86 119.705 ;
      RECT  113.15 119.5 112.97 117.795 ;
      RECT  114.98 119.705 114.77 119.5 ;
      RECT  115.19 120.085 114.98 119.705 ;
      POLYGON  112.58 118.42 112.58 118.01 112.325 118.01 112.325 118.34 112.405 118.42 112.58 118.42 ;
      RECT  114.59 120.415 114.41 119.5 ;
      RECT  114.98 120.415 114.77 120.085 ;
      RECT  114.98 120.085 114.77 119.705 ;
      RECT  112.79 120.38 112.58 120.79 ;
      RECT  115.19 119.375 114.98 119.705 ;
      RECT  112.145 120.29 112.07 121.995 ;
      RECT  112.23 120.875 112.145 121.285 ;
      RECT  113.15 119.375 112.97 120.29 ;
      POLYGON  112.145 119.375 112.145 119.705 112.58 119.705 112.58 120.085 112.145 120.085 112.145 120.29 112.07 120.29 112.07 119.375 112.145 119.375 ;
      RECT  112.07 120.29 111.86 121.995 ;
      POLYGON  112.58 120.38 112.58 120.79 112.405 120.79 112.325 120.71 112.325 120.38 112.58 120.38 ;
      RECT  115.19 120.29 114.98 121.995 ;
      RECT  113.51 119.375 113.33 120.29 ;
      RECT  114.59 120.29 114.41 121.995 ;
      RECT  112.79 121.37 112.58 121.78 ;
      RECT  112.07 120.085 111.86 120.29 ;
      RECT  114.98 120.29 114.77 121.995 ;
      RECT  112.79 119.705 112.58 120.085 ;
      RECT  114.23 120.29 114.05 121.995 ;
      RECT  113.51 120.29 113.33 121.995 ;
      RECT  114.23 119.375 114.05 120.29 ;
      RECT  112.07 119.375 111.86 119.705 ;
      RECT  113.87 120.29 113.69 121.995 ;
      RECT  113.87 119.375 113.69 120.29 ;
      RECT  115.19 120.085 114.98 120.29 ;
      RECT  112.07 119.705 111.86 120.085 ;
      RECT  113.15 120.29 112.97 121.995 ;
      RECT  114.98 120.085 114.77 120.29 ;
      RECT  115.19 119.705 114.98 120.085 ;
      POLYGON  112.58 121.37 112.58 121.78 112.325 121.78 112.325 121.45 112.405 121.37 112.58 121.37 ;
      RECT  114.59 119.375 114.41 120.29 ;
      RECT  114.98 119.375 114.77 119.705 ;
      RECT  114.98 119.705 114.77 120.085 ;
      RECT  112.79 123.36 112.58 122.95 ;
      RECT  115.19 124.365 114.98 124.035 ;
      RECT  112.145 123.45 112.07 121.745 ;
      RECT  112.23 122.865 112.145 122.455 ;
      RECT  113.15 124.365 112.97 123.45 ;
      POLYGON  112.145 124.365 112.145 124.035 112.58 124.035 112.58 123.655 112.145 123.655 112.145 123.45 112.07 123.45 112.07 124.365 112.145 124.365 ;
      RECT  112.07 123.45 111.86 121.745 ;
      POLYGON  112.58 123.36 112.58 122.95 112.405 122.95 112.325 123.03 112.325 123.36 112.58 123.36 ;
      RECT  115.19 123.45 114.98 121.745 ;
      RECT  113.51 124.365 113.33 123.45 ;
      RECT  114.59 123.45 114.41 121.745 ;
      RECT  112.79 122.37 112.58 121.96 ;
      RECT  112.07 123.655 111.86 123.45 ;
      RECT  114.98 123.45 114.77 121.745 ;
      RECT  112.79 124.035 112.58 123.655 ;
      RECT  114.23 123.45 114.05 121.745 ;
      RECT  113.51 123.45 113.33 121.745 ;
      RECT  114.23 124.365 114.05 123.45 ;
      RECT  112.07 124.365 111.86 124.035 ;
      RECT  113.87 123.45 113.69 121.745 ;
      RECT  113.87 124.365 113.69 123.45 ;
      RECT  115.19 123.655 114.98 123.45 ;
      RECT  112.07 124.035 111.86 123.655 ;
      RECT  113.15 123.45 112.97 121.745 ;
      RECT  114.98 123.655 114.77 123.45 ;
      RECT  115.19 124.035 114.98 123.655 ;
      POLYGON  112.58 122.37 112.58 121.96 112.325 121.96 112.325 122.29 112.405 122.37 112.58 122.37 ;
      RECT  114.59 124.365 114.41 123.45 ;
      RECT  114.98 124.365 114.77 124.035 ;
      RECT  114.98 124.035 114.77 123.655 ;
      RECT  117.17 92.73 117.38 93.14 ;
      RECT  114.77 91.725 114.98 92.055 ;
      RECT  117.815 92.64 117.89 94.345 ;
      RECT  117.73 93.225 117.815 93.635 ;
      RECT  116.81 91.725 116.99 92.64 ;
      POLYGON  117.815 91.725 117.815 92.055 117.38 92.055 117.38 92.435 117.815 92.435 117.815 92.64 117.89 92.64 117.89 91.725 117.815 91.725 ;
      RECT  117.89 92.64 118.1 94.345 ;
      POLYGON  117.38 92.73 117.38 93.14 117.555 93.14 117.635 93.06 117.635 92.73 117.38 92.73 ;
      RECT  114.77 92.64 114.98 94.345 ;
      RECT  116.45 91.725 116.63 92.64 ;
      RECT  115.37 92.64 115.55 94.345 ;
      RECT  117.17 93.72 117.38 94.13 ;
      RECT  117.89 92.435 118.1 92.64 ;
      RECT  114.98 92.64 115.19 94.345 ;
      RECT  117.17 92.055 117.38 92.435 ;
      RECT  115.73 92.64 115.91 94.345 ;
      RECT  116.45 92.64 116.63 94.345 ;
      RECT  115.73 91.725 115.91 92.64 ;
      RECT  117.89 91.725 118.1 92.055 ;
      RECT  116.09 92.64 116.27 94.345 ;
      RECT  116.09 91.725 116.27 92.64 ;
      RECT  114.77 92.435 114.98 92.64 ;
      RECT  117.89 92.055 118.1 92.435 ;
      RECT  116.81 92.64 116.99 94.345 ;
      RECT  114.98 92.435 115.19 92.64 ;
      RECT  114.77 92.055 114.98 92.435 ;
      POLYGON  117.38 93.72 117.38 94.13 117.635 94.13 117.635 93.8 117.555 93.72 117.38 93.72 ;
      RECT  115.37 91.725 115.55 92.64 ;
      RECT  114.98 91.725 115.19 92.055 ;
      RECT  114.98 92.055 115.19 92.435 ;
      RECT  117.17 95.71 117.38 95.3 ;
      RECT  114.77 96.715 114.98 96.385 ;
      RECT  117.815 95.8 117.89 94.095 ;
      RECT  117.73 95.215 117.815 94.805 ;
      RECT  116.81 96.715 116.99 95.8 ;
      POLYGON  117.815 96.715 117.815 96.385 117.38 96.385 117.38 96.005 117.815 96.005 117.815 95.8 117.89 95.8 117.89 96.715 117.815 96.715 ;
      RECT  117.89 95.8 118.1 94.095 ;
      POLYGON  117.38 95.71 117.38 95.3 117.555 95.3 117.635 95.38 117.635 95.71 117.38 95.71 ;
      RECT  114.77 95.8 114.98 94.095 ;
      RECT  116.45 96.715 116.63 95.8 ;
      RECT  115.37 95.8 115.55 94.095 ;
      RECT  117.17 94.72 117.38 94.31 ;
      RECT  117.89 96.005 118.1 95.8 ;
      RECT  114.98 95.8 115.19 94.095 ;
      RECT  117.17 96.385 117.38 96.005 ;
      RECT  115.73 95.8 115.91 94.095 ;
      RECT  116.45 95.8 116.63 94.095 ;
      RECT  115.73 96.715 115.91 95.8 ;
      RECT  117.89 96.715 118.1 96.385 ;
      RECT  116.09 95.8 116.27 94.095 ;
      RECT  116.09 96.715 116.27 95.8 ;
      RECT  114.77 96.005 114.98 95.8 ;
      RECT  117.89 96.385 118.1 96.005 ;
      RECT  116.81 95.8 116.99 94.095 ;
      RECT  114.98 96.005 115.19 95.8 ;
      RECT  114.77 96.385 114.98 96.005 ;
      POLYGON  117.38 94.72 117.38 94.31 117.635 94.31 117.635 94.64 117.555 94.72 117.38 94.72 ;
      RECT  115.37 96.715 115.55 95.8 ;
      RECT  114.98 96.715 115.19 96.385 ;
      RECT  114.98 96.385 115.19 96.005 ;
      RECT  117.17 96.68 117.38 97.09 ;
      RECT  114.77 95.675 114.98 96.005 ;
      RECT  117.815 96.59 117.89 98.295 ;
      RECT  117.73 97.175 117.815 97.585 ;
      RECT  116.81 95.675 116.99 96.59 ;
      POLYGON  117.815 95.675 117.815 96.005 117.38 96.005 117.38 96.385 117.815 96.385 117.815 96.59 117.89 96.59 117.89 95.675 117.815 95.675 ;
      RECT  117.89 96.59 118.1 98.295 ;
      POLYGON  117.38 96.68 117.38 97.09 117.555 97.09 117.635 97.01 117.635 96.68 117.38 96.68 ;
      RECT  114.77 96.59 114.98 98.295 ;
      RECT  116.45 95.675 116.63 96.59 ;
      RECT  115.37 96.59 115.55 98.295 ;
      RECT  117.17 97.67 117.38 98.08 ;
      RECT  117.89 96.385 118.1 96.59 ;
      RECT  114.98 96.59 115.19 98.295 ;
      RECT  117.17 96.005 117.38 96.385 ;
      RECT  115.73 96.59 115.91 98.295 ;
      RECT  116.45 96.59 116.63 98.295 ;
      RECT  115.73 95.675 115.91 96.59 ;
      RECT  117.89 95.675 118.1 96.005 ;
      RECT  116.09 96.59 116.27 98.295 ;
      RECT  116.09 95.675 116.27 96.59 ;
      RECT  114.77 96.385 114.98 96.59 ;
      RECT  117.89 96.005 118.1 96.385 ;
      RECT  116.81 96.59 116.99 98.295 ;
      RECT  114.98 96.385 115.19 96.59 ;
      RECT  114.77 96.005 114.98 96.385 ;
      POLYGON  117.38 97.67 117.38 98.08 117.635 98.08 117.635 97.75 117.555 97.67 117.38 97.67 ;
      RECT  115.37 95.675 115.55 96.59 ;
      RECT  114.98 95.675 115.19 96.005 ;
      RECT  114.98 96.005 115.19 96.385 ;
      RECT  117.17 99.66 117.38 99.25 ;
      RECT  114.77 100.665 114.98 100.335 ;
      RECT  117.815 99.75 117.89 98.045 ;
      RECT  117.73 99.165 117.815 98.755 ;
      RECT  116.81 100.665 116.99 99.75 ;
      POLYGON  117.815 100.665 117.815 100.335 117.38 100.335 117.38 99.955 117.815 99.955 117.815 99.75 117.89 99.75 117.89 100.665 117.815 100.665 ;
      RECT  117.89 99.75 118.1 98.045 ;
      POLYGON  117.38 99.66 117.38 99.25 117.555 99.25 117.635 99.33 117.635 99.66 117.38 99.66 ;
      RECT  114.77 99.75 114.98 98.045 ;
      RECT  116.45 100.665 116.63 99.75 ;
      RECT  115.37 99.75 115.55 98.045 ;
      RECT  117.17 98.67 117.38 98.26 ;
      RECT  117.89 99.955 118.1 99.75 ;
      RECT  114.98 99.75 115.19 98.045 ;
      RECT  117.17 100.335 117.38 99.955 ;
      RECT  115.73 99.75 115.91 98.045 ;
      RECT  116.45 99.75 116.63 98.045 ;
      RECT  115.73 100.665 115.91 99.75 ;
      RECT  117.89 100.665 118.1 100.335 ;
      RECT  116.09 99.75 116.27 98.045 ;
      RECT  116.09 100.665 116.27 99.75 ;
      RECT  114.77 99.955 114.98 99.75 ;
      RECT  117.89 100.335 118.1 99.955 ;
      RECT  116.81 99.75 116.99 98.045 ;
      RECT  114.98 99.955 115.19 99.75 ;
      RECT  114.77 100.335 114.98 99.955 ;
      POLYGON  117.38 98.67 117.38 98.26 117.635 98.26 117.635 98.59 117.555 98.67 117.38 98.67 ;
      RECT  115.37 100.665 115.55 99.75 ;
      RECT  114.98 100.665 115.19 100.335 ;
      RECT  114.98 100.335 115.19 99.955 ;
      RECT  117.17 100.63 117.38 101.04 ;
      RECT  114.77 99.625 114.98 99.955 ;
      RECT  117.815 100.54 117.89 102.245 ;
      RECT  117.73 101.125 117.815 101.535 ;
      RECT  116.81 99.625 116.99 100.54 ;
      POLYGON  117.815 99.625 117.815 99.955 117.38 99.955 117.38 100.335 117.815 100.335 117.815 100.54 117.89 100.54 117.89 99.625 117.815 99.625 ;
      RECT  117.89 100.54 118.1 102.245 ;
      POLYGON  117.38 100.63 117.38 101.04 117.555 101.04 117.635 100.96 117.635 100.63 117.38 100.63 ;
      RECT  114.77 100.54 114.98 102.245 ;
      RECT  116.45 99.625 116.63 100.54 ;
      RECT  115.37 100.54 115.55 102.245 ;
      RECT  117.17 101.62 117.38 102.03 ;
      RECT  117.89 100.335 118.1 100.54 ;
      RECT  114.98 100.54 115.19 102.245 ;
      RECT  117.17 99.955 117.38 100.335 ;
      RECT  115.73 100.54 115.91 102.245 ;
      RECT  116.45 100.54 116.63 102.245 ;
      RECT  115.73 99.625 115.91 100.54 ;
      RECT  117.89 99.625 118.1 99.955 ;
      RECT  116.09 100.54 116.27 102.245 ;
      RECT  116.09 99.625 116.27 100.54 ;
      RECT  114.77 100.335 114.98 100.54 ;
      RECT  117.89 99.955 118.1 100.335 ;
      RECT  116.81 100.54 116.99 102.245 ;
      RECT  114.98 100.335 115.19 100.54 ;
      RECT  114.77 99.955 114.98 100.335 ;
      POLYGON  117.38 101.62 117.38 102.03 117.635 102.03 117.635 101.7 117.555 101.62 117.38 101.62 ;
      RECT  115.37 99.625 115.55 100.54 ;
      RECT  114.98 99.625 115.19 99.955 ;
      RECT  114.98 99.955 115.19 100.335 ;
      RECT  117.17 103.61 117.38 103.2 ;
      RECT  114.77 104.615 114.98 104.285 ;
      RECT  117.815 103.7 117.89 101.995 ;
      RECT  117.73 103.115 117.815 102.705 ;
      RECT  116.81 104.615 116.99 103.7 ;
      POLYGON  117.815 104.615 117.815 104.285 117.38 104.285 117.38 103.905 117.815 103.905 117.815 103.7 117.89 103.7 117.89 104.615 117.815 104.615 ;
      RECT  117.89 103.7 118.1 101.995 ;
      POLYGON  117.38 103.61 117.38 103.2 117.555 103.2 117.635 103.28 117.635 103.61 117.38 103.61 ;
      RECT  114.77 103.7 114.98 101.995 ;
      RECT  116.45 104.615 116.63 103.7 ;
      RECT  115.37 103.7 115.55 101.995 ;
      RECT  117.17 102.62 117.38 102.21 ;
      RECT  117.89 103.905 118.1 103.7 ;
      RECT  114.98 103.7 115.19 101.995 ;
      RECT  117.17 104.285 117.38 103.905 ;
      RECT  115.73 103.7 115.91 101.995 ;
      RECT  116.45 103.7 116.63 101.995 ;
      RECT  115.73 104.615 115.91 103.7 ;
      RECT  117.89 104.615 118.1 104.285 ;
      RECT  116.09 103.7 116.27 101.995 ;
      RECT  116.09 104.615 116.27 103.7 ;
      RECT  114.77 103.905 114.98 103.7 ;
      RECT  117.89 104.285 118.1 103.905 ;
      RECT  116.81 103.7 116.99 101.995 ;
      RECT  114.98 103.905 115.19 103.7 ;
      RECT  114.77 104.285 114.98 103.905 ;
      POLYGON  117.38 102.62 117.38 102.21 117.635 102.21 117.635 102.54 117.555 102.62 117.38 102.62 ;
      RECT  115.37 104.615 115.55 103.7 ;
      RECT  114.98 104.615 115.19 104.285 ;
      RECT  114.98 104.285 115.19 103.905 ;
      RECT  117.17 104.58 117.38 104.99 ;
      RECT  114.77 103.575 114.98 103.905 ;
      RECT  117.815 104.49 117.89 106.195 ;
      RECT  117.73 105.075 117.815 105.485 ;
      RECT  116.81 103.575 116.99 104.49 ;
      POLYGON  117.815 103.575 117.815 103.905 117.38 103.905 117.38 104.285 117.815 104.285 117.815 104.49 117.89 104.49 117.89 103.575 117.815 103.575 ;
      RECT  117.89 104.49 118.1 106.195 ;
      POLYGON  117.38 104.58 117.38 104.99 117.555 104.99 117.635 104.91 117.635 104.58 117.38 104.58 ;
      RECT  114.77 104.49 114.98 106.195 ;
      RECT  116.45 103.575 116.63 104.49 ;
      RECT  115.37 104.49 115.55 106.195 ;
      RECT  117.17 105.57 117.38 105.98 ;
      RECT  117.89 104.285 118.1 104.49 ;
      RECT  114.98 104.49 115.19 106.195 ;
      RECT  117.17 103.905 117.38 104.285 ;
      RECT  115.73 104.49 115.91 106.195 ;
      RECT  116.45 104.49 116.63 106.195 ;
      RECT  115.73 103.575 115.91 104.49 ;
      RECT  117.89 103.575 118.1 103.905 ;
      RECT  116.09 104.49 116.27 106.195 ;
      RECT  116.09 103.575 116.27 104.49 ;
      RECT  114.77 104.285 114.98 104.49 ;
      RECT  117.89 103.905 118.1 104.285 ;
      RECT  116.81 104.49 116.99 106.195 ;
      RECT  114.98 104.285 115.19 104.49 ;
      RECT  114.77 103.905 114.98 104.285 ;
      POLYGON  117.38 105.57 117.38 105.98 117.635 105.98 117.635 105.65 117.555 105.57 117.38 105.57 ;
      RECT  115.37 103.575 115.55 104.49 ;
      RECT  114.98 103.575 115.19 103.905 ;
      RECT  114.98 103.905 115.19 104.285 ;
      RECT  117.17 107.56 117.38 107.15 ;
      RECT  114.77 108.565 114.98 108.235 ;
      RECT  117.815 107.65 117.89 105.945 ;
      RECT  117.73 107.065 117.815 106.655 ;
      RECT  116.81 108.565 116.99 107.65 ;
      POLYGON  117.815 108.565 117.815 108.235 117.38 108.235 117.38 107.855 117.815 107.855 117.815 107.65 117.89 107.65 117.89 108.565 117.815 108.565 ;
      RECT  117.89 107.65 118.1 105.945 ;
      POLYGON  117.38 107.56 117.38 107.15 117.555 107.15 117.635 107.23 117.635 107.56 117.38 107.56 ;
      RECT  114.77 107.65 114.98 105.945 ;
      RECT  116.45 108.565 116.63 107.65 ;
      RECT  115.37 107.65 115.55 105.945 ;
      RECT  117.17 106.57 117.38 106.16 ;
      RECT  117.89 107.855 118.1 107.65 ;
      RECT  114.98 107.65 115.19 105.945 ;
      RECT  117.17 108.235 117.38 107.855 ;
      RECT  115.73 107.65 115.91 105.945 ;
      RECT  116.45 107.65 116.63 105.945 ;
      RECT  115.73 108.565 115.91 107.65 ;
      RECT  117.89 108.565 118.1 108.235 ;
      RECT  116.09 107.65 116.27 105.945 ;
      RECT  116.09 108.565 116.27 107.65 ;
      RECT  114.77 107.855 114.98 107.65 ;
      RECT  117.89 108.235 118.1 107.855 ;
      RECT  116.81 107.65 116.99 105.945 ;
      RECT  114.98 107.855 115.19 107.65 ;
      RECT  114.77 108.235 114.98 107.855 ;
      POLYGON  117.38 106.57 117.38 106.16 117.635 106.16 117.635 106.49 117.555 106.57 117.38 106.57 ;
      RECT  115.37 108.565 115.55 107.65 ;
      RECT  114.98 108.565 115.19 108.235 ;
      RECT  114.98 108.235 115.19 107.855 ;
      RECT  117.17 108.53 117.38 108.94 ;
      RECT  114.77 107.525 114.98 107.855 ;
      RECT  117.815 108.44 117.89 110.145 ;
      RECT  117.73 109.025 117.815 109.435 ;
      RECT  116.81 107.525 116.99 108.44 ;
      POLYGON  117.815 107.525 117.815 107.855 117.38 107.855 117.38 108.235 117.815 108.235 117.815 108.44 117.89 108.44 117.89 107.525 117.815 107.525 ;
      RECT  117.89 108.44 118.1 110.145 ;
      POLYGON  117.38 108.53 117.38 108.94 117.555 108.94 117.635 108.86 117.635 108.53 117.38 108.53 ;
      RECT  114.77 108.44 114.98 110.145 ;
      RECT  116.45 107.525 116.63 108.44 ;
      RECT  115.37 108.44 115.55 110.145 ;
      RECT  117.17 109.52 117.38 109.93 ;
      RECT  117.89 108.235 118.1 108.44 ;
      RECT  114.98 108.44 115.19 110.145 ;
      RECT  117.17 107.855 117.38 108.235 ;
      RECT  115.73 108.44 115.91 110.145 ;
      RECT  116.45 108.44 116.63 110.145 ;
      RECT  115.73 107.525 115.91 108.44 ;
      RECT  117.89 107.525 118.1 107.855 ;
      RECT  116.09 108.44 116.27 110.145 ;
      RECT  116.09 107.525 116.27 108.44 ;
      RECT  114.77 108.235 114.98 108.44 ;
      RECT  117.89 107.855 118.1 108.235 ;
      RECT  116.81 108.44 116.99 110.145 ;
      RECT  114.98 108.235 115.19 108.44 ;
      RECT  114.77 107.855 114.98 108.235 ;
      POLYGON  117.38 109.52 117.38 109.93 117.635 109.93 117.635 109.6 117.555 109.52 117.38 109.52 ;
      RECT  115.37 107.525 115.55 108.44 ;
      RECT  114.98 107.525 115.19 107.855 ;
      RECT  114.98 107.855 115.19 108.235 ;
      RECT  117.17 111.51 117.38 111.1 ;
      RECT  114.77 112.515 114.98 112.185 ;
      RECT  117.815 111.6 117.89 109.895 ;
      RECT  117.73 111.015 117.815 110.605 ;
      RECT  116.81 112.515 116.99 111.6 ;
      POLYGON  117.815 112.515 117.815 112.185 117.38 112.185 117.38 111.805 117.815 111.805 117.815 111.6 117.89 111.6 117.89 112.515 117.815 112.515 ;
      RECT  117.89 111.6 118.1 109.895 ;
      POLYGON  117.38 111.51 117.38 111.1 117.555 111.1 117.635 111.18 117.635 111.51 117.38 111.51 ;
      RECT  114.77 111.6 114.98 109.895 ;
      RECT  116.45 112.515 116.63 111.6 ;
      RECT  115.37 111.6 115.55 109.895 ;
      RECT  117.17 110.52 117.38 110.11 ;
      RECT  117.89 111.805 118.1 111.6 ;
      RECT  114.98 111.6 115.19 109.895 ;
      RECT  117.17 112.185 117.38 111.805 ;
      RECT  115.73 111.6 115.91 109.895 ;
      RECT  116.45 111.6 116.63 109.895 ;
      RECT  115.73 112.515 115.91 111.6 ;
      RECT  117.89 112.515 118.1 112.185 ;
      RECT  116.09 111.6 116.27 109.895 ;
      RECT  116.09 112.515 116.27 111.6 ;
      RECT  114.77 111.805 114.98 111.6 ;
      RECT  117.89 112.185 118.1 111.805 ;
      RECT  116.81 111.6 116.99 109.895 ;
      RECT  114.98 111.805 115.19 111.6 ;
      RECT  114.77 112.185 114.98 111.805 ;
      POLYGON  117.38 110.52 117.38 110.11 117.635 110.11 117.635 110.44 117.555 110.52 117.38 110.52 ;
      RECT  115.37 112.515 115.55 111.6 ;
      RECT  114.98 112.515 115.19 112.185 ;
      RECT  114.98 112.185 115.19 111.805 ;
      RECT  117.17 112.48 117.38 112.89 ;
      RECT  114.77 111.475 114.98 111.805 ;
      RECT  117.815 112.39 117.89 114.095 ;
      RECT  117.73 112.975 117.815 113.385 ;
      RECT  116.81 111.475 116.99 112.39 ;
      POLYGON  117.815 111.475 117.815 111.805 117.38 111.805 117.38 112.185 117.815 112.185 117.815 112.39 117.89 112.39 117.89 111.475 117.815 111.475 ;
      RECT  117.89 112.39 118.1 114.095 ;
      POLYGON  117.38 112.48 117.38 112.89 117.555 112.89 117.635 112.81 117.635 112.48 117.38 112.48 ;
      RECT  114.77 112.39 114.98 114.095 ;
      RECT  116.45 111.475 116.63 112.39 ;
      RECT  115.37 112.39 115.55 114.095 ;
      RECT  117.17 113.47 117.38 113.88 ;
      RECT  117.89 112.185 118.1 112.39 ;
      RECT  114.98 112.39 115.19 114.095 ;
      RECT  117.17 111.805 117.38 112.185 ;
      RECT  115.73 112.39 115.91 114.095 ;
      RECT  116.45 112.39 116.63 114.095 ;
      RECT  115.73 111.475 115.91 112.39 ;
      RECT  117.89 111.475 118.1 111.805 ;
      RECT  116.09 112.39 116.27 114.095 ;
      RECT  116.09 111.475 116.27 112.39 ;
      RECT  114.77 112.185 114.98 112.39 ;
      RECT  117.89 111.805 118.1 112.185 ;
      RECT  116.81 112.39 116.99 114.095 ;
      RECT  114.98 112.185 115.19 112.39 ;
      RECT  114.77 111.805 114.98 112.185 ;
      POLYGON  117.38 113.47 117.38 113.88 117.635 113.88 117.635 113.55 117.555 113.47 117.38 113.47 ;
      RECT  115.37 111.475 115.55 112.39 ;
      RECT  114.98 111.475 115.19 111.805 ;
      RECT  114.98 111.805 115.19 112.185 ;
      RECT  117.17 115.46 117.38 115.05 ;
      RECT  114.77 116.465 114.98 116.135 ;
      RECT  117.815 115.55 117.89 113.845 ;
      RECT  117.73 114.965 117.815 114.555 ;
      RECT  116.81 116.465 116.99 115.55 ;
      POLYGON  117.815 116.465 117.815 116.135 117.38 116.135 117.38 115.755 117.815 115.755 117.815 115.55 117.89 115.55 117.89 116.465 117.815 116.465 ;
      RECT  117.89 115.55 118.1 113.845 ;
      POLYGON  117.38 115.46 117.38 115.05 117.555 115.05 117.635 115.13 117.635 115.46 117.38 115.46 ;
      RECT  114.77 115.55 114.98 113.845 ;
      RECT  116.45 116.465 116.63 115.55 ;
      RECT  115.37 115.55 115.55 113.845 ;
      RECT  117.17 114.47 117.38 114.06 ;
      RECT  117.89 115.755 118.1 115.55 ;
      RECT  114.98 115.55 115.19 113.845 ;
      RECT  117.17 116.135 117.38 115.755 ;
      RECT  115.73 115.55 115.91 113.845 ;
      RECT  116.45 115.55 116.63 113.845 ;
      RECT  115.73 116.465 115.91 115.55 ;
      RECT  117.89 116.465 118.1 116.135 ;
      RECT  116.09 115.55 116.27 113.845 ;
      RECT  116.09 116.465 116.27 115.55 ;
      RECT  114.77 115.755 114.98 115.55 ;
      RECT  117.89 116.135 118.1 115.755 ;
      RECT  116.81 115.55 116.99 113.845 ;
      RECT  114.98 115.755 115.19 115.55 ;
      RECT  114.77 116.135 114.98 115.755 ;
      POLYGON  117.38 114.47 117.38 114.06 117.635 114.06 117.635 114.39 117.555 114.47 117.38 114.47 ;
      RECT  115.37 116.465 115.55 115.55 ;
      RECT  114.98 116.465 115.19 116.135 ;
      RECT  114.98 116.135 115.19 115.755 ;
      RECT  117.17 116.43 117.38 116.84 ;
      RECT  114.77 115.425 114.98 115.755 ;
      RECT  117.815 116.34 117.89 118.045 ;
      RECT  117.73 116.925 117.815 117.335 ;
      RECT  116.81 115.425 116.99 116.34 ;
      POLYGON  117.815 115.425 117.815 115.755 117.38 115.755 117.38 116.135 117.815 116.135 117.815 116.34 117.89 116.34 117.89 115.425 117.815 115.425 ;
      RECT  117.89 116.34 118.1 118.045 ;
      POLYGON  117.38 116.43 117.38 116.84 117.555 116.84 117.635 116.76 117.635 116.43 117.38 116.43 ;
      RECT  114.77 116.34 114.98 118.045 ;
      RECT  116.45 115.425 116.63 116.34 ;
      RECT  115.37 116.34 115.55 118.045 ;
      RECT  117.17 117.42 117.38 117.83 ;
      RECT  117.89 116.135 118.1 116.34 ;
      RECT  114.98 116.34 115.19 118.045 ;
      RECT  117.17 115.755 117.38 116.135 ;
      RECT  115.73 116.34 115.91 118.045 ;
      RECT  116.45 116.34 116.63 118.045 ;
      RECT  115.73 115.425 115.91 116.34 ;
      RECT  117.89 115.425 118.1 115.755 ;
      RECT  116.09 116.34 116.27 118.045 ;
      RECT  116.09 115.425 116.27 116.34 ;
      RECT  114.77 116.135 114.98 116.34 ;
      RECT  117.89 115.755 118.1 116.135 ;
      RECT  116.81 116.34 116.99 118.045 ;
      RECT  114.98 116.135 115.19 116.34 ;
      RECT  114.77 115.755 114.98 116.135 ;
      POLYGON  117.38 117.42 117.38 117.83 117.635 117.83 117.635 117.5 117.555 117.42 117.38 117.42 ;
      RECT  115.37 115.425 115.55 116.34 ;
      RECT  114.98 115.425 115.19 115.755 ;
      RECT  114.98 115.755 115.19 116.135 ;
      RECT  117.17 119.41 117.38 119.0 ;
      RECT  114.77 120.415 114.98 120.085 ;
      RECT  117.815 119.5 117.89 117.795 ;
      RECT  117.73 118.915 117.815 118.505 ;
      RECT  116.81 120.415 116.99 119.5 ;
      POLYGON  117.815 120.415 117.815 120.085 117.38 120.085 117.38 119.705 117.815 119.705 117.815 119.5 117.89 119.5 117.89 120.415 117.815 120.415 ;
      RECT  117.89 119.5 118.1 117.795 ;
      POLYGON  117.38 119.41 117.38 119.0 117.555 119.0 117.635 119.08 117.635 119.41 117.38 119.41 ;
      RECT  114.77 119.5 114.98 117.795 ;
      RECT  116.45 120.415 116.63 119.5 ;
      RECT  115.37 119.5 115.55 117.795 ;
      RECT  117.17 118.42 117.38 118.01 ;
      RECT  117.89 119.705 118.1 119.5 ;
      RECT  114.98 119.5 115.19 117.795 ;
      RECT  117.17 120.085 117.38 119.705 ;
      RECT  115.73 119.5 115.91 117.795 ;
      RECT  116.45 119.5 116.63 117.795 ;
      RECT  115.73 120.415 115.91 119.5 ;
      RECT  117.89 120.415 118.1 120.085 ;
      RECT  116.09 119.5 116.27 117.795 ;
      RECT  116.09 120.415 116.27 119.5 ;
      RECT  114.77 119.705 114.98 119.5 ;
      RECT  117.89 120.085 118.1 119.705 ;
      RECT  116.81 119.5 116.99 117.795 ;
      RECT  114.98 119.705 115.19 119.5 ;
      RECT  114.77 120.085 114.98 119.705 ;
      POLYGON  117.38 118.42 117.38 118.01 117.635 118.01 117.635 118.34 117.555 118.42 117.38 118.42 ;
      RECT  115.37 120.415 115.55 119.5 ;
      RECT  114.98 120.415 115.19 120.085 ;
      RECT  114.98 120.085 115.19 119.705 ;
      RECT  117.17 120.38 117.38 120.79 ;
      RECT  114.77 119.375 114.98 119.705 ;
      RECT  117.815 120.29 117.89 121.995 ;
      RECT  117.73 120.875 117.815 121.285 ;
      RECT  116.81 119.375 116.99 120.29 ;
      POLYGON  117.815 119.375 117.815 119.705 117.38 119.705 117.38 120.085 117.815 120.085 117.815 120.29 117.89 120.29 117.89 119.375 117.815 119.375 ;
      RECT  117.89 120.29 118.1 121.995 ;
      POLYGON  117.38 120.38 117.38 120.79 117.555 120.79 117.635 120.71 117.635 120.38 117.38 120.38 ;
      RECT  114.77 120.29 114.98 121.995 ;
      RECT  116.45 119.375 116.63 120.29 ;
      RECT  115.37 120.29 115.55 121.995 ;
      RECT  117.17 121.37 117.38 121.78 ;
      RECT  117.89 120.085 118.1 120.29 ;
      RECT  114.98 120.29 115.19 121.995 ;
      RECT  117.17 119.705 117.38 120.085 ;
      RECT  115.73 120.29 115.91 121.995 ;
      RECT  116.45 120.29 116.63 121.995 ;
      RECT  115.73 119.375 115.91 120.29 ;
      RECT  117.89 119.375 118.1 119.705 ;
      RECT  116.09 120.29 116.27 121.995 ;
      RECT  116.09 119.375 116.27 120.29 ;
      RECT  114.77 120.085 114.98 120.29 ;
      RECT  117.89 119.705 118.1 120.085 ;
      RECT  116.81 120.29 116.99 121.995 ;
      RECT  114.98 120.085 115.19 120.29 ;
      RECT  114.77 119.705 114.98 120.085 ;
      POLYGON  117.38 121.37 117.38 121.78 117.635 121.78 117.635 121.45 117.555 121.37 117.38 121.37 ;
      RECT  115.37 119.375 115.55 120.29 ;
      RECT  114.98 119.375 115.19 119.705 ;
      RECT  114.98 119.705 115.19 120.085 ;
      RECT  117.17 123.36 117.38 122.95 ;
      RECT  114.77 124.365 114.98 124.035 ;
      RECT  117.815 123.45 117.89 121.745 ;
      RECT  117.73 122.865 117.815 122.455 ;
      RECT  116.81 124.365 116.99 123.45 ;
      POLYGON  117.815 124.365 117.815 124.035 117.38 124.035 117.38 123.655 117.815 123.655 117.815 123.45 117.89 123.45 117.89 124.365 117.815 124.365 ;
      RECT  117.89 123.45 118.1 121.745 ;
      POLYGON  117.38 123.36 117.38 122.95 117.555 122.95 117.635 123.03 117.635 123.36 117.38 123.36 ;
      RECT  114.77 123.45 114.98 121.745 ;
      RECT  116.45 124.365 116.63 123.45 ;
      RECT  115.37 123.45 115.55 121.745 ;
      RECT  117.17 122.37 117.38 121.96 ;
      RECT  117.89 123.655 118.1 123.45 ;
      RECT  114.98 123.45 115.19 121.745 ;
      RECT  117.17 124.035 117.38 123.655 ;
      RECT  115.73 123.45 115.91 121.745 ;
      RECT  116.45 123.45 116.63 121.745 ;
      RECT  115.73 124.365 115.91 123.45 ;
      RECT  117.89 124.365 118.1 124.035 ;
      RECT  116.09 123.45 116.27 121.745 ;
      RECT  116.09 124.365 116.27 123.45 ;
      RECT  114.77 123.655 114.98 123.45 ;
      RECT  117.89 124.035 118.1 123.655 ;
      RECT  116.81 123.45 116.99 121.745 ;
      RECT  114.98 123.655 115.19 123.45 ;
      RECT  114.77 124.035 114.98 123.655 ;
      POLYGON  117.38 122.37 117.38 121.96 117.635 121.96 117.635 122.29 117.555 122.37 117.38 122.37 ;
      RECT  115.37 124.365 115.55 123.45 ;
      RECT  114.98 124.365 115.19 124.035 ;
      RECT  114.98 124.035 115.19 123.655 ;
      RECT  119.03 92.73 118.82 93.14 ;
      RECT  121.43 91.725 121.22 92.055 ;
      RECT  118.385 92.64 118.31 94.345 ;
      RECT  118.47 93.225 118.385 93.635 ;
      RECT  119.39 91.725 119.21 92.64 ;
      POLYGON  118.385 91.725 118.385 92.055 118.82 92.055 118.82 92.435 118.385 92.435 118.385 92.64 118.31 92.64 118.31 91.725 118.385 91.725 ;
      RECT  118.31 92.64 118.1 94.345 ;
      POLYGON  118.82 92.73 118.82 93.14 118.645 93.14 118.565 93.06 118.565 92.73 118.82 92.73 ;
      RECT  121.43 92.64 121.22 94.345 ;
      RECT  119.75 91.725 119.57 92.64 ;
      RECT  120.83 92.64 120.65 94.345 ;
      RECT  119.03 93.72 118.82 94.13 ;
      RECT  118.31 92.435 118.1 92.64 ;
      RECT  121.22 92.64 121.01 94.345 ;
      RECT  119.03 92.055 118.82 92.435 ;
      RECT  120.47 92.64 120.29 94.345 ;
      RECT  119.75 92.64 119.57 94.345 ;
      RECT  120.47 91.725 120.29 92.64 ;
      RECT  118.31 91.725 118.1 92.055 ;
      RECT  120.11 92.64 119.93 94.345 ;
      RECT  120.11 91.725 119.93 92.64 ;
      RECT  121.43 92.435 121.22 92.64 ;
      RECT  118.31 92.055 118.1 92.435 ;
      RECT  119.39 92.64 119.21 94.345 ;
      RECT  121.22 92.435 121.01 92.64 ;
      RECT  121.43 92.055 121.22 92.435 ;
      POLYGON  118.82 93.72 118.82 94.13 118.565 94.13 118.565 93.8 118.645 93.72 118.82 93.72 ;
      RECT  120.83 91.725 120.65 92.64 ;
      RECT  121.22 91.725 121.01 92.055 ;
      RECT  121.22 92.055 121.01 92.435 ;
      RECT  119.03 95.71 118.82 95.3 ;
      RECT  121.43 96.715 121.22 96.385 ;
      RECT  118.385 95.8 118.31 94.095 ;
      RECT  118.47 95.215 118.385 94.805 ;
      RECT  119.39 96.715 119.21 95.8 ;
      POLYGON  118.385 96.715 118.385 96.385 118.82 96.385 118.82 96.005 118.385 96.005 118.385 95.8 118.31 95.8 118.31 96.715 118.385 96.715 ;
      RECT  118.31 95.8 118.1 94.095 ;
      POLYGON  118.82 95.71 118.82 95.3 118.645 95.3 118.565 95.38 118.565 95.71 118.82 95.71 ;
      RECT  121.43 95.8 121.22 94.095 ;
      RECT  119.75 96.715 119.57 95.8 ;
      RECT  120.83 95.8 120.65 94.095 ;
      RECT  119.03 94.72 118.82 94.31 ;
      RECT  118.31 96.005 118.1 95.8 ;
      RECT  121.22 95.8 121.01 94.095 ;
      RECT  119.03 96.385 118.82 96.005 ;
      RECT  120.47 95.8 120.29 94.095 ;
      RECT  119.75 95.8 119.57 94.095 ;
      RECT  120.47 96.715 120.29 95.8 ;
      RECT  118.31 96.715 118.1 96.385 ;
      RECT  120.11 95.8 119.93 94.095 ;
      RECT  120.11 96.715 119.93 95.8 ;
      RECT  121.43 96.005 121.22 95.8 ;
      RECT  118.31 96.385 118.1 96.005 ;
      RECT  119.39 95.8 119.21 94.095 ;
      RECT  121.22 96.005 121.01 95.8 ;
      RECT  121.43 96.385 121.22 96.005 ;
      POLYGON  118.82 94.72 118.82 94.31 118.565 94.31 118.565 94.64 118.645 94.72 118.82 94.72 ;
      RECT  120.83 96.715 120.65 95.8 ;
      RECT  121.22 96.715 121.01 96.385 ;
      RECT  121.22 96.385 121.01 96.005 ;
      RECT  119.03 96.68 118.82 97.09 ;
      RECT  121.43 95.675 121.22 96.005 ;
      RECT  118.385 96.59 118.31 98.295 ;
      RECT  118.47 97.175 118.385 97.585 ;
      RECT  119.39 95.675 119.21 96.59 ;
      POLYGON  118.385 95.675 118.385 96.005 118.82 96.005 118.82 96.385 118.385 96.385 118.385 96.59 118.31 96.59 118.31 95.675 118.385 95.675 ;
      RECT  118.31 96.59 118.1 98.295 ;
      POLYGON  118.82 96.68 118.82 97.09 118.645 97.09 118.565 97.01 118.565 96.68 118.82 96.68 ;
      RECT  121.43 96.59 121.22 98.295 ;
      RECT  119.75 95.675 119.57 96.59 ;
      RECT  120.83 96.59 120.65 98.295 ;
      RECT  119.03 97.67 118.82 98.08 ;
      RECT  118.31 96.385 118.1 96.59 ;
      RECT  121.22 96.59 121.01 98.295 ;
      RECT  119.03 96.005 118.82 96.385 ;
      RECT  120.47 96.59 120.29 98.295 ;
      RECT  119.75 96.59 119.57 98.295 ;
      RECT  120.47 95.675 120.29 96.59 ;
      RECT  118.31 95.675 118.1 96.005 ;
      RECT  120.11 96.59 119.93 98.295 ;
      RECT  120.11 95.675 119.93 96.59 ;
      RECT  121.43 96.385 121.22 96.59 ;
      RECT  118.31 96.005 118.1 96.385 ;
      RECT  119.39 96.59 119.21 98.295 ;
      RECT  121.22 96.385 121.01 96.59 ;
      RECT  121.43 96.005 121.22 96.385 ;
      POLYGON  118.82 97.67 118.82 98.08 118.565 98.08 118.565 97.75 118.645 97.67 118.82 97.67 ;
      RECT  120.83 95.675 120.65 96.59 ;
      RECT  121.22 95.675 121.01 96.005 ;
      RECT  121.22 96.005 121.01 96.385 ;
      RECT  119.03 99.66 118.82 99.25 ;
      RECT  121.43 100.665 121.22 100.335 ;
      RECT  118.385 99.75 118.31 98.045 ;
      RECT  118.47 99.165 118.385 98.755 ;
      RECT  119.39 100.665 119.21 99.75 ;
      POLYGON  118.385 100.665 118.385 100.335 118.82 100.335 118.82 99.955 118.385 99.955 118.385 99.75 118.31 99.75 118.31 100.665 118.385 100.665 ;
      RECT  118.31 99.75 118.1 98.045 ;
      POLYGON  118.82 99.66 118.82 99.25 118.645 99.25 118.565 99.33 118.565 99.66 118.82 99.66 ;
      RECT  121.43 99.75 121.22 98.045 ;
      RECT  119.75 100.665 119.57 99.75 ;
      RECT  120.83 99.75 120.65 98.045 ;
      RECT  119.03 98.67 118.82 98.26 ;
      RECT  118.31 99.955 118.1 99.75 ;
      RECT  121.22 99.75 121.01 98.045 ;
      RECT  119.03 100.335 118.82 99.955 ;
      RECT  120.47 99.75 120.29 98.045 ;
      RECT  119.75 99.75 119.57 98.045 ;
      RECT  120.47 100.665 120.29 99.75 ;
      RECT  118.31 100.665 118.1 100.335 ;
      RECT  120.11 99.75 119.93 98.045 ;
      RECT  120.11 100.665 119.93 99.75 ;
      RECT  121.43 99.955 121.22 99.75 ;
      RECT  118.31 100.335 118.1 99.955 ;
      RECT  119.39 99.75 119.21 98.045 ;
      RECT  121.22 99.955 121.01 99.75 ;
      RECT  121.43 100.335 121.22 99.955 ;
      POLYGON  118.82 98.67 118.82 98.26 118.565 98.26 118.565 98.59 118.645 98.67 118.82 98.67 ;
      RECT  120.83 100.665 120.65 99.75 ;
      RECT  121.22 100.665 121.01 100.335 ;
      RECT  121.22 100.335 121.01 99.955 ;
      RECT  119.03 100.63 118.82 101.04 ;
      RECT  121.43 99.625 121.22 99.955 ;
      RECT  118.385 100.54 118.31 102.245 ;
      RECT  118.47 101.125 118.385 101.535 ;
      RECT  119.39 99.625 119.21 100.54 ;
      POLYGON  118.385 99.625 118.385 99.955 118.82 99.955 118.82 100.335 118.385 100.335 118.385 100.54 118.31 100.54 118.31 99.625 118.385 99.625 ;
      RECT  118.31 100.54 118.1 102.245 ;
      POLYGON  118.82 100.63 118.82 101.04 118.645 101.04 118.565 100.96 118.565 100.63 118.82 100.63 ;
      RECT  121.43 100.54 121.22 102.245 ;
      RECT  119.75 99.625 119.57 100.54 ;
      RECT  120.83 100.54 120.65 102.245 ;
      RECT  119.03 101.62 118.82 102.03 ;
      RECT  118.31 100.335 118.1 100.54 ;
      RECT  121.22 100.54 121.01 102.245 ;
      RECT  119.03 99.955 118.82 100.335 ;
      RECT  120.47 100.54 120.29 102.245 ;
      RECT  119.75 100.54 119.57 102.245 ;
      RECT  120.47 99.625 120.29 100.54 ;
      RECT  118.31 99.625 118.1 99.955 ;
      RECT  120.11 100.54 119.93 102.245 ;
      RECT  120.11 99.625 119.93 100.54 ;
      RECT  121.43 100.335 121.22 100.54 ;
      RECT  118.31 99.955 118.1 100.335 ;
      RECT  119.39 100.54 119.21 102.245 ;
      RECT  121.22 100.335 121.01 100.54 ;
      RECT  121.43 99.955 121.22 100.335 ;
      POLYGON  118.82 101.62 118.82 102.03 118.565 102.03 118.565 101.7 118.645 101.62 118.82 101.62 ;
      RECT  120.83 99.625 120.65 100.54 ;
      RECT  121.22 99.625 121.01 99.955 ;
      RECT  121.22 99.955 121.01 100.335 ;
      RECT  119.03 103.61 118.82 103.2 ;
      RECT  121.43 104.615 121.22 104.285 ;
      RECT  118.385 103.7 118.31 101.995 ;
      RECT  118.47 103.115 118.385 102.705 ;
      RECT  119.39 104.615 119.21 103.7 ;
      POLYGON  118.385 104.615 118.385 104.285 118.82 104.285 118.82 103.905 118.385 103.905 118.385 103.7 118.31 103.7 118.31 104.615 118.385 104.615 ;
      RECT  118.31 103.7 118.1 101.995 ;
      POLYGON  118.82 103.61 118.82 103.2 118.645 103.2 118.565 103.28 118.565 103.61 118.82 103.61 ;
      RECT  121.43 103.7 121.22 101.995 ;
      RECT  119.75 104.615 119.57 103.7 ;
      RECT  120.83 103.7 120.65 101.995 ;
      RECT  119.03 102.62 118.82 102.21 ;
      RECT  118.31 103.905 118.1 103.7 ;
      RECT  121.22 103.7 121.01 101.995 ;
      RECT  119.03 104.285 118.82 103.905 ;
      RECT  120.47 103.7 120.29 101.995 ;
      RECT  119.75 103.7 119.57 101.995 ;
      RECT  120.47 104.615 120.29 103.7 ;
      RECT  118.31 104.615 118.1 104.285 ;
      RECT  120.11 103.7 119.93 101.995 ;
      RECT  120.11 104.615 119.93 103.7 ;
      RECT  121.43 103.905 121.22 103.7 ;
      RECT  118.31 104.285 118.1 103.905 ;
      RECT  119.39 103.7 119.21 101.995 ;
      RECT  121.22 103.905 121.01 103.7 ;
      RECT  121.43 104.285 121.22 103.905 ;
      POLYGON  118.82 102.62 118.82 102.21 118.565 102.21 118.565 102.54 118.645 102.62 118.82 102.62 ;
      RECT  120.83 104.615 120.65 103.7 ;
      RECT  121.22 104.615 121.01 104.285 ;
      RECT  121.22 104.285 121.01 103.905 ;
      RECT  119.03 104.58 118.82 104.99 ;
      RECT  121.43 103.575 121.22 103.905 ;
      RECT  118.385 104.49 118.31 106.195 ;
      RECT  118.47 105.075 118.385 105.485 ;
      RECT  119.39 103.575 119.21 104.49 ;
      POLYGON  118.385 103.575 118.385 103.905 118.82 103.905 118.82 104.285 118.385 104.285 118.385 104.49 118.31 104.49 118.31 103.575 118.385 103.575 ;
      RECT  118.31 104.49 118.1 106.195 ;
      POLYGON  118.82 104.58 118.82 104.99 118.645 104.99 118.565 104.91 118.565 104.58 118.82 104.58 ;
      RECT  121.43 104.49 121.22 106.195 ;
      RECT  119.75 103.575 119.57 104.49 ;
      RECT  120.83 104.49 120.65 106.195 ;
      RECT  119.03 105.57 118.82 105.98 ;
      RECT  118.31 104.285 118.1 104.49 ;
      RECT  121.22 104.49 121.01 106.195 ;
      RECT  119.03 103.905 118.82 104.285 ;
      RECT  120.47 104.49 120.29 106.195 ;
      RECT  119.75 104.49 119.57 106.195 ;
      RECT  120.47 103.575 120.29 104.49 ;
      RECT  118.31 103.575 118.1 103.905 ;
      RECT  120.11 104.49 119.93 106.195 ;
      RECT  120.11 103.575 119.93 104.49 ;
      RECT  121.43 104.285 121.22 104.49 ;
      RECT  118.31 103.905 118.1 104.285 ;
      RECT  119.39 104.49 119.21 106.195 ;
      RECT  121.22 104.285 121.01 104.49 ;
      RECT  121.43 103.905 121.22 104.285 ;
      POLYGON  118.82 105.57 118.82 105.98 118.565 105.98 118.565 105.65 118.645 105.57 118.82 105.57 ;
      RECT  120.83 103.575 120.65 104.49 ;
      RECT  121.22 103.575 121.01 103.905 ;
      RECT  121.22 103.905 121.01 104.285 ;
      RECT  119.03 107.56 118.82 107.15 ;
      RECT  121.43 108.565 121.22 108.235 ;
      RECT  118.385 107.65 118.31 105.945 ;
      RECT  118.47 107.065 118.385 106.655 ;
      RECT  119.39 108.565 119.21 107.65 ;
      POLYGON  118.385 108.565 118.385 108.235 118.82 108.235 118.82 107.855 118.385 107.855 118.385 107.65 118.31 107.65 118.31 108.565 118.385 108.565 ;
      RECT  118.31 107.65 118.1 105.945 ;
      POLYGON  118.82 107.56 118.82 107.15 118.645 107.15 118.565 107.23 118.565 107.56 118.82 107.56 ;
      RECT  121.43 107.65 121.22 105.945 ;
      RECT  119.75 108.565 119.57 107.65 ;
      RECT  120.83 107.65 120.65 105.945 ;
      RECT  119.03 106.57 118.82 106.16 ;
      RECT  118.31 107.855 118.1 107.65 ;
      RECT  121.22 107.65 121.01 105.945 ;
      RECT  119.03 108.235 118.82 107.855 ;
      RECT  120.47 107.65 120.29 105.945 ;
      RECT  119.75 107.65 119.57 105.945 ;
      RECT  120.47 108.565 120.29 107.65 ;
      RECT  118.31 108.565 118.1 108.235 ;
      RECT  120.11 107.65 119.93 105.945 ;
      RECT  120.11 108.565 119.93 107.65 ;
      RECT  121.43 107.855 121.22 107.65 ;
      RECT  118.31 108.235 118.1 107.855 ;
      RECT  119.39 107.65 119.21 105.945 ;
      RECT  121.22 107.855 121.01 107.65 ;
      RECT  121.43 108.235 121.22 107.855 ;
      POLYGON  118.82 106.57 118.82 106.16 118.565 106.16 118.565 106.49 118.645 106.57 118.82 106.57 ;
      RECT  120.83 108.565 120.65 107.65 ;
      RECT  121.22 108.565 121.01 108.235 ;
      RECT  121.22 108.235 121.01 107.855 ;
      RECT  119.03 108.53 118.82 108.94 ;
      RECT  121.43 107.525 121.22 107.855 ;
      RECT  118.385 108.44 118.31 110.145 ;
      RECT  118.47 109.025 118.385 109.435 ;
      RECT  119.39 107.525 119.21 108.44 ;
      POLYGON  118.385 107.525 118.385 107.855 118.82 107.855 118.82 108.235 118.385 108.235 118.385 108.44 118.31 108.44 118.31 107.525 118.385 107.525 ;
      RECT  118.31 108.44 118.1 110.145 ;
      POLYGON  118.82 108.53 118.82 108.94 118.645 108.94 118.565 108.86 118.565 108.53 118.82 108.53 ;
      RECT  121.43 108.44 121.22 110.145 ;
      RECT  119.75 107.525 119.57 108.44 ;
      RECT  120.83 108.44 120.65 110.145 ;
      RECT  119.03 109.52 118.82 109.93 ;
      RECT  118.31 108.235 118.1 108.44 ;
      RECT  121.22 108.44 121.01 110.145 ;
      RECT  119.03 107.855 118.82 108.235 ;
      RECT  120.47 108.44 120.29 110.145 ;
      RECT  119.75 108.44 119.57 110.145 ;
      RECT  120.47 107.525 120.29 108.44 ;
      RECT  118.31 107.525 118.1 107.855 ;
      RECT  120.11 108.44 119.93 110.145 ;
      RECT  120.11 107.525 119.93 108.44 ;
      RECT  121.43 108.235 121.22 108.44 ;
      RECT  118.31 107.855 118.1 108.235 ;
      RECT  119.39 108.44 119.21 110.145 ;
      RECT  121.22 108.235 121.01 108.44 ;
      RECT  121.43 107.855 121.22 108.235 ;
      POLYGON  118.82 109.52 118.82 109.93 118.565 109.93 118.565 109.6 118.645 109.52 118.82 109.52 ;
      RECT  120.83 107.525 120.65 108.44 ;
      RECT  121.22 107.525 121.01 107.855 ;
      RECT  121.22 107.855 121.01 108.235 ;
      RECT  119.03 111.51 118.82 111.1 ;
      RECT  121.43 112.515 121.22 112.185 ;
      RECT  118.385 111.6 118.31 109.895 ;
      RECT  118.47 111.015 118.385 110.605 ;
      RECT  119.39 112.515 119.21 111.6 ;
      POLYGON  118.385 112.515 118.385 112.185 118.82 112.185 118.82 111.805 118.385 111.805 118.385 111.6 118.31 111.6 118.31 112.515 118.385 112.515 ;
      RECT  118.31 111.6 118.1 109.895 ;
      POLYGON  118.82 111.51 118.82 111.1 118.645 111.1 118.565 111.18 118.565 111.51 118.82 111.51 ;
      RECT  121.43 111.6 121.22 109.895 ;
      RECT  119.75 112.515 119.57 111.6 ;
      RECT  120.83 111.6 120.65 109.895 ;
      RECT  119.03 110.52 118.82 110.11 ;
      RECT  118.31 111.805 118.1 111.6 ;
      RECT  121.22 111.6 121.01 109.895 ;
      RECT  119.03 112.185 118.82 111.805 ;
      RECT  120.47 111.6 120.29 109.895 ;
      RECT  119.75 111.6 119.57 109.895 ;
      RECT  120.47 112.515 120.29 111.6 ;
      RECT  118.31 112.515 118.1 112.185 ;
      RECT  120.11 111.6 119.93 109.895 ;
      RECT  120.11 112.515 119.93 111.6 ;
      RECT  121.43 111.805 121.22 111.6 ;
      RECT  118.31 112.185 118.1 111.805 ;
      RECT  119.39 111.6 119.21 109.895 ;
      RECT  121.22 111.805 121.01 111.6 ;
      RECT  121.43 112.185 121.22 111.805 ;
      POLYGON  118.82 110.52 118.82 110.11 118.565 110.11 118.565 110.44 118.645 110.52 118.82 110.52 ;
      RECT  120.83 112.515 120.65 111.6 ;
      RECT  121.22 112.515 121.01 112.185 ;
      RECT  121.22 112.185 121.01 111.805 ;
      RECT  119.03 112.48 118.82 112.89 ;
      RECT  121.43 111.475 121.22 111.805 ;
      RECT  118.385 112.39 118.31 114.095 ;
      RECT  118.47 112.975 118.385 113.385 ;
      RECT  119.39 111.475 119.21 112.39 ;
      POLYGON  118.385 111.475 118.385 111.805 118.82 111.805 118.82 112.185 118.385 112.185 118.385 112.39 118.31 112.39 118.31 111.475 118.385 111.475 ;
      RECT  118.31 112.39 118.1 114.095 ;
      POLYGON  118.82 112.48 118.82 112.89 118.645 112.89 118.565 112.81 118.565 112.48 118.82 112.48 ;
      RECT  121.43 112.39 121.22 114.095 ;
      RECT  119.75 111.475 119.57 112.39 ;
      RECT  120.83 112.39 120.65 114.095 ;
      RECT  119.03 113.47 118.82 113.88 ;
      RECT  118.31 112.185 118.1 112.39 ;
      RECT  121.22 112.39 121.01 114.095 ;
      RECT  119.03 111.805 118.82 112.185 ;
      RECT  120.47 112.39 120.29 114.095 ;
      RECT  119.75 112.39 119.57 114.095 ;
      RECT  120.47 111.475 120.29 112.39 ;
      RECT  118.31 111.475 118.1 111.805 ;
      RECT  120.11 112.39 119.93 114.095 ;
      RECT  120.11 111.475 119.93 112.39 ;
      RECT  121.43 112.185 121.22 112.39 ;
      RECT  118.31 111.805 118.1 112.185 ;
      RECT  119.39 112.39 119.21 114.095 ;
      RECT  121.22 112.185 121.01 112.39 ;
      RECT  121.43 111.805 121.22 112.185 ;
      POLYGON  118.82 113.47 118.82 113.88 118.565 113.88 118.565 113.55 118.645 113.47 118.82 113.47 ;
      RECT  120.83 111.475 120.65 112.39 ;
      RECT  121.22 111.475 121.01 111.805 ;
      RECT  121.22 111.805 121.01 112.185 ;
      RECT  119.03 115.46 118.82 115.05 ;
      RECT  121.43 116.465 121.22 116.135 ;
      RECT  118.385 115.55 118.31 113.845 ;
      RECT  118.47 114.965 118.385 114.555 ;
      RECT  119.39 116.465 119.21 115.55 ;
      POLYGON  118.385 116.465 118.385 116.135 118.82 116.135 118.82 115.755 118.385 115.755 118.385 115.55 118.31 115.55 118.31 116.465 118.385 116.465 ;
      RECT  118.31 115.55 118.1 113.845 ;
      POLYGON  118.82 115.46 118.82 115.05 118.645 115.05 118.565 115.13 118.565 115.46 118.82 115.46 ;
      RECT  121.43 115.55 121.22 113.845 ;
      RECT  119.75 116.465 119.57 115.55 ;
      RECT  120.83 115.55 120.65 113.845 ;
      RECT  119.03 114.47 118.82 114.06 ;
      RECT  118.31 115.755 118.1 115.55 ;
      RECT  121.22 115.55 121.01 113.845 ;
      RECT  119.03 116.135 118.82 115.755 ;
      RECT  120.47 115.55 120.29 113.845 ;
      RECT  119.75 115.55 119.57 113.845 ;
      RECT  120.47 116.465 120.29 115.55 ;
      RECT  118.31 116.465 118.1 116.135 ;
      RECT  120.11 115.55 119.93 113.845 ;
      RECT  120.11 116.465 119.93 115.55 ;
      RECT  121.43 115.755 121.22 115.55 ;
      RECT  118.31 116.135 118.1 115.755 ;
      RECT  119.39 115.55 119.21 113.845 ;
      RECT  121.22 115.755 121.01 115.55 ;
      RECT  121.43 116.135 121.22 115.755 ;
      POLYGON  118.82 114.47 118.82 114.06 118.565 114.06 118.565 114.39 118.645 114.47 118.82 114.47 ;
      RECT  120.83 116.465 120.65 115.55 ;
      RECT  121.22 116.465 121.01 116.135 ;
      RECT  121.22 116.135 121.01 115.755 ;
      RECT  119.03 116.43 118.82 116.84 ;
      RECT  121.43 115.425 121.22 115.755 ;
      RECT  118.385 116.34 118.31 118.045 ;
      RECT  118.47 116.925 118.385 117.335 ;
      RECT  119.39 115.425 119.21 116.34 ;
      POLYGON  118.385 115.425 118.385 115.755 118.82 115.755 118.82 116.135 118.385 116.135 118.385 116.34 118.31 116.34 118.31 115.425 118.385 115.425 ;
      RECT  118.31 116.34 118.1 118.045 ;
      POLYGON  118.82 116.43 118.82 116.84 118.645 116.84 118.565 116.76 118.565 116.43 118.82 116.43 ;
      RECT  121.43 116.34 121.22 118.045 ;
      RECT  119.75 115.425 119.57 116.34 ;
      RECT  120.83 116.34 120.65 118.045 ;
      RECT  119.03 117.42 118.82 117.83 ;
      RECT  118.31 116.135 118.1 116.34 ;
      RECT  121.22 116.34 121.01 118.045 ;
      RECT  119.03 115.755 118.82 116.135 ;
      RECT  120.47 116.34 120.29 118.045 ;
      RECT  119.75 116.34 119.57 118.045 ;
      RECT  120.47 115.425 120.29 116.34 ;
      RECT  118.31 115.425 118.1 115.755 ;
      RECT  120.11 116.34 119.93 118.045 ;
      RECT  120.11 115.425 119.93 116.34 ;
      RECT  121.43 116.135 121.22 116.34 ;
      RECT  118.31 115.755 118.1 116.135 ;
      RECT  119.39 116.34 119.21 118.045 ;
      RECT  121.22 116.135 121.01 116.34 ;
      RECT  121.43 115.755 121.22 116.135 ;
      POLYGON  118.82 117.42 118.82 117.83 118.565 117.83 118.565 117.5 118.645 117.42 118.82 117.42 ;
      RECT  120.83 115.425 120.65 116.34 ;
      RECT  121.22 115.425 121.01 115.755 ;
      RECT  121.22 115.755 121.01 116.135 ;
      RECT  119.03 119.41 118.82 119.0 ;
      RECT  121.43 120.415 121.22 120.085 ;
      RECT  118.385 119.5 118.31 117.795 ;
      RECT  118.47 118.915 118.385 118.505 ;
      RECT  119.39 120.415 119.21 119.5 ;
      POLYGON  118.385 120.415 118.385 120.085 118.82 120.085 118.82 119.705 118.385 119.705 118.385 119.5 118.31 119.5 118.31 120.415 118.385 120.415 ;
      RECT  118.31 119.5 118.1 117.795 ;
      POLYGON  118.82 119.41 118.82 119.0 118.645 119.0 118.565 119.08 118.565 119.41 118.82 119.41 ;
      RECT  121.43 119.5 121.22 117.795 ;
      RECT  119.75 120.415 119.57 119.5 ;
      RECT  120.83 119.5 120.65 117.795 ;
      RECT  119.03 118.42 118.82 118.01 ;
      RECT  118.31 119.705 118.1 119.5 ;
      RECT  121.22 119.5 121.01 117.795 ;
      RECT  119.03 120.085 118.82 119.705 ;
      RECT  120.47 119.5 120.29 117.795 ;
      RECT  119.75 119.5 119.57 117.795 ;
      RECT  120.47 120.415 120.29 119.5 ;
      RECT  118.31 120.415 118.1 120.085 ;
      RECT  120.11 119.5 119.93 117.795 ;
      RECT  120.11 120.415 119.93 119.5 ;
      RECT  121.43 119.705 121.22 119.5 ;
      RECT  118.31 120.085 118.1 119.705 ;
      RECT  119.39 119.5 119.21 117.795 ;
      RECT  121.22 119.705 121.01 119.5 ;
      RECT  121.43 120.085 121.22 119.705 ;
      POLYGON  118.82 118.42 118.82 118.01 118.565 118.01 118.565 118.34 118.645 118.42 118.82 118.42 ;
      RECT  120.83 120.415 120.65 119.5 ;
      RECT  121.22 120.415 121.01 120.085 ;
      RECT  121.22 120.085 121.01 119.705 ;
      RECT  119.03 120.38 118.82 120.79 ;
      RECT  121.43 119.375 121.22 119.705 ;
      RECT  118.385 120.29 118.31 121.995 ;
      RECT  118.47 120.875 118.385 121.285 ;
      RECT  119.39 119.375 119.21 120.29 ;
      POLYGON  118.385 119.375 118.385 119.705 118.82 119.705 118.82 120.085 118.385 120.085 118.385 120.29 118.31 120.29 118.31 119.375 118.385 119.375 ;
      RECT  118.31 120.29 118.1 121.995 ;
      POLYGON  118.82 120.38 118.82 120.79 118.645 120.79 118.565 120.71 118.565 120.38 118.82 120.38 ;
      RECT  121.43 120.29 121.22 121.995 ;
      RECT  119.75 119.375 119.57 120.29 ;
      RECT  120.83 120.29 120.65 121.995 ;
      RECT  119.03 121.37 118.82 121.78 ;
      RECT  118.31 120.085 118.1 120.29 ;
      RECT  121.22 120.29 121.01 121.995 ;
      RECT  119.03 119.705 118.82 120.085 ;
      RECT  120.47 120.29 120.29 121.995 ;
      RECT  119.75 120.29 119.57 121.995 ;
      RECT  120.47 119.375 120.29 120.29 ;
      RECT  118.31 119.375 118.1 119.705 ;
      RECT  120.11 120.29 119.93 121.995 ;
      RECT  120.11 119.375 119.93 120.29 ;
      RECT  121.43 120.085 121.22 120.29 ;
      RECT  118.31 119.705 118.1 120.085 ;
      RECT  119.39 120.29 119.21 121.995 ;
      RECT  121.22 120.085 121.01 120.29 ;
      RECT  121.43 119.705 121.22 120.085 ;
      POLYGON  118.82 121.37 118.82 121.78 118.565 121.78 118.565 121.45 118.645 121.37 118.82 121.37 ;
      RECT  120.83 119.375 120.65 120.29 ;
      RECT  121.22 119.375 121.01 119.705 ;
      RECT  121.22 119.705 121.01 120.085 ;
      RECT  119.03 123.36 118.82 122.95 ;
      RECT  121.43 124.365 121.22 124.035 ;
      RECT  118.385 123.45 118.31 121.745 ;
      RECT  118.47 122.865 118.385 122.455 ;
      RECT  119.39 124.365 119.21 123.45 ;
      POLYGON  118.385 124.365 118.385 124.035 118.82 124.035 118.82 123.655 118.385 123.655 118.385 123.45 118.31 123.45 118.31 124.365 118.385 124.365 ;
      RECT  118.31 123.45 118.1 121.745 ;
      POLYGON  118.82 123.36 118.82 122.95 118.645 122.95 118.565 123.03 118.565 123.36 118.82 123.36 ;
      RECT  121.43 123.45 121.22 121.745 ;
      RECT  119.75 124.365 119.57 123.45 ;
      RECT  120.83 123.45 120.65 121.745 ;
      RECT  119.03 122.37 118.82 121.96 ;
      RECT  118.31 123.655 118.1 123.45 ;
      RECT  121.22 123.45 121.01 121.745 ;
      RECT  119.03 124.035 118.82 123.655 ;
      RECT  120.47 123.45 120.29 121.745 ;
      RECT  119.75 123.45 119.57 121.745 ;
      RECT  120.47 124.365 120.29 123.45 ;
      RECT  118.31 124.365 118.1 124.035 ;
      RECT  120.11 123.45 119.93 121.745 ;
      RECT  120.11 124.365 119.93 123.45 ;
      RECT  121.43 123.655 121.22 123.45 ;
      RECT  118.31 124.035 118.1 123.655 ;
      RECT  119.39 123.45 119.21 121.745 ;
      RECT  121.22 123.655 121.01 123.45 ;
      RECT  121.43 124.035 121.22 123.655 ;
      POLYGON  118.82 122.37 118.82 121.96 118.565 121.96 118.565 122.29 118.645 122.37 118.82 122.37 ;
      RECT  120.83 124.365 120.65 123.45 ;
      RECT  121.22 124.365 121.01 124.035 ;
      RECT  121.22 124.035 121.01 123.655 ;
      RECT  123.41 92.73 123.62 93.14 ;
      RECT  121.01 91.725 121.22 92.055 ;
      RECT  124.055 92.64 124.13 94.345 ;
      RECT  123.97 93.225 124.055 93.635 ;
      RECT  123.05 91.725 123.23 92.64 ;
      POLYGON  124.055 91.725 124.055 92.055 123.62 92.055 123.62 92.435 124.055 92.435 124.055 92.64 124.13 92.64 124.13 91.725 124.055 91.725 ;
      RECT  124.13 92.64 124.34 94.345 ;
      POLYGON  123.62 92.73 123.62 93.14 123.795 93.14 123.875 93.06 123.875 92.73 123.62 92.73 ;
      RECT  121.01 92.64 121.22 94.345 ;
      RECT  122.69 91.725 122.87 92.64 ;
      RECT  121.61 92.64 121.79 94.345 ;
      RECT  123.41 93.72 123.62 94.13 ;
      RECT  124.13 92.435 124.34 92.64 ;
      RECT  121.22 92.64 121.43 94.345 ;
      RECT  123.41 92.055 123.62 92.435 ;
      RECT  121.97 92.64 122.15 94.345 ;
      RECT  122.69 92.64 122.87 94.345 ;
      RECT  121.97 91.725 122.15 92.64 ;
      RECT  124.13 91.725 124.34 92.055 ;
      RECT  122.33 92.64 122.51 94.345 ;
      RECT  122.33 91.725 122.51 92.64 ;
      RECT  121.01 92.435 121.22 92.64 ;
      RECT  124.13 92.055 124.34 92.435 ;
      RECT  123.05 92.64 123.23 94.345 ;
      RECT  121.22 92.435 121.43 92.64 ;
      RECT  121.01 92.055 121.22 92.435 ;
      POLYGON  123.62 93.72 123.62 94.13 123.875 94.13 123.875 93.8 123.795 93.72 123.62 93.72 ;
      RECT  121.61 91.725 121.79 92.64 ;
      RECT  121.22 91.725 121.43 92.055 ;
      RECT  121.22 92.055 121.43 92.435 ;
      RECT  123.41 95.71 123.62 95.3 ;
      RECT  121.01 96.715 121.22 96.385 ;
      RECT  124.055 95.8 124.13 94.095 ;
      RECT  123.97 95.215 124.055 94.805 ;
      RECT  123.05 96.715 123.23 95.8 ;
      POLYGON  124.055 96.715 124.055 96.385 123.62 96.385 123.62 96.005 124.055 96.005 124.055 95.8 124.13 95.8 124.13 96.715 124.055 96.715 ;
      RECT  124.13 95.8 124.34 94.095 ;
      POLYGON  123.62 95.71 123.62 95.3 123.795 95.3 123.875 95.38 123.875 95.71 123.62 95.71 ;
      RECT  121.01 95.8 121.22 94.095 ;
      RECT  122.69 96.715 122.87 95.8 ;
      RECT  121.61 95.8 121.79 94.095 ;
      RECT  123.41 94.72 123.62 94.31 ;
      RECT  124.13 96.005 124.34 95.8 ;
      RECT  121.22 95.8 121.43 94.095 ;
      RECT  123.41 96.385 123.62 96.005 ;
      RECT  121.97 95.8 122.15 94.095 ;
      RECT  122.69 95.8 122.87 94.095 ;
      RECT  121.97 96.715 122.15 95.8 ;
      RECT  124.13 96.715 124.34 96.385 ;
      RECT  122.33 95.8 122.51 94.095 ;
      RECT  122.33 96.715 122.51 95.8 ;
      RECT  121.01 96.005 121.22 95.8 ;
      RECT  124.13 96.385 124.34 96.005 ;
      RECT  123.05 95.8 123.23 94.095 ;
      RECT  121.22 96.005 121.43 95.8 ;
      RECT  121.01 96.385 121.22 96.005 ;
      POLYGON  123.62 94.72 123.62 94.31 123.875 94.31 123.875 94.64 123.795 94.72 123.62 94.72 ;
      RECT  121.61 96.715 121.79 95.8 ;
      RECT  121.22 96.715 121.43 96.385 ;
      RECT  121.22 96.385 121.43 96.005 ;
      RECT  123.41 96.68 123.62 97.09 ;
      RECT  121.01 95.675 121.22 96.005 ;
      RECT  124.055 96.59 124.13 98.295 ;
      RECT  123.97 97.175 124.055 97.585 ;
      RECT  123.05 95.675 123.23 96.59 ;
      POLYGON  124.055 95.675 124.055 96.005 123.62 96.005 123.62 96.385 124.055 96.385 124.055 96.59 124.13 96.59 124.13 95.675 124.055 95.675 ;
      RECT  124.13 96.59 124.34 98.295 ;
      POLYGON  123.62 96.68 123.62 97.09 123.795 97.09 123.875 97.01 123.875 96.68 123.62 96.68 ;
      RECT  121.01 96.59 121.22 98.295 ;
      RECT  122.69 95.675 122.87 96.59 ;
      RECT  121.61 96.59 121.79 98.295 ;
      RECT  123.41 97.67 123.62 98.08 ;
      RECT  124.13 96.385 124.34 96.59 ;
      RECT  121.22 96.59 121.43 98.295 ;
      RECT  123.41 96.005 123.62 96.385 ;
      RECT  121.97 96.59 122.15 98.295 ;
      RECT  122.69 96.59 122.87 98.295 ;
      RECT  121.97 95.675 122.15 96.59 ;
      RECT  124.13 95.675 124.34 96.005 ;
      RECT  122.33 96.59 122.51 98.295 ;
      RECT  122.33 95.675 122.51 96.59 ;
      RECT  121.01 96.385 121.22 96.59 ;
      RECT  124.13 96.005 124.34 96.385 ;
      RECT  123.05 96.59 123.23 98.295 ;
      RECT  121.22 96.385 121.43 96.59 ;
      RECT  121.01 96.005 121.22 96.385 ;
      POLYGON  123.62 97.67 123.62 98.08 123.875 98.08 123.875 97.75 123.795 97.67 123.62 97.67 ;
      RECT  121.61 95.675 121.79 96.59 ;
      RECT  121.22 95.675 121.43 96.005 ;
      RECT  121.22 96.005 121.43 96.385 ;
      RECT  123.41 99.66 123.62 99.25 ;
      RECT  121.01 100.665 121.22 100.335 ;
      RECT  124.055 99.75 124.13 98.045 ;
      RECT  123.97 99.165 124.055 98.755 ;
      RECT  123.05 100.665 123.23 99.75 ;
      POLYGON  124.055 100.665 124.055 100.335 123.62 100.335 123.62 99.955 124.055 99.955 124.055 99.75 124.13 99.75 124.13 100.665 124.055 100.665 ;
      RECT  124.13 99.75 124.34 98.045 ;
      POLYGON  123.62 99.66 123.62 99.25 123.795 99.25 123.875 99.33 123.875 99.66 123.62 99.66 ;
      RECT  121.01 99.75 121.22 98.045 ;
      RECT  122.69 100.665 122.87 99.75 ;
      RECT  121.61 99.75 121.79 98.045 ;
      RECT  123.41 98.67 123.62 98.26 ;
      RECT  124.13 99.955 124.34 99.75 ;
      RECT  121.22 99.75 121.43 98.045 ;
      RECT  123.41 100.335 123.62 99.955 ;
      RECT  121.97 99.75 122.15 98.045 ;
      RECT  122.69 99.75 122.87 98.045 ;
      RECT  121.97 100.665 122.15 99.75 ;
      RECT  124.13 100.665 124.34 100.335 ;
      RECT  122.33 99.75 122.51 98.045 ;
      RECT  122.33 100.665 122.51 99.75 ;
      RECT  121.01 99.955 121.22 99.75 ;
      RECT  124.13 100.335 124.34 99.955 ;
      RECT  123.05 99.75 123.23 98.045 ;
      RECT  121.22 99.955 121.43 99.75 ;
      RECT  121.01 100.335 121.22 99.955 ;
      POLYGON  123.62 98.67 123.62 98.26 123.875 98.26 123.875 98.59 123.795 98.67 123.62 98.67 ;
      RECT  121.61 100.665 121.79 99.75 ;
      RECT  121.22 100.665 121.43 100.335 ;
      RECT  121.22 100.335 121.43 99.955 ;
      RECT  123.41 100.63 123.62 101.04 ;
      RECT  121.01 99.625 121.22 99.955 ;
      RECT  124.055 100.54 124.13 102.245 ;
      RECT  123.97 101.125 124.055 101.535 ;
      RECT  123.05 99.625 123.23 100.54 ;
      POLYGON  124.055 99.625 124.055 99.955 123.62 99.955 123.62 100.335 124.055 100.335 124.055 100.54 124.13 100.54 124.13 99.625 124.055 99.625 ;
      RECT  124.13 100.54 124.34 102.245 ;
      POLYGON  123.62 100.63 123.62 101.04 123.795 101.04 123.875 100.96 123.875 100.63 123.62 100.63 ;
      RECT  121.01 100.54 121.22 102.245 ;
      RECT  122.69 99.625 122.87 100.54 ;
      RECT  121.61 100.54 121.79 102.245 ;
      RECT  123.41 101.62 123.62 102.03 ;
      RECT  124.13 100.335 124.34 100.54 ;
      RECT  121.22 100.54 121.43 102.245 ;
      RECT  123.41 99.955 123.62 100.335 ;
      RECT  121.97 100.54 122.15 102.245 ;
      RECT  122.69 100.54 122.87 102.245 ;
      RECT  121.97 99.625 122.15 100.54 ;
      RECT  124.13 99.625 124.34 99.955 ;
      RECT  122.33 100.54 122.51 102.245 ;
      RECT  122.33 99.625 122.51 100.54 ;
      RECT  121.01 100.335 121.22 100.54 ;
      RECT  124.13 99.955 124.34 100.335 ;
      RECT  123.05 100.54 123.23 102.245 ;
      RECT  121.22 100.335 121.43 100.54 ;
      RECT  121.01 99.955 121.22 100.335 ;
      POLYGON  123.62 101.62 123.62 102.03 123.875 102.03 123.875 101.7 123.795 101.62 123.62 101.62 ;
      RECT  121.61 99.625 121.79 100.54 ;
      RECT  121.22 99.625 121.43 99.955 ;
      RECT  121.22 99.955 121.43 100.335 ;
      RECT  123.41 103.61 123.62 103.2 ;
      RECT  121.01 104.615 121.22 104.285 ;
      RECT  124.055 103.7 124.13 101.995 ;
      RECT  123.97 103.115 124.055 102.705 ;
      RECT  123.05 104.615 123.23 103.7 ;
      POLYGON  124.055 104.615 124.055 104.285 123.62 104.285 123.62 103.905 124.055 103.905 124.055 103.7 124.13 103.7 124.13 104.615 124.055 104.615 ;
      RECT  124.13 103.7 124.34 101.995 ;
      POLYGON  123.62 103.61 123.62 103.2 123.795 103.2 123.875 103.28 123.875 103.61 123.62 103.61 ;
      RECT  121.01 103.7 121.22 101.995 ;
      RECT  122.69 104.615 122.87 103.7 ;
      RECT  121.61 103.7 121.79 101.995 ;
      RECT  123.41 102.62 123.62 102.21 ;
      RECT  124.13 103.905 124.34 103.7 ;
      RECT  121.22 103.7 121.43 101.995 ;
      RECT  123.41 104.285 123.62 103.905 ;
      RECT  121.97 103.7 122.15 101.995 ;
      RECT  122.69 103.7 122.87 101.995 ;
      RECT  121.97 104.615 122.15 103.7 ;
      RECT  124.13 104.615 124.34 104.285 ;
      RECT  122.33 103.7 122.51 101.995 ;
      RECT  122.33 104.615 122.51 103.7 ;
      RECT  121.01 103.905 121.22 103.7 ;
      RECT  124.13 104.285 124.34 103.905 ;
      RECT  123.05 103.7 123.23 101.995 ;
      RECT  121.22 103.905 121.43 103.7 ;
      RECT  121.01 104.285 121.22 103.905 ;
      POLYGON  123.62 102.62 123.62 102.21 123.875 102.21 123.875 102.54 123.795 102.62 123.62 102.62 ;
      RECT  121.61 104.615 121.79 103.7 ;
      RECT  121.22 104.615 121.43 104.285 ;
      RECT  121.22 104.285 121.43 103.905 ;
      RECT  123.41 104.58 123.62 104.99 ;
      RECT  121.01 103.575 121.22 103.905 ;
      RECT  124.055 104.49 124.13 106.195 ;
      RECT  123.97 105.075 124.055 105.485 ;
      RECT  123.05 103.575 123.23 104.49 ;
      POLYGON  124.055 103.575 124.055 103.905 123.62 103.905 123.62 104.285 124.055 104.285 124.055 104.49 124.13 104.49 124.13 103.575 124.055 103.575 ;
      RECT  124.13 104.49 124.34 106.195 ;
      POLYGON  123.62 104.58 123.62 104.99 123.795 104.99 123.875 104.91 123.875 104.58 123.62 104.58 ;
      RECT  121.01 104.49 121.22 106.195 ;
      RECT  122.69 103.575 122.87 104.49 ;
      RECT  121.61 104.49 121.79 106.195 ;
      RECT  123.41 105.57 123.62 105.98 ;
      RECT  124.13 104.285 124.34 104.49 ;
      RECT  121.22 104.49 121.43 106.195 ;
      RECT  123.41 103.905 123.62 104.285 ;
      RECT  121.97 104.49 122.15 106.195 ;
      RECT  122.69 104.49 122.87 106.195 ;
      RECT  121.97 103.575 122.15 104.49 ;
      RECT  124.13 103.575 124.34 103.905 ;
      RECT  122.33 104.49 122.51 106.195 ;
      RECT  122.33 103.575 122.51 104.49 ;
      RECT  121.01 104.285 121.22 104.49 ;
      RECT  124.13 103.905 124.34 104.285 ;
      RECT  123.05 104.49 123.23 106.195 ;
      RECT  121.22 104.285 121.43 104.49 ;
      RECT  121.01 103.905 121.22 104.285 ;
      POLYGON  123.62 105.57 123.62 105.98 123.875 105.98 123.875 105.65 123.795 105.57 123.62 105.57 ;
      RECT  121.61 103.575 121.79 104.49 ;
      RECT  121.22 103.575 121.43 103.905 ;
      RECT  121.22 103.905 121.43 104.285 ;
      RECT  123.41 107.56 123.62 107.15 ;
      RECT  121.01 108.565 121.22 108.235 ;
      RECT  124.055 107.65 124.13 105.945 ;
      RECT  123.97 107.065 124.055 106.655 ;
      RECT  123.05 108.565 123.23 107.65 ;
      POLYGON  124.055 108.565 124.055 108.235 123.62 108.235 123.62 107.855 124.055 107.855 124.055 107.65 124.13 107.65 124.13 108.565 124.055 108.565 ;
      RECT  124.13 107.65 124.34 105.945 ;
      POLYGON  123.62 107.56 123.62 107.15 123.795 107.15 123.875 107.23 123.875 107.56 123.62 107.56 ;
      RECT  121.01 107.65 121.22 105.945 ;
      RECT  122.69 108.565 122.87 107.65 ;
      RECT  121.61 107.65 121.79 105.945 ;
      RECT  123.41 106.57 123.62 106.16 ;
      RECT  124.13 107.855 124.34 107.65 ;
      RECT  121.22 107.65 121.43 105.945 ;
      RECT  123.41 108.235 123.62 107.855 ;
      RECT  121.97 107.65 122.15 105.945 ;
      RECT  122.69 107.65 122.87 105.945 ;
      RECT  121.97 108.565 122.15 107.65 ;
      RECT  124.13 108.565 124.34 108.235 ;
      RECT  122.33 107.65 122.51 105.945 ;
      RECT  122.33 108.565 122.51 107.65 ;
      RECT  121.01 107.855 121.22 107.65 ;
      RECT  124.13 108.235 124.34 107.855 ;
      RECT  123.05 107.65 123.23 105.945 ;
      RECT  121.22 107.855 121.43 107.65 ;
      RECT  121.01 108.235 121.22 107.855 ;
      POLYGON  123.62 106.57 123.62 106.16 123.875 106.16 123.875 106.49 123.795 106.57 123.62 106.57 ;
      RECT  121.61 108.565 121.79 107.65 ;
      RECT  121.22 108.565 121.43 108.235 ;
      RECT  121.22 108.235 121.43 107.855 ;
      RECT  123.41 108.53 123.62 108.94 ;
      RECT  121.01 107.525 121.22 107.855 ;
      RECT  124.055 108.44 124.13 110.145 ;
      RECT  123.97 109.025 124.055 109.435 ;
      RECT  123.05 107.525 123.23 108.44 ;
      POLYGON  124.055 107.525 124.055 107.855 123.62 107.855 123.62 108.235 124.055 108.235 124.055 108.44 124.13 108.44 124.13 107.525 124.055 107.525 ;
      RECT  124.13 108.44 124.34 110.145 ;
      POLYGON  123.62 108.53 123.62 108.94 123.795 108.94 123.875 108.86 123.875 108.53 123.62 108.53 ;
      RECT  121.01 108.44 121.22 110.145 ;
      RECT  122.69 107.525 122.87 108.44 ;
      RECT  121.61 108.44 121.79 110.145 ;
      RECT  123.41 109.52 123.62 109.93 ;
      RECT  124.13 108.235 124.34 108.44 ;
      RECT  121.22 108.44 121.43 110.145 ;
      RECT  123.41 107.855 123.62 108.235 ;
      RECT  121.97 108.44 122.15 110.145 ;
      RECT  122.69 108.44 122.87 110.145 ;
      RECT  121.97 107.525 122.15 108.44 ;
      RECT  124.13 107.525 124.34 107.855 ;
      RECT  122.33 108.44 122.51 110.145 ;
      RECT  122.33 107.525 122.51 108.44 ;
      RECT  121.01 108.235 121.22 108.44 ;
      RECT  124.13 107.855 124.34 108.235 ;
      RECT  123.05 108.44 123.23 110.145 ;
      RECT  121.22 108.235 121.43 108.44 ;
      RECT  121.01 107.855 121.22 108.235 ;
      POLYGON  123.62 109.52 123.62 109.93 123.875 109.93 123.875 109.6 123.795 109.52 123.62 109.52 ;
      RECT  121.61 107.525 121.79 108.44 ;
      RECT  121.22 107.525 121.43 107.855 ;
      RECT  121.22 107.855 121.43 108.235 ;
      RECT  123.41 111.51 123.62 111.1 ;
      RECT  121.01 112.515 121.22 112.185 ;
      RECT  124.055 111.6 124.13 109.895 ;
      RECT  123.97 111.015 124.055 110.605 ;
      RECT  123.05 112.515 123.23 111.6 ;
      POLYGON  124.055 112.515 124.055 112.185 123.62 112.185 123.62 111.805 124.055 111.805 124.055 111.6 124.13 111.6 124.13 112.515 124.055 112.515 ;
      RECT  124.13 111.6 124.34 109.895 ;
      POLYGON  123.62 111.51 123.62 111.1 123.795 111.1 123.875 111.18 123.875 111.51 123.62 111.51 ;
      RECT  121.01 111.6 121.22 109.895 ;
      RECT  122.69 112.515 122.87 111.6 ;
      RECT  121.61 111.6 121.79 109.895 ;
      RECT  123.41 110.52 123.62 110.11 ;
      RECT  124.13 111.805 124.34 111.6 ;
      RECT  121.22 111.6 121.43 109.895 ;
      RECT  123.41 112.185 123.62 111.805 ;
      RECT  121.97 111.6 122.15 109.895 ;
      RECT  122.69 111.6 122.87 109.895 ;
      RECT  121.97 112.515 122.15 111.6 ;
      RECT  124.13 112.515 124.34 112.185 ;
      RECT  122.33 111.6 122.51 109.895 ;
      RECT  122.33 112.515 122.51 111.6 ;
      RECT  121.01 111.805 121.22 111.6 ;
      RECT  124.13 112.185 124.34 111.805 ;
      RECT  123.05 111.6 123.23 109.895 ;
      RECT  121.22 111.805 121.43 111.6 ;
      RECT  121.01 112.185 121.22 111.805 ;
      POLYGON  123.62 110.52 123.62 110.11 123.875 110.11 123.875 110.44 123.795 110.52 123.62 110.52 ;
      RECT  121.61 112.515 121.79 111.6 ;
      RECT  121.22 112.515 121.43 112.185 ;
      RECT  121.22 112.185 121.43 111.805 ;
      RECT  123.41 112.48 123.62 112.89 ;
      RECT  121.01 111.475 121.22 111.805 ;
      RECT  124.055 112.39 124.13 114.095 ;
      RECT  123.97 112.975 124.055 113.385 ;
      RECT  123.05 111.475 123.23 112.39 ;
      POLYGON  124.055 111.475 124.055 111.805 123.62 111.805 123.62 112.185 124.055 112.185 124.055 112.39 124.13 112.39 124.13 111.475 124.055 111.475 ;
      RECT  124.13 112.39 124.34 114.095 ;
      POLYGON  123.62 112.48 123.62 112.89 123.795 112.89 123.875 112.81 123.875 112.48 123.62 112.48 ;
      RECT  121.01 112.39 121.22 114.095 ;
      RECT  122.69 111.475 122.87 112.39 ;
      RECT  121.61 112.39 121.79 114.095 ;
      RECT  123.41 113.47 123.62 113.88 ;
      RECT  124.13 112.185 124.34 112.39 ;
      RECT  121.22 112.39 121.43 114.095 ;
      RECT  123.41 111.805 123.62 112.185 ;
      RECT  121.97 112.39 122.15 114.095 ;
      RECT  122.69 112.39 122.87 114.095 ;
      RECT  121.97 111.475 122.15 112.39 ;
      RECT  124.13 111.475 124.34 111.805 ;
      RECT  122.33 112.39 122.51 114.095 ;
      RECT  122.33 111.475 122.51 112.39 ;
      RECT  121.01 112.185 121.22 112.39 ;
      RECT  124.13 111.805 124.34 112.185 ;
      RECT  123.05 112.39 123.23 114.095 ;
      RECT  121.22 112.185 121.43 112.39 ;
      RECT  121.01 111.805 121.22 112.185 ;
      POLYGON  123.62 113.47 123.62 113.88 123.875 113.88 123.875 113.55 123.795 113.47 123.62 113.47 ;
      RECT  121.61 111.475 121.79 112.39 ;
      RECT  121.22 111.475 121.43 111.805 ;
      RECT  121.22 111.805 121.43 112.185 ;
      RECT  123.41 115.46 123.62 115.05 ;
      RECT  121.01 116.465 121.22 116.135 ;
      RECT  124.055 115.55 124.13 113.845 ;
      RECT  123.97 114.965 124.055 114.555 ;
      RECT  123.05 116.465 123.23 115.55 ;
      POLYGON  124.055 116.465 124.055 116.135 123.62 116.135 123.62 115.755 124.055 115.755 124.055 115.55 124.13 115.55 124.13 116.465 124.055 116.465 ;
      RECT  124.13 115.55 124.34 113.845 ;
      POLYGON  123.62 115.46 123.62 115.05 123.795 115.05 123.875 115.13 123.875 115.46 123.62 115.46 ;
      RECT  121.01 115.55 121.22 113.845 ;
      RECT  122.69 116.465 122.87 115.55 ;
      RECT  121.61 115.55 121.79 113.845 ;
      RECT  123.41 114.47 123.62 114.06 ;
      RECT  124.13 115.755 124.34 115.55 ;
      RECT  121.22 115.55 121.43 113.845 ;
      RECT  123.41 116.135 123.62 115.755 ;
      RECT  121.97 115.55 122.15 113.845 ;
      RECT  122.69 115.55 122.87 113.845 ;
      RECT  121.97 116.465 122.15 115.55 ;
      RECT  124.13 116.465 124.34 116.135 ;
      RECT  122.33 115.55 122.51 113.845 ;
      RECT  122.33 116.465 122.51 115.55 ;
      RECT  121.01 115.755 121.22 115.55 ;
      RECT  124.13 116.135 124.34 115.755 ;
      RECT  123.05 115.55 123.23 113.845 ;
      RECT  121.22 115.755 121.43 115.55 ;
      RECT  121.01 116.135 121.22 115.755 ;
      POLYGON  123.62 114.47 123.62 114.06 123.875 114.06 123.875 114.39 123.795 114.47 123.62 114.47 ;
      RECT  121.61 116.465 121.79 115.55 ;
      RECT  121.22 116.465 121.43 116.135 ;
      RECT  121.22 116.135 121.43 115.755 ;
      RECT  123.41 116.43 123.62 116.84 ;
      RECT  121.01 115.425 121.22 115.755 ;
      RECT  124.055 116.34 124.13 118.045 ;
      RECT  123.97 116.925 124.055 117.335 ;
      RECT  123.05 115.425 123.23 116.34 ;
      POLYGON  124.055 115.425 124.055 115.755 123.62 115.755 123.62 116.135 124.055 116.135 124.055 116.34 124.13 116.34 124.13 115.425 124.055 115.425 ;
      RECT  124.13 116.34 124.34 118.045 ;
      POLYGON  123.62 116.43 123.62 116.84 123.795 116.84 123.875 116.76 123.875 116.43 123.62 116.43 ;
      RECT  121.01 116.34 121.22 118.045 ;
      RECT  122.69 115.425 122.87 116.34 ;
      RECT  121.61 116.34 121.79 118.045 ;
      RECT  123.41 117.42 123.62 117.83 ;
      RECT  124.13 116.135 124.34 116.34 ;
      RECT  121.22 116.34 121.43 118.045 ;
      RECT  123.41 115.755 123.62 116.135 ;
      RECT  121.97 116.34 122.15 118.045 ;
      RECT  122.69 116.34 122.87 118.045 ;
      RECT  121.97 115.425 122.15 116.34 ;
      RECT  124.13 115.425 124.34 115.755 ;
      RECT  122.33 116.34 122.51 118.045 ;
      RECT  122.33 115.425 122.51 116.34 ;
      RECT  121.01 116.135 121.22 116.34 ;
      RECT  124.13 115.755 124.34 116.135 ;
      RECT  123.05 116.34 123.23 118.045 ;
      RECT  121.22 116.135 121.43 116.34 ;
      RECT  121.01 115.755 121.22 116.135 ;
      POLYGON  123.62 117.42 123.62 117.83 123.875 117.83 123.875 117.5 123.795 117.42 123.62 117.42 ;
      RECT  121.61 115.425 121.79 116.34 ;
      RECT  121.22 115.425 121.43 115.755 ;
      RECT  121.22 115.755 121.43 116.135 ;
      RECT  123.41 119.41 123.62 119.0 ;
      RECT  121.01 120.415 121.22 120.085 ;
      RECT  124.055 119.5 124.13 117.795 ;
      RECT  123.97 118.915 124.055 118.505 ;
      RECT  123.05 120.415 123.23 119.5 ;
      POLYGON  124.055 120.415 124.055 120.085 123.62 120.085 123.62 119.705 124.055 119.705 124.055 119.5 124.13 119.5 124.13 120.415 124.055 120.415 ;
      RECT  124.13 119.5 124.34 117.795 ;
      POLYGON  123.62 119.41 123.62 119.0 123.795 119.0 123.875 119.08 123.875 119.41 123.62 119.41 ;
      RECT  121.01 119.5 121.22 117.795 ;
      RECT  122.69 120.415 122.87 119.5 ;
      RECT  121.61 119.5 121.79 117.795 ;
      RECT  123.41 118.42 123.62 118.01 ;
      RECT  124.13 119.705 124.34 119.5 ;
      RECT  121.22 119.5 121.43 117.795 ;
      RECT  123.41 120.085 123.62 119.705 ;
      RECT  121.97 119.5 122.15 117.795 ;
      RECT  122.69 119.5 122.87 117.795 ;
      RECT  121.97 120.415 122.15 119.5 ;
      RECT  124.13 120.415 124.34 120.085 ;
      RECT  122.33 119.5 122.51 117.795 ;
      RECT  122.33 120.415 122.51 119.5 ;
      RECT  121.01 119.705 121.22 119.5 ;
      RECT  124.13 120.085 124.34 119.705 ;
      RECT  123.05 119.5 123.23 117.795 ;
      RECT  121.22 119.705 121.43 119.5 ;
      RECT  121.01 120.085 121.22 119.705 ;
      POLYGON  123.62 118.42 123.62 118.01 123.875 118.01 123.875 118.34 123.795 118.42 123.62 118.42 ;
      RECT  121.61 120.415 121.79 119.5 ;
      RECT  121.22 120.415 121.43 120.085 ;
      RECT  121.22 120.085 121.43 119.705 ;
      RECT  123.41 120.38 123.62 120.79 ;
      RECT  121.01 119.375 121.22 119.705 ;
      RECT  124.055 120.29 124.13 121.995 ;
      RECT  123.97 120.875 124.055 121.285 ;
      RECT  123.05 119.375 123.23 120.29 ;
      POLYGON  124.055 119.375 124.055 119.705 123.62 119.705 123.62 120.085 124.055 120.085 124.055 120.29 124.13 120.29 124.13 119.375 124.055 119.375 ;
      RECT  124.13 120.29 124.34 121.995 ;
      POLYGON  123.62 120.38 123.62 120.79 123.795 120.79 123.875 120.71 123.875 120.38 123.62 120.38 ;
      RECT  121.01 120.29 121.22 121.995 ;
      RECT  122.69 119.375 122.87 120.29 ;
      RECT  121.61 120.29 121.79 121.995 ;
      RECT  123.41 121.37 123.62 121.78 ;
      RECT  124.13 120.085 124.34 120.29 ;
      RECT  121.22 120.29 121.43 121.995 ;
      RECT  123.41 119.705 123.62 120.085 ;
      RECT  121.97 120.29 122.15 121.995 ;
      RECT  122.69 120.29 122.87 121.995 ;
      RECT  121.97 119.375 122.15 120.29 ;
      RECT  124.13 119.375 124.34 119.705 ;
      RECT  122.33 120.29 122.51 121.995 ;
      RECT  122.33 119.375 122.51 120.29 ;
      RECT  121.01 120.085 121.22 120.29 ;
      RECT  124.13 119.705 124.34 120.085 ;
      RECT  123.05 120.29 123.23 121.995 ;
      RECT  121.22 120.085 121.43 120.29 ;
      RECT  121.01 119.705 121.22 120.085 ;
      POLYGON  123.62 121.37 123.62 121.78 123.875 121.78 123.875 121.45 123.795 121.37 123.62 121.37 ;
      RECT  121.61 119.375 121.79 120.29 ;
      RECT  121.22 119.375 121.43 119.705 ;
      RECT  121.22 119.705 121.43 120.085 ;
      RECT  123.41 123.36 123.62 122.95 ;
      RECT  121.01 124.365 121.22 124.035 ;
      RECT  124.055 123.45 124.13 121.745 ;
      RECT  123.97 122.865 124.055 122.455 ;
      RECT  123.05 124.365 123.23 123.45 ;
      POLYGON  124.055 124.365 124.055 124.035 123.62 124.035 123.62 123.655 124.055 123.655 124.055 123.45 124.13 123.45 124.13 124.365 124.055 124.365 ;
      RECT  124.13 123.45 124.34 121.745 ;
      POLYGON  123.62 123.36 123.62 122.95 123.795 122.95 123.875 123.03 123.875 123.36 123.62 123.36 ;
      RECT  121.01 123.45 121.22 121.745 ;
      RECT  122.69 124.365 122.87 123.45 ;
      RECT  121.61 123.45 121.79 121.745 ;
      RECT  123.41 122.37 123.62 121.96 ;
      RECT  124.13 123.655 124.34 123.45 ;
      RECT  121.22 123.45 121.43 121.745 ;
      RECT  123.41 124.035 123.62 123.655 ;
      RECT  121.97 123.45 122.15 121.745 ;
      RECT  122.69 123.45 122.87 121.745 ;
      RECT  121.97 124.365 122.15 123.45 ;
      RECT  124.13 124.365 124.34 124.035 ;
      RECT  122.33 123.45 122.51 121.745 ;
      RECT  122.33 124.365 122.51 123.45 ;
      RECT  121.01 123.655 121.22 123.45 ;
      RECT  124.13 124.035 124.34 123.655 ;
      RECT  123.05 123.45 123.23 121.745 ;
      RECT  121.22 123.655 121.43 123.45 ;
      RECT  121.01 124.035 121.22 123.655 ;
      POLYGON  123.62 122.37 123.62 121.96 123.875 121.96 123.875 122.29 123.795 122.37 123.62 122.37 ;
      RECT  121.61 124.365 121.79 123.45 ;
      RECT  121.22 124.365 121.43 124.035 ;
      RECT  121.22 124.035 121.43 123.655 ;
      RECT  125.27 92.73 125.06 93.14 ;
      RECT  127.67 91.725 127.46 92.055 ;
      RECT  124.625 92.64 124.55 94.345 ;
      RECT  124.71 93.225 124.625 93.635 ;
      RECT  125.63 91.725 125.45 92.64 ;
      POLYGON  124.625 91.725 124.625 92.055 125.06 92.055 125.06 92.435 124.625 92.435 124.625 92.64 124.55 92.64 124.55 91.725 124.625 91.725 ;
      RECT  124.55 92.64 124.34 94.345 ;
      POLYGON  125.06 92.73 125.06 93.14 124.885 93.14 124.805 93.06 124.805 92.73 125.06 92.73 ;
      RECT  127.67 92.64 127.46 94.345 ;
      RECT  125.99 91.725 125.81 92.64 ;
      RECT  127.07 92.64 126.89 94.345 ;
      RECT  125.27 93.72 125.06 94.13 ;
      RECT  124.55 92.435 124.34 92.64 ;
      RECT  127.46 92.64 127.25 94.345 ;
      RECT  125.27 92.055 125.06 92.435 ;
      RECT  126.71 92.64 126.53 94.345 ;
      RECT  125.99 92.64 125.81 94.345 ;
      RECT  126.71 91.725 126.53 92.64 ;
      RECT  124.55 91.725 124.34 92.055 ;
      RECT  126.35 92.64 126.17 94.345 ;
      RECT  126.35 91.725 126.17 92.64 ;
      RECT  127.67 92.435 127.46 92.64 ;
      RECT  124.55 92.055 124.34 92.435 ;
      RECT  125.63 92.64 125.45 94.345 ;
      RECT  127.46 92.435 127.25 92.64 ;
      RECT  127.67 92.055 127.46 92.435 ;
      POLYGON  125.06 93.72 125.06 94.13 124.805 94.13 124.805 93.8 124.885 93.72 125.06 93.72 ;
      RECT  127.07 91.725 126.89 92.64 ;
      RECT  127.46 91.725 127.25 92.055 ;
      RECT  127.46 92.055 127.25 92.435 ;
      RECT  125.27 95.71 125.06 95.3 ;
      RECT  127.67 96.715 127.46 96.385 ;
      RECT  124.625 95.8 124.55 94.095 ;
      RECT  124.71 95.215 124.625 94.805 ;
      RECT  125.63 96.715 125.45 95.8 ;
      POLYGON  124.625 96.715 124.625 96.385 125.06 96.385 125.06 96.005 124.625 96.005 124.625 95.8 124.55 95.8 124.55 96.715 124.625 96.715 ;
      RECT  124.55 95.8 124.34 94.095 ;
      POLYGON  125.06 95.71 125.06 95.3 124.885 95.3 124.805 95.38 124.805 95.71 125.06 95.71 ;
      RECT  127.67 95.8 127.46 94.095 ;
      RECT  125.99 96.715 125.81 95.8 ;
      RECT  127.07 95.8 126.89 94.095 ;
      RECT  125.27 94.72 125.06 94.31 ;
      RECT  124.55 96.005 124.34 95.8 ;
      RECT  127.46 95.8 127.25 94.095 ;
      RECT  125.27 96.385 125.06 96.005 ;
      RECT  126.71 95.8 126.53 94.095 ;
      RECT  125.99 95.8 125.81 94.095 ;
      RECT  126.71 96.715 126.53 95.8 ;
      RECT  124.55 96.715 124.34 96.385 ;
      RECT  126.35 95.8 126.17 94.095 ;
      RECT  126.35 96.715 126.17 95.8 ;
      RECT  127.67 96.005 127.46 95.8 ;
      RECT  124.55 96.385 124.34 96.005 ;
      RECT  125.63 95.8 125.45 94.095 ;
      RECT  127.46 96.005 127.25 95.8 ;
      RECT  127.67 96.385 127.46 96.005 ;
      POLYGON  125.06 94.72 125.06 94.31 124.805 94.31 124.805 94.64 124.885 94.72 125.06 94.72 ;
      RECT  127.07 96.715 126.89 95.8 ;
      RECT  127.46 96.715 127.25 96.385 ;
      RECT  127.46 96.385 127.25 96.005 ;
      RECT  125.27 96.68 125.06 97.09 ;
      RECT  127.67 95.675 127.46 96.005 ;
      RECT  124.625 96.59 124.55 98.295 ;
      RECT  124.71 97.175 124.625 97.585 ;
      RECT  125.63 95.675 125.45 96.59 ;
      POLYGON  124.625 95.675 124.625 96.005 125.06 96.005 125.06 96.385 124.625 96.385 124.625 96.59 124.55 96.59 124.55 95.675 124.625 95.675 ;
      RECT  124.55 96.59 124.34 98.295 ;
      POLYGON  125.06 96.68 125.06 97.09 124.885 97.09 124.805 97.01 124.805 96.68 125.06 96.68 ;
      RECT  127.67 96.59 127.46 98.295 ;
      RECT  125.99 95.675 125.81 96.59 ;
      RECT  127.07 96.59 126.89 98.295 ;
      RECT  125.27 97.67 125.06 98.08 ;
      RECT  124.55 96.385 124.34 96.59 ;
      RECT  127.46 96.59 127.25 98.295 ;
      RECT  125.27 96.005 125.06 96.385 ;
      RECT  126.71 96.59 126.53 98.295 ;
      RECT  125.99 96.59 125.81 98.295 ;
      RECT  126.71 95.675 126.53 96.59 ;
      RECT  124.55 95.675 124.34 96.005 ;
      RECT  126.35 96.59 126.17 98.295 ;
      RECT  126.35 95.675 126.17 96.59 ;
      RECT  127.67 96.385 127.46 96.59 ;
      RECT  124.55 96.005 124.34 96.385 ;
      RECT  125.63 96.59 125.45 98.295 ;
      RECT  127.46 96.385 127.25 96.59 ;
      RECT  127.67 96.005 127.46 96.385 ;
      POLYGON  125.06 97.67 125.06 98.08 124.805 98.08 124.805 97.75 124.885 97.67 125.06 97.67 ;
      RECT  127.07 95.675 126.89 96.59 ;
      RECT  127.46 95.675 127.25 96.005 ;
      RECT  127.46 96.005 127.25 96.385 ;
      RECT  125.27 99.66 125.06 99.25 ;
      RECT  127.67 100.665 127.46 100.335 ;
      RECT  124.625 99.75 124.55 98.045 ;
      RECT  124.71 99.165 124.625 98.755 ;
      RECT  125.63 100.665 125.45 99.75 ;
      POLYGON  124.625 100.665 124.625 100.335 125.06 100.335 125.06 99.955 124.625 99.955 124.625 99.75 124.55 99.75 124.55 100.665 124.625 100.665 ;
      RECT  124.55 99.75 124.34 98.045 ;
      POLYGON  125.06 99.66 125.06 99.25 124.885 99.25 124.805 99.33 124.805 99.66 125.06 99.66 ;
      RECT  127.67 99.75 127.46 98.045 ;
      RECT  125.99 100.665 125.81 99.75 ;
      RECT  127.07 99.75 126.89 98.045 ;
      RECT  125.27 98.67 125.06 98.26 ;
      RECT  124.55 99.955 124.34 99.75 ;
      RECT  127.46 99.75 127.25 98.045 ;
      RECT  125.27 100.335 125.06 99.955 ;
      RECT  126.71 99.75 126.53 98.045 ;
      RECT  125.99 99.75 125.81 98.045 ;
      RECT  126.71 100.665 126.53 99.75 ;
      RECT  124.55 100.665 124.34 100.335 ;
      RECT  126.35 99.75 126.17 98.045 ;
      RECT  126.35 100.665 126.17 99.75 ;
      RECT  127.67 99.955 127.46 99.75 ;
      RECT  124.55 100.335 124.34 99.955 ;
      RECT  125.63 99.75 125.45 98.045 ;
      RECT  127.46 99.955 127.25 99.75 ;
      RECT  127.67 100.335 127.46 99.955 ;
      POLYGON  125.06 98.67 125.06 98.26 124.805 98.26 124.805 98.59 124.885 98.67 125.06 98.67 ;
      RECT  127.07 100.665 126.89 99.75 ;
      RECT  127.46 100.665 127.25 100.335 ;
      RECT  127.46 100.335 127.25 99.955 ;
      RECT  125.27 100.63 125.06 101.04 ;
      RECT  127.67 99.625 127.46 99.955 ;
      RECT  124.625 100.54 124.55 102.245 ;
      RECT  124.71 101.125 124.625 101.535 ;
      RECT  125.63 99.625 125.45 100.54 ;
      POLYGON  124.625 99.625 124.625 99.955 125.06 99.955 125.06 100.335 124.625 100.335 124.625 100.54 124.55 100.54 124.55 99.625 124.625 99.625 ;
      RECT  124.55 100.54 124.34 102.245 ;
      POLYGON  125.06 100.63 125.06 101.04 124.885 101.04 124.805 100.96 124.805 100.63 125.06 100.63 ;
      RECT  127.67 100.54 127.46 102.245 ;
      RECT  125.99 99.625 125.81 100.54 ;
      RECT  127.07 100.54 126.89 102.245 ;
      RECT  125.27 101.62 125.06 102.03 ;
      RECT  124.55 100.335 124.34 100.54 ;
      RECT  127.46 100.54 127.25 102.245 ;
      RECT  125.27 99.955 125.06 100.335 ;
      RECT  126.71 100.54 126.53 102.245 ;
      RECT  125.99 100.54 125.81 102.245 ;
      RECT  126.71 99.625 126.53 100.54 ;
      RECT  124.55 99.625 124.34 99.955 ;
      RECT  126.35 100.54 126.17 102.245 ;
      RECT  126.35 99.625 126.17 100.54 ;
      RECT  127.67 100.335 127.46 100.54 ;
      RECT  124.55 99.955 124.34 100.335 ;
      RECT  125.63 100.54 125.45 102.245 ;
      RECT  127.46 100.335 127.25 100.54 ;
      RECT  127.67 99.955 127.46 100.335 ;
      POLYGON  125.06 101.62 125.06 102.03 124.805 102.03 124.805 101.7 124.885 101.62 125.06 101.62 ;
      RECT  127.07 99.625 126.89 100.54 ;
      RECT  127.46 99.625 127.25 99.955 ;
      RECT  127.46 99.955 127.25 100.335 ;
      RECT  125.27 103.61 125.06 103.2 ;
      RECT  127.67 104.615 127.46 104.285 ;
      RECT  124.625 103.7 124.55 101.995 ;
      RECT  124.71 103.115 124.625 102.705 ;
      RECT  125.63 104.615 125.45 103.7 ;
      POLYGON  124.625 104.615 124.625 104.285 125.06 104.285 125.06 103.905 124.625 103.905 124.625 103.7 124.55 103.7 124.55 104.615 124.625 104.615 ;
      RECT  124.55 103.7 124.34 101.995 ;
      POLYGON  125.06 103.61 125.06 103.2 124.885 103.2 124.805 103.28 124.805 103.61 125.06 103.61 ;
      RECT  127.67 103.7 127.46 101.995 ;
      RECT  125.99 104.615 125.81 103.7 ;
      RECT  127.07 103.7 126.89 101.995 ;
      RECT  125.27 102.62 125.06 102.21 ;
      RECT  124.55 103.905 124.34 103.7 ;
      RECT  127.46 103.7 127.25 101.995 ;
      RECT  125.27 104.285 125.06 103.905 ;
      RECT  126.71 103.7 126.53 101.995 ;
      RECT  125.99 103.7 125.81 101.995 ;
      RECT  126.71 104.615 126.53 103.7 ;
      RECT  124.55 104.615 124.34 104.285 ;
      RECT  126.35 103.7 126.17 101.995 ;
      RECT  126.35 104.615 126.17 103.7 ;
      RECT  127.67 103.905 127.46 103.7 ;
      RECT  124.55 104.285 124.34 103.905 ;
      RECT  125.63 103.7 125.45 101.995 ;
      RECT  127.46 103.905 127.25 103.7 ;
      RECT  127.67 104.285 127.46 103.905 ;
      POLYGON  125.06 102.62 125.06 102.21 124.805 102.21 124.805 102.54 124.885 102.62 125.06 102.62 ;
      RECT  127.07 104.615 126.89 103.7 ;
      RECT  127.46 104.615 127.25 104.285 ;
      RECT  127.46 104.285 127.25 103.905 ;
      RECT  125.27 104.58 125.06 104.99 ;
      RECT  127.67 103.575 127.46 103.905 ;
      RECT  124.625 104.49 124.55 106.195 ;
      RECT  124.71 105.075 124.625 105.485 ;
      RECT  125.63 103.575 125.45 104.49 ;
      POLYGON  124.625 103.575 124.625 103.905 125.06 103.905 125.06 104.285 124.625 104.285 124.625 104.49 124.55 104.49 124.55 103.575 124.625 103.575 ;
      RECT  124.55 104.49 124.34 106.195 ;
      POLYGON  125.06 104.58 125.06 104.99 124.885 104.99 124.805 104.91 124.805 104.58 125.06 104.58 ;
      RECT  127.67 104.49 127.46 106.195 ;
      RECT  125.99 103.575 125.81 104.49 ;
      RECT  127.07 104.49 126.89 106.195 ;
      RECT  125.27 105.57 125.06 105.98 ;
      RECT  124.55 104.285 124.34 104.49 ;
      RECT  127.46 104.49 127.25 106.195 ;
      RECT  125.27 103.905 125.06 104.285 ;
      RECT  126.71 104.49 126.53 106.195 ;
      RECT  125.99 104.49 125.81 106.195 ;
      RECT  126.71 103.575 126.53 104.49 ;
      RECT  124.55 103.575 124.34 103.905 ;
      RECT  126.35 104.49 126.17 106.195 ;
      RECT  126.35 103.575 126.17 104.49 ;
      RECT  127.67 104.285 127.46 104.49 ;
      RECT  124.55 103.905 124.34 104.285 ;
      RECT  125.63 104.49 125.45 106.195 ;
      RECT  127.46 104.285 127.25 104.49 ;
      RECT  127.67 103.905 127.46 104.285 ;
      POLYGON  125.06 105.57 125.06 105.98 124.805 105.98 124.805 105.65 124.885 105.57 125.06 105.57 ;
      RECT  127.07 103.575 126.89 104.49 ;
      RECT  127.46 103.575 127.25 103.905 ;
      RECT  127.46 103.905 127.25 104.285 ;
      RECT  125.27 107.56 125.06 107.15 ;
      RECT  127.67 108.565 127.46 108.235 ;
      RECT  124.625 107.65 124.55 105.945 ;
      RECT  124.71 107.065 124.625 106.655 ;
      RECT  125.63 108.565 125.45 107.65 ;
      POLYGON  124.625 108.565 124.625 108.235 125.06 108.235 125.06 107.855 124.625 107.855 124.625 107.65 124.55 107.65 124.55 108.565 124.625 108.565 ;
      RECT  124.55 107.65 124.34 105.945 ;
      POLYGON  125.06 107.56 125.06 107.15 124.885 107.15 124.805 107.23 124.805 107.56 125.06 107.56 ;
      RECT  127.67 107.65 127.46 105.945 ;
      RECT  125.99 108.565 125.81 107.65 ;
      RECT  127.07 107.65 126.89 105.945 ;
      RECT  125.27 106.57 125.06 106.16 ;
      RECT  124.55 107.855 124.34 107.65 ;
      RECT  127.46 107.65 127.25 105.945 ;
      RECT  125.27 108.235 125.06 107.855 ;
      RECT  126.71 107.65 126.53 105.945 ;
      RECT  125.99 107.65 125.81 105.945 ;
      RECT  126.71 108.565 126.53 107.65 ;
      RECT  124.55 108.565 124.34 108.235 ;
      RECT  126.35 107.65 126.17 105.945 ;
      RECT  126.35 108.565 126.17 107.65 ;
      RECT  127.67 107.855 127.46 107.65 ;
      RECT  124.55 108.235 124.34 107.855 ;
      RECT  125.63 107.65 125.45 105.945 ;
      RECT  127.46 107.855 127.25 107.65 ;
      RECT  127.67 108.235 127.46 107.855 ;
      POLYGON  125.06 106.57 125.06 106.16 124.805 106.16 124.805 106.49 124.885 106.57 125.06 106.57 ;
      RECT  127.07 108.565 126.89 107.65 ;
      RECT  127.46 108.565 127.25 108.235 ;
      RECT  127.46 108.235 127.25 107.855 ;
      RECT  125.27 108.53 125.06 108.94 ;
      RECT  127.67 107.525 127.46 107.855 ;
      RECT  124.625 108.44 124.55 110.145 ;
      RECT  124.71 109.025 124.625 109.435 ;
      RECT  125.63 107.525 125.45 108.44 ;
      POLYGON  124.625 107.525 124.625 107.855 125.06 107.855 125.06 108.235 124.625 108.235 124.625 108.44 124.55 108.44 124.55 107.525 124.625 107.525 ;
      RECT  124.55 108.44 124.34 110.145 ;
      POLYGON  125.06 108.53 125.06 108.94 124.885 108.94 124.805 108.86 124.805 108.53 125.06 108.53 ;
      RECT  127.67 108.44 127.46 110.145 ;
      RECT  125.99 107.525 125.81 108.44 ;
      RECT  127.07 108.44 126.89 110.145 ;
      RECT  125.27 109.52 125.06 109.93 ;
      RECT  124.55 108.235 124.34 108.44 ;
      RECT  127.46 108.44 127.25 110.145 ;
      RECT  125.27 107.855 125.06 108.235 ;
      RECT  126.71 108.44 126.53 110.145 ;
      RECT  125.99 108.44 125.81 110.145 ;
      RECT  126.71 107.525 126.53 108.44 ;
      RECT  124.55 107.525 124.34 107.855 ;
      RECT  126.35 108.44 126.17 110.145 ;
      RECT  126.35 107.525 126.17 108.44 ;
      RECT  127.67 108.235 127.46 108.44 ;
      RECT  124.55 107.855 124.34 108.235 ;
      RECT  125.63 108.44 125.45 110.145 ;
      RECT  127.46 108.235 127.25 108.44 ;
      RECT  127.67 107.855 127.46 108.235 ;
      POLYGON  125.06 109.52 125.06 109.93 124.805 109.93 124.805 109.6 124.885 109.52 125.06 109.52 ;
      RECT  127.07 107.525 126.89 108.44 ;
      RECT  127.46 107.525 127.25 107.855 ;
      RECT  127.46 107.855 127.25 108.235 ;
      RECT  125.27 111.51 125.06 111.1 ;
      RECT  127.67 112.515 127.46 112.185 ;
      RECT  124.625 111.6 124.55 109.895 ;
      RECT  124.71 111.015 124.625 110.605 ;
      RECT  125.63 112.515 125.45 111.6 ;
      POLYGON  124.625 112.515 124.625 112.185 125.06 112.185 125.06 111.805 124.625 111.805 124.625 111.6 124.55 111.6 124.55 112.515 124.625 112.515 ;
      RECT  124.55 111.6 124.34 109.895 ;
      POLYGON  125.06 111.51 125.06 111.1 124.885 111.1 124.805 111.18 124.805 111.51 125.06 111.51 ;
      RECT  127.67 111.6 127.46 109.895 ;
      RECT  125.99 112.515 125.81 111.6 ;
      RECT  127.07 111.6 126.89 109.895 ;
      RECT  125.27 110.52 125.06 110.11 ;
      RECT  124.55 111.805 124.34 111.6 ;
      RECT  127.46 111.6 127.25 109.895 ;
      RECT  125.27 112.185 125.06 111.805 ;
      RECT  126.71 111.6 126.53 109.895 ;
      RECT  125.99 111.6 125.81 109.895 ;
      RECT  126.71 112.515 126.53 111.6 ;
      RECT  124.55 112.515 124.34 112.185 ;
      RECT  126.35 111.6 126.17 109.895 ;
      RECT  126.35 112.515 126.17 111.6 ;
      RECT  127.67 111.805 127.46 111.6 ;
      RECT  124.55 112.185 124.34 111.805 ;
      RECT  125.63 111.6 125.45 109.895 ;
      RECT  127.46 111.805 127.25 111.6 ;
      RECT  127.67 112.185 127.46 111.805 ;
      POLYGON  125.06 110.52 125.06 110.11 124.805 110.11 124.805 110.44 124.885 110.52 125.06 110.52 ;
      RECT  127.07 112.515 126.89 111.6 ;
      RECT  127.46 112.515 127.25 112.185 ;
      RECT  127.46 112.185 127.25 111.805 ;
      RECT  125.27 112.48 125.06 112.89 ;
      RECT  127.67 111.475 127.46 111.805 ;
      RECT  124.625 112.39 124.55 114.095 ;
      RECT  124.71 112.975 124.625 113.385 ;
      RECT  125.63 111.475 125.45 112.39 ;
      POLYGON  124.625 111.475 124.625 111.805 125.06 111.805 125.06 112.185 124.625 112.185 124.625 112.39 124.55 112.39 124.55 111.475 124.625 111.475 ;
      RECT  124.55 112.39 124.34 114.095 ;
      POLYGON  125.06 112.48 125.06 112.89 124.885 112.89 124.805 112.81 124.805 112.48 125.06 112.48 ;
      RECT  127.67 112.39 127.46 114.095 ;
      RECT  125.99 111.475 125.81 112.39 ;
      RECT  127.07 112.39 126.89 114.095 ;
      RECT  125.27 113.47 125.06 113.88 ;
      RECT  124.55 112.185 124.34 112.39 ;
      RECT  127.46 112.39 127.25 114.095 ;
      RECT  125.27 111.805 125.06 112.185 ;
      RECT  126.71 112.39 126.53 114.095 ;
      RECT  125.99 112.39 125.81 114.095 ;
      RECT  126.71 111.475 126.53 112.39 ;
      RECT  124.55 111.475 124.34 111.805 ;
      RECT  126.35 112.39 126.17 114.095 ;
      RECT  126.35 111.475 126.17 112.39 ;
      RECT  127.67 112.185 127.46 112.39 ;
      RECT  124.55 111.805 124.34 112.185 ;
      RECT  125.63 112.39 125.45 114.095 ;
      RECT  127.46 112.185 127.25 112.39 ;
      RECT  127.67 111.805 127.46 112.185 ;
      POLYGON  125.06 113.47 125.06 113.88 124.805 113.88 124.805 113.55 124.885 113.47 125.06 113.47 ;
      RECT  127.07 111.475 126.89 112.39 ;
      RECT  127.46 111.475 127.25 111.805 ;
      RECT  127.46 111.805 127.25 112.185 ;
      RECT  125.27 115.46 125.06 115.05 ;
      RECT  127.67 116.465 127.46 116.135 ;
      RECT  124.625 115.55 124.55 113.845 ;
      RECT  124.71 114.965 124.625 114.555 ;
      RECT  125.63 116.465 125.45 115.55 ;
      POLYGON  124.625 116.465 124.625 116.135 125.06 116.135 125.06 115.755 124.625 115.755 124.625 115.55 124.55 115.55 124.55 116.465 124.625 116.465 ;
      RECT  124.55 115.55 124.34 113.845 ;
      POLYGON  125.06 115.46 125.06 115.05 124.885 115.05 124.805 115.13 124.805 115.46 125.06 115.46 ;
      RECT  127.67 115.55 127.46 113.845 ;
      RECT  125.99 116.465 125.81 115.55 ;
      RECT  127.07 115.55 126.89 113.845 ;
      RECT  125.27 114.47 125.06 114.06 ;
      RECT  124.55 115.755 124.34 115.55 ;
      RECT  127.46 115.55 127.25 113.845 ;
      RECT  125.27 116.135 125.06 115.755 ;
      RECT  126.71 115.55 126.53 113.845 ;
      RECT  125.99 115.55 125.81 113.845 ;
      RECT  126.71 116.465 126.53 115.55 ;
      RECT  124.55 116.465 124.34 116.135 ;
      RECT  126.35 115.55 126.17 113.845 ;
      RECT  126.35 116.465 126.17 115.55 ;
      RECT  127.67 115.755 127.46 115.55 ;
      RECT  124.55 116.135 124.34 115.755 ;
      RECT  125.63 115.55 125.45 113.845 ;
      RECT  127.46 115.755 127.25 115.55 ;
      RECT  127.67 116.135 127.46 115.755 ;
      POLYGON  125.06 114.47 125.06 114.06 124.805 114.06 124.805 114.39 124.885 114.47 125.06 114.47 ;
      RECT  127.07 116.465 126.89 115.55 ;
      RECT  127.46 116.465 127.25 116.135 ;
      RECT  127.46 116.135 127.25 115.755 ;
      RECT  125.27 116.43 125.06 116.84 ;
      RECT  127.67 115.425 127.46 115.755 ;
      RECT  124.625 116.34 124.55 118.045 ;
      RECT  124.71 116.925 124.625 117.335 ;
      RECT  125.63 115.425 125.45 116.34 ;
      POLYGON  124.625 115.425 124.625 115.755 125.06 115.755 125.06 116.135 124.625 116.135 124.625 116.34 124.55 116.34 124.55 115.425 124.625 115.425 ;
      RECT  124.55 116.34 124.34 118.045 ;
      POLYGON  125.06 116.43 125.06 116.84 124.885 116.84 124.805 116.76 124.805 116.43 125.06 116.43 ;
      RECT  127.67 116.34 127.46 118.045 ;
      RECT  125.99 115.425 125.81 116.34 ;
      RECT  127.07 116.34 126.89 118.045 ;
      RECT  125.27 117.42 125.06 117.83 ;
      RECT  124.55 116.135 124.34 116.34 ;
      RECT  127.46 116.34 127.25 118.045 ;
      RECT  125.27 115.755 125.06 116.135 ;
      RECT  126.71 116.34 126.53 118.045 ;
      RECT  125.99 116.34 125.81 118.045 ;
      RECT  126.71 115.425 126.53 116.34 ;
      RECT  124.55 115.425 124.34 115.755 ;
      RECT  126.35 116.34 126.17 118.045 ;
      RECT  126.35 115.425 126.17 116.34 ;
      RECT  127.67 116.135 127.46 116.34 ;
      RECT  124.55 115.755 124.34 116.135 ;
      RECT  125.63 116.34 125.45 118.045 ;
      RECT  127.46 116.135 127.25 116.34 ;
      RECT  127.67 115.755 127.46 116.135 ;
      POLYGON  125.06 117.42 125.06 117.83 124.805 117.83 124.805 117.5 124.885 117.42 125.06 117.42 ;
      RECT  127.07 115.425 126.89 116.34 ;
      RECT  127.46 115.425 127.25 115.755 ;
      RECT  127.46 115.755 127.25 116.135 ;
      RECT  125.27 119.41 125.06 119.0 ;
      RECT  127.67 120.415 127.46 120.085 ;
      RECT  124.625 119.5 124.55 117.795 ;
      RECT  124.71 118.915 124.625 118.505 ;
      RECT  125.63 120.415 125.45 119.5 ;
      POLYGON  124.625 120.415 124.625 120.085 125.06 120.085 125.06 119.705 124.625 119.705 124.625 119.5 124.55 119.5 124.55 120.415 124.625 120.415 ;
      RECT  124.55 119.5 124.34 117.795 ;
      POLYGON  125.06 119.41 125.06 119.0 124.885 119.0 124.805 119.08 124.805 119.41 125.06 119.41 ;
      RECT  127.67 119.5 127.46 117.795 ;
      RECT  125.99 120.415 125.81 119.5 ;
      RECT  127.07 119.5 126.89 117.795 ;
      RECT  125.27 118.42 125.06 118.01 ;
      RECT  124.55 119.705 124.34 119.5 ;
      RECT  127.46 119.5 127.25 117.795 ;
      RECT  125.27 120.085 125.06 119.705 ;
      RECT  126.71 119.5 126.53 117.795 ;
      RECT  125.99 119.5 125.81 117.795 ;
      RECT  126.71 120.415 126.53 119.5 ;
      RECT  124.55 120.415 124.34 120.085 ;
      RECT  126.35 119.5 126.17 117.795 ;
      RECT  126.35 120.415 126.17 119.5 ;
      RECT  127.67 119.705 127.46 119.5 ;
      RECT  124.55 120.085 124.34 119.705 ;
      RECT  125.63 119.5 125.45 117.795 ;
      RECT  127.46 119.705 127.25 119.5 ;
      RECT  127.67 120.085 127.46 119.705 ;
      POLYGON  125.06 118.42 125.06 118.01 124.805 118.01 124.805 118.34 124.885 118.42 125.06 118.42 ;
      RECT  127.07 120.415 126.89 119.5 ;
      RECT  127.46 120.415 127.25 120.085 ;
      RECT  127.46 120.085 127.25 119.705 ;
      RECT  125.27 120.38 125.06 120.79 ;
      RECT  127.67 119.375 127.46 119.705 ;
      RECT  124.625 120.29 124.55 121.995 ;
      RECT  124.71 120.875 124.625 121.285 ;
      RECT  125.63 119.375 125.45 120.29 ;
      POLYGON  124.625 119.375 124.625 119.705 125.06 119.705 125.06 120.085 124.625 120.085 124.625 120.29 124.55 120.29 124.55 119.375 124.625 119.375 ;
      RECT  124.55 120.29 124.34 121.995 ;
      POLYGON  125.06 120.38 125.06 120.79 124.885 120.79 124.805 120.71 124.805 120.38 125.06 120.38 ;
      RECT  127.67 120.29 127.46 121.995 ;
      RECT  125.99 119.375 125.81 120.29 ;
      RECT  127.07 120.29 126.89 121.995 ;
      RECT  125.27 121.37 125.06 121.78 ;
      RECT  124.55 120.085 124.34 120.29 ;
      RECT  127.46 120.29 127.25 121.995 ;
      RECT  125.27 119.705 125.06 120.085 ;
      RECT  126.71 120.29 126.53 121.995 ;
      RECT  125.99 120.29 125.81 121.995 ;
      RECT  126.71 119.375 126.53 120.29 ;
      RECT  124.55 119.375 124.34 119.705 ;
      RECT  126.35 120.29 126.17 121.995 ;
      RECT  126.35 119.375 126.17 120.29 ;
      RECT  127.67 120.085 127.46 120.29 ;
      RECT  124.55 119.705 124.34 120.085 ;
      RECT  125.63 120.29 125.45 121.995 ;
      RECT  127.46 120.085 127.25 120.29 ;
      RECT  127.67 119.705 127.46 120.085 ;
      POLYGON  125.06 121.37 125.06 121.78 124.805 121.78 124.805 121.45 124.885 121.37 125.06 121.37 ;
      RECT  127.07 119.375 126.89 120.29 ;
      RECT  127.46 119.375 127.25 119.705 ;
      RECT  127.46 119.705 127.25 120.085 ;
      RECT  125.27 123.36 125.06 122.95 ;
      RECT  127.67 124.365 127.46 124.035 ;
      RECT  124.625 123.45 124.55 121.745 ;
      RECT  124.71 122.865 124.625 122.455 ;
      RECT  125.63 124.365 125.45 123.45 ;
      POLYGON  124.625 124.365 124.625 124.035 125.06 124.035 125.06 123.655 124.625 123.655 124.625 123.45 124.55 123.45 124.55 124.365 124.625 124.365 ;
      RECT  124.55 123.45 124.34 121.745 ;
      POLYGON  125.06 123.36 125.06 122.95 124.885 122.95 124.805 123.03 124.805 123.36 125.06 123.36 ;
      RECT  127.67 123.45 127.46 121.745 ;
      RECT  125.99 124.365 125.81 123.45 ;
      RECT  127.07 123.45 126.89 121.745 ;
      RECT  125.27 122.37 125.06 121.96 ;
      RECT  124.55 123.655 124.34 123.45 ;
      RECT  127.46 123.45 127.25 121.745 ;
      RECT  125.27 124.035 125.06 123.655 ;
      RECT  126.71 123.45 126.53 121.745 ;
      RECT  125.99 123.45 125.81 121.745 ;
      RECT  126.71 124.365 126.53 123.45 ;
      RECT  124.55 124.365 124.34 124.035 ;
      RECT  126.35 123.45 126.17 121.745 ;
      RECT  126.35 124.365 126.17 123.45 ;
      RECT  127.67 123.655 127.46 123.45 ;
      RECT  124.55 124.035 124.34 123.655 ;
      RECT  125.63 123.45 125.45 121.745 ;
      RECT  127.46 123.655 127.25 123.45 ;
      RECT  127.67 124.035 127.46 123.655 ;
      POLYGON  125.06 122.37 125.06 121.96 124.805 121.96 124.805 122.29 124.885 122.37 125.06 122.37 ;
      RECT  127.07 124.365 126.89 123.45 ;
      RECT  127.46 124.365 127.25 124.035 ;
      RECT  127.46 124.035 127.25 123.655 ;
      RECT  129.65 92.73 129.86 93.14 ;
      RECT  127.25 91.725 127.46 92.055 ;
      RECT  130.295 92.64 130.37 94.345 ;
      RECT  130.21 93.225 130.295 93.635 ;
      RECT  129.29 91.725 129.47 92.64 ;
      POLYGON  130.295 91.725 130.295 92.055 129.86 92.055 129.86 92.435 130.295 92.435 130.295 92.64 130.37 92.64 130.37 91.725 130.295 91.725 ;
      RECT  130.37 92.64 130.58 94.345 ;
      POLYGON  129.86 92.73 129.86 93.14 130.035 93.14 130.115 93.06 130.115 92.73 129.86 92.73 ;
      RECT  127.25 92.64 127.46 94.345 ;
      RECT  128.93 91.725 129.11 92.64 ;
      RECT  127.85 92.64 128.03 94.345 ;
      RECT  129.65 93.72 129.86 94.13 ;
      RECT  130.37 92.435 130.58 92.64 ;
      RECT  127.46 92.64 127.67 94.345 ;
      RECT  129.65 92.055 129.86 92.435 ;
      RECT  128.21 92.64 128.39 94.345 ;
      RECT  128.93 92.64 129.11 94.345 ;
      RECT  128.21 91.725 128.39 92.64 ;
      RECT  130.37 91.725 130.58 92.055 ;
      RECT  128.57 92.64 128.75 94.345 ;
      RECT  128.57 91.725 128.75 92.64 ;
      RECT  127.25 92.435 127.46 92.64 ;
      RECT  130.37 92.055 130.58 92.435 ;
      RECT  129.29 92.64 129.47 94.345 ;
      RECT  127.46 92.435 127.67 92.64 ;
      RECT  127.25 92.055 127.46 92.435 ;
      POLYGON  129.86 93.72 129.86 94.13 130.115 94.13 130.115 93.8 130.035 93.72 129.86 93.72 ;
      RECT  127.85 91.725 128.03 92.64 ;
      RECT  127.46 91.725 127.67 92.055 ;
      RECT  127.46 92.055 127.67 92.435 ;
      RECT  129.65 95.71 129.86 95.3 ;
      RECT  127.25 96.715 127.46 96.385 ;
      RECT  130.295 95.8 130.37 94.095 ;
      RECT  130.21 95.215 130.295 94.805 ;
      RECT  129.29 96.715 129.47 95.8 ;
      POLYGON  130.295 96.715 130.295 96.385 129.86 96.385 129.86 96.005 130.295 96.005 130.295 95.8 130.37 95.8 130.37 96.715 130.295 96.715 ;
      RECT  130.37 95.8 130.58 94.095 ;
      POLYGON  129.86 95.71 129.86 95.3 130.035 95.3 130.115 95.38 130.115 95.71 129.86 95.71 ;
      RECT  127.25 95.8 127.46 94.095 ;
      RECT  128.93 96.715 129.11 95.8 ;
      RECT  127.85 95.8 128.03 94.095 ;
      RECT  129.65 94.72 129.86 94.31 ;
      RECT  130.37 96.005 130.58 95.8 ;
      RECT  127.46 95.8 127.67 94.095 ;
      RECT  129.65 96.385 129.86 96.005 ;
      RECT  128.21 95.8 128.39 94.095 ;
      RECT  128.93 95.8 129.11 94.095 ;
      RECT  128.21 96.715 128.39 95.8 ;
      RECT  130.37 96.715 130.58 96.385 ;
      RECT  128.57 95.8 128.75 94.095 ;
      RECT  128.57 96.715 128.75 95.8 ;
      RECT  127.25 96.005 127.46 95.8 ;
      RECT  130.37 96.385 130.58 96.005 ;
      RECT  129.29 95.8 129.47 94.095 ;
      RECT  127.46 96.005 127.67 95.8 ;
      RECT  127.25 96.385 127.46 96.005 ;
      POLYGON  129.86 94.72 129.86 94.31 130.115 94.31 130.115 94.64 130.035 94.72 129.86 94.72 ;
      RECT  127.85 96.715 128.03 95.8 ;
      RECT  127.46 96.715 127.67 96.385 ;
      RECT  127.46 96.385 127.67 96.005 ;
      RECT  129.65 96.68 129.86 97.09 ;
      RECT  127.25 95.675 127.46 96.005 ;
      RECT  130.295 96.59 130.37 98.295 ;
      RECT  130.21 97.175 130.295 97.585 ;
      RECT  129.29 95.675 129.47 96.59 ;
      POLYGON  130.295 95.675 130.295 96.005 129.86 96.005 129.86 96.385 130.295 96.385 130.295 96.59 130.37 96.59 130.37 95.675 130.295 95.675 ;
      RECT  130.37 96.59 130.58 98.295 ;
      POLYGON  129.86 96.68 129.86 97.09 130.035 97.09 130.115 97.01 130.115 96.68 129.86 96.68 ;
      RECT  127.25 96.59 127.46 98.295 ;
      RECT  128.93 95.675 129.11 96.59 ;
      RECT  127.85 96.59 128.03 98.295 ;
      RECT  129.65 97.67 129.86 98.08 ;
      RECT  130.37 96.385 130.58 96.59 ;
      RECT  127.46 96.59 127.67 98.295 ;
      RECT  129.65 96.005 129.86 96.385 ;
      RECT  128.21 96.59 128.39 98.295 ;
      RECT  128.93 96.59 129.11 98.295 ;
      RECT  128.21 95.675 128.39 96.59 ;
      RECT  130.37 95.675 130.58 96.005 ;
      RECT  128.57 96.59 128.75 98.295 ;
      RECT  128.57 95.675 128.75 96.59 ;
      RECT  127.25 96.385 127.46 96.59 ;
      RECT  130.37 96.005 130.58 96.385 ;
      RECT  129.29 96.59 129.47 98.295 ;
      RECT  127.46 96.385 127.67 96.59 ;
      RECT  127.25 96.005 127.46 96.385 ;
      POLYGON  129.86 97.67 129.86 98.08 130.115 98.08 130.115 97.75 130.035 97.67 129.86 97.67 ;
      RECT  127.85 95.675 128.03 96.59 ;
      RECT  127.46 95.675 127.67 96.005 ;
      RECT  127.46 96.005 127.67 96.385 ;
      RECT  129.65 99.66 129.86 99.25 ;
      RECT  127.25 100.665 127.46 100.335 ;
      RECT  130.295 99.75 130.37 98.045 ;
      RECT  130.21 99.165 130.295 98.755 ;
      RECT  129.29 100.665 129.47 99.75 ;
      POLYGON  130.295 100.665 130.295 100.335 129.86 100.335 129.86 99.955 130.295 99.955 130.295 99.75 130.37 99.75 130.37 100.665 130.295 100.665 ;
      RECT  130.37 99.75 130.58 98.045 ;
      POLYGON  129.86 99.66 129.86 99.25 130.035 99.25 130.115 99.33 130.115 99.66 129.86 99.66 ;
      RECT  127.25 99.75 127.46 98.045 ;
      RECT  128.93 100.665 129.11 99.75 ;
      RECT  127.85 99.75 128.03 98.045 ;
      RECT  129.65 98.67 129.86 98.26 ;
      RECT  130.37 99.955 130.58 99.75 ;
      RECT  127.46 99.75 127.67 98.045 ;
      RECT  129.65 100.335 129.86 99.955 ;
      RECT  128.21 99.75 128.39 98.045 ;
      RECT  128.93 99.75 129.11 98.045 ;
      RECT  128.21 100.665 128.39 99.75 ;
      RECT  130.37 100.665 130.58 100.335 ;
      RECT  128.57 99.75 128.75 98.045 ;
      RECT  128.57 100.665 128.75 99.75 ;
      RECT  127.25 99.955 127.46 99.75 ;
      RECT  130.37 100.335 130.58 99.955 ;
      RECT  129.29 99.75 129.47 98.045 ;
      RECT  127.46 99.955 127.67 99.75 ;
      RECT  127.25 100.335 127.46 99.955 ;
      POLYGON  129.86 98.67 129.86 98.26 130.115 98.26 130.115 98.59 130.035 98.67 129.86 98.67 ;
      RECT  127.85 100.665 128.03 99.75 ;
      RECT  127.46 100.665 127.67 100.335 ;
      RECT  127.46 100.335 127.67 99.955 ;
      RECT  129.65 100.63 129.86 101.04 ;
      RECT  127.25 99.625 127.46 99.955 ;
      RECT  130.295 100.54 130.37 102.245 ;
      RECT  130.21 101.125 130.295 101.535 ;
      RECT  129.29 99.625 129.47 100.54 ;
      POLYGON  130.295 99.625 130.295 99.955 129.86 99.955 129.86 100.335 130.295 100.335 130.295 100.54 130.37 100.54 130.37 99.625 130.295 99.625 ;
      RECT  130.37 100.54 130.58 102.245 ;
      POLYGON  129.86 100.63 129.86 101.04 130.035 101.04 130.115 100.96 130.115 100.63 129.86 100.63 ;
      RECT  127.25 100.54 127.46 102.245 ;
      RECT  128.93 99.625 129.11 100.54 ;
      RECT  127.85 100.54 128.03 102.245 ;
      RECT  129.65 101.62 129.86 102.03 ;
      RECT  130.37 100.335 130.58 100.54 ;
      RECT  127.46 100.54 127.67 102.245 ;
      RECT  129.65 99.955 129.86 100.335 ;
      RECT  128.21 100.54 128.39 102.245 ;
      RECT  128.93 100.54 129.11 102.245 ;
      RECT  128.21 99.625 128.39 100.54 ;
      RECT  130.37 99.625 130.58 99.955 ;
      RECT  128.57 100.54 128.75 102.245 ;
      RECT  128.57 99.625 128.75 100.54 ;
      RECT  127.25 100.335 127.46 100.54 ;
      RECT  130.37 99.955 130.58 100.335 ;
      RECT  129.29 100.54 129.47 102.245 ;
      RECT  127.46 100.335 127.67 100.54 ;
      RECT  127.25 99.955 127.46 100.335 ;
      POLYGON  129.86 101.62 129.86 102.03 130.115 102.03 130.115 101.7 130.035 101.62 129.86 101.62 ;
      RECT  127.85 99.625 128.03 100.54 ;
      RECT  127.46 99.625 127.67 99.955 ;
      RECT  127.46 99.955 127.67 100.335 ;
      RECT  129.65 103.61 129.86 103.2 ;
      RECT  127.25 104.615 127.46 104.285 ;
      RECT  130.295 103.7 130.37 101.995 ;
      RECT  130.21 103.115 130.295 102.705 ;
      RECT  129.29 104.615 129.47 103.7 ;
      POLYGON  130.295 104.615 130.295 104.285 129.86 104.285 129.86 103.905 130.295 103.905 130.295 103.7 130.37 103.7 130.37 104.615 130.295 104.615 ;
      RECT  130.37 103.7 130.58 101.995 ;
      POLYGON  129.86 103.61 129.86 103.2 130.035 103.2 130.115 103.28 130.115 103.61 129.86 103.61 ;
      RECT  127.25 103.7 127.46 101.995 ;
      RECT  128.93 104.615 129.11 103.7 ;
      RECT  127.85 103.7 128.03 101.995 ;
      RECT  129.65 102.62 129.86 102.21 ;
      RECT  130.37 103.905 130.58 103.7 ;
      RECT  127.46 103.7 127.67 101.995 ;
      RECT  129.65 104.285 129.86 103.905 ;
      RECT  128.21 103.7 128.39 101.995 ;
      RECT  128.93 103.7 129.11 101.995 ;
      RECT  128.21 104.615 128.39 103.7 ;
      RECT  130.37 104.615 130.58 104.285 ;
      RECT  128.57 103.7 128.75 101.995 ;
      RECT  128.57 104.615 128.75 103.7 ;
      RECT  127.25 103.905 127.46 103.7 ;
      RECT  130.37 104.285 130.58 103.905 ;
      RECT  129.29 103.7 129.47 101.995 ;
      RECT  127.46 103.905 127.67 103.7 ;
      RECT  127.25 104.285 127.46 103.905 ;
      POLYGON  129.86 102.62 129.86 102.21 130.115 102.21 130.115 102.54 130.035 102.62 129.86 102.62 ;
      RECT  127.85 104.615 128.03 103.7 ;
      RECT  127.46 104.615 127.67 104.285 ;
      RECT  127.46 104.285 127.67 103.905 ;
      RECT  129.65 104.58 129.86 104.99 ;
      RECT  127.25 103.575 127.46 103.905 ;
      RECT  130.295 104.49 130.37 106.195 ;
      RECT  130.21 105.075 130.295 105.485 ;
      RECT  129.29 103.575 129.47 104.49 ;
      POLYGON  130.295 103.575 130.295 103.905 129.86 103.905 129.86 104.285 130.295 104.285 130.295 104.49 130.37 104.49 130.37 103.575 130.295 103.575 ;
      RECT  130.37 104.49 130.58 106.195 ;
      POLYGON  129.86 104.58 129.86 104.99 130.035 104.99 130.115 104.91 130.115 104.58 129.86 104.58 ;
      RECT  127.25 104.49 127.46 106.195 ;
      RECT  128.93 103.575 129.11 104.49 ;
      RECT  127.85 104.49 128.03 106.195 ;
      RECT  129.65 105.57 129.86 105.98 ;
      RECT  130.37 104.285 130.58 104.49 ;
      RECT  127.46 104.49 127.67 106.195 ;
      RECT  129.65 103.905 129.86 104.285 ;
      RECT  128.21 104.49 128.39 106.195 ;
      RECT  128.93 104.49 129.11 106.195 ;
      RECT  128.21 103.575 128.39 104.49 ;
      RECT  130.37 103.575 130.58 103.905 ;
      RECT  128.57 104.49 128.75 106.195 ;
      RECT  128.57 103.575 128.75 104.49 ;
      RECT  127.25 104.285 127.46 104.49 ;
      RECT  130.37 103.905 130.58 104.285 ;
      RECT  129.29 104.49 129.47 106.195 ;
      RECT  127.46 104.285 127.67 104.49 ;
      RECT  127.25 103.905 127.46 104.285 ;
      POLYGON  129.86 105.57 129.86 105.98 130.115 105.98 130.115 105.65 130.035 105.57 129.86 105.57 ;
      RECT  127.85 103.575 128.03 104.49 ;
      RECT  127.46 103.575 127.67 103.905 ;
      RECT  127.46 103.905 127.67 104.285 ;
      RECT  129.65 107.56 129.86 107.15 ;
      RECT  127.25 108.565 127.46 108.235 ;
      RECT  130.295 107.65 130.37 105.945 ;
      RECT  130.21 107.065 130.295 106.655 ;
      RECT  129.29 108.565 129.47 107.65 ;
      POLYGON  130.295 108.565 130.295 108.235 129.86 108.235 129.86 107.855 130.295 107.855 130.295 107.65 130.37 107.65 130.37 108.565 130.295 108.565 ;
      RECT  130.37 107.65 130.58 105.945 ;
      POLYGON  129.86 107.56 129.86 107.15 130.035 107.15 130.115 107.23 130.115 107.56 129.86 107.56 ;
      RECT  127.25 107.65 127.46 105.945 ;
      RECT  128.93 108.565 129.11 107.65 ;
      RECT  127.85 107.65 128.03 105.945 ;
      RECT  129.65 106.57 129.86 106.16 ;
      RECT  130.37 107.855 130.58 107.65 ;
      RECT  127.46 107.65 127.67 105.945 ;
      RECT  129.65 108.235 129.86 107.855 ;
      RECT  128.21 107.65 128.39 105.945 ;
      RECT  128.93 107.65 129.11 105.945 ;
      RECT  128.21 108.565 128.39 107.65 ;
      RECT  130.37 108.565 130.58 108.235 ;
      RECT  128.57 107.65 128.75 105.945 ;
      RECT  128.57 108.565 128.75 107.65 ;
      RECT  127.25 107.855 127.46 107.65 ;
      RECT  130.37 108.235 130.58 107.855 ;
      RECT  129.29 107.65 129.47 105.945 ;
      RECT  127.46 107.855 127.67 107.65 ;
      RECT  127.25 108.235 127.46 107.855 ;
      POLYGON  129.86 106.57 129.86 106.16 130.115 106.16 130.115 106.49 130.035 106.57 129.86 106.57 ;
      RECT  127.85 108.565 128.03 107.65 ;
      RECT  127.46 108.565 127.67 108.235 ;
      RECT  127.46 108.235 127.67 107.855 ;
      RECT  129.65 108.53 129.86 108.94 ;
      RECT  127.25 107.525 127.46 107.855 ;
      RECT  130.295 108.44 130.37 110.145 ;
      RECT  130.21 109.025 130.295 109.435 ;
      RECT  129.29 107.525 129.47 108.44 ;
      POLYGON  130.295 107.525 130.295 107.855 129.86 107.855 129.86 108.235 130.295 108.235 130.295 108.44 130.37 108.44 130.37 107.525 130.295 107.525 ;
      RECT  130.37 108.44 130.58 110.145 ;
      POLYGON  129.86 108.53 129.86 108.94 130.035 108.94 130.115 108.86 130.115 108.53 129.86 108.53 ;
      RECT  127.25 108.44 127.46 110.145 ;
      RECT  128.93 107.525 129.11 108.44 ;
      RECT  127.85 108.44 128.03 110.145 ;
      RECT  129.65 109.52 129.86 109.93 ;
      RECT  130.37 108.235 130.58 108.44 ;
      RECT  127.46 108.44 127.67 110.145 ;
      RECT  129.65 107.855 129.86 108.235 ;
      RECT  128.21 108.44 128.39 110.145 ;
      RECT  128.93 108.44 129.11 110.145 ;
      RECT  128.21 107.525 128.39 108.44 ;
      RECT  130.37 107.525 130.58 107.855 ;
      RECT  128.57 108.44 128.75 110.145 ;
      RECT  128.57 107.525 128.75 108.44 ;
      RECT  127.25 108.235 127.46 108.44 ;
      RECT  130.37 107.855 130.58 108.235 ;
      RECT  129.29 108.44 129.47 110.145 ;
      RECT  127.46 108.235 127.67 108.44 ;
      RECT  127.25 107.855 127.46 108.235 ;
      POLYGON  129.86 109.52 129.86 109.93 130.115 109.93 130.115 109.6 130.035 109.52 129.86 109.52 ;
      RECT  127.85 107.525 128.03 108.44 ;
      RECT  127.46 107.525 127.67 107.855 ;
      RECT  127.46 107.855 127.67 108.235 ;
      RECT  129.65 111.51 129.86 111.1 ;
      RECT  127.25 112.515 127.46 112.185 ;
      RECT  130.295 111.6 130.37 109.895 ;
      RECT  130.21 111.015 130.295 110.605 ;
      RECT  129.29 112.515 129.47 111.6 ;
      POLYGON  130.295 112.515 130.295 112.185 129.86 112.185 129.86 111.805 130.295 111.805 130.295 111.6 130.37 111.6 130.37 112.515 130.295 112.515 ;
      RECT  130.37 111.6 130.58 109.895 ;
      POLYGON  129.86 111.51 129.86 111.1 130.035 111.1 130.115 111.18 130.115 111.51 129.86 111.51 ;
      RECT  127.25 111.6 127.46 109.895 ;
      RECT  128.93 112.515 129.11 111.6 ;
      RECT  127.85 111.6 128.03 109.895 ;
      RECT  129.65 110.52 129.86 110.11 ;
      RECT  130.37 111.805 130.58 111.6 ;
      RECT  127.46 111.6 127.67 109.895 ;
      RECT  129.65 112.185 129.86 111.805 ;
      RECT  128.21 111.6 128.39 109.895 ;
      RECT  128.93 111.6 129.11 109.895 ;
      RECT  128.21 112.515 128.39 111.6 ;
      RECT  130.37 112.515 130.58 112.185 ;
      RECT  128.57 111.6 128.75 109.895 ;
      RECT  128.57 112.515 128.75 111.6 ;
      RECT  127.25 111.805 127.46 111.6 ;
      RECT  130.37 112.185 130.58 111.805 ;
      RECT  129.29 111.6 129.47 109.895 ;
      RECT  127.46 111.805 127.67 111.6 ;
      RECT  127.25 112.185 127.46 111.805 ;
      POLYGON  129.86 110.52 129.86 110.11 130.115 110.11 130.115 110.44 130.035 110.52 129.86 110.52 ;
      RECT  127.85 112.515 128.03 111.6 ;
      RECT  127.46 112.515 127.67 112.185 ;
      RECT  127.46 112.185 127.67 111.805 ;
      RECT  129.65 112.48 129.86 112.89 ;
      RECT  127.25 111.475 127.46 111.805 ;
      RECT  130.295 112.39 130.37 114.095 ;
      RECT  130.21 112.975 130.295 113.385 ;
      RECT  129.29 111.475 129.47 112.39 ;
      POLYGON  130.295 111.475 130.295 111.805 129.86 111.805 129.86 112.185 130.295 112.185 130.295 112.39 130.37 112.39 130.37 111.475 130.295 111.475 ;
      RECT  130.37 112.39 130.58 114.095 ;
      POLYGON  129.86 112.48 129.86 112.89 130.035 112.89 130.115 112.81 130.115 112.48 129.86 112.48 ;
      RECT  127.25 112.39 127.46 114.095 ;
      RECT  128.93 111.475 129.11 112.39 ;
      RECT  127.85 112.39 128.03 114.095 ;
      RECT  129.65 113.47 129.86 113.88 ;
      RECT  130.37 112.185 130.58 112.39 ;
      RECT  127.46 112.39 127.67 114.095 ;
      RECT  129.65 111.805 129.86 112.185 ;
      RECT  128.21 112.39 128.39 114.095 ;
      RECT  128.93 112.39 129.11 114.095 ;
      RECT  128.21 111.475 128.39 112.39 ;
      RECT  130.37 111.475 130.58 111.805 ;
      RECT  128.57 112.39 128.75 114.095 ;
      RECT  128.57 111.475 128.75 112.39 ;
      RECT  127.25 112.185 127.46 112.39 ;
      RECT  130.37 111.805 130.58 112.185 ;
      RECT  129.29 112.39 129.47 114.095 ;
      RECT  127.46 112.185 127.67 112.39 ;
      RECT  127.25 111.805 127.46 112.185 ;
      POLYGON  129.86 113.47 129.86 113.88 130.115 113.88 130.115 113.55 130.035 113.47 129.86 113.47 ;
      RECT  127.85 111.475 128.03 112.39 ;
      RECT  127.46 111.475 127.67 111.805 ;
      RECT  127.46 111.805 127.67 112.185 ;
      RECT  129.65 115.46 129.86 115.05 ;
      RECT  127.25 116.465 127.46 116.135 ;
      RECT  130.295 115.55 130.37 113.845 ;
      RECT  130.21 114.965 130.295 114.555 ;
      RECT  129.29 116.465 129.47 115.55 ;
      POLYGON  130.295 116.465 130.295 116.135 129.86 116.135 129.86 115.755 130.295 115.755 130.295 115.55 130.37 115.55 130.37 116.465 130.295 116.465 ;
      RECT  130.37 115.55 130.58 113.845 ;
      POLYGON  129.86 115.46 129.86 115.05 130.035 115.05 130.115 115.13 130.115 115.46 129.86 115.46 ;
      RECT  127.25 115.55 127.46 113.845 ;
      RECT  128.93 116.465 129.11 115.55 ;
      RECT  127.85 115.55 128.03 113.845 ;
      RECT  129.65 114.47 129.86 114.06 ;
      RECT  130.37 115.755 130.58 115.55 ;
      RECT  127.46 115.55 127.67 113.845 ;
      RECT  129.65 116.135 129.86 115.755 ;
      RECT  128.21 115.55 128.39 113.845 ;
      RECT  128.93 115.55 129.11 113.845 ;
      RECT  128.21 116.465 128.39 115.55 ;
      RECT  130.37 116.465 130.58 116.135 ;
      RECT  128.57 115.55 128.75 113.845 ;
      RECT  128.57 116.465 128.75 115.55 ;
      RECT  127.25 115.755 127.46 115.55 ;
      RECT  130.37 116.135 130.58 115.755 ;
      RECT  129.29 115.55 129.47 113.845 ;
      RECT  127.46 115.755 127.67 115.55 ;
      RECT  127.25 116.135 127.46 115.755 ;
      POLYGON  129.86 114.47 129.86 114.06 130.115 114.06 130.115 114.39 130.035 114.47 129.86 114.47 ;
      RECT  127.85 116.465 128.03 115.55 ;
      RECT  127.46 116.465 127.67 116.135 ;
      RECT  127.46 116.135 127.67 115.755 ;
      RECT  129.65 116.43 129.86 116.84 ;
      RECT  127.25 115.425 127.46 115.755 ;
      RECT  130.295 116.34 130.37 118.045 ;
      RECT  130.21 116.925 130.295 117.335 ;
      RECT  129.29 115.425 129.47 116.34 ;
      POLYGON  130.295 115.425 130.295 115.755 129.86 115.755 129.86 116.135 130.295 116.135 130.295 116.34 130.37 116.34 130.37 115.425 130.295 115.425 ;
      RECT  130.37 116.34 130.58 118.045 ;
      POLYGON  129.86 116.43 129.86 116.84 130.035 116.84 130.115 116.76 130.115 116.43 129.86 116.43 ;
      RECT  127.25 116.34 127.46 118.045 ;
      RECT  128.93 115.425 129.11 116.34 ;
      RECT  127.85 116.34 128.03 118.045 ;
      RECT  129.65 117.42 129.86 117.83 ;
      RECT  130.37 116.135 130.58 116.34 ;
      RECT  127.46 116.34 127.67 118.045 ;
      RECT  129.65 115.755 129.86 116.135 ;
      RECT  128.21 116.34 128.39 118.045 ;
      RECT  128.93 116.34 129.11 118.045 ;
      RECT  128.21 115.425 128.39 116.34 ;
      RECT  130.37 115.425 130.58 115.755 ;
      RECT  128.57 116.34 128.75 118.045 ;
      RECT  128.57 115.425 128.75 116.34 ;
      RECT  127.25 116.135 127.46 116.34 ;
      RECT  130.37 115.755 130.58 116.135 ;
      RECT  129.29 116.34 129.47 118.045 ;
      RECT  127.46 116.135 127.67 116.34 ;
      RECT  127.25 115.755 127.46 116.135 ;
      POLYGON  129.86 117.42 129.86 117.83 130.115 117.83 130.115 117.5 130.035 117.42 129.86 117.42 ;
      RECT  127.85 115.425 128.03 116.34 ;
      RECT  127.46 115.425 127.67 115.755 ;
      RECT  127.46 115.755 127.67 116.135 ;
      RECT  129.65 119.41 129.86 119.0 ;
      RECT  127.25 120.415 127.46 120.085 ;
      RECT  130.295 119.5 130.37 117.795 ;
      RECT  130.21 118.915 130.295 118.505 ;
      RECT  129.29 120.415 129.47 119.5 ;
      POLYGON  130.295 120.415 130.295 120.085 129.86 120.085 129.86 119.705 130.295 119.705 130.295 119.5 130.37 119.5 130.37 120.415 130.295 120.415 ;
      RECT  130.37 119.5 130.58 117.795 ;
      POLYGON  129.86 119.41 129.86 119.0 130.035 119.0 130.115 119.08 130.115 119.41 129.86 119.41 ;
      RECT  127.25 119.5 127.46 117.795 ;
      RECT  128.93 120.415 129.11 119.5 ;
      RECT  127.85 119.5 128.03 117.795 ;
      RECT  129.65 118.42 129.86 118.01 ;
      RECT  130.37 119.705 130.58 119.5 ;
      RECT  127.46 119.5 127.67 117.795 ;
      RECT  129.65 120.085 129.86 119.705 ;
      RECT  128.21 119.5 128.39 117.795 ;
      RECT  128.93 119.5 129.11 117.795 ;
      RECT  128.21 120.415 128.39 119.5 ;
      RECT  130.37 120.415 130.58 120.085 ;
      RECT  128.57 119.5 128.75 117.795 ;
      RECT  128.57 120.415 128.75 119.5 ;
      RECT  127.25 119.705 127.46 119.5 ;
      RECT  130.37 120.085 130.58 119.705 ;
      RECT  129.29 119.5 129.47 117.795 ;
      RECT  127.46 119.705 127.67 119.5 ;
      RECT  127.25 120.085 127.46 119.705 ;
      POLYGON  129.86 118.42 129.86 118.01 130.115 118.01 130.115 118.34 130.035 118.42 129.86 118.42 ;
      RECT  127.85 120.415 128.03 119.5 ;
      RECT  127.46 120.415 127.67 120.085 ;
      RECT  127.46 120.085 127.67 119.705 ;
      RECT  129.65 120.38 129.86 120.79 ;
      RECT  127.25 119.375 127.46 119.705 ;
      RECT  130.295 120.29 130.37 121.995 ;
      RECT  130.21 120.875 130.295 121.285 ;
      RECT  129.29 119.375 129.47 120.29 ;
      POLYGON  130.295 119.375 130.295 119.705 129.86 119.705 129.86 120.085 130.295 120.085 130.295 120.29 130.37 120.29 130.37 119.375 130.295 119.375 ;
      RECT  130.37 120.29 130.58 121.995 ;
      POLYGON  129.86 120.38 129.86 120.79 130.035 120.79 130.115 120.71 130.115 120.38 129.86 120.38 ;
      RECT  127.25 120.29 127.46 121.995 ;
      RECT  128.93 119.375 129.11 120.29 ;
      RECT  127.85 120.29 128.03 121.995 ;
      RECT  129.65 121.37 129.86 121.78 ;
      RECT  130.37 120.085 130.58 120.29 ;
      RECT  127.46 120.29 127.67 121.995 ;
      RECT  129.65 119.705 129.86 120.085 ;
      RECT  128.21 120.29 128.39 121.995 ;
      RECT  128.93 120.29 129.11 121.995 ;
      RECT  128.21 119.375 128.39 120.29 ;
      RECT  130.37 119.375 130.58 119.705 ;
      RECT  128.57 120.29 128.75 121.995 ;
      RECT  128.57 119.375 128.75 120.29 ;
      RECT  127.25 120.085 127.46 120.29 ;
      RECT  130.37 119.705 130.58 120.085 ;
      RECT  129.29 120.29 129.47 121.995 ;
      RECT  127.46 120.085 127.67 120.29 ;
      RECT  127.25 119.705 127.46 120.085 ;
      POLYGON  129.86 121.37 129.86 121.78 130.115 121.78 130.115 121.45 130.035 121.37 129.86 121.37 ;
      RECT  127.85 119.375 128.03 120.29 ;
      RECT  127.46 119.375 127.67 119.705 ;
      RECT  127.46 119.705 127.67 120.085 ;
      RECT  129.65 123.36 129.86 122.95 ;
      RECT  127.25 124.365 127.46 124.035 ;
      RECT  130.295 123.45 130.37 121.745 ;
      RECT  130.21 122.865 130.295 122.455 ;
      RECT  129.29 124.365 129.47 123.45 ;
      POLYGON  130.295 124.365 130.295 124.035 129.86 124.035 129.86 123.655 130.295 123.655 130.295 123.45 130.37 123.45 130.37 124.365 130.295 124.365 ;
      RECT  130.37 123.45 130.58 121.745 ;
      POLYGON  129.86 123.36 129.86 122.95 130.035 122.95 130.115 123.03 130.115 123.36 129.86 123.36 ;
      RECT  127.25 123.45 127.46 121.745 ;
      RECT  128.93 124.365 129.11 123.45 ;
      RECT  127.85 123.45 128.03 121.745 ;
      RECT  129.65 122.37 129.86 121.96 ;
      RECT  130.37 123.655 130.58 123.45 ;
      RECT  127.46 123.45 127.67 121.745 ;
      RECT  129.65 124.035 129.86 123.655 ;
      RECT  128.21 123.45 128.39 121.745 ;
      RECT  128.93 123.45 129.11 121.745 ;
      RECT  128.21 124.365 128.39 123.45 ;
      RECT  130.37 124.365 130.58 124.035 ;
      RECT  128.57 123.45 128.75 121.745 ;
      RECT  128.57 124.365 128.75 123.45 ;
      RECT  127.25 123.655 127.46 123.45 ;
      RECT  130.37 124.035 130.58 123.655 ;
      RECT  129.29 123.45 129.47 121.745 ;
      RECT  127.46 123.655 127.67 123.45 ;
      RECT  127.25 124.035 127.46 123.655 ;
      POLYGON  129.86 122.37 129.86 121.96 130.115 121.96 130.115 122.29 130.035 122.37 129.86 122.37 ;
      RECT  127.85 124.365 128.03 123.45 ;
      RECT  127.46 124.365 127.67 124.035 ;
      RECT  127.46 124.035 127.67 123.655 ;
      RECT  131.51 92.73 131.3 93.14 ;
      RECT  133.91 91.725 133.7 92.055 ;
      RECT  130.865 92.64 130.79 94.345 ;
      RECT  130.95 93.225 130.865 93.635 ;
      RECT  131.87 91.725 131.69 92.64 ;
      POLYGON  130.865 91.725 130.865 92.055 131.3 92.055 131.3 92.435 130.865 92.435 130.865 92.64 130.79 92.64 130.79 91.725 130.865 91.725 ;
      RECT  130.79 92.64 130.58 94.345 ;
      POLYGON  131.3 92.73 131.3 93.14 131.125 93.14 131.045 93.06 131.045 92.73 131.3 92.73 ;
      RECT  133.91 92.64 133.7 94.345 ;
      RECT  132.23 91.725 132.05 92.64 ;
      RECT  133.31 92.64 133.13 94.345 ;
      RECT  131.51 93.72 131.3 94.13 ;
      RECT  130.79 92.435 130.58 92.64 ;
      RECT  133.7 92.64 133.49 94.345 ;
      RECT  131.51 92.055 131.3 92.435 ;
      RECT  132.95 92.64 132.77 94.345 ;
      RECT  132.23 92.64 132.05 94.345 ;
      RECT  132.95 91.725 132.77 92.64 ;
      RECT  130.79 91.725 130.58 92.055 ;
      RECT  132.59 92.64 132.41 94.345 ;
      RECT  132.59 91.725 132.41 92.64 ;
      RECT  133.91 92.435 133.7 92.64 ;
      RECT  130.79 92.055 130.58 92.435 ;
      RECT  131.87 92.64 131.69 94.345 ;
      RECT  133.7 92.435 133.49 92.64 ;
      RECT  133.91 92.055 133.7 92.435 ;
      POLYGON  131.3 93.72 131.3 94.13 131.045 94.13 131.045 93.8 131.125 93.72 131.3 93.72 ;
      RECT  133.31 91.725 133.13 92.64 ;
      RECT  133.7 91.725 133.49 92.055 ;
      RECT  133.7 92.055 133.49 92.435 ;
      RECT  131.51 95.71 131.3 95.3 ;
      RECT  133.91 96.715 133.7 96.385 ;
      RECT  130.865 95.8 130.79 94.095 ;
      RECT  130.95 95.215 130.865 94.805 ;
      RECT  131.87 96.715 131.69 95.8 ;
      POLYGON  130.865 96.715 130.865 96.385 131.3 96.385 131.3 96.005 130.865 96.005 130.865 95.8 130.79 95.8 130.79 96.715 130.865 96.715 ;
      RECT  130.79 95.8 130.58 94.095 ;
      POLYGON  131.3 95.71 131.3 95.3 131.125 95.3 131.045 95.38 131.045 95.71 131.3 95.71 ;
      RECT  133.91 95.8 133.7 94.095 ;
      RECT  132.23 96.715 132.05 95.8 ;
      RECT  133.31 95.8 133.13 94.095 ;
      RECT  131.51 94.72 131.3 94.31 ;
      RECT  130.79 96.005 130.58 95.8 ;
      RECT  133.7 95.8 133.49 94.095 ;
      RECT  131.51 96.385 131.3 96.005 ;
      RECT  132.95 95.8 132.77 94.095 ;
      RECT  132.23 95.8 132.05 94.095 ;
      RECT  132.95 96.715 132.77 95.8 ;
      RECT  130.79 96.715 130.58 96.385 ;
      RECT  132.59 95.8 132.41 94.095 ;
      RECT  132.59 96.715 132.41 95.8 ;
      RECT  133.91 96.005 133.7 95.8 ;
      RECT  130.79 96.385 130.58 96.005 ;
      RECT  131.87 95.8 131.69 94.095 ;
      RECT  133.7 96.005 133.49 95.8 ;
      RECT  133.91 96.385 133.7 96.005 ;
      POLYGON  131.3 94.72 131.3 94.31 131.045 94.31 131.045 94.64 131.125 94.72 131.3 94.72 ;
      RECT  133.31 96.715 133.13 95.8 ;
      RECT  133.7 96.715 133.49 96.385 ;
      RECT  133.7 96.385 133.49 96.005 ;
      RECT  131.51 96.68 131.3 97.09 ;
      RECT  133.91 95.675 133.7 96.005 ;
      RECT  130.865 96.59 130.79 98.295 ;
      RECT  130.95 97.175 130.865 97.585 ;
      RECT  131.87 95.675 131.69 96.59 ;
      POLYGON  130.865 95.675 130.865 96.005 131.3 96.005 131.3 96.385 130.865 96.385 130.865 96.59 130.79 96.59 130.79 95.675 130.865 95.675 ;
      RECT  130.79 96.59 130.58 98.295 ;
      POLYGON  131.3 96.68 131.3 97.09 131.125 97.09 131.045 97.01 131.045 96.68 131.3 96.68 ;
      RECT  133.91 96.59 133.7 98.295 ;
      RECT  132.23 95.675 132.05 96.59 ;
      RECT  133.31 96.59 133.13 98.295 ;
      RECT  131.51 97.67 131.3 98.08 ;
      RECT  130.79 96.385 130.58 96.59 ;
      RECT  133.7 96.59 133.49 98.295 ;
      RECT  131.51 96.005 131.3 96.385 ;
      RECT  132.95 96.59 132.77 98.295 ;
      RECT  132.23 96.59 132.05 98.295 ;
      RECT  132.95 95.675 132.77 96.59 ;
      RECT  130.79 95.675 130.58 96.005 ;
      RECT  132.59 96.59 132.41 98.295 ;
      RECT  132.59 95.675 132.41 96.59 ;
      RECT  133.91 96.385 133.7 96.59 ;
      RECT  130.79 96.005 130.58 96.385 ;
      RECT  131.87 96.59 131.69 98.295 ;
      RECT  133.7 96.385 133.49 96.59 ;
      RECT  133.91 96.005 133.7 96.385 ;
      POLYGON  131.3 97.67 131.3 98.08 131.045 98.08 131.045 97.75 131.125 97.67 131.3 97.67 ;
      RECT  133.31 95.675 133.13 96.59 ;
      RECT  133.7 95.675 133.49 96.005 ;
      RECT  133.7 96.005 133.49 96.385 ;
      RECT  131.51 99.66 131.3 99.25 ;
      RECT  133.91 100.665 133.7 100.335 ;
      RECT  130.865 99.75 130.79 98.045 ;
      RECT  130.95 99.165 130.865 98.755 ;
      RECT  131.87 100.665 131.69 99.75 ;
      POLYGON  130.865 100.665 130.865 100.335 131.3 100.335 131.3 99.955 130.865 99.955 130.865 99.75 130.79 99.75 130.79 100.665 130.865 100.665 ;
      RECT  130.79 99.75 130.58 98.045 ;
      POLYGON  131.3 99.66 131.3 99.25 131.125 99.25 131.045 99.33 131.045 99.66 131.3 99.66 ;
      RECT  133.91 99.75 133.7 98.045 ;
      RECT  132.23 100.665 132.05 99.75 ;
      RECT  133.31 99.75 133.13 98.045 ;
      RECT  131.51 98.67 131.3 98.26 ;
      RECT  130.79 99.955 130.58 99.75 ;
      RECT  133.7 99.75 133.49 98.045 ;
      RECT  131.51 100.335 131.3 99.955 ;
      RECT  132.95 99.75 132.77 98.045 ;
      RECT  132.23 99.75 132.05 98.045 ;
      RECT  132.95 100.665 132.77 99.75 ;
      RECT  130.79 100.665 130.58 100.335 ;
      RECT  132.59 99.75 132.41 98.045 ;
      RECT  132.59 100.665 132.41 99.75 ;
      RECT  133.91 99.955 133.7 99.75 ;
      RECT  130.79 100.335 130.58 99.955 ;
      RECT  131.87 99.75 131.69 98.045 ;
      RECT  133.7 99.955 133.49 99.75 ;
      RECT  133.91 100.335 133.7 99.955 ;
      POLYGON  131.3 98.67 131.3 98.26 131.045 98.26 131.045 98.59 131.125 98.67 131.3 98.67 ;
      RECT  133.31 100.665 133.13 99.75 ;
      RECT  133.7 100.665 133.49 100.335 ;
      RECT  133.7 100.335 133.49 99.955 ;
      RECT  131.51 100.63 131.3 101.04 ;
      RECT  133.91 99.625 133.7 99.955 ;
      RECT  130.865 100.54 130.79 102.245 ;
      RECT  130.95 101.125 130.865 101.535 ;
      RECT  131.87 99.625 131.69 100.54 ;
      POLYGON  130.865 99.625 130.865 99.955 131.3 99.955 131.3 100.335 130.865 100.335 130.865 100.54 130.79 100.54 130.79 99.625 130.865 99.625 ;
      RECT  130.79 100.54 130.58 102.245 ;
      POLYGON  131.3 100.63 131.3 101.04 131.125 101.04 131.045 100.96 131.045 100.63 131.3 100.63 ;
      RECT  133.91 100.54 133.7 102.245 ;
      RECT  132.23 99.625 132.05 100.54 ;
      RECT  133.31 100.54 133.13 102.245 ;
      RECT  131.51 101.62 131.3 102.03 ;
      RECT  130.79 100.335 130.58 100.54 ;
      RECT  133.7 100.54 133.49 102.245 ;
      RECT  131.51 99.955 131.3 100.335 ;
      RECT  132.95 100.54 132.77 102.245 ;
      RECT  132.23 100.54 132.05 102.245 ;
      RECT  132.95 99.625 132.77 100.54 ;
      RECT  130.79 99.625 130.58 99.955 ;
      RECT  132.59 100.54 132.41 102.245 ;
      RECT  132.59 99.625 132.41 100.54 ;
      RECT  133.91 100.335 133.7 100.54 ;
      RECT  130.79 99.955 130.58 100.335 ;
      RECT  131.87 100.54 131.69 102.245 ;
      RECT  133.7 100.335 133.49 100.54 ;
      RECT  133.91 99.955 133.7 100.335 ;
      POLYGON  131.3 101.62 131.3 102.03 131.045 102.03 131.045 101.7 131.125 101.62 131.3 101.62 ;
      RECT  133.31 99.625 133.13 100.54 ;
      RECT  133.7 99.625 133.49 99.955 ;
      RECT  133.7 99.955 133.49 100.335 ;
      RECT  131.51 103.61 131.3 103.2 ;
      RECT  133.91 104.615 133.7 104.285 ;
      RECT  130.865 103.7 130.79 101.995 ;
      RECT  130.95 103.115 130.865 102.705 ;
      RECT  131.87 104.615 131.69 103.7 ;
      POLYGON  130.865 104.615 130.865 104.285 131.3 104.285 131.3 103.905 130.865 103.905 130.865 103.7 130.79 103.7 130.79 104.615 130.865 104.615 ;
      RECT  130.79 103.7 130.58 101.995 ;
      POLYGON  131.3 103.61 131.3 103.2 131.125 103.2 131.045 103.28 131.045 103.61 131.3 103.61 ;
      RECT  133.91 103.7 133.7 101.995 ;
      RECT  132.23 104.615 132.05 103.7 ;
      RECT  133.31 103.7 133.13 101.995 ;
      RECT  131.51 102.62 131.3 102.21 ;
      RECT  130.79 103.905 130.58 103.7 ;
      RECT  133.7 103.7 133.49 101.995 ;
      RECT  131.51 104.285 131.3 103.905 ;
      RECT  132.95 103.7 132.77 101.995 ;
      RECT  132.23 103.7 132.05 101.995 ;
      RECT  132.95 104.615 132.77 103.7 ;
      RECT  130.79 104.615 130.58 104.285 ;
      RECT  132.59 103.7 132.41 101.995 ;
      RECT  132.59 104.615 132.41 103.7 ;
      RECT  133.91 103.905 133.7 103.7 ;
      RECT  130.79 104.285 130.58 103.905 ;
      RECT  131.87 103.7 131.69 101.995 ;
      RECT  133.7 103.905 133.49 103.7 ;
      RECT  133.91 104.285 133.7 103.905 ;
      POLYGON  131.3 102.62 131.3 102.21 131.045 102.21 131.045 102.54 131.125 102.62 131.3 102.62 ;
      RECT  133.31 104.615 133.13 103.7 ;
      RECT  133.7 104.615 133.49 104.285 ;
      RECT  133.7 104.285 133.49 103.905 ;
      RECT  131.51 104.58 131.3 104.99 ;
      RECT  133.91 103.575 133.7 103.905 ;
      RECT  130.865 104.49 130.79 106.195 ;
      RECT  130.95 105.075 130.865 105.485 ;
      RECT  131.87 103.575 131.69 104.49 ;
      POLYGON  130.865 103.575 130.865 103.905 131.3 103.905 131.3 104.285 130.865 104.285 130.865 104.49 130.79 104.49 130.79 103.575 130.865 103.575 ;
      RECT  130.79 104.49 130.58 106.195 ;
      POLYGON  131.3 104.58 131.3 104.99 131.125 104.99 131.045 104.91 131.045 104.58 131.3 104.58 ;
      RECT  133.91 104.49 133.7 106.195 ;
      RECT  132.23 103.575 132.05 104.49 ;
      RECT  133.31 104.49 133.13 106.195 ;
      RECT  131.51 105.57 131.3 105.98 ;
      RECT  130.79 104.285 130.58 104.49 ;
      RECT  133.7 104.49 133.49 106.195 ;
      RECT  131.51 103.905 131.3 104.285 ;
      RECT  132.95 104.49 132.77 106.195 ;
      RECT  132.23 104.49 132.05 106.195 ;
      RECT  132.95 103.575 132.77 104.49 ;
      RECT  130.79 103.575 130.58 103.905 ;
      RECT  132.59 104.49 132.41 106.195 ;
      RECT  132.59 103.575 132.41 104.49 ;
      RECT  133.91 104.285 133.7 104.49 ;
      RECT  130.79 103.905 130.58 104.285 ;
      RECT  131.87 104.49 131.69 106.195 ;
      RECT  133.7 104.285 133.49 104.49 ;
      RECT  133.91 103.905 133.7 104.285 ;
      POLYGON  131.3 105.57 131.3 105.98 131.045 105.98 131.045 105.65 131.125 105.57 131.3 105.57 ;
      RECT  133.31 103.575 133.13 104.49 ;
      RECT  133.7 103.575 133.49 103.905 ;
      RECT  133.7 103.905 133.49 104.285 ;
      RECT  131.51 107.56 131.3 107.15 ;
      RECT  133.91 108.565 133.7 108.235 ;
      RECT  130.865 107.65 130.79 105.945 ;
      RECT  130.95 107.065 130.865 106.655 ;
      RECT  131.87 108.565 131.69 107.65 ;
      POLYGON  130.865 108.565 130.865 108.235 131.3 108.235 131.3 107.855 130.865 107.855 130.865 107.65 130.79 107.65 130.79 108.565 130.865 108.565 ;
      RECT  130.79 107.65 130.58 105.945 ;
      POLYGON  131.3 107.56 131.3 107.15 131.125 107.15 131.045 107.23 131.045 107.56 131.3 107.56 ;
      RECT  133.91 107.65 133.7 105.945 ;
      RECT  132.23 108.565 132.05 107.65 ;
      RECT  133.31 107.65 133.13 105.945 ;
      RECT  131.51 106.57 131.3 106.16 ;
      RECT  130.79 107.855 130.58 107.65 ;
      RECT  133.7 107.65 133.49 105.945 ;
      RECT  131.51 108.235 131.3 107.855 ;
      RECT  132.95 107.65 132.77 105.945 ;
      RECT  132.23 107.65 132.05 105.945 ;
      RECT  132.95 108.565 132.77 107.65 ;
      RECT  130.79 108.565 130.58 108.235 ;
      RECT  132.59 107.65 132.41 105.945 ;
      RECT  132.59 108.565 132.41 107.65 ;
      RECT  133.91 107.855 133.7 107.65 ;
      RECT  130.79 108.235 130.58 107.855 ;
      RECT  131.87 107.65 131.69 105.945 ;
      RECT  133.7 107.855 133.49 107.65 ;
      RECT  133.91 108.235 133.7 107.855 ;
      POLYGON  131.3 106.57 131.3 106.16 131.045 106.16 131.045 106.49 131.125 106.57 131.3 106.57 ;
      RECT  133.31 108.565 133.13 107.65 ;
      RECT  133.7 108.565 133.49 108.235 ;
      RECT  133.7 108.235 133.49 107.855 ;
      RECT  131.51 108.53 131.3 108.94 ;
      RECT  133.91 107.525 133.7 107.855 ;
      RECT  130.865 108.44 130.79 110.145 ;
      RECT  130.95 109.025 130.865 109.435 ;
      RECT  131.87 107.525 131.69 108.44 ;
      POLYGON  130.865 107.525 130.865 107.855 131.3 107.855 131.3 108.235 130.865 108.235 130.865 108.44 130.79 108.44 130.79 107.525 130.865 107.525 ;
      RECT  130.79 108.44 130.58 110.145 ;
      POLYGON  131.3 108.53 131.3 108.94 131.125 108.94 131.045 108.86 131.045 108.53 131.3 108.53 ;
      RECT  133.91 108.44 133.7 110.145 ;
      RECT  132.23 107.525 132.05 108.44 ;
      RECT  133.31 108.44 133.13 110.145 ;
      RECT  131.51 109.52 131.3 109.93 ;
      RECT  130.79 108.235 130.58 108.44 ;
      RECT  133.7 108.44 133.49 110.145 ;
      RECT  131.51 107.855 131.3 108.235 ;
      RECT  132.95 108.44 132.77 110.145 ;
      RECT  132.23 108.44 132.05 110.145 ;
      RECT  132.95 107.525 132.77 108.44 ;
      RECT  130.79 107.525 130.58 107.855 ;
      RECT  132.59 108.44 132.41 110.145 ;
      RECT  132.59 107.525 132.41 108.44 ;
      RECT  133.91 108.235 133.7 108.44 ;
      RECT  130.79 107.855 130.58 108.235 ;
      RECT  131.87 108.44 131.69 110.145 ;
      RECT  133.7 108.235 133.49 108.44 ;
      RECT  133.91 107.855 133.7 108.235 ;
      POLYGON  131.3 109.52 131.3 109.93 131.045 109.93 131.045 109.6 131.125 109.52 131.3 109.52 ;
      RECT  133.31 107.525 133.13 108.44 ;
      RECT  133.7 107.525 133.49 107.855 ;
      RECT  133.7 107.855 133.49 108.235 ;
      RECT  131.51 111.51 131.3 111.1 ;
      RECT  133.91 112.515 133.7 112.185 ;
      RECT  130.865 111.6 130.79 109.895 ;
      RECT  130.95 111.015 130.865 110.605 ;
      RECT  131.87 112.515 131.69 111.6 ;
      POLYGON  130.865 112.515 130.865 112.185 131.3 112.185 131.3 111.805 130.865 111.805 130.865 111.6 130.79 111.6 130.79 112.515 130.865 112.515 ;
      RECT  130.79 111.6 130.58 109.895 ;
      POLYGON  131.3 111.51 131.3 111.1 131.125 111.1 131.045 111.18 131.045 111.51 131.3 111.51 ;
      RECT  133.91 111.6 133.7 109.895 ;
      RECT  132.23 112.515 132.05 111.6 ;
      RECT  133.31 111.6 133.13 109.895 ;
      RECT  131.51 110.52 131.3 110.11 ;
      RECT  130.79 111.805 130.58 111.6 ;
      RECT  133.7 111.6 133.49 109.895 ;
      RECT  131.51 112.185 131.3 111.805 ;
      RECT  132.95 111.6 132.77 109.895 ;
      RECT  132.23 111.6 132.05 109.895 ;
      RECT  132.95 112.515 132.77 111.6 ;
      RECT  130.79 112.515 130.58 112.185 ;
      RECT  132.59 111.6 132.41 109.895 ;
      RECT  132.59 112.515 132.41 111.6 ;
      RECT  133.91 111.805 133.7 111.6 ;
      RECT  130.79 112.185 130.58 111.805 ;
      RECT  131.87 111.6 131.69 109.895 ;
      RECT  133.7 111.805 133.49 111.6 ;
      RECT  133.91 112.185 133.7 111.805 ;
      POLYGON  131.3 110.52 131.3 110.11 131.045 110.11 131.045 110.44 131.125 110.52 131.3 110.52 ;
      RECT  133.31 112.515 133.13 111.6 ;
      RECT  133.7 112.515 133.49 112.185 ;
      RECT  133.7 112.185 133.49 111.805 ;
      RECT  131.51 112.48 131.3 112.89 ;
      RECT  133.91 111.475 133.7 111.805 ;
      RECT  130.865 112.39 130.79 114.095 ;
      RECT  130.95 112.975 130.865 113.385 ;
      RECT  131.87 111.475 131.69 112.39 ;
      POLYGON  130.865 111.475 130.865 111.805 131.3 111.805 131.3 112.185 130.865 112.185 130.865 112.39 130.79 112.39 130.79 111.475 130.865 111.475 ;
      RECT  130.79 112.39 130.58 114.095 ;
      POLYGON  131.3 112.48 131.3 112.89 131.125 112.89 131.045 112.81 131.045 112.48 131.3 112.48 ;
      RECT  133.91 112.39 133.7 114.095 ;
      RECT  132.23 111.475 132.05 112.39 ;
      RECT  133.31 112.39 133.13 114.095 ;
      RECT  131.51 113.47 131.3 113.88 ;
      RECT  130.79 112.185 130.58 112.39 ;
      RECT  133.7 112.39 133.49 114.095 ;
      RECT  131.51 111.805 131.3 112.185 ;
      RECT  132.95 112.39 132.77 114.095 ;
      RECT  132.23 112.39 132.05 114.095 ;
      RECT  132.95 111.475 132.77 112.39 ;
      RECT  130.79 111.475 130.58 111.805 ;
      RECT  132.59 112.39 132.41 114.095 ;
      RECT  132.59 111.475 132.41 112.39 ;
      RECT  133.91 112.185 133.7 112.39 ;
      RECT  130.79 111.805 130.58 112.185 ;
      RECT  131.87 112.39 131.69 114.095 ;
      RECT  133.7 112.185 133.49 112.39 ;
      RECT  133.91 111.805 133.7 112.185 ;
      POLYGON  131.3 113.47 131.3 113.88 131.045 113.88 131.045 113.55 131.125 113.47 131.3 113.47 ;
      RECT  133.31 111.475 133.13 112.39 ;
      RECT  133.7 111.475 133.49 111.805 ;
      RECT  133.7 111.805 133.49 112.185 ;
      RECT  131.51 115.46 131.3 115.05 ;
      RECT  133.91 116.465 133.7 116.135 ;
      RECT  130.865 115.55 130.79 113.845 ;
      RECT  130.95 114.965 130.865 114.555 ;
      RECT  131.87 116.465 131.69 115.55 ;
      POLYGON  130.865 116.465 130.865 116.135 131.3 116.135 131.3 115.755 130.865 115.755 130.865 115.55 130.79 115.55 130.79 116.465 130.865 116.465 ;
      RECT  130.79 115.55 130.58 113.845 ;
      POLYGON  131.3 115.46 131.3 115.05 131.125 115.05 131.045 115.13 131.045 115.46 131.3 115.46 ;
      RECT  133.91 115.55 133.7 113.845 ;
      RECT  132.23 116.465 132.05 115.55 ;
      RECT  133.31 115.55 133.13 113.845 ;
      RECT  131.51 114.47 131.3 114.06 ;
      RECT  130.79 115.755 130.58 115.55 ;
      RECT  133.7 115.55 133.49 113.845 ;
      RECT  131.51 116.135 131.3 115.755 ;
      RECT  132.95 115.55 132.77 113.845 ;
      RECT  132.23 115.55 132.05 113.845 ;
      RECT  132.95 116.465 132.77 115.55 ;
      RECT  130.79 116.465 130.58 116.135 ;
      RECT  132.59 115.55 132.41 113.845 ;
      RECT  132.59 116.465 132.41 115.55 ;
      RECT  133.91 115.755 133.7 115.55 ;
      RECT  130.79 116.135 130.58 115.755 ;
      RECT  131.87 115.55 131.69 113.845 ;
      RECT  133.7 115.755 133.49 115.55 ;
      RECT  133.91 116.135 133.7 115.755 ;
      POLYGON  131.3 114.47 131.3 114.06 131.045 114.06 131.045 114.39 131.125 114.47 131.3 114.47 ;
      RECT  133.31 116.465 133.13 115.55 ;
      RECT  133.7 116.465 133.49 116.135 ;
      RECT  133.7 116.135 133.49 115.755 ;
      RECT  131.51 116.43 131.3 116.84 ;
      RECT  133.91 115.425 133.7 115.755 ;
      RECT  130.865 116.34 130.79 118.045 ;
      RECT  130.95 116.925 130.865 117.335 ;
      RECT  131.87 115.425 131.69 116.34 ;
      POLYGON  130.865 115.425 130.865 115.755 131.3 115.755 131.3 116.135 130.865 116.135 130.865 116.34 130.79 116.34 130.79 115.425 130.865 115.425 ;
      RECT  130.79 116.34 130.58 118.045 ;
      POLYGON  131.3 116.43 131.3 116.84 131.125 116.84 131.045 116.76 131.045 116.43 131.3 116.43 ;
      RECT  133.91 116.34 133.7 118.045 ;
      RECT  132.23 115.425 132.05 116.34 ;
      RECT  133.31 116.34 133.13 118.045 ;
      RECT  131.51 117.42 131.3 117.83 ;
      RECT  130.79 116.135 130.58 116.34 ;
      RECT  133.7 116.34 133.49 118.045 ;
      RECT  131.51 115.755 131.3 116.135 ;
      RECT  132.95 116.34 132.77 118.045 ;
      RECT  132.23 116.34 132.05 118.045 ;
      RECT  132.95 115.425 132.77 116.34 ;
      RECT  130.79 115.425 130.58 115.755 ;
      RECT  132.59 116.34 132.41 118.045 ;
      RECT  132.59 115.425 132.41 116.34 ;
      RECT  133.91 116.135 133.7 116.34 ;
      RECT  130.79 115.755 130.58 116.135 ;
      RECT  131.87 116.34 131.69 118.045 ;
      RECT  133.7 116.135 133.49 116.34 ;
      RECT  133.91 115.755 133.7 116.135 ;
      POLYGON  131.3 117.42 131.3 117.83 131.045 117.83 131.045 117.5 131.125 117.42 131.3 117.42 ;
      RECT  133.31 115.425 133.13 116.34 ;
      RECT  133.7 115.425 133.49 115.755 ;
      RECT  133.7 115.755 133.49 116.135 ;
      RECT  131.51 119.41 131.3 119.0 ;
      RECT  133.91 120.415 133.7 120.085 ;
      RECT  130.865 119.5 130.79 117.795 ;
      RECT  130.95 118.915 130.865 118.505 ;
      RECT  131.87 120.415 131.69 119.5 ;
      POLYGON  130.865 120.415 130.865 120.085 131.3 120.085 131.3 119.705 130.865 119.705 130.865 119.5 130.79 119.5 130.79 120.415 130.865 120.415 ;
      RECT  130.79 119.5 130.58 117.795 ;
      POLYGON  131.3 119.41 131.3 119.0 131.125 119.0 131.045 119.08 131.045 119.41 131.3 119.41 ;
      RECT  133.91 119.5 133.7 117.795 ;
      RECT  132.23 120.415 132.05 119.5 ;
      RECT  133.31 119.5 133.13 117.795 ;
      RECT  131.51 118.42 131.3 118.01 ;
      RECT  130.79 119.705 130.58 119.5 ;
      RECT  133.7 119.5 133.49 117.795 ;
      RECT  131.51 120.085 131.3 119.705 ;
      RECT  132.95 119.5 132.77 117.795 ;
      RECT  132.23 119.5 132.05 117.795 ;
      RECT  132.95 120.415 132.77 119.5 ;
      RECT  130.79 120.415 130.58 120.085 ;
      RECT  132.59 119.5 132.41 117.795 ;
      RECT  132.59 120.415 132.41 119.5 ;
      RECT  133.91 119.705 133.7 119.5 ;
      RECT  130.79 120.085 130.58 119.705 ;
      RECT  131.87 119.5 131.69 117.795 ;
      RECT  133.7 119.705 133.49 119.5 ;
      RECT  133.91 120.085 133.7 119.705 ;
      POLYGON  131.3 118.42 131.3 118.01 131.045 118.01 131.045 118.34 131.125 118.42 131.3 118.42 ;
      RECT  133.31 120.415 133.13 119.5 ;
      RECT  133.7 120.415 133.49 120.085 ;
      RECT  133.7 120.085 133.49 119.705 ;
      RECT  131.51 120.38 131.3 120.79 ;
      RECT  133.91 119.375 133.7 119.705 ;
      RECT  130.865 120.29 130.79 121.995 ;
      RECT  130.95 120.875 130.865 121.285 ;
      RECT  131.87 119.375 131.69 120.29 ;
      POLYGON  130.865 119.375 130.865 119.705 131.3 119.705 131.3 120.085 130.865 120.085 130.865 120.29 130.79 120.29 130.79 119.375 130.865 119.375 ;
      RECT  130.79 120.29 130.58 121.995 ;
      POLYGON  131.3 120.38 131.3 120.79 131.125 120.79 131.045 120.71 131.045 120.38 131.3 120.38 ;
      RECT  133.91 120.29 133.7 121.995 ;
      RECT  132.23 119.375 132.05 120.29 ;
      RECT  133.31 120.29 133.13 121.995 ;
      RECT  131.51 121.37 131.3 121.78 ;
      RECT  130.79 120.085 130.58 120.29 ;
      RECT  133.7 120.29 133.49 121.995 ;
      RECT  131.51 119.705 131.3 120.085 ;
      RECT  132.95 120.29 132.77 121.995 ;
      RECT  132.23 120.29 132.05 121.995 ;
      RECT  132.95 119.375 132.77 120.29 ;
      RECT  130.79 119.375 130.58 119.705 ;
      RECT  132.59 120.29 132.41 121.995 ;
      RECT  132.59 119.375 132.41 120.29 ;
      RECT  133.91 120.085 133.7 120.29 ;
      RECT  130.79 119.705 130.58 120.085 ;
      RECT  131.87 120.29 131.69 121.995 ;
      RECT  133.7 120.085 133.49 120.29 ;
      RECT  133.91 119.705 133.7 120.085 ;
      POLYGON  131.3 121.37 131.3 121.78 131.045 121.78 131.045 121.45 131.125 121.37 131.3 121.37 ;
      RECT  133.31 119.375 133.13 120.29 ;
      RECT  133.7 119.375 133.49 119.705 ;
      RECT  133.7 119.705 133.49 120.085 ;
      RECT  131.51 123.36 131.3 122.95 ;
      RECT  133.91 124.365 133.7 124.035 ;
      RECT  130.865 123.45 130.79 121.745 ;
      RECT  130.95 122.865 130.865 122.455 ;
      RECT  131.87 124.365 131.69 123.45 ;
      POLYGON  130.865 124.365 130.865 124.035 131.3 124.035 131.3 123.655 130.865 123.655 130.865 123.45 130.79 123.45 130.79 124.365 130.865 124.365 ;
      RECT  130.79 123.45 130.58 121.745 ;
      POLYGON  131.3 123.36 131.3 122.95 131.125 122.95 131.045 123.03 131.045 123.36 131.3 123.36 ;
      RECT  133.91 123.45 133.7 121.745 ;
      RECT  132.23 124.365 132.05 123.45 ;
      RECT  133.31 123.45 133.13 121.745 ;
      RECT  131.51 122.37 131.3 121.96 ;
      RECT  130.79 123.655 130.58 123.45 ;
      RECT  133.7 123.45 133.49 121.745 ;
      RECT  131.51 124.035 131.3 123.655 ;
      RECT  132.95 123.45 132.77 121.745 ;
      RECT  132.23 123.45 132.05 121.745 ;
      RECT  132.95 124.365 132.77 123.45 ;
      RECT  130.79 124.365 130.58 124.035 ;
      RECT  132.59 123.45 132.41 121.745 ;
      RECT  132.59 124.365 132.41 123.45 ;
      RECT  133.91 123.655 133.7 123.45 ;
      RECT  130.79 124.035 130.58 123.655 ;
      RECT  131.87 123.45 131.69 121.745 ;
      RECT  133.7 123.655 133.49 123.45 ;
      RECT  133.91 124.035 133.7 123.655 ;
      POLYGON  131.3 122.37 131.3 121.96 131.045 121.96 131.045 122.29 131.125 122.37 131.3 122.37 ;
      RECT  133.31 124.365 133.13 123.45 ;
      RECT  133.7 124.365 133.49 124.035 ;
      RECT  133.7 124.035 133.49 123.655 ;
      RECT  135.89 92.73 136.1 93.14 ;
      RECT  133.49 91.725 133.7 92.055 ;
      RECT  136.535 92.64 136.61 94.345 ;
      RECT  136.45 93.225 136.535 93.635 ;
      RECT  135.53 91.725 135.71 92.64 ;
      POLYGON  136.535 91.725 136.535 92.055 136.1 92.055 136.1 92.435 136.535 92.435 136.535 92.64 136.61 92.64 136.61 91.725 136.535 91.725 ;
      RECT  136.61 92.64 136.82 94.345 ;
      POLYGON  136.1 92.73 136.1 93.14 136.275 93.14 136.355 93.06 136.355 92.73 136.1 92.73 ;
      RECT  133.49 92.64 133.7 94.345 ;
      RECT  135.17 91.725 135.35 92.64 ;
      RECT  134.09 92.64 134.27 94.345 ;
      RECT  135.89 93.72 136.1 94.13 ;
      RECT  136.61 92.435 136.82 92.64 ;
      RECT  133.7 92.64 133.91 94.345 ;
      RECT  135.89 92.055 136.1 92.435 ;
      RECT  134.45 92.64 134.63 94.345 ;
      RECT  135.17 92.64 135.35 94.345 ;
      RECT  134.45 91.725 134.63 92.64 ;
      RECT  136.61 91.725 136.82 92.055 ;
      RECT  134.81 92.64 134.99 94.345 ;
      RECT  134.81 91.725 134.99 92.64 ;
      RECT  133.49 92.435 133.7 92.64 ;
      RECT  136.61 92.055 136.82 92.435 ;
      RECT  135.53 92.64 135.71 94.345 ;
      RECT  133.7 92.435 133.91 92.64 ;
      RECT  133.49 92.055 133.7 92.435 ;
      POLYGON  136.1 93.72 136.1 94.13 136.355 94.13 136.355 93.8 136.275 93.72 136.1 93.72 ;
      RECT  134.09 91.725 134.27 92.64 ;
      RECT  133.7 91.725 133.91 92.055 ;
      RECT  133.7 92.055 133.91 92.435 ;
      RECT  135.89 95.71 136.1 95.3 ;
      RECT  133.49 96.715 133.7 96.385 ;
      RECT  136.535 95.8 136.61 94.095 ;
      RECT  136.45 95.215 136.535 94.805 ;
      RECT  135.53 96.715 135.71 95.8 ;
      POLYGON  136.535 96.715 136.535 96.385 136.1 96.385 136.1 96.005 136.535 96.005 136.535 95.8 136.61 95.8 136.61 96.715 136.535 96.715 ;
      RECT  136.61 95.8 136.82 94.095 ;
      POLYGON  136.1 95.71 136.1 95.3 136.275 95.3 136.355 95.38 136.355 95.71 136.1 95.71 ;
      RECT  133.49 95.8 133.7 94.095 ;
      RECT  135.17 96.715 135.35 95.8 ;
      RECT  134.09 95.8 134.27 94.095 ;
      RECT  135.89 94.72 136.1 94.31 ;
      RECT  136.61 96.005 136.82 95.8 ;
      RECT  133.7 95.8 133.91 94.095 ;
      RECT  135.89 96.385 136.1 96.005 ;
      RECT  134.45 95.8 134.63 94.095 ;
      RECT  135.17 95.8 135.35 94.095 ;
      RECT  134.45 96.715 134.63 95.8 ;
      RECT  136.61 96.715 136.82 96.385 ;
      RECT  134.81 95.8 134.99 94.095 ;
      RECT  134.81 96.715 134.99 95.8 ;
      RECT  133.49 96.005 133.7 95.8 ;
      RECT  136.61 96.385 136.82 96.005 ;
      RECT  135.53 95.8 135.71 94.095 ;
      RECT  133.7 96.005 133.91 95.8 ;
      RECT  133.49 96.385 133.7 96.005 ;
      POLYGON  136.1 94.72 136.1 94.31 136.355 94.31 136.355 94.64 136.275 94.72 136.1 94.72 ;
      RECT  134.09 96.715 134.27 95.8 ;
      RECT  133.7 96.715 133.91 96.385 ;
      RECT  133.7 96.385 133.91 96.005 ;
      RECT  135.89 96.68 136.1 97.09 ;
      RECT  133.49 95.675 133.7 96.005 ;
      RECT  136.535 96.59 136.61 98.295 ;
      RECT  136.45 97.175 136.535 97.585 ;
      RECT  135.53 95.675 135.71 96.59 ;
      POLYGON  136.535 95.675 136.535 96.005 136.1 96.005 136.1 96.385 136.535 96.385 136.535 96.59 136.61 96.59 136.61 95.675 136.535 95.675 ;
      RECT  136.61 96.59 136.82 98.295 ;
      POLYGON  136.1 96.68 136.1 97.09 136.275 97.09 136.355 97.01 136.355 96.68 136.1 96.68 ;
      RECT  133.49 96.59 133.7 98.295 ;
      RECT  135.17 95.675 135.35 96.59 ;
      RECT  134.09 96.59 134.27 98.295 ;
      RECT  135.89 97.67 136.1 98.08 ;
      RECT  136.61 96.385 136.82 96.59 ;
      RECT  133.7 96.59 133.91 98.295 ;
      RECT  135.89 96.005 136.1 96.385 ;
      RECT  134.45 96.59 134.63 98.295 ;
      RECT  135.17 96.59 135.35 98.295 ;
      RECT  134.45 95.675 134.63 96.59 ;
      RECT  136.61 95.675 136.82 96.005 ;
      RECT  134.81 96.59 134.99 98.295 ;
      RECT  134.81 95.675 134.99 96.59 ;
      RECT  133.49 96.385 133.7 96.59 ;
      RECT  136.61 96.005 136.82 96.385 ;
      RECT  135.53 96.59 135.71 98.295 ;
      RECT  133.7 96.385 133.91 96.59 ;
      RECT  133.49 96.005 133.7 96.385 ;
      POLYGON  136.1 97.67 136.1 98.08 136.355 98.08 136.355 97.75 136.275 97.67 136.1 97.67 ;
      RECT  134.09 95.675 134.27 96.59 ;
      RECT  133.7 95.675 133.91 96.005 ;
      RECT  133.7 96.005 133.91 96.385 ;
      RECT  135.89 99.66 136.1 99.25 ;
      RECT  133.49 100.665 133.7 100.335 ;
      RECT  136.535 99.75 136.61 98.045 ;
      RECT  136.45 99.165 136.535 98.755 ;
      RECT  135.53 100.665 135.71 99.75 ;
      POLYGON  136.535 100.665 136.535 100.335 136.1 100.335 136.1 99.955 136.535 99.955 136.535 99.75 136.61 99.75 136.61 100.665 136.535 100.665 ;
      RECT  136.61 99.75 136.82 98.045 ;
      POLYGON  136.1 99.66 136.1 99.25 136.275 99.25 136.355 99.33 136.355 99.66 136.1 99.66 ;
      RECT  133.49 99.75 133.7 98.045 ;
      RECT  135.17 100.665 135.35 99.75 ;
      RECT  134.09 99.75 134.27 98.045 ;
      RECT  135.89 98.67 136.1 98.26 ;
      RECT  136.61 99.955 136.82 99.75 ;
      RECT  133.7 99.75 133.91 98.045 ;
      RECT  135.89 100.335 136.1 99.955 ;
      RECT  134.45 99.75 134.63 98.045 ;
      RECT  135.17 99.75 135.35 98.045 ;
      RECT  134.45 100.665 134.63 99.75 ;
      RECT  136.61 100.665 136.82 100.335 ;
      RECT  134.81 99.75 134.99 98.045 ;
      RECT  134.81 100.665 134.99 99.75 ;
      RECT  133.49 99.955 133.7 99.75 ;
      RECT  136.61 100.335 136.82 99.955 ;
      RECT  135.53 99.75 135.71 98.045 ;
      RECT  133.7 99.955 133.91 99.75 ;
      RECT  133.49 100.335 133.7 99.955 ;
      POLYGON  136.1 98.67 136.1 98.26 136.355 98.26 136.355 98.59 136.275 98.67 136.1 98.67 ;
      RECT  134.09 100.665 134.27 99.75 ;
      RECT  133.7 100.665 133.91 100.335 ;
      RECT  133.7 100.335 133.91 99.955 ;
      RECT  135.89 100.63 136.1 101.04 ;
      RECT  133.49 99.625 133.7 99.955 ;
      RECT  136.535 100.54 136.61 102.245 ;
      RECT  136.45 101.125 136.535 101.535 ;
      RECT  135.53 99.625 135.71 100.54 ;
      POLYGON  136.535 99.625 136.535 99.955 136.1 99.955 136.1 100.335 136.535 100.335 136.535 100.54 136.61 100.54 136.61 99.625 136.535 99.625 ;
      RECT  136.61 100.54 136.82 102.245 ;
      POLYGON  136.1 100.63 136.1 101.04 136.275 101.04 136.355 100.96 136.355 100.63 136.1 100.63 ;
      RECT  133.49 100.54 133.7 102.245 ;
      RECT  135.17 99.625 135.35 100.54 ;
      RECT  134.09 100.54 134.27 102.245 ;
      RECT  135.89 101.62 136.1 102.03 ;
      RECT  136.61 100.335 136.82 100.54 ;
      RECT  133.7 100.54 133.91 102.245 ;
      RECT  135.89 99.955 136.1 100.335 ;
      RECT  134.45 100.54 134.63 102.245 ;
      RECT  135.17 100.54 135.35 102.245 ;
      RECT  134.45 99.625 134.63 100.54 ;
      RECT  136.61 99.625 136.82 99.955 ;
      RECT  134.81 100.54 134.99 102.245 ;
      RECT  134.81 99.625 134.99 100.54 ;
      RECT  133.49 100.335 133.7 100.54 ;
      RECT  136.61 99.955 136.82 100.335 ;
      RECT  135.53 100.54 135.71 102.245 ;
      RECT  133.7 100.335 133.91 100.54 ;
      RECT  133.49 99.955 133.7 100.335 ;
      POLYGON  136.1 101.62 136.1 102.03 136.355 102.03 136.355 101.7 136.275 101.62 136.1 101.62 ;
      RECT  134.09 99.625 134.27 100.54 ;
      RECT  133.7 99.625 133.91 99.955 ;
      RECT  133.7 99.955 133.91 100.335 ;
      RECT  135.89 103.61 136.1 103.2 ;
      RECT  133.49 104.615 133.7 104.285 ;
      RECT  136.535 103.7 136.61 101.995 ;
      RECT  136.45 103.115 136.535 102.705 ;
      RECT  135.53 104.615 135.71 103.7 ;
      POLYGON  136.535 104.615 136.535 104.285 136.1 104.285 136.1 103.905 136.535 103.905 136.535 103.7 136.61 103.7 136.61 104.615 136.535 104.615 ;
      RECT  136.61 103.7 136.82 101.995 ;
      POLYGON  136.1 103.61 136.1 103.2 136.275 103.2 136.355 103.28 136.355 103.61 136.1 103.61 ;
      RECT  133.49 103.7 133.7 101.995 ;
      RECT  135.17 104.615 135.35 103.7 ;
      RECT  134.09 103.7 134.27 101.995 ;
      RECT  135.89 102.62 136.1 102.21 ;
      RECT  136.61 103.905 136.82 103.7 ;
      RECT  133.7 103.7 133.91 101.995 ;
      RECT  135.89 104.285 136.1 103.905 ;
      RECT  134.45 103.7 134.63 101.995 ;
      RECT  135.17 103.7 135.35 101.995 ;
      RECT  134.45 104.615 134.63 103.7 ;
      RECT  136.61 104.615 136.82 104.285 ;
      RECT  134.81 103.7 134.99 101.995 ;
      RECT  134.81 104.615 134.99 103.7 ;
      RECT  133.49 103.905 133.7 103.7 ;
      RECT  136.61 104.285 136.82 103.905 ;
      RECT  135.53 103.7 135.71 101.995 ;
      RECT  133.7 103.905 133.91 103.7 ;
      RECT  133.49 104.285 133.7 103.905 ;
      POLYGON  136.1 102.62 136.1 102.21 136.355 102.21 136.355 102.54 136.275 102.62 136.1 102.62 ;
      RECT  134.09 104.615 134.27 103.7 ;
      RECT  133.7 104.615 133.91 104.285 ;
      RECT  133.7 104.285 133.91 103.905 ;
      RECT  135.89 104.58 136.1 104.99 ;
      RECT  133.49 103.575 133.7 103.905 ;
      RECT  136.535 104.49 136.61 106.195 ;
      RECT  136.45 105.075 136.535 105.485 ;
      RECT  135.53 103.575 135.71 104.49 ;
      POLYGON  136.535 103.575 136.535 103.905 136.1 103.905 136.1 104.285 136.535 104.285 136.535 104.49 136.61 104.49 136.61 103.575 136.535 103.575 ;
      RECT  136.61 104.49 136.82 106.195 ;
      POLYGON  136.1 104.58 136.1 104.99 136.275 104.99 136.355 104.91 136.355 104.58 136.1 104.58 ;
      RECT  133.49 104.49 133.7 106.195 ;
      RECT  135.17 103.575 135.35 104.49 ;
      RECT  134.09 104.49 134.27 106.195 ;
      RECT  135.89 105.57 136.1 105.98 ;
      RECT  136.61 104.285 136.82 104.49 ;
      RECT  133.7 104.49 133.91 106.195 ;
      RECT  135.89 103.905 136.1 104.285 ;
      RECT  134.45 104.49 134.63 106.195 ;
      RECT  135.17 104.49 135.35 106.195 ;
      RECT  134.45 103.575 134.63 104.49 ;
      RECT  136.61 103.575 136.82 103.905 ;
      RECT  134.81 104.49 134.99 106.195 ;
      RECT  134.81 103.575 134.99 104.49 ;
      RECT  133.49 104.285 133.7 104.49 ;
      RECT  136.61 103.905 136.82 104.285 ;
      RECT  135.53 104.49 135.71 106.195 ;
      RECT  133.7 104.285 133.91 104.49 ;
      RECT  133.49 103.905 133.7 104.285 ;
      POLYGON  136.1 105.57 136.1 105.98 136.355 105.98 136.355 105.65 136.275 105.57 136.1 105.57 ;
      RECT  134.09 103.575 134.27 104.49 ;
      RECT  133.7 103.575 133.91 103.905 ;
      RECT  133.7 103.905 133.91 104.285 ;
      RECT  135.89 107.56 136.1 107.15 ;
      RECT  133.49 108.565 133.7 108.235 ;
      RECT  136.535 107.65 136.61 105.945 ;
      RECT  136.45 107.065 136.535 106.655 ;
      RECT  135.53 108.565 135.71 107.65 ;
      POLYGON  136.535 108.565 136.535 108.235 136.1 108.235 136.1 107.855 136.535 107.855 136.535 107.65 136.61 107.65 136.61 108.565 136.535 108.565 ;
      RECT  136.61 107.65 136.82 105.945 ;
      POLYGON  136.1 107.56 136.1 107.15 136.275 107.15 136.355 107.23 136.355 107.56 136.1 107.56 ;
      RECT  133.49 107.65 133.7 105.945 ;
      RECT  135.17 108.565 135.35 107.65 ;
      RECT  134.09 107.65 134.27 105.945 ;
      RECT  135.89 106.57 136.1 106.16 ;
      RECT  136.61 107.855 136.82 107.65 ;
      RECT  133.7 107.65 133.91 105.945 ;
      RECT  135.89 108.235 136.1 107.855 ;
      RECT  134.45 107.65 134.63 105.945 ;
      RECT  135.17 107.65 135.35 105.945 ;
      RECT  134.45 108.565 134.63 107.65 ;
      RECT  136.61 108.565 136.82 108.235 ;
      RECT  134.81 107.65 134.99 105.945 ;
      RECT  134.81 108.565 134.99 107.65 ;
      RECT  133.49 107.855 133.7 107.65 ;
      RECT  136.61 108.235 136.82 107.855 ;
      RECT  135.53 107.65 135.71 105.945 ;
      RECT  133.7 107.855 133.91 107.65 ;
      RECT  133.49 108.235 133.7 107.855 ;
      POLYGON  136.1 106.57 136.1 106.16 136.355 106.16 136.355 106.49 136.275 106.57 136.1 106.57 ;
      RECT  134.09 108.565 134.27 107.65 ;
      RECT  133.7 108.565 133.91 108.235 ;
      RECT  133.7 108.235 133.91 107.855 ;
      RECT  135.89 108.53 136.1 108.94 ;
      RECT  133.49 107.525 133.7 107.855 ;
      RECT  136.535 108.44 136.61 110.145 ;
      RECT  136.45 109.025 136.535 109.435 ;
      RECT  135.53 107.525 135.71 108.44 ;
      POLYGON  136.535 107.525 136.535 107.855 136.1 107.855 136.1 108.235 136.535 108.235 136.535 108.44 136.61 108.44 136.61 107.525 136.535 107.525 ;
      RECT  136.61 108.44 136.82 110.145 ;
      POLYGON  136.1 108.53 136.1 108.94 136.275 108.94 136.355 108.86 136.355 108.53 136.1 108.53 ;
      RECT  133.49 108.44 133.7 110.145 ;
      RECT  135.17 107.525 135.35 108.44 ;
      RECT  134.09 108.44 134.27 110.145 ;
      RECT  135.89 109.52 136.1 109.93 ;
      RECT  136.61 108.235 136.82 108.44 ;
      RECT  133.7 108.44 133.91 110.145 ;
      RECT  135.89 107.855 136.1 108.235 ;
      RECT  134.45 108.44 134.63 110.145 ;
      RECT  135.17 108.44 135.35 110.145 ;
      RECT  134.45 107.525 134.63 108.44 ;
      RECT  136.61 107.525 136.82 107.855 ;
      RECT  134.81 108.44 134.99 110.145 ;
      RECT  134.81 107.525 134.99 108.44 ;
      RECT  133.49 108.235 133.7 108.44 ;
      RECT  136.61 107.855 136.82 108.235 ;
      RECT  135.53 108.44 135.71 110.145 ;
      RECT  133.7 108.235 133.91 108.44 ;
      RECT  133.49 107.855 133.7 108.235 ;
      POLYGON  136.1 109.52 136.1 109.93 136.355 109.93 136.355 109.6 136.275 109.52 136.1 109.52 ;
      RECT  134.09 107.525 134.27 108.44 ;
      RECT  133.7 107.525 133.91 107.855 ;
      RECT  133.7 107.855 133.91 108.235 ;
      RECT  135.89 111.51 136.1 111.1 ;
      RECT  133.49 112.515 133.7 112.185 ;
      RECT  136.535 111.6 136.61 109.895 ;
      RECT  136.45 111.015 136.535 110.605 ;
      RECT  135.53 112.515 135.71 111.6 ;
      POLYGON  136.535 112.515 136.535 112.185 136.1 112.185 136.1 111.805 136.535 111.805 136.535 111.6 136.61 111.6 136.61 112.515 136.535 112.515 ;
      RECT  136.61 111.6 136.82 109.895 ;
      POLYGON  136.1 111.51 136.1 111.1 136.275 111.1 136.355 111.18 136.355 111.51 136.1 111.51 ;
      RECT  133.49 111.6 133.7 109.895 ;
      RECT  135.17 112.515 135.35 111.6 ;
      RECT  134.09 111.6 134.27 109.895 ;
      RECT  135.89 110.52 136.1 110.11 ;
      RECT  136.61 111.805 136.82 111.6 ;
      RECT  133.7 111.6 133.91 109.895 ;
      RECT  135.89 112.185 136.1 111.805 ;
      RECT  134.45 111.6 134.63 109.895 ;
      RECT  135.17 111.6 135.35 109.895 ;
      RECT  134.45 112.515 134.63 111.6 ;
      RECT  136.61 112.515 136.82 112.185 ;
      RECT  134.81 111.6 134.99 109.895 ;
      RECT  134.81 112.515 134.99 111.6 ;
      RECT  133.49 111.805 133.7 111.6 ;
      RECT  136.61 112.185 136.82 111.805 ;
      RECT  135.53 111.6 135.71 109.895 ;
      RECT  133.7 111.805 133.91 111.6 ;
      RECT  133.49 112.185 133.7 111.805 ;
      POLYGON  136.1 110.52 136.1 110.11 136.355 110.11 136.355 110.44 136.275 110.52 136.1 110.52 ;
      RECT  134.09 112.515 134.27 111.6 ;
      RECT  133.7 112.515 133.91 112.185 ;
      RECT  133.7 112.185 133.91 111.805 ;
      RECT  135.89 112.48 136.1 112.89 ;
      RECT  133.49 111.475 133.7 111.805 ;
      RECT  136.535 112.39 136.61 114.095 ;
      RECT  136.45 112.975 136.535 113.385 ;
      RECT  135.53 111.475 135.71 112.39 ;
      POLYGON  136.535 111.475 136.535 111.805 136.1 111.805 136.1 112.185 136.535 112.185 136.535 112.39 136.61 112.39 136.61 111.475 136.535 111.475 ;
      RECT  136.61 112.39 136.82 114.095 ;
      POLYGON  136.1 112.48 136.1 112.89 136.275 112.89 136.355 112.81 136.355 112.48 136.1 112.48 ;
      RECT  133.49 112.39 133.7 114.095 ;
      RECT  135.17 111.475 135.35 112.39 ;
      RECT  134.09 112.39 134.27 114.095 ;
      RECT  135.89 113.47 136.1 113.88 ;
      RECT  136.61 112.185 136.82 112.39 ;
      RECT  133.7 112.39 133.91 114.095 ;
      RECT  135.89 111.805 136.1 112.185 ;
      RECT  134.45 112.39 134.63 114.095 ;
      RECT  135.17 112.39 135.35 114.095 ;
      RECT  134.45 111.475 134.63 112.39 ;
      RECT  136.61 111.475 136.82 111.805 ;
      RECT  134.81 112.39 134.99 114.095 ;
      RECT  134.81 111.475 134.99 112.39 ;
      RECT  133.49 112.185 133.7 112.39 ;
      RECT  136.61 111.805 136.82 112.185 ;
      RECT  135.53 112.39 135.71 114.095 ;
      RECT  133.7 112.185 133.91 112.39 ;
      RECT  133.49 111.805 133.7 112.185 ;
      POLYGON  136.1 113.47 136.1 113.88 136.355 113.88 136.355 113.55 136.275 113.47 136.1 113.47 ;
      RECT  134.09 111.475 134.27 112.39 ;
      RECT  133.7 111.475 133.91 111.805 ;
      RECT  133.7 111.805 133.91 112.185 ;
      RECT  135.89 115.46 136.1 115.05 ;
      RECT  133.49 116.465 133.7 116.135 ;
      RECT  136.535 115.55 136.61 113.845 ;
      RECT  136.45 114.965 136.535 114.555 ;
      RECT  135.53 116.465 135.71 115.55 ;
      POLYGON  136.535 116.465 136.535 116.135 136.1 116.135 136.1 115.755 136.535 115.755 136.535 115.55 136.61 115.55 136.61 116.465 136.535 116.465 ;
      RECT  136.61 115.55 136.82 113.845 ;
      POLYGON  136.1 115.46 136.1 115.05 136.275 115.05 136.355 115.13 136.355 115.46 136.1 115.46 ;
      RECT  133.49 115.55 133.7 113.845 ;
      RECT  135.17 116.465 135.35 115.55 ;
      RECT  134.09 115.55 134.27 113.845 ;
      RECT  135.89 114.47 136.1 114.06 ;
      RECT  136.61 115.755 136.82 115.55 ;
      RECT  133.7 115.55 133.91 113.845 ;
      RECT  135.89 116.135 136.1 115.755 ;
      RECT  134.45 115.55 134.63 113.845 ;
      RECT  135.17 115.55 135.35 113.845 ;
      RECT  134.45 116.465 134.63 115.55 ;
      RECT  136.61 116.465 136.82 116.135 ;
      RECT  134.81 115.55 134.99 113.845 ;
      RECT  134.81 116.465 134.99 115.55 ;
      RECT  133.49 115.755 133.7 115.55 ;
      RECT  136.61 116.135 136.82 115.755 ;
      RECT  135.53 115.55 135.71 113.845 ;
      RECT  133.7 115.755 133.91 115.55 ;
      RECT  133.49 116.135 133.7 115.755 ;
      POLYGON  136.1 114.47 136.1 114.06 136.355 114.06 136.355 114.39 136.275 114.47 136.1 114.47 ;
      RECT  134.09 116.465 134.27 115.55 ;
      RECT  133.7 116.465 133.91 116.135 ;
      RECT  133.7 116.135 133.91 115.755 ;
      RECT  135.89 116.43 136.1 116.84 ;
      RECT  133.49 115.425 133.7 115.755 ;
      RECT  136.535 116.34 136.61 118.045 ;
      RECT  136.45 116.925 136.535 117.335 ;
      RECT  135.53 115.425 135.71 116.34 ;
      POLYGON  136.535 115.425 136.535 115.755 136.1 115.755 136.1 116.135 136.535 116.135 136.535 116.34 136.61 116.34 136.61 115.425 136.535 115.425 ;
      RECT  136.61 116.34 136.82 118.045 ;
      POLYGON  136.1 116.43 136.1 116.84 136.275 116.84 136.355 116.76 136.355 116.43 136.1 116.43 ;
      RECT  133.49 116.34 133.7 118.045 ;
      RECT  135.17 115.425 135.35 116.34 ;
      RECT  134.09 116.34 134.27 118.045 ;
      RECT  135.89 117.42 136.1 117.83 ;
      RECT  136.61 116.135 136.82 116.34 ;
      RECT  133.7 116.34 133.91 118.045 ;
      RECT  135.89 115.755 136.1 116.135 ;
      RECT  134.45 116.34 134.63 118.045 ;
      RECT  135.17 116.34 135.35 118.045 ;
      RECT  134.45 115.425 134.63 116.34 ;
      RECT  136.61 115.425 136.82 115.755 ;
      RECT  134.81 116.34 134.99 118.045 ;
      RECT  134.81 115.425 134.99 116.34 ;
      RECT  133.49 116.135 133.7 116.34 ;
      RECT  136.61 115.755 136.82 116.135 ;
      RECT  135.53 116.34 135.71 118.045 ;
      RECT  133.7 116.135 133.91 116.34 ;
      RECT  133.49 115.755 133.7 116.135 ;
      POLYGON  136.1 117.42 136.1 117.83 136.355 117.83 136.355 117.5 136.275 117.42 136.1 117.42 ;
      RECT  134.09 115.425 134.27 116.34 ;
      RECT  133.7 115.425 133.91 115.755 ;
      RECT  133.7 115.755 133.91 116.135 ;
      RECT  135.89 119.41 136.1 119.0 ;
      RECT  133.49 120.415 133.7 120.085 ;
      RECT  136.535 119.5 136.61 117.795 ;
      RECT  136.45 118.915 136.535 118.505 ;
      RECT  135.53 120.415 135.71 119.5 ;
      POLYGON  136.535 120.415 136.535 120.085 136.1 120.085 136.1 119.705 136.535 119.705 136.535 119.5 136.61 119.5 136.61 120.415 136.535 120.415 ;
      RECT  136.61 119.5 136.82 117.795 ;
      POLYGON  136.1 119.41 136.1 119.0 136.275 119.0 136.355 119.08 136.355 119.41 136.1 119.41 ;
      RECT  133.49 119.5 133.7 117.795 ;
      RECT  135.17 120.415 135.35 119.5 ;
      RECT  134.09 119.5 134.27 117.795 ;
      RECT  135.89 118.42 136.1 118.01 ;
      RECT  136.61 119.705 136.82 119.5 ;
      RECT  133.7 119.5 133.91 117.795 ;
      RECT  135.89 120.085 136.1 119.705 ;
      RECT  134.45 119.5 134.63 117.795 ;
      RECT  135.17 119.5 135.35 117.795 ;
      RECT  134.45 120.415 134.63 119.5 ;
      RECT  136.61 120.415 136.82 120.085 ;
      RECT  134.81 119.5 134.99 117.795 ;
      RECT  134.81 120.415 134.99 119.5 ;
      RECT  133.49 119.705 133.7 119.5 ;
      RECT  136.61 120.085 136.82 119.705 ;
      RECT  135.53 119.5 135.71 117.795 ;
      RECT  133.7 119.705 133.91 119.5 ;
      RECT  133.49 120.085 133.7 119.705 ;
      POLYGON  136.1 118.42 136.1 118.01 136.355 118.01 136.355 118.34 136.275 118.42 136.1 118.42 ;
      RECT  134.09 120.415 134.27 119.5 ;
      RECT  133.7 120.415 133.91 120.085 ;
      RECT  133.7 120.085 133.91 119.705 ;
      RECT  135.89 120.38 136.1 120.79 ;
      RECT  133.49 119.375 133.7 119.705 ;
      RECT  136.535 120.29 136.61 121.995 ;
      RECT  136.45 120.875 136.535 121.285 ;
      RECT  135.53 119.375 135.71 120.29 ;
      POLYGON  136.535 119.375 136.535 119.705 136.1 119.705 136.1 120.085 136.535 120.085 136.535 120.29 136.61 120.29 136.61 119.375 136.535 119.375 ;
      RECT  136.61 120.29 136.82 121.995 ;
      POLYGON  136.1 120.38 136.1 120.79 136.275 120.79 136.355 120.71 136.355 120.38 136.1 120.38 ;
      RECT  133.49 120.29 133.7 121.995 ;
      RECT  135.17 119.375 135.35 120.29 ;
      RECT  134.09 120.29 134.27 121.995 ;
      RECT  135.89 121.37 136.1 121.78 ;
      RECT  136.61 120.085 136.82 120.29 ;
      RECT  133.7 120.29 133.91 121.995 ;
      RECT  135.89 119.705 136.1 120.085 ;
      RECT  134.45 120.29 134.63 121.995 ;
      RECT  135.17 120.29 135.35 121.995 ;
      RECT  134.45 119.375 134.63 120.29 ;
      RECT  136.61 119.375 136.82 119.705 ;
      RECT  134.81 120.29 134.99 121.995 ;
      RECT  134.81 119.375 134.99 120.29 ;
      RECT  133.49 120.085 133.7 120.29 ;
      RECT  136.61 119.705 136.82 120.085 ;
      RECT  135.53 120.29 135.71 121.995 ;
      RECT  133.7 120.085 133.91 120.29 ;
      RECT  133.49 119.705 133.7 120.085 ;
      POLYGON  136.1 121.37 136.1 121.78 136.355 121.78 136.355 121.45 136.275 121.37 136.1 121.37 ;
      RECT  134.09 119.375 134.27 120.29 ;
      RECT  133.7 119.375 133.91 119.705 ;
      RECT  133.7 119.705 133.91 120.085 ;
      RECT  135.89 123.36 136.1 122.95 ;
      RECT  133.49 124.365 133.7 124.035 ;
      RECT  136.535 123.45 136.61 121.745 ;
      RECT  136.45 122.865 136.535 122.455 ;
      RECT  135.53 124.365 135.71 123.45 ;
      POLYGON  136.535 124.365 136.535 124.035 136.1 124.035 136.1 123.655 136.535 123.655 136.535 123.45 136.61 123.45 136.61 124.365 136.535 124.365 ;
      RECT  136.61 123.45 136.82 121.745 ;
      POLYGON  136.1 123.36 136.1 122.95 136.275 122.95 136.355 123.03 136.355 123.36 136.1 123.36 ;
      RECT  133.49 123.45 133.7 121.745 ;
      RECT  135.17 124.365 135.35 123.45 ;
      RECT  134.09 123.45 134.27 121.745 ;
      RECT  135.89 122.37 136.1 121.96 ;
      RECT  136.61 123.655 136.82 123.45 ;
      RECT  133.7 123.45 133.91 121.745 ;
      RECT  135.89 124.035 136.1 123.655 ;
      RECT  134.45 123.45 134.63 121.745 ;
      RECT  135.17 123.45 135.35 121.745 ;
      RECT  134.45 124.365 134.63 123.45 ;
      RECT  136.61 124.365 136.82 124.035 ;
      RECT  134.81 123.45 134.99 121.745 ;
      RECT  134.81 124.365 134.99 123.45 ;
      RECT  133.49 123.655 133.7 123.45 ;
      RECT  136.61 124.035 136.82 123.655 ;
      RECT  135.53 123.45 135.71 121.745 ;
      RECT  133.7 123.655 133.91 123.45 ;
      RECT  133.49 124.035 133.7 123.655 ;
      POLYGON  136.1 122.37 136.1 121.96 136.355 121.96 136.355 122.29 136.275 122.37 136.1 122.37 ;
      RECT  134.09 124.365 134.27 123.45 ;
      RECT  133.7 124.365 133.91 124.035 ;
      RECT  133.7 124.035 133.91 123.655 ;
      RECT  137.75 92.73 137.54 93.14 ;
      RECT  140.15 91.725 139.94 92.055 ;
      RECT  137.105 92.64 137.03 94.345 ;
      RECT  137.19 93.225 137.105 93.635 ;
      RECT  138.11 91.725 137.93 92.64 ;
      POLYGON  137.105 91.725 137.105 92.055 137.54 92.055 137.54 92.435 137.105 92.435 137.105 92.64 137.03 92.64 137.03 91.725 137.105 91.725 ;
      RECT  137.03 92.64 136.82 94.345 ;
      POLYGON  137.54 92.73 137.54 93.14 137.365 93.14 137.285 93.06 137.285 92.73 137.54 92.73 ;
      RECT  140.15 92.64 139.94 94.345 ;
      RECT  138.47 91.725 138.29 92.64 ;
      RECT  139.55 92.64 139.37 94.345 ;
      RECT  137.75 93.72 137.54 94.13 ;
      RECT  137.03 92.435 136.82 92.64 ;
      RECT  139.94 92.64 139.73 94.345 ;
      RECT  137.75 92.055 137.54 92.435 ;
      RECT  139.19 92.64 139.01 94.345 ;
      RECT  138.47 92.64 138.29 94.345 ;
      RECT  139.19 91.725 139.01 92.64 ;
      RECT  137.03 91.725 136.82 92.055 ;
      RECT  138.83 92.64 138.65 94.345 ;
      RECT  138.83 91.725 138.65 92.64 ;
      RECT  140.15 92.435 139.94 92.64 ;
      RECT  137.03 92.055 136.82 92.435 ;
      RECT  138.11 92.64 137.93 94.345 ;
      RECT  139.94 92.435 139.73 92.64 ;
      RECT  140.15 92.055 139.94 92.435 ;
      POLYGON  137.54 93.72 137.54 94.13 137.285 94.13 137.285 93.8 137.365 93.72 137.54 93.72 ;
      RECT  139.55 91.725 139.37 92.64 ;
      RECT  139.94 91.725 139.73 92.055 ;
      RECT  139.94 92.055 139.73 92.435 ;
      RECT  137.75 95.71 137.54 95.3 ;
      RECT  140.15 96.715 139.94 96.385 ;
      RECT  137.105 95.8 137.03 94.095 ;
      RECT  137.19 95.215 137.105 94.805 ;
      RECT  138.11 96.715 137.93 95.8 ;
      POLYGON  137.105 96.715 137.105 96.385 137.54 96.385 137.54 96.005 137.105 96.005 137.105 95.8 137.03 95.8 137.03 96.715 137.105 96.715 ;
      RECT  137.03 95.8 136.82 94.095 ;
      POLYGON  137.54 95.71 137.54 95.3 137.365 95.3 137.285 95.38 137.285 95.71 137.54 95.71 ;
      RECT  140.15 95.8 139.94 94.095 ;
      RECT  138.47 96.715 138.29 95.8 ;
      RECT  139.55 95.8 139.37 94.095 ;
      RECT  137.75 94.72 137.54 94.31 ;
      RECT  137.03 96.005 136.82 95.8 ;
      RECT  139.94 95.8 139.73 94.095 ;
      RECT  137.75 96.385 137.54 96.005 ;
      RECT  139.19 95.8 139.01 94.095 ;
      RECT  138.47 95.8 138.29 94.095 ;
      RECT  139.19 96.715 139.01 95.8 ;
      RECT  137.03 96.715 136.82 96.385 ;
      RECT  138.83 95.8 138.65 94.095 ;
      RECT  138.83 96.715 138.65 95.8 ;
      RECT  140.15 96.005 139.94 95.8 ;
      RECT  137.03 96.385 136.82 96.005 ;
      RECT  138.11 95.8 137.93 94.095 ;
      RECT  139.94 96.005 139.73 95.8 ;
      RECT  140.15 96.385 139.94 96.005 ;
      POLYGON  137.54 94.72 137.54 94.31 137.285 94.31 137.285 94.64 137.365 94.72 137.54 94.72 ;
      RECT  139.55 96.715 139.37 95.8 ;
      RECT  139.94 96.715 139.73 96.385 ;
      RECT  139.94 96.385 139.73 96.005 ;
      RECT  137.75 96.68 137.54 97.09 ;
      RECT  140.15 95.675 139.94 96.005 ;
      RECT  137.105 96.59 137.03 98.295 ;
      RECT  137.19 97.175 137.105 97.585 ;
      RECT  138.11 95.675 137.93 96.59 ;
      POLYGON  137.105 95.675 137.105 96.005 137.54 96.005 137.54 96.385 137.105 96.385 137.105 96.59 137.03 96.59 137.03 95.675 137.105 95.675 ;
      RECT  137.03 96.59 136.82 98.295 ;
      POLYGON  137.54 96.68 137.54 97.09 137.365 97.09 137.285 97.01 137.285 96.68 137.54 96.68 ;
      RECT  140.15 96.59 139.94 98.295 ;
      RECT  138.47 95.675 138.29 96.59 ;
      RECT  139.55 96.59 139.37 98.295 ;
      RECT  137.75 97.67 137.54 98.08 ;
      RECT  137.03 96.385 136.82 96.59 ;
      RECT  139.94 96.59 139.73 98.295 ;
      RECT  137.75 96.005 137.54 96.385 ;
      RECT  139.19 96.59 139.01 98.295 ;
      RECT  138.47 96.59 138.29 98.295 ;
      RECT  139.19 95.675 139.01 96.59 ;
      RECT  137.03 95.675 136.82 96.005 ;
      RECT  138.83 96.59 138.65 98.295 ;
      RECT  138.83 95.675 138.65 96.59 ;
      RECT  140.15 96.385 139.94 96.59 ;
      RECT  137.03 96.005 136.82 96.385 ;
      RECT  138.11 96.59 137.93 98.295 ;
      RECT  139.94 96.385 139.73 96.59 ;
      RECT  140.15 96.005 139.94 96.385 ;
      POLYGON  137.54 97.67 137.54 98.08 137.285 98.08 137.285 97.75 137.365 97.67 137.54 97.67 ;
      RECT  139.55 95.675 139.37 96.59 ;
      RECT  139.94 95.675 139.73 96.005 ;
      RECT  139.94 96.005 139.73 96.385 ;
      RECT  137.75 99.66 137.54 99.25 ;
      RECT  140.15 100.665 139.94 100.335 ;
      RECT  137.105 99.75 137.03 98.045 ;
      RECT  137.19 99.165 137.105 98.755 ;
      RECT  138.11 100.665 137.93 99.75 ;
      POLYGON  137.105 100.665 137.105 100.335 137.54 100.335 137.54 99.955 137.105 99.955 137.105 99.75 137.03 99.75 137.03 100.665 137.105 100.665 ;
      RECT  137.03 99.75 136.82 98.045 ;
      POLYGON  137.54 99.66 137.54 99.25 137.365 99.25 137.285 99.33 137.285 99.66 137.54 99.66 ;
      RECT  140.15 99.75 139.94 98.045 ;
      RECT  138.47 100.665 138.29 99.75 ;
      RECT  139.55 99.75 139.37 98.045 ;
      RECT  137.75 98.67 137.54 98.26 ;
      RECT  137.03 99.955 136.82 99.75 ;
      RECT  139.94 99.75 139.73 98.045 ;
      RECT  137.75 100.335 137.54 99.955 ;
      RECT  139.19 99.75 139.01 98.045 ;
      RECT  138.47 99.75 138.29 98.045 ;
      RECT  139.19 100.665 139.01 99.75 ;
      RECT  137.03 100.665 136.82 100.335 ;
      RECT  138.83 99.75 138.65 98.045 ;
      RECT  138.83 100.665 138.65 99.75 ;
      RECT  140.15 99.955 139.94 99.75 ;
      RECT  137.03 100.335 136.82 99.955 ;
      RECT  138.11 99.75 137.93 98.045 ;
      RECT  139.94 99.955 139.73 99.75 ;
      RECT  140.15 100.335 139.94 99.955 ;
      POLYGON  137.54 98.67 137.54 98.26 137.285 98.26 137.285 98.59 137.365 98.67 137.54 98.67 ;
      RECT  139.55 100.665 139.37 99.75 ;
      RECT  139.94 100.665 139.73 100.335 ;
      RECT  139.94 100.335 139.73 99.955 ;
      RECT  137.75 100.63 137.54 101.04 ;
      RECT  140.15 99.625 139.94 99.955 ;
      RECT  137.105 100.54 137.03 102.245 ;
      RECT  137.19 101.125 137.105 101.535 ;
      RECT  138.11 99.625 137.93 100.54 ;
      POLYGON  137.105 99.625 137.105 99.955 137.54 99.955 137.54 100.335 137.105 100.335 137.105 100.54 137.03 100.54 137.03 99.625 137.105 99.625 ;
      RECT  137.03 100.54 136.82 102.245 ;
      POLYGON  137.54 100.63 137.54 101.04 137.365 101.04 137.285 100.96 137.285 100.63 137.54 100.63 ;
      RECT  140.15 100.54 139.94 102.245 ;
      RECT  138.47 99.625 138.29 100.54 ;
      RECT  139.55 100.54 139.37 102.245 ;
      RECT  137.75 101.62 137.54 102.03 ;
      RECT  137.03 100.335 136.82 100.54 ;
      RECT  139.94 100.54 139.73 102.245 ;
      RECT  137.75 99.955 137.54 100.335 ;
      RECT  139.19 100.54 139.01 102.245 ;
      RECT  138.47 100.54 138.29 102.245 ;
      RECT  139.19 99.625 139.01 100.54 ;
      RECT  137.03 99.625 136.82 99.955 ;
      RECT  138.83 100.54 138.65 102.245 ;
      RECT  138.83 99.625 138.65 100.54 ;
      RECT  140.15 100.335 139.94 100.54 ;
      RECT  137.03 99.955 136.82 100.335 ;
      RECT  138.11 100.54 137.93 102.245 ;
      RECT  139.94 100.335 139.73 100.54 ;
      RECT  140.15 99.955 139.94 100.335 ;
      POLYGON  137.54 101.62 137.54 102.03 137.285 102.03 137.285 101.7 137.365 101.62 137.54 101.62 ;
      RECT  139.55 99.625 139.37 100.54 ;
      RECT  139.94 99.625 139.73 99.955 ;
      RECT  139.94 99.955 139.73 100.335 ;
      RECT  137.75 103.61 137.54 103.2 ;
      RECT  140.15 104.615 139.94 104.285 ;
      RECT  137.105 103.7 137.03 101.995 ;
      RECT  137.19 103.115 137.105 102.705 ;
      RECT  138.11 104.615 137.93 103.7 ;
      POLYGON  137.105 104.615 137.105 104.285 137.54 104.285 137.54 103.905 137.105 103.905 137.105 103.7 137.03 103.7 137.03 104.615 137.105 104.615 ;
      RECT  137.03 103.7 136.82 101.995 ;
      POLYGON  137.54 103.61 137.54 103.2 137.365 103.2 137.285 103.28 137.285 103.61 137.54 103.61 ;
      RECT  140.15 103.7 139.94 101.995 ;
      RECT  138.47 104.615 138.29 103.7 ;
      RECT  139.55 103.7 139.37 101.995 ;
      RECT  137.75 102.62 137.54 102.21 ;
      RECT  137.03 103.905 136.82 103.7 ;
      RECT  139.94 103.7 139.73 101.995 ;
      RECT  137.75 104.285 137.54 103.905 ;
      RECT  139.19 103.7 139.01 101.995 ;
      RECT  138.47 103.7 138.29 101.995 ;
      RECT  139.19 104.615 139.01 103.7 ;
      RECT  137.03 104.615 136.82 104.285 ;
      RECT  138.83 103.7 138.65 101.995 ;
      RECT  138.83 104.615 138.65 103.7 ;
      RECT  140.15 103.905 139.94 103.7 ;
      RECT  137.03 104.285 136.82 103.905 ;
      RECT  138.11 103.7 137.93 101.995 ;
      RECT  139.94 103.905 139.73 103.7 ;
      RECT  140.15 104.285 139.94 103.905 ;
      POLYGON  137.54 102.62 137.54 102.21 137.285 102.21 137.285 102.54 137.365 102.62 137.54 102.62 ;
      RECT  139.55 104.615 139.37 103.7 ;
      RECT  139.94 104.615 139.73 104.285 ;
      RECT  139.94 104.285 139.73 103.905 ;
      RECT  137.75 104.58 137.54 104.99 ;
      RECT  140.15 103.575 139.94 103.905 ;
      RECT  137.105 104.49 137.03 106.195 ;
      RECT  137.19 105.075 137.105 105.485 ;
      RECT  138.11 103.575 137.93 104.49 ;
      POLYGON  137.105 103.575 137.105 103.905 137.54 103.905 137.54 104.285 137.105 104.285 137.105 104.49 137.03 104.49 137.03 103.575 137.105 103.575 ;
      RECT  137.03 104.49 136.82 106.195 ;
      POLYGON  137.54 104.58 137.54 104.99 137.365 104.99 137.285 104.91 137.285 104.58 137.54 104.58 ;
      RECT  140.15 104.49 139.94 106.195 ;
      RECT  138.47 103.575 138.29 104.49 ;
      RECT  139.55 104.49 139.37 106.195 ;
      RECT  137.75 105.57 137.54 105.98 ;
      RECT  137.03 104.285 136.82 104.49 ;
      RECT  139.94 104.49 139.73 106.195 ;
      RECT  137.75 103.905 137.54 104.285 ;
      RECT  139.19 104.49 139.01 106.195 ;
      RECT  138.47 104.49 138.29 106.195 ;
      RECT  139.19 103.575 139.01 104.49 ;
      RECT  137.03 103.575 136.82 103.905 ;
      RECT  138.83 104.49 138.65 106.195 ;
      RECT  138.83 103.575 138.65 104.49 ;
      RECT  140.15 104.285 139.94 104.49 ;
      RECT  137.03 103.905 136.82 104.285 ;
      RECT  138.11 104.49 137.93 106.195 ;
      RECT  139.94 104.285 139.73 104.49 ;
      RECT  140.15 103.905 139.94 104.285 ;
      POLYGON  137.54 105.57 137.54 105.98 137.285 105.98 137.285 105.65 137.365 105.57 137.54 105.57 ;
      RECT  139.55 103.575 139.37 104.49 ;
      RECT  139.94 103.575 139.73 103.905 ;
      RECT  139.94 103.905 139.73 104.285 ;
      RECT  137.75 107.56 137.54 107.15 ;
      RECT  140.15 108.565 139.94 108.235 ;
      RECT  137.105 107.65 137.03 105.945 ;
      RECT  137.19 107.065 137.105 106.655 ;
      RECT  138.11 108.565 137.93 107.65 ;
      POLYGON  137.105 108.565 137.105 108.235 137.54 108.235 137.54 107.855 137.105 107.855 137.105 107.65 137.03 107.65 137.03 108.565 137.105 108.565 ;
      RECT  137.03 107.65 136.82 105.945 ;
      POLYGON  137.54 107.56 137.54 107.15 137.365 107.15 137.285 107.23 137.285 107.56 137.54 107.56 ;
      RECT  140.15 107.65 139.94 105.945 ;
      RECT  138.47 108.565 138.29 107.65 ;
      RECT  139.55 107.65 139.37 105.945 ;
      RECT  137.75 106.57 137.54 106.16 ;
      RECT  137.03 107.855 136.82 107.65 ;
      RECT  139.94 107.65 139.73 105.945 ;
      RECT  137.75 108.235 137.54 107.855 ;
      RECT  139.19 107.65 139.01 105.945 ;
      RECT  138.47 107.65 138.29 105.945 ;
      RECT  139.19 108.565 139.01 107.65 ;
      RECT  137.03 108.565 136.82 108.235 ;
      RECT  138.83 107.65 138.65 105.945 ;
      RECT  138.83 108.565 138.65 107.65 ;
      RECT  140.15 107.855 139.94 107.65 ;
      RECT  137.03 108.235 136.82 107.855 ;
      RECT  138.11 107.65 137.93 105.945 ;
      RECT  139.94 107.855 139.73 107.65 ;
      RECT  140.15 108.235 139.94 107.855 ;
      POLYGON  137.54 106.57 137.54 106.16 137.285 106.16 137.285 106.49 137.365 106.57 137.54 106.57 ;
      RECT  139.55 108.565 139.37 107.65 ;
      RECT  139.94 108.565 139.73 108.235 ;
      RECT  139.94 108.235 139.73 107.855 ;
      RECT  137.75 108.53 137.54 108.94 ;
      RECT  140.15 107.525 139.94 107.855 ;
      RECT  137.105 108.44 137.03 110.145 ;
      RECT  137.19 109.025 137.105 109.435 ;
      RECT  138.11 107.525 137.93 108.44 ;
      POLYGON  137.105 107.525 137.105 107.855 137.54 107.855 137.54 108.235 137.105 108.235 137.105 108.44 137.03 108.44 137.03 107.525 137.105 107.525 ;
      RECT  137.03 108.44 136.82 110.145 ;
      POLYGON  137.54 108.53 137.54 108.94 137.365 108.94 137.285 108.86 137.285 108.53 137.54 108.53 ;
      RECT  140.15 108.44 139.94 110.145 ;
      RECT  138.47 107.525 138.29 108.44 ;
      RECT  139.55 108.44 139.37 110.145 ;
      RECT  137.75 109.52 137.54 109.93 ;
      RECT  137.03 108.235 136.82 108.44 ;
      RECT  139.94 108.44 139.73 110.145 ;
      RECT  137.75 107.855 137.54 108.235 ;
      RECT  139.19 108.44 139.01 110.145 ;
      RECT  138.47 108.44 138.29 110.145 ;
      RECT  139.19 107.525 139.01 108.44 ;
      RECT  137.03 107.525 136.82 107.855 ;
      RECT  138.83 108.44 138.65 110.145 ;
      RECT  138.83 107.525 138.65 108.44 ;
      RECT  140.15 108.235 139.94 108.44 ;
      RECT  137.03 107.855 136.82 108.235 ;
      RECT  138.11 108.44 137.93 110.145 ;
      RECT  139.94 108.235 139.73 108.44 ;
      RECT  140.15 107.855 139.94 108.235 ;
      POLYGON  137.54 109.52 137.54 109.93 137.285 109.93 137.285 109.6 137.365 109.52 137.54 109.52 ;
      RECT  139.55 107.525 139.37 108.44 ;
      RECT  139.94 107.525 139.73 107.855 ;
      RECT  139.94 107.855 139.73 108.235 ;
      RECT  137.75 111.51 137.54 111.1 ;
      RECT  140.15 112.515 139.94 112.185 ;
      RECT  137.105 111.6 137.03 109.895 ;
      RECT  137.19 111.015 137.105 110.605 ;
      RECT  138.11 112.515 137.93 111.6 ;
      POLYGON  137.105 112.515 137.105 112.185 137.54 112.185 137.54 111.805 137.105 111.805 137.105 111.6 137.03 111.6 137.03 112.515 137.105 112.515 ;
      RECT  137.03 111.6 136.82 109.895 ;
      POLYGON  137.54 111.51 137.54 111.1 137.365 111.1 137.285 111.18 137.285 111.51 137.54 111.51 ;
      RECT  140.15 111.6 139.94 109.895 ;
      RECT  138.47 112.515 138.29 111.6 ;
      RECT  139.55 111.6 139.37 109.895 ;
      RECT  137.75 110.52 137.54 110.11 ;
      RECT  137.03 111.805 136.82 111.6 ;
      RECT  139.94 111.6 139.73 109.895 ;
      RECT  137.75 112.185 137.54 111.805 ;
      RECT  139.19 111.6 139.01 109.895 ;
      RECT  138.47 111.6 138.29 109.895 ;
      RECT  139.19 112.515 139.01 111.6 ;
      RECT  137.03 112.515 136.82 112.185 ;
      RECT  138.83 111.6 138.65 109.895 ;
      RECT  138.83 112.515 138.65 111.6 ;
      RECT  140.15 111.805 139.94 111.6 ;
      RECT  137.03 112.185 136.82 111.805 ;
      RECT  138.11 111.6 137.93 109.895 ;
      RECT  139.94 111.805 139.73 111.6 ;
      RECT  140.15 112.185 139.94 111.805 ;
      POLYGON  137.54 110.52 137.54 110.11 137.285 110.11 137.285 110.44 137.365 110.52 137.54 110.52 ;
      RECT  139.55 112.515 139.37 111.6 ;
      RECT  139.94 112.515 139.73 112.185 ;
      RECT  139.94 112.185 139.73 111.805 ;
      RECT  137.75 112.48 137.54 112.89 ;
      RECT  140.15 111.475 139.94 111.805 ;
      RECT  137.105 112.39 137.03 114.095 ;
      RECT  137.19 112.975 137.105 113.385 ;
      RECT  138.11 111.475 137.93 112.39 ;
      POLYGON  137.105 111.475 137.105 111.805 137.54 111.805 137.54 112.185 137.105 112.185 137.105 112.39 137.03 112.39 137.03 111.475 137.105 111.475 ;
      RECT  137.03 112.39 136.82 114.095 ;
      POLYGON  137.54 112.48 137.54 112.89 137.365 112.89 137.285 112.81 137.285 112.48 137.54 112.48 ;
      RECT  140.15 112.39 139.94 114.095 ;
      RECT  138.47 111.475 138.29 112.39 ;
      RECT  139.55 112.39 139.37 114.095 ;
      RECT  137.75 113.47 137.54 113.88 ;
      RECT  137.03 112.185 136.82 112.39 ;
      RECT  139.94 112.39 139.73 114.095 ;
      RECT  137.75 111.805 137.54 112.185 ;
      RECT  139.19 112.39 139.01 114.095 ;
      RECT  138.47 112.39 138.29 114.095 ;
      RECT  139.19 111.475 139.01 112.39 ;
      RECT  137.03 111.475 136.82 111.805 ;
      RECT  138.83 112.39 138.65 114.095 ;
      RECT  138.83 111.475 138.65 112.39 ;
      RECT  140.15 112.185 139.94 112.39 ;
      RECT  137.03 111.805 136.82 112.185 ;
      RECT  138.11 112.39 137.93 114.095 ;
      RECT  139.94 112.185 139.73 112.39 ;
      RECT  140.15 111.805 139.94 112.185 ;
      POLYGON  137.54 113.47 137.54 113.88 137.285 113.88 137.285 113.55 137.365 113.47 137.54 113.47 ;
      RECT  139.55 111.475 139.37 112.39 ;
      RECT  139.94 111.475 139.73 111.805 ;
      RECT  139.94 111.805 139.73 112.185 ;
      RECT  137.75 115.46 137.54 115.05 ;
      RECT  140.15 116.465 139.94 116.135 ;
      RECT  137.105 115.55 137.03 113.845 ;
      RECT  137.19 114.965 137.105 114.555 ;
      RECT  138.11 116.465 137.93 115.55 ;
      POLYGON  137.105 116.465 137.105 116.135 137.54 116.135 137.54 115.755 137.105 115.755 137.105 115.55 137.03 115.55 137.03 116.465 137.105 116.465 ;
      RECT  137.03 115.55 136.82 113.845 ;
      POLYGON  137.54 115.46 137.54 115.05 137.365 115.05 137.285 115.13 137.285 115.46 137.54 115.46 ;
      RECT  140.15 115.55 139.94 113.845 ;
      RECT  138.47 116.465 138.29 115.55 ;
      RECT  139.55 115.55 139.37 113.845 ;
      RECT  137.75 114.47 137.54 114.06 ;
      RECT  137.03 115.755 136.82 115.55 ;
      RECT  139.94 115.55 139.73 113.845 ;
      RECT  137.75 116.135 137.54 115.755 ;
      RECT  139.19 115.55 139.01 113.845 ;
      RECT  138.47 115.55 138.29 113.845 ;
      RECT  139.19 116.465 139.01 115.55 ;
      RECT  137.03 116.465 136.82 116.135 ;
      RECT  138.83 115.55 138.65 113.845 ;
      RECT  138.83 116.465 138.65 115.55 ;
      RECT  140.15 115.755 139.94 115.55 ;
      RECT  137.03 116.135 136.82 115.755 ;
      RECT  138.11 115.55 137.93 113.845 ;
      RECT  139.94 115.755 139.73 115.55 ;
      RECT  140.15 116.135 139.94 115.755 ;
      POLYGON  137.54 114.47 137.54 114.06 137.285 114.06 137.285 114.39 137.365 114.47 137.54 114.47 ;
      RECT  139.55 116.465 139.37 115.55 ;
      RECT  139.94 116.465 139.73 116.135 ;
      RECT  139.94 116.135 139.73 115.755 ;
      RECT  137.75 116.43 137.54 116.84 ;
      RECT  140.15 115.425 139.94 115.755 ;
      RECT  137.105 116.34 137.03 118.045 ;
      RECT  137.19 116.925 137.105 117.335 ;
      RECT  138.11 115.425 137.93 116.34 ;
      POLYGON  137.105 115.425 137.105 115.755 137.54 115.755 137.54 116.135 137.105 116.135 137.105 116.34 137.03 116.34 137.03 115.425 137.105 115.425 ;
      RECT  137.03 116.34 136.82 118.045 ;
      POLYGON  137.54 116.43 137.54 116.84 137.365 116.84 137.285 116.76 137.285 116.43 137.54 116.43 ;
      RECT  140.15 116.34 139.94 118.045 ;
      RECT  138.47 115.425 138.29 116.34 ;
      RECT  139.55 116.34 139.37 118.045 ;
      RECT  137.75 117.42 137.54 117.83 ;
      RECT  137.03 116.135 136.82 116.34 ;
      RECT  139.94 116.34 139.73 118.045 ;
      RECT  137.75 115.755 137.54 116.135 ;
      RECT  139.19 116.34 139.01 118.045 ;
      RECT  138.47 116.34 138.29 118.045 ;
      RECT  139.19 115.425 139.01 116.34 ;
      RECT  137.03 115.425 136.82 115.755 ;
      RECT  138.83 116.34 138.65 118.045 ;
      RECT  138.83 115.425 138.65 116.34 ;
      RECT  140.15 116.135 139.94 116.34 ;
      RECT  137.03 115.755 136.82 116.135 ;
      RECT  138.11 116.34 137.93 118.045 ;
      RECT  139.94 116.135 139.73 116.34 ;
      RECT  140.15 115.755 139.94 116.135 ;
      POLYGON  137.54 117.42 137.54 117.83 137.285 117.83 137.285 117.5 137.365 117.42 137.54 117.42 ;
      RECT  139.55 115.425 139.37 116.34 ;
      RECT  139.94 115.425 139.73 115.755 ;
      RECT  139.94 115.755 139.73 116.135 ;
      RECT  137.75 119.41 137.54 119.0 ;
      RECT  140.15 120.415 139.94 120.085 ;
      RECT  137.105 119.5 137.03 117.795 ;
      RECT  137.19 118.915 137.105 118.505 ;
      RECT  138.11 120.415 137.93 119.5 ;
      POLYGON  137.105 120.415 137.105 120.085 137.54 120.085 137.54 119.705 137.105 119.705 137.105 119.5 137.03 119.5 137.03 120.415 137.105 120.415 ;
      RECT  137.03 119.5 136.82 117.795 ;
      POLYGON  137.54 119.41 137.54 119.0 137.365 119.0 137.285 119.08 137.285 119.41 137.54 119.41 ;
      RECT  140.15 119.5 139.94 117.795 ;
      RECT  138.47 120.415 138.29 119.5 ;
      RECT  139.55 119.5 139.37 117.795 ;
      RECT  137.75 118.42 137.54 118.01 ;
      RECT  137.03 119.705 136.82 119.5 ;
      RECT  139.94 119.5 139.73 117.795 ;
      RECT  137.75 120.085 137.54 119.705 ;
      RECT  139.19 119.5 139.01 117.795 ;
      RECT  138.47 119.5 138.29 117.795 ;
      RECT  139.19 120.415 139.01 119.5 ;
      RECT  137.03 120.415 136.82 120.085 ;
      RECT  138.83 119.5 138.65 117.795 ;
      RECT  138.83 120.415 138.65 119.5 ;
      RECT  140.15 119.705 139.94 119.5 ;
      RECT  137.03 120.085 136.82 119.705 ;
      RECT  138.11 119.5 137.93 117.795 ;
      RECT  139.94 119.705 139.73 119.5 ;
      RECT  140.15 120.085 139.94 119.705 ;
      POLYGON  137.54 118.42 137.54 118.01 137.285 118.01 137.285 118.34 137.365 118.42 137.54 118.42 ;
      RECT  139.55 120.415 139.37 119.5 ;
      RECT  139.94 120.415 139.73 120.085 ;
      RECT  139.94 120.085 139.73 119.705 ;
      RECT  137.75 120.38 137.54 120.79 ;
      RECT  140.15 119.375 139.94 119.705 ;
      RECT  137.105 120.29 137.03 121.995 ;
      RECT  137.19 120.875 137.105 121.285 ;
      RECT  138.11 119.375 137.93 120.29 ;
      POLYGON  137.105 119.375 137.105 119.705 137.54 119.705 137.54 120.085 137.105 120.085 137.105 120.29 137.03 120.29 137.03 119.375 137.105 119.375 ;
      RECT  137.03 120.29 136.82 121.995 ;
      POLYGON  137.54 120.38 137.54 120.79 137.365 120.79 137.285 120.71 137.285 120.38 137.54 120.38 ;
      RECT  140.15 120.29 139.94 121.995 ;
      RECT  138.47 119.375 138.29 120.29 ;
      RECT  139.55 120.29 139.37 121.995 ;
      RECT  137.75 121.37 137.54 121.78 ;
      RECT  137.03 120.085 136.82 120.29 ;
      RECT  139.94 120.29 139.73 121.995 ;
      RECT  137.75 119.705 137.54 120.085 ;
      RECT  139.19 120.29 139.01 121.995 ;
      RECT  138.47 120.29 138.29 121.995 ;
      RECT  139.19 119.375 139.01 120.29 ;
      RECT  137.03 119.375 136.82 119.705 ;
      RECT  138.83 120.29 138.65 121.995 ;
      RECT  138.83 119.375 138.65 120.29 ;
      RECT  140.15 120.085 139.94 120.29 ;
      RECT  137.03 119.705 136.82 120.085 ;
      RECT  138.11 120.29 137.93 121.995 ;
      RECT  139.94 120.085 139.73 120.29 ;
      RECT  140.15 119.705 139.94 120.085 ;
      POLYGON  137.54 121.37 137.54 121.78 137.285 121.78 137.285 121.45 137.365 121.37 137.54 121.37 ;
      RECT  139.55 119.375 139.37 120.29 ;
      RECT  139.94 119.375 139.73 119.705 ;
      RECT  139.94 119.705 139.73 120.085 ;
      RECT  137.75 123.36 137.54 122.95 ;
      RECT  140.15 124.365 139.94 124.035 ;
      RECT  137.105 123.45 137.03 121.745 ;
      RECT  137.19 122.865 137.105 122.455 ;
      RECT  138.11 124.365 137.93 123.45 ;
      POLYGON  137.105 124.365 137.105 124.035 137.54 124.035 137.54 123.655 137.105 123.655 137.105 123.45 137.03 123.45 137.03 124.365 137.105 124.365 ;
      RECT  137.03 123.45 136.82 121.745 ;
      POLYGON  137.54 123.36 137.54 122.95 137.365 122.95 137.285 123.03 137.285 123.36 137.54 123.36 ;
      RECT  140.15 123.45 139.94 121.745 ;
      RECT  138.47 124.365 138.29 123.45 ;
      RECT  139.55 123.45 139.37 121.745 ;
      RECT  137.75 122.37 137.54 121.96 ;
      RECT  137.03 123.655 136.82 123.45 ;
      RECT  139.94 123.45 139.73 121.745 ;
      RECT  137.75 124.035 137.54 123.655 ;
      RECT  139.19 123.45 139.01 121.745 ;
      RECT  138.47 123.45 138.29 121.745 ;
      RECT  139.19 124.365 139.01 123.45 ;
      RECT  137.03 124.365 136.82 124.035 ;
      RECT  138.83 123.45 138.65 121.745 ;
      RECT  138.83 124.365 138.65 123.45 ;
      RECT  140.15 123.655 139.94 123.45 ;
      RECT  137.03 124.035 136.82 123.655 ;
      RECT  138.11 123.45 137.93 121.745 ;
      RECT  139.94 123.655 139.73 123.45 ;
      RECT  140.15 124.035 139.94 123.655 ;
      POLYGON  137.54 122.37 137.54 121.96 137.285 121.96 137.285 122.29 137.365 122.37 137.54 122.37 ;
      RECT  139.55 124.365 139.37 123.45 ;
      RECT  139.94 124.365 139.73 124.035 ;
      RECT  139.94 124.035 139.73 123.655 ;
      RECT  142.13 92.73 142.34 93.14 ;
      RECT  139.73 91.725 139.94 92.055 ;
      RECT  142.775 92.64 142.85 94.345 ;
      RECT  142.69 93.225 142.775 93.635 ;
      RECT  141.77 91.725 141.95 92.64 ;
      POLYGON  142.775 91.725 142.775 92.055 142.34 92.055 142.34 92.435 142.775 92.435 142.775 92.64 142.85 92.64 142.85 91.725 142.775 91.725 ;
      RECT  142.85 92.64 143.06 94.345 ;
      POLYGON  142.34 92.73 142.34 93.14 142.515 93.14 142.595 93.06 142.595 92.73 142.34 92.73 ;
      RECT  139.73 92.64 139.94 94.345 ;
      RECT  141.41 91.725 141.59 92.64 ;
      RECT  140.33 92.64 140.51 94.345 ;
      RECT  142.13 93.72 142.34 94.13 ;
      RECT  142.85 92.435 143.06 92.64 ;
      RECT  139.94 92.64 140.15 94.345 ;
      RECT  142.13 92.055 142.34 92.435 ;
      RECT  140.69 92.64 140.87 94.345 ;
      RECT  141.41 92.64 141.59 94.345 ;
      RECT  140.69 91.725 140.87 92.64 ;
      RECT  142.85 91.725 143.06 92.055 ;
      RECT  141.05 92.64 141.23 94.345 ;
      RECT  141.05 91.725 141.23 92.64 ;
      RECT  139.73 92.435 139.94 92.64 ;
      RECT  142.85 92.055 143.06 92.435 ;
      RECT  141.77 92.64 141.95 94.345 ;
      RECT  139.94 92.435 140.15 92.64 ;
      RECT  139.73 92.055 139.94 92.435 ;
      POLYGON  142.34 93.72 142.34 94.13 142.595 94.13 142.595 93.8 142.515 93.72 142.34 93.72 ;
      RECT  140.33 91.725 140.51 92.64 ;
      RECT  139.94 91.725 140.15 92.055 ;
      RECT  139.94 92.055 140.15 92.435 ;
      RECT  142.13 95.71 142.34 95.3 ;
      RECT  139.73 96.715 139.94 96.385 ;
      RECT  142.775 95.8 142.85 94.095 ;
      RECT  142.69 95.215 142.775 94.805 ;
      RECT  141.77 96.715 141.95 95.8 ;
      POLYGON  142.775 96.715 142.775 96.385 142.34 96.385 142.34 96.005 142.775 96.005 142.775 95.8 142.85 95.8 142.85 96.715 142.775 96.715 ;
      RECT  142.85 95.8 143.06 94.095 ;
      POLYGON  142.34 95.71 142.34 95.3 142.515 95.3 142.595 95.38 142.595 95.71 142.34 95.71 ;
      RECT  139.73 95.8 139.94 94.095 ;
      RECT  141.41 96.715 141.59 95.8 ;
      RECT  140.33 95.8 140.51 94.095 ;
      RECT  142.13 94.72 142.34 94.31 ;
      RECT  142.85 96.005 143.06 95.8 ;
      RECT  139.94 95.8 140.15 94.095 ;
      RECT  142.13 96.385 142.34 96.005 ;
      RECT  140.69 95.8 140.87 94.095 ;
      RECT  141.41 95.8 141.59 94.095 ;
      RECT  140.69 96.715 140.87 95.8 ;
      RECT  142.85 96.715 143.06 96.385 ;
      RECT  141.05 95.8 141.23 94.095 ;
      RECT  141.05 96.715 141.23 95.8 ;
      RECT  139.73 96.005 139.94 95.8 ;
      RECT  142.85 96.385 143.06 96.005 ;
      RECT  141.77 95.8 141.95 94.095 ;
      RECT  139.94 96.005 140.15 95.8 ;
      RECT  139.73 96.385 139.94 96.005 ;
      POLYGON  142.34 94.72 142.34 94.31 142.595 94.31 142.595 94.64 142.515 94.72 142.34 94.72 ;
      RECT  140.33 96.715 140.51 95.8 ;
      RECT  139.94 96.715 140.15 96.385 ;
      RECT  139.94 96.385 140.15 96.005 ;
      RECT  142.13 96.68 142.34 97.09 ;
      RECT  139.73 95.675 139.94 96.005 ;
      RECT  142.775 96.59 142.85 98.295 ;
      RECT  142.69 97.175 142.775 97.585 ;
      RECT  141.77 95.675 141.95 96.59 ;
      POLYGON  142.775 95.675 142.775 96.005 142.34 96.005 142.34 96.385 142.775 96.385 142.775 96.59 142.85 96.59 142.85 95.675 142.775 95.675 ;
      RECT  142.85 96.59 143.06 98.295 ;
      POLYGON  142.34 96.68 142.34 97.09 142.515 97.09 142.595 97.01 142.595 96.68 142.34 96.68 ;
      RECT  139.73 96.59 139.94 98.295 ;
      RECT  141.41 95.675 141.59 96.59 ;
      RECT  140.33 96.59 140.51 98.295 ;
      RECT  142.13 97.67 142.34 98.08 ;
      RECT  142.85 96.385 143.06 96.59 ;
      RECT  139.94 96.59 140.15 98.295 ;
      RECT  142.13 96.005 142.34 96.385 ;
      RECT  140.69 96.59 140.87 98.295 ;
      RECT  141.41 96.59 141.59 98.295 ;
      RECT  140.69 95.675 140.87 96.59 ;
      RECT  142.85 95.675 143.06 96.005 ;
      RECT  141.05 96.59 141.23 98.295 ;
      RECT  141.05 95.675 141.23 96.59 ;
      RECT  139.73 96.385 139.94 96.59 ;
      RECT  142.85 96.005 143.06 96.385 ;
      RECT  141.77 96.59 141.95 98.295 ;
      RECT  139.94 96.385 140.15 96.59 ;
      RECT  139.73 96.005 139.94 96.385 ;
      POLYGON  142.34 97.67 142.34 98.08 142.595 98.08 142.595 97.75 142.515 97.67 142.34 97.67 ;
      RECT  140.33 95.675 140.51 96.59 ;
      RECT  139.94 95.675 140.15 96.005 ;
      RECT  139.94 96.005 140.15 96.385 ;
      RECT  142.13 99.66 142.34 99.25 ;
      RECT  139.73 100.665 139.94 100.335 ;
      RECT  142.775 99.75 142.85 98.045 ;
      RECT  142.69 99.165 142.775 98.755 ;
      RECT  141.77 100.665 141.95 99.75 ;
      POLYGON  142.775 100.665 142.775 100.335 142.34 100.335 142.34 99.955 142.775 99.955 142.775 99.75 142.85 99.75 142.85 100.665 142.775 100.665 ;
      RECT  142.85 99.75 143.06 98.045 ;
      POLYGON  142.34 99.66 142.34 99.25 142.515 99.25 142.595 99.33 142.595 99.66 142.34 99.66 ;
      RECT  139.73 99.75 139.94 98.045 ;
      RECT  141.41 100.665 141.59 99.75 ;
      RECT  140.33 99.75 140.51 98.045 ;
      RECT  142.13 98.67 142.34 98.26 ;
      RECT  142.85 99.955 143.06 99.75 ;
      RECT  139.94 99.75 140.15 98.045 ;
      RECT  142.13 100.335 142.34 99.955 ;
      RECT  140.69 99.75 140.87 98.045 ;
      RECT  141.41 99.75 141.59 98.045 ;
      RECT  140.69 100.665 140.87 99.75 ;
      RECT  142.85 100.665 143.06 100.335 ;
      RECT  141.05 99.75 141.23 98.045 ;
      RECT  141.05 100.665 141.23 99.75 ;
      RECT  139.73 99.955 139.94 99.75 ;
      RECT  142.85 100.335 143.06 99.955 ;
      RECT  141.77 99.75 141.95 98.045 ;
      RECT  139.94 99.955 140.15 99.75 ;
      RECT  139.73 100.335 139.94 99.955 ;
      POLYGON  142.34 98.67 142.34 98.26 142.595 98.26 142.595 98.59 142.515 98.67 142.34 98.67 ;
      RECT  140.33 100.665 140.51 99.75 ;
      RECT  139.94 100.665 140.15 100.335 ;
      RECT  139.94 100.335 140.15 99.955 ;
      RECT  142.13 100.63 142.34 101.04 ;
      RECT  139.73 99.625 139.94 99.955 ;
      RECT  142.775 100.54 142.85 102.245 ;
      RECT  142.69 101.125 142.775 101.535 ;
      RECT  141.77 99.625 141.95 100.54 ;
      POLYGON  142.775 99.625 142.775 99.955 142.34 99.955 142.34 100.335 142.775 100.335 142.775 100.54 142.85 100.54 142.85 99.625 142.775 99.625 ;
      RECT  142.85 100.54 143.06 102.245 ;
      POLYGON  142.34 100.63 142.34 101.04 142.515 101.04 142.595 100.96 142.595 100.63 142.34 100.63 ;
      RECT  139.73 100.54 139.94 102.245 ;
      RECT  141.41 99.625 141.59 100.54 ;
      RECT  140.33 100.54 140.51 102.245 ;
      RECT  142.13 101.62 142.34 102.03 ;
      RECT  142.85 100.335 143.06 100.54 ;
      RECT  139.94 100.54 140.15 102.245 ;
      RECT  142.13 99.955 142.34 100.335 ;
      RECT  140.69 100.54 140.87 102.245 ;
      RECT  141.41 100.54 141.59 102.245 ;
      RECT  140.69 99.625 140.87 100.54 ;
      RECT  142.85 99.625 143.06 99.955 ;
      RECT  141.05 100.54 141.23 102.245 ;
      RECT  141.05 99.625 141.23 100.54 ;
      RECT  139.73 100.335 139.94 100.54 ;
      RECT  142.85 99.955 143.06 100.335 ;
      RECT  141.77 100.54 141.95 102.245 ;
      RECT  139.94 100.335 140.15 100.54 ;
      RECT  139.73 99.955 139.94 100.335 ;
      POLYGON  142.34 101.62 142.34 102.03 142.595 102.03 142.595 101.7 142.515 101.62 142.34 101.62 ;
      RECT  140.33 99.625 140.51 100.54 ;
      RECT  139.94 99.625 140.15 99.955 ;
      RECT  139.94 99.955 140.15 100.335 ;
      RECT  142.13 103.61 142.34 103.2 ;
      RECT  139.73 104.615 139.94 104.285 ;
      RECT  142.775 103.7 142.85 101.995 ;
      RECT  142.69 103.115 142.775 102.705 ;
      RECT  141.77 104.615 141.95 103.7 ;
      POLYGON  142.775 104.615 142.775 104.285 142.34 104.285 142.34 103.905 142.775 103.905 142.775 103.7 142.85 103.7 142.85 104.615 142.775 104.615 ;
      RECT  142.85 103.7 143.06 101.995 ;
      POLYGON  142.34 103.61 142.34 103.2 142.515 103.2 142.595 103.28 142.595 103.61 142.34 103.61 ;
      RECT  139.73 103.7 139.94 101.995 ;
      RECT  141.41 104.615 141.59 103.7 ;
      RECT  140.33 103.7 140.51 101.995 ;
      RECT  142.13 102.62 142.34 102.21 ;
      RECT  142.85 103.905 143.06 103.7 ;
      RECT  139.94 103.7 140.15 101.995 ;
      RECT  142.13 104.285 142.34 103.905 ;
      RECT  140.69 103.7 140.87 101.995 ;
      RECT  141.41 103.7 141.59 101.995 ;
      RECT  140.69 104.615 140.87 103.7 ;
      RECT  142.85 104.615 143.06 104.285 ;
      RECT  141.05 103.7 141.23 101.995 ;
      RECT  141.05 104.615 141.23 103.7 ;
      RECT  139.73 103.905 139.94 103.7 ;
      RECT  142.85 104.285 143.06 103.905 ;
      RECT  141.77 103.7 141.95 101.995 ;
      RECT  139.94 103.905 140.15 103.7 ;
      RECT  139.73 104.285 139.94 103.905 ;
      POLYGON  142.34 102.62 142.34 102.21 142.595 102.21 142.595 102.54 142.515 102.62 142.34 102.62 ;
      RECT  140.33 104.615 140.51 103.7 ;
      RECT  139.94 104.615 140.15 104.285 ;
      RECT  139.94 104.285 140.15 103.905 ;
      RECT  142.13 104.58 142.34 104.99 ;
      RECT  139.73 103.575 139.94 103.905 ;
      RECT  142.775 104.49 142.85 106.195 ;
      RECT  142.69 105.075 142.775 105.485 ;
      RECT  141.77 103.575 141.95 104.49 ;
      POLYGON  142.775 103.575 142.775 103.905 142.34 103.905 142.34 104.285 142.775 104.285 142.775 104.49 142.85 104.49 142.85 103.575 142.775 103.575 ;
      RECT  142.85 104.49 143.06 106.195 ;
      POLYGON  142.34 104.58 142.34 104.99 142.515 104.99 142.595 104.91 142.595 104.58 142.34 104.58 ;
      RECT  139.73 104.49 139.94 106.195 ;
      RECT  141.41 103.575 141.59 104.49 ;
      RECT  140.33 104.49 140.51 106.195 ;
      RECT  142.13 105.57 142.34 105.98 ;
      RECT  142.85 104.285 143.06 104.49 ;
      RECT  139.94 104.49 140.15 106.195 ;
      RECT  142.13 103.905 142.34 104.285 ;
      RECT  140.69 104.49 140.87 106.195 ;
      RECT  141.41 104.49 141.59 106.195 ;
      RECT  140.69 103.575 140.87 104.49 ;
      RECT  142.85 103.575 143.06 103.905 ;
      RECT  141.05 104.49 141.23 106.195 ;
      RECT  141.05 103.575 141.23 104.49 ;
      RECT  139.73 104.285 139.94 104.49 ;
      RECT  142.85 103.905 143.06 104.285 ;
      RECT  141.77 104.49 141.95 106.195 ;
      RECT  139.94 104.285 140.15 104.49 ;
      RECT  139.73 103.905 139.94 104.285 ;
      POLYGON  142.34 105.57 142.34 105.98 142.595 105.98 142.595 105.65 142.515 105.57 142.34 105.57 ;
      RECT  140.33 103.575 140.51 104.49 ;
      RECT  139.94 103.575 140.15 103.905 ;
      RECT  139.94 103.905 140.15 104.285 ;
      RECT  142.13 107.56 142.34 107.15 ;
      RECT  139.73 108.565 139.94 108.235 ;
      RECT  142.775 107.65 142.85 105.945 ;
      RECT  142.69 107.065 142.775 106.655 ;
      RECT  141.77 108.565 141.95 107.65 ;
      POLYGON  142.775 108.565 142.775 108.235 142.34 108.235 142.34 107.855 142.775 107.855 142.775 107.65 142.85 107.65 142.85 108.565 142.775 108.565 ;
      RECT  142.85 107.65 143.06 105.945 ;
      POLYGON  142.34 107.56 142.34 107.15 142.515 107.15 142.595 107.23 142.595 107.56 142.34 107.56 ;
      RECT  139.73 107.65 139.94 105.945 ;
      RECT  141.41 108.565 141.59 107.65 ;
      RECT  140.33 107.65 140.51 105.945 ;
      RECT  142.13 106.57 142.34 106.16 ;
      RECT  142.85 107.855 143.06 107.65 ;
      RECT  139.94 107.65 140.15 105.945 ;
      RECT  142.13 108.235 142.34 107.855 ;
      RECT  140.69 107.65 140.87 105.945 ;
      RECT  141.41 107.65 141.59 105.945 ;
      RECT  140.69 108.565 140.87 107.65 ;
      RECT  142.85 108.565 143.06 108.235 ;
      RECT  141.05 107.65 141.23 105.945 ;
      RECT  141.05 108.565 141.23 107.65 ;
      RECT  139.73 107.855 139.94 107.65 ;
      RECT  142.85 108.235 143.06 107.855 ;
      RECT  141.77 107.65 141.95 105.945 ;
      RECT  139.94 107.855 140.15 107.65 ;
      RECT  139.73 108.235 139.94 107.855 ;
      POLYGON  142.34 106.57 142.34 106.16 142.595 106.16 142.595 106.49 142.515 106.57 142.34 106.57 ;
      RECT  140.33 108.565 140.51 107.65 ;
      RECT  139.94 108.565 140.15 108.235 ;
      RECT  139.94 108.235 140.15 107.855 ;
      RECT  142.13 108.53 142.34 108.94 ;
      RECT  139.73 107.525 139.94 107.855 ;
      RECT  142.775 108.44 142.85 110.145 ;
      RECT  142.69 109.025 142.775 109.435 ;
      RECT  141.77 107.525 141.95 108.44 ;
      POLYGON  142.775 107.525 142.775 107.855 142.34 107.855 142.34 108.235 142.775 108.235 142.775 108.44 142.85 108.44 142.85 107.525 142.775 107.525 ;
      RECT  142.85 108.44 143.06 110.145 ;
      POLYGON  142.34 108.53 142.34 108.94 142.515 108.94 142.595 108.86 142.595 108.53 142.34 108.53 ;
      RECT  139.73 108.44 139.94 110.145 ;
      RECT  141.41 107.525 141.59 108.44 ;
      RECT  140.33 108.44 140.51 110.145 ;
      RECT  142.13 109.52 142.34 109.93 ;
      RECT  142.85 108.235 143.06 108.44 ;
      RECT  139.94 108.44 140.15 110.145 ;
      RECT  142.13 107.855 142.34 108.235 ;
      RECT  140.69 108.44 140.87 110.145 ;
      RECT  141.41 108.44 141.59 110.145 ;
      RECT  140.69 107.525 140.87 108.44 ;
      RECT  142.85 107.525 143.06 107.855 ;
      RECT  141.05 108.44 141.23 110.145 ;
      RECT  141.05 107.525 141.23 108.44 ;
      RECT  139.73 108.235 139.94 108.44 ;
      RECT  142.85 107.855 143.06 108.235 ;
      RECT  141.77 108.44 141.95 110.145 ;
      RECT  139.94 108.235 140.15 108.44 ;
      RECT  139.73 107.855 139.94 108.235 ;
      POLYGON  142.34 109.52 142.34 109.93 142.595 109.93 142.595 109.6 142.515 109.52 142.34 109.52 ;
      RECT  140.33 107.525 140.51 108.44 ;
      RECT  139.94 107.525 140.15 107.855 ;
      RECT  139.94 107.855 140.15 108.235 ;
      RECT  142.13 111.51 142.34 111.1 ;
      RECT  139.73 112.515 139.94 112.185 ;
      RECT  142.775 111.6 142.85 109.895 ;
      RECT  142.69 111.015 142.775 110.605 ;
      RECT  141.77 112.515 141.95 111.6 ;
      POLYGON  142.775 112.515 142.775 112.185 142.34 112.185 142.34 111.805 142.775 111.805 142.775 111.6 142.85 111.6 142.85 112.515 142.775 112.515 ;
      RECT  142.85 111.6 143.06 109.895 ;
      POLYGON  142.34 111.51 142.34 111.1 142.515 111.1 142.595 111.18 142.595 111.51 142.34 111.51 ;
      RECT  139.73 111.6 139.94 109.895 ;
      RECT  141.41 112.515 141.59 111.6 ;
      RECT  140.33 111.6 140.51 109.895 ;
      RECT  142.13 110.52 142.34 110.11 ;
      RECT  142.85 111.805 143.06 111.6 ;
      RECT  139.94 111.6 140.15 109.895 ;
      RECT  142.13 112.185 142.34 111.805 ;
      RECT  140.69 111.6 140.87 109.895 ;
      RECT  141.41 111.6 141.59 109.895 ;
      RECT  140.69 112.515 140.87 111.6 ;
      RECT  142.85 112.515 143.06 112.185 ;
      RECT  141.05 111.6 141.23 109.895 ;
      RECT  141.05 112.515 141.23 111.6 ;
      RECT  139.73 111.805 139.94 111.6 ;
      RECT  142.85 112.185 143.06 111.805 ;
      RECT  141.77 111.6 141.95 109.895 ;
      RECT  139.94 111.805 140.15 111.6 ;
      RECT  139.73 112.185 139.94 111.805 ;
      POLYGON  142.34 110.52 142.34 110.11 142.595 110.11 142.595 110.44 142.515 110.52 142.34 110.52 ;
      RECT  140.33 112.515 140.51 111.6 ;
      RECT  139.94 112.515 140.15 112.185 ;
      RECT  139.94 112.185 140.15 111.805 ;
      RECT  142.13 112.48 142.34 112.89 ;
      RECT  139.73 111.475 139.94 111.805 ;
      RECT  142.775 112.39 142.85 114.095 ;
      RECT  142.69 112.975 142.775 113.385 ;
      RECT  141.77 111.475 141.95 112.39 ;
      POLYGON  142.775 111.475 142.775 111.805 142.34 111.805 142.34 112.185 142.775 112.185 142.775 112.39 142.85 112.39 142.85 111.475 142.775 111.475 ;
      RECT  142.85 112.39 143.06 114.095 ;
      POLYGON  142.34 112.48 142.34 112.89 142.515 112.89 142.595 112.81 142.595 112.48 142.34 112.48 ;
      RECT  139.73 112.39 139.94 114.095 ;
      RECT  141.41 111.475 141.59 112.39 ;
      RECT  140.33 112.39 140.51 114.095 ;
      RECT  142.13 113.47 142.34 113.88 ;
      RECT  142.85 112.185 143.06 112.39 ;
      RECT  139.94 112.39 140.15 114.095 ;
      RECT  142.13 111.805 142.34 112.185 ;
      RECT  140.69 112.39 140.87 114.095 ;
      RECT  141.41 112.39 141.59 114.095 ;
      RECT  140.69 111.475 140.87 112.39 ;
      RECT  142.85 111.475 143.06 111.805 ;
      RECT  141.05 112.39 141.23 114.095 ;
      RECT  141.05 111.475 141.23 112.39 ;
      RECT  139.73 112.185 139.94 112.39 ;
      RECT  142.85 111.805 143.06 112.185 ;
      RECT  141.77 112.39 141.95 114.095 ;
      RECT  139.94 112.185 140.15 112.39 ;
      RECT  139.73 111.805 139.94 112.185 ;
      POLYGON  142.34 113.47 142.34 113.88 142.595 113.88 142.595 113.55 142.515 113.47 142.34 113.47 ;
      RECT  140.33 111.475 140.51 112.39 ;
      RECT  139.94 111.475 140.15 111.805 ;
      RECT  139.94 111.805 140.15 112.185 ;
      RECT  142.13 115.46 142.34 115.05 ;
      RECT  139.73 116.465 139.94 116.135 ;
      RECT  142.775 115.55 142.85 113.845 ;
      RECT  142.69 114.965 142.775 114.555 ;
      RECT  141.77 116.465 141.95 115.55 ;
      POLYGON  142.775 116.465 142.775 116.135 142.34 116.135 142.34 115.755 142.775 115.755 142.775 115.55 142.85 115.55 142.85 116.465 142.775 116.465 ;
      RECT  142.85 115.55 143.06 113.845 ;
      POLYGON  142.34 115.46 142.34 115.05 142.515 115.05 142.595 115.13 142.595 115.46 142.34 115.46 ;
      RECT  139.73 115.55 139.94 113.845 ;
      RECT  141.41 116.465 141.59 115.55 ;
      RECT  140.33 115.55 140.51 113.845 ;
      RECT  142.13 114.47 142.34 114.06 ;
      RECT  142.85 115.755 143.06 115.55 ;
      RECT  139.94 115.55 140.15 113.845 ;
      RECT  142.13 116.135 142.34 115.755 ;
      RECT  140.69 115.55 140.87 113.845 ;
      RECT  141.41 115.55 141.59 113.845 ;
      RECT  140.69 116.465 140.87 115.55 ;
      RECT  142.85 116.465 143.06 116.135 ;
      RECT  141.05 115.55 141.23 113.845 ;
      RECT  141.05 116.465 141.23 115.55 ;
      RECT  139.73 115.755 139.94 115.55 ;
      RECT  142.85 116.135 143.06 115.755 ;
      RECT  141.77 115.55 141.95 113.845 ;
      RECT  139.94 115.755 140.15 115.55 ;
      RECT  139.73 116.135 139.94 115.755 ;
      POLYGON  142.34 114.47 142.34 114.06 142.595 114.06 142.595 114.39 142.515 114.47 142.34 114.47 ;
      RECT  140.33 116.465 140.51 115.55 ;
      RECT  139.94 116.465 140.15 116.135 ;
      RECT  139.94 116.135 140.15 115.755 ;
      RECT  142.13 116.43 142.34 116.84 ;
      RECT  139.73 115.425 139.94 115.755 ;
      RECT  142.775 116.34 142.85 118.045 ;
      RECT  142.69 116.925 142.775 117.335 ;
      RECT  141.77 115.425 141.95 116.34 ;
      POLYGON  142.775 115.425 142.775 115.755 142.34 115.755 142.34 116.135 142.775 116.135 142.775 116.34 142.85 116.34 142.85 115.425 142.775 115.425 ;
      RECT  142.85 116.34 143.06 118.045 ;
      POLYGON  142.34 116.43 142.34 116.84 142.515 116.84 142.595 116.76 142.595 116.43 142.34 116.43 ;
      RECT  139.73 116.34 139.94 118.045 ;
      RECT  141.41 115.425 141.59 116.34 ;
      RECT  140.33 116.34 140.51 118.045 ;
      RECT  142.13 117.42 142.34 117.83 ;
      RECT  142.85 116.135 143.06 116.34 ;
      RECT  139.94 116.34 140.15 118.045 ;
      RECT  142.13 115.755 142.34 116.135 ;
      RECT  140.69 116.34 140.87 118.045 ;
      RECT  141.41 116.34 141.59 118.045 ;
      RECT  140.69 115.425 140.87 116.34 ;
      RECT  142.85 115.425 143.06 115.755 ;
      RECT  141.05 116.34 141.23 118.045 ;
      RECT  141.05 115.425 141.23 116.34 ;
      RECT  139.73 116.135 139.94 116.34 ;
      RECT  142.85 115.755 143.06 116.135 ;
      RECT  141.77 116.34 141.95 118.045 ;
      RECT  139.94 116.135 140.15 116.34 ;
      RECT  139.73 115.755 139.94 116.135 ;
      POLYGON  142.34 117.42 142.34 117.83 142.595 117.83 142.595 117.5 142.515 117.42 142.34 117.42 ;
      RECT  140.33 115.425 140.51 116.34 ;
      RECT  139.94 115.425 140.15 115.755 ;
      RECT  139.94 115.755 140.15 116.135 ;
      RECT  142.13 119.41 142.34 119.0 ;
      RECT  139.73 120.415 139.94 120.085 ;
      RECT  142.775 119.5 142.85 117.795 ;
      RECT  142.69 118.915 142.775 118.505 ;
      RECT  141.77 120.415 141.95 119.5 ;
      POLYGON  142.775 120.415 142.775 120.085 142.34 120.085 142.34 119.705 142.775 119.705 142.775 119.5 142.85 119.5 142.85 120.415 142.775 120.415 ;
      RECT  142.85 119.5 143.06 117.795 ;
      POLYGON  142.34 119.41 142.34 119.0 142.515 119.0 142.595 119.08 142.595 119.41 142.34 119.41 ;
      RECT  139.73 119.5 139.94 117.795 ;
      RECT  141.41 120.415 141.59 119.5 ;
      RECT  140.33 119.5 140.51 117.795 ;
      RECT  142.13 118.42 142.34 118.01 ;
      RECT  142.85 119.705 143.06 119.5 ;
      RECT  139.94 119.5 140.15 117.795 ;
      RECT  142.13 120.085 142.34 119.705 ;
      RECT  140.69 119.5 140.87 117.795 ;
      RECT  141.41 119.5 141.59 117.795 ;
      RECT  140.69 120.415 140.87 119.5 ;
      RECT  142.85 120.415 143.06 120.085 ;
      RECT  141.05 119.5 141.23 117.795 ;
      RECT  141.05 120.415 141.23 119.5 ;
      RECT  139.73 119.705 139.94 119.5 ;
      RECT  142.85 120.085 143.06 119.705 ;
      RECT  141.77 119.5 141.95 117.795 ;
      RECT  139.94 119.705 140.15 119.5 ;
      RECT  139.73 120.085 139.94 119.705 ;
      POLYGON  142.34 118.42 142.34 118.01 142.595 118.01 142.595 118.34 142.515 118.42 142.34 118.42 ;
      RECT  140.33 120.415 140.51 119.5 ;
      RECT  139.94 120.415 140.15 120.085 ;
      RECT  139.94 120.085 140.15 119.705 ;
      RECT  142.13 120.38 142.34 120.79 ;
      RECT  139.73 119.375 139.94 119.705 ;
      RECT  142.775 120.29 142.85 121.995 ;
      RECT  142.69 120.875 142.775 121.285 ;
      RECT  141.77 119.375 141.95 120.29 ;
      POLYGON  142.775 119.375 142.775 119.705 142.34 119.705 142.34 120.085 142.775 120.085 142.775 120.29 142.85 120.29 142.85 119.375 142.775 119.375 ;
      RECT  142.85 120.29 143.06 121.995 ;
      POLYGON  142.34 120.38 142.34 120.79 142.515 120.79 142.595 120.71 142.595 120.38 142.34 120.38 ;
      RECT  139.73 120.29 139.94 121.995 ;
      RECT  141.41 119.375 141.59 120.29 ;
      RECT  140.33 120.29 140.51 121.995 ;
      RECT  142.13 121.37 142.34 121.78 ;
      RECT  142.85 120.085 143.06 120.29 ;
      RECT  139.94 120.29 140.15 121.995 ;
      RECT  142.13 119.705 142.34 120.085 ;
      RECT  140.69 120.29 140.87 121.995 ;
      RECT  141.41 120.29 141.59 121.995 ;
      RECT  140.69 119.375 140.87 120.29 ;
      RECT  142.85 119.375 143.06 119.705 ;
      RECT  141.05 120.29 141.23 121.995 ;
      RECT  141.05 119.375 141.23 120.29 ;
      RECT  139.73 120.085 139.94 120.29 ;
      RECT  142.85 119.705 143.06 120.085 ;
      RECT  141.77 120.29 141.95 121.995 ;
      RECT  139.94 120.085 140.15 120.29 ;
      RECT  139.73 119.705 139.94 120.085 ;
      POLYGON  142.34 121.37 142.34 121.78 142.595 121.78 142.595 121.45 142.515 121.37 142.34 121.37 ;
      RECT  140.33 119.375 140.51 120.29 ;
      RECT  139.94 119.375 140.15 119.705 ;
      RECT  139.94 119.705 140.15 120.085 ;
      RECT  142.13 123.36 142.34 122.95 ;
      RECT  139.73 124.365 139.94 124.035 ;
      RECT  142.775 123.45 142.85 121.745 ;
      RECT  142.69 122.865 142.775 122.455 ;
      RECT  141.77 124.365 141.95 123.45 ;
      POLYGON  142.775 124.365 142.775 124.035 142.34 124.035 142.34 123.655 142.775 123.655 142.775 123.45 142.85 123.45 142.85 124.365 142.775 124.365 ;
      RECT  142.85 123.45 143.06 121.745 ;
      POLYGON  142.34 123.36 142.34 122.95 142.515 122.95 142.595 123.03 142.595 123.36 142.34 123.36 ;
      RECT  139.73 123.45 139.94 121.745 ;
      RECT  141.41 124.365 141.59 123.45 ;
      RECT  140.33 123.45 140.51 121.745 ;
      RECT  142.13 122.37 142.34 121.96 ;
      RECT  142.85 123.655 143.06 123.45 ;
      RECT  139.94 123.45 140.15 121.745 ;
      RECT  142.13 124.035 142.34 123.655 ;
      RECT  140.69 123.45 140.87 121.745 ;
      RECT  141.41 123.45 141.59 121.745 ;
      RECT  140.69 124.365 140.87 123.45 ;
      RECT  142.85 124.365 143.06 124.035 ;
      RECT  141.05 123.45 141.23 121.745 ;
      RECT  141.05 124.365 141.23 123.45 ;
      RECT  139.73 123.655 139.94 123.45 ;
      RECT  142.85 124.035 143.06 123.655 ;
      RECT  141.77 123.45 141.95 121.745 ;
      RECT  139.94 123.655 140.15 123.45 ;
      RECT  139.73 124.035 139.94 123.655 ;
      POLYGON  142.34 122.37 142.34 121.96 142.595 121.96 142.595 122.29 142.515 122.37 142.34 122.37 ;
      RECT  140.33 124.365 140.51 123.45 ;
      RECT  139.94 124.365 140.15 124.035 ;
      RECT  139.94 124.035 140.15 123.655 ;
      RECT  143.99 92.73 143.78 93.14 ;
      RECT  146.39 91.725 146.18 92.055 ;
      RECT  143.345 92.64 143.27 94.345 ;
      RECT  143.43 93.225 143.345 93.635 ;
      RECT  144.35 91.725 144.17 92.64 ;
      POLYGON  143.345 91.725 143.345 92.055 143.78 92.055 143.78 92.435 143.345 92.435 143.345 92.64 143.27 92.64 143.27 91.725 143.345 91.725 ;
      RECT  143.27 92.64 143.06 94.345 ;
      POLYGON  143.78 92.73 143.78 93.14 143.605 93.14 143.525 93.06 143.525 92.73 143.78 92.73 ;
      RECT  146.39 92.64 146.18 94.345 ;
      RECT  144.71 91.725 144.53 92.64 ;
      RECT  145.79 92.64 145.61 94.345 ;
      RECT  143.99 93.72 143.78 94.13 ;
      RECT  143.27 92.435 143.06 92.64 ;
      RECT  146.18 92.64 145.97 94.345 ;
      RECT  143.99 92.055 143.78 92.435 ;
      RECT  145.43 92.64 145.25 94.345 ;
      RECT  144.71 92.64 144.53 94.345 ;
      RECT  145.43 91.725 145.25 92.64 ;
      RECT  143.27 91.725 143.06 92.055 ;
      RECT  145.07 92.64 144.89 94.345 ;
      RECT  145.07 91.725 144.89 92.64 ;
      RECT  146.39 92.435 146.18 92.64 ;
      RECT  143.27 92.055 143.06 92.435 ;
      RECT  144.35 92.64 144.17 94.345 ;
      RECT  146.18 92.435 145.97 92.64 ;
      RECT  146.39 92.055 146.18 92.435 ;
      POLYGON  143.78 93.72 143.78 94.13 143.525 94.13 143.525 93.8 143.605 93.72 143.78 93.72 ;
      RECT  145.79 91.725 145.61 92.64 ;
      RECT  146.18 91.725 145.97 92.055 ;
      RECT  146.18 92.055 145.97 92.435 ;
      RECT  143.99 95.71 143.78 95.3 ;
      RECT  146.39 96.715 146.18 96.385 ;
      RECT  143.345 95.8 143.27 94.095 ;
      RECT  143.43 95.215 143.345 94.805 ;
      RECT  144.35 96.715 144.17 95.8 ;
      POLYGON  143.345 96.715 143.345 96.385 143.78 96.385 143.78 96.005 143.345 96.005 143.345 95.8 143.27 95.8 143.27 96.715 143.345 96.715 ;
      RECT  143.27 95.8 143.06 94.095 ;
      POLYGON  143.78 95.71 143.78 95.3 143.605 95.3 143.525 95.38 143.525 95.71 143.78 95.71 ;
      RECT  146.39 95.8 146.18 94.095 ;
      RECT  144.71 96.715 144.53 95.8 ;
      RECT  145.79 95.8 145.61 94.095 ;
      RECT  143.99 94.72 143.78 94.31 ;
      RECT  143.27 96.005 143.06 95.8 ;
      RECT  146.18 95.8 145.97 94.095 ;
      RECT  143.99 96.385 143.78 96.005 ;
      RECT  145.43 95.8 145.25 94.095 ;
      RECT  144.71 95.8 144.53 94.095 ;
      RECT  145.43 96.715 145.25 95.8 ;
      RECT  143.27 96.715 143.06 96.385 ;
      RECT  145.07 95.8 144.89 94.095 ;
      RECT  145.07 96.715 144.89 95.8 ;
      RECT  146.39 96.005 146.18 95.8 ;
      RECT  143.27 96.385 143.06 96.005 ;
      RECT  144.35 95.8 144.17 94.095 ;
      RECT  146.18 96.005 145.97 95.8 ;
      RECT  146.39 96.385 146.18 96.005 ;
      POLYGON  143.78 94.72 143.78 94.31 143.525 94.31 143.525 94.64 143.605 94.72 143.78 94.72 ;
      RECT  145.79 96.715 145.61 95.8 ;
      RECT  146.18 96.715 145.97 96.385 ;
      RECT  146.18 96.385 145.97 96.005 ;
      RECT  143.99 96.68 143.78 97.09 ;
      RECT  146.39 95.675 146.18 96.005 ;
      RECT  143.345 96.59 143.27 98.295 ;
      RECT  143.43 97.175 143.345 97.585 ;
      RECT  144.35 95.675 144.17 96.59 ;
      POLYGON  143.345 95.675 143.345 96.005 143.78 96.005 143.78 96.385 143.345 96.385 143.345 96.59 143.27 96.59 143.27 95.675 143.345 95.675 ;
      RECT  143.27 96.59 143.06 98.295 ;
      POLYGON  143.78 96.68 143.78 97.09 143.605 97.09 143.525 97.01 143.525 96.68 143.78 96.68 ;
      RECT  146.39 96.59 146.18 98.295 ;
      RECT  144.71 95.675 144.53 96.59 ;
      RECT  145.79 96.59 145.61 98.295 ;
      RECT  143.99 97.67 143.78 98.08 ;
      RECT  143.27 96.385 143.06 96.59 ;
      RECT  146.18 96.59 145.97 98.295 ;
      RECT  143.99 96.005 143.78 96.385 ;
      RECT  145.43 96.59 145.25 98.295 ;
      RECT  144.71 96.59 144.53 98.295 ;
      RECT  145.43 95.675 145.25 96.59 ;
      RECT  143.27 95.675 143.06 96.005 ;
      RECT  145.07 96.59 144.89 98.295 ;
      RECT  145.07 95.675 144.89 96.59 ;
      RECT  146.39 96.385 146.18 96.59 ;
      RECT  143.27 96.005 143.06 96.385 ;
      RECT  144.35 96.59 144.17 98.295 ;
      RECT  146.18 96.385 145.97 96.59 ;
      RECT  146.39 96.005 146.18 96.385 ;
      POLYGON  143.78 97.67 143.78 98.08 143.525 98.08 143.525 97.75 143.605 97.67 143.78 97.67 ;
      RECT  145.79 95.675 145.61 96.59 ;
      RECT  146.18 95.675 145.97 96.005 ;
      RECT  146.18 96.005 145.97 96.385 ;
      RECT  143.99 99.66 143.78 99.25 ;
      RECT  146.39 100.665 146.18 100.335 ;
      RECT  143.345 99.75 143.27 98.045 ;
      RECT  143.43 99.165 143.345 98.755 ;
      RECT  144.35 100.665 144.17 99.75 ;
      POLYGON  143.345 100.665 143.345 100.335 143.78 100.335 143.78 99.955 143.345 99.955 143.345 99.75 143.27 99.75 143.27 100.665 143.345 100.665 ;
      RECT  143.27 99.75 143.06 98.045 ;
      POLYGON  143.78 99.66 143.78 99.25 143.605 99.25 143.525 99.33 143.525 99.66 143.78 99.66 ;
      RECT  146.39 99.75 146.18 98.045 ;
      RECT  144.71 100.665 144.53 99.75 ;
      RECT  145.79 99.75 145.61 98.045 ;
      RECT  143.99 98.67 143.78 98.26 ;
      RECT  143.27 99.955 143.06 99.75 ;
      RECT  146.18 99.75 145.97 98.045 ;
      RECT  143.99 100.335 143.78 99.955 ;
      RECT  145.43 99.75 145.25 98.045 ;
      RECT  144.71 99.75 144.53 98.045 ;
      RECT  145.43 100.665 145.25 99.75 ;
      RECT  143.27 100.665 143.06 100.335 ;
      RECT  145.07 99.75 144.89 98.045 ;
      RECT  145.07 100.665 144.89 99.75 ;
      RECT  146.39 99.955 146.18 99.75 ;
      RECT  143.27 100.335 143.06 99.955 ;
      RECT  144.35 99.75 144.17 98.045 ;
      RECT  146.18 99.955 145.97 99.75 ;
      RECT  146.39 100.335 146.18 99.955 ;
      POLYGON  143.78 98.67 143.78 98.26 143.525 98.26 143.525 98.59 143.605 98.67 143.78 98.67 ;
      RECT  145.79 100.665 145.61 99.75 ;
      RECT  146.18 100.665 145.97 100.335 ;
      RECT  146.18 100.335 145.97 99.955 ;
      RECT  143.99 100.63 143.78 101.04 ;
      RECT  146.39 99.625 146.18 99.955 ;
      RECT  143.345 100.54 143.27 102.245 ;
      RECT  143.43 101.125 143.345 101.535 ;
      RECT  144.35 99.625 144.17 100.54 ;
      POLYGON  143.345 99.625 143.345 99.955 143.78 99.955 143.78 100.335 143.345 100.335 143.345 100.54 143.27 100.54 143.27 99.625 143.345 99.625 ;
      RECT  143.27 100.54 143.06 102.245 ;
      POLYGON  143.78 100.63 143.78 101.04 143.605 101.04 143.525 100.96 143.525 100.63 143.78 100.63 ;
      RECT  146.39 100.54 146.18 102.245 ;
      RECT  144.71 99.625 144.53 100.54 ;
      RECT  145.79 100.54 145.61 102.245 ;
      RECT  143.99 101.62 143.78 102.03 ;
      RECT  143.27 100.335 143.06 100.54 ;
      RECT  146.18 100.54 145.97 102.245 ;
      RECT  143.99 99.955 143.78 100.335 ;
      RECT  145.43 100.54 145.25 102.245 ;
      RECT  144.71 100.54 144.53 102.245 ;
      RECT  145.43 99.625 145.25 100.54 ;
      RECT  143.27 99.625 143.06 99.955 ;
      RECT  145.07 100.54 144.89 102.245 ;
      RECT  145.07 99.625 144.89 100.54 ;
      RECT  146.39 100.335 146.18 100.54 ;
      RECT  143.27 99.955 143.06 100.335 ;
      RECT  144.35 100.54 144.17 102.245 ;
      RECT  146.18 100.335 145.97 100.54 ;
      RECT  146.39 99.955 146.18 100.335 ;
      POLYGON  143.78 101.62 143.78 102.03 143.525 102.03 143.525 101.7 143.605 101.62 143.78 101.62 ;
      RECT  145.79 99.625 145.61 100.54 ;
      RECT  146.18 99.625 145.97 99.955 ;
      RECT  146.18 99.955 145.97 100.335 ;
      RECT  143.99 103.61 143.78 103.2 ;
      RECT  146.39 104.615 146.18 104.285 ;
      RECT  143.345 103.7 143.27 101.995 ;
      RECT  143.43 103.115 143.345 102.705 ;
      RECT  144.35 104.615 144.17 103.7 ;
      POLYGON  143.345 104.615 143.345 104.285 143.78 104.285 143.78 103.905 143.345 103.905 143.345 103.7 143.27 103.7 143.27 104.615 143.345 104.615 ;
      RECT  143.27 103.7 143.06 101.995 ;
      POLYGON  143.78 103.61 143.78 103.2 143.605 103.2 143.525 103.28 143.525 103.61 143.78 103.61 ;
      RECT  146.39 103.7 146.18 101.995 ;
      RECT  144.71 104.615 144.53 103.7 ;
      RECT  145.79 103.7 145.61 101.995 ;
      RECT  143.99 102.62 143.78 102.21 ;
      RECT  143.27 103.905 143.06 103.7 ;
      RECT  146.18 103.7 145.97 101.995 ;
      RECT  143.99 104.285 143.78 103.905 ;
      RECT  145.43 103.7 145.25 101.995 ;
      RECT  144.71 103.7 144.53 101.995 ;
      RECT  145.43 104.615 145.25 103.7 ;
      RECT  143.27 104.615 143.06 104.285 ;
      RECT  145.07 103.7 144.89 101.995 ;
      RECT  145.07 104.615 144.89 103.7 ;
      RECT  146.39 103.905 146.18 103.7 ;
      RECT  143.27 104.285 143.06 103.905 ;
      RECT  144.35 103.7 144.17 101.995 ;
      RECT  146.18 103.905 145.97 103.7 ;
      RECT  146.39 104.285 146.18 103.905 ;
      POLYGON  143.78 102.62 143.78 102.21 143.525 102.21 143.525 102.54 143.605 102.62 143.78 102.62 ;
      RECT  145.79 104.615 145.61 103.7 ;
      RECT  146.18 104.615 145.97 104.285 ;
      RECT  146.18 104.285 145.97 103.905 ;
      RECT  143.99 104.58 143.78 104.99 ;
      RECT  146.39 103.575 146.18 103.905 ;
      RECT  143.345 104.49 143.27 106.195 ;
      RECT  143.43 105.075 143.345 105.485 ;
      RECT  144.35 103.575 144.17 104.49 ;
      POLYGON  143.345 103.575 143.345 103.905 143.78 103.905 143.78 104.285 143.345 104.285 143.345 104.49 143.27 104.49 143.27 103.575 143.345 103.575 ;
      RECT  143.27 104.49 143.06 106.195 ;
      POLYGON  143.78 104.58 143.78 104.99 143.605 104.99 143.525 104.91 143.525 104.58 143.78 104.58 ;
      RECT  146.39 104.49 146.18 106.195 ;
      RECT  144.71 103.575 144.53 104.49 ;
      RECT  145.79 104.49 145.61 106.195 ;
      RECT  143.99 105.57 143.78 105.98 ;
      RECT  143.27 104.285 143.06 104.49 ;
      RECT  146.18 104.49 145.97 106.195 ;
      RECT  143.99 103.905 143.78 104.285 ;
      RECT  145.43 104.49 145.25 106.195 ;
      RECT  144.71 104.49 144.53 106.195 ;
      RECT  145.43 103.575 145.25 104.49 ;
      RECT  143.27 103.575 143.06 103.905 ;
      RECT  145.07 104.49 144.89 106.195 ;
      RECT  145.07 103.575 144.89 104.49 ;
      RECT  146.39 104.285 146.18 104.49 ;
      RECT  143.27 103.905 143.06 104.285 ;
      RECT  144.35 104.49 144.17 106.195 ;
      RECT  146.18 104.285 145.97 104.49 ;
      RECT  146.39 103.905 146.18 104.285 ;
      POLYGON  143.78 105.57 143.78 105.98 143.525 105.98 143.525 105.65 143.605 105.57 143.78 105.57 ;
      RECT  145.79 103.575 145.61 104.49 ;
      RECT  146.18 103.575 145.97 103.905 ;
      RECT  146.18 103.905 145.97 104.285 ;
      RECT  143.99 107.56 143.78 107.15 ;
      RECT  146.39 108.565 146.18 108.235 ;
      RECT  143.345 107.65 143.27 105.945 ;
      RECT  143.43 107.065 143.345 106.655 ;
      RECT  144.35 108.565 144.17 107.65 ;
      POLYGON  143.345 108.565 143.345 108.235 143.78 108.235 143.78 107.855 143.345 107.855 143.345 107.65 143.27 107.65 143.27 108.565 143.345 108.565 ;
      RECT  143.27 107.65 143.06 105.945 ;
      POLYGON  143.78 107.56 143.78 107.15 143.605 107.15 143.525 107.23 143.525 107.56 143.78 107.56 ;
      RECT  146.39 107.65 146.18 105.945 ;
      RECT  144.71 108.565 144.53 107.65 ;
      RECT  145.79 107.65 145.61 105.945 ;
      RECT  143.99 106.57 143.78 106.16 ;
      RECT  143.27 107.855 143.06 107.65 ;
      RECT  146.18 107.65 145.97 105.945 ;
      RECT  143.99 108.235 143.78 107.855 ;
      RECT  145.43 107.65 145.25 105.945 ;
      RECT  144.71 107.65 144.53 105.945 ;
      RECT  145.43 108.565 145.25 107.65 ;
      RECT  143.27 108.565 143.06 108.235 ;
      RECT  145.07 107.65 144.89 105.945 ;
      RECT  145.07 108.565 144.89 107.65 ;
      RECT  146.39 107.855 146.18 107.65 ;
      RECT  143.27 108.235 143.06 107.855 ;
      RECT  144.35 107.65 144.17 105.945 ;
      RECT  146.18 107.855 145.97 107.65 ;
      RECT  146.39 108.235 146.18 107.855 ;
      POLYGON  143.78 106.57 143.78 106.16 143.525 106.16 143.525 106.49 143.605 106.57 143.78 106.57 ;
      RECT  145.79 108.565 145.61 107.65 ;
      RECT  146.18 108.565 145.97 108.235 ;
      RECT  146.18 108.235 145.97 107.855 ;
      RECT  143.99 108.53 143.78 108.94 ;
      RECT  146.39 107.525 146.18 107.855 ;
      RECT  143.345 108.44 143.27 110.145 ;
      RECT  143.43 109.025 143.345 109.435 ;
      RECT  144.35 107.525 144.17 108.44 ;
      POLYGON  143.345 107.525 143.345 107.855 143.78 107.855 143.78 108.235 143.345 108.235 143.345 108.44 143.27 108.44 143.27 107.525 143.345 107.525 ;
      RECT  143.27 108.44 143.06 110.145 ;
      POLYGON  143.78 108.53 143.78 108.94 143.605 108.94 143.525 108.86 143.525 108.53 143.78 108.53 ;
      RECT  146.39 108.44 146.18 110.145 ;
      RECT  144.71 107.525 144.53 108.44 ;
      RECT  145.79 108.44 145.61 110.145 ;
      RECT  143.99 109.52 143.78 109.93 ;
      RECT  143.27 108.235 143.06 108.44 ;
      RECT  146.18 108.44 145.97 110.145 ;
      RECT  143.99 107.855 143.78 108.235 ;
      RECT  145.43 108.44 145.25 110.145 ;
      RECT  144.71 108.44 144.53 110.145 ;
      RECT  145.43 107.525 145.25 108.44 ;
      RECT  143.27 107.525 143.06 107.855 ;
      RECT  145.07 108.44 144.89 110.145 ;
      RECT  145.07 107.525 144.89 108.44 ;
      RECT  146.39 108.235 146.18 108.44 ;
      RECT  143.27 107.855 143.06 108.235 ;
      RECT  144.35 108.44 144.17 110.145 ;
      RECT  146.18 108.235 145.97 108.44 ;
      RECT  146.39 107.855 146.18 108.235 ;
      POLYGON  143.78 109.52 143.78 109.93 143.525 109.93 143.525 109.6 143.605 109.52 143.78 109.52 ;
      RECT  145.79 107.525 145.61 108.44 ;
      RECT  146.18 107.525 145.97 107.855 ;
      RECT  146.18 107.855 145.97 108.235 ;
      RECT  143.99 111.51 143.78 111.1 ;
      RECT  146.39 112.515 146.18 112.185 ;
      RECT  143.345 111.6 143.27 109.895 ;
      RECT  143.43 111.015 143.345 110.605 ;
      RECT  144.35 112.515 144.17 111.6 ;
      POLYGON  143.345 112.515 143.345 112.185 143.78 112.185 143.78 111.805 143.345 111.805 143.345 111.6 143.27 111.6 143.27 112.515 143.345 112.515 ;
      RECT  143.27 111.6 143.06 109.895 ;
      POLYGON  143.78 111.51 143.78 111.1 143.605 111.1 143.525 111.18 143.525 111.51 143.78 111.51 ;
      RECT  146.39 111.6 146.18 109.895 ;
      RECT  144.71 112.515 144.53 111.6 ;
      RECT  145.79 111.6 145.61 109.895 ;
      RECT  143.99 110.52 143.78 110.11 ;
      RECT  143.27 111.805 143.06 111.6 ;
      RECT  146.18 111.6 145.97 109.895 ;
      RECT  143.99 112.185 143.78 111.805 ;
      RECT  145.43 111.6 145.25 109.895 ;
      RECT  144.71 111.6 144.53 109.895 ;
      RECT  145.43 112.515 145.25 111.6 ;
      RECT  143.27 112.515 143.06 112.185 ;
      RECT  145.07 111.6 144.89 109.895 ;
      RECT  145.07 112.515 144.89 111.6 ;
      RECT  146.39 111.805 146.18 111.6 ;
      RECT  143.27 112.185 143.06 111.805 ;
      RECT  144.35 111.6 144.17 109.895 ;
      RECT  146.18 111.805 145.97 111.6 ;
      RECT  146.39 112.185 146.18 111.805 ;
      POLYGON  143.78 110.52 143.78 110.11 143.525 110.11 143.525 110.44 143.605 110.52 143.78 110.52 ;
      RECT  145.79 112.515 145.61 111.6 ;
      RECT  146.18 112.515 145.97 112.185 ;
      RECT  146.18 112.185 145.97 111.805 ;
      RECT  143.99 112.48 143.78 112.89 ;
      RECT  146.39 111.475 146.18 111.805 ;
      RECT  143.345 112.39 143.27 114.095 ;
      RECT  143.43 112.975 143.345 113.385 ;
      RECT  144.35 111.475 144.17 112.39 ;
      POLYGON  143.345 111.475 143.345 111.805 143.78 111.805 143.78 112.185 143.345 112.185 143.345 112.39 143.27 112.39 143.27 111.475 143.345 111.475 ;
      RECT  143.27 112.39 143.06 114.095 ;
      POLYGON  143.78 112.48 143.78 112.89 143.605 112.89 143.525 112.81 143.525 112.48 143.78 112.48 ;
      RECT  146.39 112.39 146.18 114.095 ;
      RECT  144.71 111.475 144.53 112.39 ;
      RECT  145.79 112.39 145.61 114.095 ;
      RECT  143.99 113.47 143.78 113.88 ;
      RECT  143.27 112.185 143.06 112.39 ;
      RECT  146.18 112.39 145.97 114.095 ;
      RECT  143.99 111.805 143.78 112.185 ;
      RECT  145.43 112.39 145.25 114.095 ;
      RECT  144.71 112.39 144.53 114.095 ;
      RECT  145.43 111.475 145.25 112.39 ;
      RECT  143.27 111.475 143.06 111.805 ;
      RECT  145.07 112.39 144.89 114.095 ;
      RECT  145.07 111.475 144.89 112.39 ;
      RECT  146.39 112.185 146.18 112.39 ;
      RECT  143.27 111.805 143.06 112.185 ;
      RECT  144.35 112.39 144.17 114.095 ;
      RECT  146.18 112.185 145.97 112.39 ;
      RECT  146.39 111.805 146.18 112.185 ;
      POLYGON  143.78 113.47 143.78 113.88 143.525 113.88 143.525 113.55 143.605 113.47 143.78 113.47 ;
      RECT  145.79 111.475 145.61 112.39 ;
      RECT  146.18 111.475 145.97 111.805 ;
      RECT  146.18 111.805 145.97 112.185 ;
      RECT  143.99 115.46 143.78 115.05 ;
      RECT  146.39 116.465 146.18 116.135 ;
      RECT  143.345 115.55 143.27 113.845 ;
      RECT  143.43 114.965 143.345 114.555 ;
      RECT  144.35 116.465 144.17 115.55 ;
      POLYGON  143.345 116.465 143.345 116.135 143.78 116.135 143.78 115.755 143.345 115.755 143.345 115.55 143.27 115.55 143.27 116.465 143.345 116.465 ;
      RECT  143.27 115.55 143.06 113.845 ;
      POLYGON  143.78 115.46 143.78 115.05 143.605 115.05 143.525 115.13 143.525 115.46 143.78 115.46 ;
      RECT  146.39 115.55 146.18 113.845 ;
      RECT  144.71 116.465 144.53 115.55 ;
      RECT  145.79 115.55 145.61 113.845 ;
      RECT  143.99 114.47 143.78 114.06 ;
      RECT  143.27 115.755 143.06 115.55 ;
      RECT  146.18 115.55 145.97 113.845 ;
      RECT  143.99 116.135 143.78 115.755 ;
      RECT  145.43 115.55 145.25 113.845 ;
      RECT  144.71 115.55 144.53 113.845 ;
      RECT  145.43 116.465 145.25 115.55 ;
      RECT  143.27 116.465 143.06 116.135 ;
      RECT  145.07 115.55 144.89 113.845 ;
      RECT  145.07 116.465 144.89 115.55 ;
      RECT  146.39 115.755 146.18 115.55 ;
      RECT  143.27 116.135 143.06 115.755 ;
      RECT  144.35 115.55 144.17 113.845 ;
      RECT  146.18 115.755 145.97 115.55 ;
      RECT  146.39 116.135 146.18 115.755 ;
      POLYGON  143.78 114.47 143.78 114.06 143.525 114.06 143.525 114.39 143.605 114.47 143.78 114.47 ;
      RECT  145.79 116.465 145.61 115.55 ;
      RECT  146.18 116.465 145.97 116.135 ;
      RECT  146.18 116.135 145.97 115.755 ;
      RECT  143.99 116.43 143.78 116.84 ;
      RECT  146.39 115.425 146.18 115.755 ;
      RECT  143.345 116.34 143.27 118.045 ;
      RECT  143.43 116.925 143.345 117.335 ;
      RECT  144.35 115.425 144.17 116.34 ;
      POLYGON  143.345 115.425 143.345 115.755 143.78 115.755 143.78 116.135 143.345 116.135 143.345 116.34 143.27 116.34 143.27 115.425 143.345 115.425 ;
      RECT  143.27 116.34 143.06 118.045 ;
      POLYGON  143.78 116.43 143.78 116.84 143.605 116.84 143.525 116.76 143.525 116.43 143.78 116.43 ;
      RECT  146.39 116.34 146.18 118.045 ;
      RECT  144.71 115.425 144.53 116.34 ;
      RECT  145.79 116.34 145.61 118.045 ;
      RECT  143.99 117.42 143.78 117.83 ;
      RECT  143.27 116.135 143.06 116.34 ;
      RECT  146.18 116.34 145.97 118.045 ;
      RECT  143.99 115.755 143.78 116.135 ;
      RECT  145.43 116.34 145.25 118.045 ;
      RECT  144.71 116.34 144.53 118.045 ;
      RECT  145.43 115.425 145.25 116.34 ;
      RECT  143.27 115.425 143.06 115.755 ;
      RECT  145.07 116.34 144.89 118.045 ;
      RECT  145.07 115.425 144.89 116.34 ;
      RECT  146.39 116.135 146.18 116.34 ;
      RECT  143.27 115.755 143.06 116.135 ;
      RECT  144.35 116.34 144.17 118.045 ;
      RECT  146.18 116.135 145.97 116.34 ;
      RECT  146.39 115.755 146.18 116.135 ;
      POLYGON  143.78 117.42 143.78 117.83 143.525 117.83 143.525 117.5 143.605 117.42 143.78 117.42 ;
      RECT  145.79 115.425 145.61 116.34 ;
      RECT  146.18 115.425 145.97 115.755 ;
      RECT  146.18 115.755 145.97 116.135 ;
      RECT  143.99 119.41 143.78 119.0 ;
      RECT  146.39 120.415 146.18 120.085 ;
      RECT  143.345 119.5 143.27 117.795 ;
      RECT  143.43 118.915 143.345 118.505 ;
      RECT  144.35 120.415 144.17 119.5 ;
      POLYGON  143.345 120.415 143.345 120.085 143.78 120.085 143.78 119.705 143.345 119.705 143.345 119.5 143.27 119.5 143.27 120.415 143.345 120.415 ;
      RECT  143.27 119.5 143.06 117.795 ;
      POLYGON  143.78 119.41 143.78 119.0 143.605 119.0 143.525 119.08 143.525 119.41 143.78 119.41 ;
      RECT  146.39 119.5 146.18 117.795 ;
      RECT  144.71 120.415 144.53 119.5 ;
      RECT  145.79 119.5 145.61 117.795 ;
      RECT  143.99 118.42 143.78 118.01 ;
      RECT  143.27 119.705 143.06 119.5 ;
      RECT  146.18 119.5 145.97 117.795 ;
      RECT  143.99 120.085 143.78 119.705 ;
      RECT  145.43 119.5 145.25 117.795 ;
      RECT  144.71 119.5 144.53 117.795 ;
      RECT  145.43 120.415 145.25 119.5 ;
      RECT  143.27 120.415 143.06 120.085 ;
      RECT  145.07 119.5 144.89 117.795 ;
      RECT  145.07 120.415 144.89 119.5 ;
      RECT  146.39 119.705 146.18 119.5 ;
      RECT  143.27 120.085 143.06 119.705 ;
      RECT  144.35 119.5 144.17 117.795 ;
      RECT  146.18 119.705 145.97 119.5 ;
      RECT  146.39 120.085 146.18 119.705 ;
      POLYGON  143.78 118.42 143.78 118.01 143.525 118.01 143.525 118.34 143.605 118.42 143.78 118.42 ;
      RECT  145.79 120.415 145.61 119.5 ;
      RECT  146.18 120.415 145.97 120.085 ;
      RECT  146.18 120.085 145.97 119.705 ;
      RECT  143.99 120.38 143.78 120.79 ;
      RECT  146.39 119.375 146.18 119.705 ;
      RECT  143.345 120.29 143.27 121.995 ;
      RECT  143.43 120.875 143.345 121.285 ;
      RECT  144.35 119.375 144.17 120.29 ;
      POLYGON  143.345 119.375 143.345 119.705 143.78 119.705 143.78 120.085 143.345 120.085 143.345 120.29 143.27 120.29 143.27 119.375 143.345 119.375 ;
      RECT  143.27 120.29 143.06 121.995 ;
      POLYGON  143.78 120.38 143.78 120.79 143.605 120.79 143.525 120.71 143.525 120.38 143.78 120.38 ;
      RECT  146.39 120.29 146.18 121.995 ;
      RECT  144.71 119.375 144.53 120.29 ;
      RECT  145.79 120.29 145.61 121.995 ;
      RECT  143.99 121.37 143.78 121.78 ;
      RECT  143.27 120.085 143.06 120.29 ;
      RECT  146.18 120.29 145.97 121.995 ;
      RECT  143.99 119.705 143.78 120.085 ;
      RECT  145.43 120.29 145.25 121.995 ;
      RECT  144.71 120.29 144.53 121.995 ;
      RECT  145.43 119.375 145.25 120.29 ;
      RECT  143.27 119.375 143.06 119.705 ;
      RECT  145.07 120.29 144.89 121.995 ;
      RECT  145.07 119.375 144.89 120.29 ;
      RECT  146.39 120.085 146.18 120.29 ;
      RECT  143.27 119.705 143.06 120.085 ;
      RECT  144.35 120.29 144.17 121.995 ;
      RECT  146.18 120.085 145.97 120.29 ;
      RECT  146.39 119.705 146.18 120.085 ;
      POLYGON  143.78 121.37 143.78 121.78 143.525 121.78 143.525 121.45 143.605 121.37 143.78 121.37 ;
      RECT  145.79 119.375 145.61 120.29 ;
      RECT  146.18 119.375 145.97 119.705 ;
      RECT  146.18 119.705 145.97 120.085 ;
      RECT  143.99 123.36 143.78 122.95 ;
      RECT  146.39 124.365 146.18 124.035 ;
      RECT  143.345 123.45 143.27 121.745 ;
      RECT  143.43 122.865 143.345 122.455 ;
      RECT  144.35 124.365 144.17 123.45 ;
      POLYGON  143.345 124.365 143.345 124.035 143.78 124.035 143.78 123.655 143.345 123.655 143.345 123.45 143.27 123.45 143.27 124.365 143.345 124.365 ;
      RECT  143.27 123.45 143.06 121.745 ;
      POLYGON  143.78 123.36 143.78 122.95 143.605 122.95 143.525 123.03 143.525 123.36 143.78 123.36 ;
      RECT  146.39 123.45 146.18 121.745 ;
      RECT  144.71 124.365 144.53 123.45 ;
      RECT  145.79 123.45 145.61 121.745 ;
      RECT  143.99 122.37 143.78 121.96 ;
      RECT  143.27 123.655 143.06 123.45 ;
      RECT  146.18 123.45 145.97 121.745 ;
      RECT  143.99 124.035 143.78 123.655 ;
      RECT  145.43 123.45 145.25 121.745 ;
      RECT  144.71 123.45 144.53 121.745 ;
      RECT  145.43 124.365 145.25 123.45 ;
      RECT  143.27 124.365 143.06 124.035 ;
      RECT  145.07 123.45 144.89 121.745 ;
      RECT  145.07 124.365 144.89 123.45 ;
      RECT  146.39 123.655 146.18 123.45 ;
      RECT  143.27 124.035 143.06 123.655 ;
      RECT  144.35 123.45 144.17 121.745 ;
      RECT  146.18 123.655 145.97 123.45 ;
      RECT  146.39 124.035 146.18 123.655 ;
      POLYGON  143.78 122.37 143.78 121.96 143.525 121.96 143.525 122.29 143.605 122.37 143.78 122.37 ;
      RECT  145.79 124.365 145.61 123.45 ;
      RECT  146.18 124.365 145.97 124.035 ;
      RECT  146.18 124.035 145.97 123.655 ;
      RECT  96.65 92.245 96.83 123.845 ;
      RECT  97.01 92.245 97.19 123.845 ;
      RECT  97.73 92.245 97.91 123.845 ;
      RECT  98.09 92.245 98.27 123.845 ;
      RECT  101.93 92.245 102.11 123.845 ;
      RECT  101.57 92.245 101.75 123.845 ;
      RECT  100.85 92.245 101.03 123.845 ;
      RECT  100.49 92.245 100.67 123.845 ;
      RECT  102.89 92.245 103.07 123.845 ;
      RECT  103.25 92.245 103.43 123.845 ;
      RECT  103.97 92.245 104.15 123.845 ;
      RECT  104.33 92.245 104.51 123.845 ;
      RECT  108.17 92.245 108.35 123.845 ;
      RECT  107.81 92.245 107.99 123.845 ;
      RECT  107.09 92.245 107.27 123.845 ;
      RECT  106.73 92.245 106.91 123.845 ;
      RECT  109.13 92.245 109.31 123.845 ;
      RECT  109.49 92.245 109.67 123.845 ;
      RECT  110.21 92.245 110.39 123.845 ;
      RECT  110.57 92.245 110.75 123.845 ;
      RECT  114.41 92.245 114.59 123.845 ;
      RECT  114.05 92.245 114.23 123.845 ;
      RECT  113.33 92.245 113.51 123.845 ;
      RECT  112.97 92.245 113.15 123.845 ;
      RECT  115.37 92.245 115.55 123.845 ;
      RECT  115.73 92.245 115.91 123.845 ;
      RECT  116.45 92.245 116.63 123.845 ;
      RECT  116.81 92.245 116.99 123.845 ;
      RECT  120.65 92.245 120.83 123.845 ;
      RECT  120.29 92.245 120.47 123.845 ;
      RECT  119.57 92.245 119.75 123.845 ;
      RECT  119.21 92.245 119.39 123.845 ;
      RECT  121.61 92.245 121.79 123.845 ;
      RECT  121.97 92.245 122.15 123.845 ;
      RECT  122.69 92.245 122.87 123.845 ;
      RECT  123.05 92.245 123.23 123.845 ;
      RECT  126.89 92.245 127.07 123.845 ;
      RECT  126.53 92.245 126.71 123.845 ;
      RECT  125.81 92.245 125.99 123.845 ;
      RECT  125.45 92.245 125.63 123.845 ;
      RECT  127.85 92.245 128.03 123.845 ;
      RECT  128.21 92.245 128.39 123.845 ;
      RECT  128.93 92.245 129.11 123.845 ;
      RECT  129.29 92.245 129.47 123.845 ;
      RECT  133.13 92.245 133.31 123.845 ;
      RECT  132.77 92.245 132.95 123.845 ;
      RECT  132.05 92.245 132.23 123.845 ;
      RECT  131.69 92.245 131.87 123.845 ;
      RECT  134.09 92.245 134.27 123.845 ;
      RECT  134.45 92.245 134.63 123.845 ;
      RECT  135.17 92.245 135.35 123.845 ;
      RECT  135.53 92.245 135.71 123.845 ;
      RECT  139.37 92.245 139.55 123.845 ;
      RECT  139.01 92.245 139.19 123.845 ;
      RECT  138.29 92.245 138.47 123.845 ;
      RECT  137.93 92.245 138.11 123.845 ;
      RECT  140.33 92.245 140.51 123.845 ;
      RECT  140.69 92.245 140.87 123.845 ;
      RECT  141.41 92.245 141.59 123.845 ;
      RECT  141.77 92.245 141.95 123.845 ;
      RECT  145.61 92.245 145.79 123.845 ;
      RECT  145.25 92.245 145.43 123.845 ;
      RECT  144.53 92.245 144.71 123.845 ;
      RECT  144.17 92.245 144.35 123.845 ;
      RECT  138.65 105.945 138.83 107.65 ;
      RECT  128.57 113.845 128.75 115.55 ;
      RECT  119.93 117.795 120.11 119.5 ;
      RECT  116.09 121.745 116.27 123.45 ;
      RECT  116.09 113.845 116.27 115.55 ;
      RECT  109.85 109.895 110.03 111.6 ;
      RECT  138.65 98.045 138.83 99.75 ;
      RECT  101.21 94.095 101.39 95.8 ;
      RECT  119.93 109.895 120.11 111.6 ;
      RECT  144.89 120.29 145.07 121.995 ;
      RECT  122.33 96.59 122.51 98.295 ;
      RECT  126.17 109.895 126.35 111.6 ;
      RECT  116.09 98.045 116.27 99.75 ;
      RECT  122.33 113.845 122.51 115.55 ;
      RECT  144.89 117.795 145.07 119.5 ;
      RECT  113.69 113.845 113.87 115.55 ;
      RECT  97.37 113.845 97.55 115.55 ;
      RECT  107.45 117.795 107.63 119.5 ;
      RECT  97.37 120.29 97.55 121.995 ;
      RECT  103.61 120.29 103.79 121.995 ;
      RECT  134.81 120.29 134.99 121.995 ;
      RECT  109.85 112.39 110.03 114.095 ;
      RECT  126.17 100.54 126.35 102.245 ;
      RECT  116.09 112.39 116.27 114.095 ;
      RECT  119.93 112.39 120.11 114.095 ;
      RECT  132.41 121.745 132.59 123.45 ;
      RECT  119.93 98.045 120.11 99.75 ;
      RECT  138.65 94.095 138.83 95.8 ;
      RECT  103.61 96.59 103.79 98.295 ;
      RECT  113.69 116.34 113.87 118.045 ;
      RECT  116.09 109.895 116.27 111.6 ;
      RECT  128.57 117.795 128.75 119.5 ;
      RECT  138.65 92.64 138.83 94.345 ;
      RECT  109.85 105.945 110.03 107.65 ;
      RECT  97.37 98.045 97.55 99.75 ;
      RECT  97.37 108.44 97.55 110.145 ;
      RECT  101.21 109.895 101.39 111.6 ;
      RECT  107.45 92.64 107.63 94.345 ;
      RECT  134.81 98.045 134.99 99.75 ;
      RECT  122.33 105.945 122.51 107.65 ;
      RECT  101.21 120.29 101.39 121.995 ;
      RECT  128.57 112.39 128.75 114.095 ;
      RECT  109.85 120.29 110.03 121.995 ;
      RECT  101.21 116.34 101.39 118.045 ;
      RECT  144.89 94.095 145.07 95.8 ;
      RECT  113.69 98.045 113.87 99.75 ;
      RECT  132.41 113.845 132.59 115.55 ;
      RECT  103.61 108.44 103.79 110.145 ;
      RECT  119.93 108.44 120.11 110.145 ;
      RECT  144.89 100.54 145.07 102.245 ;
      RECT  97.37 104.49 97.55 106.195 ;
      RECT  122.33 108.44 122.51 110.145 ;
      RECT  116.09 101.995 116.27 103.7 ;
      RECT  103.61 112.39 103.79 114.095 ;
      RECT  128.57 92.64 128.75 94.345 ;
      RECT  141.05 112.39 141.23 114.095 ;
      RECT  119.93 105.945 120.11 107.65 ;
      RECT  132.41 116.34 132.59 118.045 ;
      RECT  144.89 121.745 145.07 123.45 ;
      RECT  126.17 120.29 126.35 121.995 ;
      RECT  107.45 120.29 107.63 121.995 ;
      RECT  122.33 117.795 122.51 119.5 ;
      RECT  134.81 104.49 134.99 106.195 ;
      RECT  128.57 120.29 128.75 121.995 ;
      RECT  101.21 113.845 101.39 115.55 ;
      RECT  97.37 112.39 97.55 114.095 ;
      RECT  132.41 101.995 132.59 103.7 ;
      RECT  126.17 121.745 126.35 123.45 ;
      RECT  103.61 117.795 103.79 119.5 ;
      RECT  119.93 121.745 120.11 123.45 ;
      RECT  109.85 116.34 110.03 118.045 ;
      RECT  97.37 109.895 97.55 111.6 ;
      RECT  141.05 98.045 141.23 99.75 ;
      RECT  141.05 109.895 141.23 111.6 ;
      RECT  119.93 96.59 120.11 98.295 ;
      RECT  141.05 120.29 141.23 121.995 ;
      RECT  132.41 98.045 132.59 99.75 ;
      RECT  116.09 120.29 116.27 121.995 ;
      RECT  107.45 101.995 107.63 103.7 ;
      RECT  132.41 92.64 132.59 94.345 ;
      RECT  97.37 117.795 97.55 119.5 ;
      RECT  138.65 117.795 138.83 119.5 ;
      RECT  119.93 120.29 120.11 121.995 ;
      RECT  134.81 113.845 134.99 115.55 ;
      RECT  138.65 116.34 138.83 118.045 ;
      RECT  107.45 105.945 107.63 107.65 ;
      RECT  144.89 101.995 145.07 103.7 ;
      RECT  103.61 104.49 103.79 106.195 ;
      RECT  119.93 100.54 120.11 102.245 ;
      RECT  113.69 117.795 113.87 119.5 ;
      RECT  109.85 100.54 110.03 102.245 ;
      RECT  122.33 121.745 122.51 123.45 ;
      RECT  113.69 109.895 113.87 111.6 ;
      RECT  141.05 104.49 141.23 106.195 ;
      RECT  126.17 113.845 126.35 115.55 ;
      RECT  122.33 94.095 122.51 95.8 ;
      RECT  113.69 108.44 113.87 110.145 ;
      RECT  126.17 94.095 126.35 95.8 ;
      RECT  141.05 94.095 141.23 95.8 ;
      RECT  101.21 96.59 101.39 98.295 ;
      RECT  141.05 101.995 141.23 103.7 ;
      RECT  116.09 108.44 116.27 110.145 ;
      RECT  97.37 121.745 97.55 123.45 ;
      RECT  97.37 96.59 97.55 98.295 ;
      RECT  122.33 109.895 122.51 111.6 ;
      RECT  132.41 96.59 132.59 98.295 ;
      RECT  141.05 96.59 141.23 98.295 ;
      RECT  116.09 104.49 116.27 106.195 ;
      RECT  132.41 112.39 132.59 114.095 ;
      RECT  144.89 96.59 145.07 98.295 ;
      RECT  126.17 112.39 126.35 114.095 ;
      RECT  101.21 104.49 101.39 106.195 ;
      RECT  144.89 92.64 145.07 94.345 ;
      RECT  103.61 100.54 103.79 102.245 ;
      RECT  103.61 105.945 103.79 107.65 ;
      RECT  103.61 113.845 103.79 115.55 ;
      RECT  116.09 100.54 116.27 102.245 ;
      RECT  134.81 109.895 134.99 111.6 ;
      RECT  101.21 98.045 101.39 99.75 ;
      RECT  138.65 101.995 138.83 103.7 ;
      RECT  141.05 105.945 141.23 107.65 ;
      RECT  109.85 108.44 110.03 110.145 ;
      RECT  141.05 117.795 141.23 119.5 ;
      RECT  128.57 100.54 128.75 102.245 ;
      RECT  134.81 101.995 134.99 103.7 ;
      RECT  103.61 109.895 103.79 111.6 ;
      RECT  97.37 94.095 97.55 95.8 ;
      RECT  103.61 98.045 103.79 99.75 ;
      RECT  101.21 100.54 101.39 102.245 ;
      RECT  138.65 96.59 138.83 98.295 ;
      RECT  122.33 112.39 122.51 114.095 ;
      RECT  107.45 112.39 107.63 114.095 ;
      RECT  144.89 108.44 145.07 110.145 ;
      RECT  126.17 105.945 126.35 107.65 ;
      RECT  134.81 94.095 134.99 95.8 ;
      RECT  103.61 101.995 103.79 103.7 ;
      RECT  126.17 92.64 126.35 94.345 ;
      RECT  134.81 92.64 134.99 94.345 ;
      RECT  126.17 108.44 126.35 110.145 ;
      RECT  113.69 121.745 113.87 123.45 ;
      RECT  144.89 98.045 145.07 99.75 ;
      RECT  119.93 113.845 120.11 115.55 ;
      RECT  97.37 92.64 97.55 94.345 ;
      RECT  107.45 100.54 107.63 102.245 ;
      RECT  128.57 101.995 128.75 103.7 ;
      RECT  134.81 105.945 134.99 107.65 ;
      RECT  126.17 116.34 126.35 118.045 ;
      RECT  128.57 96.59 128.75 98.295 ;
      RECT  119.93 101.995 120.11 103.7 ;
      RECT  97.37 100.54 97.55 102.245 ;
      RECT  107.45 113.845 107.63 115.55 ;
      RECT  113.69 92.64 113.87 94.345 ;
      RECT  132.41 100.54 132.59 102.245 ;
      RECT  119.93 104.49 120.11 106.195 ;
      RECT  97.37 105.945 97.55 107.65 ;
      RECT  101.21 108.44 101.39 110.145 ;
      RECT  138.65 109.895 138.83 111.6 ;
      RECT  113.69 105.945 113.87 107.65 ;
      RECT  138.65 120.29 138.83 121.995 ;
      RECT  109.85 96.59 110.03 98.295 ;
      RECT  109.85 98.045 110.03 99.75 ;
      RECT  109.85 113.845 110.03 115.55 ;
      RECT  138.65 112.39 138.83 114.095 ;
      RECT  144.89 113.845 145.07 115.55 ;
      RECT  113.69 100.54 113.87 102.245 ;
      RECT  107.45 98.045 107.63 99.75 ;
      RECT  109.85 94.095 110.03 95.8 ;
      RECT  144.89 105.945 145.07 107.65 ;
      RECT  134.81 116.34 134.99 118.045 ;
      RECT  107.45 116.34 107.63 118.045 ;
      RECT  116.09 105.945 116.27 107.65 ;
      RECT  134.81 100.54 134.99 102.245 ;
      RECT  116.09 117.795 116.27 119.5 ;
      RECT  126.17 117.795 126.35 119.5 ;
      RECT  119.93 94.095 120.11 95.8 ;
      RECT  126.17 98.045 126.35 99.75 ;
      RECT  97.37 116.34 97.55 118.045 ;
      RECT  132.41 109.895 132.59 111.6 ;
      RECT  122.33 92.64 122.51 94.345 ;
      RECT  141.05 121.745 141.23 123.45 ;
      RECT  101.21 101.995 101.39 103.7 ;
      RECT  122.33 98.045 122.51 99.75 ;
      RECT  132.41 105.945 132.59 107.65 ;
      RECT  107.45 109.895 107.63 111.6 ;
      RECT  126.17 101.995 126.35 103.7 ;
      RECT  128.57 108.44 128.75 110.145 ;
      RECT  101.21 105.945 101.39 107.65 ;
      RECT  103.61 116.34 103.79 118.045 ;
      RECT  113.69 94.095 113.87 95.8 ;
      RECT  138.65 100.54 138.83 102.245 ;
      RECT  101.21 117.795 101.39 119.5 ;
      RECT  126.17 104.49 126.35 106.195 ;
      RECT  128.57 105.945 128.75 107.65 ;
      RECT  138.65 108.44 138.83 110.145 ;
      RECT  128.57 94.095 128.75 95.8 ;
      RECT  119.93 116.34 120.11 118.045 ;
      RECT  103.61 121.745 103.79 123.45 ;
      RECT  141.05 100.54 141.23 102.245 ;
      RECT  132.41 104.49 132.59 106.195 ;
      RECT  109.85 121.745 110.03 123.45 ;
      RECT  109.85 117.795 110.03 119.5 ;
      RECT  138.65 121.745 138.83 123.45 ;
      RECT  122.33 100.54 122.51 102.245 ;
      RECT  126.17 96.59 126.35 98.295 ;
      RECT  144.89 104.49 145.07 106.195 ;
      RECT  101.21 121.745 101.39 123.45 ;
      RECT  113.69 101.995 113.87 103.7 ;
      RECT  132.41 117.795 132.59 119.5 ;
      RECT  128.57 121.745 128.75 123.45 ;
      RECT  134.81 96.59 134.99 98.295 ;
      RECT  113.69 104.49 113.87 106.195 ;
      RECT  113.69 120.29 113.87 121.995 ;
      RECT  119.93 92.64 120.11 94.345 ;
      RECT  141.05 108.44 141.23 110.145 ;
      RECT  107.45 94.095 107.63 95.8 ;
      RECT  113.69 96.59 113.87 98.295 ;
      RECT  101.21 112.39 101.39 114.095 ;
      RECT  113.69 112.39 113.87 114.095 ;
      RECT  128.57 104.49 128.75 106.195 ;
      RECT  128.57 116.34 128.75 118.045 ;
      RECT  141.05 116.34 141.23 118.045 ;
      RECT  128.57 109.895 128.75 111.6 ;
      RECT  116.09 94.095 116.27 95.8 ;
      RECT  144.89 109.895 145.07 111.6 ;
      RECT  109.85 92.64 110.03 94.345 ;
      RECT  103.61 94.095 103.79 95.8 ;
      RECT  144.89 112.39 145.07 114.095 ;
      RECT  107.45 104.49 107.63 106.195 ;
      RECT  134.81 108.44 134.99 110.145 ;
      RECT  107.45 108.44 107.63 110.145 ;
      RECT  116.09 96.59 116.27 98.295 ;
      RECT  132.41 108.44 132.59 110.145 ;
      RECT  144.89 116.34 145.07 118.045 ;
      RECT  116.09 92.64 116.27 94.345 ;
      RECT  132.41 94.095 132.59 95.8 ;
      RECT  103.61 92.64 103.79 94.345 ;
      RECT  109.85 101.995 110.03 103.7 ;
      RECT  141.05 113.845 141.23 115.55 ;
      RECT  122.33 104.49 122.51 106.195 ;
      RECT  122.33 101.995 122.51 103.7 ;
      RECT  122.33 120.29 122.51 121.995 ;
      RECT  132.41 120.29 132.59 121.995 ;
      RECT  134.81 117.795 134.99 119.5 ;
      RECT  116.09 116.34 116.27 118.045 ;
      RECT  107.45 121.745 107.63 123.45 ;
      RECT  134.81 121.745 134.99 123.45 ;
      RECT  128.57 98.045 128.75 99.75 ;
      RECT  109.85 104.49 110.03 106.195 ;
      RECT  101.21 92.64 101.39 94.345 ;
      RECT  97.37 101.995 97.55 103.7 ;
      RECT  138.65 104.49 138.83 106.195 ;
      RECT  122.33 116.34 122.51 118.045 ;
      RECT  141.05 92.64 141.23 94.345 ;
      RECT  107.45 96.59 107.63 98.295 ;
      RECT  134.81 112.39 134.99 114.095 ;
      RECT  138.65 113.845 138.83 115.55 ;
      RECT  94.79 89.085 94.61 90.665 ;
      RECT  95.15 88.295 94.97 89.085 ;
      RECT  95.19 89.085 95.06 89.795 ;
      RECT  95.51 88.295 95.33 89.085 ;
      RECT  94.43 89.085 94.25 90.665 ;
      RECT  94.79 88.295 94.61 89.085 ;
      RECT  94.43 88.295 94.25 89.085 ;
      RECT  95.87 89.085 95.69 90.665 ;
      RECT  95.87 88.295 95.69 89.085 ;
      RECT  95.51 89.085 95.33 90.665 ;
      RECT  95.06 89.085 94.93 89.795 ;
      RECT  95.15 89.085 94.97 90.665 ;
      RECT  94.07 91.76 93.86 91.35 ;
      RECT  96.47 92.765 96.26 92.435 ;
      RECT  93.425 91.85 93.35 90.145 ;
      RECT  93.51 91.265 93.425 90.855 ;
      RECT  94.43 92.765 94.25 91.85 ;
      POLYGON  93.425 92.765 93.425 92.435 93.86 92.435 93.86 92.055 93.425 92.055 93.425 91.85 93.35 91.85 93.35 92.765 93.425 92.765 ;
      RECT  93.35 91.85 93.14 90.145 ;
      POLYGON  93.86 91.76 93.86 91.35 93.685 91.35 93.605 91.43 93.605 91.76 93.86 91.76 ;
      RECT  96.47 91.85 96.26 90.145 ;
      RECT  94.79 92.765 94.61 91.85 ;
      RECT  95.87 91.85 95.69 90.145 ;
      RECT  94.07 90.77 93.86 90.36 ;
      RECT  93.35 92.055 93.14 91.85 ;
      RECT  96.26 91.85 96.05 90.145 ;
      RECT  94.07 92.435 93.86 92.055 ;
      RECT  95.51 91.85 95.33 90.145 ;
      RECT  94.79 91.85 94.61 90.145 ;
      RECT  95.51 92.765 95.33 91.85 ;
      RECT  93.35 92.765 93.14 92.435 ;
      RECT  95.15 91.85 94.97 90.145 ;
      RECT  95.15 92.765 94.97 91.85 ;
      RECT  96.47 92.055 96.26 91.85 ;
      RECT  93.35 92.435 93.14 92.055 ;
      RECT  94.43 91.85 94.25 90.145 ;
      RECT  96.26 92.055 96.05 91.85 ;
      RECT  96.47 92.435 96.26 92.055 ;
      POLYGON  93.86 90.77 93.86 90.36 93.605 90.36 93.605 90.69 93.685 90.77 93.86 90.77 ;
      RECT  95.87 92.765 95.69 91.85 ;
      RECT  96.26 92.765 96.05 92.435 ;
      RECT  96.26 92.435 96.05 92.055 ;
      RECT  94.07 92.73 93.86 93.14 ;
      RECT  96.47 91.725 96.26 92.055 ;
      RECT  93.425 92.64 93.35 94.345 ;
      RECT  93.51 93.225 93.425 93.635 ;
      RECT  94.43 91.725 94.25 92.64 ;
      POLYGON  93.425 91.725 93.425 92.055 93.86 92.055 93.86 92.435 93.425 92.435 93.425 92.64 93.35 92.64 93.35 91.725 93.425 91.725 ;
      RECT  93.35 92.64 93.14 94.345 ;
      POLYGON  93.86 92.73 93.86 93.14 93.685 93.14 93.605 93.06 93.605 92.73 93.86 92.73 ;
      RECT  96.47 92.64 96.26 94.345 ;
      RECT  94.79 91.725 94.61 92.64 ;
      RECT  95.87 92.64 95.69 94.345 ;
      RECT  94.07 93.72 93.86 94.13 ;
      RECT  93.35 92.435 93.14 92.64 ;
      RECT  96.26 92.64 96.05 94.345 ;
      RECT  94.07 92.055 93.86 92.435 ;
      RECT  95.51 92.64 95.33 94.345 ;
      RECT  94.79 92.64 94.61 94.345 ;
      RECT  95.51 91.725 95.33 92.64 ;
      RECT  93.35 91.725 93.14 92.055 ;
      RECT  95.15 92.64 94.97 94.345 ;
      RECT  95.15 91.725 94.97 92.64 ;
      RECT  96.47 92.435 96.26 92.64 ;
      RECT  93.35 92.055 93.14 92.435 ;
      RECT  94.43 92.64 94.25 94.345 ;
      RECT  96.26 92.435 96.05 92.64 ;
      RECT  96.47 92.055 96.26 92.435 ;
      POLYGON  93.86 93.72 93.86 94.13 93.605 94.13 93.605 93.8 93.685 93.72 93.86 93.72 ;
      RECT  95.87 91.725 95.69 92.64 ;
      RECT  96.26 91.725 96.05 92.055 ;
      RECT  96.26 92.055 96.05 92.435 ;
      RECT  94.07 95.71 93.86 95.3 ;
      RECT  96.47 96.715 96.26 96.385 ;
      RECT  93.425 95.8 93.35 94.095 ;
      RECT  93.51 95.215 93.425 94.805 ;
      RECT  94.43 96.715 94.25 95.8 ;
      POLYGON  93.425 96.715 93.425 96.385 93.86 96.385 93.86 96.005 93.425 96.005 93.425 95.8 93.35 95.8 93.35 96.715 93.425 96.715 ;
      RECT  93.35 95.8 93.14 94.095 ;
      POLYGON  93.86 95.71 93.86 95.3 93.685 95.3 93.605 95.38 93.605 95.71 93.86 95.71 ;
      RECT  96.47 95.8 96.26 94.095 ;
      RECT  94.79 96.715 94.61 95.8 ;
      RECT  95.87 95.8 95.69 94.095 ;
      RECT  94.07 94.72 93.86 94.31 ;
      RECT  93.35 96.005 93.14 95.8 ;
      RECT  96.26 95.8 96.05 94.095 ;
      RECT  94.07 96.385 93.86 96.005 ;
      RECT  95.51 95.8 95.33 94.095 ;
      RECT  94.79 95.8 94.61 94.095 ;
      RECT  95.51 96.715 95.33 95.8 ;
      RECT  93.35 96.715 93.14 96.385 ;
      RECT  95.15 95.8 94.97 94.095 ;
      RECT  95.15 96.715 94.97 95.8 ;
      RECT  96.47 96.005 96.26 95.8 ;
      RECT  93.35 96.385 93.14 96.005 ;
      RECT  94.43 95.8 94.25 94.095 ;
      RECT  96.26 96.005 96.05 95.8 ;
      RECT  96.47 96.385 96.26 96.005 ;
      POLYGON  93.86 94.72 93.86 94.31 93.605 94.31 93.605 94.64 93.685 94.72 93.86 94.72 ;
      RECT  95.87 96.715 95.69 95.8 ;
      RECT  96.26 96.715 96.05 96.385 ;
      RECT  96.26 96.385 96.05 96.005 ;
      RECT  94.07 96.68 93.86 97.09 ;
      RECT  96.47 95.675 96.26 96.005 ;
      RECT  93.425 96.59 93.35 98.295 ;
      RECT  93.51 97.175 93.425 97.585 ;
      RECT  94.43 95.675 94.25 96.59 ;
      POLYGON  93.425 95.675 93.425 96.005 93.86 96.005 93.86 96.385 93.425 96.385 93.425 96.59 93.35 96.59 93.35 95.675 93.425 95.675 ;
      RECT  93.35 96.59 93.14 98.295 ;
      POLYGON  93.86 96.68 93.86 97.09 93.685 97.09 93.605 97.01 93.605 96.68 93.86 96.68 ;
      RECT  96.47 96.59 96.26 98.295 ;
      RECT  94.79 95.675 94.61 96.59 ;
      RECT  95.87 96.59 95.69 98.295 ;
      RECT  94.07 97.67 93.86 98.08 ;
      RECT  93.35 96.385 93.14 96.59 ;
      RECT  96.26 96.59 96.05 98.295 ;
      RECT  94.07 96.005 93.86 96.385 ;
      RECT  95.51 96.59 95.33 98.295 ;
      RECT  94.79 96.59 94.61 98.295 ;
      RECT  95.51 95.675 95.33 96.59 ;
      RECT  93.35 95.675 93.14 96.005 ;
      RECT  95.15 96.59 94.97 98.295 ;
      RECT  95.15 95.675 94.97 96.59 ;
      RECT  96.47 96.385 96.26 96.59 ;
      RECT  93.35 96.005 93.14 96.385 ;
      RECT  94.43 96.59 94.25 98.295 ;
      RECT  96.26 96.385 96.05 96.59 ;
      RECT  96.47 96.005 96.26 96.385 ;
      POLYGON  93.86 97.67 93.86 98.08 93.605 98.08 93.605 97.75 93.685 97.67 93.86 97.67 ;
      RECT  95.87 95.675 95.69 96.59 ;
      RECT  96.26 95.675 96.05 96.005 ;
      RECT  96.26 96.005 96.05 96.385 ;
      RECT  94.07 99.66 93.86 99.25 ;
      RECT  96.47 100.665 96.26 100.335 ;
      RECT  93.425 99.75 93.35 98.045 ;
      RECT  93.51 99.165 93.425 98.755 ;
      RECT  94.43 100.665 94.25 99.75 ;
      POLYGON  93.425 100.665 93.425 100.335 93.86 100.335 93.86 99.955 93.425 99.955 93.425 99.75 93.35 99.75 93.35 100.665 93.425 100.665 ;
      RECT  93.35 99.75 93.14 98.045 ;
      POLYGON  93.86 99.66 93.86 99.25 93.685 99.25 93.605 99.33 93.605 99.66 93.86 99.66 ;
      RECT  96.47 99.75 96.26 98.045 ;
      RECT  94.79 100.665 94.61 99.75 ;
      RECT  95.87 99.75 95.69 98.045 ;
      RECT  94.07 98.67 93.86 98.26 ;
      RECT  93.35 99.955 93.14 99.75 ;
      RECT  96.26 99.75 96.05 98.045 ;
      RECT  94.07 100.335 93.86 99.955 ;
      RECT  95.51 99.75 95.33 98.045 ;
      RECT  94.79 99.75 94.61 98.045 ;
      RECT  95.51 100.665 95.33 99.75 ;
      RECT  93.35 100.665 93.14 100.335 ;
      RECT  95.15 99.75 94.97 98.045 ;
      RECT  95.15 100.665 94.97 99.75 ;
      RECT  96.47 99.955 96.26 99.75 ;
      RECT  93.35 100.335 93.14 99.955 ;
      RECT  94.43 99.75 94.25 98.045 ;
      RECT  96.26 99.955 96.05 99.75 ;
      RECT  96.47 100.335 96.26 99.955 ;
      POLYGON  93.86 98.67 93.86 98.26 93.605 98.26 93.605 98.59 93.685 98.67 93.86 98.67 ;
      RECT  95.87 100.665 95.69 99.75 ;
      RECT  96.26 100.665 96.05 100.335 ;
      RECT  96.26 100.335 96.05 99.955 ;
      RECT  94.07 100.63 93.86 101.04 ;
      RECT  96.47 99.625 96.26 99.955 ;
      RECT  93.425 100.54 93.35 102.245 ;
      RECT  93.51 101.125 93.425 101.535 ;
      RECT  94.43 99.625 94.25 100.54 ;
      POLYGON  93.425 99.625 93.425 99.955 93.86 99.955 93.86 100.335 93.425 100.335 93.425 100.54 93.35 100.54 93.35 99.625 93.425 99.625 ;
      RECT  93.35 100.54 93.14 102.245 ;
      POLYGON  93.86 100.63 93.86 101.04 93.685 101.04 93.605 100.96 93.605 100.63 93.86 100.63 ;
      RECT  96.47 100.54 96.26 102.245 ;
      RECT  94.79 99.625 94.61 100.54 ;
      RECT  95.87 100.54 95.69 102.245 ;
      RECT  94.07 101.62 93.86 102.03 ;
      RECT  93.35 100.335 93.14 100.54 ;
      RECT  96.26 100.54 96.05 102.245 ;
      RECT  94.07 99.955 93.86 100.335 ;
      RECT  95.51 100.54 95.33 102.245 ;
      RECT  94.79 100.54 94.61 102.245 ;
      RECT  95.51 99.625 95.33 100.54 ;
      RECT  93.35 99.625 93.14 99.955 ;
      RECT  95.15 100.54 94.97 102.245 ;
      RECT  95.15 99.625 94.97 100.54 ;
      RECT  96.47 100.335 96.26 100.54 ;
      RECT  93.35 99.955 93.14 100.335 ;
      RECT  94.43 100.54 94.25 102.245 ;
      RECT  96.26 100.335 96.05 100.54 ;
      RECT  96.47 99.955 96.26 100.335 ;
      POLYGON  93.86 101.62 93.86 102.03 93.605 102.03 93.605 101.7 93.685 101.62 93.86 101.62 ;
      RECT  95.87 99.625 95.69 100.54 ;
      RECT  96.26 99.625 96.05 99.955 ;
      RECT  96.26 99.955 96.05 100.335 ;
      RECT  94.07 103.61 93.86 103.2 ;
      RECT  96.47 104.615 96.26 104.285 ;
      RECT  93.425 103.7 93.35 101.995 ;
      RECT  93.51 103.115 93.425 102.705 ;
      RECT  94.43 104.615 94.25 103.7 ;
      POLYGON  93.425 104.615 93.425 104.285 93.86 104.285 93.86 103.905 93.425 103.905 93.425 103.7 93.35 103.7 93.35 104.615 93.425 104.615 ;
      RECT  93.35 103.7 93.14 101.995 ;
      POLYGON  93.86 103.61 93.86 103.2 93.685 103.2 93.605 103.28 93.605 103.61 93.86 103.61 ;
      RECT  96.47 103.7 96.26 101.995 ;
      RECT  94.79 104.615 94.61 103.7 ;
      RECT  95.87 103.7 95.69 101.995 ;
      RECT  94.07 102.62 93.86 102.21 ;
      RECT  93.35 103.905 93.14 103.7 ;
      RECT  96.26 103.7 96.05 101.995 ;
      RECT  94.07 104.285 93.86 103.905 ;
      RECT  95.51 103.7 95.33 101.995 ;
      RECT  94.79 103.7 94.61 101.995 ;
      RECT  95.51 104.615 95.33 103.7 ;
      RECT  93.35 104.615 93.14 104.285 ;
      RECT  95.15 103.7 94.97 101.995 ;
      RECT  95.15 104.615 94.97 103.7 ;
      RECT  96.47 103.905 96.26 103.7 ;
      RECT  93.35 104.285 93.14 103.905 ;
      RECT  94.43 103.7 94.25 101.995 ;
      RECT  96.26 103.905 96.05 103.7 ;
      RECT  96.47 104.285 96.26 103.905 ;
      POLYGON  93.86 102.62 93.86 102.21 93.605 102.21 93.605 102.54 93.685 102.62 93.86 102.62 ;
      RECT  95.87 104.615 95.69 103.7 ;
      RECT  96.26 104.615 96.05 104.285 ;
      RECT  96.26 104.285 96.05 103.905 ;
      RECT  94.07 104.58 93.86 104.99 ;
      RECT  96.47 103.575 96.26 103.905 ;
      RECT  93.425 104.49 93.35 106.195 ;
      RECT  93.51 105.075 93.425 105.485 ;
      RECT  94.43 103.575 94.25 104.49 ;
      POLYGON  93.425 103.575 93.425 103.905 93.86 103.905 93.86 104.285 93.425 104.285 93.425 104.49 93.35 104.49 93.35 103.575 93.425 103.575 ;
      RECT  93.35 104.49 93.14 106.195 ;
      POLYGON  93.86 104.58 93.86 104.99 93.685 104.99 93.605 104.91 93.605 104.58 93.86 104.58 ;
      RECT  96.47 104.49 96.26 106.195 ;
      RECT  94.79 103.575 94.61 104.49 ;
      RECT  95.87 104.49 95.69 106.195 ;
      RECT  94.07 105.57 93.86 105.98 ;
      RECT  93.35 104.285 93.14 104.49 ;
      RECT  96.26 104.49 96.05 106.195 ;
      RECT  94.07 103.905 93.86 104.285 ;
      RECT  95.51 104.49 95.33 106.195 ;
      RECT  94.79 104.49 94.61 106.195 ;
      RECT  95.51 103.575 95.33 104.49 ;
      RECT  93.35 103.575 93.14 103.905 ;
      RECT  95.15 104.49 94.97 106.195 ;
      RECT  95.15 103.575 94.97 104.49 ;
      RECT  96.47 104.285 96.26 104.49 ;
      RECT  93.35 103.905 93.14 104.285 ;
      RECT  94.43 104.49 94.25 106.195 ;
      RECT  96.26 104.285 96.05 104.49 ;
      RECT  96.47 103.905 96.26 104.285 ;
      POLYGON  93.86 105.57 93.86 105.98 93.605 105.98 93.605 105.65 93.685 105.57 93.86 105.57 ;
      RECT  95.87 103.575 95.69 104.49 ;
      RECT  96.26 103.575 96.05 103.905 ;
      RECT  96.26 103.905 96.05 104.285 ;
      RECT  94.07 107.56 93.86 107.15 ;
      RECT  96.47 108.565 96.26 108.235 ;
      RECT  93.425 107.65 93.35 105.945 ;
      RECT  93.51 107.065 93.425 106.655 ;
      RECT  94.43 108.565 94.25 107.65 ;
      POLYGON  93.425 108.565 93.425 108.235 93.86 108.235 93.86 107.855 93.425 107.855 93.425 107.65 93.35 107.65 93.35 108.565 93.425 108.565 ;
      RECT  93.35 107.65 93.14 105.945 ;
      POLYGON  93.86 107.56 93.86 107.15 93.685 107.15 93.605 107.23 93.605 107.56 93.86 107.56 ;
      RECT  96.47 107.65 96.26 105.945 ;
      RECT  94.79 108.565 94.61 107.65 ;
      RECT  95.87 107.65 95.69 105.945 ;
      RECT  94.07 106.57 93.86 106.16 ;
      RECT  93.35 107.855 93.14 107.65 ;
      RECT  96.26 107.65 96.05 105.945 ;
      RECT  94.07 108.235 93.86 107.855 ;
      RECT  95.51 107.65 95.33 105.945 ;
      RECT  94.79 107.65 94.61 105.945 ;
      RECT  95.51 108.565 95.33 107.65 ;
      RECT  93.35 108.565 93.14 108.235 ;
      RECT  95.15 107.65 94.97 105.945 ;
      RECT  95.15 108.565 94.97 107.65 ;
      RECT  96.47 107.855 96.26 107.65 ;
      RECT  93.35 108.235 93.14 107.855 ;
      RECT  94.43 107.65 94.25 105.945 ;
      RECT  96.26 107.855 96.05 107.65 ;
      RECT  96.47 108.235 96.26 107.855 ;
      POLYGON  93.86 106.57 93.86 106.16 93.605 106.16 93.605 106.49 93.685 106.57 93.86 106.57 ;
      RECT  95.87 108.565 95.69 107.65 ;
      RECT  96.26 108.565 96.05 108.235 ;
      RECT  96.26 108.235 96.05 107.855 ;
      RECT  94.07 108.53 93.86 108.94 ;
      RECT  96.47 107.525 96.26 107.855 ;
      RECT  93.425 108.44 93.35 110.145 ;
      RECT  93.51 109.025 93.425 109.435 ;
      RECT  94.43 107.525 94.25 108.44 ;
      POLYGON  93.425 107.525 93.425 107.855 93.86 107.855 93.86 108.235 93.425 108.235 93.425 108.44 93.35 108.44 93.35 107.525 93.425 107.525 ;
      RECT  93.35 108.44 93.14 110.145 ;
      POLYGON  93.86 108.53 93.86 108.94 93.685 108.94 93.605 108.86 93.605 108.53 93.86 108.53 ;
      RECT  96.47 108.44 96.26 110.145 ;
      RECT  94.79 107.525 94.61 108.44 ;
      RECT  95.87 108.44 95.69 110.145 ;
      RECT  94.07 109.52 93.86 109.93 ;
      RECT  93.35 108.235 93.14 108.44 ;
      RECT  96.26 108.44 96.05 110.145 ;
      RECT  94.07 107.855 93.86 108.235 ;
      RECT  95.51 108.44 95.33 110.145 ;
      RECT  94.79 108.44 94.61 110.145 ;
      RECT  95.51 107.525 95.33 108.44 ;
      RECT  93.35 107.525 93.14 107.855 ;
      RECT  95.15 108.44 94.97 110.145 ;
      RECT  95.15 107.525 94.97 108.44 ;
      RECT  96.47 108.235 96.26 108.44 ;
      RECT  93.35 107.855 93.14 108.235 ;
      RECT  94.43 108.44 94.25 110.145 ;
      RECT  96.26 108.235 96.05 108.44 ;
      RECT  96.47 107.855 96.26 108.235 ;
      POLYGON  93.86 109.52 93.86 109.93 93.605 109.93 93.605 109.6 93.685 109.52 93.86 109.52 ;
      RECT  95.87 107.525 95.69 108.44 ;
      RECT  96.26 107.525 96.05 107.855 ;
      RECT  96.26 107.855 96.05 108.235 ;
      RECT  94.07 111.51 93.86 111.1 ;
      RECT  96.47 112.515 96.26 112.185 ;
      RECT  93.425 111.6 93.35 109.895 ;
      RECT  93.51 111.015 93.425 110.605 ;
      RECT  94.43 112.515 94.25 111.6 ;
      POLYGON  93.425 112.515 93.425 112.185 93.86 112.185 93.86 111.805 93.425 111.805 93.425 111.6 93.35 111.6 93.35 112.515 93.425 112.515 ;
      RECT  93.35 111.6 93.14 109.895 ;
      POLYGON  93.86 111.51 93.86 111.1 93.685 111.1 93.605 111.18 93.605 111.51 93.86 111.51 ;
      RECT  96.47 111.6 96.26 109.895 ;
      RECT  94.79 112.515 94.61 111.6 ;
      RECT  95.87 111.6 95.69 109.895 ;
      RECT  94.07 110.52 93.86 110.11 ;
      RECT  93.35 111.805 93.14 111.6 ;
      RECT  96.26 111.6 96.05 109.895 ;
      RECT  94.07 112.185 93.86 111.805 ;
      RECT  95.51 111.6 95.33 109.895 ;
      RECT  94.79 111.6 94.61 109.895 ;
      RECT  95.51 112.515 95.33 111.6 ;
      RECT  93.35 112.515 93.14 112.185 ;
      RECT  95.15 111.6 94.97 109.895 ;
      RECT  95.15 112.515 94.97 111.6 ;
      RECT  96.47 111.805 96.26 111.6 ;
      RECT  93.35 112.185 93.14 111.805 ;
      RECT  94.43 111.6 94.25 109.895 ;
      RECT  96.26 111.805 96.05 111.6 ;
      RECT  96.47 112.185 96.26 111.805 ;
      POLYGON  93.86 110.52 93.86 110.11 93.605 110.11 93.605 110.44 93.685 110.52 93.86 110.52 ;
      RECT  95.87 112.515 95.69 111.6 ;
      RECT  96.26 112.515 96.05 112.185 ;
      RECT  96.26 112.185 96.05 111.805 ;
      RECT  94.07 112.48 93.86 112.89 ;
      RECT  96.47 111.475 96.26 111.805 ;
      RECT  93.425 112.39 93.35 114.095 ;
      RECT  93.51 112.975 93.425 113.385 ;
      RECT  94.43 111.475 94.25 112.39 ;
      POLYGON  93.425 111.475 93.425 111.805 93.86 111.805 93.86 112.185 93.425 112.185 93.425 112.39 93.35 112.39 93.35 111.475 93.425 111.475 ;
      RECT  93.35 112.39 93.14 114.095 ;
      POLYGON  93.86 112.48 93.86 112.89 93.685 112.89 93.605 112.81 93.605 112.48 93.86 112.48 ;
      RECT  96.47 112.39 96.26 114.095 ;
      RECT  94.79 111.475 94.61 112.39 ;
      RECT  95.87 112.39 95.69 114.095 ;
      RECT  94.07 113.47 93.86 113.88 ;
      RECT  93.35 112.185 93.14 112.39 ;
      RECT  96.26 112.39 96.05 114.095 ;
      RECT  94.07 111.805 93.86 112.185 ;
      RECT  95.51 112.39 95.33 114.095 ;
      RECT  94.79 112.39 94.61 114.095 ;
      RECT  95.51 111.475 95.33 112.39 ;
      RECT  93.35 111.475 93.14 111.805 ;
      RECT  95.15 112.39 94.97 114.095 ;
      RECT  95.15 111.475 94.97 112.39 ;
      RECT  96.47 112.185 96.26 112.39 ;
      RECT  93.35 111.805 93.14 112.185 ;
      RECT  94.43 112.39 94.25 114.095 ;
      RECT  96.26 112.185 96.05 112.39 ;
      RECT  96.47 111.805 96.26 112.185 ;
      POLYGON  93.86 113.47 93.86 113.88 93.605 113.88 93.605 113.55 93.685 113.47 93.86 113.47 ;
      RECT  95.87 111.475 95.69 112.39 ;
      RECT  96.26 111.475 96.05 111.805 ;
      RECT  96.26 111.805 96.05 112.185 ;
      RECT  94.07 115.46 93.86 115.05 ;
      RECT  96.47 116.465 96.26 116.135 ;
      RECT  93.425 115.55 93.35 113.845 ;
      RECT  93.51 114.965 93.425 114.555 ;
      RECT  94.43 116.465 94.25 115.55 ;
      POLYGON  93.425 116.465 93.425 116.135 93.86 116.135 93.86 115.755 93.425 115.755 93.425 115.55 93.35 115.55 93.35 116.465 93.425 116.465 ;
      RECT  93.35 115.55 93.14 113.845 ;
      POLYGON  93.86 115.46 93.86 115.05 93.685 115.05 93.605 115.13 93.605 115.46 93.86 115.46 ;
      RECT  96.47 115.55 96.26 113.845 ;
      RECT  94.79 116.465 94.61 115.55 ;
      RECT  95.87 115.55 95.69 113.845 ;
      RECT  94.07 114.47 93.86 114.06 ;
      RECT  93.35 115.755 93.14 115.55 ;
      RECT  96.26 115.55 96.05 113.845 ;
      RECT  94.07 116.135 93.86 115.755 ;
      RECT  95.51 115.55 95.33 113.845 ;
      RECT  94.79 115.55 94.61 113.845 ;
      RECT  95.51 116.465 95.33 115.55 ;
      RECT  93.35 116.465 93.14 116.135 ;
      RECT  95.15 115.55 94.97 113.845 ;
      RECT  95.15 116.465 94.97 115.55 ;
      RECT  96.47 115.755 96.26 115.55 ;
      RECT  93.35 116.135 93.14 115.755 ;
      RECT  94.43 115.55 94.25 113.845 ;
      RECT  96.26 115.755 96.05 115.55 ;
      RECT  96.47 116.135 96.26 115.755 ;
      POLYGON  93.86 114.47 93.86 114.06 93.605 114.06 93.605 114.39 93.685 114.47 93.86 114.47 ;
      RECT  95.87 116.465 95.69 115.55 ;
      RECT  96.26 116.465 96.05 116.135 ;
      RECT  96.26 116.135 96.05 115.755 ;
      RECT  94.07 116.43 93.86 116.84 ;
      RECT  96.47 115.425 96.26 115.755 ;
      RECT  93.425 116.34 93.35 118.045 ;
      RECT  93.51 116.925 93.425 117.335 ;
      RECT  94.43 115.425 94.25 116.34 ;
      POLYGON  93.425 115.425 93.425 115.755 93.86 115.755 93.86 116.135 93.425 116.135 93.425 116.34 93.35 116.34 93.35 115.425 93.425 115.425 ;
      RECT  93.35 116.34 93.14 118.045 ;
      POLYGON  93.86 116.43 93.86 116.84 93.685 116.84 93.605 116.76 93.605 116.43 93.86 116.43 ;
      RECT  96.47 116.34 96.26 118.045 ;
      RECT  94.79 115.425 94.61 116.34 ;
      RECT  95.87 116.34 95.69 118.045 ;
      RECT  94.07 117.42 93.86 117.83 ;
      RECT  93.35 116.135 93.14 116.34 ;
      RECT  96.26 116.34 96.05 118.045 ;
      RECT  94.07 115.755 93.86 116.135 ;
      RECT  95.51 116.34 95.33 118.045 ;
      RECT  94.79 116.34 94.61 118.045 ;
      RECT  95.51 115.425 95.33 116.34 ;
      RECT  93.35 115.425 93.14 115.755 ;
      RECT  95.15 116.34 94.97 118.045 ;
      RECT  95.15 115.425 94.97 116.34 ;
      RECT  96.47 116.135 96.26 116.34 ;
      RECT  93.35 115.755 93.14 116.135 ;
      RECT  94.43 116.34 94.25 118.045 ;
      RECT  96.26 116.135 96.05 116.34 ;
      RECT  96.47 115.755 96.26 116.135 ;
      POLYGON  93.86 117.42 93.86 117.83 93.605 117.83 93.605 117.5 93.685 117.42 93.86 117.42 ;
      RECT  95.87 115.425 95.69 116.34 ;
      RECT  96.26 115.425 96.05 115.755 ;
      RECT  96.26 115.755 96.05 116.135 ;
      RECT  94.07 119.41 93.86 119.0 ;
      RECT  96.47 120.415 96.26 120.085 ;
      RECT  93.425 119.5 93.35 117.795 ;
      RECT  93.51 118.915 93.425 118.505 ;
      RECT  94.43 120.415 94.25 119.5 ;
      POLYGON  93.425 120.415 93.425 120.085 93.86 120.085 93.86 119.705 93.425 119.705 93.425 119.5 93.35 119.5 93.35 120.415 93.425 120.415 ;
      RECT  93.35 119.5 93.14 117.795 ;
      POLYGON  93.86 119.41 93.86 119.0 93.685 119.0 93.605 119.08 93.605 119.41 93.86 119.41 ;
      RECT  96.47 119.5 96.26 117.795 ;
      RECT  94.79 120.415 94.61 119.5 ;
      RECT  95.87 119.5 95.69 117.795 ;
      RECT  94.07 118.42 93.86 118.01 ;
      RECT  93.35 119.705 93.14 119.5 ;
      RECT  96.26 119.5 96.05 117.795 ;
      RECT  94.07 120.085 93.86 119.705 ;
      RECT  95.51 119.5 95.33 117.795 ;
      RECT  94.79 119.5 94.61 117.795 ;
      RECT  95.51 120.415 95.33 119.5 ;
      RECT  93.35 120.415 93.14 120.085 ;
      RECT  95.15 119.5 94.97 117.795 ;
      RECT  95.15 120.415 94.97 119.5 ;
      RECT  96.47 119.705 96.26 119.5 ;
      RECT  93.35 120.085 93.14 119.705 ;
      RECT  94.43 119.5 94.25 117.795 ;
      RECT  96.26 119.705 96.05 119.5 ;
      RECT  96.47 120.085 96.26 119.705 ;
      POLYGON  93.86 118.42 93.86 118.01 93.605 118.01 93.605 118.34 93.685 118.42 93.86 118.42 ;
      RECT  95.87 120.415 95.69 119.5 ;
      RECT  96.26 120.415 96.05 120.085 ;
      RECT  96.26 120.085 96.05 119.705 ;
      RECT  94.07 120.38 93.86 120.79 ;
      RECT  96.47 119.375 96.26 119.705 ;
      RECT  93.425 120.29 93.35 121.995 ;
      RECT  93.51 120.875 93.425 121.285 ;
      RECT  94.43 119.375 94.25 120.29 ;
      POLYGON  93.425 119.375 93.425 119.705 93.86 119.705 93.86 120.085 93.425 120.085 93.425 120.29 93.35 120.29 93.35 119.375 93.425 119.375 ;
      RECT  93.35 120.29 93.14 121.995 ;
      POLYGON  93.86 120.38 93.86 120.79 93.685 120.79 93.605 120.71 93.605 120.38 93.86 120.38 ;
      RECT  96.47 120.29 96.26 121.995 ;
      RECT  94.79 119.375 94.61 120.29 ;
      RECT  95.87 120.29 95.69 121.995 ;
      RECT  94.07 121.37 93.86 121.78 ;
      RECT  93.35 120.085 93.14 120.29 ;
      RECT  96.26 120.29 96.05 121.995 ;
      RECT  94.07 119.705 93.86 120.085 ;
      RECT  95.51 120.29 95.33 121.995 ;
      RECT  94.79 120.29 94.61 121.995 ;
      RECT  95.51 119.375 95.33 120.29 ;
      RECT  93.35 119.375 93.14 119.705 ;
      RECT  95.15 120.29 94.97 121.995 ;
      RECT  95.15 119.375 94.97 120.29 ;
      RECT  96.47 120.085 96.26 120.29 ;
      RECT  93.35 119.705 93.14 120.085 ;
      RECT  94.43 120.29 94.25 121.995 ;
      RECT  96.26 120.085 96.05 120.29 ;
      RECT  96.47 119.705 96.26 120.085 ;
      POLYGON  93.86 121.37 93.86 121.78 93.605 121.78 93.605 121.45 93.685 121.37 93.86 121.37 ;
      RECT  95.87 119.375 95.69 120.29 ;
      RECT  96.26 119.375 96.05 119.705 ;
      RECT  96.26 119.705 96.05 120.085 ;
      RECT  94.07 123.36 93.86 122.95 ;
      RECT  96.47 124.365 96.26 124.035 ;
      RECT  93.425 123.45 93.35 121.745 ;
      RECT  93.51 122.865 93.425 122.455 ;
      RECT  94.43 124.365 94.25 123.45 ;
      POLYGON  93.425 124.365 93.425 124.035 93.86 124.035 93.86 123.655 93.425 123.655 93.425 123.45 93.35 123.45 93.35 124.365 93.425 124.365 ;
      RECT  93.35 123.45 93.14 121.745 ;
      POLYGON  93.86 123.36 93.86 122.95 93.685 122.95 93.605 123.03 93.605 123.36 93.86 123.36 ;
      RECT  96.47 123.45 96.26 121.745 ;
      RECT  94.79 124.365 94.61 123.45 ;
      RECT  95.87 123.45 95.69 121.745 ;
      RECT  94.07 122.37 93.86 121.96 ;
      RECT  93.35 123.655 93.14 123.45 ;
      RECT  96.26 123.45 96.05 121.745 ;
      RECT  94.07 124.035 93.86 123.655 ;
      RECT  95.51 123.45 95.33 121.745 ;
      RECT  94.79 123.45 94.61 121.745 ;
      RECT  95.51 124.365 95.33 123.45 ;
      RECT  93.35 124.365 93.14 124.035 ;
      RECT  95.15 123.45 94.97 121.745 ;
      RECT  95.15 124.365 94.97 123.45 ;
      RECT  96.47 123.655 96.26 123.45 ;
      RECT  93.35 124.035 93.14 123.655 ;
      RECT  94.43 123.45 94.25 121.745 ;
      RECT  96.26 123.655 96.05 123.45 ;
      RECT  96.47 124.035 96.26 123.655 ;
      POLYGON  93.86 122.37 93.86 121.96 93.605 121.96 93.605 122.29 93.685 122.37 93.86 122.37 ;
      RECT  95.87 124.365 95.69 123.45 ;
      RECT  96.26 124.365 96.05 124.035 ;
      RECT  96.26 124.035 96.05 123.655 ;
      RECT  94.07 124.33 93.86 124.74 ;
      RECT  96.47 123.325 96.26 123.655 ;
      RECT  93.425 124.24 93.35 125.945 ;
      RECT  93.51 124.825 93.425 125.235 ;
      RECT  94.43 123.325 94.25 124.24 ;
      POLYGON  93.425 123.325 93.425 123.655 93.86 123.655 93.86 124.035 93.425 124.035 93.425 124.24 93.35 124.24 93.35 123.325 93.425 123.325 ;
      RECT  93.35 124.24 93.14 125.945 ;
      POLYGON  93.86 124.33 93.86 124.74 93.685 124.74 93.605 124.66 93.605 124.33 93.86 124.33 ;
      RECT  96.47 124.24 96.26 125.945 ;
      RECT  94.79 123.325 94.61 124.24 ;
      RECT  95.87 124.24 95.69 125.945 ;
      RECT  94.07 125.32 93.86 125.73 ;
      RECT  93.35 124.035 93.14 124.24 ;
      RECT  96.26 124.24 96.05 125.945 ;
      RECT  94.07 123.655 93.86 124.035 ;
      RECT  95.51 124.24 95.33 125.945 ;
      RECT  94.79 124.24 94.61 125.945 ;
      RECT  95.51 123.325 95.33 124.24 ;
      RECT  93.35 123.325 93.14 123.655 ;
      RECT  95.15 124.24 94.97 125.945 ;
      RECT  95.15 123.325 94.97 124.24 ;
      RECT  96.47 124.035 96.26 124.24 ;
      RECT  93.35 123.655 93.14 124.035 ;
      RECT  94.43 124.24 94.25 125.945 ;
      RECT  96.26 124.035 96.05 124.24 ;
      RECT  96.47 123.655 96.26 124.035 ;
      POLYGON  93.86 125.32 93.86 125.73 93.605 125.73 93.605 125.4 93.685 125.32 93.86 125.32 ;
      RECT  95.87 123.325 95.69 124.24 ;
      RECT  96.26 123.325 96.05 123.655 ;
      RECT  96.26 123.655 96.05 124.035 ;
      RECT  94.79 127.005 94.61 125.425 ;
      RECT  95.15 127.795 94.97 127.005 ;
      RECT  95.19 127.005 95.06 126.295 ;
      RECT  95.51 127.795 95.33 127.005 ;
      RECT  94.43 127.005 94.25 125.425 ;
      RECT  94.79 127.795 94.61 127.005 ;
      RECT  94.43 127.795 94.25 127.005 ;
      RECT  95.87 127.005 95.69 125.425 ;
      RECT  95.87 127.795 95.69 127.005 ;
      RECT  95.51 127.005 95.33 125.425 ;
      RECT  95.06 127.005 94.93 126.295 ;
      RECT  95.15 127.005 94.97 125.425 ;
      RECT  94.97 124.24 95.15 125.945 ;
      RECT  94.97 96.59 95.15 98.295 ;
      RECT  94.97 92.64 95.15 94.345 ;
      RECT  94.97 101.995 95.15 103.7 ;
      RECT  94.97 117.795 95.15 119.5 ;
      RECT  94.97 105.945 95.15 107.65 ;
      RECT  94.97 121.745 95.15 123.45 ;
      RECT  94.97 94.095 95.15 95.8 ;
      RECT  94.97 109.895 95.15 111.6 ;
      RECT  94.97 108.44 95.15 110.145 ;
      RECT  94.97 90.145 95.15 91.85 ;
      RECT  94.97 104.49 95.15 106.195 ;
      RECT  94.97 98.045 95.15 99.75 ;
      RECT  94.97 116.34 95.15 118.045 ;
      RECT  94.97 112.39 95.15 114.095 ;
      RECT  94.97 120.29 95.15 121.995 ;
      RECT  94.97 100.54 95.15 102.245 ;
      RECT  94.97 113.845 95.15 115.55 ;
      RECT  147.65 89.085 147.83 90.665 ;
      RECT  147.29 88.295 147.47 89.085 ;
      RECT  147.25 89.085 147.38 89.795 ;
      RECT  146.93 88.295 147.11 89.085 ;
      RECT  148.01 89.085 148.19 90.665 ;
      RECT  147.65 88.295 147.83 89.085 ;
      RECT  148.01 88.295 148.19 89.085 ;
      RECT  146.57 89.085 146.75 90.665 ;
      RECT  146.57 88.295 146.75 89.085 ;
      RECT  146.93 89.085 147.11 90.665 ;
      RECT  147.38 89.085 147.51 89.795 ;
      RECT  147.29 89.085 147.47 90.665 ;
      RECT  148.37 91.76 148.58 91.35 ;
      RECT  145.97 92.765 146.18 92.435 ;
      RECT  149.015 91.85 149.09 90.145 ;
      RECT  148.93 91.265 149.015 90.855 ;
      RECT  148.01 92.765 148.19 91.85 ;
      POLYGON  149.015 92.765 149.015 92.435 148.58 92.435 148.58 92.055 149.015 92.055 149.015 91.85 149.09 91.85 149.09 92.765 149.015 92.765 ;
      RECT  149.09 91.85 149.3 90.145 ;
      POLYGON  148.58 91.76 148.58 91.35 148.755 91.35 148.835 91.43 148.835 91.76 148.58 91.76 ;
      RECT  145.97 91.85 146.18 90.145 ;
      RECT  147.65 92.765 147.83 91.85 ;
      RECT  146.57 91.85 146.75 90.145 ;
      RECT  148.37 90.77 148.58 90.36 ;
      RECT  149.09 92.055 149.3 91.85 ;
      RECT  146.18 91.85 146.39 90.145 ;
      RECT  148.37 92.435 148.58 92.055 ;
      RECT  146.93 91.85 147.11 90.145 ;
      RECT  147.65 91.85 147.83 90.145 ;
      RECT  146.93 92.765 147.11 91.85 ;
      RECT  149.09 92.765 149.3 92.435 ;
      RECT  147.29 91.85 147.47 90.145 ;
      RECT  147.29 92.765 147.47 91.85 ;
      RECT  145.97 92.055 146.18 91.85 ;
      RECT  149.09 92.435 149.3 92.055 ;
      RECT  148.01 91.85 148.19 90.145 ;
      RECT  146.18 92.055 146.39 91.85 ;
      RECT  145.97 92.435 146.18 92.055 ;
      POLYGON  148.58 90.77 148.58 90.36 148.835 90.36 148.835 90.69 148.755 90.77 148.58 90.77 ;
      RECT  146.57 92.765 146.75 91.85 ;
      RECT  146.18 92.765 146.39 92.435 ;
      RECT  146.18 92.435 146.39 92.055 ;
      RECT  148.37 92.73 148.58 93.14 ;
      RECT  145.97 91.725 146.18 92.055 ;
      RECT  149.015 92.64 149.09 94.345 ;
      RECT  148.93 93.225 149.015 93.635 ;
      RECT  148.01 91.725 148.19 92.64 ;
      POLYGON  149.015 91.725 149.015 92.055 148.58 92.055 148.58 92.435 149.015 92.435 149.015 92.64 149.09 92.64 149.09 91.725 149.015 91.725 ;
      RECT  149.09 92.64 149.3 94.345 ;
      POLYGON  148.58 92.73 148.58 93.14 148.755 93.14 148.835 93.06 148.835 92.73 148.58 92.73 ;
      RECT  145.97 92.64 146.18 94.345 ;
      RECT  147.65 91.725 147.83 92.64 ;
      RECT  146.57 92.64 146.75 94.345 ;
      RECT  148.37 93.72 148.58 94.13 ;
      RECT  149.09 92.435 149.3 92.64 ;
      RECT  146.18 92.64 146.39 94.345 ;
      RECT  148.37 92.055 148.58 92.435 ;
      RECT  146.93 92.64 147.11 94.345 ;
      RECT  147.65 92.64 147.83 94.345 ;
      RECT  146.93 91.725 147.11 92.64 ;
      RECT  149.09 91.725 149.3 92.055 ;
      RECT  147.29 92.64 147.47 94.345 ;
      RECT  147.29 91.725 147.47 92.64 ;
      RECT  145.97 92.435 146.18 92.64 ;
      RECT  149.09 92.055 149.3 92.435 ;
      RECT  148.01 92.64 148.19 94.345 ;
      RECT  146.18 92.435 146.39 92.64 ;
      RECT  145.97 92.055 146.18 92.435 ;
      POLYGON  148.58 93.72 148.58 94.13 148.835 94.13 148.835 93.8 148.755 93.72 148.58 93.72 ;
      RECT  146.57 91.725 146.75 92.64 ;
      RECT  146.18 91.725 146.39 92.055 ;
      RECT  146.18 92.055 146.39 92.435 ;
      RECT  148.37 95.71 148.58 95.3 ;
      RECT  145.97 96.715 146.18 96.385 ;
      RECT  149.015 95.8 149.09 94.095 ;
      RECT  148.93 95.215 149.015 94.805 ;
      RECT  148.01 96.715 148.19 95.8 ;
      POLYGON  149.015 96.715 149.015 96.385 148.58 96.385 148.58 96.005 149.015 96.005 149.015 95.8 149.09 95.8 149.09 96.715 149.015 96.715 ;
      RECT  149.09 95.8 149.3 94.095 ;
      POLYGON  148.58 95.71 148.58 95.3 148.755 95.3 148.835 95.38 148.835 95.71 148.58 95.71 ;
      RECT  145.97 95.8 146.18 94.095 ;
      RECT  147.65 96.715 147.83 95.8 ;
      RECT  146.57 95.8 146.75 94.095 ;
      RECT  148.37 94.72 148.58 94.31 ;
      RECT  149.09 96.005 149.3 95.8 ;
      RECT  146.18 95.8 146.39 94.095 ;
      RECT  148.37 96.385 148.58 96.005 ;
      RECT  146.93 95.8 147.11 94.095 ;
      RECT  147.65 95.8 147.83 94.095 ;
      RECT  146.93 96.715 147.11 95.8 ;
      RECT  149.09 96.715 149.3 96.385 ;
      RECT  147.29 95.8 147.47 94.095 ;
      RECT  147.29 96.715 147.47 95.8 ;
      RECT  145.97 96.005 146.18 95.8 ;
      RECT  149.09 96.385 149.3 96.005 ;
      RECT  148.01 95.8 148.19 94.095 ;
      RECT  146.18 96.005 146.39 95.8 ;
      RECT  145.97 96.385 146.18 96.005 ;
      POLYGON  148.58 94.72 148.58 94.31 148.835 94.31 148.835 94.64 148.755 94.72 148.58 94.72 ;
      RECT  146.57 96.715 146.75 95.8 ;
      RECT  146.18 96.715 146.39 96.385 ;
      RECT  146.18 96.385 146.39 96.005 ;
      RECT  148.37 96.68 148.58 97.09 ;
      RECT  145.97 95.675 146.18 96.005 ;
      RECT  149.015 96.59 149.09 98.295 ;
      RECT  148.93 97.175 149.015 97.585 ;
      RECT  148.01 95.675 148.19 96.59 ;
      POLYGON  149.015 95.675 149.015 96.005 148.58 96.005 148.58 96.385 149.015 96.385 149.015 96.59 149.09 96.59 149.09 95.675 149.015 95.675 ;
      RECT  149.09 96.59 149.3 98.295 ;
      POLYGON  148.58 96.68 148.58 97.09 148.755 97.09 148.835 97.01 148.835 96.68 148.58 96.68 ;
      RECT  145.97 96.59 146.18 98.295 ;
      RECT  147.65 95.675 147.83 96.59 ;
      RECT  146.57 96.59 146.75 98.295 ;
      RECT  148.37 97.67 148.58 98.08 ;
      RECT  149.09 96.385 149.3 96.59 ;
      RECT  146.18 96.59 146.39 98.295 ;
      RECT  148.37 96.005 148.58 96.385 ;
      RECT  146.93 96.59 147.11 98.295 ;
      RECT  147.65 96.59 147.83 98.295 ;
      RECT  146.93 95.675 147.11 96.59 ;
      RECT  149.09 95.675 149.3 96.005 ;
      RECT  147.29 96.59 147.47 98.295 ;
      RECT  147.29 95.675 147.47 96.59 ;
      RECT  145.97 96.385 146.18 96.59 ;
      RECT  149.09 96.005 149.3 96.385 ;
      RECT  148.01 96.59 148.19 98.295 ;
      RECT  146.18 96.385 146.39 96.59 ;
      RECT  145.97 96.005 146.18 96.385 ;
      POLYGON  148.58 97.67 148.58 98.08 148.835 98.08 148.835 97.75 148.755 97.67 148.58 97.67 ;
      RECT  146.57 95.675 146.75 96.59 ;
      RECT  146.18 95.675 146.39 96.005 ;
      RECT  146.18 96.005 146.39 96.385 ;
      RECT  148.37 99.66 148.58 99.25 ;
      RECT  145.97 100.665 146.18 100.335 ;
      RECT  149.015 99.75 149.09 98.045 ;
      RECT  148.93 99.165 149.015 98.755 ;
      RECT  148.01 100.665 148.19 99.75 ;
      POLYGON  149.015 100.665 149.015 100.335 148.58 100.335 148.58 99.955 149.015 99.955 149.015 99.75 149.09 99.75 149.09 100.665 149.015 100.665 ;
      RECT  149.09 99.75 149.3 98.045 ;
      POLYGON  148.58 99.66 148.58 99.25 148.755 99.25 148.835 99.33 148.835 99.66 148.58 99.66 ;
      RECT  145.97 99.75 146.18 98.045 ;
      RECT  147.65 100.665 147.83 99.75 ;
      RECT  146.57 99.75 146.75 98.045 ;
      RECT  148.37 98.67 148.58 98.26 ;
      RECT  149.09 99.955 149.3 99.75 ;
      RECT  146.18 99.75 146.39 98.045 ;
      RECT  148.37 100.335 148.58 99.955 ;
      RECT  146.93 99.75 147.11 98.045 ;
      RECT  147.65 99.75 147.83 98.045 ;
      RECT  146.93 100.665 147.11 99.75 ;
      RECT  149.09 100.665 149.3 100.335 ;
      RECT  147.29 99.75 147.47 98.045 ;
      RECT  147.29 100.665 147.47 99.75 ;
      RECT  145.97 99.955 146.18 99.75 ;
      RECT  149.09 100.335 149.3 99.955 ;
      RECT  148.01 99.75 148.19 98.045 ;
      RECT  146.18 99.955 146.39 99.75 ;
      RECT  145.97 100.335 146.18 99.955 ;
      POLYGON  148.58 98.67 148.58 98.26 148.835 98.26 148.835 98.59 148.755 98.67 148.58 98.67 ;
      RECT  146.57 100.665 146.75 99.75 ;
      RECT  146.18 100.665 146.39 100.335 ;
      RECT  146.18 100.335 146.39 99.955 ;
      RECT  148.37 100.63 148.58 101.04 ;
      RECT  145.97 99.625 146.18 99.955 ;
      RECT  149.015 100.54 149.09 102.245 ;
      RECT  148.93 101.125 149.015 101.535 ;
      RECT  148.01 99.625 148.19 100.54 ;
      POLYGON  149.015 99.625 149.015 99.955 148.58 99.955 148.58 100.335 149.015 100.335 149.015 100.54 149.09 100.54 149.09 99.625 149.015 99.625 ;
      RECT  149.09 100.54 149.3 102.245 ;
      POLYGON  148.58 100.63 148.58 101.04 148.755 101.04 148.835 100.96 148.835 100.63 148.58 100.63 ;
      RECT  145.97 100.54 146.18 102.245 ;
      RECT  147.65 99.625 147.83 100.54 ;
      RECT  146.57 100.54 146.75 102.245 ;
      RECT  148.37 101.62 148.58 102.03 ;
      RECT  149.09 100.335 149.3 100.54 ;
      RECT  146.18 100.54 146.39 102.245 ;
      RECT  148.37 99.955 148.58 100.335 ;
      RECT  146.93 100.54 147.11 102.245 ;
      RECT  147.65 100.54 147.83 102.245 ;
      RECT  146.93 99.625 147.11 100.54 ;
      RECT  149.09 99.625 149.3 99.955 ;
      RECT  147.29 100.54 147.47 102.245 ;
      RECT  147.29 99.625 147.47 100.54 ;
      RECT  145.97 100.335 146.18 100.54 ;
      RECT  149.09 99.955 149.3 100.335 ;
      RECT  148.01 100.54 148.19 102.245 ;
      RECT  146.18 100.335 146.39 100.54 ;
      RECT  145.97 99.955 146.18 100.335 ;
      POLYGON  148.58 101.62 148.58 102.03 148.835 102.03 148.835 101.7 148.755 101.62 148.58 101.62 ;
      RECT  146.57 99.625 146.75 100.54 ;
      RECT  146.18 99.625 146.39 99.955 ;
      RECT  146.18 99.955 146.39 100.335 ;
      RECT  148.37 103.61 148.58 103.2 ;
      RECT  145.97 104.615 146.18 104.285 ;
      RECT  149.015 103.7 149.09 101.995 ;
      RECT  148.93 103.115 149.015 102.705 ;
      RECT  148.01 104.615 148.19 103.7 ;
      POLYGON  149.015 104.615 149.015 104.285 148.58 104.285 148.58 103.905 149.015 103.905 149.015 103.7 149.09 103.7 149.09 104.615 149.015 104.615 ;
      RECT  149.09 103.7 149.3 101.995 ;
      POLYGON  148.58 103.61 148.58 103.2 148.755 103.2 148.835 103.28 148.835 103.61 148.58 103.61 ;
      RECT  145.97 103.7 146.18 101.995 ;
      RECT  147.65 104.615 147.83 103.7 ;
      RECT  146.57 103.7 146.75 101.995 ;
      RECT  148.37 102.62 148.58 102.21 ;
      RECT  149.09 103.905 149.3 103.7 ;
      RECT  146.18 103.7 146.39 101.995 ;
      RECT  148.37 104.285 148.58 103.905 ;
      RECT  146.93 103.7 147.11 101.995 ;
      RECT  147.65 103.7 147.83 101.995 ;
      RECT  146.93 104.615 147.11 103.7 ;
      RECT  149.09 104.615 149.3 104.285 ;
      RECT  147.29 103.7 147.47 101.995 ;
      RECT  147.29 104.615 147.47 103.7 ;
      RECT  145.97 103.905 146.18 103.7 ;
      RECT  149.09 104.285 149.3 103.905 ;
      RECT  148.01 103.7 148.19 101.995 ;
      RECT  146.18 103.905 146.39 103.7 ;
      RECT  145.97 104.285 146.18 103.905 ;
      POLYGON  148.58 102.62 148.58 102.21 148.835 102.21 148.835 102.54 148.755 102.62 148.58 102.62 ;
      RECT  146.57 104.615 146.75 103.7 ;
      RECT  146.18 104.615 146.39 104.285 ;
      RECT  146.18 104.285 146.39 103.905 ;
      RECT  148.37 104.58 148.58 104.99 ;
      RECT  145.97 103.575 146.18 103.905 ;
      RECT  149.015 104.49 149.09 106.195 ;
      RECT  148.93 105.075 149.015 105.485 ;
      RECT  148.01 103.575 148.19 104.49 ;
      POLYGON  149.015 103.575 149.015 103.905 148.58 103.905 148.58 104.285 149.015 104.285 149.015 104.49 149.09 104.49 149.09 103.575 149.015 103.575 ;
      RECT  149.09 104.49 149.3 106.195 ;
      POLYGON  148.58 104.58 148.58 104.99 148.755 104.99 148.835 104.91 148.835 104.58 148.58 104.58 ;
      RECT  145.97 104.49 146.18 106.195 ;
      RECT  147.65 103.575 147.83 104.49 ;
      RECT  146.57 104.49 146.75 106.195 ;
      RECT  148.37 105.57 148.58 105.98 ;
      RECT  149.09 104.285 149.3 104.49 ;
      RECT  146.18 104.49 146.39 106.195 ;
      RECT  148.37 103.905 148.58 104.285 ;
      RECT  146.93 104.49 147.11 106.195 ;
      RECT  147.65 104.49 147.83 106.195 ;
      RECT  146.93 103.575 147.11 104.49 ;
      RECT  149.09 103.575 149.3 103.905 ;
      RECT  147.29 104.49 147.47 106.195 ;
      RECT  147.29 103.575 147.47 104.49 ;
      RECT  145.97 104.285 146.18 104.49 ;
      RECT  149.09 103.905 149.3 104.285 ;
      RECT  148.01 104.49 148.19 106.195 ;
      RECT  146.18 104.285 146.39 104.49 ;
      RECT  145.97 103.905 146.18 104.285 ;
      POLYGON  148.58 105.57 148.58 105.98 148.835 105.98 148.835 105.65 148.755 105.57 148.58 105.57 ;
      RECT  146.57 103.575 146.75 104.49 ;
      RECT  146.18 103.575 146.39 103.905 ;
      RECT  146.18 103.905 146.39 104.285 ;
      RECT  148.37 107.56 148.58 107.15 ;
      RECT  145.97 108.565 146.18 108.235 ;
      RECT  149.015 107.65 149.09 105.945 ;
      RECT  148.93 107.065 149.015 106.655 ;
      RECT  148.01 108.565 148.19 107.65 ;
      POLYGON  149.015 108.565 149.015 108.235 148.58 108.235 148.58 107.855 149.015 107.855 149.015 107.65 149.09 107.65 149.09 108.565 149.015 108.565 ;
      RECT  149.09 107.65 149.3 105.945 ;
      POLYGON  148.58 107.56 148.58 107.15 148.755 107.15 148.835 107.23 148.835 107.56 148.58 107.56 ;
      RECT  145.97 107.65 146.18 105.945 ;
      RECT  147.65 108.565 147.83 107.65 ;
      RECT  146.57 107.65 146.75 105.945 ;
      RECT  148.37 106.57 148.58 106.16 ;
      RECT  149.09 107.855 149.3 107.65 ;
      RECT  146.18 107.65 146.39 105.945 ;
      RECT  148.37 108.235 148.58 107.855 ;
      RECT  146.93 107.65 147.11 105.945 ;
      RECT  147.65 107.65 147.83 105.945 ;
      RECT  146.93 108.565 147.11 107.65 ;
      RECT  149.09 108.565 149.3 108.235 ;
      RECT  147.29 107.65 147.47 105.945 ;
      RECT  147.29 108.565 147.47 107.65 ;
      RECT  145.97 107.855 146.18 107.65 ;
      RECT  149.09 108.235 149.3 107.855 ;
      RECT  148.01 107.65 148.19 105.945 ;
      RECT  146.18 107.855 146.39 107.65 ;
      RECT  145.97 108.235 146.18 107.855 ;
      POLYGON  148.58 106.57 148.58 106.16 148.835 106.16 148.835 106.49 148.755 106.57 148.58 106.57 ;
      RECT  146.57 108.565 146.75 107.65 ;
      RECT  146.18 108.565 146.39 108.235 ;
      RECT  146.18 108.235 146.39 107.855 ;
      RECT  148.37 108.53 148.58 108.94 ;
      RECT  145.97 107.525 146.18 107.855 ;
      RECT  149.015 108.44 149.09 110.145 ;
      RECT  148.93 109.025 149.015 109.435 ;
      RECT  148.01 107.525 148.19 108.44 ;
      POLYGON  149.015 107.525 149.015 107.855 148.58 107.855 148.58 108.235 149.015 108.235 149.015 108.44 149.09 108.44 149.09 107.525 149.015 107.525 ;
      RECT  149.09 108.44 149.3 110.145 ;
      POLYGON  148.58 108.53 148.58 108.94 148.755 108.94 148.835 108.86 148.835 108.53 148.58 108.53 ;
      RECT  145.97 108.44 146.18 110.145 ;
      RECT  147.65 107.525 147.83 108.44 ;
      RECT  146.57 108.44 146.75 110.145 ;
      RECT  148.37 109.52 148.58 109.93 ;
      RECT  149.09 108.235 149.3 108.44 ;
      RECT  146.18 108.44 146.39 110.145 ;
      RECT  148.37 107.855 148.58 108.235 ;
      RECT  146.93 108.44 147.11 110.145 ;
      RECT  147.65 108.44 147.83 110.145 ;
      RECT  146.93 107.525 147.11 108.44 ;
      RECT  149.09 107.525 149.3 107.855 ;
      RECT  147.29 108.44 147.47 110.145 ;
      RECT  147.29 107.525 147.47 108.44 ;
      RECT  145.97 108.235 146.18 108.44 ;
      RECT  149.09 107.855 149.3 108.235 ;
      RECT  148.01 108.44 148.19 110.145 ;
      RECT  146.18 108.235 146.39 108.44 ;
      RECT  145.97 107.855 146.18 108.235 ;
      POLYGON  148.58 109.52 148.58 109.93 148.835 109.93 148.835 109.6 148.755 109.52 148.58 109.52 ;
      RECT  146.57 107.525 146.75 108.44 ;
      RECT  146.18 107.525 146.39 107.855 ;
      RECT  146.18 107.855 146.39 108.235 ;
      RECT  148.37 111.51 148.58 111.1 ;
      RECT  145.97 112.515 146.18 112.185 ;
      RECT  149.015 111.6 149.09 109.895 ;
      RECT  148.93 111.015 149.015 110.605 ;
      RECT  148.01 112.515 148.19 111.6 ;
      POLYGON  149.015 112.515 149.015 112.185 148.58 112.185 148.58 111.805 149.015 111.805 149.015 111.6 149.09 111.6 149.09 112.515 149.015 112.515 ;
      RECT  149.09 111.6 149.3 109.895 ;
      POLYGON  148.58 111.51 148.58 111.1 148.755 111.1 148.835 111.18 148.835 111.51 148.58 111.51 ;
      RECT  145.97 111.6 146.18 109.895 ;
      RECT  147.65 112.515 147.83 111.6 ;
      RECT  146.57 111.6 146.75 109.895 ;
      RECT  148.37 110.52 148.58 110.11 ;
      RECT  149.09 111.805 149.3 111.6 ;
      RECT  146.18 111.6 146.39 109.895 ;
      RECT  148.37 112.185 148.58 111.805 ;
      RECT  146.93 111.6 147.11 109.895 ;
      RECT  147.65 111.6 147.83 109.895 ;
      RECT  146.93 112.515 147.11 111.6 ;
      RECT  149.09 112.515 149.3 112.185 ;
      RECT  147.29 111.6 147.47 109.895 ;
      RECT  147.29 112.515 147.47 111.6 ;
      RECT  145.97 111.805 146.18 111.6 ;
      RECT  149.09 112.185 149.3 111.805 ;
      RECT  148.01 111.6 148.19 109.895 ;
      RECT  146.18 111.805 146.39 111.6 ;
      RECT  145.97 112.185 146.18 111.805 ;
      POLYGON  148.58 110.52 148.58 110.11 148.835 110.11 148.835 110.44 148.755 110.52 148.58 110.52 ;
      RECT  146.57 112.515 146.75 111.6 ;
      RECT  146.18 112.515 146.39 112.185 ;
      RECT  146.18 112.185 146.39 111.805 ;
      RECT  148.37 112.48 148.58 112.89 ;
      RECT  145.97 111.475 146.18 111.805 ;
      RECT  149.015 112.39 149.09 114.095 ;
      RECT  148.93 112.975 149.015 113.385 ;
      RECT  148.01 111.475 148.19 112.39 ;
      POLYGON  149.015 111.475 149.015 111.805 148.58 111.805 148.58 112.185 149.015 112.185 149.015 112.39 149.09 112.39 149.09 111.475 149.015 111.475 ;
      RECT  149.09 112.39 149.3 114.095 ;
      POLYGON  148.58 112.48 148.58 112.89 148.755 112.89 148.835 112.81 148.835 112.48 148.58 112.48 ;
      RECT  145.97 112.39 146.18 114.095 ;
      RECT  147.65 111.475 147.83 112.39 ;
      RECT  146.57 112.39 146.75 114.095 ;
      RECT  148.37 113.47 148.58 113.88 ;
      RECT  149.09 112.185 149.3 112.39 ;
      RECT  146.18 112.39 146.39 114.095 ;
      RECT  148.37 111.805 148.58 112.185 ;
      RECT  146.93 112.39 147.11 114.095 ;
      RECT  147.65 112.39 147.83 114.095 ;
      RECT  146.93 111.475 147.11 112.39 ;
      RECT  149.09 111.475 149.3 111.805 ;
      RECT  147.29 112.39 147.47 114.095 ;
      RECT  147.29 111.475 147.47 112.39 ;
      RECT  145.97 112.185 146.18 112.39 ;
      RECT  149.09 111.805 149.3 112.185 ;
      RECT  148.01 112.39 148.19 114.095 ;
      RECT  146.18 112.185 146.39 112.39 ;
      RECT  145.97 111.805 146.18 112.185 ;
      POLYGON  148.58 113.47 148.58 113.88 148.835 113.88 148.835 113.55 148.755 113.47 148.58 113.47 ;
      RECT  146.57 111.475 146.75 112.39 ;
      RECT  146.18 111.475 146.39 111.805 ;
      RECT  146.18 111.805 146.39 112.185 ;
      RECT  148.37 115.46 148.58 115.05 ;
      RECT  145.97 116.465 146.18 116.135 ;
      RECT  149.015 115.55 149.09 113.845 ;
      RECT  148.93 114.965 149.015 114.555 ;
      RECT  148.01 116.465 148.19 115.55 ;
      POLYGON  149.015 116.465 149.015 116.135 148.58 116.135 148.58 115.755 149.015 115.755 149.015 115.55 149.09 115.55 149.09 116.465 149.015 116.465 ;
      RECT  149.09 115.55 149.3 113.845 ;
      POLYGON  148.58 115.46 148.58 115.05 148.755 115.05 148.835 115.13 148.835 115.46 148.58 115.46 ;
      RECT  145.97 115.55 146.18 113.845 ;
      RECT  147.65 116.465 147.83 115.55 ;
      RECT  146.57 115.55 146.75 113.845 ;
      RECT  148.37 114.47 148.58 114.06 ;
      RECT  149.09 115.755 149.3 115.55 ;
      RECT  146.18 115.55 146.39 113.845 ;
      RECT  148.37 116.135 148.58 115.755 ;
      RECT  146.93 115.55 147.11 113.845 ;
      RECT  147.65 115.55 147.83 113.845 ;
      RECT  146.93 116.465 147.11 115.55 ;
      RECT  149.09 116.465 149.3 116.135 ;
      RECT  147.29 115.55 147.47 113.845 ;
      RECT  147.29 116.465 147.47 115.55 ;
      RECT  145.97 115.755 146.18 115.55 ;
      RECT  149.09 116.135 149.3 115.755 ;
      RECT  148.01 115.55 148.19 113.845 ;
      RECT  146.18 115.755 146.39 115.55 ;
      RECT  145.97 116.135 146.18 115.755 ;
      POLYGON  148.58 114.47 148.58 114.06 148.835 114.06 148.835 114.39 148.755 114.47 148.58 114.47 ;
      RECT  146.57 116.465 146.75 115.55 ;
      RECT  146.18 116.465 146.39 116.135 ;
      RECT  146.18 116.135 146.39 115.755 ;
      RECT  148.37 116.43 148.58 116.84 ;
      RECT  145.97 115.425 146.18 115.755 ;
      RECT  149.015 116.34 149.09 118.045 ;
      RECT  148.93 116.925 149.015 117.335 ;
      RECT  148.01 115.425 148.19 116.34 ;
      POLYGON  149.015 115.425 149.015 115.755 148.58 115.755 148.58 116.135 149.015 116.135 149.015 116.34 149.09 116.34 149.09 115.425 149.015 115.425 ;
      RECT  149.09 116.34 149.3 118.045 ;
      POLYGON  148.58 116.43 148.58 116.84 148.755 116.84 148.835 116.76 148.835 116.43 148.58 116.43 ;
      RECT  145.97 116.34 146.18 118.045 ;
      RECT  147.65 115.425 147.83 116.34 ;
      RECT  146.57 116.34 146.75 118.045 ;
      RECT  148.37 117.42 148.58 117.83 ;
      RECT  149.09 116.135 149.3 116.34 ;
      RECT  146.18 116.34 146.39 118.045 ;
      RECT  148.37 115.755 148.58 116.135 ;
      RECT  146.93 116.34 147.11 118.045 ;
      RECT  147.65 116.34 147.83 118.045 ;
      RECT  146.93 115.425 147.11 116.34 ;
      RECT  149.09 115.425 149.3 115.755 ;
      RECT  147.29 116.34 147.47 118.045 ;
      RECT  147.29 115.425 147.47 116.34 ;
      RECT  145.97 116.135 146.18 116.34 ;
      RECT  149.09 115.755 149.3 116.135 ;
      RECT  148.01 116.34 148.19 118.045 ;
      RECT  146.18 116.135 146.39 116.34 ;
      RECT  145.97 115.755 146.18 116.135 ;
      POLYGON  148.58 117.42 148.58 117.83 148.835 117.83 148.835 117.5 148.755 117.42 148.58 117.42 ;
      RECT  146.57 115.425 146.75 116.34 ;
      RECT  146.18 115.425 146.39 115.755 ;
      RECT  146.18 115.755 146.39 116.135 ;
      RECT  148.37 119.41 148.58 119.0 ;
      RECT  145.97 120.415 146.18 120.085 ;
      RECT  149.015 119.5 149.09 117.795 ;
      RECT  148.93 118.915 149.015 118.505 ;
      RECT  148.01 120.415 148.19 119.5 ;
      POLYGON  149.015 120.415 149.015 120.085 148.58 120.085 148.58 119.705 149.015 119.705 149.015 119.5 149.09 119.5 149.09 120.415 149.015 120.415 ;
      RECT  149.09 119.5 149.3 117.795 ;
      POLYGON  148.58 119.41 148.58 119.0 148.755 119.0 148.835 119.08 148.835 119.41 148.58 119.41 ;
      RECT  145.97 119.5 146.18 117.795 ;
      RECT  147.65 120.415 147.83 119.5 ;
      RECT  146.57 119.5 146.75 117.795 ;
      RECT  148.37 118.42 148.58 118.01 ;
      RECT  149.09 119.705 149.3 119.5 ;
      RECT  146.18 119.5 146.39 117.795 ;
      RECT  148.37 120.085 148.58 119.705 ;
      RECT  146.93 119.5 147.11 117.795 ;
      RECT  147.65 119.5 147.83 117.795 ;
      RECT  146.93 120.415 147.11 119.5 ;
      RECT  149.09 120.415 149.3 120.085 ;
      RECT  147.29 119.5 147.47 117.795 ;
      RECT  147.29 120.415 147.47 119.5 ;
      RECT  145.97 119.705 146.18 119.5 ;
      RECT  149.09 120.085 149.3 119.705 ;
      RECT  148.01 119.5 148.19 117.795 ;
      RECT  146.18 119.705 146.39 119.5 ;
      RECT  145.97 120.085 146.18 119.705 ;
      POLYGON  148.58 118.42 148.58 118.01 148.835 118.01 148.835 118.34 148.755 118.42 148.58 118.42 ;
      RECT  146.57 120.415 146.75 119.5 ;
      RECT  146.18 120.415 146.39 120.085 ;
      RECT  146.18 120.085 146.39 119.705 ;
      RECT  148.37 120.38 148.58 120.79 ;
      RECT  145.97 119.375 146.18 119.705 ;
      RECT  149.015 120.29 149.09 121.995 ;
      RECT  148.93 120.875 149.015 121.285 ;
      RECT  148.01 119.375 148.19 120.29 ;
      POLYGON  149.015 119.375 149.015 119.705 148.58 119.705 148.58 120.085 149.015 120.085 149.015 120.29 149.09 120.29 149.09 119.375 149.015 119.375 ;
      RECT  149.09 120.29 149.3 121.995 ;
      POLYGON  148.58 120.38 148.58 120.79 148.755 120.79 148.835 120.71 148.835 120.38 148.58 120.38 ;
      RECT  145.97 120.29 146.18 121.995 ;
      RECT  147.65 119.375 147.83 120.29 ;
      RECT  146.57 120.29 146.75 121.995 ;
      RECT  148.37 121.37 148.58 121.78 ;
      RECT  149.09 120.085 149.3 120.29 ;
      RECT  146.18 120.29 146.39 121.995 ;
      RECT  148.37 119.705 148.58 120.085 ;
      RECT  146.93 120.29 147.11 121.995 ;
      RECT  147.65 120.29 147.83 121.995 ;
      RECT  146.93 119.375 147.11 120.29 ;
      RECT  149.09 119.375 149.3 119.705 ;
      RECT  147.29 120.29 147.47 121.995 ;
      RECT  147.29 119.375 147.47 120.29 ;
      RECT  145.97 120.085 146.18 120.29 ;
      RECT  149.09 119.705 149.3 120.085 ;
      RECT  148.01 120.29 148.19 121.995 ;
      RECT  146.18 120.085 146.39 120.29 ;
      RECT  145.97 119.705 146.18 120.085 ;
      POLYGON  148.58 121.37 148.58 121.78 148.835 121.78 148.835 121.45 148.755 121.37 148.58 121.37 ;
      RECT  146.57 119.375 146.75 120.29 ;
      RECT  146.18 119.375 146.39 119.705 ;
      RECT  146.18 119.705 146.39 120.085 ;
      RECT  148.37 123.36 148.58 122.95 ;
      RECT  145.97 124.365 146.18 124.035 ;
      RECT  149.015 123.45 149.09 121.745 ;
      RECT  148.93 122.865 149.015 122.455 ;
      RECT  148.01 124.365 148.19 123.45 ;
      POLYGON  149.015 124.365 149.015 124.035 148.58 124.035 148.58 123.655 149.015 123.655 149.015 123.45 149.09 123.45 149.09 124.365 149.015 124.365 ;
      RECT  149.09 123.45 149.3 121.745 ;
      POLYGON  148.58 123.36 148.58 122.95 148.755 122.95 148.835 123.03 148.835 123.36 148.58 123.36 ;
      RECT  145.97 123.45 146.18 121.745 ;
      RECT  147.65 124.365 147.83 123.45 ;
      RECT  146.57 123.45 146.75 121.745 ;
      RECT  148.37 122.37 148.58 121.96 ;
      RECT  149.09 123.655 149.3 123.45 ;
      RECT  146.18 123.45 146.39 121.745 ;
      RECT  148.37 124.035 148.58 123.655 ;
      RECT  146.93 123.45 147.11 121.745 ;
      RECT  147.65 123.45 147.83 121.745 ;
      RECT  146.93 124.365 147.11 123.45 ;
      RECT  149.09 124.365 149.3 124.035 ;
      RECT  147.29 123.45 147.47 121.745 ;
      RECT  147.29 124.365 147.47 123.45 ;
      RECT  145.97 123.655 146.18 123.45 ;
      RECT  149.09 124.035 149.3 123.655 ;
      RECT  148.01 123.45 148.19 121.745 ;
      RECT  146.18 123.655 146.39 123.45 ;
      RECT  145.97 124.035 146.18 123.655 ;
      POLYGON  148.58 122.37 148.58 121.96 148.835 121.96 148.835 122.29 148.755 122.37 148.58 122.37 ;
      RECT  146.57 124.365 146.75 123.45 ;
      RECT  146.18 124.365 146.39 124.035 ;
      RECT  146.18 124.035 146.39 123.655 ;
      RECT  148.37 124.33 148.58 124.74 ;
      RECT  145.97 123.325 146.18 123.655 ;
      RECT  149.015 124.24 149.09 125.945 ;
      RECT  148.93 124.825 149.015 125.235 ;
      RECT  148.01 123.325 148.19 124.24 ;
      POLYGON  149.015 123.325 149.015 123.655 148.58 123.655 148.58 124.035 149.015 124.035 149.015 124.24 149.09 124.24 149.09 123.325 149.015 123.325 ;
      RECT  149.09 124.24 149.3 125.945 ;
      POLYGON  148.58 124.33 148.58 124.74 148.755 124.74 148.835 124.66 148.835 124.33 148.58 124.33 ;
      RECT  145.97 124.24 146.18 125.945 ;
      RECT  147.65 123.325 147.83 124.24 ;
      RECT  146.57 124.24 146.75 125.945 ;
      RECT  148.37 125.32 148.58 125.73 ;
      RECT  149.09 124.035 149.3 124.24 ;
      RECT  146.18 124.24 146.39 125.945 ;
      RECT  148.37 123.655 148.58 124.035 ;
      RECT  146.93 124.24 147.11 125.945 ;
      RECT  147.65 124.24 147.83 125.945 ;
      RECT  146.93 123.325 147.11 124.24 ;
      RECT  149.09 123.325 149.3 123.655 ;
      RECT  147.29 124.24 147.47 125.945 ;
      RECT  147.29 123.325 147.47 124.24 ;
      RECT  145.97 124.035 146.18 124.24 ;
      RECT  149.09 123.655 149.3 124.035 ;
      RECT  148.01 124.24 148.19 125.945 ;
      RECT  146.18 124.035 146.39 124.24 ;
      RECT  145.97 123.655 146.18 124.035 ;
      POLYGON  148.58 125.32 148.58 125.73 148.835 125.73 148.835 125.4 148.755 125.32 148.58 125.32 ;
      RECT  146.57 123.325 146.75 124.24 ;
      RECT  146.18 123.325 146.39 123.655 ;
      RECT  146.18 123.655 146.39 124.035 ;
      RECT  147.65 127.005 147.83 125.425 ;
      RECT  147.29 127.795 147.47 127.005 ;
      RECT  147.25 127.005 147.38 126.295 ;
      RECT  146.93 127.795 147.11 127.005 ;
      RECT  148.01 127.005 148.19 125.425 ;
      RECT  147.65 127.795 147.83 127.005 ;
      RECT  148.01 127.795 148.19 127.005 ;
      RECT  146.57 127.005 146.75 125.425 ;
      RECT  146.57 127.795 146.75 127.005 ;
      RECT  146.93 127.005 147.11 125.425 ;
      RECT  147.38 127.005 147.51 126.295 ;
      RECT  147.29 127.005 147.47 125.425 ;
      RECT  147.29 124.24 147.47 125.945 ;
      RECT  147.29 120.29 147.47 121.995 ;
      RECT  147.29 108.44 147.47 110.145 ;
      RECT  147.29 90.145 147.47 91.85 ;
      RECT  147.29 105.945 147.47 107.65 ;
      RECT  147.29 121.745 147.47 123.45 ;
      RECT  147.29 109.895 147.47 111.6 ;
      RECT  147.29 116.34 147.47 118.045 ;
      RECT  147.29 113.845 147.47 115.55 ;
      RECT  147.29 96.59 147.47 98.295 ;
      RECT  147.29 101.995 147.47 103.7 ;
      RECT  147.29 94.095 147.47 95.8 ;
      RECT  147.29 104.49 147.47 106.195 ;
      RECT  147.29 117.795 147.47 119.5 ;
      RECT  147.29 92.64 147.47 94.345 ;
      RECT  147.29 100.54 147.47 102.245 ;
      RECT  147.29 98.045 147.47 99.75 ;
      RECT  147.29 112.39 147.47 114.095 ;
      RECT  98.45 91.76 98.66 91.35 ;
      RECT  96.05 92.765 96.26 92.435 ;
      RECT  99.095 91.85 99.17 90.145 ;
      RECT  99.01 91.265 99.095 90.855 ;
      RECT  98.09 92.765 98.27 91.85 ;
      POLYGON  99.095 92.765 99.095 92.435 98.66 92.435 98.66 92.055 99.095 92.055 99.095 91.85 99.17 91.85 99.17 92.765 99.095 92.765 ;
      RECT  99.17 91.85 99.38 90.145 ;
      POLYGON  98.66 91.76 98.66 91.35 98.835 91.35 98.915 91.43 98.915 91.76 98.66 91.76 ;
      RECT  96.05 91.85 96.26 90.145 ;
      RECT  97.73 92.765 97.91 91.85 ;
      RECT  96.65 91.85 96.83 90.145 ;
      RECT  98.45 90.77 98.66 90.36 ;
      RECT  99.17 92.055 99.38 91.85 ;
      RECT  96.26 91.85 96.47 90.145 ;
      RECT  98.45 92.435 98.66 92.055 ;
      RECT  97.01 91.85 97.19 90.145 ;
      RECT  97.73 91.85 97.91 90.145 ;
      RECT  97.01 92.765 97.19 91.85 ;
      RECT  99.17 92.765 99.38 92.435 ;
      RECT  97.37 91.85 97.55 90.145 ;
      RECT  97.37 92.765 97.55 91.85 ;
      RECT  96.05 92.055 96.26 91.85 ;
      RECT  99.17 92.435 99.38 92.055 ;
      RECT  98.09 91.85 98.27 90.145 ;
      RECT  96.26 92.055 96.47 91.85 ;
      RECT  96.05 92.435 96.26 92.055 ;
      POLYGON  98.66 90.77 98.66 90.36 98.915 90.36 98.915 90.69 98.835 90.77 98.66 90.77 ;
      RECT  96.65 92.765 96.83 91.85 ;
      RECT  96.26 92.765 96.47 92.435 ;
      RECT  96.26 92.435 96.47 92.055 ;
      RECT  100.31 91.76 100.1 91.35 ;
      RECT  102.71 92.765 102.5 92.435 ;
      RECT  99.665 91.85 99.59 90.145 ;
      RECT  99.75 91.265 99.665 90.855 ;
      RECT  100.67 92.765 100.49 91.85 ;
      POLYGON  99.665 92.765 99.665 92.435 100.1 92.435 100.1 92.055 99.665 92.055 99.665 91.85 99.59 91.85 99.59 92.765 99.665 92.765 ;
      RECT  99.59 91.85 99.38 90.145 ;
      POLYGON  100.1 91.76 100.1 91.35 99.925 91.35 99.845 91.43 99.845 91.76 100.1 91.76 ;
      RECT  102.71 91.85 102.5 90.145 ;
      RECT  101.03 92.765 100.85 91.85 ;
      RECT  102.11 91.85 101.93 90.145 ;
      RECT  100.31 90.77 100.1 90.36 ;
      RECT  99.59 92.055 99.38 91.85 ;
      RECT  102.5 91.85 102.29 90.145 ;
      RECT  100.31 92.435 100.1 92.055 ;
      RECT  101.75 91.85 101.57 90.145 ;
      RECT  101.03 91.85 100.85 90.145 ;
      RECT  101.75 92.765 101.57 91.85 ;
      RECT  99.59 92.765 99.38 92.435 ;
      RECT  101.39 91.85 101.21 90.145 ;
      RECT  101.39 92.765 101.21 91.85 ;
      RECT  102.71 92.055 102.5 91.85 ;
      RECT  99.59 92.435 99.38 92.055 ;
      RECT  100.67 91.85 100.49 90.145 ;
      RECT  102.5 92.055 102.29 91.85 ;
      RECT  102.71 92.435 102.5 92.055 ;
      POLYGON  100.1 90.77 100.1 90.36 99.845 90.36 99.845 90.69 99.925 90.77 100.1 90.77 ;
      RECT  102.11 92.765 101.93 91.85 ;
      RECT  102.5 92.765 102.29 92.435 ;
      RECT  102.5 92.435 102.29 92.055 ;
      RECT  104.69 91.76 104.9 91.35 ;
      RECT  102.29 92.765 102.5 92.435 ;
      RECT  105.335 91.85 105.41 90.145 ;
      RECT  105.25 91.265 105.335 90.855 ;
      RECT  104.33 92.765 104.51 91.85 ;
      POLYGON  105.335 92.765 105.335 92.435 104.9 92.435 104.9 92.055 105.335 92.055 105.335 91.85 105.41 91.85 105.41 92.765 105.335 92.765 ;
      RECT  105.41 91.85 105.62 90.145 ;
      POLYGON  104.9 91.76 104.9 91.35 105.075 91.35 105.155 91.43 105.155 91.76 104.9 91.76 ;
      RECT  102.29 91.85 102.5 90.145 ;
      RECT  103.97 92.765 104.15 91.85 ;
      RECT  102.89 91.85 103.07 90.145 ;
      RECT  104.69 90.77 104.9 90.36 ;
      RECT  105.41 92.055 105.62 91.85 ;
      RECT  102.5 91.85 102.71 90.145 ;
      RECT  104.69 92.435 104.9 92.055 ;
      RECT  103.25 91.85 103.43 90.145 ;
      RECT  103.97 91.85 104.15 90.145 ;
      RECT  103.25 92.765 103.43 91.85 ;
      RECT  105.41 92.765 105.62 92.435 ;
      RECT  103.61 91.85 103.79 90.145 ;
      RECT  103.61 92.765 103.79 91.85 ;
      RECT  102.29 92.055 102.5 91.85 ;
      RECT  105.41 92.435 105.62 92.055 ;
      RECT  104.33 91.85 104.51 90.145 ;
      RECT  102.5 92.055 102.71 91.85 ;
      RECT  102.29 92.435 102.5 92.055 ;
      POLYGON  104.9 90.77 104.9 90.36 105.155 90.36 105.155 90.69 105.075 90.77 104.9 90.77 ;
      RECT  102.89 92.765 103.07 91.85 ;
      RECT  102.5 92.765 102.71 92.435 ;
      RECT  102.5 92.435 102.71 92.055 ;
      RECT  106.55 91.76 106.34 91.35 ;
      RECT  108.95 92.765 108.74 92.435 ;
      RECT  105.905 91.85 105.83 90.145 ;
      RECT  105.99 91.265 105.905 90.855 ;
      RECT  106.91 92.765 106.73 91.85 ;
      POLYGON  105.905 92.765 105.905 92.435 106.34 92.435 106.34 92.055 105.905 92.055 105.905 91.85 105.83 91.85 105.83 92.765 105.905 92.765 ;
      RECT  105.83 91.85 105.62 90.145 ;
      POLYGON  106.34 91.76 106.34 91.35 106.165 91.35 106.085 91.43 106.085 91.76 106.34 91.76 ;
      RECT  108.95 91.85 108.74 90.145 ;
      RECT  107.27 92.765 107.09 91.85 ;
      RECT  108.35 91.85 108.17 90.145 ;
      RECT  106.55 90.77 106.34 90.36 ;
      RECT  105.83 92.055 105.62 91.85 ;
      RECT  108.74 91.85 108.53 90.145 ;
      RECT  106.55 92.435 106.34 92.055 ;
      RECT  107.99 91.85 107.81 90.145 ;
      RECT  107.27 91.85 107.09 90.145 ;
      RECT  107.99 92.765 107.81 91.85 ;
      RECT  105.83 92.765 105.62 92.435 ;
      RECT  107.63 91.85 107.45 90.145 ;
      RECT  107.63 92.765 107.45 91.85 ;
      RECT  108.95 92.055 108.74 91.85 ;
      RECT  105.83 92.435 105.62 92.055 ;
      RECT  106.91 91.85 106.73 90.145 ;
      RECT  108.74 92.055 108.53 91.85 ;
      RECT  108.95 92.435 108.74 92.055 ;
      POLYGON  106.34 90.77 106.34 90.36 106.085 90.36 106.085 90.69 106.165 90.77 106.34 90.77 ;
      RECT  108.35 92.765 108.17 91.85 ;
      RECT  108.74 92.765 108.53 92.435 ;
      RECT  108.74 92.435 108.53 92.055 ;
      RECT  110.93 91.76 111.14 91.35 ;
      RECT  108.53 92.765 108.74 92.435 ;
      RECT  111.575 91.85 111.65 90.145 ;
      RECT  111.49 91.265 111.575 90.855 ;
      RECT  110.57 92.765 110.75 91.85 ;
      POLYGON  111.575 92.765 111.575 92.435 111.14 92.435 111.14 92.055 111.575 92.055 111.575 91.85 111.65 91.85 111.65 92.765 111.575 92.765 ;
      RECT  111.65 91.85 111.86 90.145 ;
      POLYGON  111.14 91.76 111.14 91.35 111.315 91.35 111.395 91.43 111.395 91.76 111.14 91.76 ;
      RECT  108.53 91.85 108.74 90.145 ;
      RECT  110.21 92.765 110.39 91.85 ;
      RECT  109.13 91.85 109.31 90.145 ;
      RECT  110.93 90.77 111.14 90.36 ;
      RECT  111.65 92.055 111.86 91.85 ;
      RECT  108.74 91.85 108.95 90.145 ;
      RECT  110.93 92.435 111.14 92.055 ;
      RECT  109.49 91.85 109.67 90.145 ;
      RECT  110.21 91.85 110.39 90.145 ;
      RECT  109.49 92.765 109.67 91.85 ;
      RECT  111.65 92.765 111.86 92.435 ;
      RECT  109.85 91.85 110.03 90.145 ;
      RECT  109.85 92.765 110.03 91.85 ;
      RECT  108.53 92.055 108.74 91.85 ;
      RECT  111.65 92.435 111.86 92.055 ;
      RECT  110.57 91.85 110.75 90.145 ;
      RECT  108.74 92.055 108.95 91.85 ;
      RECT  108.53 92.435 108.74 92.055 ;
      POLYGON  111.14 90.77 111.14 90.36 111.395 90.36 111.395 90.69 111.315 90.77 111.14 90.77 ;
      RECT  109.13 92.765 109.31 91.85 ;
      RECT  108.74 92.765 108.95 92.435 ;
      RECT  108.74 92.435 108.95 92.055 ;
      RECT  112.79 91.76 112.58 91.35 ;
      RECT  115.19 92.765 114.98 92.435 ;
      RECT  112.145 91.85 112.07 90.145 ;
      RECT  112.23 91.265 112.145 90.855 ;
      RECT  113.15 92.765 112.97 91.85 ;
      POLYGON  112.145 92.765 112.145 92.435 112.58 92.435 112.58 92.055 112.145 92.055 112.145 91.85 112.07 91.85 112.07 92.765 112.145 92.765 ;
      RECT  112.07 91.85 111.86 90.145 ;
      POLYGON  112.58 91.76 112.58 91.35 112.405 91.35 112.325 91.43 112.325 91.76 112.58 91.76 ;
      RECT  115.19 91.85 114.98 90.145 ;
      RECT  113.51 92.765 113.33 91.85 ;
      RECT  114.59 91.85 114.41 90.145 ;
      RECT  112.79 90.77 112.58 90.36 ;
      RECT  112.07 92.055 111.86 91.85 ;
      RECT  114.98 91.85 114.77 90.145 ;
      RECT  112.79 92.435 112.58 92.055 ;
      RECT  114.23 91.85 114.05 90.145 ;
      RECT  113.51 91.85 113.33 90.145 ;
      RECT  114.23 92.765 114.05 91.85 ;
      RECT  112.07 92.765 111.86 92.435 ;
      RECT  113.87 91.85 113.69 90.145 ;
      RECT  113.87 92.765 113.69 91.85 ;
      RECT  115.19 92.055 114.98 91.85 ;
      RECT  112.07 92.435 111.86 92.055 ;
      RECT  113.15 91.85 112.97 90.145 ;
      RECT  114.98 92.055 114.77 91.85 ;
      RECT  115.19 92.435 114.98 92.055 ;
      POLYGON  112.58 90.77 112.58 90.36 112.325 90.36 112.325 90.69 112.405 90.77 112.58 90.77 ;
      RECT  114.59 92.765 114.41 91.85 ;
      RECT  114.98 92.765 114.77 92.435 ;
      RECT  114.98 92.435 114.77 92.055 ;
      RECT  117.17 91.76 117.38 91.35 ;
      RECT  114.77 92.765 114.98 92.435 ;
      RECT  117.815 91.85 117.89 90.145 ;
      RECT  117.73 91.265 117.815 90.855 ;
      RECT  116.81 92.765 116.99 91.85 ;
      POLYGON  117.815 92.765 117.815 92.435 117.38 92.435 117.38 92.055 117.815 92.055 117.815 91.85 117.89 91.85 117.89 92.765 117.815 92.765 ;
      RECT  117.89 91.85 118.1 90.145 ;
      POLYGON  117.38 91.76 117.38 91.35 117.555 91.35 117.635 91.43 117.635 91.76 117.38 91.76 ;
      RECT  114.77 91.85 114.98 90.145 ;
      RECT  116.45 92.765 116.63 91.85 ;
      RECT  115.37 91.85 115.55 90.145 ;
      RECT  117.17 90.77 117.38 90.36 ;
      RECT  117.89 92.055 118.1 91.85 ;
      RECT  114.98 91.85 115.19 90.145 ;
      RECT  117.17 92.435 117.38 92.055 ;
      RECT  115.73 91.85 115.91 90.145 ;
      RECT  116.45 91.85 116.63 90.145 ;
      RECT  115.73 92.765 115.91 91.85 ;
      RECT  117.89 92.765 118.1 92.435 ;
      RECT  116.09 91.85 116.27 90.145 ;
      RECT  116.09 92.765 116.27 91.85 ;
      RECT  114.77 92.055 114.98 91.85 ;
      RECT  117.89 92.435 118.1 92.055 ;
      RECT  116.81 91.85 116.99 90.145 ;
      RECT  114.98 92.055 115.19 91.85 ;
      RECT  114.77 92.435 114.98 92.055 ;
      POLYGON  117.38 90.77 117.38 90.36 117.635 90.36 117.635 90.69 117.555 90.77 117.38 90.77 ;
      RECT  115.37 92.765 115.55 91.85 ;
      RECT  114.98 92.765 115.19 92.435 ;
      RECT  114.98 92.435 115.19 92.055 ;
      RECT  119.03 91.76 118.82 91.35 ;
      RECT  121.43 92.765 121.22 92.435 ;
      RECT  118.385 91.85 118.31 90.145 ;
      RECT  118.47 91.265 118.385 90.855 ;
      RECT  119.39 92.765 119.21 91.85 ;
      POLYGON  118.385 92.765 118.385 92.435 118.82 92.435 118.82 92.055 118.385 92.055 118.385 91.85 118.31 91.85 118.31 92.765 118.385 92.765 ;
      RECT  118.31 91.85 118.1 90.145 ;
      POLYGON  118.82 91.76 118.82 91.35 118.645 91.35 118.565 91.43 118.565 91.76 118.82 91.76 ;
      RECT  121.43 91.85 121.22 90.145 ;
      RECT  119.75 92.765 119.57 91.85 ;
      RECT  120.83 91.85 120.65 90.145 ;
      RECT  119.03 90.77 118.82 90.36 ;
      RECT  118.31 92.055 118.1 91.85 ;
      RECT  121.22 91.85 121.01 90.145 ;
      RECT  119.03 92.435 118.82 92.055 ;
      RECT  120.47 91.85 120.29 90.145 ;
      RECT  119.75 91.85 119.57 90.145 ;
      RECT  120.47 92.765 120.29 91.85 ;
      RECT  118.31 92.765 118.1 92.435 ;
      RECT  120.11 91.85 119.93 90.145 ;
      RECT  120.11 92.765 119.93 91.85 ;
      RECT  121.43 92.055 121.22 91.85 ;
      RECT  118.31 92.435 118.1 92.055 ;
      RECT  119.39 91.85 119.21 90.145 ;
      RECT  121.22 92.055 121.01 91.85 ;
      RECT  121.43 92.435 121.22 92.055 ;
      POLYGON  118.82 90.77 118.82 90.36 118.565 90.36 118.565 90.69 118.645 90.77 118.82 90.77 ;
      RECT  120.83 92.765 120.65 91.85 ;
      RECT  121.22 92.765 121.01 92.435 ;
      RECT  121.22 92.435 121.01 92.055 ;
      RECT  123.41 91.76 123.62 91.35 ;
      RECT  121.01 92.765 121.22 92.435 ;
      RECT  124.055 91.85 124.13 90.145 ;
      RECT  123.97 91.265 124.055 90.855 ;
      RECT  123.05 92.765 123.23 91.85 ;
      POLYGON  124.055 92.765 124.055 92.435 123.62 92.435 123.62 92.055 124.055 92.055 124.055 91.85 124.13 91.85 124.13 92.765 124.055 92.765 ;
      RECT  124.13 91.85 124.34 90.145 ;
      POLYGON  123.62 91.76 123.62 91.35 123.795 91.35 123.875 91.43 123.875 91.76 123.62 91.76 ;
      RECT  121.01 91.85 121.22 90.145 ;
      RECT  122.69 92.765 122.87 91.85 ;
      RECT  121.61 91.85 121.79 90.145 ;
      RECT  123.41 90.77 123.62 90.36 ;
      RECT  124.13 92.055 124.34 91.85 ;
      RECT  121.22 91.85 121.43 90.145 ;
      RECT  123.41 92.435 123.62 92.055 ;
      RECT  121.97 91.85 122.15 90.145 ;
      RECT  122.69 91.85 122.87 90.145 ;
      RECT  121.97 92.765 122.15 91.85 ;
      RECT  124.13 92.765 124.34 92.435 ;
      RECT  122.33 91.85 122.51 90.145 ;
      RECT  122.33 92.765 122.51 91.85 ;
      RECT  121.01 92.055 121.22 91.85 ;
      RECT  124.13 92.435 124.34 92.055 ;
      RECT  123.05 91.85 123.23 90.145 ;
      RECT  121.22 92.055 121.43 91.85 ;
      RECT  121.01 92.435 121.22 92.055 ;
      POLYGON  123.62 90.77 123.62 90.36 123.875 90.36 123.875 90.69 123.795 90.77 123.62 90.77 ;
      RECT  121.61 92.765 121.79 91.85 ;
      RECT  121.22 92.765 121.43 92.435 ;
      RECT  121.22 92.435 121.43 92.055 ;
      RECT  125.27 91.76 125.06 91.35 ;
      RECT  127.67 92.765 127.46 92.435 ;
      RECT  124.625 91.85 124.55 90.145 ;
      RECT  124.71 91.265 124.625 90.855 ;
      RECT  125.63 92.765 125.45 91.85 ;
      POLYGON  124.625 92.765 124.625 92.435 125.06 92.435 125.06 92.055 124.625 92.055 124.625 91.85 124.55 91.85 124.55 92.765 124.625 92.765 ;
      RECT  124.55 91.85 124.34 90.145 ;
      POLYGON  125.06 91.76 125.06 91.35 124.885 91.35 124.805 91.43 124.805 91.76 125.06 91.76 ;
      RECT  127.67 91.85 127.46 90.145 ;
      RECT  125.99 92.765 125.81 91.85 ;
      RECT  127.07 91.85 126.89 90.145 ;
      RECT  125.27 90.77 125.06 90.36 ;
      RECT  124.55 92.055 124.34 91.85 ;
      RECT  127.46 91.85 127.25 90.145 ;
      RECT  125.27 92.435 125.06 92.055 ;
      RECT  126.71 91.85 126.53 90.145 ;
      RECT  125.99 91.85 125.81 90.145 ;
      RECT  126.71 92.765 126.53 91.85 ;
      RECT  124.55 92.765 124.34 92.435 ;
      RECT  126.35 91.85 126.17 90.145 ;
      RECT  126.35 92.765 126.17 91.85 ;
      RECT  127.67 92.055 127.46 91.85 ;
      RECT  124.55 92.435 124.34 92.055 ;
      RECT  125.63 91.85 125.45 90.145 ;
      RECT  127.46 92.055 127.25 91.85 ;
      RECT  127.67 92.435 127.46 92.055 ;
      POLYGON  125.06 90.77 125.06 90.36 124.805 90.36 124.805 90.69 124.885 90.77 125.06 90.77 ;
      RECT  127.07 92.765 126.89 91.85 ;
      RECT  127.46 92.765 127.25 92.435 ;
      RECT  127.46 92.435 127.25 92.055 ;
      RECT  129.65 91.76 129.86 91.35 ;
      RECT  127.25 92.765 127.46 92.435 ;
      RECT  130.295 91.85 130.37 90.145 ;
      RECT  130.21 91.265 130.295 90.855 ;
      RECT  129.29 92.765 129.47 91.85 ;
      POLYGON  130.295 92.765 130.295 92.435 129.86 92.435 129.86 92.055 130.295 92.055 130.295 91.85 130.37 91.85 130.37 92.765 130.295 92.765 ;
      RECT  130.37 91.85 130.58 90.145 ;
      POLYGON  129.86 91.76 129.86 91.35 130.035 91.35 130.115 91.43 130.115 91.76 129.86 91.76 ;
      RECT  127.25 91.85 127.46 90.145 ;
      RECT  128.93 92.765 129.11 91.85 ;
      RECT  127.85 91.85 128.03 90.145 ;
      RECT  129.65 90.77 129.86 90.36 ;
      RECT  130.37 92.055 130.58 91.85 ;
      RECT  127.46 91.85 127.67 90.145 ;
      RECT  129.65 92.435 129.86 92.055 ;
      RECT  128.21 91.85 128.39 90.145 ;
      RECT  128.93 91.85 129.11 90.145 ;
      RECT  128.21 92.765 128.39 91.85 ;
      RECT  130.37 92.765 130.58 92.435 ;
      RECT  128.57 91.85 128.75 90.145 ;
      RECT  128.57 92.765 128.75 91.85 ;
      RECT  127.25 92.055 127.46 91.85 ;
      RECT  130.37 92.435 130.58 92.055 ;
      RECT  129.29 91.85 129.47 90.145 ;
      RECT  127.46 92.055 127.67 91.85 ;
      RECT  127.25 92.435 127.46 92.055 ;
      POLYGON  129.86 90.77 129.86 90.36 130.115 90.36 130.115 90.69 130.035 90.77 129.86 90.77 ;
      RECT  127.85 92.765 128.03 91.85 ;
      RECT  127.46 92.765 127.67 92.435 ;
      RECT  127.46 92.435 127.67 92.055 ;
      RECT  131.51 91.76 131.3 91.35 ;
      RECT  133.91 92.765 133.7 92.435 ;
      RECT  130.865 91.85 130.79 90.145 ;
      RECT  130.95 91.265 130.865 90.855 ;
      RECT  131.87 92.765 131.69 91.85 ;
      POLYGON  130.865 92.765 130.865 92.435 131.3 92.435 131.3 92.055 130.865 92.055 130.865 91.85 130.79 91.85 130.79 92.765 130.865 92.765 ;
      RECT  130.79 91.85 130.58 90.145 ;
      POLYGON  131.3 91.76 131.3 91.35 131.125 91.35 131.045 91.43 131.045 91.76 131.3 91.76 ;
      RECT  133.91 91.85 133.7 90.145 ;
      RECT  132.23 92.765 132.05 91.85 ;
      RECT  133.31 91.85 133.13 90.145 ;
      RECT  131.51 90.77 131.3 90.36 ;
      RECT  130.79 92.055 130.58 91.85 ;
      RECT  133.7 91.85 133.49 90.145 ;
      RECT  131.51 92.435 131.3 92.055 ;
      RECT  132.95 91.85 132.77 90.145 ;
      RECT  132.23 91.85 132.05 90.145 ;
      RECT  132.95 92.765 132.77 91.85 ;
      RECT  130.79 92.765 130.58 92.435 ;
      RECT  132.59 91.85 132.41 90.145 ;
      RECT  132.59 92.765 132.41 91.85 ;
      RECT  133.91 92.055 133.7 91.85 ;
      RECT  130.79 92.435 130.58 92.055 ;
      RECT  131.87 91.85 131.69 90.145 ;
      RECT  133.7 92.055 133.49 91.85 ;
      RECT  133.91 92.435 133.7 92.055 ;
      POLYGON  131.3 90.77 131.3 90.36 131.045 90.36 131.045 90.69 131.125 90.77 131.3 90.77 ;
      RECT  133.31 92.765 133.13 91.85 ;
      RECT  133.7 92.765 133.49 92.435 ;
      RECT  133.7 92.435 133.49 92.055 ;
      RECT  135.89 91.76 136.1 91.35 ;
      RECT  133.49 92.765 133.7 92.435 ;
      RECT  136.535 91.85 136.61 90.145 ;
      RECT  136.45 91.265 136.535 90.855 ;
      RECT  135.53 92.765 135.71 91.85 ;
      POLYGON  136.535 92.765 136.535 92.435 136.1 92.435 136.1 92.055 136.535 92.055 136.535 91.85 136.61 91.85 136.61 92.765 136.535 92.765 ;
      RECT  136.61 91.85 136.82 90.145 ;
      POLYGON  136.1 91.76 136.1 91.35 136.275 91.35 136.355 91.43 136.355 91.76 136.1 91.76 ;
      RECT  133.49 91.85 133.7 90.145 ;
      RECT  135.17 92.765 135.35 91.85 ;
      RECT  134.09 91.85 134.27 90.145 ;
      RECT  135.89 90.77 136.1 90.36 ;
      RECT  136.61 92.055 136.82 91.85 ;
      RECT  133.7 91.85 133.91 90.145 ;
      RECT  135.89 92.435 136.1 92.055 ;
      RECT  134.45 91.85 134.63 90.145 ;
      RECT  135.17 91.85 135.35 90.145 ;
      RECT  134.45 92.765 134.63 91.85 ;
      RECT  136.61 92.765 136.82 92.435 ;
      RECT  134.81 91.85 134.99 90.145 ;
      RECT  134.81 92.765 134.99 91.85 ;
      RECT  133.49 92.055 133.7 91.85 ;
      RECT  136.61 92.435 136.82 92.055 ;
      RECT  135.53 91.85 135.71 90.145 ;
      RECT  133.7 92.055 133.91 91.85 ;
      RECT  133.49 92.435 133.7 92.055 ;
      POLYGON  136.1 90.77 136.1 90.36 136.355 90.36 136.355 90.69 136.275 90.77 136.1 90.77 ;
      RECT  134.09 92.765 134.27 91.85 ;
      RECT  133.7 92.765 133.91 92.435 ;
      RECT  133.7 92.435 133.91 92.055 ;
      RECT  137.75 91.76 137.54 91.35 ;
      RECT  140.15 92.765 139.94 92.435 ;
      RECT  137.105 91.85 137.03 90.145 ;
      RECT  137.19 91.265 137.105 90.855 ;
      RECT  138.11 92.765 137.93 91.85 ;
      POLYGON  137.105 92.765 137.105 92.435 137.54 92.435 137.54 92.055 137.105 92.055 137.105 91.85 137.03 91.85 137.03 92.765 137.105 92.765 ;
      RECT  137.03 91.85 136.82 90.145 ;
      POLYGON  137.54 91.76 137.54 91.35 137.365 91.35 137.285 91.43 137.285 91.76 137.54 91.76 ;
      RECT  140.15 91.85 139.94 90.145 ;
      RECT  138.47 92.765 138.29 91.85 ;
      RECT  139.55 91.85 139.37 90.145 ;
      RECT  137.75 90.77 137.54 90.36 ;
      RECT  137.03 92.055 136.82 91.85 ;
      RECT  139.94 91.85 139.73 90.145 ;
      RECT  137.75 92.435 137.54 92.055 ;
      RECT  139.19 91.85 139.01 90.145 ;
      RECT  138.47 91.85 138.29 90.145 ;
      RECT  139.19 92.765 139.01 91.85 ;
      RECT  137.03 92.765 136.82 92.435 ;
      RECT  138.83 91.85 138.65 90.145 ;
      RECT  138.83 92.765 138.65 91.85 ;
      RECT  140.15 92.055 139.94 91.85 ;
      RECT  137.03 92.435 136.82 92.055 ;
      RECT  138.11 91.85 137.93 90.145 ;
      RECT  139.94 92.055 139.73 91.85 ;
      RECT  140.15 92.435 139.94 92.055 ;
      POLYGON  137.54 90.77 137.54 90.36 137.285 90.36 137.285 90.69 137.365 90.77 137.54 90.77 ;
      RECT  139.55 92.765 139.37 91.85 ;
      RECT  139.94 92.765 139.73 92.435 ;
      RECT  139.94 92.435 139.73 92.055 ;
      RECT  142.13 91.76 142.34 91.35 ;
      RECT  139.73 92.765 139.94 92.435 ;
      RECT  142.775 91.85 142.85 90.145 ;
      RECT  142.69 91.265 142.775 90.855 ;
      RECT  141.77 92.765 141.95 91.85 ;
      POLYGON  142.775 92.765 142.775 92.435 142.34 92.435 142.34 92.055 142.775 92.055 142.775 91.85 142.85 91.85 142.85 92.765 142.775 92.765 ;
      RECT  142.85 91.85 143.06 90.145 ;
      POLYGON  142.34 91.76 142.34 91.35 142.515 91.35 142.595 91.43 142.595 91.76 142.34 91.76 ;
      RECT  139.73 91.85 139.94 90.145 ;
      RECT  141.41 92.765 141.59 91.85 ;
      RECT  140.33 91.85 140.51 90.145 ;
      RECT  142.13 90.77 142.34 90.36 ;
      RECT  142.85 92.055 143.06 91.85 ;
      RECT  139.94 91.85 140.15 90.145 ;
      RECT  142.13 92.435 142.34 92.055 ;
      RECT  140.69 91.85 140.87 90.145 ;
      RECT  141.41 91.85 141.59 90.145 ;
      RECT  140.69 92.765 140.87 91.85 ;
      RECT  142.85 92.765 143.06 92.435 ;
      RECT  141.05 91.85 141.23 90.145 ;
      RECT  141.05 92.765 141.23 91.85 ;
      RECT  139.73 92.055 139.94 91.85 ;
      RECT  142.85 92.435 143.06 92.055 ;
      RECT  141.77 91.85 141.95 90.145 ;
      RECT  139.94 92.055 140.15 91.85 ;
      RECT  139.73 92.435 139.94 92.055 ;
      POLYGON  142.34 90.77 142.34 90.36 142.595 90.36 142.595 90.69 142.515 90.77 142.34 90.77 ;
      RECT  140.33 92.765 140.51 91.85 ;
      RECT  139.94 92.765 140.15 92.435 ;
      RECT  139.94 92.435 140.15 92.055 ;
      RECT  143.99 91.76 143.78 91.35 ;
      RECT  146.39 92.765 146.18 92.435 ;
      RECT  143.345 91.85 143.27 90.145 ;
      RECT  143.43 91.265 143.345 90.855 ;
      RECT  144.35 92.765 144.17 91.85 ;
      POLYGON  143.345 92.765 143.345 92.435 143.78 92.435 143.78 92.055 143.345 92.055 143.345 91.85 143.27 91.85 143.27 92.765 143.345 92.765 ;
      RECT  143.27 91.85 143.06 90.145 ;
      POLYGON  143.78 91.76 143.78 91.35 143.605 91.35 143.525 91.43 143.525 91.76 143.78 91.76 ;
      RECT  146.39 91.85 146.18 90.145 ;
      RECT  144.71 92.765 144.53 91.85 ;
      RECT  145.79 91.85 145.61 90.145 ;
      RECT  143.99 90.77 143.78 90.36 ;
      RECT  143.27 92.055 143.06 91.85 ;
      RECT  146.18 91.85 145.97 90.145 ;
      RECT  143.99 92.435 143.78 92.055 ;
      RECT  145.43 91.85 145.25 90.145 ;
      RECT  144.71 91.85 144.53 90.145 ;
      RECT  145.43 92.765 145.25 91.85 ;
      RECT  143.27 92.765 143.06 92.435 ;
      RECT  145.07 91.85 144.89 90.145 ;
      RECT  145.07 92.765 144.89 91.85 ;
      RECT  146.39 92.055 146.18 91.85 ;
      RECT  143.27 92.435 143.06 92.055 ;
      RECT  144.35 91.85 144.17 90.145 ;
      RECT  146.18 92.055 145.97 91.85 ;
      RECT  146.39 92.435 146.18 92.055 ;
      POLYGON  143.78 90.77 143.78 90.36 143.525 90.36 143.525 90.69 143.605 90.77 143.78 90.77 ;
      RECT  145.79 92.765 145.61 91.85 ;
      RECT  146.18 92.765 145.97 92.435 ;
      RECT  146.18 92.435 145.97 92.055 ;
      RECT  96.65 92.245 96.83 90.27 ;
      RECT  97.01 92.245 97.19 90.27 ;
      RECT  97.73 92.245 97.91 90.27 ;
      RECT  98.09 92.245 98.27 90.27 ;
      RECT  101.93 92.245 102.11 90.27 ;
      RECT  101.57 92.245 101.75 90.27 ;
      RECT  100.85 92.245 101.03 90.27 ;
      RECT  100.49 92.245 100.67 90.27 ;
      RECT  102.89 92.245 103.07 90.27 ;
      RECT  103.25 92.245 103.43 90.27 ;
      RECT  103.97 92.245 104.15 90.27 ;
      RECT  104.33 92.245 104.51 90.27 ;
      RECT  108.17 92.245 108.35 90.27 ;
      RECT  107.81 92.245 107.99 90.27 ;
      RECT  107.09 92.245 107.27 90.27 ;
      RECT  106.73 92.245 106.91 90.27 ;
      RECT  109.13 92.245 109.31 90.27 ;
      RECT  109.49 92.245 109.67 90.27 ;
      RECT  110.21 92.245 110.39 90.27 ;
      RECT  110.57 92.245 110.75 90.27 ;
      RECT  114.41 92.245 114.59 90.27 ;
      RECT  114.05 92.245 114.23 90.27 ;
      RECT  113.33 92.245 113.51 90.27 ;
      RECT  112.97 92.245 113.15 90.27 ;
      RECT  115.37 92.245 115.55 90.27 ;
      RECT  115.73 92.245 115.91 90.27 ;
      RECT  116.45 92.245 116.63 90.27 ;
      RECT  116.81 92.245 116.99 90.27 ;
      RECT  120.65 92.245 120.83 90.27 ;
      RECT  120.29 92.245 120.47 90.27 ;
      RECT  119.57 92.245 119.75 90.27 ;
      RECT  119.21 92.245 119.39 90.27 ;
      RECT  121.61 92.245 121.79 90.27 ;
      RECT  121.97 92.245 122.15 90.27 ;
      RECT  122.69 92.245 122.87 90.27 ;
      RECT  123.05 92.245 123.23 90.27 ;
      RECT  126.89 92.245 127.07 90.27 ;
      RECT  126.53 92.245 126.71 90.27 ;
      RECT  125.81 92.245 125.99 90.27 ;
      RECT  125.45 92.245 125.63 90.27 ;
      RECT  127.85 92.245 128.03 90.27 ;
      RECT  128.21 92.245 128.39 90.27 ;
      RECT  128.93 92.245 129.11 90.27 ;
      RECT  129.29 92.245 129.47 90.27 ;
      RECT  133.13 92.245 133.31 90.27 ;
      RECT  132.77 92.245 132.95 90.27 ;
      RECT  132.05 92.245 132.23 90.27 ;
      RECT  131.69 92.245 131.87 90.27 ;
      RECT  134.09 92.245 134.27 90.27 ;
      RECT  134.45 92.245 134.63 90.27 ;
      RECT  135.17 92.245 135.35 90.27 ;
      RECT  135.53 92.245 135.71 90.27 ;
      RECT  139.37 92.245 139.55 90.27 ;
      RECT  139.01 92.245 139.19 90.27 ;
      RECT  138.29 92.245 138.47 90.27 ;
      RECT  137.93 92.245 138.11 90.27 ;
      RECT  140.33 92.245 140.51 90.27 ;
      RECT  140.69 92.245 140.87 90.27 ;
      RECT  141.41 92.245 141.59 90.27 ;
      RECT  141.77 92.245 141.95 90.27 ;
      RECT  145.61 92.245 145.79 90.27 ;
      RECT  145.25 92.245 145.43 90.27 ;
      RECT  144.53 92.245 144.71 90.27 ;
      RECT  144.17 92.245 144.35 90.27 ;
      RECT  109.85 91.85 110.03 90.145 ;
      RECT  144.89 91.85 145.07 90.145 ;
      RECT  113.69 91.85 113.87 90.145 ;
      RECT  138.65 91.85 138.83 90.145 ;
      RECT  126.17 91.85 126.35 90.145 ;
      RECT  107.45 91.85 107.63 90.145 ;
      RECT  101.21 91.85 101.39 90.145 ;
      RECT  116.09 91.85 116.27 90.145 ;
      RECT  119.93 91.85 120.11 90.145 ;
      RECT  134.81 91.85 134.99 90.145 ;
      RECT  103.61 91.85 103.79 90.145 ;
      RECT  122.33 91.85 122.51 90.145 ;
      RECT  97.37 91.85 97.55 90.145 ;
      RECT  132.41 91.85 132.59 90.145 ;
      RECT  128.57 91.85 128.75 90.145 ;
      RECT  141.05 91.85 141.23 90.145 ;
      RECT  98.45 124.33 98.66 124.74 ;
      RECT  96.05 123.325 96.26 123.655 ;
      RECT  99.095 124.24 99.17 125.945 ;
      RECT  99.01 124.825 99.095 125.235 ;
      RECT  98.09 123.325 98.27 124.24 ;
      POLYGON  99.095 123.325 99.095 123.655 98.66 123.655 98.66 124.035 99.095 124.035 99.095 124.24 99.17 124.24 99.17 123.325 99.095 123.325 ;
      RECT  99.17 124.24 99.38 125.945 ;
      POLYGON  98.66 124.33 98.66 124.74 98.835 124.74 98.915 124.66 98.915 124.33 98.66 124.33 ;
      RECT  96.05 124.24 96.26 125.945 ;
      RECT  97.73 123.325 97.91 124.24 ;
      RECT  96.65 124.24 96.83 125.945 ;
      RECT  98.45 125.32 98.66 125.73 ;
      RECT  99.17 124.035 99.38 124.24 ;
      RECT  96.26 124.24 96.47 125.945 ;
      RECT  98.45 123.655 98.66 124.035 ;
      RECT  97.01 124.24 97.19 125.945 ;
      RECT  97.73 124.24 97.91 125.945 ;
      RECT  97.01 123.325 97.19 124.24 ;
      RECT  99.17 123.325 99.38 123.655 ;
      RECT  97.37 124.24 97.55 125.945 ;
      RECT  97.37 123.325 97.55 124.24 ;
      RECT  96.05 124.035 96.26 124.24 ;
      RECT  99.17 123.655 99.38 124.035 ;
      RECT  98.09 124.24 98.27 125.945 ;
      RECT  96.26 124.035 96.47 124.24 ;
      RECT  96.05 123.655 96.26 124.035 ;
      POLYGON  98.66 125.32 98.66 125.73 98.915 125.73 98.915 125.4 98.835 125.32 98.66 125.32 ;
      RECT  96.65 123.325 96.83 124.24 ;
      RECT  96.26 123.325 96.47 123.655 ;
      RECT  96.26 123.655 96.47 124.035 ;
      RECT  100.31 124.33 100.1 124.74 ;
      RECT  102.71 123.325 102.5 123.655 ;
      RECT  99.665 124.24 99.59 125.945 ;
      RECT  99.75 124.825 99.665 125.235 ;
      RECT  100.67 123.325 100.49 124.24 ;
      POLYGON  99.665 123.325 99.665 123.655 100.1 123.655 100.1 124.035 99.665 124.035 99.665 124.24 99.59 124.24 99.59 123.325 99.665 123.325 ;
      RECT  99.59 124.24 99.38 125.945 ;
      POLYGON  100.1 124.33 100.1 124.74 99.925 124.74 99.845 124.66 99.845 124.33 100.1 124.33 ;
      RECT  102.71 124.24 102.5 125.945 ;
      RECT  101.03 123.325 100.85 124.24 ;
      RECT  102.11 124.24 101.93 125.945 ;
      RECT  100.31 125.32 100.1 125.73 ;
      RECT  99.59 124.035 99.38 124.24 ;
      RECT  102.5 124.24 102.29 125.945 ;
      RECT  100.31 123.655 100.1 124.035 ;
      RECT  101.75 124.24 101.57 125.945 ;
      RECT  101.03 124.24 100.85 125.945 ;
      RECT  101.75 123.325 101.57 124.24 ;
      RECT  99.59 123.325 99.38 123.655 ;
      RECT  101.39 124.24 101.21 125.945 ;
      RECT  101.39 123.325 101.21 124.24 ;
      RECT  102.71 124.035 102.5 124.24 ;
      RECT  99.59 123.655 99.38 124.035 ;
      RECT  100.67 124.24 100.49 125.945 ;
      RECT  102.5 124.035 102.29 124.24 ;
      RECT  102.71 123.655 102.5 124.035 ;
      POLYGON  100.1 125.32 100.1 125.73 99.845 125.73 99.845 125.4 99.925 125.32 100.1 125.32 ;
      RECT  102.11 123.325 101.93 124.24 ;
      RECT  102.5 123.325 102.29 123.655 ;
      RECT  102.5 123.655 102.29 124.035 ;
      RECT  104.69 124.33 104.9 124.74 ;
      RECT  102.29 123.325 102.5 123.655 ;
      RECT  105.335 124.24 105.41 125.945 ;
      RECT  105.25 124.825 105.335 125.235 ;
      RECT  104.33 123.325 104.51 124.24 ;
      POLYGON  105.335 123.325 105.335 123.655 104.9 123.655 104.9 124.035 105.335 124.035 105.335 124.24 105.41 124.24 105.41 123.325 105.335 123.325 ;
      RECT  105.41 124.24 105.62 125.945 ;
      POLYGON  104.9 124.33 104.9 124.74 105.075 124.74 105.155 124.66 105.155 124.33 104.9 124.33 ;
      RECT  102.29 124.24 102.5 125.945 ;
      RECT  103.97 123.325 104.15 124.24 ;
      RECT  102.89 124.24 103.07 125.945 ;
      RECT  104.69 125.32 104.9 125.73 ;
      RECT  105.41 124.035 105.62 124.24 ;
      RECT  102.5 124.24 102.71 125.945 ;
      RECT  104.69 123.655 104.9 124.035 ;
      RECT  103.25 124.24 103.43 125.945 ;
      RECT  103.97 124.24 104.15 125.945 ;
      RECT  103.25 123.325 103.43 124.24 ;
      RECT  105.41 123.325 105.62 123.655 ;
      RECT  103.61 124.24 103.79 125.945 ;
      RECT  103.61 123.325 103.79 124.24 ;
      RECT  102.29 124.035 102.5 124.24 ;
      RECT  105.41 123.655 105.62 124.035 ;
      RECT  104.33 124.24 104.51 125.945 ;
      RECT  102.5 124.035 102.71 124.24 ;
      RECT  102.29 123.655 102.5 124.035 ;
      POLYGON  104.9 125.32 104.9 125.73 105.155 125.73 105.155 125.4 105.075 125.32 104.9 125.32 ;
      RECT  102.89 123.325 103.07 124.24 ;
      RECT  102.5 123.325 102.71 123.655 ;
      RECT  102.5 123.655 102.71 124.035 ;
      RECT  106.55 124.33 106.34 124.74 ;
      RECT  108.95 123.325 108.74 123.655 ;
      RECT  105.905 124.24 105.83 125.945 ;
      RECT  105.99 124.825 105.905 125.235 ;
      RECT  106.91 123.325 106.73 124.24 ;
      POLYGON  105.905 123.325 105.905 123.655 106.34 123.655 106.34 124.035 105.905 124.035 105.905 124.24 105.83 124.24 105.83 123.325 105.905 123.325 ;
      RECT  105.83 124.24 105.62 125.945 ;
      POLYGON  106.34 124.33 106.34 124.74 106.165 124.74 106.085 124.66 106.085 124.33 106.34 124.33 ;
      RECT  108.95 124.24 108.74 125.945 ;
      RECT  107.27 123.325 107.09 124.24 ;
      RECT  108.35 124.24 108.17 125.945 ;
      RECT  106.55 125.32 106.34 125.73 ;
      RECT  105.83 124.035 105.62 124.24 ;
      RECT  108.74 124.24 108.53 125.945 ;
      RECT  106.55 123.655 106.34 124.035 ;
      RECT  107.99 124.24 107.81 125.945 ;
      RECT  107.27 124.24 107.09 125.945 ;
      RECT  107.99 123.325 107.81 124.24 ;
      RECT  105.83 123.325 105.62 123.655 ;
      RECT  107.63 124.24 107.45 125.945 ;
      RECT  107.63 123.325 107.45 124.24 ;
      RECT  108.95 124.035 108.74 124.24 ;
      RECT  105.83 123.655 105.62 124.035 ;
      RECT  106.91 124.24 106.73 125.945 ;
      RECT  108.74 124.035 108.53 124.24 ;
      RECT  108.95 123.655 108.74 124.035 ;
      POLYGON  106.34 125.32 106.34 125.73 106.085 125.73 106.085 125.4 106.165 125.32 106.34 125.32 ;
      RECT  108.35 123.325 108.17 124.24 ;
      RECT  108.74 123.325 108.53 123.655 ;
      RECT  108.74 123.655 108.53 124.035 ;
      RECT  110.93 124.33 111.14 124.74 ;
      RECT  108.53 123.325 108.74 123.655 ;
      RECT  111.575 124.24 111.65 125.945 ;
      RECT  111.49 124.825 111.575 125.235 ;
      RECT  110.57 123.325 110.75 124.24 ;
      POLYGON  111.575 123.325 111.575 123.655 111.14 123.655 111.14 124.035 111.575 124.035 111.575 124.24 111.65 124.24 111.65 123.325 111.575 123.325 ;
      RECT  111.65 124.24 111.86 125.945 ;
      POLYGON  111.14 124.33 111.14 124.74 111.315 124.74 111.395 124.66 111.395 124.33 111.14 124.33 ;
      RECT  108.53 124.24 108.74 125.945 ;
      RECT  110.21 123.325 110.39 124.24 ;
      RECT  109.13 124.24 109.31 125.945 ;
      RECT  110.93 125.32 111.14 125.73 ;
      RECT  111.65 124.035 111.86 124.24 ;
      RECT  108.74 124.24 108.95 125.945 ;
      RECT  110.93 123.655 111.14 124.035 ;
      RECT  109.49 124.24 109.67 125.945 ;
      RECT  110.21 124.24 110.39 125.945 ;
      RECT  109.49 123.325 109.67 124.24 ;
      RECT  111.65 123.325 111.86 123.655 ;
      RECT  109.85 124.24 110.03 125.945 ;
      RECT  109.85 123.325 110.03 124.24 ;
      RECT  108.53 124.035 108.74 124.24 ;
      RECT  111.65 123.655 111.86 124.035 ;
      RECT  110.57 124.24 110.75 125.945 ;
      RECT  108.74 124.035 108.95 124.24 ;
      RECT  108.53 123.655 108.74 124.035 ;
      POLYGON  111.14 125.32 111.14 125.73 111.395 125.73 111.395 125.4 111.315 125.32 111.14 125.32 ;
      RECT  109.13 123.325 109.31 124.24 ;
      RECT  108.74 123.325 108.95 123.655 ;
      RECT  108.74 123.655 108.95 124.035 ;
      RECT  112.79 124.33 112.58 124.74 ;
      RECT  115.19 123.325 114.98 123.655 ;
      RECT  112.145 124.24 112.07 125.945 ;
      RECT  112.23 124.825 112.145 125.235 ;
      RECT  113.15 123.325 112.97 124.24 ;
      POLYGON  112.145 123.325 112.145 123.655 112.58 123.655 112.58 124.035 112.145 124.035 112.145 124.24 112.07 124.24 112.07 123.325 112.145 123.325 ;
      RECT  112.07 124.24 111.86 125.945 ;
      POLYGON  112.58 124.33 112.58 124.74 112.405 124.74 112.325 124.66 112.325 124.33 112.58 124.33 ;
      RECT  115.19 124.24 114.98 125.945 ;
      RECT  113.51 123.325 113.33 124.24 ;
      RECT  114.59 124.24 114.41 125.945 ;
      RECT  112.79 125.32 112.58 125.73 ;
      RECT  112.07 124.035 111.86 124.24 ;
      RECT  114.98 124.24 114.77 125.945 ;
      RECT  112.79 123.655 112.58 124.035 ;
      RECT  114.23 124.24 114.05 125.945 ;
      RECT  113.51 124.24 113.33 125.945 ;
      RECT  114.23 123.325 114.05 124.24 ;
      RECT  112.07 123.325 111.86 123.655 ;
      RECT  113.87 124.24 113.69 125.945 ;
      RECT  113.87 123.325 113.69 124.24 ;
      RECT  115.19 124.035 114.98 124.24 ;
      RECT  112.07 123.655 111.86 124.035 ;
      RECT  113.15 124.24 112.97 125.945 ;
      RECT  114.98 124.035 114.77 124.24 ;
      RECT  115.19 123.655 114.98 124.035 ;
      POLYGON  112.58 125.32 112.58 125.73 112.325 125.73 112.325 125.4 112.405 125.32 112.58 125.32 ;
      RECT  114.59 123.325 114.41 124.24 ;
      RECT  114.98 123.325 114.77 123.655 ;
      RECT  114.98 123.655 114.77 124.035 ;
      RECT  117.17 124.33 117.38 124.74 ;
      RECT  114.77 123.325 114.98 123.655 ;
      RECT  117.815 124.24 117.89 125.945 ;
      RECT  117.73 124.825 117.815 125.235 ;
      RECT  116.81 123.325 116.99 124.24 ;
      POLYGON  117.815 123.325 117.815 123.655 117.38 123.655 117.38 124.035 117.815 124.035 117.815 124.24 117.89 124.24 117.89 123.325 117.815 123.325 ;
      RECT  117.89 124.24 118.1 125.945 ;
      POLYGON  117.38 124.33 117.38 124.74 117.555 124.74 117.635 124.66 117.635 124.33 117.38 124.33 ;
      RECT  114.77 124.24 114.98 125.945 ;
      RECT  116.45 123.325 116.63 124.24 ;
      RECT  115.37 124.24 115.55 125.945 ;
      RECT  117.17 125.32 117.38 125.73 ;
      RECT  117.89 124.035 118.1 124.24 ;
      RECT  114.98 124.24 115.19 125.945 ;
      RECT  117.17 123.655 117.38 124.035 ;
      RECT  115.73 124.24 115.91 125.945 ;
      RECT  116.45 124.24 116.63 125.945 ;
      RECT  115.73 123.325 115.91 124.24 ;
      RECT  117.89 123.325 118.1 123.655 ;
      RECT  116.09 124.24 116.27 125.945 ;
      RECT  116.09 123.325 116.27 124.24 ;
      RECT  114.77 124.035 114.98 124.24 ;
      RECT  117.89 123.655 118.1 124.035 ;
      RECT  116.81 124.24 116.99 125.945 ;
      RECT  114.98 124.035 115.19 124.24 ;
      RECT  114.77 123.655 114.98 124.035 ;
      POLYGON  117.38 125.32 117.38 125.73 117.635 125.73 117.635 125.4 117.555 125.32 117.38 125.32 ;
      RECT  115.37 123.325 115.55 124.24 ;
      RECT  114.98 123.325 115.19 123.655 ;
      RECT  114.98 123.655 115.19 124.035 ;
      RECT  119.03 124.33 118.82 124.74 ;
      RECT  121.43 123.325 121.22 123.655 ;
      RECT  118.385 124.24 118.31 125.945 ;
      RECT  118.47 124.825 118.385 125.235 ;
      RECT  119.39 123.325 119.21 124.24 ;
      POLYGON  118.385 123.325 118.385 123.655 118.82 123.655 118.82 124.035 118.385 124.035 118.385 124.24 118.31 124.24 118.31 123.325 118.385 123.325 ;
      RECT  118.31 124.24 118.1 125.945 ;
      POLYGON  118.82 124.33 118.82 124.74 118.645 124.74 118.565 124.66 118.565 124.33 118.82 124.33 ;
      RECT  121.43 124.24 121.22 125.945 ;
      RECT  119.75 123.325 119.57 124.24 ;
      RECT  120.83 124.24 120.65 125.945 ;
      RECT  119.03 125.32 118.82 125.73 ;
      RECT  118.31 124.035 118.1 124.24 ;
      RECT  121.22 124.24 121.01 125.945 ;
      RECT  119.03 123.655 118.82 124.035 ;
      RECT  120.47 124.24 120.29 125.945 ;
      RECT  119.75 124.24 119.57 125.945 ;
      RECT  120.47 123.325 120.29 124.24 ;
      RECT  118.31 123.325 118.1 123.655 ;
      RECT  120.11 124.24 119.93 125.945 ;
      RECT  120.11 123.325 119.93 124.24 ;
      RECT  121.43 124.035 121.22 124.24 ;
      RECT  118.31 123.655 118.1 124.035 ;
      RECT  119.39 124.24 119.21 125.945 ;
      RECT  121.22 124.035 121.01 124.24 ;
      RECT  121.43 123.655 121.22 124.035 ;
      POLYGON  118.82 125.32 118.82 125.73 118.565 125.73 118.565 125.4 118.645 125.32 118.82 125.32 ;
      RECT  120.83 123.325 120.65 124.24 ;
      RECT  121.22 123.325 121.01 123.655 ;
      RECT  121.22 123.655 121.01 124.035 ;
      RECT  123.41 124.33 123.62 124.74 ;
      RECT  121.01 123.325 121.22 123.655 ;
      RECT  124.055 124.24 124.13 125.945 ;
      RECT  123.97 124.825 124.055 125.235 ;
      RECT  123.05 123.325 123.23 124.24 ;
      POLYGON  124.055 123.325 124.055 123.655 123.62 123.655 123.62 124.035 124.055 124.035 124.055 124.24 124.13 124.24 124.13 123.325 124.055 123.325 ;
      RECT  124.13 124.24 124.34 125.945 ;
      POLYGON  123.62 124.33 123.62 124.74 123.795 124.74 123.875 124.66 123.875 124.33 123.62 124.33 ;
      RECT  121.01 124.24 121.22 125.945 ;
      RECT  122.69 123.325 122.87 124.24 ;
      RECT  121.61 124.24 121.79 125.945 ;
      RECT  123.41 125.32 123.62 125.73 ;
      RECT  124.13 124.035 124.34 124.24 ;
      RECT  121.22 124.24 121.43 125.945 ;
      RECT  123.41 123.655 123.62 124.035 ;
      RECT  121.97 124.24 122.15 125.945 ;
      RECT  122.69 124.24 122.87 125.945 ;
      RECT  121.97 123.325 122.15 124.24 ;
      RECT  124.13 123.325 124.34 123.655 ;
      RECT  122.33 124.24 122.51 125.945 ;
      RECT  122.33 123.325 122.51 124.24 ;
      RECT  121.01 124.035 121.22 124.24 ;
      RECT  124.13 123.655 124.34 124.035 ;
      RECT  123.05 124.24 123.23 125.945 ;
      RECT  121.22 124.035 121.43 124.24 ;
      RECT  121.01 123.655 121.22 124.035 ;
      POLYGON  123.62 125.32 123.62 125.73 123.875 125.73 123.875 125.4 123.795 125.32 123.62 125.32 ;
      RECT  121.61 123.325 121.79 124.24 ;
      RECT  121.22 123.325 121.43 123.655 ;
      RECT  121.22 123.655 121.43 124.035 ;
      RECT  125.27 124.33 125.06 124.74 ;
      RECT  127.67 123.325 127.46 123.655 ;
      RECT  124.625 124.24 124.55 125.945 ;
      RECT  124.71 124.825 124.625 125.235 ;
      RECT  125.63 123.325 125.45 124.24 ;
      POLYGON  124.625 123.325 124.625 123.655 125.06 123.655 125.06 124.035 124.625 124.035 124.625 124.24 124.55 124.24 124.55 123.325 124.625 123.325 ;
      RECT  124.55 124.24 124.34 125.945 ;
      POLYGON  125.06 124.33 125.06 124.74 124.885 124.74 124.805 124.66 124.805 124.33 125.06 124.33 ;
      RECT  127.67 124.24 127.46 125.945 ;
      RECT  125.99 123.325 125.81 124.24 ;
      RECT  127.07 124.24 126.89 125.945 ;
      RECT  125.27 125.32 125.06 125.73 ;
      RECT  124.55 124.035 124.34 124.24 ;
      RECT  127.46 124.24 127.25 125.945 ;
      RECT  125.27 123.655 125.06 124.035 ;
      RECT  126.71 124.24 126.53 125.945 ;
      RECT  125.99 124.24 125.81 125.945 ;
      RECT  126.71 123.325 126.53 124.24 ;
      RECT  124.55 123.325 124.34 123.655 ;
      RECT  126.35 124.24 126.17 125.945 ;
      RECT  126.35 123.325 126.17 124.24 ;
      RECT  127.67 124.035 127.46 124.24 ;
      RECT  124.55 123.655 124.34 124.035 ;
      RECT  125.63 124.24 125.45 125.945 ;
      RECT  127.46 124.035 127.25 124.24 ;
      RECT  127.67 123.655 127.46 124.035 ;
      POLYGON  125.06 125.32 125.06 125.73 124.805 125.73 124.805 125.4 124.885 125.32 125.06 125.32 ;
      RECT  127.07 123.325 126.89 124.24 ;
      RECT  127.46 123.325 127.25 123.655 ;
      RECT  127.46 123.655 127.25 124.035 ;
      RECT  129.65 124.33 129.86 124.74 ;
      RECT  127.25 123.325 127.46 123.655 ;
      RECT  130.295 124.24 130.37 125.945 ;
      RECT  130.21 124.825 130.295 125.235 ;
      RECT  129.29 123.325 129.47 124.24 ;
      POLYGON  130.295 123.325 130.295 123.655 129.86 123.655 129.86 124.035 130.295 124.035 130.295 124.24 130.37 124.24 130.37 123.325 130.295 123.325 ;
      RECT  130.37 124.24 130.58 125.945 ;
      POLYGON  129.86 124.33 129.86 124.74 130.035 124.74 130.115 124.66 130.115 124.33 129.86 124.33 ;
      RECT  127.25 124.24 127.46 125.945 ;
      RECT  128.93 123.325 129.11 124.24 ;
      RECT  127.85 124.24 128.03 125.945 ;
      RECT  129.65 125.32 129.86 125.73 ;
      RECT  130.37 124.035 130.58 124.24 ;
      RECT  127.46 124.24 127.67 125.945 ;
      RECT  129.65 123.655 129.86 124.035 ;
      RECT  128.21 124.24 128.39 125.945 ;
      RECT  128.93 124.24 129.11 125.945 ;
      RECT  128.21 123.325 128.39 124.24 ;
      RECT  130.37 123.325 130.58 123.655 ;
      RECT  128.57 124.24 128.75 125.945 ;
      RECT  128.57 123.325 128.75 124.24 ;
      RECT  127.25 124.035 127.46 124.24 ;
      RECT  130.37 123.655 130.58 124.035 ;
      RECT  129.29 124.24 129.47 125.945 ;
      RECT  127.46 124.035 127.67 124.24 ;
      RECT  127.25 123.655 127.46 124.035 ;
      POLYGON  129.86 125.32 129.86 125.73 130.115 125.73 130.115 125.4 130.035 125.32 129.86 125.32 ;
      RECT  127.85 123.325 128.03 124.24 ;
      RECT  127.46 123.325 127.67 123.655 ;
      RECT  127.46 123.655 127.67 124.035 ;
      RECT  131.51 124.33 131.3 124.74 ;
      RECT  133.91 123.325 133.7 123.655 ;
      RECT  130.865 124.24 130.79 125.945 ;
      RECT  130.95 124.825 130.865 125.235 ;
      RECT  131.87 123.325 131.69 124.24 ;
      POLYGON  130.865 123.325 130.865 123.655 131.3 123.655 131.3 124.035 130.865 124.035 130.865 124.24 130.79 124.24 130.79 123.325 130.865 123.325 ;
      RECT  130.79 124.24 130.58 125.945 ;
      POLYGON  131.3 124.33 131.3 124.74 131.125 124.74 131.045 124.66 131.045 124.33 131.3 124.33 ;
      RECT  133.91 124.24 133.7 125.945 ;
      RECT  132.23 123.325 132.05 124.24 ;
      RECT  133.31 124.24 133.13 125.945 ;
      RECT  131.51 125.32 131.3 125.73 ;
      RECT  130.79 124.035 130.58 124.24 ;
      RECT  133.7 124.24 133.49 125.945 ;
      RECT  131.51 123.655 131.3 124.035 ;
      RECT  132.95 124.24 132.77 125.945 ;
      RECT  132.23 124.24 132.05 125.945 ;
      RECT  132.95 123.325 132.77 124.24 ;
      RECT  130.79 123.325 130.58 123.655 ;
      RECT  132.59 124.24 132.41 125.945 ;
      RECT  132.59 123.325 132.41 124.24 ;
      RECT  133.91 124.035 133.7 124.24 ;
      RECT  130.79 123.655 130.58 124.035 ;
      RECT  131.87 124.24 131.69 125.945 ;
      RECT  133.7 124.035 133.49 124.24 ;
      RECT  133.91 123.655 133.7 124.035 ;
      POLYGON  131.3 125.32 131.3 125.73 131.045 125.73 131.045 125.4 131.125 125.32 131.3 125.32 ;
      RECT  133.31 123.325 133.13 124.24 ;
      RECT  133.7 123.325 133.49 123.655 ;
      RECT  133.7 123.655 133.49 124.035 ;
      RECT  135.89 124.33 136.1 124.74 ;
      RECT  133.49 123.325 133.7 123.655 ;
      RECT  136.535 124.24 136.61 125.945 ;
      RECT  136.45 124.825 136.535 125.235 ;
      RECT  135.53 123.325 135.71 124.24 ;
      POLYGON  136.535 123.325 136.535 123.655 136.1 123.655 136.1 124.035 136.535 124.035 136.535 124.24 136.61 124.24 136.61 123.325 136.535 123.325 ;
      RECT  136.61 124.24 136.82 125.945 ;
      POLYGON  136.1 124.33 136.1 124.74 136.275 124.74 136.355 124.66 136.355 124.33 136.1 124.33 ;
      RECT  133.49 124.24 133.7 125.945 ;
      RECT  135.17 123.325 135.35 124.24 ;
      RECT  134.09 124.24 134.27 125.945 ;
      RECT  135.89 125.32 136.1 125.73 ;
      RECT  136.61 124.035 136.82 124.24 ;
      RECT  133.7 124.24 133.91 125.945 ;
      RECT  135.89 123.655 136.1 124.035 ;
      RECT  134.45 124.24 134.63 125.945 ;
      RECT  135.17 124.24 135.35 125.945 ;
      RECT  134.45 123.325 134.63 124.24 ;
      RECT  136.61 123.325 136.82 123.655 ;
      RECT  134.81 124.24 134.99 125.945 ;
      RECT  134.81 123.325 134.99 124.24 ;
      RECT  133.49 124.035 133.7 124.24 ;
      RECT  136.61 123.655 136.82 124.035 ;
      RECT  135.53 124.24 135.71 125.945 ;
      RECT  133.7 124.035 133.91 124.24 ;
      RECT  133.49 123.655 133.7 124.035 ;
      POLYGON  136.1 125.32 136.1 125.73 136.355 125.73 136.355 125.4 136.275 125.32 136.1 125.32 ;
      RECT  134.09 123.325 134.27 124.24 ;
      RECT  133.7 123.325 133.91 123.655 ;
      RECT  133.7 123.655 133.91 124.035 ;
      RECT  137.75 124.33 137.54 124.74 ;
      RECT  140.15 123.325 139.94 123.655 ;
      RECT  137.105 124.24 137.03 125.945 ;
      RECT  137.19 124.825 137.105 125.235 ;
      RECT  138.11 123.325 137.93 124.24 ;
      POLYGON  137.105 123.325 137.105 123.655 137.54 123.655 137.54 124.035 137.105 124.035 137.105 124.24 137.03 124.24 137.03 123.325 137.105 123.325 ;
      RECT  137.03 124.24 136.82 125.945 ;
      POLYGON  137.54 124.33 137.54 124.74 137.365 124.74 137.285 124.66 137.285 124.33 137.54 124.33 ;
      RECT  140.15 124.24 139.94 125.945 ;
      RECT  138.47 123.325 138.29 124.24 ;
      RECT  139.55 124.24 139.37 125.945 ;
      RECT  137.75 125.32 137.54 125.73 ;
      RECT  137.03 124.035 136.82 124.24 ;
      RECT  139.94 124.24 139.73 125.945 ;
      RECT  137.75 123.655 137.54 124.035 ;
      RECT  139.19 124.24 139.01 125.945 ;
      RECT  138.47 124.24 138.29 125.945 ;
      RECT  139.19 123.325 139.01 124.24 ;
      RECT  137.03 123.325 136.82 123.655 ;
      RECT  138.83 124.24 138.65 125.945 ;
      RECT  138.83 123.325 138.65 124.24 ;
      RECT  140.15 124.035 139.94 124.24 ;
      RECT  137.03 123.655 136.82 124.035 ;
      RECT  138.11 124.24 137.93 125.945 ;
      RECT  139.94 124.035 139.73 124.24 ;
      RECT  140.15 123.655 139.94 124.035 ;
      POLYGON  137.54 125.32 137.54 125.73 137.285 125.73 137.285 125.4 137.365 125.32 137.54 125.32 ;
      RECT  139.55 123.325 139.37 124.24 ;
      RECT  139.94 123.325 139.73 123.655 ;
      RECT  139.94 123.655 139.73 124.035 ;
      RECT  142.13 124.33 142.34 124.74 ;
      RECT  139.73 123.325 139.94 123.655 ;
      RECT  142.775 124.24 142.85 125.945 ;
      RECT  142.69 124.825 142.775 125.235 ;
      RECT  141.77 123.325 141.95 124.24 ;
      POLYGON  142.775 123.325 142.775 123.655 142.34 123.655 142.34 124.035 142.775 124.035 142.775 124.24 142.85 124.24 142.85 123.325 142.775 123.325 ;
      RECT  142.85 124.24 143.06 125.945 ;
      POLYGON  142.34 124.33 142.34 124.74 142.515 124.74 142.595 124.66 142.595 124.33 142.34 124.33 ;
      RECT  139.73 124.24 139.94 125.945 ;
      RECT  141.41 123.325 141.59 124.24 ;
      RECT  140.33 124.24 140.51 125.945 ;
      RECT  142.13 125.32 142.34 125.73 ;
      RECT  142.85 124.035 143.06 124.24 ;
      RECT  139.94 124.24 140.15 125.945 ;
      RECT  142.13 123.655 142.34 124.035 ;
      RECT  140.69 124.24 140.87 125.945 ;
      RECT  141.41 124.24 141.59 125.945 ;
      RECT  140.69 123.325 140.87 124.24 ;
      RECT  142.85 123.325 143.06 123.655 ;
      RECT  141.05 124.24 141.23 125.945 ;
      RECT  141.05 123.325 141.23 124.24 ;
      RECT  139.73 124.035 139.94 124.24 ;
      RECT  142.85 123.655 143.06 124.035 ;
      RECT  141.77 124.24 141.95 125.945 ;
      RECT  139.94 124.035 140.15 124.24 ;
      RECT  139.73 123.655 139.94 124.035 ;
      POLYGON  142.34 125.32 142.34 125.73 142.595 125.73 142.595 125.4 142.515 125.32 142.34 125.32 ;
      RECT  140.33 123.325 140.51 124.24 ;
      RECT  139.94 123.325 140.15 123.655 ;
      RECT  139.94 123.655 140.15 124.035 ;
      RECT  143.99 124.33 143.78 124.74 ;
      RECT  146.39 123.325 146.18 123.655 ;
      RECT  143.345 124.24 143.27 125.945 ;
      RECT  143.43 124.825 143.345 125.235 ;
      RECT  144.35 123.325 144.17 124.24 ;
      POLYGON  143.345 123.325 143.345 123.655 143.78 123.655 143.78 124.035 143.345 124.035 143.345 124.24 143.27 124.24 143.27 123.325 143.345 123.325 ;
      RECT  143.27 124.24 143.06 125.945 ;
      POLYGON  143.78 124.33 143.78 124.74 143.605 124.74 143.525 124.66 143.525 124.33 143.78 124.33 ;
      RECT  146.39 124.24 146.18 125.945 ;
      RECT  144.71 123.325 144.53 124.24 ;
      RECT  145.79 124.24 145.61 125.945 ;
      RECT  143.99 125.32 143.78 125.73 ;
      RECT  143.27 124.035 143.06 124.24 ;
      RECT  146.18 124.24 145.97 125.945 ;
      RECT  143.99 123.655 143.78 124.035 ;
      RECT  145.43 124.24 145.25 125.945 ;
      RECT  144.71 124.24 144.53 125.945 ;
      RECT  145.43 123.325 145.25 124.24 ;
      RECT  143.27 123.325 143.06 123.655 ;
      RECT  145.07 124.24 144.89 125.945 ;
      RECT  145.07 123.325 144.89 124.24 ;
      RECT  146.39 124.035 146.18 124.24 ;
      RECT  143.27 123.655 143.06 124.035 ;
      RECT  144.35 124.24 144.17 125.945 ;
      RECT  146.18 124.035 145.97 124.24 ;
      RECT  146.39 123.655 146.18 124.035 ;
      POLYGON  143.78 125.32 143.78 125.73 143.525 125.73 143.525 125.4 143.605 125.32 143.78 125.32 ;
      RECT  145.79 123.325 145.61 124.24 ;
      RECT  146.18 123.325 145.97 123.655 ;
      RECT  146.18 123.655 145.97 124.035 ;
      RECT  96.65 123.845 96.83 125.82 ;
      RECT  97.01 123.845 97.19 125.82 ;
      RECT  97.73 123.845 97.91 125.82 ;
      RECT  98.09 123.845 98.27 125.82 ;
      RECT  101.93 123.845 102.11 125.82 ;
      RECT  101.57 123.845 101.75 125.82 ;
      RECT  100.85 123.845 101.03 125.82 ;
      RECT  100.49 123.845 100.67 125.82 ;
      RECT  102.89 123.845 103.07 125.82 ;
      RECT  103.25 123.845 103.43 125.82 ;
      RECT  103.97 123.845 104.15 125.82 ;
      RECT  104.33 123.845 104.51 125.82 ;
      RECT  108.17 123.845 108.35 125.82 ;
      RECT  107.81 123.845 107.99 125.82 ;
      RECT  107.09 123.845 107.27 125.82 ;
      RECT  106.73 123.845 106.91 125.82 ;
      RECT  109.13 123.845 109.31 125.82 ;
      RECT  109.49 123.845 109.67 125.82 ;
      RECT  110.21 123.845 110.39 125.82 ;
      RECT  110.57 123.845 110.75 125.82 ;
      RECT  114.41 123.845 114.59 125.82 ;
      RECT  114.05 123.845 114.23 125.82 ;
      RECT  113.33 123.845 113.51 125.82 ;
      RECT  112.97 123.845 113.15 125.82 ;
      RECT  115.37 123.845 115.55 125.82 ;
      RECT  115.73 123.845 115.91 125.82 ;
      RECT  116.45 123.845 116.63 125.82 ;
      RECT  116.81 123.845 116.99 125.82 ;
      RECT  120.65 123.845 120.83 125.82 ;
      RECT  120.29 123.845 120.47 125.82 ;
      RECT  119.57 123.845 119.75 125.82 ;
      RECT  119.21 123.845 119.39 125.82 ;
      RECT  121.61 123.845 121.79 125.82 ;
      RECT  121.97 123.845 122.15 125.82 ;
      RECT  122.69 123.845 122.87 125.82 ;
      RECT  123.05 123.845 123.23 125.82 ;
      RECT  126.89 123.845 127.07 125.82 ;
      RECT  126.53 123.845 126.71 125.82 ;
      RECT  125.81 123.845 125.99 125.82 ;
      RECT  125.45 123.845 125.63 125.82 ;
      RECT  127.85 123.845 128.03 125.82 ;
      RECT  128.21 123.845 128.39 125.82 ;
      RECT  128.93 123.845 129.11 125.82 ;
      RECT  129.29 123.845 129.47 125.82 ;
      RECT  133.13 123.845 133.31 125.82 ;
      RECT  132.77 123.845 132.95 125.82 ;
      RECT  132.05 123.845 132.23 125.82 ;
      RECT  131.69 123.845 131.87 125.82 ;
      RECT  134.09 123.845 134.27 125.82 ;
      RECT  134.45 123.845 134.63 125.82 ;
      RECT  135.17 123.845 135.35 125.82 ;
      RECT  135.53 123.845 135.71 125.82 ;
      RECT  139.37 123.845 139.55 125.82 ;
      RECT  139.01 123.845 139.19 125.82 ;
      RECT  138.29 123.845 138.47 125.82 ;
      RECT  137.93 123.845 138.11 125.82 ;
      RECT  140.33 123.845 140.51 125.82 ;
      RECT  140.69 123.845 140.87 125.82 ;
      RECT  141.41 123.845 141.59 125.82 ;
      RECT  141.77 123.845 141.95 125.82 ;
      RECT  145.61 123.845 145.79 125.82 ;
      RECT  145.25 123.845 145.43 125.82 ;
      RECT  144.53 123.845 144.71 125.82 ;
      RECT  144.17 123.845 144.35 125.82 ;
      RECT  109.85 124.24 110.03 125.945 ;
      RECT  144.89 124.24 145.07 125.945 ;
      RECT  113.69 124.24 113.87 125.945 ;
      RECT  138.65 124.24 138.83 125.945 ;
      RECT  126.17 124.24 126.35 125.945 ;
      RECT  107.45 124.24 107.63 125.945 ;
      RECT  101.21 124.24 101.39 125.945 ;
      RECT  116.09 124.24 116.27 125.945 ;
      RECT  119.93 124.24 120.11 125.945 ;
      RECT  134.81 124.24 134.99 125.945 ;
      RECT  103.61 124.24 103.79 125.945 ;
      RECT  122.33 124.24 122.51 125.945 ;
      RECT  97.37 124.24 97.55 125.945 ;
      RECT  132.41 124.24 132.59 125.945 ;
      RECT  128.57 124.24 128.75 125.945 ;
      RECT  141.05 124.24 141.23 125.945 ;
      RECT  97.73 89.085 97.91 90.665 ;
      RECT  97.37 88.295 97.55 89.085 ;
      RECT  97.33 89.085 97.46 89.795 ;
      RECT  97.01 88.295 97.19 89.085 ;
      RECT  98.09 89.085 98.27 90.665 ;
      RECT  97.73 88.295 97.91 89.085 ;
      RECT  98.09 88.295 98.27 89.085 ;
      RECT  96.65 89.085 96.83 90.665 ;
      RECT  96.65 88.295 96.83 89.085 ;
      RECT  97.01 89.085 97.19 90.665 ;
      RECT  97.46 89.085 97.59 89.795 ;
      RECT  97.37 89.085 97.55 90.665 ;
      RECT  101.03 89.085 100.85 90.665 ;
      RECT  101.39 88.295 101.21 89.085 ;
      RECT  101.43 89.085 101.3 89.795 ;
      RECT  101.75 88.295 101.57 89.085 ;
      RECT  100.67 89.085 100.49 90.665 ;
      RECT  101.03 88.295 100.85 89.085 ;
      RECT  100.67 88.295 100.49 89.085 ;
      RECT  102.11 89.085 101.93 90.665 ;
      RECT  102.11 88.295 101.93 89.085 ;
      RECT  101.75 89.085 101.57 90.665 ;
      RECT  101.3 89.085 101.17 89.795 ;
      RECT  101.39 89.085 101.21 90.665 ;
      RECT  103.97 89.085 104.15 90.665 ;
      RECT  103.61 88.295 103.79 89.085 ;
      RECT  103.57 89.085 103.7 89.795 ;
      RECT  103.25 88.295 103.43 89.085 ;
      RECT  104.33 89.085 104.51 90.665 ;
      RECT  103.97 88.295 104.15 89.085 ;
      RECT  104.33 88.295 104.51 89.085 ;
      RECT  102.89 89.085 103.07 90.665 ;
      RECT  102.89 88.295 103.07 89.085 ;
      RECT  103.25 89.085 103.43 90.665 ;
      RECT  103.7 89.085 103.83 89.795 ;
      RECT  103.61 89.085 103.79 90.665 ;
      RECT  107.27 89.085 107.09 90.665 ;
      RECT  107.63 88.295 107.45 89.085 ;
      RECT  107.67 89.085 107.54 89.795 ;
      RECT  107.99 88.295 107.81 89.085 ;
      RECT  106.91 89.085 106.73 90.665 ;
      RECT  107.27 88.295 107.09 89.085 ;
      RECT  106.91 88.295 106.73 89.085 ;
      RECT  108.35 89.085 108.17 90.665 ;
      RECT  108.35 88.295 108.17 89.085 ;
      RECT  107.99 89.085 107.81 90.665 ;
      RECT  107.54 89.085 107.41 89.795 ;
      RECT  107.63 89.085 107.45 90.665 ;
      RECT  110.21 89.085 110.39 90.665 ;
      RECT  109.85 88.295 110.03 89.085 ;
      RECT  109.81 89.085 109.94 89.795 ;
      RECT  109.49 88.295 109.67 89.085 ;
      RECT  110.57 89.085 110.75 90.665 ;
      RECT  110.21 88.295 110.39 89.085 ;
      RECT  110.57 88.295 110.75 89.085 ;
      RECT  109.13 89.085 109.31 90.665 ;
      RECT  109.13 88.295 109.31 89.085 ;
      RECT  109.49 89.085 109.67 90.665 ;
      RECT  109.94 89.085 110.07 89.795 ;
      RECT  109.85 89.085 110.03 90.665 ;
      RECT  113.51 89.085 113.33 90.665 ;
      RECT  113.87 88.295 113.69 89.085 ;
      RECT  113.91 89.085 113.78 89.795 ;
      RECT  114.23 88.295 114.05 89.085 ;
      RECT  113.15 89.085 112.97 90.665 ;
      RECT  113.51 88.295 113.33 89.085 ;
      RECT  113.15 88.295 112.97 89.085 ;
      RECT  114.59 89.085 114.41 90.665 ;
      RECT  114.59 88.295 114.41 89.085 ;
      RECT  114.23 89.085 114.05 90.665 ;
      RECT  113.78 89.085 113.65 89.795 ;
      RECT  113.87 89.085 113.69 90.665 ;
      RECT  116.45 89.085 116.63 90.665 ;
      RECT  116.09 88.295 116.27 89.085 ;
      RECT  116.05 89.085 116.18 89.795 ;
      RECT  115.73 88.295 115.91 89.085 ;
      RECT  116.81 89.085 116.99 90.665 ;
      RECT  116.45 88.295 116.63 89.085 ;
      RECT  116.81 88.295 116.99 89.085 ;
      RECT  115.37 89.085 115.55 90.665 ;
      RECT  115.37 88.295 115.55 89.085 ;
      RECT  115.73 89.085 115.91 90.665 ;
      RECT  116.18 89.085 116.31 89.795 ;
      RECT  116.09 89.085 116.27 90.665 ;
      RECT  119.75 89.085 119.57 90.665 ;
      RECT  120.11 88.295 119.93 89.085 ;
      RECT  120.15 89.085 120.02 89.795 ;
      RECT  120.47 88.295 120.29 89.085 ;
      RECT  119.39 89.085 119.21 90.665 ;
      RECT  119.75 88.295 119.57 89.085 ;
      RECT  119.39 88.295 119.21 89.085 ;
      RECT  120.83 89.085 120.65 90.665 ;
      RECT  120.83 88.295 120.65 89.085 ;
      RECT  120.47 89.085 120.29 90.665 ;
      RECT  120.02 89.085 119.89 89.795 ;
      RECT  120.11 89.085 119.93 90.665 ;
      RECT  122.69 89.085 122.87 90.665 ;
      RECT  122.33 88.295 122.51 89.085 ;
      RECT  122.29 89.085 122.42 89.795 ;
      RECT  121.97 88.295 122.15 89.085 ;
      RECT  123.05 89.085 123.23 90.665 ;
      RECT  122.69 88.295 122.87 89.085 ;
      RECT  123.05 88.295 123.23 89.085 ;
      RECT  121.61 89.085 121.79 90.665 ;
      RECT  121.61 88.295 121.79 89.085 ;
      RECT  121.97 89.085 122.15 90.665 ;
      RECT  122.42 89.085 122.55 89.795 ;
      RECT  122.33 89.085 122.51 90.665 ;
      RECT  125.99 89.085 125.81 90.665 ;
      RECT  126.35 88.295 126.17 89.085 ;
      RECT  126.39 89.085 126.26 89.795 ;
      RECT  126.71 88.295 126.53 89.085 ;
      RECT  125.63 89.085 125.45 90.665 ;
      RECT  125.99 88.295 125.81 89.085 ;
      RECT  125.63 88.295 125.45 89.085 ;
      RECT  127.07 89.085 126.89 90.665 ;
      RECT  127.07 88.295 126.89 89.085 ;
      RECT  126.71 89.085 126.53 90.665 ;
      RECT  126.26 89.085 126.13 89.795 ;
      RECT  126.35 89.085 126.17 90.665 ;
      RECT  128.93 89.085 129.11 90.665 ;
      RECT  128.57 88.295 128.75 89.085 ;
      RECT  128.53 89.085 128.66 89.795 ;
      RECT  128.21 88.295 128.39 89.085 ;
      RECT  129.29 89.085 129.47 90.665 ;
      RECT  128.93 88.295 129.11 89.085 ;
      RECT  129.29 88.295 129.47 89.085 ;
      RECT  127.85 89.085 128.03 90.665 ;
      RECT  127.85 88.295 128.03 89.085 ;
      RECT  128.21 89.085 128.39 90.665 ;
      RECT  128.66 89.085 128.79 89.795 ;
      RECT  128.57 89.085 128.75 90.665 ;
      RECT  132.23 89.085 132.05 90.665 ;
      RECT  132.59 88.295 132.41 89.085 ;
      RECT  132.63 89.085 132.5 89.795 ;
      RECT  132.95 88.295 132.77 89.085 ;
      RECT  131.87 89.085 131.69 90.665 ;
      RECT  132.23 88.295 132.05 89.085 ;
      RECT  131.87 88.295 131.69 89.085 ;
      RECT  133.31 89.085 133.13 90.665 ;
      RECT  133.31 88.295 133.13 89.085 ;
      RECT  132.95 89.085 132.77 90.665 ;
      RECT  132.5 89.085 132.37 89.795 ;
      RECT  132.59 89.085 132.41 90.665 ;
      RECT  135.17 89.085 135.35 90.665 ;
      RECT  134.81 88.295 134.99 89.085 ;
      RECT  134.77 89.085 134.9 89.795 ;
      RECT  134.45 88.295 134.63 89.085 ;
      RECT  135.53 89.085 135.71 90.665 ;
      RECT  135.17 88.295 135.35 89.085 ;
      RECT  135.53 88.295 135.71 89.085 ;
      RECT  134.09 89.085 134.27 90.665 ;
      RECT  134.09 88.295 134.27 89.085 ;
      RECT  134.45 89.085 134.63 90.665 ;
      RECT  134.9 89.085 135.03 89.795 ;
      RECT  134.81 89.085 134.99 90.665 ;
      RECT  138.47 89.085 138.29 90.665 ;
      RECT  138.83 88.295 138.65 89.085 ;
      RECT  138.87 89.085 138.74 89.795 ;
      RECT  139.19 88.295 139.01 89.085 ;
      RECT  138.11 89.085 137.93 90.665 ;
      RECT  138.47 88.295 138.29 89.085 ;
      RECT  138.11 88.295 137.93 89.085 ;
      RECT  139.55 89.085 139.37 90.665 ;
      RECT  139.55 88.295 139.37 89.085 ;
      RECT  139.19 89.085 139.01 90.665 ;
      RECT  138.74 89.085 138.61 89.795 ;
      RECT  138.83 89.085 138.65 90.665 ;
      RECT  141.41 89.085 141.59 90.665 ;
      RECT  141.05 88.295 141.23 89.085 ;
      RECT  141.01 89.085 141.14 89.795 ;
      RECT  140.69 88.295 140.87 89.085 ;
      RECT  141.77 89.085 141.95 90.665 ;
      RECT  141.41 88.295 141.59 89.085 ;
      RECT  141.77 88.295 141.95 89.085 ;
      RECT  140.33 89.085 140.51 90.665 ;
      RECT  140.33 88.295 140.51 89.085 ;
      RECT  140.69 89.085 140.87 90.665 ;
      RECT  141.14 89.085 141.27 89.795 ;
      RECT  141.05 89.085 141.23 90.665 ;
      RECT  144.71 89.085 144.53 90.665 ;
      RECT  145.07 88.295 144.89 89.085 ;
      RECT  145.11 89.085 144.98 89.795 ;
      RECT  145.43 88.295 145.25 89.085 ;
      RECT  144.35 89.085 144.17 90.665 ;
      RECT  144.71 88.295 144.53 89.085 ;
      RECT  144.35 88.295 144.17 89.085 ;
      RECT  145.79 89.085 145.61 90.665 ;
      RECT  145.79 88.295 145.61 89.085 ;
      RECT  145.43 89.085 145.25 90.665 ;
      RECT  144.98 89.085 144.85 89.795 ;
      RECT  145.07 89.085 144.89 90.665 ;
      RECT  96.65 88.295 96.83 90.27 ;
      RECT  97.01 88.295 97.19 90.27 ;
      RECT  97.73 88.295 97.91 90.27 ;
      RECT  98.09 88.295 98.27 90.27 ;
      RECT  101.93 88.295 102.11 90.27 ;
      RECT  101.57 88.295 101.75 90.27 ;
      RECT  100.85 88.295 101.03 90.27 ;
      RECT  100.49 88.295 100.67 90.27 ;
      RECT  102.89 88.295 103.07 90.27 ;
      RECT  103.25 88.295 103.43 90.27 ;
      RECT  103.97 88.295 104.15 90.27 ;
      RECT  104.33 88.295 104.51 90.27 ;
      RECT  108.17 88.295 108.35 90.27 ;
      RECT  107.81 88.295 107.99 90.27 ;
      RECT  107.09 88.295 107.27 90.27 ;
      RECT  106.73 88.295 106.91 90.27 ;
      RECT  109.13 88.295 109.31 90.27 ;
      RECT  109.49 88.295 109.67 90.27 ;
      RECT  110.21 88.295 110.39 90.27 ;
      RECT  110.57 88.295 110.75 90.27 ;
      RECT  114.41 88.295 114.59 90.27 ;
      RECT  114.05 88.295 114.23 90.27 ;
      RECT  113.33 88.295 113.51 90.27 ;
      RECT  112.97 88.295 113.15 90.27 ;
      RECT  115.37 88.295 115.55 90.27 ;
      RECT  115.73 88.295 115.91 90.27 ;
      RECT  116.45 88.295 116.63 90.27 ;
      RECT  116.81 88.295 116.99 90.27 ;
      RECT  120.65 88.295 120.83 90.27 ;
      RECT  120.29 88.295 120.47 90.27 ;
      RECT  119.57 88.295 119.75 90.27 ;
      RECT  119.21 88.295 119.39 90.27 ;
      RECT  121.61 88.295 121.79 90.27 ;
      RECT  121.97 88.295 122.15 90.27 ;
      RECT  122.69 88.295 122.87 90.27 ;
      RECT  123.05 88.295 123.23 90.27 ;
      RECT  126.89 88.295 127.07 90.27 ;
      RECT  126.53 88.295 126.71 90.27 ;
      RECT  125.81 88.295 125.99 90.27 ;
      RECT  125.45 88.295 125.63 90.27 ;
      RECT  127.85 88.295 128.03 90.27 ;
      RECT  128.21 88.295 128.39 90.27 ;
      RECT  128.93 88.295 129.11 90.27 ;
      RECT  129.29 88.295 129.47 90.27 ;
      RECT  133.13 88.295 133.31 90.27 ;
      RECT  132.77 88.295 132.95 90.27 ;
      RECT  132.05 88.295 132.23 90.27 ;
      RECT  131.69 88.295 131.87 90.27 ;
      RECT  134.09 88.295 134.27 90.27 ;
      RECT  134.45 88.295 134.63 90.27 ;
      RECT  135.17 88.295 135.35 90.27 ;
      RECT  135.53 88.295 135.71 90.27 ;
      RECT  139.37 88.295 139.55 90.27 ;
      RECT  139.01 88.295 139.19 90.27 ;
      RECT  138.29 88.295 138.47 90.27 ;
      RECT  137.93 88.295 138.11 90.27 ;
      RECT  140.33 88.295 140.51 90.27 ;
      RECT  140.69 88.295 140.87 90.27 ;
      RECT  141.41 88.295 141.59 90.27 ;
      RECT  141.77 88.295 141.95 90.27 ;
      RECT  145.61 88.295 145.79 90.27 ;
      RECT  145.25 88.295 145.43 90.27 ;
      RECT  144.53 88.295 144.71 90.27 ;
      RECT  144.17 88.295 144.35 90.27 ;
      RECT  97.73 127.005 97.91 125.425 ;
      RECT  97.37 127.795 97.55 127.005 ;
      RECT  97.33 127.005 97.46 126.295 ;
      RECT  97.01 127.795 97.19 127.005 ;
      RECT  98.09 127.005 98.27 125.425 ;
      RECT  97.73 127.795 97.91 127.005 ;
      RECT  98.09 127.795 98.27 127.005 ;
      RECT  96.65 127.005 96.83 125.425 ;
      RECT  96.65 127.795 96.83 127.005 ;
      RECT  97.01 127.005 97.19 125.425 ;
      RECT  97.46 127.005 97.59 126.295 ;
      RECT  97.37 127.005 97.55 125.425 ;
      RECT  101.03 127.005 100.85 125.425 ;
      RECT  101.39 127.795 101.21 127.005 ;
      RECT  101.43 127.005 101.3 126.295 ;
      RECT  101.75 127.795 101.57 127.005 ;
      RECT  100.67 127.005 100.49 125.425 ;
      RECT  101.03 127.795 100.85 127.005 ;
      RECT  100.67 127.795 100.49 127.005 ;
      RECT  102.11 127.005 101.93 125.425 ;
      RECT  102.11 127.795 101.93 127.005 ;
      RECT  101.75 127.005 101.57 125.425 ;
      RECT  101.3 127.005 101.17 126.295 ;
      RECT  101.39 127.005 101.21 125.425 ;
      RECT  103.97 127.005 104.15 125.425 ;
      RECT  103.61 127.795 103.79 127.005 ;
      RECT  103.57 127.005 103.7 126.295 ;
      RECT  103.25 127.795 103.43 127.005 ;
      RECT  104.33 127.005 104.51 125.425 ;
      RECT  103.97 127.795 104.15 127.005 ;
      RECT  104.33 127.795 104.51 127.005 ;
      RECT  102.89 127.005 103.07 125.425 ;
      RECT  102.89 127.795 103.07 127.005 ;
      RECT  103.25 127.005 103.43 125.425 ;
      RECT  103.7 127.005 103.83 126.295 ;
      RECT  103.61 127.005 103.79 125.425 ;
      RECT  107.27 127.005 107.09 125.425 ;
      RECT  107.63 127.795 107.45 127.005 ;
      RECT  107.67 127.005 107.54 126.295 ;
      RECT  107.99 127.795 107.81 127.005 ;
      RECT  106.91 127.005 106.73 125.425 ;
      RECT  107.27 127.795 107.09 127.005 ;
      RECT  106.91 127.795 106.73 127.005 ;
      RECT  108.35 127.005 108.17 125.425 ;
      RECT  108.35 127.795 108.17 127.005 ;
      RECT  107.99 127.005 107.81 125.425 ;
      RECT  107.54 127.005 107.41 126.295 ;
      RECT  107.63 127.005 107.45 125.425 ;
      RECT  110.21 127.005 110.39 125.425 ;
      RECT  109.85 127.795 110.03 127.005 ;
      RECT  109.81 127.005 109.94 126.295 ;
      RECT  109.49 127.795 109.67 127.005 ;
      RECT  110.57 127.005 110.75 125.425 ;
      RECT  110.21 127.795 110.39 127.005 ;
      RECT  110.57 127.795 110.75 127.005 ;
      RECT  109.13 127.005 109.31 125.425 ;
      RECT  109.13 127.795 109.31 127.005 ;
      RECT  109.49 127.005 109.67 125.425 ;
      RECT  109.94 127.005 110.07 126.295 ;
      RECT  109.85 127.005 110.03 125.425 ;
      RECT  113.51 127.005 113.33 125.425 ;
      RECT  113.87 127.795 113.69 127.005 ;
      RECT  113.91 127.005 113.78 126.295 ;
      RECT  114.23 127.795 114.05 127.005 ;
      RECT  113.15 127.005 112.97 125.425 ;
      RECT  113.51 127.795 113.33 127.005 ;
      RECT  113.15 127.795 112.97 127.005 ;
      RECT  114.59 127.005 114.41 125.425 ;
      RECT  114.59 127.795 114.41 127.005 ;
      RECT  114.23 127.005 114.05 125.425 ;
      RECT  113.78 127.005 113.65 126.295 ;
      RECT  113.87 127.005 113.69 125.425 ;
      RECT  116.45 127.005 116.63 125.425 ;
      RECT  116.09 127.795 116.27 127.005 ;
      RECT  116.05 127.005 116.18 126.295 ;
      RECT  115.73 127.795 115.91 127.005 ;
      RECT  116.81 127.005 116.99 125.425 ;
      RECT  116.45 127.795 116.63 127.005 ;
      RECT  116.81 127.795 116.99 127.005 ;
      RECT  115.37 127.005 115.55 125.425 ;
      RECT  115.37 127.795 115.55 127.005 ;
      RECT  115.73 127.005 115.91 125.425 ;
      RECT  116.18 127.005 116.31 126.295 ;
      RECT  116.09 127.005 116.27 125.425 ;
      RECT  119.75 127.005 119.57 125.425 ;
      RECT  120.11 127.795 119.93 127.005 ;
      RECT  120.15 127.005 120.02 126.295 ;
      RECT  120.47 127.795 120.29 127.005 ;
      RECT  119.39 127.005 119.21 125.425 ;
      RECT  119.75 127.795 119.57 127.005 ;
      RECT  119.39 127.795 119.21 127.005 ;
      RECT  120.83 127.005 120.65 125.425 ;
      RECT  120.83 127.795 120.65 127.005 ;
      RECT  120.47 127.005 120.29 125.425 ;
      RECT  120.02 127.005 119.89 126.295 ;
      RECT  120.11 127.005 119.93 125.425 ;
      RECT  122.69 127.005 122.87 125.425 ;
      RECT  122.33 127.795 122.51 127.005 ;
      RECT  122.29 127.005 122.42 126.295 ;
      RECT  121.97 127.795 122.15 127.005 ;
      RECT  123.05 127.005 123.23 125.425 ;
      RECT  122.69 127.795 122.87 127.005 ;
      RECT  123.05 127.795 123.23 127.005 ;
      RECT  121.61 127.005 121.79 125.425 ;
      RECT  121.61 127.795 121.79 127.005 ;
      RECT  121.97 127.005 122.15 125.425 ;
      RECT  122.42 127.005 122.55 126.295 ;
      RECT  122.33 127.005 122.51 125.425 ;
      RECT  125.99 127.005 125.81 125.425 ;
      RECT  126.35 127.795 126.17 127.005 ;
      RECT  126.39 127.005 126.26 126.295 ;
      RECT  126.71 127.795 126.53 127.005 ;
      RECT  125.63 127.005 125.45 125.425 ;
      RECT  125.99 127.795 125.81 127.005 ;
      RECT  125.63 127.795 125.45 127.005 ;
      RECT  127.07 127.005 126.89 125.425 ;
      RECT  127.07 127.795 126.89 127.005 ;
      RECT  126.71 127.005 126.53 125.425 ;
      RECT  126.26 127.005 126.13 126.295 ;
      RECT  126.35 127.005 126.17 125.425 ;
      RECT  128.93 127.005 129.11 125.425 ;
      RECT  128.57 127.795 128.75 127.005 ;
      RECT  128.53 127.005 128.66 126.295 ;
      RECT  128.21 127.795 128.39 127.005 ;
      RECT  129.29 127.005 129.47 125.425 ;
      RECT  128.93 127.795 129.11 127.005 ;
      RECT  129.29 127.795 129.47 127.005 ;
      RECT  127.85 127.005 128.03 125.425 ;
      RECT  127.85 127.795 128.03 127.005 ;
      RECT  128.21 127.005 128.39 125.425 ;
      RECT  128.66 127.005 128.79 126.295 ;
      RECT  128.57 127.005 128.75 125.425 ;
      RECT  132.23 127.005 132.05 125.425 ;
      RECT  132.59 127.795 132.41 127.005 ;
      RECT  132.63 127.005 132.5 126.295 ;
      RECT  132.95 127.795 132.77 127.005 ;
      RECT  131.87 127.005 131.69 125.425 ;
      RECT  132.23 127.795 132.05 127.005 ;
      RECT  131.87 127.795 131.69 127.005 ;
      RECT  133.31 127.005 133.13 125.425 ;
      RECT  133.31 127.795 133.13 127.005 ;
      RECT  132.95 127.005 132.77 125.425 ;
      RECT  132.5 127.005 132.37 126.295 ;
      RECT  132.59 127.005 132.41 125.425 ;
      RECT  135.17 127.005 135.35 125.425 ;
      RECT  134.81 127.795 134.99 127.005 ;
      RECT  134.77 127.005 134.9 126.295 ;
      RECT  134.45 127.795 134.63 127.005 ;
      RECT  135.53 127.005 135.71 125.425 ;
      RECT  135.17 127.795 135.35 127.005 ;
      RECT  135.53 127.795 135.71 127.005 ;
      RECT  134.09 127.005 134.27 125.425 ;
      RECT  134.09 127.795 134.27 127.005 ;
      RECT  134.45 127.005 134.63 125.425 ;
      RECT  134.9 127.005 135.03 126.295 ;
      RECT  134.81 127.005 134.99 125.425 ;
      RECT  138.47 127.005 138.29 125.425 ;
      RECT  138.83 127.795 138.65 127.005 ;
      RECT  138.87 127.005 138.74 126.295 ;
      RECT  139.19 127.795 139.01 127.005 ;
      RECT  138.11 127.005 137.93 125.425 ;
      RECT  138.47 127.795 138.29 127.005 ;
      RECT  138.11 127.795 137.93 127.005 ;
      RECT  139.55 127.005 139.37 125.425 ;
      RECT  139.55 127.795 139.37 127.005 ;
      RECT  139.19 127.005 139.01 125.425 ;
      RECT  138.74 127.005 138.61 126.295 ;
      RECT  138.83 127.005 138.65 125.425 ;
      RECT  141.41 127.005 141.59 125.425 ;
      RECT  141.05 127.795 141.23 127.005 ;
      RECT  141.01 127.005 141.14 126.295 ;
      RECT  140.69 127.795 140.87 127.005 ;
      RECT  141.77 127.005 141.95 125.425 ;
      RECT  141.41 127.795 141.59 127.005 ;
      RECT  141.77 127.795 141.95 127.005 ;
      RECT  140.33 127.005 140.51 125.425 ;
      RECT  140.33 127.795 140.51 127.005 ;
      RECT  140.69 127.005 140.87 125.425 ;
      RECT  141.14 127.005 141.27 126.295 ;
      RECT  141.05 127.005 141.23 125.425 ;
      RECT  144.71 127.005 144.53 125.425 ;
      RECT  145.07 127.795 144.89 127.005 ;
      RECT  145.11 127.005 144.98 126.295 ;
      RECT  145.43 127.795 145.25 127.005 ;
      RECT  144.35 127.005 144.17 125.425 ;
      RECT  144.71 127.795 144.53 127.005 ;
      RECT  144.35 127.795 144.17 127.005 ;
      RECT  145.79 127.005 145.61 125.425 ;
      RECT  145.79 127.795 145.61 127.005 ;
      RECT  145.43 127.005 145.25 125.425 ;
      RECT  144.98 127.005 144.85 126.295 ;
      RECT  145.07 127.005 144.89 125.425 ;
      RECT  96.65 127.795 96.83 125.82 ;
      RECT  97.01 127.795 97.19 125.82 ;
      RECT  97.73 127.795 97.91 125.82 ;
      RECT  98.09 127.795 98.27 125.82 ;
      RECT  101.93 127.795 102.11 125.82 ;
      RECT  101.57 127.795 101.75 125.82 ;
      RECT  100.85 127.795 101.03 125.82 ;
      RECT  100.49 127.795 100.67 125.82 ;
      RECT  102.89 127.795 103.07 125.82 ;
      RECT  103.25 127.795 103.43 125.82 ;
      RECT  103.97 127.795 104.15 125.82 ;
      RECT  104.33 127.795 104.51 125.82 ;
      RECT  108.17 127.795 108.35 125.82 ;
      RECT  107.81 127.795 107.99 125.82 ;
      RECT  107.09 127.795 107.27 125.82 ;
      RECT  106.73 127.795 106.91 125.82 ;
      RECT  109.13 127.795 109.31 125.82 ;
      RECT  109.49 127.795 109.67 125.82 ;
      RECT  110.21 127.795 110.39 125.82 ;
      RECT  110.57 127.795 110.75 125.82 ;
      RECT  114.41 127.795 114.59 125.82 ;
      RECT  114.05 127.795 114.23 125.82 ;
      RECT  113.33 127.795 113.51 125.82 ;
      RECT  112.97 127.795 113.15 125.82 ;
      RECT  115.37 127.795 115.55 125.82 ;
      RECT  115.73 127.795 115.91 125.82 ;
      RECT  116.45 127.795 116.63 125.82 ;
      RECT  116.81 127.795 116.99 125.82 ;
      RECT  120.65 127.795 120.83 125.82 ;
      RECT  120.29 127.795 120.47 125.82 ;
      RECT  119.57 127.795 119.75 125.82 ;
      RECT  119.21 127.795 119.39 125.82 ;
      RECT  121.61 127.795 121.79 125.82 ;
      RECT  121.97 127.795 122.15 125.82 ;
      RECT  122.69 127.795 122.87 125.82 ;
      RECT  123.05 127.795 123.23 125.82 ;
      RECT  126.89 127.795 127.07 125.82 ;
      RECT  126.53 127.795 126.71 125.82 ;
      RECT  125.81 127.795 125.99 125.82 ;
      RECT  125.45 127.795 125.63 125.82 ;
      RECT  127.85 127.795 128.03 125.82 ;
      RECT  128.21 127.795 128.39 125.82 ;
      RECT  128.93 127.795 129.11 125.82 ;
      RECT  129.29 127.795 129.47 125.82 ;
      RECT  133.13 127.795 133.31 125.82 ;
      RECT  132.77 127.795 132.95 125.82 ;
      RECT  132.05 127.795 132.23 125.82 ;
      RECT  131.69 127.795 131.87 125.82 ;
      RECT  134.09 127.795 134.27 125.82 ;
      RECT  134.45 127.795 134.63 125.82 ;
      RECT  135.17 127.795 135.35 125.82 ;
      RECT  135.53 127.795 135.71 125.82 ;
      RECT  139.37 127.795 139.55 125.82 ;
      RECT  139.01 127.795 139.19 125.82 ;
      RECT  138.29 127.795 138.47 125.82 ;
      RECT  137.93 127.795 138.11 125.82 ;
      RECT  140.33 127.795 140.51 125.82 ;
      RECT  140.69 127.795 140.87 125.82 ;
      RECT  141.41 127.795 141.59 125.82 ;
      RECT  141.77 127.795 141.95 125.82 ;
      RECT  145.61 127.795 145.79 125.82 ;
      RECT  145.25 127.795 145.43 125.82 ;
      RECT  144.53 127.795 144.71 125.82 ;
      RECT  144.17 127.795 144.35 125.82 ;
      RECT  96.65 88.295 96.83 127.795 ;
      RECT  97.01 88.295 97.19 127.795 ;
      RECT  97.73 88.295 97.91 127.795 ;
      RECT  98.09 88.295 98.27 127.795 ;
      RECT  101.93 88.295 102.11 127.795 ;
      RECT  101.57 88.295 101.75 127.795 ;
      RECT  100.85 88.295 101.03 127.795 ;
      RECT  100.49 88.295 100.67 127.795 ;
      RECT  102.89 88.295 103.07 127.795 ;
      RECT  103.25 88.295 103.43 127.795 ;
      RECT  103.97 88.295 104.15 127.795 ;
      RECT  104.33 88.295 104.51 127.795 ;
      RECT  108.17 88.295 108.35 127.795 ;
      RECT  107.81 88.295 107.99 127.795 ;
      RECT  107.09 88.295 107.27 127.795 ;
      RECT  106.73 88.295 106.91 127.795 ;
      RECT  109.13 88.295 109.31 127.795 ;
      RECT  109.49 88.295 109.67 127.795 ;
      RECT  110.21 88.295 110.39 127.795 ;
      RECT  110.57 88.295 110.75 127.795 ;
      RECT  114.41 88.295 114.59 127.795 ;
      RECT  114.05 88.295 114.23 127.795 ;
      RECT  113.33 88.295 113.51 127.795 ;
      RECT  112.97 88.295 113.15 127.795 ;
      RECT  115.37 88.295 115.55 127.795 ;
      RECT  115.73 88.295 115.91 127.795 ;
      RECT  116.45 88.295 116.63 127.795 ;
      RECT  116.81 88.295 116.99 127.795 ;
      RECT  120.65 88.295 120.83 127.795 ;
      RECT  120.29 88.295 120.47 127.795 ;
      RECT  119.57 88.295 119.75 127.795 ;
      RECT  119.21 88.295 119.39 127.795 ;
      RECT  121.61 88.295 121.79 127.795 ;
      RECT  121.97 88.295 122.15 127.795 ;
      RECT  122.69 88.295 122.87 127.795 ;
      RECT  123.05 88.295 123.23 127.795 ;
      RECT  126.89 88.295 127.07 127.795 ;
      RECT  126.53 88.295 126.71 127.795 ;
      RECT  125.81 88.295 125.99 127.795 ;
      RECT  125.45 88.295 125.63 127.795 ;
      RECT  127.85 88.295 128.03 127.795 ;
      RECT  128.21 88.295 128.39 127.795 ;
      RECT  128.93 88.295 129.11 127.795 ;
      RECT  129.29 88.295 129.47 127.795 ;
      RECT  133.13 88.295 133.31 127.795 ;
      RECT  132.77 88.295 132.95 127.795 ;
      RECT  132.05 88.295 132.23 127.795 ;
      RECT  131.69 88.295 131.87 127.795 ;
      RECT  134.09 88.295 134.27 127.795 ;
      RECT  134.45 88.295 134.63 127.795 ;
      RECT  135.17 88.295 135.35 127.795 ;
      RECT  135.53 88.295 135.71 127.795 ;
      RECT  139.37 88.295 139.55 127.795 ;
      RECT  139.01 88.295 139.19 127.795 ;
      RECT  138.29 88.295 138.47 127.795 ;
      RECT  137.93 88.295 138.11 127.795 ;
      RECT  140.33 88.295 140.51 127.795 ;
      RECT  140.69 88.295 140.87 127.795 ;
      RECT  141.41 88.295 141.59 127.795 ;
      RECT  141.77 88.295 141.95 127.795 ;
      RECT  145.61 88.295 145.79 127.795 ;
      RECT  145.25 88.295 145.43 127.795 ;
      RECT  144.53 88.295 144.71 127.795 ;
      RECT  144.17 88.295 144.35 127.795 ;
      RECT  95.69 88.295 95.87 127.795 ;
      RECT  95.33 88.295 95.51 127.795 ;
      RECT  147.65 88.295 147.83 127.795 ;
      RECT  148.01 88.295 148.19 127.795 ;
      RECT  147.29 112.39 147.47 114.095 ;
      RECT  94.97 101.995 95.15 103.7 ;
      RECT  94.97 113.845 95.15 115.55 ;
      RECT  94.97 121.745 95.15 123.45 ;
      RECT  147.29 117.795 147.47 119.5 ;
      RECT  94.97 94.095 95.15 95.8 ;
      RECT  94.97 109.895 95.15 111.6 ;
      RECT  147.29 98.045 147.47 99.75 ;
      RECT  94.97 90.145 95.15 91.85 ;
      RECT  94.97 124.24 95.15 125.945 ;
      RECT  147.29 90.145 147.47 91.85 ;
      RECT  147.29 92.64 147.47 94.345 ;
      RECT  147.29 113.845 147.47 115.55 ;
      RECT  94.97 96.59 95.15 98.295 ;
      RECT  94.97 117.795 95.15 119.5 ;
      RECT  147.29 120.29 147.47 121.995 ;
      RECT  147.29 116.34 147.47 118.045 ;
      RECT  147.29 124.24 147.47 125.945 ;
      RECT  94.97 108.44 95.15 110.145 ;
      RECT  147.29 101.995 147.47 103.7 ;
      RECT  94.97 120.29 95.15 121.995 ;
      RECT  147.29 105.945 147.47 107.65 ;
      RECT  94.97 100.54 95.15 102.245 ;
      RECT  94.97 105.945 95.15 107.65 ;
      RECT  94.97 104.49 95.15 106.195 ;
      RECT  147.29 108.44 147.47 110.145 ;
      RECT  147.29 109.895 147.47 111.6 ;
      RECT  94.97 116.34 95.15 118.045 ;
      RECT  94.97 112.39 95.15 114.095 ;
      RECT  147.29 121.745 147.47 123.45 ;
      RECT  94.97 92.64 95.15 94.345 ;
      RECT  147.29 94.095 147.47 95.8 ;
      RECT  147.29 100.54 147.47 102.245 ;
      RECT  147.29 104.49 147.47 106.195 ;
      RECT  147.29 96.59 147.47 98.295 ;
      RECT  94.97 98.045 95.15 99.75 ;
      RECT  95.93 83.265 95.79 87.035 ;
      RECT  93.61 83.265 93.47 87.035 ;
      RECT  96.59 83.265 96.73 87.035 ;
      RECT  98.91 83.265 99.05 87.035 ;
      RECT  102.17 83.265 102.03 87.035 ;
      RECT  99.85 83.265 99.71 87.035 ;
      RECT  102.83 83.265 102.97 87.035 ;
      RECT  105.15 83.265 105.29 87.035 ;
      RECT  108.41 83.265 108.27 87.035 ;
      RECT  106.09 83.265 105.95 87.035 ;
      RECT  109.07 83.265 109.21 87.035 ;
      RECT  111.39 83.265 111.53 87.035 ;
      RECT  114.65 83.265 114.51 87.035 ;
      RECT  112.33 83.265 112.19 87.035 ;
      RECT  115.31 83.265 115.45 87.035 ;
      RECT  117.63 83.265 117.77 87.035 ;
      RECT  120.89 83.265 120.75 87.035 ;
      RECT  118.57 83.265 118.43 87.035 ;
      RECT  121.55 83.265 121.69 87.035 ;
      RECT  123.87 83.265 124.01 87.035 ;
      RECT  127.13 83.265 126.99 87.035 ;
      RECT  124.81 83.265 124.67 87.035 ;
      RECT  127.79 83.265 127.93 87.035 ;
      RECT  130.11 83.265 130.25 87.035 ;
      RECT  133.37 83.265 133.23 87.035 ;
      RECT  131.05 83.265 130.91 87.035 ;
      RECT  134.03 83.265 134.17 87.035 ;
      RECT  136.35 83.265 136.49 87.035 ;
      RECT  139.61 83.265 139.47 87.035 ;
      RECT  137.29 83.265 137.15 87.035 ;
      RECT  140.27 83.265 140.41 87.035 ;
      RECT  142.59 83.265 142.73 87.035 ;
      RECT  145.85 83.265 145.71 87.035 ;
      RECT  143.53 83.265 143.39 87.035 ;
      RECT  95.79 83.265 95.93 87.035 ;
      RECT  93.47 83.265 93.61 87.035 ;
      RECT  96.59 83.265 96.73 87.035 ;
      RECT  98.91 83.265 99.05 87.035 ;
      RECT  102.03 83.265 102.17 87.035 ;
      RECT  99.71 83.265 99.85 87.035 ;
      RECT  102.83 83.265 102.97 87.035 ;
      RECT  105.15 83.265 105.29 87.035 ;
      RECT  108.27 83.265 108.41 87.035 ;
      RECT  105.95 83.265 106.09 87.035 ;
      RECT  109.07 83.265 109.21 87.035 ;
      RECT  111.39 83.265 111.53 87.035 ;
      RECT  114.51 83.265 114.65 87.035 ;
      RECT  112.19 83.265 112.33 87.035 ;
      RECT  115.31 83.265 115.45 87.035 ;
      RECT  117.63 83.265 117.77 87.035 ;
      RECT  120.75 83.265 120.89 87.035 ;
      RECT  118.43 83.265 118.57 87.035 ;
      RECT  121.55 83.265 121.69 87.035 ;
      RECT  123.87 83.265 124.01 87.035 ;
      RECT  126.99 83.265 127.13 87.035 ;
      RECT  124.67 83.265 124.81 87.035 ;
      RECT  127.79 83.265 127.93 87.035 ;
      RECT  130.11 83.265 130.25 87.035 ;
      RECT  133.23 83.265 133.37 87.035 ;
      RECT  130.91 83.265 131.05 87.035 ;
      RECT  134.03 83.265 134.17 87.035 ;
      RECT  136.35 83.265 136.49 87.035 ;
      RECT  139.47 83.265 139.61 87.035 ;
      RECT  137.15 83.265 137.29 87.035 ;
      RECT  140.27 83.265 140.41 87.035 ;
      RECT  142.59 83.265 142.73 87.035 ;
      RECT  145.71 83.265 145.85 87.035 ;
      RECT  143.39 83.265 143.53 87.035 ;
      RECT  97.62 76.435 97.76 82.005 ;
      RECT  97.62 76.145 97.96 76.435 ;
      RECT  97.24 76.375 97.41 82.005 ;
      RECT  98.4 80.75 98.63 81.12 ;
      RECT  96.73 81.545 97.02 81.845 ;
      RECT  97.95 76.895 98.26 77.235 ;
      RECT  98.05 72.685 98.28 73.065 ;
      RECT  98.05 71.08 98.28 71.45 ;
      RECT  96.78 70.725 97.01 71.995 ;
      RECT  97.24 70.725 97.41 76.145 ;
      RECT  97.18 76.145 97.47 76.375 ;
      RECT  97.62 70.725 97.76 76.145 ;
      RECT  100.52 76.435 100.38 82.005 ;
      RECT  100.52 76.145 100.18 76.435 ;
      RECT  100.9 76.375 100.73 82.005 ;
      RECT  99.74 80.75 99.51 81.12 ;
      RECT  101.41 81.545 101.12 81.845 ;
      RECT  100.19 76.895 99.88 77.235 ;
      RECT  100.09 72.685 99.86 73.065 ;
      RECT  100.09 71.08 99.86 71.45 ;
      RECT  101.36 70.725 101.13 71.995 ;
      RECT  100.9 70.725 100.73 76.145 ;
      RECT  100.96 76.145 100.67 76.375 ;
      RECT  100.52 70.725 100.38 76.145 ;
      RECT  103.86 76.435 104.0 82.005 ;
      RECT  103.86 76.145 104.2 76.435 ;
      RECT  103.48 76.375 103.65 82.005 ;
      RECT  104.64 80.75 104.87 81.12 ;
      RECT  102.97 81.545 103.26 81.845 ;
      RECT  104.19 76.895 104.5 77.235 ;
      RECT  104.29 72.685 104.52 73.065 ;
      RECT  104.29 71.08 104.52 71.45 ;
      RECT  103.02 70.725 103.25 71.995 ;
      RECT  103.48 70.725 103.65 76.145 ;
      RECT  103.42 76.145 103.71 76.375 ;
      RECT  103.86 70.725 104.0 76.145 ;
      RECT  106.76 76.435 106.62 82.005 ;
      RECT  106.76 76.145 106.42 76.435 ;
      RECT  107.14 76.375 106.97 82.005 ;
      RECT  105.98 80.75 105.75 81.12 ;
      RECT  107.65 81.545 107.36 81.845 ;
      RECT  106.43 76.895 106.12 77.235 ;
      RECT  106.33 72.685 106.1 73.065 ;
      RECT  106.33 71.08 106.1 71.45 ;
      RECT  107.6 70.725 107.37 71.995 ;
      RECT  107.14 70.725 106.97 76.145 ;
      RECT  107.2 76.145 106.91 76.375 ;
      RECT  106.76 70.725 106.62 76.145 ;
      RECT  110.1 76.435 110.24 82.005 ;
      RECT  110.1 76.145 110.44 76.435 ;
      RECT  109.72 76.375 109.89 82.005 ;
      RECT  110.88 80.75 111.11 81.12 ;
      RECT  109.21 81.545 109.5 81.845 ;
      RECT  110.43 76.895 110.74 77.235 ;
      RECT  110.53 72.685 110.76 73.065 ;
      RECT  110.53 71.08 110.76 71.45 ;
      RECT  109.26 70.725 109.49 71.995 ;
      RECT  109.72 70.725 109.89 76.145 ;
      RECT  109.66 76.145 109.95 76.375 ;
      RECT  110.1 70.725 110.24 76.145 ;
      RECT  113.0 76.435 112.86 82.005 ;
      RECT  113.0 76.145 112.66 76.435 ;
      RECT  113.38 76.375 113.21 82.005 ;
      RECT  112.22 80.75 111.99 81.12 ;
      RECT  113.89 81.545 113.6 81.845 ;
      RECT  112.67 76.895 112.36 77.235 ;
      RECT  112.57 72.685 112.34 73.065 ;
      RECT  112.57 71.08 112.34 71.45 ;
      RECT  113.84 70.725 113.61 71.995 ;
      RECT  113.38 70.725 113.21 76.145 ;
      RECT  113.44 76.145 113.15 76.375 ;
      RECT  113.0 70.725 112.86 76.145 ;
      RECT  116.34 76.435 116.48 82.005 ;
      RECT  116.34 76.145 116.68 76.435 ;
      RECT  115.96 76.375 116.13 82.005 ;
      RECT  117.12 80.75 117.35 81.12 ;
      RECT  115.45 81.545 115.74 81.845 ;
      RECT  116.67 76.895 116.98 77.235 ;
      RECT  116.77 72.685 117.0 73.065 ;
      RECT  116.77 71.08 117.0 71.45 ;
      RECT  115.5 70.725 115.73 71.995 ;
      RECT  115.96 70.725 116.13 76.145 ;
      RECT  115.9 76.145 116.19 76.375 ;
      RECT  116.34 70.725 116.48 76.145 ;
      RECT  119.24 76.435 119.1 82.005 ;
      RECT  119.24 76.145 118.9 76.435 ;
      RECT  119.62 76.375 119.45 82.005 ;
      RECT  118.46 80.75 118.23 81.12 ;
      RECT  120.13 81.545 119.84 81.845 ;
      RECT  118.91 76.895 118.6 77.235 ;
      RECT  118.81 72.685 118.58 73.065 ;
      RECT  118.81 71.08 118.58 71.45 ;
      RECT  120.08 70.725 119.85 71.995 ;
      RECT  119.62 70.725 119.45 76.145 ;
      RECT  119.68 76.145 119.39 76.375 ;
      RECT  119.24 70.725 119.1 76.145 ;
      RECT  122.58 76.435 122.72 82.005 ;
      RECT  122.58 76.145 122.92 76.435 ;
      RECT  122.2 76.375 122.37 82.005 ;
      RECT  123.36 80.75 123.59 81.12 ;
      RECT  121.69 81.545 121.98 81.845 ;
      RECT  122.91 76.895 123.22 77.235 ;
      RECT  123.01 72.685 123.24 73.065 ;
      RECT  123.01 71.08 123.24 71.45 ;
      RECT  121.74 70.725 121.97 71.995 ;
      RECT  122.2 70.725 122.37 76.145 ;
      RECT  122.14 76.145 122.43 76.375 ;
      RECT  122.58 70.725 122.72 76.145 ;
      RECT  125.48 76.435 125.34 82.005 ;
      RECT  125.48 76.145 125.14 76.435 ;
      RECT  125.86 76.375 125.69 82.005 ;
      RECT  124.7 80.75 124.47 81.12 ;
      RECT  126.37 81.545 126.08 81.845 ;
      RECT  125.15 76.895 124.84 77.235 ;
      RECT  125.05 72.685 124.82 73.065 ;
      RECT  125.05 71.08 124.82 71.45 ;
      RECT  126.32 70.725 126.09 71.995 ;
      RECT  125.86 70.725 125.69 76.145 ;
      RECT  125.92 76.145 125.63 76.375 ;
      RECT  125.48 70.725 125.34 76.145 ;
      RECT  128.82 76.435 128.96 82.005 ;
      RECT  128.82 76.145 129.16 76.435 ;
      RECT  128.44 76.375 128.61 82.005 ;
      RECT  129.6 80.75 129.83 81.12 ;
      RECT  127.93 81.545 128.22 81.845 ;
      RECT  129.15 76.895 129.46 77.235 ;
      RECT  129.25 72.685 129.48 73.065 ;
      RECT  129.25 71.08 129.48 71.45 ;
      RECT  127.98 70.725 128.21 71.995 ;
      RECT  128.44 70.725 128.61 76.145 ;
      RECT  128.38 76.145 128.67 76.375 ;
      RECT  128.82 70.725 128.96 76.145 ;
      RECT  131.72 76.435 131.58 82.005 ;
      RECT  131.72 76.145 131.38 76.435 ;
      RECT  132.1 76.375 131.93 82.005 ;
      RECT  130.94 80.75 130.71 81.12 ;
      RECT  132.61 81.545 132.32 81.845 ;
      RECT  131.39 76.895 131.08 77.235 ;
      RECT  131.29 72.685 131.06 73.065 ;
      RECT  131.29 71.08 131.06 71.45 ;
      RECT  132.56 70.725 132.33 71.995 ;
      RECT  132.1 70.725 131.93 76.145 ;
      RECT  132.16 76.145 131.87 76.375 ;
      RECT  131.72 70.725 131.58 76.145 ;
      RECT  135.06 76.435 135.2 82.005 ;
      RECT  135.06 76.145 135.4 76.435 ;
      RECT  134.68 76.375 134.85 82.005 ;
      RECT  135.84 80.75 136.07 81.12 ;
      RECT  134.17 81.545 134.46 81.845 ;
      RECT  135.39 76.895 135.7 77.235 ;
      RECT  135.49 72.685 135.72 73.065 ;
      RECT  135.49 71.08 135.72 71.45 ;
      RECT  134.22 70.725 134.45 71.995 ;
      RECT  134.68 70.725 134.85 76.145 ;
      RECT  134.62 76.145 134.91 76.375 ;
      RECT  135.06 70.725 135.2 76.145 ;
      RECT  137.96 76.435 137.82 82.005 ;
      RECT  137.96 76.145 137.62 76.435 ;
      RECT  138.34 76.375 138.17 82.005 ;
      RECT  137.18 80.75 136.95 81.12 ;
      RECT  138.85 81.545 138.56 81.845 ;
      RECT  137.63 76.895 137.32 77.235 ;
      RECT  137.53 72.685 137.3 73.065 ;
      RECT  137.53 71.08 137.3 71.45 ;
      RECT  138.8 70.725 138.57 71.995 ;
      RECT  138.34 70.725 138.17 76.145 ;
      RECT  138.4 76.145 138.11 76.375 ;
      RECT  137.96 70.725 137.82 76.145 ;
      RECT  141.3 76.435 141.44 82.005 ;
      RECT  141.3 76.145 141.64 76.435 ;
      RECT  140.92 76.375 141.09 82.005 ;
      RECT  142.08 80.75 142.31 81.12 ;
      RECT  140.41 81.545 140.7 81.845 ;
      RECT  141.63 76.895 141.94 77.235 ;
      RECT  141.73 72.685 141.96 73.065 ;
      RECT  141.73 71.08 141.96 71.45 ;
      RECT  140.46 70.725 140.69 71.995 ;
      RECT  140.92 70.725 141.09 76.145 ;
      RECT  140.86 76.145 141.15 76.375 ;
      RECT  141.3 70.725 141.44 76.145 ;
      RECT  144.2 76.435 144.06 82.005 ;
      RECT  144.2 76.145 143.86 76.435 ;
      RECT  144.58 76.375 144.41 82.005 ;
      RECT  143.42 80.75 143.19 81.12 ;
      RECT  145.09 81.545 144.8 81.845 ;
      RECT  143.87 76.895 143.56 77.235 ;
      RECT  143.77 72.685 143.54 73.065 ;
      RECT  143.77 71.08 143.54 71.45 ;
      RECT  145.04 70.725 144.81 71.995 ;
      RECT  144.58 70.725 144.41 76.145 ;
      RECT  144.64 76.145 144.35 76.375 ;
      RECT  144.2 70.725 144.06 76.145 ;
      RECT  96.78 70.725 97.01 71.995 ;
      RECT  97.24 76.375 97.41 82.005 ;
      RECT  97.62 76.435 97.76 82.005 ;
      RECT  101.13 70.725 101.36 71.995 ;
      RECT  100.73 76.375 100.9 82.005 ;
      RECT  100.38 76.435 100.52 82.005 ;
      RECT  103.02 70.725 103.25 71.995 ;
      RECT  103.48 76.375 103.65 82.005 ;
      RECT  103.86 76.435 104.0 82.005 ;
      RECT  107.37 70.725 107.6 71.995 ;
      RECT  106.97 76.375 107.14 82.005 ;
      RECT  106.62 76.435 106.76 82.005 ;
      RECT  109.26 70.725 109.49 71.995 ;
      RECT  109.72 76.375 109.89 82.005 ;
      RECT  110.1 76.435 110.24 82.005 ;
      RECT  113.61 70.725 113.84 71.995 ;
      RECT  113.21 76.375 113.38 82.005 ;
      RECT  112.86 76.435 113.0 82.005 ;
      RECT  115.5 70.725 115.73 71.995 ;
      RECT  115.96 76.375 116.13 82.005 ;
      RECT  116.34 76.435 116.48 82.005 ;
      RECT  119.85 70.725 120.08 71.995 ;
      RECT  119.45 76.375 119.62 82.005 ;
      RECT  119.1 76.435 119.24 82.005 ;
      RECT  121.74 70.725 121.97 71.995 ;
      RECT  122.2 76.375 122.37 82.005 ;
      RECT  122.58 76.435 122.72 82.005 ;
      RECT  126.09 70.725 126.32 71.995 ;
      RECT  125.69 76.375 125.86 82.005 ;
      RECT  125.34 76.435 125.48 82.005 ;
      RECT  127.98 70.725 128.21 71.995 ;
      RECT  128.44 76.375 128.61 82.005 ;
      RECT  128.82 76.435 128.96 82.005 ;
      RECT  132.33 70.725 132.56 71.995 ;
      RECT  131.93 76.375 132.1 82.005 ;
      RECT  131.58 76.435 131.72 82.005 ;
      RECT  134.22 70.725 134.45 71.995 ;
      RECT  134.68 76.375 134.85 82.005 ;
      RECT  135.06 76.435 135.2 82.005 ;
      RECT  138.57 70.725 138.8 71.995 ;
      RECT  138.17 76.375 138.34 82.005 ;
      RECT  137.82 76.435 137.96 82.005 ;
      RECT  140.46 70.725 140.69 71.995 ;
      RECT  140.92 76.375 141.09 82.005 ;
      RECT  141.3 76.435 141.44 82.005 ;
      RECT  144.81 70.725 145.04 71.995 ;
      RECT  144.41 76.375 144.58 82.005 ;
      RECT  144.06 76.435 144.2 82.005 ;
      RECT  97.995 63.33 98.36 63.355 ;
      RECT  97.325 67.185 97.755 67.215 ;
      RECT  97.77 68.915 98.055 69.205 ;
      RECT  97.9 69.205 98.05 69.465 ;
      RECT  96.755 59.88 98.76 60.05 ;
      RECT  96.755 60.05 97.045 60.19 ;
      RECT  97.325 65.0 97.755 65.23 ;
      RECT  97.355 62.33 97.785 62.56 ;
      RECT  97.325 67.215 97.865 67.385 ;
      RECT  97.425 60.25 97.855 60.48 ;
      RECT  97.535 59.43 97.835 59.71 ;
      RECT  96.89 69.205 97.04 69.465 ;
      RECT  97.93 63.355 98.36 63.56 ;
      RECT  96.885 68.915 97.17 69.205 ;
      RECT  97.325 67.385 97.755 67.415 ;
      RECT  100.145 63.33 99.78 63.355 ;
      RECT  100.815 67.185 100.385 67.215 ;
      RECT  100.37 68.915 100.085 69.205 ;
      RECT  100.24 69.205 100.09 69.465 ;
      RECT  101.385 59.88 99.38 60.05 ;
      RECT  101.385 60.05 101.095 60.19 ;
      RECT  100.815 65.0 100.385 65.23 ;
      RECT  100.785 62.33 100.355 62.56 ;
      RECT  100.815 67.215 100.275 67.385 ;
      RECT  100.715 60.25 100.285 60.48 ;
      RECT  100.605 59.43 100.305 59.71 ;
      RECT  101.25 69.205 101.1 69.465 ;
      RECT  100.21 63.355 99.78 63.56 ;
      RECT  101.255 68.915 100.97 69.205 ;
      RECT  100.815 67.385 100.385 67.415 ;
      RECT  104.235 63.33 104.6 63.355 ;
      RECT  103.565 67.185 103.995 67.215 ;
      RECT  104.01 68.915 104.295 69.205 ;
      RECT  104.14 69.205 104.29 69.465 ;
      RECT  102.995 59.88 105.0 60.05 ;
      RECT  102.995 60.05 103.285 60.19 ;
      RECT  103.565 65.0 103.995 65.23 ;
      RECT  103.595 62.33 104.025 62.56 ;
      RECT  103.565 67.215 104.105 67.385 ;
      RECT  103.665 60.25 104.095 60.48 ;
      RECT  103.775 59.43 104.075 59.71 ;
      RECT  103.13 69.205 103.28 69.465 ;
      RECT  104.17 63.355 104.6 63.56 ;
      RECT  103.125 68.915 103.41 69.205 ;
      RECT  103.565 67.385 103.995 67.415 ;
      RECT  106.385 63.33 106.02 63.355 ;
      RECT  107.055 67.185 106.625 67.215 ;
      RECT  106.61 68.915 106.325 69.205 ;
      RECT  106.48 69.205 106.33 69.465 ;
      RECT  107.625 59.88 105.62 60.05 ;
      RECT  107.625 60.05 107.335 60.19 ;
      RECT  107.055 65.0 106.625 65.23 ;
      RECT  107.025 62.33 106.595 62.56 ;
      RECT  107.055 67.215 106.515 67.385 ;
      RECT  106.955 60.25 106.525 60.48 ;
      RECT  106.845 59.43 106.545 59.71 ;
      RECT  107.49 69.205 107.34 69.465 ;
      RECT  106.45 63.355 106.02 63.56 ;
      RECT  107.495 68.915 107.21 69.205 ;
      RECT  107.055 67.385 106.625 67.415 ;
      RECT  110.475 63.33 110.84 63.355 ;
      RECT  109.805 67.185 110.235 67.215 ;
      RECT  110.25 68.915 110.535 69.205 ;
      RECT  110.38 69.205 110.53 69.465 ;
      RECT  109.235 59.88 111.24 60.05 ;
      RECT  109.235 60.05 109.525 60.19 ;
      RECT  109.805 65.0 110.235 65.23 ;
      RECT  109.835 62.33 110.265 62.56 ;
      RECT  109.805 67.215 110.345 67.385 ;
      RECT  109.905 60.25 110.335 60.48 ;
      RECT  110.015 59.43 110.315 59.71 ;
      RECT  109.37 69.205 109.52 69.465 ;
      RECT  110.41 63.355 110.84 63.56 ;
      RECT  109.365 68.915 109.65 69.205 ;
      RECT  109.805 67.385 110.235 67.415 ;
      RECT  112.625 63.33 112.26 63.355 ;
      RECT  113.295 67.185 112.865 67.215 ;
      RECT  112.85 68.915 112.565 69.205 ;
      RECT  112.72 69.205 112.57 69.465 ;
      RECT  113.865 59.88 111.86 60.05 ;
      RECT  113.865 60.05 113.575 60.19 ;
      RECT  113.295 65.0 112.865 65.23 ;
      RECT  113.265 62.33 112.835 62.56 ;
      RECT  113.295 67.215 112.755 67.385 ;
      RECT  113.195 60.25 112.765 60.48 ;
      RECT  113.085 59.43 112.785 59.71 ;
      RECT  113.73 69.205 113.58 69.465 ;
      RECT  112.69 63.355 112.26 63.56 ;
      RECT  113.735 68.915 113.45 69.205 ;
      RECT  113.295 67.385 112.865 67.415 ;
      RECT  116.715 63.33 117.08 63.355 ;
      RECT  116.045 67.185 116.475 67.215 ;
      RECT  116.49 68.915 116.775 69.205 ;
      RECT  116.62 69.205 116.77 69.465 ;
      RECT  115.475 59.88 117.48 60.05 ;
      RECT  115.475 60.05 115.765 60.19 ;
      RECT  116.045 65.0 116.475 65.23 ;
      RECT  116.075 62.33 116.505 62.56 ;
      RECT  116.045 67.215 116.585 67.385 ;
      RECT  116.145 60.25 116.575 60.48 ;
      RECT  116.255 59.43 116.555 59.71 ;
      RECT  115.61 69.205 115.76 69.465 ;
      RECT  116.65 63.355 117.08 63.56 ;
      RECT  115.605 68.915 115.89 69.205 ;
      RECT  116.045 67.385 116.475 67.415 ;
      RECT  118.865 63.33 118.5 63.355 ;
      RECT  119.535 67.185 119.105 67.215 ;
      RECT  119.09 68.915 118.805 69.205 ;
      RECT  118.96 69.205 118.81 69.465 ;
      RECT  120.105 59.88 118.1 60.05 ;
      RECT  120.105 60.05 119.815 60.19 ;
      RECT  119.535 65.0 119.105 65.23 ;
      RECT  119.505 62.33 119.075 62.56 ;
      RECT  119.535 67.215 118.995 67.385 ;
      RECT  119.435 60.25 119.005 60.48 ;
      RECT  119.325 59.43 119.025 59.71 ;
      RECT  119.97 69.205 119.82 69.465 ;
      RECT  118.93 63.355 118.5 63.56 ;
      RECT  119.975 68.915 119.69 69.205 ;
      RECT  119.535 67.385 119.105 67.415 ;
      RECT  122.955 63.33 123.32 63.355 ;
      RECT  122.285 67.185 122.715 67.215 ;
      RECT  122.73 68.915 123.015 69.205 ;
      RECT  122.86 69.205 123.01 69.465 ;
      RECT  121.715 59.88 123.72 60.05 ;
      RECT  121.715 60.05 122.005 60.19 ;
      RECT  122.285 65.0 122.715 65.23 ;
      RECT  122.315 62.33 122.745 62.56 ;
      RECT  122.285 67.215 122.825 67.385 ;
      RECT  122.385 60.25 122.815 60.48 ;
      RECT  122.495 59.43 122.795 59.71 ;
      RECT  121.85 69.205 122.0 69.465 ;
      RECT  122.89 63.355 123.32 63.56 ;
      RECT  121.845 68.915 122.13 69.205 ;
      RECT  122.285 67.385 122.715 67.415 ;
      RECT  125.105 63.33 124.74 63.355 ;
      RECT  125.775 67.185 125.345 67.215 ;
      RECT  125.33 68.915 125.045 69.205 ;
      RECT  125.2 69.205 125.05 69.465 ;
      RECT  126.345 59.88 124.34 60.05 ;
      RECT  126.345 60.05 126.055 60.19 ;
      RECT  125.775 65.0 125.345 65.23 ;
      RECT  125.745 62.33 125.315 62.56 ;
      RECT  125.775 67.215 125.235 67.385 ;
      RECT  125.675 60.25 125.245 60.48 ;
      RECT  125.565 59.43 125.265 59.71 ;
      RECT  126.21 69.205 126.06 69.465 ;
      RECT  125.17 63.355 124.74 63.56 ;
      RECT  126.215 68.915 125.93 69.205 ;
      RECT  125.775 67.385 125.345 67.415 ;
      RECT  129.195 63.33 129.56 63.355 ;
      RECT  128.525 67.185 128.955 67.215 ;
      RECT  128.97 68.915 129.255 69.205 ;
      RECT  129.1 69.205 129.25 69.465 ;
      RECT  127.955 59.88 129.96 60.05 ;
      RECT  127.955 60.05 128.245 60.19 ;
      RECT  128.525 65.0 128.955 65.23 ;
      RECT  128.555 62.33 128.985 62.56 ;
      RECT  128.525 67.215 129.065 67.385 ;
      RECT  128.625 60.25 129.055 60.48 ;
      RECT  128.735 59.43 129.035 59.71 ;
      RECT  128.09 69.205 128.24 69.465 ;
      RECT  129.13 63.355 129.56 63.56 ;
      RECT  128.085 68.915 128.37 69.205 ;
      RECT  128.525 67.385 128.955 67.415 ;
      RECT  131.345 63.33 130.98 63.355 ;
      RECT  132.015 67.185 131.585 67.215 ;
      RECT  131.57 68.915 131.285 69.205 ;
      RECT  131.44 69.205 131.29 69.465 ;
      RECT  132.585 59.88 130.58 60.05 ;
      RECT  132.585 60.05 132.295 60.19 ;
      RECT  132.015 65.0 131.585 65.23 ;
      RECT  131.985 62.33 131.555 62.56 ;
      RECT  132.015 67.215 131.475 67.385 ;
      RECT  131.915 60.25 131.485 60.48 ;
      RECT  131.805 59.43 131.505 59.71 ;
      RECT  132.45 69.205 132.3 69.465 ;
      RECT  131.41 63.355 130.98 63.56 ;
      RECT  132.455 68.915 132.17 69.205 ;
      RECT  132.015 67.385 131.585 67.415 ;
      RECT  135.435 63.33 135.8 63.355 ;
      RECT  134.765 67.185 135.195 67.215 ;
      RECT  135.21 68.915 135.495 69.205 ;
      RECT  135.34 69.205 135.49 69.465 ;
      RECT  134.195 59.88 136.2 60.05 ;
      RECT  134.195 60.05 134.485 60.19 ;
      RECT  134.765 65.0 135.195 65.23 ;
      RECT  134.795 62.33 135.225 62.56 ;
      RECT  134.765 67.215 135.305 67.385 ;
      RECT  134.865 60.25 135.295 60.48 ;
      RECT  134.975 59.43 135.275 59.71 ;
      RECT  134.33 69.205 134.48 69.465 ;
      RECT  135.37 63.355 135.8 63.56 ;
      RECT  134.325 68.915 134.61 69.205 ;
      RECT  134.765 67.385 135.195 67.415 ;
      RECT  137.585 63.33 137.22 63.355 ;
      RECT  138.255 67.185 137.825 67.215 ;
      RECT  137.81 68.915 137.525 69.205 ;
      RECT  137.68 69.205 137.53 69.465 ;
      RECT  138.825 59.88 136.82 60.05 ;
      RECT  138.825 60.05 138.535 60.19 ;
      RECT  138.255 65.0 137.825 65.23 ;
      RECT  138.225 62.33 137.795 62.56 ;
      RECT  138.255 67.215 137.715 67.385 ;
      RECT  138.155 60.25 137.725 60.48 ;
      RECT  138.045 59.43 137.745 59.71 ;
      RECT  138.69 69.205 138.54 69.465 ;
      RECT  137.65 63.355 137.22 63.56 ;
      RECT  138.695 68.915 138.41 69.205 ;
      RECT  138.255 67.385 137.825 67.415 ;
      RECT  141.675 63.33 142.04 63.355 ;
      RECT  141.005 67.185 141.435 67.215 ;
      RECT  141.45 68.915 141.735 69.205 ;
      RECT  141.58 69.205 141.73 69.465 ;
      RECT  140.435 59.88 142.44 60.05 ;
      RECT  140.435 60.05 140.725 60.19 ;
      RECT  141.005 65.0 141.435 65.23 ;
      RECT  141.035 62.33 141.465 62.56 ;
      RECT  141.005 67.215 141.545 67.385 ;
      RECT  141.105 60.25 141.535 60.48 ;
      RECT  141.215 59.43 141.515 59.71 ;
      RECT  140.57 69.205 140.72 69.465 ;
      RECT  141.61 63.355 142.04 63.56 ;
      RECT  140.565 68.915 140.85 69.205 ;
      RECT  141.005 67.385 141.435 67.415 ;
      RECT  143.825 63.33 143.46 63.355 ;
      RECT  144.495 67.185 144.065 67.215 ;
      RECT  144.05 68.915 143.765 69.205 ;
      RECT  143.92 69.205 143.77 69.465 ;
      RECT  145.065 59.88 143.06 60.05 ;
      RECT  145.065 60.05 144.775 60.19 ;
      RECT  144.495 65.0 144.065 65.23 ;
      RECT  144.465 62.33 144.035 62.56 ;
      RECT  144.495 67.215 143.955 67.385 ;
      RECT  144.395 60.25 143.965 60.48 ;
      RECT  144.285 59.43 143.985 59.71 ;
      RECT  144.93 69.205 144.78 69.465 ;
      RECT  143.89 63.355 143.46 63.56 ;
      RECT  144.935 68.915 144.65 69.205 ;
      RECT  144.495 67.385 144.065 67.415 ;
      RECT  97.535 59.43 97.835 59.71 ;
      RECT  100.305 59.43 100.605 59.71 ;
      RECT  103.775 59.43 104.075 59.71 ;
      RECT  106.545 59.43 106.845 59.71 ;
      RECT  110.015 59.43 110.315 59.71 ;
      RECT  112.785 59.43 113.085 59.71 ;
      RECT  116.255 59.43 116.555 59.71 ;
      RECT  119.025 59.43 119.325 59.71 ;
      RECT  122.495 59.43 122.795 59.71 ;
      RECT  125.265 59.43 125.565 59.71 ;
      RECT  128.735 59.43 129.035 59.71 ;
      RECT  131.505 59.43 131.805 59.71 ;
      RECT  134.975 59.43 135.275 59.71 ;
      RECT  137.745 59.43 138.045 59.71 ;
      RECT  141.215 59.43 141.515 59.71 ;
      RECT  143.985 59.43 144.285 59.71 ;
      RECT  96.89 69.205 97.04 69.465 ;
      RECT  97.9 69.205 98.05 69.465 ;
      RECT  101.1 69.205 101.25 69.465 ;
      RECT  100.09 69.205 100.24 69.465 ;
      RECT  103.13 69.205 103.28 69.465 ;
      RECT  104.14 69.205 104.29 69.465 ;
      RECT  107.34 69.205 107.49 69.465 ;
      RECT  106.33 69.205 106.48 69.465 ;
      RECT  109.37 69.205 109.52 69.465 ;
      RECT  110.38 69.205 110.53 69.465 ;
      RECT  113.58 69.205 113.73 69.465 ;
      RECT  112.57 69.205 112.72 69.465 ;
      RECT  115.61 69.205 115.76 69.465 ;
      RECT  116.62 69.205 116.77 69.465 ;
      RECT  119.82 69.205 119.97 69.465 ;
      RECT  118.81 69.205 118.96 69.465 ;
      RECT  121.85 69.205 122.0 69.465 ;
      RECT  122.86 69.205 123.01 69.465 ;
      RECT  126.06 69.205 126.21 69.465 ;
      RECT  125.05 69.205 125.2 69.465 ;
      RECT  128.09 69.205 128.24 69.465 ;
      RECT  129.1 69.205 129.25 69.465 ;
      RECT  132.3 69.205 132.45 69.465 ;
      RECT  131.29 69.205 131.44 69.465 ;
      RECT  134.33 69.205 134.48 69.465 ;
      RECT  135.34 69.205 135.49 69.465 ;
      RECT  138.54 69.205 138.69 69.465 ;
      RECT  137.53 69.205 137.68 69.465 ;
      RECT  140.57 69.205 140.72 69.465 ;
      RECT  141.58 69.205 141.73 69.465 ;
      RECT  144.78 69.205 144.93 69.465 ;
      RECT  143.77 69.205 143.92 69.465 ;
      RECT  96.755 59.88 120.6 60.05 ;
      RECT  121.715 59.88 145.56 60.05 ;
      RECT  95.79 87.035 95.93 83.265 ;
      RECT  93.47 87.035 93.61 83.265 ;
      RECT  96.78 71.995 97.01 70.725 ;
      RECT  101.13 71.995 101.36 70.725 ;
      RECT  103.02 71.995 103.25 70.725 ;
      RECT  107.37 71.995 107.6 70.725 ;
      RECT  109.26 71.995 109.49 70.725 ;
      RECT  113.61 71.995 113.84 70.725 ;
      RECT  115.5 71.995 115.73 70.725 ;
      RECT  119.85 71.995 120.08 70.725 ;
      RECT  121.74 71.995 121.97 70.725 ;
      RECT  126.09 71.995 126.32 70.725 ;
      RECT  127.98 71.995 128.21 70.725 ;
      RECT  132.33 71.995 132.56 70.725 ;
      RECT  134.22 71.995 134.45 70.725 ;
      RECT  138.57 71.995 138.8 70.725 ;
      RECT  140.46 71.995 140.69 70.725 ;
      RECT  144.81 71.995 145.04 70.725 ;
      RECT  97.535 59.71 97.835 59.43 ;
      RECT  100.305 59.71 100.605 59.43 ;
      RECT  103.775 59.71 104.075 59.43 ;
      RECT  106.545 59.71 106.845 59.43 ;
      RECT  110.015 59.71 110.315 59.43 ;
      RECT  112.785 59.71 113.085 59.43 ;
      RECT  116.255 59.71 116.555 59.43 ;
      RECT  119.025 59.71 119.325 59.43 ;
      RECT  122.495 59.71 122.795 59.43 ;
      RECT  125.265 59.71 125.565 59.43 ;
      RECT  128.735 59.71 129.035 59.43 ;
      RECT  131.505 59.71 131.805 59.43 ;
      RECT  134.975 59.71 135.275 59.43 ;
      RECT  137.745 59.71 138.045 59.43 ;
      RECT  141.215 59.71 141.515 59.43 ;
      RECT  143.985 59.71 144.285 59.43 ;
      RECT  96.59 132.825 96.73 129.055 ;
      RECT  98.91 132.825 99.05 129.055 ;
      RECT  102.17 132.825 102.03 129.055 ;
      RECT  99.85 132.825 99.71 129.055 ;
      RECT  102.83 132.825 102.97 129.055 ;
      RECT  105.15 132.825 105.29 129.055 ;
      RECT  108.41 132.825 108.27 129.055 ;
      RECT  106.09 132.825 105.95 129.055 ;
      RECT  109.07 132.825 109.21 129.055 ;
      RECT  111.39 132.825 111.53 129.055 ;
      RECT  114.65 132.825 114.51 129.055 ;
      RECT  112.33 132.825 112.19 129.055 ;
      RECT  115.31 132.825 115.45 129.055 ;
      RECT  117.63 132.825 117.77 129.055 ;
      RECT  120.89 132.825 120.75 129.055 ;
      RECT  118.57 132.825 118.43 129.055 ;
      RECT  121.55 132.825 121.69 129.055 ;
      RECT  123.87 132.825 124.01 129.055 ;
      RECT  127.13 132.825 126.99 129.055 ;
      RECT  124.81 132.825 124.67 129.055 ;
      RECT  127.79 132.825 127.93 129.055 ;
      RECT  130.11 132.825 130.25 129.055 ;
      RECT  133.37 132.825 133.23 129.055 ;
      RECT  131.05 132.825 130.91 129.055 ;
      RECT  134.03 132.825 134.17 129.055 ;
      RECT  136.35 132.825 136.49 129.055 ;
      RECT  139.61 132.825 139.47 129.055 ;
      RECT  137.29 132.825 137.15 129.055 ;
      RECT  140.27 132.825 140.41 129.055 ;
      RECT  142.59 132.825 142.73 129.055 ;
      RECT  145.85 132.825 145.71 129.055 ;
      RECT  143.53 132.825 143.39 129.055 ;
      RECT  146.51 132.825 146.65 129.055 ;
      RECT  148.83 132.825 148.97 129.055 ;
      RECT  96.59 132.825 96.73 129.055 ;
      RECT  98.91 132.825 99.05 129.055 ;
      RECT  102.03 132.825 102.17 129.055 ;
      RECT  99.71 132.825 99.85 129.055 ;
      RECT  102.83 132.825 102.97 129.055 ;
      RECT  105.15 132.825 105.29 129.055 ;
      RECT  108.27 132.825 108.41 129.055 ;
      RECT  105.95 132.825 106.09 129.055 ;
      RECT  109.07 132.825 109.21 129.055 ;
      RECT  111.39 132.825 111.53 129.055 ;
      RECT  114.51 132.825 114.65 129.055 ;
      RECT  112.19 132.825 112.33 129.055 ;
      RECT  115.31 132.825 115.45 129.055 ;
      RECT  117.63 132.825 117.77 129.055 ;
      RECT  120.75 132.825 120.89 129.055 ;
      RECT  118.43 132.825 118.57 129.055 ;
      RECT  121.55 132.825 121.69 129.055 ;
      RECT  123.87 132.825 124.01 129.055 ;
      RECT  126.99 132.825 127.13 129.055 ;
      RECT  124.67 132.825 124.81 129.055 ;
      RECT  127.79 132.825 127.93 129.055 ;
      RECT  130.11 132.825 130.25 129.055 ;
      RECT  133.23 132.825 133.37 129.055 ;
      RECT  130.91 132.825 131.05 129.055 ;
      RECT  134.03 132.825 134.17 129.055 ;
      RECT  136.35 132.825 136.49 129.055 ;
      RECT  139.47 132.825 139.61 129.055 ;
      RECT  137.15 132.825 137.29 129.055 ;
      RECT  140.27 132.825 140.41 129.055 ;
      RECT  142.59 132.825 142.73 129.055 ;
      RECT  145.71 132.825 145.85 129.055 ;
      RECT  143.39 132.825 143.53 129.055 ;
      RECT  146.51 132.825 146.65 129.055 ;
      RECT  148.83 132.825 148.97 129.055 ;
      RECT  97.62 139.655 97.76 134.085 ;
      RECT  97.62 139.945 97.96 139.655 ;
      RECT  97.24 139.715 97.41 134.085 ;
      RECT  98.4 135.34 98.63 134.97 ;
      RECT  96.73 134.545 97.02 134.245 ;
      RECT  97.95 139.195 98.26 138.855 ;
      RECT  98.05 143.405 98.28 143.025 ;
      RECT  98.05 145.01 98.28 144.64 ;
      RECT  96.78 145.365 97.01 144.095 ;
      RECT  97.24 145.365 97.41 139.945 ;
      RECT  97.18 139.945 97.47 139.715 ;
      RECT  97.62 145.365 97.76 139.945 ;
      RECT  100.52 139.655 100.38 134.085 ;
      RECT  100.52 139.945 100.18 139.655 ;
      RECT  100.9 139.715 100.73 134.085 ;
      RECT  99.74 135.34 99.51 134.97 ;
      RECT  101.41 134.545 101.12 134.245 ;
      RECT  100.19 139.195 99.88 138.855 ;
      RECT  100.09 143.405 99.86 143.025 ;
      RECT  100.09 145.01 99.86 144.64 ;
      RECT  101.36 145.365 101.13 144.095 ;
      RECT  100.9 145.365 100.73 139.945 ;
      RECT  100.96 139.945 100.67 139.715 ;
      RECT  100.52 145.365 100.38 139.945 ;
      RECT  103.86 139.655 104.0 134.085 ;
      RECT  103.86 139.945 104.2 139.655 ;
      RECT  103.48 139.715 103.65 134.085 ;
      RECT  104.64 135.34 104.87 134.97 ;
      RECT  102.97 134.545 103.26 134.245 ;
      RECT  104.19 139.195 104.5 138.855 ;
      RECT  104.29 143.405 104.52 143.025 ;
      RECT  104.29 145.01 104.52 144.64 ;
      RECT  103.02 145.365 103.25 144.095 ;
      RECT  103.48 145.365 103.65 139.945 ;
      RECT  103.42 139.945 103.71 139.715 ;
      RECT  103.86 145.365 104.0 139.945 ;
      RECT  106.76 139.655 106.62 134.085 ;
      RECT  106.76 139.945 106.42 139.655 ;
      RECT  107.14 139.715 106.97 134.085 ;
      RECT  105.98 135.34 105.75 134.97 ;
      RECT  107.65 134.545 107.36 134.245 ;
      RECT  106.43 139.195 106.12 138.855 ;
      RECT  106.33 143.405 106.1 143.025 ;
      RECT  106.33 145.01 106.1 144.64 ;
      RECT  107.6 145.365 107.37 144.095 ;
      RECT  107.14 145.365 106.97 139.945 ;
      RECT  107.2 139.945 106.91 139.715 ;
      RECT  106.76 145.365 106.62 139.945 ;
      RECT  110.1 139.655 110.24 134.085 ;
      RECT  110.1 139.945 110.44 139.655 ;
      RECT  109.72 139.715 109.89 134.085 ;
      RECT  110.88 135.34 111.11 134.97 ;
      RECT  109.21 134.545 109.5 134.245 ;
      RECT  110.43 139.195 110.74 138.855 ;
      RECT  110.53 143.405 110.76 143.025 ;
      RECT  110.53 145.01 110.76 144.64 ;
      RECT  109.26 145.365 109.49 144.095 ;
      RECT  109.72 145.365 109.89 139.945 ;
      RECT  109.66 139.945 109.95 139.715 ;
      RECT  110.1 145.365 110.24 139.945 ;
      RECT  113.0 139.655 112.86 134.085 ;
      RECT  113.0 139.945 112.66 139.655 ;
      RECT  113.38 139.715 113.21 134.085 ;
      RECT  112.22 135.34 111.99 134.97 ;
      RECT  113.89 134.545 113.6 134.245 ;
      RECT  112.67 139.195 112.36 138.855 ;
      RECT  112.57 143.405 112.34 143.025 ;
      RECT  112.57 145.01 112.34 144.64 ;
      RECT  113.84 145.365 113.61 144.095 ;
      RECT  113.38 145.365 113.21 139.945 ;
      RECT  113.44 139.945 113.15 139.715 ;
      RECT  113.0 145.365 112.86 139.945 ;
      RECT  116.34 139.655 116.48 134.085 ;
      RECT  116.34 139.945 116.68 139.655 ;
      RECT  115.96 139.715 116.13 134.085 ;
      RECT  117.12 135.34 117.35 134.97 ;
      RECT  115.45 134.545 115.74 134.245 ;
      RECT  116.67 139.195 116.98 138.855 ;
      RECT  116.77 143.405 117.0 143.025 ;
      RECT  116.77 145.01 117.0 144.64 ;
      RECT  115.5 145.365 115.73 144.095 ;
      RECT  115.96 145.365 116.13 139.945 ;
      RECT  115.9 139.945 116.19 139.715 ;
      RECT  116.34 145.365 116.48 139.945 ;
      RECT  119.24 139.655 119.1 134.085 ;
      RECT  119.24 139.945 118.9 139.655 ;
      RECT  119.62 139.715 119.45 134.085 ;
      RECT  118.46 135.34 118.23 134.97 ;
      RECT  120.13 134.545 119.84 134.245 ;
      RECT  118.91 139.195 118.6 138.855 ;
      RECT  118.81 143.405 118.58 143.025 ;
      RECT  118.81 145.01 118.58 144.64 ;
      RECT  120.08 145.365 119.85 144.095 ;
      RECT  119.62 145.365 119.45 139.945 ;
      RECT  119.68 139.945 119.39 139.715 ;
      RECT  119.24 145.365 119.1 139.945 ;
      RECT  122.58 139.655 122.72 134.085 ;
      RECT  122.58 139.945 122.92 139.655 ;
      RECT  122.2 139.715 122.37 134.085 ;
      RECT  123.36 135.34 123.59 134.97 ;
      RECT  121.69 134.545 121.98 134.245 ;
      RECT  122.91 139.195 123.22 138.855 ;
      RECT  123.01 143.405 123.24 143.025 ;
      RECT  123.01 145.01 123.24 144.64 ;
      RECT  121.74 145.365 121.97 144.095 ;
      RECT  122.2 145.365 122.37 139.945 ;
      RECT  122.14 139.945 122.43 139.715 ;
      RECT  122.58 145.365 122.72 139.945 ;
      RECT  125.48 139.655 125.34 134.085 ;
      RECT  125.48 139.945 125.14 139.655 ;
      RECT  125.86 139.715 125.69 134.085 ;
      RECT  124.7 135.34 124.47 134.97 ;
      RECT  126.37 134.545 126.08 134.245 ;
      RECT  125.15 139.195 124.84 138.855 ;
      RECT  125.05 143.405 124.82 143.025 ;
      RECT  125.05 145.01 124.82 144.64 ;
      RECT  126.32 145.365 126.09 144.095 ;
      RECT  125.86 145.365 125.69 139.945 ;
      RECT  125.92 139.945 125.63 139.715 ;
      RECT  125.48 145.365 125.34 139.945 ;
      RECT  128.82 139.655 128.96 134.085 ;
      RECT  128.82 139.945 129.16 139.655 ;
      RECT  128.44 139.715 128.61 134.085 ;
      RECT  129.6 135.34 129.83 134.97 ;
      RECT  127.93 134.545 128.22 134.245 ;
      RECT  129.15 139.195 129.46 138.855 ;
      RECT  129.25 143.405 129.48 143.025 ;
      RECT  129.25 145.01 129.48 144.64 ;
      RECT  127.98 145.365 128.21 144.095 ;
      RECT  128.44 145.365 128.61 139.945 ;
      RECT  128.38 139.945 128.67 139.715 ;
      RECT  128.82 145.365 128.96 139.945 ;
      RECT  131.72 139.655 131.58 134.085 ;
      RECT  131.72 139.945 131.38 139.655 ;
      RECT  132.1 139.715 131.93 134.085 ;
      RECT  130.94 135.34 130.71 134.97 ;
      RECT  132.61 134.545 132.32 134.245 ;
      RECT  131.39 139.195 131.08 138.855 ;
      RECT  131.29 143.405 131.06 143.025 ;
      RECT  131.29 145.01 131.06 144.64 ;
      RECT  132.56 145.365 132.33 144.095 ;
      RECT  132.1 145.365 131.93 139.945 ;
      RECT  132.16 139.945 131.87 139.715 ;
      RECT  131.72 145.365 131.58 139.945 ;
      RECT  135.06 139.655 135.2 134.085 ;
      RECT  135.06 139.945 135.4 139.655 ;
      RECT  134.68 139.715 134.85 134.085 ;
      RECT  135.84 135.34 136.07 134.97 ;
      RECT  134.17 134.545 134.46 134.245 ;
      RECT  135.39 139.195 135.7 138.855 ;
      RECT  135.49 143.405 135.72 143.025 ;
      RECT  135.49 145.01 135.72 144.64 ;
      RECT  134.22 145.365 134.45 144.095 ;
      RECT  134.68 145.365 134.85 139.945 ;
      RECT  134.62 139.945 134.91 139.715 ;
      RECT  135.06 145.365 135.2 139.945 ;
      RECT  137.96 139.655 137.82 134.085 ;
      RECT  137.96 139.945 137.62 139.655 ;
      RECT  138.34 139.715 138.17 134.085 ;
      RECT  137.18 135.34 136.95 134.97 ;
      RECT  138.85 134.545 138.56 134.245 ;
      RECT  137.63 139.195 137.32 138.855 ;
      RECT  137.53 143.405 137.3 143.025 ;
      RECT  137.53 145.01 137.3 144.64 ;
      RECT  138.8 145.365 138.57 144.095 ;
      RECT  138.34 145.365 138.17 139.945 ;
      RECT  138.4 139.945 138.11 139.715 ;
      RECT  137.96 145.365 137.82 139.945 ;
      RECT  141.3 139.655 141.44 134.085 ;
      RECT  141.3 139.945 141.64 139.655 ;
      RECT  140.92 139.715 141.09 134.085 ;
      RECT  142.08 135.34 142.31 134.97 ;
      RECT  140.41 134.545 140.7 134.245 ;
      RECT  141.63 139.195 141.94 138.855 ;
      RECT  141.73 143.405 141.96 143.025 ;
      RECT  141.73 145.01 141.96 144.64 ;
      RECT  140.46 145.365 140.69 144.095 ;
      RECT  140.92 145.365 141.09 139.945 ;
      RECT  140.86 139.945 141.15 139.715 ;
      RECT  141.3 145.365 141.44 139.945 ;
      RECT  144.2 139.655 144.06 134.085 ;
      RECT  144.2 139.945 143.86 139.655 ;
      RECT  144.58 139.715 144.41 134.085 ;
      RECT  143.42 135.34 143.19 134.97 ;
      RECT  145.09 134.545 144.8 134.245 ;
      RECT  143.87 139.195 143.56 138.855 ;
      RECT  143.77 143.405 143.54 143.025 ;
      RECT  143.77 145.01 143.54 144.64 ;
      RECT  145.04 145.365 144.81 144.095 ;
      RECT  144.58 145.365 144.41 139.945 ;
      RECT  144.64 139.945 144.35 139.715 ;
      RECT  144.2 145.365 144.06 139.945 ;
      RECT  96.78 145.365 97.01 144.095 ;
      RECT  97.24 139.715 97.41 134.085 ;
      RECT  97.62 139.655 97.76 134.085 ;
      RECT  101.13 145.365 101.36 144.095 ;
      RECT  100.73 139.715 100.9 134.085 ;
      RECT  100.38 139.655 100.52 134.085 ;
      RECT  103.02 145.365 103.25 144.095 ;
      RECT  103.48 139.715 103.65 134.085 ;
      RECT  103.86 139.655 104.0 134.085 ;
      RECT  107.37 145.365 107.6 144.095 ;
      RECT  106.97 139.715 107.14 134.085 ;
      RECT  106.62 139.655 106.76 134.085 ;
      RECT  109.26 145.365 109.49 144.095 ;
      RECT  109.72 139.715 109.89 134.085 ;
      RECT  110.1 139.655 110.24 134.085 ;
      RECT  113.61 145.365 113.84 144.095 ;
      RECT  113.21 139.715 113.38 134.085 ;
      RECT  112.86 139.655 113.0 134.085 ;
      RECT  115.5 145.365 115.73 144.095 ;
      RECT  115.96 139.715 116.13 134.085 ;
      RECT  116.34 139.655 116.48 134.085 ;
      RECT  119.85 145.365 120.08 144.095 ;
      RECT  119.45 139.715 119.62 134.085 ;
      RECT  119.1 139.655 119.24 134.085 ;
      RECT  121.74 145.365 121.97 144.095 ;
      RECT  122.2 139.715 122.37 134.085 ;
      RECT  122.58 139.655 122.72 134.085 ;
      RECT  126.09 145.365 126.32 144.095 ;
      RECT  125.69 139.715 125.86 134.085 ;
      RECT  125.34 139.655 125.48 134.085 ;
      RECT  127.98 145.365 128.21 144.095 ;
      RECT  128.44 139.715 128.61 134.085 ;
      RECT  128.82 139.655 128.96 134.085 ;
      RECT  132.33 145.365 132.56 144.095 ;
      RECT  131.93 139.715 132.1 134.085 ;
      RECT  131.58 139.655 131.72 134.085 ;
      RECT  134.22 145.365 134.45 144.095 ;
      RECT  134.68 139.715 134.85 134.085 ;
      RECT  135.06 139.655 135.2 134.085 ;
      RECT  138.57 145.365 138.8 144.095 ;
      RECT  138.17 139.715 138.34 134.085 ;
      RECT  137.82 139.655 137.96 134.085 ;
      RECT  140.46 145.365 140.69 144.095 ;
      RECT  140.92 139.715 141.09 134.085 ;
      RECT  141.3 139.655 141.44 134.085 ;
      RECT  144.81 145.365 145.04 144.095 ;
      RECT  144.41 139.715 144.58 134.085 ;
      RECT  144.06 139.655 144.2 134.085 ;
      RECT  146.51 129.055 146.65 132.825 ;
      RECT  148.83 129.055 148.97 132.825 ;
      RECT  96.78 144.095 97.01 145.365 ;
      RECT  101.13 144.095 101.36 145.365 ;
      RECT  103.02 144.095 103.25 145.365 ;
      RECT  107.37 144.095 107.6 145.365 ;
      RECT  109.26 144.095 109.49 145.365 ;
      RECT  113.61 144.095 113.84 145.365 ;
      RECT  115.5 144.095 115.73 145.365 ;
      RECT  119.85 144.095 120.08 145.365 ;
      RECT  121.74 144.095 121.97 145.365 ;
      RECT  126.09 144.095 126.32 145.365 ;
      RECT  127.98 144.095 128.21 145.365 ;
      RECT  132.33 144.095 132.56 145.365 ;
      RECT  134.22 144.095 134.45 145.365 ;
      RECT  138.57 144.095 138.8 145.365 ;
      RECT  140.46 144.095 140.69 145.365 ;
      RECT  144.81 144.095 145.04 145.365 ;
      RECT  46.7 92.39 46.84 94.365 ;
      RECT  45.34 92.39 45.48 94.365 ;
      RECT  46.7 96.34 46.84 94.365 ;
      RECT  45.34 96.34 45.48 94.365 ;
      RECT  53.26 92.23 53.51 94.4 ;
      RECT  51.14 92.24 51.38 94.4 ;
      RECT  56.57 92.39 56.71 94.365 ;
      RECT  55.21 92.39 55.35 94.365 ;
      RECT  56.57 92.39 56.71 94.365 ;
      RECT  53.26 92.23 53.51 94.4 ;
      RECT  55.21 92.39 55.35 94.365 ;
      RECT  51.14 92.24 51.38 94.4 ;
      RECT  53.26 96.5 53.51 94.33 ;
      RECT  51.14 96.49 51.38 94.33 ;
      RECT  56.57 96.34 56.71 94.365 ;
      RECT  55.21 96.34 55.35 94.365 ;
      RECT  56.57 96.34 56.71 94.365 ;
      RECT  53.26 96.5 53.51 94.33 ;
      RECT  55.21 96.34 55.35 94.365 ;
      RECT  51.14 96.49 51.38 94.33 ;
      RECT  53.26 96.18 53.51 98.35 ;
      RECT  51.14 96.19 51.38 98.35 ;
      RECT  56.57 96.34 56.71 98.315 ;
      RECT  55.21 96.34 55.35 98.315 ;
      RECT  56.57 96.34 56.71 98.315 ;
      RECT  53.26 96.18 53.51 98.35 ;
      RECT  55.21 96.34 55.35 98.315 ;
      RECT  51.14 96.19 51.38 98.35 ;
      RECT  53.26 100.45 53.51 98.28 ;
      RECT  51.14 100.44 51.38 98.28 ;
      RECT  56.57 100.29 56.71 98.315 ;
      RECT  55.21 100.29 55.35 98.315 ;
      RECT  56.57 100.29 56.71 98.315 ;
      RECT  53.26 100.45 53.51 98.28 ;
      RECT  55.21 100.29 55.35 98.315 ;
      RECT  51.14 100.44 51.38 98.28 ;
      RECT  43.16 93.215 43.42 93.535 ;
      RECT  43.56 95.195 43.82 95.515 ;
      RECT  46.7 104.24 46.84 106.215 ;
      RECT  45.34 104.24 45.48 106.215 ;
      RECT  46.7 108.19 46.84 106.215 ;
      RECT  45.34 108.19 45.48 106.215 ;
      RECT  53.26 104.08 53.51 106.25 ;
      RECT  51.14 104.09 51.38 106.25 ;
      RECT  56.57 104.24 56.71 106.215 ;
      RECT  55.21 104.24 55.35 106.215 ;
      RECT  56.57 104.24 56.71 106.215 ;
      RECT  53.26 104.08 53.51 106.25 ;
      RECT  55.21 104.24 55.35 106.215 ;
      RECT  51.14 104.09 51.38 106.25 ;
      RECT  53.26 108.35 53.51 106.18 ;
      RECT  51.14 108.34 51.38 106.18 ;
      RECT  56.57 108.19 56.71 106.215 ;
      RECT  55.21 108.19 55.35 106.215 ;
      RECT  56.57 108.19 56.71 106.215 ;
      RECT  53.26 108.35 53.51 106.18 ;
      RECT  55.21 108.19 55.35 106.215 ;
      RECT  51.14 108.34 51.38 106.18 ;
      RECT  53.26 108.03 53.51 110.2 ;
      RECT  51.14 108.04 51.38 110.2 ;
      RECT  56.57 108.19 56.71 110.165 ;
      RECT  55.21 108.19 55.35 110.165 ;
      RECT  56.57 108.19 56.71 110.165 ;
      RECT  53.26 108.03 53.51 110.2 ;
      RECT  55.21 108.19 55.35 110.165 ;
      RECT  51.14 108.04 51.38 110.2 ;
      RECT  53.26 112.3 53.51 110.13 ;
      RECT  51.14 112.29 51.38 110.13 ;
      RECT  56.57 112.14 56.71 110.165 ;
      RECT  55.21 112.14 55.35 110.165 ;
      RECT  56.57 112.14 56.71 110.165 ;
      RECT  53.26 112.3 53.51 110.13 ;
      RECT  55.21 112.14 55.35 110.165 ;
      RECT  51.14 112.29 51.38 110.13 ;
      RECT  43.16 105.065 43.42 105.385 ;
      RECT  43.56 107.045 43.82 107.365 ;
      RECT  64.33 92.23 64.58 94.4 ;
      RECT  62.21 92.24 62.45 94.4 ;
      RECT  67.64 92.39 67.78 94.365 ;
      RECT  66.28 92.39 66.42 94.365 ;
      RECT  67.64 92.39 67.78 94.365 ;
      RECT  64.33 92.23 64.58 94.4 ;
      RECT  66.28 92.39 66.42 94.365 ;
      RECT  62.21 92.24 62.45 94.4 ;
      RECT  64.33 96.5 64.58 94.33 ;
      RECT  62.21 96.49 62.45 94.33 ;
      RECT  67.64 96.34 67.78 94.365 ;
      RECT  66.28 96.34 66.42 94.365 ;
      RECT  67.64 96.34 67.78 94.365 ;
      RECT  64.33 96.5 64.58 94.33 ;
      RECT  66.28 96.34 66.42 94.365 ;
      RECT  62.21 96.49 62.45 94.33 ;
      RECT  64.33 96.18 64.58 98.35 ;
      RECT  62.21 96.19 62.45 98.35 ;
      RECT  67.64 96.34 67.78 98.315 ;
      RECT  66.28 96.34 66.42 98.315 ;
      RECT  67.64 96.34 67.78 98.315 ;
      RECT  64.33 96.18 64.58 98.35 ;
      RECT  66.28 96.34 66.42 98.315 ;
      RECT  62.21 96.19 62.45 98.35 ;
      RECT  64.33 100.45 64.58 98.28 ;
      RECT  62.21 100.44 62.45 98.28 ;
      RECT  67.64 100.29 67.78 98.315 ;
      RECT  66.28 100.29 66.42 98.315 ;
      RECT  67.64 100.29 67.78 98.315 ;
      RECT  64.33 100.45 64.58 98.28 ;
      RECT  66.28 100.29 66.42 98.315 ;
      RECT  62.21 100.44 62.45 98.28 ;
      RECT  64.33 100.13 64.58 102.3 ;
      RECT  62.21 100.14 62.45 102.3 ;
      RECT  67.64 100.29 67.78 102.265 ;
      RECT  66.28 100.29 66.42 102.265 ;
      RECT  67.64 100.29 67.78 102.265 ;
      RECT  64.33 100.13 64.58 102.3 ;
      RECT  66.28 100.29 66.42 102.265 ;
      RECT  62.21 100.14 62.45 102.3 ;
      RECT  64.33 104.4 64.58 102.23 ;
      RECT  62.21 104.39 62.45 102.23 ;
      RECT  67.64 104.24 67.78 102.265 ;
      RECT  66.28 104.24 66.42 102.265 ;
      RECT  67.64 104.24 67.78 102.265 ;
      RECT  64.33 104.4 64.58 102.23 ;
      RECT  66.28 104.24 66.42 102.265 ;
      RECT  62.21 104.39 62.45 102.23 ;
      RECT  64.33 104.08 64.58 106.25 ;
      RECT  62.21 104.09 62.45 106.25 ;
      RECT  67.64 104.24 67.78 106.215 ;
      RECT  66.28 104.24 66.42 106.215 ;
      RECT  67.64 104.24 67.78 106.215 ;
      RECT  64.33 104.08 64.58 106.25 ;
      RECT  66.28 104.24 66.42 106.215 ;
      RECT  62.21 104.09 62.45 106.25 ;
      RECT  64.33 108.35 64.58 106.18 ;
      RECT  62.21 108.34 62.45 106.18 ;
      RECT  67.64 108.19 67.78 106.215 ;
      RECT  66.28 108.19 66.42 106.215 ;
      RECT  67.64 108.19 67.78 106.215 ;
      RECT  64.33 108.35 64.58 106.18 ;
      RECT  66.28 108.19 66.42 106.215 ;
      RECT  62.21 108.34 62.45 106.18 ;
      RECT  64.33 108.03 64.58 110.2 ;
      RECT  62.21 108.04 62.45 110.2 ;
      RECT  67.64 108.19 67.78 110.165 ;
      RECT  66.28 108.19 66.42 110.165 ;
      RECT  67.64 108.19 67.78 110.165 ;
      RECT  64.33 108.03 64.58 110.2 ;
      RECT  66.28 108.19 66.42 110.165 ;
      RECT  62.21 108.04 62.45 110.2 ;
      RECT  64.33 112.3 64.58 110.13 ;
      RECT  62.21 112.29 62.45 110.13 ;
      RECT  67.64 112.14 67.78 110.165 ;
      RECT  66.28 112.14 66.42 110.165 ;
      RECT  67.64 112.14 67.78 110.165 ;
      RECT  64.33 112.3 64.58 110.13 ;
      RECT  66.28 112.14 66.42 110.165 ;
      RECT  62.21 112.29 62.45 110.13 ;
      RECT  64.33 111.98 64.58 114.15 ;
      RECT  62.21 111.99 62.45 114.15 ;
      RECT  67.64 112.14 67.78 114.115 ;
      RECT  66.28 112.14 66.42 114.115 ;
      RECT  67.64 112.14 67.78 114.115 ;
      RECT  64.33 111.98 64.58 114.15 ;
      RECT  66.28 112.14 66.42 114.115 ;
      RECT  62.21 111.99 62.45 114.15 ;
      RECT  64.33 116.25 64.58 114.08 ;
      RECT  62.21 116.24 62.45 114.08 ;
      RECT  67.64 116.09 67.78 114.115 ;
      RECT  66.28 116.09 66.42 114.115 ;
      RECT  67.64 116.09 67.78 114.115 ;
      RECT  64.33 116.25 64.58 114.08 ;
      RECT  66.28 116.09 66.42 114.115 ;
      RECT  62.21 116.24 62.45 114.08 ;
      RECT  64.33 115.93 64.58 118.1 ;
      RECT  62.21 115.94 62.45 118.1 ;
      RECT  67.64 116.09 67.78 118.065 ;
      RECT  66.28 116.09 66.42 118.065 ;
      RECT  67.64 116.09 67.78 118.065 ;
      RECT  64.33 115.93 64.58 118.1 ;
      RECT  66.28 116.09 66.42 118.065 ;
      RECT  62.21 115.94 62.45 118.1 ;
      RECT  64.33 120.2 64.58 118.03 ;
      RECT  62.21 120.19 62.45 118.03 ;
      RECT  67.64 120.04 67.78 118.065 ;
      RECT  66.28 120.04 66.42 118.065 ;
      RECT  67.64 120.04 67.78 118.065 ;
      RECT  64.33 120.2 64.58 118.03 ;
      RECT  66.28 120.04 66.42 118.065 ;
      RECT  62.21 120.19 62.45 118.03 ;
      RECT  64.33 119.88 64.58 122.05 ;
      RECT  62.21 119.89 62.45 122.05 ;
      RECT  67.64 120.04 67.78 122.015 ;
      RECT  66.28 120.04 66.42 122.015 ;
      RECT  67.64 120.04 67.78 122.015 ;
      RECT  64.33 119.88 64.58 122.05 ;
      RECT  66.28 120.04 66.42 122.015 ;
      RECT  62.21 119.89 62.45 122.05 ;
      RECT  64.33 124.15 64.58 121.98 ;
      RECT  62.21 124.14 62.45 121.98 ;
      RECT  67.64 123.99 67.78 122.015 ;
      RECT  66.28 123.99 66.42 122.015 ;
      RECT  67.64 123.99 67.78 122.015 ;
      RECT  64.33 124.15 64.58 121.98 ;
      RECT  66.28 123.99 66.42 122.015 ;
      RECT  62.21 124.14 62.45 121.98 ;
      RECT  41.08 92.39 41.22 112.14 ;
      RECT  41.48 92.39 41.62 112.14 ;
      RECT  41.88 92.39 42.02 112.14 ;
      RECT  42.28 92.39 42.42 112.14 ;
      RECT  71.94 92.085 72.19 94.255 ;
      RECT  69.82 92.095 70.06 94.255 ;
      RECT  84.83 92.245 84.97 94.22 ;
      RECT  77.21 92.245 77.35 94.22 ;
      RECT  84.83 92.245 84.97 94.22 ;
      RECT  71.94 92.085 72.19 94.255 ;
      RECT  77.21 92.245 77.35 94.22 ;
      RECT  69.82 92.095 70.06 94.255 ;
      RECT  71.94 96.355 72.19 94.185 ;
      RECT  69.82 96.345 70.06 94.185 ;
      RECT  84.83 96.195 84.97 94.22 ;
      RECT  77.21 96.195 77.35 94.22 ;
      RECT  84.83 96.195 84.97 94.22 ;
      RECT  71.94 96.355 72.19 94.185 ;
      RECT  77.21 96.195 77.35 94.22 ;
      RECT  69.82 96.345 70.06 94.185 ;
      RECT  71.94 96.035 72.19 98.205 ;
      RECT  69.82 96.045 70.06 98.205 ;
      RECT  84.83 96.195 84.97 98.17 ;
      RECT  77.21 96.195 77.35 98.17 ;
      RECT  84.83 96.195 84.97 98.17 ;
      RECT  71.94 96.035 72.19 98.205 ;
      RECT  77.21 96.195 77.35 98.17 ;
      RECT  69.82 96.045 70.06 98.205 ;
      RECT  71.94 100.305 72.19 98.135 ;
      RECT  69.82 100.295 70.06 98.135 ;
      RECT  84.83 100.145 84.97 98.17 ;
      RECT  77.21 100.145 77.35 98.17 ;
      RECT  84.83 100.145 84.97 98.17 ;
      RECT  71.94 100.305 72.19 98.135 ;
      RECT  77.21 100.145 77.35 98.17 ;
      RECT  69.82 100.295 70.06 98.135 ;
      RECT  71.94 99.985 72.19 102.155 ;
      RECT  69.82 99.995 70.06 102.155 ;
      RECT  84.83 100.145 84.97 102.12 ;
      RECT  77.21 100.145 77.35 102.12 ;
      RECT  84.83 100.145 84.97 102.12 ;
      RECT  71.94 99.985 72.19 102.155 ;
      RECT  77.21 100.145 77.35 102.12 ;
      RECT  69.82 99.995 70.06 102.155 ;
      RECT  71.94 104.255 72.19 102.085 ;
      RECT  69.82 104.245 70.06 102.085 ;
      RECT  84.83 104.095 84.97 102.12 ;
      RECT  77.21 104.095 77.35 102.12 ;
      RECT  84.83 104.095 84.97 102.12 ;
      RECT  71.94 104.255 72.19 102.085 ;
      RECT  77.21 104.095 77.35 102.12 ;
      RECT  69.82 104.245 70.06 102.085 ;
      RECT  71.94 103.935 72.19 106.105 ;
      RECT  69.82 103.945 70.06 106.105 ;
      RECT  84.83 104.095 84.97 106.07 ;
      RECT  77.21 104.095 77.35 106.07 ;
      RECT  84.83 104.095 84.97 106.07 ;
      RECT  71.94 103.935 72.19 106.105 ;
      RECT  77.21 104.095 77.35 106.07 ;
      RECT  69.82 103.945 70.06 106.105 ;
      RECT  71.94 108.205 72.19 106.035 ;
      RECT  69.82 108.195 70.06 106.035 ;
      RECT  84.83 108.045 84.97 106.07 ;
      RECT  77.21 108.045 77.35 106.07 ;
      RECT  84.83 108.045 84.97 106.07 ;
      RECT  71.94 108.205 72.19 106.035 ;
      RECT  77.21 108.045 77.35 106.07 ;
      RECT  69.82 108.195 70.06 106.035 ;
      RECT  71.94 107.885 72.19 110.055 ;
      RECT  69.82 107.895 70.06 110.055 ;
      RECT  84.83 108.045 84.97 110.02 ;
      RECT  77.21 108.045 77.35 110.02 ;
      RECT  84.83 108.045 84.97 110.02 ;
      RECT  71.94 107.885 72.19 110.055 ;
      RECT  77.21 108.045 77.35 110.02 ;
      RECT  69.82 107.895 70.06 110.055 ;
      RECT  71.94 112.155 72.19 109.985 ;
      RECT  69.82 112.145 70.06 109.985 ;
      RECT  84.83 111.995 84.97 110.02 ;
      RECT  77.21 111.995 77.35 110.02 ;
      RECT  84.83 111.995 84.97 110.02 ;
      RECT  71.94 112.155 72.19 109.985 ;
      RECT  77.21 111.995 77.35 110.02 ;
      RECT  69.82 112.145 70.06 109.985 ;
      RECT  71.94 111.835 72.19 114.005 ;
      RECT  69.82 111.845 70.06 114.005 ;
      RECT  84.83 111.995 84.97 113.97 ;
      RECT  77.21 111.995 77.35 113.97 ;
      RECT  84.83 111.995 84.97 113.97 ;
      RECT  71.94 111.835 72.19 114.005 ;
      RECT  77.21 111.995 77.35 113.97 ;
      RECT  69.82 111.845 70.06 114.005 ;
      RECT  71.94 116.105 72.19 113.935 ;
      RECT  69.82 116.095 70.06 113.935 ;
      RECT  84.83 115.945 84.97 113.97 ;
      RECT  77.21 115.945 77.35 113.97 ;
      RECT  84.83 115.945 84.97 113.97 ;
      RECT  71.94 116.105 72.19 113.935 ;
      RECT  77.21 115.945 77.35 113.97 ;
      RECT  69.82 116.095 70.06 113.935 ;
      RECT  71.94 115.785 72.19 117.955 ;
      RECT  69.82 115.795 70.06 117.955 ;
      RECT  84.83 115.945 84.97 117.92 ;
      RECT  77.21 115.945 77.35 117.92 ;
      RECT  84.83 115.945 84.97 117.92 ;
      RECT  71.94 115.785 72.19 117.955 ;
      RECT  77.21 115.945 77.35 117.92 ;
      RECT  69.82 115.795 70.06 117.955 ;
      RECT  71.94 120.055 72.19 117.885 ;
      RECT  69.82 120.045 70.06 117.885 ;
      RECT  84.83 119.895 84.97 117.92 ;
      RECT  77.21 119.895 77.35 117.92 ;
      RECT  84.83 119.895 84.97 117.92 ;
      RECT  71.94 120.055 72.19 117.885 ;
      RECT  77.21 119.895 77.35 117.92 ;
      RECT  69.82 120.045 70.06 117.885 ;
      RECT  71.94 119.735 72.19 121.905 ;
      RECT  69.82 119.745 70.06 121.905 ;
      RECT  84.83 119.895 84.97 121.87 ;
      RECT  77.21 119.895 77.35 121.87 ;
      RECT  84.83 119.895 84.97 121.87 ;
      RECT  71.94 119.735 72.19 121.905 ;
      RECT  77.21 119.895 77.35 121.87 ;
      RECT  69.82 119.745 70.06 121.905 ;
      RECT  71.94 124.005 72.19 121.835 ;
      RECT  69.82 123.995 70.06 121.835 ;
      RECT  84.83 123.845 84.97 121.87 ;
      RECT  77.21 123.845 77.35 121.87 ;
      RECT  84.83 123.845 84.97 121.87 ;
      RECT  71.94 124.005 72.19 121.835 ;
      RECT  77.21 123.845 77.35 121.87 ;
      RECT  69.82 123.995 70.06 121.835 ;
      RECT  71.995 92.085 72.135 123.845 ;
      RECT  84.83 92.245 84.97 123.845 ;
      RECT  77.21 92.245 77.35 123.845 ;
      RECT  69.87 92.095 70.01 123.845 ;
      RECT  41.08 92.39 41.22 112.14 ;
      RECT  41.48 92.39 41.62 112.14 ;
      RECT  41.88 92.39 42.02 112.14 ;
      RECT  42.28 92.39 42.42 112.14 ;
      RECT  195.74 92.39 195.6 94.365 ;
      RECT  197.1 92.39 196.96 94.365 ;
      RECT  195.74 96.34 195.6 94.365 ;
      RECT  197.1 96.34 196.96 94.365 ;
      RECT  189.18 92.23 188.93 94.4 ;
      RECT  191.3 92.24 191.06 94.4 ;
      RECT  185.87 92.39 185.73 94.365 ;
      RECT  187.23 92.39 187.09 94.365 ;
      RECT  185.87 92.39 185.73 94.365 ;
      RECT  189.18 92.23 188.93 94.4 ;
      RECT  187.23 92.39 187.09 94.365 ;
      RECT  191.3 92.24 191.06 94.4 ;
      RECT  189.18 96.5 188.93 94.33 ;
      RECT  191.3 96.49 191.06 94.33 ;
      RECT  185.87 96.34 185.73 94.365 ;
      RECT  187.23 96.34 187.09 94.365 ;
      RECT  185.87 96.34 185.73 94.365 ;
      RECT  189.18 96.5 188.93 94.33 ;
      RECT  187.23 96.34 187.09 94.365 ;
      RECT  191.3 96.49 191.06 94.33 ;
      RECT  189.18 96.18 188.93 98.35 ;
      RECT  191.3 96.19 191.06 98.35 ;
      RECT  185.87 96.34 185.73 98.315 ;
      RECT  187.23 96.34 187.09 98.315 ;
      RECT  185.87 96.34 185.73 98.315 ;
      RECT  189.18 96.18 188.93 98.35 ;
      RECT  187.23 96.34 187.09 98.315 ;
      RECT  191.3 96.19 191.06 98.35 ;
      RECT  189.18 100.45 188.93 98.28 ;
      RECT  191.3 100.44 191.06 98.28 ;
      RECT  185.87 100.29 185.73 98.315 ;
      RECT  187.23 100.29 187.09 98.315 ;
      RECT  185.87 100.29 185.73 98.315 ;
      RECT  189.18 100.45 188.93 98.28 ;
      RECT  187.23 100.29 187.09 98.315 ;
      RECT  191.3 100.44 191.06 98.28 ;
      RECT  199.28 93.215 199.02 93.535 ;
      RECT  198.88 95.195 198.62 95.515 ;
      RECT  195.74 104.24 195.6 106.215 ;
      RECT  197.1 104.24 196.96 106.215 ;
      RECT  195.74 108.19 195.6 106.215 ;
      RECT  197.1 108.19 196.96 106.215 ;
      RECT  189.18 104.08 188.93 106.25 ;
      RECT  191.3 104.09 191.06 106.25 ;
      RECT  185.87 104.24 185.73 106.215 ;
      RECT  187.23 104.24 187.09 106.215 ;
      RECT  185.87 104.24 185.73 106.215 ;
      RECT  189.18 104.08 188.93 106.25 ;
      RECT  187.23 104.24 187.09 106.215 ;
      RECT  191.3 104.09 191.06 106.25 ;
      RECT  189.18 108.35 188.93 106.18 ;
      RECT  191.3 108.34 191.06 106.18 ;
      RECT  185.87 108.19 185.73 106.215 ;
      RECT  187.23 108.19 187.09 106.215 ;
      RECT  185.87 108.19 185.73 106.215 ;
      RECT  189.18 108.35 188.93 106.18 ;
      RECT  187.23 108.19 187.09 106.215 ;
      RECT  191.3 108.34 191.06 106.18 ;
      RECT  189.18 108.03 188.93 110.2 ;
      RECT  191.3 108.04 191.06 110.2 ;
      RECT  185.87 108.19 185.73 110.165 ;
      RECT  187.23 108.19 187.09 110.165 ;
      RECT  185.87 108.19 185.73 110.165 ;
      RECT  189.18 108.03 188.93 110.2 ;
      RECT  187.23 108.19 187.09 110.165 ;
      RECT  191.3 108.04 191.06 110.2 ;
      RECT  189.18 112.3 188.93 110.13 ;
      RECT  191.3 112.29 191.06 110.13 ;
      RECT  185.87 112.14 185.73 110.165 ;
      RECT  187.23 112.14 187.09 110.165 ;
      RECT  185.87 112.14 185.73 110.165 ;
      RECT  189.18 112.3 188.93 110.13 ;
      RECT  187.23 112.14 187.09 110.165 ;
      RECT  191.3 112.29 191.06 110.13 ;
      RECT  199.28 105.065 199.02 105.385 ;
      RECT  198.88 107.045 198.62 107.365 ;
      RECT  178.11 92.23 177.86 94.4 ;
      RECT  180.23 92.24 179.99 94.4 ;
      RECT  174.8 92.39 174.66 94.365 ;
      RECT  176.16 92.39 176.02 94.365 ;
      RECT  174.8 92.39 174.66 94.365 ;
      RECT  178.11 92.23 177.86 94.4 ;
      RECT  176.16 92.39 176.02 94.365 ;
      RECT  180.23 92.24 179.99 94.4 ;
      RECT  178.11 96.5 177.86 94.33 ;
      RECT  180.23 96.49 179.99 94.33 ;
      RECT  174.8 96.34 174.66 94.365 ;
      RECT  176.16 96.34 176.02 94.365 ;
      RECT  174.8 96.34 174.66 94.365 ;
      RECT  178.11 96.5 177.86 94.33 ;
      RECT  176.16 96.34 176.02 94.365 ;
      RECT  180.23 96.49 179.99 94.33 ;
      RECT  178.11 96.18 177.86 98.35 ;
      RECT  180.23 96.19 179.99 98.35 ;
      RECT  174.8 96.34 174.66 98.315 ;
      RECT  176.16 96.34 176.02 98.315 ;
      RECT  174.8 96.34 174.66 98.315 ;
      RECT  178.11 96.18 177.86 98.35 ;
      RECT  176.16 96.34 176.02 98.315 ;
      RECT  180.23 96.19 179.99 98.35 ;
      RECT  178.11 100.45 177.86 98.28 ;
      RECT  180.23 100.44 179.99 98.28 ;
      RECT  174.8 100.29 174.66 98.315 ;
      RECT  176.16 100.29 176.02 98.315 ;
      RECT  174.8 100.29 174.66 98.315 ;
      RECT  178.11 100.45 177.86 98.28 ;
      RECT  176.16 100.29 176.02 98.315 ;
      RECT  180.23 100.44 179.99 98.28 ;
      RECT  178.11 100.13 177.86 102.3 ;
      RECT  180.23 100.14 179.99 102.3 ;
      RECT  174.8 100.29 174.66 102.265 ;
      RECT  176.16 100.29 176.02 102.265 ;
      RECT  174.8 100.29 174.66 102.265 ;
      RECT  178.11 100.13 177.86 102.3 ;
      RECT  176.16 100.29 176.02 102.265 ;
      RECT  180.23 100.14 179.99 102.3 ;
      RECT  178.11 104.4 177.86 102.23 ;
      RECT  180.23 104.39 179.99 102.23 ;
      RECT  174.8 104.24 174.66 102.265 ;
      RECT  176.16 104.24 176.02 102.265 ;
      RECT  174.8 104.24 174.66 102.265 ;
      RECT  178.11 104.4 177.86 102.23 ;
      RECT  176.16 104.24 176.02 102.265 ;
      RECT  180.23 104.39 179.99 102.23 ;
      RECT  178.11 104.08 177.86 106.25 ;
      RECT  180.23 104.09 179.99 106.25 ;
      RECT  174.8 104.24 174.66 106.215 ;
      RECT  176.16 104.24 176.02 106.215 ;
      RECT  174.8 104.24 174.66 106.215 ;
      RECT  178.11 104.08 177.86 106.25 ;
      RECT  176.16 104.24 176.02 106.215 ;
      RECT  180.23 104.09 179.99 106.25 ;
      RECT  178.11 108.35 177.86 106.18 ;
      RECT  180.23 108.34 179.99 106.18 ;
      RECT  174.8 108.19 174.66 106.215 ;
      RECT  176.16 108.19 176.02 106.215 ;
      RECT  174.8 108.19 174.66 106.215 ;
      RECT  178.11 108.35 177.86 106.18 ;
      RECT  176.16 108.19 176.02 106.215 ;
      RECT  180.23 108.34 179.99 106.18 ;
      RECT  178.11 108.03 177.86 110.2 ;
      RECT  180.23 108.04 179.99 110.2 ;
      RECT  174.8 108.19 174.66 110.165 ;
      RECT  176.16 108.19 176.02 110.165 ;
      RECT  174.8 108.19 174.66 110.165 ;
      RECT  178.11 108.03 177.86 110.2 ;
      RECT  176.16 108.19 176.02 110.165 ;
      RECT  180.23 108.04 179.99 110.2 ;
      RECT  178.11 112.3 177.86 110.13 ;
      RECT  180.23 112.29 179.99 110.13 ;
      RECT  174.8 112.14 174.66 110.165 ;
      RECT  176.16 112.14 176.02 110.165 ;
      RECT  174.8 112.14 174.66 110.165 ;
      RECT  178.11 112.3 177.86 110.13 ;
      RECT  176.16 112.14 176.02 110.165 ;
      RECT  180.23 112.29 179.99 110.13 ;
      RECT  178.11 111.98 177.86 114.15 ;
      RECT  180.23 111.99 179.99 114.15 ;
      RECT  174.8 112.14 174.66 114.115 ;
      RECT  176.16 112.14 176.02 114.115 ;
      RECT  174.8 112.14 174.66 114.115 ;
      RECT  178.11 111.98 177.86 114.15 ;
      RECT  176.16 112.14 176.02 114.115 ;
      RECT  180.23 111.99 179.99 114.15 ;
      RECT  178.11 116.25 177.86 114.08 ;
      RECT  180.23 116.24 179.99 114.08 ;
      RECT  174.8 116.09 174.66 114.115 ;
      RECT  176.16 116.09 176.02 114.115 ;
      RECT  174.8 116.09 174.66 114.115 ;
      RECT  178.11 116.25 177.86 114.08 ;
      RECT  176.16 116.09 176.02 114.115 ;
      RECT  180.23 116.24 179.99 114.08 ;
      RECT  178.11 115.93 177.86 118.1 ;
      RECT  180.23 115.94 179.99 118.1 ;
      RECT  174.8 116.09 174.66 118.065 ;
      RECT  176.16 116.09 176.02 118.065 ;
      RECT  174.8 116.09 174.66 118.065 ;
      RECT  178.11 115.93 177.86 118.1 ;
      RECT  176.16 116.09 176.02 118.065 ;
      RECT  180.23 115.94 179.99 118.1 ;
      RECT  178.11 120.2 177.86 118.03 ;
      RECT  180.23 120.19 179.99 118.03 ;
      RECT  174.8 120.04 174.66 118.065 ;
      RECT  176.16 120.04 176.02 118.065 ;
      RECT  174.8 120.04 174.66 118.065 ;
      RECT  178.11 120.2 177.86 118.03 ;
      RECT  176.16 120.04 176.02 118.065 ;
      RECT  180.23 120.19 179.99 118.03 ;
      RECT  178.11 119.88 177.86 122.05 ;
      RECT  180.23 119.89 179.99 122.05 ;
      RECT  174.8 120.04 174.66 122.015 ;
      RECT  176.16 120.04 176.02 122.015 ;
      RECT  174.8 120.04 174.66 122.015 ;
      RECT  178.11 119.88 177.86 122.05 ;
      RECT  176.16 120.04 176.02 122.015 ;
      RECT  180.23 119.89 179.99 122.05 ;
      RECT  178.11 124.15 177.86 121.98 ;
      RECT  180.23 124.14 179.99 121.98 ;
      RECT  174.8 123.99 174.66 122.015 ;
      RECT  176.16 123.99 176.02 122.015 ;
      RECT  174.8 123.99 174.66 122.015 ;
      RECT  178.11 124.15 177.86 121.98 ;
      RECT  176.16 123.99 176.02 122.015 ;
      RECT  180.23 124.14 179.99 121.98 ;
      RECT  201.36 92.39 201.22 112.14 ;
      RECT  200.96 92.39 200.82 112.14 ;
      RECT  200.56 92.39 200.42 112.14 ;
      RECT  200.16 92.39 200.02 112.14 ;
      RECT  170.5 92.085 170.25 94.255 ;
      RECT  172.62 92.095 172.38 94.255 ;
      RECT  157.61 92.245 157.47 94.22 ;
      RECT  165.23 92.245 165.09 94.22 ;
      RECT  157.61 92.245 157.47 94.22 ;
      RECT  170.5 92.085 170.25 94.255 ;
      RECT  165.23 92.245 165.09 94.22 ;
      RECT  172.62 92.095 172.38 94.255 ;
      RECT  170.5 96.355 170.25 94.185 ;
      RECT  172.62 96.345 172.38 94.185 ;
      RECT  157.61 96.195 157.47 94.22 ;
      RECT  165.23 96.195 165.09 94.22 ;
      RECT  157.61 96.195 157.47 94.22 ;
      RECT  170.5 96.355 170.25 94.185 ;
      RECT  165.23 96.195 165.09 94.22 ;
      RECT  172.62 96.345 172.38 94.185 ;
      RECT  170.5 96.035 170.25 98.205 ;
      RECT  172.62 96.045 172.38 98.205 ;
      RECT  157.61 96.195 157.47 98.17 ;
      RECT  165.23 96.195 165.09 98.17 ;
      RECT  157.61 96.195 157.47 98.17 ;
      RECT  170.5 96.035 170.25 98.205 ;
      RECT  165.23 96.195 165.09 98.17 ;
      RECT  172.62 96.045 172.38 98.205 ;
      RECT  170.5 100.305 170.25 98.135 ;
      RECT  172.62 100.295 172.38 98.135 ;
      RECT  157.61 100.145 157.47 98.17 ;
      RECT  165.23 100.145 165.09 98.17 ;
      RECT  157.61 100.145 157.47 98.17 ;
      RECT  170.5 100.305 170.25 98.135 ;
      RECT  165.23 100.145 165.09 98.17 ;
      RECT  172.62 100.295 172.38 98.135 ;
      RECT  170.5 99.985 170.25 102.155 ;
      RECT  172.62 99.995 172.38 102.155 ;
      RECT  157.61 100.145 157.47 102.12 ;
      RECT  165.23 100.145 165.09 102.12 ;
      RECT  157.61 100.145 157.47 102.12 ;
      RECT  170.5 99.985 170.25 102.155 ;
      RECT  165.23 100.145 165.09 102.12 ;
      RECT  172.62 99.995 172.38 102.155 ;
      RECT  170.5 104.255 170.25 102.085 ;
      RECT  172.62 104.245 172.38 102.085 ;
      RECT  157.61 104.095 157.47 102.12 ;
      RECT  165.23 104.095 165.09 102.12 ;
      RECT  157.61 104.095 157.47 102.12 ;
      RECT  170.5 104.255 170.25 102.085 ;
      RECT  165.23 104.095 165.09 102.12 ;
      RECT  172.62 104.245 172.38 102.085 ;
      RECT  170.5 103.935 170.25 106.105 ;
      RECT  172.62 103.945 172.38 106.105 ;
      RECT  157.61 104.095 157.47 106.07 ;
      RECT  165.23 104.095 165.09 106.07 ;
      RECT  157.61 104.095 157.47 106.07 ;
      RECT  170.5 103.935 170.25 106.105 ;
      RECT  165.23 104.095 165.09 106.07 ;
      RECT  172.62 103.945 172.38 106.105 ;
      RECT  170.5 108.205 170.25 106.035 ;
      RECT  172.62 108.195 172.38 106.035 ;
      RECT  157.61 108.045 157.47 106.07 ;
      RECT  165.23 108.045 165.09 106.07 ;
      RECT  157.61 108.045 157.47 106.07 ;
      RECT  170.5 108.205 170.25 106.035 ;
      RECT  165.23 108.045 165.09 106.07 ;
      RECT  172.62 108.195 172.38 106.035 ;
      RECT  170.5 107.885 170.25 110.055 ;
      RECT  172.62 107.895 172.38 110.055 ;
      RECT  157.61 108.045 157.47 110.02 ;
      RECT  165.23 108.045 165.09 110.02 ;
      RECT  157.61 108.045 157.47 110.02 ;
      RECT  170.5 107.885 170.25 110.055 ;
      RECT  165.23 108.045 165.09 110.02 ;
      RECT  172.62 107.895 172.38 110.055 ;
      RECT  170.5 112.155 170.25 109.985 ;
      RECT  172.62 112.145 172.38 109.985 ;
      RECT  157.61 111.995 157.47 110.02 ;
      RECT  165.23 111.995 165.09 110.02 ;
      RECT  157.61 111.995 157.47 110.02 ;
      RECT  170.5 112.155 170.25 109.985 ;
      RECT  165.23 111.995 165.09 110.02 ;
      RECT  172.62 112.145 172.38 109.985 ;
      RECT  170.5 111.835 170.25 114.005 ;
      RECT  172.62 111.845 172.38 114.005 ;
      RECT  157.61 111.995 157.47 113.97 ;
      RECT  165.23 111.995 165.09 113.97 ;
      RECT  157.61 111.995 157.47 113.97 ;
      RECT  170.5 111.835 170.25 114.005 ;
      RECT  165.23 111.995 165.09 113.97 ;
      RECT  172.62 111.845 172.38 114.005 ;
      RECT  170.5 116.105 170.25 113.935 ;
      RECT  172.62 116.095 172.38 113.935 ;
      RECT  157.61 115.945 157.47 113.97 ;
      RECT  165.23 115.945 165.09 113.97 ;
      RECT  157.61 115.945 157.47 113.97 ;
      RECT  170.5 116.105 170.25 113.935 ;
      RECT  165.23 115.945 165.09 113.97 ;
      RECT  172.62 116.095 172.38 113.935 ;
      RECT  170.5 115.785 170.25 117.955 ;
      RECT  172.62 115.795 172.38 117.955 ;
      RECT  157.61 115.945 157.47 117.92 ;
      RECT  165.23 115.945 165.09 117.92 ;
      RECT  157.61 115.945 157.47 117.92 ;
      RECT  170.5 115.785 170.25 117.955 ;
      RECT  165.23 115.945 165.09 117.92 ;
      RECT  172.62 115.795 172.38 117.955 ;
      RECT  170.5 120.055 170.25 117.885 ;
      RECT  172.62 120.045 172.38 117.885 ;
      RECT  157.61 119.895 157.47 117.92 ;
      RECT  165.23 119.895 165.09 117.92 ;
      RECT  157.61 119.895 157.47 117.92 ;
      RECT  170.5 120.055 170.25 117.885 ;
      RECT  165.23 119.895 165.09 117.92 ;
      RECT  172.62 120.045 172.38 117.885 ;
      RECT  170.5 119.735 170.25 121.905 ;
      RECT  172.62 119.745 172.38 121.905 ;
      RECT  157.61 119.895 157.47 121.87 ;
      RECT  165.23 119.895 165.09 121.87 ;
      RECT  157.61 119.895 157.47 121.87 ;
      RECT  170.5 119.735 170.25 121.905 ;
      RECT  165.23 119.895 165.09 121.87 ;
      RECT  172.62 119.745 172.38 121.905 ;
      RECT  170.5 124.005 170.25 121.835 ;
      RECT  172.62 123.995 172.38 121.835 ;
      RECT  157.61 123.845 157.47 121.87 ;
      RECT  165.23 123.845 165.09 121.87 ;
      RECT  157.61 123.845 157.47 121.87 ;
      RECT  170.5 124.005 170.25 121.835 ;
      RECT  165.23 123.845 165.09 121.87 ;
      RECT  172.62 123.995 172.38 121.835 ;
      RECT  170.445 92.085 170.305 123.845 ;
      RECT  157.61 92.245 157.47 123.845 ;
      RECT  165.23 92.245 165.09 123.845 ;
      RECT  172.57 92.095 172.43 123.845 ;
      RECT  201.36 92.39 201.22 112.14 ;
      RECT  200.96 92.39 200.82 112.14 ;
      RECT  200.56 92.39 200.42 112.14 ;
      RECT  200.16 92.39 200.02 112.14 ;
      RECT  96.78 70.725 97.01 71.995 ;
      RECT  101.13 70.725 101.36 71.995 ;
      RECT  103.02 70.725 103.25 71.995 ;
      RECT  107.37 70.725 107.6 71.995 ;
      RECT  109.26 70.725 109.49 71.995 ;
      RECT  113.61 70.725 113.84 71.995 ;
      RECT  115.5 70.725 115.73 71.995 ;
      RECT  119.85 70.725 120.08 71.995 ;
      RECT  121.74 70.725 121.97 71.995 ;
      RECT  126.09 70.725 126.32 71.995 ;
      RECT  127.98 70.725 128.21 71.995 ;
      RECT  132.33 70.725 132.56 71.995 ;
      RECT  134.22 70.725 134.45 71.995 ;
      RECT  138.57 70.725 138.8 71.995 ;
      RECT  140.46 70.725 140.69 71.995 ;
      RECT  144.81 70.725 145.04 71.995 ;
      RECT  96.78 144.095 97.01 145.365 ;
      RECT  101.13 144.095 101.36 145.365 ;
      RECT  103.02 144.095 103.25 145.365 ;
      RECT  107.37 144.095 107.6 145.365 ;
      RECT  109.26 144.095 109.49 145.365 ;
      RECT  113.61 144.095 113.84 145.365 ;
      RECT  115.5 144.095 115.73 145.365 ;
      RECT  119.85 144.095 120.08 145.365 ;
      RECT  121.74 144.095 121.97 145.365 ;
      RECT  126.09 144.095 126.32 145.365 ;
      RECT  127.98 144.095 128.21 145.365 ;
      RECT  132.33 144.095 132.56 145.365 ;
      RECT  134.22 144.095 134.45 145.365 ;
      RECT  138.57 144.095 138.8 145.365 ;
      RECT  140.46 144.095 140.69 145.365 ;
      RECT  144.81 144.095 145.04 145.365 ;
      RECT  97.535 59.43 97.835 59.71 ;
      RECT  100.305 59.43 100.605 59.71 ;
      RECT  103.775 59.43 104.075 59.71 ;
      RECT  106.545 59.43 106.845 59.71 ;
      RECT  110.015 59.43 110.315 59.71 ;
      RECT  112.785 59.43 113.085 59.71 ;
      RECT  116.255 59.43 116.555 59.71 ;
      RECT  119.025 59.43 119.325 59.71 ;
      RECT  122.495 59.43 122.795 59.71 ;
      RECT  125.265 59.43 125.565 59.71 ;
      RECT  128.735 59.43 129.035 59.71 ;
      RECT  131.505 59.43 131.805 59.71 ;
      RECT  134.975 59.43 135.275 59.71 ;
      RECT  137.745 59.43 138.045 59.71 ;
      RECT  141.215 59.43 141.515 59.71 ;
      RECT  143.985 59.43 144.285 59.71 ;
      RECT  41.08 92.39 41.22 112.14 ;
      RECT  41.48 92.39 41.62 112.14 ;
      RECT  41.88 92.39 42.02 112.14 ;
      RECT  42.28 92.39 42.42 112.14 ;
      RECT  201.22 92.39 201.36 112.14 ;
      RECT  200.82 92.39 200.96 112.14 ;
      RECT  200.42 92.39 200.56 112.14 ;
      RECT  200.02 92.39 200.16 112.14 ;
      RECT  0.74 33.24 1.03 33.47 ;
      RECT  5.16 32.27 5.33 33.24 ;
      RECT  6.11 32.27 6.28 33.98 ;
      RECT  3.855 32.27 4.025 34.84 ;
      RECT  0.8 32.27 0.97 33.24 ;
      RECT  2.515 33.115 2.685 34.395 ;
      RECT  2.455 32.84 2.745 33.07 ;
      RECT  2.455 34.44 2.745 34.67 ;
      RECT  2.465 32.795 2.735 32.84 ;
      RECT  5.1 34.84 5.39 35.07 ;
      RECT  2.045 34.84 2.335 35.07 ;
      RECT  5.1 33.24 5.39 33.47 ;
      RECT  1.125 34.07 2.275 34.24 ;
      RECT  6.05 34.84 6.34 35.07 ;
      RECT  0.74 34.84 1.03 35.07 ;
      RECT  2.045 32.04 2.335 32.27 ;
      RECT  6.03 33.98 6.36 34.24 ;
      RECT  1.125 34.04 1.415 34.07 ;
      RECT  0.8 33.47 0.97 34.84 ;
      RECT  2.105 32.27 2.275 34.07 ;
      RECT  2.465 34.395 2.735 34.44 ;
      RECT  5.64 33.225 5.97 33.485 ;
      RECT  5.16 33.47 5.33 34.84 ;
      RECT  6.11 34.24 6.28 34.84 ;
      RECT  1.125 34.24 1.415 34.27 ;
      RECT  2.465 34.67 2.735 34.715 ;
      RECT  3.795 32.04 4.085 32.27 ;
      RECT  2.105 34.24 2.275 34.84 ;
      RECT  3.795 34.84 4.085 35.07 ;
      RECT  5.1 32.04 5.39 32.27 ;
      RECT  2.465 33.07 2.735 33.115 ;
      RECT  0.74 32.04 1.03 32.27 ;
      RECT  1.305 33.625 1.635 33.885 ;
      RECT  6.05 32.04 6.34 32.27 ;
      RECT  0.74 42.77 1.03 42.54 ;
      RECT  5.16 43.74 5.33 42.77 ;
      RECT  6.11 43.74 6.28 42.03 ;
      RECT  3.855 43.74 4.025 41.17 ;
      RECT  0.8 43.74 0.97 42.77 ;
      RECT  2.515 42.895 2.685 41.615 ;
      RECT  2.455 43.17 2.745 42.94 ;
      RECT  2.455 41.57 2.745 41.34 ;
      RECT  2.465 43.215 2.735 43.17 ;
      RECT  5.1 41.17 5.39 40.94 ;
      RECT  2.045 41.17 2.335 40.94 ;
      RECT  5.1 42.77 5.39 42.54 ;
      RECT  1.125 41.94 2.275 41.77 ;
      RECT  6.05 41.17 6.34 40.94 ;
      RECT  0.74 41.17 1.03 40.94 ;
      RECT  2.045 43.97 2.335 43.74 ;
      RECT  6.03 42.03 6.36 41.77 ;
      RECT  1.125 41.97 1.415 41.94 ;
      RECT  0.8 42.54 0.97 41.17 ;
      RECT  2.105 43.74 2.275 41.94 ;
      RECT  2.465 41.615 2.735 41.57 ;
      RECT  5.64 42.785 5.97 42.525 ;
      RECT  5.16 42.54 5.33 41.17 ;
      RECT  6.11 41.77 6.28 41.17 ;
      RECT  1.125 41.77 1.415 41.74 ;
      RECT  2.465 41.34 2.735 41.295 ;
      RECT  3.795 43.97 4.085 43.74 ;
      RECT  2.105 41.77 2.275 41.17 ;
      RECT  3.795 41.17 4.085 40.94 ;
      RECT  5.1 43.97 5.39 43.74 ;
      RECT  2.465 42.94 2.735 42.895 ;
      RECT  0.74 43.97 1.03 43.74 ;
      RECT  1.305 42.385 1.635 42.125 ;
      RECT  6.05 43.97 6.34 43.74 ;
      RECT  240.62 168.71 240.33 168.48 ;
      RECT  236.2 169.68 236.03 168.71 ;
      RECT  235.25 169.68 235.08 167.97 ;
      RECT  237.505 169.68 237.335 167.11 ;
      RECT  240.56 169.68 240.39 168.71 ;
      RECT  238.845 168.835 238.675 167.555 ;
      RECT  238.905 169.11 238.615 168.88 ;
      RECT  238.905 167.51 238.615 167.28 ;
      RECT  238.895 169.155 238.625 169.11 ;
      RECT  236.26 167.11 235.97 166.88 ;
      RECT  239.315 167.11 239.025 166.88 ;
      RECT  236.26 168.71 235.97 168.48 ;
      RECT  240.235 167.88 239.085 167.71 ;
      RECT  235.31 167.11 235.02 166.88 ;
      RECT  240.62 167.11 240.33 166.88 ;
      RECT  239.315 169.91 239.025 169.68 ;
      RECT  235.33 167.97 235.0 167.71 ;
      RECT  240.235 167.91 239.945 167.88 ;
      RECT  240.56 168.48 240.39 167.11 ;
      RECT  239.255 169.68 239.085 167.88 ;
      RECT  238.895 167.555 238.625 167.51 ;
      RECT  235.72 168.725 235.39 168.465 ;
      RECT  236.2 168.48 236.03 167.11 ;
      RECT  235.25 167.71 235.08 167.11 ;
      RECT  240.235 167.71 239.945 167.68 ;
      RECT  238.895 167.28 238.625 167.235 ;
      RECT  237.565 169.91 237.275 169.68 ;
      RECT  239.255 167.71 239.085 167.11 ;
      RECT  237.565 167.11 237.275 166.88 ;
      RECT  236.26 169.91 235.97 169.68 ;
      RECT  238.895 168.88 238.625 168.835 ;
      RECT  240.62 169.91 240.33 169.68 ;
      RECT  240.055 168.325 239.725 168.065 ;
      RECT  235.31 169.91 235.02 169.68 ;
      RECT  34.43 141.8 34.72 142.03 ;
      RECT  38.85 140.83 39.02 141.8 ;
      RECT  39.8 140.83 39.97 142.54 ;
      RECT  37.545 140.83 37.715 143.4 ;
      RECT  34.49 140.83 34.66 141.8 ;
      RECT  36.205 141.675 36.375 142.955 ;
      RECT  36.145 141.4 36.435 141.63 ;
      RECT  36.145 143.0 36.435 143.23 ;
      RECT  36.155 141.355 36.425 141.4 ;
      RECT  38.79 143.4 39.08 143.63 ;
      RECT  35.735 143.4 36.025 143.63 ;
      RECT  38.79 141.8 39.08 142.03 ;
      RECT  34.815 142.63 35.965 142.8 ;
      RECT  39.74 143.4 40.03 143.63 ;
      RECT  34.43 143.4 34.72 143.63 ;
      RECT  35.735 140.6 36.025 140.83 ;
      RECT  39.72 142.54 40.05 142.8 ;
      RECT  34.815 142.6 35.105 142.63 ;
      RECT  34.49 142.03 34.66 143.4 ;
      RECT  35.795 140.83 35.965 142.63 ;
      RECT  36.155 142.955 36.425 143.0 ;
      RECT  39.33 141.785 39.66 142.045 ;
      RECT  38.85 142.03 39.02 143.4 ;
      RECT  39.8 142.8 39.97 143.4 ;
      RECT  34.815 142.8 35.105 142.83 ;
      RECT  36.155 143.23 36.425 143.275 ;
      RECT  37.485 140.6 37.775 140.83 ;
      RECT  35.795 142.8 35.965 143.4 ;
      RECT  37.485 143.4 37.775 143.63 ;
      RECT  38.79 140.6 39.08 140.83 ;
      RECT  36.155 141.63 36.425 141.675 ;
      RECT  34.43 140.6 34.72 140.83 ;
      RECT  34.995 142.185 35.325 142.445 ;
      RECT  39.74 140.6 40.03 140.83 ;
      RECT  34.43 151.33 34.72 151.1 ;
      RECT  38.85 152.3 39.02 151.33 ;
      RECT  39.8 152.3 39.97 150.59 ;
      RECT  37.545 152.3 37.715 149.73 ;
      RECT  34.49 152.3 34.66 151.33 ;
      RECT  36.205 151.455 36.375 150.175 ;
      RECT  36.145 151.73 36.435 151.5 ;
      RECT  36.145 150.13 36.435 149.9 ;
      RECT  36.155 151.775 36.425 151.73 ;
      RECT  38.79 149.73 39.08 149.5 ;
      RECT  35.735 149.73 36.025 149.5 ;
      RECT  38.79 151.33 39.08 151.1 ;
      RECT  34.815 150.5 35.965 150.33 ;
      RECT  39.74 149.73 40.03 149.5 ;
      RECT  34.43 149.73 34.72 149.5 ;
      RECT  35.735 152.53 36.025 152.3 ;
      RECT  39.72 150.59 40.05 150.33 ;
      RECT  34.815 150.53 35.105 150.5 ;
      RECT  34.49 151.1 34.66 149.73 ;
      RECT  35.795 152.3 35.965 150.5 ;
      RECT  36.155 150.175 36.425 150.13 ;
      RECT  39.33 151.345 39.66 151.085 ;
      RECT  38.85 151.1 39.02 149.73 ;
      RECT  39.8 150.33 39.97 149.73 ;
      RECT  34.815 150.33 35.105 150.3 ;
      RECT  36.155 149.9 36.425 149.855 ;
      RECT  37.485 152.53 37.775 152.3 ;
      RECT  35.795 150.33 35.965 149.73 ;
      RECT  37.485 149.73 37.775 149.5 ;
      RECT  38.79 152.53 39.08 152.3 ;
      RECT  36.155 151.5 36.425 151.455 ;
      RECT  34.43 152.53 34.72 152.3 ;
      RECT  34.995 150.945 35.325 150.685 ;
      RECT  39.74 152.53 40.03 152.3 ;
      RECT  34.43 155.94 34.72 156.17 ;
      RECT  38.85 154.97 39.02 155.94 ;
      RECT  39.8 154.97 39.97 156.68 ;
      RECT  37.545 154.97 37.715 157.54 ;
      RECT  34.49 154.97 34.66 155.94 ;
      RECT  36.205 155.815 36.375 157.095 ;
      RECT  36.145 155.54 36.435 155.77 ;
      RECT  36.145 157.14 36.435 157.37 ;
      RECT  36.155 155.495 36.425 155.54 ;
      RECT  38.79 157.54 39.08 157.77 ;
      RECT  35.735 157.54 36.025 157.77 ;
      RECT  38.79 155.94 39.08 156.17 ;
      RECT  34.815 156.77 35.965 156.94 ;
      RECT  39.74 157.54 40.03 157.77 ;
      RECT  34.43 157.54 34.72 157.77 ;
      RECT  35.735 154.74 36.025 154.97 ;
      RECT  39.72 156.68 40.05 156.94 ;
      RECT  34.815 156.74 35.105 156.77 ;
      RECT  34.49 156.17 34.66 157.54 ;
      RECT  35.795 154.97 35.965 156.77 ;
      RECT  36.155 157.095 36.425 157.14 ;
      RECT  39.33 155.925 39.66 156.185 ;
      RECT  38.85 156.17 39.02 157.54 ;
      RECT  39.8 156.94 39.97 157.54 ;
      RECT  34.815 156.94 35.105 156.97 ;
      RECT  36.155 157.37 36.425 157.415 ;
      RECT  37.485 154.74 37.775 154.97 ;
      RECT  35.795 156.94 35.965 157.54 ;
      RECT  37.485 157.54 37.775 157.77 ;
      RECT  38.79 154.74 39.08 154.97 ;
      RECT  36.155 155.77 36.425 155.815 ;
      RECT  34.43 154.74 34.72 154.97 ;
      RECT  34.995 156.325 35.325 156.585 ;
      RECT  39.74 154.74 40.03 154.97 ;
      RECT  34.43 165.47 34.72 165.24 ;
      RECT  38.85 166.44 39.02 165.47 ;
      RECT  39.8 166.44 39.97 164.73 ;
      RECT  37.545 166.44 37.715 163.87 ;
      RECT  34.49 166.44 34.66 165.47 ;
      RECT  36.205 165.595 36.375 164.315 ;
      RECT  36.145 165.87 36.435 165.64 ;
      RECT  36.145 164.27 36.435 164.04 ;
      RECT  36.155 165.915 36.425 165.87 ;
      RECT  38.79 163.87 39.08 163.64 ;
      RECT  35.735 163.87 36.025 163.64 ;
      RECT  38.79 165.47 39.08 165.24 ;
      RECT  34.815 164.64 35.965 164.47 ;
      RECT  39.74 163.87 40.03 163.64 ;
      RECT  34.43 163.87 34.72 163.64 ;
      RECT  35.735 166.67 36.025 166.44 ;
      RECT  39.72 164.73 40.05 164.47 ;
      RECT  34.815 164.67 35.105 164.64 ;
      RECT  34.49 165.24 34.66 163.87 ;
      RECT  35.795 166.44 35.965 164.64 ;
      RECT  36.155 164.315 36.425 164.27 ;
      RECT  39.33 165.485 39.66 165.225 ;
      RECT  38.85 165.24 39.02 163.87 ;
      RECT  39.8 164.47 39.97 163.87 ;
      RECT  34.815 164.47 35.105 164.44 ;
      RECT  36.155 164.04 36.425 163.995 ;
      RECT  37.485 166.67 37.775 166.44 ;
      RECT  35.795 164.47 35.965 163.87 ;
      RECT  37.485 163.87 37.775 163.64 ;
      RECT  38.79 166.67 39.08 166.44 ;
      RECT  36.155 165.64 36.425 165.595 ;
      RECT  34.43 166.67 34.72 166.44 ;
      RECT  34.995 165.085 35.325 164.825 ;
      RECT  39.74 166.67 40.03 166.44 ;
      RECT  208.43 74.29 208.14 74.06 ;
      RECT  204.01 75.26 203.84 74.29 ;
      RECT  203.06 75.26 202.89 73.55 ;
      RECT  205.315 75.26 205.145 72.69 ;
      RECT  208.37 75.26 208.2 74.29 ;
      RECT  206.655 74.415 206.485 73.135 ;
      RECT  206.715 74.69 206.425 74.46 ;
      RECT  206.715 73.09 206.425 72.86 ;
      RECT  206.705 74.735 206.435 74.69 ;
      RECT  204.07 72.69 203.78 72.46 ;
      RECT  207.125 72.69 206.835 72.46 ;
      RECT  204.07 74.29 203.78 74.06 ;
      RECT  208.045 73.46 206.895 73.29 ;
      RECT  203.12 72.69 202.83 72.46 ;
      RECT  208.43 72.69 208.14 72.46 ;
      RECT  207.125 75.49 206.835 75.26 ;
      RECT  203.14 73.55 202.81 73.29 ;
      RECT  208.045 73.49 207.755 73.46 ;
      RECT  208.37 74.06 208.2 72.69 ;
      RECT  207.065 75.26 206.895 73.46 ;
      RECT  206.705 73.135 206.435 73.09 ;
      RECT  203.53 74.305 203.2 74.045 ;
      RECT  204.01 74.06 203.84 72.69 ;
      RECT  203.06 73.29 202.89 72.69 ;
      RECT  208.045 73.29 207.755 73.26 ;
      RECT  206.705 72.86 206.435 72.815 ;
      RECT  205.375 75.49 205.085 75.26 ;
      RECT  207.065 73.29 206.895 72.69 ;
      RECT  205.375 72.69 205.085 72.46 ;
      RECT  204.07 75.49 203.78 75.26 ;
      RECT  206.705 74.46 206.435 74.415 ;
      RECT  208.43 75.49 208.14 75.26 ;
      RECT  207.865 73.905 207.535 73.645 ;
      RECT  203.12 75.49 202.83 75.26 ;
      RECT  208.43 64.76 208.14 64.99 ;
      RECT  204.01 63.79 203.84 64.76 ;
      RECT  203.06 63.79 202.89 65.5 ;
      RECT  205.315 63.79 205.145 66.36 ;
      RECT  208.37 63.79 208.2 64.76 ;
      RECT  206.655 64.635 206.485 65.915 ;
      RECT  206.715 64.36 206.425 64.59 ;
      RECT  206.715 65.96 206.425 66.19 ;
      RECT  206.705 64.315 206.435 64.36 ;
      RECT  204.07 66.36 203.78 66.59 ;
      RECT  207.125 66.36 206.835 66.59 ;
      RECT  204.07 64.76 203.78 64.99 ;
      RECT  208.045 65.59 206.895 65.76 ;
      RECT  203.12 66.36 202.83 66.59 ;
      RECT  208.43 66.36 208.14 66.59 ;
      RECT  207.125 63.56 206.835 63.79 ;
      RECT  203.14 65.5 202.81 65.76 ;
      RECT  208.045 65.56 207.755 65.59 ;
      RECT  208.37 64.99 208.2 66.36 ;
      RECT  207.065 63.79 206.895 65.59 ;
      RECT  206.705 65.915 206.435 65.96 ;
      RECT  203.53 64.745 203.2 65.005 ;
      RECT  204.01 64.99 203.84 66.36 ;
      RECT  203.06 65.76 202.89 66.36 ;
      RECT  208.045 65.76 207.755 65.79 ;
      RECT  206.705 66.19 206.435 66.235 ;
      RECT  205.375 63.56 205.085 63.79 ;
      RECT  207.065 65.76 206.895 66.36 ;
      RECT  205.375 66.36 205.085 66.59 ;
      RECT  204.07 63.56 203.78 63.79 ;
      RECT  206.705 64.59 206.435 64.635 ;
      RECT  208.43 63.56 208.14 63.79 ;
      RECT  207.865 65.145 207.535 65.405 ;
      RECT  203.12 63.56 202.83 63.79 ;
      RECT  208.43 60.15 208.14 59.92 ;
      RECT  204.01 61.12 203.84 60.15 ;
      RECT  203.06 61.12 202.89 59.41 ;
      RECT  205.315 61.12 205.145 58.55 ;
      RECT  208.37 61.12 208.2 60.15 ;
      RECT  206.655 60.275 206.485 58.995 ;
      RECT  206.715 60.55 206.425 60.32 ;
      RECT  206.715 58.95 206.425 58.72 ;
      RECT  206.705 60.595 206.435 60.55 ;
      RECT  204.07 58.55 203.78 58.32 ;
      RECT  207.125 58.55 206.835 58.32 ;
      RECT  204.07 60.15 203.78 59.92 ;
      RECT  208.045 59.32 206.895 59.15 ;
      RECT  203.12 58.55 202.83 58.32 ;
      RECT  208.43 58.55 208.14 58.32 ;
      RECT  207.125 61.35 206.835 61.12 ;
      RECT  203.14 59.41 202.81 59.15 ;
      RECT  208.045 59.35 207.755 59.32 ;
      RECT  208.37 59.92 208.2 58.55 ;
      RECT  207.065 61.12 206.895 59.32 ;
      RECT  206.705 58.995 206.435 58.95 ;
      RECT  203.53 60.165 203.2 59.905 ;
      RECT  204.01 59.92 203.84 58.55 ;
      RECT  203.06 59.15 202.89 58.55 ;
      RECT  208.045 59.15 207.755 59.12 ;
      RECT  206.705 58.72 206.435 58.675 ;
      RECT  205.375 61.35 205.085 61.12 ;
      RECT  207.065 59.15 206.895 58.55 ;
      RECT  205.375 58.55 205.085 58.32 ;
      RECT  204.07 61.35 203.78 61.12 ;
      RECT  206.705 60.32 206.435 60.275 ;
      RECT  208.43 61.35 208.14 61.12 ;
      RECT  207.865 59.765 207.535 59.505 ;
      RECT  203.12 61.35 202.83 61.12 ;
      RECT  208.43 50.62 208.14 50.85 ;
      RECT  204.01 49.65 203.84 50.62 ;
      RECT  203.06 49.65 202.89 51.36 ;
      RECT  205.315 49.65 205.145 52.22 ;
      RECT  208.37 49.65 208.2 50.62 ;
      RECT  206.655 50.495 206.485 51.775 ;
      RECT  206.715 50.22 206.425 50.45 ;
      RECT  206.715 51.82 206.425 52.05 ;
      RECT  206.705 50.175 206.435 50.22 ;
      RECT  204.07 52.22 203.78 52.45 ;
      RECT  207.125 52.22 206.835 52.45 ;
      RECT  204.07 50.62 203.78 50.85 ;
      RECT  208.045 51.45 206.895 51.62 ;
      RECT  203.12 52.22 202.83 52.45 ;
      RECT  208.43 52.22 208.14 52.45 ;
      RECT  207.125 49.42 206.835 49.65 ;
      RECT  203.14 51.36 202.81 51.62 ;
      RECT  208.045 51.42 207.755 51.45 ;
      RECT  208.37 50.85 208.2 52.22 ;
      RECT  207.065 49.65 206.895 51.45 ;
      RECT  206.705 51.775 206.435 51.82 ;
      RECT  203.53 50.605 203.2 50.865 ;
      RECT  204.01 50.85 203.84 52.22 ;
      RECT  203.06 51.62 202.89 52.22 ;
      RECT  208.045 51.62 207.755 51.65 ;
      RECT  206.705 52.05 206.435 52.095 ;
      RECT  205.375 49.42 205.085 49.65 ;
      RECT  207.065 51.62 206.895 52.22 ;
      RECT  205.375 52.22 205.085 52.45 ;
      RECT  204.07 49.42 203.78 49.65 ;
      RECT  206.705 50.45 206.435 50.495 ;
      RECT  208.43 49.42 208.14 49.65 ;
      RECT  207.865 51.005 207.535 51.265 ;
      RECT  203.12 49.42 202.83 49.65 ;
      RECT  46.11 2.645 46.4 2.875 ;
      RECT  50.53 1.675 50.7 2.645 ;
      RECT  51.48 1.675 51.65 3.385 ;
      RECT  49.225 1.675 49.395 4.245 ;
      RECT  46.17 1.675 46.34 2.645 ;
      RECT  47.885 2.52 48.055 3.8 ;
      RECT  47.825 2.245 48.115 2.475 ;
      RECT  47.825 3.845 48.115 4.075 ;
      RECT  47.835 2.2 48.105 2.245 ;
      RECT  50.47 4.245 50.76 4.475 ;
      RECT  47.415 4.245 47.705 4.475 ;
      RECT  50.47 2.645 50.76 2.875 ;
      RECT  46.495 3.475 47.645 3.645 ;
      RECT  51.42 4.245 51.71 4.475 ;
      RECT  46.11 4.245 46.4 4.475 ;
      RECT  47.415 1.445 47.705 1.675 ;
      RECT  51.4 3.385 51.73 3.645 ;
      RECT  46.495 3.445 46.785 3.475 ;
      RECT  46.17 2.875 46.34 4.245 ;
      RECT  47.475 1.675 47.645 3.475 ;
      RECT  47.835 3.8 48.105 3.845 ;
      RECT  51.01 2.63 51.34 2.89 ;
      RECT  50.53 2.875 50.7 4.245 ;
      RECT  51.48 3.645 51.65 4.245 ;
      RECT  46.495 3.645 46.785 3.675 ;
      RECT  47.835 4.075 48.105 4.12 ;
      RECT  49.165 1.445 49.455 1.675 ;
      RECT  47.475 3.645 47.645 4.245 ;
      RECT  49.165 4.245 49.455 4.475 ;
      RECT  50.47 1.445 50.76 1.675 ;
      RECT  47.835 2.475 48.105 2.52 ;
      RECT  46.11 1.445 46.4 1.675 ;
      RECT  46.675 3.03 47.005 3.29 ;
      RECT  51.42 1.445 51.71 1.675 ;
      RECT  51.95 2.645 52.24 2.875 ;
      RECT  56.37 1.675 56.54 2.645 ;
      RECT  57.32 1.675 57.49 3.385 ;
      RECT  55.065 1.675 55.235 4.245 ;
      RECT  52.01 1.675 52.18 2.645 ;
      RECT  53.725 2.52 53.895 3.8 ;
      RECT  53.665 2.245 53.955 2.475 ;
      RECT  53.665 3.845 53.955 4.075 ;
      RECT  53.675 2.2 53.945 2.245 ;
      RECT  56.31 4.245 56.6 4.475 ;
      RECT  53.255 4.245 53.545 4.475 ;
      RECT  56.31 2.645 56.6 2.875 ;
      RECT  52.335 3.475 53.485 3.645 ;
      RECT  57.26 4.245 57.55 4.475 ;
      RECT  51.95 4.245 52.24 4.475 ;
      RECT  53.255 1.445 53.545 1.675 ;
      RECT  57.24 3.385 57.57 3.645 ;
      RECT  52.335 3.445 52.625 3.475 ;
      RECT  52.01 2.875 52.18 4.245 ;
      RECT  53.315 1.675 53.485 3.475 ;
      RECT  53.675 3.8 53.945 3.845 ;
      RECT  56.85 2.63 57.18 2.89 ;
      RECT  56.37 2.875 56.54 4.245 ;
      RECT  57.32 3.645 57.49 4.245 ;
      RECT  52.335 3.645 52.625 3.675 ;
      RECT  53.675 4.075 53.945 4.12 ;
      RECT  55.005 1.445 55.295 1.675 ;
      RECT  53.315 3.645 53.485 4.245 ;
      RECT  55.005 4.245 55.295 4.475 ;
      RECT  56.31 1.445 56.6 1.675 ;
      RECT  53.675 2.475 53.945 2.52 ;
      RECT  51.95 1.445 52.24 1.675 ;
      RECT  52.515 3.03 52.845 3.29 ;
      RECT  57.26 1.445 57.55 1.675 ;
      RECT  57.79 2.645 58.08 2.875 ;
      RECT  62.21 1.675 62.38 2.645 ;
      RECT  63.16 1.675 63.33 3.385 ;
      RECT  60.905 1.675 61.075 4.245 ;
      RECT  57.85 1.675 58.02 2.645 ;
      RECT  59.565 2.52 59.735 3.8 ;
      RECT  59.505 2.245 59.795 2.475 ;
      RECT  59.505 3.845 59.795 4.075 ;
      RECT  59.515 2.2 59.785 2.245 ;
      RECT  62.15 4.245 62.44 4.475 ;
      RECT  59.095 4.245 59.385 4.475 ;
      RECT  62.15 2.645 62.44 2.875 ;
      RECT  58.175 3.475 59.325 3.645 ;
      RECT  63.1 4.245 63.39 4.475 ;
      RECT  57.79 4.245 58.08 4.475 ;
      RECT  59.095 1.445 59.385 1.675 ;
      RECT  63.08 3.385 63.41 3.645 ;
      RECT  58.175 3.445 58.465 3.475 ;
      RECT  57.85 2.875 58.02 4.245 ;
      RECT  59.155 1.675 59.325 3.475 ;
      RECT  59.515 3.8 59.785 3.845 ;
      RECT  62.69 2.63 63.02 2.89 ;
      RECT  62.21 2.875 62.38 4.245 ;
      RECT  63.16 3.645 63.33 4.245 ;
      RECT  58.175 3.645 58.465 3.675 ;
      RECT  59.515 4.075 59.785 4.12 ;
      RECT  60.845 1.445 61.135 1.675 ;
      RECT  59.155 3.645 59.325 4.245 ;
      RECT  60.845 4.245 61.135 4.475 ;
      RECT  62.15 1.445 62.44 1.675 ;
      RECT  59.515 2.475 59.785 2.52 ;
      RECT  57.79 1.445 58.08 1.675 ;
      RECT  58.355 3.03 58.685 3.29 ;
      RECT  63.1 1.445 63.39 1.675 ;
      RECT  63.63 2.645 63.92 2.875 ;
      RECT  68.05 1.675 68.22 2.645 ;
      RECT  69.0 1.675 69.17 3.385 ;
      RECT  66.745 1.675 66.915 4.245 ;
      RECT  63.69 1.675 63.86 2.645 ;
      RECT  65.405 2.52 65.575 3.8 ;
      RECT  65.345 2.245 65.635 2.475 ;
      RECT  65.345 3.845 65.635 4.075 ;
      RECT  65.355 2.2 65.625 2.245 ;
      RECT  67.99 4.245 68.28 4.475 ;
      RECT  64.935 4.245 65.225 4.475 ;
      RECT  67.99 2.645 68.28 2.875 ;
      RECT  64.015 3.475 65.165 3.645 ;
      RECT  68.94 4.245 69.23 4.475 ;
      RECT  63.63 4.245 63.92 4.475 ;
      RECT  64.935 1.445 65.225 1.675 ;
      RECT  68.92 3.385 69.25 3.645 ;
      RECT  64.015 3.445 64.305 3.475 ;
      RECT  63.69 2.875 63.86 4.245 ;
      RECT  64.995 1.675 65.165 3.475 ;
      RECT  65.355 3.8 65.625 3.845 ;
      RECT  68.53 2.63 68.86 2.89 ;
      RECT  68.05 2.875 68.22 4.245 ;
      RECT  69.0 3.645 69.17 4.245 ;
      RECT  64.015 3.645 64.305 3.675 ;
      RECT  65.355 4.075 65.625 4.12 ;
      RECT  66.685 1.445 66.975 1.675 ;
      RECT  64.995 3.645 65.165 4.245 ;
      RECT  66.685 4.245 66.975 4.475 ;
      RECT  67.99 1.445 68.28 1.675 ;
      RECT  65.355 2.475 65.625 2.52 ;
      RECT  63.63 1.445 63.92 1.675 ;
      RECT  64.195 3.03 64.525 3.29 ;
      RECT  68.94 1.445 69.23 1.675 ;
      RECT  69.47 2.645 69.76 2.875 ;
      RECT  73.89 1.675 74.06 2.645 ;
      RECT  74.84 1.675 75.01 3.385 ;
      RECT  72.585 1.675 72.755 4.245 ;
      RECT  69.53 1.675 69.7 2.645 ;
      RECT  71.245 2.52 71.415 3.8 ;
      RECT  71.185 2.245 71.475 2.475 ;
      RECT  71.185 3.845 71.475 4.075 ;
      RECT  71.195 2.2 71.465 2.245 ;
      RECT  73.83 4.245 74.12 4.475 ;
      RECT  70.775 4.245 71.065 4.475 ;
      RECT  73.83 2.645 74.12 2.875 ;
      RECT  69.855 3.475 71.005 3.645 ;
      RECT  74.78 4.245 75.07 4.475 ;
      RECT  69.47 4.245 69.76 4.475 ;
      RECT  70.775 1.445 71.065 1.675 ;
      RECT  74.76 3.385 75.09 3.645 ;
      RECT  69.855 3.445 70.145 3.475 ;
      RECT  69.53 2.875 69.7 4.245 ;
      RECT  70.835 1.675 71.005 3.475 ;
      RECT  71.195 3.8 71.465 3.845 ;
      RECT  74.37 2.63 74.7 2.89 ;
      RECT  73.89 2.875 74.06 4.245 ;
      RECT  74.84 3.645 75.01 4.245 ;
      RECT  69.855 3.645 70.145 3.675 ;
      RECT  71.195 4.075 71.465 4.12 ;
      RECT  72.525 1.445 72.815 1.675 ;
      RECT  70.835 3.645 71.005 4.245 ;
      RECT  72.525 4.245 72.815 4.475 ;
      RECT  73.83 1.445 74.12 1.675 ;
      RECT  71.195 2.475 71.465 2.52 ;
      RECT  69.47 1.445 69.76 1.675 ;
      RECT  70.035 3.03 70.365 3.29 ;
      RECT  74.78 1.445 75.07 1.675 ;
      RECT  75.31 2.645 75.6 2.875 ;
      RECT  79.73 1.675 79.9 2.645 ;
      RECT  80.68 1.675 80.85 3.385 ;
      RECT  78.425 1.675 78.595 4.245 ;
      RECT  75.37 1.675 75.54 2.645 ;
      RECT  77.085 2.52 77.255 3.8 ;
      RECT  77.025 2.245 77.315 2.475 ;
      RECT  77.025 3.845 77.315 4.075 ;
      RECT  77.035 2.2 77.305 2.245 ;
      RECT  79.67 4.245 79.96 4.475 ;
      RECT  76.615 4.245 76.905 4.475 ;
      RECT  79.67 2.645 79.96 2.875 ;
      RECT  75.695 3.475 76.845 3.645 ;
      RECT  80.62 4.245 80.91 4.475 ;
      RECT  75.31 4.245 75.6 4.475 ;
      RECT  76.615 1.445 76.905 1.675 ;
      RECT  80.6 3.385 80.93 3.645 ;
      RECT  75.695 3.445 75.985 3.475 ;
      RECT  75.37 2.875 75.54 4.245 ;
      RECT  76.675 1.675 76.845 3.475 ;
      RECT  77.035 3.8 77.305 3.845 ;
      RECT  80.21 2.63 80.54 2.89 ;
      RECT  79.73 2.875 79.9 4.245 ;
      RECT  80.68 3.645 80.85 4.245 ;
      RECT  75.695 3.645 75.985 3.675 ;
      RECT  77.035 4.075 77.305 4.12 ;
      RECT  78.365 1.445 78.655 1.675 ;
      RECT  76.675 3.645 76.845 4.245 ;
      RECT  78.365 4.245 78.655 4.475 ;
      RECT  79.67 1.445 79.96 1.675 ;
      RECT  77.035 2.475 77.305 2.52 ;
      RECT  75.31 1.445 75.6 1.675 ;
      RECT  75.875 3.03 76.205 3.29 ;
      RECT  80.62 1.445 80.91 1.675 ;
      RECT  81.15 2.645 81.44 2.875 ;
      RECT  85.57 1.675 85.74 2.645 ;
      RECT  86.52 1.675 86.69 3.385 ;
      RECT  84.265 1.675 84.435 4.245 ;
      RECT  81.21 1.675 81.38 2.645 ;
      RECT  82.925 2.52 83.095 3.8 ;
      RECT  82.865 2.245 83.155 2.475 ;
      RECT  82.865 3.845 83.155 4.075 ;
      RECT  82.875 2.2 83.145 2.245 ;
      RECT  85.51 4.245 85.8 4.475 ;
      RECT  82.455 4.245 82.745 4.475 ;
      RECT  85.51 2.645 85.8 2.875 ;
      RECT  81.535 3.475 82.685 3.645 ;
      RECT  86.46 4.245 86.75 4.475 ;
      RECT  81.15 4.245 81.44 4.475 ;
      RECT  82.455 1.445 82.745 1.675 ;
      RECT  86.44 3.385 86.77 3.645 ;
      RECT  81.535 3.445 81.825 3.475 ;
      RECT  81.21 2.875 81.38 4.245 ;
      RECT  82.515 1.675 82.685 3.475 ;
      RECT  82.875 3.8 83.145 3.845 ;
      RECT  86.05 2.63 86.38 2.89 ;
      RECT  85.57 2.875 85.74 4.245 ;
      RECT  86.52 3.645 86.69 4.245 ;
      RECT  81.535 3.645 81.825 3.675 ;
      RECT  82.875 4.075 83.145 4.12 ;
      RECT  84.205 1.445 84.495 1.675 ;
      RECT  82.515 3.645 82.685 4.245 ;
      RECT  84.205 4.245 84.495 4.475 ;
      RECT  85.51 1.445 85.8 1.675 ;
      RECT  82.875 2.475 83.145 2.52 ;
      RECT  81.15 1.445 81.44 1.675 ;
      RECT  81.715 3.03 82.045 3.29 ;
      RECT  86.46 1.445 86.75 1.675 ;
      RECT  86.99 2.645 87.28 2.875 ;
      RECT  91.41 1.675 91.58 2.645 ;
      RECT  92.36 1.675 92.53 3.385 ;
      RECT  90.105 1.675 90.275 4.245 ;
      RECT  87.05 1.675 87.22 2.645 ;
      RECT  88.765 2.52 88.935 3.8 ;
      RECT  88.705 2.245 88.995 2.475 ;
      RECT  88.705 3.845 88.995 4.075 ;
      RECT  88.715 2.2 88.985 2.245 ;
      RECT  91.35 4.245 91.64 4.475 ;
      RECT  88.295 4.245 88.585 4.475 ;
      RECT  91.35 2.645 91.64 2.875 ;
      RECT  87.375 3.475 88.525 3.645 ;
      RECT  92.3 4.245 92.59 4.475 ;
      RECT  86.99 4.245 87.28 4.475 ;
      RECT  88.295 1.445 88.585 1.675 ;
      RECT  92.28 3.385 92.61 3.645 ;
      RECT  87.375 3.445 87.665 3.475 ;
      RECT  87.05 2.875 87.22 4.245 ;
      RECT  88.355 1.675 88.525 3.475 ;
      RECT  88.715 3.8 88.985 3.845 ;
      RECT  91.89 2.63 92.22 2.89 ;
      RECT  91.41 2.875 91.58 4.245 ;
      RECT  92.36 3.645 92.53 4.245 ;
      RECT  87.375 3.645 87.665 3.675 ;
      RECT  88.715 4.075 88.985 4.12 ;
      RECT  90.045 1.445 90.335 1.675 ;
      RECT  88.355 3.645 88.525 4.245 ;
      RECT  90.045 4.245 90.335 4.475 ;
      RECT  91.35 1.445 91.64 1.675 ;
      RECT  88.715 2.475 88.985 2.52 ;
      RECT  86.99 1.445 87.28 1.675 ;
      RECT  87.555 3.03 87.885 3.29 ;
      RECT  92.3 1.445 92.59 1.675 ;
      RECT  92.83 2.645 93.12 2.875 ;
      RECT  97.25 1.675 97.42 2.645 ;
      RECT  98.2 1.675 98.37 3.385 ;
      RECT  95.945 1.675 96.115 4.245 ;
      RECT  92.89 1.675 93.06 2.645 ;
      RECT  94.605 2.52 94.775 3.8 ;
      RECT  94.545 2.245 94.835 2.475 ;
      RECT  94.545 3.845 94.835 4.075 ;
      RECT  94.555 2.2 94.825 2.245 ;
      RECT  97.19 4.245 97.48 4.475 ;
      RECT  94.135 4.245 94.425 4.475 ;
      RECT  97.19 2.645 97.48 2.875 ;
      RECT  93.215 3.475 94.365 3.645 ;
      RECT  98.14 4.245 98.43 4.475 ;
      RECT  92.83 4.245 93.12 4.475 ;
      RECT  94.135 1.445 94.425 1.675 ;
      RECT  98.12 3.385 98.45 3.645 ;
      RECT  93.215 3.445 93.505 3.475 ;
      RECT  92.89 2.875 93.06 4.245 ;
      RECT  94.195 1.675 94.365 3.475 ;
      RECT  94.555 3.8 94.825 3.845 ;
      RECT  97.73 2.63 98.06 2.89 ;
      RECT  97.25 2.875 97.42 4.245 ;
      RECT  98.2 3.645 98.37 4.245 ;
      RECT  93.215 3.645 93.505 3.675 ;
      RECT  94.555 4.075 94.825 4.12 ;
      RECT  95.885 1.445 96.175 1.675 ;
      RECT  94.195 3.645 94.365 4.245 ;
      RECT  95.885 4.245 96.175 4.475 ;
      RECT  97.19 1.445 97.48 1.675 ;
      RECT  94.555 2.475 94.825 2.52 ;
      RECT  92.83 1.445 93.12 1.675 ;
      RECT  93.395 3.03 93.725 3.29 ;
      RECT  98.14 1.445 98.43 1.675 ;
      RECT  98.67 2.645 98.96 2.875 ;
      RECT  103.09 1.675 103.26 2.645 ;
      RECT  104.04 1.675 104.21 3.385 ;
      RECT  101.785 1.675 101.955 4.245 ;
      RECT  98.73 1.675 98.9 2.645 ;
      RECT  100.445 2.52 100.615 3.8 ;
      RECT  100.385 2.245 100.675 2.475 ;
      RECT  100.385 3.845 100.675 4.075 ;
      RECT  100.395 2.2 100.665 2.245 ;
      RECT  103.03 4.245 103.32 4.475 ;
      RECT  99.975 4.245 100.265 4.475 ;
      RECT  103.03 2.645 103.32 2.875 ;
      RECT  99.055 3.475 100.205 3.645 ;
      RECT  103.98 4.245 104.27 4.475 ;
      RECT  98.67 4.245 98.96 4.475 ;
      RECT  99.975 1.445 100.265 1.675 ;
      RECT  103.96 3.385 104.29 3.645 ;
      RECT  99.055 3.445 99.345 3.475 ;
      RECT  98.73 2.875 98.9 4.245 ;
      RECT  100.035 1.675 100.205 3.475 ;
      RECT  100.395 3.8 100.665 3.845 ;
      RECT  103.57 2.63 103.9 2.89 ;
      RECT  103.09 2.875 103.26 4.245 ;
      RECT  104.04 3.645 104.21 4.245 ;
      RECT  99.055 3.645 99.345 3.675 ;
      RECT  100.395 4.075 100.665 4.12 ;
      RECT  101.725 1.445 102.015 1.675 ;
      RECT  100.035 3.645 100.205 4.245 ;
      RECT  101.725 4.245 102.015 4.475 ;
      RECT  103.03 1.445 103.32 1.675 ;
      RECT  100.395 2.475 100.665 2.52 ;
      RECT  98.67 1.445 98.96 1.675 ;
      RECT  99.235 3.03 99.565 3.29 ;
      RECT  103.98 1.445 104.27 1.675 ;
      RECT  104.51 2.645 104.8 2.875 ;
      RECT  108.93 1.675 109.1 2.645 ;
      RECT  109.88 1.675 110.05 3.385 ;
      RECT  107.625 1.675 107.795 4.245 ;
      RECT  104.57 1.675 104.74 2.645 ;
      RECT  106.285 2.52 106.455 3.8 ;
      RECT  106.225 2.245 106.515 2.475 ;
      RECT  106.225 3.845 106.515 4.075 ;
      RECT  106.235 2.2 106.505 2.245 ;
      RECT  108.87 4.245 109.16 4.475 ;
      RECT  105.815 4.245 106.105 4.475 ;
      RECT  108.87 2.645 109.16 2.875 ;
      RECT  104.895 3.475 106.045 3.645 ;
      RECT  109.82 4.245 110.11 4.475 ;
      RECT  104.51 4.245 104.8 4.475 ;
      RECT  105.815 1.445 106.105 1.675 ;
      RECT  109.8 3.385 110.13 3.645 ;
      RECT  104.895 3.445 105.185 3.475 ;
      RECT  104.57 2.875 104.74 4.245 ;
      RECT  105.875 1.675 106.045 3.475 ;
      RECT  106.235 3.8 106.505 3.845 ;
      RECT  109.41 2.63 109.74 2.89 ;
      RECT  108.93 2.875 109.1 4.245 ;
      RECT  109.88 3.645 110.05 4.245 ;
      RECT  104.895 3.645 105.185 3.675 ;
      RECT  106.235 4.075 106.505 4.12 ;
      RECT  107.565 1.445 107.855 1.675 ;
      RECT  105.875 3.645 106.045 4.245 ;
      RECT  107.565 4.245 107.855 4.475 ;
      RECT  108.87 1.445 109.16 1.675 ;
      RECT  106.235 2.475 106.505 2.52 ;
      RECT  104.51 1.445 104.8 1.675 ;
      RECT  105.075 3.03 105.405 3.29 ;
      RECT  109.82 1.445 110.11 1.675 ;
      RECT  110.35 2.645 110.64 2.875 ;
      RECT  114.77 1.675 114.94 2.645 ;
      RECT  115.72 1.675 115.89 3.385 ;
      RECT  113.465 1.675 113.635 4.245 ;
      RECT  110.41 1.675 110.58 2.645 ;
      RECT  112.125 2.52 112.295 3.8 ;
      RECT  112.065 2.245 112.355 2.475 ;
      RECT  112.065 3.845 112.355 4.075 ;
      RECT  112.075 2.2 112.345 2.245 ;
      RECT  114.71 4.245 115.0 4.475 ;
      RECT  111.655 4.245 111.945 4.475 ;
      RECT  114.71 2.645 115.0 2.875 ;
      RECT  110.735 3.475 111.885 3.645 ;
      RECT  115.66 4.245 115.95 4.475 ;
      RECT  110.35 4.245 110.64 4.475 ;
      RECT  111.655 1.445 111.945 1.675 ;
      RECT  115.64 3.385 115.97 3.645 ;
      RECT  110.735 3.445 111.025 3.475 ;
      RECT  110.41 2.875 110.58 4.245 ;
      RECT  111.715 1.675 111.885 3.475 ;
      RECT  112.075 3.8 112.345 3.845 ;
      RECT  115.25 2.63 115.58 2.89 ;
      RECT  114.77 2.875 114.94 4.245 ;
      RECT  115.72 3.645 115.89 4.245 ;
      RECT  110.735 3.645 111.025 3.675 ;
      RECT  112.075 4.075 112.345 4.12 ;
      RECT  113.405 1.445 113.695 1.675 ;
      RECT  111.715 3.645 111.885 4.245 ;
      RECT  113.405 4.245 113.695 4.475 ;
      RECT  114.71 1.445 115.0 1.675 ;
      RECT  112.075 2.475 112.345 2.52 ;
      RECT  110.35 1.445 110.64 1.675 ;
      RECT  110.915 3.03 111.245 3.29 ;
      RECT  115.66 1.445 115.95 1.675 ;
      RECT  116.19 2.645 116.48 2.875 ;
      RECT  120.61 1.675 120.78 2.645 ;
      RECT  121.56 1.675 121.73 3.385 ;
      RECT  119.305 1.675 119.475 4.245 ;
      RECT  116.25 1.675 116.42 2.645 ;
      RECT  117.965 2.52 118.135 3.8 ;
      RECT  117.905 2.245 118.195 2.475 ;
      RECT  117.905 3.845 118.195 4.075 ;
      RECT  117.915 2.2 118.185 2.245 ;
      RECT  120.55 4.245 120.84 4.475 ;
      RECT  117.495 4.245 117.785 4.475 ;
      RECT  120.55 2.645 120.84 2.875 ;
      RECT  116.575 3.475 117.725 3.645 ;
      RECT  121.5 4.245 121.79 4.475 ;
      RECT  116.19 4.245 116.48 4.475 ;
      RECT  117.495 1.445 117.785 1.675 ;
      RECT  121.48 3.385 121.81 3.645 ;
      RECT  116.575 3.445 116.865 3.475 ;
      RECT  116.25 2.875 116.42 4.245 ;
      RECT  117.555 1.675 117.725 3.475 ;
      RECT  117.915 3.8 118.185 3.845 ;
      RECT  121.09 2.63 121.42 2.89 ;
      RECT  120.61 2.875 120.78 4.245 ;
      RECT  121.56 3.645 121.73 4.245 ;
      RECT  116.575 3.645 116.865 3.675 ;
      RECT  117.915 4.075 118.185 4.12 ;
      RECT  119.245 1.445 119.535 1.675 ;
      RECT  117.555 3.645 117.725 4.245 ;
      RECT  119.245 4.245 119.535 4.475 ;
      RECT  120.55 1.445 120.84 1.675 ;
      RECT  117.915 2.475 118.185 2.52 ;
      RECT  116.19 1.445 116.48 1.675 ;
      RECT  116.755 3.03 117.085 3.29 ;
      RECT  121.5 1.445 121.79 1.675 ;
      RECT  122.03 2.645 122.32 2.875 ;
      RECT  126.45 1.675 126.62 2.645 ;
      RECT  127.4 1.675 127.57 3.385 ;
      RECT  125.145 1.675 125.315 4.245 ;
      RECT  122.09 1.675 122.26 2.645 ;
      RECT  123.805 2.52 123.975 3.8 ;
      RECT  123.745 2.245 124.035 2.475 ;
      RECT  123.745 3.845 124.035 4.075 ;
      RECT  123.755 2.2 124.025 2.245 ;
      RECT  126.39 4.245 126.68 4.475 ;
      RECT  123.335 4.245 123.625 4.475 ;
      RECT  126.39 2.645 126.68 2.875 ;
      RECT  122.415 3.475 123.565 3.645 ;
      RECT  127.34 4.245 127.63 4.475 ;
      RECT  122.03 4.245 122.32 4.475 ;
      RECT  123.335 1.445 123.625 1.675 ;
      RECT  127.32 3.385 127.65 3.645 ;
      RECT  122.415 3.445 122.705 3.475 ;
      RECT  122.09 2.875 122.26 4.245 ;
      RECT  123.395 1.675 123.565 3.475 ;
      RECT  123.755 3.8 124.025 3.845 ;
      RECT  126.93 2.63 127.26 2.89 ;
      RECT  126.45 2.875 126.62 4.245 ;
      RECT  127.4 3.645 127.57 4.245 ;
      RECT  122.415 3.645 122.705 3.675 ;
      RECT  123.755 4.075 124.025 4.12 ;
      RECT  125.085 1.445 125.375 1.675 ;
      RECT  123.395 3.645 123.565 4.245 ;
      RECT  125.085 4.245 125.375 4.475 ;
      RECT  126.39 1.445 126.68 1.675 ;
      RECT  123.755 2.475 124.025 2.52 ;
      RECT  122.03 1.445 122.32 1.675 ;
      RECT  122.595 3.03 122.925 3.29 ;
      RECT  127.34 1.445 127.63 1.675 ;
      RECT  127.87 2.645 128.16 2.875 ;
      RECT  132.29 1.675 132.46 2.645 ;
      RECT  133.24 1.675 133.41 3.385 ;
      RECT  130.985 1.675 131.155 4.245 ;
      RECT  127.93 1.675 128.1 2.645 ;
      RECT  129.645 2.52 129.815 3.8 ;
      RECT  129.585 2.245 129.875 2.475 ;
      RECT  129.585 3.845 129.875 4.075 ;
      RECT  129.595 2.2 129.865 2.245 ;
      RECT  132.23 4.245 132.52 4.475 ;
      RECT  129.175 4.245 129.465 4.475 ;
      RECT  132.23 2.645 132.52 2.875 ;
      RECT  128.255 3.475 129.405 3.645 ;
      RECT  133.18 4.245 133.47 4.475 ;
      RECT  127.87 4.245 128.16 4.475 ;
      RECT  129.175 1.445 129.465 1.675 ;
      RECT  133.16 3.385 133.49 3.645 ;
      RECT  128.255 3.445 128.545 3.475 ;
      RECT  127.93 2.875 128.1 4.245 ;
      RECT  129.235 1.675 129.405 3.475 ;
      RECT  129.595 3.8 129.865 3.845 ;
      RECT  132.77 2.63 133.1 2.89 ;
      RECT  132.29 2.875 132.46 4.245 ;
      RECT  133.24 3.645 133.41 4.245 ;
      RECT  128.255 3.645 128.545 3.675 ;
      RECT  129.595 4.075 129.865 4.12 ;
      RECT  130.925 1.445 131.215 1.675 ;
      RECT  129.235 3.645 129.405 4.245 ;
      RECT  130.925 4.245 131.215 4.475 ;
      RECT  132.23 1.445 132.52 1.675 ;
      RECT  129.595 2.475 129.865 2.52 ;
      RECT  127.87 1.445 128.16 1.675 ;
      RECT  128.435 3.03 128.765 3.29 ;
      RECT  133.18 1.445 133.47 1.675 ;
      RECT  133.71 2.645 134.0 2.875 ;
      RECT  138.13 1.675 138.3 2.645 ;
      RECT  139.08 1.675 139.25 3.385 ;
      RECT  136.825 1.675 136.995 4.245 ;
      RECT  133.77 1.675 133.94 2.645 ;
      RECT  135.485 2.52 135.655 3.8 ;
      RECT  135.425 2.245 135.715 2.475 ;
      RECT  135.425 3.845 135.715 4.075 ;
      RECT  135.435 2.2 135.705 2.245 ;
      RECT  138.07 4.245 138.36 4.475 ;
      RECT  135.015 4.245 135.305 4.475 ;
      RECT  138.07 2.645 138.36 2.875 ;
      RECT  134.095 3.475 135.245 3.645 ;
      RECT  139.02 4.245 139.31 4.475 ;
      RECT  133.71 4.245 134.0 4.475 ;
      RECT  135.015 1.445 135.305 1.675 ;
      RECT  139.0 3.385 139.33 3.645 ;
      RECT  134.095 3.445 134.385 3.475 ;
      RECT  133.77 2.875 133.94 4.245 ;
      RECT  135.075 1.675 135.245 3.475 ;
      RECT  135.435 3.8 135.705 3.845 ;
      RECT  138.61 2.63 138.94 2.89 ;
      RECT  138.13 2.875 138.3 4.245 ;
      RECT  139.08 3.645 139.25 4.245 ;
      RECT  134.095 3.645 134.385 3.675 ;
      RECT  135.435 4.075 135.705 4.12 ;
      RECT  136.765 1.445 137.055 1.675 ;
      RECT  135.075 3.645 135.245 4.245 ;
      RECT  136.765 4.245 137.055 4.475 ;
      RECT  138.07 1.445 138.36 1.675 ;
      RECT  135.435 2.475 135.705 2.52 ;
      RECT  133.71 1.445 134.0 1.675 ;
      RECT  134.275 3.03 134.605 3.29 ;
      RECT  139.02 1.445 139.31 1.675 ;
      RECT  139.55 2.645 139.84 2.875 ;
      RECT  143.97 1.675 144.14 2.645 ;
      RECT  144.92 1.675 145.09 3.385 ;
      RECT  142.665 1.675 142.835 4.245 ;
      RECT  139.61 1.675 139.78 2.645 ;
      RECT  141.325 2.52 141.495 3.8 ;
      RECT  141.265 2.245 141.555 2.475 ;
      RECT  141.265 3.845 141.555 4.075 ;
      RECT  141.275 2.2 141.545 2.245 ;
      RECT  143.91 4.245 144.2 4.475 ;
      RECT  140.855 4.245 141.145 4.475 ;
      RECT  143.91 2.645 144.2 2.875 ;
      RECT  139.935 3.475 141.085 3.645 ;
      RECT  144.86 4.245 145.15 4.475 ;
      RECT  139.55 4.245 139.84 4.475 ;
      RECT  140.855 1.445 141.145 1.675 ;
      RECT  144.84 3.385 145.17 3.645 ;
      RECT  139.935 3.445 140.225 3.475 ;
      RECT  139.61 2.875 139.78 4.245 ;
      RECT  140.915 1.675 141.085 3.475 ;
      RECT  141.275 3.8 141.545 3.845 ;
      RECT  144.45 2.63 144.78 2.89 ;
      RECT  143.97 2.875 144.14 4.245 ;
      RECT  144.92 3.645 145.09 4.245 ;
      RECT  139.935 3.645 140.225 3.675 ;
      RECT  141.275 4.075 141.545 4.12 ;
      RECT  142.605 1.445 142.895 1.675 ;
      RECT  140.915 3.645 141.085 4.245 ;
      RECT  142.605 4.245 142.895 4.475 ;
      RECT  143.91 1.445 144.2 1.675 ;
      RECT  141.275 2.475 141.545 2.52 ;
      RECT  139.55 1.445 139.84 1.675 ;
      RECT  140.115 3.03 140.445 3.29 ;
      RECT  144.86 1.445 145.15 1.675 ;
      RECT  145.39 2.645 145.68 2.875 ;
      RECT  149.81 1.675 149.98 2.645 ;
      RECT  150.76 1.675 150.93 3.385 ;
      RECT  148.505 1.675 148.675 4.245 ;
      RECT  145.45 1.675 145.62 2.645 ;
      RECT  147.165 2.52 147.335 3.8 ;
      RECT  147.105 2.245 147.395 2.475 ;
      RECT  147.105 3.845 147.395 4.075 ;
      RECT  147.115 2.2 147.385 2.245 ;
      RECT  149.75 4.245 150.04 4.475 ;
      RECT  146.695 4.245 146.985 4.475 ;
      RECT  149.75 2.645 150.04 2.875 ;
      RECT  145.775 3.475 146.925 3.645 ;
      RECT  150.7 4.245 150.99 4.475 ;
      RECT  145.39 4.245 145.68 4.475 ;
      RECT  146.695 1.445 146.985 1.675 ;
      RECT  150.68 3.385 151.01 3.645 ;
      RECT  145.775 3.445 146.065 3.475 ;
      RECT  145.45 2.875 145.62 4.245 ;
      RECT  146.755 1.675 146.925 3.475 ;
      RECT  147.115 3.8 147.385 3.845 ;
      RECT  150.29 2.63 150.62 2.89 ;
      RECT  149.81 2.875 149.98 4.245 ;
      RECT  150.76 3.645 150.93 4.245 ;
      RECT  145.775 3.645 146.065 3.675 ;
      RECT  147.115 4.075 147.385 4.12 ;
      RECT  148.445 1.445 148.735 1.675 ;
      RECT  146.755 3.645 146.925 4.245 ;
      RECT  148.445 4.245 148.735 4.475 ;
      RECT  149.75 1.445 150.04 1.675 ;
      RECT  147.115 2.475 147.385 2.52 ;
      RECT  145.39 1.445 145.68 1.675 ;
      RECT  145.955 3.03 146.285 3.29 ;
      RECT  150.7 1.445 150.99 1.675 ;
   LAYER  m2 ;
      RECT  96.05 93.24 97.19 93.62 ;
      RECT  98.45 93.0 98.66 93.07 ;
      RECT  98.66 93.86 99.17 94.1 ;
      RECT  96.26 92.76 98.66 93.0 ;
      RECT  98.66 93.0 98.86 93.07 ;
      RECT  98.45 93.79 98.66 93.86 ;
      RECT  99.17 92.76 99.38 93.0 ;
      POLYGON  97.73 93.24 97.73 93.62 98.28 93.62 98.28 93.55 98.66 93.55 98.66 93.31 98.28 93.31 98.28 93.24 97.73 93.24 ;
      RECT  99.17 93.24 99.38 93.62 ;
      RECT  96.05 91.97 96.26 92.52 ;
      RECT  96.26 91.97 97.19 92.52 ;
      RECT  97.19 93.24 97.73 93.62 ;
      RECT  99.17 93.86 99.38 94.1 ;
      RECT  97.73 91.97 99.38 92.52 ;
      RECT  96.05 92.76 96.26 93.0 ;
      RECT  98.66 93.79 98.86 93.86 ;
      POLYGON  99.03 93.24 99.03 93.31 98.66 93.31 98.66 93.55 99.03 93.55 99.03 93.62 99.17 93.62 99.17 93.24 99.03 93.24 ;
      RECT  96.05 93.86 96.26 94.1 ;
      RECT  96.26 93.86 98.66 94.1 ;
      RECT  98.66 92.76 99.17 93.0 ;
      RECT  97.19 91.97 97.73 92.52 ;
      RECT  96.05 95.2 97.19 94.82 ;
      RECT  98.45 95.44 98.66 95.37 ;
      RECT  98.66 94.58 99.17 94.34 ;
      RECT  96.26 95.68 98.66 95.44 ;
      RECT  98.66 95.44 98.86 95.37 ;
      RECT  98.45 94.65 98.66 94.58 ;
      RECT  99.17 95.68 99.38 95.44 ;
      POLYGON  97.73 95.2 97.73 94.82 98.28 94.82 98.28 94.89 98.66 94.89 98.66 95.13 98.28 95.13 98.28 95.2 97.73 95.2 ;
      RECT  99.17 95.2 99.38 94.82 ;
      RECT  96.05 96.47 96.26 95.92 ;
      RECT  96.26 96.47 97.19 95.92 ;
      RECT  97.19 95.2 97.73 94.82 ;
      RECT  99.17 94.58 99.38 94.34 ;
      RECT  97.73 96.47 99.38 95.92 ;
      RECT  96.05 95.68 96.26 95.44 ;
      RECT  98.66 94.65 98.86 94.58 ;
      POLYGON  99.03 95.2 99.03 95.13 98.66 95.13 98.66 94.89 99.03 94.89 99.03 94.82 99.17 94.82 99.17 95.2 99.03 95.2 ;
      RECT  96.05 94.58 96.26 94.34 ;
      RECT  96.26 94.58 98.66 94.34 ;
      RECT  98.66 95.68 99.17 95.44 ;
      RECT  97.19 96.47 97.73 95.92 ;
      RECT  96.05 97.19 97.19 97.57 ;
      RECT  98.45 96.95 98.66 97.02 ;
      RECT  98.66 97.81 99.17 98.05 ;
      RECT  96.26 96.71 98.66 96.95 ;
      RECT  98.66 96.95 98.86 97.02 ;
      RECT  98.45 97.74 98.66 97.81 ;
      RECT  99.17 96.71 99.38 96.95 ;
      POLYGON  97.73 97.19 97.73 97.57 98.28 97.57 98.28 97.5 98.66 97.5 98.66 97.26 98.28 97.26 98.28 97.19 97.73 97.19 ;
      RECT  99.17 97.19 99.38 97.57 ;
      RECT  96.05 95.92 96.26 96.47 ;
      RECT  96.26 95.92 97.19 96.47 ;
      RECT  97.19 97.19 97.73 97.57 ;
      RECT  99.17 97.81 99.38 98.05 ;
      RECT  97.73 95.92 99.38 96.47 ;
      RECT  96.05 96.71 96.26 96.95 ;
      RECT  98.66 97.74 98.86 97.81 ;
      POLYGON  99.03 97.19 99.03 97.26 98.66 97.26 98.66 97.5 99.03 97.5 99.03 97.57 99.17 97.57 99.17 97.19 99.03 97.19 ;
      RECT  96.05 97.81 96.26 98.05 ;
      RECT  96.26 97.81 98.66 98.05 ;
      RECT  98.66 96.71 99.17 96.95 ;
      RECT  97.19 95.92 97.73 96.47 ;
      RECT  96.05 99.15 97.19 98.77 ;
      RECT  98.45 99.39 98.66 99.32 ;
      RECT  98.66 98.53 99.17 98.29 ;
      RECT  96.26 99.63 98.66 99.39 ;
      RECT  98.66 99.39 98.86 99.32 ;
      RECT  98.45 98.6 98.66 98.53 ;
      RECT  99.17 99.63 99.38 99.39 ;
      POLYGON  97.73 99.15 97.73 98.77 98.28 98.77 98.28 98.84 98.66 98.84 98.66 99.08 98.28 99.08 98.28 99.15 97.73 99.15 ;
      RECT  99.17 99.15 99.38 98.77 ;
      RECT  96.05 100.42 96.26 99.87 ;
      RECT  96.26 100.42 97.19 99.87 ;
      RECT  97.19 99.15 97.73 98.77 ;
      RECT  99.17 98.53 99.38 98.29 ;
      RECT  97.73 100.42 99.38 99.87 ;
      RECT  96.05 99.63 96.26 99.39 ;
      RECT  98.66 98.6 98.86 98.53 ;
      POLYGON  99.03 99.15 99.03 99.08 98.66 99.08 98.66 98.84 99.03 98.84 99.03 98.77 99.17 98.77 99.17 99.15 99.03 99.15 ;
      RECT  96.05 98.53 96.26 98.29 ;
      RECT  96.26 98.53 98.66 98.29 ;
      RECT  98.66 99.63 99.17 99.39 ;
      RECT  97.19 100.42 97.73 99.87 ;
      RECT  96.05 101.14 97.19 101.52 ;
      RECT  98.45 100.9 98.66 100.97 ;
      RECT  98.66 101.76 99.17 102.0 ;
      RECT  96.26 100.66 98.66 100.9 ;
      RECT  98.66 100.9 98.86 100.97 ;
      RECT  98.45 101.69 98.66 101.76 ;
      RECT  99.17 100.66 99.38 100.9 ;
      POLYGON  97.73 101.14 97.73 101.52 98.28 101.52 98.28 101.45 98.66 101.45 98.66 101.21 98.28 101.21 98.28 101.14 97.73 101.14 ;
      RECT  99.17 101.14 99.38 101.52 ;
      RECT  96.05 99.87 96.26 100.42 ;
      RECT  96.26 99.87 97.19 100.42 ;
      RECT  97.19 101.14 97.73 101.52 ;
      RECT  99.17 101.76 99.38 102.0 ;
      RECT  97.73 99.87 99.38 100.42 ;
      RECT  96.05 100.66 96.26 100.9 ;
      RECT  98.66 101.69 98.86 101.76 ;
      POLYGON  99.03 101.14 99.03 101.21 98.66 101.21 98.66 101.45 99.03 101.45 99.03 101.52 99.17 101.52 99.17 101.14 99.03 101.14 ;
      RECT  96.05 101.76 96.26 102.0 ;
      RECT  96.26 101.76 98.66 102.0 ;
      RECT  98.66 100.66 99.17 100.9 ;
      RECT  97.19 99.87 97.73 100.42 ;
      RECT  96.05 103.1 97.19 102.72 ;
      RECT  98.45 103.34 98.66 103.27 ;
      RECT  98.66 102.48 99.17 102.24 ;
      RECT  96.26 103.58 98.66 103.34 ;
      RECT  98.66 103.34 98.86 103.27 ;
      RECT  98.45 102.55 98.66 102.48 ;
      RECT  99.17 103.58 99.38 103.34 ;
      POLYGON  97.73 103.1 97.73 102.72 98.28 102.72 98.28 102.79 98.66 102.79 98.66 103.03 98.28 103.03 98.28 103.1 97.73 103.1 ;
      RECT  99.17 103.1 99.38 102.72 ;
      RECT  96.05 104.37 96.26 103.82 ;
      RECT  96.26 104.37 97.19 103.82 ;
      RECT  97.19 103.1 97.73 102.72 ;
      RECT  99.17 102.48 99.38 102.24 ;
      RECT  97.73 104.37 99.38 103.82 ;
      RECT  96.05 103.58 96.26 103.34 ;
      RECT  98.66 102.55 98.86 102.48 ;
      POLYGON  99.03 103.1 99.03 103.03 98.66 103.03 98.66 102.79 99.03 102.79 99.03 102.72 99.17 102.72 99.17 103.1 99.03 103.1 ;
      RECT  96.05 102.48 96.26 102.24 ;
      RECT  96.26 102.48 98.66 102.24 ;
      RECT  98.66 103.58 99.17 103.34 ;
      RECT  97.19 104.37 97.73 103.82 ;
      RECT  96.05 105.09 97.19 105.47 ;
      RECT  98.45 104.85 98.66 104.92 ;
      RECT  98.66 105.71 99.17 105.95 ;
      RECT  96.26 104.61 98.66 104.85 ;
      RECT  98.66 104.85 98.86 104.92 ;
      RECT  98.45 105.64 98.66 105.71 ;
      RECT  99.17 104.61 99.38 104.85 ;
      POLYGON  97.73 105.09 97.73 105.47 98.28 105.47 98.28 105.4 98.66 105.4 98.66 105.16 98.28 105.16 98.28 105.09 97.73 105.09 ;
      RECT  99.17 105.09 99.38 105.47 ;
      RECT  96.05 103.82 96.26 104.37 ;
      RECT  96.26 103.82 97.19 104.37 ;
      RECT  97.19 105.09 97.73 105.47 ;
      RECT  99.17 105.71 99.38 105.95 ;
      RECT  97.73 103.82 99.38 104.37 ;
      RECT  96.05 104.61 96.26 104.85 ;
      RECT  98.66 105.64 98.86 105.71 ;
      POLYGON  99.03 105.09 99.03 105.16 98.66 105.16 98.66 105.4 99.03 105.4 99.03 105.47 99.17 105.47 99.17 105.09 99.03 105.09 ;
      RECT  96.05 105.71 96.26 105.95 ;
      RECT  96.26 105.71 98.66 105.95 ;
      RECT  98.66 104.61 99.17 104.85 ;
      RECT  97.19 103.82 97.73 104.37 ;
      RECT  96.05 107.05 97.19 106.67 ;
      RECT  98.45 107.29 98.66 107.22 ;
      RECT  98.66 106.43 99.17 106.19 ;
      RECT  96.26 107.53 98.66 107.29 ;
      RECT  98.66 107.29 98.86 107.22 ;
      RECT  98.45 106.5 98.66 106.43 ;
      RECT  99.17 107.53 99.38 107.29 ;
      POLYGON  97.73 107.05 97.73 106.67 98.28 106.67 98.28 106.74 98.66 106.74 98.66 106.98 98.28 106.98 98.28 107.05 97.73 107.05 ;
      RECT  99.17 107.05 99.38 106.67 ;
      RECT  96.05 108.32 96.26 107.77 ;
      RECT  96.26 108.32 97.19 107.77 ;
      RECT  97.19 107.05 97.73 106.67 ;
      RECT  99.17 106.43 99.38 106.19 ;
      RECT  97.73 108.32 99.38 107.77 ;
      RECT  96.05 107.53 96.26 107.29 ;
      RECT  98.66 106.5 98.86 106.43 ;
      POLYGON  99.03 107.05 99.03 106.98 98.66 106.98 98.66 106.74 99.03 106.74 99.03 106.67 99.17 106.67 99.17 107.05 99.03 107.05 ;
      RECT  96.05 106.43 96.26 106.19 ;
      RECT  96.26 106.43 98.66 106.19 ;
      RECT  98.66 107.53 99.17 107.29 ;
      RECT  97.19 108.32 97.73 107.77 ;
      RECT  96.05 109.04 97.19 109.42 ;
      RECT  98.45 108.8 98.66 108.87 ;
      RECT  98.66 109.66 99.17 109.9 ;
      RECT  96.26 108.56 98.66 108.8 ;
      RECT  98.66 108.8 98.86 108.87 ;
      RECT  98.45 109.59 98.66 109.66 ;
      RECT  99.17 108.56 99.38 108.8 ;
      POLYGON  97.73 109.04 97.73 109.42 98.28 109.42 98.28 109.35 98.66 109.35 98.66 109.11 98.28 109.11 98.28 109.04 97.73 109.04 ;
      RECT  99.17 109.04 99.38 109.42 ;
      RECT  96.05 107.77 96.26 108.32 ;
      RECT  96.26 107.77 97.19 108.32 ;
      RECT  97.19 109.04 97.73 109.42 ;
      RECT  99.17 109.66 99.38 109.9 ;
      RECT  97.73 107.77 99.38 108.32 ;
      RECT  96.05 108.56 96.26 108.8 ;
      RECT  98.66 109.59 98.86 109.66 ;
      POLYGON  99.03 109.04 99.03 109.11 98.66 109.11 98.66 109.35 99.03 109.35 99.03 109.42 99.17 109.42 99.17 109.04 99.03 109.04 ;
      RECT  96.05 109.66 96.26 109.9 ;
      RECT  96.26 109.66 98.66 109.9 ;
      RECT  98.66 108.56 99.17 108.8 ;
      RECT  97.19 107.77 97.73 108.32 ;
      RECT  96.05 111.0 97.19 110.62 ;
      RECT  98.45 111.24 98.66 111.17 ;
      RECT  98.66 110.38 99.17 110.14 ;
      RECT  96.26 111.48 98.66 111.24 ;
      RECT  98.66 111.24 98.86 111.17 ;
      RECT  98.45 110.45 98.66 110.38 ;
      RECT  99.17 111.48 99.38 111.24 ;
      POLYGON  97.73 111.0 97.73 110.62 98.28 110.62 98.28 110.69 98.66 110.69 98.66 110.93 98.28 110.93 98.28 111.0 97.73 111.0 ;
      RECT  99.17 111.0 99.38 110.62 ;
      RECT  96.05 112.27 96.26 111.72 ;
      RECT  96.26 112.27 97.19 111.72 ;
      RECT  97.19 111.0 97.73 110.62 ;
      RECT  99.17 110.38 99.38 110.14 ;
      RECT  97.73 112.27 99.38 111.72 ;
      RECT  96.05 111.48 96.26 111.24 ;
      RECT  98.66 110.45 98.86 110.38 ;
      POLYGON  99.03 111.0 99.03 110.93 98.66 110.93 98.66 110.69 99.03 110.69 99.03 110.62 99.17 110.62 99.17 111.0 99.03 111.0 ;
      RECT  96.05 110.38 96.26 110.14 ;
      RECT  96.26 110.38 98.66 110.14 ;
      RECT  98.66 111.48 99.17 111.24 ;
      RECT  97.19 112.27 97.73 111.72 ;
      RECT  96.05 112.99 97.19 113.37 ;
      RECT  98.45 112.75 98.66 112.82 ;
      RECT  98.66 113.61 99.17 113.85 ;
      RECT  96.26 112.51 98.66 112.75 ;
      RECT  98.66 112.75 98.86 112.82 ;
      RECT  98.45 113.54 98.66 113.61 ;
      RECT  99.17 112.51 99.38 112.75 ;
      POLYGON  97.73 112.99 97.73 113.37 98.28 113.37 98.28 113.3 98.66 113.3 98.66 113.06 98.28 113.06 98.28 112.99 97.73 112.99 ;
      RECT  99.17 112.99 99.38 113.37 ;
      RECT  96.05 111.72 96.26 112.27 ;
      RECT  96.26 111.72 97.19 112.27 ;
      RECT  97.19 112.99 97.73 113.37 ;
      RECT  99.17 113.61 99.38 113.85 ;
      RECT  97.73 111.72 99.38 112.27 ;
      RECT  96.05 112.51 96.26 112.75 ;
      RECT  98.66 113.54 98.86 113.61 ;
      POLYGON  99.03 112.99 99.03 113.06 98.66 113.06 98.66 113.3 99.03 113.3 99.03 113.37 99.17 113.37 99.17 112.99 99.03 112.99 ;
      RECT  96.05 113.61 96.26 113.85 ;
      RECT  96.26 113.61 98.66 113.85 ;
      RECT  98.66 112.51 99.17 112.75 ;
      RECT  97.19 111.72 97.73 112.27 ;
      RECT  96.05 114.95 97.19 114.57 ;
      RECT  98.45 115.19 98.66 115.12 ;
      RECT  98.66 114.33 99.17 114.09 ;
      RECT  96.26 115.43 98.66 115.19 ;
      RECT  98.66 115.19 98.86 115.12 ;
      RECT  98.45 114.4 98.66 114.33 ;
      RECT  99.17 115.43 99.38 115.19 ;
      POLYGON  97.73 114.95 97.73 114.57 98.28 114.57 98.28 114.64 98.66 114.64 98.66 114.88 98.28 114.88 98.28 114.95 97.73 114.95 ;
      RECT  99.17 114.95 99.38 114.57 ;
      RECT  96.05 116.22 96.26 115.67 ;
      RECT  96.26 116.22 97.19 115.67 ;
      RECT  97.19 114.95 97.73 114.57 ;
      RECT  99.17 114.33 99.38 114.09 ;
      RECT  97.73 116.22 99.38 115.67 ;
      RECT  96.05 115.43 96.26 115.19 ;
      RECT  98.66 114.4 98.86 114.33 ;
      POLYGON  99.03 114.95 99.03 114.88 98.66 114.88 98.66 114.64 99.03 114.64 99.03 114.57 99.17 114.57 99.17 114.95 99.03 114.95 ;
      RECT  96.05 114.33 96.26 114.09 ;
      RECT  96.26 114.33 98.66 114.09 ;
      RECT  98.66 115.43 99.17 115.19 ;
      RECT  97.19 116.22 97.73 115.67 ;
      RECT  96.05 116.94 97.19 117.32 ;
      RECT  98.45 116.7 98.66 116.77 ;
      RECT  98.66 117.56 99.17 117.8 ;
      RECT  96.26 116.46 98.66 116.7 ;
      RECT  98.66 116.7 98.86 116.77 ;
      RECT  98.45 117.49 98.66 117.56 ;
      RECT  99.17 116.46 99.38 116.7 ;
      POLYGON  97.73 116.94 97.73 117.32 98.28 117.32 98.28 117.25 98.66 117.25 98.66 117.01 98.28 117.01 98.28 116.94 97.73 116.94 ;
      RECT  99.17 116.94 99.38 117.32 ;
      RECT  96.05 115.67 96.26 116.22 ;
      RECT  96.26 115.67 97.19 116.22 ;
      RECT  97.19 116.94 97.73 117.32 ;
      RECT  99.17 117.56 99.38 117.8 ;
      RECT  97.73 115.67 99.38 116.22 ;
      RECT  96.05 116.46 96.26 116.7 ;
      RECT  98.66 117.49 98.86 117.56 ;
      POLYGON  99.03 116.94 99.03 117.01 98.66 117.01 98.66 117.25 99.03 117.25 99.03 117.32 99.17 117.32 99.17 116.94 99.03 116.94 ;
      RECT  96.05 117.56 96.26 117.8 ;
      RECT  96.26 117.56 98.66 117.8 ;
      RECT  98.66 116.46 99.17 116.7 ;
      RECT  97.19 115.67 97.73 116.22 ;
      RECT  96.05 118.9 97.19 118.52 ;
      RECT  98.45 119.14 98.66 119.07 ;
      RECT  98.66 118.28 99.17 118.04 ;
      RECT  96.26 119.38 98.66 119.14 ;
      RECT  98.66 119.14 98.86 119.07 ;
      RECT  98.45 118.35 98.66 118.28 ;
      RECT  99.17 119.38 99.38 119.14 ;
      POLYGON  97.73 118.9 97.73 118.52 98.28 118.52 98.28 118.59 98.66 118.59 98.66 118.83 98.28 118.83 98.28 118.9 97.73 118.9 ;
      RECT  99.17 118.9 99.38 118.52 ;
      RECT  96.05 120.17 96.26 119.62 ;
      RECT  96.26 120.17 97.19 119.62 ;
      RECT  97.19 118.9 97.73 118.52 ;
      RECT  99.17 118.28 99.38 118.04 ;
      RECT  97.73 120.17 99.38 119.62 ;
      RECT  96.05 119.38 96.26 119.14 ;
      RECT  98.66 118.35 98.86 118.28 ;
      POLYGON  99.03 118.9 99.03 118.83 98.66 118.83 98.66 118.59 99.03 118.59 99.03 118.52 99.17 118.52 99.17 118.9 99.03 118.9 ;
      RECT  96.05 118.28 96.26 118.04 ;
      RECT  96.26 118.28 98.66 118.04 ;
      RECT  98.66 119.38 99.17 119.14 ;
      RECT  97.19 120.17 97.73 119.62 ;
      RECT  96.05 120.89 97.19 121.27 ;
      RECT  98.45 120.65 98.66 120.72 ;
      RECT  98.66 121.51 99.17 121.75 ;
      RECT  96.26 120.41 98.66 120.65 ;
      RECT  98.66 120.65 98.86 120.72 ;
      RECT  98.45 121.44 98.66 121.51 ;
      RECT  99.17 120.41 99.38 120.65 ;
      POLYGON  97.73 120.89 97.73 121.27 98.28 121.27 98.28 121.2 98.66 121.2 98.66 120.96 98.28 120.96 98.28 120.89 97.73 120.89 ;
      RECT  99.17 120.89 99.38 121.27 ;
      RECT  96.05 119.62 96.26 120.17 ;
      RECT  96.26 119.62 97.19 120.17 ;
      RECT  97.19 120.89 97.73 121.27 ;
      RECT  99.17 121.51 99.38 121.75 ;
      RECT  97.73 119.62 99.38 120.17 ;
      RECT  96.05 120.41 96.26 120.65 ;
      RECT  98.66 121.44 98.86 121.51 ;
      POLYGON  99.03 120.89 99.03 120.96 98.66 120.96 98.66 121.2 99.03 121.2 99.03 121.27 99.17 121.27 99.17 120.89 99.03 120.89 ;
      RECT  96.05 121.51 96.26 121.75 ;
      RECT  96.26 121.51 98.66 121.75 ;
      RECT  98.66 120.41 99.17 120.65 ;
      RECT  97.19 119.62 97.73 120.17 ;
      RECT  96.05 122.85 97.19 122.47 ;
      RECT  98.45 123.09 98.66 123.02 ;
      RECT  98.66 122.23 99.17 121.99 ;
      RECT  96.26 123.33 98.66 123.09 ;
      RECT  98.66 123.09 98.86 123.02 ;
      RECT  98.45 122.3 98.66 122.23 ;
      RECT  99.17 123.33 99.38 123.09 ;
      POLYGON  97.73 122.85 97.73 122.47 98.28 122.47 98.28 122.54 98.66 122.54 98.66 122.78 98.28 122.78 98.28 122.85 97.73 122.85 ;
      RECT  99.17 122.85 99.38 122.47 ;
      RECT  96.05 124.12 96.26 123.57 ;
      RECT  96.26 124.12 97.19 123.57 ;
      RECT  97.19 122.85 97.73 122.47 ;
      RECT  99.17 122.23 99.38 121.99 ;
      RECT  97.73 124.12 99.38 123.57 ;
      RECT  96.05 123.33 96.26 123.09 ;
      RECT  98.66 122.3 98.86 122.23 ;
      POLYGON  99.03 122.85 99.03 122.78 98.66 122.78 98.66 122.54 99.03 122.54 99.03 122.47 99.17 122.47 99.17 122.85 99.03 122.85 ;
      RECT  96.05 122.23 96.26 121.99 ;
      RECT  96.26 122.23 98.66 121.99 ;
      RECT  98.66 123.33 99.17 123.09 ;
      RECT  97.19 124.12 97.73 123.57 ;
      RECT  102.71 93.24 101.57 93.62 ;
      RECT  100.31 93.0 100.1 93.07 ;
      RECT  100.1 93.86 99.59 94.1 ;
      RECT  102.5 92.76 100.1 93.0 ;
      RECT  100.1 93.0 99.9 93.07 ;
      RECT  100.31 93.79 100.1 93.86 ;
      RECT  99.59 92.76 99.38 93.0 ;
      POLYGON  101.03 93.24 101.03 93.62 100.48 93.62 100.48 93.55 100.1 93.55 100.1 93.31 100.48 93.31 100.48 93.24 101.03 93.24 ;
      RECT  99.59 93.24 99.38 93.62 ;
      RECT  102.71 91.97 102.5 92.52 ;
      RECT  102.5 91.97 101.57 92.52 ;
      RECT  101.57 93.24 101.03 93.62 ;
      RECT  99.59 93.86 99.38 94.1 ;
      RECT  101.03 91.97 99.38 92.52 ;
      RECT  102.71 92.76 102.5 93.0 ;
      RECT  100.1 93.79 99.9 93.86 ;
      POLYGON  99.73 93.24 99.73 93.31 100.1 93.31 100.1 93.55 99.73 93.55 99.73 93.62 99.59 93.62 99.59 93.24 99.73 93.24 ;
      RECT  102.71 93.86 102.5 94.1 ;
      RECT  102.5 93.86 100.1 94.1 ;
      RECT  100.1 92.76 99.59 93.0 ;
      RECT  101.57 91.97 101.03 92.52 ;
      RECT  102.71 95.2 101.57 94.82 ;
      RECT  100.31 95.44 100.1 95.37 ;
      RECT  100.1 94.58 99.59 94.34 ;
      RECT  102.5 95.68 100.1 95.44 ;
      RECT  100.1 95.44 99.9 95.37 ;
      RECT  100.31 94.65 100.1 94.58 ;
      RECT  99.59 95.68 99.38 95.44 ;
      POLYGON  101.03 95.2 101.03 94.82 100.48 94.82 100.48 94.89 100.1 94.89 100.1 95.13 100.48 95.13 100.48 95.2 101.03 95.2 ;
      RECT  99.59 95.2 99.38 94.82 ;
      RECT  102.71 96.47 102.5 95.92 ;
      RECT  102.5 96.47 101.57 95.92 ;
      RECT  101.57 95.2 101.03 94.82 ;
      RECT  99.59 94.58 99.38 94.34 ;
      RECT  101.03 96.47 99.38 95.92 ;
      RECT  102.71 95.68 102.5 95.44 ;
      RECT  100.1 94.65 99.9 94.58 ;
      POLYGON  99.73 95.2 99.73 95.13 100.1 95.13 100.1 94.89 99.73 94.89 99.73 94.82 99.59 94.82 99.59 95.2 99.73 95.2 ;
      RECT  102.71 94.58 102.5 94.34 ;
      RECT  102.5 94.58 100.1 94.34 ;
      RECT  100.1 95.68 99.59 95.44 ;
      RECT  101.57 96.47 101.03 95.92 ;
      RECT  102.71 97.19 101.57 97.57 ;
      RECT  100.31 96.95 100.1 97.02 ;
      RECT  100.1 97.81 99.59 98.05 ;
      RECT  102.5 96.71 100.1 96.95 ;
      RECT  100.1 96.95 99.9 97.02 ;
      RECT  100.31 97.74 100.1 97.81 ;
      RECT  99.59 96.71 99.38 96.95 ;
      POLYGON  101.03 97.19 101.03 97.57 100.48 97.57 100.48 97.5 100.1 97.5 100.1 97.26 100.48 97.26 100.48 97.19 101.03 97.19 ;
      RECT  99.59 97.19 99.38 97.57 ;
      RECT  102.71 95.92 102.5 96.47 ;
      RECT  102.5 95.92 101.57 96.47 ;
      RECT  101.57 97.19 101.03 97.57 ;
      RECT  99.59 97.81 99.38 98.05 ;
      RECT  101.03 95.92 99.38 96.47 ;
      RECT  102.71 96.71 102.5 96.95 ;
      RECT  100.1 97.74 99.9 97.81 ;
      POLYGON  99.73 97.19 99.73 97.26 100.1 97.26 100.1 97.5 99.73 97.5 99.73 97.57 99.59 97.57 99.59 97.19 99.73 97.19 ;
      RECT  102.71 97.81 102.5 98.05 ;
      RECT  102.5 97.81 100.1 98.05 ;
      RECT  100.1 96.71 99.59 96.95 ;
      RECT  101.57 95.92 101.03 96.47 ;
      RECT  102.71 99.15 101.57 98.77 ;
      RECT  100.31 99.39 100.1 99.32 ;
      RECT  100.1 98.53 99.59 98.29 ;
      RECT  102.5 99.63 100.1 99.39 ;
      RECT  100.1 99.39 99.9 99.32 ;
      RECT  100.31 98.6 100.1 98.53 ;
      RECT  99.59 99.63 99.38 99.39 ;
      POLYGON  101.03 99.15 101.03 98.77 100.48 98.77 100.48 98.84 100.1 98.84 100.1 99.08 100.48 99.08 100.48 99.15 101.03 99.15 ;
      RECT  99.59 99.15 99.38 98.77 ;
      RECT  102.71 100.42 102.5 99.87 ;
      RECT  102.5 100.42 101.57 99.87 ;
      RECT  101.57 99.15 101.03 98.77 ;
      RECT  99.59 98.53 99.38 98.29 ;
      RECT  101.03 100.42 99.38 99.87 ;
      RECT  102.71 99.63 102.5 99.39 ;
      RECT  100.1 98.6 99.9 98.53 ;
      POLYGON  99.73 99.15 99.73 99.08 100.1 99.08 100.1 98.84 99.73 98.84 99.73 98.77 99.59 98.77 99.59 99.15 99.73 99.15 ;
      RECT  102.71 98.53 102.5 98.29 ;
      RECT  102.5 98.53 100.1 98.29 ;
      RECT  100.1 99.63 99.59 99.39 ;
      RECT  101.57 100.42 101.03 99.87 ;
      RECT  102.71 101.14 101.57 101.52 ;
      RECT  100.31 100.9 100.1 100.97 ;
      RECT  100.1 101.76 99.59 102.0 ;
      RECT  102.5 100.66 100.1 100.9 ;
      RECT  100.1 100.9 99.9 100.97 ;
      RECT  100.31 101.69 100.1 101.76 ;
      RECT  99.59 100.66 99.38 100.9 ;
      POLYGON  101.03 101.14 101.03 101.52 100.48 101.52 100.48 101.45 100.1 101.45 100.1 101.21 100.48 101.21 100.48 101.14 101.03 101.14 ;
      RECT  99.59 101.14 99.38 101.52 ;
      RECT  102.71 99.87 102.5 100.42 ;
      RECT  102.5 99.87 101.57 100.42 ;
      RECT  101.57 101.14 101.03 101.52 ;
      RECT  99.59 101.76 99.38 102.0 ;
      RECT  101.03 99.87 99.38 100.42 ;
      RECT  102.71 100.66 102.5 100.9 ;
      RECT  100.1 101.69 99.9 101.76 ;
      POLYGON  99.73 101.14 99.73 101.21 100.1 101.21 100.1 101.45 99.73 101.45 99.73 101.52 99.59 101.52 99.59 101.14 99.73 101.14 ;
      RECT  102.71 101.76 102.5 102.0 ;
      RECT  102.5 101.76 100.1 102.0 ;
      RECT  100.1 100.66 99.59 100.9 ;
      RECT  101.57 99.87 101.03 100.42 ;
      RECT  102.71 103.1 101.57 102.72 ;
      RECT  100.31 103.34 100.1 103.27 ;
      RECT  100.1 102.48 99.59 102.24 ;
      RECT  102.5 103.58 100.1 103.34 ;
      RECT  100.1 103.34 99.9 103.27 ;
      RECT  100.31 102.55 100.1 102.48 ;
      RECT  99.59 103.58 99.38 103.34 ;
      POLYGON  101.03 103.1 101.03 102.72 100.48 102.72 100.48 102.79 100.1 102.79 100.1 103.03 100.48 103.03 100.48 103.1 101.03 103.1 ;
      RECT  99.59 103.1 99.38 102.72 ;
      RECT  102.71 104.37 102.5 103.82 ;
      RECT  102.5 104.37 101.57 103.82 ;
      RECT  101.57 103.1 101.03 102.72 ;
      RECT  99.59 102.48 99.38 102.24 ;
      RECT  101.03 104.37 99.38 103.82 ;
      RECT  102.71 103.58 102.5 103.34 ;
      RECT  100.1 102.55 99.9 102.48 ;
      POLYGON  99.73 103.1 99.73 103.03 100.1 103.03 100.1 102.79 99.73 102.79 99.73 102.72 99.59 102.72 99.59 103.1 99.73 103.1 ;
      RECT  102.71 102.48 102.5 102.24 ;
      RECT  102.5 102.48 100.1 102.24 ;
      RECT  100.1 103.58 99.59 103.34 ;
      RECT  101.57 104.37 101.03 103.82 ;
      RECT  102.71 105.09 101.57 105.47 ;
      RECT  100.31 104.85 100.1 104.92 ;
      RECT  100.1 105.71 99.59 105.95 ;
      RECT  102.5 104.61 100.1 104.85 ;
      RECT  100.1 104.85 99.9 104.92 ;
      RECT  100.31 105.64 100.1 105.71 ;
      RECT  99.59 104.61 99.38 104.85 ;
      POLYGON  101.03 105.09 101.03 105.47 100.48 105.47 100.48 105.4 100.1 105.4 100.1 105.16 100.48 105.16 100.48 105.09 101.03 105.09 ;
      RECT  99.59 105.09 99.38 105.47 ;
      RECT  102.71 103.82 102.5 104.37 ;
      RECT  102.5 103.82 101.57 104.37 ;
      RECT  101.57 105.09 101.03 105.47 ;
      RECT  99.59 105.71 99.38 105.95 ;
      RECT  101.03 103.82 99.38 104.37 ;
      RECT  102.71 104.61 102.5 104.85 ;
      RECT  100.1 105.64 99.9 105.71 ;
      POLYGON  99.73 105.09 99.73 105.16 100.1 105.16 100.1 105.4 99.73 105.4 99.73 105.47 99.59 105.47 99.59 105.09 99.73 105.09 ;
      RECT  102.71 105.71 102.5 105.95 ;
      RECT  102.5 105.71 100.1 105.95 ;
      RECT  100.1 104.61 99.59 104.85 ;
      RECT  101.57 103.82 101.03 104.37 ;
      RECT  102.71 107.05 101.57 106.67 ;
      RECT  100.31 107.29 100.1 107.22 ;
      RECT  100.1 106.43 99.59 106.19 ;
      RECT  102.5 107.53 100.1 107.29 ;
      RECT  100.1 107.29 99.9 107.22 ;
      RECT  100.31 106.5 100.1 106.43 ;
      RECT  99.59 107.53 99.38 107.29 ;
      POLYGON  101.03 107.05 101.03 106.67 100.48 106.67 100.48 106.74 100.1 106.74 100.1 106.98 100.48 106.98 100.48 107.05 101.03 107.05 ;
      RECT  99.59 107.05 99.38 106.67 ;
      RECT  102.71 108.32 102.5 107.77 ;
      RECT  102.5 108.32 101.57 107.77 ;
      RECT  101.57 107.05 101.03 106.67 ;
      RECT  99.59 106.43 99.38 106.19 ;
      RECT  101.03 108.32 99.38 107.77 ;
      RECT  102.71 107.53 102.5 107.29 ;
      RECT  100.1 106.5 99.9 106.43 ;
      POLYGON  99.73 107.05 99.73 106.98 100.1 106.98 100.1 106.74 99.73 106.74 99.73 106.67 99.59 106.67 99.59 107.05 99.73 107.05 ;
      RECT  102.71 106.43 102.5 106.19 ;
      RECT  102.5 106.43 100.1 106.19 ;
      RECT  100.1 107.53 99.59 107.29 ;
      RECT  101.57 108.32 101.03 107.77 ;
      RECT  102.71 109.04 101.57 109.42 ;
      RECT  100.31 108.8 100.1 108.87 ;
      RECT  100.1 109.66 99.59 109.9 ;
      RECT  102.5 108.56 100.1 108.8 ;
      RECT  100.1 108.8 99.9 108.87 ;
      RECT  100.31 109.59 100.1 109.66 ;
      RECT  99.59 108.56 99.38 108.8 ;
      POLYGON  101.03 109.04 101.03 109.42 100.48 109.42 100.48 109.35 100.1 109.35 100.1 109.11 100.48 109.11 100.48 109.04 101.03 109.04 ;
      RECT  99.59 109.04 99.38 109.42 ;
      RECT  102.71 107.77 102.5 108.32 ;
      RECT  102.5 107.77 101.57 108.32 ;
      RECT  101.57 109.04 101.03 109.42 ;
      RECT  99.59 109.66 99.38 109.9 ;
      RECT  101.03 107.77 99.38 108.32 ;
      RECT  102.71 108.56 102.5 108.8 ;
      RECT  100.1 109.59 99.9 109.66 ;
      POLYGON  99.73 109.04 99.73 109.11 100.1 109.11 100.1 109.35 99.73 109.35 99.73 109.42 99.59 109.42 99.59 109.04 99.73 109.04 ;
      RECT  102.71 109.66 102.5 109.9 ;
      RECT  102.5 109.66 100.1 109.9 ;
      RECT  100.1 108.56 99.59 108.8 ;
      RECT  101.57 107.77 101.03 108.32 ;
      RECT  102.71 111.0 101.57 110.62 ;
      RECT  100.31 111.24 100.1 111.17 ;
      RECT  100.1 110.38 99.59 110.14 ;
      RECT  102.5 111.48 100.1 111.24 ;
      RECT  100.1 111.24 99.9 111.17 ;
      RECT  100.31 110.45 100.1 110.38 ;
      RECT  99.59 111.48 99.38 111.24 ;
      POLYGON  101.03 111.0 101.03 110.62 100.48 110.62 100.48 110.69 100.1 110.69 100.1 110.93 100.48 110.93 100.48 111.0 101.03 111.0 ;
      RECT  99.59 111.0 99.38 110.62 ;
      RECT  102.71 112.27 102.5 111.72 ;
      RECT  102.5 112.27 101.57 111.72 ;
      RECT  101.57 111.0 101.03 110.62 ;
      RECT  99.59 110.38 99.38 110.14 ;
      RECT  101.03 112.27 99.38 111.72 ;
      RECT  102.71 111.48 102.5 111.24 ;
      RECT  100.1 110.45 99.9 110.38 ;
      POLYGON  99.73 111.0 99.73 110.93 100.1 110.93 100.1 110.69 99.73 110.69 99.73 110.62 99.59 110.62 99.59 111.0 99.73 111.0 ;
      RECT  102.71 110.38 102.5 110.14 ;
      RECT  102.5 110.38 100.1 110.14 ;
      RECT  100.1 111.48 99.59 111.24 ;
      RECT  101.57 112.27 101.03 111.72 ;
      RECT  102.71 112.99 101.57 113.37 ;
      RECT  100.31 112.75 100.1 112.82 ;
      RECT  100.1 113.61 99.59 113.85 ;
      RECT  102.5 112.51 100.1 112.75 ;
      RECT  100.1 112.75 99.9 112.82 ;
      RECT  100.31 113.54 100.1 113.61 ;
      RECT  99.59 112.51 99.38 112.75 ;
      POLYGON  101.03 112.99 101.03 113.37 100.48 113.37 100.48 113.3 100.1 113.3 100.1 113.06 100.48 113.06 100.48 112.99 101.03 112.99 ;
      RECT  99.59 112.99 99.38 113.37 ;
      RECT  102.71 111.72 102.5 112.27 ;
      RECT  102.5 111.72 101.57 112.27 ;
      RECT  101.57 112.99 101.03 113.37 ;
      RECT  99.59 113.61 99.38 113.85 ;
      RECT  101.03 111.72 99.38 112.27 ;
      RECT  102.71 112.51 102.5 112.75 ;
      RECT  100.1 113.54 99.9 113.61 ;
      POLYGON  99.73 112.99 99.73 113.06 100.1 113.06 100.1 113.3 99.73 113.3 99.73 113.37 99.59 113.37 99.59 112.99 99.73 112.99 ;
      RECT  102.71 113.61 102.5 113.85 ;
      RECT  102.5 113.61 100.1 113.85 ;
      RECT  100.1 112.51 99.59 112.75 ;
      RECT  101.57 111.72 101.03 112.27 ;
      RECT  102.71 114.95 101.57 114.57 ;
      RECT  100.31 115.19 100.1 115.12 ;
      RECT  100.1 114.33 99.59 114.09 ;
      RECT  102.5 115.43 100.1 115.19 ;
      RECT  100.1 115.19 99.9 115.12 ;
      RECT  100.31 114.4 100.1 114.33 ;
      RECT  99.59 115.43 99.38 115.19 ;
      POLYGON  101.03 114.95 101.03 114.57 100.48 114.57 100.48 114.64 100.1 114.64 100.1 114.88 100.48 114.88 100.48 114.95 101.03 114.95 ;
      RECT  99.59 114.95 99.38 114.57 ;
      RECT  102.71 116.22 102.5 115.67 ;
      RECT  102.5 116.22 101.57 115.67 ;
      RECT  101.57 114.95 101.03 114.57 ;
      RECT  99.59 114.33 99.38 114.09 ;
      RECT  101.03 116.22 99.38 115.67 ;
      RECT  102.71 115.43 102.5 115.19 ;
      RECT  100.1 114.4 99.9 114.33 ;
      POLYGON  99.73 114.95 99.73 114.88 100.1 114.88 100.1 114.64 99.73 114.64 99.73 114.57 99.59 114.57 99.59 114.95 99.73 114.95 ;
      RECT  102.71 114.33 102.5 114.09 ;
      RECT  102.5 114.33 100.1 114.09 ;
      RECT  100.1 115.43 99.59 115.19 ;
      RECT  101.57 116.22 101.03 115.67 ;
      RECT  102.71 116.94 101.57 117.32 ;
      RECT  100.31 116.7 100.1 116.77 ;
      RECT  100.1 117.56 99.59 117.8 ;
      RECT  102.5 116.46 100.1 116.7 ;
      RECT  100.1 116.7 99.9 116.77 ;
      RECT  100.31 117.49 100.1 117.56 ;
      RECT  99.59 116.46 99.38 116.7 ;
      POLYGON  101.03 116.94 101.03 117.32 100.48 117.32 100.48 117.25 100.1 117.25 100.1 117.01 100.48 117.01 100.48 116.94 101.03 116.94 ;
      RECT  99.59 116.94 99.38 117.32 ;
      RECT  102.71 115.67 102.5 116.22 ;
      RECT  102.5 115.67 101.57 116.22 ;
      RECT  101.57 116.94 101.03 117.32 ;
      RECT  99.59 117.56 99.38 117.8 ;
      RECT  101.03 115.67 99.38 116.22 ;
      RECT  102.71 116.46 102.5 116.7 ;
      RECT  100.1 117.49 99.9 117.56 ;
      POLYGON  99.73 116.94 99.73 117.01 100.1 117.01 100.1 117.25 99.73 117.25 99.73 117.32 99.59 117.32 99.59 116.94 99.73 116.94 ;
      RECT  102.71 117.56 102.5 117.8 ;
      RECT  102.5 117.56 100.1 117.8 ;
      RECT  100.1 116.46 99.59 116.7 ;
      RECT  101.57 115.67 101.03 116.22 ;
      RECT  102.71 118.9 101.57 118.52 ;
      RECT  100.31 119.14 100.1 119.07 ;
      RECT  100.1 118.28 99.59 118.04 ;
      RECT  102.5 119.38 100.1 119.14 ;
      RECT  100.1 119.14 99.9 119.07 ;
      RECT  100.31 118.35 100.1 118.28 ;
      RECT  99.59 119.38 99.38 119.14 ;
      POLYGON  101.03 118.9 101.03 118.52 100.48 118.52 100.48 118.59 100.1 118.59 100.1 118.83 100.48 118.83 100.48 118.9 101.03 118.9 ;
      RECT  99.59 118.9 99.38 118.52 ;
      RECT  102.71 120.17 102.5 119.62 ;
      RECT  102.5 120.17 101.57 119.62 ;
      RECT  101.57 118.9 101.03 118.52 ;
      RECT  99.59 118.28 99.38 118.04 ;
      RECT  101.03 120.17 99.38 119.62 ;
      RECT  102.71 119.38 102.5 119.14 ;
      RECT  100.1 118.35 99.9 118.28 ;
      POLYGON  99.73 118.9 99.73 118.83 100.1 118.83 100.1 118.59 99.73 118.59 99.73 118.52 99.59 118.52 99.59 118.9 99.73 118.9 ;
      RECT  102.71 118.28 102.5 118.04 ;
      RECT  102.5 118.28 100.1 118.04 ;
      RECT  100.1 119.38 99.59 119.14 ;
      RECT  101.57 120.17 101.03 119.62 ;
      RECT  102.71 120.89 101.57 121.27 ;
      RECT  100.31 120.65 100.1 120.72 ;
      RECT  100.1 121.51 99.59 121.75 ;
      RECT  102.5 120.41 100.1 120.65 ;
      RECT  100.1 120.65 99.9 120.72 ;
      RECT  100.31 121.44 100.1 121.51 ;
      RECT  99.59 120.41 99.38 120.65 ;
      POLYGON  101.03 120.89 101.03 121.27 100.48 121.27 100.48 121.2 100.1 121.2 100.1 120.96 100.48 120.96 100.48 120.89 101.03 120.89 ;
      RECT  99.59 120.89 99.38 121.27 ;
      RECT  102.71 119.62 102.5 120.17 ;
      RECT  102.5 119.62 101.57 120.17 ;
      RECT  101.57 120.89 101.03 121.27 ;
      RECT  99.59 121.51 99.38 121.75 ;
      RECT  101.03 119.62 99.38 120.17 ;
      RECT  102.71 120.41 102.5 120.65 ;
      RECT  100.1 121.44 99.9 121.51 ;
      POLYGON  99.73 120.89 99.73 120.96 100.1 120.96 100.1 121.2 99.73 121.2 99.73 121.27 99.59 121.27 99.59 120.89 99.73 120.89 ;
      RECT  102.71 121.51 102.5 121.75 ;
      RECT  102.5 121.51 100.1 121.75 ;
      RECT  100.1 120.41 99.59 120.65 ;
      RECT  101.57 119.62 101.03 120.17 ;
      RECT  102.71 122.85 101.57 122.47 ;
      RECT  100.31 123.09 100.1 123.02 ;
      RECT  100.1 122.23 99.59 121.99 ;
      RECT  102.5 123.33 100.1 123.09 ;
      RECT  100.1 123.09 99.9 123.02 ;
      RECT  100.31 122.3 100.1 122.23 ;
      RECT  99.59 123.33 99.38 123.09 ;
      POLYGON  101.03 122.85 101.03 122.47 100.48 122.47 100.48 122.54 100.1 122.54 100.1 122.78 100.48 122.78 100.48 122.85 101.03 122.85 ;
      RECT  99.59 122.85 99.38 122.47 ;
      RECT  102.71 124.12 102.5 123.57 ;
      RECT  102.5 124.12 101.57 123.57 ;
      RECT  101.57 122.85 101.03 122.47 ;
      RECT  99.59 122.23 99.38 121.99 ;
      RECT  101.03 124.12 99.38 123.57 ;
      RECT  102.71 123.33 102.5 123.09 ;
      RECT  100.1 122.3 99.9 122.23 ;
      POLYGON  99.73 122.85 99.73 122.78 100.1 122.78 100.1 122.54 99.73 122.54 99.73 122.47 99.59 122.47 99.59 122.85 99.73 122.85 ;
      RECT  102.71 122.23 102.5 121.99 ;
      RECT  102.5 122.23 100.1 121.99 ;
      RECT  100.1 123.33 99.59 123.09 ;
      RECT  101.57 124.12 101.03 123.57 ;
      RECT  102.29 93.24 103.43 93.62 ;
      RECT  104.69 93.0 104.9 93.07 ;
      RECT  104.9 93.86 105.41 94.1 ;
      RECT  102.5 92.76 104.9 93.0 ;
      RECT  104.9 93.0 105.1 93.07 ;
      RECT  104.69 93.79 104.9 93.86 ;
      RECT  105.41 92.76 105.62 93.0 ;
      POLYGON  103.97 93.24 103.97 93.62 104.52 93.62 104.52 93.55 104.9 93.55 104.9 93.31 104.52 93.31 104.52 93.24 103.97 93.24 ;
      RECT  105.41 93.24 105.62 93.62 ;
      RECT  102.29 91.97 102.5 92.52 ;
      RECT  102.5 91.97 103.43 92.52 ;
      RECT  103.43 93.24 103.97 93.62 ;
      RECT  105.41 93.86 105.62 94.1 ;
      RECT  103.97 91.97 105.62 92.52 ;
      RECT  102.29 92.76 102.5 93.0 ;
      RECT  104.9 93.79 105.1 93.86 ;
      POLYGON  105.27 93.24 105.27 93.31 104.9 93.31 104.9 93.55 105.27 93.55 105.27 93.62 105.41 93.62 105.41 93.24 105.27 93.24 ;
      RECT  102.29 93.86 102.5 94.1 ;
      RECT  102.5 93.86 104.9 94.1 ;
      RECT  104.9 92.76 105.41 93.0 ;
      RECT  103.43 91.97 103.97 92.52 ;
      RECT  102.29 95.2 103.43 94.82 ;
      RECT  104.69 95.44 104.9 95.37 ;
      RECT  104.9 94.58 105.41 94.34 ;
      RECT  102.5 95.68 104.9 95.44 ;
      RECT  104.9 95.44 105.1 95.37 ;
      RECT  104.69 94.65 104.9 94.58 ;
      RECT  105.41 95.68 105.62 95.44 ;
      POLYGON  103.97 95.2 103.97 94.82 104.52 94.82 104.52 94.89 104.9 94.89 104.9 95.13 104.52 95.13 104.52 95.2 103.97 95.2 ;
      RECT  105.41 95.2 105.62 94.82 ;
      RECT  102.29 96.47 102.5 95.92 ;
      RECT  102.5 96.47 103.43 95.92 ;
      RECT  103.43 95.2 103.97 94.82 ;
      RECT  105.41 94.58 105.62 94.34 ;
      RECT  103.97 96.47 105.62 95.92 ;
      RECT  102.29 95.68 102.5 95.44 ;
      RECT  104.9 94.65 105.1 94.58 ;
      POLYGON  105.27 95.2 105.27 95.13 104.9 95.13 104.9 94.89 105.27 94.89 105.27 94.82 105.41 94.82 105.41 95.2 105.27 95.2 ;
      RECT  102.29 94.58 102.5 94.34 ;
      RECT  102.5 94.58 104.9 94.34 ;
      RECT  104.9 95.68 105.41 95.44 ;
      RECT  103.43 96.47 103.97 95.92 ;
      RECT  102.29 97.19 103.43 97.57 ;
      RECT  104.69 96.95 104.9 97.02 ;
      RECT  104.9 97.81 105.41 98.05 ;
      RECT  102.5 96.71 104.9 96.95 ;
      RECT  104.9 96.95 105.1 97.02 ;
      RECT  104.69 97.74 104.9 97.81 ;
      RECT  105.41 96.71 105.62 96.95 ;
      POLYGON  103.97 97.19 103.97 97.57 104.52 97.57 104.52 97.5 104.9 97.5 104.9 97.26 104.52 97.26 104.52 97.19 103.97 97.19 ;
      RECT  105.41 97.19 105.62 97.57 ;
      RECT  102.29 95.92 102.5 96.47 ;
      RECT  102.5 95.92 103.43 96.47 ;
      RECT  103.43 97.19 103.97 97.57 ;
      RECT  105.41 97.81 105.62 98.05 ;
      RECT  103.97 95.92 105.62 96.47 ;
      RECT  102.29 96.71 102.5 96.95 ;
      RECT  104.9 97.74 105.1 97.81 ;
      POLYGON  105.27 97.19 105.27 97.26 104.9 97.26 104.9 97.5 105.27 97.5 105.27 97.57 105.41 97.57 105.41 97.19 105.27 97.19 ;
      RECT  102.29 97.81 102.5 98.05 ;
      RECT  102.5 97.81 104.9 98.05 ;
      RECT  104.9 96.71 105.41 96.95 ;
      RECT  103.43 95.92 103.97 96.47 ;
      RECT  102.29 99.15 103.43 98.77 ;
      RECT  104.69 99.39 104.9 99.32 ;
      RECT  104.9 98.53 105.41 98.29 ;
      RECT  102.5 99.63 104.9 99.39 ;
      RECT  104.9 99.39 105.1 99.32 ;
      RECT  104.69 98.6 104.9 98.53 ;
      RECT  105.41 99.63 105.62 99.39 ;
      POLYGON  103.97 99.15 103.97 98.77 104.52 98.77 104.52 98.84 104.9 98.84 104.9 99.08 104.52 99.08 104.52 99.15 103.97 99.15 ;
      RECT  105.41 99.15 105.62 98.77 ;
      RECT  102.29 100.42 102.5 99.87 ;
      RECT  102.5 100.42 103.43 99.87 ;
      RECT  103.43 99.15 103.97 98.77 ;
      RECT  105.41 98.53 105.62 98.29 ;
      RECT  103.97 100.42 105.62 99.87 ;
      RECT  102.29 99.63 102.5 99.39 ;
      RECT  104.9 98.6 105.1 98.53 ;
      POLYGON  105.27 99.15 105.27 99.08 104.9 99.08 104.9 98.84 105.27 98.84 105.27 98.77 105.41 98.77 105.41 99.15 105.27 99.15 ;
      RECT  102.29 98.53 102.5 98.29 ;
      RECT  102.5 98.53 104.9 98.29 ;
      RECT  104.9 99.63 105.41 99.39 ;
      RECT  103.43 100.42 103.97 99.87 ;
      RECT  102.29 101.14 103.43 101.52 ;
      RECT  104.69 100.9 104.9 100.97 ;
      RECT  104.9 101.76 105.41 102.0 ;
      RECT  102.5 100.66 104.9 100.9 ;
      RECT  104.9 100.9 105.1 100.97 ;
      RECT  104.69 101.69 104.9 101.76 ;
      RECT  105.41 100.66 105.62 100.9 ;
      POLYGON  103.97 101.14 103.97 101.52 104.52 101.52 104.52 101.45 104.9 101.45 104.9 101.21 104.52 101.21 104.52 101.14 103.97 101.14 ;
      RECT  105.41 101.14 105.62 101.52 ;
      RECT  102.29 99.87 102.5 100.42 ;
      RECT  102.5 99.87 103.43 100.42 ;
      RECT  103.43 101.14 103.97 101.52 ;
      RECT  105.41 101.76 105.62 102.0 ;
      RECT  103.97 99.87 105.62 100.42 ;
      RECT  102.29 100.66 102.5 100.9 ;
      RECT  104.9 101.69 105.1 101.76 ;
      POLYGON  105.27 101.14 105.27 101.21 104.9 101.21 104.9 101.45 105.27 101.45 105.27 101.52 105.41 101.52 105.41 101.14 105.27 101.14 ;
      RECT  102.29 101.76 102.5 102.0 ;
      RECT  102.5 101.76 104.9 102.0 ;
      RECT  104.9 100.66 105.41 100.9 ;
      RECT  103.43 99.87 103.97 100.42 ;
      RECT  102.29 103.1 103.43 102.72 ;
      RECT  104.69 103.34 104.9 103.27 ;
      RECT  104.9 102.48 105.41 102.24 ;
      RECT  102.5 103.58 104.9 103.34 ;
      RECT  104.9 103.34 105.1 103.27 ;
      RECT  104.69 102.55 104.9 102.48 ;
      RECT  105.41 103.58 105.62 103.34 ;
      POLYGON  103.97 103.1 103.97 102.72 104.52 102.72 104.52 102.79 104.9 102.79 104.9 103.03 104.52 103.03 104.52 103.1 103.97 103.1 ;
      RECT  105.41 103.1 105.62 102.72 ;
      RECT  102.29 104.37 102.5 103.82 ;
      RECT  102.5 104.37 103.43 103.82 ;
      RECT  103.43 103.1 103.97 102.72 ;
      RECT  105.41 102.48 105.62 102.24 ;
      RECT  103.97 104.37 105.62 103.82 ;
      RECT  102.29 103.58 102.5 103.34 ;
      RECT  104.9 102.55 105.1 102.48 ;
      POLYGON  105.27 103.1 105.27 103.03 104.9 103.03 104.9 102.79 105.27 102.79 105.27 102.72 105.41 102.72 105.41 103.1 105.27 103.1 ;
      RECT  102.29 102.48 102.5 102.24 ;
      RECT  102.5 102.48 104.9 102.24 ;
      RECT  104.9 103.58 105.41 103.34 ;
      RECT  103.43 104.37 103.97 103.82 ;
      RECT  102.29 105.09 103.43 105.47 ;
      RECT  104.69 104.85 104.9 104.92 ;
      RECT  104.9 105.71 105.41 105.95 ;
      RECT  102.5 104.61 104.9 104.85 ;
      RECT  104.9 104.85 105.1 104.92 ;
      RECT  104.69 105.64 104.9 105.71 ;
      RECT  105.41 104.61 105.62 104.85 ;
      POLYGON  103.97 105.09 103.97 105.47 104.52 105.47 104.52 105.4 104.9 105.4 104.9 105.16 104.52 105.16 104.52 105.09 103.97 105.09 ;
      RECT  105.41 105.09 105.62 105.47 ;
      RECT  102.29 103.82 102.5 104.37 ;
      RECT  102.5 103.82 103.43 104.37 ;
      RECT  103.43 105.09 103.97 105.47 ;
      RECT  105.41 105.71 105.62 105.95 ;
      RECT  103.97 103.82 105.62 104.37 ;
      RECT  102.29 104.61 102.5 104.85 ;
      RECT  104.9 105.64 105.1 105.71 ;
      POLYGON  105.27 105.09 105.27 105.16 104.9 105.16 104.9 105.4 105.27 105.4 105.27 105.47 105.41 105.47 105.41 105.09 105.27 105.09 ;
      RECT  102.29 105.71 102.5 105.95 ;
      RECT  102.5 105.71 104.9 105.95 ;
      RECT  104.9 104.61 105.41 104.85 ;
      RECT  103.43 103.82 103.97 104.37 ;
      RECT  102.29 107.05 103.43 106.67 ;
      RECT  104.69 107.29 104.9 107.22 ;
      RECT  104.9 106.43 105.41 106.19 ;
      RECT  102.5 107.53 104.9 107.29 ;
      RECT  104.9 107.29 105.1 107.22 ;
      RECT  104.69 106.5 104.9 106.43 ;
      RECT  105.41 107.53 105.62 107.29 ;
      POLYGON  103.97 107.05 103.97 106.67 104.52 106.67 104.52 106.74 104.9 106.74 104.9 106.98 104.52 106.98 104.52 107.05 103.97 107.05 ;
      RECT  105.41 107.05 105.62 106.67 ;
      RECT  102.29 108.32 102.5 107.77 ;
      RECT  102.5 108.32 103.43 107.77 ;
      RECT  103.43 107.05 103.97 106.67 ;
      RECT  105.41 106.43 105.62 106.19 ;
      RECT  103.97 108.32 105.62 107.77 ;
      RECT  102.29 107.53 102.5 107.29 ;
      RECT  104.9 106.5 105.1 106.43 ;
      POLYGON  105.27 107.05 105.27 106.98 104.9 106.98 104.9 106.74 105.27 106.74 105.27 106.67 105.41 106.67 105.41 107.05 105.27 107.05 ;
      RECT  102.29 106.43 102.5 106.19 ;
      RECT  102.5 106.43 104.9 106.19 ;
      RECT  104.9 107.53 105.41 107.29 ;
      RECT  103.43 108.32 103.97 107.77 ;
      RECT  102.29 109.04 103.43 109.42 ;
      RECT  104.69 108.8 104.9 108.87 ;
      RECT  104.9 109.66 105.41 109.9 ;
      RECT  102.5 108.56 104.9 108.8 ;
      RECT  104.9 108.8 105.1 108.87 ;
      RECT  104.69 109.59 104.9 109.66 ;
      RECT  105.41 108.56 105.62 108.8 ;
      POLYGON  103.97 109.04 103.97 109.42 104.52 109.42 104.52 109.35 104.9 109.35 104.9 109.11 104.52 109.11 104.52 109.04 103.97 109.04 ;
      RECT  105.41 109.04 105.62 109.42 ;
      RECT  102.29 107.77 102.5 108.32 ;
      RECT  102.5 107.77 103.43 108.32 ;
      RECT  103.43 109.04 103.97 109.42 ;
      RECT  105.41 109.66 105.62 109.9 ;
      RECT  103.97 107.77 105.62 108.32 ;
      RECT  102.29 108.56 102.5 108.8 ;
      RECT  104.9 109.59 105.1 109.66 ;
      POLYGON  105.27 109.04 105.27 109.11 104.9 109.11 104.9 109.35 105.27 109.35 105.27 109.42 105.41 109.42 105.41 109.04 105.27 109.04 ;
      RECT  102.29 109.66 102.5 109.9 ;
      RECT  102.5 109.66 104.9 109.9 ;
      RECT  104.9 108.56 105.41 108.8 ;
      RECT  103.43 107.77 103.97 108.32 ;
      RECT  102.29 111.0 103.43 110.62 ;
      RECT  104.69 111.24 104.9 111.17 ;
      RECT  104.9 110.38 105.41 110.14 ;
      RECT  102.5 111.48 104.9 111.24 ;
      RECT  104.9 111.24 105.1 111.17 ;
      RECT  104.69 110.45 104.9 110.38 ;
      RECT  105.41 111.48 105.62 111.24 ;
      POLYGON  103.97 111.0 103.97 110.62 104.52 110.62 104.52 110.69 104.9 110.69 104.9 110.93 104.52 110.93 104.52 111.0 103.97 111.0 ;
      RECT  105.41 111.0 105.62 110.62 ;
      RECT  102.29 112.27 102.5 111.72 ;
      RECT  102.5 112.27 103.43 111.72 ;
      RECT  103.43 111.0 103.97 110.62 ;
      RECT  105.41 110.38 105.62 110.14 ;
      RECT  103.97 112.27 105.62 111.72 ;
      RECT  102.29 111.48 102.5 111.24 ;
      RECT  104.9 110.45 105.1 110.38 ;
      POLYGON  105.27 111.0 105.27 110.93 104.9 110.93 104.9 110.69 105.27 110.69 105.27 110.62 105.41 110.62 105.41 111.0 105.27 111.0 ;
      RECT  102.29 110.38 102.5 110.14 ;
      RECT  102.5 110.38 104.9 110.14 ;
      RECT  104.9 111.48 105.41 111.24 ;
      RECT  103.43 112.27 103.97 111.72 ;
      RECT  102.29 112.99 103.43 113.37 ;
      RECT  104.69 112.75 104.9 112.82 ;
      RECT  104.9 113.61 105.41 113.85 ;
      RECT  102.5 112.51 104.9 112.75 ;
      RECT  104.9 112.75 105.1 112.82 ;
      RECT  104.69 113.54 104.9 113.61 ;
      RECT  105.41 112.51 105.62 112.75 ;
      POLYGON  103.97 112.99 103.97 113.37 104.52 113.37 104.52 113.3 104.9 113.3 104.9 113.06 104.52 113.06 104.52 112.99 103.97 112.99 ;
      RECT  105.41 112.99 105.62 113.37 ;
      RECT  102.29 111.72 102.5 112.27 ;
      RECT  102.5 111.72 103.43 112.27 ;
      RECT  103.43 112.99 103.97 113.37 ;
      RECT  105.41 113.61 105.62 113.85 ;
      RECT  103.97 111.72 105.62 112.27 ;
      RECT  102.29 112.51 102.5 112.75 ;
      RECT  104.9 113.54 105.1 113.61 ;
      POLYGON  105.27 112.99 105.27 113.06 104.9 113.06 104.9 113.3 105.27 113.3 105.27 113.37 105.41 113.37 105.41 112.99 105.27 112.99 ;
      RECT  102.29 113.61 102.5 113.85 ;
      RECT  102.5 113.61 104.9 113.85 ;
      RECT  104.9 112.51 105.41 112.75 ;
      RECT  103.43 111.72 103.97 112.27 ;
      RECT  102.29 114.95 103.43 114.57 ;
      RECT  104.69 115.19 104.9 115.12 ;
      RECT  104.9 114.33 105.41 114.09 ;
      RECT  102.5 115.43 104.9 115.19 ;
      RECT  104.9 115.19 105.1 115.12 ;
      RECT  104.69 114.4 104.9 114.33 ;
      RECT  105.41 115.43 105.62 115.19 ;
      POLYGON  103.97 114.95 103.97 114.57 104.52 114.57 104.52 114.64 104.9 114.64 104.9 114.88 104.52 114.88 104.52 114.95 103.97 114.95 ;
      RECT  105.41 114.95 105.62 114.57 ;
      RECT  102.29 116.22 102.5 115.67 ;
      RECT  102.5 116.22 103.43 115.67 ;
      RECT  103.43 114.95 103.97 114.57 ;
      RECT  105.41 114.33 105.62 114.09 ;
      RECT  103.97 116.22 105.62 115.67 ;
      RECT  102.29 115.43 102.5 115.19 ;
      RECT  104.9 114.4 105.1 114.33 ;
      POLYGON  105.27 114.95 105.27 114.88 104.9 114.88 104.9 114.64 105.27 114.64 105.27 114.57 105.41 114.57 105.41 114.95 105.27 114.95 ;
      RECT  102.29 114.33 102.5 114.09 ;
      RECT  102.5 114.33 104.9 114.09 ;
      RECT  104.9 115.43 105.41 115.19 ;
      RECT  103.43 116.22 103.97 115.67 ;
      RECT  102.29 116.94 103.43 117.32 ;
      RECT  104.69 116.7 104.9 116.77 ;
      RECT  104.9 117.56 105.41 117.8 ;
      RECT  102.5 116.46 104.9 116.7 ;
      RECT  104.9 116.7 105.1 116.77 ;
      RECT  104.69 117.49 104.9 117.56 ;
      RECT  105.41 116.46 105.62 116.7 ;
      POLYGON  103.97 116.94 103.97 117.32 104.52 117.32 104.52 117.25 104.9 117.25 104.9 117.01 104.52 117.01 104.52 116.94 103.97 116.94 ;
      RECT  105.41 116.94 105.62 117.32 ;
      RECT  102.29 115.67 102.5 116.22 ;
      RECT  102.5 115.67 103.43 116.22 ;
      RECT  103.43 116.94 103.97 117.32 ;
      RECT  105.41 117.56 105.62 117.8 ;
      RECT  103.97 115.67 105.62 116.22 ;
      RECT  102.29 116.46 102.5 116.7 ;
      RECT  104.9 117.49 105.1 117.56 ;
      POLYGON  105.27 116.94 105.27 117.01 104.9 117.01 104.9 117.25 105.27 117.25 105.27 117.32 105.41 117.32 105.41 116.94 105.27 116.94 ;
      RECT  102.29 117.56 102.5 117.8 ;
      RECT  102.5 117.56 104.9 117.8 ;
      RECT  104.9 116.46 105.41 116.7 ;
      RECT  103.43 115.67 103.97 116.22 ;
      RECT  102.29 118.9 103.43 118.52 ;
      RECT  104.69 119.14 104.9 119.07 ;
      RECT  104.9 118.28 105.41 118.04 ;
      RECT  102.5 119.38 104.9 119.14 ;
      RECT  104.9 119.14 105.1 119.07 ;
      RECT  104.69 118.35 104.9 118.28 ;
      RECT  105.41 119.38 105.62 119.14 ;
      POLYGON  103.97 118.9 103.97 118.52 104.52 118.52 104.52 118.59 104.9 118.59 104.9 118.83 104.52 118.83 104.52 118.9 103.97 118.9 ;
      RECT  105.41 118.9 105.62 118.52 ;
      RECT  102.29 120.17 102.5 119.62 ;
      RECT  102.5 120.17 103.43 119.62 ;
      RECT  103.43 118.9 103.97 118.52 ;
      RECT  105.41 118.28 105.62 118.04 ;
      RECT  103.97 120.17 105.62 119.62 ;
      RECT  102.29 119.38 102.5 119.14 ;
      RECT  104.9 118.35 105.1 118.28 ;
      POLYGON  105.27 118.9 105.27 118.83 104.9 118.83 104.9 118.59 105.27 118.59 105.27 118.52 105.41 118.52 105.41 118.9 105.27 118.9 ;
      RECT  102.29 118.28 102.5 118.04 ;
      RECT  102.5 118.28 104.9 118.04 ;
      RECT  104.9 119.38 105.41 119.14 ;
      RECT  103.43 120.17 103.97 119.62 ;
      RECT  102.29 120.89 103.43 121.27 ;
      RECT  104.69 120.65 104.9 120.72 ;
      RECT  104.9 121.51 105.41 121.75 ;
      RECT  102.5 120.41 104.9 120.65 ;
      RECT  104.9 120.65 105.1 120.72 ;
      RECT  104.69 121.44 104.9 121.51 ;
      RECT  105.41 120.41 105.62 120.65 ;
      POLYGON  103.97 120.89 103.97 121.27 104.52 121.27 104.52 121.2 104.9 121.2 104.9 120.96 104.52 120.96 104.52 120.89 103.97 120.89 ;
      RECT  105.41 120.89 105.62 121.27 ;
      RECT  102.29 119.62 102.5 120.17 ;
      RECT  102.5 119.62 103.43 120.17 ;
      RECT  103.43 120.89 103.97 121.27 ;
      RECT  105.41 121.51 105.62 121.75 ;
      RECT  103.97 119.62 105.62 120.17 ;
      RECT  102.29 120.41 102.5 120.65 ;
      RECT  104.9 121.44 105.1 121.51 ;
      POLYGON  105.27 120.89 105.27 120.96 104.9 120.96 104.9 121.2 105.27 121.2 105.27 121.27 105.41 121.27 105.41 120.89 105.27 120.89 ;
      RECT  102.29 121.51 102.5 121.75 ;
      RECT  102.5 121.51 104.9 121.75 ;
      RECT  104.9 120.41 105.41 120.65 ;
      RECT  103.43 119.62 103.97 120.17 ;
      RECT  102.29 122.85 103.43 122.47 ;
      RECT  104.69 123.09 104.9 123.02 ;
      RECT  104.9 122.23 105.41 121.99 ;
      RECT  102.5 123.33 104.9 123.09 ;
      RECT  104.9 123.09 105.1 123.02 ;
      RECT  104.69 122.3 104.9 122.23 ;
      RECT  105.41 123.33 105.62 123.09 ;
      POLYGON  103.97 122.85 103.97 122.47 104.52 122.47 104.52 122.54 104.9 122.54 104.9 122.78 104.52 122.78 104.52 122.85 103.97 122.85 ;
      RECT  105.41 122.85 105.62 122.47 ;
      RECT  102.29 124.12 102.5 123.57 ;
      RECT  102.5 124.12 103.43 123.57 ;
      RECT  103.43 122.85 103.97 122.47 ;
      RECT  105.41 122.23 105.62 121.99 ;
      RECT  103.97 124.12 105.62 123.57 ;
      RECT  102.29 123.33 102.5 123.09 ;
      RECT  104.9 122.3 105.1 122.23 ;
      POLYGON  105.27 122.85 105.27 122.78 104.9 122.78 104.9 122.54 105.27 122.54 105.27 122.47 105.41 122.47 105.41 122.85 105.27 122.85 ;
      RECT  102.29 122.23 102.5 121.99 ;
      RECT  102.5 122.23 104.9 121.99 ;
      RECT  104.9 123.33 105.41 123.09 ;
      RECT  103.43 124.12 103.97 123.57 ;
      RECT  108.95 93.24 107.81 93.62 ;
      RECT  106.55 93.0 106.34 93.07 ;
      RECT  106.34 93.86 105.83 94.1 ;
      RECT  108.74 92.76 106.34 93.0 ;
      RECT  106.34 93.0 106.14 93.07 ;
      RECT  106.55 93.79 106.34 93.86 ;
      RECT  105.83 92.76 105.62 93.0 ;
      POLYGON  107.27 93.24 107.27 93.62 106.72 93.62 106.72 93.55 106.34 93.55 106.34 93.31 106.72 93.31 106.72 93.24 107.27 93.24 ;
      RECT  105.83 93.24 105.62 93.62 ;
      RECT  108.95 91.97 108.74 92.52 ;
      RECT  108.74 91.97 107.81 92.52 ;
      RECT  107.81 93.24 107.27 93.62 ;
      RECT  105.83 93.86 105.62 94.1 ;
      RECT  107.27 91.97 105.62 92.52 ;
      RECT  108.95 92.76 108.74 93.0 ;
      RECT  106.34 93.79 106.14 93.86 ;
      POLYGON  105.97 93.24 105.97 93.31 106.34 93.31 106.34 93.55 105.97 93.55 105.97 93.62 105.83 93.62 105.83 93.24 105.97 93.24 ;
      RECT  108.95 93.86 108.74 94.1 ;
      RECT  108.74 93.86 106.34 94.1 ;
      RECT  106.34 92.76 105.83 93.0 ;
      RECT  107.81 91.97 107.27 92.52 ;
      RECT  108.95 95.2 107.81 94.82 ;
      RECT  106.55 95.44 106.34 95.37 ;
      RECT  106.34 94.58 105.83 94.34 ;
      RECT  108.74 95.68 106.34 95.44 ;
      RECT  106.34 95.44 106.14 95.37 ;
      RECT  106.55 94.65 106.34 94.58 ;
      RECT  105.83 95.68 105.62 95.44 ;
      POLYGON  107.27 95.2 107.27 94.82 106.72 94.82 106.72 94.89 106.34 94.89 106.34 95.13 106.72 95.13 106.72 95.2 107.27 95.2 ;
      RECT  105.83 95.2 105.62 94.82 ;
      RECT  108.95 96.47 108.74 95.92 ;
      RECT  108.74 96.47 107.81 95.92 ;
      RECT  107.81 95.2 107.27 94.82 ;
      RECT  105.83 94.58 105.62 94.34 ;
      RECT  107.27 96.47 105.62 95.92 ;
      RECT  108.95 95.68 108.74 95.44 ;
      RECT  106.34 94.65 106.14 94.58 ;
      POLYGON  105.97 95.2 105.97 95.13 106.34 95.13 106.34 94.89 105.97 94.89 105.97 94.82 105.83 94.82 105.83 95.2 105.97 95.2 ;
      RECT  108.95 94.58 108.74 94.34 ;
      RECT  108.74 94.58 106.34 94.34 ;
      RECT  106.34 95.68 105.83 95.44 ;
      RECT  107.81 96.47 107.27 95.92 ;
      RECT  108.95 97.19 107.81 97.57 ;
      RECT  106.55 96.95 106.34 97.02 ;
      RECT  106.34 97.81 105.83 98.05 ;
      RECT  108.74 96.71 106.34 96.95 ;
      RECT  106.34 96.95 106.14 97.02 ;
      RECT  106.55 97.74 106.34 97.81 ;
      RECT  105.83 96.71 105.62 96.95 ;
      POLYGON  107.27 97.19 107.27 97.57 106.72 97.57 106.72 97.5 106.34 97.5 106.34 97.26 106.72 97.26 106.72 97.19 107.27 97.19 ;
      RECT  105.83 97.19 105.62 97.57 ;
      RECT  108.95 95.92 108.74 96.47 ;
      RECT  108.74 95.92 107.81 96.47 ;
      RECT  107.81 97.19 107.27 97.57 ;
      RECT  105.83 97.81 105.62 98.05 ;
      RECT  107.27 95.92 105.62 96.47 ;
      RECT  108.95 96.71 108.74 96.95 ;
      RECT  106.34 97.74 106.14 97.81 ;
      POLYGON  105.97 97.19 105.97 97.26 106.34 97.26 106.34 97.5 105.97 97.5 105.97 97.57 105.83 97.57 105.83 97.19 105.97 97.19 ;
      RECT  108.95 97.81 108.74 98.05 ;
      RECT  108.74 97.81 106.34 98.05 ;
      RECT  106.34 96.71 105.83 96.95 ;
      RECT  107.81 95.92 107.27 96.47 ;
      RECT  108.95 99.15 107.81 98.77 ;
      RECT  106.55 99.39 106.34 99.32 ;
      RECT  106.34 98.53 105.83 98.29 ;
      RECT  108.74 99.63 106.34 99.39 ;
      RECT  106.34 99.39 106.14 99.32 ;
      RECT  106.55 98.6 106.34 98.53 ;
      RECT  105.83 99.63 105.62 99.39 ;
      POLYGON  107.27 99.15 107.27 98.77 106.72 98.77 106.72 98.84 106.34 98.84 106.34 99.08 106.72 99.08 106.72 99.15 107.27 99.15 ;
      RECT  105.83 99.15 105.62 98.77 ;
      RECT  108.95 100.42 108.74 99.87 ;
      RECT  108.74 100.42 107.81 99.87 ;
      RECT  107.81 99.15 107.27 98.77 ;
      RECT  105.83 98.53 105.62 98.29 ;
      RECT  107.27 100.42 105.62 99.87 ;
      RECT  108.95 99.63 108.74 99.39 ;
      RECT  106.34 98.6 106.14 98.53 ;
      POLYGON  105.97 99.15 105.97 99.08 106.34 99.08 106.34 98.84 105.97 98.84 105.97 98.77 105.83 98.77 105.83 99.15 105.97 99.15 ;
      RECT  108.95 98.53 108.74 98.29 ;
      RECT  108.74 98.53 106.34 98.29 ;
      RECT  106.34 99.63 105.83 99.39 ;
      RECT  107.81 100.42 107.27 99.87 ;
      RECT  108.95 101.14 107.81 101.52 ;
      RECT  106.55 100.9 106.34 100.97 ;
      RECT  106.34 101.76 105.83 102.0 ;
      RECT  108.74 100.66 106.34 100.9 ;
      RECT  106.34 100.9 106.14 100.97 ;
      RECT  106.55 101.69 106.34 101.76 ;
      RECT  105.83 100.66 105.62 100.9 ;
      POLYGON  107.27 101.14 107.27 101.52 106.72 101.52 106.72 101.45 106.34 101.45 106.34 101.21 106.72 101.21 106.72 101.14 107.27 101.14 ;
      RECT  105.83 101.14 105.62 101.52 ;
      RECT  108.95 99.87 108.74 100.42 ;
      RECT  108.74 99.87 107.81 100.42 ;
      RECT  107.81 101.14 107.27 101.52 ;
      RECT  105.83 101.76 105.62 102.0 ;
      RECT  107.27 99.87 105.62 100.42 ;
      RECT  108.95 100.66 108.74 100.9 ;
      RECT  106.34 101.69 106.14 101.76 ;
      POLYGON  105.97 101.14 105.97 101.21 106.34 101.21 106.34 101.45 105.97 101.45 105.97 101.52 105.83 101.52 105.83 101.14 105.97 101.14 ;
      RECT  108.95 101.76 108.74 102.0 ;
      RECT  108.74 101.76 106.34 102.0 ;
      RECT  106.34 100.66 105.83 100.9 ;
      RECT  107.81 99.87 107.27 100.42 ;
      RECT  108.95 103.1 107.81 102.72 ;
      RECT  106.55 103.34 106.34 103.27 ;
      RECT  106.34 102.48 105.83 102.24 ;
      RECT  108.74 103.58 106.34 103.34 ;
      RECT  106.34 103.34 106.14 103.27 ;
      RECT  106.55 102.55 106.34 102.48 ;
      RECT  105.83 103.58 105.62 103.34 ;
      POLYGON  107.27 103.1 107.27 102.72 106.72 102.72 106.72 102.79 106.34 102.79 106.34 103.03 106.72 103.03 106.72 103.1 107.27 103.1 ;
      RECT  105.83 103.1 105.62 102.72 ;
      RECT  108.95 104.37 108.74 103.82 ;
      RECT  108.74 104.37 107.81 103.82 ;
      RECT  107.81 103.1 107.27 102.72 ;
      RECT  105.83 102.48 105.62 102.24 ;
      RECT  107.27 104.37 105.62 103.82 ;
      RECT  108.95 103.58 108.74 103.34 ;
      RECT  106.34 102.55 106.14 102.48 ;
      POLYGON  105.97 103.1 105.97 103.03 106.34 103.03 106.34 102.79 105.97 102.79 105.97 102.72 105.83 102.72 105.83 103.1 105.97 103.1 ;
      RECT  108.95 102.48 108.74 102.24 ;
      RECT  108.74 102.48 106.34 102.24 ;
      RECT  106.34 103.58 105.83 103.34 ;
      RECT  107.81 104.37 107.27 103.82 ;
      RECT  108.95 105.09 107.81 105.47 ;
      RECT  106.55 104.85 106.34 104.92 ;
      RECT  106.34 105.71 105.83 105.95 ;
      RECT  108.74 104.61 106.34 104.85 ;
      RECT  106.34 104.85 106.14 104.92 ;
      RECT  106.55 105.64 106.34 105.71 ;
      RECT  105.83 104.61 105.62 104.85 ;
      POLYGON  107.27 105.09 107.27 105.47 106.72 105.47 106.72 105.4 106.34 105.4 106.34 105.16 106.72 105.16 106.72 105.09 107.27 105.09 ;
      RECT  105.83 105.09 105.62 105.47 ;
      RECT  108.95 103.82 108.74 104.37 ;
      RECT  108.74 103.82 107.81 104.37 ;
      RECT  107.81 105.09 107.27 105.47 ;
      RECT  105.83 105.71 105.62 105.95 ;
      RECT  107.27 103.82 105.62 104.37 ;
      RECT  108.95 104.61 108.74 104.85 ;
      RECT  106.34 105.64 106.14 105.71 ;
      POLYGON  105.97 105.09 105.97 105.16 106.34 105.16 106.34 105.4 105.97 105.4 105.97 105.47 105.83 105.47 105.83 105.09 105.97 105.09 ;
      RECT  108.95 105.71 108.74 105.95 ;
      RECT  108.74 105.71 106.34 105.95 ;
      RECT  106.34 104.61 105.83 104.85 ;
      RECT  107.81 103.82 107.27 104.37 ;
      RECT  108.95 107.05 107.81 106.67 ;
      RECT  106.55 107.29 106.34 107.22 ;
      RECT  106.34 106.43 105.83 106.19 ;
      RECT  108.74 107.53 106.34 107.29 ;
      RECT  106.34 107.29 106.14 107.22 ;
      RECT  106.55 106.5 106.34 106.43 ;
      RECT  105.83 107.53 105.62 107.29 ;
      POLYGON  107.27 107.05 107.27 106.67 106.72 106.67 106.72 106.74 106.34 106.74 106.34 106.98 106.72 106.98 106.72 107.05 107.27 107.05 ;
      RECT  105.83 107.05 105.62 106.67 ;
      RECT  108.95 108.32 108.74 107.77 ;
      RECT  108.74 108.32 107.81 107.77 ;
      RECT  107.81 107.05 107.27 106.67 ;
      RECT  105.83 106.43 105.62 106.19 ;
      RECT  107.27 108.32 105.62 107.77 ;
      RECT  108.95 107.53 108.74 107.29 ;
      RECT  106.34 106.5 106.14 106.43 ;
      POLYGON  105.97 107.05 105.97 106.98 106.34 106.98 106.34 106.74 105.97 106.74 105.97 106.67 105.83 106.67 105.83 107.05 105.97 107.05 ;
      RECT  108.95 106.43 108.74 106.19 ;
      RECT  108.74 106.43 106.34 106.19 ;
      RECT  106.34 107.53 105.83 107.29 ;
      RECT  107.81 108.32 107.27 107.77 ;
      RECT  108.95 109.04 107.81 109.42 ;
      RECT  106.55 108.8 106.34 108.87 ;
      RECT  106.34 109.66 105.83 109.9 ;
      RECT  108.74 108.56 106.34 108.8 ;
      RECT  106.34 108.8 106.14 108.87 ;
      RECT  106.55 109.59 106.34 109.66 ;
      RECT  105.83 108.56 105.62 108.8 ;
      POLYGON  107.27 109.04 107.27 109.42 106.72 109.42 106.72 109.35 106.34 109.35 106.34 109.11 106.72 109.11 106.72 109.04 107.27 109.04 ;
      RECT  105.83 109.04 105.62 109.42 ;
      RECT  108.95 107.77 108.74 108.32 ;
      RECT  108.74 107.77 107.81 108.32 ;
      RECT  107.81 109.04 107.27 109.42 ;
      RECT  105.83 109.66 105.62 109.9 ;
      RECT  107.27 107.77 105.62 108.32 ;
      RECT  108.95 108.56 108.74 108.8 ;
      RECT  106.34 109.59 106.14 109.66 ;
      POLYGON  105.97 109.04 105.97 109.11 106.34 109.11 106.34 109.35 105.97 109.35 105.97 109.42 105.83 109.42 105.83 109.04 105.97 109.04 ;
      RECT  108.95 109.66 108.74 109.9 ;
      RECT  108.74 109.66 106.34 109.9 ;
      RECT  106.34 108.56 105.83 108.8 ;
      RECT  107.81 107.77 107.27 108.32 ;
      RECT  108.95 111.0 107.81 110.62 ;
      RECT  106.55 111.24 106.34 111.17 ;
      RECT  106.34 110.38 105.83 110.14 ;
      RECT  108.74 111.48 106.34 111.24 ;
      RECT  106.34 111.24 106.14 111.17 ;
      RECT  106.55 110.45 106.34 110.38 ;
      RECT  105.83 111.48 105.62 111.24 ;
      POLYGON  107.27 111.0 107.27 110.62 106.72 110.62 106.72 110.69 106.34 110.69 106.34 110.93 106.72 110.93 106.72 111.0 107.27 111.0 ;
      RECT  105.83 111.0 105.62 110.62 ;
      RECT  108.95 112.27 108.74 111.72 ;
      RECT  108.74 112.27 107.81 111.72 ;
      RECT  107.81 111.0 107.27 110.62 ;
      RECT  105.83 110.38 105.62 110.14 ;
      RECT  107.27 112.27 105.62 111.72 ;
      RECT  108.95 111.48 108.74 111.24 ;
      RECT  106.34 110.45 106.14 110.38 ;
      POLYGON  105.97 111.0 105.97 110.93 106.34 110.93 106.34 110.69 105.97 110.69 105.97 110.62 105.83 110.62 105.83 111.0 105.97 111.0 ;
      RECT  108.95 110.38 108.74 110.14 ;
      RECT  108.74 110.38 106.34 110.14 ;
      RECT  106.34 111.48 105.83 111.24 ;
      RECT  107.81 112.27 107.27 111.72 ;
      RECT  108.95 112.99 107.81 113.37 ;
      RECT  106.55 112.75 106.34 112.82 ;
      RECT  106.34 113.61 105.83 113.85 ;
      RECT  108.74 112.51 106.34 112.75 ;
      RECT  106.34 112.75 106.14 112.82 ;
      RECT  106.55 113.54 106.34 113.61 ;
      RECT  105.83 112.51 105.62 112.75 ;
      POLYGON  107.27 112.99 107.27 113.37 106.72 113.37 106.72 113.3 106.34 113.3 106.34 113.06 106.72 113.06 106.72 112.99 107.27 112.99 ;
      RECT  105.83 112.99 105.62 113.37 ;
      RECT  108.95 111.72 108.74 112.27 ;
      RECT  108.74 111.72 107.81 112.27 ;
      RECT  107.81 112.99 107.27 113.37 ;
      RECT  105.83 113.61 105.62 113.85 ;
      RECT  107.27 111.72 105.62 112.27 ;
      RECT  108.95 112.51 108.74 112.75 ;
      RECT  106.34 113.54 106.14 113.61 ;
      POLYGON  105.97 112.99 105.97 113.06 106.34 113.06 106.34 113.3 105.97 113.3 105.97 113.37 105.83 113.37 105.83 112.99 105.97 112.99 ;
      RECT  108.95 113.61 108.74 113.85 ;
      RECT  108.74 113.61 106.34 113.85 ;
      RECT  106.34 112.51 105.83 112.75 ;
      RECT  107.81 111.72 107.27 112.27 ;
      RECT  108.95 114.95 107.81 114.57 ;
      RECT  106.55 115.19 106.34 115.12 ;
      RECT  106.34 114.33 105.83 114.09 ;
      RECT  108.74 115.43 106.34 115.19 ;
      RECT  106.34 115.19 106.14 115.12 ;
      RECT  106.55 114.4 106.34 114.33 ;
      RECT  105.83 115.43 105.62 115.19 ;
      POLYGON  107.27 114.95 107.27 114.57 106.72 114.57 106.72 114.64 106.34 114.64 106.34 114.88 106.72 114.88 106.72 114.95 107.27 114.95 ;
      RECT  105.83 114.95 105.62 114.57 ;
      RECT  108.95 116.22 108.74 115.67 ;
      RECT  108.74 116.22 107.81 115.67 ;
      RECT  107.81 114.95 107.27 114.57 ;
      RECT  105.83 114.33 105.62 114.09 ;
      RECT  107.27 116.22 105.62 115.67 ;
      RECT  108.95 115.43 108.74 115.19 ;
      RECT  106.34 114.4 106.14 114.33 ;
      POLYGON  105.97 114.95 105.97 114.88 106.34 114.88 106.34 114.64 105.97 114.64 105.97 114.57 105.83 114.57 105.83 114.95 105.97 114.95 ;
      RECT  108.95 114.33 108.74 114.09 ;
      RECT  108.74 114.33 106.34 114.09 ;
      RECT  106.34 115.43 105.83 115.19 ;
      RECT  107.81 116.22 107.27 115.67 ;
      RECT  108.95 116.94 107.81 117.32 ;
      RECT  106.55 116.7 106.34 116.77 ;
      RECT  106.34 117.56 105.83 117.8 ;
      RECT  108.74 116.46 106.34 116.7 ;
      RECT  106.34 116.7 106.14 116.77 ;
      RECT  106.55 117.49 106.34 117.56 ;
      RECT  105.83 116.46 105.62 116.7 ;
      POLYGON  107.27 116.94 107.27 117.32 106.72 117.32 106.72 117.25 106.34 117.25 106.34 117.01 106.72 117.01 106.72 116.94 107.27 116.94 ;
      RECT  105.83 116.94 105.62 117.32 ;
      RECT  108.95 115.67 108.74 116.22 ;
      RECT  108.74 115.67 107.81 116.22 ;
      RECT  107.81 116.94 107.27 117.32 ;
      RECT  105.83 117.56 105.62 117.8 ;
      RECT  107.27 115.67 105.62 116.22 ;
      RECT  108.95 116.46 108.74 116.7 ;
      RECT  106.34 117.49 106.14 117.56 ;
      POLYGON  105.97 116.94 105.97 117.01 106.34 117.01 106.34 117.25 105.97 117.25 105.97 117.32 105.83 117.32 105.83 116.94 105.97 116.94 ;
      RECT  108.95 117.56 108.74 117.8 ;
      RECT  108.74 117.56 106.34 117.8 ;
      RECT  106.34 116.46 105.83 116.7 ;
      RECT  107.81 115.67 107.27 116.22 ;
      RECT  108.95 118.9 107.81 118.52 ;
      RECT  106.55 119.14 106.34 119.07 ;
      RECT  106.34 118.28 105.83 118.04 ;
      RECT  108.74 119.38 106.34 119.14 ;
      RECT  106.34 119.14 106.14 119.07 ;
      RECT  106.55 118.35 106.34 118.28 ;
      RECT  105.83 119.38 105.62 119.14 ;
      POLYGON  107.27 118.9 107.27 118.52 106.72 118.52 106.72 118.59 106.34 118.59 106.34 118.83 106.72 118.83 106.72 118.9 107.27 118.9 ;
      RECT  105.83 118.9 105.62 118.52 ;
      RECT  108.95 120.17 108.74 119.62 ;
      RECT  108.74 120.17 107.81 119.62 ;
      RECT  107.81 118.9 107.27 118.52 ;
      RECT  105.83 118.28 105.62 118.04 ;
      RECT  107.27 120.17 105.62 119.62 ;
      RECT  108.95 119.38 108.74 119.14 ;
      RECT  106.34 118.35 106.14 118.28 ;
      POLYGON  105.97 118.9 105.97 118.83 106.34 118.83 106.34 118.59 105.97 118.59 105.97 118.52 105.83 118.52 105.83 118.9 105.97 118.9 ;
      RECT  108.95 118.28 108.74 118.04 ;
      RECT  108.74 118.28 106.34 118.04 ;
      RECT  106.34 119.38 105.83 119.14 ;
      RECT  107.81 120.17 107.27 119.62 ;
      RECT  108.95 120.89 107.81 121.27 ;
      RECT  106.55 120.65 106.34 120.72 ;
      RECT  106.34 121.51 105.83 121.75 ;
      RECT  108.74 120.41 106.34 120.65 ;
      RECT  106.34 120.65 106.14 120.72 ;
      RECT  106.55 121.44 106.34 121.51 ;
      RECT  105.83 120.41 105.62 120.65 ;
      POLYGON  107.27 120.89 107.27 121.27 106.72 121.27 106.72 121.2 106.34 121.2 106.34 120.96 106.72 120.96 106.72 120.89 107.27 120.89 ;
      RECT  105.83 120.89 105.62 121.27 ;
      RECT  108.95 119.62 108.74 120.17 ;
      RECT  108.74 119.62 107.81 120.17 ;
      RECT  107.81 120.89 107.27 121.27 ;
      RECT  105.83 121.51 105.62 121.75 ;
      RECT  107.27 119.62 105.62 120.17 ;
      RECT  108.95 120.41 108.74 120.65 ;
      RECT  106.34 121.44 106.14 121.51 ;
      POLYGON  105.97 120.89 105.97 120.96 106.34 120.96 106.34 121.2 105.97 121.2 105.97 121.27 105.83 121.27 105.83 120.89 105.97 120.89 ;
      RECT  108.95 121.51 108.74 121.75 ;
      RECT  108.74 121.51 106.34 121.75 ;
      RECT  106.34 120.41 105.83 120.65 ;
      RECT  107.81 119.62 107.27 120.17 ;
      RECT  108.95 122.85 107.81 122.47 ;
      RECT  106.55 123.09 106.34 123.02 ;
      RECT  106.34 122.23 105.83 121.99 ;
      RECT  108.74 123.33 106.34 123.09 ;
      RECT  106.34 123.09 106.14 123.02 ;
      RECT  106.55 122.3 106.34 122.23 ;
      RECT  105.83 123.33 105.62 123.09 ;
      POLYGON  107.27 122.85 107.27 122.47 106.72 122.47 106.72 122.54 106.34 122.54 106.34 122.78 106.72 122.78 106.72 122.85 107.27 122.85 ;
      RECT  105.83 122.85 105.62 122.47 ;
      RECT  108.95 124.12 108.74 123.57 ;
      RECT  108.74 124.12 107.81 123.57 ;
      RECT  107.81 122.85 107.27 122.47 ;
      RECT  105.83 122.23 105.62 121.99 ;
      RECT  107.27 124.12 105.62 123.57 ;
      RECT  108.95 123.33 108.74 123.09 ;
      RECT  106.34 122.3 106.14 122.23 ;
      POLYGON  105.97 122.85 105.97 122.78 106.34 122.78 106.34 122.54 105.97 122.54 105.97 122.47 105.83 122.47 105.83 122.85 105.97 122.85 ;
      RECT  108.95 122.23 108.74 121.99 ;
      RECT  108.74 122.23 106.34 121.99 ;
      RECT  106.34 123.33 105.83 123.09 ;
      RECT  107.81 124.12 107.27 123.57 ;
      RECT  108.53 93.24 109.67 93.62 ;
      RECT  110.93 93.0 111.14 93.07 ;
      RECT  111.14 93.86 111.65 94.1 ;
      RECT  108.74 92.76 111.14 93.0 ;
      RECT  111.14 93.0 111.34 93.07 ;
      RECT  110.93 93.79 111.14 93.86 ;
      RECT  111.65 92.76 111.86 93.0 ;
      POLYGON  110.21 93.24 110.21 93.62 110.76 93.62 110.76 93.55 111.14 93.55 111.14 93.31 110.76 93.31 110.76 93.24 110.21 93.24 ;
      RECT  111.65 93.24 111.86 93.62 ;
      RECT  108.53 91.97 108.74 92.52 ;
      RECT  108.74 91.97 109.67 92.52 ;
      RECT  109.67 93.24 110.21 93.62 ;
      RECT  111.65 93.86 111.86 94.1 ;
      RECT  110.21 91.97 111.86 92.52 ;
      RECT  108.53 92.76 108.74 93.0 ;
      RECT  111.14 93.79 111.34 93.86 ;
      POLYGON  111.51 93.24 111.51 93.31 111.14 93.31 111.14 93.55 111.51 93.55 111.51 93.62 111.65 93.62 111.65 93.24 111.51 93.24 ;
      RECT  108.53 93.86 108.74 94.1 ;
      RECT  108.74 93.86 111.14 94.1 ;
      RECT  111.14 92.76 111.65 93.0 ;
      RECT  109.67 91.97 110.21 92.52 ;
      RECT  108.53 95.2 109.67 94.82 ;
      RECT  110.93 95.44 111.14 95.37 ;
      RECT  111.14 94.58 111.65 94.34 ;
      RECT  108.74 95.68 111.14 95.44 ;
      RECT  111.14 95.44 111.34 95.37 ;
      RECT  110.93 94.65 111.14 94.58 ;
      RECT  111.65 95.68 111.86 95.44 ;
      POLYGON  110.21 95.2 110.21 94.82 110.76 94.82 110.76 94.89 111.14 94.89 111.14 95.13 110.76 95.13 110.76 95.2 110.21 95.2 ;
      RECT  111.65 95.2 111.86 94.82 ;
      RECT  108.53 96.47 108.74 95.92 ;
      RECT  108.74 96.47 109.67 95.92 ;
      RECT  109.67 95.2 110.21 94.82 ;
      RECT  111.65 94.58 111.86 94.34 ;
      RECT  110.21 96.47 111.86 95.92 ;
      RECT  108.53 95.68 108.74 95.44 ;
      RECT  111.14 94.65 111.34 94.58 ;
      POLYGON  111.51 95.2 111.51 95.13 111.14 95.13 111.14 94.89 111.51 94.89 111.51 94.82 111.65 94.82 111.65 95.2 111.51 95.2 ;
      RECT  108.53 94.58 108.74 94.34 ;
      RECT  108.74 94.58 111.14 94.34 ;
      RECT  111.14 95.68 111.65 95.44 ;
      RECT  109.67 96.47 110.21 95.92 ;
      RECT  108.53 97.19 109.67 97.57 ;
      RECT  110.93 96.95 111.14 97.02 ;
      RECT  111.14 97.81 111.65 98.05 ;
      RECT  108.74 96.71 111.14 96.95 ;
      RECT  111.14 96.95 111.34 97.02 ;
      RECT  110.93 97.74 111.14 97.81 ;
      RECT  111.65 96.71 111.86 96.95 ;
      POLYGON  110.21 97.19 110.21 97.57 110.76 97.57 110.76 97.5 111.14 97.5 111.14 97.26 110.76 97.26 110.76 97.19 110.21 97.19 ;
      RECT  111.65 97.19 111.86 97.57 ;
      RECT  108.53 95.92 108.74 96.47 ;
      RECT  108.74 95.92 109.67 96.47 ;
      RECT  109.67 97.19 110.21 97.57 ;
      RECT  111.65 97.81 111.86 98.05 ;
      RECT  110.21 95.92 111.86 96.47 ;
      RECT  108.53 96.71 108.74 96.95 ;
      RECT  111.14 97.74 111.34 97.81 ;
      POLYGON  111.51 97.19 111.51 97.26 111.14 97.26 111.14 97.5 111.51 97.5 111.51 97.57 111.65 97.57 111.65 97.19 111.51 97.19 ;
      RECT  108.53 97.81 108.74 98.05 ;
      RECT  108.74 97.81 111.14 98.05 ;
      RECT  111.14 96.71 111.65 96.95 ;
      RECT  109.67 95.92 110.21 96.47 ;
      RECT  108.53 99.15 109.67 98.77 ;
      RECT  110.93 99.39 111.14 99.32 ;
      RECT  111.14 98.53 111.65 98.29 ;
      RECT  108.74 99.63 111.14 99.39 ;
      RECT  111.14 99.39 111.34 99.32 ;
      RECT  110.93 98.6 111.14 98.53 ;
      RECT  111.65 99.63 111.86 99.39 ;
      POLYGON  110.21 99.15 110.21 98.77 110.76 98.77 110.76 98.84 111.14 98.84 111.14 99.08 110.76 99.08 110.76 99.15 110.21 99.15 ;
      RECT  111.65 99.15 111.86 98.77 ;
      RECT  108.53 100.42 108.74 99.87 ;
      RECT  108.74 100.42 109.67 99.87 ;
      RECT  109.67 99.15 110.21 98.77 ;
      RECT  111.65 98.53 111.86 98.29 ;
      RECT  110.21 100.42 111.86 99.87 ;
      RECT  108.53 99.63 108.74 99.39 ;
      RECT  111.14 98.6 111.34 98.53 ;
      POLYGON  111.51 99.15 111.51 99.08 111.14 99.08 111.14 98.84 111.51 98.84 111.51 98.77 111.65 98.77 111.65 99.15 111.51 99.15 ;
      RECT  108.53 98.53 108.74 98.29 ;
      RECT  108.74 98.53 111.14 98.29 ;
      RECT  111.14 99.63 111.65 99.39 ;
      RECT  109.67 100.42 110.21 99.87 ;
      RECT  108.53 101.14 109.67 101.52 ;
      RECT  110.93 100.9 111.14 100.97 ;
      RECT  111.14 101.76 111.65 102.0 ;
      RECT  108.74 100.66 111.14 100.9 ;
      RECT  111.14 100.9 111.34 100.97 ;
      RECT  110.93 101.69 111.14 101.76 ;
      RECT  111.65 100.66 111.86 100.9 ;
      POLYGON  110.21 101.14 110.21 101.52 110.76 101.52 110.76 101.45 111.14 101.45 111.14 101.21 110.76 101.21 110.76 101.14 110.21 101.14 ;
      RECT  111.65 101.14 111.86 101.52 ;
      RECT  108.53 99.87 108.74 100.42 ;
      RECT  108.74 99.87 109.67 100.42 ;
      RECT  109.67 101.14 110.21 101.52 ;
      RECT  111.65 101.76 111.86 102.0 ;
      RECT  110.21 99.87 111.86 100.42 ;
      RECT  108.53 100.66 108.74 100.9 ;
      RECT  111.14 101.69 111.34 101.76 ;
      POLYGON  111.51 101.14 111.51 101.21 111.14 101.21 111.14 101.45 111.51 101.45 111.51 101.52 111.65 101.52 111.65 101.14 111.51 101.14 ;
      RECT  108.53 101.76 108.74 102.0 ;
      RECT  108.74 101.76 111.14 102.0 ;
      RECT  111.14 100.66 111.65 100.9 ;
      RECT  109.67 99.87 110.21 100.42 ;
      RECT  108.53 103.1 109.67 102.72 ;
      RECT  110.93 103.34 111.14 103.27 ;
      RECT  111.14 102.48 111.65 102.24 ;
      RECT  108.74 103.58 111.14 103.34 ;
      RECT  111.14 103.34 111.34 103.27 ;
      RECT  110.93 102.55 111.14 102.48 ;
      RECT  111.65 103.58 111.86 103.34 ;
      POLYGON  110.21 103.1 110.21 102.72 110.76 102.72 110.76 102.79 111.14 102.79 111.14 103.03 110.76 103.03 110.76 103.1 110.21 103.1 ;
      RECT  111.65 103.1 111.86 102.72 ;
      RECT  108.53 104.37 108.74 103.82 ;
      RECT  108.74 104.37 109.67 103.82 ;
      RECT  109.67 103.1 110.21 102.72 ;
      RECT  111.65 102.48 111.86 102.24 ;
      RECT  110.21 104.37 111.86 103.82 ;
      RECT  108.53 103.58 108.74 103.34 ;
      RECT  111.14 102.55 111.34 102.48 ;
      POLYGON  111.51 103.1 111.51 103.03 111.14 103.03 111.14 102.79 111.51 102.79 111.51 102.72 111.65 102.72 111.65 103.1 111.51 103.1 ;
      RECT  108.53 102.48 108.74 102.24 ;
      RECT  108.74 102.48 111.14 102.24 ;
      RECT  111.14 103.58 111.65 103.34 ;
      RECT  109.67 104.37 110.21 103.82 ;
      RECT  108.53 105.09 109.67 105.47 ;
      RECT  110.93 104.85 111.14 104.92 ;
      RECT  111.14 105.71 111.65 105.95 ;
      RECT  108.74 104.61 111.14 104.85 ;
      RECT  111.14 104.85 111.34 104.92 ;
      RECT  110.93 105.64 111.14 105.71 ;
      RECT  111.65 104.61 111.86 104.85 ;
      POLYGON  110.21 105.09 110.21 105.47 110.76 105.47 110.76 105.4 111.14 105.4 111.14 105.16 110.76 105.16 110.76 105.09 110.21 105.09 ;
      RECT  111.65 105.09 111.86 105.47 ;
      RECT  108.53 103.82 108.74 104.37 ;
      RECT  108.74 103.82 109.67 104.37 ;
      RECT  109.67 105.09 110.21 105.47 ;
      RECT  111.65 105.71 111.86 105.95 ;
      RECT  110.21 103.82 111.86 104.37 ;
      RECT  108.53 104.61 108.74 104.85 ;
      RECT  111.14 105.64 111.34 105.71 ;
      POLYGON  111.51 105.09 111.51 105.16 111.14 105.16 111.14 105.4 111.51 105.4 111.51 105.47 111.65 105.47 111.65 105.09 111.51 105.09 ;
      RECT  108.53 105.71 108.74 105.95 ;
      RECT  108.74 105.71 111.14 105.95 ;
      RECT  111.14 104.61 111.65 104.85 ;
      RECT  109.67 103.82 110.21 104.37 ;
      RECT  108.53 107.05 109.67 106.67 ;
      RECT  110.93 107.29 111.14 107.22 ;
      RECT  111.14 106.43 111.65 106.19 ;
      RECT  108.74 107.53 111.14 107.29 ;
      RECT  111.14 107.29 111.34 107.22 ;
      RECT  110.93 106.5 111.14 106.43 ;
      RECT  111.65 107.53 111.86 107.29 ;
      POLYGON  110.21 107.05 110.21 106.67 110.76 106.67 110.76 106.74 111.14 106.74 111.14 106.98 110.76 106.98 110.76 107.05 110.21 107.05 ;
      RECT  111.65 107.05 111.86 106.67 ;
      RECT  108.53 108.32 108.74 107.77 ;
      RECT  108.74 108.32 109.67 107.77 ;
      RECT  109.67 107.05 110.21 106.67 ;
      RECT  111.65 106.43 111.86 106.19 ;
      RECT  110.21 108.32 111.86 107.77 ;
      RECT  108.53 107.53 108.74 107.29 ;
      RECT  111.14 106.5 111.34 106.43 ;
      POLYGON  111.51 107.05 111.51 106.98 111.14 106.98 111.14 106.74 111.51 106.74 111.51 106.67 111.65 106.67 111.65 107.05 111.51 107.05 ;
      RECT  108.53 106.43 108.74 106.19 ;
      RECT  108.74 106.43 111.14 106.19 ;
      RECT  111.14 107.53 111.65 107.29 ;
      RECT  109.67 108.32 110.21 107.77 ;
      RECT  108.53 109.04 109.67 109.42 ;
      RECT  110.93 108.8 111.14 108.87 ;
      RECT  111.14 109.66 111.65 109.9 ;
      RECT  108.74 108.56 111.14 108.8 ;
      RECT  111.14 108.8 111.34 108.87 ;
      RECT  110.93 109.59 111.14 109.66 ;
      RECT  111.65 108.56 111.86 108.8 ;
      POLYGON  110.21 109.04 110.21 109.42 110.76 109.42 110.76 109.35 111.14 109.35 111.14 109.11 110.76 109.11 110.76 109.04 110.21 109.04 ;
      RECT  111.65 109.04 111.86 109.42 ;
      RECT  108.53 107.77 108.74 108.32 ;
      RECT  108.74 107.77 109.67 108.32 ;
      RECT  109.67 109.04 110.21 109.42 ;
      RECT  111.65 109.66 111.86 109.9 ;
      RECT  110.21 107.77 111.86 108.32 ;
      RECT  108.53 108.56 108.74 108.8 ;
      RECT  111.14 109.59 111.34 109.66 ;
      POLYGON  111.51 109.04 111.51 109.11 111.14 109.11 111.14 109.35 111.51 109.35 111.51 109.42 111.65 109.42 111.65 109.04 111.51 109.04 ;
      RECT  108.53 109.66 108.74 109.9 ;
      RECT  108.74 109.66 111.14 109.9 ;
      RECT  111.14 108.56 111.65 108.8 ;
      RECT  109.67 107.77 110.21 108.32 ;
      RECT  108.53 111.0 109.67 110.62 ;
      RECT  110.93 111.24 111.14 111.17 ;
      RECT  111.14 110.38 111.65 110.14 ;
      RECT  108.74 111.48 111.14 111.24 ;
      RECT  111.14 111.24 111.34 111.17 ;
      RECT  110.93 110.45 111.14 110.38 ;
      RECT  111.65 111.48 111.86 111.24 ;
      POLYGON  110.21 111.0 110.21 110.62 110.76 110.62 110.76 110.69 111.14 110.69 111.14 110.93 110.76 110.93 110.76 111.0 110.21 111.0 ;
      RECT  111.65 111.0 111.86 110.62 ;
      RECT  108.53 112.27 108.74 111.72 ;
      RECT  108.74 112.27 109.67 111.72 ;
      RECT  109.67 111.0 110.21 110.62 ;
      RECT  111.65 110.38 111.86 110.14 ;
      RECT  110.21 112.27 111.86 111.72 ;
      RECT  108.53 111.48 108.74 111.24 ;
      RECT  111.14 110.45 111.34 110.38 ;
      POLYGON  111.51 111.0 111.51 110.93 111.14 110.93 111.14 110.69 111.51 110.69 111.51 110.62 111.65 110.62 111.65 111.0 111.51 111.0 ;
      RECT  108.53 110.38 108.74 110.14 ;
      RECT  108.74 110.38 111.14 110.14 ;
      RECT  111.14 111.48 111.65 111.24 ;
      RECT  109.67 112.27 110.21 111.72 ;
      RECT  108.53 112.99 109.67 113.37 ;
      RECT  110.93 112.75 111.14 112.82 ;
      RECT  111.14 113.61 111.65 113.85 ;
      RECT  108.74 112.51 111.14 112.75 ;
      RECT  111.14 112.75 111.34 112.82 ;
      RECT  110.93 113.54 111.14 113.61 ;
      RECT  111.65 112.51 111.86 112.75 ;
      POLYGON  110.21 112.99 110.21 113.37 110.76 113.37 110.76 113.3 111.14 113.3 111.14 113.06 110.76 113.06 110.76 112.99 110.21 112.99 ;
      RECT  111.65 112.99 111.86 113.37 ;
      RECT  108.53 111.72 108.74 112.27 ;
      RECT  108.74 111.72 109.67 112.27 ;
      RECT  109.67 112.99 110.21 113.37 ;
      RECT  111.65 113.61 111.86 113.85 ;
      RECT  110.21 111.72 111.86 112.27 ;
      RECT  108.53 112.51 108.74 112.75 ;
      RECT  111.14 113.54 111.34 113.61 ;
      POLYGON  111.51 112.99 111.51 113.06 111.14 113.06 111.14 113.3 111.51 113.3 111.51 113.37 111.65 113.37 111.65 112.99 111.51 112.99 ;
      RECT  108.53 113.61 108.74 113.85 ;
      RECT  108.74 113.61 111.14 113.85 ;
      RECT  111.14 112.51 111.65 112.75 ;
      RECT  109.67 111.72 110.21 112.27 ;
      RECT  108.53 114.95 109.67 114.57 ;
      RECT  110.93 115.19 111.14 115.12 ;
      RECT  111.14 114.33 111.65 114.09 ;
      RECT  108.74 115.43 111.14 115.19 ;
      RECT  111.14 115.19 111.34 115.12 ;
      RECT  110.93 114.4 111.14 114.33 ;
      RECT  111.65 115.43 111.86 115.19 ;
      POLYGON  110.21 114.95 110.21 114.57 110.76 114.57 110.76 114.64 111.14 114.64 111.14 114.88 110.76 114.88 110.76 114.95 110.21 114.95 ;
      RECT  111.65 114.95 111.86 114.57 ;
      RECT  108.53 116.22 108.74 115.67 ;
      RECT  108.74 116.22 109.67 115.67 ;
      RECT  109.67 114.95 110.21 114.57 ;
      RECT  111.65 114.33 111.86 114.09 ;
      RECT  110.21 116.22 111.86 115.67 ;
      RECT  108.53 115.43 108.74 115.19 ;
      RECT  111.14 114.4 111.34 114.33 ;
      POLYGON  111.51 114.95 111.51 114.88 111.14 114.88 111.14 114.64 111.51 114.64 111.51 114.57 111.65 114.57 111.65 114.95 111.51 114.95 ;
      RECT  108.53 114.33 108.74 114.09 ;
      RECT  108.74 114.33 111.14 114.09 ;
      RECT  111.14 115.43 111.65 115.19 ;
      RECT  109.67 116.22 110.21 115.67 ;
      RECT  108.53 116.94 109.67 117.32 ;
      RECT  110.93 116.7 111.14 116.77 ;
      RECT  111.14 117.56 111.65 117.8 ;
      RECT  108.74 116.46 111.14 116.7 ;
      RECT  111.14 116.7 111.34 116.77 ;
      RECT  110.93 117.49 111.14 117.56 ;
      RECT  111.65 116.46 111.86 116.7 ;
      POLYGON  110.21 116.94 110.21 117.32 110.76 117.32 110.76 117.25 111.14 117.25 111.14 117.01 110.76 117.01 110.76 116.94 110.21 116.94 ;
      RECT  111.65 116.94 111.86 117.32 ;
      RECT  108.53 115.67 108.74 116.22 ;
      RECT  108.74 115.67 109.67 116.22 ;
      RECT  109.67 116.94 110.21 117.32 ;
      RECT  111.65 117.56 111.86 117.8 ;
      RECT  110.21 115.67 111.86 116.22 ;
      RECT  108.53 116.46 108.74 116.7 ;
      RECT  111.14 117.49 111.34 117.56 ;
      POLYGON  111.51 116.94 111.51 117.01 111.14 117.01 111.14 117.25 111.51 117.25 111.51 117.32 111.65 117.32 111.65 116.94 111.51 116.94 ;
      RECT  108.53 117.56 108.74 117.8 ;
      RECT  108.74 117.56 111.14 117.8 ;
      RECT  111.14 116.46 111.65 116.7 ;
      RECT  109.67 115.67 110.21 116.22 ;
      RECT  108.53 118.9 109.67 118.52 ;
      RECT  110.93 119.14 111.14 119.07 ;
      RECT  111.14 118.28 111.65 118.04 ;
      RECT  108.74 119.38 111.14 119.14 ;
      RECT  111.14 119.14 111.34 119.07 ;
      RECT  110.93 118.35 111.14 118.28 ;
      RECT  111.65 119.38 111.86 119.14 ;
      POLYGON  110.21 118.9 110.21 118.52 110.76 118.52 110.76 118.59 111.14 118.59 111.14 118.83 110.76 118.83 110.76 118.9 110.21 118.9 ;
      RECT  111.65 118.9 111.86 118.52 ;
      RECT  108.53 120.17 108.74 119.62 ;
      RECT  108.74 120.17 109.67 119.62 ;
      RECT  109.67 118.9 110.21 118.52 ;
      RECT  111.65 118.28 111.86 118.04 ;
      RECT  110.21 120.17 111.86 119.62 ;
      RECT  108.53 119.38 108.74 119.14 ;
      RECT  111.14 118.35 111.34 118.28 ;
      POLYGON  111.51 118.9 111.51 118.83 111.14 118.83 111.14 118.59 111.51 118.59 111.51 118.52 111.65 118.52 111.65 118.9 111.51 118.9 ;
      RECT  108.53 118.28 108.74 118.04 ;
      RECT  108.74 118.28 111.14 118.04 ;
      RECT  111.14 119.38 111.65 119.14 ;
      RECT  109.67 120.17 110.21 119.62 ;
      RECT  108.53 120.89 109.67 121.27 ;
      RECT  110.93 120.65 111.14 120.72 ;
      RECT  111.14 121.51 111.65 121.75 ;
      RECT  108.74 120.41 111.14 120.65 ;
      RECT  111.14 120.65 111.34 120.72 ;
      RECT  110.93 121.44 111.14 121.51 ;
      RECT  111.65 120.41 111.86 120.65 ;
      POLYGON  110.21 120.89 110.21 121.27 110.76 121.27 110.76 121.2 111.14 121.2 111.14 120.96 110.76 120.96 110.76 120.89 110.21 120.89 ;
      RECT  111.65 120.89 111.86 121.27 ;
      RECT  108.53 119.62 108.74 120.17 ;
      RECT  108.74 119.62 109.67 120.17 ;
      RECT  109.67 120.89 110.21 121.27 ;
      RECT  111.65 121.51 111.86 121.75 ;
      RECT  110.21 119.62 111.86 120.17 ;
      RECT  108.53 120.41 108.74 120.65 ;
      RECT  111.14 121.44 111.34 121.51 ;
      POLYGON  111.51 120.89 111.51 120.96 111.14 120.96 111.14 121.2 111.51 121.2 111.51 121.27 111.65 121.27 111.65 120.89 111.51 120.89 ;
      RECT  108.53 121.51 108.74 121.75 ;
      RECT  108.74 121.51 111.14 121.75 ;
      RECT  111.14 120.41 111.65 120.65 ;
      RECT  109.67 119.62 110.21 120.17 ;
      RECT  108.53 122.85 109.67 122.47 ;
      RECT  110.93 123.09 111.14 123.02 ;
      RECT  111.14 122.23 111.65 121.99 ;
      RECT  108.74 123.33 111.14 123.09 ;
      RECT  111.14 123.09 111.34 123.02 ;
      RECT  110.93 122.3 111.14 122.23 ;
      RECT  111.65 123.33 111.86 123.09 ;
      POLYGON  110.21 122.85 110.21 122.47 110.76 122.47 110.76 122.54 111.14 122.54 111.14 122.78 110.76 122.78 110.76 122.85 110.21 122.85 ;
      RECT  111.65 122.85 111.86 122.47 ;
      RECT  108.53 124.12 108.74 123.57 ;
      RECT  108.74 124.12 109.67 123.57 ;
      RECT  109.67 122.85 110.21 122.47 ;
      RECT  111.65 122.23 111.86 121.99 ;
      RECT  110.21 124.12 111.86 123.57 ;
      RECT  108.53 123.33 108.74 123.09 ;
      RECT  111.14 122.3 111.34 122.23 ;
      POLYGON  111.51 122.85 111.51 122.78 111.14 122.78 111.14 122.54 111.51 122.54 111.51 122.47 111.65 122.47 111.65 122.85 111.51 122.85 ;
      RECT  108.53 122.23 108.74 121.99 ;
      RECT  108.74 122.23 111.14 121.99 ;
      RECT  111.14 123.33 111.65 123.09 ;
      RECT  109.67 124.12 110.21 123.57 ;
      RECT  115.19 93.24 114.05 93.62 ;
      RECT  112.79 93.0 112.58 93.07 ;
      RECT  112.58 93.86 112.07 94.1 ;
      RECT  114.98 92.76 112.58 93.0 ;
      RECT  112.58 93.0 112.38 93.07 ;
      RECT  112.79 93.79 112.58 93.86 ;
      RECT  112.07 92.76 111.86 93.0 ;
      POLYGON  113.51 93.24 113.51 93.62 112.96 93.62 112.96 93.55 112.58 93.55 112.58 93.31 112.96 93.31 112.96 93.24 113.51 93.24 ;
      RECT  112.07 93.24 111.86 93.62 ;
      RECT  115.19 91.97 114.98 92.52 ;
      RECT  114.98 91.97 114.05 92.52 ;
      RECT  114.05 93.24 113.51 93.62 ;
      RECT  112.07 93.86 111.86 94.1 ;
      RECT  113.51 91.97 111.86 92.52 ;
      RECT  115.19 92.76 114.98 93.0 ;
      RECT  112.58 93.79 112.38 93.86 ;
      POLYGON  112.21 93.24 112.21 93.31 112.58 93.31 112.58 93.55 112.21 93.55 112.21 93.62 112.07 93.62 112.07 93.24 112.21 93.24 ;
      RECT  115.19 93.86 114.98 94.1 ;
      RECT  114.98 93.86 112.58 94.1 ;
      RECT  112.58 92.76 112.07 93.0 ;
      RECT  114.05 91.97 113.51 92.52 ;
      RECT  115.19 95.2 114.05 94.82 ;
      RECT  112.79 95.44 112.58 95.37 ;
      RECT  112.58 94.58 112.07 94.34 ;
      RECT  114.98 95.68 112.58 95.44 ;
      RECT  112.58 95.44 112.38 95.37 ;
      RECT  112.79 94.65 112.58 94.58 ;
      RECT  112.07 95.68 111.86 95.44 ;
      POLYGON  113.51 95.2 113.51 94.82 112.96 94.82 112.96 94.89 112.58 94.89 112.58 95.13 112.96 95.13 112.96 95.2 113.51 95.2 ;
      RECT  112.07 95.2 111.86 94.82 ;
      RECT  115.19 96.47 114.98 95.92 ;
      RECT  114.98 96.47 114.05 95.92 ;
      RECT  114.05 95.2 113.51 94.82 ;
      RECT  112.07 94.58 111.86 94.34 ;
      RECT  113.51 96.47 111.86 95.92 ;
      RECT  115.19 95.68 114.98 95.44 ;
      RECT  112.58 94.65 112.38 94.58 ;
      POLYGON  112.21 95.2 112.21 95.13 112.58 95.13 112.58 94.89 112.21 94.89 112.21 94.82 112.07 94.82 112.07 95.2 112.21 95.2 ;
      RECT  115.19 94.58 114.98 94.34 ;
      RECT  114.98 94.58 112.58 94.34 ;
      RECT  112.58 95.68 112.07 95.44 ;
      RECT  114.05 96.47 113.51 95.92 ;
      RECT  115.19 97.19 114.05 97.57 ;
      RECT  112.79 96.95 112.58 97.02 ;
      RECT  112.58 97.81 112.07 98.05 ;
      RECT  114.98 96.71 112.58 96.95 ;
      RECT  112.58 96.95 112.38 97.02 ;
      RECT  112.79 97.74 112.58 97.81 ;
      RECT  112.07 96.71 111.86 96.95 ;
      POLYGON  113.51 97.19 113.51 97.57 112.96 97.57 112.96 97.5 112.58 97.5 112.58 97.26 112.96 97.26 112.96 97.19 113.51 97.19 ;
      RECT  112.07 97.19 111.86 97.57 ;
      RECT  115.19 95.92 114.98 96.47 ;
      RECT  114.98 95.92 114.05 96.47 ;
      RECT  114.05 97.19 113.51 97.57 ;
      RECT  112.07 97.81 111.86 98.05 ;
      RECT  113.51 95.92 111.86 96.47 ;
      RECT  115.19 96.71 114.98 96.95 ;
      RECT  112.58 97.74 112.38 97.81 ;
      POLYGON  112.21 97.19 112.21 97.26 112.58 97.26 112.58 97.5 112.21 97.5 112.21 97.57 112.07 97.57 112.07 97.19 112.21 97.19 ;
      RECT  115.19 97.81 114.98 98.05 ;
      RECT  114.98 97.81 112.58 98.05 ;
      RECT  112.58 96.71 112.07 96.95 ;
      RECT  114.05 95.92 113.51 96.47 ;
      RECT  115.19 99.15 114.05 98.77 ;
      RECT  112.79 99.39 112.58 99.32 ;
      RECT  112.58 98.53 112.07 98.29 ;
      RECT  114.98 99.63 112.58 99.39 ;
      RECT  112.58 99.39 112.38 99.32 ;
      RECT  112.79 98.6 112.58 98.53 ;
      RECT  112.07 99.63 111.86 99.39 ;
      POLYGON  113.51 99.15 113.51 98.77 112.96 98.77 112.96 98.84 112.58 98.84 112.58 99.08 112.96 99.08 112.96 99.15 113.51 99.15 ;
      RECT  112.07 99.15 111.86 98.77 ;
      RECT  115.19 100.42 114.98 99.87 ;
      RECT  114.98 100.42 114.05 99.87 ;
      RECT  114.05 99.15 113.51 98.77 ;
      RECT  112.07 98.53 111.86 98.29 ;
      RECT  113.51 100.42 111.86 99.87 ;
      RECT  115.19 99.63 114.98 99.39 ;
      RECT  112.58 98.6 112.38 98.53 ;
      POLYGON  112.21 99.15 112.21 99.08 112.58 99.08 112.58 98.84 112.21 98.84 112.21 98.77 112.07 98.77 112.07 99.15 112.21 99.15 ;
      RECT  115.19 98.53 114.98 98.29 ;
      RECT  114.98 98.53 112.58 98.29 ;
      RECT  112.58 99.63 112.07 99.39 ;
      RECT  114.05 100.42 113.51 99.87 ;
      RECT  115.19 101.14 114.05 101.52 ;
      RECT  112.79 100.9 112.58 100.97 ;
      RECT  112.58 101.76 112.07 102.0 ;
      RECT  114.98 100.66 112.58 100.9 ;
      RECT  112.58 100.9 112.38 100.97 ;
      RECT  112.79 101.69 112.58 101.76 ;
      RECT  112.07 100.66 111.86 100.9 ;
      POLYGON  113.51 101.14 113.51 101.52 112.96 101.52 112.96 101.45 112.58 101.45 112.58 101.21 112.96 101.21 112.96 101.14 113.51 101.14 ;
      RECT  112.07 101.14 111.86 101.52 ;
      RECT  115.19 99.87 114.98 100.42 ;
      RECT  114.98 99.87 114.05 100.42 ;
      RECT  114.05 101.14 113.51 101.52 ;
      RECT  112.07 101.76 111.86 102.0 ;
      RECT  113.51 99.87 111.86 100.42 ;
      RECT  115.19 100.66 114.98 100.9 ;
      RECT  112.58 101.69 112.38 101.76 ;
      POLYGON  112.21 101.14 112.21 101.21 112.58 101.21 112.58 101.45 112.21 101.45 112.21 101.52 112.07 101.52 112.07 101.14 112.21 101.14 ;
      RECT  115.19 101.76 114.98 102.0 ;
      RECT  114.98 101.76 112.58 102.0 ;
      RECT  112.58 100.66 112.07 100.9 ;
      RECT  114.05 99.87 113.51 100.42 ;
      RECT  115.19 103.1 114.05 102.72 ;
      RECT  112.79 103.34 112.58 103.27 ;
      RECT  112.58 102.48 112.07 102.24 ;
      RECT  114.98 103.58 112.58 103.34 ;
      RECT  112.58 103.34 112.38 103.27 ;
      RECT  112.79 102.55 112.58 102.48 ;
      RECT  112.07 103.58 111.86 103.34 ;
      POLYGON  113.51 103.1 113.51 102.72 112.96 102.72 112.96 102.79 112.58 102.79 112.58 103.03 112.96 103.03 112.96 103.1 113.51 103.1 ;
      RECT  112.07 103.1 111.86 102.72 ;
      RECT  115.19 104.37 114.98 103.82 ;
      RECT  114.98 104.37 114.05 103.82 ;
      RECT  114.05 103.1 113.51 102.72 ;
      RECT  112.07 102.48 111.86 102.24 ;
      RECT  113.51 104.37 111.86 103.82 ;
      RECT  115.19 103.58 114.98 103.34 ;
      RECT  112.58 102.55 112.38 102.48 ;
      POLYGON  112.21 103.1 112.21 103.03 112.58 103.03 112.58 102.79 112.21 102.79 112.21 102.72 112.07 102.72 112.07 103.1 112.21 103.1 ;
      RECT  115.19 102.48 114.98 102.24 ;
      RECT  114.98 102.48 112.58 102.24 ;
      RECT  112.58 103.58 112.07 103.34 ;
      RECT  114.05 104.37 113.51 103.82 ;
      RECT  115.19 105.09 114.05 105.47 ;
      RECT  112.79 104.85 112.58 104.92 ;
      RECT  112.58 105.71 112.07 105.95 ;
      RECT  114.98 104.61 112.58 104.85 ;
      RECT  112.58 104.85 112.38 104.92 ;
      RECT  112.79 105.64 112.58 105.71 ;
      RECT  112.07 104.61 111.86 104.85 ;
      POLYGON  113.51 105.09 113.51 105.47 112.96 105.47 112.96 105.4 112.58 105.4 112.58 105.16 112.96 105.16 112.96 105.09 113.51 105.09 ;
      RECT  112.07 105.09 111.86 105.47 ;
      RECT  115.19 103.82 114.98 104.37 ;
      RECT  114.98 103.82 114.05 104.37 ;
      RECT  114.05 105.09 113.51 105.47 ;
      RECT  112.07 105.71 111.86 105.95 ;
      RECT  113.51 103.82 111.86 104.37 ;
      RECT  115.19 104.61 114.98 104.85 ;
      RECT  112.58 105.64 112.38 105.71 ;
      POLYGON  112.21 105.09 112.21 105.16 112.58 105.16 112.58 105.4 112.21 105.4 112.21 105.47 112.07 105.47 112.07 105.09 112.21 105.09 ;
      RECT  115.19 105.71 114.98 105.95 ;
      RECT  114.98 105.71 112.58 105.95 ;
      RECT  112.58 104.61 112.07 104.85 ;
      RECT  114.05 103.82 113.51 104.37 ;
      RECT  115.19 107.05 114.05 106.67 ;
      RECT  112.79 107.29 112.58 107.22 ;
      RECT  112.58 106.43 112.07 106.19 ;
      RECT  114.98 107.53 112.58 107.29 ;
      RECT  112.58 107.29 112.38 107.22 ;
      RECT  112.79 106.5 112.58 106.43 ;
      RECT  112.07 107.53 111.86 107.29 ;
      POLYGON  113.51 107.05 113.51 106.67 112.96 106.67 112.96 106.74 112.58 106.74 112.58 106.98 112.96 106.98 112.96 107.05 113.51 107.05 ;
      RECT  112.07 107.05 111.86 106.67 ;
      RECT  115.19 108.32 114.98 107.77 ;
      RECT  114.98 108.32 114.05 107.77 ;
      RECT  114.05 107.05 113.51 106.67 ;
      RECT  112.07 106.43 111.86 106.19 ;
      RECT  113.51 108.32 111.86 107.77 ;
      RECT  115.19 107.53 114.98 107.29 ;
      RECT  112.58 106.5 112.38 106.43 ;
      POLYGON  112.21 107.05 112.21 106.98 112.58 106.98 112.58 106.74 112.21 106.74 112.21 106.67 112.07 106.67 112.07 107.05 112.21 107.05 ;
      RECT  115.19 106.43 114.98 106.19 ;
      RECT  114.98 106.43 112.58 106.19 ;
      RECT  112.58 107.53 112.07 107.29 ;
      RECT  114.05 108.32 113.51 107.77 ;
      RECT  115.19 109.04 114.05 109.42 ;
      RECT  112.79 108.8 112.58 108.87 ;
      RECT  112.58 109.66 112.07 109.9 ;
      RECT  114.98 108.56 112.58 108.8 ;
      RECT  112.58 108.8 112.38 108.87 ;
      RECT  112.79 109.59 112.58 109.66 ;
      RECT  112.07 108.56 111.86 108.8 ;
      POLYGON  113.51 109.04 113.51 109.42 112.96 109.42 112.96 109.35 112.58 109.35 112.58 109.11 112.96 109.11 112.96 109.04 113.51 109.04 ;
      RECT  112.07 109.04 111.86 109.42 ;
      RECT  115.19 107.77 114.98 108.32 ;
      RECT  114.98 107.77 114.05 108.32 ;
      RECT  114.05 109.04 113.51 109.42 ;
      RECT  112.07 109.66 111.86 109.9 ;
      RECT  113.51 107.77 111.86 108.32 ;
      RECT  115.19 108.56 114.98 108.8 ;
      RECT  112.58 109.59 112.38 109.66 ;
      POLYGON  112.21 109.04 112.21 109.11 112.58 109.11 112.58 109.35 112.21 109.35 112.21 109.42 112.07 109.42 112.07 109.04 112.21 109.04 ;
      RECT  115.19 109.66 114.98 109.9 ;
      RECT  114.98 109.66 112.58 109.9 ;
      RECT  112.58 108.56 112.07 108.8 ;
      RECT  114.05 107.77 113.51 108.32 ;
      RECT  115.19 111.0 114.05 110.62 ;
      RECT  112.79 111.24 112.58 111.17 ;
      RECT  112.58 110.38 112.07 110.14 ;
      RECT  114.98 111.48 112.58 111.24 ;
      RECT  112.58 111.24 112.38 111.17 ;
      RECT  112.79 110.45 112.58 110.38 ;
      RECT  112.07 111.48 111.86 111.24 ;
      POLYGON  113.51 111.0 113.51 110.62 112.96 110.62 112.96 110.69 112.58 110.69 112.58 110.93 112.96 110.93 112.96 111.0 113.51 111.0 ;
      RECT  112.07 111.0 111.86 110.62 ;
      RECT  115.19 112.27 114.98 111.72 ;
      RECT  114.98 112.27 114.05 111.72 ;
      RECT  114.05 111.0 113.51 110.62 ;
      RECT  112.07 110.38 111.86 110.14 ;
      RECT  113.51 112.27 111.86 111.72 ;
      RECT  115.19 111.48 114.98 111.24 ;
      RECT  112.58 110.45 112.38 110.38 ;
      POLYGON  112.21 111.0 112.21 110.93 112.58 110.93 112.58 110.69 112.21 110.69 112.21 110.62 112.07 110.62 112.07 111.0 112.21 111.0 ;
      RECT  115.19 110.38 114.98 110.14 ;
      RECT  114.98 110.38 112.58 110.14 ;
      RECT  112.58 111.48 112.07 111.24 ;
      RECT  114.05 112.27 113.51 111.72 ;
      RECT  115.19 112.99 114.05 113.37 ;
      RECT  112.79 112.75 112.58 112.82 ;
      RECT  112.58 113.61 112.07 113.85 ;
      RECT  114.98 112.51 112.58 112.75 ;
      RECT  112.58 112.75 112.38 112.82 ;
      RECT  112.79 113.54 112.58 113.61 ;
      RECT  112.07 112.51 111.86 112.75 ;
      POLYGON  113.51 112.99 113.51 113.37 112.96 113.37 112.96 113.3 112.58 113.3 112.58 113.06 112.96 113.06 112.96 112.99 113.51 112.99 ;
      RECT  112.07 112.99 111.86 113.37 ;
      RECT  115.19 111.72 114.98 112.27 ;
      RECT  114.98 111.72 114.05 112.27 ;
      RECT  114.05 112.99 113.51 113.37 ;
      RECT  112.07 113.61 111.86 113.85 ;
      RECT  113.51 111.72 111.86 112.27 ;
      RECT  115.19 112.51 114.98 112.75 ;
      RECT  112.58 113.54 112.38 113.61 ;
      POLYGON  112.21 112.99 112.21 113.06 112.58 113.06 112.58 113.3 112.21 113.3 112.21 113.37 112.07 113.37 112.07 112.99 112.21 112.99 ;
      RECT  115.19 113.61 114.98 113.85 ;
      RECT  114.98 113.61 112.58 113.85 ;
      RECT  112.58 112.51 112.07 112.75 ;
      RECT  114.05 111.72 113.51 112.27 ;
      RECT  115.19 114.95 114.05 114.57 ;
      RECT  112.79 115.19 112.58 115.12 ;
      RECT  112.58 114.33 112.07 114.09 ;
      RECT  114.98 115.43 112.58 115.19 ;
      RECT  112.58 115.19 112.38 115.12 ;
      RECT  112.79 114.4 112.58 114.33 ;
      RECT  112.07 115.43 111.86 115.19 ;
      POLYGON  113.51 114.95 113.51 114.57 112.96 114.57 112.96 114.64 112.58 114.64 112.58 114.88 112.96 114.88 112.96 114.95 113.51 114.95 ;
      RECT  112.07 114.95 111.86 114.57 ;
      RECT  115.19 116.22 114.98 115.67 ;
      RECT  114.98 116.22 114.05 115.67 ;
      RECT  114.05 114.95 113.51 114.57 ;
      RECT  112.07 114.33 111.86 114.09 ;
      RECT  113.51 116.22 111.86 115.67 ;
      RECT  115.19 115.43 114.98 115.19 ;
      RECT  112.58 114.4 112.38 114.33 ;
      POLYGON  112.21 114.95 112.21 114.88 112.58 114.88 112.58 114.64 112.21 114.64 112.21 114.57 112.07 114.57 112.07 114.95 112.21 114.95 ;
      RECT  115.19 114.33 114.98 114.09 ;
      RECT  114.98 114.33 112.58 114.09 ;
      RECT  112.58 115.43 112.07 115.19 ;
      RECT  114.05 116.22 113.51 115.67 ;
      RECT  115.19 116.94 114.05 117.32 ;
      RECT  112.79 116.7 112.58 116.77 ;
      RECT  112.58 117.56 112.07 117.8 ;
      RECT  114.98 116.46 112.58 116.7 ;
      RECT  112.58 116.7 112.38 116.77 ;
      RECT  112.79 117.49 112.58 117.56 ;
      RECT  112.07 116.46 111.86 116.7 ;
      POLYGON  113.51 116.94 113.51 117.32 112.96 117.32 112.96 117.25 112.58 117.25 112.58 117.01 112.96 117.01 112.96 116.94 113.51 116.94 ;
      RECT  112.07 116.94 111.86 117.32 ;
      RECT  115.19 115.67 114.98 116.22 ;
      RECT  114.98 115.67 114.05 116.22 ;
      RECT  114.05 116.94 113.51 117.32 ;
      RECT  112.07 117.56 111.86 117.8 ;
      RECT  113.51 115.67 111.86 116.22 ;
      RECT  115.19 116.46 114.98 116.7 ;
      RECT  112.58 117.49 112.38 117.56 ;
      POLYGON  112.21 116.94 112.21 117.01 112.58 117.01 112.58 117.25 112.21 117.25 112.21 117.32 112.07 117.32 112.07 116.94 112.21 116.94 ;
      RECT  115.19 117.56 114.98 117.8 ;
      RECT  114.98 117.56 112.58 117.8 ;
      RECT  112.58 116.46 112.07 116.7 ;
      RECT  114.05 115.67 113.51 116.22 ;
      RECT  115.19 118.9 114.05 118.52 ;
      RECT  112.79 119.14 112.58 119.07 ;
      RECT  112.58 118.28 112.07 118.04 ;
      RECT  114.98 119.38 112.58 119.14 ;
      RECT  112.58 119.14 112.38 119.07 ;
      RECT  112.79 118.35 112.58 118.28 ;
      RECT  112.07 119.38 111.86 119.14 ;
      POLYGON  113.51 118.9 113.51 118.52 112.96 118.52 112.96 118.59 112.58 118.59 112.58 118.83 112.96 118.83 112.96 118.9 113.51 118.9 ;
      RECT  112.07 118.9 111.86 118.52 ;
      RECT  115.19 120.17 114.98 119.62 ;
      RECT  114.98 120.17 114.05 119.62 ;
      RECT  114.05 118.9 113.51 118.52 ;
      RECT  112.07 118.28 111.86 118.04 ;
      RECT  113.51 120.17 111.86 119.62 ;
      RECT  115.19 119.38 114.98 119.14 ;
      RECT  112.58 118.35 112.38 118.28 ;
      POLYGON  112.21 118.9 112.21 118.83 112.58 118.83 112.58 118.59 112.21 118.59 112.21 118.52 112.07 118.52 112.07 118.9 112.21 118.9 ;
      RECT  115.19 118.28 114.98 118.04 ;
      RECT  114.98 118.28 112.58 118.04 ;
      RECT  112.58 119.38 112.07 119.14 ;
      RECT  114.05 120.17 113.51 119.62 ;
      RECT  115.19 120.89 114.05 121.27 ;
      RECT  112.79 120.65 112.58 120.72 ;
      RECT  112.58 121.51 112.07 121.75 ;
      RECT  114.98 120.41 112.58 120.65 ;
      RECT  112.58 120.65 112.38 120.72 ;
      RECT  112.79 121.44 112.58 121.51 ;
      RECT  112.07 120.41 111.86 120.65 ;
      POLYGON  113.51 120.89 113.51 121.27 112.96 121.27 112.96 121.2 112.58 121.2 112.58 120.96 112.96 120.96 112.96 120.89 113.51 120.89 ;
      RECT  112.07 120.89 111.86 121.27 ;
      RECT  115.19 119.62 114.98 120.17 ;
      RECT  114.98 119.62 114.05 120.17 ;
      RECT  114.05 120.89 113.51 121.27 ;
      RECT  112.07 121.51 111.86 121.75 ;
      RECT  113.51 119.62 111.86 120.17 ;
      RECT  115.19 120.41 114.98 120.65 ;
      RECT  112.58 121.44 112.38 121.51 ;
      POLYGON  112.21 120.89 112.21 120.96 112.58 120.96 112.58 121.2 112.21 121.2 112.21 121.27 112.07 121.27 112.07 120.89 112.21 120.89 ;
      RECT  115.19 121.51 114.98 121.75 ;
      RECT  114.98 121.51 112.58 121.75 ;
      RECT  112.58 120.41 112.07 120.65 ;
      RECT  114.05 119.62 113.51 120.17 ;
      RECT  115.19 122.85 114.05 122.47 ;
      RECT  112.79 123.09 112.58 123.02 ;
      RECT  112.58 122.23 112.07 121.99 ;
      RECT  114.98 123.33 112.58 123.09 ;
      RECT  112.58 123.09 112.38 123.02 ;
      RECT  112.79 122.3 112.58 122.23 ;
      RECT  112.07 123.33 111.86 123.09 ;
      POLYGON  113.51 122.85 113.51 122.47 112.96 122.47 112.96 122.54 112.58 122.54 112.58 122.78 112.96 122.78 112.96 122.85 113.51 122.85 ;
      RECT  112.07 122.85 111.86 122.47 ;
      RECT  115.19 124.12 114.98 123.57 ;
      RECT  114.98 124.12 114.05 123.57 ;
      RECT  114.05 122.85 113.51 122.47 ;
      RECT  112.07 122.23 111.86 121.99 ;
      RECT  113.51 124.12 111.86 123.57 ;
      RECT  115.19 123.33 114.98 123.09 ;
      RECT  112.58 122.3 112.38 122.23 ;
      POLYGON  112.21 122.85 112.21 122.78 112.58 122.78 112.58 122.54 112.21 122.54 112.21 122.47 112.07 122.47 112.07 122.85 112.21 122.85 ;
      RECT  115.19 122.23 114.98 121.99 ;
      RECT  114.98 122.23 112.58 121.99 ;
      RECT  112.58 123.33 112.07 123.09 ;
      RECT  114.05 124.12 113.51 123.57 ;
      RECT  114.77 93.24 115.91 93.62 ;
      RECT  117.17 93.0 117.38 93.07 ;
      RECT  117.38 93.86 117.89 94.1 ;
      RECT  114.98 92.76 117.38 93.0 ;
      RECT  117.38 93.0 117.58 93.07 ;
      RECT  117.17 93.79 117.38 93.86 ;
      RECT  117.89 92.76 118.1 93.0 ;
      POLYGON  116.45 93.24 116.45 93.62 117.0 93.62 117.0 93.55 117.38 93.55 117.38 93.31 117.0 93.31 117.0 93.24 116.45 93.24 ;
      RECT  117.89 93.24 118.1 93.62 ;
      RECT  114.77 91.97 114.98 92.52 ;
      RECT  114.98 91.97 115.91 92.52 ;
      RECT  115.91 93.24 116.45 93.62 ;
      RECT  117.89 93.86 118.1 94.1 ;
      RECT  116.45 91.97 118.1 92.52 ;
      RECT  114.77 92.76 114.98 93.0 ;
      RECT  117.38 93.79 117.58 93.86 ;
      POLYGON  117.75 93.24 117.75 93.31 117.38 93.31 117.38 93.55 117.75 93.55 117.75 93.62 117.89 93.62 117.89 93.24 117.75 93.24 ;
      RECT  114.77 93.86 114.98 94.1 ;
      RECT  114.98 93.86 117.38 94.1 ;
      RECT  117.38 92.76 117.89 93.0 ;
      RECT  115.91 91.97 116.45 92.52 ;
      RECT  114.77 95.2 115.91 94.82 ;
      RECT  117.17 95.44 117.38 95.37 ;
      RECT  117.38 94.58 117.89 94.34 ;
      RECT  114.98 95.68 117.38 95.44 ;
      RECT  117.38 95.44 117.58 95.37 ;
      RECT  117.17 94.65 117.38 94.58 ;
      RECT  117.89 95.68 118.1 95.44 ;
      POLYGON  116.45 95.2 116.45 94.82 117.0 94.82 117.0 94.89 117.38 94.89 117.38 95.13 117.0 95.13 117.0 95.2 116.45 95.2 ;
      RECT  117.89 95.2 118.1 94.82 ;
      RECT  114.77 96.47 114.98 95.92 ;
      RECT  114.98 96.47 115.91 95.92 ;
      RECT  115.91 95.2 116.45 94.82 ;
      RECT  117.89 94.58 118.1 94.34 ;
      RECT  116.45 96.47 118.1 95.92 ;
      RECT  114.77 95.68 114.98 95.44 ;
      RECT  117.38 94.65 117.58 94.58 ;
      POLYGON  117.75 95.2 117.75 95.13 117.38 95.13 117.38 94.89 117.75 94.89 117.75 94.82 117.89 94.82 117.89 95.2 117.75 95.2 ;
      RECT  114.77 94.58 114.98 94.34 ;
      RECT  114.98 94.58 117.38 94.34 ;
      RECT  117.38 95.68 117.89 95.44 ;
      RECT  115.91 96.47 116.45 95.92 ;
      RECT  114.77 97.19 115.91 97.57 ;
      RECT  117.17 96.95 117.38 97.02 ;
      RECT  117.38 97.81 117.89 98.05 ;
      RECT  114.98 96.71 117.38 96.95 ;
      RECT  117.38 96.95 117.58 97.02 ;
      RECT  117.17 97.74 117.38 97.81 ;
      RECT  117.89 96.71 118.1 96.95 ;
      POLYGON  116.45 97.19 116.45 97.57 117.0 97.57 117.0 97.5 117.38 97.5 117.38 97.26 117.0 97.26 117.0 97.19 116.45 97.19 ;
      RECT  117.89 97.19 118.1 97.57 ;
      RECT  114.77 95.92 114.98 96.47 ;
      RECT  114.98 95.92 115.91 96.47 ;
      RECT  115.91 97.19 116.45 97.57 ;
      RECT  117.89 97.81 118.1 98.05 ;
      RECT  116.45 95.92 118.1 96.47 ;
      RECT  114.77 96.71 114.98 96.95 ;
      RECT  117.38 97.74 117.58 97.81 ;
      POLYGON  117.75 97.19 117.75 97.26 117.38 97.26 117.38 97.5 117.75 97.5 117.75 97.57 117.89 97.57 117.89 97.19 117.75 97.19 ;
      RECT  114.77 97.81 114.98 98.05 ;
      RECT  114.98 97.81 117.38 98.05 ;
      RECT  117.38 96.71 117.89 96.95 ;
      RECT  115.91 95.92 116.45 96.47 ;
      RECT  114.77 99.15 115.91 98.77 ;
      RECT  117.17 99.39 117.38 99.32 ;
      RECT  117.38 98.53 117.89 98.29 ;
      RECT  114.98 99.63 117.38 99.39 ;
      RECT  117.38 99.39 117.58 99.32 ;
      RECT  117.17 98.6 117.38 98.53 ;
      RECT  117.89 99.63 118.1 99.39 ;
      POLYGON  116.45 99.15 116.45 98.77 117.0 98.77 117.0 98.84 117.38 98.84 117.38 99.08 117.0 99.08 117.0 99.15 116.45 99.15 ;
      RECT  117.89 99.15 118.1 98.77 ;
      RECT  114.77 100.42 114.98 99.87 ;
      RECT  114.98 100.42 115.91 99.87 ;
      RECT  115.91 99.15 116.45 98.77 ;
      RECT  117.89 98.53 118.1 98.29 ;
      RECT  116.45 100.42 118.1 99.87 ;
      RECT  114.77 99.63 114.98 99.39 ;
      RECT  117.38 98.6 117.58 98.53 ;
      POLYGON  117.75 99.15 117.75 99.08 117.38 99.08 117.38 98.84 117.75 98.84 117.75 98.77 117.89 98.77 117.89 99.15 117.75 99.15 ;
      RECT  114.77 98.53 114.98 98.29 ;
      RECT  114.98 98.53 117.38 98.29 ;
      RECT  117.38 99.63 117.89 99.39 ;
      RECT  115.91 100.42 116.45 99.87 ;
      RECT  114.77 101.14 115.91 101.52 ;
      RECT  117.17 100.9 117.38 100.97 ;
      RECT  117.38 101.76 117.89 102.0 ;
      RECT  114.98 100.66 117.38 100.9 ;
      RECT  117.38 100.9 117.58 100.97 ;
      RECT  117.17 101.69 117.38 101.76 ;
      RECT  117.89 100.66 118.1 100.9 ;
      POLYGON  116.45 101.14 116.45 101.52 117.0 101.52 117.0 101.45 117.38 101.45 117.38 101.21 117.0 101.21 117.0 101.14 116.45 101.14 ;
      RECT  117.89 101.14 118.1 101.52 ;
      RECT  114.77 99.87 114.98 100.42 ;
      RECT  114.98 99.87 115.91 100.42 ;
      RECT  115.91 101.14 116.45 101.52 ;
      RECT  117.89 101.76 118.1 102.0 ;
      RECT  116.45 99.87 118.1 100.42 ;
      RECT  114.77 100.66 114.98 100.9 ;
      RECT  117.38 101.69 117.58 101.76 ;
      POLYGON  117.75 101.14 117.75 101.21 117.38 101.21 117.38 101.45 117.75 101.45 117.75 101.52 117.89 101.52 117.89 101.14 117.75 101.14 ;
      RECT  114.77 101.76 114.98 102.0 ;
      RECT  114.98 101.76 117.38 102.0 ;
      RECT  117.38 100.66 117.89 100.9 ;
      RECT  115.91 99.87 116.45 100.42 ;
      RECT  114.77 103.1 115.91 102.72 ;
      RECT  117.17 103.34 117.38 103.27 ;
      RECT  117.38 102.48 117.89 102.24 ;
      RECT  114.98 103.58 117.38 103.34 ;
      RECT  117.38 103.34 117.58 103.27 ;
      RECT  117.17 102.55 117.38 102.48 ;
      RECT  117.89 103.58 118.1 103.34 ;
      POLYGON  116.45 103.1 116.45 102.72 117.0 102.72 117.0 102.79 117.38 102.79 117.38 103.03 117.0 103.03 117.0 103.1 116.45 103.1 ;
      RECT  117.89 103.1 118.1 102.72 ;
      RECT  114.77 104.37 114.98 103.82 ;
      RECT  114.98 104.37 115.91 103.82 ;
      RECT  115.91 103.1 116.45 102.72 ;
      RECT  117.89 102.48 118.1 102.24 ;
      RECT  116.45 104.37 118.1 103.82 ;
      RECT  114.77 103.58 114.98 103.34 ;
      RECT  117.38 102.55 117.58 102.48 ;
      POLYGON  117.75 103.1 117.75 103.03 117.38 103.03 117.38 102.79 117.75 102.79 117.75 102.72 117.89 102.72 117.89 103.1 117.75 103.1 ;
      RECT  114.77 102.48 114.98 102.24 ;
      RECT  114.98 102.48 117.38 102.24 ;
      RECT  117.38 103.58 117.89 103.34 ;
      RECT  115.91 104.37 116.45 103.82 ;
      RECT  114.77 105.09 115.91 105.47 ;
      RECT  117.17 104.85 117.38 104.92 ;
      RECT  117.38 105.71 117.89 105.95 ;
      RECT  114.98 104.61 117.38 104.85 ;
      RECT  117.38 104.85 117.58 104.92 ;
      RECT  117.17 105.64 117.38 105.71 ;
      RECT  117.89 104.61 118.1 104.85 ;
      POLYGON  116.45 105.09 116.45 105.47 117.0 105.47 117.0 105.4 117.38 105.4 117.38 105.16 117.0 105.16 117.0 105.09 116.45 105.09 ;
      RECT  117.89 105.09 118.1 105.47 ;
      RECT  114.77 103.82 114.98 104.37 ;
      RECT  114.98 103.82 115.91 104.37 ;
      RECT  115.91 105.09 116.45 105.47 ;
      RECT  117.89 105.71 118.1 105.95 ;
      RECT  116.45 103.82 118.1 104.37 ;
      RECT  114.77 104.61 114.98 104.85 ;
      RECT  117.38 105.64 117.58 105.71 ;
      POLYGON  117.75 105.09 117.75 105.16 117.38 105.16 117.38 105.4 117.75 105.4 117.75 105.47 117.89 105.47 117.89 105.09 117.75 105.09 ;
      RECT  114.77 105.71 114.98 105.95 ;
      RECT  114.98 105.71 117.38 105.95 ;
      RECT  117.38 104.61 117.89 104.85 ;
      RECT  115.91 103.82 116.45 104.37 ;
      RECT  114.77 107.05 115.91 106.67 ;
      RECT  117.17 107.29 117.38 107.22 ;
      RECT  117.38 106.43 117.89 106.19 ;
      RECT  114.98 107.53 117.38 107.29 ;
      RECT  117.38 107.29 117.58 107.22 ;
      RECT  117.17 106.5 117.38 106.43 ;
      RECT  117.89 107.53 118.1 107.29 ;
      POLYGON  116.45 107.05 116.45 106.67 117.0 106.67 117.0 106.74 117.38 106.74 117.38 106.98 117.0 106.98 117.0 107.05 116.45 107.05 ;
      RECT  117.89 107.05 118.1 106.67 ;
      RECT  114.77 108.32 114.98 107.77 ;
      RECT  114.98 108.32 115.91 107.77 ;
      RECT  115.91 107.05 116.45 106.67 ;
      RECT  117.89 106.43 118.1 106.19 ;
      RECT  116.45 108.32 118.1 107.77 ;
      RECT  114.77 107.53 114.98 107.29 ;
      RECT  117.38 106.5 117.58 106.43 ;
      POLYGON  117.75 107.05 117.75 106.98 117.38 106.98 117.38 106.74 117.75 106.74 117.75 106.67 117.89 106.67 117.89 107.05 117.75 107.05 ;
      RECT  114.77 106.43 114.98 106.19 ;
      RECT  114.98 106.43 117.38 106.19 ;
      RECT  117.38 107.53 117.89 107.29 ;
      RECT  115.91 108.32 116.45 107.77 ;
      RECT  114.77 109.04 115.91 109.42 ;
      RECT  117.17 108.8 117.38 108.87 ;
      RECT  117.38 109.66 117.89 109.9 ;
      RECT  114.98 108.56 117.38 108.8 ;
      RECT  117.38 108.8 117.58 108.87 ;
      RECT  117.17 109.59 117.38 109.66 ;
      RECT  117.89 108.56 118.1 108.8 ;
      POLYGON  116.45 109.04 116.45 109.42 117.0 109.42 117.0 109.35 117.38 109.35 117.38 109.11 117.0 109.11 117.0 109.04 116.45 109.04 ;
      RECT  117.89 109.04 118.1 109.42 ;
      RECT  114.77 107.77 114.98 108.32 ;
      RECT  114.98 107.77 115.91 108.32 ;
      RECT  115.91 109.04 116.45 109.42 ;
      RECT  117.89 109.66 118.1 109.9 ;
      RECT  116.45 107.77 118.1 108.32 ;
      RECT  114.77 108.56 114.98 108.8 ;
      RECT  117.38 109.59 117.58 109.66 ;
      POLYGON  117.75 109.04 117.75 109.11 117.38 109.11 117.38 109.35 117.75 109.35 117.75 109.42 117.89 109.42 117.89 109.04 117.75 109.04 ;
      RECT  114.77 109.66 114.98 109.9 ;
      RECT  114.98 109.66 117.38 109.9 ;
      RECT  117.38 108.56 117.89 108.8 ;
      RECT  115.91 107.77 116.45 108.32 ;
      RECT  114.77 111.0 115.91 110.62 ;
      RECT  117.17 111.24 117.38 111.17 ;
      RECT  117.38 110.38 117.89 110.14 ;
      RECT  114.98 111.48 117.38 111.24 ;
      RECT  117.38 111.24 117.58 111.17 ;
      RECT  117.17 110.45 117.38 110.38 ;
      RECT  117.89 111.48 118.1 111.24 ;
      POLYGON  116.45 111.0 116.45 110.62 117.0 110.62 117.0 110.69 117.38 110.69 117.38 110.93 117.0 110.93 117.0 111.0 116.45 111.0 ;
      RECT  117.89 111.0 118.1 110.62 ;
      RECT  114.77 112.27 114.98 111.72 ;
      RECT  114.98 112.27 115.91 111.72 ;
      RECT  115.91 111.0 116.45 110.62 ;
      RECT  117.89 110.38 118.1 110.14 ;
      RECT  116.45 112.27 118.1 111.72 ;
      RECT  114.77 111.48 114.98 111.24 ;
      RECT  117.38 110.45 117.58 110.38 ;
      POLYGON  117.75 111.0 117.75 110.93 117.38 110.93 117.38 110.69 117.75 110.69 117.75 110.62 117.89 110.62 117.89 111.0 117.75 111.0 ;
      RECT  114.77 110.38 114.98 110.14 ;
      RECT  114.98 110.38 117.38 110.14 ;
      RECT  117.38 111.48 117.89 111.24 ;
      RECT  115.91 112.27 116.45 111.72 ;
      RECT  114.77 112.99 115.91 113.37 ;
      RECT  117.17 112.75 117.38 112.82 ;
      RECT  117.38 113.61 117.89 113.85 ;
      RECT  114.98 112.51 117.38 112.75 ;
      RECT  117.38 112.75 117.58 112.82 ;
      RECT  117.17 113.54 117.38 113.61 ;
      RECT  117.89 112.51 118.1 112.75 ;
      POLYGON  116.45 112.99 116.45 113.37 117.0 113.37 117.0 113.3 117.38 113.3 117.38 113.06 117.0 113.06 117.0 112.99 116.45 112.99 ;
      RECT  117.89 112.99 118.1 113.37 ;
      RECT  114.77 111.72 114.98 112.27 ;
      RECT  114.98 111.72 115.91 112.27 ;
      RECT  115.91 112.99 116.45 113.37 ;
      RECT  117.89 113.61 118.1 113.85 ;
      RECT  116.45 111.72 118.1 112.27 ;
      RECT  114.77 112.51 114.98 112.75 ;
      RECT  117.38 113.54 117.58 113.61 ;
      POLYGON  117.75 112.99 117.75 113.06 117.38 113.06 117.38 113.3 117.75 113.3 117.75 113.37 117.89 113.37 117.89 112.99 117.75 112.99 ;
      RECT  114.77 113.61 114.98 113.85 ;
      RECT  114.98 113.61 117.38 113.85 ;
      RECT  117.38 112.51 117.89 112.75 ;
      RECT  115.91 111.72 116.45 112.27 ;
      RECT  114.77 114.95 115.91 114.57 ;
      RECT  117.17 115.19 117.38 115.12 ;
      RECT  117.38 114.33 117.89 114.09 ;
      RECT  114.98 115.43 117.38 115.19 ;
      RECT  117.38 115.19 117.58 115.12 ;
      RECT  117.17 114.4 117.38 114.33 ;
      RECT  117.89 115.43 118.1 115.19 ;
      POLYGON  116.45 114.95 116.45 114.57 117.0 114.57 117.0 114.64 117.38 114.64 117.38 114.88 117.0 114.88 117.0 114.95 116.45 114.95 ;
      RECT  117.89 114.95 118.1 114.57 ;
      RECT  114.77 116.22 114.98 115.67 ;
      RECT  114.98 116.22 115.91 115.67 ;
      RECT  115.91 114.95 116.45 114.57 ;
      RECT  117.89 114.33 118.1 114.09 ;
      RECT  116.45 116.22 118.1 115.67 ;
      RECT  114.77 115.43 114.98 115.19 ;
      RECT  117.38 114.4 117.58 114.33 ;
      POLYGON  117.75 114.95 117.75 114.88 117.38 114.88 117.38 114.64 117.75 114.64 117.75 114.57 117.89 114.57 117.89 114.95 117.75 114.95 ;
      RECT  114.77 114.33 114.98 114.09 ;
      RECT  114.98 114.33 117.38 114.09 ;
      RECT  117.38 115.43 117.89 115.19 ;
      RECT  115.91 116.22 116.45 115.67 ;
      RECT  114.77 116.94 115.91 117.32 ;
      RECT  117.17 116.7 117.38 116.77 ;
      RECT  117.38 117.56 117.89 117.8 ;
      RECT  114.98 116.46 117.38 116.7 ;
      RECT  117.38 116.7 117.58 116.77 ;
      RECT  117.17 117.49 117.38 117.56 ;
      RECT  117.89 116.46 118.1 116.7 ;
      POLYGON  116.45 116.94 116.45 117.32 117.0 117.32 117.0 117.25 117.38 117.25 117.38 117.01 117.0 117.01 117.0 116.94 116.45 116.94 ;
      RECT  117.89 116.94 118.1 117.32 ;
      RECT  114.77 115.67 114.98 116.22 ;
      RECT  114.98 115.67 115.91 116.22 ;
      RECT  115.91 116.94 116.45 117.32 ;
      RECT  117.89 117.56 118.1 117.8 ;
      RECT  116.45 115.67 118.1 116.22 ;
      RECT  114.77 116.46 114.98 116.7 ;
      RECT  117.38 117.49 117.58 117.56 ;
      POLYGON  117.75 116.94 117.75 117.01 117.38 117.01 117.38 117.25 117.75 117.25 117.75 117.32 117.89 117.32 117.89 116.94 117.75 116.94 ;
      RECT  114.77 117.56 114.98 117.8 ;
      RECT  114.98 117.56 117.38 117.8 ;
      RECT  117.38 116.46 117.89 116.7 ;
      RECT  115.91 115.67 116.45 116.22 ;
      RECT  114.77 118.9 115.91 118.52 ;
      RECT  117.17 119.14 117.38 119.07 ;
      RECT  117.38 118.28 117.89 118.04 ;
      RECT  114.98 119.38 117.38 119.14 ;
      RECT  117.38 119.14 117.58 119.07 ;
      RECT  117.17 118.35 117.38 118.28 ;
      RECT  117.89 119.38 118.1 119.14 ;
      POLYGON  116.45 118.9 116.45 118.52 117.0 118.52 117.0 118.59 117.38 118.59 117.38 118.83 117.0 118.83 117.0 118.9 116.45 118.9 ;
      RECT  117.89 118.9 118.1 118.52 ;
      RECT  114.77 120.17 114.98 119.62 ;
      RECT  114.98 120.17 115.91 119.62 ;
      RECT  115.91 118.9 116.45 118.52 ;
      RECT  117.89 118.28 118.1 118.04 ;
      RECT  116.45 120.17 118.1 119.62 ;
      RECT  114.77 119.38 114.98 119.14 ;
      RECT  117.38 118.35 117.58 118.28 ;
      POLYGON  117.75 118.9 117.75 118.83 117.38 118.83 117.38 118.59 117.75 118.59 117.75 118.52 117.89 118.52 117.89 118.9 117.75 118.9 ;
      RECT  114.77 118.28 114.98 118.04 ;
      RECT  114.98 118.28 117.38 118.04 ;
      RECT  117.38 119.38 117.89 119.14 ;
      RECT  115.91 120.17 116.45 119.62 ;
      RECT  114.77 120.89 115.91 121.27 ;
      RECT  117.17 120.65 117.38 120.72 ;
      RECT  117.38 121.51 117.89 121.75 ;
      RECT  114.98 120.41 117.38 120.65 ;
      RECT  117.38 120.65 117.58 120.72 ;
      RECT  117.17 121.44 117.38 121.51 ;
      RECT  117.89 120.41 118.1 120.65 ;
      POLYGON  116.45 120.89 116.45 121.27 117.0 121.27 117.0 121.2 117.38 121.2 117.38 120.96 117.0 120.96 117.0 120.89 116.45 120.89 ;
      RECT  117.89 120.89 118.1 121.27 ;
      RECT  114.77 119.62 114.98 120.17 ;
      RECT  114.98 119.62 115.91 120.17 ;
      RECT  115.91 120.89 116.45 121.27 ;
      RECT  117.89 121.51 118.1 121.75 ;
      RECT  116.45 119.62 118.1 120.17 ;
      RECT  114.77 120.41 114.98 120.65 ;
      RECT  117.38 121.44 117.58 121.51 ;
      POLYGON  117.75 120.89 117.75 120.96 117.38 120.96 117.38 121.2 117.75 121.2 117.75 121.27 117.89 121.27 117.89 120.89 117.75 120.89 ;
      RECT  114.77 121.51 114.98 121.75 ;
      RECT  114.98 121.51 117.38 121.75 ;
      RECT  117.38 120.41 117.89 120.65 ;
      RECT  115.91 119.62 116.45 120.17 ;
      RECT  114.77 122.85 115.91 122.47 ;
      RECT  117.17 123.09 117.38 123.02 ;
      RECT  117.38 122.23 117.89 121.99 ;
      RECT  114.98 123.33 117.38 123.09 ;
      RECT  117.38 123.09 117.58 123.02 ;
      RECT  117.17 122.3 117.38 122.23 ;
      RECT  117.89 123.33 118.1 123.09 ;
      POLYGON  116.45 122.85 116.45 122.47 117.0 122.47 117.0 122.54 117.38 122.54 117.38 122.78 117.0 122.78 117.0 122.85 116.45 122.85 ;
      RECT  117.89 122.85 118.1 122.47 ;
      RECT  114.77 124.12 114.98 123.57 ;
      RECT  114.98 124.12 115.91 123.57 ;
      RECT  115.91 122.85 116.45 122.47 ;
      RECT  117.89 122.23 118.1 121.99 ;
      RECT  116.45 124.12 118.1 123.57 ;
      RECT  114.77 123.33 114.98 123.09 ;
      RECT  117.38 122.3 117.58 122.23 ;
      POLYGON  117.75 122.85 117.75 122.78 117.38 122.78 117.38 122.54 117.75 122.54 117.75 122.47 117.89 122.47 117.89 122.85 117.75 122.85 ;
      RECT  114.77 122.23 114.98 121.99 ;
      RECT  114.98 122.23 117.38 121.99 ;
      RECT  117.38 123.33 117.89 123.09 ;
      RECT  115.91 124.12 116.45 123.57 ;
      RECT  121.43 93.24 120.29 93.62 ;
      RECT  119.03 93.0 118.82 93.07 ;
      RECT  118.82 93.86 118.31 94.1 ;
      RECT  121.22 92.76 118.82 93.0 ;
      RECT  118.82 93.0 118.62 93.07 ;
      RECT  119.03 93.79 118.82 93.86 ;
      RECT  118.31 92.76 118.1 93.0 ;
      POLYGON  119.75 93.24 119.75 93.62 119.2 93.62 119.2 93.55 118.82 93.55 118.82 93.31 119.2 93.31 119.2 93.24 119.75 93.24 ;
      RECT  118.31 93.24 118.1 93.62 ;
      RECT  121.43 91.97 121.22 92.52 ;
      RECT  121.22 91.97 120.29 92.52 ;
      RECT  120.29 93.24 119.75 93.62 ;
      RECT  118.31 93.86 118.1 94.1 ;
      RECT  119.75 91.97 118.1 92.52 ;
      RECT  121.43 92.76 121.22 93.0 ;
      RECT  118.82 93.79 118.62 93.86 ;
      POLYGON  118.45 93.24 118.45 93.31 118.82 93.31 118.82 93.55 118.45 93.55 118.45 93.62 118.31 93.62 118.31 93.24 118.45 93.24 ;
      RECT  121.43 93.86 121.22 94.1 ;
      RECT  121.22 93.86 118.82 94.1 ;
      RECT  118.82 92.76 118.31 93.0 ;
      RECT  120.29 91.97 119.75 92.52 ;
      RECT  121.43 95.2 120.29 94.82 ;
      RECT  119.03 95.44 118.82 95.37 ;
      RECT  118.82 94.58 118.31 94.34 ;
      RECT  121.22 95.68 118.82 95.44 ;
      RECT  118.82 95.44 118.62 95.37 ;
      RECT  119.03 94.65 118.82 94.58 ;
      RECT  118.31 95.68 118.1 95.44 ;
      POLYGON  119.75 95.2 119.75 94.82 119.2 94.82 119.2 94.89 118.82 94.89 118.82 95.13 119.2 95.13 119.2 95.2 119.75 95.2 ;
      RECT  118.31 95.2 118.1 94.82 ;
      RECT  121.43 96.47 121.22 95.92 ;
      RECT  121.22 96.47 120.29 95.92 ;
      RECT  120.29 95.2 119.75 94.82 ;
      RECT  118.31 94.58 118.1 94.34 ;
      RECT  119.75 96.47 118.1 95.92 ;
      RECT  121.43 95.68 121.22 95.44 ;
      RECT  118.82 94.65 118.62 94.58 ;
      POLYGON  118.45 95.2 118.45 95.13 118.82 95.13 118.82 94.89 118.45 94.89 118.45 94.82 118.31 94.82 118.31 95.2 118.45 95.2 ;
      RECT  121.43 94.58 121.22 94.34 ;
      RECT  121.22 94.58 118.82 94.34 ;
      RECT  118.82 95.68 118.31 95.44 ;
      RECT  120.29 96.47 119.75 95.92 ;
      RECT  121.43 97.19 120.29 97.57 ;
      RECT  119.03 96.95 118.82 97.02 ;
      RECT  118.82 97.81 118.31 98.05 ;
      RECT  121.22 96.71 118.82 96.95 ;
      RECT  118.82 96.95 118.62 97.02 ;
      RECT  119.03 97.74 118.82 97.81 ;
      RECT  118.31 96.71 118.1 96.95 ;
      POLYGON  119.75 97.19 119.75 97.57 119.2 97.57 119.2 97.5 118.82 97.5 118.82 97.26 119.2 97.26 119.2 97.19 119.75 97.19 ;
      RECT  118.31 97.19 118.1 97.57 ;
      RECT  121.43 95.92 121.22 96.47 ;
      RECT  121.22 95.92 120.29 96.47 ;
      RECT  120.29 97.19 119.75 97.57 ;
      RECT  118.31 97.81 118.1 98.05 ;
      RECT  119.75 95.92 118.1 96.47 ;
      RECT  121.43 96.71 121.22 96.95 ;
      RECT  118.82 97.74 118.62 97.81 ;
      POLYGON  118.45 97.19 118.45 97.26 118.82 97.26 118.82 97.5 118.45 97.5 118.45 97.57 118.31 97.57 118.31 97.19 118.45 97.19 ;
      RECT  121.43 97.81 121.22 98.05 ;
      RECT  121.22 97.81 118.82 98.05 ;
      RECT  118.82 96.71 118.31 96.95 ;
      RECT  120.29 95.92 119.75 96.47 ;
      RECT  121.43 99.15 120.29 98.77 ;
      RECT  119.03 99.39 118.82 99.32 ;
      RECT  118.82 98.53 118.31 98.29 ;
      RECT  121.22 99.63 118.82 99.39 ;
      RECT  118.82 99.39 118.62 99.32 ;
      RECT  119.03 98.6 118.82 98.53 ;
      RECT  118.31 99.63 118.1 99.39 ;
      POLYGON  119.75 99.15 119.75 98.77 119.2 98.77 119.2 98.84 118.82 98.84 118.82 99.08 119.2 99.08 119.2 99.15 119.75 99.15 ;
      RECT  118.31 99.15 118.1 98.77 ;
      RECT  121.43 100.42 121.22 99.87 ;
      RECT  121.22 100.42 120.29 99.87 ;
      RECT  120.29 99.15 119.75 98.77 ;
      RECT  118.31 98.53 118.1 98.29 ;
      RECT  119.75 100.42 118.1 99.87 ;
      RECT  121.43 99.63 121.22 99.39 ;
      RECT  118.82 98.6 118.62 98.53 ;
      POLYGON  118.45 99.15 118.45 99.08 118.82 99.08 118.82 98.84 118.45 98.84 118.45 98.77 118.31 98.77 118.31 99.15 118.45 99.15 ;
      RECT  121.43 98.53 121.22 98.29 ;
      RECT  121.22 98.53 118.82 98.29 ;
      RECT  118.82 99.63 118.31 99.39 ;
      RECT  120.29 100.42 119.75 99.87 ;
      RECT  121.43 101.14 120.29 101.52 ;
      RECT  119.03 100.9 118.82 100.97 ;
      RECT  118.82 101.76 118.31 102.0 ;
      RECT  121.22 100.66 118.82 100.9 ;
      RECT  118.82 100.9 118.62 100.97 ;
      RECT  119.03 101.69 118.82 101.76 ;
      RECT  118.31 100.66 118.1 100.9 ;
      POLYGON  119.75 101.14 119.75 101.52 119.2 101.52 119.2 101.45 118.82 101.45 118.82 101.21 119.2 101.21 119.2 101.14 119.75 101.14 ;
      RECT  118.31 101.14 118.1 101.52 ;
      RECT  121.43 99.87 121.22 100.42 ;
      RECT  121.22 99.87 120.29 100.42 ;
      RECT  120.29 101.14 119.75 101.52 ;
      RECT  118.31 101.76 118.1 102.0 ;
      RECT  119.75 99.87 118.1 100.42 ;
      RECT  121.43 100.66 121.22 100.9 ;
      RECT  118.82 101.69 118.62 101.76 ;
      POLYGON  118.45 101.14 118.45 101.21 118.82 101.21 118.82 101.45 118.45 101.45 118.45 101.52 118.31 101.52 118.31 101.14 118.45 101.14 ;
      RECT  121.43 101.76 121.22 102.0 ;
      RECT  121.22 101.76 118.82 102.0 ;
      RECT  118.82 100.66 118.31 100.9 ;
      RECT  120.29 99.87 119.75 100.42 ;
      RECT  121.43 103.1 120.29 102.72 ;
      RECT  119.03 103.34 118.82 103.27 ;
      RECT  118.82 102.48 118.31 102.24 ;
      RECT  121.22 103.58 118.82 103.34 ;
      RECT  118.82 103.34 118.62 103.27 ;
      RECT  119.03 102.55 118.82 102.48 ;
      RECT  118.31 103.58 118.1 103.34 ;
      POLYGON  119.75 103.1 119.75 102.72 119.2 102.72 119.2 102.79 118.82 102.79 118.82 103.03 119.2 103.03 119.2 103.1 119.75 103.1 ;
      RECT  118.31 103.1 118.1 102.72 ;
      RECT  121.43 104.37 121.22 103.82 ;
      RECT  121.22 104.37 120.29 103.82 ;
      RECT  120.29 103.1 119.75 102.72 ;
      RECT  118.31 102.48 118.1 102.24 ;
      RECT  119.75 104.37 118.1 103.82 ;
      RECT  121.43 103.58 121.22 103.34 ;
      RECT  118.82 102.55 118.62 102.48 ;
      POLYGON  118.45 103.1 118.45 103.03 118.82 103.03 118.82 102.79 118.45 102.79 118.45 102.72 118.31 102.72 118.31 103.1 118.45 103.1 ;
      RECT  121.43 102.48 121.22 102.24 ;
      RECT  121.22 102.48 118.82 102.24 ;
      RECT  118.82 103.58 118.31 103.34 ;
      RECT  120.29 104.37 119.75 103.82 ;
      RECT  121.43 105.09 120.29 105.47 ;
      RECT  119.03 104.85 118.82 104.92 ;
      RECT  118.82 105.71 118.31 105.95 ;
      RECT  121.22 104.61 118.82 104.85 ;
      RECT  118.82 104.85 118.62 104.92 ;
      RECT  119.03 105.64 118.82 105.71 ;
      RECT  118.31 104.61 118.1 104.85 ;
      POLYGON  119.75 105.09 119.75 105.47 119.2 105.47 119.2 105.4 118.82 105.4 118.82 105.16 119.2 105.16 119.2 105.09 119.75 105.09 ;
      RECT  118.31 105.09 118.1 105.47 ;
      RECT  121.43 103.82 121.22 104.37 ;
      RECT  121.22 103.82 120.29 104.37 ;
      RECT  120.29 105.09 119.75 105.47 ;
      RECT  118.31 105.71 118.1 105.95 ;
      RECT  119.75 103.82 118.1 104.37 ;
      RECT  121.43 104.61 121.22 104.85 ;
      RECT  118.82 105.64 118.62 105.71 ;
      POLYGON  118.45 105.09 118.45 105.16 118.82 105.16 118.82 105.4 118.45 105.4 118.45 105.47 118.31 105.47 118.31 105.09 118.45 105.09 ;
      RECT  121.43 105.71 121.22 105.95 ;
      RECT  121.22 105.71 118.82 105.95 ;
      RECT  118.82 104.61 118.31 104.85 ;
      RECT  120.29 103.82 119.75 104.37 ;
      RECT  121.43 107.05 120.29 106.67 ;
      RECT  119.03 107.29 118.82 107.22 ;
      RECT  118.82 106.43 118.31 106.19 ;
      RECT  121.22 107.53 118.82 107.29 ;
      RECT  118.82 107.29 118.62 107.22 ;
      RECT  119.03 106.5 118.82 106.43 ;
      RECT  118.31 107.53 118.1 107.29 ;
      POLYGON  119.75 107.05 119.75 106.67 119.2 106.67 119.2 106.74 118.82 106.74 118.82 106.98 119.2 106.98 119.2 107.05 119.75 107.05 ;
      RECT  118.31 107.05 118.1 106.67 ;
      RECT  121.43 108.32 121.22 107.77 ;
      RECT  121.22 108.32 120.29 107.77 ;
      RECT  120.29 107.05 119.75 106.67 ;
      RECT  118.31 106.43 118.1 106.19 ;
      RECT  119.75 108.32 118.1 107.77 ;
      RECT  121.43 107.53 121.22 107.29 ;
      RECT  118.82 106.5 118.62 106.43 ;
      POLYGON  118.45 107.05 118.45 106.98 118.82 106.98 118.82 106.74 118.45 106.74 118.45 106.67 118.31 106.67 118.31 107.05 118.45 107.05 ;
      RECT  121.43 106.43 121.22 106.19 ;
      RECT  121.22 106.43 118.82 106.19 ;
      RECT  118.82 107.53 118.31 107.29 ;
      RECT  120.29 108.32 119.75 107.77 ;
      RECT  121.43 109.04 120.29 109.42 ;
      RECT  119.03 108.8 118.82 108.87 ;
      RECT  118.82 109.66 118.31 109.9 ;
      RECT  121.22 108.56 118.82 108.8 ;
      RECT  118.82 108.8 118.62 108.87 ;
      RECT  119.03 109.59 118.82 109.66 ;
      RECT  118.31 108.56 118.1 108.8 ;
      POLYGON  119.75 109.04 119.75 109.42 119.2 109.42 119.2 109.35 118.82 109.35 118.82 109.11 119.2 109.11 119.2 109.04 119.75 109.04 ;
      RECT  118.31 109.04 118.1 109.42 ;
      RECT  121.43 107.77 121.22 108.32 ;
      RECT  121.22 107.77 120.29 108.32 ;
      RECT  120.29 109.04 119.75 109.42 ;
      RECT  118.31 109.66 118.1 109.9 ;
      RECT  119.75 107.77 118.1 108.32 ;
      RECT  121.43 108.56 121.22 108.8 ;
      RECT  118.82 109.59 118.62 109.66 ;
      POLYGON  118.45 109.04 118.45 109.11 118.82 109.11 118.82 109.35 118.45 109.35 118.45 109.42 118.31 109.42 118.31 109.04 118.45 109.04 ;
      RECT  121.43 109.66 121.22 109.9 ;
      RECT  121.22 109.66 118.82 109.9 ;
      RECT  118.82 108.56 118.31 108.8 ;
      RECT  120.29 107.77 119.75 108.32 ;
      RECT  121.43 111.0 120.29 110.62 ;
      RECT  119.03 111.24 118.82 111.17 ;
      RECT  118.82 110.38 118.31 110.14 ;
      RECT  121.22 111.48 118.82 111.24 ;
      RECT  118.82 111.24 118.62 111.17 ;
      RECT  119.03 110.45 118.82 110.38 ;
      RECT  118.31 111.48 118.1 111.24 ;
      POLYGON  119.75 111.0 119.75 110.62 119.2 110.62 119.2 110.69 118.82 110.69 118.82 110.93 119.2 110.93 119.2 111.0 119.75 111.0 ;
      RECT  118.31 111.0 118.1 110.62 ;
      RECT  121.43 112.27 121.22 111.72 ;
      RECT  121.22 112.27 120.29 111.72 ;
      RECT  120.29 111.0 119.75 110.62 ;
      RECT  118.31 110.38 118.1 110.14 ;
      RECT  119.75 112.27 118.1 111.72 ;
      RECT  121.43 111.48 121.22 111.24 ;
      RECT  118.82 110.45 118.62 110.38 ;
      POLYGON  118.45 111.0 118.45 110.93 118.82 110.93 118.82 110.69 118.45 110.69 118.45 110.62 118.31 110.62 118.31 111.0 118.45 111.0 ;
      RECT  121.43 110.38 121.22 110.14 ;
      RECT  121.22 110.38 118.82 110.14 ;
      RECT  118.82 111.48 118.31 111.24 ;
      RECT  120.29 112.27 119.75 111.72 ;
      RECT  121.43 112.99 120.29 113.37 ;
      RECT  119.03 112.75 118.82 112.82 ;
      RECT  118.82 113.61 118.31 113.85 ;
      RECT  121.22 112.51 118.82 112.75 ;
      RECT  118.82 112.75 118.62 112.82 ;
      RECT  119.03 113.54 118.82 113.61 ;
      RECT  118.31 112.51 118.1 112.75 ;
      POLYGON  119.75 112.99 119.75 113.37 119.2 113.37 119.2 113.3 118.82 113.3 118.82 113.06 119.2 113.06 119.2 112.99 119.75 112.99 ;
      RECT  118.31 112.99 118.1 113.37 ;
      RECT  121.43 111.72 121.22 112.27 ;
      RECT  121.22 111.72 120.29 112.27 ;
      RECT  120.29 112.99 119.75 113.37 ;
      RECT  118.31 113.61 118.1 113.85 ;
      RECT  119.75 111.72 118.1 112.27 ;
      RECT  121.43 112.51 121.22 112.75 ;
      RECT  118.82 113.54 118.62 113.61 ;
      POLYGON  118.45 112.99 118.45 113.06 118.82 113.06 118.82 113.3 118.45 113.3 118.45 113.37 118.31 113.37 118.31 112.99 118.45 112.99 ;
      RECT  121.43 113.61 121.22 113.85 ;
      RECT  121.22 113.61 118.82 113.85 ;
      RECT  118.82 112.51 118.31 112.75 ;
      RECT  120.29 111.72 119.75 112.27 ;
      RECT  121.43 114.95 120.29 114.57 ;
      RECT  119.03 115.19 118.82 115.12 ;
      RECT  118.82 114.33 118.31 114.09 ;
      RECT  121.22 115.43 118.82 115.19 ;
      RECT  118.82 115.19 118.62 115.12 ;
      RECT  119.03 114.4 118.82 114.33 ;
      RECT  118.31 115.43 118.1 115.19 ;
      POLYGON  119.75 114.95 119.75 114.57 119.2 114.57 119.2 114.64 118.82 114.64 118.82 114.88 119.2 114.88 119.2 114.95 119.75 114.95 ;
      RECT  118.31 114.95 118.1 114.57 ;
      RECT  121.43 116.22 121.22 115.67 ;
      RECT  121.22 116.22 120.29 115.67 ;
      RECT  120.29 114.95 119.75 114.57 ;
      RECT  118.31 114.33 118.1 114.09 ;
      RECT  119.75 116.22 118.1 115.67 ;
      RECT  121.43 115.43 121.22 115.19 ;
      RECT  118.82 114.4 118.62 114.33 ;
      POLYGON  118.45 114.95 118.45 114.88 118.82 114.88 118.82 114.64 118.45 114.64 118.45 114.57 118.31 114.57 118.31 114.95 118.45 114.95 ;
      RECT  121.43 114.33 121.22 114.09 ;
      RECT  121.22 114.33 118.82 114.09 ;
      RECT  118.82 115.43 118.31 115.19 ;
      RECT  120.29 116.22 119.75 115.67 ;
      RECT  121.43 116.94 120.29 117.32 ;
      RECT  119.03 116.7 118.82 116.77 ;
      RECT  118.82 117.56 118.31 117.8 ;
      RECT  121.22 116.46 118.82 116.7 ;
      RECT  118.82 116.7 118.62 116.77 ;
      RECT  119.03 117.49 118.82 117.56 ;
      RECT  118.31 116.46 118.1 116.7 ;
      POLYGON  119.75 116.94 119.75 117.32 119.2 117.32 119.2 117.25 118.82 117.25 118.82 117.01 119.2 117.01 119.2 116.94 119.75 116.94 ;
      RECT  118.31 116.94 118.1 117.32 ;
      RECT  121.43 115.67 121.22 116.22 ;
      RECT  121.22 115.67 120.29 116.22 ;
      RECT  120.29 116.94 119.75 117.32 ;
      RECT  118.31 117.56 118.1 117.8 ;
      RECT  119.75 115.67 118.1 116.22 ;
      RECT  121.43 116.46 121.22 116.7 ;
      RECT  118.82 117.49 118.62 117.56 ;
      POLYGON  118.45 116.94 118.45 117.01 118.82 117.01 118.82 117.25 118.45 117.25 118.45 117.32 118.31 117.32 118.31 116.94 118.45 116.94 ;
      RECT  121.43 117.56 121.22 117.8 ;
      RECT  121.22 117.56 118.82 117.8 ;
      RECT  118.82 116.46 118.31 116.7 ;
      RECT  120.29 115.67 119.75 116.22 ;
      RECT  121.43 118.9 120.29 118.52 ;
      RECT  119.03 119.14 118.82 119.07 ;
      RECT  118.82 118.28 118.31 118.04 ;
      RECT  121.22 119.38 118.82 119.14 ;
      RECT  118.82 119.14 118.62 119.07 ;
      RECT  119.03 118.35 118.82 118.28 ;
      RECT  118.31 119.38 118.1 119.14 ;
      POLYGON  119.75 118.9 119.75 118.52 119.2 118.52 119.2 118.59 118.82 118.59 118.82 118.83 119.2 118.83 119.2 118.9 119.75 118.9 ;
      RECT  118.31 118.9 118.1 118.52 ;
      RECT  121.43 120.17 121.22 119.62 ;
      RECT  121.22 120.17 120.29 119.62 ;
      RECT  120.29 118.9 119.75 118.52 ;
      RECT  118.31 118.28 118.1 118.04 ;
      RECT  119.75 120.17 118.1 119.62 ;
      RECT  121.43 119.38 121.22 119.14 ;
      RECT  118.82 118.35 118.62 118.28 ;
      POLYGON  118.45 118.9 118.45 118.83 118.82 118.83 118.82 118.59 118.45 118.59 118.45 118.52 118.31 118.52 118.31 118.9 118.45 118.9 ;
      RECT  121.43 118.28 121.22 118.04 ;
      RECT  121.22 118.28 118.82 118.04 ;
      RECT  118.82 119.38 118.31 119.14 ;
      RECT  120.29 120.17 119.75 119.62 ;
      RECT  121.43 120.89 120.29 121.27 ;
      RECT  119.03 120.65 118.82 120.72 ;
      RECT  118.82 121.51 118.31 121.75 ;
      RECT  121.22 120.41 118.82 120.65 ;
      RECT  118.82 120.65 118.62 120.72 ;
      RECT  119.03 121.44 118.82 121.51 ;
      RECT  118.31 120.41 118.1 120.65 ;
      POLYGON  119.75 120.89 119.75 121.27 119.2 121.27 119.2 121.2 118.82 121.2 118.82 120.96 119.2 120.96 119.2 120.89 119.75 120.89 ;
      RECT  118.31 120.89 118.1 121.27 ;
      RECT  121.43 119.62 121.22 120.17 ;
      RECT  121.22 119.62 120.29 120.17 ;
      RECT  120.29 120.89 119.75 121.27 ;
      RECT  118.31 121.51 118.1 121.75 ;
      RECT  119.75 119.62 118.1 120.17 ;
      RECT  121.43 120.41 121.22 120.65 ;
      RECT  118.82 121.44 118.62 121.51 ;
      POLYGON  118.45 120.89 118.45 120.96 118.82 120.96 118.82 121.2 118.45 121.2 118.45 121.27 118.31 121.27 118.31 120.89 118.45 120.89 ;
      RECT  121.43 121.51 121.22 121.75 ;
      RECT  121.22 121.51 118.82 121.75 ;
      RECT  118.82 120.41 118.31 120.65 ;
      RECT  120.29 119.62 119.75 120.17 ;
      RECT  121.43 122.85 120.29 122.47 ;
      RECT  119.03 123.09 118.82 123.02 ;
      RECT  118.82 122.23 118.31 121.99 ;
      RECT  121.22 123.33 118.82 123.09 ;
      RECT  118.82 123.09 118.62 123.02 ;
      RECT  119.03 122.3 118.82 122.23 ;
      RECT  118.31 123.33 118.1 123.09 ;
      POLYGON  119.75 122.85 119.75 122.47 119.2 122.47 119.2 122.54 118.82 122.54 118.82 122.78 119.2 122.78 119.2 122.85 119.75 122.85 ;
      RECT  118.31 122.85 118.1 122.47 ;
      RECT  121.43 124.12 121.22 123.57 ;
      RECT  121.22 124.12 120.29 123.57 ;
      RECT  120.29 122.85 119.75 122.47 ;
      RECT  118.31 122.23 118.1 121.99 ;
      RECT  119.75 124.12 118.1 123.57 ;
      RECT  121.43 123.33 121.22 123.09 ;
      RECT  118.82 122.3 118.62 122.23 ;
      POLYGON  118.45 122.85 118.45 122.78 118.82 122.78 118.82 122.54 118.45 122.54 118.45 122.47 118.31 122.47 118.31 122.85 118.45 122.85 ;
      RECT  121.43 122.23 121.22 121.99 ;
      RECT  121.22 122.23 118.82 121.99 ;
      RECT  118.82 123.33 118.31 123.09 ;
      RECT  120.29 124.12 119.75 123.57 ;
      RECT  121.01 93.24 122.15 93.62 ;
      RECT  123.41 93.0 123.62 93.07 ;
      RECT  123.62 93.86 124.13 94.1 ;
      RECT  121.22 92.76 123.62 93.0 ;
      RECT  123.62 93.0 123.82 93.07 ;
      RECT  123.41 93.79 123.62 93.86 ;
      RECT  124.13 92.76 124.34 93.0 ;
      POLYGON  122.69 93.24 122.69 93.62 123.24 93.62 123.24 93.55 123.62 93.55 123.62 93.31 123.24 93.31 123.24 93.24 122.69 93.24 ;
      RECT  124.13 93.24 124.34 93.62 ;
      RECT  121.01 91.97 121.22 92.52 ;
      RECT  121.22 91.97 122.15 92.52 ;
      RECT  122.15 93.24 122.69 93.62 ;
      RECT  124.13 93.86 124.34 94.1 ;
      RECT  122.69 91.97 124.34 92.52 ;
      RECT  121.01 92.76 121.22 93.0 ;
      RECT  123.62 93.79 123.82 93.86 ;
      POLYGON  123.99 93.24 123.99 93.31 123.62 93.31 123.62 93.55 123.99 93.55 123.99 93.62 124.13 93.62 124.13 93.24 123.99 93.24 ;
      RECT  121.01 93.86 121.22 94.1 ;
      RECT  121.22 93.86 123.62 94.1 ;
      RECT  123.62 92.76 124.13 93.0 ;
      RECT  122.15 91.97 122.69 92.52 ;
      RECT  121.01 95.2 122.15 94.82 ;
      RECT  123.41 95.44 123.62 95.37 ;
      RECT  123.62 94.58 124.13 94.34 ;
      RECT  121.22 95.68 123.62 95.44 ;
      RECT  123.62 95.44 123.82 95.37 ;
      RECT  123.41 94.65 123.62 94.58 ;
      RECT  124.13 95.68 124.34 95.44 ;
      POLYGON  122.69 95.2 122.69 94.82 123.24 94.82 123.24 94.89 123.62 94.89 123.62 95.13 123.24 95.13 123.24 95.2 122.69 95.2 ;
      RECT  124.13 95.2 124.34 94.82 ;
      RECT  121.01 96.47 121.22 95.92 ;
      RECT  121.22 96.47 122.15 95.92 ;
      RECT  122.15 95.2 122.69 94.82 ;
      RECT  124.13 94.58 124.34 94.34 ;
      RECT  122.69 96.47 124.34 95.92 ;
      RECT  121.01 95.68 121.22 95.44 ;
      RECT  123.62 94.65 123.82 94.58 ;
      POLYGON  123.99 95.2 123.99 95.13 123.62 95.13 123.62 94.89 123.99 94.89 123.99 94.82 124.13 94.82 124.13 95.2 123.99 95.2 ;
      RECT  121.01 94.58 121.22 94.34 ;
      RECT  121.22 94.58 123.62 94.34 ;
      RECT  123.62 95.68 124.13 95.44 ;
      RECT  122.15 96.47 122.69 95.92 ;
      RECT  121.01 97.19 122.15 97.57 ;
      RECT  123.41 96.95 123.62 97.02 ;
      RECT  123.62 97.81 124.13 98.05 ;
      RECT  121.22 96.71 123.62 96.95 ;
      RECT  123.62 96.95 123.82 97.02 ;
      RECT  123.41 97.74 123.62 97.81 ;
      RECT  124.13 96.71 124.34 96.95 ;
      POLYGON  122.69 97.19 122.69 97.57 123.24 97.57 123.24 97.5 123.62 97.5 123.62 97.26 123.24 97.26 123.24 97.19 122.69 97.19 ;
      RECT  124.13 97.19 124.34 97.57 ;
      RECT  121.01 95.92 121.22 96.47 ;
      RECT  121.22 95.92 122.15 96.47 ;
      RECT  122.15 97.19 122.69 97.57 ;
      RECT  124.13 97.81 124.34 98.05 ;
      RECT  122.69 95.92 124.34 96.47 ;
      RECT  121.01 96.71 121.22 96.95 ;
      RECT  123.62 97.74 123.82 97.81 ;
      POLYGON  123.99 97.19 123.99 97.26 123.62 97.26 123.62 97.5 123.99 97.5 123.99 97.57 124.13 97.57 124.13 97.19 123.99 97.19 ;
      RECT  121.01 97.81 121.22 98.05 ;
      RECT  121.22 97.81 123.62 98.05 ;
      RECT  123.62 96.71 124.13 96.95 ;
      RECT  122.15 95.92 122.69 96.47 ;
      RECT  121.01 99.15 122.15 98.77 ;
      RECT  123.41 99.39 123.62 99.32 ;
      RECT  123.62 98.53 124.13 98.29 ;
      RECT  121.22 99.63 123.62 99.39 ;
      RECT  123.62 99.39 123.82 99.32 ;
      RECT  123.41 98.6 123.62 98.53 ;
      RECT  124.13 99.63 124.34 99.39 ;
      POLYGON  122.69 99.15 122.69 98.77 123.24 98.77 123.24 98.84 123.62 98.84 123.62 99.08 123.24 99.08 123.24 99.15 122.69 99.15 ;
      RECT  124.13 99.15 124.34 98.77 ;
      RECT  121.01 100.42 121.22 99.87 ;
      RECT  121.22 100.42 122.15 99.87 ;
      RECT  122.15 99.15 122.69 98.77 ;
      RECT  124.13 98.53 124.34 98.29 ;
      RECT  122.69 100.42 124.34 99.87 ;
      RECT  121.01 99.63 121.22 99.39 ;
      RECT  123.62 98.6 123.82 98.53 ;
      POLYGON  123.99 99.15 123.99 99.08 123.62 99.08 123.62 98.84 123.99 98.84 123.99 98.77 124.13 98.77 124.13 99.15 123.99 99.15 ;
      RECT  121.01 98.53 121.22 98.29 ;
      RECT  121.22 98.53 123.62 98.29 ;
      RECT  123.62 99.63 124.13 99.39 ;
      RECT  122.15 100.42 122.69 99.87 ;
      RECT  121.01 101.14 122.15 101.52 ;
      RECT  123.41 100.9 123.62 100.97 ;
      RECT  123.62 101.76 124.13 102.0 ;
      RECT  121.22 100.66 123.62 100.9 ;
      RECT  123.62 100.9 123.82 100.97 ;
      RECT  123.41 101.69 123.62 101.76 ;
      RECT  124.13 100.66 124.34 100.9 ;
      POLYGON  122.69 101.14 122.69 101.52 123.24 101.52 123.24 101.45 123.62 101.45 123.62 101.21 123.24 101.21 123.24 101.14 122.69 101.14 ;
      RECT  124.13 101.14 124.34 101.52 ;
      RECT  121.01 99.87 121.22 100.42 ;
      RECT  121.22 99.87 122.15 100.42 ;
      RECT  122.15 101.14 122.69 101.52 ;
      RECT  124.13 101.76 124.34 102.0 ;
      RECT  122.69 99.87 124.34 100.42 ;
      RECT  121.01 100.66 121.22 100.9 ;
      RECT  123.62 101.69 123.82 101.76 ;
      POLYGON  123.99 101.14 123.99 101.21 123.62 101.21 123.62 101.45 123.99 101.45 123.99 101.52 124.13 101.52 124.13 101.14 123.99 101.14 ;
      RECT  121.01 101.76 121.22 102.0 ;
      RECT  121.22 101.76 123.62 102.0 ;
      RECT  123.62 100.66 124.13 100.9 ;
      RECT  122.15 99.87 122.69 100.42 ;
      RECT  121.01 103.1 122.15 102.72 ;
      RECT  123.41 103.34 123.62 103.27 ;
      RECT  123.62 102.48 124.13 102.24 ;
      RECT  121.22 103.58 123.62 103.34 ;
      RECT  123.62 103.34 123.82 103.27 ;
      RECT  123.41 102.55 123.62 102.48 ;
      RECT  124.13 103.58 124.34 103.34 ;
      POLYGON  122.69 103.1 122.69 102.72 123.24 102.72 123.24 102.79 123.62 102.79 123.62 103.03 123.24 103.03 123.24 103.1 122.69 103.1 ;
      RECT  124.13 103.1 124.34 102.72 ;
      RECT  121.01 104.37 121.22 103.82 ;
      RECT  121.22 104.37 122.15 103.82 ;
      RECT  122.15 103.1 122.69 102.72 ;
      RECT  124.13 102.48 124.34 102.24 ;
      RECT  122.69 104.37 124.34 103.82 ;
      RECT  121.01 103.58 121.22 103.34 ;
      RECT  123.62 102.55 123.82 102.48 ;
      POLYGON  123.99 103.1 123.99 103.03 123.62 103.03 123.62 102.79 123.99 102.79 123.99 102.72 124.13 102.72 124.13 103.1 123.99 103.1 ;
      RECT  121.01 102.48 121.22 102.24 ;
      RECT  121.22 102.48 123.62 102.24 ;
      RECT  123.62 103.58 124.13 103.34 ;
      RECT  122.15 104.37 122.69 103.82 ;
      RECT  121.01 105.09 122.15 105.47 ;
      RECT  123.41 104.85 123.62 104.92 ;
      RECT  123.62 105.71 124.13 105.95 ;
      RECT  121.22 104.61 123.62 104.85 ;
      RECT  123.62 104.85 123.82 104.92 ;
      RECT  123.41 105.64 123.62 105.71 ;
      RECT  124.13 104.61 124.34 104.85 ;
      POLYGON  122.69 105.09 122.69 105.47 123.24 105.47 123.24 105.4 123.62 105.4 123.62 105.16 123.24 105.16 123.24 105.09 122.69 105.09 ;
      RECT  124.13 105.09 124.34 105.47 ;
      RECT  121.01 103.82 121.22 104.37 ;
      RECT  121.22 103.82 122.15 104.37 ;
      RECT  122.15 105.09 122.69 105.47 ;
      RECT  124.13 105.71 124.34 105.95 ;
      RECT  122.69 103.82 124.34 104.37 ;
      RECT  121.01 104.61 121.22 104.85 ;
      RECT  123.62 105.64 123.82 105.71 ;
      POLYGON  123.99 105.09 123.99 105.16 123.62 105.16 123.62 105.4 123.99 105.4 123.99 105.47 124.13 105.47 124.13 105.09 123.99 105.09 ;
      RECT  121.01 105.71 121.22 105.95 ;
      RECT  121.22 105.71 123.62 105.95 ;
      RECT  123.62 104.61 124.13 104.85 ;
      RECT  122.15 103.82 122.69 104.37 ;
      RECT  121.01 107.05 122.15 106.67 ;
      RECT  123.41 107.29 123.62 107.22 ;
      RECT  123.62 106.43 124.13 106.19 ;
      RECT  121.22 107.53 123.62 107.29 ;
      RECT  123.62 107.29 123.82 107.22 ;
      RECT  123.41 106.5 123.62 106.43 ;
      RECT  124.13 107.53 124.34 107.29 ;
      POLYGON  122.69 107.05 122.69 106.67 123.24 106.67 123.24 106.74 123.62 106.74 123.62 106.98 123.24 106.98 123.24 107.05 122.69 107.05 ;
      RECT  124.13 107.05 124.34 106.67 ;
      RECT  121.01 108.32 121.22 107.77 ;
      RECT  121.22 108.32 122.15 107.77 ;
      RECT  122.15 107.05 122.69 106.67 ;
      RECT  124.13 106.43 124.34 106.19 ;
      RECT  122.69 108.32 124.34 107.77 ;
      RECT  121.01 107.53 121.22 107.29 ;
      RECT  123.62 106.5 123.82 106.43 ;
      POLYGON  123.99 107.05 123.99 106.98 123.62 106.98 123.62 106.74 123.99 106.74 123.99 106.67 124.13 106.67 124.13 107.05 123.99 107.05 ;
      RECT  121.01 106.43 121.22 106.19 ;
      RECT  121.22 106.43 123.62 106.19 ;
      RECT  123.62 107.53 124.13 107.29 ;
      RECT  122.15 108.32 122.69 107.77 ;
      RECT  121.01 109.04 122.15 109.42 ;
      RECT  123.41 108.8 123.62 108.87 ;
      RECT  123.62 109.66 124.13 109.9 ;
      RECT  121.22 108.56 123.62 108.8 ;
      RECT  123.62 108.8 123.82 108.87 ;
      RECT  123.41 109.59 123.62 109.66 ;
      RECT  124.13 108.56 124.34 108.8 ;
      POLYGON  122.69 109.04 122.69 109.42 123.24 109.42 123.24 109.35 123.62 109.35 123.62 109.11 123.24 109.11 123.24 109.04 122.69 109.04 ;
      RECT  124.13 109.04 124.34 109.42 ;
      RECT  121.01 107.77 121.22 108.32 ;
      RECT  121.22 107.77 122.15 108.32 ;
      RECT  122.15 109.04 122.69 109.42 ;
      RECT  124.13 109.66 124.34 109.9 ;
      RECT  122.69 107.77 124.34 108.32 ;
      RECT  121.01 108.56 121.22 108.8 ;
      RECT  123.62 109.59 123.82 109.66 ;
      POLYGON  123.99 109.04 123.99 109.11 123.62 109.11 123.62 109.35 123.99 109.35 123.99 109.42 124.13 109.42 124.13 109.04 123.99 109.04 ;
      RECT  121.01 109.66 121.22 109.9 ;
      RECT  121.22 109.66 123.62 109.9 ;
      RECT  123.62 108.56 124.13 108.8 ;
      RECT  122.15 107.77 122.69 108.32 ;
      RECT  121.01 111.0 122.15 110.62 ;
      RECT  123.41 111.24 123.62 111.17 ;
      RECT  123.62 110.38 124.13 110.14 ;
      RECT  121.22 111.48 123.62 111.24 ;
      RECT  123.62 111.24 123.82 111.17 ;
      RECT  123.41 110.45 123.62 110.38 ;
      RECT  124.13 111.48 124.34 111.24 ;
      POLYGON  122.69 111.0 122.69 110.62 123.24 110.62 123.24 110.69 123.62 110.69 123.62 110.93 123.24 110.93 123.24 111.0 122.69 111.0 ;
      RECT  124.13 111.0 124.34 110.62 ;
      RECT  121.01 112.27 121.22 111.72 ;
      RECT  121.22 112.27 122.15 111.72 ;
      RECT  122.15 111.0 122.69 110.62 ;
      RECT  124.13 110.38 124.34 110.14 ;
      RECT  122.69 112.27 124.34 111.72 ;
      RECT  121.01 111.48 121.22 111.24 ;
      RECT  123.62 110.45 123.82 110.38 ;
      POLYGON  123.99 111.0 123.99 110.93 123.62 110.93 123.62 110.69 123.99 110.69 123.99 110.62 124.13 110.62 124.13 111.0 123.99 111.0 ;
      RECT  121.01 110.38 121.22 110.14 ;
      RECT  121.22 110.38 123.62 110.14 ;
      RECT  123.62 111.48 124.13 111.24 ;
      RECT  122.15 112.27 122.69 111.72 ;
      RECT  121.01 112.99 122.15 113.37 ;
      RECT  123.41 112.75 123.62 112.82 ;
      RECT  123.62 113.61 124.13 113.85 ;
      RECT  121.22 112.51 123.62 112.75 ;
      RECT  123.62 112.75 123.82 112.82 ;
      RECT  123.41 113.54 123.62 113.61 ;
      RECT  124.13 112.51 124.34 112.75 ;
      POLYGON  122.69 112.99 122.69 113.37 123.24 113.37 123.24 113.3 123.62 113.3 123.62 113.06 123.24 113.06 123.24 112.99 122.69 112.99 ;
      RECT  124.13 112.99 124.34 113.37 ;
      RECT  121.01 111.72 121.22 112.27 ;
      RECT  121.22 111.72 122.15 112.27 ;
      RECT  122.15 112.99 122.69 113.37 ;
      RECT  124.13 113.61 124.34 113.85 ;
      RECT  122.69 111.72 124.34 112.27 ;
      RECT  121.01 112.51 121.22 112.75 ;
      RECT  123.62 113.54 123.82 113.61 ;
      POLYGON  123.99 112.99 123.99 113.06 123.62 113.06 123.62 113.3 123.99 113.3 123.99 113.37 124.13 113.37 124.13 112.99 123.99 112.99 ;
      RECT  121.01 113.61 121.22 113.85 ;
      RECT  121.22 113.61 123.62 113.85 ;
      RECT  123.62 112.51 124.13 112.75 ;
      RECT  122.15 111.72 122.69 112.27 ;
      RECT  121.01 114.95 122.15 114.57 ;
      RECT  123.41 115.19 123.62 115.12 ;
      RECT  123.62 114.33 124.13 114.09 ;
      RECT  121.22 115.43 123.62 115.19 ;
      RECT  123.62 115.19 123.82 115.12 ;
      RECT  123.41 114.4 123.62 114.33 ;
      RECT  124.13 115.43 124.34 115.19 ;
      POLYGON  122.69 114.95 122.69 114.57 123.24 114.57 123.24 114.64 123.62 114.64 123.62 114.88 123.24 114.88 123.24 114.95 122.69 114.95 ;
      RECT  124.13 114.95 124.34 114.57 ;
      RECT  121.01 116.22 121.22 115.67 ;
      RECT  121.22 116.22 122.15 115.67 ;
      RECT  122.15 114.95 122.69 114.57 ;
      RECT  124.13 114.33 124.34 114.09 ;
      RECT  122.69 116.22 124.34 115.67 ;
      RECT  121.01 115.43 121.22 115.19 ;
      RECT  123.62 114.4 123.82 114.33 ;
      POLYGON  123.99 114.95 123.99 114.88 123.62 114.88 123.62 114.64 123.99 114.64 123.99 114.57 124.13 114.57 124.13 114.95 123.99 114.95 ;
      RECT  121.01 114.33 121.22 114.09 ;
      RECT  121.22 114.33 123.62 114.09 ;
      RECT  123.62 115.43 124.13 115.19 ;
      RECT  122.15 116.22 122.69 115.67 ;
      RECT  121.01 116.94 122.15 117.32 ;
      RECT  123.41 116.7 123.62 116.77 ;
      RECT  123.62 117.56 124.13 117.8 ;
      RECT  121.22 116.46 123.62 116.7 ;
      RECT  123.62 116.7 123.82 116.77 ;
      RECT  123.41 117.49 123.62 117.56 ;
      RECT  124.13 116.46 124.34 116.7 ;
      POLYGON  122.69 116.94 122.69 117.32 123.24 117.32 123.24 117.25 123.62 117.25 123.62 117.01 123.24 117.01 123.24 116.94 122.69 116.94 ;
      RECT  124.13 116.94 124.34 117.32 ;
      RECT  121.01 115.67 121.22 116.22 ;
      RECT  121.22 115.67 122.15 116.22 ;
      RECT  122.15 116.94 122.69 117.32 ;
      RECT  124.13 117.56 124.34 117.8 ;
      RECT  122.69 115.67 124.34 116.22 ;
      RECT  121.01 116.46 121.22 116.7 ;
      RECT  123.62 117.49 123.82 117.56 ;
      POLYGON  123.99 116.94 123.99 117.01 123.62 117.01 123.62 117.25 123.99 117.25 123.99 117.32 124.13 117.32 124.13 116.94 123.99 116.94 ;
      RECT  121.01 117.56 121.22 117.8 ;
      RECT  121.22 117.56 123.62 117.8 ;
      RECT  123.62 116.46 124.13 116.7 ;
      RECT  122.15 115.67 122.69 116.22 ;
      RECT  121.01 118.9 122.15 118.52 ;
      RECT  123.41 119.14 123.62 119.07 ;
      RECT  123.62 118.28 124.13 118.04 ;
      RECT  121.22 119.38 123.62 119.14 ;
      RECT  123.62 119.14 123.82 119.07 ;
      RECT  123.41 118.35 123.62 118.28 ;
      RECT  124.13 119.38 124.34 119.14 ;
      POLYGON  122.69 118.9 122.69 118.52 123.24 118.52 123.24 118.59 123.62 118.59 123.62 118.83 123.24 118.83 123.24 118.9 122.69 118.9 ;
      RECT  124.13 118.9 124.34 118.52 ;
      RECT  121.01 120.17 121.22 119.62 ;
      RECT  121.22 120.17 122.15 119.62 ;
      RECT  122.15 118.9 122.69 118.52 ;
      RECT  124.13 118.28 124.34 118.04 ;
      RECT  122.69 120.17 124.34 119.62 ;
      RECT  121.01 119.38 121.22 119.14 ;
      RECT  123.62 118.35 123.82 118.28 ;
      POLYGON  123.99 118.9 123.99 118.83 123.62 118.83 123.62 118.59 123.99 118.59 123.99 118.52 124.13 118.52 124.13 118.9 123.99 118.9 ;
      RECT  121.01 118.28 121.22 118.04 ;
      RECT  121.22 118.28 123.62 118.04 ;
      RECT  123.62 119.38 124.13 119.14 ;
      RECT  122.15 120.17 122.69 119.62 ;
      RECT  121.01 120.89 122.15 121.27 ;
      RECT  123.41 120.65 123.62 120.72 ;
      RECT  123.62 121.51 124.13 121.75 ;
      RECT  121.22 120.41 123.62 120.65 ;
      RECT  123.62 120.65 123.82 120.72 ;
      RECT  123.41 121.44 123.62 121.51 ;
      RECT  124.13 120.41 124.34 120.65 ;
      POLYGON  122.69 120.89 122.69 121.27 123.24 121.27 123.24 121.2 123.62 121.2 123.62 120.96 123.24 120.96 123.24 120.89 122.69 120.89 ;
      RECT  124.13 120.89 124.34 121.27 ;
      RECT  121.01 119.62 121.22 120.17 ;
      RECT  121.22 119.62 122.15 120.17 ;
      RECT  122.15 120.89 122.69 121.27 ;
      RECT  124.13 121.51 124.34 121.75 ;
      RECT  122.69 119.62 124.34 120.17 ;
      RECT  121.01 120.41 121.22 120.65 ;
      RECT  123.62 121.44 123.82 121.51 ;
      POLYGON  123.99 120.89 123.99 120.96 123.62 120.96 123.62 121.2 123.99 121.2 123.99 121.27 124.13 121.27 124.13 120.89 123.99 120.89 ;
      RECT  121.01 121.51 121.22 121.75 ;
      RECT  121.22 121.51 123.62 121.75 ;
      RECT  123.62 120.41 124.13 120.65 ;
      RECT  122.15 119.62 122.69 120.17 ;
      RECT  121.01 122.85 122.15 122.47 ;
      RECT  123.41 123.09 123.62 123.02 ;
      RECT  123.62 122.23 124.13 121.99 ;
      RECT  121.22 123.33 123.62 123.09 ;
      RECT  123.62 123.09 123.82 123.02 ;
      RECT  123.41 122.3 123.62 122.23 ;
      RECT  124.13 123.33 124.34 123.09 ;
      POLYGON  122.69 122.85 122.69 122.47 123.24 122.47 123.24 122.54 123.62 122.54 123.62 122.78 123.24 122.78 123.24 122.85 122.69 122.85 ;
      RECT  124.13 122.85 124.34 122.47 ;
      RECT  121.01 124.12 121.22 123.57 ;
      RECT  121.22 124.12 122.15 123.57 ;
      RECT  122.15 122.85 122.69 122.47 ;
      RECT  124.13 122.23 124.34 121.99 ;
      RECT  122.69 124.12 124.34 123.57 ;
      RECT  121.01 123.33 121.22 123.09 ;
      RECT  123.62 122.3 123.82 122.23 ;
      POLYGON  123.99 122.85 123.99 122.78 123.62 122.78 123.62 122.54 123.99 122.54 123.99 122.47 124.13 122.47 124.13 122.85 123.99 122.85 ;
      RECT  121.01 122.23 121.22 121.99 ;
      RECT  121.22 122.23 123.62 121.99 ;
      RECT  123.62 123.33 124.13 123.09 ;
      RECT  122.15 124.12 122.69 123.57 ;
      RECT  127.67 93.24 126.53 93.62 ;
      RECT  125.27 93.0 125.06 93.07 ;
      RECT  125.06 93.86 124.55 94.1 ;
      RECT  127.46 92.76 125.06 93.0 ;
      RECT  125.06 93.0 124.86 93.07 ;
      RECT  125.27 93.79 125.06 93.86 ;
      RECT  124.55 92.76 124.34 93.0 ;
      POLYGON  125.99 93.24 125.99 93.62 125.44 93.62 125.44 93.55 125.06 93.55 125.06 93.31 125.44 93.31 125.44 93.24 125.99 93.24 ;
      RECT  124.55 93.24 124.34 93.62 ;
      RECT  127.67 91.97 127.46 92.52 ;
      RECT  127.46 91.97 126.53 92.52 ;
      RECT  126.53 93.24 125.99 93.62 ;
      RECT  124.55 93.86 124.34 94.1 ;
      RECT  125.99 91.97 124.34 92.52 ;
      RECT  127.67 92.76 127.46 93.0 ;
      RECT  125.06 93.79 124.86 93.86 ;
      POLYGON  124.69 93.24 124.69 93.31 125.06 93.31 125.06 93.55 124.69 93.55 124.69 93.62 124.55 93.62 124.55 93.24 124.69 93.24 ;
      RECT  127.67 93.86 127.46 94.1 ;
      RECT  127.46 93.86 125.06 94.1 ;
      RECT  125.06 92.76 124.55 93.0 ;
      RECT  126.53 91.97 125.99 92.52 ;
      RECT  127.67 95.2 126.53 94.82 ;
      RECT  125.27 95.44 125.06 95.37 ;
      RECT  125.06 94.58 124.55 94.34 ;
      RECT  127.46 95.68 125.06 95.44 ;
      RECT  125.06 95.44 124.86 95.37 ;
      RECT  125.27 94.65 125.06 94.58 ;
      RECT  124.55 95.68 124.34 95.44 ;
      POLYGON  125.99 95.2 125.99 94.82 125.44 94.82 125.44 94.89 125.06 94.89 125.06 95.13 125.44 95.13 125.44 95.2 125.99 95.2 ;
      RECT  124.55 95.2 124.34 94.82 ;
      RECT  127.67 96.47 127.46 95.92 ;
      RECT  127.46 96.47 126.53 95.92 ;
      RECT  126.53 95.2 125.99 94.82 ;
      RECT  124.55 94.58 124.34 94.34 ;
      RECT  125.99 96.47 124.34 95.92 ;
      RECT  127.67 95.68 127.46 95.44 ;
      RECT  125.06 94.65 124.86 94.58 ;
      POLYGON  124.69 95.2 124.69 95.13 125.06 95.13 125.06 94.89 124.69 94.89 124.69 94.82 124.55 94.82 124.55 95.2 124.69 95.2 ;
      RECT  127.67 94.58 127.46 94.34 ;
      RECT  127.46 94.58 125.06 94.34 ;
      RECT  125.06 95.68 124.55 95.44 ;
      RECT  126.53 96.47 125.99 95.92 ;
      RECT  127.67 97.19 126.53 97.57 ;
      RECT  125.27 96.95 125.06 97.02 ;
      RECT  125.06 97.81 124.55 98.05 ;
      RECT  127.46 96.71 125.06 96.95 ;
      RECT  125.06 96.95 124.86 97.02 ;
      RECT  125.27 97.74 125.06 97.81 ;
      RECT  124.55 96.71 124.34 96.95 ;
      POLYGON  125.99 97.19 125.99 97.57 125.44 97.57 125.44 97.5 125.06 97.5 125.06 97.26 125.44 97.26 125.44 97.19 125.99 97.19 ;
      RECT  124.55 97.19 124.34 97.57 ;
      RECT  127.67 95.92 127.46 96.47 ;
      RECT  127.46 95.92 126.53 96.47 ;
      RECT  126.53 97.19 125.99 97.57 ;
      RECT  124.55 97.81 124.34 98.05 ;
      RECT  125.99 95.92 124.34 96.47 ;
      RECT  127.67 96.71 127.46 96.95 ;
      RECT  125.06 97.74 124.86 97.81 ;
      POLYGON  124.69 97.19 124.69 97.26 125.06 97.26 125.06 97.5 124.69 97.5 124.69 97.57 124.55 97.57 124.55 97.19 124.69 97.19 ;
      RECT  127.67 97.81 127.46 98.05 ;
      RECT  127.46 97.81 125.06 98.05 ;
      RECT  125.06 96.71 124.55 96.95 ;
      RECT  126.53 95.92 125.99 96.47 ;
      RECT  127.67 99.15 126.53 98.77 ;
      RECT  125.27 99.39 125.06 99.32 ;
      RECT  125.06 98.53 124.55 98.29 ;
      RECT  127.46 99.63 125.06 99.39 ;
      RECT  125.06 99.39 124.86 99.32 ;
      RECT  125.27 98.6 125.06 98.53 ;
      RECT  124.55 99.63 124.34 99.39 ;
      POLYGON  125.99 99.15 125.99 98.77 125.44 98.77 125.44 98.84 125.06 98.84 125.06 99.08 125.44 99.08 125.44 99.15 125.99 99.15 ;
      RECT  124.55 99.15 124.34 98.77 ;
      RECT  127.67 100.42 127.46 99.87 ;
      RECT  127.46 100.42 126.53 99.87 ;
      RECT  126.53 99.15 125.99 98.77 ;
      RECT  124.55 98.53 124.34 98.29 ;
      RECT  125.99 100.42 124.34 99.87 ;
      RECT  127.67 99.63 127.46 99.39 ;
      RECT  125.06 98.6 124.86 98.53 ;
      POLYGON  124.69 99.15 124.69 99.08 125.06 99.08 125.06 98.84 124.69 98.84 124.69 98.77 124.55 98.77 124.55 99.15 124.69 99.15 ;
      RECT  127.67 98.53 127.46 98.29 ;
      RECT  127.46 98.53 125.06 98.29 ;
      RECT  125.06 99.63 124.55 99.39 ;
      RECT  126.53 100.42 125.99 99.87 ;
      RECT  127.67 101.14 126.53 101.52 ;
      RECT  125.27 100.9 125.06 100.97 ;
      RECT  125.06 101.76 124.55 102.0 ;
      RECT  127.46 100.66 125.06 100.9 ;
      RECT  125.06 100.9 124.86 100.97 ;
      RECT  125.27 101.69 125.06 101.76 ;
      RECT  124.55 100.66 124.34 100.9 ;
      POLYGON  125.99 101.14 125.99 101.52 125.44 101.52 125.44 101.45 125.06 101.45 125.06 101.21 125.44 101.21 125.44 101.14 125.99 101.14 ;
      RECT  124.55 101.14 124.34 101.52 ;
      RECT  127.67 99.87 127.46 100.42 ;
      RECT  127.46 99.87 126.53 100.42 ;
      RECT  126.53 101.14 125.99 101.52 ;
      RECT  124.55 101.76 124.34 102.0 ;
      RECT  125.99 99.87 124.34 100.42 ;
      RECT  127.67 100.66 127.46 100.9 ;
      RECT  125.06 101.69 124.86 101.76 ;
      POLYGON  124.69 101.14 124.69 101.21 125.06 101.21 125.06 101.45 124.69 101.45 124.69 101.52 124.55 101.52 124.55 101.14 124.69 101.14 ;
      RECT  127.67 101.76 127.46 102.0 ;
      RECT  127.46 101.76 125.06 102.0 ;
      RECT  125.06 100.66 124.55 100.9 ;
      RECT  126.53 99.87 125.99 100.42 ;
      RECT  127.67 103.1 126.53 102.72 ;
      RECT  125.27 103.34 125.06 103.27 ;
      RECT  125.06 102.48 124.55 102.24 ;
      RECT  127.46 103.58 125.06 103.34 ;
      RECT  125.06 103.34 124.86 103.27 ;
      RECT  125.27 102.55 125.06 102.48 ;
      RECT  124.55 103.58 124.34 103.34 ;
      POLYGON  125.99 103.1 125.99 102.72 125.44 102.72 125.44 102.79 125.06 102.79 125.06 103.03 125.44 103.03 125.44 103.1 125.99 103.1 ;
      RECT  124.55 103.1 124.34 102.72 ;
      RECT  127.67 104.37 127.46 103.82 ;
      RECT  127.46 104.37 126.53 103.82 ;
      RECT  126.53 103.1 125.99 102.72 ;
      RECT  124.55 102.48 124.34 102.24 ;
      RECT  125.99 104.37 124.34 103.82 ;
      RECT  127.67 103.58 127.46 103.34 ;
      RECT  125.06 102.55 124.86 102.48 ;
      POLYGON  124.69 103.1 124.69 103.03 125.06 103.03 125.06 102.79 124.69 102.79 124.69 102.72 124.55 102.72 124.55 103.1 124.69 103.1 ;
      RECT  127.67 102.48 127.46 102.24 ;
      RECT  127.46 102.48 125.06 102.24 ;
      RECT  125.06 103.58 124.55 103.34 ;
      RECT  126.53 104.37 125.99 103.82 ;
      RECT  127.67 105.09 126.53 105.47 ;
      RECT  125.27 104.85 125.06 104.92 ;
      RECT  125.06 105.71 124.55 105.95 ;
      RECT  127.46 104.61 125.06 104.85 ;
      RECT  125.06 104.85 124.86 104.92 ;
      RECT  125.27 105.64 125.06 105.71 ;
      RECT  124.55 104.61 124.34 104.85 ;
      POLYGON  125.99 105.09 125.99 105.47 125.44 105.47 125.44 105.4 125.06 105.4 125.06 105.16 125.44 105.16 125.44 105.09 125.99 105.09 ;
      RECT  124.55 105.09 124.34 105.47 ;
      RECT  127.67 103.82 127.46 104.37 ;
      RECT  127.46 103.82 126.53 104.37 ;
      RECT  126.53 105.09 125.99 105.47 ;
      RECT  124.55 105.71 124.34 105.95 ;
      RECT  125.99 103.82 124.34 104.37 ;
      RECT  127.67 104.61 127.46 104.85 ;
      RECT  125.06 105.64 124.86 105.71 ;
      POLYGON  124.69 105.09 124.69 105.16 125.06 105.16 125.06 105.4 124.69 105.4 124.69 105.47 124.55 105.47 124.55 105.09 124.69 105.09 ;
      RECT  127.67 105.71 127.46 105.95 ;
      RECT  127.46 105.71 125.06 105.95 ;
      RECT  125.06 104.61 124.55 104.85 ;
      RECT  126.53 103.82 125.99 104.37 ;
      RECT  127.67 107.05 126.53 106.67 ;
      RECT  125.27 107.29 125.06 107.22 ;
      RECT  125.06 106.43 124.55 106.19 ;
      RECT  127.46 107.53 125.06 107.29 ;
      RECT  125.06 107.29 124.86 107.22 ;
      RECT  125.27 106.5 125.06 106.43 ;
      RECT  124.55 107.53 124.34 107.29 ;
      POLYGON  125.99 107.05 125.99 106.67 125.44 106.67 125.44 106.74 125.06 106.74 125.06 106.98 125.44 106.98 125.44 107.05 125.99 107.05 ;
      RECT  124.55 107.05 124.34 106.67 ;
      RECT  127.67 108.32 127.46 107.77 ;
      RECT  127.46 108.32 126.53 107.77 ;
      RECT  126.53 107.05 125.99 106.67 ;
      RECT  124.55 106.43 124.34 106.19 ;
      RECT  125.99 108.32 124.34 107.77 ;
      RECT  127.67 107.53 127.46 107.29 ;
      RECT  125.06 106.5 124.86 106.43 ;
      POLYGON  124.69 107.05 124.69 106.98 125.06 106.98 125.06 106.74 124.69 106.74 124.69 106.67 124.55 106.67 124.55 107.05 124.69 107.05 ;
      RECT  127.67 106.43 127.46 106.19 ;
      RECT  127.46 106.43 125.06 106.19 ;
      RECT  125.06 107.53 124.55 107.29 ;
      RECT  126.53 108.32 125.99 107.77 ;
      RECT  127.67 109.04 126.53 109.42 ;
      RECT  125.27 108.8 125.06 108.87 ;
      RECT  125.06 109.66 124.55 109.9 ;
      RECT  127.46 108.56 125.06 108.8 ;
      RECT  125.06 108.8 124.86 108.87 ;
      RECT  125.27 109.59 125.06 109.66 ;
      RECT  124.55 108.56 124.34 108.8 ;
      POLYGON  125.99 109.04 125.99 109.42 125.44 109.42 125.44 109.35 125.06 109.35 125.06 109.11 125.44 109.11 125.44 109.04 125.99 109.04 ;
      RECT  124.55 109.04 124.34 109.42 ;
      RECT  127.67 107.77 127.46 108.32 ;
      RECT  127.46 107.77 126.53 108.32 ;
      RECT  126.53 109.04 125.99 109.42 ;
      RECT  124.55 109.66 124.34 109.9 ;
      RECT  125.99 107.77 124.34 108.32 ;
      RECT  127.67 108.56 127.46 108.8 ;
      RECT  125.06 109.59 124.86 109.66 ;
      POLYGON  124.69 109.04 124.69 109.11 125.06 109.11 125.06 109.35 124.69 109.35 124.69 109.42 124.55 109.42 124.55 109.04 124.69 109.04 ;
      RECT  127.67 109.66 127.46 109.9 ;
      RECT  127.46 109.66 125.06 109.9 ;
      RECT  125.06 108.56 124.55 108.8 ;
      RECT  126.53 107.77 125.99 108.32 ;
      RECT  127.67 111.0 126.53 110.62 ;
      RECT  125.27 111.24 125.06 111.17 ;
      RECT  125.06 110.38 124.55 110.14 ;
      RECT  127.46 111.48 125.06 111.24 ;
      RECT  125.06 111.24 124.86 111.17 ;
      RECT  125.27 110.45 125.06 110.38 ;
      RECT  124.55 111.48 124.34 111.24 ;
      POLYGON  125.99 111.0 125.99 110.62 125.44 110.62 125.44 110.69 125.06 110.69 125.06 110.93 125.44 110.93 125.44 111.0 125.99 111.0 ;
      RECT  124.55 111.0 124.34 110.62 ;
      RECT  127.67 112.27 127.46 111.72 ;
      RECT  127.46 112.27 126.53 111.72 ;
      RECT  126.53 111.0 125.99 110.62 ;
      RECT  124.55 110.38 124.34 110.14 ;
      RECT  125.99 112.27 124.34 111.72 ;
      RECT  127.67 111.48 127.46 111.24 ;
      RECT  125.06 110.45 124.86 110.38 ;
      POLYGON  124.69 111.0 124.69 110.93 125.06 110.93 125.06 110.69 124.69 110.69 124.69 110.62 124.55 110.62 124.55 111.0 124.69 111.0 ;
      RECT  127.67 110.38 127.46 110.14 ;
      RECT  127.46 110.38 125.06 110.14 ;
      RECT  125.06 111.48 124.55 111.24 ;
      RECT  126.53 112.27 125.99 111.72 ;
      RECT  127.67 112.99 126.53 113.37 ;
      RECT  125.27 112.75 125.06 112.82 ;
      RECT  125.06 113.61 124.55 113.85 ;
      RECT  127.46 112.51 125.06 112.75 ;
      RECT  125.06 112.75 124.86 112.82 ;
      RECT  125.27 113.54 125.06 113.61 ;
      RECT  124.55 112.51 124.34 112.75 ;
      POLYGON  125.99 112.99 125.99 113.37 125.44 113.37 125.44 113.3 125.06 113.3 125.06 113.06 125.44 113.06 125.44 112.99 125.99 112.99 ;
      RECT  124.55 112.99 124.34 113.37 ;
      RECT  127.67 111.72 127.46 112.27 ;
      RECT  127.46 111.72 126.53 112.27 ;
      RECT  126.53 112.99 125.99 113.37 ;
      RECT  124.55 113.61 124.34 113.85 ;
      RECT  125.99 111.72 124.34 112.27 ;
      RECT  127.67 112.51 127.46 112.75 ;
      RECT  125.06 113.54 124.86 113.61 ;
      POLYGON  124.69 112.99 124.69 113.06 125.06 113.06 125.06 113.3 124.69 113.3 124.69 113.37 124.55 113.37 124.55 112.99 124.69 112.99 ;
      RECT  127.67 113.61 127.46 113.85 ;
      RECT  127.46 113.61 125.06 113.85 ;
      RECT  125.06 112.51 124.55 112.75 ;
      RECT  126.53 111.72 125.99 112.27 ;
      RECT  127.67 114.95 126.53 114.57 ;
      RECT  125.27 115.19 125.06 115.12 ;
      RECT  125.06 114.33 124.55 114.09 ;
      RECT  127.46 115.43 125.06 115.19 ;
      RECT  125.06 115.19 124.86 115.12 ;
      RECT  125.27 114.4 125.06 114.33 ;
      RECT  124.55 115.43 124.34 115.19 ;
      POLYGON  125.99 114.95 125.99 114.57 125.44 114.57 125.44 114.64 125.06 114.64 125.06 114.88 125.44 114.88 125.44 114.95 125.99 114.95 ;
      RECT  124.55 114.95 124.34 114.57 ;
      RECT  127.67 116.22 127.46 115.67 ;
      RECT  127.46 116.22 126.53 115.67 ;
      RECT  126.53 114.95 125.99 114.57 ;
      RECT  124.55 114.33 124.34 114.09 ;
      RECT  125.99 116.22 124.34 115.67 ;
      RECT  127.67 115.43 127.46 115.19 ;
      RECT  125.06 114.4 124.86 114.33 ;
      POLYGON  124.69 114.95 124.69 114.88 125.06 114.88 125.06 114.64 124.69 114.64 124.69 114.57 124.55 114.57 124.55 114.95 124.69 114.95 ;
      RECT  127.67 114.33 127.46 114.09 ;
      RECT  127.46 114.33 125.06 114.09 ;
      RECT  125.06 115.43 124.55 115.19 ;
      RECT  126.53 116.22 125.99 115.67 ;
      RECT  127.67 116.94 126.53 117.32 ;
      RECT  125.27 116.7 125.06 116.77 ;
      RECT  125.06 117.56 124.55 117.8 ;
      RECT  127.46 116.46 125.06 116.7 ;
      RECT  125.06 116.7 124.86 116.77 ;
      RECT  125.27 117.49 125.06 117.56 ;
      RECT  124.55 116.46 124.34 116.7 ;
      POLYGON  125.99 116.94 125.99 117.32 125.44 117.32 125.44 117.25 125.06 117.25 125.06 117.01 125.44 117.01 125.44 116.94 125.99 116.94 ;
      RECT  124.55 116.94 124.34 117.32 ;
      RECT  127.67 115.67 127.46 116.22 ;
      RECT  127.46 115.67 126.53 116.22 ;
      RECT  126.53 116.94 125.99 117.32 ;
      RECT  124.55 117.56 124.34 117.8 ;
      RECT  125.99 115.67 124.34 116.22 ;
      RECT  127.67 116.46 127.46 116.7 ;
      RECT  125.06 117.49 124.86 117.56 ;
      POLYGON  124.69 116.94 124.69 117.01 125.06 117.01 125.06 117.25 124.69 117.25 124.69 117.32 124.55 117.32 124.55 116.94 124.69 116.94 ;
      RECT  127.67 117.56 127.46 117.8 ;
      RECT  127.46 117.56 125.06 117.8 ;
      RECT  125.06 116.46 124.55 116.7 ;
      RECT  126.53 115.67 125.99 116.22 ;
      RECT  127.67 118.9 126.53 118.52 ;
      RECT  125.27 119.14 125.06 119.07 ;
      RECT  125.06 118.28 124.55 118.04 ;
      RECT  127.46 119.38 125.06 119.14 ;
      RECT  125.06 119.14 124.86 119.07 ;
      RECT  125.27 118.35 125.06 118.28 ;
      RECT  124.55 119.38 124.34 119.14 ;
      POLYGON  125.99 118.9 125.99 118.52 125.44 118.52 125.44 118.59 125.06 118.59 125.06 118.83 125.44 118.83 125.44 118.9 125.99 118.9 ;
      RECT  124.55 118.9 124.34 118.52 ;
      RECT  127.67 120.17 127.46 119.62 ;
      RECT  127.46 120.17 126.53 119.62 ;
      RECT  126.53 118.9 125.99 118.52 ;
      RECT  124.55 118.28 124.34 118.04 ;
      RECT  125.99 120.17 124.34 119.62 ;
      RECT  127.67 119.38 127.46 119.14 ;
      RECT  125.06 118.35 124.86 118.28 ;
      POLYGON  124.69 118.9 124.69 118.83 125.06 118.83 125.06 118.59 124.69 118.59 124.69 118.52 124.55 118.52 124.55 118.9 124.69 118.9 ;
      RECT  127.67 118.28 127.46 118.04 ;
      RECT  127.46 118.28 125.06 118.04 ;
      RECT  125.06 119.38 124.55 119.14 ;
      RECT  126.53 120.17 125.99 119.62 ;
      RECT  127.67 120.89 126.53 121.27 ;
      RECT  125.27 120.65 125.06 120.72 ;
      RECT  125.06 121.51 124.55 121.75 ;
      RECT  127.46 120.41 125.06 120.65 ;
      RECT  125.06 120.65 124.86 120.72 ;
      RECT  125.27 121.44 125.06 121.51 ;
      RECT  124.55 120.41 124.34 120.65 ;
      POLYGON  125.99 120.89 125.99 121.27 125.44 121.27 125.44 121.2 125.06 121.2 125.06 120.96 125.44 120.96 125.44 120.89 125.99 120.89 ;
      RECT  124.55 120.89 124.34 121.27 ;
      RECT  127.67 119.62 127.46 120.17 ;
      RECT  127.46 119.62 126.53 120.17 ;
      RECT  126.53 120.89 125.99 121.27 ;
      RECT  124.55 121.51 124.34 121.75 ;
      RECT  125.99 119.62 124.34 120.17 ;
      RECT  127.67 120.41 127.46 120.65 ;
      RECT  125.06 121.44 124.86 121.51 ;
      POLYGON  124.69 120.89 124.69 120.96 125.06 120.96 125.06 121.2 124.69 121.2 124.69 121.27 124.55 121.27 124.55 120.89 124.69 120.89 ;
      RECT  127.67 121.51 127.46 121.75 ;
      RECT  127.46 121.51 125.06 121.75 ;
      RECT  125.06 120.41 124.55 120.65 ;
      RECT  126.53 119.62 125.99 120.17 ;
      RECT  127.67 122.85 126.53 122.47 ;
      RECT  125.27 123.09 125.06 123.02 ;
      RECT  125.06 122.23 124.55 121.99 ;
      RECT  127.46 123.33 125.06 123.09 ;
      RECT  125.06 123.09 124.86 123.02 ;
      RECT  125.27 122.3 125.06 122.23 ;
      RECT  124.55 123.33 124.34 123.09 ;
      POLYGON  125.99 122.85 125.99 122.47 125.44 122.47 125.44 122.54 125.06 122.54 125.06 122.78 125.44 122.78 125.44 122.85 125.99 122.85 ;
      RECT  124.55 122.85 124.34 122.47 ;
      RECT  127.67 124.12 127.46 123.57 ;
      RECT  127.46 124.12 126.53 123.57 ;
      RECT  126.53 122.85 125.99 122.47 ;
      RECT  124.55 122.23 124.34 121.99 ;
      RECT  125.99 124.12 124.34 123.57 ;
      RECT  127.67 123.33 127.46 123.09 ;
      RECT  125.06 122.3 124.86 122.23 ;
      POLYGON  124.69 122.85 124.69 122.78 125.06 122.78 125.06 122.54 124.69 122.54 124.69 122.47 124.55 122.47 124.55 122.85 124.69 122.85 ;
      RECT  127.67 122.23 127.46 121.99 ;
      RECT  127.46 122.23 125.06 121.99 ;
      RECT  125.06 123.33 124.55 123.09 ;
      RECT  126.53 124.12 125.99 123.57 ;
      RECT  127.25 93.24 128.39 93.62 ;
      RECT  129.65 93.0 129.86 93.07 ;
      RECT  129.86 93.86 130.37 94.1 ;
      RECT  127.46 92.76 129.86 93.0 ;
      RECT  129.86 93.0 130.06 93.07 ;
      RECT  129.65 93.79 129.86 93.86 ;
      RECT  130.37 92.76 130.58 93.0 ;
      POLYGON  128.93 93.24 128.93 93.62 129.48 93.62 129.48 93.55 129.86 93.55 129.86 93.31 129.48 93.31 129.48 93.24 128.93 93.24 ;
      RECT  130.37 93.24 130.58 93.62 ;
      RECT  127.25 91.97 127.46 92.52 ;
      RECT  127.46 91.97 128.39 92.52 ;
      RECT  128.39 93.24 128.93 93.62 ;
      RECT  130.37 93.86 130.58 94.1 ;
      RECT  128.93 91.97 130.58 92.52 ;
      RECT  127.25 92.76 127.46 93.0 ;
      RECT  129.86 93.79 130.06 93.86 ;
      POLYGON  130.23 93.24 130.23 93.31 129.86 93.31 129.86 93.55 130.23 93.55 130.23 93.62 130.37 93.62 130.37 93.24 130.23 93.24 ;
      RECT  127.25 93.86 127.46 94.1 ;
      RECT  127.46 93.86 129.86 94.1 ;
      RECT  129.86 92.76 130.37 93.0 ;
      RECT  128.39 91.97 128.93 92.52 ;
      RECT  127.25 95.2 128.39 94.82 ;
      RECT  129.65 95.44 129.86 95.37 ;
      RECT  129.86 94.58 130.37 94.34 ;
      RECT  127.46 95.68 129.86 95.44 ;
      RECT  129.86 95.44 130.06 95.37 ;
      RECT  129.65 94.65 129.86 94.58 ;
      RECT  130.37 95.68 130.58 95.44 ;
      POLYGON  128.93 95.2 128.93 94.82 129.48 94.82 129.48 94.89 129.86 94.89 129.86 95.13 129.48 95.13 129.48 95.2 128.93 95.2 ;
      RECT  130.37 95.2 130.58 94.82 ;
      RECT  127.25 96.47 127.46 95.92 ;
      RECT  127.46 96.47 128.39 95.92 ;
      RECT  128.39 95.2 128.93 94.82 ;
      RECT  130.37 94.58 130.58 94.34 ;
      RECT  128.93 96.47 130.58 95.92 ;
      RECT  127.25 95.68 127.46 95.44 ;
      RECT  129.86 94.65 130.06 94.58 ;
      POLYGON  130.23 95.2 130.23 95.13 129.86 95.13 129.86 94.89 130.23 94.89 130.23 94.82 130.37 94.82 130.37 95.2 130.23 95.2 ;
      RECT  127.25 94.58 127.46 94.34 ;
      RECT  127.46 94.58 129.86 94.34 ;
      RECT  129.86 95.68 130.37 95.44 ;
      RECT  128.39 96.47 128.93 95.92 ;
      RECT  127.25 97.19 128.39 97.57 ;
      RECT  129.65 96.95 129.86 97.02 ;
      RECT  129.86 97.81 130.37 98.05 ;
      RECT  127.46 96.71 129.86 96.95 ;
      RECT  129.86 96.95 130.06 97.02 ;
      RECT  129.65 97.74 129.86 97.81 ;
      RECT  130.37 96.71 130.58 96.95 ;
      POLYGON  128.93 97.19 128.93 97.57 129.48 97.57 129.48 97.5 129.86 97.5 129.86 97.26 129.48 97.26 129.48 97.19 128.93 97.19 ;
      RECT  130.37 97.19 130.58 97.57 ;
      RECT  127.25 95.92 127.46 96.47 ;
      RECT  127.46 95.92 128.39 96.47 ;
      RECT  128.39 97.19 128.93 97.57 ;
      RECT  130.37 97.81 130.58 98.05 ;
      RECT  128.93 95.92 130.58 96.47 ;
      RECT  127.25 96.71 127.46 96.95 ;
      RECT  129.86 97.74 130.06 97.81 ;
      POLYGON  130.23 97.19 130.23 97.26 129.86 97.26 129.86 97.5 130.23 97.5 130.23 97.57 130.37 97.57 130.37 97.19 130.23 97.19 ;
      RECT  127.25 97.81 127.46 98.05 ;
      RECT  127.46 97.81 129.86 98.05 ;
      RECT  129.86 96.71 130.37 96.95 ;
      RECT  128.39 95.92 128.93 96.47 ;
      RECT  127.25 99.15 128.39 98.77 ;
      RECT  129.65 99.39 129.86 99.32 ;
      RECT  129.86 98.53 130.37 98.29 ;
      RECT  127.46 99.63 129.86 99.39 ;
      RECT  129.86 99.39 130.06 99.32 ;
      RECT  129.65 98.6 129.86 98.53 ;
      RECT  130.37 99.63 130.58 99.39 ;
      POLYGON  128.93 99.15 128.93 98.77 129.48 98.77 129.48 98.84 129.86 98.84 129.86 99.08 129.48 99.08 129.48 99.15 128.93 99.15 ;
      RECT  130.37 99.15 130.58 98.77 ;
      RECT  127.25 100.42 127.46 99.87 ;
      RECT  127.46 100.42 128.39 99.87 ;
      RECT  128.39 99.15 128.93 98.77 ;
      RECT  130.37 98.53 130.58 98.29 ;
      RECT  128.93 100.42 130.58 99.87 ;
      RECT  127.25 99.63 127.46 99.39 ;
      RECT  129.86 98.6 130.06 98.53 ;
      POLYGON  130.23 99.15 130.23 99.08 129.86 99.08 129.86 98.84 130.23 98.84 130.23 98.77 130.37 98.77 130.37 99.15 130.23 99.15 ;
      RECT  127.25 98.53 127.46 98.29 ;
      RECT  127.46 98.53 129.86 98.29 ;
      RECT  129.86 99.63 130.37 99.39 ;
      RECT  128.39 100.42 128.93 99.87 ;
      RECT  127.25 101.14 128.39 101.52 ;
      RECT  129.65 100.9 129.86 100.97 ;
      RECT  129.86 101.76 130.37 102.0 ;
      RECT  127.46 100.66 129.86 100.9 ;
      RECT  129.86 100.9 130.06 100.97 ;
      RECT  129.65 101.69 129.86 101.76 ;
      RECT  130.37 100.66 130.58 100.9 ;
      POLYGON  128.93 101.14 128.93 101.52 129.48 101.52 129.48 101.45 129.86 101.45 129.86 101.21 129.48 101.21 129.48 101.14 128.93 101.14 ;
      RECT  130.37 101.14 130.58 101.52 ;
      RECT  127.25 99.87 127.46 100.42 ;
      RECT  127.46 99.87 128.39 100.42 ;
      RECT  128.39 101.14 128.93 101.52 ;
      RECT  130.37 101.76 130.58 102.0 ;
      RECT  128.93 99.87 130.58 100.42 ;
      RECT  127.25 100.66 127.46 100.9 ;
      RECT  129.86 101.69 130.06 101.76 ;
      POLYGON  130.23 101.14 130.23 101.21 129.86 101.21 129.86 101.45 130.23 101.45 130.23 101.52 130.37 101.52 130.37 101.14 130.23 101.14 ;
      RECT  127.25 101.76 127.46 102.0 ;
      RECT  127.46 101.76 129.86 102.0 ;
      RECT  129.86 100.66 130.37 100.9 ;
      RECT  128.39 99.87 128.93 100.42 ;
      RECT  127.25 103.1 128.39 102.72 ;
      RECT  129.65 103.34 129.86 103.27 ;
      RECT  129.86 102.48 130.37 102.24 ;
      RECT  127.46 103.58 129.86 103.34 ;
      RECT  129.86 103.34 130.06 103.27 ;
      RECT  129.65 102.55 129.86 102.48 ;
      RECT  130.37 103.58 130.58 103.34 ;
      POLYGON  128.93 103.1 128.93 102.72 129.48 102.72 129.48 102.79 129.86 102.79 129.86 103.03 129.48 103.03 129.48 103.1 128.93 103.1 ;
      RECT  130.37 103.1 130.58 102.72 ;
      RECT  127.25 104.37 127.46 103.82 ;
      RECT  127.46 104.37 128.39 103.82 ;
      RECT  128.39 103.1 128.93 102.72 ;
      RECT  130.37 102.48 130.58 102.24 ;
      RECT  128.93 104.37 130.58 103.82 ;
      RECT  127.25 103.58 127.46 103.34 ;
      RECT  129.86 102.55 130.06 102.48 ;
      POLYGON  130.23 103.1 130.23 103.03 129.86 103.03 129.86 102.79 130.23 102.79 130.23 102.72 130.37 102.72 130.37 103.1 130.23 103.1 ;
      RECT  127.25 102.48 127.46 102.24 ;
      RECT  127.46 102.48 129.86 102.24 ;
      RECT  129.86 103.58 130.37 103.34 ;
      RECT  128.39 104.37 128.93 103.82 ;
      RECT  127.25 105.09 128.39 105.47 ;
      RECT  129.65 104.85 129.86 104.92 ;
      RECT  129.86 105.71 130.37 105.95 ;
      RECT  127.46 104.61 129.86 104.85 ;
      RECT  129.86 104.85 130.06 104.92 ;
      RECT  129.65 105.64 129.86 105.71 ;
      RECT  130.37 104.61 130.58 104.85 ;
      POLYGON  128.93 105.09 128.93 105.47 129.48 105.47 129.48 105.4 129.86 105.4 129.86 105.16 129.48 105.16 129.48 105.09 128.93 105.09 ;
      RECT  130.37 105.09 130.58 105.47 ;
      RECT  127.25 103.82 127.46 104.37 ;
      RECT  127.46 103.82 128.39 104.37 ;
      RECT  128.39 105.09 128.93 105.47 ;
      RECT  130.37 105.71 130.58 105.95 ;
      RECT  128.93 103.82 130.58 104.37 ;
      RECT  127.25 104.61 127.46 104.85 ;
      RECT  129.86 105.64 130.06 105.71 ;
      POLYGON  130.23 105.09 130.23 105.16 129.86 105.16 129.86 105.4 130.23 105.4 130.23 105.47 130.37 105.47 130.37 105.09 130.23 105.09 ;
      RECT  127.25 105.71 127.46 105.95 ;
      RECT  127.46 105.71 129.86 105.95 ;
      RECT  129.86 104.61 130.37 104.85 ;
      RECT  128.39 103.82 128.93 104.37 ;
      RECT  127.25 107.05 128.39 106.67 ;
      RECT  129.65 107.29 129.86 107.22 ;
      RECT  129.86 106.43 130.37 106.19 ;
      RECT  127.46 107.53 129.86 107.29 ;
      RECT  129.86 107.29 130.06 107.22 ;
      RECT  129.65 106.5 129.86 106.43 ;
      RECT  130.37 107.53 130.58 107.29 ;
      POLYGON  128.93 107.05 128.93 106.67 129.48 106.67 129.48 106.74 129.86 106.74 129.86 106.98 129.48 106.98 129.48 107.05 128.93 107.05 ;
      RECT  130.37 107.05 130.58 106.67 ;
      RECT  127.25 108.32 127.46 107.77 ;
      RECT  127.46 108.32 128.39 107.77 ;
      RECT  128.39 107.05 128.93 106.67 ;
      RECT  130.37 106.43 130.58 106.19 ;
      RECT  128.93 108.32 130.58 107.77 ;
      RECT  127.25 107.53 127.46 107.29 ;
      RECT  129.86 106.5 130.06 106.43 ;
      POLYGON  130.23 107.05 130.23 106.98 129.86 106.98 129.86 106.74 130.23 106.74 130.23 106.67 130.37 106.67 130.37 107.05 130.23 107.05 ;
      RECT  127.25 106.43 127.46 106.19 ;
      RECT  127.46 106.43 129.86 106.19 ;
      RECT  129.86 107.53 130.37 107.29 ;
      RECT  128.39 108.32 128.93 107.77 ;
      RECT  127.25 109.04 128.39 109.42 ;
      RECT  129.65 108.8 129.86 108.87 ;
      RECT  129.86 109.66 130.37 109.9 ;
      RECT  127.46 108.56 129.86 108.8 ;
      RECT  129.86 108.8 130.06 108.87 ;
      RECT  129.65 109.59 129.86 109.66 ;
      RECT  130.37 108.56 130.58 108.8 ;
      POLYGON  128.93 109.04 128.93 109.42 129.48 109.42 129.48 109.35 129.86 109.35 129.86 109.11 129.48 109.11 129.48 109.04 128.93 109.04 ;
      RECT  130.37 109.04 130.58 109.42 ;
      RECT  127.25 107.77 127.46 108.32 ;
      RECT  127.46 107.77 128.39 108.32 ;
      RECT  128.39 109.04 128.93 109.42 ;
      RECT  130.37 109.66 130.58 109.9 ;
      RECT  128.93 107.77 130.58 108.32 ;
      RECT  127.25 108.56 127.46 108.8 ;
      RECT  129.86 109.59 130.06 109.66 ;
      POLYGON  130.23 109.04 130.23 109.11 129.86 109.11 129.86 109.35 130.23 109.35 130.23 109.42 130.37 109.42 130.37 109.04 130.23 109.04 ;
      RECT  127.25 109.66 127.46 109.9 ;
      RECT  127.46 109.66 129.86 109.9 ;
      RECT  129.86 108.56 130.37 108.8 ;
      RECT  128.39 107.77 128.93 108.32 ;
      RECT  127.25 111.0 128.39 110.62 ;
      RECT  129.65 111.24 129.86 111.17 ;
      RECT  129.86 110.38 130.37 110.14 ;
      RECT  127.46 111.48 129.86 111.24 ;
      RECT  129.86 111.24 130.06 111.17 ;
      RECT  129.65 110.45 129.86 110.38 ;
      RECT  130.37 111.48 130.58 111.24 ;
      POLYGON  128.93 111.0 128.93 110.62 129.48 110.62 129.48 110.69 129.86 110.69 129.86 110.93 129.48 110.93 129.48 111.0 128.93 111.0 ;
      RECT  130.37 111.0 130.58 110.62 ;
      RECT  127.25 112.27 127.46 111.72 ;
      RECT  127.46 112.27 128.39 111.72 ;
      RECT  128.39 111.0 128.93 110.62 ;
      RECT  130.37 110.38 130.58 110.14 ;
      RECT  128.93 112.27 130.58 111.72 ;
      RECT  127.25 111.48 127.46 111.24 ;
      RECT  129.86 110.45 130.06 110.38 ;
      POLYGON  130.23 111.0 130.23 110.93 129.86 110.93 129.86 110.69 130.23 110.69 130.23 110.62 130.37 110.62 130.37 111.0 130.23 111.0 ;
      RECT  127.25 110.38 127.46 110.14 ;
      RECT  127.46 110.38 129.86 110.14 ;
      RECT  129.86 111.48 130.37 111.24 ;
      RECT  128.39 112.27 128.93 111.72 ;
      RECT  127.25 112.99 128.39 113.37 ;
      RECT  129.65 112.75 129.86 112.82 ;
      RECT  129.86 113.61 130.37 113.85 ;
      RECT  127.46 112.51 129.86 112.75 ;
      RECT  129.86 112.75 130.06 112.82 ;
      RECT  129.65 113.54 129.86 113.61 ;
      RECT  130.37 112.51 130.58 112.75 ;
      POLYGON  128.93 112.99 128.93 113.37 129.48 113.37 129.48 113.3 129.86 113.3 129.86 113.06 129.48 113.06 129.48 112.99 128.93 112.99 ;
      RECT  130.37 112.99 130.58 113.37 ;
      RECT  127.25 111.72 127.46 112.27 ;
      RECT  127.46 111.72 128.39 112.27 ;
      RECT  128.39 112.99 128.93 113.37 ;
      RECT  130.37 113.61 130.58 113.85 ;
      RECT  128.93 111.72 130.58 112.27 ;
      RECT  127.25 112.51 127.46 112.75 ;
      RECT  129.86 113.54 130.06 113.61 ;
      POLYGON  130.23 112.99 130.23 113.06 129.86 113.06 129.86 113.3 130.23 113.3 130.23 113.37 130.37 113.37 130.37 112.99 130.23 112.99 ;
      RECT  127.25 113.61 127.46 113.85 ;
      RECT  127.46 113.61 129.86 113.85 ;
      RECT  129.86 112.51 130.37 112.75 ;
      RECT  128.39 111.72 128.93 112.27 ;
      RECT  127.25 114.95 128.39 114.57 ;
      RECT  129.65 115.19 129.86 115.12 ;
      RECT  129.86 114.33 130.37 114.09 ;
      RECT  127.46 115.43 129.86 115.19 ;
      RECT  129.86 115.19 130.06 115.12 ;
      RECT  129.65 114.4 129.86 114.33 ;
      RECT  130.37 115.43 130.58 115.19 ;
      POLYGON  128.93 114.95 128.93 114.57 129.48 114.57 129.48 114.64 129.86 114.64 129.86 114.88 129.48 114.88 129.48 114.95 128.93 114.95 ;
      RECT  130.37 114.95 130.58 114.57 ;
      RECT  127.25 116.22 127.46 115.67 ;
      RECT  127.46 116.22 128.39 115.67 ;
      RECT  128.39 114.95 128.93 114.57 ;
      RECT  130.37 114.33 130.58 114.09 ;
      RECT  128.93 116.22 130.58 115.67 ;
      RECT  127.25 115.43 127.46 115.19 ;
      RECT  129.86 114.4 130.06 114.33 ;
      POLYGON  130.23 114.95 130.23 114.88 129.86 114.88 129.86 114.64 130.23 114.64 130.23 114.57 130.37 114.57 130.37 114.95 130.23 114.95 ;
      RECT  127.25 114.33 127.46 114.09 ;
      RECT  127.46 114.33 129.86 114.09 ;
      RECT  129.86 115.43 130.37 115.19 ;
      RECT  128.39 116.22 128.93 115.67 ;
      RECT  127.25 116.94 128.39 117.32 ;
      RECT  129.65 116.7 129.86 116.77 ;
      RECT  129.86 117.56 130.37 117.8 ;
      RECT  127.46 116.46 129.86 116.7 ;
      RECT  129.86 116.7 130.06 116.77 ;
      RECT  129.65 117.49 129.86 117.56 ;
      RECT  130.37 116.46 130.58 116.7 ;
      POLYGON  128.93 116.94 128.93 117.32 129.48 117.32 129.48 117.25 129.86 117.25 129.86 117.01 129.48 117.01 129.48 116.94 128.93 116.94 ;
      RECT  130.37 116.94 130.58 117.32 ;
      RECT  127.25 115.67 127.46 116.22 ;
      RECT  127.46 115.67 128.39 116.22 ;
      RECT  128.39 116.94 128.93 117.32 ;
      RECT  130.37 117.56 130.58 117.8 ;
      RECT  128.93 115.67 130.58 116.22 ;
      RECT  127.25 116.46 127.46 116.7 ;
      RECT  129.86 117.49 130.06 117.56 ;
      POLYGON  130.23 116.94 130.23 117.01 129.86 117.01 129.86 117.25 130.23 117.25 130.23 117.32 130.37 117.32 130.37 116.94 130.23 116.94 ;
      RECT  127.25 117.56 127.46 117.8 ;
      RECT  127.46 117.56 129.86 117.8 ;
      RECT  129.86 116.46 130.37 116.7 ;
      RECT  128.39 115.67 128.93 116.22 ;
      RECT  127.25 118.9 128.39 118.52 ;
      RECT  129.65 119.14 129.86 119.07 ;
      RECT  129.86 118.28 130.37 118.04 ;
      RECT  127.46 119.38 129.86 119.14 ;
      RECT  129.86 119.14 130.06 119.07 ;
      RECT  129.65 118.35 129.86 118.28 ;
      RECT  130.37 119.38 130.58 119.14 ;
      POLYGON  128.93 118.9 128.93 118.52 129.48 118.52 129.48 118.59 129.86 118.59 129.86 118.83 129.48 118.83 129.48 118.9 128.93 118.9 ;
      RECT  130.37 118.9 130.58 118.52 ;
      RECT  127.25 120.17 127.46 119.62 ;
      RECT  127.46 120.17 128.39 119.62 ;
      RECT  128.39 118.9 128.93 118.52 ;
      RECT  130.37 118.28 130.58 118.04 ;
      RECT  128.93 120.17 130.58 119.62 ;
      RECT  127.25 119.38 127.46 119.14 ;
      RECT  129.86 118.35 130.06 118.28 ;
      POLYGON  130.23 118.9 130.23 118.83 129.86 118.83 129.86 118.59 130.23 118.59 130.23 118.52 130.37 118.52 130.37 118.9 130.23 118.9 ;
      RECT  127.25 118.28 127.46 118.04 ;
      RECT  127.46 118.28 129.86 118.04 ;
      RECT  129.86 119.38 130.37 119.14 ;
      RECT  128.39 120.17 128.93 119.62 ;
      RECT  127.25 120.89 128.39 121.27 ;
      RECT  129.65 120.65 129.86 120.72 ;
      RECT  129.86 121.51 130.37 121.75 ;
      RECT  127.46 120.41 129.86 120.65 ;
      RECT  129.86 120.65 130.06 120.72 ;
      RECT  129.65 121.44 129.86 121.51 ;
      RECT  130.37 120.41 130.58 120.65 ;
      POLYGON  128.93 120.89 128.93 121.27 129.48 121.27 129.48 121.2 129.86 121.2 129.86 120.96 129.48 120.96 129.48 120.89 128.93 120.89 ;
      RECT  130.37 120.89 130.58 121.27 ;
      RECT  127.25 119.62 127.46 120.17 ;
      RECT  127.46 119.62 128.39 120.17 ;
      RECT  128.39 120.89 128.93 121.27 ;
      RECT  130.37 121.51 130.58 121.75 ;
      RECT  128.93 119.62 130.58 120.17 ;
      RECT  127.25 120.41 127.46 120.65 ;
      RECT  129.86 121.44 130.06 121.51 ;
      POLYGON  130.23 120.89 130.23 120.96 129.86 120.96 129.86 121.2 130.23 121.2 130.23 121.27 130.37 121.27 130.37 120.89 130.23 120.89 ;
      RECT  127.25 121.51 127.46 121.75 ;
      RECT  127.46 121.51 129.86 121.75 ;
      RECT  129.86 120.41 130.37 120.65 ;
      RECT  128.39 119.62 128.93 120.17 ;
      RECT  127.25 122.85 128.39 122.47 ;
      RECT  129.65 123.09 129.86 123.02 ;
      RECT  129.86 122.23 130.37 121.99 ;
      RECT  127.46 123.33 129.86 123.09 ;
      RECT  129.86 123.09 130.06 123.02 ;
      RECT  129.65 122.3 129.86 122.23 ;
      RECT  130.37 123.33 130.58 123.09 ;
      POLYGON  128.93 122.85 128.93 122.47 129.48 122.47 129.48 122.54 129.86 122.54 129.86 122.78 129.48 122.78 129.48 122.85 128.93 122.85 ;
      RECT  130.37 122.85 130.58 122.47 ;
      RECT  127.25 124.12 127.46 123.57 ;
      RECT  127.46 124.12 128.39 123.57 ;
      RECT  128.39 122.85 128.93 122.47 ;
      RECT  130.37 122.23 130.58 121.99 ;
      RECT  128.93 124.12 130.58 123.57 ;
      RECT  127.25 123.33 127.46 123.09 ;
      RECT  129.86 122.3 130.06 122.23 ;
      POLYGON  130.23 122.85 130.23 122.78 129.86 122.78 129.86 122.54 130.23 122.54 130.23 122.47 130.37 122.47 130.37 122.85 130.23 122.85 ;
      RECT  127.25 122.23 127.46 121.99 ;
      RECT  127.46 122.23 129.86 121.99 ;
      RECT  129.86 123.33 130.37 123.09 ;
      RECT  128.39 124.12 128.93 123.57 ;
      RECT  133.91 93.24 132.77 93.62 ;
      RECT  131.51 93.0 131.3 93.07 ;
      RECT  131.3 93.86 130.79 94.1 ;
      RECT  133.7 92.76 131.3 93.0 ;
      RECT  131.3 93.0 131.1 93.07 ;
      RECT  131.51 93.79 131.3 93.86 ;
      RECT  130.79 92.76 130.58 93.0 ;
      POLYGON  132.23 93.24 132.23 93.62 131.68 93.62 131.68 93.55 131.3 93.55 131.3 93.31 131.68 93.31 131.68 93.24 132.23 93.24 ;
      RECT  130.79 93.24 130.58 93.62 ;
      RECT  133.91 91.97 133.7 92.52 ;
      RECT  133.7 91.97 132.77 92.52 ;
      RECT  132.77 93.24 132.23 93.62 ;
      RECT  130.79 93.86 130.58 94.1 ;
      RECT  132.23 91.97 130.58 92.52 ;
      RECT  133.91 92.76 133.7 93.0 ;
      RECT  131.3 93.79 131.1 93.86 ;
      POLYGON  130.93 93.24 130.93 93.31 131.3 93.31 131.3 93.55 130.93 93.55 130.93 93.62 130.79 93.62 130.79 93.24 130.93 93.24 ;
      RECT  133.91 93.86 133.7 94.1 ;
      RECT  133.7 93.86 131.3 94.1 ;
      RECT  131.3 92.76 130.79 93.0 ;
      RECT  132.77 91.97 132.23 92.52 ;
      RECT  133.91 95.2 132.77 94.82 ;
      RECT  131.51 95.44 131.3 95.37 ;
      RECT  131.3 94.58 130.79 94.34 ;
      RECT  133.7 95.68 131.3 95.44 ;
      RECT  131.3 95.44 131.1 95.37 ;
      RECT  131.51 94.65 131.3 94.58 ;
      RECT  130.79 95.68 130.58 95.44 ;
      POLYGON  132.23 95.2 132.23 94.82 131.68 94.82 131.68 94.89 131.3 94.89 131.3 95.13 131.68 95.13 131.68 95.2 132.23 95.2 ;
      RECT  130.79 95.2 130.58 94.82 ;
      RECT  133.91 96.47 133.7 95.92 ;
      RECT  133.7 96.47 132.77 95.92 ;
      RECT  132.77 95.2 132.23 94.82 ;
      RECT  130.79 94.58 130.58 94.34 ;
      RECT  132.23 96.47 130.58 95.92 ;
      RECT  133.91 95.68 133.7 95.44 ;
      RECT  131.3 94.65 131.1 94.58 ;
      POLYGON  130.93 95.2 130.93 95.13 131.3 95.13 131.3 94.89 130.93 94.89 130.93 94.82 130.79 94.82 130.79 95.2 130.93 95.2 ;
      RECT  133.91 94.58 133.7 94.34 ;
      RECT  133.7 94.58 131.3 94.34 ;
      RECT  131.3 95.68 130.79 95.44 ;
      RECT  132.77 96.47 132.23 95.92 ;
      RECT  133.91 97.19 132.77 97.57 ;
      RECT  131.51 96.95 131.3 97.02 ;
      RECT  131.3 97.81 130.79 98.05 ;
      RECT  133.7 96.71 131.3 96.95 ;
      RECT  131.3 96.95 131.1 97.02 ;
      RECT  131.51 97.74 131.3 97.81 ;
      RECT  130.79 96.71 130.58 96.95 ;
      POLYGON  132.23 97.19 132.23 97.57 131.68 97.57 131.68 97.5 131.3 97.5 131.3 97.26 131.68 97.26 131.68 97.19 132.23 97.19 ;
      RECT  130.79 97.19 130.58 97.57 ;
      RECT  133.91 95.92 133.7 96.47 ;
      RECT  133.7 95.92 132.77 96.47 ;
      RECT  132.77 97.19 132.23 97.57 ;
      RECT  130.79 97.81 130.58 98.05 ;
      RECT  132.23 95.92 130.58 96.47 ;
      RECT  133.91 96.71 133.7 96.95 ;
      RECT  131.3 97.74 131.1 97.81 ;
      POLYGON  130.93 97.19 130.93 97.26 131.3 97.26 131.3 97.5 130.93 97.5 130.93 97.57 130.79 97.57 130.79 97.19 130.93 97.19 ;
      RECT  133.91 97.81 133.7 98.05 ;
      RECT  133.7 97.81 131.3 98.05 ;
      RECT  131.3 96.71 130.79 96.95 ;
      RECT  132.77 95.92 132.23 96.47 ;
      RECT  133.91 99.15 132.77 98.77 ;
      RECT  131.51 99.39 131.3 99.32 ;
      RECT  131.3 98.53 130.79 98.29 ;
      RECT  133.7 99.63 131.3 99.39 ;
      RECT  131.3 99.39 131.1 99.32 ;
      RECT  131.51 98.6 131.3 98.53 ;
      RECT  130.79 99.63 130.58 99.39 ;
      POLYGON  132.23 99.15 132.23 98.77 131.68 98.77 131.68 98.84 131.3 98.84 131.3 99.08 131.68 99.08 131.68 99.15 132.23 99.15 ;
      RECT  130.79 99.15 130.58 98.77 ;
      RECT  133.91 100.42 133.7 99.87 ;
      RECT  133.7 100.42 132.77 99.87 ;
      RECT  132.77 99.15 132.23 98.77 ;
      RECT  130.79 98.53 130.58 98.29 ;
      RECT  132.23 100.42 130.58 99.87 ;
      RECT  133.91 99.63 133.7 99.39 ;
      RECT  131.3 98.6 131.1 98.53 ;
      POLYGON  130.93 99.15 130.93 99.08 131.3 99.08 131.3 98.84 130.93 98.84 130.93 98.77 130.79 98.77 130.79 99.15 130.93 99.15 ;
      RECT  133.91 98.53 133.7 98.29 ;
      RECT  133.7 98.53 131.3 98.29 ;
      RECT  131.3 99.63 130.79 99.39 ;
      RECT  132.77 100.42 132.23 99.87 ;
      RECT  133.91 101.14 132.77 101.52 ;
      RECT  131.51 100.9 131.3 100.97 ;
      RECT  131.3 101.76 130.79 102.0 ;
      RECT  133.7 100.66 131.3 100.9 ;
      RECT  131.3 100.9 131.1 100.97 ;
      RECT  131.51 101.69 131.3 101.76 ;
      RECT  130.79 100.66 130.58 100.9 ;
      POLYGON  132.23 101.14 132.23 101.52 131.68 101.52 131.68 101.45 131.3 101.45 131.3 101.21 131.68 101.21 131.68 101.14 132.23 101.14 ;
      RECT  130.79 101.14 130.58 101.52 ;
      RECT  133.91 99.87 133.7 100.42 ;
      RECT  133.7 99.87 132.77 100.42 ;
      RECT  132.77 101.14 132.23 101.52 ;
      RECT  130.79 101.76 130.58 102.0 ;
      RECT  132.23 99.87 130.58 100.42 ;
      RECT  133.91 100.66 133.7 100.9 ;
      RECT  131.3 101.69 131.1 101.76 ;
      POLYGON  130.93 101.14 130.93 101.21 131.3 101.21 131.3 101.45 130.93 101.45 130.93 101.52 130.79 101.52 130.79 101.14 130.93 101.14 ;
      RECT  133.91 101.76 133.7 102.0 ;
      RECT  133.7 101.76 131.3 102.0 ;
      RECT  131.3 100.66 130.79 100.9 ;
      RECT  132.77 99.87 132.23 100.42 ;
      RECT  133.91 103.1 132.77 102.72 ;
      RECT  131.51 103.34 131.3 103.27 ;
      RECT  131.3 102.48 130.79 102.24 ;
      RECT  133.7 103.58 131.3 103.34 ;
      RECT  131.3 103.34 131.1 103.27 ;
      RECT  131.51 102.55 131.3 102.48 ;
      RECT  130.79 103.58 130.58 103.34 ;
      POLYGON  132.23 103.1 132.23 102.72 131.68 102.72 131.68 102.79 131.3 102.79 131.3 103.03 131.68 103.03 131.68 103.1 132.23 103.1 ;
      RECT  130.79 103.1 130.58 102.72 ;
      RECT  133.91 104.37 133.7 103.82 ;
      RECT  133.7 104.37 132.77 103.82 ;
      RECT  132.77 103.1 132.23 102.72 ;
      RECT  130.79 102.48 130.58 102.24 ;
      RECT  132.23 104.37 130.58 103.82 ;
      RECT  133.91 103.58 133.7 103.34 ;
      RECT  131.3 102.55 131.1 102.48 ;
      POLYGON  130.93 103.1 130.93 103.03 131.3 103.03 131.3 102.79 130.93 102.79 130.93 102.72 130.79 102.72 130.79 103.1 130.93 103.1 ;
      RECT  133.91 102.48 133.7 102.24 ;
      RECT  133.7 102.48 131.3 102.24 ;
      RECT  131.3 103.58 130.79 103.34 ;
      RECT  132.77 104.37 132.23 103.82 ;
      RECT  133.91 105.09 132.77 105.47 ;
      RECT  131.51 104.85 131.3 104.92 ;
      RECT  131.3 105.71 130.79 105.95 ;
      RECT  133.7 104.61 131.3 104.85 ;
      RECT  131.3 104.85 131.1 104.92 ;
      RECT  131.51 105.64 131.3 105.71 ;
      RECT  130.79 104.61 130.58 104.85 ;
      POLYGON  132.23 105.09 132.23 105.47 131.68 105.47 131.68 105.4 131.3 105.4 131.3 105.16 131.68 105.16 131.68 105.09 132.23 105.09 ;
      RECT  130.79 105.09 130.58 105.47 ;
      RECT  133.91 103.82 133.7 104.37 ;
      RECT  133.7 103.82 132.77 104.37 ;
      RECT  132.77 105.09 132.23 105.47 ;
      RECT  130.79 105.71 130.58 105.95 ;
      RECT  132.23 103.82 130.58 104.37 ;
      RECT  133.91 104.61 133.7 104.85 ;
      RECT  131.3 105.64 131.1 105.71 ;
      POLYGON  130.93 105.09 130.93 105.16 131.3 105.16 131.3 105.4 130.93 105.4 130.93 105.47 130.79 105.47 130.79 105.09 130.93 105.09 ;
      RECT  133.91 105.71 133.7 105.95 ;
      RECT  133.7 105.71 131.3 105.95 ;
      RECT  131.3 104.61 130.79 104.85 ;
      RECT  132.77 103.82 132.23 104.37 ;
      RECT  133.91 107.05 132.77 106.67 ;
      RECT  131.51 107.29 131.3 107.22 ;
      RECT  131.3 106.43 130.79 106.19 ;
      RECT  133.7 107.53 131.3 107.29 ;
      RECT  131.3 107.29 131.1 107.22 ;
      RECT  131.51 106.5 131.3 106.43 ;
      RECT  130.79 107.53 130.58 107.29 ;
      POLYGON  132.23 107.05 132.23 106.67 131.68 106.67 131.68 106.74 131.3 106.74 131.3 106.98 131.68 106.98 131.68 107.05 132.23 107.05 ;
      RECT  130.79 107.05 130.58 106.67 ;
      RECT  133.91 108.32 133.7 107.77 ;
      RECT  133.7 108.32 132.77 107.77 ;
      RECT  132.77 107.05 132.23 106.67 ;
      RECT  130.79 106.43 130.58 106.19 ;
      RECT  132.23 108.32 130.58 107.77 ;
      RECT  133.91 107.53 133.7 107.29 ;
      RECT  131.3 106.5 131.1 106.43 ;
      POLYGON  130.93 107.05 130.93 106.98 131.3 106.98 131.3 106.74 130.93 106.74 130.93 106.67 130.79 106.67 130.79 107.05 130.93 107.05 ;
      RECT  133.91 106.43 133.7 106.19 ;
      RECT  133.7 106.43 131.3 106.19 ;
      RECT  131.3 107.53 130.79 107.29 ;
      RECT  132.77 108.32 132.23 107.77 ;
      RECT  133.91 109.04 132.77 109.42 ;
      RECT  131.51 108.8 131.3 108.87 ;
      RECT  131.3 109.66 130.79 109.9 ;
      RECT  133.7 108.56 131.3 108.8 ;
      RECT  131.3 108.8 131.1 108.87 ;
      RECT  131.51 109.59 131.3 109.66 ;
      RECT  130.79 108.56 130.58 108.8 ;
      POLYGON  132.23 109.04 132.23 109.42 131.68 109.42 131.68 109.35 131.3 109.35 131.3 109.11 131.68 109.11 131.68 109.04 132.23 109.04 ;
      RECT  130.79 109.04 130.58 109.42 ;
      RECT  133.91 107.77 133.7 108.32 ;
      RECT  133.7 107.77 132.77 108.32 ;
      RECT  132.77 109.04 132.23 109.42 ;
      RECT  130.79 109.66 130.58 109.9 ;
      RECT  132.23 107.77 130.58 108.32 ;
      RECT  133.91 108.56 133.7 108.8 ;
      RECT  131.3 109.59 131.1 109.66 ;
      POLYGON  130.93 109.04 130.93 109.11 131.3 109.11 131.3 109.35 130.93 109.35 130.93 109.42 130.79 109.42 130.79 109.04 130.93 109.04 ;
      RECT  133.91 109.66 133.7 109.9 ;
      RECT  133.7 109.66 131.3 109.9 ;
      RECT  131.3 108.56 130.79 108.8 ;
      RECT  132.77 107.77 132.23 108.32 ;
      RECT  133.91 111.0 132.77 110.62 ;
      RECT  131.51 111.24 131.3 111.17 ;
      RECT  131.3 110.38 130.79 110.14 ;
      RECT  133.7 111.48 131.3 111.24 ;
      RECT  131.3 111.24 131.1 111.17 ;
      RECT  131.51 110.45 131.3 110.38 ;
      RECT  130.79 111.48 130.58 111.24 ;
      POLYGON  132.23 111.0 132.23 110.62 131.68 110.62 131.68 110.69 131.3 110.69 131.3 110.93 131.68 110.93 131.68 111.0 132.23 111.0 ;
      RECT  130.79 111.0 130.58 110.62 ;
      RECT  133.91 112.27 133.7 111.72 ;
      RECT  133.7 112.27 132.77 111.72 ;
      RECT  132.77 111.0 132.23 110.62 ;
      RECT  130.79 110.38 130.58 110.14 ;
      RECT  132.23 112.27 130.58 111.72 ;
      RECT  133.91 111.48 133.7 111.24 ;
      RECT  131.3 110.45 131.1 110.38 ;
      POLYGON  130.93 111.0 130.93 110.93 131.3 110.93 131.3 110.69 130.93 110.69 130.93 110.62 130.79 110.62 130.79 111.0 130.93 111.0 ;
      RECT  133.91 110.38 133.7 110.14 ;
      RECT  133.7 110.38 131.3 110.14 ;
      RECT  131.3 111.48 130.79 111.24 ;
      RECT  132.77 112.27 132.23 111.72 ;
      RECT  133.91 112.99 132.77 113.37 ;
      RECT  131.51 112.75 131.3 112.82 ;
      RECT  131.3 113.61 130.79 113.85 ;
      RECT  133.7 112.51 131.3 112.75 ;
      RECT  131.3 112.75 131.1 112.82 ;
      RECT  131.51 113.54 131.3 113.61 ;
      RECT  130.79 112.51 130.58 112.75 ;
      POLYGON  132.23 112.99 132.23 113.37 131.68 113.37 131.68 113.3 131.3 113.3 131.3 113.06 131.68 113.06 131.68 112.99 132.23 112.99 ;
      RECT  130.79 112.99 130.58 113.37 ;
      RECT  133.91 111.72 133.7 112.27 ;
      RECT  133.7 111.72 132.77 112.27 ;
      RECT  132.77 112.99 132.23 113.37 ;
      RECT  130.79 113.61 130.58 113.85 ;
      RECT  132.23 111.72 130.58 112.27 ;
      RECT  133.91 112.51 133.7 112.75 ;
      RECT  131.3 113.54 131.1 113.61 ;
      POLYGON  130.93 112.99 130.93 113.06 131.3 113.06 131.3 113.3 130.93 113.3 130.93 113.37 130.79 113.37 130.79 112.99 130.93 112.99 ;
      RECT  133.91 113.61 133.7 113.85 ;
      RECT  133.7 113.61 131.3 113.85 ;
      RECT  131.3 112.51 130.79 112.75 ;
      RECT  132.77 111.72 132.23 112.27 ;
      RECT  133.91 114.95 132.77 114.57 ;
      RECT  131.51 115.19 131.3 115.12 ;
      RECT  131.3 114.33 130.79 114.09 ;
      RECT  133.7 115.43 131.3 115.19 ;
      RECT  131.3 115.19 131.1 115.12 ;
      RECT  131.51 114.4 131.3 114.33 ;
      RECT  130.79 115.43 130.58 115.19 ;
      POLYGON  132.23 114.95 132.23 114.57 131.68 114.57 131.68 114.64 131.3 114.64 131.3 114.88 131.68 114.88 131.68 114.95 132.23 114.95 ;
      RECT  130.79 114.95 130.58 114.57 ;
      RECT  133.91 116.22 133.7 115.67 ;
      RECT  133.7 116.22 132.77 115.67 ;
      RECT  132.77 114.95 132.23 114.57 ;
      RECT  130.79 114.33 130.58 114.09 ;
      RECT  132.23 116.22 130.58 115.67 ;
      RECT  133.91 115.43 133.7 115.19 ;
      RECT  131.3 114.4 131.1 114.33 ;
      POLYGON  130.93 114.95 130.93 114.88 131.3 114.88 131.3 114.64 130.93 114.64 130.93 114.57 130.79 114.57 130.79 114.95 130.93 114.95 ;
      RECT  133.91 114.33 133.7 114.09 ;
      RECT  133.7 114.33 131.3 114.09 ;
      RECT  131.3 115.43 130.79 115.19 ;
      RECT  132.77 116.22 132.23 115.67 ;
      RECT  133.91 116.94 132.77 117.32 ;
      RECT  131.51 116.7 131.3 116.77 ;
      RECT  131.3 117.56 130.79 117.8 ;
      RECT  133.7 116.46 131.3 116.7 ;
      RECT  131.3 116.7 131.1 116.77 ;
      RECT  131.51 117.49 131.3 117.56 ;
      RECT  130.79 116.46 130.58 116.7 ;
      POLYGON  132.23 116.94 132.23 117.32 131.68 117.32 131.68 117.25 131.3 117.25 131.3 117.01 131.68 117.01 131.68 116.94 132.23 116.94 ;
      RECT  130.79 116.94 130.58 117.32 ;
      RECT  133.91 115.67 133.7 116.22 ;
      RECT  133.7 115.67 132.77 116.22 ;
      RECT  132.77 116.94 132.23 117.32 ;
      RECT  130.79 117.56 130.58 117.8 ;
      RECT  132.23 115.67 130.58 116.22 ;
      RECT  133.91 116.46 133.7 116.7 ;
      RECT  131.3 117.49 131.1 117.56 ;
      POLYGON  130.93 116.94 130.93 117.01 131.3 117.01 131.3 117.25 130.93 117.25 130.93 117.32 130.79 117.32 130.79 116.94 130.93 116.94 ;
      RECT  133.91 117.56 133.7 117.8 ;
      RECT  133.7 117.56 131.3 117.8 ;
      RECT  131.3 116.46 130.79 116.7 ;
      RECT  132.77 115.67 132.23 116.22 ;
      RECT  133.91 118.9 132.77 118.52 ;
      RECT  131.51 119.14 131.3 119.07 ;
      RECT  131.3 118.28 130.79 118.04 ;
      RECT  133.7 119.38 131.3 119.14 ;
      RECT  131.3 119.14 131.1 119.07 ;
      RECT  131.51 118.35 131.3 118.28 ;
      RECT  130.79 119.38 130.58 119.14 ;
      POLYGON  132.23 118.9 132.23 118.52 131.68 118.52 131.68 118.59 131.3 118.59 131.3 118.83 131.68 118.83 131.68 118.9 132.23 118.9 ;
      RECT  130.79 118.9 130.58 118.52 ;
      RECT  133.91 120.17 133.7 119.62 ;
      RECT  133.7 120.17 132.77 119.62 ;
      RECT  132.77 118.9 132.23 118.52 ;
      RECT  130.79 118.28 130.58 118.04 ;
      RECT  132.23 120.17 130.58 119.62 ;
      RECT  133.91 119.38 133.7 119.14 ;
      RECT  131.3 118.35 131.1 118.28 ;
      POLYGON  130.93 118.9 130.93 118.83 131.3 118.83 131.3 118.59 130.93 118.59 130.93 118.52 130.79 118.52 130.79 118.9 130.93 118.9 ;
      RECT  133.91 118.28 133.7 118.04 ;
      RECT  133.7 118.28 131.3 118.04 ;
      RECT  131.3 119.38 130.79 119.14 ;
      RECT  132.77 120.17 132.23 119.62 ;
      RECT  133.91 120.89 132.77 121.27 ;
      RECT  131.51 120.65 131.3 120.72 ;
      RECT  131.3 121.51 130.79 121.75 ;
      RECT  133.7 120.41 131.3 120.65 ;
      RECT  131.3 120.65 131.1 120.72 ;
      RECT  131.51 121.44 131.3 121.51 ;
      RECT  130.79 120.41 130.58 120.65 ;
      POLYGON  132.23 120.89 132.23 121.27 131.68 121.27 131.68 121.2 131.3 121.2 131.3 120.96 131.68 120.96 131.68 120.89 132.23 120.89 ;
      RECT  130.79 120.89 130.58 121.27 ;
      RECT  133.91 119.62 133.7 120.17 ;
      RECT  133.7 119.62 132.77 120.17 ;
      RECT  132.77 120.89 132.23 121.27 ;
      RECT  130.79 121.51 130.58 121.75 ;
      RECT  132.23 119.62 130.58 120.17 ;
      RECT  133.91 120.41 133.7 120.65 ;
      RECT  131.3 121.44 131.1 121.51 ;
      POLYGON  130.93 120.89 130.93 120.96 131.3 120.96 131.3 121.2 130.93 121.2 130.93 121.27 130.79 121.27 130.79 120.89 130.93 120.89 ;
      RECT  133.91 121.51 133.7 121.75 ;
      RECT  133.7 121.51 131.3 121.75 ;
      RECT  131.3 120.41 130.79 120.65 ;
      RECT  132.77 119.62 132.23 120.17 ;
      RECT  133.91 122.85 132.77 122.47 ;
      RECT  131.51 123.09 131.3 123.02 ;
      RECT  131.3 122.23 130.79 121.99 ;
      RECT  133.7 123.33 131.3 123.09 ;
      RECT  131.3 123.09 131.1 123.02 ;
      RECT  131.51 122.3 131.3 122.23 ;
      RECT  130.79 123.33 130.58 123.09 ;
      POLYGON  132.23 122.85 132.23 122.47 131.68 122.47 131.68 122.54 131.3 122.54 131.3 122.78 131.68 122.78 131.68 122.85 132.23 122.85 ;
      RECT  130.79 122.85 130.58 122.47 ;
      RECT  133.91 124.12 133.7 123.57 ;
      RECT  133.7 124.12 132.77 123.57 ;
      RECT  132.77 122.85 132.23 122.47 ;
      RECT  130.79 122.23 130.58 121.99 ;
      RECT  132.23 124.12 130.58 123.57 ;
      RECT  133.91 123.33 133.7 123.09 ;
      RECT  131.3 122.3 131.1 122.23 ;
      POLYGON  130.93 122.85 130.93 122.78 131.3 122.78 131.3 122.54 130.93 122.54 130.93 122.47 130.79 122.47 130.79 122.85 130.93 122.85 ;
      RECT  133.91 122.23 133.7 121.99 ;
      RECT  133.7 122.23 131.3 121.99 ;
      RECT  131.3 123.33 130.79 123.09 ;
      RECT  132.77 124.12 132.23 123.57 ;
      RECT  133.49 93.24 134.63 93.62 ;
      RECT  135.89 93.0 136.1 93.07 ;
      RECT  136.1 93.86 136.61 94.1 ;
      RECT  133.7 92.76 136.1 93.0 ;
      RECT  136.1 93.0 136.3 93.07 ;
      RECT  135.89 93.79 136.1 93.86 ;
      RECT  136.61 92.76 136.82 93.0 ;
      POLYGON  135.17 93.24 135.17 93.62 135.72 93.62 135.72 93.55 136.1 93.55 136.1 93.31 135.72 93.31 135.72 93.24 135.17 93.24 ;
      RECT  136.61 93.24 136.82 93.62 ;
      RECT  133.49 91.97 133.7 92.52 ;
      RECT  133.7 91.97 134.63 92.52 ;
      RECT  134.63 93.24 135.17 93.62 ;
      RECT  136.61 93.86 136.82 94.1 ;
      RECT  135.17 91.97 136.82 92.52 ;
      RECT  133.49 92.76 133.7 93.0 ;
      RECT  136.1 93.79 136.3 93.86 ;
      POLYGON  136.47 93.24 136.47 93.31 136.1 93.31 136.1 93.55 136.47 93.55 136.47 93.62 136.61 93.62 136.61 93.24 136.47 93.24 ;
      RECT  133.49 93.86 133.7 94.1 ;
      RECT  133.7 93.86 136.1 94.1 ;
      RECT  136.1 92.76 136.61 93.0 ;
      RECT  134.63 91.97 135.17 92.52 ;
      RECT  133.49 95.2 134.63 94.82 ;
      RECT  135.89 95.44 136.1 95.37 ;
      RECT  136.1 94.58 136.61 94.34 ;
      RECT  133.7 95.68 136.1 95.44 ;
      RECT  136.1 95.44 136.3 95.37 ;
      RECT  135.89 94.65 136.1 94.58 ;
      RECT  136.61 95.68 136.82 95.44 ;
      POLYGON  135.17 95.2 135.17 94.82 135.72 94.82 135.72 94.89 136.1 94.89 136.1 95.13 135.72 95.13 135.72 95.2 135.17 95.2 ;
      RECT  136.61 95.2 136.82 94.82 ;
      RECT  133.49 96.47 133.7 95.92 ;
      RECT  133.7 96.47 134.63 95.92 ;
      RECT  134.63 95.2 135.17 94.82 ;
      RECT  136.61 94.58 136.82 94.34 ;
      RECT  135.17 96.47 136.82 95.92 ;
      RECT  133.49 95.68 133.7 95.44 ;
      RECT  136.1 94.65 136.3 94.58 ;
      POLYGON  136.47 95.2 136.47 95.13 136.1 95.13 136.1 94.89 136.47 94.89 136.47 94.82 136.61 94.82 136.61 95.2 136.47 95.2 ;
      RECT  133.49 94.58 133.7 94.34 ;
      RECT  133.7 94.58 136.1 94.34 ;
      RECT  136.1 95.68 136.61 95.44 ;
      RECT  134.63 96.47 135.17 95.92 ;
      RECT  133.49 97.19 134.63 97.57 ;
      RECT  135.89 96.95 136.1 97.02 ;
      RECT  136.1 97.81 136.61 98.05 ;
      RECT  133.7 96.71 136.1 96.95 ;
      RECT  136.1 96.95 136.3 97.02 ;
      RECT  135.89 97.74 136.1 97.81 ;
      RECT  136.61 96.71 136.82 96.95 ;
      POLYGON  135.17 97.19 135.17 97.57 135.72 97.57 135.72 97.5 136.1 97.5 136.1 97.26 135.72 97.26 135.72 97.19 135.17 97.19 ;
      RECT  136.61 97.19 136.82 97.57 ;
      RECT  133.49 95.92 133.7 96.47 ;
      RECT  133.7 95.92 134.63 96.47 ;
      RECT  134.63 97.19 135.17 97.57 ;
      RECT  136.61 97.81 136.82 98.05 ;
      RECT  135.17 95.92 136.82 96.47 ;
      RECT  133.49 96.71 133.7 96.95 ;
      RECT  136.1 97.74 136.3 97.81 ;
      POLYGON  136.47 97.19 136.47 97.26 136.1 97.26 136.1 97.5 136.47 97.5 136.47 97.57 136.61 97.57 136.61 97.19 136.47 97.19 ;
      RECT  133.49 97.81 133.7 98.05 ;
      RECT  133.7 97.81 136.1 98.05 ;
      RECT  136.1 96.71 136.61 96.95 ;
      RECT  134.63 95.92 135.17 96.47 ;
      RECT  133.49 99.15 134.63 98.77 ;
      RECT  135.89 99.39 136.1 99.32 ;
      RECT  136.1 98.53 136.61 98.29 ;
      RECT  133.7 99.63 136.1 99.39 ;
      RECT  136.1 99.39 136.3 99.32 ;
      RECT  135.89 98.6 136.1 98.53 ;
      RECT  136.61 99.63 136.82 99.39 ;
      POLYGON  135.17 99.15 135.17 98.77 135.72 98.77 135.72 98.84 136.1 98.84 136.1 99.08 135.72 99.08 135.72 99.15 135.17 99.15 ;
      RECT  136.61 99.15 136.82 98.77 ;
      RECT  133.49 100.42 133.7 99.87 ;
      RECT  133.7 100.42 134.63 99.87 ;
      RECT  134.63 99.15 135.17 98.77 ;
      RECT  136.61 98.53 136.82 98.29 ;
      RECT  135.17 100.42 136.82 99.87 ;
      RECT  133.49 99.63 133.7 99.39 ;
      RECT  136.1 98.6 136.3 98.53 ;
      POLYGON  136.47 99.15 136.47 99.08 136.1 99.08 136.1 98.84 136.47 98.84 136.47 98.77 136.61 98.77 136.61 99.15 136.47 99.15 ;
      RECT  133.49 98.53 133.7 98.29 ;
      RECT  133.7 98.53 136.1 98.29 ;
      RECT  136.1 99.63 136.61 99.39 ;
      RECT  134.63 100.42 135.17 99.87 ;
      RECT  133.49 101.14 134.63 101.52 ;
      RECT  135.89 100.9 136.1 100.97 ;
      RECT  136.1 101.76 136.61 102.0 ;
      RECT  133.7 100.66 136.1 100.9 ;
      RECT  136.1 100.9 136.3 100.97 ;
      RECT  135.89 101.69 136.1 101.76 ;
      RECT  136.61 100.66 136.82 100.9 ;
      POLYGON  135.17 101.14 135.17 101.52 135.72 101.52 135.72 101.45 136.1 101.45 136.1 101.21 135.72 101.21 135.72 101.14 135.17 101.14 ;
      RECT  136.61 101.14 136.82 101.52 ;
      RECT  133.49 99.87 133.7 100.42 ;
      RECT  133.7 99.87 134.63 100.42 ;
      RECT  134.63 101.14 135.17 101.52 ;
      RECT  136.61 101.76 136.82 102.0 ;
      RECT  135.17 99.87 136.82 100.42 ;
      RECT  133.49 100.66 133.7 100.9 ;
      RECT  136.1 101.69 136.3 101.76 ;
      POLYGON  136.47 101.14 136.47 101.21 136.1 101.21 136.1 101.45 136.47 101.45 136.47 101.52 136.61 101.52 136.61 101.14 136.47 101.14 ;
      RECT  133.49 101.76 133.7 102.0 ;
      RECT  133.7 101.76 136.1 102.0 ;
      RECT  136.1 100.66 136.61 100.9 ;
      RECT  134.63 99.87 135.17 100.42 ;
      RECT  133.49 103.1 134.63 102.72 ;
      RECT  135.89 103.34 136.1 103.27 ;
      RECT  136.1 102.48 136.61 102.24 ;
      RECT  133.7 103.58 136.1 103.34 ;
      RECT  136.1 103.34 136.3 103.27 ;
      RECT  135.89 102.55 136.1 102.48 ;
      RECT  136.61 103.58 136.82 103.34 ;
      POLYGON  135.17 103.1 135.17 102.72 135.72 102.72 135.72 102.79 136.1 102.79 136.1 103.03 135.72 103.03 135.72 103.1 135.17 103.1 ;
      RECT  136.61 103.1 136.82 102.72 ;
      RECT  133.49 104.37 133.7 103.82 ;
      RECT  133.7 104.37 134.63 103.82 ;
      RECT  134.63 103.1 135.17 102.72 ;
      RECT  136.61 102.48 136.82 102.24 ;
      RECT  135.17 104.37 136.82 103.82 ;
      RECT  133.49 103.58 133.7 103.34 ;
      RECT  136.1 102.55 136.3 102.48 ;
      POLYGON  136.47 103.1 136.47 103.03 136.1 103.03 136.1 102.79 136.47 102.79 136.47 102.72 136.61 102.72 136.61 103.1 136.47 103.1 ;
      RECT  133.49 102.48 133.7 102.24 ;
      RECT  133.7 102.48 136.1 102.24 ;
      RECT  136.1 103.58 136.61 103.34 ;
      RECT  134.63 104.37 135.17 103.82 ;
      RECT  133.49 105.09 134.63 105.47 ;
      RECT  135.89 104.85 136.1 104.92 ;
      RECT  136.1 105.71 136.61 105.95 ;
      RECT  133.7 104.61 136.1 104.85 ;
      RECT  136.1 104.85 136.3 104.92 ;
      RECT  135.89 105.64 136.1 105.71 ;
      RECT  136.61 104.61 136.82 104.85 ;
      POLYGON  135.17 105.09 135.17 105.47 135.72 105.47 135.72 105.4 136.1 105.4 136.1 105.16 135.72 105.16 135.72 105.09 135.17 105.09 ;
      RECT  136.61 105.09 136.82 105.47 ;
      RECT  133.49 103.82 133.7 104.37 ;
      RECT  133.7 103.82 134.63 104.37 ;
      RECT  134.63 105.09 135.17 105.47 ;
      RECT  136.61 105.71 136.82 105.95 ;
      RECT  135.17 103.82 136.82 104.37 ;
      RECT  133.49 104.61 133.7 104.85 ;
      RECT  136.1 105.64 136.3 105.71 ;
      POLYGON  136.47 105.09 136.47 105.16 136.1 105.16 136.1 105.4 136.47 105.4 136.47 105.47 136.61 105.47 136.61 105.09 136.47 105.09 ;
      RECT  133.49 105.71 133.7 105.95 ;
      RECT  133.7 105.71 136.1 105.95 ;
      RECT  136.1 104.61 136.61 104.85 ;
      RECT  134.63 103.82 135.17 104.37 ;
      RECT  133.49 107.05 134.63 106.67 ;
      RECT  135.89 107.29 136.1 107.22 ;
      RECT  136.1 106.43 136.61 106.19 ;
      RECT  133.7 107.53 136.1 107.29 ;
      RECT  136.1 107.29 136.3 107.22 ;
      RECT  135.89 106.5 136.1 106.43 ;
      RECT  136.61 107.53 136.82 107.29 ;
      POLYGON  135.17 107.05 135.17 106.67 135.72 106.67 135.72 106.74 136.1 106.74 136.1 106.98 135.72 106.98 135.72 107.05 135.17 107.05 ;
      RECT  136.61 107.05 136.82 106.67 ;
      RECT  133.49 108.32 133.7 107.77 ;
      RECT  133.7 108.32 134.63 107.77 ;
      RECT  134.63 107.05 135.17 106.67 ;
      RECT  136.61 106.43 136.82 106.19 ;
      RECT  135.17 108.32 136.82 107.77 ;
      RECT  133.49 107.53 133.7 107.29 ;
      RECT  136.1 106.5 136.3 106.43 ;
      POLYGON  136.47 107.05 136.47 106.98 136.1 106.98 136.1 106.74 136.47 106.74 136.47 106.67 136.61 106.67 136.61 107.05 136.47 107.05 ;
      RECT  133.49 106.43 133.7 106.19 ;
      RECT  133.7 106.43 136.1 106.19 ;
      RECT  136.1 107.53 136.61 107.29 ;
      RECT  134.63 108.32 135.17 107.77 ;
      RECT  133.49 109.04 134.63 109.42 ;
      RECT  135.89 108.8 136.1 108.87 ;
      RECT  136.1 109.66 136.61 109.9 ;
      RECT  133.7 108.56 136.1 108.8 ;
      RECT  136.1 108.8 136.3 108.87 ;
      RECT  135.89 109.59 136.1 109.66 ;
      RECT  136.61 108.56 136.82 108.8 ;
      POLYGON  135.17 109.04 135.17 109.42 135.72 109.42 135.72 109.35 136.1 109.35 136.1 109.11 135.72 109.11 135.72 109.04 135.17 109.04 ;
      RECT  136.61 109.04 136.82 109.42 ;
      RECT  133.49 107.77 133.7 108.32 ;
      RECT  133.7 107.77 134.63 108.32 ;
      RECT  134.63 109.04 135.17 109.42 ;
      RECT  136.61 109.66 136.82 109.9 ;
      RECT  135.17 107.77 136.82 108.32 ;
      RECT  133.49 108.56 133.7 108.8 ;
      RECT  136.1 109.59 136.3 109.66 ;
      POLYGON  136.47 109.04 136.47 109.11 136.1 109.11 136.1 109.35 136.47 109.35 136.47 109.42 136.61 109.42 136.61 109.04 136.47 109.04 ;
      RECT  133.49 109.66 133.7 109.9 ;
      RECT  133.7 109.66 136.1 109.9 ;
      RECT  136.1 108.56 136.61 108.8 ;
      RECT  134.63 107.77 135.17 108.32 ;
      RECT  133.49 111.0 134.63 110.62 ;
      RECT  135.89 111.24 136.1 111.17 ;
      RECT  136.1 110.38 136.61 110.14 ;
      RECT  133.7 111.48 136.1 111.24 ;
      RECT  136.1 111.24 136.3 111.17 ;
      RECT  135.89 110.45 136.1 110.38 ;
      RECT  136.61 111.48 136.82 111.24 ;
      POLYGON  135.17 111.0 135.17 110.62 135.72 110.62 135.72 110.69 136.1 110.69 136.1 110.93 135.72 110.93 135.72 111.0 135.17 111.0 ;
      RECT  136.61 111.0 136.82 110.62 ;
      RECT  133.49 112.27 133.7 111.72 ;
      RECT  133.7 112.27 134.63 111.72 ;
      RECT  134.63 111.0 135.17 110.62 ;
      RECT  136.61 110.38 136.82 110.14 ;
      RECT  135.17 112.27 136.82 111.72 ;
      RECT  133.49 111.48 133.7 111.24 ;
      RECT  136.1 110.45 136.3 110.38 ;
      POLYGON  136.47 111.0 136.47 110.93 136.1 110.93 136.1 110.69 136.47 110.69 136.47 110.62 136.61 110.62 136.61 111.0 136.47 111.0 ;
      RECT  133.49 110.38 133.7 110.14 ;
      RECT  133.7 110.38 136.1 110.14 ;
      RECT  136.1 111.48 136.61 111.24 ;
      RECT  134.63 112.27 135.17 111.72 ;
      RECT  133.49 112.99 134.63 113.37 ;
      RECT  135.89 112.75 136.1 112.82 ;
      RECT  136.1 113.61 136.61 113.85 ;
      RECT  133.7 112.51 136.1 112.75 ;
      RECT  136.1 112.75 136.3 112.82 ;
      RECT  135.89 113.54 136.1 113.61 ;
      RECT  136.61 112.51 136.82 112.75 ;
      POLYGON  135.17 112.99 135.17 113.37 135.72 113.37 135.72 113.3 136.1 113.3 136.1 113.06 135.72 113.06 135.72 112.99 135.17 112.99 ;
      RECT  136.61 112.99 136.82 113.37 ;
      RECT  133.49 111.72 133.7 112.27 ;
      RECT  133.7 111.72 134.63 112.27 ;
      RECT  134.63 112.99 135.17 113.37 ;
      RECT  136.61 113.61 136.82 113.85 ;
      RECT  135.17 111.72 136.82 112.27 ;
      RECT  133.49 112.51 133.7 112.75 ;
      RECT  136.1 113.54 136.3 113.61 ;
      POLYGON  136.47 112.99 136.47 113.06 136.1 113.06 136.1 113.3 136.47 113.3 136.47 113.37 136.61 113.37 136.61 112.99 136.47 112.99 ;
      RECT  133.49 113.61 133.7 113.85 ;
      RECT  133.7 113.61 136.1 113.85 ;
      RECT  136.1 112.51 136.61 112.75 ;
      RECT  134.63 111.72 135.17 112.27 ;
      RECT  133.49 114.95 134.63 114.57 ;
      RECT  135.89 115.19 136.1 115.12 ;
      RECT  136.1 114.33 136.61 114.09 ;
      RECT  133.7 115.43 136.1 115.19 ;
      RECT  136.1 115.19 136.3 115.12 ;
      RECT  135.89 114.4 136.1 114.33 ;
      RECT  136.61 115.43 136.82 115.19 ;
      POLYGON  135.17 114.95 135.17 114.57 135.72 114.57 135.72 114.64 136.1 114.64 136.1 114.88 135.72 114.88 135.72 114.95 135.17 114.95 ;
      RECT  136.61 114.95 136.82 114.57 ;
      RECT  133.49 116.22 133.7 115.67 ;
      RECT  133.7 116.22 134.63 115.67 ;
      RECT  134.63 114.95 135.17 114.57 ;
      RECT  136.61 114.33 136.82 114.09 ;
      RECT  135.17 116.22 136.82 115.67 ;
      RECT  133.49 115.43 133.7 115.19 ;
      RECT  136.1 114.4 136.3 114.33 ;
      POLYGON  136.47 114.95 136.47 114.88 136.1 114.88 136.1 114.64 136.47 114.64 136.47 114.57 136.61 114.57 136.61 114.95 136.47 114.95 ;
      RECT  133.49 114.33 133.7 114.09 ;
      RECT  133.7 114.33 136.1 114.09 ;
      RECT  136.1 115.43 136.61 115.19 ;
      RECT  134.63 116.22 135.17 115.67 ;
      RECT  133.49 116.94 134.63 117.32 ;
      RECT  135.89 116.7 136.1 116.77 ;
      RECT  136.1 117.56 136.61 117.8 ;
      RECT  133.7 116.46 136.1 116.7 ;
      RECT  136.1 116.7 136.3 116.77 ;
      RECT  135.89 117.49 136.1 117.56 ;
      RECT  136.61 116.46 136.82 116.7 ;
      POLYGON  135.17 116.94 135.17 117.32 135.72 117.32 135.72 117.25 136.1 117.25 136.1 117.01 135.72 117.01 135.72 116.94 135.17 116.94 ;
      RECT  136.61 116.94 136.82 117.32 ;
      RECT  133.49 115.67 133.7 116.22 ;
      RECT  133.7 115.67 134.63 116.22 ;
      RECT  134.63 116.94 135.17 117.32 ;
      RECT  136.61 117.56 136.82 117.8 ;
      RECT  135.17 115.67 136.82 116.22 ;
      RECT  133.49 116.46 133.7 116.7 ;
      RECT  136.1 117.49 136.3 117.56 ;
      POLYGON  136.47 116.94 136.47 117.01 136.1 117.01 136.1 117.25 136.47 117.25 136.47 117.32 136.61 117.32 136.61 116.94 136.47 116.94 ;
      RECT  133.49 117.56 133.7 117.8 ;
      RECT  133.7 117.56 136.1 117.8 ;
      RECT  136.1 116.46 136.61 116.7 ;
      RECT  134.63 115.67 135.17 116.22 ;
      RECT  133.49 118.9 134.63 118.52 ;
      RECT  135.89 119.14 136.1 119.07 ;
      RECT  136.1 118.28 136.61 118.04 ;
      RECT  133.7 119.38 136.1 119.14 ;
      RECT  136.1 119.14 136.3 119.07 ;
      RECT  135.89 118.35 136.1 118.28 ;
      RECT  136.61 119.38 136.82 119.14 ;
      POLYGON  135.17 118.9 135.17 118.52 135.72 118.52 135.72 118.59 136.1 118.59 136.1 118.83 135.72 118.83 135.72 118.9 135.17 118.9 ;
      RECT  136.61 118.9 136.82 118.52 ;
      RECT  133.49 120.17 133.7 119.62 ;
      RECT  133.7 120.17 134.63 119.62 ;
      RECT  134.63 118.9 135.17 118.52 ;
      RECT  136.61 118.28 136.82 118.04 ;
      RECT  135.17 120.17 136.82 119.62 ;
      RECT  133.49 119.38 133.7 119.14 ;
      RECT  136.1 118.35 136.3 118.28 ;
      POLYGON  136.47 118.9 136.47 118.83 136.1 118.83 136.1 118.59 136.47 118.59 136.47 118.52 136.61 118.52 136.61 118.9 136.47 118.9 ;
      RECT  133.49 118.28 133.7 118.04 ;
      RECT  133.7 118.28 136.1 118.04 ;
      RECT  136.1 119.38 136.61 119.14 ;
      RECT  134.63 120.17 135.17 119.62 ;
      RECT  133.49 120.89 134.63 121.27 ;
      RECT  135.89 120.65 136.1 120.72 ;
      RECT  136.1 121.51 136.61 121.75 ;
      RECT  133.7 120.41 136.1 120.65 ;
      RECT  136.1 120.65 136.3 120.72 ;
      RECT  135.89 121.44 136.1 121.51 ;
      RECT  136.61 120.41 136.82 120.65 ;
      POLYGON  135.17 120.89 135.17 121.27 135.72 121.27 135.72 121.2 136.1 121.2 136.1 120.96 135.72 120.96 135.72 120.89 135.17 120.89 ;
      RECT  136.61 120.89 136.82 121.27 ;
      RECT  133.49 119.62 133.7 120.17 ;
      RECT  133.7 119.62 134.63 120.17 ;
      RECT  134.63 120.89 135.17 121.27 ;
      RECT  136.61 121.51 136.82 121.75 ;
      RECT  135.17 119.62 136.82 120.17 ;
      RECT  133.49 120.41 133.7 120.65 ;
      RECT  136.1 121.44 136.3 121.51 ;
      POLYGON  136.47 120.89 136.47 120.96 136.1 120.96 136.1 121.2 136.47 121.2 136.47 121.27 136.61 121.27 136.61 120.89 136.47 120.89 ;
      RECT  133.49 121.51 133.7 121.75 ;
      RECT  133.7 121.51 136.1 121.75 ;
      RECT  136.1 120.41 136.61 120.65 ;
      RECT  134.63 119.62 135.17 120.17 ;
      RECT  133.49 122.85 134.63 122.47 ;
      RECT  135.89 123.09 136.1 123.02 ;
      RECT  136.1 122.23 136.61 121.99 ;
      RECT  133.7 123.33 136.1 123.09 ;
      RECT  136.1 123.09 136.3 123.02 ;
      RECT  135.89 122.3 136.1 122.23 ;
      RECT  136.61 123.33 136.82 123.09 ;
      POLYGON  135.17 122.85 135.17 122.47 135.72 122.47 135.72 122.54 136.1 122.54 136.1 122.78 135.72 122.78 135.72 122.85 135.17 122.85 ;
      RECT  136.61 122.85 136.82 122.47 ;
      RECT  133.49 124.12 133.7 123.57 ;
      RECT  133.7 124.12 134.63 123.57 ;
      RECT  134.63 122.85 135.17 122.47 ;
      RECT  136.61 122.23 136.82 121.99 ;
      RECT  135.17 124.12 136.82 123.57 ;
      RECT  133.49 123.33 133.7 123.09 ;
      RECT  136.1 122.3 136.3 122.23 ;
      POLYGON  136.47 122.85 136.47 122.78 136.1 122.78 136.1 122.54 136.47 122.54 136.47 122.47 136.61 122.47 136.61 122.85 136.47 122.85 ;
      RECT  133.49 122.23 133.7 121.99 ;
      RECT  133.7 122.23 136.1 121.99 ;
      RECT  136.1 123.33 136.61 123.09 ;
      RECT  134.63 124.12 135.17 123.57 ;
      RECT  140.15 93.24 139.01 93.62 ;
      RECT  137.75 93.0 137.54 93.07 ;
      RECT  137.54 93.86 137.03 94.1 ;
      RECT  139.94 92.76 137.54 93.0 ;
      RECT  137.54 93.0 137.34 93.07 ;
      RECT  137.75 93.79 137.54 93.86 ;
      RECT  137.03 92.76 136.82 93.0 ;
      POLYGON  138.47 93.24 138.47 93.62 137.92 93.62 137.92 93.55 137.54 93.55 137.54 93.31 137.92 93.31 137.92 93.24 138.47 93.24 ;
      RECT  137.03 93.24 136.82 93.62 ;
      RECT  140.15 91.97 139.94 92.52 ;
      RECT  139.94 91.97 139.01 92.52 ;
      RECT  139.01 93.24 138.47 93.62 ;
      RECT  137.03 93.86 136.82 94.1 ;
      RECT  138.47 91.97 136.82 92.52 ;
      RECT  140.15 92.76 139.94 93.0 ;
      RECT  137.54 93.79 137.34 93.86 ;
      POLYGON  137.17 93.24 137.17 93.31 137.54 93.31 137.54 93.55 137.17 93.55 137.17 93.62 137.03 93.62 137.03 93.24 137.17 93.24 ;
      RECT  140.15 93.86 139.94 94.1 ;
      RECT  139.94 93.86 137.54 94.1 ;
      RECT  137.54 92.76 137.03 93.0 ;
      RECT  139.01 91.97 138.47 92.52 ;
      RECT  140.15 95.2 139.01 94.82 ;
      RECT  137.75 95.44 137.54 95.37 ;
      RECT  137.54 94.58 137.03 94.34 ;
      RECT  139.94 95.68 137.54 95.44 ;
      RECT  137.54 95.44 137.34 95.37 ;
      RECT  137.75 94.65 137.54 94.58 ;
      RECT  137.03 95.68 136.82 95.44 ;
      POLYGON  138.47 95.2 138.47 94.82 137.92 94.82 137.92 94.89 137.54 94.89 137.54 95.13 137.92 95.13 137.92 95.2 138.47 95.2 ;
      RECT  137.03 95.2 136.82 94.82 ;
      RECT  140.15 96.47 139.94 95.92 ;
      RECT  139.94 96.47 139.01 95.92 ;
      RECT  139.01 95.2 138.47 94.82 ;
      RECT  137.03 94.58 136.82 94.34 ;
      RECT  138.47 96.47 136.82 95.92 ;
      RECT  140.15 95.68 139.94 95.44 ;
      RECT  137.54 94.65 137.34 94.58 ;
      POLYGON  137.17 95.2 137.17 95.13 137.54 95.13 137.54 94.89 137.17 94.89 137.17 94.82 137.03 94.82 137.03 95.2 137.17 95.2 ;
      RECT  140.15 94.58 139.94 94.34 ;
      RECT  139.94 94.58 137.54 94.34 ;
      RECT  137.54 95.68 137.03 95.44 ;
      RECT  139.01 96.47 138.47 95.92 ;
      RECT  140.15 97.19 139.01 97.57 ;
      RECT  137.75 96.95 137.54 97.02 ;
      RECT  137.54 97.81 137.03 98.05 ;
      RECT  139.94 96.71 137.54 96.95 ;
      RECT  137.54 96.95 137.34 97.02 ;
      RECT  137.75 97.74 137.54 97.81 ;
      RECT  137.03 96.71 136.82 96.95 ;
      POLYGON  138.47 97.19 138.47 97.57 137.92 97.57 137.92 97.5 137.54 97.5 137.54 97.26 137.92 97.26 137.92 97.19 138.47 97.19 ;
      RECT  137.03 97.19 136.82 97.57 ;
      RECT  140.15 95.92 139.94 96.47 ;
      RECT  139.94 95.92 139.01 96.47 ;
      RECT  139.01 97.19 138.47 97.57 ;
      RECT  137.03 97.81 136.82 98.05 ;
      RECT  138.47 95.92 136.82 96.47 ;
      RECT  140.15 96.71 139.94 96.95 ;
      RECT  137.54 97.74 137.34 97.81 ;
      POLYGON  137.17 97.19 137.17 97.26 137.54 97.26 137.54 97.5 137.17 97.5 137.17 97.57 137.03 97.57 137.03 97.19 137.17 97.19 ;
      RECT  140.15 97.81 139.94 98.05 ;
      RECT  139.94 97.81 137.54 98.05 ;
      RECT  137.54 96.71 137.03 96.95 ;
      RECT  139.01 95.92 138.47 96.47 ;
      RECT  140.15 99.15 139.01 98.77 ;
      RECT  137.75 99.39 137.54 99.32 ;
      RECT  137.54 98.53 137.03 98.29 ;
      RECT  139.94 99.63 137.54 99.39 ;
      RECT  137.54 99.39 137.34 99.32 ;
      RECT  137.75 98.6 137.54 98.53 ;
      RECT  137.03 99.63 136.82 99.39 ;
      POLYGON  138.47 99.15 138.47 98.77 137.92 98.77 137.92 98.84 137.54 98.84 137.54 99.08 137.92 99.08 137.92 99.15 138.47 99.15 ;
      RECT  137.03 99.15 136.82 98.77 ;
      RECT  140.15 100.42 139.94 99.87 ;
      RECT  139.94 100.42 139.01 99.87 ;
      RECT  139.01 99.15 138.47 98.77 ;
      RECT  137.03 98.53 136.82 98.29 ;
      RECT  138.47 100.42 136.82 99.87 ;
      RECT  140.15 99.63 139.94 99.39 ;
      RECT  137.54 98.6 137.34 98.53 ;
      POLYGON  137.17 99.15 137.17 99.08 137.54 99.08 137.54 98.84 137.17 98.84 137.17 98.77 137.03 98.77 137.03 99.15 137.17 99.15 ;
      RECT  140.15 98.53 139.94 98.29 ;
      RECT  139.94 98.53 137.54 98.29 ;
      RECT  137.54 99.63 137.03 99.39 ;
      RECT  139.01 100.42 138.47 99.87 ;
      RECT  140.15 101.14 139.01 101.52 ;
      RECT  137.75 100.9 137.54 100.97 ;
      RECT  137.54 101.76 137.03 102.0 ;
      RECT  139.94 100.66 137.54 100.9 ;
      RECT  137.54 100.9 137.34 100.97 ;
      RECT  137.75 101.69 137.54 101.76 ;
      RECT  137.03 100.66 136.82 100.9 ;
      POLYGON  138.47 101.14 138.47 101.52 137.92 101.52 137.92 101.45 137.54 101.45 137.54 101.21 137.92 101.21 137.92 101.14 138.47 101.14 ;
      RECT  137.03 101.14 136.82 101.52 ;
      RECT  140.15 99.87 139.94 100.42 ;
      RECT  139.94 99.87 139.01 100.42 ;
      RECT  139.01 101.14 138.47 101.52 ;
      RECT  137.03 101.76 136.82 102.0 ;
      RECT  138.47 99.87 136.82 100.42 ;
      RECT  140.15 100.66 139.94 100.9 ;
      RECT  137.54 101.69 137.34 101.76 ;
      POLYGON  137.17 101.14 137.17 101.21 137.54 101.21 137.54 101.45 137.17 101.45 137.17 101.52 137.03 101.52 137.03 101.14 137.17 101.14 ;
      RECT  140.15 101.76 139.94 102.0 ;
      RECT  139.94 101.76 137.54 102.0 ;
      RECT  137.54 100.66 137.03 100.9 ;
      RECT  139.01 99.87 138.47 100.42 ;
      RECT  140.15 103.1 139.01 102.72 ;
      RECT  137.75 103.34 137.54 103.27 ;
      RECT  137.54 102.48 137.03 102.24 ;
      RECT  139.94 103.58 137.54 103.34 ;
      RECT  137.54 103.34 137.34 103.27 ;
      RECT  137.75 102.55 137.54 102.48 ;
      RECT  137.03 103.58 136.82 103.34 ;
      POLYGON  138.47 103.1 138.47 102.72 137.92 102.72 137.92 102.79 137.54 102.79 137.54 103.03 137.92 103.03 137.92 103.1 138.47 103.1 ;
      RECT  137.03 103.1 136.82 102.72 ;
      RECT  140.15 104.37 139.94 103.82 ;
      RECT  139.94 104.37 139.01 103.82 ;
      RECT  139.01 103.1 138.47 102.72 ;
      RECT  137.03 102.48 136.82 102.24 ;
      RECT  138.47 104.37 136.82 103.82 ;
      RECT  140.15 103.58 139.94 103.34 ;
      RECT  137.54 102.55 137.34 102.48 ;
      POLYGON  137.17 103.1 137.17 103.03 137.54 103.03 137.54 102.79 137.17 102.79 137.17 102.72 137.03 102.72 137.03 103.1 137.17 103.1 ;
      RECT  140.15 102.48 139.94 102.24 ;
      RECT  139.94 102.48 137.54 102.24 ;
      RECT  137.54 103.58 137.03 103.34 ;
      RECT  139.01 104.37 138.47 103.82 ;
      RECT  140.15 105.09 139.01 105.47 ;
      RECT  137.75 104.85 137.54 104.92 ;
      RECT  137.54 105.71 137.03 105.95 ;
      RECT  139.94 104.61 137.54 104.85 ;
      RECT  137.54 104.85 137.34 104.92 ;
      RECT  137.75 105.64 137.54 105.71 ;
      RECT  137.03 104.61 136.82 104.85 ;
      POLYGON  138.47 105.09 138.47 105.47 137.92 105.47 137.92 105.4 137.54 105.4 137.54 105.16 137.92 105.16 137.92 105.09 138.47 105.09 ;
      RECT  137.03 105.09 136.82 105.47 ;
      RECT  140.15 103.82 139.94 104.37 ;
      RECT  139.94 103.82 139.01 104.37 ;
      RECT  139.01 105.09 138.47 105.47 ;
      RECT  137.03 105.71 136.82 105.95 ;
      RECT  138.47 103.82 136.82 104.37 ;
      RECT  140.15 104.61 139.94 104.85 ;
      RECT  137.54 105.64 137.34 105.71 ;
      POLYGON  137.17 105.09 137.17 105.16 137.54 105.16 137.54 105.4 137.17 105.4 137.17 105.47 137.03 105.47 137.03 105.09 137.17 105.09 ;
      RECT  140.15 105.71 139.94 105.95 ;
      RECT  139.94 105.71 137.54 105.95 ;
      RECT  137.54 104.61 137.03 104.85 ;
      RECT  139.01 103.82 138.47 104.37 ;
      RECT  140.15 107.05 139.01 106.67 ;
      RECT  137.75 107.29 137.54 107.22 ;
      RECT  137.54 106.43 137.03 106.19 ;
      RECT  139.94 107.53 137.54 107.29 ;
      RECT  137.54 107.29 137.34 107.22 ;
      RECT  137.75 106.5 137.54 106.43 ;
      RECT  137.03 107.53 136.82 107.29 ;
      POLYGON  138.47 107.05 138.47 106.67 137.92 106.67 137.92 106.74 137.54 106.74 137.54 106.98 137.92 106.98 137.92 107.05 138.47 107.05 ;
      RECT  137.03 107.05 136.82 106.67 ;
      RECT  140.15 108.32 139.94 107.77 ;
      RECT  139.94 108.32 139.01 107.77 ;
      RECT  139.01 107.05 138.47 106.67 ;
      RECT  137.03 106.43 136.82 106.19 ;
      RECT  138.47 108.32 136.82 107.77 ;
      RECT  140.15 107.53 139.94 107.29 ;
      RECT  137.54 106.5 137.34 106.43 ;
      POLYGON  137.17 107.05 137.17 106.98 137.54 106.98 137.54 106.74 137.17 106.74 137.17 106.67 137.03 106.67 137.03 107.05 137.17 107.05 ;
      RECT  140.15 106.43 139.94 106.19 ;
      RECT  139.94 106.43 137.54 106.19 ;
      RECT  137.54 107.53 137.03 107.29 ;
      RECT  139.01 108.32 138.47 107.77 ;
      RECT  140.15 109.04 139.01 109.42 ;
      RECT  137.75 108.8 137.54 108.87 ;
      RECT  137.54 109.66 137.03 109.9 ;
      RECT  139.94 108.56 137.54 108.8 ;
      RECT  137.54 108.8 137.34 108.87 ;
      RECT  137.75 109.59 137.54 109.66 ;
      RECT  137.03 108.56 136.82 108.8 ;
      POLYGON  138.47 109.04 138.47 109.42 137.92 109.42 137.92 109.35 137.54 109.35 137.54 109.11 137.92 109.11 137.92 109.04 138.47 109.04 ;
      RECT  137.03 109.04 136.82 109.42 ;
      RECT  140.15 107.77 139.94 108.32 ;
      RECT  139.94 107.77 139.01 108.32 ;
      RECT  139.01 109.04 138.47 109.42 ;
      RECT  137.03 109.66 136.82 109.9 ;
      RECT  138.47 107.77 136.82 108.32 ;
      RECT  140.15 108.56 139.94 108.8 ;
      RECT  137.54 109.59 137.34 109.66 ;
      POLYGON  137.17 109.04 137.17 109.11 137.54 109.11 137.54 109.35 137.17 109.35 137.17 109.42 137.03 109.42 137.03 109.04 137.17 109.04 ;
      RECT  140.15 109.66 139.94 109.9 ;
      RECT  139.94 109.66 137.54 109.9 ;
      RECT  137.54 108.56 137.03 108.8 ;
      RECT  139.01 107.77 138.47 108.32 ;
      RECT  140.15 111.0 139.01 110.62 ;
      RECT  137.75 111.24 137.54 111.17 ;
      RECT  137.54 110.38 137.03 110.14 ;
      RECT  139.94 111.48 137.54 111.24 ;
      RECT  137.54 111.24 137.34 111.17 ;
      RECT  137.75 110.45 137.54 110.38 ;
      RECT  137.03 111.48 136.82 111.24 ;
      POLYGON  138.47 111.0 138.47 110.62 137.92 110.62 137.92 110.69 137.54 110.69 137.54 110.93 137.92 110.93 137.92 111.0 138.47 111.0 ;
      RECT  137.03 111.0 136.82 110.62 ;
      RECT  140.15 112.27 139.94 111.72 ;
      RECT  139.94 112.27 139.01 111.72 ;
      RECT  139.01 111.0 138.47 110.62 ;
      RECT  137.03 110.38 136.82 110.14 ;
      RECT  138.47 112.27 136.82 111.72 ;
      RECT  140.15 111.48 139.94 111.24 ;
      RECT  137.54 110.45 137.34 110.38 ;
      POLYGON  137.17 111.0 137.17 110.93 137.54 110.93 137.54 110.69 137.17 110.69 137.17 110.62 137.03 110.62 137.03 111.0 137.17 111.0 ;
      RECT  140.15 110.38 139.94 110.14 ;
      RECT  139.94 110.38 137.54 110.14 ;
      RECT  137.54 111.48 137.03 111.24 ;
      RECT  139.01 112.27 138.47 111.72 ;
      RECT  140.15 112.99 139.01 113.37 ;
      RECT  137.75 112.75 137.54 112.82 ;
      RECT  137.54 113.61 137.03 113.85 ;
      RECT  139.94 112.51 137.54 112.75 ;
      RECT  137.54 112.75 137.34 112.82 ;
      RECT  137.75 113.54 137.54 113.61 ;
      RECT  137.03 112.51 136.82 112.75 ;
      POLYGON  138.47 112.99 138.47 113.37 137.92 113.37 137.92 113.3 137.54 113.3 137.54 113.06 137.92 113.06 137.92 112.99 138.47 112.99 ;
      RECT  137.03 112.99 136.82 113.37 ;
      RECT  140.15 111.72 139.94 112.27 ;
      RECT  139.94 111.72 139.01 112.27 ;
      RECT  139.01 112.99 138.47 113.37 ;
      RECT  137.03 113.61 136.82 113.85 ;
      RECT  138.47 111.72 136.82 112.27 ;
      RECT  140.15 112.51 139.94 112.75 ;
      RECT  137.54 113.54 137.34 113.61 ;
      POLYGON  137.17 112.99 137.17 113.06 137.54 113.06 137.54 113.3 137.17 113.3 137.17 113.37 137.03 113.37 137.03 112.99 137.17 112.99 ;
      RECT  140.15 113.61 139.94 113.85 ;
      RECT  139.94 113.61 137.54 113.85 ;
      RECT  137.54 112.51 137.03 112.75 ;
      RECT  139.01 111.72 138.47 112.27 ;
      RECT  140.15 114.95 139.01 114.57 ;
      RECT  137.75 115.19 137.54 115.12 ;
      RECT  137.54 114.33 137.03 114.09 ;
      RECT  139.94 115.43 137.54 115.19 ;
      RECT  137.54 115.19 137.34 115.12 ;
      RECT  137.75 114.4 137.54 114.33 ;
      RECT  137.03 115.43 136.82 115.19 ;
      POLYGON  138.47 114.95 138.47 114.57 137.92 114.57 137.92 114.64 137.54 114.64 137.54 114.88 137.92 114.88 137.92 114.95 138.47 114.95 ;
      RECT  137.03 114.95 136.82 114.57 ;
      RECT  140.15 116.22 139.94 115.67 ;
      RECT  139.94 116.22 139.01 115.67 ;
      RECT  139.01 114.95 138.47 114.57 ;
      RECT  137.03 114.33 136.82 114.09 ;
      RECT  138.47 116.22 136.82 115.67 ;
      RECT  140.15 115.43 139.94 115.19 ;
      RECT  137.54 114.4 137.34 114.33 ;
      POLYGON  137.17 114.95 137.17 114.88 137.54 114.88 137.54 114.64 137.17 114.64 137.17 114.57 137.03 114.57 137.03 114.95 137.17 114.95 ;
      RECT  140.15 114.33 139.94 114.09 ;
      RECT  139.94 114.33 137.54 114.09 ;
      RECT  137.54 115.43 137.03 115.19 ;
      RECT  139.01 116.22 138.47 115.67 ;
      RECT  140.15 116.94 139.01 117.32 ;
      RECT  137.75 116.7 137.54 116.77 ;
      RECT  137.54 117.56 137.03 117.8 ;
      RECT  139.94 116.46 137.54 116.7 ;
      RECT  137.54 116.7 137.34 116.77 ;
      RECT  137.75 117.49 137.54 117.56 ;
      RECT  137.03 116.46 136.82 116.7 ;
      POLYGON  138.47 116.94 138.47 117.32 137.92 117.32 137.92 117.25 137.54 117.25 137.54 117.01 137.92 117.01 137.92 116.94 138.47 116.94 ;
      RECT  137.03 116.94 136.82 117.32 ;
      RECT  140.15 115.67 139.94 116.22 ;
      RECT  139.94 115.67 139.01 116.22 ;
      RECT  139.01 116.94 138.47 117.32 ;
      RECT  137.03 117.56 136.82 117.8 ;
      RECT  138.47 115.67 136.82 116.22 ;
      RECT  140.15 116.46 139.94 116.7 ;
      RECT  137.54 117.49 137.34 117.56 ;
      POLYGON  137.17 116.94 137.17 117.01 137.54 117.01 137.54 117.25 137.17 117.25 137.17 117.32 137.03 117.32 137.03 116.94 137.17 116.94 ;
      RECT  140.15 117.56 139.94 117.8 ;
      RECT  139.94 117.56 137.54 117.8 ;
      RECT  137.54 116.46 137.03 116.7 ;
      RECT  139.01 115.67 138.47 116.22 ;
      RECT  140.15 118.9 139.01 118.52 ;
      RECT  137.75 119.14 137.54 119.07 ;
      RECT  137.54 118.28 137.03 118.04 ;
      RECT  139.94 119.38 137.54 119.14 ;
      RECT  137.54 119.14 137.34 119.07 ;
      RECT  137.75 118.35 137.54 118.28 ;
      RECT  137.03 119.38 136.82 119.14 ;
      POLYGON  138.47 118.9 138.47 118.52 137.92 118.52 137.92 118.59 137.54 118.59 137.54 118.83 137.92 118.83 137.92 118.9 138.47 118.9 ;
      RECT  137.03 118.9 136.82 118.52 ;
      RECT  140.15 120.17 139.94 119.62 ;
      RECT  139.94 120.17 139.01 119.62 ;
      RECT  139.01 118.9 138.47 118.52 ;
      RECT  137.03 118.28 136.82 118.04 ;
      RECT  138.47 120.17 136.82 119.62 ;
      RECT  140.15 119.38 139.94 119.14 ;
      RECT  137.54 118.35 137.34 118.28 ;
      POLYGON  137.17 118.9 137.17 118.83 137.54 118.83 137.54 118.59 137.17 118.59 137.17 118.52 137.03 118.52 137.03 118.9 137.17 118.9 ;
      RECT  140.15 118.28 139.94 118.04 ;
      RECT  139.94 118.28 137.54 118.04 ;
      RECT  137.54 119.38 137.03 119.14 ;
      RECT  139.01 120.17 138.47 119.62 ;
      RECT  140.15 120.89 139.01 121.27 ;
      RECT  137.75 120.65 137.54 120.72 ;
      RECT  137.54 121.51 137.03 121.75 ;
      RECT  139.94 120.41 137.54 120.65 ;
      RECT  137.54 120.65 137.34 120.72 ;
      RECT  137.75 121.44 137.54 121.51 ;
      RECT  137.03 120.41 136.82 120.65 ;
      POLYGON  138.47 120.89 138.47 121.27 137.92 121.27 137.92 121.2 137.54 121.2 137.54 120.96 137.92 120.96 137.92 120.89 138.47 120.89 ;
      RECT  137.03 120.89 136.82 121.27 ;
      RECT  140.15 119.62 139.94 120.17 ;
      RECT  139.94 119.62 139.01 120.17 ;
      RECT  139.01 120.89 138.47 121.27 ;
      RECT  137.03 121.51 136.82 121.75 ;
      RECT  138.47 119.62 136.82 120.17 ;
      RECT  140.15 120.41 139.94 120.65 ;
      RECT  137.54 121.44 137.34 121.51 ;
      POLYGON  137.17 120.89 137.17 120.96 137.54 120.96 137.54 121.2 137.17 121.2 137.17 121.27 137.03 121.27 137.03 120.89 137.17 120.89 ;
      RECT  140.15 121.51 139.94 121.75 ;
      RECT  139.94 121.51 137.54 121.75 ;
      RECT  137.54 120.41 137.03 120.65 ;
      RECT  139.01 119.62 138.47 120.17 ;
      RECT  140.15 122.85 139.01 122.47 ;
      RECT  137.75 123.09 137.54 123.02 ;
      RECT  137.54 122.23 137.03 121.99 ;
      RECT  139.94 123.33 137.54 123.09 ;
      RECT  137.54 123.09 137.34 123.02 ;
      RECT  137.75 122.3 137.54 122.23 ;
      RECT  137.03 123.33 136.82 123.09 ;
      POLYGON  138.47 122.85 138.47 122.47 137.92 122.47 137.92 122.54 137.54 122.54 137.54 122.78 137.92 122.78 137.92 122.85 138.47 122.85 ;
      RECT  137.03 122.85 136.82 122.47 ;
      RECT  140.15 124.12 139.94 123.57 ;
      RECT  139.94 124.12 139.01 123.57 ;
      RECT  139.01 122.85 138.47 122.47 ;
      RECT  137.03 122.23 136.82 121.99 ;
      RECT  138.47 124.12 136.82 123.57 ;
      RECT  140.15 123.33 139.94 123.09 ;
      RECT  137.54 122.3 137.34 122.23 ;
      POLYGON  137.17 122.85 137.17 122.78 137.54 122.78 137.54 122.54 137.17 122.54 137.17 122.47 137.03 122.47 137.03 122.85 137.17 122.85 ;
      RECT  140.15 122.23 139.94 121.99 ;
      RECT  139.94 122.23 137.54 121.99 ;
      RECT  137.54 123.33 137.03 123.09 ;
      RECT  139.01 124.12 138.47 123.57 ;
      RECT  139.73 93.24 140.87 93.62 ;
      RECT  142.13 93.0 142.34 93.07 ;
      RECT  142.34 93.86 142.85 94.1 ;
      RECT  139.94 92.76 142.34 93.0 ;
      RECT  142.34 93.0 142.54 93.07 ;
      RECT  142.13 93.79 142.34 93.86 ;
      RECT  142.85 92.76 143.06 93.0 ;
      POLYGON  141.41 93.24 141.41 93.62 141.96 93.62 141.96 93.55 142.34 93.55 142.34 93.31 141.96 93.31 141.96 93.24 141.41 93.24 ;
      RECT  142.85 93.24 143.06 93.62 ;
      RECT  139.73 91.97 139.94 92.52 ;
      RECT  139.94 91.97 140.87 92.52 ;
      RECT  140.87 93.24 141.41 93.62 ;
      RECT  142.85 93.86 143.06 94.1 ;
      RECT  141.41 91.97 143.06 92.52 ;
      RECT  139.73 92.76 139.94 93.0 ;
      RECT  142.34 93.79 142.54 93.86 ;
      POLYGON  142.71 93.24 142.71 93.31 142.34 93.31 142.34 93.55 142.71 93.55 142.71 93.62 142.85 93.62 142.85 93.24 142.71 93.24 ;
      RECT  139.73 93.86 139.94 94.1 ;
      RECT  139.94 93.86 142.34 94.1 ;
      RECT  142.34 92.76 142.85 93.0 ;
      RECT  140.87 91.97 141.41 92.52 ;
      RECT  139.73 95.2 140.87 94.82 ;
      RECT  142.13 95.44 142.34 95.37 ;
      RECT  142.34 94.58 142.85 94.34 ;
      RECT  139.94 95.68 142.34 95.44 ;
      RECT  142.34 95.44 142.54 95.37 ;
      RECT  142.13 94.65 142.34 94.58 ;
      RECT  142.85 95.68 143.06 95.44 ;
      POLYGON  141.41 95.2 141.41 94.82 141.96 94.82 141.96 94.89 142.34 94.89 142.34 95.13 141.96 95.13 141.96 95.2 141.41 95.2 ;
      RECT  142.85 95.2 143.06 94.82 ;
      RECT  139.73 96.47 139.94 95.92 ;
      RECT  139.94 96.47 140.87 95.92 ;
      RECT  140.87 95.2 141.41 94.82 ;
      RECT  142.85 94.58 143.06 94.34 ;
      RECT  141.41 96.47 143.06 95.92 ;
      RECT  139.73 95.68 139.94 95.44 ;
      RECT  142.34 94.65 142.54 94.58 ;
      POLYGON  142.71 95.2 142.71 95.13 142.34 95.13 142.34 94.89 142.71 94.89 142.71 94.82 142.85 94.82 142.85 95.2 142.71 95.2 ;
      RECT  139.73 94.58 139.94 94.34 ;
      RECT  139.94 94.58 142.34 94.34 ;
      RECT  142.34 95.68 142.85 95.44 ;
      RECT  140.87 96.47 141.41 95.92 ;
      RECT  139.73 97.19 140.87 97.57 ;
      RECT  142.13 96.95 142.34 97.02 ;
      RECT  142.34 97.81 142.85 98.05 ;
      RECT  139.94 96.71 142.34 96.95 ;
      RECT  142.34 96.95 142.54 97.02 ;
      RECT  142.13 97.74 142.34 97.81 ;
      RECT  142.85 96.71 143.06 96.95 ;
      POLYGON  141.41 97.19 141.41 97.57 141.96 97.57 141.96 97.5 142.34 97.5 142.34 97.26 141.96 97.26 141.96 97.19 141.41 97.19 ;
      RECT  142.85 97.19 143.06 97.57 ;
      RECT  139.73 95.92 139.94 96.47 ;
      RECT  139.94 95.92 140.87 96.47 ;
      RECT  140.87 97.19 141.41 97.57 ;
      RECT  142.85 97.81 143.06 98.05 ;
      RECT  141.41 95.92 143.06 96.47 ;
      RECT  139.73 96.71 139.94 96.95 ;
      RECT  142.34 97.74 142.54 97.81 ;
      POLYGON  142.71 97.19 142.71 97.26 142.34 97.26 142.34 97.5 142.71 97.5 142.71 97.57 142.85 97.57 142.85 97.19 142.71 97.19 ;
      RECT  139.73 97.81 139.94 98.05 ;
      RECT  139.94 97.81 142.34 98.05 ;
      RECT  142.34 96.71 142.85 96.95 ;
      RECT  140.87 95.92 141.41 96.47 ;
      RECT  139.73 99.15 140.87 98.77 ;
      RECT  142.13 99.39 142.34 99.32 ;
      RECT  142.34 98.53 142.85 98.29 ;
      RECT  139.94 99.63 142.34 99.39 ;
      RECT  142.34 99.39 142.54 99.32 ;
      RECT  142.13 98.6 142.34 98.53 ;
      RECT  142.85 99.63 143.06 99.39 ;
      POLYGON  141.41 99.15 141.41 98.77 141.96 98.77 141.96 98.84 142.34 98.84 142.34 99.08 141.96 99.08 141.96 99.15 141.41 99.15 ;
      RECT  142.85 99.15 143.06 98.77 ;
      RECT  139.73 100.42 139.94 99.87 ;
      RECT  139.94 100.42 140.87 99.87 ;
      RECT  140.87 99.15 141.41 98.77 ;
      RECT  142.85 98.53 143.06 98.29 ;
      RECT  141.41 100.42 143.06 99.87 ;
      RECT  139.73 99.63 139.94 99.39 ;
      RECT  142.34 98.6 142.54 98.53 ;
      POLYGON  142.71 99.15 142.71 99.08 142.34 99.08 142.34 98.84 142.71 98.84 142.71 98.77 142.85 98.77 142.85 99.15 142.71 99.15 ;
      RECT  139.73 98.53 139.94 98.29 ;
      RECT  139.94 98.53 142.34 98.29 ;
      RECT  142.34 99.63 142.85 99.39 ;
      RECT  140.87 100.42 141.41 99.87 ;
      RECT  139.73 101.14 140.87 101.52 ;
      RECT  142.13 100.9 142.34 100.97 ;
      RECT  142.34 101.76 142.85 102.0 ;
      RECT  139.94 100.66 142.34 100.9 ;
      RECT  142.34 100.9 142.54 100.97 ;
      RECT  142.13 101.69 142.34 101.76 ;
      RECT  142.85 100.66 143.06 100.9 ;
      POLYGON  141.41 101.14 141.41 101.52 141.96 101.52 141.96 101.45 142.34 101.45 142.34 101.21 141.96 101.21 141.96 101.14 141.41 101.14 ;
      RECT  142.85 101.14 143.06 101.52 ;
      RECT  139.73 99.87 139.94 100.42 ;
      RECT  139.94 99.87 140.87 100.42 ;
      RECT  140.87 101.14 141.41 101.52 ;
      RECT  142.85 101.76 143.06 102.0 ;
      RECT  141.41 99.87 143.06 100.42 ;
      RECT  139.73 100.66 139.94 100.9 ;
      RECT  142.34 101.69 142.54 101.76 ;
      POLYGON  142.71 101.14 142.71 101.21 142.34 101.21 142.34 101.45 142.71 101.45 142.71 101.52 142.85 101.52 142.85 101.14 142.71 101.14 ;
      RECT  139.73 101.76 139.94 102.0 ;
      RECT  139.94 101.76 142.34 102.0 ;
      RECT  142.34 100.66 142.85 100.9 ;
      RECT  140.87 99.87 141.41 100.42 ;
      RECT  139.73 103.1 140.87 102.72 ;
      RECT  142.13 103.34 142.34 103.27 ;
      RECT  142.34 102.48 142.85 102.24 ;
      RECT  139.94 103.58 142.34 103.34 ;
      RECT  142.34 103.34 142.54 103.27 ;
      RECT  142.13 102.55 142.34 102.48 ;
      RECT  142.85 103.58 143.06 103.34 ;
      POLYGON  141.41 103.1 141.41 102.72 141.96 102.72 141.96 102.79 142.34 102.79 142.34 103.03 141.96 103.03 141.96 103.1 141.41 103.1 ;
      RECT  142.85 103.1 143.06 102.72 ;
      RECT  139.73 104.37 139.94 103.82 ;
      RECT  139.94 104.37 140.87 103.82 ;
      RECT  140.87 103.1 141.41 102.72 ;
      RECT  142.85 102.48 143.06 102.24 ;
      RECT  141.41 104.37 143.06 103.82 ;
      RECT  139.73 103.58 139.94 103.34 ;
      RECT  142.34 102.55 142.54 102.48 ;
      POLYGON  142.71 103.1 142.71 103.03 142.34 103.03 142.34 102.79 142.71 102.79 142.71 102.72 142.85 102.72 142.85 103.1 142.71 103.1 ;
      RECT  139.73 102.48 139.94 102.24 ;
      RECT  139.94 102.48 142.34 102.24 ;
      RECT  142.34 103.58 142.85 103.34 ;
      RECT  140.87 104.37 141.41 103.82 ;
      RECT  139.73 105.09 140.87 105.47 ;
      RECT  142.13 104.85 142.34 104.92 ;
      RECT  142.34 105.71 142.85 105.95 ;
      RECT  139.94 104.61 142.34 104.85 ;
      RECT  142.34 104.85 142.54 104.92 ;
      RECT  142.13 105.64 142.34 105.71 ;
      RECT  142.85 104.61 143.06 104.85 ;
      POLYGON  141.41 105.09 141.41 105.47 141.96 105.47 141.96 105.4 142.34 105.4 142.34 105.16 141.96 105.16 141.96 105.09 141.41 105.09 ;
      RECT  142.85 105.09 143.06 105.47 ;
      RECT  139.73 103.82 139.94 104.37 ;
      RECT  139.94 103.82 140.87 104.37 ;
      RECT  140.87 105.09 141.41 105.47 ;
      RECT  142.85 105.71 143.06 105.95 ;
      RECT  141.41 103.82 143.06 104.37 ;
      RECT  139.73 104.61 139.94 104.85 ;
      RECT  142.34 105.64 142.54 105.71 ;
      POLYGON  142.71 105.09 142.71 105.16 142.34 105.16 142.34 105.4 142.71 105.4 142.71 105.47 142.85 105.47 142.85 105.09 142.71 105.09 ;
      RECT  139.73 105.71 139.94 105.95 ;
      RECT  139.94 105.71 142.34 105.95 ;
      RECT  142.34 104.61 142.85 104.85 ;
      RECT  140.87 103.82 141.41 104.37 ;
      RECT  139.73 107.05 140.87 106.67 ;
      RECT  142.13 107.29 142.34 107.22 ;
      RECT  142.34 106.43 142.85 106.19 ;
      RECT  139.94 107.53 142.34 107.29 ;
      RECT  142.34 107.29 142.54 107.22 ;
      RECT  142.13 106.5 142.34 106.43 ;
      RECT  142.85 107.53 143.06 107.29 ;
      POLYGON  141.41 107.05 141.41 106.67 141.96 106.67 141.96 106.74 142.34 106.74 142.34 106.98 141.96 106.98 141.96 107.05 141.41 107.05 ;
      RECT  142.85 107.05 143.06 106.67 ;
      RECT  139.73 108.32 139.94 107.77 ;
      RECT  139.94 108.32 140.87 107.77 ;
      RECT  140.87 107.05 141.41 106.67 ;
      RECT  142.85 106.43 143.06 106.19 ;
      RECT  141.41 108.32 143.06 107.77 ;
      RECT  139.73 107.53 139.94 107.29 ;
      RECT  142.34 106.5 142.54 106.43 ;
      POLYGON  142.71 107.05 142.71 106.98 142.34 106.98 142.34 106.74 142.71 106.74 142.71 106.67 142.85 106.67 142.85 107.05 142.71 107.05 ;
      RECT  139.73 106.43 139.94 106.19 ;
      RECT  139.94 106.43 142.34 106.19 ;
      RECT  142.34 107.53 142.85 107.29 ;
      RECT  140.87 108.32 141.41 107.77 ;
      RECT  139.73 109.04 140.87 109.42 ;
      RECT  142.13 108.8 142.34 108.87 ;
      RECT  142.34 109.66 142.85 109.9 ;
      RECT  139.94 108.56 142.34 108.8 ;
      RECT  142.34 108.8 142.54 108.87 ;
      RECT  142.13 109.59 142.34 109.66 ;
      RECT  142.85 108.56 143.06 108.8 ;
      POLYGON  141.41 109.04 141.41 109.42 141.96 109.42 141.96 109.35 142.34 109.35 142.34 109.11 141.96 109.11 141.96 109.04 141.41 109.04 ;
      RECT  142.85 109.04 143.06 109.42 ;
      RECT  139.73 107.77 139.94 108.32 ;
      RECT  139.94 107.77 140.87 108.32 ;
      RECT  140.87 109.04 141.41 109.42 ;
      RECT  142.85 109.66 143.06 109.9 ;
      RECT  141.41 107.77 143.06 108.32 ;
      RECT  139.73 108.56 139.94 108.8 ;
      RECT  142.34 109.59 142.54 109.66 ;
      POLYGON  142.71 109.04 142.71 109.11 142.34 109.11 142.34 109.35 142.71 109.35 142.71 109.42 142.85 109.42 142.85 109.04 142.71 109.04 ;
      RECT  139.73 109.66 139.94 109.9 ;
      RECT  139.94 109.66 142.34 109.9 ;
      RECT  142.34 108.56 142.85 108.8 ;
      RECT  140.87 107.77 141.41 108.32 ;
      RECT  139.73 111.0 140.87 110.62 ;
      RECT  142.13 111.24 142.34 111.17 ;
      RECT  142.34 110.38 142.85 110.14 ;
      RECT  139.94 111.48 142.34 111.24 ;
      RECT  142.34 111.24 142.54 111.17 ;
      RECT  142.13 110.45 142.34 110.38 ;
      RECT  142.85 111.48 143.06 111.24 ;
      POLYGON  141.41 111.0 141.41 110.62 141.96 110.62 141.96 110.69 142.34 110.69 142.34 110.93 141.96 110.93 141.96 111.0 141.41 111.0 ;
      RECT  142.85 111.0 143.06 110.62 ;
      RECT  139.73 112.27 139.94 111.72 ;
      RECT  139.94 112.27 140.87 111.72 ;
      RECT  140.87 111.0 141.41 110.62 ;
      RECT  142.85 110.38 143.06 110.14 ;
      RECT  141.41 112.27 143.06 111.72 ;
      RECT  139.73 111.48 139.94 111.24 ;
      RECT  142.34 110.45 142.54 110.38 ;
      POLYGON  142.71 111.0 142.71 110.93 142.34 110.93 142.34 110.69 142.71 110.69 142.71 110.62 142.85 110.62 142.85 111.0 142.71 111.0 ;
      RECT  139.73 110.38 139.94 110.14 ;
      RECT  139.94 110.38 142.34 110.14 ;
      RECT  142.34 111.48 142.85 111.24 ;
      RECT  140.87 112.27 141.41 111.72 ;
      RECT  139.73 112.99 140.87 113.37 ;
      RECT  142.13 112.75 142.34 112.82 ;
      RECT  142.34 113.61 142.85 113.85 ;
      RECT  139.94 112.51 142.34 112.75 ;
      RECT  142.34 112.75 142.54 112.82 ;
      RECT  142.13 113.54 142.34 113.61 ;
      RECT  142.85 112.51 143.06 112.75 ;
      POLYGON  141.41 112.99 141.41 113.37 141.96 113.37 141.96 113.3 142.34 113.3 142.34 113.06 141.96 113.06 141.96 112.99 141.41 112.99 ;
      RECT  142.85 112.99 143.06 113.37 ;
      RECT  139.73 111.72 139.94 112.27 ;
      RECT  139.94 111.72 140.87 112.27 ;
      RECT  140.87 112.99 141.41 113.37 ;
      RECT  142.85 113.61 143.06 113.85 ;
      RECT  141.41 111.72 143.06 112.27 ;
      RECT  139.73 112.51 139.94 112.75 ;
      RECT  142.34 113.54 142.54 113.61 ;
      POLYGON  142.71 112.99 142.71 113.06 142.34 113.06 142.34 113.3 142.71 113.3 142.71 113.37 142.85 113.37 142.85 112.99 142.71 112.99 ;
      RECT  139.73 113.61 139.94 113.85 ;
      RECT  139.94 113.61 142.34 113.85 ;
      RECT  142.34 112.51 142.85 112.75 ;
      RECT  140.87 111.72 141.41 112.27 ;
      RECT  139.73 114.95 140.87 114.57 ;
      RECT  142.13 115.19 142.34 115.12 ;
      RECT  142.34 114.33 142.85 114.09 ;
      RECT  139.94 115.43 142.34 115.19 ;
      RECT  142.34 115.19 142.54 115.12 ;
      RECT  142.13 114.4 142.34 114.33 ;
      RECT  142.85 115.43 143.06 115.19 ;
      POLYGON  141.41 114.95 141.41 114.57 141.96 114.57 141.96 114.64 142.34 114.64 142.34 114.88 141.96 114.88 141.96 114.95 141.41 114.95 ;
      RECT  142.85 114.95 143.06 114.57 ;
      RECT  139.73 116.22 139.94 115.67 ;
      RECT  139.94 116.22 140.87 115.67 ;
      RECT  140.87 114.95 141.41 114.57 ;
      RECT  142.85 114.33 143.06 114.09 ;
      RECT  141.41 116.22 143.06 115.67 ;
      RECT  139.73 115.43 139.94 115.19 ;
      RECT  142.34 114.4 142.54 114.33 ;
      POLYGON  142.71 114.95 142.71 114.88 142.34 114.88 142.34 114.64 142.71 114.64 142.71 114.57 142.85 114.57 142.85 114.95 142.71 114.95 ;
      RECT  139.73 114.33 139.94 114.09 ;
      RECT  139.94 114.33 142.34 114.09 ;
      RECT  142.34 115.43 142.85 115.19 ;
      RECT  140.87 116.22 141.41 115.67 ;
      RECT  139.73 116.94 140.87 117.32 ;
      RECT  142.13 116.7 142.34 116.77 ;
      RECT  142.34 117.56 142.85 117.8 ;
      RECT  139.94 116.46 142.34 116.7 ;
      RECT  142.34 116.7 142.54 116.77 ;
      RECT  142.13 117.49 142.34 117.56 ;
      RECT  142.85 116.46 143.06 116.7 ;
      POLYGON  141.41 116.94 141.41 117.32 141.96 117.32 141.96 117.25 142.34 117.25 142.34 117.01 141.96 117.01 141.96 116.94 141.41 116.94 ;
      RECT  142.85 116.94 143.06 117.32 ;
      RECT  139.73 115.67 139.94 116.22 ;
      RECT  139.94 115.67 140.87 116.22 ;
      RECT  140.87 116.94 141.41 117.32 ;
      RECT  142.85 117.56 143.06 117.8 ;
      RECT  141.41 115.67 143.06 116.22 ;
      RECT  139.73 116.46 139.94 116.7 ;
      RECT  142.34 117.49 142.54 117.56 ;
      POLYGON  142.71 116.94 142.71 117.01 142.34 117.01 142.34 117.25 142.71 117.25 142.71 117.32 142.85 117.32 142.85 116.94 142.71 116.94 ;
      RECT  139.73 117.56 139.94 117.8 ;
      RECT  139.94 117.56 142.34 117.8 ;
      RECT  142.34 116.46 142.85 116.7 ;
      RECT  140.87 115.67 141.41 116.22 ;
      RECT  139.73 118.9 140.87 118.52 ;
      RECT  142.13 119.14 142.34 119.07 ;
      RECT  142.34 118.28 142.85 118.04 ;
      RECT  139.94 119.38 142.34 119.14 ;
      RECT  142.34 119.14 142.54 119.07 ;
      RECT  142.13 118.35 142.34 118.28 ;
      RECT  142.85 119.38 143.06 119.14 ;
      POLYGON  141.41 118.9 141.41 118.52 141.96 118.52 141.96 118.59 142.34 118.59 142.34 118.83 141.96 118.83 141.96 118.9 141.41 118.9 ;
      RECT  142.85 118.9 143.06 118.52 ;
      RECT  139.73 120.17 139.94 119.62 ;
      RECT  139.94 120.17 140.87 119.62 ;
      RECT  140.87 118.9 141.41 118.52 ;
      RECT  142.85 118.28 143.06 118.04 ;
      RECT  141.41 120.17 143.06 119.62 ;
      RECT  139.73 119.38 139.94 119.14 ;
      RECT  142.34 118.35 142.54 118.28 ;
      POLYGON  142.71 118.9 142.71 118.83 142.34 118.83 142.34 118.59 142.71 118.59 142.71 118.52 142.85 118.52 142.85 118.9 142.71 118.9 ;
      RECT  139.73 118.28 139.94 118.04 ;
      RECT  139.94 118.28 142.34 118.04 ;
      RECT  142.34 119.38 142.85 119.14 ;
      RECT  140.87 120.17 141.41 119.62 ;
      RECT  139.73 120.89 140.87 121.27 ;
      RECT  142.13 120.65 142.34 120.72 ;
      RECT  142.34 121.51 142.85 121.75 ;
      RECT  139.94 120.41 142.34 120.65 ;
      RECT  142.34 120.65 142.54 120.72 ;
      RECT  142.13 121.44 142.34 121.51 ;
      RECT  142.85 120.41 143.06 120.65 ;
      POLYGON  141.41 120.89 141.41 121.27 141.96 121.27 141.96 121.2 142.34 121.2 142.34 120.96 141.96 120.96 141.96 120.89 141.41 120.89 ;
      RECT  142.85 120.89 143.06 121.27 ;
      RECT  139.73 119.62 139.94 120.17 ;
      RECT  139.94 119.62 140.87 120.17 ;
      RECT  140.87 120.89 141.41 121.27 ;
      RECT  142.85 121.51 143.06 121.75 ;
      RECT  141.41 119.62 143.06 120.17 ;
      RECT  139.73 120.41 139.94 120.65 ;
      RECT  142.34 121.44 142.54 121.51 ;
      POLYGON  142.71 120.89 142.71 120.96 142.34 120.96 142.34 121.2 142.71 121.2 142.71 121.27 142.85 121.27 142.85 120.89 142.71 120.89 ;
      RECT  139.73 121.51 139.94 121.75 ;
      RECT  139.94 121.51 142.34 121.75 ;
      RECT  142.34 120.41 142.85 120.65 ;
      RECT  140.87 119.62 141.41 120.17 ;
      RECT  139.73 122.85 140.87 122.47 ;
      RECT  142.13 123.09 142.34 123.02 ;
      RECT  142.34 122.23 142.85 121.99 ;
      RECT  139.94 123.33 142.34 123.09 ;
      RECT  142.34 123.09 142.54 123.02 ;
      RECT  142.13 122.3 142.34 122.23 ;
      RECT  142.85 123.33 143.06 123.09 ;
      POLYGON  141.41 122.85 141.41 122.47 141.96 122.47 141.96 122.54 142.34 122.54 142.34 122.78 141.96 122.78 141.96 122.85 141.41 122.85 ;
      RECT  142.85 122.85 143.06 122.47 ;
      RECT  139.73 124.12 139.94 123.57 ;
      RECT  139.94 124.12 140.87 123.57 ;
      RECT  140.87 122.85 141.41 122.47 ;
      RECT  142.85 122.23 143.06 121.99 ;
      RECT  141.41 124.12 143.06 123.57 ;
      RECT  139.73 123.33 139.94 123.09 ;
      RECT  142.34 122.3 142.54 122.23 ;
      POLYGON  142.71 122.85 142.71 122.78 142.34 122.78 142.34 122.54 142.71 122.54 142.71 122.47 142.85 122.47 142.85 122.85 142.71 122.85 ;
      RECT  139.73 122.23 139.94 121.99 ;
      RECT  139.94 122.23 142.34 121.99 ;
      RECT  142.34 123.33 142.85 123.09 ;
      RECT  140.87 124.12 141.41 123.57 ;
      RECT  146.39 93.24 145.25 93.62 ;
      RECT  143.99 93.0 143.78 93.07 ;
      RECT  143.78 93.86 143.27 94.1 ;
      RECT  146.18 92.76 143.78 93.0 ;
      RECT  143.78 93.0 143.58 93.07 ;
      RECT  143.99 93.79 143.78 93.86 ;
      RECT  143.27 92.76 143.06 93.0 ;
      POLYGON  144.71 93.24 144.71 93.62 144.16 93.62 144.16 93.55 143.78 93.55 143.78 93.31 144.16 93.31 144.16 93.24 144.71 93.24 ;
      RECT  143.27 93.24 143.06 93.62 ;
      RECT  146.39 91.97 146.18 92.52 ;
      RECT  146.18 91.97 145.25 92.52 ;
      RECT  145.25 93.24 144.71 93.62 ;
      RECT  143.27 93.86 143.06 94.1 ;
      RECT  144.71 91.97 143.06 92.52 ;
      RECT  146.39 92.76 146.18 93.0 ;
      RECT  143.78 93.79 143.58 93.86 ;
      POLYGON  143.41 93.24 143.41 93.31 143.78 93.31 143.78 93.55 143.41 93.55 143.41 93.62 143.27 93.62 143.27 93.24 143.41 93.24 ;
      RECT  146.39 93.86 146.18 94.1 ;
      RECT  146.18 93.86 143.78 94.1 ;
      RECT  143.78 92.76 143.27 93.0 ;
      RECT  145.25 91.97 144.71 92.52 ;
      RECT  146.39 95.2 145.25 94.82 ;
      RECT  143.99 95.44 143.78 95.37 ;
      RECT  143.78 94.58 143.27 94.34 ;
      RECT  146.18 95.68 143.78 95.44 ;
      RECT  143.78 95.44 143.58 95.37 ;
      RECT  143.99 94.65 143.78 94.58 ;
      RECT  143.27 95.68 143.06 95.44 ;
      POLYGON  144.71 95.2 144.71 94.82 144.16 94.82 144.16 94.89 143.78 94.89 143.78 95.13 144.16 95.13 144.16 95.2 144.71 95.2 ;
      RECT  143.27 95.2 143.06 94.82 ;
      RECT  146.39 96.47 146.18 95.92 ;
      RECT  146.18 96.47 145.25 95.92 ;
      RECT  145.25 95.2 144.71 94.82 ;
      RECT  143.27 94.58 143.06 94.34 ;
      RECT  144.71 96.47 143.06 95.92 ;
      RECT  146.39 95.68 146.18 95.44 ;
      RECT  143.78 94.65 143.58 94.58 ;
      POLYGON  143.41 95.2 143.41 95.13 143.78 95.13 143.78 94.89 143.41 94.89 143.41 94.82 143.27 94.82 143.27 95.2 143.41 95.2 ;
      RECT  146.39 94.58 146.18 94.34 ;
      RECT  146.18 94.58 143.78 94.34 ;
      RECT  143.78 95.68 143.27 95.44 ;
      RECT  145.25 96.47 144.71 95.92 ;
      RECT  146.39 97.19 145.25 97.57 ;
      RECT  143.99 96.95 143.78 97.02 ;
      RECT  143.78 97.81 143.27 98.05 ;
      RECT  146.18 96.71 143.78 96.95 ;
      RECT  143.78 96.95 143.58 97.02 ;
      RECT  143.99 97.74 143.78 97.81 ;
      RECT  143.27 96.71 143.06 96.95 ;
      POLYGON  144.71 97.19 144.71 97.57 144.16 97.57 144.16 97.5 143.78 97.5 143.78 97.26 144.16 97.26 144.16 97.19 144.71 97.19 ;
      RECT  143.27 97.19 143.06 97.57 ;
      RECT  146.39 95.92 146.18 96.47 ;
      RECT  146.18 95.92 145.25 96.47 ;
      RECT  145.25 97.19 144.71 97.57 ;
      RECT  143.27 97.81 143.06 98.05 ;
      RECT  144.71 95.92 143.06 96.47 ;
      RECT  146.39 96.71 146.18 96.95 ;
      RECT  143.78 97.74 143.58 97.81 ;
      POLYGON  143.41 97.19 143.41 97.26 143.78 97.26 143.78 97.5 143.41 97.5 143.41 97.57 143.27 97.57 143.27 97.19 143.41 97.19 ;
      RECT  146.39 97.81 146.18 98.05 ;
      RECT  146.18 97.81 143.78 98.05 ;
      RECT  143.78 96.71 143.27 96.95 ;
      RECT  145.25 95.92 144.71 96.47 ;
      RECT  146.39 99.15 145.25 98.77 ;
      RECT  143.99 99.39 143.78 99.32 ;
      RECT  143.78 98.53 143.27 98.29 ;
      RECT  146.18 99.63 143.78 99.39 ;
      RECT  143.78 99.39 143.58 99.32 ;
      RECT  143.99 98.6 143.78 98.53 ;
      RECT  143.27 99.63 143.06 99.39 ;
      POLYGON  144.71 99.15 144.71 98.77 144.16 98.77 144.16 98.84 143.78 98.84 143.78 99.08 144.16 99.08 144.16 99.15 144.71 99.15 ;
      RECT  143.27 99.15 143.06 98.77 ;
      RECT  146.39 100.42 146.18 99.87 ;
      RECT  146.18 100.42 145.25 99.87 ;
      RECT  145.25 99.15 144.71 98.77 ;
      RECT  143.27 98.53 143.06 98.29 ;
      RECT  144.71 100.42 143.06 99.87 ;
      RECT  146.39 99.63 146.18 99.39 ;
      RECT  143.78 98.6 143.58 98.53 ;
      POLYGON  143.41 99.15 143.41 99.08 143.78 99.08 143.78 98.84 143.41 98.84 143.41 98.77 143.27 98.77 143.27 99.15 143.41 99.15 ;
      RECT  146.39 98.53 146.18 98.29 ;
      RECT  146.18 98.53 143.78 98.29 ;
      RECT  143.78 99.63 143.27 99.39 ;
      RECT  145.25 100.42 144.71 99.87 ;
      RECT  146.39 101.14 145.25 101.52 ;
      RECT  143.99 100.9 143.78 100.97 ;
      RECT  143.78 101.76 143.27 102.0 ;
      RECT  146.18 100.66 143.78 100.9 ;
      RECT  143.78 100.9 143.58 100.97 ;
      RECT  143.99 101.69 143.78 101.76 ;
      RECT  143.27 100.66 143.06 100.9 ;
      POLYGON  144.71 101.14 144.71 101.52 144.16 101.52 144.16 101.45 143.78 101.45 143.78 101.21 144.16 101.21 144.16 101.14 144.71 101.14 ;
      RECT  143.27 101.14 143.06 101.52 ;
      RECT  146.39 99.87 146.18 100.42 ;
      RECT  146.18 99.87 145.25 100.42 ;
      RECT  145.25 101.14 144.71 101.52 ;
      RECT  143.27 101.76 143.06 102.0 ;
      RECT  144.71 99.87 143.06 100.42 ;
      RECT  146.39 100.66 146.18 100.9 ;
      RECT  143.78 101.69 143.58 101.76 ;
      POLYGON  143.41 101.14 143.41 101.21 143.78 101.21 143.78 101.45 143.41 101.45 143.41 101.52 143.27 101.52 143.27 101.14 143.41 101.14 ;
      RECT  146.39 101.76 146.18 102.0 ;
      RECT  146.18 101.76 143.78 102.0 ;
      RECT  143.78 100.66 143.27 100.9 ;
      RECT  145.25 99.87 144.71 100.42 ;
      RECT  146.39 103.1 145.25 102.72 ;
      RECT  143.99 103.34 143.78 103.27 ;
      RECT  143.78 102.48 143.27 102.24 ;
      RECT  146.18 103.58 143.78 103.34 ;
      RECT  143.78 103.34 143.58 103.27 ;
      RECT  143.99 102.55 143.78 102.48 ;
      RECT  143.27 103.58 143.06 103.34 ;
      POLYGON  144.71 103.1 144.71 102.72 144.16 102.72 144.16 102.79 143.78 102.79 143.78 103.03 144.16 103.03 144.16 103.1 144.71 103.1 ;
      RECT  143.27 103.1 143.06 102.72 ;
      RECT  146.39 104.37 146.18 103.82 ;
      RECT  146.18 104.37 145.25 103.82 ;
      RECT  145.25 103.1 144.71 102.72 ;
      RECT  143.27 102.48 143.06 102.24 ;
      RECT  144.71 104.37 143.06 103.82 ;
      RECT  146.39 103.58 146.18 103.34 ;
      RECT  143.78 102.55 143.58 102.48 ;
      POLYGON  143.41 103.1 143.41 103.03 143.78 103.03 143.78 102.79 143.41 102.79 143.41 102.72 143.27 102.72 143.27 103.1 143.41 103.1 ;
      RECT  146.39 102.48 146.18 102.24 ;
      RECT  146.18 102.48 143.78 102.24 ;
      RECT  143.78 103.58 143.27 103.34 ;
      RECT  145.25 104.37 144.71 103.82 ;
      RECT  146.39 105.09 145.25 105.47 ;
      RECT  143.99 104.85 143.78 104.92 ;
      RECT  143.78 105.71 143.27 105.95 ;
      RECT  146.18 104.61 143.78 104.85 ;
      RECT  143.78 104.85 143.58 104.92 ;
      RECT  143.99 105.64 143.78 105.71 ;
      RECT  143.27 104.61 143.06 104.85 ;
      POLYGON  144.71 105.09 144.71 105.47 144.16 105.47 144.16 105.4 143.78 105.4 143.78 105.16 144.16 105.16 144.16 105.09 144.71 105.09 ;
      RECT  143.27 105.09 143.06 105.47 ;
      RECT  146.39 103.82 146.18 104.37 ;
      RECT  146.18 103.82 145.25 104.37 ;
      RECT  145.25 105.09 144.71 105.47 ;
      RECT  143.27 105.71 143.06 105.95 ;
      RECT  144.71 103.82 143.06 104.37 ;
      RECT  146.39 104.61 146.18 104.85 ;
      RECT  143.78 105.64 143.58 105.71 ;
      POLYGON  143.41 105.09 143.41 105.16 143.78 105.16 143.78 105.4 143.41 105.4 143.41 105.47 143.27 105.47 143.27 105.09 143.41 105.09 ;
      RECT  146.39 105.71 146.18 105.95 ;
      RECT  146.18 105.71 143.78 105.95 ;
      RECT  143.78 104.61 143.27 104.85 ;
      RECT  145.25 103.82 144.71 104.37 ;
      RECT  146.39 107.05 145.25 106.67 ;
      RECT  143.99 107.29 143.78 107.22 ;
      RECT  143.78 106.43 143.27 106.19 ;
      RECT  146.18 107.53 143.78 107.29 ;
      RECT  143.78 107.29 143.58 107.22 ;
      RECT  143.99 106.5 143.78 106.43 ;
      RECT  143.27 107.53 143.06 107.29 ;
      POLYGON  144.71 107.05 144.71 106.67 144.16 106.67 144.16 106.74 143.78 106.74 143.78 106.98 144.16 106.98 144.16 107.05 144.71 107.05 ;
      RECT  143.27 107.05 143.06 106.67 ;
      RECT  146.39 108.32 146.18 107.77 ;
      RECT  146.18 108.32 145.25 107.77 ;
      RECT  145.25 107.05 144.71 106.67 ;
      RECT  143.27 106.43 143.06 106.19 ;
      RECT  144.71 108.32 143.06 107.77 ;
      RECT  146.39 107.53 146.18 107.29 ;
      RECT  143.78 106.5 143.58 106.43 ;
      POLYGON  143.41 107.05 143.41 106.98 143.78 106.98 143.78 106.74 143.41 106.74 143.41 106.67 143.27 106.67 143.27 107.05 143.41 107.05 ;
      RECT  146.39 106.43 146.18 106.19 ;
      RECT  146.18 106.43 143.78 106.19 ;
      RECT  143.78 107.53 143.27 107.29 ;
      RECT  145.25 108.32 144.71 107.77 ;
      RECT  146.39 109.04 145.25 109.42 ;
      RECT  143.99 108.8 143.78 108.87 ;
      RECT  143.78 109.66 143.27 109.9 ;
      RECT  146.18 108.56 143.78 108.8 ;
      RECT  143.78 108.8 143.58 108.87 ;
      RECT  143.99 109.59 143.78 109.66 ;
      RECT  143.27 108.56 143.06 108.8 ;
      POLYGON  144.71 109.04 144.71 109.42 144.16 109.42 144.16 109.35 143.78 109.35 143.78 109.11 144.16 109.11 144.16 109.04 144.71 109.04 ;
      RECT  143.27 109.04 143.06 109.42 ;
      RECT  146.39 107.77 146.18 108.32 ;
      RECT  146.18 107.77 145.25 108.32 ;
      RECT  145.25 109.04 144.71 109.42 ;
      RECT  143.27 109.66 143.06 109.9 ;
      RECT  144.71 107.77 143.06 108.32 ;
      RECT  146.39 108.56 146.18 108.8 ;
      RECT  143.78 109.59 143.58 109.66 ;
      POLYGON  143.41 109.04 143.41 109.11 143.78 109.11 143.78 109.35 143.41 109.35 143.41 109.42 143.27 109.42 143.27 109.04 143.41 109.04 ;
      RECT  146.39 109.66 146.18 109.9 ;
      RECT  146.18 109.66 143.78 109.9 ;
      RECT  143.78 108.56 143.27 108.8 ;
      RECT  145.25 107.77 144.71 108.32 ;
      RECT  146.39 111.0 145.25 110.62 ;
      RECT  143.99 111.24 143.78 111.17 ;
      RECT  143.78 110.38 143.27 110.14 ;
      RECT  146.18 111.48 143.78 111.24 ;
      RECT  143.78 111.24 143.58 111.17 ;
      RECT  143.99 110.45 143.78 110.38 ;
      RECT  143.27 111.48 143.06 111.24 ;
      POLYGON  144.71 111.0 144.71 110.62 144.16 110.62 144.16 110.69 143.78 110.69 143.78 110.93 144.16 110.93 144.16 111.0 144.71 111.0 ;
      RECT  143.27 111.0 143.06 110.62 ;
      RECT  146.39 112.27 146.18 111.72 ;
      RECT  146.18 112.27 145.25 111.72 ;
      RECT  145.25 111.0 144.71 110.62 ;
      RECT  143.27 110.38 143.06 110.14 ;
      RECT  144.71 112.27 143.06 111.72 ;
      RECT  146.39 111.48 146.18 111.24 ;
      RECT  143.78 110.45 143.58 110.38 ;
      POLYGON  143.41 111.0 143.41 110.93 143.78 110.93 143.78 110.69 143.41 110.69 143.41 110.62 143.27 110.62 143.27 111.0 143.41 111.0 ;
      RECT  146.39 110.38 146.18 110.14 ;
      RECT  146.18 110.38 143.78 110.14 ;
      RECT  143.78 111.48 143.27 111.24 ;
      RECT  145.25 112.27 144.71 111.72 ;
      RECT  146.39 112.99 145.25 113.37 ;
      RECT  143.99 112.75 143.78 112.82 ;
      RECT  143.78 113.61 143.27 113.85 ;
      RECT  146.18 112.51 143.78 112.75 ;
      RECT  143.78 112.75 143.58 112.82 ;
      RECT  143.99 113.54 143.78 113.61 ;
      RECT  143.27 112.51 143.06 112.75 ;
      POLYGON  144.71 112.99 144.71 113.37 144.16 113.37 144.16 113.3 143.78 113.3 143.78 113.06 144.16 113.06 144.16 112.99 144.71 112.99 ;
      RECT  143.27 112.99 143.06 113.37 ;
      RECT  146.39 111.72 146.18 112.27 ;
      RECT  146.18 111.72 145.25 112.27 ;
      RECT  145.25 112.99 144.71 113.37 ;
      RECT  143.27 113.61 143.06 113.85 ;
      RECT  144.71 111.72 143.06 112.27 ;
      RECT  146.39 112.51 146.18 112.75 ;
      RECT  143.78 113.54 143.58 113.61 ;
      POLYGON  143.41 112.99 143.41 113.06 143.78 113.06 143.78 113.3 143.41 113.3 143.41 113.37 143.27 113.37 143.27 112.99 143.41 112.99 ;
      RECT  146.39 113.61 146.18 113.85 ;
      RECT  146.18 113.61 143.78 113.85 ;
      RECT  143.78 112.51 143.27 112.75 ;
      RECT  145.25 111.72 144.71 112.27 ;
      RECT  146.39 114.95 145.25 114.57 ;
      RECT  143.99 115.19 143.78 115.12 ;
      RECT  143.78 114.33 143.27 114.09 ;
      RECT  146.18 115.43 143.78 115.19 ;
      RECT  143.78 115.19 143.58 115.12 ;
      RECT  143.99 114.4 143.78 114.33 ;
      RECT  143.27 115.43 143.06 115.19 ;
      POLYGON  144.71 114.95 144.71 114.57 144.16 114.57 144.16 114.64 143.78 114.64 143.78 114.88 144.16 114.88 144.16 114.95 144.71 114.95 ;
      RECT  143.27 114.95 143.06 114.57 ;
      RECT  146.39 116.22 146.18 115.67 ;
      RECT  146.18 116.22 145.25 115.67 ;
      RECT  145.25 114.95 144.71 114.57 ;
      RECT  143.27 114.33 143.06 114.09 ;
      RECT  144.71 116.22 143.06 115.67 ;
      RECT  146.39 115.43 146.18 115.19 ;
      RECT  143.78 114.4 143.58 114.33 ;
      POLYGON  143.41 114.95 143.41 114.88 143.78 114.88 143.78 114.64 143.41 114.64 143.41 114.57 143.27 114.57 143.27 114.95 143.41 114.95 ;
      RECT  146.39 114.33 146.18 114.09 ;
      RECT  146.18 114.33 143.78 114.09 ;
      RECT  143.78 115.43 143.27 115.19 ;
      RECT  145.25 116.22 144.71 115.67 ;
      RECT  146.39 116.94 145.25 117.32 ;
      RECT  143.99 116.7 143.78 116.77 ;
      RECT  143.78 117.56 143.27 117.8 ;
      RECT  146.18 116.46 143.78 116.7 ;
      RECT  143.78 116.7 143.58 116.77 ;
      RECT  143.99 117.49 143.78 117.56 ;
      RECT  143.27 116.46 143.06 116.7 ;
      POLYGON  144.71 116.94 144.71 117.32 144.16 117.32 144.16 117.25 143.78 117.25 143.78 117.01 144.16 117.01 144.16 116.94 144.71 116.94 ;
      RECT  143.27 116.94 143.06 117.32 ;
      RECT  146.39 115.67 146.18 116.22 ;
      RECT  146.18 115.67 145.25 116.22 ;
      RECT  145.25 116.94 144.71 117.32 ;
      RECT  143.27 117.56 143.06 117.8 ;
      RECT  144.71 115.67 143.06 116.22 ;
      RECT  146.39 116.46 146.18 116.7 ;
      RECT  143.78 117.49 143.58 117.56 ;
      POLYGON  143.41 116.94 143.41 117.01 143.78 117.01 143.78 117.25 143.41 117.25 143.41 117.32 143.27 117.32 143.27 116.94 143.41 116.94 ;
      RECT  146.39 117.56 146.18 117.8 ;
      RECT  146.18 117.56 143.78 117.8 ;
      RECT  143.78 116.46 143.27 116.7 ;
      RECT  145.25 115.67 144.71 116.22 ;
      RECT  146.39 118.9 145.25 118.52 ;
      RECT  143.99 119.14 143.78 119.07 ;
      RECT  143.78 118.28 143.27 118.04 ;
      RECT  146.18 119.38 143.78 119.14 ;
      RECT  143.78 119.14 143.58 119.07 ;
      RECT  143.99 118.35 143.78 118.28 ;
      RECT  143.27 119.38 143.06 119.14 ;
      POLYGON  144.71 118.9 144.71 118.52 144.16 118.52 144.16 118.59 143.78 118.59 143.78 118.83 144.16 118.83 144.16 118.9 144.71 118.9 ;
      RECT  143.27 118.9 143.06 118.52 ;
      RECT  146.39 120.17 146.18 119.62 ;
      RECT  146.18 120.17 145.25 119.62 ;
      RECT  145.25 118.9 144.71 118.52 ;
      RECT  143.27 118.28 143.06 118.04 ;
      RECT  144.71 120.17 143.06 119.62 ;
      RECT  146.39 119.38 146.18 119.14 ;
      RECT  143.78 118.35 143.58 118.28 ;
      POLYGON  143.41 118.9 143.41 118.83 143.78 118.83 143.78 118.59 143.41 118.59 143.41 118.52 143.27 118.52 143.27 118.9 143.41 118.9 ;
      RECT  146.39 118.28 146.18 118.04 ;
      RECT  146.18 118.28 143.78 118.04 ;
      RECT  143.78 119.38 143.27 119.14 ;
      RECT  145.25 120.17 144.71 119.62 ;
      RECT  146.39 120.89 145.25 121.27 ;
      RECT  143.99 120.65 143.78 120.72 ;
      RECT  143.78 121.51 143.27 121.75 ;
      RECT  146.18 120.41 143.78 120.65 ;
      RECT  143.78 120.65 143.58 120.72 ;
      RECT  143.99 121.44 143.78 121.51 ;
      RECT  143.27 120.41 143.06 120.65 ;
      POLYGON  144.71 120.89 144.71 121.27 144.16 121.27 144.16 121.2 143.78 121.2 143.78 120.96 144.16 120.96 144.16 120.89 144.71 120.89 ;
      RECT  143.27 120.89 143.06 121.27 ;
      RECT  146.39 119.62 146.18 120.17 ;
      RECT  146.18 119.62 145.25 120.17 ;
      RECT  145.25 120.89 144.71 121.27 ;
      RECT  143.27 121.51 143.06 121.75 ;
      RECT  144.71 119.62 143.06 120.17 ;
      RECT  146.39 120.41 146.18 120.65 ;
      RECT  143.78 121.44 143.58 121.51 ;
      POLYGON  143.41 120.89 143.41 120.96 143.78 120.96 143.78 121.2 143.41 121.2 143.41 121.27 143.27 121.27 143.27 120.89 143.41 120.89 ;
      RECT  146.39 121.51 146.18 121.75 ;
      RECT  146.18 121.51 143.78 121.75 ;
      RECT  143.78 120.41 143.27 120.65 ;
      RECT  145.25 119.62 144.71 120.17 ;
      RECT  146.39 122.85 145.25 122.47 ;
      RECT  143.99 123.09 143.78 123.02 ;
      RECT  143.78 122.23 143.27 121.99 ;
      RECT  146.18 123.33 143.78 123.09 ;
      RECT  143.78 123.09 143.58 123.02 ;
      RECT  143.99 122.3 143.78 122.23 ;
      RECT  143.27 123.33 143.06 123.09 ;
      POLYGON  144.71 122.85 144.71 122.47 144.16 122.47 144.16 122.54 143.78 122.54 143.78 122.78 144.16 122.78 144.16 122.85 144.71 122.85 ;
      RECT  143.27 122.85 143.06 122.47 ;
      RECT  146.39 124.12 146.18 123.57 ;
      RECT  146.18 124.12 145.25 123.57 ;
      RECT  145.25 122.85 144.71 122.47 ;
      RECT  143.27 122.23 143.06 121.99 ;
      RECT  144.71 124.12 143.06 123.57 ;
      RECT  146.39 123.33 146.18 123.09 ;
      RECT  143.78 122.3 143.58 122.23 ;
      POLYGON  143.41 122.85 143.41 122.78 143.78 122.78 143.78 122.54 143.41 122.54 143.41 122.47 143.27 122.47 143.27 122.85 143.41 122.85 ;
      RECT  146.39 122.23 146.18 121.99 ;
      RECT  146.18 122.23 143.78 121.99 ;
      RECT  143.78 123.33 143.27 123.09 ;
      RECT  145.25 124.12 144.71 123.57 ;
      RECT  96.26 93.86 146.18 94.1 ;
      RECT  96.26 92.76 146.18 93.0 ;
      RECT  96.26 94.34 146.18 94.58 ;
      RECT  96.26 95.44 146.18 95.68 ;
      RECT  96.26 97.81 146.18 98.05 ;
      RECT  96.26 96.71 146.18 96.95 ;
      RECT  96.26 98.29 146.18 98.53 ;
      RECT  96.26 99.39 146.18 99.63 ;
      RECT  96.26 101.76 146.18 102.0 ;
      RECT  96.26 100.66 146.18 100.9 ;
      RECT  96.26 102.24 146.18 102.48 ;
      RECT  96.26 103.34 146.18 103.58 ;
      RECT  96.26 105.71 146.18 105.95 ;
      RECT  96.26 104.61 146.18 104.85 ;
      RECT  96.26 106.19 146.18 106.43 ;
      RECT  96.26 107.29 146.18 107.53 ;
      RECT  96.26 109.66 146.18 109.9 ;
      RECT  96.26 108.56 146.18 108.8 ;
      RECT  96.26 110.14 146.18 110.38 ;
      RECT  96.26 111.24 146.18 111.48 ;
      RECT  96.26 113.61 146.18 113.85 ;
      RECT  96.26 112.51 146.18 112.75 ;
      RECT  96.26 114.09 146.18 114.33 ;
      RECT  96.26 115.19 146.18 115.43 ;
      RECT  96.26 117.56 146.18 117.8 ;
      RECT  96.26 116.46 146.18 116.7 ;
      RECT  96.26 118.04 146.18 118.28 ;
      RECT  96.26 119.14 146.18 119.38 ;
      RECT  96.26 121.51 146.18 121.75 ;
      RECT  96.26 120.41 146.18 120.65 ;
      RECT  96.26 121.99 146.18 122.23 ;
      RECT  96.26 123.09 146.18 123.33 ;
      RECT  144.71 118.52 145.25 118.9 ;
      RECT  113.51 115.67 114.05 116.22 ;
      RECT  122.15 95.92 122.69 96.47 ;
      RECT  97.19 95.92 97.73 96.47 ;
      RECT  119.75 118.52 120.29 118.9 ;
      RECT  103.43 115.67 103.97 116.22 ;
      RECT  140.87 99.87 141.41 100.42 ;
      RECT  122.15 122.47 122.69 122.85 ;
      RECT  113.51 123.57 114.05 124.12 ;
      RECT  109.67 93.24 110.21 93.62 ;
      RECT  132.23 103.82 132.77 104.37 ;
      RECT  122.15 115.67 122.69 116.22 ;
      RECT  132.23 109.04 132.77 109.42 ;
      RECT  109.67 110.62 110.21 111.0 ;
      RECT  109.67 118.52 110.21 118.9 ;
      RECT  138.47 122.47 139.01 122.85 ;
      RECT  101.03 97.19 101.57 97.57 ;
      RECT  101.03 106.67 101.57 107.05 ;
      RECT  119.75 119.62 120.29 120.17 ;
      RECT  107.27 99.87 107.81 100.42 ;
      RECT  113.51 98.77 114.05 99.15 ;
      RECT  97.19 110.62 97.73 111.0 ;
      RECT  144.71 123.57 145.25 124.12 ;
      RECT  113.51 120.89 114.05 121.27 ;
      RECT  109.67 91.97 110.21 92.52 ;
      RECT  113.51 94.82 114.05 95.2 ;
      RECT  125.99 107.77 126.53 108.32 ;
      RECT  122.15 102.72 122.69 103.1 ;
      RECT  115.91 98.77 116.45 99.15 ;
      RECT  119.75 123.57 120.29 124.12 ;
      RECT  122.15 93.24 122.69 93.62 ;
      RECT  103.43 116.94 103.97 117.32 ;
      RECT  97.19 123.57 97.73 124.12 ;
      RECT  97.19 109.04 97.73 109.42 ;
      RECT  144.71 114.57 145.25 114.95 ;
      RECT  109.67 97.19 110.21 97.57 ;
      RECT  101.03 119.62 101.57 120.17 ;
      RECT  138.47 105.09 139.01 105.47 ;
      RECT  140.87 105.09 141.41 105.47 ;
      RECT  115.91 116.94 116.45 117.32 ;
      RECT  134.63 111.72 135.17 112.27 ;
      RECT  128.39 111.72 128.93 112.27 ;
      RECT  115.91 105.09 116.45 105.47 ;
      RECT  134.63 97.19 135.17 97.57 ;
      RECT  134.63 94.82 135.17 95.2 ;
      RECT  107.27 118.52 107.81 118.9 ;
      RECT  140.87 115.67 141.41 116.22 ;
      RECT  138.47 116.94 139.01 117.32 ;
      RECT  115.91 109.04 116.45 109.42 ;
      RECT  138.47 99.87 139.01 100.42 ;
      RECT  125.99 111.72 126.53 112.27 ;
      RECT  122.15 114.57 122.69 114.95 ;
      RECT  125.99 115.67 126.53 116.22 ;
      RECT  101.03 107.77 101.57 108.32 ;
      RECT  119.75 101.14 120.29 101.52 ;
      RECT  138.47 115.67 139.01 116.22 ;
      RECT  134.63 119.62 135.17 120.17 ;
      RECT  122.15 106.67 122.69 107.05 ;
      RECT  109.67 98.77 110.21 99.15 ;
      RECT  144.71 119.62 145.25 120.17 ;
      RECT  119.75 95.92 120.29 96.47 ;
      RECT  125.99 98.77 126.53 99.15 ;
      RECT  115.91 91.97 116.45 92.52 ;
      RECT  113.51 110.62 114.05 111.0 ;
      RECT  144.71 111.72 145.25 112.27 ;
      RECT  107.27 119.62 107.81 120.17 ;
      RECT  103.43 120.89 103.97 121.27 ;
      RECT  134.63 98.77 135.17 99.15 ;
      RECT  140.87 118.52 141.41 118.9 ;
      RECT  119.75 91.97 120.29 92.52 ;
      RECT  113.51 111.72 114.05 112.27 ;
      RECT  144.71 110.62 145.25 111.0 ;
      RECT  101.03 102.72 101.57 103.1 ;
      RECT  138.47 110.62 139.01 111.0 ;
      RECT  97.19 91.97 97.73 92.52 ;
      RECT  125.99 93.24 126.53 93.62 ;
      RECT  101.03 101.14 101.57 101.52 ;
      RECT  115.91 97.19 116.45 97.57 ;
      RECT  109.67 105.09 110.21 105.47 ;
      RECT  128.39 118.52 128.93 118.9 ;
      RECT  122.15 98.77 122.69 99.15 ;
      RECT  113.51 114.57 114.05 114.95 ;
      RECT  125.99 105.09 126.53 105.47 ;
      RECT  140.87 123.57 141.41 124.12 ;
      RECT  138.47 101.14 139.01 101.52 ;
      RECT  113.51 105.09 114.05 105.47 ;
      RECT  140.87 94.82 141.41 95.2 ;
      RECT  132.23 111.72 132.77 112.27 ;
      RECT  103.43 122.47 103.97 122.85 ;
      RECT  113.51 95.92 114.05 96.47 ;
      RECT  109.67 111.72 110.21 112.27 ;
      RECT  132.23 107.77 132.77 108.32 ;
      RECT  101.03 118.52 101.57 118.9 ;
      RECT  113.51 109.04 114.05 109.42 ;
      RECT  119.75 99.87 120.29 100.42 ;
      RECT  134.63 112.99 135.17 113.37 ;
      RECT  134.63 115.67 135.17 116.22 ;
      RECT  140.87 116.94 141.41 117.32 ;
      RECT  109.67 102.72 110.21 103.1 ;
      RECT  103.43 102.72 103.97 103.1 ;
      RECT  113.51 97.19 114.05 97.57 ;
      RECT  128.39 114.57 128.93 114.95 ;
      RECT  107.27 107.77 107.81 108.32 ;
      RECT  97.19 94.82 97.73 95.2 ;
      RECT  115.91 118.52 116.45 118.9 ;
      RECT  138.47 120.89 139.01 121.27 ;
      RECT  103.43 110.62 103.97 111.0 ;
      RECT  109.67 99.87 110.21 100.42 ;
      RECT  97.19 102.72 97.73 103.1 ;
      RECT  115.91 101.14 116.45 101.52 ;
      RECT  119.75 114.57 120.29 114.95 ;
      RECT  138.47 112.99 139.01 113.37 ;
      RECT  122.15 123.57 122.69 124.12 ;
      RECT  128.39 95.92 128.93 96.47 ;
      RECT  128.39 102.72 128.93 103.1 ;
      RECT  115.91 93.24 116.45 93.62 ;
      RECT  119.75 98.77 120.29 99.15 ;
      RECT  103.43 109.04 103.97 109.42 ;
      RECT  109.67 123.57 110.21 124.12 ;
      RECT  122.15 94.82 122.69 95.2 ;
      RECT  140.87 91.97 141.41 92.52 ;
      RECT  125.99 103.82 126.53 104.37 ;
      RECT  103.43 103.82 103.97 104.37 ;
      RECT  97.19 103.82 97.73 104.37 ;
      RECT  134.63 118.52 135.17 118.9 ;
      RECT  103.43 112.99 103.97 113.37 ;
      RECT  128.39 106.67 128.93 107.05 ;
      RECT  119.75 120.89 120.29 121.27 ;
      RECT  103.43 123.57 103.97 124.12 ;
      RECT  107.27 101.14 107.81 101.52 ;
      RECT  103.43 98.77 103.97 99.15 ;
      RECT  140.87 119.62 141.41 120.17 ;
      RECT  115.91 102.72 116.45 103.1 ;
      RECT  97.19 101.14 97.73 101.52 ;
      RECT  97.19 119.62 97.73 120.17 ;
      RECT  122.15 119.62 122.69 120.17 ;
      RECT  144.71 112.99 145.25 113.37 ;
      RECT  119.75 107.77 120.29 108.32 ;
      RECT  115.91 123.57 116.45 124.12 ;
      RECT  128.39 99.87 128.93 100.42 ;
      RECT  132.23 99.87 132.77 100.42 ;
      RECT  103.43 101.14 103.97 101.52 ;
      RECT  144.71 99.87 145.25 100.42 ;
      RECT  125.99 95.92 126.53 96.47 ;
      RECT  101.03 99.87 101.57 100.42 ;
      RECT  144.71 103.82 145.25 104.37 ;
      RECT  125.99 116.94 126.53 117.32 ;
      RECT  113.51 116.94 114.05 117.32 ;
      RECT  128.39 105.09 128.93 105.47 ;
      RECT  107.27 91.97 107.81 92.52 ;
      RECT  132.23 105.09 132.77 105.47 ;
      RECT  122.15 91.97 122.69 92.52 ;
      RECT  144.71 95.92 145.25 96.47 ;
      RECT  119.75 105.09 120.29 105.47 ;
      RECT  134.63 101.14 135.17 101.52 ;
      RECT  122.15 110.62 122.69 111.0 ;
      RECT  138.47 94.82 139.01 95.2 ;
      RECT  134.63 102.72 135.17 103.1 ;
      RECT  97.19 105.09 97.73 105.47 ;
      RECT  103.43 91.97 103.97 92.52 ;
      RECT  119.75 111.72 120.29 112.27 ;
      RECT  122.15 118.52 122.69 118.9 ;
      RECT  132.23 106.67 132.77 107.05 ;
      RECT  134.63 105.09 135.17 105.47 ;
      RECT  119.75 102.72 120.29 103.1 ;
      RECT  97.19 116.94 97.73 117.32 ;
      RECT  125.99 114.57 126.53 114.95 ;
      RECT  107.27 110.62 107.81 111.0 ;
      RECT  138.47 95.92 139.01 96.47 ;
      RECT  134.63 91.97 135.17 92.52 ;
      RECT  140.87 112.99 141.41 113.37 ;
      RECT  122.15 105.09 122.69 105.47 ;
      RECT  115.91 111.72 116.45 112.27 ;
      RECT  103.43 106.67 103.97 107.05 ;
      RECT  113.51 101.14 114.05 101.52 ;
      RECT  107.27 95.92 107.81 96.47 ;
      RECT  132.23 112.99 132.77 113.37 ;
      RECT  122.15 112.99 122.69 113.37 ;
      RECT  115.91 119.62 116.45 120.17 ;
      RECT  140.87 103.82 141.41 104.37 ;
      RECT  138.47 102.72 139.01 103.1 ;
      RECT  134.63 103.82 135.17 104.37 ;
      RECT  132.23 116.94 132.77 117.32 ;
      RECT  109.67 109.04 110.21 109.42 ;
      RECT  144.71 106.67 145.25 107.05 ;
      RECT  132.23 115.67 132.77 116.22 ;
      RECT  107.27 109.04 107.81 109.42 ;
      RECT  107.27 120.89 107.81 121.27 ;
      RECT  125.99 112.99 126.53 113.37 ;
      RECT  122.15 101.14 122.69 101.52 ;
      RECT  132.23 91.97 132.77 92.52 ;
      RECT  107.27 97.19 107.81 97.57 ;
      RECT  103.43 107.77 103.97 108.32 ;
      RECT  101.03 91.97 101.57 92.52 ;
      RECT  107.27 94.82 107.81 95.2 ;
      RECT  115.91 122.47 116.45 122.85 ;
      RECT  128.39 94.82 128.93 95.2 ;
      RECT  97.19 93.24 97.73 93.62 ;
      RECT  144.71 120.89 145.25 121.27 ;
      RECT  119.75 109.04 120.29 109.42 ;
      RECT  101.03 110.62 101.57 111.0 ;
      RECT  115.91 103.82 116.45 104.37 ;
      RECT  109.67 101.14 110.21 101.52 ;
      RECT  107.27 122.47 107.81 122.85 ;
      RECT  125.99 97.19 126.53 97.57 ;
      RECT  128.39 116.94 128.93 117.32 ;
      RECT  109.67 120.89 110.21 121.27 ;
      RECT  113.51 91.97 114.05 92.52 ;
      RECT  122.15 97.19 122.69 97.57 ;
      RECT  109.67 103.82 110.21 104.37 ;
      RECT  144.71 98.77 145.25 99.15 ;
      RECT  134.63 114.57 135.17 114.95 ;
      RECT  119.75 110.62 120.29 111.0 ;
      RECT  107.27 102.72 107.81 103.1 ;
      RECT  134.63 99.87 135.17 100.42 ;
      RECT  101.03 95.92 101.57 96.47 ;
      RECT  101.03 123.57 101.57 124.12 ;
      RECT  107.27 115.67 107.81 116.22 ;
      RECT  144.71 94.82 145.25 95.2 ;
      RECT  113.51 106.67 114.05 107.05 ;
      RECT  138.47 97.19 139.01 97.57 ;
      RECT  140.87 98.77 141.41 99.15 ;
      RECT  122.15 109.04 122.69 109.42 ;
      RECT  138.47 111.72 139.01 112.27 ;
      RECT  101.03 94.82 101.57 95.2 ;
      RECT  138.47 106.67 139.01 107.05 ;
      RECT  125.99 119.62 126.53 120.17 ;
      RECT  132.23 118.52 132.77 118.9 ;
      RECT  115.91 114.57 116.45 114.95 ;
      RECT  109.67 106.67 110.21 107.05 ;
      RECT  119.75 94.82 120.29 95.2 ;
      RECT  97.19 106.67 97.73 107.05 ;
      RECT  144.71 91.97 145.25 92.52 ;
      RECT  109.67 119.62 110.21 120.17 ;
      RECT  134.63 123.57 135.17 124.12 ;
      RECT  113.51 118.52 114.05 118.9 ;
      RECT  140.87 120.89 141.41 121.27 ;
      RECT  132.23 101.14 132.77 101.52 ;
      RECT  119.75 112.99 120.29 113.37 ;
      RECT  140.87 102.72 141.41 103.1 ;
      RECT  144.71 93.24 145.25 93.62 ;
      RECT  134.63 93.24 135.17 93.62 ;
      RECT  101.03 114.57 101.57 114.95 ;
      RECT  115.91 120.89 116.45 121.27 ;
      RECT  128.39 122.47 128.93 122.85 ;
      RECT  132.23 110.62 132.77 111.0 ;
      RECT  101.03 103.82 101.57 104.37 ;
      RECT  97.19 114.57 97.73 114.95 ;
      RECT  101.03 120.89 101.57 121.27 ;
      RECT  119.75 93.24 120.29 93.62 ;
      RECT  107.27 106.67 107.81 107.05 ;
      RECT  115.91 112.99 116.45 113.37 ;
      RECT  101.03 93.24 101.57 93.62 ;
      RECT  144.71 105.09 145.25 105.47 ;
      RECT  132.23 114.57 132.77 114.95 ;
      RECT  140.87 95.92 141.41 96.47 ;
      RECT  132.23 120.89 132.77 121.27 ;
      RECT  140.87 106.67 141.41 107.05 ;
      RECT  113.51 112.99 114.05 113.37 ;
      RECT  144.71 107.77 145.25 108.32 ;
      RECT  103.43 119.62 103.97 120.17 ;
      RECT  125.99 91.97 126.53 92.52 ;
      RECT  107.27 98.77 107.81 99.15 ;
      RECT  122.15 116.94 122.69 117.32 ;
      RECT  128.39 107.77 128.93 108.32 ;
      RECT  101.03 115.67 101.57 116.22 ;
      RECT  132.23 95.92 132.77 96.47 ;
      RECT  140.87 109.04 141.41 109.42 ;
      RECT  125.99 94.82 126.53 95.2 ;
      RECT  138.47 93.24 139.01 93.62 ;
      RECT  115.91 94.82 116.45 95.2 ;
      RECT  103.43 99.87 103.97 100.42 ;
      RECT  119.75 116.94 120.29 117.32 ;
      RECT  128.39 120.89 128.93 121.27 ;
      RECT  113.51 93.24 114.05 93.62 ;
      RECT  97.19 122.47 97.73 122.85 ;
      RECT  128.39 115.67 128.93 116.22 ;
      RECT  103.43 114.57 103.97 114.95 ;
      RECT  132.23 98.77 132.77 99.15 ;
      RECT  140.87 107.77 141.41 108.32 ;
      RECT  138.47 118.52 139.01 118.9 ;
      RECT  119.75 97.19 120.29 97.57 ;
      RECT  125.99 122.47 126.53 122.85 ;
      RECT  138.47 123.57 139.01 124.12 ;
      RECT  113.51 99.87 114.05 100.42 ;
      RECT  97.19 120.89 97.73 121.27 ;
      RECT  109.67 115.67 110.21 116.22 ;
      RECT  144.71 115.67 145.25 116.22 ;
      RECT  103.43 111.72 103.97 112.27 ;
      RECT  132.23 93.24 132.77 93.62 ;
      RECT  138.47 119.62 139.01 120.17 ;
      RECT  122.15 103.82 122.69 104.37 ;
      RECT  125.99 120.89 126.53 121.27 ;
      RECT  128.39 103.82 128.93 104.37 ;
      RECT  122.15 107.77 122.69 108.32 ;
      RECT  134.63 106.67 135.17 107.05 ;
      RECT  115.91 110.62 116.45 111.0 ;
      RECT  125.99 106.67 126.53 107.05 ;
      RECT  125.99 123.57 126.53 124.12 ;
      RECT  134.63 116.94 135.17 117.32 ;
      RECT  119.75 106.67 120.29 107.05 ;
      RECT  134.63 95.92 135.17 96.47 ;
      RECT  125.99 110.62 126.53 111.0 ;
      RECT  101.03 116.94 101.57 117.32 ;
      RECT  107.27 114.57 107.81 114.95 ;
      RECT  101.03 105.09 101.57 105.47 ;
      RECT  144.71 97.19 145.25 97.57 ;
      RECT  128.39 109.04 128.93 109.42 ;
      RECT  103.43 97.19 103.97 97.57 ;
      RECT  140.87 101.14 141.41 101.52 ;
      RECT  103.43 95.92 103.97 96.47 ;
      RECT  97.19 111.72 97.73 112.27 ;
      RECT  109.67 95.92 110.21 96.47 ;
      RECT  122.15 120.89 122.69 121.27 ;
      RECT  109.67 112.99 110.21 113.37 ;
      RECT  138.47 109.04 139.01 109.42 ;
      RECT  128.39 97.19 128.93 97.57 ;
      RECT  97.19 97.19 97.73 97.57 ;
      RECT  144.71 122.47 145.25 122.85 ;
      RECT  128.39 93.24 128.93 93.62 ;
      RECT  103.43 118.52 103.97 118.9 ;
      RECT  128.39 101.14 128.93 101.52 ;
      RECT  113.51 102.72 114.05 103.1 ;
      RECT  109.67 114.57 110.21 114.95 ;
      RECT  128.39 112.99 128.93 113.37 ;
      RECT  101.03 111.72 101.57 112.27 ;
      RECT  132.23 119.62 132.77 120.17 ;
      RECT  132.23 102.72 132.77 103.1 ;
      RECT  144.71 102.72 145.25 103.1 ;
      RECT  134.63 122.47 135.17 122.85 ;
      RECT  138.47 103.82 139.01 104.37 ;
      RECT  140.87 93.24 141.41 93.62 ;
      RECT  113.51 122.47 114.05 122.85 ;
      RECT  119.75 103.82 120.29 104.37 ;
      RECT  101.03 109.04 101.57 109.42 ;
      RECT  101.03 112.99 101.57 113.37 ;
      RECT  109.67 107.77 110.21 108.32 ;
      RECT  109.67 94.82 110.21 95.2 ;
      RECT  101.03 122.47 101.57 122.85 ;
      RECT  115.91 106.67 116.45 107.05 ;
      RECT  115.91 95.92 116.45 96.47 ;
      RECT  97.19 112.99 97.73 113.37 ;
      RECT  103.43 93.24 103.97 93.62 ;
      RECT  107.27 123.57 107.81 124.12 ;
      RECT  113.51 107.77 114.05 108.32 ;
      RECT  103.43 105.09 103.97 105.47 ;
      RECT  128.39 119.62 128.93 120.17 ;
      RECT  97.19 98.77 97.73 99.15 ;
      RECT  128.39 98.77 128.93 99.15 ;
      RECT  107.27 93.24 107.81 93.62 ;
      RECT  115.91 107.77 116.45 108.32 ;
      RECT  132.23 123.57 132.77 124.12 ;
      RECT  132.23 122.47 132.77 122.85 ;
      RECT  113.51 103.82 114.05 104.37 ;
      RECT  140.87 114.57 141.41 114.95 ;
      RECT  115.91 99.87 116.45 100.42 ;
      RECT  138.47 91.97 139.01 92.52 ;
      RECT  107.27 103.82 107.81 104.37 ;
      RECT  125.99 99.87 126.53 100.42 ;
      RECT  134.63 110.62 135.17 111.0 ;
      RECT  107.27 116.94 107.81 117.32 ;
      RECT  144.71 116.94 145.25 117.32 ;
      RECT  125.99 118.52 126.53 118.9 ;
      RECT  107.27 105.09 107.81 105.47 ;
      RECT  97.19 115.67 97.73 116.22 ;
      RECT  125.99 101.14 126.53 101.52 ;
      RECT  134.63 107.77 135.17 108.32 ;
      RECT  134.63 120.89 135.17 121.27 ;
      RECT  125.99 102.72 126.53 103.1 ;
      RECT  109.67 116.94 110.21 117.32 ;
      RECT  128.39 110.62 128.93 111.0 ;
      RECT  119.75 115.67 120.29 116.22 ;
      RECT  128.39 91.97 128.93 92.52 ;
      RECT  144.71 109.04 145.25 109.42 ;
      RECT  97.19 118.52 97.73 118.9 ;
      RECT  132.23 94.82 132.77 95.2 ;
      RECT  144.71 101.14 145.25 101.52 ;
      RECT  107.27 111.72 107.81 112.27 ;
      RECT  128.39 123.57 128.93 124.12 ;
      RECT  101.03 98.77 101.57 99.15 ;
      RECT  125.99 109.04 126.53 109.42 ;
      RECT  122.15 111.72 122.69 112.27 ;
      RECT  138.47 107.77 139.01 108.32 ;
      RECT  140.87 122.47 141.41 122.85 ;
      RECT  134.63 109.04 135.17 109.42 ;
      RECT  103.43 94.82 103.97 95.2 ;
      RECT  97.19 99.87 97.73 100.42 ;
      RECT  107.27 112.99 107.81 113.37 ;
      RECT  109.67 122.47 110.21 122.85 ;
      RECT  138.47 98.77 139.01 99.15 ;
      RECT  132.23 97.19 132.77 97.57 ;
      RECT  140.87 97.19 141.41 97.57 ;
      RECT  140.87 111.72 141.41 112.27 ;
      RECT  140.87 110.62 141.41 111.0 ;
      RECT  113.51 119.62 114.05 120.17 ;
      RECT  122.15 99.87 122.69 100.42 ;
      RECT  97.19 107.77 97.73 108.32 ;
      RECT  115.91 115.67 116.45 116.22 ;
      RECT  119.75 122.47 120.29 122.85 ;
      RECT  138.47 114.57 139.01 114.95 ;
      RECT  96.26 89.165 93.14 89.715 ;
      RECT  96.47 91.25 95.33 90.87 ;
      RECT  94.07 91.49 93.86 91.42 ;
      RECT  93.86 90.63 93.35 90.39 ;
      RECT  96.26 91.73 93.86 91.49 ;
      RECT  93.86 91.49 93.66 91.42 ;
      RECT  94.07 90.7 93.86 90.63 ;
      RECT  93.35 91.73 93.14 91.49 ;
      POLYGON  94.79 91.25 94.79 90.87 94.24 90.87 94.24 90.94 93.86 90.94 93.86 91.18 94.24 91.18 94.24 91.25 94.79 91.25 ;
      RECT  93.35 91.25 93.14 90.87 ;
      RECT  96.47 92.52 96.26 91.97 ;
      RECT  96.26 92.52 95.33 91.97 ;
      RECT  95.33 91.25 94.79 90.87 ;
      RECT  93.35 90.63 93.14 90.39 ;
      RECT  94.79 92.52 93.14 91.97 ;
      RECT  96.47 91.73 96.26 91.49 ;
      RECT  93.86 90.7 93.66 90.63 ;
      POLYGON  93.49 91.25 93.49 91.18 93.86 91.18 93.86 90.94 93.49 90.94 93.49 90.87 93.35 90.87 93.35 91.25 93.49 91.25 ;
      RECT  96.47 90.63 96.26 90.39 ;
      RECT  96.26 90.63 93.86 90.39 ;
      RECT  93.86 91.73 93.35 91.49 ;
      RECT  95.33 92.52 94.79 91.97 ;
      RECT  96.47 93.24 95.33 93.62 ;
      RECT  94.07 93.0 93.86 93.07 ;
      RECT  93.86 93.86 93.35 94.1 ;
      RECT  96.26 92.76 93.86 93.0 ;
      RECT  93.86 93.0 93.66 93.07 ;
      RECT  94.07 93.79 93.86 93.86 ;
      RECT  93.35 92.76 93.14 93.0 ;
      POLYGON  94.79 93.24 94.79 93.62 94.24 93.62 94.24 93.55 93.86 93.55 93.86 93.31 94.24 93.31 94.24 93.24 94.79 93.24 ;
      RECT  93.35 93.24 93.14 93.62 ;
      RECT  96.47 91.97 96.26 92.52 ;
      RECT  96.26 91.97 95.33 92.52 ;
      RECT  95.33 93.24 94.79 93.62 ;
      RECT  93.35 93.86 93.14 94.1 ;
      RECT  94.79 91.97 93.14 92.52 ;
      RECT  96.47 92.76 96.26 93.0 ;
      RECT  93.86 93.79 93.66 93.86 ;
      POLYGON  93.49 93.24 93.49 93.31 93.86 93.31 93.86 93.55 93.49 93.55 93.49 93.62 93.35 93.62 93.35 93.24 93.49 93.24 ;
      RECT  96.47 93.86 96.26 94.1 ;
      RECT  96.26 93.86 93.86 94.1 ;
      RECT  93.86 92.76 93.35 93.0 ;
      RECT  95.33 91.97 94.79 92.52 ;
      RECT  96.47 95.2 95.33 94.82 ;
      RECT  94.07 95.44 93.86 95.37 ;
      RECT  93.86 94.58 93.35 94.34 ;
      RECT  96.26 95.68 93.86 95.44 ;
      RECT  93.86 95.44 93.66 95.37 ;
      RECT  94.07 94.65 93.86 94.58 ;
      RECT  93.35 95.68 93.14 95.44 ;
      POLYGON  94.79 95.2 94.79 94.82 94.24 94.82 94.24 94.89 93.86 94.89 93.86 95.13 94.24 95.13 94.24 95.2 94.79 95.2 ;
      RECT  93.35 95.2 93.14 94.82 ;
      RECT  96.47 96.47 96.26 95.92 ;
      RECT  96.26 96.47 95.33 95.92 ;
      RECT  95.33 95.2 94.79 94.82 ;
      RECT  93.35 94.58 93.14 94.34 ;
      RECT  94.79 96.47 93.14 95.92 ;
      RECT  96.47 95.68 96.26 95.44 ;
      RECT  93.86 94.65 93.66 94.58 ;
      POLYGON  93.49 95.2 93.49 95.13 93.86 95.13 93.86 94.89 93.49 94.89 93.49 94.82 93.35 94.82 93.35 95.2 93.49 95.2 ;
      RECT  96.47 94.58 96.26 94.34 ;
      RECT  96.26 94.58 93.86 94.34 ;
      RECT  93.86 95.68 93.35 95.44 ;
      RECT  95.33 96.47 94.79 95.92 ;
      RECT  96.47 97.19 95.33 97.57 ;
      RECT  94.07 96.95 93.86 97.02 ;
      RECT  93.86 97.81 93.35 98.05 ;
      RECT  96.26 96.71 93.86 96.95 ;
      RECT  93.86 96.95 93.66 97.02 ;
      RECT  94.07 97.74 93.86 97.81 ;
      RECT  93.35 96.71 93.14 96.95 ;
      POLYGON  94.79 97.19 94.79 97.57 94.24 97.57 94.24 97.5 93.86 97.5 93.86 97.26 94.24 97.26 94.24 97.19 94.79 97.19 ;
      RECT  93.35 97.19 93.14 97.57 ;
      RECT  96.47 95.92 96.26 96.47 ;
      RECT  96.26 95.92 95.33 96.47 ;
      RECT  95.33 97.19 94.79 97.57 ;
      RECT  93.35 97.81 93.14 98.05 ;
      RECT  94.79 95.92 93.14 96.47 ;
      RECT  96.47 96.71 96.26 96.95 ;
      RECT  93.86 97.74 93.66 97.81 ;
      POLYGON  93.49 97.19 93.49 97.26 93.86 97.26 93.86 97.5 93.49 97.5 93.49 97.57 93.35 97.57 93.35 97.19 93.49 97.19 ;
      RECT  96.47 97.81 96.26 98.05 ;
      RECT  96.26 97.81 93.86 98.05 ;
      RECT  93.86 96.71 93.35 96.95 ;
      RECT  95.33 95.92 94.79 96.47 ;
      RECT  96.47 99.15 95.33 98.77 ;
      RECT  94.07 99.39 93.86 99.32 ;
      RECT  93.86 98.53 93.35 98.29 ;
      RECT  96.26 99.63 93.86 99.39 ;
      RECT  93.86 99.39 93.66 99.32 ;
      RECT  94.07 98.6 93.86 98.53 ;
      RECT  93.35 99.63 93.14 99.39 ;
      POLYGON  94.79 99.15 94.79 98.77 94.24 98.77 94.24 98.84 93.86 98.84 93.86 99.08 94.24 99.08 94.24 99.15 94.79 99.15 ;
      RECT  93.35 99.15 93.14 98.77 ;
      RECT  96.47 100.42 96.26 99.87 ;
      RECT  96.26 100.42 95.33 99.87 ;
      RECT  95.33 99.15 94.79 98.77 ;
      RECT  93.35 98.53 93.14 98.29 ;
      RECT  94.79 100.42 93.14 99.87 ;
      RECT  96.47 99.63 96.26 99.39 ;
      RECT  93.86 98.6 93.66 98.53 ;
      POLYGON  93.49 99.15 93.49 99.08 93.86 99.08 93.86 98.84 93.49 98.84 93.49 98.77 93.35 98.77 93.35 99.15 93.49 99.15 ;
      RECT  96.47 98.53 96.26 98.29 ;
      RECT  96.26 98.53 93.86 98.29 ;
      RECT  93.86 99.63 93.35 99.39 ;
      RECT  95.33 100.42 94.79 99.87 ;
      RECT  96.47 101.14 95.33 101.52 ;
      RECT  94.07 100.9 93.86 100.97 ;
      RECT  93.86 101.76 93.35 102.0 ;
      RECT  96.26 100.66 93.86 100.9 ;
      RECT  93.86 100.9 93.66 100.97 ;
      RECT  94.07 101.69 93.86 101.76 ;
      RECT  93.35 100.66 93.14 100.9 ;
      POLYGON  94.79 101.14 94.79 101.52 94.24 101.52 94.24 101.45 93.86 101.45 93.86 101.21 94.24 101.21 94.24 101.14 94.79 101.14 ;
      RECT  93.35 101.14 93.14 101.52 ;
      RECT  96.47 99.87 96.26 100.42 ;
      RECT  96.26 99.87 95.33 100.42 ;
      RECT  95.33 101.14 94.79 101.52 ;
      RECT  93.35 101.76 93.14 102.0 ;
      RECT  94.79 99.87 93.14 100.42 ;
      RECT  96.47 100.66 96.26 100.9 ;
      RECT  93.86 101.69 93.66 101.76 ;
      POLYGON  93.49 101.14 93.49 101.21 93.86 101.21 93.86 101.45 93.49 101.45 93.49 101.52 93.35 101.52 93.35 101.14 93.49 101.14 ;
      RECT  96.47 101.76 96.26 102.0 ;
      RECT  96.26 101.76 93.86 102.0 ;
      RECT  93.86 100.66 93.35 100.9 ;
      RECT  95.33 99.87 94.79 100.42 ;
      RECT  96.47 103.1 95.33 102.72 ;
      RECT  94.07 103.34 93.86 103.27 ;
      RECT  93.86 102.48 93.35 102.24 ;
      RECT  96.26 103.58 93.86 103.34 ;
      RECT  93.86 103.34 93.66 103.27 ;
      RECT  94.07 102.55 93.86 102.48 ;
      RECT  93.35 103.58 93.14 103.34 ;
      POLYGON  94.79 103.1 94.79 102.72 94.24 102.72 94.24 102.79 93.86 102.79 93.86 103.03 94.24 103.03 94.24 103.1 94.79 103.1 ;
      RECT  93.35 103.1 93.14 102.72 ;
      RECT  96.47 104.37 96.26 103.82 ;
      RECT  96.26 104.37 95.33 103.82 ;
      RECT  95.33 103.1 94.79 102.72 ;
      RECT  93.35 102.48 93.14 102.24 ;
      RECT  94.79 104.37 93.14 103.82 ;
      RECT  96.47 103.58 96.26 103.34 ;
      RECT  93.86 102.55 93.66 102.48 ;
      POLYGON  93.49 103.1 93.49 103.03 93.86 103.03 93.86 102.79 93.49 102.79 93.49 102.72 93.35 102.72 93.35 103.1 93.49 103.1 ;
      RECT  96.47 102.48 96.26 102.24 ;
      RECT  96.26 102.48 93.86 102.24 ;
      RECT  93.86 103.58 93.35 103.34 ;
      RECT  95.33 104.37 94.79 103.82 ;
      RECT  96.47 105.09 95.33 105.47 ;
      RECT  94.07 104.85 93.86 104.92 ;
      RECT  93.86 105.71 93.35 105.95 ;
      RECT  96.26 104.61 93.86 104.85 ;
      RECT  93.86 104.85 93.66 104.92 ;
      RECT  94.07 105.64 93.86 105.71 ;
      RECT  93.35 104.61 93.14 104.85 ;
      POLYGON  94.79 105.09 94.79 105.47 94.24 105.47 94.24 105.4 93.86 105.4 93.86 105.16 94.24 105.16 94.24 105.09 94.79 105.09 ;
      RECT  93.35 105.09 93.14 105.47 ;
      RECT  96.47 103.82 96.26 104.37 ;
      RECT  96.26 103.82 95.33 104.37 ;
      RECT  95.33 105.09 94.79 105.47 ;
      RECT  93.35 105.71 93.14 105.95 ;
      RECT  94.79 103.82 93.14 104.37 ;
      RECT  96.47 104.61 96.26 104.85 ;
      RECT  93.86 105.64 93.66 105.71 ;
      POLYGON  93.49 105.09 93.49 105.16 93.86 105.16 93.86 105.4 93.49 105.4 93.49 105.47 93.35 105.47 93.35 105.09 93.49 105.09 ;
      RECT  96.47 105.71 96.26 105.95 ;
      RECT  96.26 105.71 93.86 105.95 ;
      RECT  93.86 104.61 93.35 104.85 ;
      RECT  95.33 103.82 94.79 104.37 ;
      RECT  96.47 107.05 95.33 106.67 ;
      RECT  94.07 107.29 93.86 107.22 ;
      RECT  93.86 106.43 93.35 106.19 ;
      RECT  96.26 107.53 93.86 107.29 ;
      RECT  93.86 107.29 93.66 107.22 ;
      RECT  94.07 106.5 93.86 106.43 ;
      RECT  93.35 107.53 93.14 107.29 ;
      POLYGON  94.79 107.05 94.79 106.67 94.24 106.67 94.24 106.74 93.86 106.74 93.86 106.98 94.24 106.98 94.24 107.05 94.79 107.05 ;
      RECT  93.35 107.05 93.14 106.67 ;
      RECT  96.47 108.32 96.26 107.77 ;
      RECT  96.26 108.32 95.33 107.77 ;
      RECT  95.33 107.05 94.79 106.67 ;
      RECT  93.35 106.43 93.14 106.19 ;
      RECT  94.79 108.32 93.14 107.77 ;
      RECT  96.47 107.53 96.26 107.29 ;
      RECT  93.86 106.5 93.66 106.43 ;
      POLYGON  93.49 107.05 93.49 106.98 93.86 106.98 93.86 106.74 93.49 106.74 93.49 106.67 93.35 106.67 93.35 107.05 93.49 107.05 ;
      RECT  96.47 106.43 96.26 106.19 ;
      RECT  96.26 106.43 93.86 106.19 ;
      RECT  93.86 107.53 93.35 107.29 ;
      RECT  95.33 108.32 94.79 107.77 ;
      RECT  96.47 109.04 95.33 109.42 ;
      RECT  94.07 108.8 93.86 108.87 ;
      RECT  93.86 109.66 93.35 109.9 ;
      RECT  96.26 108.56 93.86 108.8 ;
      RECT  93.86 108.8 93.66 108.87 ;
      RECT  94.07 109.59 93.86 109.66 ;
      RECT  93.35 108.56 93.14 108.8 ;
      POLYGON  94.79 109.04 94.79 109.42 94.24 109.42 94.24 109.35 93.86 109.35 93.86 109.11 94.24 109.11 94.24 109.04 94.79 109.04 ;
      RECT  93.35 109.04 93.14 109.42 ;
      RECT  96.47 107.77 96.26 108.32 ;
      RECT  96.26 107.77 95.33 108.32 ;
      RECT  95.33 109.04 94.79 109.42 ;
      RECT  93.35 109.66 93.14 109.9 ;
      RECT  94.79 107.77 93.14 108.32 ;
      RECT  96.47 108.56 96.26 108.8 ;
      RECT  93.86 109.59 93.66 109.66 ;
      POLYGON  93.49 109.04 93.49 109.11 93.86 109.11 93.86 109.35 93.49 109.35 93.49 109.42 93.35 109.42 93.35 109.04 93.49 109.04 ;
      RECT  96.47 109.66 96.26 109.9 ;
      RECT  96.26 109.66 93.86 109.9 ;
      RECT  93.86 108.56 93.35 108.8 ;
      RECT  95.33 107.77 94.79 108.32 ;
      RECT  96.47 111.0 95.33 110.62 ;
      RECT  94.07 111.24 93.86 111.17 ;
      RECT  93.86 110.38 93.35 110.14 ;
      RECT  96.26 111.48 93.86 111.24 ;
      RECT  93.86 111.24 93.66 111.17 ;
      RECT  94.07 110.45 93.86 110.38 ;
      RECT  93.35 111.48 93.14 111.24 ;
      POLYGON  94.79 111.0 94.79 110.62 94.24 110.62 94.24 110.69 93.86 110.69 93.86 110.93 94.24 110.93 94.24 111.0 94.79 111.0 ;
      RECT  93.35 111.0 93.14 110.62 ;
      RECT  96.47 112.27 96.26 111.72 ;
      RECT  96.26 112.27 95.33 111.72 ;
      RECT  95.33 111.0 94.79 110.62 ;
      RECT  93.35 110.38 93.14 110.14 ;
      RECT  94.79 112.27 93.14 111.72 ;
      RECT  96.47 111.48 96.26 111.24 ;
      RECT  93.86 110.45 93.66 110.38 ;
      POLYGON  93.49 111.0 93.49 110.93 93.86 110.93 93.86 110.69 93.49 110.69 93.49 110.62 93.35 110.62 93.35 111.0 93.49 111.0 ;
      RECT  96.47 110.38 96.26 110.14 ;
      RECT  96.26 110.38 93.86 110.14 ;
      RECT  93.86 111.48 93.35 111.24 ;
      RECT  95.33 112.27 94.79 111.72 ;
      RECT  96.47 112.99 95.33 113.37 ;
      RECT  94.07 112.75 93.86 112.82 ;
      RECT  93.86 113.61 93.35 113.85 ;
      RECT  96.26 112.51 93.86 112.75 ;
      RECT  93.86 112.75 93.66 112.82 ;
      RECT  94.07 113.54 93.86 113.61 ;
      RECT  93.35 112.51 93.14 112.75 ;
      POLYGON  94.79 112.99 94.79 113.37 94.24 113.37 94.24 113.3 93.86 113.3 93.86 113.06 94.24 113.06 94.24 112.99 94.79 112.99 ;
      RECT  93.35 112.99 93.14 113.37 ;
      RECT  96.47 111.72 96.26 112.27 ;
      RECT  96.26 111.72 95.33 112.27 ;
      RECT  95.33 112.99 94.79 113.37 ;
      RECT  93.35 113.61 93.14 113.85 ;
      RECT  94.79 111.72 93.14 112.27 ;
      RECT  96.47 112.51 96.26 112.75 ;
      RECT  93.86 113.54 93.66 113.61 ;
      POLYGON  93.49 112.99 93.49 113.06 93.86 113.06 93.86 113.3 93.49 113.3 93.49 113.37 93.35 113.37 93.35 112.99 93.49 112.99 ;
      RECT  96.47 113.61 96.26 113.85 ;
      RECT  96.26 113.61 93.86 113.85 ;
      RECT  93.86 112.51 93.35 112.75 ;
      RECT  95.33 111.72 94.79 112.27 ;
      RECT  96.47 114.95 95.33 114.57 ;
      RECT  94.07 115.19 93.86 115.12 ;
      RECT  93.86 114.33 93.35 114.09 ;
      RECT  96.26 115.43 93.86 115.19 ;
      RECT  93.86 115.19 93.66 115.12 ;
      RECT  94.07 114.4 93.86 114.33 ;
      RECT  93.35 115.43 93.14 115.19 ;
      POLYGON  94.79 114.95 94.79 114.57 94.24 114.57 94.24 114.64 93.86 114.64 93.86 114.88 94.24 114.88 94.24 114.95 94.79 114.95 ;
      RECT  93.35 114.95 93.14 114.57 ;
      RECT  96.47 116.22 96.26 115.67 ;
      RECT  96.26 116.22 95.33 115.67 ;
      RECT  95.33 114.95 94.79 114.57 ;
      RECT  93.35 114.33 93.14 114.09 ;
      RECT  94.79 116.22 93.14 115.67 ;
      RECT  96.47 115.43 96.26 115.19 ;
      RECT  93.86 114.4 93.66 114.33 ;
      POLYGON  93.49 114.95 93.49 114.88 93.86 114.88 93.86 114.64 93.49 114.64 93.49 114.57 93.35 114.57 93.35 114.95 93.49 114.95 ;
      RECT  96.47 114.33 96.26 114.09 ;
      RECT  96.26 114.33 93.86 114.09 ;
      RECT  93.86 115.43 93.35 115.19 ;
      RECT  95.33 116.22 94.79 115.67 ;
      RECT  96.47 116.94 95.33 117.32 ;
      RECT  94.07 116.7 93.86 116.77 ;
      RECT  93.86 117.56 93.35 117.8 ;
      RECT  96.26 116.46 93.86 116.7 ;
      RECT  93.86 116.7 93.66 116.77 ;
      RECT  94.07 117.49 93.86 117.56 ;
      RECT  93.35 116.46 93.14 116.7 ;
      POLYGON  94.79 116.94 94.79 117.32 94.24 117.32 94.24 117.25 93.86 117.25 93.86 117.01 94.24 117.01 94.24 116.94 94.79 116.94 ;
      RECT  93.35 116.94 93.14 117.32 ;
      RECT  96.47 115.67 96.26 116.22 ;
      RECT  96.26 115.67 95.33 116.22 ;
      RECT  95.33 116.94 94.79 117.32 ;
      RECT  93.35 117.56 93.14 117.8 ;
      RECT  94.79 115.67 93.14 116.22 ;
      RECT  96.47 116.46 96.26 116.7 ;
      RECT  93.86 117.49 93.66 117.56 ;
      POLYGON  93.49 116.94 93.49 117.01 93.86 117.01 93.86 117.25 93.49 117.25 93.49 117.32 93.35 117.32 93.35 116.94 93.49 116.94 ;
      RECT  96.47 117.56 96.26 117.8 ;
      RECT  96.26 117.56 93.86 117.8 ;
      RECT  93.86 116.46 93.35 116.7 ;
      RECT  95.33 115.67 94.79 116.22 ;
      RECT  96.47 118.9 95.33 118.52 ;
      RECT  94.07 119.14 93.86 119.07 ;
      RECT  93.86 118.28 93.35 118.04 ;
      RECT  96.26 119.38 93.86 119.14 ;
      RECT  93.86 119.14 93.66 119.07 ;
      RECT  94.07 118.35 93.86 118.28 ;
      RECT  93.35 119.38 93.14 119.14 ;
      POLYGON  94.79 118.9 94.79 118.52 94.24 118.52 94.24 118.59 93.86 118.59 93.86 118.83 94.24 118.83 94.24 118.9 94.79 118.9 ;
      RECT  93.35 118.9 93.14 118.52 ;
      RECT  96.47 120.17 96.26 119.62 ;
      RECT  96.26 120.17 95.33 119.62 ;
      RECT  95.33 118.9 94.79 118.52 ;
      RECT  93.35 118.28 93.14 118.04 ;
      RECT  94.79 120.17 93.14 119.62 ;
      RECT  96.47 119.38 96.26 119.14 ;
      RECT  93.86 118.35 93.66 118.28 ;
      POLYGON  93.49 118.9 93.49 118.83 93.86 118.83 93.86 118.59 93.49 118.59 93.49 118.52 93.35 118.52 93.35 118.9 93.49 118.9 ;
      RECT  96.47 118.28 96.26 118.04 ;
      RECT  96.26 118.28 93.86 118.04 ;
      RECT  93.86 119.38 93.35 119.14 ;
      RECT  95.33 120.17 94.79 119.62 ;
      RECT  96.47 120.89 95.33 121.27 ;
      RECT  94.07 120.65 93.86 120.72 ;
      RECT  93.86 121.51 93.35 121.75 ;
      RECT  96.26 120.41 93.86 120.65 ;
      RECT  93.86 120.65 93.66 120.72 ;
      RECT  94.07 121.44 93.86 121.51 ;
      RECT  93.35 120.41 93.14 120.65 ;
      POLYGON  94.79 120.89 94.79 121.27 94.24 121.27 94.24 121.2 93.86 121.2 93.86 120.96 94.24 120.96 94.24 120.89 94.79 120.89 ;
      RECT  93.35 120.89 93.14 121.27 ;
      RECT  96.47 119.62 96.26 120.17 ;
      RECT  96.26 119.62 95.33 120.17 ;
      RECT  95.33 120.89 94.79 121.27 ;
      RECT  93.35 121.51 93.14 121.75 ;
      RECT  94.79 119.62 93.14 120.17 ;
      RECT  96.47 120.41 96.26 120.65 ;
      RECT  93.86 121.44 93.66 121.51 ;
      POLYGON  93.49 120.89 93.49 120.96 93.86 120.96 93.86 121.2 93.49 121.2 93.49 121.27 93.35 121.27 93.35 120.89 93.49 120.89 ;
      RECT  96.47 121.51 96.26 121.75 ;
      RECT  96.26 121.51 93.86 121.75 ;
      RECT  93.86 120.41 93.35 120.65 ;
      RECT  95.33 119.62 94.79 120.17 ;
      RECT  96.47 122.85 95.33 122.47 ;
      RECT  94.07 123.09 93.86 123.02 ;
      RECT  93.86 122.23 93.35 121.99 ;
      RECT  96.26 123.33 93.86 123.09 ;
      RECT  93.86 123.09 93.66 123.02 ;
      RECT  94.07 122.3 93.86 122.23 ;
      RECT  93.35 123.33 93.14 123.09 ;
      POLYGON  94.79 122.85 94.79 122.47 94.24 122.47 94.24 122.54 93.86 122.54 93.86 122.78 94.24 122.78 94.24 122.85 94.79 122.85 ;
      RECT  93.35 122.85 93.14 122.47 ;
      RECT  96.47 124.12 96.26 123.57 ;
      RECT  96.26 124.12 95.33 123.57 ;
      RECT  95.33 122.85 94.79 122.47 ;
      RECT  93.35 122.23 93.14 121.99 ;
      RECT  94.79 124.12 93.14 123.57 ;
      RECT  96.47 123.33 96.26 123.09 ;
      RECT  93.86 122.3 93.66 122.23 ;
      POLYGON  93.49 122.85 93.49 122.78 93.86 122.78 93.86 122.54 93.49 122.54 93.49 122.47 93.35 122.47 93.35 122.85 93.49 122.85 ;
      RECT  96.47 122.23 96.26 121.99 ;
      RECT  96.26 122.23 93.86 121.99 ;
      RECT  93.86 123.33 93.35 123.09 ;
      RECT  95.33 124.12 94.79 123.57 ;
      RECT  96.47 124.84 95.33 125.22 ;
      RECT  94.07 124.6 93.86 124.67 ;
      RECT  93.86 125.46 93.35 125.7 ;
      RECT  96.26 124.36 93.86 124.6 ;
      RECT  93.86 124.6 93.66 124.67 ;
      RECT  94.07 125.39 93.86 125.46 ;
      RECT  93.35 124.36 93.14 124.6 ;
      POLYGON  94.79 124.84 94.79 125.22 94.24 125.22 94.24 125.15 93.86 125.15 93.86 124.91 94.24 124.91 94.24 124.84 94.79 124.84 ;
      RECT  93.35 124.84 93.14 125.22 ;
      RECT  96.47 123.57 96.26 124.12 ;
      RECT  96.26 123.57 95.33 124.12 ;
      RECT  95.33 124.84 94.79 125.22 ;
      RECT  93.35 125.46 93.14 125.7 ;
      RECT  94.79 123.57 93.14 124.12 ;
      RECT  96.47 124.36 96.26 124.6 ;
      RECT  93.86 125.39 93.66 125.46 ;
      POLYGON  93.49 124.84 93.49 124.91 93.86 124.91 93.86 125.15 93.49 125.15 93.49 125.22 93.35 125.22 93.35 124.84 93.49 124.84 ;
      RECT  96.47 125.46 96.26 125.7 ;
      RECT  96.26 125.46 93.86 125.7 ;
      RECT  93.86 124.36 93.35 124.6 ;
      RECT  95.33 123.57 94.79 124.12 ;
      RECT  96.26 126.925 93.14 126.375 ;
      RECT  93.14 90.39 96.26 90.63 ;
      RECT  93.14 91.49 96.26 91.73 ;
      RECT  93.14 93.86 96.26 94.1 ;
      RECT  93.14 92.76 96.26 93.0 ;
      RECT  93.14 94.34 96.26 94.58 ;
      RECT  93.14 95.44 96.26 95.68 ;
      RECT  93.14 97.81 96.26 98.05 ;
      RECT  93.14 96.71 96.26 96.95 ;
      RECT  93.14 98.29 96.26 98.53 ;
      RECT  93.14 99.39 96.26 99.63 ;
      RECT  93.14 101.76 96.26 102.0 ;
      RECT  93.14 100.66 96.26 100.9 ;
      RECT  93.14 102.24 96.26 102.48 ;
      RECT  93.14 103.34 96.26 103.58 ;
      RECT  93.14 105.71 96.26 105.95 ;
      RECT  93.14 104.61 96.26 104.85 ;
      RECT  93.14 106.19 96.26 106.43 ;
      RECT  93.14 107.29 96.26 107.53 ;
      RECT  93.14 109.66 96.26 109.9 ;
      RECT  93.14 108.56 96.26 108.8 ;
      RECT  93.14 110.14 96.26 110.38 ;
      RECT  93.14 111.24 96.26 111.48 ;
      RECT  93.14 113.61 96.26 113.85 ;
      RECT  93.14 112.51 96.26 112.75 ;
      RECT  93.14 114.09 96.26 114.33 ;
      RECT  93.14 115.19 96.26 115.43 ;
      RECT  93.14 117.56 96.26 117.8 ;
      RECT  93.14 116.46 96.26 116.7 ;
      RECT  93.14 118.04 96.26 118.28 ;
      RECT  93.14 119.14 96.26 119.38 ;
      RECT  93.14 121.51 96.26 121.75 ;
      RECT  93.14 120.41 96.26 120.65 ;
      RECT  93.14 121.99 96.26 122.23 ;
      RECT  93.14 123.09 96.26 123.33 ;
      RECT  93.14 125.46 96.26 125.7 ;
      RECT  93.14 124.36 96.26 124.6 ;
      RECT  94.79 124.84 95.33 125.22 ;
      RECT  94.79 112.99 95.33 113.37 ;
      RECT  94.79 109.04 95.33 109.42 ;
      RECT  94.79 97.19 95.33 97.57 ;
      RECT  94.79 119.62 95.33 120.17 ;
      RECT  94.79 118.52 95.33 118.9 ;
      RECT  94.79 99.87 95.33 100.42 ;
      RECT  94.79 91.97 95.33 92.52 ;
      RECT  94.79 111.72 95.33 112.27 ;
      RECT  94.79 101.14 95.33 101.52 ;
      RECT  94.79 122.47 95.33 122.85 ;
      RECT  94.79 94.82 95.33 95.2 ;
      RECT  94.79 102.72 95.33 103.1 ;
      RECT  94.79 93.24 95.33 93.62 ;
      RECT  94.79 98.77 95.33 99.15 ;
      RECT  94.79 115.67 95.33 116.22 ;
      RECT  94.79 116.94 95.33 117.32 ;
      RECT  94.79 107.77 95.33 108.32 ;
      RECT  94.79 95.92 95.33 96.47 ;
      RECT  94.79 105.09 95.33 105.47 ;
      RECT  94.79 123.57 95.33 124.12 ;
      RECT  94.79 106.67 95.33 107.05 ;
      RECT  94.79 90.87 95.33 91.25 ;
      RECT  94.79 110.62 95.33 111.0 ;
      RECT  94.79 114.57 95.33 114.95 ;
      RECT  94.79 120.89 95.33 121.27 ;
      RECT  94.79 103.82 95.33 104.37 ;
      RECT  146.18 89.165 149.3 89.715 ;
      RECT  145.97 91.25 147.11 90.87 ;
      RECT  148.37 91.49 148.58 91.42 ;
      RECT  148.58 90.63 149.09 90.39 ;
      RECT  146.18 91.73 148.58 91.49 ;
      RECT  148.58 91.49 148.78 91.42 ;
      RECT  148.37 90.7 148.58 90.63 ;
      RECT  149.09 91.73 149.3 91.49 ;
      POLYGON  147.65 91.25 147.65 90.87 148.2 90.87 148.2 90.94 148.58 90.94 148.58 91.18 148.2 91.18 148.2 91.25 147.65 91.25 ;
      RECT  149.09 91.25 149.3 90.87 ;
      RECT  145.97 92.52 146.18 91.97 ;
      RECT  146.18 92.52 147.11 91.97 ;
      RECT  147.11 91.25 147.65 90.87 ;
      RECT  149.09 90.63 149.3 90.39 ;
      RECT  147.65 92.52 149.3 91.97 ;
      RECT  145.97 91.73 146.18 91.49 ;
      RECT  148.58 90.7 148.78 90.63 ;
      POLYGON  148.95 91.25 148.95 91.18 148.58 91.18 148.58 90.94 148.95 90.94 148.95 90.87 149.09 90.87 149.09 91.25 148.95 91.25 ;
      RECT  145.97 90.63 146.18 90.39 ;
      RECT  146.18 90.63 148.58 90.39 ;
      RECT  148.58 91.73 149.09 91.49 ;
      RECT  147.11 92.52 147.65 91.97 ;
      RECT  145.97 93.24 147.11 93.62 ;
      RECT  148.37 93.0 148.58 93.07 ;
      RECT  148.58 93.86 149.09 94.1 ;
      RECT  146.18 92.76 148.58 93.0 ;
      RECT  148.58 93.0 148.78 93.07 ;
      RECT  148.37 93.79 148.58 93.86 ;
      RECT  149.09 92.76 149.3 93.0 ;
      POLYGON  147.65 93.24 147.65 93.62 148.2 93.62 148.2 93.55 148.58 93.55 148.58 93.31 148.2 93.31 148.2 93.24 147.65 93.24 ;
      RECT  149.09 93.24 149.3 93.62 ;
      RECT  145.97 91.97 146.18 92.52 ;
      RECT  146.18 91.97 147.11 92.52 ;
      RECT  147.11 93.24 147.65 93.62 ;
      RECT  149.09 93.86 149.3 94.1 ;
      RECT  147.65 91.97 149.3 92.52 ;
      RECT  145.97 92.76 146.18 93.0 ;
      RECT  148.58 93.79 148.78 93.86 ;
      POLYGON  148.95 93.24 148.95 93.31 148.58 93.31 148.58 93.55 148.95 93.55 148.95 93.62 149.09 93.62 149.09 93.24 148.95 93.24 ;
      RECT  145.97 93.86 146.18 94.1 ;
      RECT  146.18 93.86 148.58 94.1 ;
      RECT  148.58 92.76 149.09 93.0 ;
      RECT  147.11 91.97 147.65 92.52 ;
      RECT  145.97 95.2 147.11 94.82 ;
      RECT  148.37 95.44 148.58 95.37 ;
      RECT  148.58 94.58 149.09 94.34 ;
      RECT  146.18 95.68 148.58 95.44 ;
      RECT  148.58 95.44 148.78 95.37 ;
      RECT  148.37 94.65 148.58 94.58 ;
      RECT  149.09 95.68 149.3 95.44 ;
      POLYGON  147.65 95.2 147.65 94.82 148.2 94.82 148.2 94.89 148.58 94.89 148.58 95.13 148.2 95.13 148.2 95.2 147.65 95.2 ;
      RECT  149.09 95.2 149.3 94.82 ;
      RECT  145.97 96.47 146.18 95.92 ;
      RECT  146.18 96.47 147.11 95.92 ;
      RECT  147.11 95.2 147.65 94.82 ;
      RECT  149.09 94.58 149.3 94.34 ;
      RECT  147.65 96.47 149.3 95.92 ;
      RECT  145.97 95.68 146.18 95.44 ;
      RECT  148.58 94.65 148.78 94.58 ;
      POLYGON  148.95 95.2 148.95 95.13 148.58 95.13 148.58 94.89 148.95 94.89 148.95 94.82 149.09 94.82 149.09 95.2 148.95 95.2 ;
      RECT  145.97 94.58 146.18 94.34 ;
      RECT  146.18 94.58 148.58 94.34 ;
      RECT  148.58 95.68 149.09 95.44 ;
      RECT  147.11 96.47 147.65 95.92 ;
      RECT  145.97 97.19 147.11 97.57 ;
      RECT  148.37 96.95 148.58 97.02 ;
      RECT  148.58 97.81 149.09 98.05 ;
      RECT  146.18 96.71 148.58 96.95 ;
      RECT  148.58 96.95 148.78 97.02 ;
      RECT  148.37 97.74 148.58 97.81 ;
      RECT  149.09 96.71 149.3 96.95 ;
      POLYGON  147.65 97.19 147.65 97.57 148.2 97.57 148.2 97.5 148.58 97.5 148.58 97.26 148.2 97.26 148.2 97.19 147.65 97.19 ;
      RECT  149.09 97.19 149.3 97.57 ;
      RECT  145.97 95.92 146.18 96.47 ;
      RECT  146.18 95.92 147.11 96.47 ;
      RECT  147.11 97.19 147.65 97.57 ;
      RECT  149.09 97.81 149.3 98.05 ;
      RECT  147.65 95.92 149.3 96.47 ;
      RECT  145.97 96.71 146.18 96.95 ;
      RECT  148.58 97.74 148.78 97.81 ;
      POLYGON  148.95 97.19 148.95 97.26 148.58 97.26 148.58 97.5 148.95 97.5 148.95 97.57 149.09 97.57 149.09 97.19 148.95 97.19 ;
      RECT  145.97 97.81 146.18 98.05 ;
      RECT  146.18 97.81 148.58 98.05 ;
      RECT  148.58 96.71 149.09 96.95 ;
      RECT  147.11 95.92 147.65 96.47 ;
      RECT  145.97 99.15 147.11 98.77 ;
      RECT  148.37 99.39 148.58 99.32 ;
      RECT  148.58 98.53 149.09 98.29 ;
      RECT  146.18 99.63 148.58 99.39 ;
      RECT  148.58 99.39 148.78 99.32 ;
      RECT  148.37 98.6 148.58 98.53 ;
      RECT  149.09 99.63 149.3 99.39 ;
      POLYGON  147.65 99.15 147.65 98.77 148.2 98.77 148.2 98.84 148.58 98.84 148.58 99.08 148.2 99.08 148.2 99.15 147.65 99.15 ;
      RECT  149.09 99.15 149.3 98.77 ;
      RECT  145.97 100.42 146.18 99.87 ;
      RECT  146.18 100.42 147.11 99.87 ;
      RECT  147.11 99.15 147.65 98.77 ;
      RECT  149.09 98.53 149.3 98.29 ;
      RECT  147.65 100.42 149.3 99.87 ;
      RECT  145.97 99.63 146.18 99.39 ;
      RECT  148.58 98.6 148.78 98.53 ;
      POLYGON  148.95 99.15 148.95 99.08 148.58 99.08 148.58 98.84 148.95 98.84 148.95 98.77 149.09 98.77 149.09 99.15 148.95 99.15 ;
      RECT  145.97 98.53 146.18 98.29 ;
      RECT  146.18 98.53 148.58 98.29 ;
      RECT  148.58 99.63 149.09 99.39 ;
      RECT  147.11 100.42 147.65 99.87 ;
      RECT  145.97 101.14 147.11 101.52 ;
      RECT  148.37 100.9 148.58 100.97 ;
      RECT  148.58 101.76 149.09 102.0 ;
      RECT  146.18 100.66 148.58 100.9 ;
      RECT  148.58 100.9 148.78 100.97 ;
      RECT  148.37 101.69 148.58 101.76 ;
      RECT  149.09 100.66 149.3 100.9 ;
      POLYGON  147.65 101.14 147.65 101.52 148.2 101.52 148.2 101.45 148.58 101.45 148.58 101.21 148.2 101.21 148.2 101.14 147.65 101.14 ;
      RECT  149.09 101.14 149.3 101.52 ;
      RECT  145.97 99.87 146.18 100.42 ;
      RECT  146.18 99.87 147.11 100.42 ;
      RECT  147.11 101.14 147.65 101.52 ;
      RECT  149.09 101.76 149.3 102.0 ;
      RECT  147.65 99.87 149.3 100.42 ;
      RECT  145.97 100.66 146.18 100.9 ;
      RECT  148.58 101.69 148.78 101.76 ;
      POLYGON  148.95 101.14 148.95 101.21 148.58 101.21 148.58 101.45 148.95 101.45 148.95 101.52 149.09 101.52 149.09 101.14 148.95 101.14 ;
      RECT  145.97 101.76 146.18 102.0 ;
      RECT  146.18 101.76 148.58 102.0 ;
      RECT  148.58 100.66 149.09 100.9 ;
      RECT  147.11 99.87 147.65 100.42 ;
      RECT  145.97 103.1 147.11 102.72 ;
      RECT  148.37 103.34 148.58 103.27 ;
      RECT  148.58 102.48 149.09 102.24 ;
      RECT  146.18 103.58 148.58 103.34 ;
      RECT  148.58 103.34 148.78 103.27 ;
      RECT  148.37 102.55 148.58 102.48 ;
      RECT  149.09 103.58 149.3 103.34 ;
      POLYGON  147.65 103.1 147.65 102.72 148.2 102.72 148.2 102.79 148.58 102.79 148.58 103.03 148.2 103.03 148.2 103.1 147.65 103.1 ;
      RECT  149.09 103.1 149.3 102.72 ;
      RECT  145.97 104.37 146.18 103.82 ;
      RECT  146.18 104.37 147.11 103.82 ;
      RECT  147.11 103.1 147.65 102.72 ;
      RECT  149.09 102.48 149.3 102.24 ;
      RECT  147.65 104.37 149.3 103.82 ;
      RECT  145.97 103.58 146.18 103.34 ;
      RECT  148.58 102.55 148.78 102.48 ;
      POLYGON  148.95 103.1 148.95 103.03 148.58 103.03 148.58 102.79 148.95 102.79 148.95 102.72 149.09 102.72 149.09 103.1 148.95 103.1 ;
      RECT  145.97 102.48 146.18 102.24 ;
      RECT  146.18 102.48 148.58 102.24 ;
      RECT  148.58 103.58 149.09 103.34 ;
      RECT  147.11 104.37 147.65 103.82 ;
      RECT  145.97 105.09 147.11 105.47 ;
      RECT  148.37 104.85 148.58 104.92 ;
      RECT  148.58 105.71 149.09 105.95 ;
      RECT  146.18 104.61 148.58 104.85 ;
      RECT  148.58 104.85 148.78 104.92 ;
      RECT  148.37 105.64 148.58 105.71 ;
      RECT  149.09 104.61 149.3 104.85 ;
      POLYGON  147.65 105.09 147.65 105.47 148.2 105.47 148.2 105.4 148.58 105.4 148.58 105.16 148.2 105.16 148.2 105.09 147.65 105.09 ;
      RECT  149.09 105.09 149.3 105.47 ;
      RECT  145.97 103.82 146.18 104.37 ;
      RECT  146.18 103.82 147.11 104.37 ;
      RECT  147.11 105.09 147.65 105.47 ;
      RECT  149.09 105.71 149.3 105.95 ;
      RECT  147.65 103.82 149.3 104.37 ;
      RECT  145.97 104.61 146.18 104.85 ;
      RECT  148.58 105.64 148.78 105.71 ;
      POLYGON  148.95 105.09 148.95 105.16 148.58 105.16 148.58 105.4 148.95 105.4 148.95 105.47 149.09 105.47 149.09 105.09 148.95 105.09 ;
      RECT  145.97 105.71 146.18 105.95 ;
      RECT  146.18 105.71 148.58 105.95 ;
      RECT  148.58 104.61 149.09 104.85 ;
      RECT  147.11 103.82 147.65 104.37 ;
      RECT  145.97 107.05 147.11 106.67 ;
      RECT  148.37 107.29 148.58 107.22 ;
      RECT  148.58 106.43 149.09 106.19 ;
      RECT  146.18 107.53 148.58 107.29 ;
      RECT  148.58 107.29 148.78 107.22 ;
      RECT  148.37 106.5 148.58 106.43 ;
      RECT  149.09 107.53 149.3 107.29 ;
      POLYGON  147.65 107.05 147.65 106.67 148.2 106.67 148.2 106.74 148.58 106.74 148.58 106.98 148.2 106.98 148.2 107.05 147.65 107.05 ;
      RECT  149.09 107.05 149.3 106.67 ;
      RECT  145.97 108.32 146.18 107.77 ;
      RECT  146.18 108.32 147.11 107.77 ;
      RECT  147.11 107.05 147.65 106.67 ;
      RECT  149.09 106.43 149.3 106.19 ;
      RECT  147.65 108.32 149.3 107.77 ;
      RECT  145.97 107.53 146.18 107.29 ;
      RECT  148.58 106.5 148.78 106.43 ;
      POLYGON  148.95 107.05 148.95 106.98 148.58 106.98 148.58 106.74 148.95 106.74 148.95 106.67 149.09 106.67 149.09 107.05 148.95 107.05 ;
      RECT  145.97 106.43 146.18 106.19 ;
      RECT  146.18 106.43 148.58 106.19 ;
      RECT  148.58 107.53 149.09 107.29 ;
      RECT  147.11 108.32 147.65 107.77 ;
      RECT  145.97 109.04 147.11 109.42 ;
      RECT  148.37 108.8 148.58 108.87 ;
      RECT  148.58 109.66 149.09 109.9 ;
      RECT  146.18 108.56 148.58 108.8 ;
      RECT  148.58 108.8 148.78 108.87 ;
      RECT  148.37 109.59 148.58 109.66 ;
      RECT  149.09 108.56 149.3 108.8 ;
      POLYGON  147.65 109.04 147.65 109.42 148.2 109.42 148.2 109.35 148.58 109.35 148.58 109.11 148.2 109.11 148.2 109.04 147.65 109.04 ;
      RECT  149.09 109.04 149.3 109.42 ;
      RECT  145.97 107.77 146.18 108.32 ;
      RECT  146.18 107.77 147.11 108.32 ;
      RECT  147.11 109.04 147.65 109.42 ;
      RECT  149.09 109.66 149.3 109.9 ;
      RECT  147.65 107.77 149.3 108.32 ;
      RECT  145.97 108.56 146.18 108.8 ;
      RECT  148.58 109.59 148.78 109.66 ;
      POLYGON  148.95 109.04 148.95 109.11 148.58 109.11 148.58 109.35 148.95 109.35 148.95 109.42 149.09 109.42 149.09 109.04 148.95 109.04 ;
      RECT  145.97 109.66 146.18 109.9 ;
      RECT  146.18 109.66 148.58 109.9 ;
      RECT  148.58 108.56 149.09 108.8 ;
      RECT  147.11 107.77 147.65 108.32 ;
      RECT  145.97 111.0 147.11 110.62 ;
      RECT  148.37 111.24 148.58 111.17 ;
      RECT  148.58 110.38 149.09 110.14 ;
      RECT  146.18 111.48 148.58 111.24 ;
      RECT  148.58 111.24 148.78 111.17 ;
      RECT  148.37 110.45 148.58 110.38 ;
      RECT  149.09 111.48 149.3 111.24 ;
      POLYGON  147.65 111.0 147.65 110.62 148.2 110.62 148.2 110.69 148.58 110.69 148.58 110.93 148.2 110.93 148.2 111.0 147.65 111.0 ;
      RECT  149.09 111.0 149.3 110.62 ;
      RECT  145.97 112.27 146.18 111.72 ;
      RECT  146.18 112.27 147.11 111.72 ;
      RECT  147.11 111.0 147.65 110.62 ;
      RECT  149.09 110.38 149.3 110.14 ;
      RECT  147.65 112.27 149.3 111.72 ;
      RECT  145.97 111.48 146.18 111.24 ;
      RECT  148.58 110.45 148.78 110.38 ;
      POLYGON  148.95 111.0 148.95 110.93 148.58 110.93 148.58 110.69 148.95 110.69 148.95 110.62 149.09 110.62 149.09 111.0 148.95 111.0 ;
      RECT  145.97 110.38 146.18 110.14 ;
      RECT  146.18 110.38 148.58 110.14 ;
      RECT  148.58 111.48 149.09 111.24 ;
      RECT  147.11 112.27 147.65 111.72 ;
      RECT  145.97 112.99 147.11 113.37 ;
      RECT  148.37 112.75 148.58 112.82 ;
      RECT  148.58 113.61 149.09 113.85 ;
      RECT  146.18 112.51 148.58 112.75 ;
      RECT  148.58 112.75 148.78 112.82 ;
      RECT  148.37 113.54 148.58 113.61 ;
      RECT  149.09 112.51 149.3 112.75 ;
      POLYGON  147.65 112.99 147.65 113.37 148.2 113.37 148.2 113.3 148.58 113.3 148.58 113.06 148.2 113.06 148.2 112.99 147.65 112.99 ;
      RECT  149.09 112.99 149.3 113.37 ;
      RECT  145.97 111.72 146.18 112.27 ;
      RECT  146.18 111.72 147.11 112.27 ;
      RECT  147.11 112.99 147.65 113.37 ;
      RECT  149.09 113.61 149.3 113.85 ;
      RECT  147.65 111.72 149.3 112.27 ;
      RECT  145.97 112.51 146.18 112.75 ;
      RECT  148.58 113.54 148.78 113.61 ;
      POLYGON  148.95 112.99 148.95 113.06 148.58 113.06 148.58 113.3 148.95 113.3 148.95 113.37 149.09 113.37 149.09 112.99 148.95 112.99 ;
      RECT  145.97 113.61 146.18 113.85 ;
      RECT  146.18 113.61 148.58 113.85 ;
      RECT  148.58 112.51 149.09 112.75 ;
      RECT  147.11 111.72 147.65 112.27 ;
      RECT  145.97 114.95 147.11 114.57 ;
      RECT  148.37 115.19 148.58 115.12 ;
      RECT  148.58 114.33 149.09 114.09 ;
      RECT  146.18 115.43 148.58 115.19 ;
      RECT  148.58 115.19 148.78 115.12 ;
      RECT  148.37 114.4 148.58 114.33 ;
      RECT  149.09 115.43 149.3 115.19 ;
      POLYGON  147.65 114.95 147.65 114.57 148.2 114.57 148.2 114.64 148.58 114.64 148.58 114.88 148.2 114.88 148.2 114.95 147.65 114.95 ;
      RECT  149.09 114.95 149.3 114.57 ;
      RECT  145.97 116.22 146.18 115.67 ;
      RECT  146.18 116.22 147.11 115.67 ;
      RECT  147.11 114.95 147.65 114.57 ;
      RECT  149.09 114.33 149.3 114.09 ;
      RECT  147.65 116.22 149.3 115.67 ;
      RECT  145.97 115.43 146.18 115.19 ;
      RECT  148.58 114.4 148.78 114.33 ;
      POLYGON  148.95 114.95 148.95 114.88 148.58 114.88 148.58 114.64 148.95 114.64 148.95 114.57 149.09 114.57 149.09 114.95 148.95 114.95 ;
      RECT  145.97 114.33 146.18 114.09 ;
      RECT  146.18 114.33 148.58 114.09 ;
      RECT  148.58 115.43 149.09 115.19 ;
      RECT  147.11 116.22 147.65 115.67 ;
      RECT  145.97 116.94 147.11 117.32 ;
      RECT  148.37 116.7 148.58 116.77 ;
      RECT  148.58 117.56 149.09 117.8 ;
      RECT  146.18 116.46 148.58 116.7 ;
      RECT  148.58 116.7 148.78 116.77 ;
      RECT  148.37 117.49 148.58 117.56 ;
      RECT  149.09 116.46 149.3 116.7 ;
      POLYGON  147.65 116.94 147.65 117.32 148.2 117.32 148.2 117.25 148.58 117.25 148.58 117.01 148.2 117.01 148.2 116.94 147.65 116.94 ;
      RECT  149.09 116.94 149.3 117.32 ;
      RECT  145.97 115.67 146.18 116.22 ;
      RECT  146.18 115.67 147.11 116.22 ;
      RECT  147.11 116.94 147.65 117.32 ;
      RECT  149.09 117.56 149.3 117.8 ;
      RECT  147.65 115.67 149.3 116.22 ;
      RECT  145.97 116.46 146.18 116.7 ;
      RECT  148.58 117.49 148.78 117.56 ;
      POLYGON  148.95 116.94 148.95 117.01 148.58 117.01 148.58 117.25 148.95 117.25 148.95 117.32 149.09 117.32 149.09 116.94 148.95 116.94 ;
      RECT  145.97 117.56 146.18 117.8 ;
      RECT  146.18 117.56 148.58 117.8 ;
      RECT  148.58 116.46 149.09 116.7 ;
      RECT  147.11 115.67 147.65 116.22 ;
      RECT  145.97 118.9 147.11 118.52 ;
      RECT  148.37 119.14 148.58 119.07 ;
      RECT  148.58 118.28 149.09 118.04 ;
      RECT  146.18 119.38 148.58 119.14 ;
      RECT  148.58 119.14 148.78 119.07 ;
      RECT  148.37 118.35 148.58 118.28 ;
      RECT  149.09 119.38 149.3 119.14 ;
      POLYGON  147.65 118.9 147.65 118.52 148.2 118.52 148.2 118.59 148.58 118.59 148.58 118.83 148.2 118.83 148.2 118.9 147.65 118.9 ;
      RECT  149.09 118.9 149.3 118.52 ;
      RECT  145.97 120.17 146.18 119.62 ;
      RECT  146.18 120.17 147.11 119.62 ;
      RECT  147.11 118.9 147.65 118.52 ;
      RECT  149.09 118.28 149.3 118.04 ;
      RECT  147.65 120.17 149.3 119.62 ;
      RECT  145.97 119.38 146.18 119.14 ;
      RECT  148.58 118.35 148.78 118.28 ;
      POLYGON  148.95 118.9 148.95 118.83 148.58 118.83 148.58 118.59 148.95 118.59 148.95 118.52 149.09 118.52 149.09 118.9 148.95 118.9 ;
      RECT  145.97 118.28 146.18 118.04 ;
      RECT  146.18 118.28 148.58 118.04 ;
      RECT  148.58 119.38 149.09 119.14 ;
      RECT  147.11 120.17 147.65 119.62 ;
      RECT  145.97 120.89 147.11 121.27 ;
      RECT  148.37 120.65 148.58 120.72 ;
      RECT  148.58 121.51 149.09 121.75 ;
      RECT  146.18 120.41 148.58 120.65 ;
      RECT  148.58 120.65 148.78 120.72 ;
      RECT  148.37 121.44 148.58 121.51 ;
      RECT  149.09 120.41 149.3 120.65 ;
      POLYGON  147.65 120.89 147.65 121.27 148.2 121.27 148.2 121.2 148.58 121.2 148.58 120.96 148.2 120.96 148.2 120.89 147.65 120.89 ;
      RECT  149.09 120.89 149.3 121.27 ;
      RECT  145.97 119.62 146.18 120.17 ;
      RECT  146.18 119.62 147.11 120.17 ;
      RECT  147.11 120.89 147.65 121.27 ;
      RECT  149.09 121.51 149.3 121.75 ;
      RECT  147.65 119.62 149.3 120.17 ;
      RECT  145.97 120.41 146.18 120.65 ;
      RECT  148.58 121.44 148.78 121.51 ;
      POLYGON  148.95 120.89 148.95 120.96 148.58 120.96 148.58 121.2 148.95 121.2 148.95 121.27 149.09 121.27 149.09 120.89 148.95 120.89 ;
      RECT  145.97 121.51 146.18 121.75 ;
      RECT  146.18 121.51 148.58 121.75 ;
      RECT  148.58 120.41 149.09 120.65 ;
      RECT  147.11 119.62 147.65 120.17 ;
      RECT  145.97 122.85 147.11 122.47 ;
      RECT  148.37 123.09 148.58 123.02 ;
      RECT  148.58 122.23 149.09 121.99 ;
      RECT  146.18 123.33 148.58 123.09 ;
      RECT  148.58 123.09 148.78 123.02 ;
      RECT  148.37 122.3 148.58 122.23 ;
      RECT  149.09 123.33 149.3 123.09 ;
      POLYGON  147.65 122.85 147.65 122.47 148.2 122.47 148.2 122.54 148.58 122.54 148.58 122.78 148.2 122.78 148.2 122.85 147.65 122.85 ;
      RECT  149.09 122.85 149.3 122.47 ;
      RECT  145.97 124.12 146.18 123.57 ;
      RECT  146.18 124.12 147.11 123.57 ;
      RECT  147.11 122.85 147.65 122.47 ;
      RECT  149.09 122.23 149.3 121.99 ;
      RECT  147.65 124.12 149.3 123.57 ;
      RECT  145.97 123.33 146.18 123.09 ;
      RECT  148.58 122.3 148.78 122.23 ;
      POLYGON  148.95 122.85 148.95 122.78 148.58 122.78 148.58 122.54 148.95 122.54 148.95 122.47 149.09 122.47 149.09 122.85 148.95 122.85 ;
      RECT  145.97 122.23 146.18 121.99 ;
      RECT  146.18 122.23 148.58 121.99 ;
      RECT  148.58 123.33 149.09 123.09 ;
      RECT  147.11 124.12 147.65 123.57 ;
      RECT  145.97 124.84 147.11 125.22 ;
      RECT  148.37 124.6 148.58 124.67 ;
      RECT  148.58 125.46 149.09 125.7 ;
      RECT  146.18 124.36 148.58 124.6 ;
      RECT  148.58 124.6 148.78 124.67 ;
      RECT  148.37 125.39 148.58 125.46 ;
      RECT  149.09 124.36 149.3 124.6 ;
      POLYGON  147.65 124.84 147.65 125.22 148.2 125.22 148.2 125.15 148.58 125.15 148.58 124.91 148.2 124.91 148.2 124.84 147.65 124.84 ;
      RECT  149.09 124.84 149.3 125.22 ;
      RECT  145.97 123.57 146.18 124.12 ;
      RECT  146.18 123.57 147.11 124.12 ;
      RECT  147.11 124.84 147.65 125.22 ;
      RECT  149.09 125.46 149.3 125.7 ;
      RECT  147.65 123.57 149.3 124.12 ;
      RECT  145.97 124.36 146.18 124.6 ;
      RECT  148.58 125.39 148.78 125.46 ;
      POLYGON  148.95 124.84 148.95 124.91 148.58 124.91 148.58 125.15 148.95 125.15 148.95 125.22 149.09 125.22 149.09 124.84 148.95 124.84 ;
      RECT  145.97 125.46 146.18 125.7 ;
      RECT  146.18 125.46 148.58 125.7 ;
      RECT  148.58 124.36 149.09 124.6 ;
      RECT  147.11 123.57 147.65 124.12 ;
      RECT  146.18 126.925 149.3 126.375 ;
      RECT  146.18 90.39 149.3 90.63 ;
      RECT  146.18 91.49 149.3 91.73 ;
      RECT  146.18 93.86 149.3 94.1 ;
      RECT  146.18 92.76 149.3 93.0 ;
      RECT  146.18 94.34 149.3 94.58 ;
      RECT  146.18 95.44 149.3 95.68 ;
      RECT  146.18 97.81 149.3 98.05 ;
      RECT  146.18 96.71 149.3 96.95 ;
      RECT  146.18 98.29 149.3 98.53 ;
      RECT  146.18 99.39 149.3 99.63 ;
      RECT  146.18 101.76 149.3 102.0 ;
      RECT  146.18 100.66 149.3 100.9 ;
      RECT  146.18 102.24 149.3 102.48 ;
      RECT  146.18 103.34 149.3 103.58 ;
      RECT  146.18 105.71 149.3 105.95 ;
      RECT  146.18 104.61 149.3 104.85 ;
      RECT  146.18 106.19 149.3 106.43 ;
      RECT  146.18 107.29 149.3 107.53 ;
      RECT  146.18 109.66 149.3 109.9 ;
      RECT  146.18 108.56 149.3 108.8 ;
      RECT  146.18 110.14 149.3 110.38 ;
      RECT  146.18 111.24 149.3 111.48 ;
      RECT  146.18 113.61 149.3 113.85 ;
      RECT  146.18 112.51 149.3 112.75 ;
      RECT  146.18 114.09 149.3 114.33 ;
      RECT  146.18 115.19 149.3 115.43 ;
      RECT  146.18 117.56 149.3 117.8 ;
      RECT  146.18 116.46 149.3 116.7 ;
      RECT  146.18 118.04 149.3 118.28 ;
      RECT  146.18 119.14 149.3 119.38 ;
      RECT  146.18 121.51 149.3 121.75 ;
      RECT  146.18 120.41 149.3 120.65 ;
      RECT  146.18 121.99 149.3 122.23 ;
      RECT  146.18 123.09 149.3 123.33 ;
      RECT  146.18 125.46 149.3 125.7 ;
      RECT  146.18 124.36 149.3 124.6 ;
      RECT  147.11 90.87 147.65 91.25 ;
      RECT  147.11 91.97 147.65 92.52 ;
      RECT  147.11 97.19 147.65 97.57 ;
      RECT  147.11 115.67 147.65 116.22 ;
      RECT  147.11 123.57 147.65 124.12 ;
      RECT  147.11 98.77 147.65 99.15 ;
      RECT  147.11 119.62 147.65 120.17 ;
      RECT  147.11 101.14 147.65 101.52 ;
      RECT  147.11 105.09 147.65 105.47 ;
      RECT  147.11 118.52 147.65 118.9 ;
      RECT  147.11 124.84 147.65 125.22 ;
      RECT  147.11 110.62 147.65 111.0 ;
      RECT  147.11 111.72 147.65 112.27 ;
      RECT  147.11 122.47 147.65 122.85 ;
      RECT  147.11 120.89 147.65 121.27 ;
      RECT  147.11 112.99 147.65 113.37 ;
      RECT  147.11 109.04 147.65 109.42 ;
      RECT  147.11 95.92 147.65 96.47 ;
      RECT  147.11 116.94 147.65 117.32 ;
      RECT  147.11 107.77 147.65 108.32 ;
      RECT  147.11 94.82 147.65 95.2 ;
      RECT  147.11 99.87 147.65 100.42 ;
      RECT  147.11 102.72 147.65 103.1 ;
      RECT  147.11 103.82 147.65 104.37 ;
      RECT  147.11 106.67 147.65 107.05 ;
      RECT  147.11 93.24 147.65 93.62 ;
      RECT  147.11 114.57 147.65 114.95 ;
      RECT  96.05 91.25 97.19 90.87 ;
      RECT  98.45 91.49 98.66 91.42 ;
      RECT  98.66 90.63 99.17 90.39 ;
      RECT  96.26 91.73 98.66 91.49 ;
      RECT  98.66 91.49 98.86 91.42 ;
      RECT  98.45 90.7 98.66 90.63 ;
      RECT  99.17 91.73 99.38 91.49 ;
      POLYGON  97.73 91.25 97.73 90.87 98.28 90.87 98.28 90.94 98.66 90.94 98.66 91.18 98.28 91.18 98.28 91.25 97.73 91.25 ;
      RECT  99.17 91.25 99.38 90.87 ;
      RECT  96.05 92.52 96.26 91.97 ;
      RECT  96.26 92.52 97.19 91.97 ;
      RECT  97.19 91.25 97.73 90.87 ;
      RECT  99.17 90.63 99.38 90.39 ;
      RECT  97.73 92.52 99.38 91.97 ;
      RECT  96.05 91.73 96.26 91.49 ;
      RECT  98.66 90.7 98.86 90.63 ;
      POLYGON  99.03 91.25 99.03 91.18 98.66 91.18 98.66 90.94 99.03 90.94 99.03 90.87 99.17 90.87 99.17 91.25 99.03 91.25 ;
      RECT  96.05 90.63 96.26 90.39 ;
      RECT  96.26 90.63 98.66 90.39 ;
      RECT  98.66 91.73 99.17 91.49 ;
      RECT  97.19 92.52 97.73 91.97 ;
      RECT  102.71 91.25 101.57 90.87 ;
      RECT  100.31 91.49 100.1 91.42 ;
      RECT  100.1 90.63 99.59 90.39 ;
      RECT  102.5 91.73 100.1 91.49 ;
      RECT  100.1 91.49 99.9 91.42 ;
      RECT  100.31 90.7 100.1 90.63 ;
      RECT  99.59 91.73 99.38 91.49 ;
      POLYGON  101.03 91.25 101.03 90.87 100.48 90.87 100.48 90.94 100.1 90.94 100.1 91.18 100.48 91.18 100.48 91.25 101.03 91.25 ;
      RECT  99.59 91.25 99.38 90.87 ;
      RECT  102.71 92.52 102.5 91.97 ;
      RECT  102.5 92.52 101.57 91.97 ;
      RECT  101.57 91.25 101.03 90.87 ;
      RECT  99.59 90.63 99.38 90.39 ;
      RECT  101.03 92.52 99.38 91.97 ;
      RECT  102.71 91.73 102.5 91.49 ;
      RECT  100.1 90.7 99.9 90.63 ;
      POLYGON  99.73 91.25 99.73 91.18 100.1 91.18 100.1 90.94 99.73 90.94 99.73 90.87 99.59 90.87 99.59 91.25 99.73 91.25 ;
      RECT  102.71 90.63 102.5 90.39 ;
      RECT  102.5 90.63 100.1 90.39 ;
      RECT  100.1 91.73 99.59 91.49 ;
      RECT  101.57 92.52 101.03 91.97 ;
      RECT  102.29 91.25 103.43 90.87 ;
      RECT  104.69 91.49 104.9 91.42 ;
      RECT  104.9 90.63 105.41 90.39 ;
      RECT  102.5 91.73 104.9 91.49 ;
      RECT  104.9 91.49 105.1 91.42 ;
      RECT  104.69 90.7 104.9 90.63 ;
      RECT  105.41 91.73 105.62 91.49 ;
      POLYGON  103.97 91.25 103.97 90.87 104.52 90.87 104.52 90.94 104.9 90.94 104.9 91.18 104.52 91.18 104.52 91.25 103.97 91.25 ;
      RECT  105.41 91.25 105.62 90.87 ;
      RECT  102.29 92.52 102.5 91.97 ;
      RECT  102.5 92.52 103.43 91.97 ;
      RECT  103.43 91.25 103.97 90.87 ;
      RECT  105.41 90.63 105.62 90.39 ;
      RECT  103.97 92.52 105.62 91.97 ;
      RECT  102.29 91.73 102.5 91.49 ;
      RECT  104.9 90.7 105.1 90.63 ;
      POLYGON  105.27 91.25 105.27 91.18 104.9 91.18 104.9 90.94 105.27 90.94 105.27 90.87 105.41 90.87 105.41 91.25 105.27 91.25 ;
      RECT  102.29 90.63 102.5 90.39 ;
      RECT  102.5 90.63 104.9 90.39 ;
      RECT  104.9 91.73 105.41 91.49 ;
      RECT  103.43 92.52 103.97 91.97 ;
      RECT  108.95 91.25 107.81 90.87 ;
      RECT  106.55 91.49 106.34 91.42 ;
      RECT  106.34 90.63 105.83 90.39 ;
      RECT  108.74 91.73 106.34 91.49 ;
      RECT  106.34 91.49 106.14 91.42 ;
      RECT  106.55 90.7 106.34 90.63 ;
      RECT  105.83 91.73 105.62 91.49 ;
      POLYGON  107.27 91.25 107.27 90.87 106.72 90.87 106.72 90.94 106.34 90.94 106.34 91.18 106.72 91.18 106.72 91.25 107.27 91.25 ;
      RECT  105.83 91.25 105.62 90.87 ;
      RECT  108.95 92.52 108.74 91.97 ;
      RECT  108.74 92.52 107.81 91.97 ;
      RECT  107.81 91.25 107.27 90.87 ;
      RECT  105.83 90.63 105.62 90.39 ;
      RECT  107.27 92.52 105.62 91.97 ;
      RECT  108.95 91.73 108.74 91.49 ;
      RECT  106.34 90.7 106.14 90.63 ;
      POLYGON  105.97 91.25 105.97 91.18 106.34 91.18 106.34 90.94 105.97 90.94 105.97 90.87 105.83 90.87 105.83 91.25 105.97 91.25 ;
      RECT  108.95 90.63 108.74 90.39 ;
      RECT  108.74 90.63 106.34 90.39 ;
      RECT  106.34 91.73 105.83 91.49 ;
      RECT  107.81 92.52 107.27 91.97 ;
      RECT  108.53 91.25 109.67 90.87 ;
      RECT  110.93 91.49 111.14 91.42 ;
      RECT  111.14 90.63 111.65 90.39 ;
      RECT  108.74 91.73 111.14 91.49 ;
      RECT  111.14 91.49 111.34 91.42 ;
      RECT  110.93 90.7 111.14 90.63 ;
      RECT  111.65 91.73 111.86 91.49 ;
      POLYGON  110.21 91.25 110.21 90.87 110.76 90.87 110.76 90.94 111.14 90.94 111.14 91.18 110.76 91.18 110.76 91.25 110.21 91.25 ;
      RECT  111.65 91.25 111.86 90.87 ;
      RECT  108.53 92.52 108.74 91.97 ;
      RECT  108.74 92.52 109.67 91.97 ;
      RECT  109.67 91.25 110.21 90.87 ;
      RECT  111.65 90.63 111.86 90.39 ;
      RECT  110.21 92.52 111.86 91.97 ;
      RECT  108.53 91.73 108.74 91.49 ;
      RECT  111.14 90.7 111.34 90.63 ;
      POLYGON  111.51 91.25 111.51 91.18 111.14 91.18 111.14 90.94 111.51 90.94 111.51 90.87 111.65 90.87 111.65 91.25 111.51 91.25 ;
      RECT  108.53 90.63 108.74 90.39 ;
      RECT  108.74 90.63 111.14 90.39 ;
      RECT  111.14 91.73 111.65 91.49 ;
      RECT  109.67 92.52 110.21 91.97 ;
      RECT  115.19 91.25 114.05 90.87 ;
      RECT  112.79 91.49 112.58 91.42 ;
      RECT  112.58 90.63 112.07 90.39 ;
      RECT  114.98 91.73 112.58 91.49 ;
      RECT  112.58 91.49 112.38 91.42 ;
      RECT  112.79 90.7 112.58 90.63 ;
      RECT  112.07 91.73 111.86 91.49 ;
      POLYGON  113.51 91.25 113.51 90.87 112.96 90.87 112.96 90.94 112.58 90.94 112.58 91.18 112.96 91.18 112.96 91.25 113.51 91.25 ;
      RECT  112.07 91.25 111.86 90.87 ;
      RECT  115.19 92.52 114.98 91.97 ;
      RECT  114.98 92.52 114.05 91.97 ;
      RECT  114.05 91.25 113.51 90.87 ;
      RECT  112.07 90.63 111.86 90.39 ;
      RECT  113.51 92.52 111.86 91.97 ;
      RECT  115.19 91.73 114.98 91.49 ;
      RECT  112.58 90.7 112.38 90.63 ;
      POLYGON  112.21 91.25 112.21 91.18 112.58 91.18 112.58 90.94 112.21 90.94 112.21 90.87 112.07 90.87 112.07 91.25 112.21 91.25 ;
      RECT  115.19 90.63 114.98 90.39 ;
      RECT  114.98 90.63 112.58 90.39 ;
      RECT  112.58 91.73 112.07 91.49 ;
      RECT  114.05 92.52 113.51 91.97 ;
      RECT  114.77 91.25 115.91 90.87 ;
      RECT  117.17 91.49 117.38 91.42 ;
      RECT  117.38 90.63 117.89 90.39 ;
      RECT  114.98 91.73 117.38 91.49 ;
      RECT  117.38 91.49 117.58 91.42 ;
      RECT  117.17 90.7 117.38 90.63 ;
      RECT  117.89 91.73 118.1 91.49 ;
      POLYGON  116.45 91.25 116.45 90.87 117.0 90.87 117.0 90.94 117.38 90.94 117.38 91.18 117.0 91.18 117.0 91.25 116.45 91.25 ;
      RECT  117.89 91.25 118.1 90.87 ;
      RECT  114.77 92.52 114.98 91.97 ;
      RECT  114.98 92.52 115.91 91.97 ;
      RECT  115.91 91.25 116.45 90.87 ;
      RECT  117.89 90.63 118.1 90.39 ;
      RECT  116.45 92.52 118.1 91.97 ;
      RECT  114.77 91.73 114.98 91.49 ;
      RECT  117.38 90.7 117.58 90.63 ;
      POLYGON  117.75 91.25 117.75 91.18 117.38 91.18 117.38 90.94 117.75 90.94 117.75 90.87 117.89 90.87 117.89 91.25 117.75 91.25 ;
      RECT  114.77 90.63 114.98 90.39 ;
      RECT  114.98 90.63 117.38 90.39 ;
      RECT  117.38 91.73 117.89 91.49 ;
      RECT  115.91 92.52 116.45 91.97 ;
      RECT  121.43 91.25 120.29 90.87 ;
      RECT  119.03 91.49 118.82 91.42 ;
      RECT  118.82 90.63 118.31 90.39 ;
      RECT  121.22 91.73 118.82 91.49 ;
      RECT  118.82 91.49 118.62 91.42 ;
      RECT  119.03 90.7 118.82 90.63 ;
      RECT  118.31 91.73 118.1 91.49 ;
      POLYGON  119.75 91.25 119.75 90.87 119.2 90.87 119.2 90.94 118.82 90.94 118.82 91.18 119.2 91.18 119.2 91.25 119.75 91.25 ;
      RECT  118.31 91.25 118.1 90.87 ;
      RECT  121.43 92.52 121.22 91.97 ;
      RECT  121.22 92.52 120.29 91.97 ;
      RECT  120.29 91.25 119.75 90.87 ;
      RECT  118.31 90.63 118.1 90.39 ;
      RECT  119.75 92.52 118.1 91.97 ;
      RECT  121.43 91.73 121.22 91.49 ;
      RECT  118.82 90.7 118.62 90.63 ;
      POLYGON  118.45 91.25 118.45 91.18 118.82 91.18 118.82 90.94 118.45 90.94 118.45 90.87 118.31 90.87 118.31 91.25 118.45 91.25 ;
      RECT  121.43 90.63 121.22 90.39 ;
      RECT  121.22 90.63 118.82 90.39 ;
      RECT  118.82 91.73 118.31 91.49 ;
      RECT  120.29 92.52 119.75 91.97 ;
      RECT  121.01 91.25 122.15 90.87 ;
      RECT  123.41 91.49 123.62 91.42 ;
      RECT  123.62 90.63 124.13 90.39 ;
      RECT  121.22 91.73 123.62 91.49 ;
      RECT  123.62 91.49 123.82 91.42 ;
      RECT  123.41 90.7 123.62 90.63 ;
      RECT  124.13 91.73 124.34 91.49 ;
      POLYGON  122.69 91.25 122.69 90.87 123.24 90.87 123.24 90.94 123.62 90.94 123.62 91.18 123.24 91.18 123.24 91.25 122.69 91.25 ;
      RECT  124.13 91.25 124.34 90.87 ;
      RECT  121.01 92.52 121.22 91.97 ;
      RECT  121.22 92.52 122.15 91.97 ;
      RECT  122.15 91.25 122.69 90.87 ;
      RECT  124.13 90.63 124.34 90.39 ;
      RECT  122.69 92.52 124.34 91.97 ;
      RECT  121.01 91.73 121.22 91.49 ;
      RECT  123.62 90.7 123.82 90.63 ;
      POLYGON  123.99 91.25 123.99 91.18 123.62 91.18 123.62 90.94 123.99 90.94 123.99 90.87 124.13 90.87 124.13 91.25 123.99 91.25 ;
      RECT  121.01 90.63 121.22 90.39 ;
      RECT  121.22 90.63 123.62 90.39 ;
      RECT  123.62 91.73 124.13 91.49 ;
      RECT  122.15 92.52 122.69 91.97 ;
      RECT  127.67 91.25 126.53 90.87 ;
      RECT  125.27 91.49 125.06 91.42 ;
      RECT  125.06 90.63 124.55 90.39 ;
      RECT  127.46 91.73 125.06 91.49 ;
      RECT  125.06 91.49 124.86 91.42 ;
      RECT  125.27 90.7 125.06 90.63 ;
      RECT  124.55 91.73 124.34 91.49 ;
      POLYGON  125.99 91.25 125.99 90.87 125.44 90.87 125.44 90.94 125.06 90.94 125.06 91.18 125.44 91.18 125.44 91.25 125.99 91.25 ;
      RECT  124.55 91.25 124.34 90.87 ;
      RECT  127.67 92.52 127.46 91.97 ;
      RECT  127.46 92.52 126.53 91.97 ;
      RECT  126.53 91.25 125.99 90.87 ;
      RECT  124.55 90.63 124.34 90.39 ;
      RECT  125.99 92.52 124.34 91.97 ;
      RECT  127.67 91.73 127.46 91.49 ;
      RECT  125.06 90.7 124.86 90.63 ;
      POLYGON  124.69 91.25 124.69 91.18 125.06 91.18 125.06 90.94 124.69 90.94 124.69 90.87 124.55 90.87 124.55 91.25 124.69 91.25 ;
      RECT  127.67 90.63 127.46 90.39 ;
      RECT  127.46 90.63 125.06 90.39 ;
      RECT  125.06 91.73 124.55 91.49 ;
      RECT  126.53 92.52 125.99 91.97 ;
      RECT  127.25 91.25 128.39 90.87 ;
      RECT  129.65 91.49 129.86 91.42 ;
      RECT  129.86 90.63 130.37 90.39 ;
      RECT  127.46 91.73 129.86 91.49 ;
      RECT  129.86 91.49 130.06 91.42 ;
      RECT  129.65 90.7 129.86 90.63 ;
      RECT  130.37 91.73 130.58 91.49 ;
      POLYGON  128.93 91.25 128.93 90.87 129.48 90.87 129.48 90.94 129.86 90.94 129.86 91.18 129.48 91.18 129.48 91.25 128.93 91.25 ;
      RECT  130.37 91.25 130.58 90.87 ;
      RECT  127.25 92.52 127.46 91.97 ;
      RECT  127.46 92.52 128.39 91.97 ;
      RECT  128.39 91.25 128.93 90.87 ;
      RECT  130.37 90.63 130.58 90.39 ;
      RECT  128.93 92.52 130.58 91.97 ;
      RECT  127.25 91.73 127.46 91.49 ;
      RECT  129.86 90.7 130.06 90.63 ;
      POLYGON  130.23 91.25 130.23 91.18 129.86 91.18 129.86 90.94 130.23 90.94 130.23 90.87 130.37 90.87 130.37 91.25 130.23 91.25 ;
      RECT  127.25 90.63 127.46 90.39 ;
      RECT  127.46 90.63 129.86 90.39 ;
      RECT  129.86 91.73 130.37 91.49 ;
      RECT  128.39 92.52 128.93 91.97 ;
      RECT  133.91 91.25 132.77 90.87 ;
      RECT  131.51 91.49 131.3 91.42 ;
      RECT  131.3 90.63 130.79 90.39 ;
      RECT  133.7 91.73 131.3 91.49 ;
      RECT  131.3 91.49 131.1 91.42 ;
      RECT  131.51 90.7 131.3 90.63 ;
      RECT  130.79 91.73 130.58 91.49 ;
      POLYGON  132.23 91.25 132.23 90.87 131.68 90.87 131.68 90.94 131.3 90.94 131.3 91.18 131.68 91.18 131.68 91.25 132.23 91.25 ;
      RECT  130.79 91.25 130.58 90.87 ;
      RECT  133.91 92.52 133.7 91.97 ;
      RECT  133.7 92.52 132.77 91.97 ;
      RECT  132.77 91.25 132.23 90.87 ;
      RECT  130.79 90.63 130.58 90.39 ;
      RECT  132.23 92.52 130.58 91.97 ;
      RECT  133.91 91.73 133.7 91.49 ;
      RECT  131.3 90.7 131.1 90.63 ;
      POLYGON  130.93 91.25 130.93 91.18 131.3 91.18 131.3 90.94 130.93 90.94 130.93 90.87 130.79 90.87 130.79 91.25 130.93 91.25 ;
      RECT  133.91 90.63 133.7 90.39 ;
      RECT  133.7 90.63 131.3 90.39 ;
      RECT  131.3 91.73 130.79 91.49 ;
      RECT  132.77 92.52 132.23 91.97 ;
      RECT  133.49 91.25 134.63 90.87 ;
      RECT  135.89 91.49 136.1 91.42 ;
      RECT  136.1 90.63 136.61 90.39 ;
      RECT  133.7 91.73 136.1 91.49 ;
      RECT  136.1 91.49 136.3 91.42 ;
      RECT  135.89 90.7 136.1 90.63 ;
      RECT  136.61 91.73 136.82 91.49 ;
      POLYGON  135.17 91.25 135.17 90.87 135.72 90.87 135.72 90.94 136.1 90.94 136.1 91.18 135.72 91.18 135.72 91.25 135.17 91.25 ;
      RECT  136.61 91.25 136.82 90.87 ;
      RECT  133.49 92.52 133.7 91.97 ;
      RECT  133.7 92.52 134.63 91.97 ;
      RECT  134.63 91.25 135.17 90.87 ;
      RECT  136.61 90.63 136.82 90.39 ;
      RECT  135.17 92.52 136.82 91.97 ;
      RECT  133.49 91.73 133.7 91.49 ;
      RECT  136.1 90.7 136.3 90.63 ;
      POLYGON  136.47 91.25 136.47 91.18 136.1 91.18 136.1 90.94 136.47 90.94 136.47 90.87 136.61 90.87 136.61 91.25 136.47 91.25 ;
      RECT  133.49 90.63 133.7 90.39 ;
      RECT  133.7 90.63 136.1 90.39 ;
      RECT  136.1 91.73 136.61 91.49 ;
      RECT  134.63 92.52 135.17 91.97 ;
      RECT  140.15 91.25 139.01 90.87 ;
      RECT  137.75 91.49 137.54 91.42 ;
      RECT  137.54 90.63 137.03 90.39 ;
      RECT  139.94 91.73 137.54 91.49 ;
      RECT  137.54 91.49 137.34 91.42 ;
      RECT  137.75 90.7 137.54 90.63 ;
      RECT  137.03 91.73 136.82 91.49 ;
      POLYGON  138.47 91.25 138.47 90.87 137.92 90.87 137.92 90.94 137.54 90.94 137.54 91.18 137.92 91.18 137.92 91.25 138.47 91.25 ;
      RECT  137.03 91.25 136.82 90.87 ;
      RECT  140.15 92.52 139.94 91.97 ;
      RECT  139.94 92.52 139.01 91.97 ;
      RECT  139.01 91.25 138.47 90.87 ;
      RECT  137.03 90.63 136.82 90.39 ;
      RECT  138.47 92.52 136.82 91.97 ;
      RECT  140.15 91.73 139.94 91.49 ;
      RECT  137.54 90.7 137.34 90.63 ;
      POLYGON  137.17 91.25 137.17 91.18 137.54 91.18 137.54 90.94 137.17 90.94 137.17 90.87 137.03 90.87 137.03 91.25 137.17 91.25 ;
      RECT  140.15 90.63 139.94 90.39 ;
      RECT  139.94 90.63 137.54 90.39 ;
      RECT  137.54 91.73 137.03 91.49 ;
      RECT  139.01 92.52 138.47 91.97 ;
      RECT  139.73 91.25 140.87 90.87 ;
      RECT  142.13 91.49 142.34 91.42 ;
      RECT  142.34 90.63 142.85 90.39 ;
      RECT  139.94 91.73 142.34 91.49 ;
      RECT  142.34 91.49 142.54 91.42 ;
      RECT  142.13 90.7 142.34 90.63 ;
      RECT  142.85 91.73 143.06 91.49 ;
      POLYGON  141.41 91.25 141.41 90.87 141.96 90.87 141.96 90.94 142.34 90.94 142.34 91.18 141.96 91.18 141.96 91.25 141.41 91.25 ;
      RECT  142.85 91.25 143.06 90.87 ;
      RECT  139.73 92.52 139.94 91.97 ;
      RECT  139.94 92.52 140.87 91.97 ;
      RECT  140.87 91.25 141.41 90.87 ;
      RECT  142.85 90.63 143.06 90.39 ;
      RECT  141.41 92.52 143.06 91.97 ;
      RECT  139.73 91.73 139.94 91.49 ;
      RECT  142.34 90.7 142.54 90.63 ;
      POLYGON  142.71 91.25 142.71 91.18 142.34 91.18 142.34 90.94 142.71 90.94 142.71 90.87 142.85 90.87 142.85 91.25 142.71 91.25 ;
      RECT  139.73 90.63 139.94 90.39 ;
      RECT  139.94 90.63 142.34 90.39 ;
      RECT  142.34 91.73 142.85 91.49 ;
      RECT  140.87 92.52 141.41 91.97 ;
      RECT  146.39 91.25 145.25 90.87 ;
      RECT  143.99 91.49 143.78 91.42 ;
      RECT  143.78 90.63 143.27 90.39 ;
      RECT  146.18 91.73 143.78 91.49 ;
      RECT  143.78 91.49 143.58 91.42 ;
      RECT  143.99 90.7 143.78 90.63 ;
      RECT  143.27 91.73 143.06 91.49 ;
      POLYGON  144.71 91.25 144.71 90.87 144.16 90.87 144.16 90.94 143.78 90.94 143.78 91.18 144.16 91.18 144.16 91.25 144.71 91.25 ;
      RECT  143.27 91.25 143.06 90.87 ;
      RECT  146.39 92.52 146.18 91.97 ;
      RECT  146.18 92.52 145.25 91.97 ;
      RECT  145.25 91.25 144.71 90.87 ;
      RECT  143.27 90.63 143.06 90.39 ;
      RECT  144.71 92.52 143.06 91.97 ;
      RECT  146.39 91.73 146.18 91.49 ;
      RECT  143.78 90.7 143.58 90.63 ;
      POLYGON  143.41 91.25 143.41 91.18 143.78 91.18 143.78 90.94 143.41 90.94 143.41 90.87 143.27 90.87 143.27 91.25 143.41 91.25 ;
      RECT  146.39 90.63 146.18 90.39 ;
      RECT  146.18 90.63 143.78 90.39 ;
      RECT  143.78 91.73 143.27 91.49 ;
      RECT  145.25 92.52 144.71 91.97 ;
      RECT  96.26 90.63 146.18 90.39 ;
      RECT  96.26 91.73 146.18 91.49 ;
      RECT  107.27 92.52 107.81 91.97 ;
      RECT  97.19 91.25 97.73 90.87 ;
      RECT  122.15 92.52 122.69 91.97 ;
      RECT  138.47 91.25 139.01 90.87 ;
      RECT  97.19 92.52 97.73 91.97 ;
      RECT  125.99 91.25 126.53 90.87 ;
      RECT  138.47 92.52 139.01 91.97 ;
      RECT  122.15 91.25 122.69 90.87 ;
      RECT  144.71 91.25 145.25 90.87 ;
      RECT  134.63 91.25 135.17 90.87 ;
      RECT  113.51 91.25 114.05 90.87 ;
      RECT  103.43 92.52 103.97 91.97 ;
      RECT  140.87 91.25 141.41 90.87 ;
      RECT  115.91 91.25 116.45 90.87 ;
      RECT  109.67 91.25 110.21 90.87 ;
      RECT  119.75 91.25 120.29 90.87 ;
      RECT  140.87 92.52 141.41 91.97 ;
      RECT  103.43 91.25 103.97 90.87 ;
      RECT  115.91 92.52 116.45 91.97 ;
      RECT  101.03 91.25 101.57 90.87 ;
      RECT  113.51 92.52 114.05 91.97 ;
      RECT  132.23 92.52 132.77 91.97 ;
      RECT  132.23 91.25 132.77 90.87 ;
      RECT  101.03 92.52 101.57 91.97 ;
      RECT  128.39 92.52 128.93 91.97 ;
      RECT  144.71 92.52 145.25 91.97 ;
      RECT  119.75 92.52 120.29 91.97 ;
      RECT  128.39 91.25 128.93 90.87 ;
      RECT  107.27 91.25 107.81 90.87 ;
      RECT  134.63 92.52 135.17 91.97 ;
      RECT  109.67 92.52 110.21 91.97 ;
      RECT  125.99 92.52 126.53 91.97 ;
      RECT  96.05 124.84 97.19 125.22 ;
      RECT  98.45 124.6 98.66 124.67 ;
      RECT  98.66 125.46 99.17 125.7 ;
      RECT  96.26 124.36 98.66 124.6 ;
      RECT  98.66 124.6 98.86 124.67 ;
      RECT  98.45 125.39 98.66 125.46 ;
      RECT  99.17 124.36 99.38 124.6 ;
      POLYGON  97.73 124.84 97.73 125.22 98.28 125.22 98.28 125.15 98.66 125.15 98.66 124.91 98.28 124.91 98.28 124.84 97.73 124.84 ;
      RECT  99.17 124.84 99.38 125.22 ;
      RECT  96.05 123.57 96.26 124.12 ;
      RECT  96.26 123.57 97.19 124.12 ;
      RECT  97.19 124.84 97.73 125.22 ;
      RECT  99.17 125.46 99.38 125.7 ;
      RECT  97.73 123.57 99.38 124.12 ;
      RECT  96.05 124.36 96.26 124.6 ;
      RECT  98.66 125.39 98.86 125.46 ;
      POLYGON  99.03 124.84 99.03 124.91 98.66 124.91 98.66 125.15 99.03 125.15 99.03 125.22 99.17 125.22 99.17 124.84 99.03 124.84 ;
      RECT  96.05 125.46 96.26 125.7 ;
      RECT  96.26 125.46 98.66 125.7 ;
      RECT  98.66 124.36 99.17 124.6 ;
      RECT  97.19 123.57 97.73 124.12 ;
      RECT  102.71 124.84 101.57 125.22 ;
      RECT  100.31 124.6 100.1 124.67 ;
      RECT  100.1 125.46 99.59 125.7 ;
      RECT  102.5 124.36 100.1 124.6 ;
      RECT  100.1 124.6 99.9 124.67 ;
      RECT  100.31 125.39 100.1 125.46 ;
      RECT  99.59 124.36 99.38 124.6 ;
      POLYGON  101.03 124.84 101.03 125.22 100.48 125.22 100.48 125.15 100.1 125.15 100.1 124.91 100.48 124.91 100.48 124.84 101.03 124.84 ;
      RECT  99.59 124.84 99.38 125.22 ;
      RECT  102.71 123.57 102.5 124.12 ;
      RECT  102.5 123.57 101.57 124.12 ;
      RECT  101.57 124.84 101.03 125.22 ;
      RECT  99.59 125.46 99.38 125.7 ;
      RECT  101.03 123.57 99.38 124.12 ;
      RECT  102.71 124.36 102.5 124.6 ;
      RECT  100.1 125.39 99.9 125.46 ;
      POLYGON  99.73 124.84 99.73 124.91 100.1 124.91 100.1 125.15 99.73 125.15 99.73 125.22 99.59 125.22 99.59 124.84 99.73 124.84 ;
      RECT  102.71 125.46 102.5 125.7 ;
      RECT  102.5 125.46 100.1 125.7 ;
      RECT  100.1 124.36 99.59 124.6 ;
      RECT  101.57 123.57 101.03 124.12 ;
      RECT  102.29 124.84 103.43 125.22 ;
      RECT  104.69 124.6 104.9 124.67 ;
      RECT  104.9 125.46 105.41 125.7 ;
      RECT  102.5 124.36 104.9 124.6 ;
      RECT  104.9 124.6 105.1 124.67 ;
      RECT  104.69 125.39 104.9 125.46 ;
      RECT  105.41 124.36 105.62 124.6 ;
      POLYGON  103.97 124.84 103.97 125.22 104.52 125.22 104.52 125.15 104.9 125.15 104.9 124.91 104.52 124.91 104.52 124.84 103.97 124.84 ;
      RECT  105.41 124.84 105.62 125.22 ;
      RECT  102.29 123.57 102.5 124.12 ;
      RECT  102.5 123.57 103.43 124.12 ;
      RECT  103.43 124.84 103.97 125.22 ;
      RECT  105.41 125.46 105.62 125.7 ;
      RECT  103.97 123.57 105.62 124.12 ;
      RECT  102.29 124.36 102.5 124.6 ;
      RECT  104.9 125.39 105.1 125.46 ;
      POLYGON  105.27 124.84 105.27 124.91 104.9 124.91 104.9 125.15 105.27 125.15 105.27 125.22 105.41 125.22 105.41 124.84 105.27 124.84 ;
      RECT  102.29 125.46 102.5 125.7 ;
      RECT  102.5 125.46 104.9 125.7 ;
      RECT  104.9 124.36 105.41 124.6 ;
      RECT  103.43 123.57 103.97 124.12 ;
      RECT  108.95 124.84 107.81 125.22 ;
      RECT  106.55 124.6 106.34 124.67 ;
      RECT  106.34 125.46 105.83 125.7 ;
      RECT  108.74 124.36 106.34 124.6 ;
      RECT  106.34 124.6 106.14 124.67 ;
      RECT  106.55 125.39 106.34 125.46 ;
      RECT  105.83 124.36 105.62 124.6 ;
      POLYGON  107.27 124.84 107.27 125.22 106.72 125.22 106.72 125.15 106.34 125.15 106.34 124.91 106.72 124.91 106.72 124.84 107.27 124.84 ;
      RECT  105.83 124.84 105.62 125.22 ;
      RECT  108.95 123.57 108.74 124.12 ;
      RECT  108.74 123.57 107.81 124.12 ;
      RECT  107.81 124.84 107.27 125.22 ;
      RECT  105.83 125.46 105.62 125.7 ;
      RECT  107.27 123.57 105.62 124.12 ;
      RECT  108.95 124.36 108.74 124.6 ;
      RECT  106.34 125.39 106.14 125.46 ;
      POLYGON  105.97 124.84 105.97 124.91 106.34 124.91 106.34 125.15 105.97 125.15 105.97 125.22 105.83 125.22 105.83 124.84 105.97 124.84 ;
      RECT  108.95 125.46 108.74 125.7 ;
      RECT  108.74 125.46 106.34 125.7 ;
      RECT  106.34 124.36 105.83 124.6 ;
      RECT  107.81 123.57 107.27 124.12 ;
      RECT  108.53 124.84 109.67 125.22 ;
      RECT  110.93 124.6 111.14 124.67 ;
      RECT  111.14 125.46 111.65 125.7 ;
      RECT  108.74 124.36 111.14 124.6 ;
      RECT  111.14 124.6 111.34 124.67 ;
      RECT  110.93 125.39 111.14 125.46 ;
      RECT  111.65 124.36 111.86 124.6 ;
      POLYGON  110.21 124.84 110.21 125.22 110.76 125.22 110.76 125.15 111.14 125.15 111.14 124.91 110.76 124.91 110.76 124.84 110.21 124.84 ;
      RECT  111.65 124.84 111.86 125.22 ;
      RECT  108.53 123.57 108.74 124.12 ;
      RECT  108.74 123.57 109.67 124.12 ;
      RECT  109.67 124.84 110.21 125.22 ;
      RECT  111.65 125.46 111.86 125.7 ;
      RECT  110.21 123.57 111.86 124.12 ;
      RECT  108.53 124.36 108.74 124.6 ;
      RECT  111.14 125.39 111.34 125.46 ;
      POLYGON  111.51 124.84 111.51 124.91 111.14 124.91 111.14 125.15 111.51 125.15 111.51 125.22 111.65 125.22 111.65 124.84 111.51 124.84 ;
      RECT  108.53 125.46 108.74 125.7 ;
      RECT  108.74 125.46 111.14 125.7 ;
      RECT  111.14 124.36 111.65 124.6 ;
      RECT  109.67 123.57 110.21 124.12 ;
      RECT  115.19 124.84 114.05 125.22 ;
      RECT  112.79 124.6 112.58 124.67 ;
      RECT  112.58 125.46 112.07 125.7 ;
      RECT  114.98 124.36 112.58 124.6 ;
      RECT  112.58 124.6 112.38 124.67 ;
      RECT  112.79 125.39 112.58 125.46 ;
      RECT  112.07 124.36 111.86 124.6 ;
      POLYGON  113.51 124.84 113.51 125.22 112.96 125.22 112.96 125.15 112.58 125.15 112.58 124.91 112.96 124.91 112.96 124.84 113.51 124.84 ;
      RECT  112.07 124.84 111.86 125.22 ;
      RECT  115.19 123.57 114.98 124.12 ;
      RECT  114.98 123.57 114.05 124.12 ;
      RECT  114.05 124.84 113.51 125.22 ;
      RECT  112.07 125.46 111.86 125.7 ;
      RECT  113.51 123.57 111.86 124.12 ;
      RECT  115.19 124.36 114.98 124.6 ;
      RECT  112.58 125.39 112.38 125.46 ;
      POLYGON  112.21 124.84 112.21 124.91 112.58 124.91 112.58 125.15 112.21 125.15 112.21 125.22 112.07 125.22 112.07 124.84 112.21 124.84 ;
      RECT  115.19 125.46 114.98 125.7 ;
      RECT  114.98 125.46 112.58 125.7 ;
      RECT  112.58 124.36 112.07 124.6 ;
      RECT  114.05 123.57 113.51 124.12 ;
      RECT  114.77 124.84 115.91 125.22 ;
      RECT  117.17 124.6 117.38 124.67 ;
      RECT  117.38 125.46 117.89 125.7 ;
      RECT  114.98 124.36 117.38 124.6 ;
      RECT  117.38 124.6 117.58 124.67 ;
      RECT  117.17 125.39 117.38 125.46 ;
      RECT  117.89 124.36 118.1 124.6 ;
      POLYGON  116.45 124.84 116.45 125.22 117.0 125.22 117.0 125.15 117.38 125.15 117.38 124.91 117.0 124.91 117.0 124.84 116.45 124.84 ;
      RECT  117.89 124.84 118.1 125.22 ;
      RECT  114.77 123.57 114.98 124.12 ;
      RECT  114.98 123.57 115.91 124.12 ;
      RECT  115.91 124.84 116.45 125.22 ;
      RECT  117.89 125.46 118.1 125.7 ;
      RECT  116.45 123.57 118.1 124.12 ;
      RECT  114.77 124.36 114.98 124.6 ;
      RECT  117.38 125.39 117.58 125.46 ;
      POLYGON  117.75 124.84 117.75 124.91 117.38 124.91 117.38 125.15 117.75 125.15 117.75 125.22 117.89 125.22 117.89 124.84 117.75 124.84 ;
      RECT  114.77 125.46 114.98 125.7 ;
      RECT  114.98 125.46 117.38 125.7 ;
      RECT  117.38 124.36 117.89 124.6 ;
      RECT  115.91 123.57 116.45 124.12 ;
      RECT  121.43 124.84 120.29 125.22 ;
      RECT  119.03 124.6 118.82 124.67 ;
      RECT  118.82 125.46 118.31 125.7 ;
      RECT  121.22 124.36 118.82 124.6 ;
      RECT  118.82 124.6 118.62 124.67 ;
      RECT  119.03 125.39 118.82 125.46 ;
      RECT  118.31 124.36 118.1 124.6 ;
      POLYGON  119.75 124.84 119.75 125.22 119.2 125.22 119.2 125.15 118.82 125.15 118.82 124.91 119.2 124.91 119.2 124.84 119.75 124.84 ;
      RECT  118.31 124.84 118.1 125.22 ;
      RECT  121.43 123.57 121.22 124.12 ;
      RECT  121.22 123.57 120.29 124.12 ;
      RECT  120.29 124.84 119.75 125.22 ;
      RECT  118.31 125.46 118.1 125.7 ;
      RECT  119.75 123.57 118.1 124.12 ;
      RECT  121.43 124.36 121.22 124.6 ;
      RECT  118.82 125.39 118.62 125.46 ;
      POLYGON  118.45 124.84 118.45 124.91 118.82 124.91 118.82 125.15 118.45 125.15 118.45 125.22 118.31 125.22 118.31 124.84 118.45 124.84 ;
      RECT  121.43 125.46 121.22 125.7 ;
      RECT  121.22 125.46 118.82 125.7 ;
      RECT  118.82 124.36 118.31 124.6 ;
      RECT  120.29 123.57 119.75 124.12 ;
      RECT  121.01 124.84 122.15 125.22 ;
      RECT  123.41 124.6 123.62 124.67 ;
      RECT  123.62 125.46 124.13 125.7 ;
      RECT  121.22 124.36 123.62 124.6 ;
      RECT  123.62 124.6 123.82 124.67 ;
      RECT  123.41 125.39 123.62 125.46 ;
      RECT  124.13 124.36 124.34 124.6 ;
      POLYGON  122.69 124.84 122.69 125.22 123.24 125.22 123.24 125.15 123.62 125.15 123.62 124.91 123.24 124.91 123.24 124.84 122.69 124.84 ;
      RECT  124.13 124.84 124.34 125.22 ;
      RECT  121.01 123.57 121.22 124.12 ;
      RECT  121.22 123.57 122.15 124.12 ;
      RECT  122.15 124.84 122.69 125.22 ;
      RECT  124.13 125.46 124.34 125.7 ;
      RECT  122.69 123.57 124.34 124.12 ;
      RECT  121.01 124.36 121.22 124.6 ;
      RECT  123.62 125.39 123.82 125.46 ;
      POLYGON  123.99 124.84 123.99 124.91 123.62 124.91 123.62 125.15 123.99 125.15 123.99 125.22 124.13 125.22 124.13 124.84 123.99 124.84 ;
      RECT  121.01 125.46 121.22 125.7 ;
      RECT  121.22 125.46 123.62 125.7 ;
      RECT  123.62 124.36 124.13 124.6 ;
      RECT  122.15 123.57 122.69 124.12 ;
      RECT  127.67 124.84 126.53 125.22 ;
      RECT  125.27 124.6 125.06 124.67 ;
      RECT  125.06 125.46 124.55 125.7 ;
      RECT  127.46 124.36 125.06 124.6 ;
      RECT  125.06 124.6 124.86 124.67 ;
      RECT  125.27 125.39 125.06 125.46 ;
      RECT  124.55 124.36 124.34 124.6 ;
      POLYGON  125.99 124.84 125.99 125.22 125.44 125.22 125.44 125.15 125.06 125.15 125.06 124.91 125.44 124.91 125.44 124.84 125.99 124.84 ;
      RECT  124.55 124.84 124.34 125.22 ;
      RECT  127.67 123.57 127.46 124.12 ;
      RECT  127.46 123.57 126.53 124.12 ;
      RECT  126.53 124.84 125.99 125.22 ;
      RECT  124.55 125.46 124.34 125.7 ;
      RECT  125.99 123.57 124.34 124.12 ;
      RECT  127.67 124.36 127.46 124.6 ;
      RECT  125.06 125.39 124.86 125.46 ;
      POLYGON  124.69 124.84 124.69 124.91 125.06 124.91 125.06 125.15 124.69 125.15 124.69 125.22 124.55 125.22 124.55 124.84 124.69 124.84 ;
      RECT  127.67 125.46 127.46 125.7 ;
      RECT  127.46 125.46 125.06 125.7 ;
      RECT  125.06 124.36 124.55 124.6 ;
      RECT  126.53 123.57 125.99 124.12 ;
      RECT  127.25 124.84 128.39 125.22 ;
      RECT  129.65 124.6 129.86 124.67 ;
      RECT  129.86 125.46 130.37 125.7 ;
      RECT  127.46 124.36 129.86 124.6 ;
      RECT  129.86 124.6 130.06 124.67 ;
      RECT  129.65 125.39 129.86 125.46 ;
      RECT  130.37 124.36 130.58 124.6 ;
      POLYGON  128.93 124.84 128.93 125.22 129.48 125.22 129.48 125.15 129.86 125.15 129.86 124.91 129.48 124.91 129.48 124.84 128.93 124.84 ;
      RECT  130.37 124.84 130.58 125.22 ;
      RECT  127.25 123.57 127.46 124.12 ;
      RECT  127.46 123.57 128.39 124.12 ;
      RECT  128.39 124.84 128.93 125.22 ;
      RECT  130.37 125.46 130.58 125.7 ;
      RECT  128.93 123.57 130.58 124.12 ;
      RECT  127.25 124.36 127.46 124.6 ;
      RECT  129.86 125.39 130.06 125.46 ;
      POLYGON  130.23 124.84 130.23 124.91 129.86 124.91 129.86 125.15 130.23 125.15 130.23 125.22 130.37 125.22 130.37 124.84 130.23 124.84 ;
      RECT  127.25 125.46 127.46 125.7 ;
      RECT  127.46 125.46 129.86 125.7 ;
      RECT  129.86 124.36 130.37 124.6 ;
      RECT  128.39 123.57 128.93 124.12 ;
      RECT  133.91 124.84 132.77 125.22 ;
      RECT  131.51 124.6 131.3 124.67 ;
      RECT  131.3 125.46 130.79 125.7 ;
      RECT  133.7 124.36 131.3 124.6 ;
      RECT  131.3 124.6 131.1 124.67 ;
      RECT  131.51 125.39 131.3 125.46 ;
      RECT  130.79 124.36 130.58 124.6 ;
      POLYGON  132.23 124.84 132.23 125.22 131.68 125.22 131.68 125.15 131.3 125.15 131.3 124.91 131.68 124.91 131.68 124.84 132.23 124.84 ;
      RECT  130.79 124.84 130.58 125.22 ;
      RECT  133.91 123.57 133.7 124.12 ;
      RECT  133.7 123.57 132.77 124.12 ;
      RECT  132.77 124.84 132.23 125.22 ;
      RECT  130.79 125.46 130.58 125.7 ;
      RECT  132.23 123.57 130.58 124.12 ;
      RECT  133.91 124.36 133.7 124.6 ;
      RECT  131.3 125.39 131.1 125.46 ;
      POLYGON  130.93 124.84 130.93 124.91 131.3 124.91 131.3 125.15 130.93 125.15 130.93 125.22 130.79 125.22 130.79 124.84 130.93 124.84 ;
      RECT  133.91 125.46 133.7 125.7 ;
      RECT  133.7 125.46 131.3 125.7 ;
      RECT  131.3 124.36 130.79 124.6 ;
      RECT  132.77 123.57 132.23 124.12 ;
      RECT  133.49 124.84 134.63 125.22 ;
      RECT  135.89 124.6 136.1 124.67 ;
      RECT  136.1 125.46 136.61 125.7 ;
      RECT  133.7 124.36 136.1 124.6 ;
      RECT  136.1 124.6 136.3 124.67 ;
      RECT  135.89 125.39 136.1 125.46 ;
      RECT  136.61 124.36 136.82 124.6 ;
      POLYGON  135.17 124.84 135.17 125.22 135.72 125.22 135.72 125.15 136.1 125.15 136.1 124.91 135.72 124.91 135.72 124.84 135.17 124.84 ;
      RECT  136.61 124.84 136.82 125.22 ;
      RECT  133.49 123.57 133.7 124.12 ;
      RECT  133.7 123.57 134.63 124.12 ;
      RECT  134.63 124.84 135.17 125.22 ;
      RECT  136.61 125.46 136.82 125.7 ;
      RECT  135.17 123.57 136.82 124.12 ;
      RECT  133.49 124.36 133.7 124.6 ;
      RECT  136.1 125.39 136.3 125.46 ;
      POLYGON  136.47 124.84 136.47 124.91 136.1 124.91 136.1 125.15 136.47 125.15 136.47 125.22 136.61 125.22 136.61 124.84 136.47 124.84 ;
      RECT  133.49 125.46 133.7 125.7 ;
      RECT  133.7 125.46 136.1 125.7 ;
      RECT  136.1 124.36 136.61 124.6 ;
      RECT  134.63 123.57 135.17 124.12 ;
      RECT  140.15 124.84 139.01 125.22 ;
      RECT  137.75 124.6 137.54 124.67 ;
      RECT  137.54 125.46 137.03 125.7 ;
      RECT  139.94 124.36 137.54 124.6 ;
      RECT  137.54 124.6 137.34 124.67 ;
      RECT  137.75 125.39 137.54 125.46 ;
      RECT  137.03 124.36 136.82 124.6 ;
      POLYGON  138.47 124.84 138.47 125.22 137.92 125.22 137.92 125.15 137.54 125.15 137.54 124.91 137.92 124.91 137.92 124.84 138.47 124.84 ;
      RECT  137.03 124.84 136.82 125.22 ;
      RECT  140.15 123.57 139.94 124.12 ;
      RECT  139.94 123.57 139.01 124.12 ;
      RECT  139.01 124.84 138.47 125.22 ;
      RECT  137.03 125.46 136.82 125.7 ;
      RECT  138.47 123.57 136.82 124.12 ;
      RECT  140.15 124.36 139.94 124.6 ;
      RECT  137.54 125.39 137.34 125.46 ;
      POLYGON  137.17 124.84 137.17 124.91 137.54 124.91 137.54 125.15 137.17 125.15 137.17 125.22 137.03 125.22 137.03 124.84 137.17 124.84 ;
      RECT  140.15 125.46 139.94 125.7 ;
      RECT  139.94 125.46 137.54 125.7 ;
      RECT  137.54 124.36 137.03 124.6 ;
      RECT  139.01 123.57 138.47 124.12 ;
      RECT  139.73 124.84 140.87 125.22 ;
      RECT  142.13 124.6 142.34 124.67 ;
      RECT  142.34 125.46 142.85 125.7 ;
      RECT  139.94 124.36 142.34 124.6 ;
      RECT  142.34 124.6 142.54 124.67 ;
      RECT  142.13 125.39 142.34 125.46 ;
      RECT  142.85 124.36 143.06 124.6 ;
      POLYGON  141.41 124.84 141.41 125.22 141.96 125.22 141.96 125.15 142.34 125.15 142.34 124.91 141.96 124.91 141.96 124.84 141.41 124.84 ;
      RECT  142.85 124.84 143.06 125.22 ;
      RECT  139.73 123.57 139.94 124.12 ;
      RECT  139.94 123.57 140.87 124.12 ;
      RECT  140.87 124.84 141.41 125.22 ;
      RECT  142.85 125.46 143.06 125.7 ;
      RECT  141.41 123.57 143.06 124.12 ;
      RECT  139.73 124.36 139.94 124.6 ;
      RECT  142.34 125.39 142.54 125.46 ;
      POLYGON  142.71 124.84 142.71 124.91 142.34 124.91 142.34 125.15 142.71 125.15 142.71 125.22 142.85 125.22 142.85 124.84 142.71 124.84 ;
      RECT  139.73 125.46 139.94 125.7 ;
      RECT  139.94 125.46 142.34 125.7 ;
      RECT  142.34 124.36 142.85 124.6 ;
      RECT  140.87 123.57 141.41 124.12 ;
      RECT  146.39 124.84 145.25 125.22 ;
      RECT  143.99 124.6 143.78 124.67 ;
      RECT  143.78 125.46 143.27 125.7 ;
      RECT  146.18 124.36 143.78 124.6 ;
      RECT  143.78 124.6 143.58 124.67 ;
      RECT  143.99 125.39 143.78 125.46 ;
      RECT  143.27 124.36 143.06 124.6 ;
      POLYGON  144.71 124.84 144.71 125.22 144.16 125.22 144.16 125.15 143.78 125.15 143.78 124.91 144.16 124.91 144.16 124.84 144.71 124.84 ;
      RECT  143.27 124.84 143.06 125.22 ;
      RECT  146.39 123.57 146.18 124.12 ;
      RECT  146.18 123.57 145.25 124.12 ;
      RECT  145.25 124.84 144.71 125.22 ;
      RECT  143.27 125.46 143.06 125.7 ;
      RECT  144.71 123.57 143.06 124.12 ;
      RECT  146.39 124.36 146.18 124.6 ;
      RECT  143.78 125.39 143.58 125.46 ;
      POLYGON  143.41 124.84 143.41 124.91 143.78 124.91 143.78 125.15 143.41 125.15 143.41 125.22 143.27 125.22 143.27 124.84 143.41 124.84 ;
      RECT  146.39 125.46 146.18 125.7 ;
      RECT  146.18 125.46 143.78 125.7 ;
      RECT  143.78 124.36 143.27 124.6 ;
      RECT  145.25 123.57 144.71 124.12 ;
      RECT  96.26 125.46 146.18 125.7 ;
      RECT  96.26 124.36 146.18 124.6 ;
      RECT  107.27 123.57 107.81 124.12 ;
      RECT  97.19 124.84 97.73 125.22 ;
      RECT  122.15 123.57 122.69 124.12 ;
      RECT  138.47 124.84 139.01 125.22 ;
      RECT  97.19 123.57 97.73 124.12 ;
      RECT  125.99 124.84 126.53 125.22 ;
      RECT  138.47 123.57 139.01 124.12 ;
      RECT  122.15 124.84 122.69 125.22 ;
      RECT  144.71 124.84 145.25 125.22 ;
      RECT  134.63 124.84 135.17 125.22 ;
      RECT  113.51 124.84 114.05 125.22 ;
      RECT  103.43 123.57 103.97 124.12 ;
      RECT  140.87 124.84 141.41 125.22 ;
      RECT  115.91 124.84 116.45 125.22 ;
      RECT  109.67 124.84 110.21 125.22 ;
      RECT  119.75 124.84 120.29 125.22 ;
      RECT  140.87 123.57 141.41 124.12 ;
      RECT  103.43 124.84 103.97 125.22 ;
      RECT  115.91 123.57 116.45 124.12 ;
      RECT  101.03 124.84 101.57 125.22 ;
      RECT  113.51 123.57 114.05 124.12 ;
      RECT  132.23 123.57 132.77 124.12 ;
      RECT  132.23 124.84 132.77 125.22 ;
      RECT  101.03 123.57 101.57 124.12 ;
      RECT  128.39 123.57 128.93 124.12 ;
      RECT  144.71 123.57 145.25 124.12 ;
      RECT  119.75 123.57 120.29 124.12 ;
      RECT  128.39 124.84 128.93 125.22 ;
      RECT  107.27 124.84 107.81 125.22 ;
      RECT  134.63 123.57 135.17 124.12 ;
      RECT  109.67 123.57 110.21 124.12 ;
      RECT  125.99 123.57 126.53 124.12 ;
      RECT  96.26 89.165 99.38 89.715 ;
      RECT  102.5 89.165 99.38 89.715 ;
      RECT  102.5 89.165 105.62 89.715 ;
      RECT  108.74 89.165 105.62 89.715 ;
      RECT  108.74 89.165 111.86 89.715 ;
      RECT  114.98 89.165 111.86 89.715 ;
      RECT  114.98 89.165 118.1 89.715 ;
      RECT  121.22 89.165 118.1 89.715 ;
      RECT  121.22 89.165 124.34 89.715 ;
      RECT  127.46 89.165 124.34 89.715 ;
      RECT  127.46 89.165 130.58 89.715 ;
      RECT  133.7 89.165 130.58 89.715 ;
      RECT  133.7 89.165 136.82 89.715 ;
      RECT  139.94 89.165 136.82 89.715 ;
      RECT  139.94 89.165 143.06 89.715 ;
      RECT  146.18 89.165 143.06 89.715 ;
      RECT  96.26 126.925 99.38 126.375 ;
      RECT  102.5 126.925 99.38 126.375 ;
      RECT  102.5 126.925 105.62 126.375 ;
      RECT  108.74 126.925 105.62 126.375 ;
      RECT  108.74 126.925 111.86 126.375 ;
      RECT  114.98 126.925 111.86 126.375 ;
      RECT  114.98 126.925 118.1 126.375 ;
      RECT  121.22 126.925 118.1 126.375 ;
      RECT  121.22 126.925 124.34 126.375 ;
      RECT  127.46 126.925 124.34 126.375 ;
      RECT  127.46 126.925 130.58 126.375 ;
      RECT  133.7 126.925 130.58 126.375 ;
      RECT  133.7 126.925 136.82 126.375 ;
      RECT  139.94 126.925 136.82 126.375 ;
      RECT  139.94 126.925 143.06 126.375 ;
      RECT  146.18 126.925 143.06 126.375 ;
      RECT  89.81 91.25 90.95 90.87 ;
      RECT  92.21 91.49 92.42 91.42 ;
      RECT  92.42 90.63 92.93 90.39 ;
      RECT  90.02 91.73 92.42 91.49 ;
      RECT  92.42 91.49 92.62 91.42 ;
      RECT  92.21 90.7 92.42 90.63 ;
      RECT  92.93 91.73 93.14 91.49 ;
      POLYGON  91.49 91.25 91.49 90.87 92.04 90.87 92.04 90.94 92.42 90.94 92.42 91.18 92.04 91.18 92.04 91.25 91.49 91.25 ;
      RECT  92.93 91.25 93.14 90.87 ;
      RECT  89.81 92.52 90.02 91.97 ;
      RECT  90.02 92.52 90.95 91.97 ;
      RECT  90.95 91.25 91.49 90.87 ;
      RECT  92.93 90.63 93.14 90.39 ;
      RECT  91.49 92.52 93.14 91.97 ;
      RECT  89.81 91.73 90.02 91.49 ;
      RECT  92.42 90.7 92.62 90.63 ;
      POLYGON  92.79 91.25 92.79 91.18 92.42 91.18 92.42 90.94 92.79 90.94 92.79 90.87 92.93 90.87 92.93 91.25 92.79 91.25 ;
      RECT  89.81 90.63 90.02 90.39 ;
      RECT  90.02 90.63 92.42 90.39 ;
      RECT  92.42 91.73 92.93 91.49 ;
      RECT  90.95 92.52 91.49 91.97 ;
      RECT  89.81 93.24 90.95 93.62 ;
      RECT  92.21 93.0 92.42 93.07 ;
      RECT  92.42 93.86 92.93 94.1 ;
      RECT  90.02 92.76 92.42 93.0 ;
      RECT  92.42 93.0 92.62 93.07 ;
      RECT  92.21 93.79 92.42 93.86 ;
      RECT  92.93 92.76 93.14 93.0 ;
      POLYGON  91.49 93.24 91.49 93.62 92.04 93.62 92.04 93.55 92.42 93.55 92.42 93.31 92.04 93.31 92.04 93.24 91.49 93.24 ;
      RECT  92.93 93.24 93.14 93.62 ;
      RECT  89.81 91.97 90.02 92.52 ;
      RECT  90.02 91.97 90.95 92.52 ;
      RECT  90.95 93.24 91.49 93.62 ;
      RECT  92.93 93.86 93.14 94.1 ;
      RECT  91.49 91.97 93.14 92.52 ;
      RECT  89.81 92.76 90.02 93.0 ;
      RECT  92.42 93.79 92.62 93.86 ;
      POLYGON  92.79 93.24 92.79 93.31 92.42 93.31 92.42 93.55 92.79 93.55 92.79 93.62 92.93 93.62 92.93 93.24 92.79 93.24 ;
      RECT  89.81 93.86 90.02 94.1 ;
      RECT  90.02 93.86 92.42 94.1 ;
      RECT  92.42 92.76 92.93 93.0 ;
      RECT  90.95 91.97 91.49 92.52 ;
      RECT  89.81 95.2 90.95 94.82 ;
      RECT  92.21 95.44 92.42 95.37 ;
      RECT  92.42 94.58 92.93 94.34 ;
      RECT  90.02 95.68 92.42 95.44 ;
      RECT  92.42 95.44 92.62 95.37 ;
      RECT  92.21 94.65 92.42 94.58 ;
      RECT  92.93 95.68 93.14 95.44 ;
      POLYGON  91.49 95.2 91.49 94.82 92.04 94.82 92.04 94.89 92.42 94.89 92.42 95.13 92.04 95.13 92.04 95.2 91.49 95.2 ;
      RECT  92.93 95.2 93.14 94.82 ;
      RECT  89.81 96.47 90.02 95.92 ;
      RECT  90.02 96.47 90.95 95.92 ;
      RECT  90.95 95.2 91.49 94.82 ;
      RECT  92.93 94.58 93.14 94.34 ;
      RECT  91.49 96.47 93.14 95.92 ;
      RECT  89.81 95.68 90.02 95.44 ;
      RECT  92.42 94.65 92.62 94.58 ;
      POLYGON  92.79 95.2 92.79 95.13 92.42 95.13 92.42 94.89 92.79 94.89 92.79 94.82 92.93 94.82 92.93 95.2 92.79 95.2 ;
      RECT  89.81 94.58 90.02 94.34 ;
      RECT  90.02 94.58 92.42 94.34 ;
      RECT  92.42 95.68 92.93 95.44 ;
      RECT  90.95 96.47 91.49 95.92 ;
      RECT  89.81 97.19 90.95 97.57 ;
      RECT  92.21 96.95 92.42 97.02 ;
      RECT  92.42 97.81 92.93 98.05 ;
      RECT  90.02 96.71 92.42 96.95 ;
      RECT  92.42 96.95 92.62 97.02 ;
      RECT  92.21 97.74 92.42 97.81 ;
      RECT  92.93 96.71 93.14 96.95 ;
      POLYGON  91.49 97.19 91.49 97.57 92.04 97.57 92.04 97.5 92.42 97.5 92.42 97.26 92.04 97.26 92.04 97.19 91.49 97.19 ;
      RECT  92.93 97.19 93.14 97.57 ;
      RECT  89.81 95.92 90.02 96.47 ;
      RECT  90.02 95.92 90.95 96.47 ;
      RECT  90.95 97.19 91.49 97.57 ;
      RECT  92.93 97.81 93.14 98.05 ;
      RECT  91.49 95.92 93.14 96.47 ;
      RECT  89.81 96.71 90.02 96.95 ;
      RECT  92.42 97.74 92.62 97.81 ;
      POLYGON  92.79 97.19 92.79 97.26 92.42 97.26 92.42 97.5 92.79 97.5 92.79 97.57 92.93 97.57 92.93 97.19 92.79 97.19 ;
      RECT  89.81 97.81 90.02 98.05 ;
      RECT  90.02 97.81 92.42 98.05 ;
      RECT  92.42 96.71 92.93 96.95 ;
      RECT  90.95 95.92 91.49 96.47 ;
      RECT  89.81 99.15 90.95 98.77 ;
      RECT  92.21 99.39 92.42 99.32 ;
      RECT  92.42 98.53 92.93 98.29 ;
      RECT  90.02 99.63 92.42 99.39 ;
      RECT  92.42 99.39 92.62 99.32 ;
      RECT  92.21 98.6 92.42 98.53 ;
      RECT  92.93 99.63 93.14 99.39 ;
      POLYGON  91.49 99.15 91.49 98.77 92.04 98.77 92.04 98.84 92.42 98.84 92.42 99.08 92.04 99.08 92.04 99.15 91.49 99.15 ;
      RECT  92.93 99.15 93.14 98.77 ;
      RECT  89.81 100.42 90.02 99.87 ;
      RECT  90.02 100.42 90.95 99.87 ;
      RECT  90.95 99.15 91.49 98.77 ;
      RECT  92.93 98.53 93.14 98.29 ;
      RECT  91.49 100.42 93.14 99.87 ;
      RECT  89.81 99.63 90.02 99.39 ;
      RECT  92.42 98.6 92.62 98.53 ;
      POLYGON  92.79 99.15 92.79 99.08 92.42 99.08 92.42 98.84 92.79 98.84 92.79 98.77 92.93 98.77 92.93 99.15 92.79 99.15 ;
      RECT  89.81 98.53 90.02 98.29 ;
      RECT  90.02 98.53 92.42 98.29 ;
      RECT  92.42 99.63 92.93 99.39 ;
      RECT  90.95 100.42 91.49 99.87 ;
      RECT  89.81 101.14 90.95 101.52 ;
      RECT  92.21 100.9 92.42 100.97 ;
      RECT  92.42 101.76 92.93 102.0 ;
      RECT  90.02 100.66 92.42 100.9 ;
      RECT  92.42 100.9 92.62 100.97 ;
      RECT  92.21 101.69 92.42 101.76 ;
      RECT  92.93 100.66 93.14 100.9 ;
      POLYGON  91.49 101.14 91.49 101.52 92.04 101.52 92.04 101.45 92.42 101.45 92.42 101.21 92.04 101.21 92.04 101.14 91.49 101.14 ;
      RECT  92.93 101.14 93.14 101.52 ;
      RECT  89.81 99.87 90.02 100.42 ;
      RECT  90.02 99.87 90.95 100.42 ;
      RECT  90.95 101.14 91.49 101.52 ;
      RECT  92.93 101.76 93.14 102.0 ;
      RECT  91.49 99.87 93.14 100.42 ;
      RECT  89.81 100.66 90.02 100.9 ;
      RECT  92.42 101.69 92.62 101.76 ;
      POLYGON  92.79 101.14 92.79 101.21 92.42 101.21 92.42 101.45 92.79 101.45 92.79 101.52 92.93 101.52 92.93 101.14 92.79 101.14 ;
      RECT  89.81 101.76 90.02 102.0 ;
      RECT  90.02 101.76 92.42 102.0 ;
      RECT  92.42 100.66 92.93 100.9 ;
      RECT  90.95 99.87 91.49 100.42 ;
      RECT  89.81 103.1 90.95 102.72 ;
      RECT  92.21 103.34 92.42 103.27 ;
      RECT  92.42 102.48 92.93 102.24 ;
      RECT  90.02 103.58 92.42 103.34 ;
      RECT  92.42 103.34 92.62 103.27 ;
      RECT  92.21 102.55 92.42 102.48 ;
      RECT  92.93 103.58 93.14 103.34 ;
      POLYGON  91.49 103.1 91.49 102.72 92.04 102.72 92.04 102.79 92.42 102.79 92.42 103.03 92.04 103.03 92.04 103.1 91.49 103.1 ;
      RECT  92.93 103.1 93.14 102.72 ;
      RECT  89.81 104.37 90.02 103.82 ;
      RECT  90.02 104.37 90.95 103.82 ;
      RECT  90.95 103.1 91.49 102.72 ;
      RECT  92.93 102.48 93.14 102.24 ;
      RECT  91.49 104.37 93.14 103.82 ;
      RECT  89.81 103.58 90.02 103.34 ;
      RECT  92.42 102.55 92.62 102.48 ;
      POLYGON  92.79 103.1 92.79 103.03 92.42 103.03 92.42 102.79 92.79 102.79 92.79 102.72 92.93 102.72 92.93 103.1 92.79 103.1 ;
      RECT  89.81 102.48 90.02 102.24 ;
      RECT  90.02 102.48 92.42 102.24 ;
      RECT  92.42 103.58 92.93 103.34 ;
      RECT  90.95 104.37 91.49 103.82 ;
      RECT  89.81 105.09 90.95 105.47 ;
      RECT  92.21 104.85 92.42 104.92 ;
      RECT  92.42 105.71 92.93 105.95 ;
      RECT  90.02 104.61 92.42 104.85 ;
      RECT  92.42 104.85 92.62 104.92 ;
      RECT  92.21 105.64 92.42 105.71 ;
      RECT  92.93 104.61 93.14 104.85 ;
      POLYGON  91.49 105.09 91.49 105.47 92.04 105.47 92.04 105.4 92.42 105.4 92.42 105.16 92.04 105.16 92.04 105.09 91.49 105.09 ;
      RECT  92.93 105.09 93.14 105.47 ;
      RECT  89.81 103.82 90.02 104.37 ;
      RECT  90.02 103.82 90.95 104.37 ;
      RECT  90.95 105.09 91.49 105.47 ;
      RECT  92.93 105.71 93.14 105.95 ;
      RECT  91.49 103.82 93.14 104.37 ;
      RECT  89.81 104.61 90.02 104.85 ;
      RECT  92.42 105.64 92.62 105.71 ;
      POLYGON  92.79 105.09 92.79 105.16 92.42 105.16 92.42 105.4 92.79 105.4 92.79 105.47 92.93 105.47 92.93 105.09 92.79 105.09 ;
      RECT  89.81 105.71 90.02 105.95 ;
      RECT  90.02 105.71 92.42 105.95 ;
      RECT  92.42 104.61 92.93 104.85 ;
      RECT  90.95 103.82 91.49 104.37 ;
      RECT  89.81 107.05 90.95 106.67 ;
      RECT  92.21 107.29 92.42 107.22 ;
      RECT  92.42 106.43 92.93 106.19 ;
      RECT  90.02 107.53 92.42 107.29 ;
      RECT  92.42 107.29 92.62 107.22 ;
      RECT  92.21 106.5 92.42 106.43 ;
      RECT  92.93 107.53 93.14 107.29 ;
      POLYGON  91.49 107.05 91.49 106.67 92.04 106.67 92.04 106.74 92.42 106.74 92.42 106.98 92.04 106.98 92.04 107.05 91.49 107.05 ;
      RECT  92.93 107.05 93.14 106.67 ;
      RECT  89.81 108.32 90.02 107.77 ;
      RECT  90.02 108.32 90.95 107.77 ;
      RECT  90.95 107.05 91.49 106.67 ;
      RECT  92.93 106.43 93.14 106.19 ;
      RECT  91.49 108.32 93.14 107.77 ;
      RECT  89.81 107.53 90.02 107.29 ;
      RECT  92.42 106.5 92.62 106.43 ;
      POLYGON  92.79 107.05 92.79 106.98 92.42 106.98 92.42 106.74 92.79 106.74 92.79 106.67 92.93 106.67 92.93 107.05 92.79 107.05 ;
      RECT  89.81 106.43 90.02 106.19 ;
      RECT  90.02 106.43 92.42 106.19 ;
      RECT  92.42 107.53 92.93 107.29 ;
      RECT  90.95 108.32 91.49 107.77 ;
      RECT  89.81 109.04 90.95 109.42 ;
      RECT  92.21 108.8 92.42 108.87 ;
      RECT  92.42 109.66 92.93 109.9 ;
      RECT  90.02 108.56 92.42 108.8 ;
      RECT  92.42 108.8 92.62 108.87 ;
      RECT  92.21 109.59 92.42 109.66 ;
      RECT  92.93 108.56 93.14 108.8 ;
      POLYGON  91.49 109.04 91.49 109.42 92.04 109.42 92.04 109.35 92.42 109.35 92.42 109.11 92.04 109.11 92.04 109.04 91.49 109.04 ;
      RECT  92.93 109.04 93.14 109.42 ;
      RECT  89.81 107.77 90.02 108.32 ;
      RECT  90.02 107.77 90.95 108.32 ;
      RECT  90.95 109.04 91.49 109.42 ;
      RECT  92.93 109.66 93.14 109.9 ;
      RECT  91.49 107.77 93.14 108.32 ;
      RECT  89.81 108.56 90.02 108.8 ;
      RECT  92.42 109.59 92.62 109.66 ;
      POLYGON  92.79 109.04 92.79 109.11 92.42 109.11 92.42 109.35 92.79 109.35 92.79 109.42 92.93 109.42 92.93 109.04 92.79 109.04 ;
      RECT  89.81 109.66 90.02 109.9 ;
      RECT  90.02 109.66 92.42 109.9 ;
      RECT  92.42 108.56 92.93 108.8 ;
      RECT  90.95 107.77 91.49 108.32 ;
      RECT  89.81 111.0 90.95 110.62 ;
      RECT  92.21 111.24 92.42 111.17 ;
      RECT  92.42 110.38 92.93 110.14 ;
      RECT  90.02 111.48 92.42 111.24 ;
      RECT  92.42 111.24 92.62 111.17 ;
      RECT  92.21 110.45 92.42 110.38 ;
      RECT  92.93 111.48 93.14 111.24 ;
      POLYGON  91.49 111.0 91.49 110.62 92.04 110.62 92.04 110.69 92.42 110.69 92.42 110.93 92.04 110.93 92.04 111.0 91.49 111.0 ;
      RECT  92.93 111.0 93.14 110.62 ;
      RECT  89.81 112.27 90.02 111.72 ;
      RECT  90.02 112.27 90.95 111.72 ;
      RECT  90.95 111.0 91.49 110.62 ;
      RECT  92.93 110.38 93.14 110.14 ;
      RECT  91.49 112.27 93.14 111.72 ;
      RECT  89.81 111.48 90.02 111.24 ;
      RECT  92.42 110.45 92.62 110.38 ;
      POLYGON  92.79 111.0 92.79 110.93 92.42 110.93 92.42 110.69 92.79 110.69 92.79 110.62 92.93 110.62 92.93 111.0 92.79 111.0 ;
      RECT  89.81 110.38 90.02 110.14 ;
      RECT  90.02 110.38 92.42 110.14 ;
      RECT  92.42 111.48 92.93 111.24 ;
      RECT  90.95 112.27 91.49 111.72 ;
      RECT  89.81 112.99 90.95 113.37 ;
      RECT  92.21 112.75 92.42 112.82 ;
      RECT  92.42 113.61 92.93 113.85 ;
      RECT  90.02 112.51 92.42 112.75 ;
      RECT  92.42 112.75 92.62 112.82 ;
      RECT  92.21 113.54 92.42 113.61 ;
      RECT  92.93 112.51 93.14 112.75 ;
      POLYGON  91.49 112.99 91.49 113.37 92.04 113.37 92.04 113.3 92.42 113.3 92.42 113.06 92.04 113.06 92.04 112.99 91.49 112.99 ;
      RECT  92.93 112.99 93.14 113.37 ;
      RECT  89.81 111.72 90.02 112.27 ;
      RECT  90.02 111.72 90.95 112.27 ;
      RECT  90.95 112.99 91.49 113.37 ;
      RECT  92.93 113.61 93.14 113.85 ;
      RECT  91.49 111.72 93.14 112.27 ;
      RECT  89.81 112.51 90.02 112.75 ;
      RECT  92.42 113.54 92.62 113.61 ;
      POLYGON  92.79 112.99 92.79 113.06 92.42 113.06 92.42 113.3 92.79 113.3 92.79 113.37 92.93 113.37 92.93 112.99 92.79 112.99 ;
      RECT  89.81 113.61 90.02 113.85 ;
      RECT  90.02 113.61 92.42 113.85 ;
      RECT  92.42 112.51 92.93 112.75 ;
      RECT  90.95 111.72 91.49 112.27 ;
      RECT  89.81 114.95 90.95 114.57 ;
      RECT  92.21 115.19 92.42 115.12 ;
      RECT  92.42 114.33 92.93 114.09 ;
      RECT  90.02 115.43 92.42 115.19 ;
      RECT  92.42 115.19 92.62 115.12 ;
      RECT  92.21 114.4 92.42 114.33 ;
      RECT  92.93 115.43 93.14 115.19 ;
      POLYGON  91.49 114.95 91.49 114.57 92.04 114.57 92.04 114.64 92.42 114.64 92.42 114.88 92.04 114.88 92.04 114.95 91.49 114.95 ;
      RECT  92.93 114.95 93.14 114.57 ;
      RECT  89.81 116.22 90.02 115.67 ;
      RECT  90.02 116.22 90.95 115.67 ;
      RECT  90.95 114.95 91.49 114.57 ;
      RECT  92.93 114.33 93.14 114.09 ;
      RECT  91.49 116.22 93.14 115.67 ;
      RECT  89.81 115.43 90.02 115.19 ;
      RECT  92.42 114.4 92.62 114.33 ;
      POLYGON  92.79 114.95 92.79 114.88 92.42 114.88 92.42 114.64 92.79 114.64 92.79 114.57 92.93 114.57 92.93 114.95 92.79 114.95 ;
      RECT  89.81 114.33 90.02 114.09 ;
      RECT  90.02 114.33 92.42 114.09 ;
      RECT  92.42 115.43 92.93 115.19 ;
      RECT  90.95 116.22 91.49 115.67 ;
      RECT  89.81 116.94 90.95 117.32 ;
      RECT  92.21 116.7 92.42 116.77 ;
      RECT  92.42 117.56 92.93 117.8 ;
      RECT  90.02 116.46 92.42 116.7 ;
      RECT  92.42 116.7 92.62 116.77 ;
      RECT  92.21 117.49 92.42 117.56 ;
      RECT  92.93 116.46 93.14 116.7 ;
      POLYGON  91.49 116.94 91.49 117.32 92.04 117.32 92.04 117.25 92.42 117.25 92.42 117.01 92.04 117.01 92.04 116.94 91.49 116.94 ;
      RECT  92.93 116.94 93.14 117.32 ;
      RECT  89.81 115.67 90.02 116.22 ;
      RECT  90.02 115.67 90.95 116.22 ;
      RECT  90.95 116.94 91.49 117.32 ;
      RECT  92.93 117.56 93.14 117.8 ;
      RECT  91.49 115.67 93.14 116.22 ;
      RECT  89.81 116.46 90.02 116.7 ;
      RECT  92.42 117.49 92.62 117.56 ;
      POLYGON  92.79 116.94 92.79 117.01 92.42 117.01 92.42 117.25 92.79 117.25 92.79 117.32 92.93 117.32 92.93 116.94 92.79 116.94 ;
      RECT  89.81 117.56 90.02 117.8 ;
      RECT  90.02 117.56 92.42 117.8 ;
      RECT  92.42 116.46 92.93 116.7 ;
      RECT  90.95 115.67 91.49 116.22 ;
      RECT  89.81 118.9 90.95 118.52 ;
      RECT  92.21 119.14 92.42 119.07 ;
      RECT  92.42 118.28 92.93 118.04 ;
      RECT  90.02 119.38 92.42 119.14 ;
      RECT  92.42 119.14 92.62 119.07 ;
      RECT  92.21 118.35 92.42 118.28 ;
      RECT  92.93 119.38 93.14 119.14 ;
      POLYGON  91.49 118.9 91.49 118.52 92.04 118.52 92.04 118.59 92.42 118.59 92.42 118.83 92.04 118.83 92.04 118.9 91.49 118.9 ;
      RECT  92.93 118.9 93.14 118.52 ;
      RECT  89.81 120.17 90.02 119.62 ;
      RECT  90.02 120.17 90.95 119.62 ;
      RECT  90.95 118.9 91.49 118.52 ;
      RECT  92.93 118.28 93.14 118.04 ;
      RECT  91.49 120.17 93.14 119.62 ;
      RECT  89.81 119.38 90.02 119.14 ;
      RECT  92.42 118.35 92.62 118.28 ;
      POLYGON  92.79 118.9 92.79 118.83 92.42 118.83 92.42 118.59 92.79 118.59 92.79 118.52 92.93 118.52 92.93 118.9 92.79 118.9 ;
      RECT  89.81 118.28 90.02 118.04 ;
      RECT  90.02 118.28 92.42 118.04 ;
      RECT  92.42 119.38 92.93 119.14 ;
      RECT  90.95 120.17 91.49 119.62 ;
      RECT  89.81 120.89 90.95 121.27 ;
      RECT  92.21 120.65 92.42 120.72 ;
      RECT  92.42 121.51 92.93 121.75 ;
      RECT  90.02 120.41 92.42 120.65 ;
      RECT  92.42 120.65 92.62 120.72 ;
      RECT  92.21 121.44 92.42 121.51 ;
      RECT  92.93 120.41 93.14 120.65 ;
      POLYGON  91.49 120.89 91.49 121.27 92.04 121.27 92.04 121.2 92.42 121.2 92.42 120.96 92.04 120.96 92.04 120.89 91.49 120.89 ;
      RECT  92.93 120.89 93.14 121.27 ;
      RECT  89.81 119.62 90.02 120.17 ;
      RECT  90.02 119.62 90.95 120.17 ;
      RECT  90.95 120.89 91.49 121.27 ;
      RECT  92.93 121.51 93.14 121.75 ;
      RECT  91.49 119.62 93.14 120.17 ;
      RECT  89.81 120.41 90.02 120.65 ;
      RECT  92.42 121.44 92.62 121.51 ;
      POLYGON  92.79 120.89 92.79 120.96 92.42 120.96 92.42 121.2 92.79 121.2 92.79 121.27 92.93 121.27 92.93 120.89 92.79 120.89 ;
      RECT  89.81 121.51 90.02 121.75 ;
      RECT  90.02 121.51 92.42 121.75 ;
      RECT  92.42 120.41 92.93 120.65 ;
      RECT  90.95 119.62 91.49 120.17 ;
      RECT  89.81 122.85 90.95 122.47 ;
      RECT  92.21 123.09 92.42 123.02 ;
      RECT  92.42 122.23 92.93 121.99 ;
      RECT  90.02 123.33 92.42 123.09 ;
      RECT  92.42 123.09 92.62 123.02 ;
      RECT  92.21 122.3 92.42 122.23 ;
      RECT  92.93 123.33 93.14 123.09 ;
      POLYGON  91.49 122.85 91.49 122.47 92.04 122.47 92.04 122.54 92.42 122.54 92.42 122.78 92.04 122.78 92.04 122.85 91.49 122.85 ;
      RECT  92.93 122.85 93.14 122.47 ;
      RECT  89.81 124.12 90.02 123.57 ;
      RECT  90.02 124.12 90.95 123.57 ;
      RECT  90.95 122.85 91.49 122.47 ;
      RECT  92.93 122.23 93.14 121.99 ;
      RECT  91.49 124.12 93.14 123.57 ;
      RECT  89.81 123.33 90.02 123.09 ;
      RECT  92.42 122.3 92.62 122.23 ;
      POLYGON  92.79 122.85 92.79 122.78 92.42 122.78 92.42 122.54 92.79 122.54 92.79 122.47 92.93 122.47 92.93 122.85 92.79 122.85 ;
      RECT  89.81 122.23 90.02 121.99 ;
      RECT  90.02 122.23 92.42 121.99 ;
      RECT  92.42 123.33 92.93 123.09 ;
      RECT  90.95 124.12 91.49 123.57 ;
      RECT  89.81 124.84 90.95 125.22 ;
      RECT  92.21 124.6 92.42 124.67 ;
      RECT  92.42 125.46 92.93 125.7 ;
      RECT  90.02 124.36 92.42 124.6 ;
      RECT  92.42 124.6 92.62 124.67 ;
      RECT  92.21 125.39 92.42 125.46 ;
      RECT  92.93 124.36 93.14 124.6 ;
      POLYGON  91.49 124.84 91.49 125.22 92.04 125.22 92.04 125.15 92.42 125.15 92.42 124.91 92.04 124.91 92.04 124.84 91.49 124.84 ;
      RECT  92.93 124.84 93.14 125.22 ;
      RECT  89.81 123.57 90.02 124.12 ;
      RECT  90.02 123.57 90.95 124.12 ;
      RECT  90.95 124.84 91.49 125.22 ;
      RECT  92.93 125.46 93.14 125.7 ;
      RECT  91.49 123.57 93.14 124.12 ;
      RECT  89.81 124.36 90.02 124.6 ;
      RECT  92.42 125.39 92.62 125.46 ;
      POLYGON  92.79 124.84 92.79 124.91 92.42 124.91 92.42 125.15 92.79 125.15 92.79 125.22 92.93 125.22 92.93 124.84 92.79 124.84 ;
      RECT  89.81 125.46 90.02 125.7 ;
      RECT  90.02 125.46 92.42 125.7 ;
      RECT  92.42 124.36 92.93 124.6 ;
      RECT  90.95 123.57 91.49 124.12 ;
      RECT  90.02 90.39 93.14 90.63 ;
      RECT  90.02 91.49 93.14 91.73 ;
      RECT  90.02 93.86 93.14 94.1 ;
      RECT  90.02 92.76 93.14 93.0 ;
      RECT  90.02 94.34 93.14 94.58 ;
      RECT  90.02 95.44 93.14 95.68 ;
      RECT  90.02 97.81 93.14 98.05 ;
      RECT  90.02 96.71 93.14 96.95 ;
      RECT  90.02 98.29 93.14 98.53 ;
      RECT  90.02 99.39 93.14 99.63 ;
      RECT  90.02 101.76 93.14 102.0 ;
      RECT  90.02 100.66 93.14 100.9 ;
      RECT  90.02 102.24 93.14 102.48 ;
      RECT  90.02 103.34 93.14 103.58 ;
      RECT  90.02 105.71 93.14 105.95 ;
      RECT  90.02 104.61 93.14 104.85 ;
      RECT  90.02 106.19 93.14 106.43 ;
      RECT  90.02 107.29 93.14 107.53 ;
      RECT  90.02 109.66 93.14 109.9 ;
      RECT  90.02 108.56 93.14 108.8 ;
      RECT  90.02 110.14 93.14 110.38 ;
      RECT  90.02 111.24 93.14 111.48 ;
      RECT  90.02 113.61 93.14 113.85 ;
      RECT  90.02 112.51 93.14 112.75 ;
      RECT  90.02 114.09 93.14 114.33 ;
      RECT  90.02 115.19 93.14 115.43 ;
      RECT  90.02 117.56 93.14 117.8 ;
      RECT  90.02 116.46 93.14 116.7 ;
      RECT  90.02 118.04 93.14 118.28 ;
      RECT  90.02 119.14 93.14 119.38 ;
      RECT  90.02 121.51 93.14 121.75 ;
      RECT  90.02 120.41 93.14 120.65 ;
      RECT  90.02 121.99 93.14 122.23 ;
      RECT  90.02 123.09 93.14 123.33 ;
      RECT  90.02 125.46 93.14 125.7 ;
      RECT  90.02 124.36 93.14 124.6 ;
      RECT  152.63 91.25 151.49 90.87 ;
      RECT  150.23 91.49 150.02 91.42 ;
      RECT  150.02 90.63 149.51 90.39 ;
      RECT  152.42 91.73 150.02 91.49 ;
      RECT  150.02 91.49 149.82 91.42 ;
      RECT  150.23 90.7 150.02 90.63 ;
      RECT  149.51 91.73 149.3 91.49 ;
      POLYGON  150.95 91.25 150.95 90.87 150.4 90.87 150.4 90.94 150.02 90.94 150.02 91.18 150.4 91.18 150.4 91.25 150.95 91.25 ;
      RECT  149.51 91.25 149.3 90.87 ;
      RECT  152.63 92.52 152.42 91.97 ;
      RECT  152.42 92.52 151.49 91.97 ;
      RECT  151.49 91.25 150.95 90.87 ;
      RECT  149.51 90.63 149.3 90.39 ;
      RECT  150.95 92.52 149.3 91.97 ;
      RECT  152.63 91.73 152.42 91.49 ;
      RECT  150.02 90.7 149.82 90.63 ;
      POLYGON  149.65 91.25 149.65 91.18 150.02 91.18 150.02 90.94 149.65 90.94 149.65 90.87 149.51 90.87 149.51 91.25 149.65 91.25 ;
      RECT  152.63 90.63 152.42 90.39 ;
      RECT  152.42 90.63 150.02 90.39 ;
      RECT  150.02 91.73 149.51 91.49 ;
      RECT  151.49 92.52 150.95 91.97 ;
      RECT  152.63 93.24 151.49 93.62 ;
      RECT  150.23 93.0 150.02 93.07 ;
      RECT  150.02 93.86 149.51 94.1 ;
      RECT  152.42 92.76 150.02 93.0 ;
      RECT  150.02 93.0 149.82 93.07 ;
      RECT  150.23 93.79 150.02 93.86 ;
      RECT  149.51 92.76 149.3 93.0 ;
      POLYGON  150.95 93.24 150.95 93.62 150.4 93.62 150.4 93.55 150.02 93.55 150.02 93.31 150.4 93.31 150.4 93.24 150.95 93.24 ;
      RECT  149.51 93.24 149.3 93.62 ;
      RECT  152.63 91.97 152.42 92.52 ;
      RECT  152.42 91.97 151.49 92.52 ;
      RECT  151.49 93.24 150.95 93.62 ;
      RECT  149.51 93.86 149.3 94.1 ;
      RECT  150.95 91.97 149.3 92.52 ;
      RECT  152.63 92.76 152.42 93.0 ;
      RECT  150.02 93.79 149.82 93.86 ;
      POLYGON  149.65 93.24 149.65 93.31 150.02 93.31 150.02 93.55 149.65 93.55 149.65 93.62 149.51 93.62 149.51 93.24 149.65 93.24 ;
      RECT  152.63 93.86 152.42 94.1 ;
      RECT  152.42 93.86 150.02 94.1 ;
      RECT  150.02 92.76 149.51 93.0 ;
      RECT  151.49 91.97 150.95 92.52 ;
      RECT  152.63 95.2 151.49 94.82 ;
      RECT  150.23 95.44 150.02 95.37 ;
      RECT  150.02 94.58 149.51 94.34 ;
      RECT  152.42 95.68 150.02 95.44 ;
      RECT  150.02 95.44 149.82 95.37 ;
      RECT  150.23 94.65 150.02 94.58 ;
      RECT  149.51 95.68 149.3 95.44 ;
      POLYGON  150.95 95.2 150.95 94.82 150.4 94.82 150.4 94.89 150.02 94.89 150.02 95.13 150.4 95.13 150.4 95.2 150.95 95.2 ;
      RECT  149.51 95.2 149.3 94.82 ;
      RECT  152.63 96.47 152.42 95.92 ;
      RECT  152.42 96.47 151.49 95.92 ;
      RECT  151.49 95.2 150.95 94.82 ;
      RECT  149.51 94.58 149.3 94.34 ;
      RECT  150.95 96.47 149.3 95.92 ;
      RECT  152.63 95.68 152.42 95.44 ;
      RECT  150.02 94.65 149.82 94.58 ;
      POLYGON  149.65 95.2 149.65 95.13 150.02 95.13 150.02 94.89 149.65 94.89 149.65 94.82 149.51 94.82 149.51 95.2 149.65 95.2 ;
      RECT  152.63 94.58 152.42 94.34 ;
      RECT  152.42 94.58 150.02 94.34 ;
      RECT  150.02 95.68 149.51 95.44 ;
      RECT  151.49 96.47 150.95 95.92 ;
      RECT  152.63 97.19 151.49 97.57 ;
      RECT  150.23 96.95 150.02 97.02 ;
      RECT  150.02 97.81 149.51 98.05 ;
      RECT  152.42 96.71 150.02 96.95 ;
      RECT  150.02 96.95 149.82 97.02 ;
      RECT  150.23 97.74 150.02 97.81 ;
      RECT  149.51 96.71 149.3 96.95 ;
      POLYGON  150.95 97.19 150.95 97.57 150.4 97.57 150.4 97.5 150.02 97.5 150.02 97.26 150.4 97.26 150.4 97.19 150.95 97.19 ;
      RECT  149.51 97.19 149.3 97.57 ;
      RECT  152.63 95.92 152.42 96.47 ;
      RECT  152.42 95.92 151.49 96.47 ;
      RECT  151.49 97.19 150.95 97.57 ;
      RECT  149.51 97.81 149.3 98.05 ;
      RECT  150.95 95.92 149.3 96.47 ;
      RECT  152.63 96.71 152.42 96.95 ;
      RECT  150.02 97.74 149.82 97.81 ;
      POLYGON  149.65 97.19 149.65 97.26 150.02 97.26 150.02 97.5 149.65 97.5 149.65 97.57 149.51 97.57 149.51 97.19 149.65 97.19 ;
      RECT  152.63 97.81 152.42 98.05 ;
      RECT  152.42 97.81 150.02 98.05 ;
      RECT  150.02 96.71 149.51 96.95 ;
      RECT  151.49 95.92 150.95 96.47 ;
      RECT  152.63 99.15 151.49 98.77 ;
      RECT  150.23 99.39 150.02 99.32 ;
      RECT  150.02 98.53 149.51 98.29 ;
      RECT  152.42 99.63 150.02 99.39 ;
      RECT  150.02 99.39 149.82 99.32 ;
      RECT  150.23 98.6 150.02 98.53 ;
      RECT  149.51 99.63 149.3 99.39 ;
      POLYGON  150.95 99.15 150.95 98.77 150.4 98.77 150.4 98.84 150.02 98.84 150.02 99.08 150.4 99.08 150.4 99.15 150.95 99.15 ;
      RECT  149.51 99.15 149.3 98.77 ;
      RECT  152.63 100.42 152.42 99.87 ;
      RECT  152.42 100.42 151.49 99.87 ;
      RECT  151.49 99.15 150.95 98.77 ;
      RECT  149.51 98.53 149.3 98.29 ;
      RECT  150.95 100.42 149.3 99.87 ;
      RECT  152.63 99.63 152.42 99.39 ;
      RECT  150.02 98.6 149.82 98.53 ;
      POLYGON  149.65 99.15 149.65 99.08 150.02 99.08 150.02 98.84 149.65 98.84 149.65 98.77 149.51 98.77 149.51 99.15 149.65 99.15 ;
      RECT  152.63 98.53 152.42 98.29 ;
      RECT  152.42 98.53 150.02 98.29 ;
      RECT  150.02 99.63 149.51 99.39 ;
      RECT  151.49 100.42 150.95 99.87 ;
      RECT  152.63 101.14 151.49 101.52 ;
      RECT  150.23 100.9 150.02 100.97 ;
      RECT  150.02 101.76 149.51 102.0 ;
      RECT  152.42 100.66 150.02 100.9 ;
      RECT  150.02 100.9 149.82 100.97 ;
      RECT  150.23 101.69 150.02 101.76 ;
      RECT  149.51 100.66 149.3 100.9 ;
      POLYGON  150.95 101.14 150.95 101.52 150.4 101.52 150.4 101.45 150.02 101.45 150.02 101.21 150.4 101.21 150.4 101.14 150.95 101.14 ;
      RECT  149.51 101.14 149.3 101.52 ;
      RECT  152.63 99.87 152.42 100.42 ;
      RECT  152.42 99.87 151.49 100.42 ;
      RECT  151.49 101.14 150.95 101.52 ;
      RECT  149.51 101.76 149.3 102.0 ;
      RECT  150.95 99.87 149.3 100.42 ;
      RECT  152.63 100.66 152.42 100.9 ;
      RECT  150.02 101.69 149.82 101.76 ;
      POLYGON  149.65 101.14 149.65 101.21 150.02 101.21 150.02 101.45 149.65 101.45 149.65 101.52 149.51 101.52 149.51 101.14 149.65 101.14 ;
      RECT  152.63 101.76 152.42 102.0 ;
      RECT  152.42 101.76 150.02 102.0 ;
      RECT  150.02 100.66 149.51 100.9 ;
      RECT  151.49 99.87 150.95 100.42 ;
      RECT  152.63 103.1 151.49 102.72 ;
      RECT  150.23 103.34 150.02 103.27 ;
      RECT  150.02 102.48 149.51 102.24 ;
      RECT  152.42 103.58 150.02 103.34 ;
      RECT  150.02 103.34 149.82 103.27 ;
      RECT  150.23 102.55 150.02 102.48 ;
      RECT  149.51 103.58 149.3 103.34 ;
      POLYGON  150.95 103.1 150.95 102.72 150.4 102.72 150.4 102.79 150.02 102.79 150.02 103.03 150.4 103.03 150.4 103.1 150.95 103.1 ;
      RECT  149.51 103.1 149.3 102.72 ;
      RECT  152.63 104.37 152.42 103.82 ;
      RECT  152.42 104.37 151.49 103.82 ;
      RECT  151.49 103.1 150.95 102.72 ;
      RECT  149.51 102.48 149.3 102.24 ;
      RECT  150.95 104.37 149.3 103.82 ;
      RECT  152.63 103.58 152.42 103.34 ;
      RECT  150.02 102.55 149.82 102.48 ;
      POLYGON  149.65 103.1 149.65 103.03 150.02 103.03 150.02 102.79 149.65 102.79 149.65 102.72 149.51 102.72 149.51 103.1 149.65 103.1 ;
      RECT  152.63 102.48 152.42 102.24 ;
      RECT  152.42 102.48 150.02 102.24 ;
      RECT  150.02 103.58 149.51 103.34 ;
      RECT  151.49 104.37 150.95 103.82 ;
      RECT  152.63 105.09 151.49 105.47 ;
      RECT  150.23 104.85 150.02 104.92 ;
      RECT  150.02 105.71 149.51 105.95 ;
      RECT  152.42 104.61 150.02 104.85 ;
      RECT  150.02 104.85 149.82 104.92 ;
      RECT  150.23 105.64 150.02 105.71 ;
      RECT  149.51 104.61 149.3 104.85 ;
      POLYGON  150.95 105.09 150.95 105.47 150.4 105.47 150.4 105.4 150.02 105.4 150.02 105.16 150.4 105.16 150.4 105.09 150.95 105.09 ;
      RECT  149.51 105.09 149.3 105.47 ;
      RECT  152.63 103.82 152.42 104.37 ;
      RECT  152.42 103.82 151.49 104.37 ;
      RECT  151.49 105.09 150.95 105.47 ;
      RECT  149.51 105.71 149.3 105.95 ;
      RECT  150.95 103.82 149.3 104.37 ;
      RECT  152.63 104.61 152.42 104.85 ;
      RECT  150.02 105.64 149.82 105.71 ;
      POLYGON  149.65 105.09 149.65 105.16 150.02 105.16 150.02 105.4 149.65 105.4 149.65 105.47 149.51 105.47 149.51 105.09 149.65 105.09 ;
      RECT  152.63 105.71 152.42 105.95 ;
      RECT  152.42 105.71 150.02 105.95 ;
      RECT  150.02 104.61 149.51 104.85 ;
      RECT  151.49 103.82 150.95 104.37 ;
      RECT  152.63 107.05 151.49 106.67 ;
      RECT  150.23 107.29 150.02 107.22 ;
      RECT  150.02 106.43 149.51 106.19 ;
      RECT  152.42 107.53 150.02 107.29 ;
      RECT  150.02 107.29 149.82 107.22 ;
      RECT  150.23 106.5 150.02 106.43 ;
      RECT  149.51 107.53 149.3 107.29 ;
      POLYGON  150.95 107.05 150.95 106.67 150.4 106.67 150.4 106.74 150.02 106.74 150.02 106.98 150.4 106.98 150.4 107.05 150.95 107.05 ;
      RECT  149.51 107.05 149.3 106.67 ;
      RECT  152.63 108.32 152.42 107.77 ;
      RECT  152.42 108.32 151.49 107.77 ;
      RECT  151.49 107.05 150.95 106.67 ;
      RECT  149.51 106.43 149.3 106.19 ;
      RECT  150.95 108.32 149.3 107.77 ;
      RECT  152.63 107.53 152.42 107.29 ;
      RECT  150.02 106.5 149.82 106.43 ;
      POLYGON  149.65 107.05 149.65 106.98 150.02 106.98 150.02 106.74 149.65 106.74 149.65 106.67 149.51 106.67 149.51 107.05 149.65 107.05 ;
      RECT  152.63 106.43 152.42 106.19 ;
      RECT  152.42 106.43 150.02 106.19 ;
      RECT  150.02 107.53 149.51 107.29 ;
      RECT  151.49 108.32 150.95 107.77 ;
      RECT  152.63 109.04 151.49 109.42 ;
      RECT  150.23 108.8 150.02 108.87 ;
      RECT  150.02 109.66 149.51 109.9 ;
      RECT  152.42 108.56 150.02 108.8 ;
      RECT  150.02 108.8 149.82 108.87 ;
      RECT  150.23 109.59 150.02 109.66 ;
      RECT  149.51 108.56 149.3 108.8 ;
      POLYGON  150.95 109.04 150.95 109.42 150.4 109.42 150.4 109.35 150.02 109.35 150.02 109.11 150.4 109.11 150.4 109.04 150.95 109.04 ;
      RECT  149.51 109.04 149.3 109.42 ;
      RECT  152.63 107.77 152.42 108.32 ;
      RECT  152.42 107.77 151.49 108.32 ;
      RECT  151.49 109.04 150.95 109.42 ;
      RECT  149.51 109.66 149.3 109.9 ;
      RECT  150.95 107.77 149.3 108.32 ;
      RECT  152.63 108.56 152.42 108.8 ;
      RECT  150.02 109.59 149.82 109.66 ;
      POLYGON  149.65 109.04 149.65 109.11 150.02 109.11 150.02 109.35 149.65 109.35 149.65 109.42 149.51 109.42 149.51 109.04 149.65 109.04 ;
      RECT  152.63 109.66 152.42 109.9 ;
      RECT  152.42 109.66 150.02 109.9 ;
      RECT  150.02 108.56 149.51 108.8 ;
      RECT  151.49 107.77 150.95 108.32 ;
      RECT  152.63 111.0 151.49 110.62 ;
      RECT  150.23 111.24 150.02 111.17 ;
      RECT  150.02 110.38 149.51 110.14 ;
      RECT  152.42 111.48 150.02 111.24 ;
      RECT  150.02 111.24 149.82 111.17 ;
      RECT  150.23 110.45 150.02 110.38 ;
      RECT  149.51 111.48 149.3 111.24 ;
      POLYGON  150.95 111.0 150.95 110.62 150.4 110.62 150.4 110.69 150.02 110.69 150.02 110.93 150.4 110.93 150.4 111.0 150.95 111.0 ;
      RECT  149.51 111.0 149.3 110.62 ;
      RECT  152.63 112.27 152.42 111.72 ;
      RECT  152.42 112.27 151.49 111.72 ;
      RECT  151.49 111.0 150.95 110.62 ;
      RECT  149.51 110.38 149.3 110.14 ;
      RECT  150.95 112.27 149.3 111.72 ;
      RECT  152.63 111.48 152.42 111.24 ;
      RECT  150.02 110.45 149.82 110.38 ;
      POLYGON  149.65 111.0 149.65 110.93 150.02 110.93 150.02 110.69 149.65 110.69 149.65 110.62 149.51 110.62 149.51 111.0 149.65 111.0 ;
      RECT  152.63 110.38 152.42 110.14 ;
      RECT  152.42 110.38 150.02 110.14 ;
      RECT  150.02 111.48 149.51 111.24 ;
      RECT  151.49 112.27 150.95 111.72 ;
      RECT  152.63 112.99 151.49 113.37 ;
      RECT  150.23 112.75 150.02 112.82 ;
      RECT  150.02 113.61 149.51 113.85 ;
      RECT  152.42 112.51 150.02 112.75 ;
      RECT  150.02 112.75 149.82 112.82 ;
      RECT  150.23 113.54 150.02 113.61 ;
      RECT  149.51 112.51 149.3 112.75 ;
      POLYGON  150.95 112.99 150.95 113.37 150.4 113.37 150.4 113.3 150.02 113.3 150.02 113.06 150.4 113.06 150.4 112.99 150.95 112.99 ;
      RECT  149.51 112.99 149.3 113.37 ;
      RECT  152.63 111.72 152.42 112.27 ;
      RECT  152.42 111.72 151.49 112.27 ;
      RECT  151.49 112.99 150.95 113.37 ;
      RECT  149.51 113.61 149.3 113.85 ;
      RECT  150.95 111.72 149.3 112.27 ;
      RECT  152.63 112.51 152.42 112.75 ;
      RECT  150.02 113.54 149.82 113.61 ;
      POLYGON  149.65 112.99 149.65 113.06 150.02 113.06 150.02 113.3 149.65 113.3 149.65 113.37 149.51 113.37 149.51 112.99 149.65 112.99 ;
      RECT  152.63 113.61 152.42 113.85 ;
      RECT  152.42 113.61 150.02 113.85 ;
      RECT  150.02 112.51 149.51 112.75 ;
      RECT  151.49 111.72 150.95 112.27 ;
      RECT  152.63 114.95 151.49 114.57 ;
      RECT  150.23 115.19 150.02 115.12 ;
      RECT  150.02 114.33 149.51 114.09 ;
      RECT  152.42 115.43 150.02 115.19 ;
      RECT  150.02 115.19 149.82 115.12 ;
      RECT  150.23 114.4 150.02 114.33 ;
      RECT  149.51 115.43 149.3 115.19 ;
      POLYGON  150.95 114.95 150.95 114.57 150.4 114.57 150.4 114.64 150.02 114.64 150.02 114.88 150.4 114.88 150.4 114.95 150.95 114.95 ;
      RECT  149.51 114.95 149.3 114.57 ;
      RECT  152.63 116.22 152.42 115.67 ;
      RECT  152.42 116.22 151.49 115.67 ;
      RECT  151.49 114.95 150.95 114.57 ;
      RECT  149.51 114.33 149.3 114.09 ;
      RECT  150.95 116.22 149.3 115.67 ;
      RECT  152.63 115.43 152.42 115.19 ;
      RECT  150.02 114.4 149.82 114.33 ;
      POLYGON  149.65 114.95 149.65 114.88 150.02 114.88 150.02 114.64 149.65 114.64 149.65 114.57 149.51 114.57 149.51 114.95 149.65 114.95 ;
      RECT  152.63 114.33 152.42 114.09 ;
      RECT  152.42 114.33 150.02 114.09 ;
      RECT  150.02 115.43 149.51 115.19 ;
      RECT  151.49 116.22 150.95 115.67 ;
      RECT  152.63 116.94 151.49 117.32 ;
      RECT  150.23 116.7 150.02 116.77 ;
      RECT  150.02 117.56 149.51 117.8 ;
      RECT  152.42 116.46 150.02 116.7 ;
      RECT  150.02 116.7 149.82 116.77 ;
      RECT  150.23 117.49 150.02 117.56 ;
      RECT  149.51 116.46 149.3 116.7 ;
      POLYGON  150.95 116.94 150.95 117.32 150.4 117.32 150.4 117.25 150.02 117.25 150.02 117.01 150.4 117.01 150.4 116.94 150.95 116.94 ;
      RECT  149.51 116.94 149.3 117.32 ;
      RECT  152.63 115.67 152.42 116.22 ;
      RECT  152.42 115.67 151.49 116.22 ;
      RECT  151.49 116.94 150.95 117.32 ;
      RECT  149.51 117.56 149.3 117.8 ;
      RECT  150.95 115.67 149.3 116.22 ;
      RECT  152.63 116.46 152.42 116.7 ;
      RECT  150.02 117.49 149.82 117.56 ;
      POLYGON  149.65 116.94 149.65 117.01 150.02 117.01 150.02 117.25 149.65 117.25 149.65 117.32 149.51 117.32 149.51 116.94 149.65 116.94 ;
      RECT  152.63 117.56 152.42 117.8 ;
      RECT  152.42 117.56 150.02 117.8 ;
      RECT  150.02 116.46 149.51 116.7 ;
      RECT  151.49 115.67 150.95 116.22 ;
      RECT  152.63 118.9 151.49 118.52 ;
      RECT  150.23 119.14 150.02 119.07 ;
      RECT  150.02 118.28 149.51 118.04 ;
      RECT  152.42 119.38 150.02 119.14 ;
      RECT  150.02 119.14 149.82 119.07 ;
      RECT  150.23 118.35 150.02 118.28 ;
      RECT  149.51 119.38 149.3 119.14 ;
      POLYGON  150.95 118.9 150.95 118.52 150.4 118.52 150.4 118.59 150.02 118.59 150.02 118.83 150.4 118.83 150.4 118.9 150.95 118.9 ;
      RECT  149.51 118.9 149.3 118.52 ;
      RECT  152.63 120.17 152.42 119.62 ;
      RECT  152.42 120.17 151.49 119.62 ;
      RECT  151.49 118.9 150.95 118.52 ;
      RECT  149.51 118.28 149.3 118.04 ;
      RECT  150.95 120.17 149.3 119.62 ;
      RECT  152.63 119.38 152.42 119.14 ;
      RECT  150.02 118.35 149.82 118.28 ;
      POLYGON  149.65 118.9 149.65 118.83 150.02 118.83 150.02 118.59 149.65 118.59 149.65 118.52 149.51 118.52 149.51 118.9 149.65 118.9 ;
      RECT  152.63 118.28 152.42 118.04 ;
      RECT  152.42 118.28 150.02 118.04 ;
      RECT  150.02 119.38 149.51 119.14 ;
      RECT  151.49 120.17 150.95 119.62 ;
      RECT  152.63 120.89 151.49 121.27 ;
      RECT  150.23 120.65 150.02 120.72 ;
      RECT  150.02 121.51 149.51 121.75 ;
      RECT  152.42 120.41 150.02 120.65 ;
      RECT  150.02 120.65 149.82 120.72 ;
      RECT  150.23 121.44 150.02 121.51 ;
      RECT  149.51 120.41 149.3 120.65 ;
      POLYGON  150.95 120.89 150.95 121.27 150.4 121.27 150.4 121.2 150.02 121.2 150.02 120.96 150.4 120.96 150.4 120.89 150.95 120.89 ;
      RECT  149.51 120.89 149.3 121.27 ;
      RECT  152.63 119.62 152.42 120.17 ;
      RECT  152.42 119.62 151.49 120.17 ;
      RECT  151.49 120.89 150.95 121.27 ;
      RECT  149.51 121.51 149.3 121.75 ;
      RECT  150.95 119.62 149.3 120.17 ;
      RECT  152.63 120.41 152.42 120.65 ;
      RECT  150.02 121.44 149.82 121.51 ;
      POLYGON  149.65 120.89 149.65 120.96 150.02 120.96 150.02 121.2 149.65 121.2 149.65 121.27 149.51 121.27 149.51 120.89 149.65 120.89 ;
      RECT  152.63 121.51 152.42 121.75 ;
      RECT  152.42 121.51 150.02 121.75 ;
      RECT  150.02 120.41 149.51 120.65 ;
      RECT  151.49 119.62 150.95 120.17 ;
      RECT  152.63 122.85 151.49 122.47 ;
      RECT  150.23 123.09 150.02 123.02 ;
      RECT  150.02 122.23 149.51 121.99 ;
      RECT  152.42 123.33 150.02 123.09 ;
      RECT  150.02 123.09 149.82 123.02 ;
      RECT  150.23 122.3 150.02 122.23 ;
      RECT  149.51 123.33 149.3 123.09 ;
      POLYGON  150.95 122.85 150.95 122.47 150.4 122.47 150.4 122.54 150.02 122.54 150.02 122.78 150.4 122.78 150.4 122.85 150.95 122.85 ;
      RECT  149.51 122.85 149.3 122.47 ;
      RECT  152.63 124.12 152.42 123.57 ;
      RECT  152.42 124.12 151.49 123.57 ;
      RECT  151.49 122.85 150.95 122.47 ;
      RECT  149.51 122.23 149.3 121.99 ;
      RECT  150.95 124.12 149.3 123.57 ;
      RECT  152.63 123.33 152.42 123.09 ;
      RECT  150.02 122.3 149.82 122.23 ;
      POLYGON  149.65 122.85 149.65 122.78 150.02 122.78 150.02 122.54 149.65 122.54 149.65 122.47 149.51 122.47 149.51 122.85 149.65 122.85 ;
      RECT  152.63 122.23 152.42 121.99 ;
      RECT  152.42 122.23 150.02 121.99 ;
      RECT  150.02 123.33 149.51 123.09 ;
      RECT  151.49 124.12 150.95 123.57 ;
      RECT  152.63 124.84 151.49 125.22 ;
      RECT  150.23 124.6 150.02 124.67 ;
      RECT  150.02 125.46 149.51 125.7 ;
      RECT  152.42 124.36 150.02 124.6 ;
      RECT  150.02 124.6 149.82 124.67 ;
      RECT  150.23 125.39 150.02 125.46 ;
      RECT  149.51 124.36 149.3 124.6 ;
      POLYGON  150.95 124.84 150.95 125.22 150.4 125.22 150.4 125.15 150.02 125.15 150.02 124.91 150.4 124.91 150.4 124.84 150.95 124.84 ;
      RECT  149.51 124.84 149.3 125.22 ;
      RECT  152.63 123.57 152.42 124.12 ;
      RECT  152.42 123.57 151.49 124.12 ;
      RECT  151.49 124.84 150.95 125.22 ;
      RECT  149.51 125.46 149.3 125.7 ;
      RECT  150.95 123.57 149.3 124.12 ;
      RECT  152.63 124.36 152.42 124.6 ;
      RECT  150.02 125.39 149.82 125.46 ;
      POLYGON  149.65 124.84 149.65 124.91 150.02 124.91 150.02 125.15 149.65 125.15 149.65 125.22 149.51 125.22 149.51 124.84 149.65 124.84 ;
      RECT  152.63 125.46 152.42 125.7 ;
      RECT  152.42 125.46 150.02 125.7 ;
      RECT  150.02 124.36 149.51 124.6 ;
      RECT  151.49 123.57 150.95 124.12 ;
      RECT  149.3 90.39 152.42 90.63 ;
      RECT  149.3 91.49 152.42 91.73 ;
      RECT  149.3 93.86 152.42 94.1 ;
      RECT  149.3 92.76 152.42 93.0 ;
      RECT  149.3 94.34 152.42 94.58 ;
      RECT  149.3 95.44 152.42 95.68 ;
      RECT  149.3 97.81 152.42 98.05 ;
      RECT  149.3 96.71 152.42 96.95 ;
      RECT  149.3 98.29 152.42 98.53 ;
      RECT  149.3 99.39 152.42 99.63 ;
      RECT  149.3 101.76 152.42 102.0 ;
      RECT  149.3 100.66 152.42 100.9 ;
      RECT  149.3 102.24 152.42 102.48 ;
      RECT  149.3 103.34 152.42 103.58 ;
      RECT  149.3 105.71 152.42 105.95 ;
      RECT  149.3 104.61 152.42 104.85 ;
      RECT  149.3 106.19 152.42 106.43 ;
      RECT  149.3 107.29 152.42 107.53 ;
      RECT  149.3 109.66 152.42 109.9 ;
      RECT  149.3 108.56 152.42 108.8 ;
      RECT  149.3 110.14 152.42 110.38 ;
      RECT  149.3 111.24 152.42 111.48 ;
      RECT  149.3 113.61 152.42 113.85 ;
      RECT  149.3 112.51 152.42 112.75 ;
      RECT  149.3 114.09 152.42 114.33 ;
      RECT  149.3 115.19 152.42 115.43 ;
      RECT  149.3 117.56 152.42 117.8 ;
      RECT  149.3 116.46 152.42 116.7 ;
      RECT  149.3 118.04 152.42 118.28 ;
      RECT  149.3 119.14 152.42 119.38 ;
      RECT  149.3 121.51 152.42 121.75 ;
      RECT  149.3 120.41 152.42 120.65 ;
      RECT  149.3 121.99 152.42 122.23 ;
      RECT  149.3 123.09 152.42 123.33 ;
      RECT  149.3 125.46 152.42 125.7 ;
      RECT  149.3 124.36 152.42 124.6 ;
      RECT  90.02 93.86 152.42 94.1 ;
      RECT  90.02 92.76 152.42 93.0 ;
      RECT  90.02 94.34 152.42 94.58 ;
      RECT  90.02 95.44 152.42 95.68 ;
      RECT  90.02 97.81 152.42 98.05 ;
      RECT  90.02 96.71 152.42 96.95 ;
      RECT  90.02 98.29 152.42 98.53 ;
      RECT  90.02 99.39 152.42 99.63 ;
      RECT  90.02 101.76 152.42 102.0 ;
      RECT  90.02 100.66 152.42 100.9 ;
      RECT  90.02 102.24 152.42 102.48 ;
      RECT  90.02 103.34 152.42 103.58 ;
      RECT  90.02 105.71 152.42 105.95 ;
      RECT  90.02 104.61 152.42 104.85 ;
      RECT  90.02 106.19 152.42 106.43 ;
      RECT  90.02 107.29 152.42 107.53 ;
      RECT  90.02 109.66 152.42 109.9 ;
      RECT  90.02 108.56 152.42 108.8 ;
      RECT  90.02 110.14 152.42 110.38 ;
      RECT  90.02 111.24 152.42 111.48 ;
      RECT  90.02 113.61 152.42 113.85 ;
      RECT  90.02 112.51 152.42 112.75 ;
      RECT  90.02 114.09 152.42 114.33 ;
      RECT  90.02 115.19 152.42 115.43 ;
      RECT  90.02 117.56 152.42 117.8 ;
      RECT  90.02 116.46 152.42 116.7 ;
      RECT  90.02 118.04 152.42 118.28 ;
      RECT  90.02 119.14 152.42 119.38 ;
      RECT  90.02 121.51 152.42 121.75 ;
      RECT  90.02 120.41 152.42 120.65 ;
      RECT  90.02 121.99 152.42 122.23 ;
      RECT  90.02 123.09 152.42 123.33 ;
      RECT  90.02 90.39 152.42 90.63 ;
      RECT  90.02 124.36 152.42 124.6 ;
      RECT  94.79 106.67 95.33 107.05 ;
      RECT  147.11 101.14 147.65 101.52 ;
      RECT  94.79 123.57 95.33 124.12 ;
      RECT  147.11 103.82 147.65 104.37 ;
      RECT  94.79 112.99 95.33 113.37 ;
      RECT  147.11 122.47 147.65 122.85 ;
      RECT  94.79 101.14 95.33 101.52 ;
      RECT  147.11 118.52 147.65 118.9 ;
      RECT  94.79 93.24 95.33 93.62 ;
      RECT  94.79 102.72 95.33 103.1 ;
      RECT  147.11 102.72 147.65 103.1 ;
      RECT  147.11 94.82 147.65 95.2 ;
      RECT  147.11 90.87 147.65 91.25 ;
      RECT  147.11 93.24 147.65 93.62 ;
      RECT  147.11 112.99 147.65 113.37 ;
      RECT  147.11 106.67 147.65 107.05 ;
      RECT  94.79 107.77 95.33 108.32 ;
      RECT  94.79 119.62 95.33 120.17 ;
      RECT  94.79 91.97 95.33 92.52 ;
      RECT  147.11 123.57 147.65 124.12 ;
      RECT  94.79 105.09 95.33 105.47 ;
      RECT  94.79 115.67 95.33 116.22 ;
      RECT  94.79 109.04 95.33 109.42 ;
      RECT  94.79 95.92 95.33 96.47 ;
      RECT  94.79 118.52 95.33 118.9 ;
      RECT  94.79 90.87 95.33 91.25 ;
      RECT  147.11 109.04 147.65 109.42 ;
      RECT  94.79 122.47 95.33 122.85 ;
      RECT  147.11 114.57 147.65 114.95 ;
      RECT  147.11 116.94 147.65 117.32 ;
      RECT  147.11 120.89 147.65 121.27 ;
      RECT  147.11 119.62 147.65 120.17 ;
      RECT  94.79 103.82 95.33 104.37 ;
      RECT  147.11 95.92 147.65 96.47 ;
      RECT  94.79 110.62 95.33 111.0 ;
      RECT  94.79 99.87 95.33 100.42 ;
      RECT  94.79 116.94 95.33 117.32 ;
      RECT  147.11 91.97 147.65 92.52 ;
      RECT  147.11 98.77 147.65 99.15 ;
      RECT  94.79 111.72 95.33 112.27 ;
      RECT  94.79 98.77 95.33 99.15 ;
      RECT  147.11 111.72 147.65 112.27 ;
      RECT  94.79 120.89 95.33 121.27 ;
      RECT  94.79 97.19 95.33 97.57 ;
      RECT  94.79 94.82 95.33 95.2 ;
      RECT  147.11 97.19 147.65 97.57 ;
      RECT  147.11 110.62 147.65 111.0 ;
      RECT  94.79 124.84 95.33 125.22 ;
      RECT  94.79 114.57 95.33 114.95 ;
      RECT  147.11 124.84 147.65 125.22 ;
      RECT  147.11 99.87 147.65 100.42 ;
      RECT  147.11 115.67 147.65 116.22 ;
      RECT  147.11 105.09 147.65 105.47 ;
      RECT  147.11 107.77 147.65 108.32 ;
      RECT  96.26 83.32 93.14 83.46 ;
      RECT  96.26 83.32 99.38 83.46 ;
      RECT  102.5 83.32 99.38 83.46 ;
      RECT  102.5 83.32 105.62 83.46 ;
      RECT  108.74 83.32 105.62 83.46 ;
      RECT  108.74 83.32 111.86 83.46 ;
      RECT  114.98 83.32 111.86 83.46 ;
      RECT  114.98 83.32 118.1 83.46 ;
      RECT  121.22 83.32 118.1 83.46 ;
      RECT  121.22 83.32 124.34 83.46 ;
      RECT  127.46 83.32 124.34 83.46 ;
      RECT  127.46 83.32 130.58 83.46 ;
      RECT  133.7 83.32 130.58 83.46 ;
      RECT  133.7 83.32 136.82 83.46 ;
      RECT  139.94 83.32 136.82 83.46 ;
      RECT  139.94 83.32 143.06 83.46 ;
      RECT  146.18 83.32 143.06 83.46 ;
      RECT  96.19 53.83 96.33 53.97 ;
      RECT  121.15 53.83 121.29 53.97 ;
      RECT  96.19 53.97 96.33 53.83 ;
      RECT  121.15 53.97 121.29 53.83 ;
      RECT  96.26 132.77 99.38 132.63 ;
      RECT  102.5 132.77 99.38 132.63 ;
      RECT  102.5 132.77 105.62 132.63 ;
      RECT  108.74 132.77 105.62 132.63 ;
      RECT  108.74 132.77 111.86 132.63 ;
      RECT  114.98 132.77 111.86 132.63 ;
      RECT  114.98 132.77 118.1 132.63 ;
      RECT  121.22 132.77 118.1 132.63 ;
      RECT  121.22 132.77 124.34 132.63 ;
      RECT  127.46 132.77 124.34 132.63 ;
      RECT  127.46 132.77 130.58 132.63 ;
      RECT  133.7 132.77 130.58 132.63 ;
      RECT  133.7 132.77 136.82 132.63 ;
      RECT  139.94 132.77 136.82 132.63 ;
      RECT  139.94 132.77 143.06 132.63 ;
      RECT  146.18 132.77 143.06 132.63 ;
      RECT  146.18 132.77 149.3 132.63 ;
      RECT  68.94 92.245 69.08 123.845 ;
      RECT  68.94 92.245 69.08 123.845 ;
      RECT  173.5 92.245 173.36 123.845 ;
      RECT  173.5 92.245 173.36 123.845 ;
      RECT  86.92 52.55 87.06 91.445 ;
      RECT  154.28 124.645 154.42 145.785 ;
      RECT  88.16 52.55 88.3 91.445 ;
      RECT  153.66 124.645 153.8 145.785 ;
      RECT  87.54 52.55 87.68 91.445 ;
      RECT  96.19 53.83 96.33 53.97 ;
      RECT  121.15 53.83 121.29 53.97 ;
      RECT  88.78 52.55 88.92 91.445 ;
      RECT  153.04 124.645 153.18 145.785 ;
      RECT  1.305 33.625 1.635 33.885 ;
      RECT  6.03 33.98 6.36 34.24 ;
      RECT  5.64 33.225 5.97 33.485 ;
      RECT  2.465 34.395 2.735 34.715 ;
      RECT  1.305 33.625 1.635 33.885 ;
      RECT  10.99 33.3 11.13 33.44 ;
      RECT  8.46 35.105 8.6 35.245 ;
      RECT  2.465 34.395 2.735 34.715 ;
      RECT  1.305 42.385 1.635 42.125 ;
      RECT  6.03 42.03 6.36 41.77 ;
      RECT  5.64 42.785 5.97 42.525 ;
      RECT  2.465 41.615 2.735 41.295 ;
      RECT  1.305 42.385 1.635 42.125 ;
      RECT  10.99 42.71 11.13 42.57 ;
      RECT  8.46 40.905 8.6 40.765 ;
      RECT  2.465 41.615 2.735 41.295 ;
      RECT  1.305 33.625 1.635 33.885 ;
      RECT  1.305 42.125 1.635 42.385 ;
      RECT  10.99 33.3 11.13 33.44 ;
      RECT  8.46 35.105 8.6 35.245 ;
      RECT  10.99 42.57 11.13 42.71 ;
      RECT  8.46 40.765 8.6 40.905 ;
      RECT  2.465 30.935 2.605 45.075 ;
      RECT  9.5 88.295 9.36 90.905 ;
      RECT  1.705 88.295 1.565 135.705 ;
      RECT  1.305 33.625 1.635 33.885 ;
      RECT  1.305 42.125 1.635 42.385 ;
      RECT  16.055 34.21 16.195 34.35 ;
      RECT  9.36 88.295 9.5 90.905 ;
      RECT  21.26 83.89 40.15 84.03 ;
      RECT  22.34 62.68 40.15 62.82 ;
      RECT  24.55 69.75 40.15 69.89 ;
      RECT  22.21 55.61 40.15 55.75 ;
      RECT  34.0 34.4 40.15 34.54 ;
      RECT  240.055 168.325 239.725 168.065 ;
      RECT  235.33 167.97 235.0 167.71 ;
      RECT  235.72 168.725 235.39 168.465 ;
      RECT  238.895 167.555 238.625 167.235 ;
      RECT  240.055 168.325 239.725 168.065 ;
      RECT  230.37 168.65 230.23 168.51 ;
      RECT  232.9 166.845 232.76 166.705 ;
      RECT  238.895 167.555 238.625 167.235 ;
      RECT  240.055 168.325 239.725 168.065 ;
      RECT  230.37 168.65 230.23 168.51 ;
      RECT  232.9 166.845 232.76 166.705 ;
      RECT  238.895 171.015 238.755 163.945 ;
      RECT  231.86 127.795 232.0 125.185 ;
      RECT  239.655 127.795 239.795 80.385 ;
      RECT  240.055 168.325 239.725 168.065 ;
      RECT  225.725 167.74 225.585 167.6 ;
      RECT  232.0 127.795 231.86 125.185 ;
      RECT  220.52 132.2 202.71 132.06 ;
      RECT  217.23 139.27 202.71 139.13 ;
      RECT  219.57 146.34 202.71 146.2 ;
      RECT  208.82 167.55 202.71 167.41 ;
      RECT  34.995 142.185 35.325 142.445 ;
      RECT  39.72 142.54 40.05 142.8 ;
      RECT  39.33 141.785 39.66 142.045 ;
      RECT  36.155 142.955 36.425 143.275 ;
      RECT  34.995 150.945 35.325 150.685 ;
      RECT  39.72 150.59 40.05 150.33 ;
      RECT  39.33 151.345 39.66 151.085 ;
      RECT  36.155 150.175 36.425 149.855 ;
      RECT  34.995 156.325 35.325 156.585 ;
      RECT  39.72 156.68 40.05 156.94 ;
      RECT  39.33 155.925 39.66 156.185 ;
      RECT  36.155 157.095 36.425 157.415 ;
      RECT  34.995 165.085 35.325 164.825 ;
      RECT  39.72 164.73 40.05 164.47 ;
      RECT  39.33 165.485 39.66 165.225 ;
      RECT  36.155 164.315 36.425 163.995 ;
      RECT  34.995 142.185 35.325 142.445 ;
      RECT  34.995 150.685 35.325 150.945 ;
      RECT  34.995 156.325 35.325 156.585 ;
      RECT  34.995 164.825 35.325 165.085 ;
      RECT  39.72 142.54 40.05 142.8 ;
      RECT  39.72 150.33 40.05 150.59 ;
      RECT  39.72 156.68 40.05 156.94 ;
      RECT  39.72 164.47 40.05 164.73 ;
      RECT  207.865 73.905 207.535 73.645 ;
      RECT  203.14 73.55 202.81 73.29 ;
      RECT  203.53 74.305 203.2 74.045 ;
      RECT  206.705 73.135 206.435 72.815 ;
      RECT  207.865 65.145 207.535 65.405 ;
      RECT  203.14 65.5 202.81 65.76 ;
      RECT  203.53 64.745 203.2 65.005 ;
      RECT  206.705 65.915 206.435 66.235 ;
      RECT  207.865 59.765 207.535 59.505 ;
      RECT  203.14 59.41 202.81 59.15 ;
      RECT  203.53 60.165 203.2 59.905 ;
      RECT  206.705 58.995 206.435 58.675 ;
      RECT  207.865 51.005 207.535 51.265 ;
      RECT  203.14 51.36 202.81 51.62 ;
      RECT  203.53 50.605 203.2 50.865 ;
      RECT  206.705 51.775 206.435 52.095 ;
      RECT  207.865 73.905 207.535 73.645 ;
      RECT  207.865 65.405 207.535 65.145 ;
      RECT  207.865 59.765 207.535 59.505 ;
      RECT  207.865 51.265 207.535 51.005 ;
      RECT  203.14 73.55 202.81 73.29 ;
      RECT  203.14 65.76 202.81 65.5 ;
      RECT  203.14 59.41 202.81 59.15 ;
      RECT  203.14 51.62 202.81 51.36 ;
      RECT  46.675 3.03 47.005 3.29 ;
      RECT  51.4 3.385 51.73 3.645 ;
      RECT  51.01 2.63 51.34 2.89 ;
      RECT  47.835 3.8 48.105 4.12 ;
      RECT  52.515 3.03 52.845 3.29 ;
      RECT  57.24 3.385 57.57 3.645 ;
      RECT  56.85 2.63 57.18 2.89 ;
      RECT  53.675 3.8 53.945 4.12 ;
      RECT  46.675 3.03 47.005 3.29 ;
      RECT  52.515 3.03 52.845 3.29 ;
      RECT  51.4 3.385 51.73 3.645 ;
      RECT  57.24 3.385 57.57 3.645 ;
      RECT  58.355 3.03 58.685 3.29 ;
      RECT  63.08 3.385 63.41 3.645 ;
      RECT  62.69 2.63 63.02 2.89 ;
      RECT  59.515 3.8 59.785 4.12 ;
      RECT  64.195 3.03 64.525 3.29 ;
      RECT  68.92 3.385 69.25 3.645 ;
      RECT  68.53 2.63 68.86 2.89 ;
      RECT  65.355 3.8 65.625 4.12 ;
      RECT  70.035 3.03 70.365 3.29 ;
      RECT  74.76 3.385 75.09 3.645 ;
      RECT  74.37 2.63 74.7 2.89 ;
      RECT  71.195 3.8 71.465 4.12 ;
      RECT  75.875 3.03 76.205 3.29 ;
      RECT  80.6 3.385 80.93 3.645 ;
      RECT  80.21 2.63 80.54 2.89 ;
      RECT  77.035 3.8 77.305 4.12 ;
      RECT  81.715 3.03 82.045 3.29 ;
      RECT  86.44 3.385 86.77 3.645 ;
      RECT  86.05 2.63 86.38 2.89 ;
      RECT  82.875 3.8 83.145 4.12 ;
      RECT  87.555 3.03 87.885 3.29 ;
      RECT  92.28 3.385 92.61 3.645 ;
      RECT  91.89 2.63 92.22 2.89 ;
      RECT  88.715 3.8 88.985 4.12 ;
      RECT  93.395 3.03 93.725 3.29 ;
      RECT  98.12 3.385 98.45 3.645 ;
      RECT  97.73 2.63 98.06 2.89 ;
      RECT  94.555 3.8 94.825 4.12 ;
      RECT  99.235 3.03 99.565 3.29 ;
      RECT  103.96 3.385 104.29 3.645 ;
      RECT  103.57 2.63 103.9 2.89 ;
      RECT  100.395 3.8 100.665 4.12 ;
      RECT  105.075 3.03 105.405 3.29 ;
      RECT  109.8 3.385 110.13 3.645 ;
      RECT  109.41 2.63 109.74 2.89 ;
      RECT  106.235 3.8 106.505 4.12 ;
      RECT  110.915 3.03 111.245 3.29 ;
      RECT  115.64 3.385 115.97 3.645 ;
      RECT  115.25 2.63 115.58 2.89 ;
      RECT  112.075 3.8 112.345 4.12 ;
      RECT  116.755 3.03 117.085 3.29 ;
      RECT  121.48 3.385 121.81 3.645 ;
      RECT  121.09 2.63 121.42 2.89 ;
      RECT  117.915 3.8 118.185 4.12 ;
      RECT  122.595 3.03 122.925 3.29 ;
      RECT  127.32 3.385 127.65 3.645 ;
      RECT  126.93 2.63 127.26 2.89 ;
      RECT  123.755 3.8 124.025 4.12 ;
      RECT  128.435 3.03 128.765 3.29 ;
      RECT  133.16 3.385 133.49 3.645 ;
      RECT  132.77 2.63 133.1 2.89 ;
      RECT  129.595 3.8 129.865 4.12 ;
      RECT  134.275 3.03 134.605 3.29 ;
      RECT  139.0 3.385 139.33 3.645 ;
      RECT  138.61 2.63 138.94 2.89 ;
      RECT  135.435 3.8 135.705 4.12 ;
      RECT  140.115 3.03 140.445 3.29 ;
      RECT  144.84 3.385 145.17 3.645 ;
      RECT  144.45 2.63 144.78 2.89 ;
      RECT  141.275 3.8 141.545 4.12 ;
      RECT  145.955 3.03 146.285 3.29 ;
      RECT  150.68 3.385 151.01 3.645 ;
      RECT  150.29 2.63 150.62 2.89 ;
      RECT  147.115 3.8 147.385 4.12 ;
      RECT  58.355 3.03 58.685 3.29 ;
      RECT  64.195 3.03 64.525 3.29 ;
      RECT  70.035 3.03 70.365 3.29 ;
      RECT  75.875 3.03 76.205 3.29 ;
      RECT  81.715 3.03 82.045 3.29 ;
      RECT  87.555 3.03 87.885 3.29 ;
      RECT  93.395 3.03 93.725 3.29 ;
      RECT  99.235 3.03 99.565 3.29 ;
      RECT  105.075 3.03 105.405 3.29 ;
      RECT  110.915 3.03 111.245 3.29 ;
      RECT  116.755 3.03 117.085 3.29 ;
      RECT  122.595 3.03 122.925 3.29 ;
      RECT  128.435 3.03 128.765 3.29 ;
      RECT  134.275 3.03 134.605 3.29 ;
      RECT  140.115 3.03 140.445 3.29 ;
      RECT  145.955 3.03 146.285 3.29 ;
      RECT  63.08 3.385 63.41 3.645 ;
      RECT  68.92 3.385 69.25 3.645 ;
      RECT  74.76 3.385 75.09 3.645 ;
      RECT  80.6 3.385 80.93 3.645 ;
      RECT  86.44 3.385 86.77 3.645 ;
      RECT  92.28 3.385 92.61 3.645 ;
      RECT  98.12 3.385 98.45 3.645 ;
      RECT  103.96 3.385 104.29 3.645 ;
      RECT  109.8 3.385 110.13 3.645 ;
      RECT  115.64 3.385 115.97 3.645 ;
      RECT  121.48 3.385 121.81 3.645 ;
      RECT  127.32 3.385 127.65 3.645 ;
      RECT  133.16 3.385 133.49 3.645 ;
      RECT  139.0 3.385 139.33 3.645 ;
      RECT  144.84 3.385 145.17 3.645 ;
      RECT  150.68 3.385 151.01 3.645 ;
   LAYER  m3 ;
      RECT  94.455 126.405 94.945 126.895 ;
      RECT  94.455 89.195 94.945 89.685 ;
      RECT  147.495 126.405 147.985 126.895 ;
      RECT  147.495 89.195 147.985 89.685 ;
      RECT  103.815 89.195 104.305 89.685 ;
      RECT  106.935 89.195 107.425 89.685 ;
      RECT  128.775 89.195 129.265 89.685 ;
      RECT  138.135 89.195 138.625 89.685 ;
      RECT  141.255 89.195 141.745 89.685 ;
      RECT  135.015 89.195 135.505 89.685 ;
      RECT  125.655 89.195 126.145 89.685 ;
      RECT  144.375 89.195 144.865 89.685 ;
      RECT  97.575 89.195 98.065 89.685 ;
      RECT  110.055 89.195 110.545 89.685 ;
      RECT  119.415 89.195 119.905 89.685 ;
      RECT  100.695 89.195 101.185 89.685 ;
      RECT  131.895 89.195 132.385 89.685 ;
      RECT  113.175 89.195 113.665 89.685 ;
      RECT  116.295 89.195 116.785 89.685 ;
      RECT  122.535 89.195 123.025 89.685 ;
      RECT  103.815 126.895 104.305 126.405 ;
      RECT  106.935 126.895 107.425 126.405 ;
      RECT  128.775 126.895 129.265 126.405 ;
      RECT  138.135 126.895 138.625 126.405 ;
      RECT  141.255 126.895 141.745 126.405 ;
      RECT  135.015 126.895 135.505 126.405 ;
      RECT  125.655 126.895 126.145 126.405 ;
      RECT  144.375 126.895 144.865 126.405 ;
      RECT  97.575 126.895 98.065 126.405 ;
      RECT  110.055 126.895 110.545 126.405 ;
      RECT  119.415 126.895 119.905 126.405 ;
      RECT  100.695 126.895 101.185 126.405 ;
      RECT  131.895 126.895 132.385 126.405 ;
      RECT  113.175 126.895 113.665 126.405 ;
      RECT  116.295 126.895 116.785 126.405 ;
      RECT  122.535 126.895 123.025 126.405 ;
      RECT  90.975 119.65 91.465 120.14 ;
      RECT  90.975 105.035 91.465 105.525 ;
      RECT  90.975 98.715 91.465 99.205 ;
      RECT  90.975 99.9 91.465 100.39 ;
      RECT  90.975 112.935 91.465 113.425 ;
      RECT  90.975 101.085 91.465 101.575 ;
      RECT  90.975 124.785 91.465 125.275 ;
      RECT  90.975 111.75 91.465 112.24 ;
      RECT  90.975 116.885 91.465 117.375 ;
      RECT  90.975 95.95 91.465 96.44 ;
      RECT  90.975 102.665 91.465 103.155 ;
      RECT  90.975 107.8 91.465 108.29 ;
      RECT  90.975 94.765 91.465 95.255 ;
      RECT  90.975 90.815 91.465 91.305 ;
      RECT  90.975 93.185 91.465 93.675 ;
      RECT  90.975 108.985 91.465 109.475 ;
      RECT  90.975 103.85 91.465 104.34 ;
      RECT  90.975 97.135 91.465 97.625 ;
      RECT  90.975 118.465 91.465 118.955 ;
      RECT  90.975 120.835 91.465 121.325 ;
      RECT  90.975 106.615 91.465 107.105 ;
      RECT  90.975 114.515 91.465 115.005 ;
      RECT  90.975 122.415 91.465 122.905 ;
      RECT  90.975 123.6 91.465 124.09 ;
      RECT  90.975 110.565 91.465 111.055 ;
      RECT  90.975 115.7 91.465 116.19 ;
      RECT  90.975 92.0 91.465 92.49 ;
      RECT  150.975 98.715 151.465 99.205 ;
      RECT  150.975 107.8 151.465 108.29 ;
      RECT  150.975 119.65 151.465 120.14 ;
      RECT  150.975 103.85 151.465 104.34 ;
      RECT  150.975 118.465 151.465 118.955 ;
      RECT  150.975 116.885 151.465 117.375 ;
      RECT  150.975 92.0 151.465 92.49 ;
      RECT  150.975 108.985 151.465 109.475 ;
      RECT  150.975 93.185 151.465 93.675 ;
      RECT  150.975 120.835 151.465 121.325 ;
      RECT  150.975 112.935 151.465 113.425 ;
      RECT  150.975 97.135 151.465 97.625 ;
      RECT  150.975 124.785 151.465 125.275 ;
      RECT  150.975 94.765 151.465 95.255 ;
      RECT  150.975 99.9 151.465 100.39 ;
      RECT  150.975 106.615 151.465 107.105 ;
      RECT  150.975 115.7 151.465 116.19 ;
      RECT  150.975 123.6 151.465 124.09 ;
      RECT  150.975 101.085 151.465 101.575 ;
      RECT  150.975 102.665 151.465 103.155 ;
      RECT  150.975 114.515 151.465 115.005 ;
      RECT  150.975 105.035 151.465 105.525 ;
      RECT  150.975 111.75 151.465 112.24 ;
      RECT  150.975 122.415 151.465 122.905 ;
      RECT  150.975 90.815 151.465 91.305 ;
      RECT  150.975 110.565 151.465 111.055 ;
      RECT  150.975 95.95 151.465 96.44 ;
      RECT  141.35 126.5 141.65 126.8 ;
      RECT  100.79 89.29 101.09 89.59 ;
      RECT  122.63 126.5 122.93 126.8 ;
      RECT  110.15 89.29 110.45 89.59 ;
      RECT  97.67 126.5 97.97 126.8 ;
      RECT  107.03 126.5 107.33 126.8 ;
      RECT  138.23 89.29 138.53 89.59 ;
      RECT  138.23 126.5 138.53 126.8 ;
      RECT  116.39 89.29 116.69 89.59 ;
      RECT  144.47 126.5 144.77 126.8 ;
      RECT  141.35 89.29 141.65 89.59 ;
      RECT  131.99 89.29 132.29 89.59 ;
      RECT  135.11 89.29 135.41 89.59 ;
      RECT  147.495 89.195 147.985 89.685 ;
      RECT  147.495 126.405 147.985 126.895 ;
      RECT  128.87 89.29 129.17 89.59 ;
      RECT  128.87 126.5 129.17 126.8 ;
      RECT  119.51 126.5 119.81 126.8 ;
      RECT  135.11 126.5 135.41 126.8 ;
      RECT  103.91 126.5 104.21 126.8 ;
      RECT  119.51 89.29 119.81 89.59 ;
      RECT  94.455 126.405 94.945 126.895 ;
      RECT  113.27 89.29 113.57 89.59 ;
      RECT  97.67 89.29 97.97 89.59 ;
      RECT  100.79 126.5 101.09 126.8 ;
      RECT  94.455 89.195 94.945 89.685 ;
      RECT  125.75 89.29 126.05 89.59 ;
      RECT  113.27 126.5 113.57 126.8 ;
      RECT  144.47 89.29 144.77 89.59 ;
      RECT  122.63 89.29 122.93 89.59 ;
      RECT  116.39 126.5 116.69 126.8 ;
      RECT  110.15 126.5 110.45 126.8 ;
      RECT  125.75 126.5 126.05 126.8 ;
      RECT  131.99 126.5 132.29 126.8 ;
      RECT  107.03 89.29 107.33 89.59 ;
      RECT  103.91 89.29 104.21 89.59 ;
      RECT  91.07 122.51 91.37 122.81 ;
      RECT  151.07 122.51 151.37 122.81 ;
      RECT  151.07 109.08 151.37 109.38 ;
      RECT  91.07 94.86 91.37 95.16 ;
      RECT  151.07 120.93 151.37 121.23 ;
      RECT  151.07 103.945 151.37 104.245 ;
      RECT  91.07 99.995 91.37 100.295 ;
      RECT  151.07 94.86 151.37 95.16 ;
      RECT  151.07 106.71 151.37 107.01 ;
      RECT  151.07 118.56 151.37 118.86 ;
      RECT  151.07 115.795 151.37 116.095 ;
      RECT  91.07 118.56 91.37 118.86 ;
      RECT  91.07 98.81 91.37 99.11 ;
      RECT  151.07 113.03 151.37 113.33 ;
      RECT  91.07 116.98 91.37 117.28 ;
      RECT  151.07 92.095 151.37 92.395 ;
      RECT  151.07 114.61 151.37 114.91 ;
      RECT  151.07 119.745 151.37 120.045 ;
      RECT  91.07 92.095 91.37 92.395 ;
      RECT  151.07 116.98 151.37 117.28 ;
      RECT  91.07 103.945 91.37 104.245 ;
      RECT  91.07 105.13 91.37 105.43 ;
      RECT  91.07 111.845 91.37 112.145 ;
      RECT  91.07 114.61 91.37 114.91 ;
      RECT  91.07 96.045 91.37 96.345 ;
      RECT  91.07 97.23 91.37 97.53 ;
      RECT  151.07 111.845 151.37 112.145 ;
      RECT  151.07 97.23 151.37 97.53 ;
      RECT  151.07 90.91 151.37 91.21 ;
      RECT  91.07 119.745 91.37 120.045 ;
      RECT  91.07 90.91 91.37 91.21 ;
      RECT  151.07 105.13 151.37 105.43 ;
      RECT  91.07 107.895 91.37 108.195 ;
      RECT  151.07 96.045 151.37 96.345 ;
      RECT  151.07 102.76 151.37 103.06 ;
      RECT  151.07 110.66 151.37 110.96 ;
      RECT  91.07 101.18 91.37 101.48 ;
      RECT  151.07 93.28 151.37 93.58 ;
      RECT  91.07 109.08 91.37 109.38 ;
      RECT  91.07 106.71 91.37 107.01 ;
      RECT  91.07 120.93 91.37 121.23 ;
      RECT  91.07 124.88 91.37 125.18 ;
      RECT  151.07 123.695 151.37 123.995 ;
      RECT  91.07 93.28 91.37 93.58 ;
      RECT  91.07 113.03 91.37 113.33 ;
      RECT  91.07 102.76 91.37 103.06 ;
      RECT  151.07 101.18 151.37 101.48 ;
      RECT  151.07 99.995 151.37 100.295 ;
      RECT  91.07 123.695 91.37 123.995 ;
      RECT  91.07 110.66 91.37 110.96 ;
      RECT  91.07 115.795 91.37 116.095 ;
      RECT  151.07 107.895 151.37 108.195 ;
      RECT  151.07 98.81 151.37 99.11 ;
      RECT  151.07 124.88 151.37 125.18 ;
      RECT  95.54 86.24 95.05 86.73 ;
      RECT  96.98 86.24 97.47 86.73 ;
      RECT  101.78 86.24 101.29 86.73 ;
      RECT  103.22 86.24 103.71 86.73 ;
      RECT  108.02 86.24 107.53 86.73 ;
      RECT  109.46 86.24 109.95 86.73 ;
      RECT  114.26 86.24 113.77 86.73 ;
      RECT  115.7 86.24 116.19 86.73 ;
      RECT  120.5 86.24 120.01 86.73 ;
      RECT  121.94 86.24 122.43 86.73 ;
      RECT  126.74 86.24 126.25 86.73 ;
      RECT  128.18 86.24 128.67 86.73 ;
      RECT  132.98 86.24 132.49 86.73 ;
      RECT  134.42 86.24 134.91 86.73 ;
      RECT  139.22 86.24 138.73 86.73 ;
      RECT  140.66 86.24 141.15 86.73 ;
      RECT  145.46 86.24 144.97 86.73 ;
      RECT  93.14 83.24 146.18 83.54 ;
      RECT  134.42 86.24 134.91 86.73 ;
      RECT  95.05 86.24 95.54 86.73 ;
      RECT  101.29 86.24 101.78 86.73 ;
      RECT  103.22 86.24 103.71 86.73 ;
      RECT  113.77 86.24 114.26 86.73 ;
      RECT  144.97 86.24 145.46 86.73 ;
      RECT  126.25 86.24 126.74 86.73 ;
      RECT  121.94 86.24 122.43 86.73 ;
      RECT  96.98 86.24 97.47 86.73 ;
      RECT  109.46 86.24 109.95 86.73 ;
      RECT  115.7 86.24 116.19 86.73 ;
      RECT  120.01 86.24 120.5 86.73 ;
      RECT  107.53 86.24 108.02 86.73 ;
      RECT  132.49 86.24 132.98 86.73 ;
      RECT  140.66 86.24 141.15 86.73 ;
      RECT  138.73 86.24 139.22 86.73 ;
      RECT  128.18 86.24 128.67 86.73 ;
      RECT  96.26 81.545 146.18 81.845 ;
      RECT  124.69 72.63 125.18 73.12 ;
      RECT  141.54 76.82 142.03 77.31 ;
      RECT  130.99 76.82 131.48 77.31 ;
      RECT  124.75 76.82 125.24 77.31 ;
      RECT  135.36 72.63 135.85 73.12 ;
      RECT  106.03 76.82 106.52 77.31 ;
      RECT  137.23 76.82 137.72 77.31 ;
      RECT  99.73 72.63 100.22 73.12 ;
      RECT  122.88 72.63 123.37 73.12 ;
      RECT  137.17 72.63 137.66 73.12 ;
      RECT  143.47 76.82 143.96 77.31 ;
      RECT  118.51 76.82 119.0 77.31 ;
      RECT  116.64 72.63 117.13 73.12 ;
      RECT  118.45 72.63 118.94 73.12 ;
      RECT  130.93 72.63 131.42 73.12 ;
      RECT  129.06 76.82 129.55 77.31 ;
      RECT  97.86 76.82 98.35 77.31 ;
      RECT  110.34 76.82 110.83 77.31 ;
      RECT  135.3 76.82 135.79 77.31 ;
      RECT  122.82 76.82 123.31 77.31 ;
      RECT  141.6 72.63 142.09 73.12 ;
      RECT  97.92 72.63 98.41 73.12 ;
      RECT  112.21 72.63 112.7 73.12 ;
      RECT  104.1 76.82 104.59 77.31 ;
      RECT  105.97 72.63 106.46 73.12 ;
      RECT  112.27 76.82 112.76 77.31 ;
      RECT  99.79 76.82 100.28 77.31 ;
      RECT  143.41 72.63 143.9 73.12 ;
      RECT  104.16 72.63 104.65 73.12 ;
      RECT  129.12 72.63 129.61 73.12 ;
      RECT  116.58 76.82 117.07 77.31 ;
      RECT  110.4 72.63 110.89 73.12 ;
      RECT  105.62 80.69 106.11 81.18 ;
      RECT  111.86 80.69 112.35 81.18 ;
      RECT  99.38 80.69 99.87 81.18 ;
      RECT  124.34 80.69 124.83 81.18 ;
      RECT  104.16 71.02 104.65 71.51 ;
      RECT  137.17 71.02 137.66 71.51 ;
      RECT  104.51 80.69 105.0 81.18 ;
      RECT  129.12 71.02 129.61 71.51 ;
      RECT  118.1 80.69 118.59 81.18 ;
      RECT  135.36 71.02 135.85 71.51 ;
      RECT  135.71 80.69 136.2 81.18 ;
      RECT  116.64 71.02 117.13 71.51 ;
      RECT  129.47 80.69 129.96 81.18 ;
      RECT  124.69 71.02 125.18 71.51 ;
      RECT  122.88 71.02 123.37 71.51 ;
      RECT  130.93 71.02 131.42 71.51 ;
      RECT  141.95 80.69 142.44 81.18 ;
      RECT  143.06 80.69 143.55 81.18 ;
      RECT  97.92 71.02 98.41 71.51 ;
      RECT  110.4 71.02 110.89 71.51 ;
      RECT  112.21 71.02 112.7 71.51 ;
      RECT  123.23 80.69 123.72 81.18 ;
      RECT  116.99 80.69 117.48 81.18 ;
      RECT  130.58 80.69 131.07 81.18 ;
      RECT  143.41 71.02 143.9 71.51 ;
      RECT  110.75 80.69 111.24 81.18 ;
      RECT  98.27 80.69 98.76 81.18 ;
      RECT  136.82 80.69 137.31 81.18 ;
      RECT  105.97 71.02 106.46 71.51 ;
      RECT  99.73 71.02 100.22 71.51 ;
      RECT  141.6 71.02 142.09 71.51 ;
      RECT  118.45 71.02 118.94 71.51 ;
      RECT  109.875 60.12 110.365 60.61 ;
      RECT  141.075 60.12 141.565 60.61 ;
      RECT  131.555 64.87 132.045 65.36 ;
      RECT  109.775 64.87 110.265 65.36 ;
      RECT  134.835 60.12 135.325 60.61 ;
      RECT  131.455 60.12 131.945 60.61 ;
      RECT  144.035 64.87 144.525 65.36 ;
      RECT  137.795 64.87 138.285 65.36 ;
      RECT  116.115 60.12 116.605 60.61 ;
      RECT  128.595 60.12 129.085 60.61 ;
      RECT  128.495 64.87 128.985 65.36 ;
      RECT  100.255 60.12 100.745 60.61 ;
      RECT  103.635 60.12 104.125 60.61 ;
      RECT  122.355 60.12 122.845 60.61 ;
      RECT  106.595 64.87 107.085 65.36 ;
      RECT  97.395 60.12 97.885 60.61 ;
      RECT  125.315 64.87 125.805 65.36 ;
      RECT  125.215 60.12 125.705 60.61 ;
      RECT  103.535 64.87 104.025 65.36 ;
      RECT  106.495 60.12 106.985 60.61 ;
      RECT  112.835 64.87 113.325 65.36 ;
      RECT  116.015 64.87 116.505 65.36 ;
      RECT  143.935 60.12 144.425 60.61 ;
      RECT  137.695 60.12 138.185 60.61 ;
      RECT  118.975 60.12 119.465 60.61 ;
      RECT  112.735 60.12 113.225 60.61 ;
      RECT  140.975 64.87 141.465 65.36 ;
      RECT  122.255 64.87 122.745 65.36 ;
      RECT  100.355 64.87 100.845 65.36 ;
      RECT  134.735 64.87 135.225 65.36 ;
      RECT  97.295 64.87 97.785 65.36 ;
      RECT  119.075 64.87 119.565 65.36 ;
      RECT  130.95 63.21 131.44 63.7 ;
      RECT  116.07 67.055 116.56 67.545 ;
      RECT  112.805 62.2 113.295 62.69 ;
      RECT  137.19 63.21 137.68 63.7 ;
      RECT  143.43 63.21 143.92 63.7 ;
      RECT  106.54 67.055 107.03 67.545 ;
      RECT  116.045 62.2 116.535 62.69 ;
      RECT  122.86 63.21 123.35 63.7 ;
      RECT  129.1 63.21 129.59 63.7 ;
      RECT  131.525 62.2 132.015 62.69 ;
      RECT  134.79 67.055 135.28 67.545 ;
      RECT  143.98 67.055 144.47 67.545 ;
      RECT  141.58 63.21 142.07 63.7 ;
      RECT  131.5 67.055 131.99 67.545 ;
      RECT  97.35 67.055 97.84 67.545 ;
      RECT  128.55 67.055 129.04 67.545 ;
      RECT  141.005 62.2 141.495 62.69 ;
      RECT  119.045 62.2 119.535 62.69 ;
      RECT  116.62 63.21 117.11 63.7 ;
      RECT  128.525 62.2 129.015 62.69 ;
      RECT  144.005 62.2 144.495 62.69 ;
      RECT  125.26 67.055 125.75 67.545 ;
      RECT  135.34 63.21 135.83 63.7 ;
      RECT  109.83 67.055 110.32 67.545 ;
      RECT  105.99 63.21 106.48 63.7 ;
      RECT  134.765 62.2 135.255 62.69 ;
      RECT  99.75 63.21 100.24 63.7 ;
      RECT  104.14 63.21 104.63 63.7 ;
      RECT  141.03 67.055 141.52 67.545 ;
      RECT  110.38 63.21 110.87 63.7 ;
      RECT  97.325 62.2 97.815 62.69 ;
      RECT  103.59 67.055 104.08 67.545 ;
      RECT  119.02 67.055 119.51 67.545 ;
      RECT  106.565 62.2 107.055 62.69 ;
      RECT  103.565 62.2 104.055 62.69 ;
      RECT  100.3 67.055 100.79 67.545 ;
      RECT  122.285 62.2 122.775 62.69 ;
      RECT  125.285 62.2 125.775 62.69 ;
      RECT  112.23 63.21 112.72 63.7 ;
      RECT  122.31 67.055 122.8 67.545 ;
      RECT  124.71 63.21 125.2 63.7 ;
      RECT  97.9 63.21 98.39 63.7 ;
      RECT  100.325 62.2 100.815 62.69 ;
      RECT  109.805 62.2 110.295 62.69 ;
      RECT  112.78 67.055 113.27 67.545 ;
      RECT  137.74 67.055 138.23 67.545 ;
      RECT  137.765 62.2 138.255 62.69 ;
      RECT  118.47 63.21 118.96 63.7 ;
      RECT  96.26 54.99 146.18 55.29 ;
      RECT  123.11 57.905 123.6 58.395 ;
      RECT  98.15 57.905 98.64 58.395 ;
      RECT  98.15 52.305 98.64 52.795 ;
      RECT  123.11 52.305 123.6 52.795 ;
      RECT  96.26 81.845 146.18 81.545 ;
      RECT  93.14 83.54 146.18 83.24 ;
      RECT  96.26 55.29 146.18 54.99 ;
      RECT  109.775 65.36 110.265 64.87 ;
      RECT  116.115 60.61 116.605 60.12 ;
      RECT  121.94 86.73 122.43 86.24 ;
      RECT  141.6 73.12 142.09 72.63 ;
      RECT  99.73 73.12 100.22 72.63 ;
      RECT  104.1 77.31 104.59 76.82 ;
      RECT  132.49 86.73 132.98 86.24 ;
      RECT  128.595 60.61 129.085 60.12 ;
      RECT  97.295 65.36 97.785 64.87 ;
      RECT  118.975 60.61 119.465 60.12 ;
      RECT  128.18 86.73 128.67 86.24 ;
      RECT  113.77 86.73 114.26 86.24 ;
      RECT  126.25 86.73 126.74 86.24 ;
      RECT  143.47 77.31 143.96 76.82 ;
      RECT  106.595 65.36 107.085 64.87 ;
      RECT  116.015 65.36 116.505 64.87 ;
      RECT  125.315 65.36 125.805 64.87 ;
      RECT  124.69 73.12 125.18 72.63 ;
      RECT  104.16 73.12 104.65 72.63 ;
      RECT  134.42 86.73 134.91 86.24 ;
      RECT  103.22 86.73 103.71 86.24 ;
      RECT  95.05 86.73 95.54 86.24 ;
      RECT  118.51 77.31 119.0 76.82 ;
      RECT  125.215 60.61 125.705 60.12 ;
      RECT  124.75 77.31 125.24 76.82 ;
      RECT  131.555 65.36 132.045 64.87 ;
      RECT  100.255 60.61 100.745 60.12 ;
      RECT  109.875 60.61 110.365 60.12 ;
      RECT  115.7 86.73 116.19 86.24 ;
      RECT  123.11 58.395 123.6 57.905 ;
      RECT  129.06 77.31 129.55 76.82 ;
      RECT  141.075 60.61 141.565 60.12 ;
      RECT  120.01 86.73 120.5 86.24 ;
      RECT  143.41 73.12 143.9 72.63 ;
      RECT  140.975 65.36 141.465 64.87 ;
      RECT  119.075 65.36 119.565 64.87 ;
      RECT  137.17 73.12 137.66 72.63 ;
      RECT  106.03 77.31 106.52 76.82 ;
      RECT  110.4 73.12 110.89 72.63 ;
      RECT  107.53 86.73 108.02 86.24 ;
      RECT  103.635 60.61 104.125 60.12 ;
      RECT  141.54 77.31 142.03 76.82 ;
      RECT  110.34 77.31 110.83 76.82 ;
      RECT  97.86 77.31 98.35 76.82 ;
      RECT  105.97 73.12 106.46 72.63 ;
      RECT  129.12 73.12 129.61 72.63 ;
      RECT  116.64 73.12 117.13 72.63 ;
      RECT  116.58 77.31 117.07 76.82 ;
      RECT  138.73 86.73 139.22 86.24 ;
      RECT  97.92 73.12 98.41 72.63 ;
      RECT  134.835 60.61 135.325 60.12 ;
      RECT  112.835 65.36 113.325 64.87 ;
      RECT  103.535 65.36 104.025 64.87 ;
      RECT  109.46 86.73 109.95 86.24 ;
      RECT  112.21 73.12 112.7 72.63 ;
      RECT  137.795 65.36 138.285 64.87 ;
      RECT  137.23 77.31 137.72 76.82 ;
      RECT  143.935 60.61 144.425 60.12 ;
      RECT  118.45 73.12 118.94 72.63 ;
      RECT  97.395 60.61 97.885 60.12 ;
      RECT  137.695 60.61 138.185 60.12 ;
      RECT  101.29 86.73 101.78 86.24 ;
      RECT  106.495 60.61 106.985 60.12 ;
      RECT  144.97 86.73 145.46 86.24 ;
      RECT  112.27 77.31 112.76 76.82 ;
      RECT  112.735 60.61 113.225 60.12 ;
      RECT  122.255 65.36 122.745 64.87 ;
      RECT  135.3 77.31 135.79 76.82 ;
      RECT  130.99 77.31 131.48 76.82 ;
      RECT  128.495 65.36 128.985 64.87 ;
      RECT  122.355 60.61 122.845 60.12 ;
      RECT  140.66 86.73 141.15 86.24 ;
      RECT  98.15 58.395 98.64 57.905 ;
      RECT  122.88 73.12 123.37 72.63 ;
      RECT  122.82 77.31 123.31 76.82 ;
      RECT  96.98 86.73 97.47 86.24 ;
      RECT  135.36 73.12 135.85 72.63 ;
      RECT  131.455 60.61 131.945 60.12 ;
      RECT  134.735 65.36 135.225 64.87 ;
      RECT  130.93 73.12 131.42 72.63 ;
      RECT  144.035 65.36 144.525 64.87 ;
      RECT  99.79 77.31 100.28 76.82 ;
      RECT  100.355 65.36 100.845 64.87 ;
      RECT  116.64 71.51 117.13 71.02 ;
      RECT  143.06 81.18 143.55 80.69 ;
      RECT  99.73 71.51 100.22 71.02 ;
      RECT  134.79 67.545 135.28 67.055 ;
      RECT  141.95 81.18 142.44 80.69 ;
      RECT  100.325 62.69 100.815 62.2 ;
      RECT  135.36 71.51 135.85 71.02 ;
      RECT  111.86 81.18 112.35 80.69 ;
      RECT  116.045 62.69 116.535 62.2 ;
      RECT  134.765 62.69 135.255 62.2 ;
      RECT  98.15 52.795 98.64 52.305 ;
      RECT  137.74 67.545 138.23 67.055 ;
      RECT  122.88 71.51 123.37 71.02 ;
      RECT  122.86 63.7 123.35 63.21 ;
      RECT  103.565 62.69 104.055 62.2 ;
      RECT  118.1 81.18 118.59 80.69 ;
      RECT  143.41 71.51 143.9 71.02 ;
      RECT  97.35 67.545 97.84 67.055 ;
      RECT  135.34 63.7 135.83 63.21 ;
      RECT  122.285 62.69 122.775 62.2 ;
      RECT  104.16 71.51 104.65 71.02 ;
      RECT  112.21 71.51 112.7 71.02 ;
      RECT  118.47 63.7 118.96 63.21 ;
      RECT  112.805 62.69 113.295 62.2 ;
      RECT  144.005 62.69 144.495 62.2 ;
      RECT  130.58 81.18 131.07 80.69 ;
      RECT  97.9 63.7 98.39 63.21 ;
      RECT  124.71 63.7 125.2 63.21 ;
      RECT  104.14 63.7 104.63 63.21 ;
      RECT  129.47 81.18 129.96 80.69 ;
      RECT  110.4 71.51 110.89 71.02 ;
      RECT  129.1 63.7 129.59 63.21 ;
      RECT  129.12 71.51 129.61 71.02 ;
      RECT  124.34 81.18 124.83 80.69 ;
      RECT  105.99 63.7 106.48 63.21 ;
      RECT  141.58 63.7 142.07 63.21 ;
      RECT  137.17 71.51 137.66 71.02 ;
      RECT  119.045 62.69 119.535 62.2 ;
      RECT  131.5 67.545 131.99 67.055 ;
      RECT  143.98 67.545 144.47 67.055 ;
      RECT  141.03 67.545 141.52 67.055 ;
      RECT  106.565 62.69 107.055 62.2 ;
      RECT  119.02 67.545 119.51 67.055 ;
      RECT  116.07 67.545 116.56 67.055 ;
      RECT  137.19 63.7 137.68 63.21 ;
      RECT  135.71 81.18 136.2 80.69 ;
      RECT  136.82 81.18 137.31 80.69 ;
      RECT  105.97 71.51 106.46 71.02 ;
      RECT  110.38 63.7 110.87 63.21 ;
      RECT  98.27 81.18 98.76 80.69 ;
      RECT  105.62 81.18 106.11 80.69 ;
      RECT  122.31 67.545 122.8 67.055 ;
      RECT  99.75 63.7 100.24 63.21 ;
      RECT  141.6 71.51 142.09 71.02 ;
      RECT  130.93 71.51 131.42 71.02 ;
      RECT  109.83 67.545 110.32 67.055 ;
      RECT  123.11 52.795 123.6 52.305 ;
      RECT  118.45 71.51 118.94 71.02 ;
      RECT  131.525 62.69 132.015 62.2 ;
      RECT  130.95 63.7 131.44 63.21 ;
      RECT  123.23 81.18 123.72 80.69 ;
      RECT  128.55 67.545 129.04 67.055 ;
      RECT  112.78 67.545 113.27 67.055 ;
      RECT  100.3 67.545 100.79 67.055 ;
      RECT  141.005 62.69 141.495 62.2 ;
      RECT  128.525 62.69 129.015 62.2 ;
      RECT  97.325 62.69 97.815 62.2 ;
      RECT  143.43 63.7 143.92 63.21 ;
      RECT  112.23 63.7 112.72 63.21 ;
      RECT  110.75 81.18 111.24 80.69 ;
      RECT  104.51 81.18 105.0 80.69 ;
      RECT  109.805 62.69 110.295 62.2 ;
      RECT  125.26 67.545 125.75 67.055 ;
      RECT  97.92 71.51 98.41 71.02 ;
      RECT  116.62 63.7 117.11 63.21 ;
      RECT  124.69 71.51 125.18 71.02 ;
      RECT  99.38 81.18 99.87 80.69 ;
      RECT  125.285 62.69 125.775 62.2 ;
      RECT  116.99 81.18 117.48 80.69 ;
      RECT  106.54 67.545 107.03 67.055 ;
      RECT  103.59 67.545 104.08 67.055 ;
      RECT  137.765 62.69 138.255 62.2 ;
      RECT  96.98 129.85 97.47 129.36 ;
      RECT  101.78 129.85 101.29 129.36 ;
      RECT  103.22 129.85 103.71 129.36 ;
      RECT  108.02 129.85 107.53 129.36 ;
      RECT  109.46 129.85 109.95 129.36 ;
      RECT  114.26 129.85 113.77 129.36 ;
      RECT  115.7 129.85 116.19 129.36 ;
      RECT  120.5 129.85 120.01 129.36 ;
      RECT  121.94 129.85 122.43 129.36 ;
      RECT  126.74 129.85 126.25 129.36 ;
      RECT  128.18 129.85 128.67 129.36 ;
      RECT  132.98 129.85 132.49 129.36 ;
      RECT  134.42 129.85 134.91 129.36 ;
      RECT  139.22 129.85 138.73 129.36 ;
      RECT  140.66 129.85 141.15 129.36 ;
      RECT  145.46 129.85 144.97 129.36 ;
      RECT  146.9 129.85 147.39 129.36 ;
      RECT  96.26 132.85 149.3 132.55 ;
      RECT  115.7 129.85 116.19 129.36 ;
      RECT  109.46 129.85 109.95 129.36 ;
      RECT  138.73 129.85 139.22 129.36 ;
      RECT  126.25 129.85 126.74 129.36 ;
      RECT  101.29 129.85 101.78 129.36 ;
      RECT  120.01 129.85 120.5 129.36 ;
      RECT  128.18 129.85 128.67 129.36 ;
      RECT  146.9 129.85 147.39 129.36 ;
      RECT  96.98 129.85 97.47 129.36 ;
      RECT  113.77 129.85 114.26 129.36 ;
      RECT  140.66 129.85 141.15 129.36 ;
      RECT  121.94 129.85 122.43 129.36 ;
      RECT  103.22 129.85 103.71 129.36 ;
      RECT  132.49 129.85 132.98 129.36 ;
      RECT  107.53 129.85 108.02 129.36 ;
      RECT  134.42 129.85 134.91 129.36 ;
      RECT  144.97 129.85 145.46 129.36 ;
      RECT  96.26 134.545 146.18 134.245 ;
      RECT  124.69 143.46 125.18 142.97 ;
      RECT  141.54 139.27 142.03 138.78 ;
      RECT  130.99 139.27 131.48 138.78 ;
      RECT  124.75 139.27 125.24 138.78 ;
      RECT  135.36 143.46 135.85 142.97 ;
      RECT  106.03 139.27 106.52 138.78 ;
      RECT  137.23 139.27 137.72 138.78 ;
      RECT  99.73 143.46 100.22 142.97 ;
      RECT  122.88 143.46 123.37 142.97 ;
      RECT  137.17 143.46 137.66 142.97 ;
      RECT  143.47 139.27 143.96 138.78 ;
      RECT  118.51 139.27 119.0 138.78 ;
      RECT  116.64 143.46 117.13 142.97 ;
      RECT  118.45 143.46 118.94 142.97 ;
      RECT  130.93 143.46 131.42 142.97 ;
      RECT  129.06 139.27 129.55 138.78 ;
      RECT  97.86 139.27 98.35 138.78 ;
      RECT  110.34 139.27 110.83 138.78 ;
      RECT  135.3 139.27 135.79 138.78 ;
      RECT  122.82 139.27 123.31 138.78 ;
      RECT  141.6 143.46 142.09 142.97 ;
      RECT  97.92 143.46 98.41 142.97 ;
      RECT  112.21 143.46 112.7 142.97 ;
      RECT  104.1 139.27 104.59 138.78 ;
      RECT  105.97 143.46 106.46 142.97 ;
      RECT  112.27 139.27 112.76 138.78 ;
      RECT  99.79 139.27 100.28 138.78 ;
      RECT  143.41 143.46 143.9 142.97 ;
      RECT  104.16 143.46 104.65 142.97 ;
      RECT  129.12 143.46 129.61 142.97 ;
      RECT  116.58 139.27 117.07 138.78 ;
      RECT  110.4 143.46 110.89 142.97 ;
      RECT  105.62 135.4 106.11 134.91 ;
      RECT  111.86 135.4 112.35 134.91 ;
      RECT  99.38 135.4 99.87 134.91 ;
      RECT  124.34 135.4 124.83 134.91 ;
      RECT  104.16 145.07 104.65 144.58 ;
      RECT  137.17 145.07 137.66 144.58 ;
      RECT  104.51 135.4 105.0 134.91 ;
      RECT  129.12 145.07 129.61 144.58 ;
      RECT  118.1 135.4 118.59 134.91 ;
      RECT  135.36 145.07 135.85 144.58 ;
      RECT  135.71 135.4 136.2 134.91 ;
      RECT  116.64 145.07 117.13 144.58 ;
      RECT  129.47 135.4 129.96 134.91 ;
      RECT  124.69 145.07 125.18 144.58 ;
      RECT  122.88 145.07 123.37 144.58 ;
      RECT  130.93 145.07 131.42 144.58 ;
      RECT  141.95 135.4 142.44 134.91 ;
      RECT  143.06 135.4 143.55 134.91 ;
      RECT  97.92 145.07 98.41 144.58 ;
      RECT  110.4 145.07 110.89 144.58 ;
      RECT  112.21 145.07 112.7 144.58 ;
      RECT  123.23 135.4 123.72 134.91 ;
      RECT  116.99 135.4 117.48 134.91 ;
      RECT  130.58 135.4 131.07 134.91 ;
      RECT  143.41 145.07 143.9 144.58 ;
      RECT  110.75 135.4 111.24 134.91 ;
      RECT  98.27 135.4 98.76 134.91 ;
      RECT  136.82 135.4 137.31 134.91 ;
      RECT  105.97 145.07 106.46 144.58 ;
      RECT  99.73 145.07 100.22 144.58 ;
      RECT  141.6 145.07 142.09 144.58 ;
      RECT  118.45 145.07 118.94 144.58 ;
      RECT  96.26 134.245 146.18 134.545 ;
      RECT  96.26 132.55 149.3 132.85 ;
      RECT  121.94 129.36 122.43 129.85 ;
      RECT  140.66 129.36 141.15 129.85 ;
      RECT  137.23 138.78 137.72 139.27 ;
      RECT  134.42 129.36 134.91 129.85 ;
      RECT  124.69 142.97 125.18 143.46 ;
      RECT  132.49 129.36 132.98 129.85 ;
      RECT  99.73 142.97 100.22 143.46 ;
      RECT  107.53 129.36 108.02 129.85 ;
      RECT  113.77 129.36 114.26 129.85 ;
      RECT  129.06 138.78 129.55 139.27 ;
      RECT  110.4 142.97 110.89 143.46 ;
      RECT  112.27 138.78 112.76 139.27 ;
      RECT  122.82 138.78 123.31 139.27 ;
      RECT  103.22 129.36 103.71 129.85 ;
      RECT  115.7 129.36 116.19 129.85 ;
      RECT  118.51 138.78 119.0 139.27 ;
      RECT  138.73 129.36 139.22 129.85 ;
      RECT  143.41 142.97 143.9 143.46 ;
      RECT  135.3 138.78 135.79 139.27 ;
      RECT  110.34 138.78 110.83 139.27 ;
      RECT  137.17 142.97 137.66 143.46 ;
      RECT  130.93 142.97 131.42 143.46 ;
      RECT  118.45 142.97 118.94 143.46 ;
      RECT  101.29 129.36 101.78 129.85 ;
      RECT  116.58 138.78 117.07 139.27 ;
      RECT  144.97 129.36 145.46 129.85 ;
      RECT  106.03 138.78 106.52 139.27 ;
      RECT  129.12 142.97 129.61 143.46 ;
      RECT  96.98 129.36 97.47 129.85 ;
      RECT  146.9 129.36 147.39 129.85 ;
      RECT  124.75 138.78 125.24 139.27 ;
      RECT  141.6 142.97 142.09 143.46 ;
      RECT  135.36 142.97 135.85 143.46 ;
      RECT  128.18 129.36 128.67 129.85 ;
      RECT  116.64 142.97 117.13 143.46 ;
      RECT  109.46 129.36 109.95 129.85 ;
      RECT  112.21 142.97 112.7 143.46 ;
      RECT  97.92 142.97 98.41 143.46 ;
      RECT  105.97 142.97 106.46 143.46 ;
      RECT  120.01 129.36 120.5 129.85 ;
      RECT  143.47 138.78 143.96 139.27 ;
      RECT  130.99 138.78 131.48 139.27 ;
      RECT  99.79 138.78 100.28 139.27 ;
      RECT  126.25 129.36 126.74 129.85 ;
      RECT  141.54 138.78 142.03 139.27 ;
      RECT  97.86 138.78 98.35 139.27 ;
      RECT  104.1 138.78 104.59 139.27 ;
      RECT  104.16 142.97 104.65 143.46 ;
      RECT  122.88 142.97 123.37 143.46 ;
      RECT  112.21 144.58 112.7 145.07 ;
      RECT  143.41 144.58 143.9 145.07 ;
      RECT  122.88 144.58 123.37 145.07 ;
      RECT  143.06 134.91 143.55 135.4 ;
      RECT  110.75 134.91 111.24 135.4 ;
      RECT  141.95 134.91 142.44 135.4 ;
      RECT  104.16 144.58 104.65 145.07 ;
      RECT  104.51 134.91 105.0 135.4 ;
      RECT  118.45 144.58 118.94 145.07 ;
      RECT  105.62 134.91 106.11 135.4 ;
      RECT  99.73 144.58 100.22 145.07 ;
      RECT  130.93 144.58 131.42 145.07 ;
      RECT  116.64 144.58 117.13 145.07 ;
      RECT  105.97 144.58 106.46 145.07 ;
      RECT  124.34 134.91 124.83 135.4 ;
      RECT  129.47 134.91 129.96 135.4 ;
      RECT  111.86 134.91 112.35 135.4 ;
      RECT  123.23 134.91 123.72 135.4 ;
      RECT  136.82 134.91 137.31 135.4 ;
      RECT  135.71 134.91 136.2 135.4 ;
      RECT  137.17 144.58 137.66 145.07 ;
      RECT  130.58 134.91 131.07 135.4 ;
      RECT  116.99 134.91 117.48 135.4 ;
      RECT  99.38 134.91 99.87 135.4 ;
      RECT  97.92 144.58 98.41 145.07 ;
      RECT  129.12 144.58 129.61 145.07 ;
      RECT  98.27 134.91 98.76 135.4 ;
      RECT  135.36 144.58 135.85 145.07 ;
      RECT  110.4 144.58 110.89 145.07 ;
      RECT  124.69 144.58 125.18 145.07 ;
      RECT  141.6 144.58 142.09 145.07 ;
      RECT  118.1 134.91 118.59 135.4 ;
      RECT  53.14 94.155 53.63 94.645 ;
      RECT  53.14 98.105 53.63 98.595 ;
      RECT  46.525 94.12 47.015 94.61 ;
      RECT  56.395 94.12 56.885 94.61 ;
      RECT  56.395 98.07 56.885 98.56 ;
      RECT  51.015 98.105 51.505 98.595 ;
      RECT  45.165 94.12 45.655 94.61 ;
      RECT  55.035 98.07 55.525 98.56 ;
      RECT  51.015 94.155 51.505 94.645 ;
      RECT  55.035 94.12 55.525 94.61 ;
      RECT  53.14 106.005 53.63 106.495 ;
      RECT  53.14 109.955 53.63 110.445 ;
      RECT  46.525 105.97 47.015 106.46 ;
      RECT  56.395 105.97 56.885 106.46 ;
      RECT  56.395 109.92 56.885 110.41 ;
      RECT  51.015 109.955 51.505 110.445 ;
      RECT  45.165 105.97 45.655 106.46 ;
      RECT  55.035 109.92 55.525 110.41 ;
      RECT  51.015 106.005 51.505 106.495 ;
      RECT  55.035 105.97 55.525 106.46 ;
      RECT  67.465 94.12 67.955 94.61 ;
      RECT  67.465 98.07 67.955 98.56 ;
      RECT  64.21 121.805 64.7 122.295 ;
      RECT  64.21 96.255 64.7 96.745 ;
      RECT  64.21 98.105 64.7 98.595 ;
      RECT  53.14 106.005 53.63 106.495 ;
      RECT  67.465 103.995 67.955 104.485 ;
      RECT  67.465 119.795 67.955 120.285 ;
      RECT  64.21 117.855 64.7 118.345 ;
      RECT  67.465 102.02 67.955 102.51 ;
      RECT  64.21 102.055 64.7 102.545 ;
      RECT  64.21 113.905 64.7 114.395 ;
      RECT  67.465 117.82 67.955 118.31 ;
      RECT  56.395 94.12 56.885 94.61 ;
      RECT  56.395 98.07 56.885 98.56 ;
      RECT  53.14 94.155 53.63 94.645 ;
      RECT  64.21 109.955 64.7 110.445 ;
      RECT  67.465 113.87 67.955 114.36 ;
      RECT  67.465 121.77 67.955 122.26 ;
      RECT  53.14 109.955 53.63 110.445 ;
      RECT  56.395 105.97 56.885 106.46 ;
      RECT  64.21 94.155 64.7 94.645 ;
      RECT  67.465 96.095 67.955 96.585 ;
      RECT  56.395 109.92 56.885 110.41 ;
      RECT  64.21 108.105 64.7 108.595 ;
      RECT  67.465 107.945 67.955 108.435 ;
      RECT  46.525 105.97 47.015 106.46 ;
      RECT  64.21 119.955 64.7 120.445 ;
      RECT  53.14 98.105 53.63 98.595 ;
      RECT  64.21 100.205 64.7 100.695 ;
      RECT  46.525 94.12 47.015 94.61 ;
      RECT  67.465 111.895 67.955 112.385 ;
      RECT  67.465 100.045 67.955 100.535 ;
      RECT  64.21 112.055 64.7 112.545 ;
      RECT  67.465 109.92 67.955 110.41 ;
      RECT  67.465 115.845 67.955 116.335 ;
      RECT  67.465 105.97 67.955 106.46 ;
      RECT  64.21 106.005 64.7 106.495 ;
      RECT  64.21 116.005 64.7 116.495 ;
      RECT  64.21 104.155 64.7 104.645 ;
      RECT  66.105 111.895 66.595 112.385 ;
      RECT  66.105 119.795 66.595 120.285 ;
      RECT  55.035 109.92 55.525 110.41 ;
      RECT  66.105 115.845 66.595 116.335 ;
      RECT  62.085 94.155 62.575 94.645 ;
      RECT  62.085 100.195 62.575 100.685 ;
      RECT  62.085 102.055 62.575 102.545 ;
      RECT  66.105 107.945 66.595 108.435 ;
      RECT  45.165 105.97 45.655 106.46 ;
      RECT  62.085 108.095 62.575 108.585 ;
      RECT  55.035 105.97 55.525 106.46 ;
      RECT  62.085 112.045 62.575 112.535 ;
      RECT  66.105 96.095 66.595 96.585 ;
      RECT  66.105 121.77 66.595 122.26 ;
      RECT  55.035 98.07 55.525 98.56 ;
      RECT  62.085 113.905 62.575 114.395 ;
      RECT  66.105 109.92 66.595 110.41 ;
      RECT  51.015 94.155 51.505 94.645 ;
      RECT  55.035 94.12 55.525 94.61 ;
      RECT  51.015 106.005 51.505 106.495 ;
      RECT  66.105 103.995 66.595 104.485 ;
      RECT  62.085 98.105 62.575 98.595 ;
      RECT  66.105 117.82 66.595 118.31 ;
      RECT  62.085 104.145 62.575 104.635 ;
      RECT  62.085 109.955 62.575 110.445 ;
      RECT  62.085 106.005 62.575 106.495 ;
      RECT  66.105 100.045 66.595 100.535 ;
      RECT  62.085 117.855 62.575 118.345 ;
      RECT  62.085 121.805 62.575 122.295 ;
      RECT  66.105 98.07 66.595 98.56 ;
      RECT  45.165 94.12 45.655 94.61 ;
      RECT  62.085 119.945 62.575 120.435 ;
      RECT  62.085 96.245 62.575 96.735 ;
      RECT  62.085 115.995 62.575 116.485 ;
      RECT  66.105 94.12 66.595 94.61 ;
      RECT  66.105 102.02 66.595 102.51 ;
      RECT  51.015 98.105 51.505 98.595 ;
      RECT  66.105 105.97 66.595 106.46 ;
      RECT  51.015 109.955 51.505 110.445 ;
      RECT  66.105 113.87 66.595 114.36 ;
      RECT  64.21 108.105 64.7 108.595 ;
      RECT  64.21 119.955 64.7 120.445 ;
      RECT  67.465 96.095 67.955 96.585 ;
      RECT  64.21 102.055 64.7 102.545 ;
      RECT  64.21 94.155 64.7 94.645 ;
      RECT  67.465 100.045 67.955 100.535 ;
      RECT  64.21 113.905 64.7 114.395 ;
      RECT  67.465 117.82 67.955 118.31 ;
      RECT  67.465 105.97 67.955 106.46 ;
      RECT  53.14 109.955 53.63 110.445 ;
      RECT  64.21 106.005 64.7 106.495 ;
      RECT  56.395 94.12 56.885 94.61 ;
      RECT  64.21 109.955 64.7 110.445 ;
      RECT  67.465 103.995 67.955 104.485 ;
      RECT  64.21 121.805 64.7 122.295 ;
      RECT  67.465 102.02 67.955 102.51 ;
      RECT  67.465 115.845 67.955 116.335 ;
      RECT  53.14 98.105 53.63 98.595 ;
      RECT  71.82 107.72 72.31 108.21 ;
      RECT  67.465 121.77 67.955 122.26 ;
      RECT  67.465 94.12 67.955 94.61 ;
      RECT  64.21 112.055 64.7 112.545 ;
      RECT  64.21 117.855 64.7 118.345 ;
      RECT  67.465 111.895 67.955 112.385 ;
      RECT  67.465 107.945 67.955 108.435 ;
      RECT  67.465 113.87 67.955 114.36 ;
      RECT  64.21 116.005 64.7 116.495 ;
      RECT  56.395 109.92 56.885 110.41 ;
      RECT  64.21 100.205 64.7 100.695 ;
      RECT  67.465 109.92 67.955 110.41 ;
      RECT  64.21 104.155 64.7 104.645 ;
      RECT  53.14 106.005 53.63 106.495 ;
      RECT  67.465 98.07 67.955 98.56 ;
      RECT  56.395 98.07 56.885 98.56 ;
      RECT  53.14 94.155 53.63 94.645 ;
      RECT  46.525 94.12 47.015 94.61 ;
      RECT  67.465 119.795 67.955 120.285 ;
      RECT  84.655 107.8 85.145 108.29 ;
      RECT  64.21 96.255 64.7 96.745 ;
      RECT  56.395 105.97 56.885 106.46 ;
      RECT  46.525 105.97 47.015 106.46 ;
      RECT  64.21 98.105 64.7 98.595 ;
      RECT  55.035 94.12 55.525 94.61 ;
      RECT  66.105 117.82 66.595 118.31 ;
      RECT  66.105 103.995 66.595 104.485 ;
      RECT  62.085 100.195 62.575 100.685 ;
      RECT  62.085 121.805 62.575 122.295 ;
      RECT  66.105 119.795 66.595 120.285 ;
      RECT  66.105 107.945 66.595 108.435 ;
      RECT  66.105 105.97 66.595 106.46 ;
      RECT  66.105 100.045 66.595 100.535 ;
      RECT  51.015 98.105 51.505 98.595 ;
      RECT  62.085 96.245 62.575 96.735 ;
      RECT  66.105 113.87 66.595 114.36 ;
      RECT  66.105 98.07 66.595 98.56 ;
      RECT  45.165 105.97 45.655 106.46 ;
      RECT  62.085 119.945 62.575 120.435 ;
      RECT  62.085 106.005 62.575 106.495 ;
      RECT  51.015 94.155 51.505 94.645 ;
      RECT  51.015 106.005 51.505 106.495 ;
      RECT  66.105 111.895 66.595 112.385 ;
      RECT  51.015 109.955 51.505 110.445 ;
      RECT  62.085 113.905 62.575 114.395 ;
      RECT  77.035 107.8 77.525 108.29 ;
      RECT  62.085 94.155 62.575 94.645 ;
      RECT  62.085 104.145 62.575 104.635 ;
      RECT  69.695 107.725 70.185 108.215 ;
      RECT  55.035 98.07 55.525 98.56 ;
      RECT  66.105 115.845 66.595 116.335 ;
      RECT  66.105 121.77 66.595 122.26 ;
      RECT  62.085 109.955 62.575 110.445 ;
      RECT  62.085 98.105 62.575 98.595 ;
      RECT  62.085 115.995 62.575 116.485 ;
      RECT  62.085 117.855 62.575 118.345 ;
      RECT  62.085 112.045 62.575 112.535 ;
      RECT  62.085 108.095 62.575 108.585 ;
      RECT  66.105 94.12 66.595 94.61 ;
      RECT  55.035 109.92 55.525 110.41 ;
      RECT  45.165 94.12 45.655 94.61 ;
      RECT  66.105 102.02 66.595 102.51 ;
      RECT  66.105 96.095 66.595 96.585 ;
      RECT  62.085 102.055 62.575 102.545 ;
      RECT  66.105 109.92 66.595 110.41 ;
      RECT  55.035 105.97 55.525 106.46 ;
      RECT  189.3 94.155 188.81 94.645 ;
      RECT  189.3 98.105 188.81 98.595 ;
      RECT  195.915 94.12 195.425 94.61 ;
      RECT  186.045 94.12 185.555 94.61 ;
      RECT  186.045 98.07 185.555 98.56 ;
      RECT  191.425 98.105 190.935 98.595 ;
      RECT  197.275 94.12 196.785 94.61 ;
      RECT  187.405 98.07 186.915 98.56 ;
      RECT  191.425 94.155 190.935 94.645 ;
      RECT  187.405 94.12 186.915 94.61 ;
      RECT  189.3 106.005 188.81 106.495 ;
      RECT  189.3 109.955 188.81 110.445 ;
      RECT  195.915 105.97 195.425 106.46 ;
      RECT  186.045 105.97 185.555 106.46 ;
      RECT  186.045 109.92 185.555 110.41 ;
      RECT  191.425 109.955 190.935 110.445 ;
      RECT  197.275 105.97 196.785 106.46 ;
      RECT  187.405 109.92 186.915 110.41 ;
      RECT  191.425 106.005 190.935 106.495 ;
      RECT  187.405 105.97 186.915 106.46 ;
      RECT  174.975 94.12 174.485 94.61 ;
      RECT  174.975 98.07 174.485 98.56 ;
      RECT  178.23 121.805 177.74 122.295 ;
      RECT  178.23 96.255 177.74 96.745 ;
      RECT  178.23 98.105 177.74 98.595 ;
      RECT  189.3 106.005 188.81 106.495 ;
      RECT  174.975 103.995 174.485 104.485 ;
      RECT  174.975 119.795 174.485 120.285 ;
      RECT  178.23 117.855 177.74 118.345 ;
      RECT  174.975 102.02 174.485 102.51 ;
      RECT  178.23 102.055 177.74 102.545 ;
      RECT  178.23 113.905 177.74 114.395 ;
      RECT  174.975 117.82 174.485 118.31 ;
      RECT  186.045 94.12 185.555 94.61 ;
      RECT  186.045 98.07 185.555 98.56 ;
      RECT  189.3 94.155 188.81 94.645 ;
      RECT  178.23 109.955 177.74 110.445 ;
      RECT  174.975 113.87 174.485 114.36 ;
      RECT  174.975 121.77 174.485 122.26 ;
      RECT  189.3 109.955 188.81 110.445 ;
      RECT  186.045 105.97 185.555 106.46 ;
      RECT  178.23 94.155 177.74 94.645 ;
      RECT  174.975 96.095 174.485 96.585 ;
      RECT  186.045 109.92 185.555 110.41 ;
      RECT  178.23 108.105 177.74 108.595 ;
      RECT  174.975 107.945 174.485 108.435 ;
      RECT  195.915 105.97 195.425 106.46 ;
      RECT  178.23 119.955 177.74 120.445 ;
      RECT  189.3 98.105 188.81 98.595 ;
      RECT  178.23 100.205 177.74 100.695 ;
      RECT  195.915 94.12 195.425 94.61 ;
      RECT  174.975 111.895 174.485 112.385 ;
      RECT  174.975 100.045 174.485 100.535 ;
      RECT  178.23 112.055 177.74 112.545 ;
      RECT  174.975 109.92 174.485 110.41 ;
      RECT  174.975 115.845 174.485 116.335 ;
      RECT  174.975 105.97 174.485 106.46 ;
      RECT  178.23 106.005 177.74 106.495 ;
      RECT  178.23 116.005 177.74 116.495 ;
      RECT  178.23 104.155 177.74 104.645 ;
      RECT  176.335 111.895 175.845 112.385 ;
      RECT  176.335 119.795 175.845 120.285 ;
      RECT  187.405 109.92 186.915 110.41 ;
      RECT  176.335 115.845 175.845 116.335 ;
      RECT  180.355 94.155 179.865 94.645 ;
      RECT  180.355 100.195 179.865 100.685 ;
      RECT  180.355 102.055 179.865 102.545 ;
      RECT  176.335 107.945 175.845 108.435 ;
      RECT  197.275 105.97 196.785 106.46 ;
      RECT  180.355 108.095 179.865 108.585 ;
      RECT  187.405 105.97 186.915 106.46 ;
      RECT  180.355 112.045 179.865 112.535 ;
      RECT  176.335 96.095 175.845 96.585 ;
      RECT  176.335 121.77 175.845 122.26 ;
      RECT  187.405 98.07 186.915 98.56 ;
      RECT  180.355 113.905 179.865 114.395 ;
      RECT  176.335 109.92 175.845 110.41 ;
      RECT  191.425 94.155 190.935 94.645 ;
      RECT  187.405 94.12 186.915 94.61 ;
      RECT  191.425 106.005 190.935 106.495 ;
      RECT  176.335 103.995 175.845 104.485 ;
      RECT  180.355 98.105 179.865 98.595 ;
      RECT  176.335 117.82 175.845 118.31 ;
      RECT  180.355 104.145 179.865 104.635 ;
      RECT  180.355 109.955 179.865 110.445 ;
      RECT  180.355 106.005 179.865 106.495 ;
      RECT  176.335 100.045 175.845 100.535 ;
      RECT  180.355 117.855 179.865 118.345 ;
      RECT  180.355 121.805 179.865 122.295 ;
      RECT  176.335 98.07 175.845 98.56 ;
      RECT  197.275 94.12 196.785 94.61 ;
      RECT  180.355 119.945 179.865 120.435 ;
      RECT  180.355 96.245 179.865 96.735 ;
      RECT  180.355 115.995 179.865 116.485 ;
      RECT  176.335 94.12 175.845 94.61 ;
      RECT  176.335 102.02 175.845 102.51 ;
      RECT  191.425 98.105 190.935 98.595 ;
      RECT  176.335 105.97 175.845 106.46 ;
      RECT  191.425 109.955 190.935 110.445 ;
      RECT  176.335 113.87 175.845 114.36 ;
      RECT  178.23 108.105 177.74 108.595 ;
      RECT  178.23 119.955 177.74 120.445 ;
      RECT  174.975 96.095 174.485 96.585 ;
      RECT  178.23 102.055 177.74 102.545 ;
      RECT  178.23 94.155 177.74 94.645 ;
      RECT  174.975 100.045 174.485 100.535 ;
      RECT  178.23 113.905 177.74 114.395 ;
      RECT  174.975 117.82 174.485 118.31 ;
      RECT  174.975 105.97 174.485 106.46 ;
      RECT  189.3 109.955 188.81 110.445 ;
      RECT  178.23 106.005 177.74 106.495 ;
      RECT  186.045 94.12 185.555 94.61 ;
      RECT  178.23 109.955 177.74 110.445 ;
      RECT  174.975 103.995 174.485 104.485 ;
      RECT  178.23 121.805 177.74 122.295 ;
      RECT  174.975 102.02 174.485 102.51 ;
      RECT  174.975 115.845 174.485 116.335 ;
      RECT  189.3 98.105 188.81 98.595 ;
      RECT  170.62 107.72 170.13 108.21 ;
      RECT  174.975 121.77 174.485 122.26 ;
      RECT  174.975 94.12 174.485 94.61 ;
      RECT  178.23 112.055 177.74 112.545 ;
      RECT  178.23 117.855 177.74 118.345 ;
      RECT  174.975 111.895 174.485 112.385 ;
      RECT  174.975 107.945 174.485 108.435 ;
      RECT  174.975 113.87 174.485 114.36 ;
      RECT  178.23 116.005 177.74 116.495 ;
      RECT  186.045 109.92 185.555 110.41 ;
      RECT  178.23 100.205 177.74 100.695 ;
      RECT  174.975 109.92 174.485 110.41 ;
      RECT  178.23 104.155 177.74 104.645 ;
      RECT  189.3 106.005 188.81 106.495 ;
      RECT  174.975 98.07 174.485 98.56 ;
      RECT  186.045 98.07 185.555 98.56 ;
      RECT  189.3 94.155 188.81 94.645 ;
      RECT  195.915 94.12 195.425 94.61 ;
      RECT  174.975 119.795 174.485 120.285 ;
      RECT  157.785 107.8 157.295 108.29 ;
      RECT  178.23 96.255 177.74 96.745 ;
      RECT  186.045 105.97 185.555 106.46 ;
      RECT  195.915 105.97 195.425 106.46 ;
      RECT  178.23 98.105 177.74 98.595 ;
      RECT  187.405 94.12 186.915 94.61 ;
      RECT  176.335 117.82 175.845 118.31 ;
      RECT  176.335 103.995 175.845 104.485 ;
      RECT  180.355 100.195 179.865 100.685 ;
      RECT  180.355 121.805 179.865 122.295 ;
      RECT  176.335 119.795 175.845 120.285 ;
      RECT  176.335 107.945 175.845 108.435 ;
      RECT  176.335 105.97 175.845 106.46 ;
      RECT  176.335 100.045 175.845 100.535 ;
      RECT  191.425 98.105 190.935 98.595 ;
      RECT  180.355 96.245 179.865 96.735 ;
      RECT  176.335 113.87 175.845 114.36 ;
      RECT  176.335 98.07 175.845 98.56 ;
      RECT  197.275 105.97 196.785 106.46 ;
      RECT  180.355 119.945 179.865 120.435 ;
      RECT  180.355 106.005 179.865 106.495 ;
      RECT  191.425 94.155 190.935 94.645 ;
      RECT  191.425 106.005 190.935 106.495 ;
      RECT  176.335 111.895 175.845 112.385 ;
      RECT  191.425 109.955 190.935 110.445 ;
      RECT  180.355 113.905 179.865 114.395 ;
      RECT  165.405 107.8 164.915 108.29 ;
      RECT  180.355 94.155 179.865 94.645 ;
      RECT  180.355 104.145 179.865 104.635 ;
      RECT  172.745 107.725 172.255 108.215 ;
      RECT  187.405 98.07 186.915 98.56 ;
      RECT  176.335 115.845 175.845 116.335 ;
      RECT  176.335 121.77 175.845 122.26 ;
      RECT  180.355 109.955 179.865 110.445 ;
      RECT  180.355 98.105 179.865 98.595 ;
      RECT  180.355 115.995 179.865 116.485 ;
      RECT  180.355 117.855 179.865 118.345 ;
      RECT  180.355 112.045 179.865 112.535 ;
      RECT  180.355 108.095 179.865 108.585 ;
      RECT  176.335 94.12 175.845 94.61 ;
      RECT  187.405 109.92 186.915 110.41 ;
      RECT  197.275 94.12 196.785 94.61 ;
      RECT  176.335 102.02 175.845 102.51 ;
      RECT  176.335 96.095 175.845 96.585 ;
      RECT  180.355 102.055 179.865 102.545 ;
      RECT  176.335 109.92 175.845 110.41 ;
      RECT  187.405 105.97 186.915 106.46 ;
      RECT  97.395 60.12 97.885 60.61 ;
      RECT  103.535 64.87 104.025 65.36 ;
      RECT  129.06 76.82 129.55 77.31 ;
      RECT  53.14 94.155 53.63 94.645 ;
      RECT  138.73 86.24 139.22 86.73 ;
      RECT  177.74 94.155 178.23 94.645 ;
      RECT  101.29 129.36 101.78 129.85 ;
      RECT  177.74 112.055 178.23 112.545 ;
      RECT  138.23 89.29 138.53 89.59 ;
      RECT  53.14 98.105 53.63 98.595 ;
      RECT  170.13 107.72 170.62 108.21 ;
      RECT  104.1 138.78 104.59 139.27 ;
      RECT  125.215 60.12 125.705 60.61 ;
      RECT  144.47 126.5 144.77 126.8 ;
      RECT  141.35 89.29 141.65 89.59 ;
      RECT  131.99 89.29 132.29 89.59 ;
      RECT  177.74 102.055 178.23 102.545 ;
      RECT  185.555 94.12 186.045 94.61 ;
      RECT  112.735 60.12 113.225 60.61 ;
      RECT  104.16 142.97 104.65 143.46 ;
      RECT  147.495 126.405 147.985 126.895 ;
      RECT  64.21 102.055 64.7 102.545 ;
      RECT  128.87 89.29 129.17 89.59 ;
      RECT  128.595 60.12 129.085 60.61 ;
      RECT  67.465 115.845 67.955 116.335 ;
      RECT  67.465 107.945 67.955 108.435 ;
      RECT  174.485 105.97 174.975 106.46 ;
      RECT  113.77 86.24 114.26 86.73 ;
      RECT  109.46 86.24 109.95 86.73 ;
      RECT  124.75 138.78 125.24 139.27 ;
      RECT  67.465 96.095 67.955 96.585 ;
      RECT  129.12 142.97 129.61 143.46 ;
      RECT  126.25 129.36 126.74 129.85 ;
      RECT  134.735 64.87 135.225 65.36 ;
      RECT  94.455 89.195 94.945 89.685 ;
      RECT  122.82 138.78 123.31 139.27 ;
      RECT  174.485 119.795 174.975 120.285 ;
      RECT  185.555 105.97 186.045 106.46 ;
      RECT  124.69 72.63 125.18 73.12 ;
      RECT  134.42 86.24 134.91 86.73 ;
      RECT  122.63 89.29 122.93 89.59 ;
      RECT  64.21 104.155 64.7 104.645 ;
      RECT  112.21 72.63 112.7 73.12 ;
      RECT  188.81 106.005 189.3 106.495 ;
      RECT  116.39 126.5 116.69 126.8 ;
      RECT  116.58 138.78 117.07 139.27 ;
      RECT  134.835 60.12 135.325 60.61 ;
      RECT  177.74 116.005 178.23 116.495 ;
      RECT  120.01 129.36 120.5 129.85 ;
      RECT  131.455 60.12 131.945 60.61 ;
      RECT  125.315 64.87 125.805 65.36 ;
      RECT  177.74 106.005 178.23 106.495 ;
      RECT  116.64 72.63 117.13 73.12 ;
      RECT  99.79 76.82 100.28 77.31 ;
      RECT  64.21 98.105 64.7 98.595 ;
      RECT  131.555 64.87 132.045 65.36 ;
      RECT  188.81 109.955 189.3 110.445 ;
      RECT  100.79 89.29 101.09 89.59 ;
      RECT  115.7 129.36 116.19 129.85 ;
      RECT  177.74 98.105 178.23 98.595 ;
      RECT  143.935 60.12 144.425 60.61 ;
      RECT  177.74 100.205 178.23 100.695 ;
      RECT  174.485 121.77 174.975 122.26 ;
      RECT  129.06 138.78 129.55 139.27 ;
      RECT  64.21 116.005 64.7 116.495 ;
      RECT  135.36 72.63 135.85 73.12 ;
      RECT  104.1 76.82 104.59 77.31 ;
      RECT  106.495 60.12 106.985 60.61 ;
      RECT  64.21 109.955 64.7 110.445 ;
      RECT  140.975 64.87 141.465 65.36 ;
      RECT  174.485 96.095 174.975 96.585 ;
      RECT  107.03 126.5 107.33 126.8 ;
      RECT  174.485 102.02 174.975 102.51 ;
      RECT  195.425 94.12 195.915 94.61 ;
      RECT  174.485 107.945 174.975 108.435 ;
      RECT  138.23 126.5 138.53 126.8 ;
      RECT  99.73 72.63 100.22 73.12 ;
      RECT  116.39 89.29 116.69 89.59 ;
      RECT  124.69 142.97 125.18 143.46 ;
      RECT  130.99 138.78 131.48 139.27 ;
      RECT  64.21 113.905 64.7 114.395 ;
      RECT  147.495 89.195 147.985 89.685 ;
      RECT  174.485 111.895 174.975 112.385 ;
      RECT  106.595 64.87 107.085 65.36 ;
      RECT  124.75 76.82 125.24 77.31 ;
      RECT  137.23 138.78 137.72 139.27 ;
      RECT  103.91 126.5 104.21 126.8 ;
      RECT  185.555 98.07 186.045 98.56 ;
      RECT  112.27 76.82 112.76 77.31 ;
      RECT  97.92 142.97 98.41 143.46 ;
      RECT  56.395 98.07 56.885 98.56 ;
      RECT  185.555 109.92 186.045 110.41 ;
      RECT  107.53 86.24 108.02 86.73 ;
      RECT  188.81 98.105 189.3 98.595 ;
      RECT  137.17 142.97 137.66 143.46 ;
      RECT  97.67 89.29 97.97 89.59 ;
      RECT  104.16 72.63 104.65 73.12 ;
      RECT  103.635 60.12 104.125 60.61 ;
      RECT  116.58 76.82 117.07 77.31 ;
      RECT  100.355 64.87 100.845 65.36 ;
      RECT  64.21 117.855 64.7 118.345 ;
      RECT  177.74 121.805 178.23 122.295 ;
      RECT  118.45 142.97 118.94 143.46 ;
      RECT  195.425 105.97 195.915 106.46 ;
      RECT  118.51 76.82 119.0 77.31 ;
      RECT  67.465 109.92 67.955 110.41 ;
      RECT  143.41 72.63 143.9 73.12 ;
      RECT  143.47 138.78 143.96 139.27 ;
      RECT  97.295 64.87 97.785 65.36 ;
      RECT  137.23 76.82 137.72 77.31 ;
      RECT  135.3 76.82 135.79 77.31 ;
      RECT  103.22 129.36 103.71 129.85 ;
      RECT  99.79 138.78 100.28 139.27 ;
      RECT  67.465 94.12 67.955 94.61 ;
      RECT  64.21 96.255 64.7 96.745 ;
      RECT  110.15 126.5 110.45 126.8 ;
      RECT  177.74 108.105 178.23 108.595 ;
      RECT  56.395 94.12 56.885 94.61 ;
      RECT  131.99 126.5 132.29 126.8 ;
      RECT  99.73 142.97 100.22 143.46 ;
      RECT  100.255 60.12 100.745 60.61 ;
      RECT  107.53 129.36 108.02 129.85 ;
      RECT  107.03 89.29 107.33 89.59 ;
      RECT  67.465 111.895 67.955 112.385 ;
      RECT  97.86 138.78 98.35 139.27 ;
      RECT  103.91 89.29 104.21 89.59 ;
      RECT  105.97 72.63 106.46 73.12 ;
      RECT  116.015 64.87 116.505 65.36 ;
      RECT  143.41 142.97 143.9 143.46 ;
      RECT  141.54 138.78 142.03 139.27 ;
      RECT  121.94 86.24 122.43 86.73 ;
      RECT  135.3 138.78 135.79 139.27 ;
      RECT  64.21 94.155 64.7 94.645 ;
      RECT  67.465 121.77 67.955 122.26 ;
      RECT  67.465 103.995 67.955 104.485 ;
      RECT  109.775 64.87 110.265 65.36 ;
      RECT  174.485 115.845 174.975 116.335 ;
      RECT  98.15 57.905 98.64 58.395 ;
      RECT  140.66 86.24 141.15 86.73 ;
      RECT  97.67 126.5 97.97 126.8 ;
      RECT  132.49 86.24 132.98 86.73 ;
      RECT  188.81 94.155 189.3 94.645 ;
      RECT  96.98 86.24 97.47 86.73 ;
      RECT  122.88 72.63 123.37 73.12 ;
      RECT  128.495 64.87 128.985 65.36 ;
      RECT  97.92 72.63 98.41 73.12 ;
      RECT  174.485 94.12 174.975 94.61 ;
      RECT  135.11 89.29 135.41 89.59 ;
      RECT  122.255 64.87 122.745 65.36 ;
      RECT  119.51 89.29 119.81 89.59 ;
      RECT  174.485 109.92 174.975 110.41 ;
      RECT  141.6 72.63 142.09 73.12 ;
      RECT  119.075 64.87 119.565 65.36 ;
      RECT  110.34 138.78 110.83 139.27 ;
      RECT  115.7 86.24 116.19 86.73 ;
      RECT  144.97 86.24 145.46 86.73 ;
      RECT  122.82 76.82 123.31 77.31 ;
      RECT  105.97 142.97 106.46 143.46 ;
      RECT  113.77 129.36 114.26 129.85 ;
      RECT  138.73 129.36 139.22 129.85 ;
      RECT  53.14 109.955 53.63 110.445 ;
      RECT  157.295 107.8 157.785 108.29 ;
      RECT  125.75 89.29 126.05 89.59 ;
      RECT  95.05 86.24 95.54 86.73 ;
      RECT  144.47 89.29 144.77 89.59 ;
      RECT  177.74 119.955 178.23 120.445 ;
      RECT  67.465 98.07 67.955 98.56 ;
      RECT  97.86 76.82 98.35 77.31 ;
      RECT  141.075 60.12 141.565 60.61 ;
      RECT  177.74 113.905 178.23 114.395 ;
      RECT  96.98 129.36 97.47 129.85 ;
      RECT  118.51 138.78 119.0 139.27 ;
      RECT  112.21 142.97 112.7 143.46 ;
      RECT  140.66 129.36 141.15 129.85 ;
      RECT  106.03 138.78 106.52 139.27 ;
      RECT  112.835 64.87 113.325 65.36 ;
      RECT  101.29 86.24 101.78 86.73 ;
      RECT  118.975 60.12 119.465 60.61 ;
      RECT  128.18 129.36 128.67 129.85 ;
      RECT  177.74 117.855 178.23 118.345 ;
      RECT  46.525 94.12 47.015 94.61 ;
      RECT  174.485 98.07 174.975 98.56 ;
      RECT  46.525 105.97 47.015 106.46 ;
      RECT  110.4 72.63 110.89 73.12 ;
      RECT  67.465 102.02 67.955 102.51 ;
      RECT  143.47 76.82 143.96 77.31 ;
      RECT  141.35 126.5 141.65 126.8 ;
      RECT  130.93 72.63 131.42 73.12 ;
      RECT  174.485 100.045 174.975 100.535 ;
      RECT  177.74 104.155 178.23 104.645 ;
      RECT  103.22 86.24 103.71 86.73 ;
      RECT  118.45 72.63 118.94 73.12 ;
      RECT  64.21 121.805 64.7 122.295 ;
      RECT  53.14 106.005 53.63 106.495 ;
      RECT  67.465 105.97 67.955 106.46 ;
      RECT  122.63 126.5 122.93 126.8 ;
      RECT  134.42 129.36 134.91 129.85 ;
      RECT  110.15 89.29 110.45 89.59 ;
      RECT  144.97 129.36 145.46 129.85 ;
      RECT  174.485 117.82 174.975 118.31 ;
      RECT  174.485 103.995 174.975 104.485 ;
      RECT  126.25 86.24 126.74 86.73 ;
      RECT  120.01 86.24 120.5 86.73 ;
      RECT  67.465 117.82 67.955 118.31 ;
      RECT  67.465 119.795 67.955 120.285 ;
      RECT  130.99 76.82 131.48 77.31 ;
      RECT  141.54 76.82 142.03 77.31 ;
      RECT  132.49 129.36 132.98 129.85 ;
      RECT  106.03 76.82 106.52 77.31 ;
      RECT  67.465 113.87 67.955 114.36 ;
      RECT  128.87 126.5 129.17 126.8 ;
      RECT  119.51 126.5 119.81 126.8 ;
      RECT  135.11 126.5 135.41 126.8 ;
      RECT  129.12 72.63 129.61 73.12 ;
      RECT  94.455 126.405 94.945 126.895 ;
      RECT  121.94 129.36 122.43 129.85 ;
      RECT  112.27 138.78 112.76 139.27 ;
      RECT  113.27 89.29 113.57 89.59 ;
      RECT  56.395 109.92 56.885 110.41 ;
      RECT  110.34 76.82 110.83 77.31 ;
      RECT  64.21 112.055 64.7 112.545 ;
      RECT  71.82 107.72 72.31 108.21 ;
      RECT  116.115 60.12 116.605 60.61 ;
      RECT  137.695 60.12 138.185 60.61 ;
      RECT  122.355 60.12 122.845 60.61 ;
      RECT  64.21 106.005 64.7 106.495 ;
      RECT  137.17 72.63 137.66 73.12 ;
      RECT  109.46 129.36 109.95 129.85 ;
      RECT  64.21 108.105 64.7 108.595 ;
      RECT  64.21 100.205 64.7 100.695 ;
      RECT  100.79 126.5 101.09 126.8 ;
      RECT  130.93 142.97 131.42 143.46 ;
      RECT  135.36 142.97 135.85 143.46 ;
      RECT  64.21 119.955 64.7 120.445 ;
      RECT  113.27 126.5 113.57 126.8 ;
      RECT  67.465 100.045 67.955 100.535 ;
      RECT  128.18 86.24 128.67 86.73 ;
      RECT  141.6 142.97 142.09 143.46 ;
      RECT  110.4 142.97 110.89 143.46 ;
      RECT  137.795 64.87 138.285 65.36 ;
      RECT  125.75 126.5 126.05 126.8 ;
      RECT  177.74 109.955 178.23 110.445 ;
      RECT  144.035 64.87 144.525 65.36 ;
      RECT  109.875 60.12 110.365 60.61 ;
      RECT  146.9 129.36 147.39 129.85 ;
      RECT  56.395 105.97 56.885 106.46 ;
      RECT  174.485 113.87 174.975 114.36 ;
      RECT  122.88 142.97 123.37 143.46 ;
      RECT  84.655 107.8 85.145 108.29 ;
      RECT  123.11 57.905 123.6 58.395 ;
      RECT  177.74 96.255 178.23 96.745 ;
      RECT  116.64 142.97 117.13 143.46 ;
      RECT  91.07 122.51 91.37 122.81 ;
      RECT  104.14 63.21 104.63 63.7 ;
      RECT  66.105 117.82 66.595 118.31 ;
      RECT  175.845 121.77 176.335 122.26 ;
      RECT  136.82 80.69 137.31 81.18 ;
      RECT  124.69 144.58 125.18 145.07 ;
      RECT  128.55 67.055 129.04 67.545 ;
      RECT  151.07 122.51 151.37 122.81 ;
      RECT  130.95 63.21 131.44 63.7 ;
      RECT  62.085 106.005 62.575 106.495 ;
      RECT  66.105 94.12 66.595 94.61 ;
      RECT  175.845 94.12 176.335 94.61 ;
      RECT  99.38 80.69 99.87 81.18 ;
      RECT  135.71 134.91 136.2 135.4 ;
      RECT  123.11 52.305 123.6 52.795 ;
      RECT  119.02 67.055 119.51 67.545 ;
      RECT  97.9 63.21 98.39 63.7 ;
      RECT  151.07 109.08 151.37 109.38 ;
      RECT  104.51 80.69 105.0 81.18 ;
      RECT  91.07 94.86 91.37 95.16 ;
      RECT  55.035 94.12 55.525 94.61 ;
      RECT  105.97 144.58 106.46 145.07 ;
      RECT  51.015 106.005 51.505 106.495 ;
      RECT  66.105 121.77 66.595 122.26 ;
      RECT  186.915 98.07 187.405 98.56 ;
      RECT  110.4 71.02 110.89 71.51 ;
      RECT  151.07 120.93 151.37 121.23 ;
      RECT  105.62 134.91 106.11 135.4 ;
      RECT  129.47 80.69 129.96 81.18 ;
      RECT  143.06 80.69 143.55 81.18 ;
      RECT  122.285 62.2 122.775 62.69 ;
      RECT  186.915 94.12 187.405 94.61 ;
      RECT  116.99 134.91 117.48 135.4 ;
      RECT  122.88 144.58 123.37 145.07 ;
      RECT  97.35 67.055 97.84 67.545 ;
      RECT  130.58 80.69 131.07 81.18 ;
      RECT  98.27 80.69 98.76 81.18 ;
      RECT  151.07 103.945 151.37 104.245 ;
      RECT  175.845 113.87 176.335 114.36 ;
      RECT  123.23 80.69 123.72 81.18 ;
      RECT  129.47 134.91 129.96 135.4 ;
      RECT  190.935 94.155 191.425 94.645 ;
      RECT  137.17 144.58 137.66 145.07 ;
      RECT  112.21 144.58 112.7 145.07 ;
      RECT  97.325 62.2 97.815 62.69 ;
      RECT  91.07 99.995 91.37 100.295 ;
      RECT  116.62 63.21 117.11 63.7 ;
      RECT  151.07 94.86 151.37 95.16 ;
      RECT  151.07 106.71 151.37 107.01 ;
      RECT  62.085 121.805 62.575 122.295 ;
      RECT  99.73 144.58 100.22 145.07 ;
      RECT  66.105 113.87 66.595 114.36 ;
      RECT  99.38 134.91 99.87 135.4 ;
      RECT  62.085 115.995 62.575 116.485 ;
      RECT  190.935 106.005 191.425 106.495 ;
      RECT  125.285 62.2 125.775 62.69 ;
      RECT  172.255 107.725 172.745 108.215 ;
      RECT  141.95 134.91 142.44 135.4 ;
      RECT  116.045 62.2 116.535 62.69 ;
      RECT  151.07 118.56 151.37 118.86 ;
      RECT  105.99 63.21 106.48 63.7 ;
      RECT  151.07 115.795 151.37 116.095 ;
      RECT  91.07 118.56 91.37 118.86 ;
      RECT  112.23 63.21 112.72 63.7 ;
      RECT  175.845 98.07 176.335 98.56 ;
      RECT  135.71 80.69 136.2 81.18 ;
      RECT  175.845 117.82 176.335 118.31 ;
      RECT  99.75 63.21 100.24 63.7 ;
      RECT  179.865 104.145 180.355 104.635 ;
      RECT  143.98 67.055 144.47 67.545 ;
      RECT  119.045 62.2 119.535 62.69 ;
      RECT  110.38 63.21 110.87 63.7 ;
      RECT  45.165 105.97 45.655 106.46 ;
      RECT  179.865 115.995 180.355 116.485 ;
      RECT  66.105 115.845 66.595 116.335 ;
      RECT  103.565 62.2 104.055 62.69 ;
      RECT  62.085 112.045 62.575 112.535 ;
      RECT  141.005 62.2 141.495 62.69 ;
      RECT  99.73 71.02 100.22 71.51 ;
      RECT  136.82 134.91 137.31 135.4 ;
      RECT  91.07 98.81 91.37 99.11 ;
      RECT  151.07 113.03 151.37 113.33 ;
      RECT  112.805 62.2 113.295 62.69 ;
      RECT  135.36 71.02 135.85 71.51 ;
      RECT  179.865 108.095 180.355 108.585 ;
      RECT  91.07 116.98 91.37 117.28 ;
      RECT  143.06 134.91 143.55 135.4 ;
      RECT  151.07 92.095 151.37 92.395 ;
      RECT  118.47 63.21 118.96 63.7 ;
      RECT  141.6 144.58 142.09 145.07 ;
      RECT  151.07 114.61 151.37 114.91 ;
      RECT  110.75 80.69 111.24 81.18 ;
      RECT  112.21 71.02 112.7 71.51 ;
      RECT  55.035 105.97 55.525 106.46 ;
      RECT  105.97 71.02 106.46 71.51 ;
      RECT  62.085 119.945 62.575 120.435 ;
      RECT  179.865 119.945 180.355 120.435 ;
      RECT  151.07 119.745 151.37 120.045 ;
      RECT  91.07 92.095 91.37 92.395 ;
      RECT  151.07 116.98 151.37 117.28 ;
      RECT  118.45 144.58 118.94 145.07 ;
      RECT  62.085 98.105 62.575 98.595 ;
      RECT  66.105 111.895 66.595 112.385 ;
      RECT  110.75 134.91 111.24 135.4 ;
      RECT  116.07 67.055 116.56 67.545 ;
      RECT  179.865 94.155 180.355 94.645 ;
      RECT  122.86 63.21 123.35 63.7 ;
      RECT  91.07 103.945 91.37 104.245 ;
      RECT  116.64 144.58 117.13 145.07 ;
      RECT  91.07 105.13 91.37 105.43 ;
      RECT  112.78 67.055 113.27 67.545 ;
      RECT  125.26 67.055 125.75 67.545 ;
      RECT  129.12 144.58 129.61 145.07 ;
      RECT  91.07 111.845 91.37 112.145 ;
      RECT  66.105 105.97 66.595 106.46 ;
      RECT  141.6 71.02 142.09 71.51 ;
      RECT  179.865 106.005 180.355 106.495 ;
      RECT  104.16 144.58 104.65 145.07 ;
      RECT  131.525 62.2 132.015 62.69 ;
      RECT  129.12 71.02 129.61 71.51 ;
      RECT  69.695 107.725 70.185 108.215 ;
      RECT  62.085 100.195 62.575 100.685 ;
      RECT  143.41 144.58 143.9 145.07 ;
      RECT  91.07 114.61 91.37 114.91 ;
      RECT  175.845 111.895 176.335 112.385 ;
      RECT  179.865 96.245 180.355 96.735 ;
      RECT  66.105 102.02 66.595 102.51 ;
      RECT  66.105 103.995 66.595 104.485 ;
      RECT  141.03 67.055 141.52 67.545 ;
      RECT  179.865 112.045 180.355 112.535 ;
      RECT  118.1 80.69 118.59 81.18 ;
      RECT  116.99 80.69 117.48 81.18 ;
      RECT  135.34 63.21 135.83 63.7 ;
      RECT  51.015 98.105 51.505 98.595 ;
      RECT  118.1 134.91 118.59 135.4 ;
      RECT  144.005 62.2 144.495 62.69 ;
      RECT  109.83 67.055 110.32 67.545 ;
      RECT  179.865 98.105 180.355 98.595 ;
      RECT  122.88 71.02 123.37 71.51 ;
      RECT  100.325 62.2 100.815 62.69 ;
      RECT  116.64 71.02 117.13 71.51 ;
      RECT  124.71 63.21 125.2 63.7 ;
      RECT  103.59 67.055 104.08 67.545 ;
      RECT  141.95 80.69 142.44 81.18 ;
      RECT  66.105 100.045 66.595 100.535 ;
      RECT  91.07 96.045 91.37 96.345 ;
      RECT  62.085 104.145 62.575 104.635 ;
      RECT  124.69 71.02 125.18 71.51 ;
      RECT  151.07 111.845 151.37 112.145 ;
      RECT  91.07 97.23 91.37 97.53 ;
      RECT  186.915 109.92 187.405 110.41 ;
      RECT  151.07 97.23 151.37 97.53 ;
      RECT  106.54 67.055 107.03 67.545 ;
      RECT  118.45 71.02 118.94 71.51 ;
      RECT  55.035 98.07 55.525 98.56 ;
      RECT  151.07 90.91 151.37 91.21 ;
      RECT  104.16 71.02 104.65 71.51 ;
      RECT  137.17 71.02 137.66 71.51 ;
      RECT  97.92 144.58 98.41 145.07 ;
      RECT  91.07 119.745 91.37 120.045 ;
      RECT  190.935 109.955 191.425 110.445 ;
      RECT  91.07 90.91 91.37 91.21 ;
      RECT  179.865 102.055 180.355 102.545 ;
      RECT  66.105 119.795 66.595 120.285 ;
      RECT  134.765 62.2 135.255 62.69 ;
      RECT  123.23 134.91 123.72 135.4 ;
      RECT  62.085 109.955 62.575 110.445 ;
      RECT  105.62 80.69 106.11 81.18 ;
      RECT  151.07 105.13 151.37 105.43 ;
      RECT  104.51 134.91 105.0 135.4 ;
      RECT  124.34 134.91 124.83 135.4 ;
      RECT  111.86 80.69 112.35 81.18 ;
      RECT  110.4 144.58 110.89 145.07 ;
      RECT  62.085 102.055 62.575 102.545 ;
      RECT  55.035 109.92 55.525 110.41 ;
      RECT  77.035 107.8 77.525 108.29 ;
      RECT  62.085 96.245 62.575 96.735 ;
      RECT  179.865 109.955 180.355 110.445 ;
      RECT  179.865 113.905 180.355 114.395 ;
      RECT  175.845 115.845 176.335 116.335 ;
      RECT  141.58 63.21 142.07 63.7 ;
      RECT  66.105 107.945 66.595 108.435 ;
      RECT  179.865 100.195 180.355 100.685 ;
      RECT  175.845 105.97 176.335 106.46 ;
      RECT  175.845 100.045 176.335 100.535 ;
      RECT  91.07 107.895 91.37 108.195 ;
      RECT  100.3 67.055 100.79 67.545 ;
      RECT  122.31 67.055 122.8 67.545 ;
      RECT  151.07 96.045 151.37 96.345 ;
      RECT  130.93 144.58 131.42 145.07 ;
      RECT  186.915 105.97 187.405 106.46 ;
      RECT  97.92 71.02 98.41 71.51 ;
      RECT  151.07 102.76 151.37 103.06 ;
      RECT  62.085 113.905 62.575 114.395 ;
      RECT  175.845 119.795 176.335 120.285 ;
      RECT  111.86 134.91 112.35 135.4 ;
      RECT  129.1 63.21 129.59 63.7 ;
      RECT  175.845 102.02 176.335 102.51 ;
      RECT  151.07 110.66 151.37 110.96 ;
      RECT  128.525 62.2 129.015 62.69 ;
      RECT  91.07 101.18 91.37 101.48 ;
      RECT  151.07 93.28 151.37 93.58 ;
      RECT  98.15 52.305 98.64 52.795 ;
      RECT  51.015 109.955 51.505 110.445 ;
      RECT  98.27 134.91 98.76 135.4 ;
      RECT  143.43 63.21 143.92 63.7 ;
      RECT  137.765 62.2 138.255 62.69 ;
      RECT  175.845 107.945 176.335 108.435 ;
      RECT  190.935 98.105 191.425 98.595 ;
      RECT  164.915 107.8 165.405 108.29 ;
      RECT  91.07 109.08 91.37 109.38 ;
      RECT  91.07 106.71 91.37 107.01 ;
      RECT  137.74 67.055 138.23 67.545 ;
      RECT  62.085 108.095 62.575 108.585 ;
      RECT  134.79 67.055 135.28 67.545 ;
      RECT  91.07 120.93 91.37 121.23 ;
      RECT  137.19 63.21 137.68 63.7 ;
      RECT  62.085 117.855 62.575 118.345 ;
      RECT  175.845 96.095 176.335 96.585 ;
      RECT  91.07 124.88 91.37 125.18 ;
      RECT  66.105 98.07 66.595 98.56 ;
      RECT  151.07 123.695 151.37 123.995 ;
      RECT  91.07 93.28 91.37 93.58 ;
      RECT  91.07 113.03 91.37 113.33 ;
      RECT  143.41 71.02 143.9 71.51 ;
      RECT  130.93 71.02 131.42 71.51 ;
      RECT  124.34 80.69 124.83 81.18 ;
      RECT  51.015 94.155 51.505 94.645 ;
      RECT  91.07 102.76 91.37 103.06 ;
      RECT  151.07 101.18 151.37 101.48 ;
      RECT  131.5 67.055 131.99 67.545 ;
      RECT  135.36 144.58 135.85 145.07 ;
      RECT  62.085 94.155 62.575 94.645 ;
      RECT  175.845 103.995 176.335 104.485 ;
      RECT  179.865 121.805 180.355 122.295 ;
      RECT  151.07 99.995 151.37 100.295 ;
      RECT  106.565 62.2 107.055 62.69 ;
      RECT  66.105 109.92 66.595 110.41 ;
      RECT  91.07 123.695 91.37 123.995 ;
      RECT  91.07 110.66 91.37 110.96 ;
      RECT  179.865 117.855 180.355 118.345 ;
      RECT  91.07 115.795 91.37 116.095 ;
      RECT  196.785 105.97 197.275 106.46 ;
      RECT  109.805 62.2 110.295 62.69 ;
      RECT  45.165 94.12 45.655 94.61 ;
      RECT  151.07 107.895 151.37 108.195 ;
      RECT  130.58 134.91 131.07 135.4 ;
      RECT  196.785 94.12 197.275 94.61 ;
      RECT  175.845 109.92 176.335 110.41 ;
      RECT  151.07 98.81 151.37 99.11 ;
      RECT  66.105 96.095 66.595 96.585 ;
      RECT  151.07 124.88 151.37 125.18 ;
      RECT  0.375 37.76 0.865 38.25 ;
      RECT  0.375 30.68 0.865 31.17 ;
      RECT  0.375 44.84 0.865 45.33 ;
      RECT  3.105 127.25 2.615 127.74 ;
      RECT  6.785 138.45 6.295 138.94 ;
      RECT  3.105 116.05 2.615 116.54 ;
      RECT  3.105 138.45 2.615 138.94 ;
      RECT  3.105 104.85 2.615 105.34 ;
      RECT  3.105 104.85 2.615 105.34 ;
      RECT  6.785 93.65 6.295 94.14 ;
      RECT  3.105 93.65 2.615 94.14 ;
      RECT  6.785 104.85 6.295 105.34 ;
      RECT  6.785 104.85 6.295 105.34 ;
      RECT  6.785 116.05 6.295 116.54 ;
      RECT  6.785 93.65 6.295 94.14 ;
      RECT  3.105 93.65 2.615 94.14 ;
      RECT  6.785 127.25 6.295 127.74 ;
      RECT  3.105 88.05 2.615 88.54 ;
      RECT  3.105 110.45 2.615 110.94 ;
      RECT  6.785 99.25 6.295 99.74 ;
      RECT  6.785 132.85 6.295 133.34 ;
      RECT  6.785 88.05 6.295 88.54 ;
      RECT  3.105 132.85 2.615 133.34 ;
      RECT  6.785 110.45 6.295 110.94 ;
      RECT  3.105 121.65 2.615 122.14 ;
      RECT  6.785 121.65 6.295 122.14 ;
      RECT  3.105 99.25 2.615 99.74 ;
      RECT  6.295 93.65 6.785 94.14 ;
      RECT  39.485 37.76 39.975 38.25 ;
      RECT  6.295 116.05 6.785 116.54 ;
      RECT  39.485 80.18 39.975 80.67 ;
      RECT  6.295 138.45 6.785 138.94 ;
      RECT  2.615 116.05 3.105 116.54 ;
      RECT  6.295 127.25 6.785 127.74 ;
      RECT  2.615 93.65 3.105 94.14 ;
      RECT  39.485 66.04 39.975 66.53 ;
      RECT  6.295 104.85 6.785 105.34 ;
      RECT  2.615 104.85 3.105 105.34 ;
      RECT  0.375 37.76 0.865 38.25 ;
      RECT  39.485 51.9 39.975 52.39 ;
      RECT  2.615 138.45 3.105 138.94 ;
      RECT  2.615 127.25 3.105 127.74 ;
      RECT  6.295 132.85 6.785 133.34 ;
      RECT  39.485 58.97 39.975 59.46 ;
      RECT  6.295 99.25 6.785 99.74 ;
      RECT  6.295 110.45 6.785 110.94 ;
      RECT  0.375 30.68 0.865 31.17 ;
      RECT  2.615 121.65 3.105 122.14 ;
      RECT  6.295 88.05 6.785 88.54 ;
      RECT  6.295 121.65 6.785 122.14 ;
      RECT  2.615 110.45 3.105 110.94 ;
      RECT  0.375 44.84 0.865 45.33 ;
      RECT  2.615 99.25 3.105 99.74 ;
      RECT  39.485 44.83 39.975 45.32 ;
      RECT  39.485 87.25 39.975 87.74 ;
      RECT  39.485 30.69 39.975 31.18 ;
      RECT  39.485 73.11 39.975 73.6 ;
      RECT  2.615 88.05 3.105 88.54 ;
      RECT  2.615 132.85 3.105 133.34 ;
      RECT  240.985 164.19 240.495 163.7 ;
      RECT  240.985 171.27 240.495 170.78 ;
      RECT  238.255 88.84 238.745 88.35 ;
      RECT  234.575 77.64 235.065 77.15 ;
      RECT  238.255 100.04 238.745 99.55 ;
      RECT  238.255 77.64 238.745 77.15 ;
      RECT  238.255 111.24 238.745 110.75 ;
      RECT  238.255 111.24 238.745 110.75 ;
      RECT  234.575 122.44 235.065 121.95 ;
      RECT  238.255 122.44 238.745 121.95 ;
      RECT  234.575 111.24 235.065 110.75 ;
      RECT  234.575 111.24 235.065 110.75 ;
      RECT  234.575 100.04 235.065 99.55 ;
      RECT  234.575 122.44 235.065 121.95 ;
      RECT  238.255 122.44 238.745 121.95 ;
      RECT  234.575 88.84 235.065 88.35 ;
      RECT  238.255 128.04 238.745 127.55 ;
      RECT  238.255 105.64 238.745 105.15 ;
      RECT  234.575 116.84 235.065 116.35 ;
      RECT  234.575 83.24 235.065 82.75 ;
      RECT  234.575 128.04 235.065 127.55 ;
      RECT  238.255 83.24 238.745 82.75 ;
      RECT  234.575 105.64 235.065 105.15 ;
      RECT  238.255 94.44 238.745 93.95 ;
      RECT  234.575 94.44 235.065 93.95 ;
      RECT  238.255 116.84 238.745 116.35 ;
      RECT  203.375 164.19 202.885 163.7 ;
      RECT  238.745 111.24 238.255 110.75 ;
      RECT  235.065 88.84 234.575 88.35 ;
      RECT  235.065 111.24 234.575 110.75 ;
      RECT  235.065 122.44 234.575 121.95 ;
      RECT  235.065 77.64 234.575 77.15 ;
      RECT  203.375 150.05 202.885 149.56 ;
      RECT  238.745 100.04 238.255 99.55 ;
      RECT  240.985 164.19 240.495 163.7 ;
      RECT  235.065 100.04 234.575 99.55 ;
      RECT  238.745 88.84 238.255 88.35 ;
      RECT  203.375 135.91 202.885 135.42 ;
      RECT  238.745 77.64 238.255 77.15 ;
      RECT  238.745 122.44 238.255 121.95 ;
      RECT  238.745 116.84 238.255 116.35 ;
      RECT  238.745 83.24 238.255 82.75 ;
      RECT  235.065 116.84 234.575 116.35 ;
      RECT  235.065 105.64 234.575 105.15 ;
      RECT  235.065 94.44 234.575 93.95 ;
      RECT  203.375 128.84 202.885 128.35 ;
      RECT  203.375 142.98 202.885 142.49 ;
      RECT  235.065 83.24 234.575 82.75 ;
      RECT  238.745 94.44 238.255 93.95 ;
      RECT  238.745 128.04 238.255 127.55 ;
      RECT  240.985 171.27 240.495 170.78 ;
      RECT  238.745 105.64 238.255 105.15 ;
      RECT  203.375 171.26 202.885 170.77 ;
      RECT  235.065 128.04 234.575 127.55 ;
      RECT  203.375 157.12 202.885 156.63 ;
      RECT  34.31 140.885 40.15 141.185 ;
      RECT  36.985 146.32 37.475 146.81 ;
      RECT  36.985 160.46 37.475 160.95 ;
      RECT  36.985 167.53 37.475 168.02 ;
      RECT  36.985 139.25 37.475 139.74 ;
      RECT  36.985 153.39 37.475 153.88 ;
      RECT  208.55 75.205 202.71 74.905 ;
      RECT  205.875 69.77 205.385 69.28 ;
      RECT  205.875 55.63 205.385 55.14 ;
      RECT  205.875 48.56 205.385 48.07 ;
      RECT  205.875 76.84 205.385 76.35 ;
      RECT  205.875 62.7 205.385 62.21 ;
      RECT  45.99 1.73 57.67 2.03 ;
      RECT  48.665 7.165 49.155 7.655 ;
      RECT  54.505 7.165 54.995 7.655 ;
      RECT  54.505 0.095 54.995 0.585 ;
      RECT  48.665 0.095 49.155 0.585 ;
      RECT  57.67 1.73 151.11 2.03 ;
      RECT  136.265 7.165 136.755 7.655 ;
      RECT  142.105 7.165 142.595 7.655 ;
      RECT  147.945 7.165 148.435 7.655 ;
      RECT  72.025 7.165 72.515 7.655 ;
      RECT  118.745 7.165 119.235 7.655 ;
      RECT  130.425 7.165 130.915 7.655 ;
      RECT  89.545 7.165 90.035 7.655 ;
      RECT  107.065 7.165 107.555 7.655 ;
      RECT  124.585 7.165 125.075 7.655 ;
      RECT  66.185 7.165 66.675 7.655 ;
      RECT  101.225 7.165 101.715 7.655 ;
      RECT  60.345 7.165 60.835 7.655 ;
      RECT  112.905 7.165 113.395 7.655 ;
      RECT  95.385 7.165 95.875 7.655 ;
      RECT  77.865 7.165 78.355 7.655 ;
      RECT  83.705 7.165 84.195 7.655 ;
      RECT  83.705 0.095 84.195 0.585 ;
      RECT  118.745 0.095 119.235 0.585 ;
      RECT  77.865 0.095 78.355 0.585 ;
      RECT  60.345 0.095 60.835 0.585 ;
      RECT  107.065 0.095 107.555 0.585 ;
      RECT  72.025 0.095 72.515 0.585 ;
      RECT  112.905 0.095 113.395 0.585 ;
      RECT  124.585 0.095 125.075 0.585 ;
      RECT  89.545 0.095 90.035 0.585 ;
      RECT  142.105 0.095 142.595 0.585 ;
      RECT  66.185 0.095 66.675 0.585 ;
      RECT  95.385 0.095 95.875 0.585 ;
      RECT  101.225 0.095 101.715 0.585 ;
      RECT  147.945 0.095 148.435 0.585 ;
      RECT  136.265 0.095 136.755 0.585 ;
      RECT  130.425 0.095 130.915 0.585 ;
   LAYER  m4 ;
   END
   END    sram_16_16_sky130_0.05
END    LIBRARY
