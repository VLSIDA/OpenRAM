magic
tech sky130A
magscale 1 2
timestamp 1595931502
<< checkpaint >>
rect -1302 -1260 1884 9160
<< ndiffc >>
rect 404 7488 438 7490
rect 14 7331 17 7363
rect 463 7331 466 7363
rect 596 7331 599 7363
rect 42 7204 76 7206
rect 42 7172 76 7174
rect 42 7046 76 7048
rect 42 7014 76 7016
rect 14 6857 17 6889
rect 463 6857 466 6889
rect 596 6857 599 6889
rect 42 6698 76 6732
rect 404 6698 438 6732
rect 14 6541 17 6573
rect 463 6541 466 6573
rect 596 6541 599 6573
rect 42 6414 76 6416
rect 42 6382 76 6384
rect 42 6256 76 6258
rect 42 6224 76 6226
rect 14 6067 17 6099
rect 463 6067 466 6099
rect 596 6067 599 6099
rect 42 5908 76 5942
rect 404 5908 438 5942
rect 14 5751 17 5783
rect 463 5751 466 5783
rect 596 5751 599 5783
rect 42 5624 76 5626
rect 42 5592 76 5594
rect 42 5466 76 5468
rect 42 5434 76 5436
rect 14 5277 17 5309
rect 463 5277 466 5309
rect 596 5277 599 5309
rect 42 5118 76 5152
rect 404 5118 438 5152
rect 14 4961 17 4993
rect 463 4961 466 4993
rect 596 4961 599 4993
rect 42 4834 76 4836
rect 42 4802 76 4804
rect 42 4676 76 4678
rect 42 4644 76 4646
rect 14 4487 17 4519
rect 463 4487 466 4519
rect 596 4487 599 4519
rect 42 4328 76 4362
rect 404 4328 438 4362
rect 14 4171 17 4203
rect 463 4171 466 4203
rect 596 4171 599 4203
rect 42 4044 76 4046
rect 42 4012 76 4014
rect 42 3886 76 3888
rect 42 3854 76 3856
rect 14 3697 17 3729
rect 463 3697 466 3729
rect 596 3697 599 3729
rect 42 3538 76 3572
rect 404 3538 438 3572
rect 14 3381 17 3413
rect 463 3381 466 3413
rect 596 3381 599 3413
rect 42 3254 76 3256
rect 42 3222 76 3224
rect 42 3096 76 3098
rect 42 3064 76 3066
rect 14 2907 17 2939
rect 463 2907 466 2939
rect 596 2907 599 2939
rect 42 2748 76 2782
rect 404 2748 438 2782
rect 14 2591 17 2623
rect 463 2591 466 2623
rect 596 2591 599 2623
rect 42 2464 76 2466
rect 42 2432 76 2434
rect 42 2306 76 2308
rect 42 2274 76 2276
rect 14 2117 17 2149
rect 463 2117 466 2149
rect 596 2117 599 2149
rect 42 1958 76 1992
rect 404 1958 438 1992
rect 14 1801 17 1833
rect 463 1801 466 1833
rect 596 1801 599 1833
rect 42 1674 76 1676
rect 42 1642 76 1644
rect 42 1516 76 1518
rect 42 1484 76 1486
rect 14 1327 17 1359
rect 463 1327 466 1359
rect 596 1327 599 1359
rect 42 1168 76 1202
rect 404 1168 438 1202
rect 14 1011 17 1043
rect 463 1011 466 1043
rect 596 1011 599 1043
rect 42 884 76 886
rect 42 852 76 854
rect 42 726 76 728
rect 42 694 76 696
rect 596 537 599 569
rect 404 410 438 412
<< locali >>
rect 42 7505 76 7522
rect 404 7505 438 7520
rect 193 7411 196 7445
rect 224 7411 227 7445
rect -14 7363 14 7364
rect -14 7331 0 7363
rect -14 7330 14 7331
rect 107 7323 109 7351
rect 139 7317 141 7351
rect 193 7330 196 7364
rect 224 7330 227 7364
rect 271 7334 278 7368
rect 339 7343 341 7377
rect 371 7343 373 7371
rect 466 7363 497 7364
rect 565 7363 596 7364
rect 466 7330 497 7331
rect 565 7330 596 7331
rect 193 7249 196 7283
rect 224 7249 227 7283
rect 193 6937 196 6971
rect 224 6937 227 6971
rect -14 6889 14 6890
rect -14 6857 0 6889
rect 107 6869 109 6897
rect 139 6869 141 6903
rect -14 6856 14 6857
rect 193 6856 196 6890
rect 224 6856 227 6890
rect 466 6889 497 6890
rect 565 6889 596 6890
rect 271 6852 278 6886
rect 339 6843 341 6877
rect 371 6849 373 6877
rect 466 6856 497 6857
rect 565 6856 596 6857
rect 193 6775 196 6809
rect 224 6775 227 6809
rect 193 6621 196 6655
rect 224 6621 227 6655
rect -14 6573 14 6574
rect -14 6541 0 6573
rect -14 6540 14 6541
rect 107 6533 109 6561
rect 139 6527 141 6561
rect 193 6540 196 6574
rect 224 6540 227 6574
rect 271 6544 278 6578
rect 339 6553 341 6587
rect 371 6553 373 6581
rect 466 6573 497 6574
rect 565 6573 596 6574
rect 466 6540 497 6541
rect 565 6540 596 6541
rect 193 6459 196 6493
rect 224 6459 227 6493
rect 193 6147 196 6181
rect 224 6147 227 6181
rect -14 6099 14 6100
rect -14 6067 0 6099
rect 107 6079 109 6107
rect 139 6079 141 6113
rect -14 6066 14 6067
rect 193 6066 196 6100
rect 224 6066 227 6100
rect 466 6099 497 6100
rect 565 6099 596 6100
rect 271 6062 278 6096
rect 339 6053 341 6087
rect 371 6059 373 6087
rect 466 6066 497 6067
rect 565 6066 596 6067
rect 193 5985 196 6019
rect 224 5985 227 6019
rect 193 5831 196 5865
rect 224 5831 227 5865
rect -14 5783 14 5784
rect -14 5751 0 5783
rect -14 5750 14 5751
rect 107 5743 109 5771
rect 139 5737 141 5771
rect 193 5750 196 5784
rect 224 5750 227 5784
rect 271 5754 278 5788
rect 339 5763 341 5797
rect 371 5763 373 5791
rect 466 5783 497 5784
rect 565 5783 596 5784
rect 466 5750 497 5751
rect 565 5750 596 5751
rect 193 5669 196 5703
rect 224 5669 227 5703
rect 193 5357 196 5391
rect 224 5357 227 5391
rect -14 5309 14 5310
rect -14 5277 0 5309
rect 107 5289 109 5317
rect 139 5289 141 5323
rect -14 5276 14 5277
rect 193 5276 196 5310
rect 224 5276 227 5310
rect 466 5309 497 5310
rect 565 5309 596 5310
rect 271 5272 278 5306
rect 339 5263 341 5297
rect 371 5269 373 5297
rect 466 5276 497 5277
rect 565 5276 596 5277
rect 193 5195 196 5229
rect 224 5195 227 5229
rect 193 5041 196 5075
rect 224 5041 227 5075
rect -14 4993 14 4994
rect -14 4961 0 4993
rect -14 4960 14 4961
rect 107 4953 109 4981
rect 139 4947 141 4981
rect 193 4960 196 4994
rect 224 4960 227 4994
rect 271 4964 278 4998
rect 339 4973 341 5007
rect 371 4973 373 5001
rect 466 4993 497 4994
rect 565 4993 596 4994
rect 466 4960 497 4961
rect 565 4960 596 4961
rect 193 4879 196 4913
rect 224 4879 227 4913
rect 193 4567 196 4601
rect 224 4567 227 4601
rect -14 4519 14 4520
rect -14 4487 0 4519
rect 107 4499 109 4527
rect 139 4499 141 4533
rect -14 4486 14 4487
rect 193 4486 196 4520
rect 224 4486 227 4520
rect 466 4519 497 4520
rect 565 4519 596 4520
rect 271 4482 278 4516
rect 339 4473 341 4507
rect 371 4479 373 4507
rect 466 4486 497 4487
rect 565 4486 596 4487
rect 193 4405 196 4439
rect 224 4405 227 4439
rect 193 4251 196 4285
rect 224 4251 227 4285
rect -14 4203 14 4204
rect -14 4171 0 4203
rect -14 4170 14 4171
rect 107 4163 109 4191
rect 139 4157 141 4191
rect 193 4170 196 4204
rect 224 4170 227 4204
rect 271 4174 278 4208
rect 339 4183 341 4217
rect 371 4183 373 4211
rect 466 4203 497 4204
rect 565 4203 596 4204
rect 466 4170 497 4171
rect 565 4170 596 4171
rect 193 4089 196 4123
rect 224 4089 227 4123
rect 193 3777 196 3811
rect 224 3777 227 3811
rect -14 3729 14 3730
rect -14 3697 0 3729
rect 107 3709 109 3737
rect 139 3709 141 3743
rect -14 3696 14 3697
rect 193 3696 196 3730
rect 224 3696 227 3730
rect 466 3729 497 3730
rect 565 3729 596 3730
rect 271 3692 278 3726
rect 339 3683 341 3717
rect 371 3689 373 3717
rect 466 3696 497 3697
rect 565 3696 596 3697
rect 193 3615 196 3649
rect 224 3615 227 3649
rect 193 3461 196 3495
rect 224 3461 227 3495
rect -14 3413 14 3414
rect -14 3381 0 3413
rect -14 3380 14 3381
rect 107 3373 109 3401
rect 139 3367 141 3401
rect 193 3380 196 3414
rect 224 3380 227 3414
rect 271 3384 278 3418
rect 339 3393 341 3427
rect 371 3393 373 3421
rect 466 3413 497 3414
rect 565 3413 596 3414
rect 466 3380 497 3381
rect 565 3380 596 3381
rect 193 3299 196 3333
rect 224 3299 227 3333
rect 193 2987 196 3021
rect 224 2987 227 3021
rect -14 2939 14 2940
rect -14 2907 0 2939
rect 107 2919 109 2947
rect 139 2919 141 2953
rect -14 2906 14 2907
rect 193 2906 196 2940
rect 224 2906 227 2940
rect 466 2939 497 2940
rect 565 2939 596 2940
rect 271 2902 278 2936
rect 339 2893 341 2927
rect 371 2899 373 2927
rect 466 2906 497 2907
rect 565 2906 596 2907
rect 193 2825 196 2859
rect 224 2825 227 2859
rect 193 2671 196 2705
rect 224 2671 227 2705
rect -14 2623 14 2624
rect -14 2591 0 2623
rect -14 2590 14 2591
rect 107 2583 109 2611
rect 139 2577 141 2611
rect 193 2590 196 2624
rect 224 2590 227 2624
rect 271 2594 278 2628
rect 339 2603 341 2637
rect 371 2603 373 2631
rect 466 2623 497 2624
rect 565 2623 596 2624
rect 466 2590 497 2591
rect 565 2590 596 2591
rect 193 2509 196 2543
rect 224 2509 227 2543
rect 193 2197 196 2231
rect 224 2197 227 2231
rect -14 2149 14 2150
rect -14 2117 0 2149
rect 107 2129 109 2157
rect 139 2129 141 2163
rect -14 2116 14 2117
rect 193 2116 196 2150
rect 224 2116 227 2150
rect 466 2149 497 2150
rect 565 2149 596 2150
rect 271 2112 278 2146
rect 339 2103 341 2137
rect 371 2109 373 2137
rect 466 2116 497 2117
rect 565 2116 596 2117
rect 193 2035 196 2069
rect 224 2035 227 2069
rect 193 1881 196 1915
rect 224 1881 227 1915
rect -14 1833 14 1834
rect -14 1801 0 1833
rect -14 1800 14 1801
rect 107 1793 109 1821
rect 139 1787 141 1821
rect 193 1800 196 1834
rect 224 1800 227 1834
rect 271 1804 278 1838
rect 339 1813 341 1847
rect 371 1813 373 1841
rect 466 1833 497 1834
rect 565 1833 596 1834
rect 466 1800 497 1801
rect 565 1800 596 1801
rect 193 1719 196 1753
rect 224 1719 227 1753
rect 193 1407 196 1441
rect 224 1407 227 1441
rect -14 1359 14 1360
rect -14 1327 0 1359
rect 107 1339 109 1367
rect 139 1339 141 1373
rect -14 1326 14 1327
rect 193 1326 196 1360
rect 224 1326 227 1360
rect 466 1359 497 1360
rect 565 1359 596 1360
rect 271 1322 278 1356
rect 339 1313 341 1347
rect 371 1319 373 1347
rect 466 1326 497 1327
rect 565 1326 596 1327
rect 193 1245 196 1279
rect 224 1245 227 1279
rect 193 1091 196 1125
rect 224 1091 227 1125
rect -14 1043 14 1044
rect -14 1011 0 1043
rect -14 1010 14 1011
rect 107 1003 109 1031
rect 139 997 141 1031
rect 193 1010 196 1044
rect 224 1010 227 1044
rect 271 1014 278 1048
rect 339 1023 341 1057
rect 371 1023 373 1051
rect 466 1043 497 1044
rect 565 1043 596 1044
rect 466 1010 497 1011
rect 565 1010 596 1011
rect 193 929 196 963
rect 224 929 227 963
rect -14 569 17 570
rect -14 537 0 569
rect 107 549 109 577
rect 139 549 141 583
rect 463 569 497 570
rect 565 569 596 570
rect -14 536 17 537
rect 339 523 341 557
rect 371 529 373 557
rect 463 536 497 537
rect 565 536 596 537
rect 42 378 76 395
rect 404 380 438 395
<< metal1 >>
rect 78 0 114 7900
rect 150 0 186 7900
rect 222 7189 258 7530
rect 222 6399 258 7031
rect 222 5609 258 6241
rect 222 4819 258 5451
rect 222 4029 258 4661
rect 222 3239 258 3871
rect 222 2449 258 3081
rect 222 1659 258 2291
rect 222 869 258 1501
rect 222 370 258 711
rect 294 0 330 7900
rect 366 0 402 7900
<< metal2 >>
rect 0 7433 624 7481
rect 186 7309 294 7385
rect 0 7213 624 7261
rect 186 7055 294 7165
rect 0 6959 624 7007
rect 186 6835 294 6911
rect 0 6739 624 6787
rect 0 6643 624 6691
rect 186 6519 294 6595
rect 0 6423 624 6471
rect 186 6265 294 6375
rect 0 6169 624 6217
rect 186 6045 294 6121
rect 0 5949 624 5997
rect 0 5853 624 5901
rect 186 5729 294 5805
rect 0 5633 624 5681
rect 186 5475 294 5585
rect 0 5379 624 5427
rect 186 5255 294 5331
rect 0 5159 624 5207
rect 0 5063 624 5111
rect 186 4939 294 5015
rect 0 4843 624 4891
rect 186 4685 294 4795
rect 0 4589 624 4637
rect 186 4465 294 4541
rect 0 4369 624 4417
rect 0 4273 624 4321
rect 186 4149 294 4225
rect 0 4053 624 4101
rect 186 3895 294 4005
rect 0 3799 624 3847
rect 186 3675 294 3751
rect 0 3579 624 3627
rect 0 3483 624 3531
rect 186 3359 294 3435
rect 0 3263 624 3311
rect 186 3105 294 3215
rect 0 3009 624 3057
rect 186 2885 294 2961
rect 0 2789 624 2837
rect 0 2693 624 2741
rect 186 2569 294 2645
rect 0 2473 624 2521
rect 186 2315 294 2425
rect 0 2219 624 2267
rect 186 2095 294 2171
rect 0 1999 624 2047
rect 0 1903 624 1951
rect 186 1779 294 1855
rect 0 1683 624 1731
rect 186 1525 294 1635
rect 0 1429 624 1477
rect 186 1305 294 1381
rect 0 1209 624 1257
rect 0 1113 624 1161
rect 186 989 294 1065
rect 0 893 624 941
rect 186 735 294 845
rect 0 639 624 687
rect 186 515 294 591
rect 0 419 624 467
<< metal3 >>
rect 263 7622 361 7720
rect 263 180 361 278
use contact_9  contact_9_1
timestamp 1595931502
transform 1 0 279 0 1 192
box 0 0 66 74
use contact_9  contact_9_0
timestamp 1595931502
transform 1 0 279 0 1 7634
box 0 0 66 74
use col_cap_cell_1rw_1r  col_cap_cell_1rw_1r_0
timestamp 1595931502
transform 1 0 0 0 -1 7900
box 0 0 624 474
use replica_cell_1rw_1r  replica_cell_1rw_1r_0
timestamp 1595931502
transform 1 0 0 0 1 7110
box -42 -104 624 420
use replica_cell_1rw_1r  replica_cell_1rw_1r_1
timestamp 1595931502
transform 1 0 0 0 -1 7110
box -42 -104 624 420
use replica_cell_1rw_1r  replica_cell_1rw_1r_2
timestamp 1595931502
transform 1 0 0 0 1 6320
box -42 -104 624 420
use replica_cell_1rw_1r  replica_cell_1rw_1r_3
timestamp 1595931502
transform 1 0 0 0 -1 6320
box -42 -104 624 420
use replica_cell_1rw_1r  replica_cell_1rw_1r_4
timestamp 1595931502
transform 1 0 0 0 1 5530
box -42 -104 624 420
use replica_cell_1rw_1r  replica_cell_1rw_1r_5
timestamp 1595931502
transform 1 0 0 0 -1 5530
box -42 -104 624 420
use replica_cell_1rw_1r  replica_cell_1rw_1r_6
timestamp 1595931502
transform 1 0 0 0 1 4740
box -42 -104 624 420
use replica_cell_1rw_1r  replica_cell_1rw_1r_7
timestamp 1595931502
transform 1 0 0 0 -1 4740
box -42 -104 624 420
use replica_cell_1rw_1r  replica_cell_1rw_1r_8
timestamp 1595931502
transform 1 0 0 0 1 3950
box -42 -104 624 420
use replica_cell_1rw_1r  replica_cell_1rw_1r_9
timestamp 1595931502
transform 1 0 0 0 -1 3950
box -42 -104 624 420
use replica_cell_1rw_1r  replica_cell_1rw_1r_10
timestamp 1595931502
transform 1 0 0 0 1 3160
box -42 -104 624 420
use replica_cell_1rw_1r  replica_cell_1rw_1r_11
timestamp 1595931502
transform 1 0 0 0 -1 3160
box -42 -104 624 420
use replica_cell_1rw_1r  replica_cell_1rw_1r_12
timestamp 1595931502
transform 1 0 0 0 1 2370
box -42 -104 624 420
use replica_cell_1rw_1r  replica_cell_1rw_1r_13
timestamp 1595931502
transform 1 0 0 0 -1 2370
box -42 -104 624 420
use replica_cell_1rw_1r  replica_cell_1rw_1r_14
timestamp 1595931502
transform 1 0 0 0 1 1580
box -42 -104 624 420
use replica_cell_1rw_1r  replica_cell_1rw_1r_15
timestamp 1595931502
transform 1 0 0 0 -1 1580
box -42 -104 624 420
use replica_cell_1rw_1r  replica_cell_1rw_1r_16
timestamp 1595931502
transform 1 0 0 0 1 790
box -42 -104 624 420
use dummy_cell_1rw_1r  dummy_cell_1rw_1r_0
timestamp 1595931502
transform 1 0 0 0 -1 790
box -42 -104 624 420
use col_cap_cell_1rw_1r  col_cap_cell_1rw_1r_1
timestamp 1595931502
transform 1 0 0 0 1 0
box 0 0 624 474
<< labels >>
rlabel metal2 s 312 6667 312 6667 4 wl0_16
rlabel metal2 s 312 4613 312 4613 4 wl1_11
rlabel metal2 s 312 6193 312 6193 4 wl1_15
rlabel metal2 s 312 1927 312 1927 4 wl0_4
rlabel metal2 s 312 917 312 917 4 wl1_2
rlabel metal2 s 312 7237 312 7237 4 wl1_18
rlabel metal2 s 312 5403 312 5403 4 wl1_13
rlabel metal1 s 168 3950 168 3950 4 br0
rlabel metal2 s 312 3823 312 3823 4 wl1_9
rlabel metal2 s 312 663 312 663 4 wl1_1
rlabel metal2 s 312 1453 312 1453 4 wl1_3
rlabel metal2 s 312 3033 312 3033 4 wl1_7
rlabel metal1 s 312 3950 312 3950 4 bl1
rlabel metal2 s 312 5657 312 5657 4 wl1_14
rlabel metal2 s 312 4393 312 4393 4 wl0_11
rlabel metal2 s 312 7457 312 7457 4 wl0_18
rlabel metal2 s 312 6447 312 6447 4 wl1_16
rlabel metal2 s 312 4077 312 4077 4 wl1_10
rlabel metal2 s 312 1707 312 1707 4 wl1_4
rlabel metal2 s 312 1233 312 1233 4 wl0_3
rlabel metal2 s 240 3397 240 3397 4 gnd
rlabel metal2 s 240 1027 240 1027 4 gnd
rlabel metal2 s 240 3713 240 3713 4 gnd
rlabel metal2 s 240 553 240 553 4 gnd
rlabel metal2 s 240 3160 240 3160 4 gnd
rlabel metal2 s 240 2923 240 2923 4 gnd
rlabel metal2 s 240 4187 240 4187 4 gnd
rlabel metal2 s 240 4740 240 4740 4 gnd
rlabel metal2 s 240 5767 240 5767 4 gnd
rlabel metal2 s 240 1343 240 1343 4 gnd
rlabel metal2 s 240 2133 240 2133 4 gnd
rlabel metal2 s 240 6320 240 6320 4 gnd
rlabel metal2 s 240 2370 240 2370 4 gnd
rlabel metal2 s 240 4977 240 4977 4 gnd
rlabel metal2 s 240 6557 240 6557 4 gnd
rlabel metal2 s 240 3950 240 3950 4 gnd
rlabel metal2 s 240 2607 240 2607 4 gnd
rlabel metal2 s 240 5530 240 5530 4 gnd
rlabel metal2 s 240 790 240 790 4 gnd
rlabel metal2 s 240 6083 240 6083 4 gnd
rlabel metal2 s 240 1580 240 1580 4 gnd
rlabel metal2 s 240 5293 240 5293 4 gnd
rlabel metal2 s 240 1817 240 1817 4 gnd
rlabel metal2 s 240 4503 240 4503 4 gnd
rlabel metal2 s 240 7110 240 7110 4 gnd
rlabel metal2 s 240 7347 240 7347 4 gnd
rlabel metal2 s 240 6873 240 6873 4 gnd
rlabel metal2 s 312 2497 312 2497 4 wl1_6
rlabel metal2 s 312 2717 312 2717 4 wl0_6
rlabel metal2 s 312 6763 312 6763 4 wl0_17
rlabel metal2 s 312 3603 312 3603 4 wl0_9
rlabel metal2 s 312 2813 312 2813 4 wl0_7
rlabel metal1 s 240 2120 240 2120 4 vdd
rlabel metal1 s 240 7359 240 7359 4 vdd
rlabel metal3 s 312 229 312 229 4 vdd
rlabel metal1 s 240 4989 240 4989 4 vdd
rlabel metal1 s 240 2619 240 2619 4 vdd
rlabel metal1 s 240 540 240 540 4 vdd
rlabel metal1 s 240 6569 240 6569 4 vdd
rlabel metal1 s 240 6860 240 6860 4 vdd
rlabel metal1 s 240 3409 240 3409 4 vdd
rlabel metal1 s 240 1330 240 1330 4 vdd
rlabel metal1 s 240 2910 240 2910 4 vdd
rlabel metal1 s 240 1829 240 1829 4 vdd
rlabel metal1 s 240 4199 240 4199 4 vdd
rlabel metal1 s 240 5280 240 5280 4 vdd
rlabel metal1 s 240 5779 240 5779 4 vdd
rlabel metal1 s 240 3700 240 3700 4 vdd
rlabel metal3 s 312 7671 312 7671 4 vdd
rlabel metal1 s 240 6070 240 6070 4 vdd
rlabel metal1 s 240 1039 240 1039 4 vdd
rlabel metal1 s 240 4490 240 4490 4 vdd
rlabel metal2 s 312 5973 312 5973 4 wl0_15
rlabel metal2 s 312 3287 312 3287 4 wl1_8
rlabel metal2 s 312 5087 312 5087 4 wl0_12
rlabel metal2 s 312 4867 312 4867 4 wl1_12
rlabel metal2 s 312 5877 312 5877 4 wl0_14
rlabel metal2 s 312 2243 312 2243 4 wl1_5
rlabel metal2 s 312 6983 312 6983 4 wl1_17
rlabel metal2 s 312 2023 312 2023 4 wl0_5
rlabel metal2 s 312 5183 312 5183 4 wl0_13
rlabel metal2 s 312 443 312 443 4 wl0_1
rlabel metal2 s 312 1137 312 1137 4 wl0_2
rlabel metal1 s 384 3950 384 3950 4 br1
rlabel metal2 s 312 4297 312 4297 4 wl0_10
rlabel metal2 s 312 3507 312 3507 4 wl0_8
rlabel metal1 s 96 3950 96 3950 4 bl0
<< properties >>
string FIXED_BBOX 0 0 624 7900
<< end >>
