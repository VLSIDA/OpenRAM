**************************************************
* OpenRAM generated memory.
* Words: 1024
* Data bits: 128
* Banks: 4
* Column mux: 2:1
**************************************************

* ptx M{0} {1} n m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p

* ptx M{0} {1} p m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p

.SUBCKT pnand2_1 A B Z vdd gnd
Mpnand2_pmos1 vdd A Z vdd p m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpnand2_pmos2 Z B vdd vdd p m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpnand2_nmos1 Z B net1 gnd n m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpnand2_nmos2 net1 A gnd gnd n m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
.ENDS pnand2_1

.SUBCKT pnand3_1 A B C Z vdd gnd
Mpnand3_pmos1 vdd A Z vdd p m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpnand3_pmos2 Z B vdd vdd p m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpnand3_pmos3 Z C vdd vdd p m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpnand3_nmos1 Z C net1 gnd n m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpnand3_nmos2 net1 B net2 gnd n m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpnand3_nmos3 net2 A gnd gnd n m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
.ENDS pnand3_1

* ptx M{0} {1} n m=1 w=1.2u l=0.6u pd=3.6u ps=3.6u as=1.8p ad=1.8p

* ptx M{0} {1} p m=1 w=3.6u l=0.6u pd=8.4u ps=8.4u as=5.4p ad=5.4p

.SUBCKT pnor2_1 A B Z vdd gnd
Mpnor2_pmos1 vdd A net1 vdd p m=1 w=3.6u l=0.6u pd=8.4u ps=8.4u as=5.4p ad=5.4p
Mpnor2_pmos2 net1 B Z vdd p m=1 w=3.6u l=0.6u pd=8.4u ps=8.4u as=5.4p ad=5.4p
Mpnor2_nmos1 Z A gnd gnd n m=1 w=1.2u l=0.6u pd=3.6u ps=3.6u as=1.8p ad=1.8p
Mpnor2_nmos2 Z B gnd gnd n m=1 w=1.2u l=0.6u pd=3.6u ps=3.6u as=1.8p ad=1.8p
.ENDS pnor2_1

.SUBCKT pinv_1 A Z vdd gnd
Mpinv_pmos Z A vdd vdd p m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpinv_nmos Z A gnd gnd n m=1 w=1.2u l=0.6u pd=3.6u ps=3.6u as=1.8p ad=1.8p
.ENDS pinv_1

* ptx M{0} {1} n m=2 w=1.2u l=0.6u pd=3.6u ps=3.6u as=1.8p ad=1.8p

* ptx M{0} {1} p m=2 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p

.SUBCKT pinv_2 A Z vdd gnd
Mpinv_pmos Z A vdd vdd p m=2 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpinv_nmos Z A gnd gnd n m=2 w=1.2u l=0.6u pd=3.6u ps=3.6u as=1.8p ad=1.8p
.ENDS pinv_2

* ptx M{0} {1} n m=3 w=1.65u l=0.6u pd=4.5u ps=4.5u as=2.475p ad=2.475p

* ptx M{0} {1} p m=3 w=3.15u l=0.6u pd=7.5u ps=7.5u as=4.725p ad=4.725p

.SUBCKT pinv_3 A Z vdd gnd
Mpinv_pmos Z A vdd vdd p m=3 w=3.15u l=0.6u pd=7.5u ps=7.5u as=4.725p ad=4.725p
Mpinv_nmos Z A gnd gnd n m=3 w=1.65u l=0.6u pd=4.5u ps=4.5u as=2.475p ad=2.475p
.ENDS pinv_3

* ptx M{0} {1} n m=5 w=1.95u l=0.6u pd=5.1u ps=5.1u as=2.925p ad=2.925p

* ptx M{0} {1} p m=5 w=3.9u l=0.6u pd=9.0u ps=9.0u as=5.85p ad=5.85p

.SUBCKT pinv_4 A Z vdd gnd
Mpinv_pmos Z A vdd vdd p m=5 w=3.9u l=0.6u pd=9.0u ps=9.0u as=5.85p ad=5.85p
Mpinv_nmos Z A gnd gnd n m=5 w=1.95u l=0.6u pd=5.1u ps=5.1u as=2.925p ad=2.925p
.ENDS pinv_4

* ptx M{0} {1} n m=10 w=1.95u l=0.6u pd=5.1u ps=5.1u as=2.925p ad=2.925p

* ptx M{0} {1} p m=10 w=3.9u l=0.6u pd=9.0u ps=9.0u as=5.85p ad=5.85p

.SUBCKT pinv_5 A Z vdd gnd
Mpinv_pmos Z A vdd vdd p m=10 w=3.9u l=0.6u pd=9.0u ps=9.0u as=5.85p ad=5.85p
Mpinv_nmos Z A gnd gnd n m=10 w=1.95u l=0.6u pd=5.1u ps=5.1u as=2.925p ad=2.925p
.ENDS pinv_5
*master-slave flip-flop with both output and inverted ouput

.subckt ms_flop din dout dout_bar clk vdd gnd
xmaster din mout mout_bar clk clk_bar vdd gnd dlatch
xslave mout_bar dout_bar dout clk_bar clk_nn vdd gnd dlatch
.ends flop

.subckt dlatch din dout dout_bar clk clk_bar vdd gnd
*clk inverter
mPff1 clk_bar clk vdd vdd p W=1.8u L=0.6u m=1
mNff1 clk_bar clk gnd gnd n W=0.9u L=0.6u m=1

*transmission gate 1
mtmP1 din clk int1 vdd p W=1.8u L=0.6u m=1
mtmN1 din clk_bar int1 gnd n W=0.9u L=0.6u m=1

*foward inverter
mPff3 dout_bar int1 vdd vdd p W=1.8u L=0.6u m=1
mNff3 dout_bar int1 gnd gnd n W=0.9u L=0.6u m=1

*backward inverter
mPff4 dout dout_bar vdd vdd p W=1.8u L=0.6u m=1
mNf4 dout dout_bar gnd gnd n W=0.9u L=0.6u m=1

*transmission gate 2
mtmP2 int1 clk_bar dout vdd p W=1.8u L=0.6u m=1
mtmN2 int1 clk dout gnd n W=0.9u L=0.6u m=1
.ends dlatch


.SUBCKT msf_control din[0] din[1] din[2] dout[0] dout_bar[0] dout[1] dout_bar[1] dout[2] dout_bar[2] clk vdd gnd
XXdff0 din[0] dout[0] dout_bar[0] clk vdd gnd ms_flop
XXdff1 din[1] dout[1] dout_bar[1] clk vdd gnd ms_flop
XXdff2 din[2] dout[2] dout_bar[2] clk vdd gnd ms_flop
.ENDS msf_control

*********************** "cell_6t" ******************************
.SUBCKT replica_cell_6t bl br wl vdd gnd
M_1 gnd net_2 vdd vdd p W='0.9u' L=1.2u
M_2 net_2 gnd vdd vdd p W='0.9u' L=1.2u
M_3 br wl net_2 gnd n W='1.2u' L=0.6u
M_4 bl wl gnd gnd n W='1.2u' L=0.6u
M_5 net_2 gnd gnd gnd n W='2.4u' L=0.6u
M_6 gnd net_2 gnd gnd n W='2.4u' L=0.6u
.ENDS	$ replica_cell_6t

*********************** "cell_6t" ******************************
.SUBCKT cell_6t bl br wl vdd gnd
M_1 net_1 net_2 vdd vdd p W='0.9u' L=1.2u
M_2 net_2 net_1 vdd vdd p W='0.9u' L=1.2u
M_3 br wl net_2 gnd n W='1.2u' L=0.6u
M_4 bl wl net_1 gnd n W='1.2u' L=0.6u
M_5 net_2 net_1 gnd gnd n W='2.4u' L=0.6u
M_6 net_1 net_2 gnd gnd n W='2.4u' L=0.6u
.ENDS	$ cell_6t

.SUBCKT bitline_load bl[0] br[0] wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] vdd gnd
Xbit_r0_c0 bl[0] br[0] wl[0] vdd gnd cell_6t
Xbit_r1_c0 bl[0] br[0] wl[1] vdd gnd cell_6t
Xbit_r2_c0 bl[0] br[0] wl[2] vdd gnd cell_6t
Xbit_r3_c0 bl[0] br[0] wl[3] vdd gnd cell_6t
Xbit_r4_c0 bl[0] br[0] wl[4] vdd gnd cell_6t
Xbit_r5_c0 bl[0] br[0] wl[5] vdd gnd cell_6t
Xbit_r6_c0 bl[0] br[0] wl[6] vdd gnd cell_6t
Xbit_r7_c0 bl[0] br[0] wl[7] vdd gnd cell_6t
Xbit_r8_c0 bl[0] br[0] wl[8] vdd gnd cell_6t
Xbit_r9_c0 bl[0] br[0] wl[9] vdd gnd cell_6t
Xbit_r10_c0 bl[0] br[0] wl[10] vdd gnd cell_6t
Xbit_r11_c0 bl[0] br[0] wl[11] vdd gnd cell_6t
Xbit_r12_c0 bl[0] br[0] wl[12] vdd gnd cell_6t
Xbit_r13_c0 bl[0] br[0] wl[13] vdd gnd cell_6t
Xbit_r14_c0 bl[0] br[0] wl[14] vdd gnd cell_6t
Xbit_r15_c0 bl[0] br[0] wl[15] vdd gnd cell_6t
Xbit_r16_c0 bl[0] br[0] wl[16] vdd gnd cell_6t
Xbit_r17_c0 bl[0] br[0] wl[17] vdd gnd cell_6t
Xbit_r18_c0 bl[0] br[0] wl[18] vdd gnd cell_6t
Xbit_r19_c0 bl[0] br[0] wl[19] vdd gnd cell_6t
Xbit_r20_c0 bl[0] br[0] wl[20] vdd gnd cell_6t
Xbit_r21_c0 bl[0] br[0] wl[21] vdd gnd cell_6t
Xbit_r22_c0 bl[0] br[0] wl[22] vdd gnd cell_6t
Xbit_r23_c0 bl[0] br[0] wl[23] vdd gnd cell_6t
Xbit_r24_c0 bl[0] br[0] wl[24] vdd gnd cell_6t
Xbit_r25_c0 bl[0] br[0] wl[25] vdd gnd cell_6t
.ENDS bitline_load

.SUBCKT pinv_6 A Z vdd gnd
Mpinv_pmos Z A vdd vdd p m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpinv_nmos Z A gnd gnd n m=1 w=1.2u l=0.6u pd=3.6u ps=3.6u as=1.8p ad=1.8p
.ENDS pinv_6

.SUBCKT delay_chain in out vdd gnd
Xdinv0 in s1 vdd gnd pinv_6
Xdinv1 s1 s2n1 vdd gnd pinv_6
Xdinv2 s1 s2n2 vdd gnd pinv_6
Xdinv3 s1 s2 vdd gnd pinv_6
Xdinv4 s2 s3n1 vdd gnd pinv_6
Xdinv5 s2 s3n2 vdd gnd pinv_6
Xdinv6 s2 s3 vdd gnd pinv_6
Xdinv7 s3 s4n1 vdd gnd pinv_6
Xdinv8 s3 s4n2 vdd gnd pinv_6
Xdinv9 s3 s4 vdd gnd pinv_6
Xdinv10 s4 s5n1 vdd gnd pinv_6
Xdinv11 s4 s5n2 vdd gnd pinv_6
Xdinv12 s4 out vdd gnd pinv_6
.ENDS delay_chain

.SUBCKT pinv_7 A Z vdd gnd
Mpinv_pmos Z A vdd vdd p m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpinv_nmos Z A gnd gnd n m=1 w=1.2u l=0.6u pd=3.6u ps=3.6u as=1.8p ad=1.8p
.ENDS pinv_7

* ptx M{0} {1} p m=1 w=1.2u l=0.6u pd=3.6u ps=3.6u as=1.8p ad=1.8p

.SUBCKT replica_bitline en out vdd gnd
Xrbl_inv bl[0] out vdd gnd pinv_7
Mrbl_access_tx vdd delayed_en bl[0] vdd p m=1 w=1.2u l=0.6u pd=3.6u ps=3.6u as=1.8p ad=1.8p
Xdelay_chain en delayed_en vdd gnd delay_chain
Xbitcell bl[0] br[0] delayed_en vdd gnd replica_cell_6t
Xload bl[0] br[0] gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd vdd gnd bitline_load
.ENDS replica_bitline

.SUBCKT control_logic csb web oeb clk s_en w_en tri_en tri_en_bar clk_bar clk_buf vdd gnd
Xmsf_control oeb csb web oe_bar oe cs_bar cs we_bar we clk_buf vdd gnd msf_control
Xinv_clk1_bar clk clk1_bar vdd gnd pinv_2
Xinv_clk2 clk1_bar clk2 vdd gnd pinv_3
Xinv_clk_bar clk2 clk_bar vdd gnd pinv_4
Xinv_clk_buf clk_bar clk_buf vdd gnd pinv_5
Xnand3_rblk_bar clk_bar oe cs rblk_bar vdd gnd pnand3_1
Xinv_rblk rblk_bar rblk vdd gnd pinv_1
Xnor2_tri_en clk_buf oe_bar tri_en vdd gnd pnor2_1
Xnand2_tri_en clk_bar oe tri_en_bar vdd gnd pnand2_1
Xinv_s_en pre_s_en_bar s_en vdd gnd pinv_1
Xinv_pre_s_en_bar pre_s_en pre_s_en_bar vdd gnd pinv_1
Xnand3_w_en_bar clk_bar cs we w_en_bar vdd gnd pnand3_1
Xinv_pre_w_en w_en_bar pre_w_en vdd gnd pinv_1
Xinv_pre_w_en_bar pre_w_en pre_w_en_bar vdd gnd pinv_1
Xinv_w_en2 pre_w_en_bar w_en vdd gnd pinv_1
Xreplica_bitline rblk pre_s_en vdd gnd replica_bitline
.ENDS control_logic

.SUBCKT bitcell_array bl[0] br[0] bl[1] br[1] bl[2] br[2] bl[3] br[3] bl[4] br[4] bl[5] br[5] bl[6] br[6] bl[7] br[7] bl[8] br[8] bl[9] br[9] bl[10] br[10] bl[11] br[11] bl[12] br[12] bl[13] br[13] bl[14] br[14] bl[15] br[15] bl[16] br[16] bl[17] br[17] bl[18] br[18] bl[19] br[19] bl[20] br[20] bl[21] br[21] bl[22] br[22] bl[23] br[23] bl[24] br[24] bl[25] br[25] bl[26] br[26] bl[27] br[27] bl[28] br[28] bl[29] br[29] bl[30] br[30] bl[31] br[31] bl[32] br[32] bl[33] br[33] bl[34] br[34] bl[35] br[35] bl[36] br[36] bl[37] br[37] bl[38] br[38] bl[39] br[39] bl[40] br[40] bl[41] br[41] bl[42] br[42] bl[43] br[43] bl[44] br[44] bl[45] br[45] bl[46] br[46] bl[47] br[47] bl[48] br[48] bl[49] br[49] bl[50] br[50] bl[51] br[51] bl[52] br[52] bl[53] br[53] bl[54] br[54] bl[55] br[55] bl[56] br[56] bl[57] br[57] bl[58] br[58] bl[59] br[59] bl[60] br[60] bl[61] br[61] bl[62] br[62] bl[63] br[63] bl[64] br[64] bl[65] br[65] bl[66] br[66] bl[67] br[67] bl[68] br[68] bl[69] br[69] bl[70] br[70] bl[71] br[71] bl[72] br[72] bl[73] br[73] bl[74] br[74] bl[75] br[75] bl[76] br[76] bl[77] br[77] bl[78] br[78] bl[79] br[79] bl[80] br[80] bl[81] br[81] bl[82] br[82] bl[83] br[83] bl[84] br[84] bl[85] br[85] bl[86] br[86] bl[87] br[87] bl[88] br[88] bl[89] br[89] bl[90] br[90] bl[91] br[91] bl[92] br[92] bl[93] br[93] bl[94] br[94] bl[95] br[95] bl[96] br[96] bl[97] br[97] bl[98] br[98] bl[99] br[99] bl[100] br[100] bl[101] br[101] bl[102] br[102] bl[103] br[103] bl[104] br[104] bl[105] br[105] bl[106] br[106] bl[107] br[107] bl[108] br[108] bl[109] br[109] bl[110] br[110] bl[111] br[111] bl[112] br[112] bl[113] br[113] bl[114] br[114] bl[115] br[115] bl[116] br[116] bl[117] br[117] bl[118] br[118] bl[119] br[119] bl[120] br[120] bl[121] br[121] bl[122] br[122] bl[123] br[123] bl[124] br[124] bl[125] br[125] bl[126] br[126] bl[127] br[127] bl[128] br[128] bl[129] br[129] bl[130] br[130] bl[131] br[131] bl[132] br[132] bl[133] br[133] bl[134] br[134] bl[135] br[135] bl[136] br[136] bl[137] br[137] bl[138] br[138] bl[139] br[139] bl[140] br[140] bl[141] br[141] bl[142] br[142] bl[143] br[143] bl[144] br[144] bl[145] br[145] bl[146] br[146] bl[147] br[147] bl[148] br[148] bl[149] br[149] bl[150] br[150] bl[151] br[151] bl[152] br[152] bl[153] br[153] bl[154] br[154] bl[155] br[155] bl[156] br[156] bl[157] br[157] bl[158] br[158] bl[159] br[159] bl[160] br[160] bl[161] br[161] bl[162] br[162] bl[163] br[163] bl[164] br[164] bl[165] br[165] bl[166] br[166] bl[167] br[167] bl[168] br[168] bl[169] br[169] bl[170] br[170] bl[171] br[171] bl[172] br[172] bl[173] br[173] bl[174] br[174] bl[175] br[175] bl[176] br[176] bl[177] br[177] bl[178] br[178] bl[179] br[179] bl[180] br[180] bl[181] br[181] bl[182] br[182] bl[183] br[183] bl[184] br[184] bl[185] br[185] bl[186] br[186] bl[187] br[187] bl[188] br[188] bl[189] br[189] bl[190] br[190] bl[191] br[191] bl[192] br[192] bl[193] br[193] bl[194] br[194] bl[195] br[195] bl[196] br[196] bl[197] br[197] bl[198] br[198] bl[199] br[199] bl[200] br[200] bl[201] br[201] bl[202] br[202] bl[203] br[203] bl[204] br[204] bl[205] br[205] bl[206] br[206] bl[207] br[207] bl[208] br[208] bl[209] br[209] bl[210] br[210] bl[211] br[211] bl[212] br[212] bl[213] br[213] bl[214] br[214] bl[215] br[215] bl[216] br[216] bl[217] br[217] bl[218] br[218] bl[219] br[219] bl[220] br[220] bl[221] br[221] bl[222] br[222] bl[223] br[223] bl[224] br[224] bl[225] br[225] bl[226] br[226] bl[227] br[227] bl[228] br[228] bl[229] br[229] bl[230] br[230] bl[231] br[231] bl[232] br[232] bl[233] br[233] bl[234] br[234] bl[235] br[235] bl[236] br[236] bl[237] br[237] bl[238] br[238] bl[239] br[239] bl[240] br[240] bl[241] br[241] bl[242] br[242] bl[243] br[243] bl[244] br[244] bl[245] br[245] bl[246] br[246] bl[247] br[247] bl[248] br[248] bl[249] br[249] bl[250] br[250] bl[251] br[251] bl[252] br[252] bl[253] br[253] bl[254] br[254] bl[255] br[255] wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55] wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63] wl[64] wl[65] wl[66] wl[67] wl[68] wl[69] wl[70] wl[71] wl[72] wl[73] wl[74] wl[75] wl[76] wl[77] wl[78] wl[79] wl[80] wl[81] wl[82] wl[83] wl[84] wl[85] wl[86] wl[87] wl[88] wl[89] wl[90] wl[91] wl[92] wl[93] wl[94] wl[95] wl[96] wl[97] wl[98] wl[99] wl[100] wl[101] wl[102] wl[103] wl[104] wl[105] wl[106] wl[107] wl[108] wl[109] wl[110] wl[111] wl[112] wl[113] wl[114] wl[115] wl[116] wl[117] wl[118] wl[119] wl[120] wl[121] wl[122] wl[123] wl[124] wl[125] wl[126] wl[127] vdd gnd
Xbit_r0_c0 bl[0] br[0] wl[0] vdd gnd cell_6t
Xbit_r1_c0 bl[0] br[0] wl[1] vdd gnd cell_6t
Xbit_r2_c0 bl[0] br[0] wl[2] vdd gnd cell_6t
Xbit_r3_c0 bl[0] br[0] wl[3] vdd gnd cell_6t
Xbit_r4_c0 bl[0] br[0] wl[4] vdd gnd cell_6t
Xbit_r5_c0 bl[0] br[0] wl[5] vdd gnd cell_6t
Xbit_r6_c0 bl[0] br[0] wl[6] vdd gnd cell_6t
Xbit_r7_c0 bl[0] br[0] wl[7] vdd gnd cell_6t
Xbit_r8_c0 bl[0] br[0] wl[8] vdd gnd cell_6t
Xbit_r9_c0 bl[0] br[0] wl[9] vdd gnd cell_6t
Xbit_r10_c0 bl[0] br[0] wl[10] vdd gnd cell_6t
Xbit_r11_c0 bl[0] br[0] wl[11] vdd gnd cell_6t
Xbit_r12_c0 bl[0] br[0] wl[12] vdd gnd cell_6t
Xbit_r13_c0 bl[0] br[0] wl[13] vdd gnd cell_6t
Xbit_r14_c0 bl[0] br[0] wl[14] vdd gnd cell_6t
Xbit_r15_c0 bl[0] br[0] wl[15] vdd gnd cell_6t
Xbit_r16_c0 bl[0] br[0] wl[16] vdd gnd cell_6t
Xbit_r17_c0 bl[0] br[0] wl[17] vdd gnd cell_6t
Xbit_r18_c0 bl[0] br[0] wl[18] vdd gnd cell_6t
Xbit_r19_c0 bl[0] br[0] wl[19] vdd gnd cell_6t
Xbit_r20_c0 bl[0] br[0] wl[20] vdd gnd cell_6t
Xbit_r21_c0 bl[0] br[0] wl[21] vdd gnd cell_6t
Xbit_r22_c0 bl[0] br[0] wl[22] vdd gnd cell_6t
Xbit_r23_c0 bl[0] br[0] wl[23] vdd gnd cell_6t
Xbit_r24_c0 bl[0] br[0] wl[24] vdd gnd cell_6t
Xbit_r25_c0 bl[0] br[0] wl[25] vdd gnd cell_6t
Xbit_r26_c0 bl[0] br[0] wl[26] vdd gnd cell_6t
Xbit_r27_c0 bl[0] br[0] wl[27] vdd gnd cell_6t
Xbit_r28_c0 bl[0] br[0] wl[28] vdd gnd cell_6t
Xbit_r29_c0 bl[0] br[0] wl[29] vdd gnd cell_6t
Xbit_r30_c0 bl[0] br[0] wl[30] vdd gnd cell_6t
Xbit_r31_c0 bl[0] br[0] wl[31] vdd gnd cell_6t
Xbit_r32_c0 bl[0] br[0] wl[32] vdd gnd cell_6t
Xbit_r33_c0 bl[0] br[0] wl[33] vdd gnd cell_6t
Xbit_r34_c0 bl[0] br[0] wl[34] vdd gnd cell_6t
Xbit_r35_c0 bl[0] br[0] wl[35] vdd gnd cell_6t
Xbit_r36_c0 bl[0] br[0] wl[36] vdd gnd cell_6t
Xbit_r37_c0 bl[0] br[0] wl[37] vdd gnd cell_6t
Xbit_r38_c0 bl[0] br[0] wl[38] vdd gnd cell_6t
Xbit_r39_c0 bl[0] br[0] wl[39] vdd gnd cell_6t
Xbit_r40_c0 bl[0] br[0] wl[40] vdd gnd cell_6t
Xbit_r41_c0 bl[0] br[0] wl[41] vdd gnd cell_6t
Xbit_r42_c0 bl[0] br[0] wl[42] vdd gnd cell_6t
Xbit_r43_c0 bl[0] br[0] wl[43] vdd gnd cell_6t
Xbit_r44_c0 bl[0] br[0] wl[44] vdd gnd cell_6t
Xbit_r45_c0 bl[0] br[0] wl[45] vdd gnd cell_6t
Xbit_r46_c0 bl[0] br[0] wl[46] vdd gnd cell_6t
Xbit_r47_c0 bl[0] br[0] wl[47] vdd gnd cell_6t
Xbit_r48_c0 bl[0] br[0] wl[48] vdd gnd cell_6t
Xbit_r49_c0 bl[0] br[0] wl[49] vdd gnd cell_6t
Xbit_r50_c0 bl[0] br[0] wl[50] vdd gnd cell_6t
Xbit_r51_c0 bl[0] br[0] wl[51] vdd gnd cell_6t
Xbit_r52_c0 bl[0] br[0] wl[52] vdd gnd cell_6t
Xbit_r53_c0 bl[0] br[0] wl[53] vdd gnd cell_6t
Xbit_r54_c0 bl[0] br[0] wl[54] vdd gnd cell_6t
Xbit_r55_c0 bl[0] br[0] wl[55] vdd gnd cell_6t
Xbit_r56_c0 bl[0] br[0] wl[56] vdd gnd cell_6t
Xbit_r57_c0 bl[0] br[0] wl[57] vdd gnd cell_6t
Xbit_r58_c0 bl[0] br[0] wl[58] vdd gnd cell_6t
Xbit_r59_c0 bl[0] br[0] wl[59] vdd gnd cell_6t
Xbit_r60_c0 bl[0] br[0] wl[60] vdd gnd cell_6t
Xbit_r61_c0 bl[0] br[0] wl[61] vdd gnd cell_6t
Xbit_r62_c0 bl[0] br[0] wl[62] vdd gnd cell_6t
Xbit_r63_c0 bl[0] br[0] wl[63] vdd gnd cell_6t
Xbit_r64_c0 bl[0] br[0] wl[64] vdd gnd cell_6t
Xbit_r65_c0 bl[0] br[0] wl[65] vdd gnd cell_6t
Xbit_r66_c0 bl[0] br[0] wl[66] vdd gnd cell_6t
Xbit_r67_c0 bl[0] br[0] wl[67] vdd gnd cell_6t
Xbit_r68_c0 bl[0] br[0] wl[68] vdd gnd cell_6t
Xbit_r69_c0 bl[0] br[0] wl[69] vdd gnd cell_6t
Xbit_r70_c0 bl[0] br[0] wl[70] vdd gnd cell_6t
Xbit_r71_c0 bl[0] br[0] wl[71] vdd gnd cell_6t
Xbit_r72_c0 bl[0] br[0] wl[72] vdd gnd cell_6t
Xbit_r73_c0 bl[0] br[0] wl[73] vdd gnd cell_6t
Xbit_r74_c0 bl[0] br[0] wl[74] vdd gnd cell_6t
Xbit_r75_c0 bl[0] br[0] wl[75] vdd gnd cell_6t
Xbit_r76_c0 bl[0] br[0] wl[76] vdd gnd cell_6t
Xbit_r77_c0 bl[0] br[0] wl[77] vdd gnd cell_6t
Xbit_r78_c0 bl[0] br[0] wl[78] vdd gnd cell_6t
Xbit_r79_c0 bl[0] br[0] wl[79] vdd gnd cell_6t
Xbit_r80_c0 bl[0] br[0] wl[80] vdd gnd cell_6t
Xbit_r81_c0 bl[0] br[0] wl[81] vdd gnd cell_6t
Xbit_r82_c0 bl[0] br[0] wl[82] vdd gnd cell_6t
Xbit_r83_c0 bl[0] br[0] wl[83] vdd gnd cell_6t
Xbit_r84_c0 bl[0] br[0] wl[84] vdd gnd cell_6t
Xbit_r85_c0 bl[0] br[0] wl[85] vdd gnd cell_6t
Xbit_r86_c0 bl[0] br[0] wl[86] vdd gnd cell_6t
Xbit_r87_c0 bl[0] br[0] wl[87] vdd gnd cell_6t
Xbit_r88_c0 bl[0] br[0] wl[88] vdd gnd cell_6t
Xbit_r89_c0 bl[0] br[0] wl[89] vdd gnd cell_6t
Xbit_r90_c0 bl[0] br[0] wl[90] vdd gnd cell_6t
Xbit_r91_c0 bl[0] br[0] wl[91] vdd gnd cell_6t
Xbit_r92_c0 bl[0] br[0] wl[92] vdd gnd cell_6t
Xbit_r93_c0 bl[0] br[0] wl[93] vdd gnd cell_6t
Xbit_r94_c0 bl[0] br[0] wl[94] vdd gnd cell_6t
Xbit_r95_c0 bl[0] br[0] wl[95] vdd gnd cell_6t
Xbit_r96_c0 bl[0] br[0] wl[96] vdd gnd cell_6t
Xbit_r97_c0 bl[0] br[0] wl[97] vdd gnd cell_6t
Xbit_r98_c0 bl[0] br[0] wl[98] vdd gnd cell_6t
Xbit_r99_c0 bl[0] br[0] wl[99] vdd gnd cell_6t
Xbit_r100_c0 bl[0] br[0] wl[100] vdd gnd cell_6t
Xbit_r101_c0 bl[0] br[0] wl[101] vdd gnd cell_6t
Xbit_r102_c0 bl[0] br[0] wl[102] vdd gnd cell_6t
Xbit_r103_c0 bl[0] br[0] wl[103] vdd gnd cell_6t
Xbit_r104_c0 bl[0] br[0] wl[104] vdd gnd cell_6t
Xbit_r105_c0 bl[0] br[0] wl[105] vdd gnd cell_6t
Xbit_r106_c0 bl[0] br[0] wl[106] vdd gnd cell_6t
Xbit_r107_c0 bl[0] br[0] wl[107] vdd gnd cell_6t
Xbit_r108_c0 bl[0] br[0] wl[108] vdd gnd cell_6t
Xbit_r109_c0 bl[0] br[0] wl[109] vdd gnd cell_6t
Xbit_r110_c0 bl[0] br[0] wl[110] vdd gnd cell_6t
Xbit_r111_c0 bl[0] br[0] wl[111] vdd gnd cell_6t
Xbit_r112_c0 bl[0] br[0] wl[112] vdd gnd cell_6t
Xbit_r113_c0 bl[0] br[0] wl[113] vdd gnd cell_6t
Xbit_r114_c0 bl[0] br[0] wl[114] vdd gnd cell_6t
Xbit_r115_c0 bl[0] br[0] wl[115] vdd gnd cell_6t
Xbit_r116_c0 bl[0] br[0] wl[116] vdd gnd cell_6t
Xbit_r117_c0 bl[0] br[0] wl[117] vdd gnd cell_6t
Xbit_r118_c0 bl[0] br[0] wl[118] vdd gnd cell_6t
Xbit_r119_c0 bl[0] br[0] wl[119] vdd gnd cell_6t
Xbit_r120_c0 bl[0] br[0] wl[120] vdd gnd cell_6t
Xbit_r121_c0 bl[0] br[0] wl[121] vdd gnd cell_6t
Xbit_r122_c0 bl[0] br[0] wl[122] vdd gnd cell_6t
Xbit_r123_c0 bl[0] br[0] wl[123] vdd gnd cell_6t
Xbit_r124_c0 bl[0] br[0] wl[124] vdd gnd cell_6t
Xbit_r125_c0 bl[0] br[0] wl[125] vdd gnd cell_6t
Xbit_r126_c0 bl[0] br[0] wl[126] vdd gnd cell_6t
Xbit_r127_c0 bl[0] br[0] wl[127] vdd gnd cell_6t
Xbit_r0_c1 bl[1] br[1] wl[0] vdd gnd cell_6t
Xbit_r1_c1 bl[1] br[1] wl[1] vdd gnd cell_6t
Xbit_r2_c1 bl[1] br[1] wl[2] vdd gnd cell_6t
Xbit_r3_c1 bl[1] br[1] wl[3] vdd gnd cell_6t
Xbit_r4_c1 bl[1] br[1] wl[4] vdd gnd cell_6t
Xbit_r5_c1 bl[1] br[1] wl[5] vdd gnd cell_6t
Xbit_r6_c1 bl[1] br[1] wl[6] vdd gnd cell_6t
Xbit_r7_c1 bl[1] br[1] wl[7] vdd gnd cell_6t
Xbit_r8_c1 bl[1] br[1] wl[8] vdd gnd cell_6t
Xbit_r9_c1 bl[1] br[1] wl[9] vdd gnd cell_6t
Xbit_r10_c1 bl[1] br[1] wl[10] vdd gnd cell_6t
Xbit_r11_c1 bl[1] br[1] wl[11] vdd gnd cell_6t
Xbit_r12_c1 bl[1] br[1] wl[12] vdd gnd cell_6t
Xbit_r13_c1 bl[1] br[1] wl[13] vdd gnd cell_6t
Xbit_r14_c1 bl[1] br[1] wl[14] vdd gnd cell_6t
Xbit_r15_c1 bl[1] br[1] wl[15] vdd gnd cell_6t
Xbit_r16_c1 bl[1] br[1] wl[16] vdd gnd cell_6t
Xbit_r17_c1 bl[1] br[1] wl[17] vdd gnd cell_6t
Xbit_r18_c1 bl[1] br[1] wl[18] vdd gnd cell_6t
Xbit_r19_c1 bl[1] br[1] wl[19] vdd gnd cell_6t
Xbit_r20_c1 bl[1] br[1] wl[20] vdd gnd cell_6t
Xbit_r21_c1 bl[1] br[1] wl[21] vdd gnd cell_6t
Xbit_r22_c1 bl[1] br[1] wl[22] vdd gnd cell_6t
Xbit_r23_c1 bl[1] br[1] wl[23] vdd gnd cell_6t
Xbit_r24_c1 bl[1] br[1] wl[24] vdd gnd cell_6t
Xbit_r25_c1 bl[1] br[1] wl[25] vdd gnd cell_6t
Xbit_r26_c1 bl[1] br[1] wl[26] vdd gnd cell_6t
Xbit_r27_c1 bl[1] br[1] wl[27] vdd gnd cell_6t
Xbit_r28_c1 bl[1] br[1] wl[28] vdd gnd cell_6t
Xbit_r29_c1 bl[1] br[1] wl[29] vdd gnd cell_6t
Xbit_r30_c1 bl[1] br[1] wl[30] vdd gnd cell_6t
Xbit_r31_c1 bl[1] br[1] wl[31] vdd gnd cell_6t
Xbit_r32_c1 bl[1] br[1] wl[32] vdd gnd cell_6t
Xbit_r33_c1 bl[1] br[1] wl[33] vdd gnd cell_6t
Xbit_r34_c1 bl[1] br[1] wl[34] vdd gnd cell_6t
Xbit_r35_c1 bl[1] br[1] wl[35] vdd gnd cell_6t
Xbit_r36_c1 bl[1] br[1] wl[36] vdd gnd cell_6t
Xbit_r37_c1 bl[1] br[1] wl[37] vdd gnd cell_6t
Xbit_r38_c1 bl[1] br[1] wl[38] vdd gnd cell_6t
Xbit_r39_c1 bl[1] br[1] wl[39] vdd gnd cell_6t
Xbit_r40_c1 bl[1] br[1] wl[40] vdd gnd cell_6t
Xbit_r41_c1 bl[1] br[1] wl[41] vdd gnd cell_6t
Xbit_r42_c1 bl[1] br[1] wl[42] vdd gnd cell_6t
Xbit_r43_c1 bl[1] br[1] wl[43] vdd gnd cell_6t
Xbit_r44_c1 bl[1] br[1] wl[44] vdd gnd cell_6t
Xbit_r45_c1 bl[1] br[1] wl[45] vdd gnd cell_6t
Xbit_r46_c1 bl[1] br[1] wl[46] vdd gnd cell_6t
Xbit_r47_c1 bl[1] br[1] wl[47] vdd gnd cell_6t
Xbit_r48_c1 bl[1] br[1] wl[48] vdd gnd cell_6t
Xbit_r49_c1 bl[1] br[1] wl[49] vdd gnd cell_6t
Xbit_r50_c1 bl[1] br[1] wl[50] vdd gnd cell_6t
Xbit_r51_c1 bl[1] br[1] wl[51] vdd gnd cell_6t
Xbit_r52_c1 bl[1] br[1] wl[52] vdd gnd cell_6t
Xbit_r53_c1 bl[1] br[1] wl[53] vdd gnd cell_6t
Xbit_r54_c1 bl[1] br[1] wl[54] vdd gnd cell_6t
Xbit_r55_c1 bl[1] br[1] wl[55] vdd gnd cell_6t
Xbit_r56_c1 bl[1] br[1] wl[56] vdd gnd cell_6t
Xbit_r57_c1 bl[1] br[1] wl[57] vdd gnd cell_6t
Xbit_r58_c1 bl[1] br[1] wl[58] vdd gnd cell_6t
Xbit_r59_c1 bl[1] br[1] wl[59] vdd gnd cell_6t
Xbit_r60_c1 bl[1] br[1] wl[60] vdd gnd cell_6t
Xbit_r61_c1 bl[1] br[1] wl[61] vdd gnd cell_6t
Xbit_r62_c1 bl[1] br[1] wl[62] vdd gnd cell_6t
Xbit_r63_c1 bl[1] br[1] wl[63] vdd gnd cell_6t
Xbit_r64_c1 bl[1] br[1] wl[64] vdd gnd cell_6t
Xbit_r65_c1 bl[1] br[1] wl[65] vdd gnd cell_6t
Xbit_r66_c1 bl[1] br[1] wl[66] vdd gnd cell_6t
Xbit_r67_c1 bl[1] br[1] wl[67] vdd gnd cell_6t
Xbit_r68_c1 bl[1] br[1] wl[68] vdd gnd cell_6t
Xbit_r69_c1 bl[1] br[1] wl[69] vdd gnd cell_6t
Xbit_r70_c1 bl[1] br[1] wl[70] vdd gnd cell_6t
Xbit_r71_c1 bl[1] br[1] wl[71] vdd gnd cell_6t
Xbit_r72_c1 bl[1] br[1] wl[72] vdd gnd cell_6t
Xbit_r73_c1 bl[1] br[1] wl[73] vdd gnd cell_6t
Xbit_r74_c1 bl[1] br[1] wl[74] vdd gnd cell_6t
Xbit_r75_c1 bl[1] br[1] wl[75] vdd gnd cell_6t
Xbit_r76_c1 bl[1] br[1] wl[76] vdd gnd cell_6t
Xbit_r77_c1 bl[1] br[1] wl[77] vdd gnd cell_6t
Xbit_r78_c1 bl[1] br[1] wl[78] vdd gnd cell_6t
Xbit_r79_c1 bl[1] br[1] wl[79] vdd gnd cell_6t
Xbit_r80_c1 bl[1] br[1] wl[80] vdd gnd cell_6t
Xbit_r81_c1 bl[1] br[1] wl[81] vdd gnd cell_6t
Xbit_r82_c1 bl[1] br[1] wl[82] vdd gnd cell_6t
Xbit_r83_c1 bl[1] br[1] wl[83] vdd gnd cell_6t
Xbit_r84_c1 bl[1] br[1] wl[84] vdd gnd cell_6t
Xbit_r85_c1 bl[1] br[1] wl[85] vdd gnd cell_6t
Xbit_r86_c1 bl[1] br[1] wl[86] vdd gnd cell_6t
Xbit_r87_c1 bl[1] br[1] wl[87] vdd gnd cell_6t
Xbit_r88_c1 bl[1] br[1] wl[88] vdd gnd cell_6t
Xbit_r89_c1 bl[1] br[1] wl[89] vdd gnd cell_6t
Xbit_r90_c1 bl[1] br[1] wl[90] vdd gnd cell_6t
Xbit_r91_c1 bl[1] br[1] wl[91] vdd gnd cell_6t
Xbit_r92_c1 bl[1] br[1] wl[92] vdd gnd cell_6t
Xbit_r93_c1 bl[1] br[1] wl[93] vdd gnd cell_6t
Xbit_r94_c1 bl[1] br[1] wl[94] vdd gnd cell_6t
Xbit_r95_c1 bl[1] br[1] wl[95] vdd gnd cell_6t
Xbit_r96_c1 bl[1] br[1] wl[96] vdd gnd cell_6t
Xbit_r97_c1 bl[1] br[1] wl[97] vdd gnd cell_6t
Xbit_r98_c1 bl[1] br[1] wl[98] vdd gnd cell_6t
Xbit_r99_c1 bl[1] br[1] wl[99] vdd gnd cell_6t
Xbit_r100_c1 bl[1] br[1] wl[100] vdd gnd cell_6t
Xbit_r101_c1 bl[1] br[1] wl[101] vdd gnd cell_6t
Xbit_r102_c1 bl[1] br[1] wl[102] vdd gnd cell_6t
Xbit_r103_c1 bl[1] br[1] wl[103] vdd gnd cell_6t
Xbit_r104_c1 bl[1] br[1] wl[104] vdd gnd cell_6t
Xbit_r105_c1 bl[1] br[1] wl[105] vdd gnd cell_6t
Xbit_r106_c1 bl[1] br[1] wl[106] vdd gnd cell_6t
Xbit_r107_c1 bl[1] br[1] wl[107] vdd gnd cell_6t
Xbit_r108_c1 bl[1] br[1] wl[108] vdd gnd cell_6t
Xbit_r109_c1 bl[1] br[1] wl[109] vdd gnd cell_6t
Xbit_r110_c1 bl[1] br[1] wl[110] vdd gnd cell_6t
Xbit_r111_c1 bl[1] br[1] wl[111] vdd gnd cell_6t
Xbit_r112_c1 bl[1] br[1] wl[112] vdd gnd cell_6t
Xbit_r113_c1 bl[1] br[1] wl[113] vdd gnd cell_6t
Xbit_r114_c1 bl[1] br[1] wl[114] vdd gnd cell_6t
Xbit_r115_c1 bl[1] br[1] wl[115] vdd gnd cell_6t
Xbit_r116_c1 bl[1] br[1] wl[116] vdd gnd cell_6t
Xbit_r117_c1 bl[1] br[1] wl[117] vdd gnd cell_6t
Xbit_r118_c1 bl[1] br[1] wl[118] vdd gnd cell_6t
Xbit_r119_c1 bl[1] br[1] wl[119] vdd gnd cell_6t
Xbit_r120_c1 bl[1] br[1] wl[120] vdd gnd cell_6t
Xbit_r121_c1 bl[1] br[1] wl[121] vdd gnd cell_6t
Xbit_r122_c1 bl[1] br[1] wl[122] vdd gnd cell_6t
Xbit_r123_c1 bl[1] br[1] wl[123] vdd gnd cell_6t
Xbit_r124_c1 bl[1] br[1] wl[124] vdd gnd cell_6t
Xbit_r125_c1 bl[1] br[1] wl[125] vdd gnd cell_6t
Xbit_r126_c1 bl[1] br[1] wl[126] vdd gnd cell_6t
Xbit_r127_c1 bl[1] br[1] wl[127] vdd gnd cell_6t
Xbit_r0_c2 bl[2] br[2] wl[0] vdd gnd cell_6t
Xbit_r1_c2 bl[2] br[2] wl[1] vdd gnd cell_6t
Xbit_r2_c2 bl[2] br[2] wl[2] vdd gnd cell_6t
Xbit_r3_c2 bl[2] br[2] wl[3] vdd gnd cell_6t
Xbit_r4_c2 bl[2] br[2] wl[4] vdd gnd cell_6t
Xbit_r5_c2 bl[2] br[2] wl[5] vdd gnd cell_6t
Xbit_r6_c2 bl[2] br[2] wl[6] vdd gnd cell_6t
Xbit_r7_c2 bl[2] br[2] wl[7] vdd gnd cell_6t
Xbit_r8_c2 bl[2] br[2] wl[8] vdd gnd cell_6t
Xbit_r9_c2 bl[2] br[2] wl[9] vdd gnd cell_6t
Xbit_r10_c2 bl[2] br[2] wl[10] vdd gnd cell_6t
Xbit_r11_c2 bl[2] br[2] wl[11] vdd gnd cell_6t
Xbit_r12_c2 bl[2] br[2] wl[12] vdd gnd cell_6t
Xbit_r13_c2 bl[2] br[2] wl[13] vdd gnd cell_6t
Xbit_r14_c2 bl[2] br[2] wl[14] vdd gnd cell_6t
Xbit_r15_c2 bl[2] br[2] wl[15] vdd gnd cell_6t
Xbit_r16_c2 bl[2] br[2] wl[16] vdd gnd cell_6t
Xbit_r17_c2 bl[2] br[2] wl[17] vdd gnd cell_6t
Xbit_r18_c2 bl[2] br[2] wl[18] vdd gnd cell_6t
Xbit_r19_c2 bl[2] br[2] wl[19] vdd gnd cell_6t
Xbit_r20_c2 bl[2] br[2] wl[20] vdd gnd cell_6t
Xbit_r21_c2 bl[2] br[2] wl[21] vdd gnd cell_6t
Xbit_r22_c2 bl[2] br[2] wl[22] vdd gnd cell_6t
Xbit_r23_c2 bl[2] br[2] wl[23] vdd gnd cell_6t
Xbit_r24_c2 bl[2] br[2] wl[24] vdd gnd cell_6t
Xbit_r25_c2 bl[2] br[2] wl[25] vdd gnd cell_6t
Xbit_r26_c2 bl[2] br[2] wl[26] vdd gnd cell_6t
Xbit_r27_c2 bl[2] br[2] wl[27] vdd gnd cell_6t
Xbit_r28_c2 bl[2] br[2] wl[28] vdd gnd cell_6t
Xbit_r29_c2 bl[2] br[2] wl[29] vdd gnd cell_6t
Xbit_r30_c2 bl[2] br[2] wl[30] vdd gnd cell_6t
Xbit_r31_c2 bl[2] br[2] wl[31] vdd gnd cell_6t
Xbit_r32_c2 bl[2] br[2] wl[32] vdd gnd cell_6t
Xbit_r33_c2 bl[2] br[2] wl[33] vdd gnd cell_6t
Xbit_r34_c2 bl[2] br[2] wl[34] vdd gnd cell_6t
Xbit_r35_c2 bl[2] br[2] wl[35] vdd gnd cell_6t
Xbit_r36_c2 bl[2] br[2] wl[36] vdd gnd cell_6t
Xbit_r37_c2 bl[2] br[2] wl[37] vdd gnd cell_6t
Xbit_r38_c2 bl[2] br[2] wl[38] vdd gnd cell_6t
Xbit_r39_c2 bl[2] br[2] wl[39] vdd gnd cell_6t
Xbit_r40_c2 bl[2] br[2] wl[40] vdd gnd cell_6t
Xbit_r41_c2 bl[2] br[2] wl[41] vdd gnd cell_6t
Xbit_r42_c2 bl[2] br[2] wl[42] vdd gnd cell_6t
Xbit_r43_c2 bl[2] br[2] wl[43] vdd gnd cell_6t
Xbit_r44_c2 bl[2] br[2] wl[44] vdd gnd cell_6t
Xbit_r45_c2 bl[2] br[2] wl[45] vdd gnd cell_6t
Xbit_r46_c2 bl[2] br[2] wl[46] vdd gnd cell_6t
Xbit_r47_c2 bl[2] br[2] wl[47] vdd gnd cell_6t
Xbit_r48_c2 bl[2] br[2] wl[48] vdd gnd cell_6t
Xbit_r49_c2 bl[2] br[2] wl[49] vdd gnd cell_6t
Xbit_r50_c2 bl[2] br[2] wl[50] vdd gnd cell_6t
Xbit_r51_c2 bl[2] br[2] wl[51] vdd gnd cell_6t
Xbit_r52_c2 bl[2] br[2] wl[52] vdd gnd cell_6t
Xbit_r53_c2 bl[2] br[2] wl[53] vdd gnd cell_6t
Xbit_r54_c2 bl[2] br[2] wl[54] vdd gnd cell_6t
Xbit_r55_c2 bl[2] br[2] wl[55] vdd gnd cell_6t
Xbit_r56_c2 bl[2] br[2] wl[56] vdd gnd cell_6t
Xbit_r57_c2 bl[2] br[2] wl[57] vdd gnd cell_6t
Xbit_r58_c2 bl[2] br[2] wl[58] vdd gnd cell_6t
Xbit_r59_c2 bl[2] br[2] wl[59] vdd gnd cell_6t
Xbit_r60_c2 bl[2] br[2] wl[60] vdd gnd cell_6t
Xbit_r61_c2 bl[2] br[2] wl[61] vdd gnd cell_6t
Xbit_r62_c2 bl[2] br[2] wl[62] vdd gnd cell_6t
Xbit_r63_c2 bl[2] br[2] wl[63] vdd gnd cell_6t
Xbit_r64_c2 bl[2] br[2] wl[64] vdd gnd cell_6t
Xbit_r65_c2 bl[2] br[2] wl[65] vdd gnd cell_6t
Xbit_r66_c2 bl[2] br[2] wl[66] vdd gnd cell_6t
Xbit_r67_c2 bl[2] br[2] wl[67] vdd gnd cell_6t
Xbit_r68_c2 bl[2] br[2] wl[68] vdd gnd cell_6t
Xbit_r69_c2 bl[2] br[2] wl[69] vdd gnd cell_6t
Xbit_r70_c2 bl[2] br[2] wl[70] vdd gnd cell_6t
Xbit_r71_c2 bl[2] br[2] wl[71] vdd gnd cell_6t
Xbit_r72_c2 bl[2] br[2] wl[72] vdd gnd cell_6t
Xbit_r73_c2 bl[2] br[2] wl[73] vdd gnd cell_6t
Xbit_r74_c2 bl[2] br[2] wl[74] vdd gnd cell_6t
Xbit_r75_c2 bl[2] br[2] wl[75] vdd gnd cell_6t
Xbit_r76_c2 bl[2] br[2] wl[76] vdd gnd cell_6t
Xbit_r77_c2 bl[2] br[2] wl[77] vdd gnd cell_6t
Xbit_r78_c2 bl[2] br[2] wl[78] vdd gnd cell_6t
Xbit_r79_c2 bl[2] br[2] wl[79] vdd gnd cell_6t
Xbit_r80_c2 bl[2] br[2] wl[80] vdd gnd cell_6t
Xbit_r81_c2 bl[2] br[2] wl[81] vdd gnd cell_6t
Xbit_r82_c2 bl[2] br[2] wl[82] vdd gnd cell_6t
Xbit_r83_c2 bl[2] br[2] wl[83] vdd gnd cell_6t
Xbit_r84_c2 bl[2] br[2] wl[84] vdd gnd cell_6t
Xbit_r85_c2 bl[2] br[2] wl[85] vdd gnd cell_6t
Xbit_r86_c2 bl[2] br[2] wl[86] vdd gnd cell_6t
Xbit_r87_c2 bl[2] br[2] wl[87] vdd gnd cell_6t
Xbit_r88_c2 bl[2] br[2] wl[88] vdd gnd cell_6t
Xbit_r89_c2 bl[2] br[2] wl[89] vdd gnd cell_6t
Xbit_r90_c2 bl[2] br[2] wl[90] vdd gnd cell_6t
Xbit_r91_c2 bl[2] br[2] wl[91] vdd gnd cell_6t
Xbit_r92_c2 bl[2] br[2] wl[92] vdd gnd cell_6t
Xbit_r93_c2 bl[2] br[2] wl[93] vdd gnd cell_6t
Xbit_r94_c2 bl[2] br[2] wl[94] vdd gnd cell_6t
Xbit_r95_c2 bl[2] br[2] wl[95] vdd gnd cell_6t
Xbit_r96_c2 bl[2] br[2] wl[96] vdd gnd cell_6t
Xbit_r97_c2 bl[2] br[2] wl[97] vdd gnd cell_6t
Xbit_r98_c2 bl[2] br[2] wl[98] vdd gnd cell_6t
Xbit_r99_c2 bl[2] br[2] wl[99] vdd gnd cell_6t
Xbit_r100_c2 bl[2] br[2] wl[100] vdd gnd cell_6t
Xbit_r101_c2 bl[2] br[2] wl[101] vdd gnd cell_6t
Xbit_r102_c2 bl[2] br[2] wl[102] vdd gnd cell_6t
Xbit_r103_c2 bl[2] br[2] wl[103] vdd gnd cell_6t
Xbit_r104_c2 bl[2] br[2] wl[104] vdd gnd cell_6t
Xbit_r105_c2 bl[2] br[2] wl[105] vdd gnd cell_6t
Xbit_r106_c2 bl[2] br[2] wl[106] vdd gnd cell_6t
Xbit_r107_c2 bl[2] br[2] wl[107] vdd gnd cell_6t
Xbit_r108_c2 bl[2] br[2] wl[108] vdd gnd cell_6t
Xbit_r109_c2 bl[2] br[2] wl[109] vdd gnd cell_6t
Xbit_r110_c2 bl[2] br[2] wl[110] vdd gnd cell_6t
Xbit_r111_c2 bl[2] br[2] wl[111] vdd gnd cell_6t
Xbit_r112_c2 bl[2] br[2] wl[112] vdd gnd cell_6t
Xbit_r113_c2 bl[2] br[2] wl[113] vdd gnd cell_6t
Xbit_r114_c2 bl[2] br[2] wl[114] vdd gnd cell_6t
Xbit_r115_c2 bl[2] br[2] wl[115] vdd gnd cell_6t
Xbit_r116_c2 bl[2] br[2] wl[116] vdd gnd cell_6t
Xbit_r117_c2 bl[2] br[2] wl[117] vdd gnd cell_6t
Xbit_r118_c2 bl[2] br[2] wl[118] vdd gnd cell_6t
Xbit_r119_c2 bl[2] br[2] wl[119] vdd gnd cell_6t
Xbit_r120_c2 bl[2] br[2] wl[120] vdd gnd cell_6t
Xbit_r121_c2 bl[2] br[2] wl[121] vdd gnd cell_6t
Xbit_r122_c2 bl[2] br[2] wl[122] vdd gnd cell_6t
Xbit_r123_c2 bl[2] br[2] wl[123] vdd gnd cell_6t
Xbit_r124_c2 bl[2] br[2] wl[124] vdd gnd cell_6t
Xbit_r125_c2 bl[2] br[2] wl[125] vdd gnd cell_6t
Xbit_r126_c2 bl[2] br[2] wl[126] vdd gnd cell_6t
Xbit_r127_c2 bl[2] br[2] wl[127] vdd gnd cell_6t
Xbit_r0_c3 bl[3] br[3] wl[0] vdd gnd cell_6t
Xbit_r1_c3 bl[3] br[3] wl[1] vdd gnd cell_6t
Xbit_r2_c3 bl[3] br[3] wl[2] vdd gnd cell_6t
Xbit_r3_c3 bl[3] br[3] wl[3] vdd gnd cell_6t
Xbit_r4_c3 bl[3] br[3] wl[4] vdd gnd cell_6t
Xbit_r5_c3 bl[3] br[3] wl[5] vdd gnd cell_6t
Xbit_r6_c3 bl[3] br[3] wl[6] vdd gnd cell_6t
Xbit_r7_c3 bl[3] br[3] wl[7] vdd gnd cell_6t
Xbit_r8_c3 bl[3] br[3] wl[8] vdd gnd cell_6t
Xbit_r9_c3 bl[3] br[3] wl[9] vdd gnd cell_6t
Xbit_r10_c3 bl[3] br[3] wl[10] vdd gnd cell_6t
Xbit_r11_c3 bl[3] br[3] wl[11] vdd gnd cell_6t
Xbit_r12_c3 bl[3] br[3] wl[12] vdd gnd cell_6t
Xbit_r13_c3 bl[3] br[3] wl[13] vdd gnd cell_6t
Xbit_r14_c3 bl[3] br[3] wl[14] vdd gnd cell_6t
Xbit_r15_c3 bl[3] br[3] wl[15] vdd gnd cell_6t
Xbit_r16_c3 bl[3] br[3] wl[16] vdd gnd cell_6t
Xbit_r17_c3 bl[3] br[3] wl[17] vdd gnd cell_6t
Xbit_r18_c3 bl[3] br[3] wl[18] vdd gnd cell_6t
Xbit_r19_c3 bl[3] br[3] wl[19] vdd gnd cell_6t
Xbit_r20_c3 bl[3] br[3] wl[20] vdd gnd cell_6t
Xbit_r21_c3 bl[3] br[3] wl[21] vdd gnd cell_6t
Xbit_r22_c3 bl[3] br[3] wl[22] vdd gnd cell_6t
Xbit_r23_c3 bl[3] br[3] wl[23] vdd gnd cell_6t
Xbit_r24_c3 bl[3] br[3] wl[24] vdd gnd cell_6t
Xbit_r25_c3 bl[3] br[3] wl[25] vdd gnd cell_6t
Xbit_r26_c3 bl[3] br[3] wl[26] vdd gnd cell_6t
Xbit_r27_c3 bl[3] br[3] wl[27] vdd gnd cell_6t
Xbit_r28_c3 bl[3] br[3] wl[28] vdd gnd cell_6t
Xbit_r29_c3 bl[3] br[3] wl[29] vdd gnd cell_6t
Xbit_r30_c3 bl[3] br[3] wl[30] vdd gnd cell_6t
Xbit_r31_c3 bl[3] br[3] wl[31] vdd gnd cell_6t
Xbit_r32_c3 bl[3] br[3] wl[32] vdd gnd cell_6t
Xbit_r33_c3 bl[3] br[3] wl[33] vdd gnd cell_6t
Xbit_r34_c3 bl[3] br[3] wl[34] vdd gnd cell_6t
Xbit_r35_c3 bl[3] br[3] wl[35] vdd gnd cell_6t
Xbit_r36_c3 bl[3] br[3] wl[36] vdd gnd cell_6t
Xbit_r37_c3 bl[3] br[3] wl[37] vdd gnd cell_6t
Xbit_r38_c3 bl[3] br[3] wl[38] vdd gnd cell_6t
Xbit_r39_c3 bl[3] br[3] wl[39] vdd gnd cell_6t
Xbit_r40_c3 bl[3] br[3] wl[40] vdd gnd cell_6t
Xbit_r41_c3 bl[3] br[3] wl[41] vdd gnd cell_6t
Xbit_r42_c3 bl[3] br[3] wl[42] vdd gnd cell_6t
Xbit_r43_c3 bl[3] br[3] wl[43] vdd gnd cell_6t
Xbit_r44_c3 bl[3] br[3] wl[44] vdd gnd cell_6t
Xbit_r45_c3 bl[3] br[3] wl[45] vdd gnd cell_6t
Xbit_r46_c3 bl[3] br[3] wl[46] vdd gnd cell_6t
Xbit_r47_c3 bl[3] br[3] wl[47] vdd gnd cell_6t
Xbit_r48_c3 bl[3] br[3] wl[48] vdd gnd cell_6t
Xbit_r49_c3 bl[3] br[3] wl[49] vdd gnd cell_6t
Xbit_r50_c3 bl[3] br[3] wl[50] vdd gnd cell_6t
Xbit_r51_c3 bl[3] br[3] wl[51] vdd gnd cell_6t
Xbit_r52_c3 bl[3] br[3] wl[52] vdd gnd cell_6t
Xbit_r53_c3 bl[3] br[3] wl[53] vdd gnd cell_6t
Xbit_r54_c3 bl[3] br[3] wl[54] vdd gnd cell_6t
Xbit_r55_c3 bl[3] br[3] wl[55] vdd gnd cell_6t
Xbit_r56_c3 bl[3] br[3] wl[56] vdd gnd cell_6t
Xbit_r57_c3 bl[3] br[3] wl[57] vdd gnd cell_6t
Xbit_r58_c3 bl[3] br[3] wl[58] vdd gnd cell_6t
Xbit_r59_c3 bl[3] br[3] wl[59] vdd gnd cell_6t
Xbit_r60_c3 bl[3] br[3] wl[60] vdd gnd cell_6t
Xbit_r61_c3 bl[3] br[3] wl[61] vdd gnd cell_6t
Xbit_r62_c3 bl[3] br[3] wl[62] vdd gnd cell_6t
Xbit_r63_c3 bl[3] br[3] wl[63] vdd gnd cell_6t
Xbit_r64_c3 bl[3] br[3] wl[64] vdd gnd cell_6t
Xbit_r65_c3 bl[3] br[3] wl[65] vdd gnd cell_6t
Xbit_r66_c3 bl[3] br[3] wl[66] vdd gnd cell_6t
Xbit_r67_c3 bl[3] br[3] wl[67] vdd gnd cell_6t
Xbit_r68_c3 bl[3] br[3] wl[68] vdd gnd cell_6t
Xbit_r69_c3 bl[3] br[3] wl[69] vdd gnd cell_6t
Xbit_r70_c3 bl[3] br[3] wl[70] vdd gnd cell_6t
Xbit_r71_c3 bl[3] br[3] wl[71] vdd gnd cell_6t
Xbit_r72_c3 bl[3] br[3] wl[72] vdd gnd cell_6t
Xbit_r73_c3 bl[3] br[3] wl[73] vdd gnd cell_6t
Xbit_r74_c3 bl[3] br[3] wl[74] vdd gnd cell_6t
Xbit_r75_c3 bl[3] br[3] wl[75] vdd gnd cell_6t
Xbit_r76_c3 bl[3] br[3] wl[76] vdd gnd cell_6t
Xbit_r77_c3 bl[3] br[3] wl[77] vdd gnd cell_6t
Xbit_r78_c3 bl[3] br[3] wl[78] vdd gnd cell_6t
Xbit_r79_c3 bl[3] br[3] wl[79] vdd gnd cell_6t
Xbit_r80_c3 bl[3] br[3] wl[80] vdd gnd cell_6t
Xbit_r81_c3 bl[3] br[3] wl[81] vdd gnd cell_6t
Xbit_r82_c3 bl[3] br[3] wl[82] vdd gnd cell_6t
Xbit_r83_c3 bl[3] br[3] wl[83] vdd gnd cell_6t
Xbit_r84_c3 bl[3] br[3] wl[84] vdd gnd cell_6t
Xbit_r85_c3 bl[3] br[3] wl[85] vdd gnd cell_6t
Xbit_r86_c3 bl[3] br[3] wl[86] vdd gnd cell_6t
Xbit_r87_c3 bl[3] br[3] wl[87] vdd gnd cell_6t
Xbit_r88_c3 bl[3] br[3] wl[88] vdd gnd cell_6t
Xbit_r89_c3 bl[3] br[3] wl[89] vdd gnd cell_6t
Xbit_r90_c3 bl[3] br[3] wl[90] vdd gnd cell_6t
Xbit_r91_c3 bl[3] br[3] wl[91] vdd gnd cell_6t
Xbit_r92_c3 bl[3] br[3] wl[92] vdd gnd cell_6t
Xbit_r93_c3 bl[3] br[3] wl[93] vdd gnd cell_6t
Xbit_r94_c3 bl[3] br[3] wl[94] vdd gnd cell_6t
Xbit_r95_c3 bl[3] br[3] wl[95] vdd gnd cell_6t
Xbit_r96_c3 bl[3] br[3] wl[96] vdd gnd cell_6t
Xbit_r97_c3 bl[3] br[3] wl[97] vdd gnd cell_6t
Xbit_r98_c3 bl[3] br[3] wl[98] vdd gnd cell_6t
Xbit_r99_c3 bl[3] br[3] wl[99] vdd gnd cell_6t
Xbit_r100_c3 bl[3] br[3] wl[100] vdd gnd cell_6t
Xbit_r101_c3 bl[3] br[3] wl[101] vdd gnd cell_6t
Xbit_r102_c3 bl[3] br[3] wl[102] vdd gnd cell_6t
Xbit_r103_c3 bl[3] br[3] wl[103] vdd gnd cell_6t
Xbit_r104_c3 bl[3] br[3] wl[104] vdd gnd cell_6t
Xbit_r105_c3 bl[3] br[3] wl[105] vdd gnd cell_6t
Xbit_r106_c3 bl[3] br[3] wl[106] vdd gnd cell_6t
Xbit_r107_c3 bl[3] br[3] wl[107] vdd gnd cell_6t
Xbit_r108_c3 bl[3] br[3] wl[108] vdd gnd cell_6t
Xbit_r109_c3 bl[3] br[3] wl[109] vdd gnd cell_6t
Xbit_r110_c3 bl[3] br[3] wl[110] vdd gnd cell_6t
Xbit_r111_c3 bl[3] br[3] wl[111] vdd gnd cell_6t
Xbit_r112_c3 bl[3] br[3] wl[112] vdd gnd cell_6t
Xbit_r113_c3 bl[3] br[3] wl[113] vdd gnd cell_6t
Xbit_r114_c3 bl[3] br[3] wl[114] vdd gnd cell_6t
Xbit_r115_c3 bl[3] br[3] wl[115] vdd gnd cell_6t
Xbit_r116_c3 bl[3] br[3] wl[116] vdd gnd cell_6t
Xbit_r117_c3 bl[3] br[3] wl[117] vdd gnd cell_6t
Xbit_r118_c3 bl[3] br[3] wl[118] vdd gnd cell_6t
Xbit_r119_c3 bl[3] br[3] wl[119] vdd gnd cell_6t
Xbit_r120_c3 bl[3] br[3] wl[120] vdd gnd cell_6t
Xbit_r121_c3 bl[3] br[3] wl[121] vdd gnd cell_6t
Xbit_r122_c3 bl[3] br[3] wl[122] vdd gnd cell_6t
Xbit_r123_c3 bl[3] br[3] wl[123] vdd gnd cell_6t
Xbit_r124_c3 bl[3] br[3] wl[124] vdd gnd cell_6t
Xbit_r125_c3 bl[3] br[3] wl[125] vdd gnd cell_6t
Xbit_r126_c3 bl[3] br[3] wl[126] vdd gnd cell_6t
Xbit_r127_c3 bl[3] br[3] wl[127] vdd gnd cell_6t
Xbit_r0_c4 bl[4] br[4] wl[0] vdd gnd cell_6t
Xbit_r1_c4 bl[4] br[4] wl[1] vdd gnd cell_6t
Xbit_r2_c4 bl[4] br[4] wl[2] vdd gnd cell_6t
Xbit_r3_c4 bl[4] br[4] wl[3] vdd gnd cell_6t
Xbit_r4_c4 bl[4] br[4] wl[4] vdd gnd cell_6t
Xbit_r5_c4 bl[4] br[4] wl[5] vdd gnd cell_6t
Xbit_r6_c4 bl[4] br[4] wl[6] vdd gnd cell_6t
Xbit_r7_c4 bl[4] br[4] wl[7] vdd gnd cell_6t
Xbit_r8_c4 bl[4] br[4] wl[8] vdd gnd cell_6t
Xbit_r9_c4 bl[4] br[4] wl[9] vdd gnd cell_6t
Xbit_r10_c4 bl[4] br[4] wl[10] vdd gnd cell_6t
Xbit_r11_c4 bl[4] br[4] wl[11] vdd gnd cell_6t
Xbit_r12_c4 bl[4] br[4] wl[12] vdd gnd cell_6t
Xbit_r13_c4 bl[4] br[4] wl[13] vdd gnd cell_6t
Xbit_r14_c4 bl[4] br[4] wl[14] vdd gnd cell_6t
Xbit_r15_c4 bl[4] br[4] wl[15] vdd gnd cell_6t
Xbit_r16_c4 bl[4] br[4] wl[16] vdd gnd cell_6t
Xbit_r17_c4 bl[4] br[4] wl[17] vdd gnd cell_6t
Xbit_r18_c4 bl[4] br[4] wl[18] vdd gnd cell_6t
Xbit_r19_c4 bl[4] br[4] wl[19] vdd gnd cell_6t
Xbit_r20_c4 bl[4] br[4] wl[20] vdd gnd cell_6t
Xbit_r21_c4 bl[4] br[4] wl[21] vdd gnd cell_6t
Xbit_r22_c4 bl[4] br[4] wl[22] vdd gnd cell_6t
Xbit_r23_c4 bl[4] br[4] wl[23] vdd gnd cell_6t
Xbit_r24_c4 bl[4] br[4] wl[24] vdd gnd cell_6t
Xbit_r25_c4 bl[4] br[4] wl[25] vdd gnd cell_6t
Xbit_r26_c4 bl[4] br[4] wl[26] vdd gnd cell_6t
Xbit_r27_c4 bl[4] br[4] wl[27] vdd gnd cell_6t
Xbit_r28_c4 bl[4] br[4] wl[28] vdd gnd cell_6t
Xbit_r29_c4 bl[4] br[4] wl[29] vdd gnd cell_6t
Xbit_r30_c4 bl[4] br[4] wl[30] vdd gnd cell_6t
Xbit_r31_c4 bl[4] br[4] wl[31] vdd gnd cell_6t
Xbit_r32_c4 bl[4] br[4] wl[32] vdd gnd cell_6t
Xbit_r33_c4 bl[4] br[4] wl[33] vdd gnd cell_6t
Xbit_r34_c4 bl[4] br[4] wl[34] vdd gnd cell_6t
Xbit_r35_c4 bl[4] br[4] wl[35] vdd gnd cell_6t
Xbit_r36_c4 bl[4] br[4] wl[36] vdd gnd cell_6t
Xbit_r37_c4 bl[4] br[4] wl[37] vdd gnd cell_6t
Xbit_r38_c4 bl[4] br[4] wl[38] vdd gnd cell_6t
Xbit_r39_c4 bl[4] br[4] wl[39] vdd gnd cell_6t
Xbit_r40_c4 bl[4] br[4] wl[40] vdd gnd cell_6t
Xbit_r41_c4 bl[4] br[4] wl[41] vdd gnd cell_6t
Xbit_r42_c4 bl[4] br[4] wl[42] vdd gnd cell_6t
Xbit_r43_c4 bl[4] br[4] wl[43] vdd gnd cell_6t
Xbit_r44_c4 bl[4] br[4] wl[44] vdd gnd cell_6t
Xbit_r45_c4 bl[4] br[4] wl[45] vdd gnd cell_6t
Xbit_r46_c4 bl[4] br[4] wl[46] vdd gnd cell_6t
Xbit_r47_c4 bl[4] br[4] wl[47] vdd gnd cell_6t
Xbit_r48_c4 bl[4] br[4] wl[48] vdd gnd cell_6t
Xbit_r49_c4 bl[4] br[4] wl[49] vdd gnd cell_6t
Xbit_r50_c4 bl[4] br[4] wl[50] vdd gnd cell_6t
Xbit_r51_c4 bl[4] br[4] wl[51] vdd gnd cell_6t
Xbit_r52_c4 bl[4] br[4] wl[52] vdd gnd cell_6t
Xbit_r53_c4 bl[4] br[4] wl[53] vdd gnd cell_6t
Xbit_r54_c4 bl[4] br[4] wl[54] vdd gnd cell_6t
Xbit_r55_c4 bl[4] br[4] wl[55] vdd gnd cell_6t
Xbit_r56_c4 bl[4] br[4] wl[56] vdd gnd cell_6t
Xbit_r57_c4 bl[4] br[4] wl[57] vdd gnd cell_6t
Xbit_r58_c4 bl[4] br[4] wl[58] vdd gnd cell_6t
Xbit_r59_c4 bl[4] br[4] wl[59] vdd gnd cell_6t
Xbit_r60_c4 bl[4] br[4] wl[60] vdd gnd cell_6t
Xbit_r61_c4 bl[4] br[4] wl[61] vdd gnd cell_6t
Xbit_r62_c4 bl[4] br[4] wl[62] vdd gnd cell_6t
Xbit_r63_c4 bl[4] br[4] wl[63] vdd gnd cell_6t
Xbit_r64_c4 bl[4] br[4] wl[64] vdd gnd cell_6t
Xbit_r65_c4 bl[4] br[4] wl[65] vdd gnd cell_6t
Xbit_r66_c4 bl[4] br[4] wl[66] vdd gnd cell_6t
Xbit_r67_c4 bl[4] br[4] wl[67] vdd gnd cell_6t
Xbit_r68_c4 bl[4] br[4] wl[68] vdd gnd cell_6t
Xbit_r69_c4 bl[4] br[4] wl[69] vdd gnd cell_6t
Xbit_r70_c4 bl[4] br[4] wl[70] vdd gnd cell_6t
Xbit_r71_c4 bl[4] br[4] wl[71] vdd gnd cell_6t
Xbit_r72_c4 bl[4] br[4] wl[72] vdd gnd cell_6t
Xbit_r73_c4 bl[4] br[4] wl[73] vdd gnd cell_6t
Xbit_r74_c4 bl[4] br[4] wl[74] vdd gnd cell_6t
Xbit_r75_c4 bl[4] br[4] wl[75] vdd gnd cell_6t
Xbit_r76_c4 bl[4] br[4] wl[76] vdd gnd cell_6t
Xbit_r77_c4 bl[4] br[4] wl[77] vdd gnd cell_6t
Xbit_r78_c4 bl[4] br[4] wl[78] vdd gnd cell_6t
Xbit_r79_c4 bl[4] br[4] wl[79] vdd gnd cell_6t
Xbit_r80_c4 bl[4] br[4] wl[80] vdd gnd cell_6t
Xbit_r81_c4 bl[4] br[4] wl[81] vdd gnd cell_6t
Xbit_r82_c4 bl[4] br[4] wl[82] vdd gnd cell_6t
Xbit_r83_c4 bl[4] br[4] wl[83] vdd gnd cell_6t
Xbit_r84_c4 bl[4] br[4] wl[84] vdd gnd cell_6t
Xbit_r85_c4 bl[4] br[4] wl[85] vdd gnd cell_6t
Xbit_r86_c4 bl[4] br[4] wl[86] vdd gnd cell_6t
Xbit_r87_c4 bl[4] br[4] wl[87] vdd gnd cell_6t
Xbit_r88_c4 bl[4] br[4] wl[88] vdd gnd cell_6t
Xbit_r89_c4 bl[4] br[4] wl[89] vdd gnd cell_6t
Xbit_r90_c4 bl[4] br[4] wl[90] vdd gnd cell_6t
Xbit_r91_c4 bl[4] br[4] wl[91] vdd gnd cell_6t
Xbit_r92_c4 bl[4] br[4] wl[92] vdd gnd cell_6t
Xbit_r93_c4 bl[4] br[4] wl[93] vdd gnd cell_6t
Xbit_r94_c4 bl[4] br[4] wl[94] vdd gnd cell_6t
Xbit_r95_c4 bl[4] br[4] wl[95] vdd gnd cell_6t
Xbit_r96_c4 bl[4] br[4] wl[96] vdd gnd cell_6t
Xbit_r97_c4 bl[4] br[4] wl[97] vdd gnd cell_6t
Xbit_r98_c4 bl[4] br[4] wl[98] vdd gnd cell_6t
Xbit_r99_c4 bl[4] br[4] wl[99] vdd gnd cell_6t
Xbit_r100_c4 bl[4] br[4] wl[100] vdd gnd cell_6t
Xbit_r101_c4 bl[4] br[4] wl[101] vdd gnd cell_6t
Xbit_r102_c4 bl[4] br[4] wl[102] vdd gnd cell_6t
Xbit_r103_c4 bl[4] br[4] wl[103] vdd gnd cell_6t
Xbit_r104_c4 bl[4] br[4] wl[104] vdd gnd cell_6t
Xbit_r105_c4 bl[4] br[4] wl[105] vdd gnd cell_6t
Xbit_r106_c4 bl[4] br[4] wl[106] vdd gnd cell_6t
Xbit_r107_c4 bl[4] br[4] wl[107] vdd gnd cell_6t
Xbit_r108_c4 bl[4] br[4] wl[108] vdd gnd cell_6t
Xbit_r109_c4 bl[4] br[4] wl[109] vdd gnd cell_6t
Xbit_r110_c4 bl[4] br[4] wl[110] vdd gnd cell_6t
Xbit_r111_c4 bl[4] br[4] wl[111] vdd gnd cell_6t
Xbit_r112_c4 bl[4] br[4] wl[112] vdd gnd cell_6t
Xbit_r113_c4 bl[4] br[4] wl[113] vdd gnd cell_6t
Xbit_r114_c4 bl[4] br[4] wl[114] vdd gnd cell_6t
Xbit_r115_c4 bl[4] br[4] wl[115] vdd gnd cell_6t
Xbit_r116_c4 bl[4] br[4] wl[116] vdd gnd cell_6t
Xbit_r117_c4 bl[4] br[4] wl[117] vdd gnd cell_6t
Xbit_r118_c4 bl[4] br[4] wl[118] vdd gnd cell_6t
Xbit_r119_c4 bl[4] br[4] wl[119] vdd gnd cell_6t
Xbit_r120_c4 bl[4] br[4] wl[120] vdd gnd cell_6t
Xbit_r121_c4 bl[4] br[4] wl[121] vdd gnd cell_6t
Xbit_r122_c4 bl[4] br[4] wl[122] vdd gnd cell_6t
Xbit_r123_c4 bl[4] br[4] wl[123] vdd gnd cell_6t
Xbit_r124_c4 bl[4] br[4] wl[124] vdd gnd cell_6t
Xbit_r125_c4 bl[4] br[4] wl[125] vdd gnd cell_6t
Xbit_r126_c4 bl[4] br[4] wl[126] vdd gnd cell_6t
Xbit_r127_c4 bl[4] br[4] wl[127] vdd gnd cell_6t
Xbit_r0_c5 bl[5] br[5] wl[0] vdd gnd cell_6t
Xbit_r1_c5 bl[5] br[5] wl[1] vdd gnd cell_6t
Xbit_r2_c5 bl[5] br[5] wl[2] vdd gnd cell_6t
Xbit_r3_c5 bl[5] br[5] wl[3] vdd gnd cell_6t
Xbit_r4_c5 bl[5] br[5] wl[4] vdd gnd cell_6t
Xbit_r5_c5 bl[5] br[5] wl[5] vdd gnd cell_6t
Xbit_r6_c5 bl[5] br[5] wl[6] vdd gnd cell_6t
Xbit_r7_c5 bl[5] br[5] wl[7] vdd gnd cell_6t
Xbit_r8_c5 bl[5] br[5] wl[8] vdd gnd cell_6t
Xbit_r9_c5 bl[5] br[5] wl[9] vdd gnd cell_6t
Xbit_r10_c5 bl[5] br[5] wl[10] vdd gnd cell_6t
Xbit_r11_c5 bl[5] br[5] wl[11] vdd gnd cell_6t
Xbit_r12_c5 bl[5] br[5] wl[12] vdd gnd cell_6t
Xbit_r13_c5 bl[5] br[5] wl[13] vdd gnd cell_6t
Xbit_r14_c5 bl[5] br[5] wl[14] vdd gnd cell_6t
Xbit_r15_c5 bl[5] br[5] wl[15] vdd gnd cell_6t
Xbit_r16_c5 bl[5] br[5] wl[16] vdd gnd cell_6t
Xbit_r17_c5 bl[5] br[5] wl[17] vdd gnd cell_6t
Xbit_r18_c5 bl[5] br[5] wl[18] vdd gnd cell_6t
Xbit_r19_c5 bl[5] br[5] wl[19] vdd gnd cell_6t
Xbit_r20_c5 bl[5] br[5] wl[20] vdd gnd cell_6t
Xbit_r21_c5 bl[5] br[5] wl[21] vdd gnd cell_6t
Xbit_r22_c5 bl[5] br[5] wl[22] vdd gnd cell_6t
Xbit_r23_c5 bl[5] br[5] wl[23] vdd gnd cell_6t
Xbit_r24_c5 bl[5] br[5] wl[24] vdd gnd cell_6t
Xbit_r25_c5 bl[5] br[5] wl[25] vdd gnd cell_6t
Xbit_r26_c5 bl[5] br[5] wl[26] vdd gnd cell_6t
Xbit_r27_c5 bl[5] br[5] wl[27] vdd gnd cell_6t
Xbit_r28_c5 bl[5] br[5] wl[28] vdd gnd cell_6t
Xbit_r29_c5 bl[5] br[5] wl[29] vdd gnd cell_6t
Xbit_r30_c5 bl[5] br[5] wl[30] vdd gnd cell_6t
Xbit_r31_c5 bl[5] br[5] wl[31] vdd gnd cell_6t
Xbit_r32_c5 bl[5] br[5] wl[32] vdd gnd cell_6t
Xbit_r33_c5 bl[5] br[5] wl[33] vdd gnd cell_6t
Xbit_r34_c5 bl[5] br[5] wl[34] vdd gnd cell_6t
Xbit_r35_c5 bl[5] br[5] wl[35] vdd gnd cell_6t
Xbit_r36_c5 bl[5] br[5] wl[36] vdd gnd cell_6t
Xbit_r37_c5 bl[5] br[5] wl[37] vdd gnd cell_6t
Xbit_r38_c5 bl[5] br[5] wl[38] vdd gnd cell_6t
Xbit_r39_c5 bl[5] br[5] wl[39] vdd gnd cell_6t
Xbit_r40_c5 bl[5] br[5] wl[40] vdd gnd cell_6t
Xbit_r41_c5 bl[5] br[5] wl[41] vdd gnd cell_6t
Xbit_r42_c5 bl[5] br[5] wl[42] vdd gnd cell_6t
Xbit_r43_c5 bl[5] br[5] wl[43] vdd gnd cell_6t
Xbit_r44_c5 bl[5] br[5] wl[44] vdd gnd cell_6t
Xbit_r45_c5 bl[5] br[5] wl[45] vdd gnd cell_6t
Xbit_r46_c5 bl[5] br[5] wl[46] vdd gnd cell_6t
Xbit_r47_c5 bl[5] br[5] wl[47] vdd gnd cell_6t
Xbit_r48_c5 bl[5] br[5] wl[48] vdd gnd cell_6t
Xbit_r49_c5 bl[5] br[5] wl[49] vdd gnd cell_6t
Xbit_r50_c5 bl[5] br[5] wl[50] vdd gnd cell_6t
Xbit_r51_c5 bl[5] br[5] wl[51] vdd gnd cell_6t
Xbit_r52_c5 bl[5] br[5] wl[52] vdd gnd cell_6t
Xbit_r53_c5 bl[5] br[5] wl[53] vdd gnd cell_6t
Xbit_r54_c5 bl[5] br[5] wl[54] vdd gnd cell_6t
Xbit_r55_c5 bl[5] br[5] wl[55] vdd gnd cell_6t
Xbit_r56_c5 bl[5] br[5] wl[56] vdd gnd cell_6t
Xbit_r57_c5 bl[5] br[5] wl[57] vdd gnd cell_6t
Xbit_r58_c5 bl[5] br[5] wl[58] vdd gnd cell_6t
Xbit_r59_c5 bl[5] br[5] wl[59] vdd gnd cell_6t
Xbit_r60_c5 bl[5] br[5] wl[60] vdd gnd cell_6t
Xbit_r61_c5 bl[5] br[5] wl[61] vdd gnd cell_6t
Xbit_r62_c5 bl[5] br[5] wl[62] vdd gnd cell_6t
Xbit_r63_c5 bl[5] br[5] wl[63] vdd gnd cell_6t
Xbit_r64_c5 bl[5] br[5] wl[64] vdd gnd cell_6t
Xbit_r65_c5 bl[5] br[5] wl[65] vdd gnd cell_6t
Xbit_r66_c5 bl[5] br[5] wl[66] vdd gnd cell_6t
Xbit_r67_c5 bl[5] br[5] wl[67] vdd gnd cell_6t
Xbit_r68_c5 bl[5] br[5] wl[68] vdd gnd cell_6t
Xbit_r69_c5 bl[5] br[5] wl[69] vdd gnd cell_6t
Xbit_r70_c5 bl[5] br[5] wl[70] vdd gnd cell_6t
Xbit_r71_c5 bl[5] br[5] wl[71] vdd gnd cell_6t
Xbit_r72_c5 bl[5] br[5] wl[72] vdd gnd cell_6t
Xbit_r73_c5 bl[5] br[5] wl[73] vdd gnd cell_6t
Xbit_r74_c5 bl[5] br[5] wl[74] vdd gnd cell_6t
Xbit_r75_c5 bl[5] br[5] wl[75] vdd gnd cell_6t
Xbit_r76_c5 bl[5] br[5] wl[76] vdd gnd cell_6t
Xbit_r77_c5 bl[5] br[5] wl[77] vdd gnd cell_6t
Xbit_r78_c5 bl[5] br[5] wl[78] vdd gnd cell_6t
Xbit_r79_c5 bl[5] br[5] wl[79] vdd gnd cell_6t
Xbit_r80_c5 bl[5] br[5] wl[80] vdd gnd cell_6t
Xbit_r81_c5 bl[5] br[5] wl[81] vdd gnd cell_6t
Xbit_r82_c5 bl[5] br[5] wl[82] vdd gnd cell_6t
Xbit_r83_c5 bl[5] br[5] wl[83] vdd gnd cell_6t
Xbit_r84_c5 bl[5] br[5] wl[84] vdd gnd cell_6t
Xbit_r85_c5 bl[5] br[5] wl[85] vdd gnd cell_6t
Xbit_r86_c5 bl[5] br[5] wl[86] vdd gnd cell_6t
Xbit_r87_c5 bl[5] br[5] wl[87] vdd gnd cell_6t
Xbit_r88_c5 bl[5] br[5] wl[88] vdd gnd cell_6t
Xbit_r89_c5 bl[5] br[5] wl[89] vdd gnd cell_6t
Xbit_r90_c5 bl[5] br[5] wl[90] vdd gnd cell_6t
Xbit_r91_c5 bl[5] br[5] wl[91] vdd gnd cell_6t
Xbit_r92_c5 bl[5] br[5] wl[92] vdd gnd cell_6t
Xbit_r93_c5 bl[5] br[5] wl[93] vdd gnd cell_6t
Xbit_r94_c5 bl[5] br[5] wl[94] vdd gnd cell_6t
Xbit_r95_c5 bl[5] br[5] wl[95] vdd gnd cell_6t
Xbit_r96_c5 bl[5] br[5] wl[96] vdd gnd cell_6t
Xbit_r97_c5 bl[5] br[5] wl[97] vdd gnd cell_6t
Xbit_r98_c5 bl[5] br[5] wl[98] vdd gnd cell_6t
Xbit_r99_c5 bl[5] br[5] wl[99] vdd gnd cell_6t
Xbit_r100_c5 bl[5] br[5] wl[100] vdd gnd cell_6t
Xbit_r101_c5 bl[5] br[5] wl[101] vdd gnd cell_6t
Xbit_r102_c5 bl[5] br[5] wl[102] vdd gnd cell_6t
Xbit_r103_c5 bl[5] br[5] wl[103] vdd gnd cell_6t
Xbit_r104_c5 bl[5] br[5] wl[104] vdd gnd cell_6t
Xbit_r105_c5 bl[5] br[5] wl[105] vdd gnd cell_6t
Xbit_r106_c5 bl[5] br[5] wl[106] vdd gnd cell_6t
Xbit_r107_c5 bl[5] br[5] wl[107] vdd gnd cell_6t
Xbit_r108_c5 bl[5] br[5] wl[108] vdd gnd cell_6t
Xbit_r109_c5 bl[5] br[5] wl[109] vdd gnd cell_6t
Xbit_r110_c5 bl[5] br[5] wl[110] vdd gnd cell_6t
Xbit_r111_c5 bl[5] br[5] wl[111] vdd gnd cell_6t
Xbit_r112_c5 bl[5] br[5] wl[112] vdd gnd cell_6t
Xbit_r113_c5 bl[5] br[5] wl[113] vdd gnd cell_6t
Xbit_r114_c5 bl[5] br[5] wl[114] vdd gnd cell_6t
Xbit_r115_c5 bl[5] br[5] wl[115] vdd gnd cell_6t
Xbit_r116_c5 bl[5] br[5] wl[116] vdd gnd cell_6t
Xbit_r117_c5 bl[5] br[5] wl[117] vdd gnd cell_6t
Xbit_r118_c5 bl[5] br[5] wl[118] vdd gnd cell_6t
Xbit_r119_c5 bl[5] br[5] wl[119] vdd gnd cell_6t
Xbit_r120_c5 bl[5] br[5] wl[120] vdd gnd cell_6t
Xbit_r121_c5 bl[5] br[5] wl[121] vdd gnd cell_6t
Xbit_r122_c5 bl[5] br[5] wl[122] vdd gnd cell_6t
Xbit_r123_c5 bl[5] br[5] wl[123] vdd gnd cell_6t
Xbit_r124_c5 bl[5] br[5] wl[124] vdd gnd cell_6t
Xbit_r125_c5 bl[5] br[5] wl[125] vdd gnd cell_6t
Xbit_r126_c5 bl[5] br[5] wl[126] vdd gnd cell_6t
Xbit_r127_c5 bl[5] br[5] wl[127] vdd gnd cell_6t
Xbit_r0_c6 bl[6] br[6] wl[0] vdd gnd cell_6t
Xbit_r1_c6 bl[6] br[6] wl[1] vdd gnd cell_6t
Xbit_r2_c6 bl[6] br[6] wl[2] vdd gnd cell_6t
Xbit_r3_c6 bl[6] br[6] wl[3] vdd gnd cell_6t
Xbit_r4_c6 bl[6] br[6] wl[4] vdd gnd cell_6t
Xbit_r5_c6 bl[6] br[6] wl[5] vdd gnd cell_6t
Xbit_r6_c6 bl[6] br[6] wl[6] vdd gnd cell_6t
Xbit_r7_c6 bl[6] br[6] wl[7] vdd gnd cell_6t
Xbit_r8_c6 bl[6] br[6] wl[8] vdd gnd cell_6t
Xbit_r9_c6 bl[6] br[6] wl[9] vdd gnd cell_6t
Xbit_r10_c6 bl[6] br[6] wl[10] vdd gnd cell_6t
Xbit_r11_c6 bl[6] br[6] wl[11] vdd gnd cell_6t
Xbit_r12_c6 bl[6] br[6] wl[12] vdd gnd cell_6t
Xbit_r13_c6 bl[6] br[6] wl[13] vdd gnd cell_6t
Xbit_r14_c6 bl[6] br[6] wl[14] vdd gnd cell_6t
Xbit_r15_c6 bl[6] br[6] wl[15] vdd gnd cell_6t
Xbit_r16_c6 bl[6] br[6] wl[16] vdd gnd cell_6t
Xbit_r17_c6 bl[6] br[6] wl[17] vdd gnd cell_6t
Xbit_r18_c6 bl[6] br[6] wl[18] vdd gnd cell_6t
Xbit_r19_c6 bl[6] br[6] wl[19] vdd gnd cell_6t
Xbit_r20_c6 bl[6] br[6] wl[20] vdd gnd cell_6t
Xbit_r21_c6 bl[6] br[6] wl[21] vdd gnd cell_6t
Xbit_r22_c6 bl[6] br[6] wl[22] vdd gnd cell_6t
Xbit_r23_c6 bl[6] br[6] wl[23] vdd gnd cell_6t
Xbit_r24_c6 bl[6] br[6] wl[24] vdd gnd cell_6t
Xbit_r25_c6 bl[6] br[6] wl[25] vdd gnd cell_6t
Xbit_r26_c6 bl[6] br[6] wl[26] vdd gnd cell_6t
Xbit_r27_c6 bl[6] br[6] wl[27] vdd gnd cell_6t
Xbit_r28_c6 bl[6] br[6] wl[28] vdd gnd cell_6t
Xbit_r29_c6 bl[6] br[6] wl[29] vdd gnd cell_6t
Xbit_r30_c6 bl[6] br[6] wl[30] vdd gnd cell_6t
Xbit_r31_c6 bl[6] br[6] wl[31] vdd gnd cell_6t
Xbit_r32_c6 bl[6] br[6] wl[32] vdd gnd cell_6t
Xbit_r33_c6 bl[6] br[6] wl[33] vdd gnd cell_6t
Xbit_r34_c6 bl[6] br[6] wl[34] vdd gnd cell_6t
Xbit_r35_c6 bl[6] br[6] wl[35] vdd gnd cell_6t
Xbit_r36_c6 bl[6] br[6] wl[36] vdd gnd cell_6t
Xbit_r37_c6 bl[6] br[6] wl[37] vdd gnd cell_6t
Xbit_r38_c6 bl[6] br[6] wl[38] vdd gnd cell_6t
Xbit_r39_c6 bl[6] br[6] wl[39] vdd gnd cell_6t
Xbit_r40_c6 bl[6] br[6] wl[40] vdd gnd cell_6t
Xbit_r41_c6 bl[6] br[6] wl[41] vdd gnd cell_6t
Xbit_r42_c6 bl[6] br[6] wl[42] vdd gnd cell_6t
Xbit_r43_c6 bl[6] br[6] wl[43] vdd gnd cell_6t
Xbit_r44_c6 bl[6] br[6] wl[44] vdd gnd cell_6t
Xbit_r45_c6 bl[6] br[6] wl[45] vdd gnd cell_6t
Xbit_r46_c6 bl[6] br[6] wl[46] vdd gnd cell_6t
Xbit_r47_c6 bl[6] br[6] wl[47] vdd gnd cell_6t
Xbit_r48_c6 bl[6] br[6] wl[48] vdd gnd cell_6t
Xbit_r49_c6 bl[6] br[6] wl[49] vdd gnd cell_6t
Xbit_r50_c6 bl[6] br[6] wl[50] vdd gnd cell_6t
Xbit_r51_c6 bl[6] br[6] wl[51] vdd gnd cell_6t
Xbit_r52_c6 bl[6] br[6] wl[52] vdd gnd cell_6t
Xbit_r53_c6 bl[6] br[6] wl[53] vdd gnd cell_6t
Xbit_r54_c6 bl[6] br[6] wl[54] vdd gnd cell_6t
Xbit_r55_c6 bl[6] br[6] wl[55] vdd gnd cell_6t
Xbit_r56_c6 bl[6] br[6] wl[56] vdd gnd cell_6t
Xbit_r57_c6 bl[6] br[6] wl[57] vdd gnd cell_6t
Xbit_r58_c6 bl[6] br[6] wl[58] vdd gnd cell_6t
Xbit_r59_c6 bl[6] br[6] wl[59] vdd gnd cell_6t
Xbit_r60_c6 bl[6] br[6] wl[60] vdd gnd cell_6t
Xbit_r61_c6 bl[6] br[6] wl[61] vdd gnd cell_6t
Xbit_r62_c6 bl[6] br[6] wl[62] vdd gnd cell_6t
Xbit_r63_c6 bl[6] br[6] wl[63] vdd gnd cell_6t
Xbit_r64_c6 bl[6] br[6] wl[64] vdd gnd cell_6t
Xbit_r65_c6 bl[6] br[6] wl[65] vdd gnd cell_6t
Xbit_r66_c6 bl[6] br[6] wl[66] vdd gnd cell_6t
Xbit_r67_c6 bl[6] br[6] wl[67] vdd gnd cell_6t
Xbit_r68_c6 bl[6] br[6] wl[68] vdd gnd cell_6t
Xbit_r69_c6 bl[6] br[6] wl[69] vdd gnd cell_6t
Xbit_r70_c6 bl[6] br[6] wl[70] vdd gnd cell_6t
Xbit_r71_c6 bl[6] br[6] wl[71] vdd gnd cell_6t
Xbit_r72_c6 bl[6] br[6] wl[72] vdd gnd cell_6t
Xbit_r73_c6 bl[6] br[6] wl[73] vdd gnd cell_6t
Xbit_r74_c6 bl[6] br[6] wl[74] vdd gnd cell_6t
Xbit_r75_c6 bl[6] br[6] wl[75] vdd gnd cell_6t
Xbit_r76_c6 bl[6] br[6] wl[76] vdd gnd cell_6t
Xbit_r77_c6 bl[6] br[6] wl[77] vdd gnd cell_6t
Xbit_r78_c6 bl[6] br[6] wl[78] vdd gnd cell_6t
Xbit_r79_c6 bl[6] br[6] wl[79] vdd gnd cell_6t
Xbit_r80_c6 bl[6] br[6] wl[80] vdd gnd cell_6t
Xbit_r81_c6 bl[6] br[6] wl[81] vdd gnd cell_6t
Xbit_r82_c6 bl[6] br[6] wl[82] vdd gnd cell_6t
Xbit_r83_c6 bl[6] br[6] wl[83] vdd gnd cell_6t
Xbit_r84_c6 bl[6] br[6] wl[84] vdd gnd cell_6t
Xbit_r85_c6 bl[6] br[6] wl[85] vdd gnd cell_6t
Xbit_r86_c6 bl[6] br[6] wl[86] vdd gnd cell_6t
Xbit_r87_c6 bl[6] br[6] wl[87] vdd gnd cell_6t
Xbit_r88_c6 bl[6] br[6] wl[88] vdd gnd cell_6t
Xbit_r89_c6 bl[6] br[6] wl[89] vdd gnd cell_6t
Xbit_r90_c6 bl[6] br[6] wl[90] vdd gnd cell_6t
Xbit_r91_c6 bl[6] br[6] wl[91] vdd gnd cell_6t
Xbit_r92_c6 bl[6] br[6] wl[92] vdd gnd cell_6t
Xbit_r93_c6 bl[6] br[6] wl[93] vdd gnd cell_6t
Xbit_r94_c6 bl[6] br[6] wl[94] vdd gnd cell_6t
Xbit_r95_c6 bl[6] br[6] wl[95] vdd gnd cell_6t
Xbit_r96_c6 bl[6] br[6] wl[96] vdd gnd cell_6t
Xbit_r97_c6 bl[6] br[6] wl[97] vdd gnd cell_6t
Xbit_r98_c6 bl[6] br[6] wl[98] vdd gnd cell_6t
Xbit_r99_c6 bl[6] br[6] wl[99] vdd gnd cell_6t
Xbit_r100_c6 bl[6] br[6] wl[100] vdd gnd cell_6t
Xbit_r101_c6 bl[6] br[6] wl[101] vdd gnd cell_6t
Xbit_r102_c6 bl[6] br[6] wl[102] vdd gnd cell_6t
Xbit_r103_c6 bl[6] br[6] wl[103] vdd gnd cell_6t
Xbit_r104_c6 bl[6] br[6] wl[104] vdd gnd cell_6t
Xbit_r105_c6 bl[6] br[6] wl[105] vdd gnd cell_6t
Xbit_r106_c6 bl[6] br[6] wl[106] vdd gnd cell_6t
Xbit_r107_c6 bl[6] br[6] wl[107] vdd gnd cell_6t
Xbit_r108_c6 bl[6] br[6] wl[108] vdd gnd cell_6t
Xbit_r109_c6 bl[6] br[6] wl[109] vdd gnd cell_6t
Xbit_r110_c6 bl[6] br[6] wl[110] vdd gnd cell_6t
Xbit_r111_c6 bl[6] br[6] wl[111] vdd gnd cell_6t
Xbit_r112_c6 bl[6] br[6] wl[112] vdd gnd cell_6t
Xbit_r113_c6 bl[6] br[6] wl[113] vdd gnd cell_6t
Xbit_r114_c6 bl[6] br[6] wl[114] vdd gnd cell_6t
Xbit_r115_c6 bl[6] br[6] wl[115] vdd gnd cell_6t
Xbit_r116_c6 bl[6] br[6] wl[116] vdd gnd cell_6t
Xbit_r117_c6 bl[6] br[6] wl[117] vdd gnd cell_6t
Xbit_r118_c6 bl[6] br[6] wl[118] vdd gnd cell_6t
Xbit_r119_c6 bl[6] br[6] wl[119] vdd gnd cell_6t
Xbit_r120_c6 bl[6] br[6] wl[120] vdd gnd cell_6t
Xbit_r121_c6 bl[6] br[6] wl[121] vdd gnd cell_6t
Xbit_r122_c6 bl[6] br[6] wl[122] vdd gnd cell_6t
Xbit_r123_c6 bl[6] br[6] wl[123] vdd gnd cell_6t
Xbit_r124_c6 bl[6] br[6] wl[124] vdd gnd cell_6t
Xbit_r125_c6 bl[6] br[6] wl[125] vdd gnd cell_6t
Xbit_r126_c6 bl[6] br[6] wl[126] vdd gnd cell_6t
Xbit_r127_c6 bl[6] br[6] wl[127] vdd gnd cell_6t
Xbit_r0_c7 bl[7] br[7] wl[0] vdd gnd cell_6t
Xbit_r1_c7 bl[7] br[7] wl[1] vdd gnd cell_6t
Xbit_r2_c7 bl[7] br[7] wl[2] vdd gnd cell_6t
Xbit_r3_c7 bl[7] br[7] wl[3] vdd gnd cell_6t
Xbit_r4_c7 bl[7] br[7] wl[4] vdd gnd cell_6t
Xbit_r5_c7 bl[7] br[7] wl[5] vdd gnd cell_6t
Xbit_r6_c7 bl[7] br[7] wl[6] vdd gnd cell_6t
Xbit_r7_c7 bl[7] br[7] wl[7] vdd gnd cell_6t
Xbit_r8_c7 bl[7] br[7] wl[8] vdd gnd cell_6t
Xbit_r9_c7 bl[7] br[7] wl[9] vdd gnd cell_6t
Xbit_r10_c7 bl[7] br[7] wl[10] vdd gnd cell_6t
Xbit_r11_c7 bl[7] br[7] wl[11] vdd gnd cell_6t
Xbit_r12_c7 bl[7] br[7] wl[12] vdd gnd cell_6t
Xbit_r13_c7 bl[7] br[7] wl[13] vdd gnd cell_6t
Xbit_r14_c7 bl[7] br[7] wl[14] vdd gnd cell_6t
Xbit_r15_c7 bl[7] br[7] wl[15] vdd gnd cell_6t
Xbit_r16_c7 bl[7] br[7] wl[16] vdd gnd cell_6t
Xbit_r17_c7 bl[7] br[7] wl[17] vdd gnd cell_6t
Xbit_r18_c7 bl[7] br[7] wl[18] vdd gnd cell_6t
Xbit_r19_c7 bl[7] br[7] wl[19] vdd gnd cell_6t
Xbit_r20_c7 bl[7] br[7] wl[20] vdd gnd cell_6t
Xbit_r21_c7 bl[7] br[7] wl[21] vdd gnd cell_6t
Xbit_r22_c7 bl[7] br[7] wl[22] vdd gnd cell_6t
Xbit_r23_c7 bl[7] br[7] wl[23] vdd gnd cell_6t
Xbit_r24_c7 bl[7] br[7] wl[24] vdd gnd cell_6t
Xbit_r25_c7 bl[7] br[7] wl[25] vdd gnd cell_6t
Xbit_r26_c7 bl[7] br[7] wl[26] vdd gnd cell_6t
Xbit_r27_c7 bl[7] br[7] wl[27] vdd gnd cell_6t
Xbit_r28_c7 bl[7] br[7] wl[28] vdd gnd cell_6t
Xbit_r29_c7 bl[7] br[7] wl[29] vdd gnd cell_6t
Xbit_r30_c7 bl[7] br[7] wl[30] vdd gnd cell_6t
Xbit_r31_c7 bl[7] br[7] wl[31] vdd gnd cell_6t
Xbit_r32_c7 bl[7] br[7] wl[32] vdd gnd cell_6t
Xbit_r33_c7 bl[7] br[7] wl[33] vdd gnd cell_6t
Xbit_r34_c7 bl[7] br[7] wl[34] vdd gnd cell_6t
Xbit_r35_c7 bl[7] br[7] wl[35] vdd gnd cell_6t
Xbit_r36_c7 bl[7] br[7] wl[36] vdd gnd cell_6t
Xbit_r37_c7 bl[7] br[7] wl[37] vdd gnd cell_6t
Xbit_r38_c7 bl[7] br[7] wl[38] vdd gnd cell_6t
Xbit_r39_c7 bl[7] br[7] wl[39] vdd gnd cell_6t
Xbit_r40_c7 bl[7] br[7] wl[40] vdd gnd cell_6t
Xbit_r41_c7 bl[7] br[7] wl[41] vdd gnd cell_6t
Xbit_r42_c7 bl[7] br[7] wl[42] vdd gnd cell_6t
Xbit_r43_c7 bl[7] br[7] wl[43] vdd gnd cell_6t
Xbit_r44_c7 bl[7] br[7] wl[44] vdd gnd cell_6t
Xbit_r45_c7 bl[7] br[7] wl[45] vdd gnd cell_6t
Xbit_r46_c7 bl[7] br[7] wl[46] vdd gnd cell_6t
Xbit_r47_c7 bl[7] br[7] wl[47] vdd gnd cell_6t
Xbit_r48_c7 bl[7] br[7] wl[48] vdd gnd cell_6t
Xbit_r49_c7 bl[7] br[7] wl[49] vdd gnd cell_6t
Xbit_r50_c7 bl[7] br[7] wl[50] vdd gnd cell_6t
Xbit_r51_c7 bl[7] br[7] wl[51] vdd gnd cell_6t
Xbit_r52_c7 bl[7] br[7] wl[52] vdd gnd cell_6t
Xbit_r53_c7 bl[7] br[7] wl[53] vdd gnd cell_6t
Xbit_r54_c7 bl[7] br[7] wl[54] vdd gnd cell_6t
Xbit_r55_c7 bl[7] br[7] wl[55] vdd gnd cell_6t
Xbit_r56_c7 bl[7] br[7] wl[56] vdd gnd cell_6t
Xbit_r57_c7 bl[7] br[7] wl[57] vdd gnd cell_6t
Xbit_r58_c7 bl[7] br[7] wl[58] vdd gnd cell_6t
Xbit_r59_c7 bl[7] br[7] wl[59] vdd gnd cell_6t
Xbit_r60_c7 bl[7] br[7] wl[60] vdd gnd cell_6t
Xbit_r61_c7 bl[7] br[7] wl[61] vdd gnd cell_6t
Xbit_r62_c7 bl[7] br[7] wl[62] vdd gnd cell_6t
Xbit_r63_c7 bl[7] br[7] wl[63] vdd gnd cell_6t
Xbit_r64_c7 bl[7] br[7] wl[64] vdd gnd cell_6t
Xbit_r65_c7 bl[7] br[7] wl[65] vdd gnd cell_6t
Xbit_r66_c7 bl[7] br[7] wl[66] vdd gnd cell_6t
Xbit_r67_c7 bl[7] br[7] wl[67] vdd gnd cell_6t
Xbit_r68_c7 bl[7] br[7] wl[68] vdd gnd cell_6t
Xbit_r69_c7 bl[7] br[7] wl[69] vdd gnd cell_6t
Xbit_r70_c7 bl[7] br[7] wl[70] vdd gnd cell_6t
Xbit_r71_c7 bl[7] br[7] wl[71] vdd gnd cell_6t
Xbit_r72_c7 bl[7] br[7] wl[72] vdd gnd cell_6t
Xbit_r73_c7 bl[7] br[7] wl[73] vdd gnd cell_6t
Xbit_r74_c7 bl[7] br[7] wl[74] vdd gnd cell_6t
Xbit_r75_c7 bl[7] br[7] wl[75] vdd gnd cell_6t
Xbit_r76_c7 bl[7] br[7] wl[76] vdd gnd cell_6t
Xbit_r77_c7 bl[7] br[7] wl[77] vdd gnd cell_6t
Xbit_r78_c7 bl[7] br[7] wl[78] vdd gnd cell_6t
Xbit_r79_c7 bl[7] br[7] wl[79] vdd gnd cell_6t
Xbit_r80_c7 bl[7] br[7] wl[80] vdd gnd cell_6t
Xbit_r81_c7 bl[7] br[7] wl[81] vdd gnd cell_6t
Xbit_r82_c7 bl[7] br[7] wl[82] vdd gnd cell_6t
Xbit_r83_c7 bl[7] br[7] wl[83] vdd gnd cell_6t
Xbit_r84_c7 bl[7] br[7] wl[84] vdd gnd cell_6t
Xbit_r85_c7 bl[7] br[7] wl[85] vdd gnd cell_6t
Xbit_r86_c7 bl[7] br[7] wl[86] vdd gnd cell_6t
Xbit_r87_c7 bl[7] br[7] wl[87] vdd gnd cell_6t
Xbit_r88_c7 bl[7] br[7] wl[88] vdd gnd cell_6t
Xbit_r89_c7 bl[7] br[7] wl[89] vdd gnd cell_6t
Xbit_r90_c7 bl[7] br[7] wl[90] vdd gnd cell_6t
Xbit_r91_c7 bl[7] br[7] wl[91] vdd gnd cell_6t
Xbit_r92_c7 bl[7] br[7] wl[92] vdd gnd cell_6t
Xbit_r93_c7 bl[7] br[7] wl[93] vdd gnd cell_6t
Xbit_r94_c7 bl[7] br[7] wl[94] vdd gnd cell_6t
Xbit_r95_c7 bl[7] br[7] wl[95] vdd gnd cell_6t
Xbit_r96_c7 bl[7] br[7] wl[96] vdd gnd cell_6t
Xbit_r97_c7 bl[7] br[7] wl[97] vdd gnd cell_6t
Xbit_r98_c7 bl[7] br[7] wl[98] vdd gnd cell_6t
Xbit_r99_c7 bl[7] br[7] wl[99] vdd gnd cell_6t
Xbit_r100_c7 bl[7] br[7] wl[100] vdd gnd cell_6t
Xbit_r101_c7 bl[7] br[7] wl[101] vdd gnd cell_6t
Xbit_r102_c7 bl[7] br[7] wl[102] vdd gnd cell_6t
Xbit_r103_c7 bl[7] br[7] wl[103] vdd gnd cell_6t
Xbit_r104_c7 bl[7] br[7] wl[104] vdd gnd cell_6t
Xbit_r105_c7 bl[7] br[7] wl[105] vdd gnd cell_6t
Xbit_r106_c7 bl[7] br[7] wl[106] vdd gnd cell_6t
Xbit_r107_c7 bl[7] br[7] wl[107] vdd gnd cell_6t
Xbit_r108_c7 bl[7] br[7] wl[108] vdd gnd cell_6t
Xbit_r109_c7 bl[7] br[7] wl[109] vdd gnd cell_6t
Xbit_r110_c7 bl[7] br[7] wl[110] vdd gnd cell_6t
Xbit_r111_c7 bl[7] br[7] wl[111] vdd gnd cell_6t
Xbit_r112_c7 bl[7] br[7] wl[112] vdd gnd cell_6t
Xbit_r113_c7 bl[7] br[7] wl[113] vdd gnd cell_6t
Xbit_r114_c7 bl[7] br[7] wl[114] vdd gnd cell_6t
Xbit_r115_c7 bl[7] br[7] wl[115] vdd gnd cell_6t
Xbit_r116_c7 bl[7] br[7] wl[116] vdd gnd cell_6t
Xbit_r117_c7 bl[7] br[7] wl[117] vdd gnd cell_6t
Xbit_r118_c7 bl[7] br[7] wl[118] vdd gnd cell_6t
Xbit_r119_c7 bl[7] br[7] wl[119] vdd gnd cell_6t
Xbit_r120_c7 bl[7] br[7] wl[120] vdd gnd cell_6t
Xbit_r121_c7 bl[7] br[7] wl[121] vdd gnd cell_6t
Xbit_r122_c7 bl[7] br[7] wl[122] vdd gnd cell_6t
Xbit_r123_c7 bl[7] br[7] wl[123] vdd gnd cell_6t
Xbit_r124_c7 bl[7] br[7] wl[124] vdd gnd cell_6t
Xbit_r125_c7 bl[7] br[7] wl[125] vdd gnd cell_6t
Xbit_r126_c7 bl[7] br[7] wl[126] vdd gnd cell_6t
Xbit_r127_c7 bl[7] br[7] wl[127] vdd gnd cell_6t
Xbit_r0_c8 bl[8] br[8] wl[0] vdd gnd cell_6t
Xbit_r1_c8 bl[8] br[8] wl[1] vdd gnd cell_6t
Xbit_r2_c8 bl[8] br[8] wl[2] vdd gnd cell_6t
Xbit_r3_c8 bl[8] br[8] wl[3] vdd gnd cell_6t
Xbit_r4_c8 bl[8] br[8] wl[4] vdd gnd cell_6t
Xbit_r5_c8 bl[8] br[8] wl[5] vdd gnd cell_6t
Xbit_r6_c8 bl[8] br[8] wl[6] vdd gnd cell_6t
Xbit_r7_c8 bl[8] br[8] wl[7] vdd gnd cell_6t
Xbit_r8_c8 bl[8] br[8] wl[8] vdd gnd cell_6t
Xbit_r9_c8 bl[8] br[8] wl[9] vdd gnd cell_6t
Xbit_r10_c8 bl[8] br[8] wl[10] vdd gnd cell_6t
Xbit_r11_c8 bl[8] br[8] wl[11] vdd gnd cell_6t
Xbit_r12_c8 bl[8] br[8] wl[12] vdd gnd cell_6t
Xbit_r13_c8 bl[8] br[8] wl[13] vdd gnd cell_6t
Xbit_r14_c8 bl[8] br[8] wl[14] vdd gnd cell_6t
Xbit_r15_c8 bl[8] br[8] wl[15] vdd gnd cell_6t
Xbit_r16_c8 bl[8] br[8] wl[16] vdd gnd cell_6t
Xbit_r17_c8 bl[8] br[8] wl[17] vdd gnd cell_6t
Xbit_r18_c8 bl[8] br[8] wl[18] vdd gnd cell_6t
Xbit_r19_c8 bl[8] br[8] wl[19] vdd gnd cell_6t
Xbit_r20_c8 bl[8] br[8] wl[20] vdd gnd cell_6t
Xbit_r21_c8 bl[8] br[8] wl[21] vdd gnd cell_6t
Xbit_r22_c8 bl[8] br[8] wl[22] vdd gnd cell_6t
Xbit_r23_c8 bl[8] br[8] wl[23] vdd gnd cell_6t
Xbit_r24_c8 bl[8] br[8] wl[24] vdd gnd cell_6t
Xbit_r25_c8 bl[8] br[8] wl[25] vdd gnd cell_6t
Xbit_r26_c8 bl[8] br[8] wl[26] vdd gnd cell_6t
Xbit_r27_c8 bl[8] br[8] wl[27] vdd gnd cell_6t
Xbit_r28_c8 bl[8] br[8] wl[28] vdd gnd cell_6t
Xbit_r29_c8 bl[8] br[8] wl[29] vdd gnd cell_6t
Xbit_r30_c8 bl[8] br[8] wl[30] vdd gnd cell_6t
Xbit_r31_c8 bl[8] br[8] wl[31] vdd gnd cell_6t
Xbit_r32_c8 bl[8] br[8] wl[32] vdd gnd cell_6t
Xbit_r33_c8 bl[8] br[8] wl[33] vdd gnd cell_6t
Xbit_r34_c8 bl[8] br[8] wl[34] vdd gnd cell_6t
Xbit_r35_c8 bl[8] br[8] wl[35] vdd gnd cell_6t
Xbit_r36_c8 bl[8] br[8] wl[36] vdd gnd cell_6t
Xbit_r37_c8 bl[8] br[8] wl[37] vdd gnd cell_6t
Xbit_r38_c8 bl[8] br[8] wl[38] vdd gnd cell_6t
Xbit_r39_c8 bl[8] br[8] wl[39] vdd gnd cell_6t
Xbit_r40_c8 bl[8] br[8] wl[40] vdd gnd cell_6t
Xbit_r41_c8 bl[8] br[8] wl[41] vdd gnd cell_6t
Xbit_r42_c8 bl[8] br[8] wl[42] vdd gnd cell_6t
Xbit_r43_c8 bl[8] br[8] wl[43] vdd gnd cell_6t
Xbit_r44_c8 bl[8] br[8] wl[44] vdd gnd cell_6t
Xbit_r45_c8 bl[8] br[8] wl[45] vdd gnd cell_6t
Xbit_r46_c8 bl[8] br[8] wl[46] vdd gnd cell_6t
Xbit_r47_c8 bl[8] br[8] wl[47] vdd gnd cell_6t
Xbit_r48_c8 bl[8] br[8] wl[48] vdd gnd cell_6t
Xbit_r49_c8 bl[8] br[8] wl[49] vdd gnd cell_6t
Xbit_r50_c8 bl[8] br[8] wl[50] vdd gnd cell_6t
Xbit_r51_c8 bl[8] br[8] wl[51] vdd gnd cell_6t
Xbit_r52_c8 bl[8] br[8] wl[52] vdd gnd cell_6t
Xbit_r53_c8 bl[8] br[8] wl[53] vdd gnd cell_6t
Xbit_r54_c8 bl[8] br[8] wl[54] vdd gnd cell_6t
Xbit_r55_c8 bl[8] br[8] wl[55] vdd gnd cell_6t
Xbit_r56_c8 bl[8] br[8] wl[56] vdd gnd cell_6t
Xbit_r57_c8 bl[8] br[8] wl[57] vdd gnd cell_6t
Xbit_r58_c8 bl[8] br[8] wl[58] vdd gnd cell_6t
Xbit_r59_c8 bl[8] br[8] wl[59] vdd gnd cell_6t
Xbit_r60_c8 bl[8] br[8] wl[60] vdd gnd cell_6t
Xbit_r61_c8 bl[8] br[8] wl[61] vdd gnd cell_6t
Xbit_r62_c8 bl[8] br[8] wl[62] vdd gnd cell_6t
Xbit_r63_c8 bl[8] br[8] wl[63] vdd gnd cell_6t
Xbit_r64_c8 bl[8] br[8] wl[64] vdd gnd cell_6t
Xbit_r65_c8 bl[8] br[8] wl[65] vdd gnd cell_6t
Xbit_r66_c8 bl[8] br[8] wl[66] vdd gnd cell_6t
Xbit_r67_c8 bl[8] br[8] wl[67] vdd gnd cell_6t
Xbit_r68_c8 bl[8] br[8] wl[68] vdd gnd cell_6t
Xbit_r69_c8 bl[8] br[8] wl[69] vdd gnd cell_6t
Xbit_r70_c8 bl[8] br[8] wl[70] vdd gnd cell_6t
Xbit_r71_c8 bl[8] br[8] wl[71] vdd gnd cell_6t
Xbit_r72_c8 bl[8] br[8] wl[72] vdd gnd cell_6t
Xbit_r73_c8 bl[8] br[8] wl[73] vdd gnd cell_6t
Xbit_r74_c8 bl[8] br[8] wl[74] vdd gnd cell_6t
Xbit_r75_c8 bl[8] br[8] wl[75] vdd gnd cell_6t
Xbit_r76_c8 bl[8] br[8] wl[76] vdd gnd cell_6t
Xbit_r77_c8 bl[8] br[8] wl[77] vdd gnd cell_6t
Xbit_r78_c8 bl[8] br[8] wl[78] vdd gnd cell_6t
Xbit_r79_c8 bl[8] br[8] wl[79] vdd gnd cell_6t
Xbit_r80_c8 bl[8] br[8] wl[80] vdd gnd cell_6t
Xbit_r81_c8 bl[8] br[8] wl[81] vdd gnd cell_6t
Xbit_r82_c8 bl[8] br[8] wl[82] vdd gnd cell_6t
Xbit_r83_c8 bl[8] br[8] wl[83] vdd gnd cell_6t
Xbit_r84_c8 bl[8] br[8] wl[84] vdd gnd cell_6t
Xbit_r85_c8 bl[8] br[8] wl[85] vdd gnd cell_6t
Xbit_r86_c8 bl[8] br[8] wl[86] vdd gnd cell_6t
Xbit_r87_c8 bl[8] br[8] wl[87] vdd gnd cell_6t
Xbit_r88_c8 bl[8] br[8] wl[88] vdd gnd cell_6t
Xbit_r89_c8 bl[8] br[8] wl[89] vdd gnd cell_6t
Xbit_r90_c8 bl[8] br[8] wl[90] vdd gnd cell_6t
Xbit_r91_c8 bl[8] br[8] wl[91] vdd gnd cell_6t
Xbit_r92_c8 bl[8] br[8] wl[92] vdd gnd cell_6t
Xbit_r93_c8 bl[8] br[8] wl[93] vdd gnd cell_6t
Xbit_r94_c8 bl[8] br[8] wl[94] vdd gnd cell_6t
Xbit_r95_c8 bl[8] br[8] wl[95] vdd gnd cell_6t
Xbit_r96_c8 bl[8] br[8] wl[96] vdd gnd cell_6t
Xbit_r97_c8 bl[8] br[8] wl[97] vdd gnd cell_6t
Xbit_r98_c8 bl[8] br[8] wl[98] vdd gnd cell_6t
Xbit_r99_c8 bl[8] br[8] wl[99] vdd gnd cell_6t
Xbit_r100_c8 bl[8] br[8] wl[100] vdd gnd cell_6t
Xbit_r101_c8 bl[8] br[8] wl[101] vdd gnd cell_6t
Xbit_r102_c8 bl[8] br[8] wl[102] vdd gnd cell_6t
Xbit_r103_c8 bl[8] br[8] wl[103] vdd gnd cell_6t
Xbit_r104_c8 bl[8] br[8] wl[104] vdd gnd cell_6t
Xbit_r105_c8 bl[8] br[8] wl[105] vdd gnd cell_6t
Xbit_r106_c8 bl[8] br[8] wl[106] vdd gnd cell_6t
Xbit_r107_c8 bl[8] br[8] wl[107] vdd gnd cell_6t
Xbit_r108_c8 bl[8] br[8] wl[108] vdd gnd cell_6t
Xbit_r109_c8 bl[8] br[8] wl[109] vdd gnd cell_6t
Xbit_r110_c8 bl[8] br[8] wl[110] vdd gnd cell_6t
Xbit_r111_c8 bl[8] br[8] wl[111] vdd gnd cell_6t
Xbit_r112_c8 bl[8] br[8] wl[112] vdd gnd cell_6t
Xbit_r113_c8 bl[8] br[8] wl[113] vdd gnd cell_6t
Xbit_r114_c8 bl[8] br[8] wl[114] vdd gnd cell_6t
Xbit_r115_c8 bl[8] br[8] wl[115] vdd gnd cell_6t
Xbit_r116_c8 bl[8] br[8] wl[116] vdd gnd cell_6t
Xbit_r117_c8 bl[8] br[8] wl[117] vdd gnd cell_6t
Xbit_r118_c8 bl[8] br[8] wl[118] vdd gnd cell_6t
Xbit_r119_c8 bl[8] br[8] wl[119] vdd gnd cell_6t
Xbit_r120_c8 bl[8] br[8] wl[120] vdd gnd cell_6t
Xbit_r121_c8 bl[8] br[8] wl[121] vdd gnd cell_6t
Xbit_r122_c8 bl[8] br[8] wl[122] vdd gnd cell_6t
Xbit_r123_c8 bl[8] br[8] wl[123] vdd gnd cell_6t
Xbit_r124_c8 bl[8] br[8] wl[124] vdd gnd cell_6t
Xbit_r125_c8 bl[8] br[8] wl[125] vdd gnd cell_6t
Xbit_r126_c8 bl[8] br[8] wl[126] vdd gnd cell_6t
Xbit_r127_c8 bl[8] br[8] wl[127] vdd gnd cell_6t
Xbit_r0_c9 bl[9] br[9] wl[0] vdd gnd cell_6t
Xbit_r1_c9 bl[9] br[9] wl[1] vdd gnd cell_6t
Xbit_r2_c9 bl[9] br[9] wl[2] vdd gnd cell_6t
Xbit_r3_c9 bl[9] br[9] wl[3] vdd gnd cell_6t
Xbit_r4_c9 bl[9] br[9] wl[4] vdd gnd cell_6t
Xbit_r5_c9 bl[9] br[9] wl[5] vdd gnd cell_6t
Xbit_r6_c9 bl[9] br[9] wl[6] vdd gnd cell_6t
Xbit_r7_c9 bl[9] br[9] wl[7] vdd gnd cell_6t
Xbit_r8_c9 bl[9] br[9] wl[8] vdd gnd cell_6t
Xbit_r9_c9 bl[9] br[9] wl[9] vdd gnd cell_6t
Xbit_r10_c9 bl[9] br[9] wl[10] vdd gnd cell_6t
Xbit_r11_c9 bl[9] br[9] wl[11] vdd gnd cell_6t
Xbit_r12_c9 bl[9] br[9] wl[12] vdd gnd cell_6t
Xbit_r13_c9 bl[9] br[9] wl[13] vdd gnd cell_6t
Xbit_r14_c9 bl[9] br[9] wl[14] vdd gnd cell_6t
Xbit_r15_c9 bl[9] br[9] wl[15] vdd gnd cell_6t
Xbit_r16_c9 bl[9] br[9] wl[16] vdd gnd cell_6t
Xbit_r17_c9 bl[9] br[9] wl[17] vdd gnd cell_6t
Xbit_r18_c9 bl[9] br[9] wl[18] vdd gnd cell_6t
Xbit_r19_c9 bl[9] br[9] wl[19] vdd gnd cell_6t
Xbit_r20_c9 bl[9] br[9] wl[20] vdd gnd cell_6t
Xbit_r21_c9 bl[9] br[9] wl[21] vdd gnd cell_6t
Xbit_r22_c9 bl[9] br[9] wl[22] vdd gnd cell_6t
Xbit_r23_c9 bl[9] br[9] wl[23] vdd gnd cell_6t
Xbit_r24_c9 bl[9] br[9] wl[24] vdd gnd cell_6t
Xbit_r25_c9 bl[9] br[9] wl[25] vdd gnd cell_6t
Xbit_r26_c9 bl[9] br[9] wl[26] vdd gnd cell_6t
Xbit_r27_c9 bl[9] br[9] wl[27] vdd gnd cell_6t
Xbit_r28_c9 bl[9] br[9] wl[28] vdd gnd cell_6t
Xbit_r29_c9 bl[9] br[9] wl[29] vdd gnd cell_6t
Xbit_r30_c9 bl[9] br[9] wl[30] vdd gnd cell_6t
Xbit_r31_c9 bl[9] br[9] wl[31] vdd gnd cell_6t
Xbit_r32_c9 bl[9] br[9] wl[32] vdd gnd cell_6t
Xbit_r33_c9 bl[9] br[9] wl[33] vdd gnd cell_6t
Xbit_r34_c9 bl[9] br[9] wl[34] vdd gnd cell_6t
Xbit_r35_c9 bl[9] br[9] wl[35] vdd gnd cell_6t
Xbit_r36_c9 bl[9] br[9] wl[36] vdd gnd cell_6t
Xbit_r37_c9 bl[9] br[9] wl[37] vdd gnd cell_6t
Xbit_r38_c9 bl[9] br[9] wl[38] vdd gnd cell_6t
Xbit_r39_c9 bl[9] br[9] wl[39] vdd gnd cell_6t
Xbit_r40_c9 bl[9] br[9] wl[40] vdd gnd cell_6t
Xbit_r41_c9 bl[9] br[9] wl[41] vdd gnd cell_6t
Xbit_r42_c9 bl[9] br[9] wl[42] vdd gnd cell_6t
Xbit_r43_c9 bl[9] br[9] wl[43] vdd gnd cell_6t
Xbit_r44_c9 bl[9] br[9] wl[44] vdd gnd cell_6t
Xbit_r45_c9 bl[9] br[9] wl[45] vdd gnd cell_6t
Xbit_r46_c9 bl[9] br[9] wl[46] vdd gnd cell_6t
Xbit_r47_c9 bl[9] br[9] wl[47] vdd gnd cell_6t
Xbit_r48_c9 bl[9] br[9] wl[48] vdd gnd cell_6t
Xbit_r49_c9 bl[9] br[9] wl[49] vdd gnd cell_6t
Xbit_r50_c9 bl[9] br[9] wl[50] vdd gnd cell_6t
Xbit_r51_c9 bl[9] br[9] wl[51] vdd gnd cell_6t
Xbit_r52_c9 bl[9] br[9] wl[52] vdd gnd cell_6t
Xbit_r53_c9 bl[9] br[9] wl[53] vdd gnd cell_6t
Xbit_r54_c9 bl[9] br[9] wl[54] vdd gnd cell_6t
Xbit_r55_c9 bl[9] br[9] wl[55] vdd gnd cell_6t
Xbit_r56_c9 bl[9] br[9] wl[56] vdd gnd cell_6t
Xbit_r57_c9 bl[9] br[9] wl[57] vdd gnd cell_6t
Xbit_r58_c9 bl[9] br[9] wl[58] vdd gnd cell_6t
Xbit_r59_c9 bl[9] br[9] wl[59] vdd gnd cell_6t
Xbit_r60_c9 bl[9] br[9] wl[60] vdd gnd cell_6t
Xbit_r61_c9 bl[9] br[9] wl[61] vdd gnd cell_6t
Xbit_r62_c9 bl[9] br[9] wl[62] vdd gnd cell_6t
Xbit_r63_c9 bl[9] br[9] wl[63] vdd gnd cell_6t
Xbit_r64_c9 bl[9] br[9] wl[64] vdd gnd cell_6t
Xbit_r65_c9 bl[9] br[9] wl[65] vdd gnd cell_6t
Xbit_r66_c9 bl[9] br[9] wl[66] vdd gnd cell_6t
Xbit_r67_c9 bl[9] br[9] wl[67] vdd gnd cell_6t
Xbit_r68_c9 bl[9] br[9] wl[68] vdd gnd cell_6t
Xbit_r69_c9 bl[9] br[9] wl[69] vdd gnd cell_6t
Xbit_r70_c9 bl[9] br[9] wl[70] vdd gnd cell_6t
Xbit_r71_c9 bl[9] br[9] wl[71] vdd gnd cell_6t
Xbit_r72_c9 bl[9] br[9] wl[72] vdd gnd cell_6t
Xbit_r73_c9 bl[9] br[9] wl[73] vdd gnd cell_6t
Xbit_r74_c9 bl[9] br[9] wl[74] vdd gnd cell_6t
Xbit_r75_c9 bl[9] br[9] wl[75] vdd gnd cell_6t
Xbit_r76_c9 bl[9] br[9] wl[76] vdd gnd cell_6t
Xbit_r77_c9 bl[9] br[9] wl[77] vdd gnd cell_6t
Xbit_r78_c9 bl[9] br[9] wl[78] vdd gnd cell_6t
Xbit_r79_c9 bl[9] br[9] wl[79] vdd gnd cell_6t
Xbit_r80_c9 bl[9] br[9] wl[80] vdd gnd cell_6t
Xbit_r81_c9 bl[9] br[9] wl[81] vdd gnd cell_6t
Xbit_r82_c9 bl[9] br[9] wl[82] vdd gnd cell_6t
Xbit_r83_c9 bl[9] br[9] wl[83] vdd gnd cell_6t
Xbit_r84_c9 bl[9] br[9] wl[84] vdd gnd cell_6t
Xbit_r85_c9 bl[9] br[9] wl[85] vdd gnd cell_6t
Xbit_r86_c9 bl[9] br[9] wl[86] vdd gnd cell_6t
Xbit_r87_c9 bl[9] br[9] wl[87] vdd gnd cell_6t
Xbit_r88_c9 bl[9] br[9] wl[88] vdd gnd cell_6t
Xbit_r89_c9 bl[9] br[9] wl[89] vdd gnd cell_6t
Xbit_r90_c9 bl[9] br[9] wl[90] vdd gnd cell_6t
Xbit_r91_c9 bl[9] br[9] wl[91] vdd gnd cell_6t
Xbit_r92_c9 bl[9] br[9] wl[92] vdd gnd cell_6t
Xbit_r93_c9 bl[9] br[9] wl[93] vdd gnd cell_6t
Xbit_r94_c9 bl[9] br[9] wl[94] vdd gnd cell_6t
Xbit_r95_c9 bl[9] br[9] wl[95] vdd gnd cell_6t
Xbit_r96_c9 bl[9] br[9] wl[96] vdd gnd cell_6t
Xbit_r97_c9 bl[9] br[9] wl[97] vdd gnd cell_6t
Xbit_r98_c9 bl[9] br[9] wl[98] vdd gnd cell_6t
Xbit_r99_c9 bl[9] br[9] wl[99] vdd gnd cell_6t
Xbit_r100_c9 bl[9] br[9] wl[100] vdd gnd cell_6t
Xbit_r101_c9 bl[9] br[9] wl[101] vdd gnd cell_6t
Xbit_r102_c9 bl[9] br[9] wl[102] vdd gnd cell_6t
Xbit_r103_c9 bl[9] br[9] wl[103] vdd gnd cell_6t
Xbit_r104_c9 bl[9] br[9] wl[104] vdd gnd cell_6t
Xbit_r105_c9 bl[9] br[9] wl[105] vdd gnd cell_6t
Xbit_r106_c9 bl[9] br[9] wl[106] vdd gnd cell_6t
Xbit_r107_c9 bl[9] br[9] wl[107] vdd gnd cell_6t
Xbit_r108_c9 bl[9] br[9] wl[108] vdd gnd cell_6t
Xbit_r109_c9 bl[9] br[9] wl[109] vdd gnd cell_6t
Xbit_r110_c9 bl[9] br[9] wl[110] vdd gnd cell_6t
Xbit_r111_c9 bl[9] br[9] wl[111] vdd gnd cell_6t
Xbit_r112_c9 bl[9] br[9] wl[112] vdd gnd cell_6t
Xbit_r113_c9 bl[9] br[9] wl[113] vdd gnd cell_6t
Xbit_r114_c9 bl[9] br[9] wl[114] vdd gnd cell_6t
Xbit_r115_c9 bl[9] br[9] wl[115] vdd gnd cell_6t
Xbit_r116_c9 bl[9] br[9] wl[116] vdd gnd cell_6t
Xbit_r117_c9 bl[9] br[9] wl[117] vdd gnd cell_6t
Xbit_r118_c9 bl[9] br[9] wl[118] vdd gnd cell_6t
Xbit_r119_c9 bl[9] br[9] wl[119] vdd gnd cell_6t
Xbit_r120_c9 bl[9] br[9] wl[120] vdd gnd cell_6t
Xbit_r121_c9 bl[9] br[9] wl[121] vdd gnd cell_6t
Xbit_r122_c9 bl[9] br[9] wl[122] vdd gnd cell_6t
Xbit_r123_c9 bl[9] br[9] wl[123] vdd gnd cell_6t
Xbit_r124_c9 bl[9] br[9] wl[124] vdd gnd cell_6t
Xbit_r125_c9 bl[9] br[9] wl[125] vdd gnd cell_6t
Xbit_r126_c9 bl[9] br[9] wl[126] vdd gnd cell_6t
Xbit_r127_c9 bl[9] br[9] wl[127] vdd gnd cell_6t
Xbit_r0_c10 bl[10] br[10] wl[0] vdd gnd cell_6t
Xbit_r1_c10 bl[10] br[10] wl[1] vdd gnd cell_6t
Xbit_r2_c10 bl[10] br[10] wl[2] vdd gnd cell_6t
Xbit_r3_c10 bl[10] br[10] wl[3] vdd gnd cell_6t
Xbit_r4_c10 bl[10] br[10] wl[4] vdd gnd cell_6t
Xbit_r5_c10 bl[10] br[10] wl[5] vdd gnd cell_6t
Xbit_r6_c10 bl[10] br[10] wl[6] vdd gnd cell_6t
Xbit_r7_c10 bl[10] br[10] wl[7] vdd gnd cell_6t
Xbit_r8_c10 bl[10] br[10] wl[8] vdd gnd cell_6t
Xbit_r9_c10 bl[10] br[10] wl[9] vdd gnd cell_6t
Xbit_r10_c10 bl[10] br[10] wl[10] vdd gnd cell_6t
Xbit_r11_c10 bl[10] br[10] wl[11] vdd gnd cell_6t
Xbit_r12_c10 bl[10] br[10] wl[12] vdd gnd cell_6t
Xbit_r13_c10 bl[10] br[10] wl[13] vdd gnd cell_6t
Xbit_r14_c10 bl[10] br[10] wl[14] vdd gnd cell_6t
Xbit_r15_c10 bl[10] br[10] wl[15] vdd gnd cell_6t
Xbit_r16_c10 bl[10] br[10] wl[16] vdd gnd cell_6t
Xbit_r17_c10 bl[10] br[10] wl[17] vdd gnd cell_6t
Xbit_r18_c10 bl[10] br[10] wl[18] vdd gnd cell_6t
Xbit_r19_c10 bl[10] br[10] wl[19] vdd gnd cell_6t
Xbit_r20_c10 bl[10] br[10] wl[20] vdd gnd cell_6t
Xbit_r21_c10 bl[10] br[10] wl[21] vdd gnd cell_6t
Xbit_r22_c10 bl[10] br[10] wl[22] vdd gnd cell_6t
Xbit_r23_c10 bl[10] br[10] wl[23] vdd gnd cell_6t
Xbit_r24_c10 bl[10] br[10] wl[24] vdd gnd cell_6t
Xbit_r25_c10 bl[10] br[10] wl[25] vdd gnd cell_6t
Xbit_r26_c10 bl[10] br[10] wl[26] vdd gnd cell_6t
Xbit_r27_c10 bl[10] br[10] wl[27] vdd gnd cell_6t
Xbit_r28_c10 bl[10] br[10] wl[28] vdd gnd cell_6t
Xbit_r29_c10 bl[10] br[10] wl[29] vdd gnd cell_6t
Xbit_r30_c10 bl[10] br[10] wl[30] vdd gnd cell_6t
Xbit_r31_c10 bl[10] br[10] wl[31] vdd gnd cell_6t
Xbit_r32_c10 bl[10] br[10] wl[32] vdd gnd cell_6t
Xbit_r33_c10 bl[10] br[10] wl[33] vdd gnd cell_6t
Xbit_r34_c10 bl[10] br[10] wl[34] vdd gnd cell_6t
Xbit_r35_c10 bl[10] br[10] wl[35] vdd gnd cell_6t
Xbit_r36_c10 bl[10] br[10] wl[36] vdd gnd cell_6t
Xbit_r37_c10 bl[10] br[10] wl[37] vdd gnd cell_6t
Xbit_r38_c10 bl[10] br[10] wl[38] vdd gnd cell_6t
Xbit_r39_c10 bl[10] br[10] wl[39] vdd gnd cell_6t
Xbit_r40_c10 bl[10] br[10] wl[40] vdd gnd cell_6t
Xbit_r41_c10 bl[10] br[10] wl[41] vdd gnd cell_6t
Xbit_r42_c10 bl[10] br[10] wl[42] vdd gnd cell_6t
Xbit_r43_c10 bl[10] br[10] wl[43] vdd gnd cell_6t
Xbit_r44_c10 bl[10] br[10] wl[44] vdd gnd cell_6t
Xbit_r45_c10 bl[10] br[10] wl[45] vdd gnd cell_6t
Xbit_r46_c10 bl[10] br[10] wl[46] vdd gnd cell_6t
Xbit_r47_c10 bl[10] br[10] wl[47] vdd gnd cell_6t
Xbit_r48_c10 bl[10] br[10] wl[48] vdd gnd cell_6t
Xbit_r49_c10 bl[10] br[10] wl[49] vdd gnd cell_6t
Xbit_r50_c10 bl[10] br[10] wl[50] vdd gnd cell_6t
Xbit_r51_c10 bl[10] br[10] wl[51] vdd gnd cell_6t
Xbit_r52_c10 bl[10] br[10] wl[52] vdd gnd cell_6t
Xbit_r53_c10 bl[10] br[10] wl[53] vdd gnd cell_6t
Xbit_r54_c10 bl[10] br[10] wl[54] vdd gnd cell_6t
Xbit_r55_c10 bl[10] br[10] wl[55] vdd gnd cell_6t
Xbit_r56_c10 bl[10] br[10] wl[56] vdd gnd cell_6t
Xbit_r57_c10 bl[10] br[10] wl[57] vdd gnd cell_6t
Xbit_r58_c10 bl[10] br[10] wl[58] vdd gnd cell_6t
Xbit_r59_c10 bl[10] br[10] wl[59] vdd gnd cell_6t
Xbit_r60_c10 bl[10] br[10] wl[60] vdd gnd cell_6t
Xbit_r61_c10 bl[10] br[10] wl[61] vdd gnd cell_6t
Xbit_r62_c10 bl[10] br[10] wl[62] vdd gnd cell_6t
Xbit_r63_c10 bl[10] br[10] wl[63] vdd gnd cell_6t
Xbit_r64_c10 bl[10] br[10] wl[64] vdd gnd cell_6t
Xbit_r65_c10 bl[10] br[10] wl[65] vdd gnd cell_6t
Xbit_r66_c10 bl[10] br[10] wl[66] vdd gnd cell_6t
Xbit_r67_c10 bl[10] br[10] wl[67] vdd gnd cell_6t
Xbit_r68_c10 bl[10] br[10] wl[68] vdd gnd cell_6t
Xbit_r69_c10 bl[10] br[10] wl[69] vdd gnd cell_6t
Xbit_r70_c10 bl[10] br[10] wl[70] vdd gnd cell_6t
Xbit_r71_c10 bl[10] br[10] wl[71] vdd gnd cell_6t
Xbit_r72_c10 bl[10] br[10] wl[72] vdd gnd cell_6t
Xbit_r73_c10 bl[10] br[10] wl[73] vdd gnd cell_6t
Xbit_r74_c10 bl[10] br[10] wl[74] vdd gnd cell_6t
Xbit_r75_c10 bl[10] br[10] wl[75] vdd gnd cell_6t
Xbit_r76_c10 bl[10] br[10] wl[76] vdd gnd cell_6t
Xbit_r77_c10 bl[10] br[10] wl[77] vdd gnd cell_6t
Xbit_r78_c10 bl[10] br[10] wl[78] vdd gnd cell_6t
Xbit_r79_c10 bl[10] br[10] wl[79] vdd gnd cell_6t
Xbit_r80_c10 bl[10] br[10] wl[80] vdd gnd cell_6t
Xbit_r81_c10 bl[10] br[10] wl[81] vdd gnd cell_6t
Xbit_r82_c10 bl[10] br[10] wl[82] vdd gnd cell_6t
Xbit_r83_c10 bl[10] br[10] wl[83] vdd gnd cell_6t
Xbit_r84_c10 bl[10] br[10] wl[84] vdd gnd cell_6t
Xbit_r85_c10 bl[10] br[10] wl[85] vdd gnd cell_6t
Xbit_r86_c10 bl[10] br[10] wl[86] vdd gnd cell_6t
Xbit_r87_c10 bl[10] br[10] wl[87] vdd gnd cell_6t
Xbit_r88_c10 bl[10] br[10] wl[88] vdd gnd cell_6t
Xbit_r89_c10 bl[10] br[10] wl[89] vdd gnd cell_6t
Xbit_r90_c10 bl[10] br[10] wl[90] vdd gnd cell_6t
Xbit_r91_c10 bl[10] br[10] wl[91] vdd gnd cell_6t
Xbit_r92_c10 bl[10] br[10] wl[92] vdd gnd cell_6t
Xbit_r93_c10 bl[10] br[10] wl[93] vdd gnd cell_6t
Xbit_r94_c10 bl[10] br[10] wl[94] vdd gnd cell_6t
Xbit_r95_c10 bl[10] br[10] wl[95] vdd gnd cell_6t
Xbit_r96_c10 bl[10] br[10] wl[96] vdd gnd cell_6t
Xbit_r97_c10 bl[10] br[10] wl[97] vdd gnd cell_6t
Xbit_r98_c10 bl[10] br[10] wl[98] vdd gnd cell_6t
Xbit_r99_c10 bl[10] br[10] wl[99] vdd gnd cell_6t
Xbit_r100_c10 bl[10] br[10] wl[100] vdd gnd cell_6t
Xbit_r101_c10 bl[10] br[10] wl[101] vdd gnd cell_6t
Xbit_r102_c10 bl[10] br[10] wl[102] vdd gnd cell_6t
Xbit_r103_c10 bl[10] br[10] wl[103] vdd gnd cell_6t
Xbit_r104_c10 bl[10] br[10] wl[104] vdd gnd cell_6t
Xbit_r105_c10 bl[10] br[10] wl[105] vdd gnd cell_6t
Xbit_r106_c10 bl[10] br[10] wl[106] vdd gnd cell_6t
Xbit_r107_c10 bl[10] br[10] wl[107] vdd gnd cell_6t
Xbit_r108_c10 bl[10] br[10] wl[108] vdd gnd cell_6t
Xbit_r109_c10 bl[10] br[10] wl[109] vdd gnd cell_6t
Xbit_r110_c10 bl[10] br[10] wl[110] vdd gnd cell_6t
Xbit_r111_c10 bl[10] br[10] wl[111] vdd gnd cell_6t
Xbit_r112_c10 bl[10] br[10] wl[112] vdd gnd cell_6t
Xbit_r113_c10 bl[10] br[10] wl[113] vdd gnd cell_6t
Xbit_r114_c10 bl[10] br[10] wl[114] vdd gnd cell_6t
Xbit_r115_c10 bl[10] br[10] wl[115] vdd gnd cell_6t
Xbit_r116_c10 bl[10] br[10] wl[116] vdd gnd cell_6t
Xbit_r117_c10 bl[10] br[10] wl[117] vdd gnd cell_6t
Xbit_r118_c10 bl[10] br[10] wl[118] vdd gnd cell_6t
Xbit_r119_c10 bl[10] br[10] wl[119] vdd gnd cell_6t
Xbit_r120_c10 bl[10] br[10] wl[120] vdd gnd cell_6t
Xbit_r121_c10 bl[10] br[10] wl[121] vdd gnd cell_6t
Xbit_r122_c10 bl[10] br[10] wl[122] vdd gnd cell_6t
Xbit_r123_c10 bl[10] br[10] wl[123] vdd gnd cell_6t
Xbit_r124_c10 bl[10] br[10] wl[124] vdd gnd cell_6t
Xbit_r125_c10 bl[10] br[10] wl[125] vdd gnd cell_6t
Xbit_r126_c10 bl[10] br[10] wl[126] vdd gnd cell_6t
Xbit_r127_c10 bl[10] br[10] wl[127] vdd gnd cell_6t
Xbit_r0_c11 bl[11] br[11] wl[0] vdd gnd cell_6t
Xbit_r1_c11 bl[11] br[11] wl[1] vdd gnd cell_6t
Xbit_r2_c11 bl[11] br[11] wl[2] vdd gnd cell_6t
Xbit_r3_c11 bl[11] br[11] wl[3] vdd gnd cell_6t
Xbit_r4_c11 bl[11] br[11] wl[4] vdd gnd cell_6t
Xbit_r5_c11 bl[11] br[11] wl[5] vdd gnd cell_6t
Xbit_r6_c11 bl[11] br[11] wl[6] vdd gnd cell_6t
Xbit_r7_c11 bl[11] br[11] wl[7] vdd gnd cell_6t
Xbit_r8_c11 bl[11] br[11] wl[8] vdd gnd cell_6t
Xbit_r9_c11 bl[11] br[11] wl[9] vdd gnd cell_6t
Xbit_r10_c11 bl[11] br[11] wl[10] vdd gnd cell_6t
Xbit_r11_c11 bl[11] br[11] wl[11] vdd gnd cell_6t
Xbit_r12_c11 bl[11] br[11] wl[12] vdd gnd cell_6t
Xbit_r13_c11 bl[11] br[11] wl[13] vdd gnd cell_6t
Xbit_r14_c11 bl[11] br[11] wl[14] vdd gnd cell_6t
Xbit_r15_c11 bl[11] br[11] wl[15] vdd gnd cell_6t
Xbit_r16_c11 bl[11] br[11] wl[16] vdd gnd cell_6t
Xbit_r17_c11 bl[11] br[11] wl[17] vdd gnd cell_6t
Xbit_r18_c11 bl[11] br[11] wl[18] vdd gnd cell_6t
Xbit_r19_c11 bl[11] br[11] wl[19] vdd gnd cell_6t
Xbit_r20_c11 bl[11] br[11] wl[20] vdd gnd cell_6t
Xbit_r21_c11 bl[11] br[11] wl[21] vdd gnd cell_6t
Xbit_r22_c11 bl[11] br[11] wl[22] vdd gnd cell_6t
Xbit_r23_c11 bl[11] br[11] wl[23] vdd gnd cell_6t
Xbit_r24_c11 bl[11] br[11] wl[24] vdd gnd cell_6t
Xbit_r25_c11 bl[11] br[11] wl[25] vdd gnd cell_6t
Xbit_r26_c11 bl[11] br[11] wl[26] vdd gnd cell_6t
Xbit_r27_c11 bl[11] br[11] wl[27] vdd gnd cell_6t
Xbit_r28_c11 bl[11] br[11] wl[28] vdd gnd cell_6t
Xbit_r29_c11 bl[11] br[11] wl[29] vdd gnd cell_6t
Xbit_r30_c11 bl[11] br[11] wl[30] vdd gnd cell_6t
Xbit_r31_c11 bl[11] br[11] wl[31] vdd gnd cell_6t
Xbit_r32_c11 bl[11] br[11] wl[32] vdd gnd cell_6t
Xbit_r33_c11 bl[11] br[11] wl[33] vdd gnd cell_6t
Xbit_r34_c11 bl[11] br[11] wl[34] vdd gnd cell_6t
Xbit_r35_c11 bl[11] br[11] wl[35] vdd gnd cell_6t
Xbit_r36_c11 bl[11] br[11] wl[36] vdd gnd cell_6t
Xbit_r37_c11 bl[11] br[11] wl[37] vdd gnd cell_6t
Xbit_r38_c11 bl[11] br[11] wl[38] vdd gnd cell_6t
Xbit_r39_c11 bl[11] br[11] wl[39] vdd gnd cell_6t
Xbit_r40_c11 bl[11] br[11] wl[40] vdd gnd cell_6t
Xbit_r41_c11 bl[11] br[11] wl[41] vdd gnd cell_6t
Xbit_r42_c11 bl[11] br[11] wl[42] vdd gnd cell_6t
Xbit_r43_c11 bl[11] br[11] wl[43] vdd gnd cell_6t
Xbit_r44_c11 bl[11] br[11] wl[44] vdd gnd cell_6t
Xbit_r45_c11 bl[11] br[11] wl[45] vdd gnd cell_6t
Xbit_r46_c11 bl[11] br[11] wl[46] vdd gnd cell_6t
Xbit_r47_c11 bl[11] br[11] wl[47] vdd gnd cell_6t
Xbit_r48_c11 bl[11] br[11] wl[48] vdd gnd cell_6t
Xbit_r49_c11 bl[11] br[11] wl[49] vdd gnd cell_6t
Xbit_r50_c11 bl[11] br[11] wl[50] vdd gnd cell_6t
Xbit_r51_c11 bl[11] br[11] wl[51] vdd gnd cell_6t
Xbit_r52_c11 bl[11] br[11] wl[52] vdd gnd cell_6t
Xbit_r53_c11 bl[11] br[11] wl[53] vdd gnd cell_6t
Xbit_r54_c11 bl[11] br[11] wl[54] vdd gnd cell_6t
Xbit_r55_c11 bl[11] br[11] wl[55] vdd gnd cell_6t
Xbit_r56_c11 bl[11] br[11] wl[56] vdd gnd cell_6t
Xbit_r57_c11 bl[11] br[11] wl[57] vdd gnd cell_6t
Xbit_r58_c11 bl[11] br[11] wl[58] vdd gnd cell_6t
Xbit_r59_c11 bl[11] br[11] wl[59] vdd gnd cell_6t
Xbit_r60_c11 bl[11] br[11] wl[60] vdd gnd cell_6t
Xbit_r61_c11 bl[11] br[11] wl[61] vdd gnd cell_6t
Xbit_r62_c11 bl[11] br[11] wl[62] vdd gnd cell_6t
Xbit_r63_c11 bl[11] br[11] wl[63] vdd gnd cell_6t
Xbit_r64_c11 bl[11] br[11] wl[64] vdd gnd cell_6t
Xbit_r65_c11 bl[11] br[11] wl[65] vdd gnd cell_6t
Xbit_r66_c11 bl[11] br[11] wl[66] vdd gnd cell_6t
Xbit_r67_c11 bl[11] br[11] wl[67] vdd gnd cell_6t
Xbit_r68_c11 bl[11] br[11] wl[68] vdd gnd cell_6t
Xbit_r69_c11 bl[11] br[11] wl[69] vdd gnd cell_6t
Xbit_r70_c11 bl[11] br[11] wl[70] vdd gnd cell_6t
Xbit_r71_c11 bl[11] br[11] wl[71] vdd gnd cell_6t
Xbit_r72_c11 bl[11] br[11] wl[72] vdd gnd cell_6t
Xbit_r73_c11 bl[11] br[11] wl[73] vdd gnd cell_6t
Xbit_r74_c11 bl[11] br[11] wl[74] vdd gnd cell_6t
Xbit_r75_c11 bl[11] br[11] wl[75] vdd gnd cell_6t
Xbit_r76_c11 bl[11] br[11] wl[76] vdd gnd cell_6t
Xbit_r77_c11 bl[11] br[11] wl[77] vdd gnd cell_6t
Xbit_r78_c11 bl[11] br[11] wl[78] vdd gnd cell_6t
Xbit_r79_c11 bl[11] br[11] wl[79] vdd gnd cell_6t
Xbit_r80_c11 bl[11] br[11] wl[80] vdd gnd cell_6t
Xbit_r81_c11 bl[11] br[11] wl[81] vdd gnd cell_6t
Xbit_r82_c11 bl[11] br[11] wl[82] vdd gnd cell_6t
Xbit_r83_c11 bl[11] br[11] wl[83] vdd gnd cell_6t
Xbit_r84_c11 bl[11] br[11] wl[84] vdd gnd cell_6t
Xbit_r85_c11 bl[11] br[11] wl[85] vdd gnd cell_6t
Xbit_r86_c11 bl[11] br[11] wl[86] vdd gnd cell_6t
Xbit_r87_c11 bl[11] br[11] wl[87] vdd gnd cell_6t
Xbit_r88_c11 bl[11] br[11] wl[88] vdd gnd cell_6t
Xbit_r89_c11 bl[11] br[11] wl[89] vdd gnd cell_6t
Xbit_r90_c11 bl[11] br[11] wl[90] vdd gnd cell_6t
Xbit_r91_c11 bl[11] br[11] wl[91] vdd gnd cell_6t
Xbit_r92_c11 bl[11] br[11] wl[92] vdd gnd cell_6t
Xbit_r93_c11 bl[11] br[11] wl[93] vdd gnd cell_6t
Xbit_r94_c11 bl[11] br[11] wl[94] vdd gnd cell_6t
Xbit_r95_c11 bl[11] br[11] wl[95] vdd gnd cell_6t
Xbit_r96_c11 bl[11] br[11] wl[96] vdd gnd cell_6t
Xbit_r97_c11 bl[11] br[11] wl[97] vdd gnd cell_6t
Xbit_r98_c11 bl[11] br[11] wl[98] vdd gnd cell_6t
Xbit_r99_c11 bl[11] br[11] wl[99] vdd gnd cell_6t
Xbit_r100_c11 bl[11] br[11] wl[100] vdd gnd cell_6t
Xbit_r101_c11 bl[11] br[11] wl[101] vdd gnd cell_6t
Xbit_r102_c11 bl[11] br[11] wl[102] vdd gnd cell_6t
Xbit_r103_c11 bl[11] br[11] wl[103] vdd gnd cell_6t
Xbit_r104_c11 bl[11] br[11] wl[104] vdd gnd cell_6t
Xbit_r105_c11 bl[11] br[11] wl[105] vdd gnd cell_6t
Xbit_r106_c11 bl[11] br[11] wl[106] vdd gnd cell_6t
Xbit_r107_c11 bl[11] br[11] wl[107] vdd gnd cell_6t
Xbit_r108_c11 bl[11] br[11] wl[108] vdd gnd cell_6t
Xbit_r109_c11 bl[11] br[11] wl[109] vdd gnd cell_6t
Xbit_r110_c11 bl[11] br[11] wl[110] vdd gnd cell_6t
Xbit_r111_c11 bl[11] br[11] wl[111] vdd gnd cell_6t
Xbit_r112_c11 bl[11] br[11] wl[112] vdd gnd cell_6t
Xbit_r113_c11 bl[11] br[11] wl[113] vdd gnd cell_6t
Xbit_r114_c11 bl[11] br[11] wl[114] vdd gnd cell_6t
Xbit_r115_c11 bl[11] br[11] wl[115] vdd gnd cell_6t
Xbit_r116_c11 bl[11] br[11] wl[116] vdd gnd cell_6t
Xbit_r117_c11 bl[11] br[11] wl[117] vdd gnd cell_6t
Xbit_r118_c11 bl[11] br[11] wl[118] vdd gnd cell_6t
Xbit_r119_c11 bl[11] br[11] wl[119] vdd gnd cell_6t
Xbit_r120_c11 bl[11] br[11] wl[120] vdd gnd cell_6t
Xbit_r121_c11 bl[11] br[11] wl[121] vdd gnd cell_6t
Xbit_r122_c11 bl[11] br[11] wl[122] vdd gnd cell_6t
Xbit_r123_c11 bl[11] br[11] wl[123] vdd gnd cell_6t
Xbit_r124_c11 bl[11] br[11] wl[124] vdd gnd cell_6t
Xbit_r125_c11 bl[11] br[11] wl[125] vdd gnd cell_6t
Xbit_r126_c11 bl[11] br[11] wl[126] vdd gnd cell_6t
Xbit_r127_c11 bl[11] br[11] wl[127] vdd gnd cell_6t
Xbit_r0_c12 bl[12] br[12] wl[0] vdd gnd cell_6t
Xbit_r1_c12 bl[12] br[12] wl[1] vdd gnd cell_6t
Xbit_r2_c12 bl[12] br[12] wl[2] vdd gnd cell_6t
Xbit_r3_c12 bl[12] br[12] wl[3] vdd gnd cell_6t
Xbit_r4_c12 bl[12] br[12] wl[4] vdd gnd cell_6t
Xbit_r5_c12 bl[12] br[12] wl[5] vdd gnd cell_6t
Xbit_r6_c12 bl[12] br[12] wl[6] vdd gnd cell_6t
Xbit_r7_c12 bl[12] br[12] wl[7] vdd gnd cell_6t
Xbit_r8_c12 bl[12] br[12] wl[8] vdd gnd cell_6t
Xbit_r9_c12 bl[12] br[12] wl[9] vdd gnd cell_6t
Xbit_r10_c12 bl[12] br[12] wl[10] vdd gnd cell_6t
Xbit_r11_c12 bl[12] br[12] wl[11] vdd gnd cell_6t
Xbit_r12_c12 bl[12] br[12] wl[12] vdd gnd cell_6t
Xbit_r13_c12 bl[12] br[12] wl[13] vdd gnd cell_6t
Xbit_r14_c12 bl[12] br[12] wl[14] vdd gnd cell_6t
Xbit_r15_c12 bl[12] br[12] wl[15] vdd gnd cell_6t
Xbit_r16_c12 bl[12] br[12] wl[16] vdd gnd cell_6t
Xbit_r17_c12 bl[12] br[12] wl[17] vdd gnd cell_6t
Xbit_r18_c12 bl[12] br[12] wl[18] vdd gnd cell_6t
Xbit_r19_c12 bl[12] br[12] wl[19] vdd gnd cell_6t
Xbit_r20_c12 bl[12] br[12] wl[20] vdd gnd cell_6t
Xbit_r21_c12 bl[12] br[12] wl[21] vdd gnd cell_6t
Xbit_r22_c12 bl[12] br[12] wl[22] vdd gnd cell_6t
Xbit_r23_c12 bl[12] br[12] wl[23] vdd gnd cell_6t
Xbit_r24_c12 bl[12] br[12] wl[24] vdd gnd cell_6t
Xbit_r25_c12 bl[12] br[12] wl[25] vdd gnd cell_6t
Xbit_r26_c12 bl[12] br[12] wl[26] vdd gnd cell_6t
Xbit_r27_c12 bl[12] br[12] wl[27] vdd gnd cell_6t
Xbit_r28_c12 bl[12] br[12] wl[28] vdd gnd cell_6t
Xbit_r29_c12 bl[12] br[12] wl[29] vdd gnd cell_6t
Xbit_r30_c12 bl[12] br[12] wl[30] vdd gnd cell_6t
Xbit_r31_c12 bl[12] br[12] wl[31] vdd gnd cell_6t
Xbit_r32_c12 bl[12] br[12] wl[32] vdd gnd cell_6t
Xbit_r33_c12 bl[12] br[12] wl[33] vdd gnd cell_6t
Xbit_r34_c12 bl[12] br[12] wl[34] vdd gnd cell_6t
Xbit_r35_c12 bl[12] br[12] wl[35] vdd gnd cell_6t
Xbit_r36_c12 bl[12] br[12] wl[36] vdd gnd cell_6t
Xbit_r37_c12 bl[12] br[12] wl[37] vdd gnd cell_6t
Xbit_r38_c12 bl[12] br[12] wl[38] vdd gnd cell_6t
Xbit_r39_c12 bl[12] br[12] wl[39] vdd gnd cell_6t
Xbit_r40_c12 bl[12] br[12] wl[40] vdd gnd cell_6t
Xbit_r41_c12 bl[12] br[12] wl[41] vdd gnd cell_6t
Xbit_r42_c12 bl[12] br[12] wl[42] vdd gnd cell_6t
Xbit_r43_c12 bl[12] br[12] wl[43] vdd gnd cell_6t
Xbit_r44_c12 bl[12] br[12] wl[44] vdd gnd cell_6t
Xbit_r45_c12 bl[12] br[12] wl[45] vdd gnd cell_6t
Xbit_r46_c12 bl[12] br[12] wl[46] vdd gnd cell_6t
Xbit_r47_c12 bl[12] br[12] wl[47] vdd gnd cell_6t
Xbit_r48_c12 bl[12] br[12] wl[48] vdd gnd cell_6t
Xbit_r49_c12 bl[12] br[12] wl[49] vdd gnd cell_6t
Xbit_r50_c12 bl[12] br[12] wl[50] vdd gnd cell_6t
Xbit_r51_c12 bl[12] br[12] wl[51] vdd gnd cell_6t
Xbit_r52_c12 bl[12] br[12] wl[52] vdd gnd cell_6t
Xbit_r53_c12 bl[12] br[12] wl[53] vdd gnd cell_6t
Xbit_r54_c12 bl[12] br[12] wl[54] vdd gnd cell_6t
Xbit_r55_c12 bl[12] br[12] wl[55] vdd gnd cell_6t
Xbit_r56_c12 bl[12] br[12] wl[56] vdd gnd cell_6t
Xbit_r57_c12 bl[12] br[12] wl[57] vdd gnd cell_6t
Xbit_r58_c12 bl[12] br[12] wl[58] vdd gnd cell_6t
Xbit_r59_c12 bl[12] br[12] wl[59] vdd gnd cell_6t
Xbit_r60_c12 bl[12] br[12] wl[60] vdd gnd cell_6t
Xbit_r61_c12 bl[12] br[12] wl[61] vdd gnd cell_6t
Xbit_r62_c12 bl[12] br[12] wl[62] vdd gnd cell_6t
Xbit_r63_c12 bl[12] br[12] wl[63] vdd gnd cell_6t
Xbit_r64_c12 bl[12] br[12] wl[64] vdd gnd cell_6t
Xbit_r65_c12 bl[12] br[12] wl[65] vdd gnd cell_6t
Xbit_r66_c12 bl[12] br[12] wl[66] vdd gnd cell_6t
Xbit_r67_c12 bl[12] br[12] wl[67] vdd gnd cell_6t
Xbit_r68_c12 bl[12] br[12] wl[68] vdd gnd cell_6t
Xbit_r69_c12 bl[12] br[12] wl[69] vdd gnd cell_6t
Xbit_r70_c12 bl[12] br[12] wl[70] vdd gnd cell_6t
Xbit_r71_c12 bl[12] br[12] wl[71] vdd gnd cell_6t
Xbit_r72_c12 bl[12] br[12] wl[72] vdd gnd cell_6t
Xbit_r73_c12 bl[12] br[12] wl[73] vdd gnd cell_6t
Xbit_r74_c12 bl[12] br[12] wl[74] vdd gnd cell_6t
Xbit_r75_c12 bl[12] br[12] wl[75] vdd gnd cell_6t
Xbit_r76_c12 bl[12] br[12] wl[76] vdd gnd cell_6t
Xbit_r77_c12 bl[12] br[12] wl[77] vdd gnd cell_6t
Xbit_r78_c12 bl[12] br[12] wl[78] vdd gnd cell_6t
Xbit_r79_c12 bl[12] br[12] wl[79] vdd gnd cell_6t
Xbit_r80_c12 bl[12] br[12] wl[80] vdd gnd cell_6t
Xbit_r81_c12 bl[12] br[12] wl[81] vdd gnd cell_6t
Xbit_r82_c12 bl[12] br[12] wl[82] vdd gnd cell_6t
Xbit_r83_c12 bl[12] br[12] wl[83] vdd gnd cell_6t
Xbit_r84_c12 bl[12] br[12] wl[84] vdd gnd cell_6t
Xbit_r85_c12 bl[12] br[12] wl[85] vdd gnd cell_6t
Xbit_r86_c12 bl[12] br[12] wl[86] vdd gnd cell_6t
Xbit_r87_c12 bl[12] br[12] wl[87] vdd gnd cell_6t
Xbit_r88_c12 bl[12] br[12] wl[88] vdd gnd cell_6t
Xbit_r89_c12 bl[12] br[12] wl[89] vdd gnd cell_6t
Xbit_r90_c12 bl[12] br[12] wl[90] vdd gnd cell_6t
Xbit_r91_c12 bl[12] br[12] wl[91] vdd gnd cell_6t
Xbit_r92_c12 bl[12] br[12] wl[92] vdd gnd cell_6t
Xbit_r93_c12 bl[12] br[12] wl[93] vdd gnd cell_6t
Xbit_r94_c12 bl[12] br[12] wl[94] vdd gnd cell_6t
Xbit_r95_c12 bl[12] br[12] wl[95] vdd gnd cell_6t
Xbit_r96_c12 bl[12] br[12] wl[96] vdd gnd cell_6t
Xbit_r97_c12 bl[12] br[12] wl[97] vdd gnd cell_6t
Xbit_r98_c12 bl[12] br[12] wl[98] vdd gnd cell_6t
Xbit_r99_c12 bl[12] br[12] wl[99] vdd gnd cell_6t
Xbit_r100_c12 bl[12] br[12] wl[100] vdd gnd cell_6t
Xbit_r101_c12 bl[12] br[12] wl[101] vdd gnd cell_6t
Xbit_r102_c12 bl[12] br[12] wl[102] vdd gnd cell_6t
Xbit_r103_c12 bl[12] br[12] wl[103] vdd gnd cell_6t
Xbit_r104_c12 bl[12] br[12] wl[104] vdd gnd cell_6t
Xbit_r105_c12 bl[12] br[12] wl[105] vdd gnd cell_6t
Xbit_r106_c12 bl[12] br[12] wl[106] vdd gnd cell_6t
Xbit_r107_c12 bl[12] br[12] wl[107] vdd gnd cell_6t
Xbit_r108_c12 bl[12] br[12] wl[108] vdd gnd cell_6t
Xbit_r109_c12 bl[12] br[12] wl[109] vdd gnd cell_6t
Xbit_r110_c12 bl[12] br[12] wl[110] vdd gnd cell_6t
Xbit_r111_c12 bl[12] br[12] wl[111] vdd gnd cell_6t
Xbit_r112_c12 bl[12] br[12] wl[112] vdd gnd cell_6t
Xbit_r113_c12 bl[12] br[12] wl[113] vdd gnd cell_6t
Xbit_r114_c12 bl[12] br[12] wl[114] vdd gnd cell_6t
Xbit_r115_c12 bl[12] br[12] wl[115] vdd gnd cell_6t
Xbit_r116_c12 bl[12] br[12] wl[116] vdd gnd cell_6t
Xbit_r117_c12 bl[12] br[12] wl[117] vdd gnd cell_6t
Xbit_r118_c12 bl[12] br[12] wl[118] vdd gnd cell_6t
Xbit_r119_c12 bl[12] br[12] wl[119] vdd gnd cell_6t
Xbit_r120_c12 bl[12] br[12] wl[120] vdd gnd cell_6t
Xbit_r121_c12 bl[12] br[12] wl[121] vdd gnd cell_6t
Xbit_r122_c12 bl[12] br[12] wl[122] vdd gnd cell_6t
Xbit_r123_c12 bl[12] br[12] wl[123] vdd gnd cell_6t
Xbit_r124_c12 bl[12] br[12] wl[124] vdd gnd cell_6t
Xbit_r125_c12 bl[12] br[12] wl[125] vdd gnd cell_6t
Xbit_r126_c12 bl[12] br[12] wl[126] vdd gnd cell_6t
Xbit_r127_c12 bl[12] br[12] wl[127] vdd gnd cell_6t
Xbit_r0_c13 bl[13] br[13] wl[0] vdd gnd cell_6t
Xbit_r1_c13 bl[13] br[13] wl[1] vdd gnd cell_6t
Xbit_r2_c13 bl[13] br[13] wl[2] vdd gnd cell_6t
Xbit_r3_c13 bl[13] br[13] wl[3] vdd gnd cell_6t
Xbit_r4_c13 bl[13] br[13] wl[4] vdd gnd cell_6t
Xbit_r5_c13 bl[13] br[13] wl[5] vdd gnd cell_6t
Xbit_r6_c13 bl[13] br[13] wl[6] vdd gnd cell_6t
Xbit_r7_c13 bl[13] br[13] wl[7] vdd gnd cell_6t
Xbit_r8_c13 bl[13] br[13] wl[8] vdd gnd cell_6t
Xbit_r9_c13 bl[13] br[13] wl[9] vdd gnd cell_6t
Xbit_r10_c13 bl[13] br[13] wl[10] vdd gnd cell_6t
Xbit_r11_c13 bl[13] br[13] wl[11] vdd gnd cell_6t
Xbit_r12_c13 bl[13] br[13] wl[12] vdd gnd cell_6t
Xbit_r13_c13 bl[13] br[13] wl[13] vdd gnd cell_6t
Xbit_r14_c13 bl[13] br[13] wl[14] vdd gnd cell_6t
Xbit_r15_c13 bl[13] br[13] wl[15] vdd gnd cell_6t
Xbit_r16_c13 bl[13] br[13] wl[16] vdd gnd cell_6t
Xbit_r17_c13 bl[13] br[13] wl[17] vdd gnd cell_6t
Xbit_r18_c13 bl[13] br[13] wl[18] vdd gnd cell_6t
Xbit_r19_c13 bl[13] br[13] wl[19] vdd gnd cell_6t
Xbit_r20_c13 bl[13] br[13] wl[20] vdd gnd cell_6t
Xbit_r21_c13 bl[13] br[13] wl[21] vdd gnd cell_6t
Xbit_r22_c13 bl[13] br[13] wl[22] vdd gnd cell_6t
Xbit_r23_c13 bl[13] br[13] wl[23] vdd gnd cell_6t
Xbit_r24_c13 bl[13] br[13] wl[24] vdd gnd cell_6t
Xbit_r25_c13 bl[13] br[13] wl[25] vdd gnd cell_6t
Xbit_r26_c13 bl[13] br[13] wl[26] vdd gnd cell_6t
Xbit_r27_c13 bl[13] br[13] wl[27] vdd gnd cell_6t
Xbit_r28_c13 bl[13] br[13] wl[28] vdd gnd cell_6t
Xbit_r29_c13 bl[13] br[13] wl[29] vdd gnd cell_6t
Xbit_r30_c13 bl[13] br[13] wl[30] vdd gnd cell_6t
Xbit_r31_c13 bl[13] br[13] wl[31] vdd gnd cell_6t
Xbit_r32_c13 bl[13] br[13] wl[32] vdd gnd cell_6t
Xbit_r33_c13 bl[13] br[13] wl[33] vdd gnd cell_6t
Xbit_r34_c13 bl[13] br[13] wl[34] vdd gnd cell_6t
Xbit_r35_c13 bl[13] br[13] wl[35] vdd gnd cell_6t
Xbit_r36_c13 bl[13] br[13] wl[36] vdd gnd cell_6t
Xbit_r37_c13 bl[13] br[13] wl[37] vdd gnd cell_6t
Xbit_r38_c13 bl[13] br[13] wl[38] vdd gnd cell_6t
Xbit_r39_c13 bl[13] br[13] wl[39] vdd gnd cell_6t
Xbit_r40_c13 bl[13] br[13] wl[40] vdd gnd cell_6t
Xbit_r41_c13 bl[13] br[13] wl[41] vdd gnd cell_6t
Xbit_r42_c13 bl[13] br[13] wl[42] vdd gnd cell_6t
Xbit_r43_c13 bl[13] br[13] wl[43] vdd gnd cell_6t
Xbit_r44_c13 bl[13] br[13] wl[44] vdd gnd cell_6t
Xbit_r45_c13 bl[13] br[13] wl[45] vdd gnd cell_6t
Xbit_r46_c13 bl[13] br[13] wl[46] vdd gnd cell_6t
Xbit_r47_c13 bl[13] br[13] wl[47] vdd gnd cell_6t
Xbit_r48_c13 bl[13] br[13] wl[48] vdd gnd cell_6t
Xbit_r49_c13 bl[13] br[13] wl[49] vdd gnd cell_6t
Xbit_r50_c13 bl[13] br[13] wl[50] vdd gnd cell_6t
Xbit_r51_c13 bl[13] br[13] wl[51] vdd gnd cell_6t
Xbit_r52_c13 bl[13] br[13] wl[52] vdd gnd cell_6t
Xbit_r53_c13 bl[13] br[13] wl[53] vdd gnd cell_6t
Xbit_r54_c13 bl[13] br[13] wl[54] vdd gnd cell_6t
Xbit_r55_c13 bl[13] br[13] wl[55] vdd gnd cell_6t
Xbit_r56_c13 bl[13] br[13] wl[56] vdd gnd cell_6t
Xbit_r57_c13 bl[13] br[13] wl[57] vdd gnd cell_6t
Xbit_r58_c13 bl[13] br[13] wl[58] vdd gnd cell_6t
Xbit_r59_c13 bl[13] br[13] wl[59] vdd gnd cell_6t
Xbit_r60_c13 bl[13] br[13] wl[60] vdd gnd cell_6t
Xbit_r61_c13 bl[13] br[13] wl[61] vdd gnd cell_6t
Xbit_r62_c13 bl[13] br[13] wl[62] vdd gnd cell_6t
Xbit_r63_c13 bl[13] br[13] wl[63] vdd gnd cell_6t
Xbit_r64_c13 bl[13] br[13] wl[64] vdd gnd cell_6t
Xbit_r65_c13 bl[13] br[13] wl[65] vdd gnd cell_6t
Xbit_r66_c13 bl[13] br[13] wl[66] vdd gnd cell_6t
Xbit_r67_c13 bl[13] br[13] wl[67] vdd gnd cell_6t
Xbit_r68_c13 bl[13] br[13] wl[68] vdd gnd cell_6t
Xbit_r69_c13 bl[13] br[13] wl[69] vdd gnd cell_6t
Xbit_r70_c13 bl[13] br[13] wl[70] vdd gnd cell_6t
Xbit_r71_c13 bl[13] br[13] wl[71] vdd gnd cell_6t
Xbit_r72_c13 bl[13] br[13] wl[72] vdd gnd cell_6t
Xbit_r73_c13 bl[13] br[13] wl[73] vdd gnd cell_6t
Xbit_r74_c13 bl[13] br[13] wl[74] vdd gnd cell_6t
Xbit_r75_c13 bl[13] br[13] wl[75] vdd gnd cell_6t
Xbit_r76_c13 bl[13] br[13] wl[76] vdd gnd cell_6t
Xbit_r77_c13 bl[13] br[13] wl[77] vdd gnd cell_6t
Xbit_r78_c13 bl[13] br[13] wl[78] vdd gnd cell_6t
Xbit_r79_c13 bl[13] br[13] wl[79] vdd gnd cell_6t
Xbit_r80_c13 bl[13] br[13] wl[80] vdd gnd cell_6t
Xbit_r81_c13 bl[13] br[13] wl[81] vdd gnd cell_6t
Xbit_r82_c13 bl[13] br[13] wl[82] vdd gnd cell_6t
Xbit_r83_c13 bl[13] br[13] wl[83] vdd gnd cell_6t
Xbit_r84_c13 bl[13] br[13] wl[84] vdd gnd cell_6t
Xbit_r85_c13 bl[13] br[13] wl[85] vdd gnd cell_6t
Xbit_r86_c13 bl[13] br[13] wl[86] vdd gnd cell_6t
Xbit_r87_c13 bl[13] br[13] wl[87] vdd gnd cell_6t
Xbit_r88_c13 bl[13] br[13] wl[88] vdd gnd cell_6t
Xbit_r89_c13 bl[13] br[13] wl[89] vdd gnd cell_6t
Xbit_r90_c13 bl[13] br[13] wl[90] vdd gnd cell_6t
Xbit_r91_c13 bl[13] br[13] wl[91] vdd gnd cell_6t
Xbit_r92_c13 bl[13] br[13] wl[92] vdd gnd cell_6t
Xbit_r93_c13 bl[13] br[13] wl[93] vdd gnd cell_6t
Xbit_r94_c13 bl[13] br[13] wl[94] vdd gnd cell_6t
Xbit_r95_c13 bl[13] br[13] wl[95] vdd gnd cell_6t
Xbit_r96_c13 bl[13] br[13] wl[96] vdd gnd cell_6t
Xbit_r97_c13 bl[13] br[13] wl[97] vdd gnd cell_6t
Xbit_r98_c13 bl[13] br[13] wl[98] vdd gnd cell_6t
Xbit_r99_c13 bl[13] br[13] wl[99] vdd gnd cell_6t
Xbit_r100_c13 bl[13] br[13] wl[100] vdd gnd cell_6t
Xbit_r101_c13 bl[13] br[13] wl[101] vdd gnd cell_6t
Xbit_r102_c13 bl[13] br[13] wl[102] vdd gnd cell_6t
Xbit_r103_c13 bl[13] br[13] wl[103] vdd gnd cell_6t
Xbit_r104_c13 bl[13] br[13] wl[104] vdd gnd cell_6t
Xbit_r105_c13 bl[13] br[13] wl[105] vdd gnd cell_6t
Xbit_r106_c13 bl[13] br[13] wl[106] vdd gnd cell_6t
Xbit_r107_c13 bl[13] br[13] wl[107] vdd gnd cell_6t
Xbit_r108_c13 bl[13] br[13] wl[108] vdd gnd cell_6t
Xbit_r109_c13 bl[13] br[13] wl[109] vdd gnd cell_6t
Xbit_r110_c13 bl[13] br[13] wl[110] vdd gnd cell_6t
Xbit_r111_c13 bl[13] br[13] wl[111] vdd gnd cell_6t
Xbit_r112_c13 bl[13] br[13] wl[112] vdd gnd cell_6t
Xbit_r113_c13 bl[13] br[13] wl[113] vdd gnd cell_6t
Xbit_r114_c13 bl[13] br[13] wl[114] vdd gnd cell_6t
Xbit_r115_c13 bl[13] br[13] wl[115] vdd gnd cell_6t
Xbit_r116_c13 bl[13] br[13] wl[116] vdd gnd cell_6t
Xbit_r117_c13 bl[13] br[13] wl[117] vdd gnd cell_6t
Xbit_r118_c13 bl[13] br[13] wl[118] vdd gnd cell_6t
Xbit_r119_c13 bl[13] br[13] wl[119] vdd gnd cell_6t
Xbit_r120_c13 bl[13] br[13] wl[120] vdd gnd cell_6t
Xbit_r121_c13 bl[13] br[13] wl[121] vdd gnd cell_6t
Xbit_r122_c13 bl[13] br[13] wl[122] vdd gnd cell_6t
Xbit_r123_c13 bl[13] br[13] wl[123] vdd gnd cell_6t
Xbit_r124_c13 bl[13] br[13] wl[124] vdd gnd cell_6t
Xbit_r125_c13 bl[13] br[13] wl[125] vdd gnd cell_6t
Xbit_r126_c13 bl[13] br[13] wl[126] vdd gnd cell_6t
Xbit_r127_c13 bl[13] br[13] wl[127] vdd gnd cell_6t
Xbit_r0_c14 bl[14] br[14] wl[0] vdd gnd cell_6t
Xbit_r1_c14 bl[14] br[14] wl[1] vdd gnd cell_6t
Xbit_r2_c14 bl[14] br[14] wl[2] vdd gnd cell_6t
Xbit_r3_c14 bl[14] br[14] wl[3] vdd gnd cell_6t
Xbit_r4_c14 bl[14] br[14] wl[4] vdd gnd cell_6t
Xbit_r5_c14 bl[14] br[14] wl[5] vdd gnd cell_6t
Xbit_r6_c14 bl[14] br[14] wl[6] vdd gnd cell_6t
Xbit_r7_c14 bl[14] br[14] wl[7] vdd gnd cell_6t
Xbit_r8_c14 bl[14] br[14] wl[8] vdd gnd cell_6t
Xbit_r9_c14 bl[14] br[14] wl[9] vdd gnd cell_6t
Xbit_r10_c14 bl[14] br[14] wl[10] vdd gnd cell_6t
Xbit_r11_c14 bl[14] br[14] wl[11] vdd gnd cell_6t
Xbit_r12_c14 bl[14] br[14] wl[12] vdd gnd cell_6t
Xbit_r13_c14 bl[14] br[14] wl[13] vdd gnd cell_6t
Xbit_r14_c14 bl[14] br[14] wl[14] vdd gnd cell_6t
Xbit_r15_c14 bl[14] br[14] wl[15] vdd gnd cell_6t
Xbit_r16_c14 bl[14] br[14] wl[16] vdd gnd cell_6t
Xbit_r17_c14 bl[14] br[14] wl[17] vdd gnd cell_6t
Xbit_r18_c14 bl[14] br[14] wl[18] vdd gnd cell_6t
Xbit_r19_c14 bl[14] br[14] wl[19] vdd gnd cell_6t
Xbit_r20_c14 bl[14] br[14] wl[20] vdd gnd cell_6t
Xbit_r21_c14 bl[14] br[14] wl[21] vdd gnd cell_6t
Xbit_r22_c14 bl[14] br[14] wl[22] vdd gnd cell_6t
Xbit_r23_c14 bl[14] br[14] wl[23] vdd gnd cell_6t
Xbit_r24_c14 bl[14] br[14] wl[24] vdd gnd cell_6t
Xbit_r25_c14 bl[14] br[14] wl[25] vdd gnd cell_6t
Xbit_r26_c14 bl[14] br[14] wl[26] vdd gnd cell_6t
Xbit_r27_c14 bl[14] br[14] wl[27] vdd gnd cell_6t
Xbit_r28_c14 bl[14] br[14] wl[28] vdd gnd cell_6t
Xbit_r29_c14 bl[14] br[14] wl[29] vdd gnd cell_6t
Xbit_r30_c14 bl[14] br[14] wl[30] vdd gnd cell_6t
Xbit_r31_c14 bl[14] br[14] wl[31] vdd gnd cell_6t
Xbit_r32_c14 bl[14] br[14] wl[32] vdd gnd cell_6t
Xbit_r33_c14 bl[14] br[14] wl[33] vdd gnd cell_6t
Xbit_r34_c14 bl[14] br[14] wl[34] vdd gnd cell_6t
Xbit_r35_c14 bl[14] br[14] wl[35] vdd gnd cell_6t
Xbit_r36_c14 bl[14] br[14] wl[36] vdd gnd cell_6t
Xbit_r37_c14 bl[14] br[14] wl[37] vdd gnd cell_6t
Xbit_r38_c14 bl[14] br[14] wl[38] vdd gnd cell_6t
Xbit_r39_c14 bl[14] br[14] wl[39] vdd gnd cell_6t
Xbit_r40_c14 bl[14] br[14] wl[40] vdd gnd cell_6t
Xbit_r41_c14 bl[14] br[14] wl[41] vdd gnd cell_6t
Xbit_r42_c14 bl[14] br[14] wl[42] vdd gnd cell_6t
Xbit_r43_c14 bl[14] br[14] wl[43] vdd gnd cell_6t
Xbit_r44_c14 bl[14] br[14] wl[44] vdd gnd cell_6t
Xbit_r45_c14 bl[14] br[14] wl[45] vdd gnd cell_6t
Xbit_r46_c14 bl[14] br[14] wl[46] vdd gnd cell_6t
Xbit_r47_c14 bl[14] br[14] wl[47] vdd gnd cell_6t
Xbit_r48_c14 bl[14] br[14] wl[48] vdd gnd cell_6t
Xbit_r49_c14 bl[14] br[14] wl[49] vdd gnd cell_6t
Xbit_r50_c14 bl[14] br[14] wl[50] vdd gnd cell_6t
Xbit_r51_c14 bl[14] br[14] wl[51] vdd gnd cell_6t
Xbit_r52_c14 bl[14] br[14] wl[52] vdd gnd cell_6t
Xbit_r53_c14 bl[14] br[14] wl[53] vdd gnd cell_6t
Xbit_r54_c14 bl[14] br[14] wl[54] vdd gnd cell_6t
Xbit_r55_c14 bl[14] br[14] wl[55] vdd gnd cell_6t
Xbit_r56_c14 bl[14] br[14] wl[56] vdd gnd cell_6t
Xbit_r57_c14 bl[14] br[14] wl[57] vdd gnd cell_6t
Xbit_r58_c14 bl[14] br[14] wl[58] vdd gnd cell_6t
Xbit_r59_c14 bl[14] br[14] wl[59] vdd gnd cell_6t
Xbit_r60_c14 bl[14] br[14] wl[60] vdd gnd cell_6t
Xbit_r61_c14 bl[14] br[14] wl[61] vdd gnd cell_6t
Xbit_r62_c14 bl[14] br[14] wl[62] vdd gnd cell_6t
Xbit_r63_c14 bl[14] br[14] wl[63] vdd gnd cell_6t
Xbit_r64_c14 bl[14] br[14] wl[64] vdd gnd cell_6t
Xbit_r65_c14 bl[14] br[14] wl[65] vdd gnd cell_6t
Xbit_r66_c14 bl[14] br[14] wl[66] vdd gnd cell_6t
Xbit_r67_c14 bl[14] br[14] wl[67] vdd gnd cell_6t
Xbit_r68_c14 bl[14] br[14] wl[68] vdd gnd cell_6t
Xbit_r69_c14 bl[14] br[14] wl[69] vdd gnd cell_6t
Xbit_r70_c14 bl[14] br[14] wl[70] vdd gnd cell_6t
Xbit_r71_c14 bl[14] br[14] wl[71] vdd gnd cell_6t
Xbit_r72_c14 bl[14] br[14] wl[72] vdd gnd cell_6t
Xbit_r73_c14 bl[14] br[14] wl[73] vdd gnd cell_6t
Xbit_r74_c14 bl[14] br[14] wl[74] vdd gnd cell_6t
Xbit_r75_c14 bl[14] br[14] wl[75] vdd gnd cell_6t
Xbit_r76_c14 bl[14] br[14] wl[76] vdd gnd cell_6t
Xbit_r77_c14 bl[14] br[14] wl[77] vdd gnd cell_6t
Xbit_r78_c14 bl[14] br[14] wl[78] vdd gnd cell_6t
Xbit_r79_c14 bl[14] br[14] wl[79] vdd gnd cell_6t
Xbit_r80_c14 bl[14] br[14] wl[80] vdd gnd cell_6t
Xbit_r81_c14 bl[14] br[14] wl[81] vdd gnd cell_6t
Xbit_r82_c14 bl[14] br[14] wl[82] vdd gnd cell_6t
Xbit_r83_c14 bl[14] br[14] wl[83] vdd gnd cell_6t
Xbit_r84_c14 bl[14] br[14] wl[84] vdd gnd cell_6t
Xbit_r85_c14 bl[14] br[14] wl[85] vdd gnd cell_6t
Xbit_r86_c14 bl[14] br[14] wl[86] vdd gnd cell_6t
Xbit_r87_c14 bl[14] br[14] wl[87] vdd gnd cell_6t
Xbit_r88_c14 bl[14] br[14] wl[88] vdd gnd cell_6t
Xbit_r89_c14 bl[14] br[14] wl[89] vdd gnd cell_6t
Xbit_r90_c14 bl[14] br[14] wl[90] vdd gnd cell_6t
Xbit_r91_c14 bl[14] br[14] wl[91] vdd gnd cell_6t
Xbit_r92_c14 bl[14] br[14] wl[92] vdd gnd cell_6t
Xbit_r93_c14 bl[14] br[14] wl[93] vdd gnd cell_6t
Xbit_r94_c14 bl[14] br[14] wl[94] vdd gnd cell_6t
Xbit_r95_c14 bl[14] br[14] wl[95] vdd gnd cell_6t
Xbit_r96_c14 bl[14] br[14] wl[96] vdd gnd cell_6t
Xbit_r97_c14 bl[14] br[14] wl[97] vdd gnd cell_6t
Xbit_r98_c14 bl[14] br[14] wl[98] vdd gnd cell_6t
Xbit_r99_c14 bl[14] br[14] wl[99] vdd gnd cell_6t
Xbit_r100_c14 bl[14] br[14] wl[100] vdd gnd cell_6t
Xbit_r101_c14 bl[14] br[14] wl[101] vdd gnd cell_6t
Xbit_r102_c14 bl[14] br[14] wl[102] vdd gnd cell_6t
Xbit_r103_c14 bl[14] br[14] wl[103] vdd gnd cell_6t
Xbit_r104_c14 bl[14] br[14] wl[104] vdd gnd cell_6t
Xbit_r105_c14 bl[14] br[14] wl[105] vdd gnd cell_6t
Xbit_r106_c14 bl[14] br[14] wl[106] vdd gnd cell_6t
Xbit_r107_c14 bl[14] br[14] wl[107] vdd gnd cell_6t
Xbit_r108_c14 bl[14] br[14] wl[108] vdd gnd cell_6t
Xbit_r109_c14 bl[14] br[14] wl[109] vdd gnd cell_6t
Xbit_r110_c14 bl[14] br[14] wl[110] vdd gnd cell_6t
Xbit_r111_c14 bl[14] br[14] wl[111] vdd gnd cell_6t
Xbit_r112_c14 bl[14] br[14] wl[112] vdd gnd cell_6t
Xbit_r113_c14 bl[14] br[14] wl[113] vdd gnd cell_6t
Xbit_r114_c14 bl[14] br[14] wl[114] vdd gnd cell_6t
Xbit_r115_c14 bl[14] br[14] wl[115] vdd gnd cell_6t
Xbit_r116_c14 bl[14] br[14] wl[116] vdd gnd cell_6t
Xbit_r117_c14 bl[14] br[14] wl[117] vdd gnd cell_6t
Xbit_r118_c14 bl[14] br[14] wl[118] vdd gnd cell_6t
Xbit_r119_c14 bl[14] br[14] wl[119] vdd gnd cell_6t
Xbit_r120_c14 bl[14] br[14] wl[120] vdd gnd cell_6t
Xbit_r121_c14 bl[14] br[14] wl[121] vdd gnd cell_6t
Xbit_r122_c14 bl[14] br[14] wl[122] vdd gnd cell_6t
Xbit_r123_c14 bl[14] br[14] wl[123] vdd gnd cell_6t
Xbit_r124_c14 bl[14] br[14] wl[124] vdd gnd cell_6t
Xbit_r125_c14 bl[14] br[14] wl[125] vdd gnd cell_6t
Xbit_r126_c14 bl[14] br[14] wl[126] vdd gnd cell_6t
Xbit_r127_c14 bl[14] br[14] wl[127] vdd gnd cell_6t
Xbit_r0_c15 bl[15] br[15] wl[0] vdd gnd cell_6t
Xbit_r1_c15 bl[15] br[15] wl[1] vdd gnd cell_6t
Xbit_r2_c15 bl[15] br[15] wl[2] vdd gnd cell_6t
Xbit_r3_c15 bl[15] br[15] wl[3] vdd gnd cell_6t
Xbit_r4_c15 bl[15] br[15] wl[4] vdd gnd cell_6t
Xbit_r5_c15 bl[15] br[15] wl[5] vdd gnd cell_6t
Xbit_r6_c15 bl[15] br[15] wl[6] vdd gnd cell_6t
Xbit_r7_c15 bl[15] br[15] wl[7] vdd gnd cell_6t
Xbit_r8_c15 bl[15] br[15] wl[8] vdd gnd cell_6t
Xbit_r9_c15 bl[15] br[15] wl[9] vdd gnd cell_6t
Xbit_r10_c15 bl[15] br[15] wl[10] vdd gnd cell_6t
Xbit_r11_c15 bl[15] br[15] wl[11] vdd gnd cell_6t
Xbit_r12_c15 bl[15] br[15] wl[12] vdd gnd cell_6t
Xbit_r13_c15 bl[15] br[15] wl[13] vdd gnd cell_6t
Xbit_r14_c15 bl[15] br[15] wl[14] vdd gnd cell_6t
Xbit_r15_c15 bl[15] br[15] wl[15] vdd gnd cell_6t
Xbit_r16_c15 bl[15] br[15] wl[16] vdd gnd cell_6t
Xbit_r17_c15 bl[15] br[15] wl[17] vdd gnd cell_6t
Xbit_r18_c15 bl[15] br[15] wl[18] vdd gnd cell_6t
Xbit_r19_c15 bl[15] br[15] wl[19] vdd gnd cell_6t
Xbit_r20_c15 bl[15] br[15] wl[20] vdd gnd cell_6t
Xbit_r21_c15 bl[15] br[15] wl[21] vdd gnd cell_6t
Xbit_r22_c15 bl[15] br[15] wl[22] vdd gnd cell_6t
Xbit_r23_c15 bl[15] br[15] wl[23] vdd gnd cell_6t
Xbit_r24_c15 bl[15] br[15] wl[24] vdd gnd cell_6t
Xbit_r25_c15 bl[15] br[15] wl[25] vdd gnd cell_6t
Xbit_r26_c15 bl[15] br[15] wl[26] vdd gnd cell_6t
Xbit_r27_c15 bl[15] br[15] wl[27] vdd gnd cell_6t
Xbit_r28_c15 bl[15] br[15] wl[28] vdd gnd cell_6t
Xbit_r29_c15 bl[15] br[15] wl[29] vdd gnd cell_6t
Xbit_r30_c15 bl[15] br[15] wl[30] vdd gnd cell_6t
Xbit_r31_c15 bl[15] br[15] wl[31] vdd gnd cell_6t
Xbit_r32_c15 bl[15] br[15] wl[32] vdd gnd cell_6t
Xbit_r33_c15 bl[15] br[15] wl[33] vdd gnd cell_6t
Xbit_r34_c15 bl[15] br[15] wl[34] vdd gnd cell_6t
Xbit_r35_c15 bl[15] br[15] wl[35] vdd gnd cell_6t
Xbit_r36_c15 bl[15] br[15] wl[36] vdd gnd cell_6t
Xbit_r37_c15 bl[15] br[15] wl[37] vdd gnd cell_6t
Xbit_r38_c15 bl[15] br[15] wl[38] vdd gnd cell_6t
Xbit_r39_c15 bl[15] br[15] wl[39] vdd gnd cell_6t
Xbit_r40_c15 bl[15] br[15] wl[40] vdd gnd cell_6t
Xbit_r41_c15 bl[15] br[15] wl[41] vdd gnd cell_6t
Xbit_r42_c15 bl[15] br[15] wl[42] vdd gnd cell_6t
Xbit_r43_c15 bl[15] br[15] wl[43] vdd gnd cell_6t
Xbit_r44_c15 bl[15] br[15] wl[44] vdd gnd cell_6t
Xbit_r45_c15 bl[15] br[15] wl[45] vdd gnd cell_6t
Xbit_r46_c15 bl[15] br[15] wl[46] vdd gnd cell_6t
Xbit_r47_c15 bl[15] br[15] wl[47] vdd gnd cell_6t
Xbit_r48_c15 bl[15] br[15] wl[48] vdd gnd cell_6t
Xbit_r49_c15 bl[15] br[15] wl[49] vdd gnd cell_6t
Xbit_r50_c15 bl[15] br[15] wl[50] vdd gnd cell_6t
Xbit_r51_c15 bl[15] br[15] wl[51] vdd gnd cell_6t
Xbit_r52_c15 bl[15] br[15] wl[52] vdd gnd cell_6t
Xbit_r53_c15 bl[15] br[15] wl[53] vdd gnd cell_6t
Xbit_r54_c15 bl[15] br[15] wl[54] vdd gnd cell_6t
Xbit_r55_c15 bl[15] br[15] wl[55] vdd gnd cell_6t
Xbit_r56_c15 bl[15] br[15] wl[56] vdd gnd cell_6t
Xbit_r57_c15 bl[15] br[15] wl[57] vdd gnd cell_6t
Xbit_r58_c15 bl[15] br[15] wl[58] vdd gnd cell_6t
Xbit_r59_c15 bl[15] br[15] wl[59] vdd gnd cell_6t
Xbit_r60_c15 bl[15] br[15] wl[60] vdd gnd cell_6t
Xbit_r61_c15 bl[15] br[15] wl[61] vdd gnd cell_6t
Xbit_r62_c15 bl[15] br[15] wl[62] vdd gnd cell_6t
Xbit_r63_c15 bl[15] br[15] wl[63] vdd gnd cell_6t
Xbit_r64_c15 bl[15] br[15] wl[64] vdd gnd cell_6t
Xbit_r65_c15 bl[15] br[15] wl[65] vdd gnd cell_6t
Xbit_r66_c15 bl[15] br[15] wl[66] vdd gnd cell_6t
Xbit_r67_c15 bl[15] br[15] wl[67] vdd gnd cell_6t
Xbit_r68_c15 bl[15] br[15] wl[68] vdd gnd cell_6t
Xbit_r69_c15 bl[15] br[15] wl[69] vdd gnd cell_6t
Xbit_r70_c15 bl[15] br[15] wl[70] vdd gnd cell_6t
Xbit_r71_c15 bl[15] br[15] wl[71] vdd gnd cell_6t
Xbit_r72_c15 bl[15] br[15] wl[72] vdd gnd cell_6t
Xbit_r73_c15 bl[15] br[15] wl[73] vdd gnd cell_6t
Xbit_r74_c15 bl[15] br[15] wl[74] vdd gnd cell_6t
Xbit_r75_c15 bl[15] br[15] wl[75] vdd gnd cell_6t
Xbit_r76_c15 bl[15] br[15] wl[76] vdd gnd cell_6t
Xbit_r77_c15 bl[15] br[15] wl[77] vdd gnd cell_6t
Xbit_r78_c15 bl[15] br[15] wl[78] vdd gnd cell_6t
Xbit_r79_c15 bl[15] br[15] wl[79] vdd gnd cell_6t
Xbit_r80_c15 bl[15] br[15] wl[80] vdd gnd cell_6t
Xbit_r81_c15 bl[15] br[15] wl[81] vdd gnd cell_6t
Xbit_r82_c15 bl[15] br[15] wl[82] vdd gnd cell_6t
Xbit_r83_c15 bl[15] br[15] wl[83] vdd gnd cell_6t
Xbit_r84_c15 bl[15] br[15] wl[84] vdd gnd cell_6t
Xbit_r85_c15 bl[15] br[15] wl[85] vdd gnd cell_6t
Xbit_r86_c15 bl[15] br[15] wl[86] vdd gnd cell_6t
Xbit_r87_c15 bl[15] br[15] wl[87] vdd gnd cell_6t
Xbit_r88_c15 bl[15] br[15] wl[88] vdd gnd cell_6t
Xbit_r89_c15 bl[15] br[15] wl[89] vdd gnd cell_6t
Xbit_r90_c15 bl[15] br[15] wl[90] vdd gnd cell_6t
Xbit_r91_c15 bl[15] br[15] wl[91] vdd gnd cell_6t
Xbit_r92_c15 bl[15] br[15] wl[92] vdd gnd cell_6t
Xbit_r93_c15 bl[15] br[15] wl[93] vdd gnd cell_6t
Xbit_r94_c15 bl[15] br[15] wl[94] vdd gnd cell_6t
Xbit_r95_c15 bl[15] br[15] wl[95] vdd gnd cell_6t
Xbit_r96_c15 bl[15] br[15] wl[96] vdd gnd cell_6t
Xbit_r97_c15 bl[15] br[15] wl[97] vdd gnd cell_6t
Xbit_r98_c15 bl[15] br[15] wl[98] vdd gnd cell_6t
Xbit_r99_c15 bl[15] br[15] wl[99] vdd gnd cell_6t
Xbit_r100_c15 bl[15] br[15] wl[100] vdd gnd cell_6t
Xbit_r101_c15 bl[15] br[15] wl[101] vdd gnd cell_6t
Xbit_r102_c15 bl[15] br[15] wl[102] vdd gnd cell_6t
Xbit_r103_c15 bl[15] br[15] wl[103] vdd gnd cell_6t
Xbit_r104_c15 bl[15] br[15] wl[104] vdd gnd cell_6t
Xbit_r105_c15 bl[15] br[15] wl[105] vdd gnd cell_6t
Xbit_r106_c15 bl[15] br[15] wl[106] vdd gnd cell_6t
Xbit_r107_c15 bl[15] br[15] wl[107] vdd gnd cell_6t
Xbit_r108_c15 bl[15] br[15] wl[108] vdd gnd cell_6t
Xbit_r109_c15 bl[15] br[15] wl[109] vdd gnd cell_6t
Xbit_r110_c15 bl[15] br[15] wl[110] vdd gnd cell_6t
Xbit_r111_c15 bl[15] br[15] wl[111] vdd gnd cell_6t
Xbit_r112_c15 bl[15] br[15] wl[112] vdd gnd cell_6t
Xbit_r113_c15 bl[15] br[15] wl[113] vdd gnd cell_6t
Xbit_r114_c15 bl[15] br[15] wl[114] vdd gnd cell_6t
Xbit_r115_c15 bl[15] br[15] wl[115] vdd gnd cell_6t
Xbit_r116_c15 bl[15] br[15] wl[116] vdd gnd cell_6t
Xbit_r117_c15 bl[15] br[15] wl[117] vdd gnd cell_6t
Xbit_r118_c15 bl[15] br[15] wl[118] vdd gnd cell_6t
Xbit_r119_c15 bl[15] br[15] wl[119] vdd gnd cell_6t
Xbit_r120_c15 bl[15] br[15] wl[120] vdd gnd cell_6t
Xbit_r121_c15 bl[15] br[15] wl[121] vdd gnd cell_6t
Xbit_r122_c15 bl[15] br[15] wl[122] vdd gnd cell_6t
Xbit_r123_c15 bl[15] br[15] wl[123] vdd gnd cell_6t
Xbit_r124_c15 bl[15] br[15] wl[124] vdd gnd cell_6t
Xbit_r125_c15 bl[15] br[15] wl[125] vdd gnd cell_6t
Xbit_r126_c15 bl[15] br[15] wl[126] vdd gnd cell_6t
Xbit_r127_c15 bl[15] br[15] wl[127] vdd gnd cell_6t
Xbit_r0_c16 bl[16] br[16] wl[0] vdd gnd cell_6t
Xbit_r1_c16 bl[16] br[16] wl[1] vdd gnd cell_6t
Xbit_r2_c16 bl[16] br[16] wl[2] vdd gnd cell_6t
Xbit_r3_c16 bl[16] br[16] wl[3] vdd gnd cell_6t
Xbit_r4_c16 bl[16] br[16] wl[4] vdd gnd cell_6t
Xbit_r5_c16 bl[16] br[16] wl[5] vdd gnd cell_6t
Xbit_r6_c16 bl[16] br[16] wl[6] vdd gnd cell_6t
Xbit_r7_c16 bl[16] br[16] wl[7] vdd gnd cell_6t
Xbit_r8_c16 bl[16] br[16] wl[8] vdd gnd cell_6t
Xbit_r9_c16 bl[16] br[16] wl[9] vdd gnd cell_6t
Xbit_r10_c16 bl[16] br[16] wl[10] vdd gnd cell_6t
Xbit_r11_c16 bl[16] br[16] wl[11] vdd gnd cell_6t
Xbit_r12_c16 bl[16] br[16] wl[12] vdd gnd cell_6t
Xbit_r13_c16 bl[16] br[16] wl[13] vdd gnd cell_6t
Xbit_r14_c16 bl[16] br[16] wl[14] vdd gnd cell_6t
Xbit_r15_c16 bl[16] br[16] wl[15] vdd gnd cell_6t
Xbit_r16_c16 bl[16] br[16] wl[16] vdd gnd cell_6t
Xbit_r17_c16 bl[16] br[16] wl[17] vdd gnd cell_6t
Xbit_r18_c16 bl[16] br[16] wl[18] vdd gnd cell_6t
Xbit_r19_c16 bl[16] br[16] wl[19] vdd gnd cell_6t
Xbit_r20_c16 bl[16] br[16] wl[20] vdd gnd cell_6t
Xbit_r21_c16 bl[16] br[16] wl[21] vdd gnd cell_6t
Xbit_r22_c16 bl[16] br[16] wl[22] vdd gnd cell_6t
Xbit_r23_c16 bl[16] br[16] wl[23] vdd gnd cell_6t
Xbit_r24_c16 bl[16] br[16] wl[24] vdd gnd cell_6t
Xbit_r25_c16 bl[16] br[16] wl[25] vdd gnd cell_6t
Xbit_r26_c16 bl[16] br[16] wl[26] vdd gnd cell_6t
Xbit_r27_c16 bl[16] br[16] wl[27] vdd gnd cell_6t
Xbit_r28_c16 bl[16] br[16] wl[28] vdd gnd cell_6t
Xbit_r29_c16 bl[16] br[16] wl[29] vdd gnd cell_6t
Xbit_r30_c16 bl[16] br[16] wl[30] vdd gnd cell_6t
Xbit_r31_c16 bl[16] br[16] wl[31] vdd gnd cell_6t
Xbit_r32_c16 bl[16] br[16] wl[32] vdd gnd cell_6t
Xbit_r33_c16 bl[16] br[16] wl[33] vdd gnd cell_6t
Xbit_r34_c16 bl[16] br[16] wl[34] vdd gnd cell_6t
Xbit_r35_c16 bl[16] br[16] wl[35] vdd gnd cell_6t
Xbit_r36_c16 bl[16] br[16] wl[36] vdd gnd cell_6t
Xbit_r37_c16 bl[16] br[16] wl[37] vdd gnd cell_6t
Xbit_r38_c16 bl[16] br[16] wl[38] vdd gnd cell_6t
Xbit_r39_c16 bl[16] br[16] wl[39] vdd gnd cell_6t
Xbit_r40_c16 bl[16] br[16] wl[40] vdd gnd cell_6t
Xbit_r41_c16 bl[16] br[16] wl[41] vdd gnd cell_6t
Xbit_r42_c16 bl[16] br[16] wl[42] vdd gnd cell_6t
Xbit_r43_c16 bl[16] br[16] wl[43] vdd gnd cell_6t
Xbit_r44_c16 bl[16] br[16] wl[44] vdd gnd cell_6t
Xbit_r45_c16 bl[16] br[16] wl[45] vdd gnd cell_6t
Xbit_r46_c16 bl[16] br[16] wl[46] vdd gnd cell_6t
Xbit_r47_c16 bl[16] br[16] wl[47] vdd gnd cell_6t
Xbit_r48_c16 bl[16] br[16] wl[48] vdd gnd cell_6t
Xbit_r49_c16 bl[16] br[16] wl[49] vdd gnd cell_6t
Xbit_r50_c16 bl[16] br[16] wl[50] vdd gnd cell_6t
Xbit_r51_c16 bl[16] br[16] wl[51] vdd gnd cell_6t
Xbit_r52_c16 bl[16] br[16] wl[52] vdd gnd cell_6t
Xbit_r53_c16 bl[16] br[16] wl[53] vdd gnd cell_6t
Xbit_r54_c16 bl[16] br[16] wl[54] vdd gnd cell_6t
Xbit_r55_c16 bl[16] br[16] wl[55] vdd gnd cell_6t
Xbit_r56_c16 bl[16] br[16] wl[56] vdd gnd cell_6t
Xbit_r57_c16 bl[16] br[16] wl[57] vdd gnd cell_6t
Xbit_r58_c16 bl[16] br[16] wl[58] vdd gnd cell_6t
Xbit_r59_c16 bl[16] br[16] wl[59] vdd gnd cell_6t
Xbit_r60_c16 bl[16] br[16] wl[60] vdd gnd cell_6t
Xbit_r61_c16 bl[16] br[16] wl[61] vdd gnd cell_6t
Xbit_r62_c16 bl[16] br[16] wl[62] vdd gnd cell_6t
Xbit_r63_c16 bl[16] br[16] wl[63] vdd gnd cell_6t
Xbit_r64_c16 bl[16] br[16] wl[64] vdd gnd cell_6t
Xbit_r65_c16 bl[16] br[16] wl[65] vdd gnd cell_6t
Xbit_r66_c16 bl[16] br[16] wl[66] vdd gnd cell_6t
Xbit_r67_c16 bl[16] br[16] wl[67] vdd gnd cell_6t
Xbit_r68_c16 bl[16] br[16] wl[68] vdd gnd cell_6t
Xbit_r69_c16 bl[16] br[16] wl[69] vdd gnd cell_6t
Xbit_r70_c16 bl[16] br[16] wl[70] vdd gnd cell_6t
Xbit_r71_c16 bl[16] br[16] wl[71] vdd gnd cell_6t
Xbit_r72_c16 bl[16] br[16] wl[72] vdd gnd cell_6t
Xbit_r73_c16 bl[16] br[16] wl[73] vdd gnd cell_6t
Xbit_r74_c16 bl[16] br[16] wl[74] vdd gnd cell_6t
Xbit_r75_c16 bl[16] br[16] wl[75] vdd gnd cell_6t
Xbit_r76_c16 bl[16] br[16] wl[76] vdd gnd cell_6t
Xbit_r77_c16 bl[16] br[16] wl[77] vdd gnd cell_6t
Xbit_r78_c16 bl[16] br[16] wl[78] vdd gnd cell_6t
Xbit_r79_c16 bl[16] br[16] wl[79] vdd gnd cell_6t
Xbit_r80_c16 bl[16] br[16] wl[80] vdd gnd cell_6t
Xbit_r81_c16 bl[16] br[16] wl[81] vdd gnd cell_6t
Xbit_r82_c16 bl[16] br[16] wl[82] vdd gnd cell_6t
Xbit_r83_c16 bl[16] br[16] wl[83] vdd gnd cell_6t
Xbit_r84_c16 bl[16] br[16] wl[84] vdd gnd cell_6t
Xbit_r85_c16 bl[16] br[16] wl[85] vdd gnd cell_6t
Xbit_r86_c16 bl[16] br[16] wl[86] vdd gnd cell_6t
Xbit_r87_c16 bl[16] br[16] wl[87] vdd gnd cell_6t
Xbit_r88_c16 bl[16] br[16] wl[88] vdd gnd cell_6t
Xbit_r89_c16 bl[16] br[16] wl[89] vdd gnd cell_6t
Xbit_r90_c16 bl[16] br[16] wl[90] vdd gnd cell_6t
Xbit_r91_c16 bl[16] br[16] wl[91] vdd gnd cell_6t
Xbit_r92_c16 bl[16] br[16] wl[92] vdd gnd cell_6t
Xbit_r93_c16 bl[16] br[16] wl[93] vdd gnd cell_6t
Xbit_r94_c16 bl[16] br[16] wl[94] vdd gnd cell_6t
Xbit_r95_c16 bl[16] br[16] wl[95] vdd gnd cell_6t
Xbit_r96_c16 bl[16] br[16] wl[96] vdd gnd cell_6t
Xbit_r97_c16 bl[16] br[16] wl[97] vdd gnd cell_6t
Xbit_r98_c16 bl[16] br[16] wl[98] vdd gnd cell_6t
Xbit_r99_c16 bl[16] br[16] wl[99] vdd gnd cell_6t
Xbit_r100_c16 bl[16] br[16] wl[100] vdd gnd cell_6t
Xbit_r101_c16 bl[16] br[16] wl[101] vdd gnd cell_6t
Xbit_r102_c16 bl[16] br[16] wl[102] vdd gnd cell_6t
Xbit_r103_c16 bl[16] br[16] wl[103] vdd gnd cell_6t
Xbit_r104_c16 bl[16] br[16] wl[104] vdd gnd cell_6t
Xbit_r105_c16 bl[16] br[16] wl[105] vdd gnd cell_6t
Xbit_r106_c16 bl[16] br[16] wl[106] vdd gnd cell_6t
Xbit_r107_c16 bl[16] br[16] wl[107] vdd gnd cell_6t
Xbit_r108_c16 bl[16] br[16] wl[108] vdd gnd cell_6t
Xbit_r109_c16 bl[16] br[16] wl[109] vdd gnd cell_6t
Xbit_r110_c16 bl[16] br[16] wl[110] vdd gnd cell_6t
Xbit_r111_c16 bl[16] br[16] wl[111] vdd gnd cell_6t
Xbit_r112_c16 bl[16] br[16] wl[112] vdd gnd cell_6t
Xbit_r113_c16 bl[16] br[16] wl[113] vdd gnd cell_6t
Xbit_r114_c16 bl[16] br[16] wl[114] vdd gnd cell_6t
Xbit_r115_c16 bl[16] br[16] wl[115] vdd gnd cell_6t
Xbit_r116_c16 bl[16] br[16] wl[116] vdd gnd cell_6t
Xbit_r117_c16 bl[16] br[16] wl[117] vdd gnd cell_6t
Xbit_r118_c16 bl[16] br[16] wl[118] vdd gnd cell_6t
Xbit_r119_c16 bl[16] br[16] wl[119] vdd gnd cell_6t
Xbit_r120_c16 bl[16] br[16] wl[120] vdd gnd cell_6t
Xbit_r121_c16 bl[16] br[16] wl[121] vdd gnd cell_6t
Xbit_r122_c16 bl[16] br[16] wl[122] vdd gnd cell_6t
Xbit_r123_c16 bl[16] br[16] wl[123] vdd gnd cell_6t
Xbit_r124_c16 bl[16] br[16] wl[124] vdd gnd cell_6t
Xbit_r125_c16 bl[16] br[16] wl[125] vdd gnd cell_6t
Xbit_r126_c16 bl[16] br[16] wl[126] vdd gnd cell_6t
Xbit_r127_c16 bl[16] br[16] wl[127] vdd gnd cell_6t
Xbit_r0_c17 bl[17] br[17] wl[0] vdd gnd cell_6t
Xbit_r1_c17 bl[17] br[17] wl[1] vdd gnd cell_6t
Xbit_r2_c17 bl[17] br[17] wl[2] vdd gnd cell_6t
Xbit_r3_c17 bl[17] br[17] wl[3] vdd gnd cell_6t
Xbit_r4_c17 bl[17] br[17] wl[4] vdd gnd cell_6t
Xbit_r5_c17 bl[17] br[17] wl[5] vdd gnd cell_6t
Xbit_r6_c17 bl[17] br[17] wl[6] vdd gnd cell_6t
Xbit_r7_c17 bl[17] br[17] wl[7] vdd gnd cell_6t
Xbit_r8_c17 bl[17] br[17] wl[8] vdd gnd cell_6t
Xbit_r9_c17 bl[17] br[17] wl[9] vdd gnd cell_6t
Xbit_r10_c17 bl[17] br[17] wl[10] vdd gnd cell_6t
Xbit_r11_c17 bl[17] br[17] wl[11] vdd gnd cell_6t
Xbit_r12_c17 bl[17] br[17] wl[12] vdd gnd cell_6t
Xbit_r13_c17 bl[17] br[17] wl[13] vdd gnd cell_6t
Xbit_r14_c17 bl[17] br[17] wl[14] vdd gnd cell_6t
Xbit_r15_c17 bl[17] br[17] wl[15] vdd gnd cell_6t
Xbit_r16_c17 bl[17] br[17] wl[16] vdd gnd cell_6t
Xbit_r17_c17 bl[17] br[17] wl[17] vdd gnd cell_6t
Xbit_r18_c17 bl[17] br[17] wl[18] vdd gnd cell_6t
Xbit_r19_c17 bl[17] br[17] wl[19] vdd gnd cell_6t
Xbit_r20_c17 bl[17] br[17] wl[20] vdd gnd cell_6t
Xbit_r21_c17 bl[17] br[17] wl[21] vdd gnd cell_6t
Xbit_r22_c17 bl[17] br[17] wl[22] vdd gnd cell_6t
Xbit_r23_c17 bl[17] br[17] wl[23] vdd gnd cell_6t
Xbit_r24_c17 bl[17] br[17] wl[24] vdd gnd cell_6t
Xbit_r25_c17 bl[17] br[17] wl[25] vdd gnd cell_6t
Xbit_r26_c17 bl[17] br[17] wl[26] vdd gnd cell_6t
Xbit_r27_c17 bl[17] br[17] wl[27] vdd gnd cell_6t
Xbit_r28_c17 bl[17] br[17] wl[28] vdd gnd cell_6t
Xbit_r29_c17 bl[17] br[17] wl[29] vdd gnd cell_6t
Xbit_r30_c17 bl[17] br[17] wl[30] vdd gnd cell_6t
Xbit_r31_c17 bl[17] br[17] wl[31] vdd gnd cell_6t
Xbit_r32_c17 bl[17] br[17] wl[32] vdd gnd cell_6t
Xbit_r33_c17 bl[17] br[17] wl[33] vdd gnd cell_6t
Xbit_r34_c17 bl[17] br[17] wl[34] vdd gnd cell_6t
Xbit_r35_c17 bl[17] br[17] wl[35] vdd gnd cell_6t
Xbit_r36_c17 bl[17] br[17] wl[36] vdd gnd cell_6t
Xbit_r37_c17 bl[17] br[17] wl[37] vdd gnd cell_6t
Xbit_r38_c17 bl[17] br[17] wl[38] vdd gnd cell_6t
Xbit_r39_c17 bl[17] br[17] wl[39] vdd gnd cell_6t
Xbit_r40_c17 bl[17] br[17] wl[40] vdd gnd cell_6t
Xbit_r41_c17 bl[17] br[17] wl[41] vdd gnd cell_6t
Xbit_r42_c17 bl[17] br[17] wl[42] vdd gnd cell_6t
Xbit_r43_c17 bl[17] br[17] wl[43] vdd gnd cell_6t
Xbit_r44_c17 bl[17] br[17] wl[44] vdd gnd cell_6t
Xbit_r45_c17 bl[17] br[17] wl[45] vdd gnd cell_6t
Xbit_r46_c17 bl[17] br[17] wl[46] vdd gnd cell_6t
Xbit_r47_c17 bl[17] br[17] wl[47] vdd gnd cell_6t
Xbit_r48_c17 bl[17] br[17] wl[48] vdd gnd cell_6t
Xbit_r49_c17 bl[17] br[17] wl[49] vdd gnd cell_6t
Xbit_r50_c17 bl[17] br[17] wl[50] vdd gnd cell_6t
Xbit_r51_c17 bl[17] br[17] wl[51] vdd gnd cell_6t
Xbit_r52_c17 bl[17] br[17] wl[52] vdd gnd cell_6t
Xbit_r53_c17 bl[17] br[17] wl[53] vdd gnd cell_6t
Xbit_r54_c17 bl[17] br[17] wl[54] vdd gnd cell_6t
Xbit_r55_c17 bl[17] br[17] wl[55] vdd gnd cell_6t
Xbit_r56_c17 bl[17] br[17] wl[56] vdd gnd cell_6t
Xbit_r57_c17 bl[17] br[17] wl[57] vdd gnd cell_6t
Xbit_r58_c17 bl[17] br[17] wl[58] vdd gnd cell_6t
Xbit_r59_c17 bl[17] br[17] wl[59] vdd gnd cell_6t
Xbit_r60_c17 bl[17] br[17] wl[60] vdd gnd cell_6t
Xbit_r61_c17 bl[17] br[17] wl[61] vdd gnd cell_6t
Xbit_r62_c17 bl[17] br[17] wl[62] vdd gnd cell_6t
Xbit_r63_c17 bl[17] br[17] wl[63] vdd gnd cell_6t
Xbit_r64_c17 bl[17] br[17] wl[64] vdd gnd cell_6t
Xbit_r65_c17 bl[17] br[17] wl[65] vdd gnd cell_6t
Xbit_r66_c17 bl[17] br[17] wl[66] vdd gnd cell_6t
Xbit_r67_c17 bl[17] br[17] wl[67] vdd gnd cell_6t
Xbit_r68_c17 bl[17] br[17] wl[68] vdd gnd cell_6t
Xbit_r69_c17 bl[17] br[17] wl[69] vdd gnd cell_6t
Xbit_r70_c17 bl[17] br[17] wl[70] vdd gnd cell_6t
Xbit_r71_c17 bl[17] br[17] wl[71] vdd gnd cell_6t
Xbit_r72_c17 bl[17] br[17] wl[72] vdd gnd cell_6t
Xbit_r73_c17 bl[17] br[17] wl[73] vdd gnd cell_6t
Xbit_r74_c17 bl[17] br[17] wl[74] vdd gnd cell_6t
Xbit_r75_c17 bl[17] br[17] wl[75] vdd gnd cell_6t
Xbit_r76_c17 bl[17] br[17] wl[76] vdd gnd cell_6t
Xbit_r77_c17 bl[17] br[17] wl[77] vdd gnd cell_6t
Xbit_r78_c17 bl[17] br[17] wl[78] vdd gnd cell_6t
Xbit_r79_c17 bl[17] br[17] wl[79] vdd gnd cell_6t
Xbit_r80_c17 bl[17] br[17] wl[80] vdd gnd cell_6t
Xbit_r81_c17 bl[17] br[17] wl[81] vdd gnd cell_6t
Xbit_r82_c17 bl[17] br[17] wl[82] vdd gnd cell_6t
Xbit_r83_c17 bl[17] br[17] wl[83] vdd gnd cell_6t
Xbit_r84_c17 bl[17] br[17] wl[84] vdd gnd cell_6t
Xbit_r85_c17 bl[17] br[17] wl[85] vdd gnd cell_6t
Xbit_r86_c17 bl[17] br[17] wl[86] vdd gnd cell_6t
Xbit_r87_c17 bl[17] br[17] wl[87] vdd gnd cell_6t
Xbit_r88_c17 bl[17] br[17] wl[88] vdd gnd cell_6t
Xbit_r89_c17 bl[17] br[17] wl[89] vdd gnd cell_6t
Xbit_r90_c17 bl[17] br[17] wl[90] vdd gnd cell_6t
Xbit_r91_c17 bl[17] br[17] wl[91] vdd gnd cell_6t
Xbit_r92_c17 bl[17] br[17] wl[92] vdd gnd cell_6t
Xbit_r93_c17 bl[17] br[17] wl[93] vdd gnd cell_6t
Xbit_r94_c17 bl[17] br[17] wl[94] vdd gnd cell_6t
Xbit_r95_c17 bl[17] br[17] wl[95] vdd gnd cell_6t
Xbit_r96_c17 bl[17] br[17] wl[96] vdd gnd cell_6t
Xbit_r97_c17 bl[17] br[17] wl[97] vdd gnd cell_6t
Xbit_r98_c17 bl[17] br[17] wl[98] vdd gnd cell_6t
Xbit_r99_c17 bl[17] br[17] wl[99] vdd gnd cell_6t
Xbit_r100_c17 bl[17] br[17] wl[100] vdd gnd cell_6t
Xbit_r101_c17 bl[17] br[17] wl[101] vdd gnd cell_6t
Xbit_r102_c17 bl[17] br[17] wl[102] vdd gnd cell_6t
Xbit_r103_c17 bl[17] br[17] wl[103] vdd gnd cell_6t
Xbit_r104_c17 bl[17] br[17] wl[104] vdd gnd cell_6t
Xbit_r105_c17 bl[17] br[17] wl[105] vdd gnd cell_6t
Xbit_r106_c17 bl[17] br[17] wl[106] vdd gnd cell_6t
Xbit_r107_c17 bl[17] br[17] wl[107] vdd gnd cell_6t
Xbit_r108_c17 bl[17] br[17] wl[108] vdd gnd cell_6t
Xbit_r109_c17 bl[17] br[17] wl[109] vdd gnd cell_6t
Xbit_r110_c17 bl[17] br[17] wl[110] vdd gnd cell_6t
Xbit_r111_c17 bl[17] br[17] wl[111] vdd gnd cell_6t
Xbit_r112_c17 bl[17] br[17] wl[112] vdd gnd cell_6t
Xbit_r113_c17 bl[17] br[17] wl[113] vdd gnd cell_6t
Xbit_r114_c17 bl[17] br[17] wl[114] vdd gnd cell_6t
Xbit_r115_c17 bl[17] br[17] wl[115] vdd gnd cell_6t
Xbit_r116_c17 bl[17] br[17] wl[116] vdd gnd cell_6t
Xbit_r117_c17 bl[17] br[17] wl[117] vdd gnd cell_6t
Xbit_r118_c17 bl[17] br[17] wl[118] vdd gnd cell_6t
Xbit_r119_c17 bl[17] br[17] wl[119] vdd gnd cell_6t
Xbit_r120_c17 bl[17] br[17] wl[120] vdd gnd cell_6t
Xbit_r121_c17 bl[17] br[17] wl[121] vdd gnd cell_6t
Xbit_r122_c17 bl[17] br[17] wl[122] vdd gnd cell_6t
Xbit_r123_c17 bl[17] br[17] wl[123] vdd gnd cell_6t
Xbit_r124_c17 bl[17] br[17] wl[124] vdd gnd cell_6t
Xbit_r125_c17 bl[17] br[17] wl[125] vdd gnd cell_6t
Xbit_r126_c17 bl[17] br[17] wl[126] vdd gnd cell_6t
Xbit_r127_c17 bl[17] br[17] wl[127] vdd gnd cell_6t
Xbit_r0_c18 bl[18] br[18] wl[0] vdd gnd cell_6t
Xbit_r1_c18 bl[18] br[18] wl[1] vdd gnd cell_6t
Xbit_r2_c18 bl[18] br[18] wl[2] vdd gnd cell_6t
Xbit_r3_c18 bl[18] br[18] wl[3] vdd gnd cell_6t
Xbit_r4_c18 bl[18] br[18] wl[4] vdd gnd cell_6t
Xbit_r5_c18 bl[18] br[18] wl[5] vdd gnd cell_6t
Xbit_r6_c18 bl[18] br[18] wl[6] vdd gnd cell_6t
Xbit_r7_c18 bl[18] br[18] wl[7] vdd gnd cell_6t
Xbit_r8_c18 bl[18] br[18] wl[8] vdd gnd cell_6t
Xbit_r9_c18 bl[18] br[18] wl[9] vdd gnd cell_6t
Xbit_r10_c18 bl[18] br[18] wl[10] vdd gnd cell_6t
Xbit_r11_c18 bl[18] br[18] wl[11] vdd gnd cell_6t
Xbit_r12_c18 bl[18] br[18] wl[12] vdd gnd cell_6t
Xbit_r13_c18 bl[18] br[18] wl[13] vdd gnd cell_6t
Xbit_r14_c18 bl[18] br[18] wl[14] vdd gnd cell_6t
Xbit_r15_c18 bl[18] br[18] wl[15] vdd gnd cell_6t
Xbit_r16_c18 bl[18] br[18] wl[16] vdd gnd cell_6t
Xbit_r17_c18 bl[18] br[18] wl[17] vdd gnd cell_6t
Xbit_r18_c18 bl[18] br[18] wl[18] vdd gnd cell_6t
Xbit_r19_c18 bl[18] br[18] wl[19] vdd gnd cell_6t
Xbit_r20_c18 bl[18] br[18] wl[20] vdd gnd cell_6t
Xbit_r21_c18 bl[18] br[18] wl[21] vdd gnd cell_6t
Xbit_r22_c18 bl[18] br[18] wl[22] vdd gnd cell_6t
Xbit_r23_c18 bl[18] br[18] wl[23] vdd gnd cell_6t
Xbit_r24_c18 bl[18] br[18] wl[24] vdd gnd cell_6t
Xbit_r25_c18 bl[18] br[18] wl[25] vdd gnd cell_6t
Xbit_r26_c18 bl[18] br[18] wl[26] vdd gnd cell_6t
Xbit_r27_c18 bl[18] br[18] wl[27] vdd gnd cell_6t
Xbit_r28_c18 bl[18] br[18] wl[28] vdd gnd cell_6t
Xbit_r29_c18 bl[18] br[18] wl[29] vdd gnd cell_6t
Xbit_r30_c18 bl[18] br[18] wl[30] vdd gnd cell_6t
Xbit_r31_c18 bl[18] br[18] wl[31] vdd gnd cell_6t
Xbit_r32_c18 bl[18] br[18] wl[32] vdd gnd cell_6t
Xbit_r33_c18 bl[18] br[18] wl[33] vdd gnd cell_6t
Xbit_r34_c18 bl[18] br[18] wl[34] vdd gnd cell_6t
Xbit_r35_c18 bl[18] br[18] wl[35] vdd gnd cell_6t
Xbit_r36_c18 bl[18] br[18] wl[36] vdd gnd cell_6t
Xbit_r37_c18 bl[18] br[18] wl[37] vdd gnd cell_6t
Xbit_r38_c18 bl[18] br[18] wl[38] vdd gnd cell_6t
Xbit_r39_c18 bl[18] br[18] wl[39] vdd gnd cell_6t
Xbit_r40_c18 bl[18] br[18] wl[40] vdd gnd cell_6t
Xbit_r41_c18 bl[18] br[18] wl[41] vdd gnd cell_6t
Xbit_r42_c18 bl[18] br[18] wl[42] vdd gnd cell_6t
Xbit_r43_c18 bl[18] br[18] wl[43] vdd gnd cell_6t
Xbit_r44_c18 bl[18] br[18] wl[44] vdd gnd cell_6t
Xbit_r45_c18 bl[18] br[18] wl[45] vdd gnd cell_6t
Xbit_r46_c18 bl[18] br[18] wl[46] vdd gnd cell_6t
Xbit_r47_c18 bl[18] br[18] wl[47] vdd gnd cell_6t
Xbit_r48_c18 bl[18] br[18] wl[48] vdd gnd cell_6t
Xbit_r49_c18 bl[18] br[18] wl[49] vdd gnd cell_6t
Xbit_r50_c18 bl[18] br[18] wl[50] vdd gnd cell_6t
Xbit_r51_c18 bl[18] br[18] wl[51] vdd gnd cell_6t
Xbit_r52_c18 bl[18] br[18] wl[52] vdd gnd cell_6t
Xbit_r53_c18 bl[18] br[18] wl[53] vdd gnd cell_6t
Xbit_r54_c18 bl[18] br[18] wl[54] vdd gnd cell_6t
Xbit_r55_c18 bl[18] br[18] wl[55] vdd gnd cell_6t
Xbit_r56_c18 bl[18] br[18] wl[56] vdd gnd cell_6t
Xbit_r57_c18 bl[18] br[18] wl[57] vdd gnd cell_6t
Xbit_r58_c18 bl[18] br[18] wl[58] vdd gnd cell_6t
Xbit_r59_c18 bl[18] br[18] wl[59] vdd gnd cell_6t
Xbit_r60_c18 bl[18] br[18] wl[60] vdd gnd cell_6t
Xbit_r61_c18 bl[18] br[18] wl[61] vdd gnd cell_6t
Xbit_r62_c18 bl[18] br[18] wl[62] vdd gnd cell_6t
Xbit_r63_c18 bl[18] br[18] wl[63] vdd gnd cell_6t
Xbit_r64_c18 bl[18] br[18] wl[64] vdd gnd cell_6t
Xbit_r65_c18 bl[18] br[18] wl[65] vdd gnd cell_6t
Xbit_r66_c18 bl[18] br[18] wl[66] vdd gnd cell_6t
Xbit_r67_c18 bl[18] br[18] wl[67] vdd gnd cell_6t
Xbit_r68_c18 bl[18] br[18] wl[68] vdd gnd cell_6t
Xbit_r69_c18 bl[18] br[18] wl[69] vdd gnd cell_6t
Xbit_r70_c18 bl[18] br[18] wl[70] vdd gnd cell_6t
Xbit_r71_c18 bl[18] br[18] wl[71] vdd gnd cell_6t
Xbit_r72_c18 bl[18] br[18] wl[72] vdd gnd cell_6t
Xbit_r73_c18 bl[18] br[18] wl[73] vdd gnd cell_6t
Xbit_r74_c18 bl[18] br[18] wl[74] vdd gnd cell_6t
Xbit_r75_c18 bl[18] br[18] wl[75] vdd gnd cell_6t
Xbit_r76_c18 bl[18] br[18] wl[76] vdd gnd cell_6t
Xbit_r77_c18 bl[18] br[18] wl[77] vdd gnd cell_6t
Xbit_r78_c18 bl[18] br[18] wl[78] vdd gnd cell_6t
Xbit_r79_c18 bl[18] br[18] wl[79] vdd gnd cell_6t
Xbit_r80_c18 bl[18] br[18] wl[80] vdd gnd cell_6t
Xbit_r81_c18 bl[18] br[18] wl[81] vdd gnd cell_6t
Xbit_r82_c18 bl[18] br[18] wl[82] vdd gnd cell_6t
Xbit_r83_c18 bl[18] br[18] wl[83] vdd gnd cell_6t
Xbit_r84_c18 bl[18] br[18] wl[84] vdd gnd cell_6t
Xbit_r85_c18 bl[18] br[18] wl[85] vdd gnd cell_6t
Xbit_r86_c18 bl[18] br[18] wl[86] vdd gnd cell_6t
Xbit_r87_c18 bl[18] br[18] wl[87] vdd gnd cell_6t
Xbit_r88_c18 bl[18] br[18] wl[88] vdd gnd cell_6t
Xbit_r89_c18 bl[18] br[18] wl[89] vdd gnd cell_6t
Xbit_r90_c18 bl[18] br[18] wl[90] vdd gnd cell_6t
Xbit_r91_c18 bl[18] br[18] wl[91] vdd gnd cell_6t
Xbit_r92_c18 bl[18] br[18] wl[92] vdd gnd cell_6t
Xbit_r93_c18 bl[18] br[18] wl[93] vdd gnd cell_6t
Xbit_r94_c18 bl[18] br[18] wl[94] vdd gnd cell_6t
Xbit_r95_c18 bl[18] br[18] wl[95] vdd gnd cell_6t
Xbit_r96_c18 bl[18] br[18] wl[96] vdd gnd cell_6t
Xbit_r97_c18 bl[18] br[18] wl[97] vdd gnd cell_6t
Xbit_r98_c18 bl[18] br[18] wl[98] vdd gnd cell_6t
Xbit_r99_c18 bl[18] br[18] wl[99] vdd gnd cell_6t
Xbit_r100_c18 bl[18] br[18] wl[100] vdd gnd cell_6t
Xbit_r101_c18 bl[18] br[18] wl[101] vdd gnd cell_6t
Xbit_r102_c18 bl[18] br[18] wl[102] vdd gnd cell_6t
Xbit_r103_c18 bl[18] br[18] wl[103] vdd gnd cell_6t
Xbit_r104_c18 bl[18] br[18] wl[104] vdd gnd cell_6t
Xbit_r105_c18 bl[18] br[18] wl[105] vdd gnd cell_6t
Xbit_r106_c18 bl[18] br[18] wl[106] vdd gnd cell_6t
Xbit_r107_c18 bl[18] br[18] wl[107] vdd gnd cell_6t
Xbit_r108_c18 bl[18] br[18] wl[108] vdd gnd cell_6t
Xbit_r109_c18 bl[18] br[18] wl[109] vdd gnd cell_6t
Xbit_r110_c18 bl[18] br[18] wl[110] vdd gnd cell_6t
Xbit_r111_c18 bl[18] br[18] wl[111] vdd gnd cell_6t
Xbit_r112_c18 bl[18] br[18] wl[112] vdd gnd cell_6t
Xbit_r113_c18 bl[18] br[18] wl[113] vdd gnd cell_6t
Xbit_r114_c18 bl[18] br[18] wl[114] vdd gnd cell_6t
Xbit_r115_c18 bl[18] br[18] wl[115] vdd gnd cell_6t
Xbit_r116_c18 bl[18] br[18] wl[116] vdd gnd cell_6t
Xbit_r117_c18 bl[18] br[18] wl[117] vdd gnd cell_6t
Xbit_r118_c18 bl[18] br[18] wl[118] vdd gnd cell_6t
Xbit_r119_c18 bl[18] br[18] wl[119] vdd gnd cell_6t
Xbit_r120_c18 bl[18] br[18] wl[120] vdd gnd cell_6t
Xbit_r121_c18 bl[18] br[18] wl[121] vdd gnd cell_6t
Xbit_r122_c18 bl[18] br[18] wl[122] vdd gnd cell_6t
Xbit_r123_c18 bl[18] br[18] wl[123] vdd gnd cell_6t
Xbit_r124_c18 bl[18] br[18] wl[124] vdd gnd cell_6t
Xbit_r125_c18 bl[18] br[18] wl[125] vdd gnd cell_6t
Xbit_r126_c18 bl[18] br[18] wl[126] vdd gnd cell_6t
Xbit_r127_c18 bl[18] br[18] wl[127] vdd gnd cell_6t
Xbit_r0_c19 bl[19] br[19] wl[0] vdd gnd cell_6t
Xbit_r1_c19 bl[19] br[19] wl[1] vdd gnd cell_6t
Xbit_r2_c19 bl[19] br[19] wl[2] vdd gnd cell_6t
Xbit_r3_c19 bl[19] br[19] wl[3] vdd gnd cell_6t
Xbit_r4_c19 bl[19] br[19] wl[4] vdd gnd cell_6t
Xbit_r5_c19 bl[19] br[19] wl[5] vdd gnd cell_6t
Xbit_r6_c19 bl[19] br[19] wl[6] vdd gnd cell_6t
Xbit_r7_c19 bl[19] br[19] wl[7] vdd gnd cell_6t
Xbit_r8_c19 bl[19] br[19] wl[8] vdd gnd cell_6t
Xbit_r9_c19 bl[19] br[19] wl[9] vdd gnd cell_6t
Xbit_r10_c19 bl[19] br[19] wl[10] vdd gnd cell_6t
Xbit_r11_c19 bl[19] br[19] wl[11] vdd gnd cell_6t
Xbit_r12_c19 bl[19] br[19] wl[12] vdd gnd cell_6t
Xbit_r13_c19 bl[19] br[19] wl[13] vdd gnd cell_6t
Xbit_r14_c19 bl[19] br[19] wl[14] vdd gnd cell_6t
Xbit_r15_c19 bl[19] br[19] wl[15] vdd gnd cell_6t
Xbit_r16_c19 bl[19] br[19] wl[16] vdd gnd cell_6t
Xbit_r17_c19 bl[19] br[19] wl[17] vdd gnd cell_6t
Xbit_r18_c19 bl[19] br[19] wl[18] vdd gnd cell_6t
Xbit_r19_c19 bl[19] br[19] wl[19] vdd gnd cell_6t
Xbit_r20_c19 bl[19] br[19] wl[20] vdd gnd cell_6t
Xbit_r21_c19 bl[19] br[19] wl[21] vdd gnd cell_6t
Xbit_r22_c19 bl[19] br[19] wl[22] vdd gnd cell_6t
Xbit_r23_c19 bl[19] br[19] wl[23] vdd gnd cell_6t
Xbit_r24_c19 bl[19] br[19] wl[24] vdd gnd cell_6t
Xbit_r25_c19 bl[19] br[19] wl[25] vdd gnd cell_6t
Xbit_r26_c19 bl[19] br[19] wl[26] vdd gnd cell_6t
Xbit_r27_c19 bl[19] br[19] wl[27] vdd gnd cell_6t
Xbit_r28_c19 bl[19] br[19] wl[28] vdd gnd cell_6t
Xbit_r29_c19 bl[19] br[19] wl[29] vdd gnd cell_6t
Xbit_r30_c19 bl[19] br[19] wl[30] vdd gnd cell_6t
Xbit_r31_c19 bl[19] br[19] wl[31] vdd gnd cell_6t
Xbit_r32_c19 bl[19] br[19] wl[32] vdd gnd cell_6t
Xbit_r33_c19 bl[19] br[19] wl[33] vdd gnd cell_6t
Xbit_r34_c19 bl[19] br[19] wl[34] vdd gnd cell_6t
Xbit_r35_c19 bl[19] br[19] wl[35] vdd gnd cell_6t
Xbit_r36_c19 bl[19] br[19] wl[36] vdd gnd cell_6t
Xbit_r37_c19 bl[19] br[19] wl[37] vdd gnd cell_6t
Xbit_r38_c19 bl[19] br[19] wl[38] vdd gnd cell_6t
Xbit_r39_c19 bl[19] br[19] wl[39] vdd gnd cell_6t
Xbit_r40_c19 bl[19] br[19] wl[40] vdd gnd cell_6t
Xbit_r41_c19 bl[19] br[19] wl[41] vdd gnd cell_6t
Xbit_r42_c19 bl[19] br[19] wl[42] vdd gnd cell_6t
Xbit_r43_c19 bl[19] br[19] wl[43] vdd gnd cell_6t
Xbit_r44_c19 bl[19] br[19] wl[44] vdd gnd cell_6t
Xbit_r45_c19 bl[19] br[19] wl[45] vdd gnd cell_6t
Xbit_r46_c19 bl[19] br[19] wl[46] vdd gnd cell_6t
Xbit_r47_c19 bl[19] br[19] wl[47] vdd gnd cell_6t
Xbit_r48_c19 bl[19] br[19] wl[48] vdd gnd cell_6t
Xbit_r49_c19 bl[19] br[19] wl[49] vdd gnd cell_6t
Xbit_r50_c19 bl[19] br[19] wl[50] vdd gnd cell_6t
Xbit_r51_c19 bl[19] br[19] wl[51] vdd gnd cell_6t
Xbit_r52_c19 bl[19] br[19] wl[52] vdd gnd cell_6t
Xbit_r53_c19 bl[19] br[19] wl[53] vdd gnd cell_6t
Xbit_r54_c19 bl[19] br[19] wl[54] vdd gnd cell_6t
Xbit_r55_c19 bl[19] br[19] wl[55] vdd gnd cell_6t
Xbit_r56_c19 bl[19] br[19] wl[56] vdd gnd cell_6t
Xbit_r57_c19 bl[19] br[19] wl[57] vdd gnd cell_6t
Xbit_r58_c19 bl[19] br[19] wl[58] vdd gnd cell_6t
Xbit_r59_c19 bl[19] br[19] wl[59] vdd gnd cell_6t
Xbit_r60_c19 bl[19] br[19] wl[60] vdd gnd cell_6t
Xbit_r61_c19 bl[19] br[19] wl[61] vdd gnd cell_6t
Xbit_r62_c19 bl[19] br[19] wl[62] vdd gnd cell_6t
Xbit_r63_c19 bl[19] br[19] wl[63] vdd gnd cell_6t
Xbit_r64_c19 bl[19] br[19] wl[64] vdd gnd cell_6t
Xbit_r65_c19 bl[19] br[19] wl[65] vdd gnd cell_6t
Xbit_r66_c19 bl[19] br[19] wl[66] vdd gnd cell_6t
Xbit_r67_c19 bl[19] br[19] wl[67] vdd gnd cell_6t
Xbit_r68_c19 bl[19] br[19] wl[68] vdd gnd cell_6t
Xbit_r69_c19 bl[19] br[19] wl[69] vdd gnd cell_6t
Xbit_r70_c19 bl[19] br[19] wl[70] vdd gnd cell_6t
Xbit_r71_c19 bl[19] br[19] wl[71] vdd gnd cell_6t
Xbit_r72_c19 bl[19] br[19] wl[72] vdd gnd cell_6t
Xbit_r73_c19 bl[19] br[19] wl[73] vdd gnd cell_6t
Xbit_r74_c19 bl[19] br[19] wl[74] vdd gnd cell_6t
Xbit_r75_c19 bl[19] br[19] wl[75] vdd gnd cell_6t
Xbit_r76_c19 bl[19] br[19] wl[76] vdd gnd cell_6t
Xbit_r77_c19 bl[19] br[19] wl[77] vdd gnd cell_6t
Xbit_r78_c19 bl[19] br[19] wl[78] vdd gnd cell_6t
Xbit_r79_c19 bl[19] br[19] wl[79] vdd gnd cell_6t
Xbit_r80_c19 bl[19] br[19] wl[80] vdd gnd cell_6t
Xbit_r81_c19 bl[19] br[19] wl[81] vdd gnd cell_6t
Xbit_r82_c19 bl[19] br[19] wl[82] vdd gnd cell_6t
Xbit_r83_c19 bl[19] br[19] wl[83] vdd gnd cell_6t
Xbit_r84_c19 bl[19] br[19] wl[84] vdd gnd cell_6t
Xbit_r85_c19 bl[19] br[19] wl[85] vdd gnd cell_6t
Xbit_r86_c19 bl[19] br[19] wl[86] vdd gnd cell_6t
Xbit_r87_c19 bl[19] br[19] wl[87] vdd gnd cell_6t
Xbit_r88_c19 bl[19] br[19] wl[88] vdd gnd cell_6t
Xbit_r89_c19 bl[19] br[19] wl[89] vdd gnd cell_6t
Xbit_r90_c19 bl[19] br[19] wl[90] vdd gnd cell_6t
Xbit_r91_c19 bl[19] br[19] wl[91] vdd gnd cell_6t
Xbit_r92_c19 bl[19] br[19] wl[92] vdd gnd cell_6t
Xbit_r93_c19 bl[19] br[19] wl[93] vdd gnd cell_6t
Xbit_r94_c19 bl[19] br[19] wl[94] vdd gnd cell_6t
Xbit_r95_c19 bl[19] br[19] wl[95] vdd gnd cell_6t
Xbit_r96_c19 bl[19] br[19] wl[96] vdd gnd cell_6t
Xbit_r97_c19 bl[19] br[19] wl[97] vdd gnd cell_6t
Xbit_r98_c19 bl[19] br[19] wl[98] vdd gnd cell_6t
Xbit_r99_c19 bl[19] br[19] wl[99] vdd gnd cell_6t
Xbit_r100_c19 bl[19] br[19] wl[100] vdd gnd cell_6t
Xbit_r101_c19 bl[19] br[19] wl[101] vdd gnd cell_6t
Xbit_r102_c19 bl[19] br[19] wl[102] vdd gnd cell_6t
Xbit_r103_c19 bl[19] br[19] wl[103] vdd gnd cell_6t
Xbit_r104_c19 bl[19] br[19] wl[104] vdd gnd cell_6t
Xbit_r105_c19 bl[19] br[19] wl[105] vdd gnd cell_6t
Xbit_r106_c19 bl[19] br[19] wl[106] vdd gnd cell_6t
Xbit_r107_c19 bl[19] br[19] wl[107] vdd gnd cell_6t
Xbit_r108_c19 bl[19] br[19] wl[108] vdd gnd cell_6t
Xbit_r109_c19 bl[19] br[19] wl[109] vdd gnd cell_6t
Xbit_r110_c19 bl[19] br[19] wl[110] vdd gnd cell_6t
Xbit_r111_c19 bl[19] br[19] wl[111] vdd gnd cell_6t
Xbit_r112_c19 bl[19] br[19] wl[112] vdd gnd cell_6t
Xbit_r113_c19 bl[19] br[19] wl[113] vdd gnd cell_6t
Xbit_r114_c19 bl[19] br[19] wl[114] vdd gnd cell_6t
Xbit_r115_c19 bl[19] br[19] wl[115] vdd gnd cell_6t
Xbit_r116_c19 bl[19] br[19] wl[116] vdd gnd cell_6t
Xbit_r117_c19 bl[19] br[19] wl[117] vdd gnd cell_6t
Xbit_r118_c19 bl[19] br[19] wl[118] vdd gnd cell_6t
Xbit_r119_c19 bl[19] br[19] wl[119] vdd gnd cell_6t
Xbit_r120_c19 bl[19] br[19] wl[120] vdd gnd cell_6t
Xbit_r121_c19 bl[19] br[19] wl[121] vdd gnd cell_6t
Xbit_r122_c19 bl[19] br[19] wl[122] vdd gnd cell_6t
Xbit_r123_c19 bl[19] br[19] wl[123] vdd gnd cell_6t
Xbit_r124_c19 bl[19] br[19] wl[124] vdd gnd cell_6t
Xbit_r125_c19 bl[19] br[19] wl[125] vdd gnd cell_6t
Xbit_r126_c19 bl[19] br[19] wl[126] vdd gnd cell_6t
Xbit_r127_c19 bl[19] br[19] wl[127] vdd gnd cell_6t
Xbit_r0_c20 bl[20] br[20] wl[0] vdd gnd cell_6t
Xbit_r1_c20 bl[20] br[20] wl[1] vdd gnd cell_6t
Xbit_r2_c20 bl[20] br[20] wl[2] vdd gnd cell_6t
Xbit_r3_c20 bl[20] br[20] wl[3] vdd gnd cell_6t
Xbit_r4_c20 bl[20] br[20] wl[4] vdd gnd cell_6t
Xbit_r5_c20 bl[20] br[20] wl[5] vdd gnd cell_6t
Xbit_r6_c20 bl[20] br[20] wl[6] vdd gnd cell_6t
Xbit_r7_c20 bl[20] br[20] wl[7] vdd gnd cell_6t
Xbit_r8_c20 bl[20] br[20] wl[8] vdd gnd cell_6t
Xbit_r9_c20 bl[20] br[20] wl[9] vdd gnd cell_6t
Xbit_r10_c20 bl[20] br[20] wl[10] vdd gnd cell_6t
Xbit_r11_c20 bl[20] br[20] wl[11] vdd gnd cell_6t
Xbit_r12_c20 bl[20] br[20] wl[12] vdd gnd cell_6t
Xbit_r13_c20 bl[20] br[20] wl[13] vdd gnd cell_6t
Xbit_r14_c20 bl[20] br[20] wl[14] vdd gnd cell_6t
Xbit_r15_c20 bl[20] br[20] wl[15] vdd gnd cell_6t
Xbit_r16_c20 bl[20] br[20] wl[16] vdd gnd cell_6t
Xbit_r17_c20 bl[20] br[20] wl[17] vdd gnd cell_6t
Xbit_r18_c20 bl[20] br[20] wl[18] vdd gnd cell_6t
Xbit_r19_c20 bl[20] br[20] wl[19] vdd gnd cell_6t
Xbit_r20_c20 bl[20] br[20] wl[20] vdd gnd cell_6t
Xbit_r21_c20 bl[20] br[20] wl[21] vdd gnd cell_6t
Xbit_r22_c20 bl[20] br[20] wl[22] vdd gnd cell_6t
Xbit_r23_c20 bl[20] br[20] wl[23] vdd gnd cell_6t
Xbit_r24_c20 bl[20] br[20] wl[24] vdd gnd cell_6t
Xbit_r25_c20 bl[20] br[20] wl[25] vdd gnd cell_6t
Xbit_r26_c20 bl[20] br[20] wl[26] vdd gnd cell_6t
Xbit_r27_c20 bl[20] br[20] wl[27] vdd gnd cell_6t
Xbit_r28_c20 bl[20] br[20] wl[28] vdd gnd cell_6t
Xbit_r29_c20 bl[20] br[20] wl[29] vdd gnd cell_6t
Xbit_r30_c20 bl[20] br[20] wl[30] vdd gnd cell_6t
Xbit_r31_c20 bl[20] br[20] wl[31] vdd gnd cell_6t
Xbit_r32_c20 bl[20] br[20] wl[32] vdd gnd cell_6t
Xbit_r33_c20 bl[20] br[20] wl[33] vdd gnd cell_6t
Xbit_r34_c20 bl[20] br[20] wl[34] vdd gnd cell_6t
Xbit_r35_c20 bl[20] br[20] wl[35] vdd gnd cell_6t
Xbit_r36_c20 bl[20] br[20] wl[36] vdd gnd cell_6t
Xbit_r37_c20 bl[20] br[20] wl[37] vdd gnd cell_6t
Xbit_r38_c20 bl[20] br[20] wl[38] vdd gnd cell_6t
Xbit_r39_c20 bl[20] br[20] wl[39] vdd gnd cell_6t
Xbit_r40_c20 bl[20] br[20] wl[40] vdd gnd cell_6t
Xbit_r41_c20 bl[20] br[20] wl[41] vdd gnd cell_6t
Xbit_r42_c20 bl[20] br[20] wl[42] vdd gnd cell_6t
Xbit_r43_c20 bl[20] br[20] wl[43] vdd gnd cell_6t
Xbit_r44_c20 bl[20] br[20] wl[44] vdd gnd cell_6t
Xbit_r45_c20 bl[20] br[20] wl[45] vdd gnd cell_6t
Xbit_r46_c20 bl[20] br[20] wl[46] vdd gnd cell_6t
Xbit_r47_c20 bl[20] br[20] wl[47] vdd gnd cell_6t
Xbit_r48_c20 bl[20] br[20] wl[48] vdd gnd cell_6t
Xbit_r49_c20 bl[20] br[20] wl[49] vdd gnd cell_6t
Xbit_r50_c20 bl[20] br[20] wl[50] vdd gnd cell_6t
Xbit_r51_c20 bl[20] br[20] wl[51] vdd gnd cell_6t
Xbit_r52_c20 bl[20] br[20] wl[52] vdd gnd cell_6t
Xbit_r53_c20 bl[20] br[20] wl[53] vdd gnd cell_6t
Xbit_r54_c20 bl[20] br[20] wl[54] vdd gnd cell_6t
Xbit_r55_c20 bl[20] br[20] wl[55] vdd gnd cell_6t
Xbit_r56_c20 bl[20] br[20] wl[56] vdd gnd cell_6t
Xbit_r57_c20 bl[20] br[20] wl[57] vdd gnd cell_6t
Xbit_r58_c20 bl[20] br[20] wl[58] vdd gnd cell_6t
Xbit_r59_c20 bl[20] br[20] wl[59] vdd gnd cell_6t
Xbit_r60_c20 bl[20] br[20] wl[60] vdd gnd cell_6t
Xbit_r61_c20 bl[20] br[20] wl[61] vdd gnd cell_6t
Xbit_r62_c20 bl[20] br[20] wl[62] vdd gnd cell_6t
Xbit_r63_c20 bl[20] br[20] wl[63] vdd gnd cell_6t
Xbit_r64_c20 bl[20] br[20] wl[64] vdd gnd cell_6t
Xbit_r65_c20 bl[20] br[20] wl[65] vdd gnd cell_6t
Xbit_r66_c20 bl[20] br[20] wl[66] vdd gnd cell_6t
Xbit_r67_c20 bl[20] br[20] wl[67] vdd gnd cell_6t
Xbit_r68_c20 bl[20] br[20] wl[68] vdd gnd cell_6t
Xbit_r69_c20 bl[20] br[20] wl[69] vdd gnd cell_6t
Xbit_r70_c20 bl[20] br[20] wl[70] vdd gnd cell_6t
Xbit_r71_c20 bl[20] br[20] wl[71] vdd gnd cell_6t
Xbit_r72_c20 bl[20] br[20] wl[72] vdd gnd cell_6t
Xbit_r73_c20 bl[20] br[20] wl[73] vdd gnd cell_6t
Xbit_r74_c20 bl[20] br[20] wl[74] vdd gnd cell_6t
Xbit_r75_c20 bl[20] br[20] wl[75] vdd gnd cell_6t
Xbit_r76_c20 bl[20] br[20] wl[76] vdd gnd cell_6t
Xbit_r77_c20 bl[20] br[20] wl[77] vdd gnd cell_6t
Xbit_r78_c20 bl[20] br[20] wl[78] vdd gnd cell_6t
Xbit_r79_c20 bl[20] br[20] wl[79] vdd gnd cell_6t
Xbit_r80_c20 bl[20] br[20] wl[80] vdd gnd cell_6t
Xbit_r81_c20 bl[20] br[20] wl[81] vdd gnd cell_6t
Xbit_r82_c20 bl[20] br[20] wl[82] vdd gnd cell_6t
Xbit_r83_c20 bl[20] br[20] wl[83] vdd gnd cell_6t
Xbit_r84_c20 bl[20] br[20] wl[84] vdd gnd cell_6t
Xbit_r85_c20 bl[20] br[20] wl[85] vdd gnd cell_6t
Xbit_r86_c20 bl[20] br[20] wl[86] vdd gnd cell_6t
Xbit_r87_c20 bl[20] br[20] wl[87] vdd gnd cell_6t
Xbit_r88_c20 bl[20] br[20] wl[88] vdd gnd cell_6t
Xbit_r89_c20 bl[20] br[20] wl[89] vdd gnd cell_6t
Xbit_r90_c20 bl[20] br[20] wl[90] vdd gnd cell_6t
Xbit_r91_c20 bl[20] br[20] wl[91] vdd gnd cell_6t
Xbit_r92_c20 bl[20] br[20] wl[92] vdd gnd cell_6t
Xbit_r93_c20 bl[20] br[20] wl[93] vdd gnd cell_6t
Xbit_r94_c20 bl[20] br[20] wl[94] vdd gnd cell_6t
Xbit_r95_c20 bl[20] br[20] wl[95] vdd gnd cell_6t
Xbit_r96_c20 bl[20] br[20] wl[96] vdd gnd cell_6t
Xbit_r97_c20 bl[20] br[20] wl[97] vdd gnd cell_6t
Xbit_r98_c20 bl[20] br[20] wl[98] vdd gnd cell_6t
Xbit_r99_c20 bl[20] br[20] wl[99] vdd gnd cell_6t
Xbit_r100_c20 bl[20] br[20] wl[100] vdd gnd cell_6t
Xbit_r101_c20 bl[20] br[20] wl[101] vdd gnd cell_6t
Xbit_r102_c20 bl[20] br[20] wl[102] vdd gnd cell_6t
Xbit_r103_c20 bl[20] br[20] wl[103] vdd gnd cell_6t
Xbit_r104_c20 bl[20] br[20] wl[104] vdd gnd cell_6t
Xbit_r105_c20 bl[20] br[20] wl[105] vdd gnd cell_6t
Xbit_r106_c20 bl[20] br[20] wl[106] vdd gnd cell_6t
Xbit_r107_c20 bl[20] br[20] wl[107] vdd gnd cell_6t
Xbit_r108_c20 bl[20] br[20] wl[108] vdd gnd cell_6t
Xbit_r109_c20 bl[20] br[20] wl[109] vdd gnd cell_6t
Xbit_r110_c20 bl[20] br[20] wl[110] vdd gnd cell_6t
Xbit_r111_c20 bl[20] br[20] wl[111] vdd gnd cell_6t
Xbit_r112_c20 bl[20] br[20] wl[112] vdd gnd cell_6t
Xbit_r113_c20 bl[20] br[20] wl[113] vdd gnd cell_6t
Xbit_r114_c20 bl[20] br[20] wl[114] vdd gnd cell_6t
Xbit_r115_c20 bl[20] br[20] wl[115] vdd gnd cell_6t
Xbit_r116_c20 bl[20] br[20] wl[116] vdd gnd cell_6t
Xbit_r117_c20 bl[20] br[20] wl[117] vdd gnd cell_6t
Xbit_r118_c20 bl[20] br[20] wl[118] vdd gnd cell_6t
Xbit_r119_c20 bl[20] br[20] wl[119] vdd gnd cell_6t
Xbit_r120_c20 bl[20] br[20] wl[120] vdd gnd cell_6t
Xbit_r121_c20 bl[20] br[20] wl[121] vdd gnd cell_6t
Xbit_r122_c20 bl[20] br[20] wl[122] vdd gnd cell_6t
Xbit_r123_c20 bl[20] br[20] wl[123] vdd gnd cell_6t
Xbit_r124_c20 bl[20] br[20] wl[124] vdd gnd cell_6t
Xbit_r125_c20 bl[20] br[20] wl[125] vdd gnd cell_6t
Xbit_r126_c20 bl[20] br[20] wl[126] vdd gnd cell_6t
Xbit_r127_c20 bl[20] br[20] wl[127] vdd gnd cell_6t
Xbit_r0_c21 bl[21] br[21] wl[0] vdd gnd cell_6t
Xbit_r1_c21 bl[21] br[21] wl[1] vdd gnd cell_6t
Xbit_r2_c21 bl[21] br[21] wl[2] vdd gnd cell_6t
Xbit_r3_c21 bl[21] br[21] wl[3] vdd gnd cell_6t
Xbit_r4_c21 bl[21] br[21] wl[4] vdd gnd cell_6t
Xbit_r5_c21 bl[21] br[21] wl[5] vdd gnd cell_6t
Xbit_r6_c21 bl[21] br[21] wl[6] vdd gnd cell_6t
Xbit_r7_c21 bl[21] br[21] wl[7] vdd gnd cell_6t
Xbit_r8_c21 bl[21] br[21] wl[8] vdd gnd cell_6t
Xbit_r9_c21 bl[21] br[21] wl[9] vdd gnd cell_6t
Xbit_r10_c21 bl[21] br[21] wl[10] vdd gnd cell_6t
Xbit_r11_c21 bl[21] br[21] wl[11] vdd gnd cell_6t
Xbit_r12_c21 bl[21] br[21] wl[12] vdd gnd cell_6t
Xbit_r13_c21 bl[21] br[21] wl[13] vdd gnd cell_6t
Xbit_r14_c21 bl[21] br[21] wl[14] vdd gnd cell_6t
Xbit_r15_c21 bl[21] br[21] wl[15] vdd gnd cell_6t
Xbit_r16_c21 bl[21] br[21] wl[16] vdd gnd cell_6t
Xbit_r17_c21 bl[21] br[21] wl[17] vdd gnd cell_6t
Xbit_r18_c21 bl[21] br[21] wl[18] vdd gnd cell_6t
Xbit_r19_c21 bl[21] br[21] wl[19] vdd gnd cell_6t
Xbit_r20_c21 bl[21] br[21] wl[20] vdd gnd cell_6t
Xbit_r21_c21 bl[21] br[21] wl[21] vdd gnd cell_6t
Xbit_r22_c21 bl[21] br[21] wl[22] vdd gnd cell_6t
Xbit_r23_c21 bl[21] br[21] wl[23] vdd gnd cell_6t
Xbit_r24_c21 bl[21] br[21] wl[24] vdd gnd cell_6t
Xbit_r25_c21 bl[21] br[21] wl[25] vdd gnd cell_6t
Xbit_r26_c21 bl[21] br[21] wl[26] vdd gnd cell_6t
Xbit_r27_c21 bl[21] br[21] wl[27] vdd gnd cell_6t
Xbit_r28_c21 bl[21] br[21] wl[28] vdd gnd cell_6t
Xbit_r29_c21 bl[21] br[21] wl[29] vdd gnd cell_6t
Xbit_r30_c21 bl[21] br[21] wl[30] vdd gnd cell_6t
Xbit_r31_c21 bl[21] br[21] wl[31] vdd gnd cell_6t
Xbit_r32_c21 bl[21] br[21] wl[32] vdd gnd cell_6t
Xbit_r33_c21 bl[21] br[21] wl[33] vdd gnd cell_6t
Xbit_r34_c21 bl[21] br[21] wl[34] vdd gnd cell_6t
Xbit_r35_c21 bl[21] br[21] wl[35] vdd gnd cell_6t
Xbit_r36_c21 bl[21] br[21] wl[36] vdd gnd cell_6t
Xbit_r37_c21 bl[21] br[21] wl[37] vdd gnd cell_6t
Xbit_r38_c21 bl[21] br[21] wl[38] vdd gnd cell_6t
Xbit_r39_c21 bl[21] br[21] wl[39] vdd gnd cell_6t
Xbit_r40_c21 bl[21] br[21] wl[40] vdd gnd cell_6t
Xbit_r41_c21 bl[21] br[21] wl[41] vdd gnd cell_6t
Xbit_r42_c21 bl[21] br[21] wl[42] vdd gnd cell_6t
Xbit_r43_c21 bl[21] br[21] wl[43] vdd gnd cell_6t
Xbit_r44_c21 bl[21] br[21] wl[44] vdd gnd cell_6t
Xbit_r45_c21 bl[21] br[21] wl[45] vdd gnd cell_6t
Xbit_r46_c21 bl[21] br[21] wl[46] vdd gnd cell_6t
Xbit_r47_c21 bl[21] br[21] wl[47] vdd gnd cell_6t
Xbit_r48_c21 bl[21] br[21] wl[48] vdd gnd cell_6t
Xbit_r49_c21 bl[21] br[21] wl[49] vdd gnd cell_6t
Xbit_r50_c21 bl[21] br[21] wl[50] vdd gnd cell_6t
Xbit_r51_c21 bl[21] br[21] wl[51] vdd gnd cell_6t
Xbit_r52_c21 bl[21] br[21] wl[52] vdd gnd cell_6t
Xbit_r53_c21 bl[21] br[21] wl[53] vdd gnd cell_6t
Xbit_r54_c21 bl[21] br[21] wl[54] vdd gnd cell_6t
Xbit_r55_c21 bl[21] br[21] wl[55] vdd gnd cell_6t
Xbit_r56_c21 bl[21] br[21] wl[56] vdd gnd cell_6t
Xbit_r57_c21 bl[21] br[21] wl[57] vdd gnd cell_6t
Xbit_r58_c21 bl[21] br[21] wl[58] vdd gnd cell_6t
Xbit_r59_c21 bl[21] br[21] wl[59] vdd gnd cell_6t
Xbit_r60_c21 bl[21] br[21] wl[60] vdd gnd cell_6t
Xbit_r61_c21 bl[21] br[21] wl[61] vdd gnd cell_6t
Xbit_r62_c21 bl[21] br[21] wl[62] vdd gnd cell_6t
Xbit_r63_c21 bl[21] br[21] wl[63] vdd gnd cell_6t
Xbit_r64_c21 bl[21] br[21] wl[64] vdd gnd cell_6t
Xbit_r65_c21 bl[21] br[21] wl[65] vdd gnd cell_6t
Xbit_r66_c21 bl[21] br[21] wl[66] vdd gnd cell_6t
Xbit_r67_c21 bl[21] br[21] wl[67] vdd gnd cell_6t
Xbit_r68_c21 bl[21] br[21] wl[68] vdd gnd cell_6t
Xbit_r69_c21 bl[21] br[21] wl[69] vdd gnd cell_6t
Xbit_r70_c21 bl[21] br[21] wl[70] vdd gnd cell_6t
Xbit_r71_c21 bl[21] br[21] wl[71] vdd gnd cell_6t
Xbit_r72_c21 bl[21] br[21] wl[72] vdd gnd cell_6t
Xbit_r73_c21 bl[21] br[21] wl[73] vdd gnd cell_6t
Xbit_r74_c21 bl[21] br[21] wl[74] vdd gnd cell_6t
Xbit_r75_c21 bl[21] br[21] wl[75] vdd gnd cell_6t
Xbit_r76_c21 bl[21] br[21] wl[76] vdd gnd cell_6t
Xbit_r77_c21 bl[21] br[21] wl[77] vdd gnd cell_6t
Xbit_r78_c21 bl[21] br[21] wl[78] vdd gnd cell_6t
Xbit_r79_c21 bl[21] br[21] wl[79] vdd gnd cell_6t
Xbit_r80_c21 bl[21] br[21] wl[80] vdd gnd cell_6t
Xbit_r81_c21 bl[21] br[21] wl[81] vdd gnd cell_6t
Xbit_r82_c21 bl[21] br[21] wl[82] vdd gnd cell_6t
Xbit_r83_c21 bl[21] br[21] wl[83] vdd gnd cell_6t
Xbit_r84_c21 bl[21] br[21] wl[84] vdd gnd cell_6t
Xbit_r85_c21 bl[21] br[21] wl[85] vdd gnd cell_6t
Xbit_r86_c21 bl[21] br[21] wl[86] vdd gnd cell_6t
Xbit_r87_c21 bl[21] br[21] wl[87] vdd gnd cell_6t
Xbit_r88_c21 bl[21] br[21] wl[88] vdd gnd cell_6t
Xbit_r89_c21 bl[21] br[21] wl[89] vdd gnd cell_6t
Xbit_r90_c21 bl[21] br[21] wl[90] vdd gnd cell_6t
Xbit_r91_c21 bl[21] br[21] wl[91] vdd gnd cell_6t
Xbit_r92_c21 bl[21] br[21] wl[92] vdd gnd cell_6t
Xbit_r93_c21 bl[21] br[21] wl[93] vdd gnd cell_6t
Xbit_r94_c21 bl[21] br[21] wl[94] vdd gnd cell_6t
Xbit_r95_c21 bl[21] br[21] wl[95] vdd gnd cell_6t
Xbit_r96_c21 bl[21] br[21] wl[96] vdd gnd cell_6t
Xbit_r97_c21 bl[21] br[21] wl[97] vdd gnd cell_6t
Xbit_r98_c21 bl[21] br[21] wl[98] vdd gnd cell_6t
Xbit_r99_c21 bl[21] br[21] wl[99] vdd gnd cell_6t
Xbit_r100_c21 bl[21] br[21] wl[100] vdd gnd cell_6t
Xbit_r101_c21 bl[21] br[21] wl[101] vdd gnd cell_6t
Xbit_r102_c21 bl[21] br[21] wl[102] vdd gnd cell_6t
Xbit_r103_c21 bl[21] br[21] wl[103] vdd gnd cell_6t
Xbit_r104_c21 bl[21] br[21] wl[104] vdd gnd cell_6t
Xbit_r105_c21 bl[21] br[21] wl[105] vdd gnd cell_6t
Xbit_r106_c21 bl[21] br[21] wl[106] vdd gnd cell_6t
Xbit_r107_c21 bl[21] br[21] wl[107] vdd gnd cell_6t
Xbit_r108_c21 bl[21] br[21] wl[108] vdd gnd cell_6t
Xbit_r109_c21 bl[21] br[21] wl[109] vdd gnd cell_6t
Xbit_r110_c21 bl[21] br[21] wl[110] vdd gnd cell_6t
Xbit_r111_c21 bl[21] br[21] wl[111] vdd gnd cell_6t
Xbit_r112_c21 bl[21] br[21] wl[112] vdd gnd cell_6t
Xbit_r113_c21 bl[21] br[21] wl[113] vdd gnd cell_6t
Xbit_r114_c21 bl[21] br[21] wl[114] vdd gnd cell_6t
Xbit_r115_c21 bl[21] br[21] wl[115] vdd gnd cell_6t
Xbit_r116_c21 bl[21] br[21] wl[116] vdd gnd cell_6t
Xbit_r117_c21 bl[21] br[21] wl[117] vdd gnd cell_6t
Xbit_r118_c21 bl[21] br[21] wl[118] vdd gnd cell_6t
Xbit_r119_c21 bl[21] br[21] wl[119] vdd gnd cell_6t
Xbit_r120_c21 bl[21] br[21] wl[120] vdd gnd cell_6t
Xbit_r121_c21 bl[21] br[21] wl[121] vdd gnd cell_6t
Xbit_r122_c21 bl[21] br[21] wl[122] vdd gnd cell_6t
Xbit_r123_c21 bl[21] br[21] wl[123] vdd gnd cell_6t
Xbit_r124_c21 bl[21] br[21] wl[124] vdd gnd cell_6t
Xbit_r125_c21 bl[21] br[21] wl[125] vdd gnd cell_6t
Xbit_r126_c21 bl[21] br[21] wl[126] vdd gnd cell_6t
Xbit_r127_c21 bl[21] br[21] wl[127] vdd gnd cell_6t
Xbit_r0_c22 bl[22] br[22] wl[0] vdd gnd cell_6t
Xbit_r1_c22 bl[22] br[22] wl[1] vdd gnd cell_6t
Xbit_r2_c22 bl[22] br[22] wl[2] vdd gnd cell_6t
Xbit_r3_c22 bl[22] br[22] wl[3] vdd gnd cell_6t
Xbit_r4_c22 bl[22] br[22] wl[4] vdd gnd cell_6t
Xbit_r5_c22 bl[22] br[22] wl[5] vdd gnd cell_6t
Xbit_r6_c22 bl[22] br[22] wl[6] vdd gnd cell_6t
Xbit_r7_c22 bl[22] br[22] wl[7] vdd gnd cell_6t
Xbit_r8_c22 bl[22] br[22] wl[8] vdd gnd cell_6t
Xbit_r9_c22 bl[22] br[22] wl[9] vdd gnd cell_6t
Xbit_r10_c22 bl[22] br[22] wl[10] vdd gnd cell_6t
Xbit_r11_c22 bl[22] br[22] wl[11] vdd gnd cell_6t
Xbit_r12_c22 bl[22] br[22] wl[12] vdd gnd cell_6t
Xbit_r13_c22 bl[22] br[22] wl[13] vdd gnd cell_6t
Xbit_r14_c22 bl[22] br[22] wl[14] vdd gnd cell_6t
Xbit_r15_c22 bl[22] br[22] wl[15] vdd gnd cell_6t
Xbit_r16_c22 bl[22] br[22] wl[16] vdd gnd cell_6t
Xbit_r17_c22 bl[22] br[22] wl[17] vdd gnd cell_6t
Xbit_r18_c22 bl[22] br[22] wl[18] vdd gnd cell_6t
Xbit_r19_c22 bl[22] br[22] wl[19] vdd gnd cell_6t
Xbit_r20_c22 bl[22] br[22] wl[20] vdd gnd cell_6t
Xbit_r21_c22 bl[22] br[22] wl[21] vdd gnd cell_6t
Xbit_r22_c22 bl[22] br[22] wl[22] vdd gnd cell_6t
Xbit_r23_c22 bl[22] br[22] wl[23] vdd gnd cell_6t
Xbit_r24_c22 bl[22] br[22] wl[24] vdd gnd cell_6t
Xbit_r25_c22 bl[22] br[22] wl[25] vdd gnd cell_6t
Xbit_r26_c22 bl[22] br[22] wl[26] vdd gnd cell_6t
Xbit_r27_c22 bl[22] br[22] wl[27] vdd gnd cell_6t
Xbit_r28_c22 bl[22] br[22] wl[28] vdd gnd cell_6t
Xbit_r29_c22 bl[22] br[22] wl[29] vdd gnd cell_6t
Xbit_r30_c22 bl[22] br[22] wl[30] vdd gnd cell_6t
Xbit_r31_c22 bl[22] br[22] wl[31] vdd gnd cell_6t
Xbit_r32_c22 bl[22] br[22] wl[32] vdd gnd cell_6t
Xbit_r33_c22 bl[22] br[22] wl[33] vdd gnd cell_6t
Xbit_r34_c22 bl[22] br[22] wl[34] vdd gnd cell_6t
Xbit_r35_c22 bl[22] br[22] wl[35] vdd gnd cell_6t
Xbit_r36_c22 bl[22] br[22] wl[36] vdd gnd cell_6t
Xbit_r37_c22 bl[22] br[22] wl[37] vdd gnd cell_6t
Xbit_r38_c22 bl[22] br[22] wl[38] vdd gnd cell_6t
Xbit_r39_c22 bl[22] br[22] wl[39] vdd gnd cell_6t
Xbit_r40_c22 bl[22] br[22] wl[40] vdd gnd cell_6t
Xbit_r41_c22 bl[22] br[22] wl[41] vdd gnd cell_6t
Xbit_r42_c22 bl[22] br[22] wl[42] vdd gnd cell_6t
Xbit_r43_c22 bl[22] br[22] wl[43] vdd gnd cell_6t
Xbit_r44_c22 bl[22] br[22] wl[44] vdd gnd cell_6t
Xbit_r45_c22 bl[22] br[22] wl[45] vdd gnd cell_6t
Xbit_r46_c22 bl[22] br[22] wl[46] vdd gnd cell_6t
Xbit_r47_c22 bl[22] br[22] wl[47] vdd gnd cell_6t
Xbit_r48_c22 bl[22] br[22] wl[48] vdd gnd cell_6t
Xbit_r49_c22 bl[22] br[22] wl[49] vdd gnd cell_6t
Xbit_r50_c22 bl[22] br[22] wl[50] vdd gnd cell_6t
Xbit_r51_c22 bl[22] br[22] wl[51] vdd gnd cell_6t
Xbit_r52_c22 bl[22] br[22] wl[52] vdd gnd cell_6t
Xbit_r53_c22 bl[22] br[22] wl[53] vdd gnd cell_6t
Xbit_r54_c22 bl[22] br[22] wl[54] vdd gnd cell_6t
Xbit_r55_c22 bl[22] br[22] wl[55] vdd gnd cell_6t
Xbit_r56_c22 bl[22] br[22] wl[56] vdd gnd cell_6t
Xbit_r57_c22 bl[22] br[22] wl[57] vdd gnd cell_6t
Xbit_r58_c22 bl[22] br[22] wl[58] vdd gnd cell_6t
Xbit_r59_c22 bl[22] br[22] wl[59] vdd gnd cell_6t
Xbit_r60_c22 bl[22] br[22] wl[60] vdd gnd cell_6t
Xbit_r61_c22 bl[22] br[22] wl[61] vdd gnd cell_6t
Xbit_r62_c22 bl[22] br[22] wl[62] vdd gnd cell_6t
Xbit_r63_c22 bl[22] br[22] wl[63] vdd gnd cell_6t
Xbit_r64_c22 bl[22] br[22] wl[64] vdd gnd cell_6t
Xbit_r65_c22 bl[22] br[22] wl[65] vdd gnd cell_6t
Xbit_r66_c22 bl[22] br[22] wl[66] vdd gnd cell_6t
Xbit_r67_c22 bl[22] br[22] wl[67] vdd gnd cell_6t
Xbit_r68_c22 bl[22] br[22] wl[68] vdd gnd cell_6t
Xbit_r69_c22 bl[22] br[22] wl[69] vdd gnd cell_6t
Xbit_r70_c22 bl[22] br[22] wl[70] vdd gnd cell_6t
Xbit_r71_c22 bl[22] br[22] wl[71] vdd gnd cell_6t
Xbit_r72_c22 bl[22] br[22] wl[72] vdd gnd cell_6t
Xbit_r73_c22 bl[22] br[22] wl[73] vdd gnd cell_6t
Xbit_r74_c22 bl[22] br[22] wl[74] vdd gnd cell_6t
Xbit_r75_c22 bl[22] br[22] wl[75] vdd gnd cell_6t
Xbit_r76_c22 bl[22] br[22] wl[76] vdd gnd cell_6t
Xbit_r77_c22 bl[22] br[22] wl[77] vdd gnd cell_6t
Xbit_r78_c22 bl[22] br[22] wl[78] vdd gnd cell_6t
Xbit_r79_c22 bl[22] br[22] wl[79] vdd gnd cell_6t
Xbit_r80_c22 bl[22] br[22] wl[80] vdd gnd cell_6t
Xbit_r81_c22 bl[22] br[22] wl[81] vdd gnd cell_6t
Xbit_r82_c22 bl[22] br[22] wl[82] vdd gnd cell_6t
Xbit_r83_c22 bl[22] br[22] wl[83] vdd gnd cell_6t
Xbit_r84_c22 bl[22] br[22] wl[84] vdd gnd cell_6t
Xbit_r85_c22 bl[22] br[22] wl[85] vdd gnd cell_6t
Xbit_r86_c22 bl[22] br[22] wl[86] vdd gnd cell_6t
Xbit_r87_c22 bl[22] br[22] wl[87] vdd gnd cell_6t
Xbit_r88_c22 bl[22] br[22] wl[88] vdd gnd cell_6t
Xbit_r89_c22 bl[22] br[22] wl[89] vdd gnd cell_6t
Xbit_r90_c22 bl[22] br[22] wl[90] vdd gnd cell_6t
Xbit_r91_c22 bl[22] br[22] wl[91] vdd gnd cell_6t
Xbit_r92_c22 bl[22] br[22] wl[92] vdd gnd cell_6t
Xbit_r93_c22 bl[22] br[22] wl[93] vdd gnd cell_6t
Xbit_r94_c22 bl[22] br[22] wl[94] vdd gnd cell_6t
Xbit_r95_c22 bl[22] br[22] wl[95] vdd gnd cell_6t
Xbit_r96_c22 bl[22] br[22] wl[96] vdd gnd cell_6t
Xbit_r97_c22 bl[22] br[22] wl[97] vdd gnd cell_6t
Xbit_r98_c22 bl[22] br[22] wl[98] vdd gnd cell_6t
Xbit_r99_c22 bl[22] br[22] wl[99] vdd gnd cell_6t
Xbit_r100_c22 bl[22] br[22] wl[100] vdd gnd cell_6t
Xbit_r101_c22 bl[22] br[22] wl[101] vdd gnd cell_6t
Xbit_r102_c22 bl[22] br[22] wl[102] vdd gnd cell_6t
Xbit_r103_c22 bl[22] br[22] wl[103] vdd gnd cell_6t
Xbit_r104_c22 bl[22] br[22] wl[104] vdd gnd cell_6t
Xbit_r105_c22 bl[22] br[22] wl[105] vdd gnd cell_6t
Xbit_r106_c22 bl[22] br[22] wl[106] vdd gnd cell_6t
Xbit_r107_c22 bl[22] br[22] wl[107] vdd gnd cell_6t
Xbit_r108_c22 bl[22] br[22] wl[108] vdd gnd cell_6t
Xbit_r109_c22 bl[22] br[22] wl[109] vdd gnd cell_6t
Xbit_r110_c22 bl[22] br[22] wl[110] vdd gnd cell_6t
Xbit_r111_c22 bl[22] br[22] wl[111] vdd gnd cell_6t
Xbit_r112_c22 bl[22] br[22] wl[112] vdd gnd cell_6t
Xbit_r113_c22 bl[22] br[22] wl[113] vdd gnd cell_6t
Xbit_r114_c22 bl[22] br[22] wl[114] vdd gnd cell_6t
Xbit_r115_c22 bl[22] br[22] wl[115] vdd gnd cell_6t
Xbit_r116_c22 bl[22] br[22] wl[116] vdd gnd cell_6t
Xbit_r117_c22 bl[22] br[22] wl[117] vdd gnd cell_6t
Xbit_r118_c22 bl[22] br[22] wl[118] vdd gnd cell_6t
Xbit_r119_c22 bl[22] br[22] wl[119] vdd gnd cell_6t
Xbit_r120_c22 bl[22] br[22] wl[120] vdd gnd cell_6t
Xbit_r121_c22 bl[22] br[22] wl[121] vdd gnd cell_6t
Xbit_r122_c22 bl[22] br[22] wl[122] vdd gnd cell_6t
Xbit_r123_c22 bl[22] br[22] wl[123] vdd gnd cell_6t
Xbit_r124_c22 bl[22] br[22] wl[124] vdd gnd cell_6t
Xbit_r125_c22 bl[22] br[22] wl[125] vdd gnd cell_6t
Xbit_r126_c22 bl[22] br[22] wl[126] vdd gnd cell_6t
Xbit_r127_c22 bl[22] br[22] wl[127] vdd gnd cell_6t
Xbit_r0_c23 bl[23] br[23] wl[0] vdd gnd cell_6t
Xbit_r1_c23 bl[23] br[23] wl[1] vdd gnd cell_6t
Xbit_r2_c23 bl[23] br[23] wl[2] vdd gnd cell_6t
Xbit_r3_c23 bl[23] br[23] wl[3] vdd gnd cell_6t
Xbit_r4_c23 bl[23] br[23] wl[4] vdd gnd cell_6t
Xbit_r5_c23 bl[23] br[23] wl[5] vdd gnd cell_6t
Xbit_r6_c23 bl[23] br[23] wl[6] vdd gnd cell_6t
Xbit_r7_c23 bl[23] br[23] wl[7] vdd gnd cell_6t
Xbit_r8_c23 bl[23] br[23] wl[8] vdd gnd cell_6t
Xbit_r9_c23 bl[23] br[23] wl[9] vdd gnd cell_6t
Xbit_r10_c23 bl[23] br[23] wl[10] vdd gnd cell_6t
Xbit_r11_c23 bl[23] br[23] wl[11] vdd gnd cell_6t
Xbit_r12_c23 bl[23] br[23] wl[12] vdd gnd cell_6t
Xbit_r13_c23 bl[23] br[23] wl[13] vdd gnd cell_6t
Xbit_r14_c23 bl[23] br[23] wl[14] vdd gnd cell_6t
Xbit_r15_c23 bl[23] br[23] wl[15] vdd gnd cell_6t
Xbit_r16_c23 bl[23] br[23] wl[16] vdd gnd cell_6t
Xbit_r17_c23 bl[23] br[23] wl[17] vdd gnd cell_6t
Xbit_r18_c23 bl[23] br[23] wl[18] vdd gnd cell_6t
Xbit_r19_c23 bl[23] br[23] wl[19] vdd gnd cell_6t
Xbit_r20_c23 bl[23] br[23] wl[20] vdd gnd cell_6t
Xbit_r21_c23 bl[23] br[23] wl[21] vdd gnd cell_6t
Xbit_r22_c23 bl[23] br[23] wl[22] vdd gnd cell_6t
Xbit_r23_c23 bl[23] br[23] wl[23] vdd gnd cell_6t
Xbit_r24_c23 bl[23] br[23] wl[24] vdd gnd cell_6t
Xbit_r25_c23 bl[23] br[23] wl[25] vdd gnd cell_6t
Xbit_r26_c23 bl[23] br[23] wl[26] vdd gnd cell_6t
Xbit_r27_c23 bl[23] br[23] wl[27] vdd gnd cell_6t
Xbit_r28_c23 bl[23] br[23] wl[28] vdd gnd cell_6t
Xbit_r29_c23 bl[23] br[23] wl[29] vdd gnd cell_6t
Xbit_r30_c23 bl[23] br[23] wl[30] vdd gnd cell_6t
Xbit_r31_c23 bl[23] br[23] wl[31] vdd gnd cell_6t
Xbit_r32_c23 bl[23] br[23] wl[32] vdd gnd cell_6t
Xbit_r33_c23 bl[23] br[23] wl[33] vdd gnd cell_6t
Xbit_r34_c23 bl[23] br[23] wl[34] vdd gnd cell_6t
Xbit_r35_c23 bl[23] br[23] wl[35] vdd gnd cell_6t
Xbit_r36_c23 bl[23] br[23] wl[36] vdd gnd cell_6t
Xbit_r37_c23 bl[23] br[23] wl[37] vdd gnd cell_6t
Xbit_r38_c23 bl[23] br[23] wl[38] vdd gnd cell_6t
Xbit_r39_c23 bl[23] br[23] wl[39] vdd gnd cell_6t
Xbit_r40_c23 bl[23] br[23] wl[40] vdd gnd cell_6t
Xbit_r41_c23 bl[23] br[23] wl[41] vdd gnd cell_6t
Xbit_r42_c23 bl[23] br[23] wl[42] vdd gnd cell_6t
Xbit_r43_c23 bl[23] br[23] wl[43] vdd gnd cell_6t
Xbit_r44_c23 bl[23] br[23] wl[44] vdd gnd cell_6t
Xbit_r45_c23 bl[23] br[23] wl[45] vdd gnd cell_6t
Xbit_r46_c23 bl[23] br[23] wl[46] vdd gnd cell_6t
Xbit_r47_c23 bl[23] br[23] wl[47] vdd gnd cell_6t
Xbit_r48_c23 bl[23] br[23] wl[48] vdd gnd cell_6t
Xbit_r49_c23 bl[23] br[23] wl[49] vdd gnd cell_6t
Xbit_r50_c23 bl[23] br[23] wl[50] vdd gnd cell_6t
Xbit_r51_c23 bl[23] br[23] wl[51] vdd gnd cell_6t
Xbit_r52_c23 bl[23] br[23] wl[52] vdd gnd cell_6t
Xbit_r53_c23 bl[23] br[23] wl[53] vdd gnd cell_6t
Xbit_r54_c23 bl[23] br[23] wl[54] vdd gnd cell_6t
Xbit_r55_c23 bl[23] br[23] wl[55] vdd gnd cell_6t
Xbit_r56_c23 bl[23] br[23] wl[56] vdd gnd cell_6t
Xbit_r57_c23 bl[23] br[23] wl[57] vdd gnd cell_6t
Xbit_r58_c23 bl[23] br[23] wl[58] vdd gnd cell_6t
Xbit_r59_c23 bl[23] br[23] wl[59] vdd gnd cell_6t
Xbit_r60_c23 bl[23] br[23] wl[60] vdd gnd cell_6t
Xbit_r61_c23 bl[23] br[23] wl[61] vdd gnd cell_6t
Xbit_r62_c23 bl[23] br[23] wl[62] vdd gnd cell_6t
Xbit_r63_c23 bl[23] br[23] wl[63] vdd gnd cell_6t
Xbit_r64_c23 bl[23] br[23] wl[64] vdd gnd cell_6t
Xbit_r65_c23 bl[23] br[23] wl[65] vdd gnd cell_6t
Xbit_r66_c23 bl[23] br[23] wl[66] vdd gnd cell_6t
Xbit_r67_c23 bl[23] br[23] wl[67] vdd gnd cell_6t
Xbit_r68_c23 bl[23] br[23] wl[68] vdd gnd cell_6t
Xbit_r69_c23 bl[23] br[23] wl[69] vdd gnd cell_6t
Xbit_r70_c23 bl[23] br[23] wl[70] vdd gnd cell_6t
Xbit_r71_c23 bl[23] br[23] wl[71] vdd gnd cell_6t
Xbit_r72_c23 bl[23] br[23] wl[72] vdd gnd cell_6t
Xbit_r73_c23 bl[23] br[23] wl[73] vdd gnd cell_6t
Xbit_r74_c23 bl[23] br[23] wl[74] vdd gnd cell_6t
Xbit_r75_c23 bl[23] br[23] wl[75] vdd gnd cell_6t
Xbit_r76_c23 bl[23] br[23] wl[76] vdd gnd cell_6t
Xbit_r77_c23 bl[23] br[23] wl[77] vdd gnd cell_6t
Xbit_r78_c23 bl[23] br[23] wl[78] vdd gnd cell_6t
Xbit_r79_c23 bl[23] br[23] wl[79] vdd gnd cell_6t
Xbit_r80_c23 bl[23] br[23] wl[80] vdd gnd cell_6t
Xbit_r81_c23 bl[23] br[23] wl[81] vdd gnd cell_6t
Xbit_r82_c23 bl[23] br[23] wl[82] vdd gnd cell_6t
Xbit_r83_c23 bl[23] br[23] wl[83] vdd gnd cell_6t
Xbit_r84_c23 bl[23] br[23] wl[84] vdd gnd cell_6t
Xbit_r85_c23 bl[23] br[23] wl[85] vdd gnd cell_6t
Xbit_r86_c23 bl[23] br[23] wl[86] vdd gnd cell_6t
Xbit_r87_c23 bl[23] br[23] wl[87] vdd gnd cell_6t
Xbit_r88_c23 bl[23] br[23] wl[88] vdd gnd cell_6t
Xbit_r89_c23 bl[23] br[23] wl[89] vdd gnd cell_6t
Xbit_r90_c23 bl[23] br[23] wl[90] vdd gnd cell_6t
Xbit_r91_c23 bl[23] br[23] wl[91] vdd gnd cell_6t
Xbit_r92_c23 bl[23] br[23] wl[92] vdd gnd cell_6t
Xbit_r93_c23 bl[23] br[23] wl[93] vdd gnd cell_6t
Xbit_r94_c23 bl[23] br[23] wl[94] vdd gnd cell_6t
Xbit_r95_c23 bl[23] br[23] wl[95] vdd gnd cell_6t
Xbit_r96_c23 bl[23] br[23] wl[96] vdd gnd cell_6t
Xbit_r97_c23 bl[23] br[23] wl[97] vdd gnd cell_6t
Xbit_r98_c23 bl[23] br[23] wl[98] vdd gnd cell_6t
Xbit_r99_c23 bl[23] br[23] wl[99] vdd gnd cell_6t
Xbit_r100_c23 bl[23] br[23] wl[100] vdd gnd cell_6t
Xbit_r101_c23 bl[23] br[23] wl[101] vdd gnd cell_6t
Xbit_r102_c23 bl[23] br[23] wl[102] vdd gnd cell_6t
Xbit_r103_c23 bl[23] br[23] wl[103] vdd gnd cell_6t
Xbit_r104_c23 bl[23] br[23] wl[104] vdd gnd cell_6t
Xbit_r105_c23 bl[23] br[23] wl[105] vdd gnd cell_6t
Xbit_r106_c23 bl[23] br[23] wl[106] vdd gnd cell_6t
Xbit_r107_c23 bl[23] br[23] wl[107] vdd gnd cell_6t
Xbit_r108_c23 bl[23] br[23] wl[108] vdd gnd cell_6t
Xbit_r109_c23 bl[23] br[23] wl[109] vdd gnd cell_6t
Xbit_r110_c23 bl[23] br[23] wl[110] vdd gnd cell_6t
Xbit_r111_c23 bl[23] br[23] wl[111] vdd gnd cell_6t
Xbit_r112_c23 bl[23] br[23] wl[112] vdd gnd cell_6t
Xbit_r113_c23 bl[23] br[23] wl[113] vdd gnd cell_6t
Xbit_r114_c23 bl[23] br[23] wl[114] vdd gnd cell_6t
Xbit_r115_c23 bl[23] br[23] wl[115] vdd gnd cell_6t
Xbit_r116_c23 bl[23] br[23] wl[116] vdd gnd cell_6t
Xbit_r117_c23 bl[23] br[23] wl[117] vdd gnd cell_6t
Xbit_r118_c23 bl[23] br[23] wl[118] vdd gnd cell_6t
Xbit_r119_c23 bl[23] br[23] wl[119] vdd gnd cell_6t
Xbit_r120_c23 bl[23] br[23] wl[120] vdd gnd cell_6t
Xbit_r121_c23 bl[23] br[23] wl[121] vdd gnd cell_6t
Xbit_r122_c23 bl[23] br[23] wl[122] vdd gnd cell_6t
Xbit_r123_c23 bl[23] br[23] wl[123] vdd gnd cell_6t
Xbit_r124_c23 bl[23] br[23] wl[124] vdd gnd cell_6t
Xbit_r125_c23 bl[23] br[23] wl[125] vdd gnd cell_6t
Xbit_r126_c23 bl[23] br[23] wl[126] vdd gnd cell_6t
Xbit_r127_c23 bl[23] br[23] wl[127] vdd gnd cell_6t
Xbit_r0_c24 bl[24] br[24] wl[0] vdd gnd cell_6t
Xbit_r1_c24 bl[24] br[24] wl[1] vdd gnd cell_6t
Xbit_r2_c24 bl[24] br[24] wl[2] vdd gnd cell_6t
Xbit_r3_c24 bl[24] br[24] wl[3] vdd gnd cell_6t
Xbit_r4_c24 bl[24] br[24] wl[4] vdd gnd cell_6t
Xbit_r5_c24 bl[24] br[24] wl[5] vdd gnd cell_6t
Xbit_r6_c24 bl[24] br[24] wl[6] vdd gnd cell_6t
Xbit_r7_c24 bl[24] br[24] wl[7] vdd gnd cell_6t
Xbit_r8_c24 bl[24] br[24] wl[8] vdd gnd cell_6t
Xbit_r9_c24 bl[24] br[24] wl[9] vdd gnd cell_6t
Xbit_r10_c24 bl[24] br[24] wl[10] vdd gnd cell_6t
Xbit_r11_c24 bl[24] br[24] wl[11] vdd gnd cell_6t
Xbit_r12_c24 bl[24] br[24] wl[12] vdd gnd cell_6t
Xbit_r13_c24 bl[24] br[24] wl[13] vdd gnd cell_6t
Xbit_r14_c24 bl[24] br[24] wl[14] vdd gnd cell_6t
Xbit_r15_c24 bl[24] br[24] wl[15] vdd gnd cell_6t
Xbit_r16_c24 bl[24] br[24] wl[16] vdd gnd cell_6t
Xbit_r17_c24 bl[24] br[24] wl[17] vdd gnd cell_6t
Xbit_r18_c24 bl[24] br[24] wl[18] vdd gnd cell_6t
Xbit_r19_c24 bl[24] br[24] wl[19] vdd gnd cell_6t
Xbit_r20_c24 bl[24] br[24] wl[20] vdd gnd cell_6t
Xbit_r21_c24 bl[24] br[24] wl[21] vdd gnd cell_6t
Xbit_r22_c24 bl[24] br[24] wl[22] vdd gnd cell_6t
Xbit_r23_c24 bl[24] br[24] wl[23] vdd gnd cell_6t
Xbit_r24_c24 bl[24] br[24] wl[24] vdd gnd cell_6t
Xbit_r25_c24 bl[24] br[24] wl[25] vdd gnd cell_6t
Xbit_r26_c24 bl[24] br[24] wl[26] vdd gnd cell_6t
Xbit_r27_c24 bl[24] br[24] wl[27] vdd gnd cell_6t
Xbit_r28_c24 bl[24] br[24] wl[28] vdd gnd cell_6t
Xbit_r29_c24 bl[24] br[24] wl[29] vdd gnd cell_6t
Xbit_r30_c24 bl[24] br[24] wl[30] vdd gnd cell_6t
Xbit_r31_c24 bl[24] br[24] wl[31] vdd gnd cell_6t
Xbit_r32_c24 bl[24] br[24] wl[32] vdd gnd cell_6t
Xbit_r33_c24 bl[24] br[24] wl[33] vdd gnd cell_6t
Xbit_r34_c24 bl[24] br[24] wl[34] vdd gnd cell_6t
Xbit_r35_c24 bl[24] br[24] wl[35] vdd gnd cell_6t
Xbit_r36_c24 bl[24] br[24] wl[36] vdd gnd cell_6t
Xbit_r37_c24 bl[24] br[24] wl[37] vdd gnd cell_6t
Xbit_r38_c24 bl[24] br[24] wl[38] vdd gnd cell_6t
Xbit_r39_c24 bl[24] br[24] wl[39] vdd gnd cell_6t
Xbit_r40_c24 bl[24] br[24] wl[40] vdd gnd cell_6t
Xbit_r41_c24 bl[24] br[24] wl[41] vdd gnd cell_6t
Xbit_r42_c24 bl[24] br[24] wl[42] vdd gnd cell_6t
Xbit_r43_c24 bl[24] br[24] wl[43] vdd gnd cell_6t
Xbit_r44_c24 bl[24] br[24] wl[44] vdd gnd cell_6t
Xbit_r45_c24 bl[24] br[24] wl[45] vdd gnd cell_6t
Xbit_r46_c24 bl[24] br[24] wl[46] vdd gnd cell_6t
Xbit_r47_c24 bl[24] br[24] wl[47] vdd gnd cell_6t
Xbit_r48_c24 bl[24] br[24] wl[48] vdd gnd cell_6t
Xbit_r49_c24 bl[24] br[24] wl[49] vdd gnd cell_6t
Xbit_r50_c24 bl[24] br[24] wl[50] vdd gnd cell_6t
Xbit_r51_c24 bl[24] br[24] wl[51] vdd gnd cell_6t
Xbit_r52_c24 bl[24] br[24] wl[52] vdd gnd cell_6t
Xbit_r53_c24 bl[24] br[24] wl[53] vdd gnd cell_6t
Xbit_r54_c24 bl[24] br[24] wl[54] vdd gnd cell_6t
Xbit_r55_c24 bl[24] br[24] wl[55] vdd gnd cell_6t
Xbit_r56_c24 bl[24] br[24] wl[56] vdd gnd cell_6t
Xbit_r57_c24 bl[24] br[24] wl[57] vdd gnd cell_6t
Xbit_r58_c24 bl[24] br[24] wl[58] vdd gnd cell_6t
Xbit_r59_c24 bl[24] br[24] wl[59] vdd gnd cell_6t
Xbit_r60_c24 bl[24] br[24] wl[60] vdd gnd cell_6t
Xbit_r61_c24 bl[24] br[24] wl[61] vdd gnd cell_6t
Xbit_r62_c24 bl[24] br[24] wl[62] vdd gnd cell_6t
Xbit_r63_c24 bl[24] br[24] wl[63] vdd gnd cell_6t
Xbit_r64_c24 bl[24] br[24] wl[64] vdd gnd cell_6t
Xbit_r65_c24 bl[24] br[24] wl[65] vdd gnd cell_6t
Xbit_r66_c24 bl[24] br[24] wl[66] vdd gnd cell_6t
Xbit_r67_c24 bl[24] br[24] wl[67] vdd gnd cell_6t
Xbit_r68_c24 bl[24] br[24] wl[68] vdd gnd cell_6t
Xbit_r69_c24 bl[24] br[24] wl[69] vdd gnd cell_6t
Xbit_r70_c24 bl[24] br[24] wl[70] vdd gnd cell_6t
Xbit_r71_c24 bl[24] br[24] wl[71] vdd gnd cell_6t
Xbit_r72_c24 bl[24] br[24] wl[72] vdd gnd cell_6t
Xbit_r73_c24 bl[24] br[24] wl[73] vdd gnd cell_6t
Xbit_r74_c24 bl[24] br[24] wl[74] vdd gnd cell_6t
Xbit_r75_c24 bl[24] br[24] wl[75] vdd gnd cell_6t
Xbit_r76_c24 bl[24] br[24] wl[76] vdd gnd cell_6t
Xbit_r77_c24 bl[24] br[24] wl[77] vdd gnd cell_6t
Xbit_r78_c24 bl[24] br[24] wl[78] vdd gnd cell_6t
Xbit_r79_c24 bl[24] br[24] wl[79] vdd gnd cell_6t
Xbit_r80_c24 bl[24] br[24] wl[80] vdd gnd cell_6t
Xbit_r81_c24 bl[24] br[24] wl[81] vdd gnd cell_6t
Xbit_r82_c24 bl[24] br[24] wl[82] vdd gnd cell_6t
Xbit_r83_c24 bl[24] br[24] wl[83] vdd gnd cell_6t
Xbit_r84_c24 bl[24] br[24] wl[84] vdd gnd cell_6t
Xbit_r85_c24 bl[24] br[24] wl[85] vdd gnd cell_6t
Xbit_r86_c24 bl[24] br[24] wl[86] vdd gnd cell_6t
Xbit_r87_c24 bl[24] br[24] wl[87] vdd gnd cell_6t
Xbit_r88_c24 bl[24] br[24] wl[88] vdd gnd cell_6t
Xbit_r89_c24 bl[24] br[24] wl[89] vdd gnd cell_6t
Xbit_r90_c24 bl[24] br[24] wl[90] vdd gnd cell_6t
Xbit_r91_c24 bl[24] br[24] wl[91] vdd gnd cell_6t
Xbit_r92_c24 bl[24] br[24] wl[92] vdd gnd cell_6t
Xbit_r93_c24 bl[24] br[24] wl[93] vdd gnd cell_6t
Xbit_r94_c24 bl[24] br[24] wl[94] vdd gnd cell_6t
Xbit_r95_c24 bl[24] br[24] wl[95] vdd gnd cell_6t
Xbit_r96_c24 bl[24] br[24] wl[96] vdd gnd cell_6t
Xbit_r97_c24 bl[24] br[24] wl[97] vdd gnd cell_6t
Xbit_r98_c24 bl[24] br[24] wl[98] vdd gnd cell_6t
Xbit_r99_c24 bl[24] br[24] wl[99] vdd gnd cell_6t
Xbit_r100_c24 bl[24] br[24] wl[100] vdd gnd cell_6t
Xbit_r101_c24 bl[24] br[24] wl[101] vdd gnd cell_6t
Xbit_r102_c24 bl[24] br[24] wl[102] vdd gnd cell_6t
Xbit_r103_c24 bl[24] br[24] wl[103] vdd gnd cell_6t
Xbit_r104_c24 bl[24] br[24] wl[104] vdd gnd cell_6t
Xbit_r105_c24 bl[24] br[24] wl[105] vdd gnd cell_6t
Xbit_r106_c24 bl[24] br[24] wl[106] vdd gnd cell_6t
Xbit_r107_c24 bl[24] br[24] wl[107] vdd gnd cell_6t
Xbit_r108_c24 bl[24] br[24] wl[108] vdd gnd cell_6t
Xbit_r109_c24 bl[24] br[24] wl[109] vdd gnd cell_6t
Xbit_r110_c24 bl[24] br[24] wl[110] vdd gnd cell_6t
Xbit_r111_c24 bl[24] br[24] wl[111] vdd gnd cell_6t
Xbit_r112_c24 bl[24] br[24] wl[112] vdd gnd cell_6t
Xbit_r113_c24 bl[24] br[24] wl[113] vdd gnd cell_6t
Xbit_r114_c24 bl[24] br[24] wl[114] vdd gnd cell_6t
Xbit_r115_c24 bl[24] br[24] wl[115] vdd gnd cell_6t
Xbit_r116_c24 bl[24] br[24] wl[116] vdd gnd cell_6t
Xbit_r117_c24 bl[24] br[24] wl[117] vdd gnd cell_6t
Xbit_r118_c24 bl[24] br[24] wl[118] vdd gnd cell_6t
Xbit_r119_c24 bl[24] br[24] wl[119] vdd gnd cell_6t
Xbit_r120_c24 bl[24] br[24] wl[120] vdd gnd cell_6t
Xbit_r121_c24 bl[24] br[24] wl[121] vdd gnd cell_6t
Xbit_r122_c24 bl[24] br[24] wl[122] vdd gnd cell_6t
Xbit_r123_c24 bl[24] br[24] wl[123] vdd gnd cell_6t
Xbit_r124_c24 bl[24] br[24] wl[124] vdd gnd cell_6t
Xbit_r125_c24 bl[24] br[24] wl[125] vdd gnd cell_6t
Xbit_r126_c24 bl[24] br[24] wl[126] vdd gnd cell_6t
Xbit_r127_c24 bl[24] br[24] wl[127] vdd gnd cell_6t
Xbit_r0_c25 bl[25] br[25] wl[0] vdd gnd cell_6t
Xbit_r1_c25 bl[25] br[25] wl[1] vdd gnd cell_6t
Xbit_r2_c25 bl[25] br[25] wl[2] vdd gnd cell_6t
Xbit_r3_c25 bl[25] br[25] wl[3] vdd gnd cell_6t
Xbit_r4_c25 bl[25] br[25] wl[4] vdd gnd cell_6t
Xbit_r5_c25 bl[25] br[25] wl[5] vdd gnd cell_6t
Xbit_r6_c25 bl[25] br[25] wl[6] vdd gnd cell_6t
Xbit_r7_c25 bl[25] br[25] wl[7] vdd gnd cell_6t
Xbit_r8_c25 bl[25] br[25] wl[8] vdd gnd cell_6t
Xbit_r9_c25 bl[25] br[25] wl[9] vdd gnd cell_6t
Xbit_r10_c25 bl[25] br[25] wl[10] vdd gnd cell_6t
Xbit_r11_c25 bl[25] br[25] wl[11] vdd gnd cell_6t
Xbit_r12_c25 bl[25] br[25] wl[12] vdd gnd cell_6t
Xbit_r13_c25 bl[25] br[25] wl[13] vdd gnd cell_6t
Xbit_r14_c25 bl[25] br[25] wl[14] vdd gnd cell_6t
Xbit_r15_c25 bl[25] br[25] wl[15] vdd gnd cell_6t
Xbit_r16_c25 bl[25] br[25] wl[16] vdd gnd cell_6t
Xbit_r17_c25 bl[25] br[25] wl[17] vdd gnd cell_6t
Xbit_r18_c25 bl[25] br[25] wl[18] vdd gnd cell_6t
Xbit_r19_c25 bl[25] br[25] wl[19] vdd gnd cell_6t
Xbit_r20_c25 bl[25] br[25] wl[20] vdd gnd cell_6t
Xbit_r21_c25 bl[25] br[25] wl[21] vdd gnd cell_6t
Xbit_r22_c25 bl[25] br[25] wl[22] vdd gnd cell_6t
Xbit_r23_c25 bl[25] br[25] wl[23] vdd gnd cell_6t
Xbit_r24_c25 bl[25] br[25] wl[24] vdd gnd cell_6t
Xbit_r25_c25 bl[25] br[25] wl[25] vdd gnd cell_6t
Xbit_r26_c25 bl[25] br[25] wl[26] vdd gnd cell_6t
Xbit_r27_c25 bl[25] br[25] wl[27] vdd gnd cell_6t
Xbit_r28_c25 bl[25] br[25] wl[28] vdd gnd cell_6t
Xbit_r29_c25 bl[25] br[25] wl[29] vdd gnd cell_6t
Xbit_r30_c25 bl[25] br[25] wl[30] vdd gnd cell_6t
Xbit_r31_c25 bl[25] br[25] wl[31] vdd gnd cell_6t
Xbit_r32_c25 bl[25] br[25] wl[32] vdd gnd cell_6t
Xbit_r33_c25 bl[25] br[25] wl[33] vdd gnd cell_6t
Xbit_r34_c25 bl[25] br[25] wl[34] vdd gnd cell_6t
Xbit_r35_c25 bl[25] br[25] wl[35] vdd gnd cell_6t
Xbit_r36_c25 bl[25] br[25] wl[36] vdd gnd cell_6t
Xbit_r37_c25 bl[25] br[25] wl[37] vdd gnd cell_6t
Xbit_r38_c25 bl[25] br[25] wl[38] vdd gnd cell_6t
Xbit_r39_c25 bl[25] br[25] wl[39] vdd gnd cell_6t
Xbit_r40_c25 bl[25] br[25] wl[40] vdd gnd cell_6t
Xbit_r41_c25 bl[25] br[25] wl[41] vdd gnd cell_6t
Xbit_r42_c25 bl[25] br[25] wl[42] vdd gnd cell_6t
Xbit_r43_c25 bl[25] br[25] wl[43] vdd gnd cell_6t
Xbit_r44_c25 bl[25] br[25] wl[44] vdd gnd cell_6t
Xbit_r45_c25 bl[25] br[25] wl[45] vdd gnd cell_6t
Xbit_r46_c25 bl[25] br[25] wl[46] vdd gnd cell_6t
Xbit_r47_c25 bl[25] br[25] wl[47] vdd gnd cell_6t
Xbit_r48_c25 bl[25] br[25] wl[48] vdd gnd cell_6t
Xbit_r49_c25 bl[25] br[25] wl[49] vdd gnd cell_6t
Xbit_r50_c25 bl[25] br[25] wl[50] vdd gnd cell_6t
Xbit_r51_c25 bl[25] br[25] wl[51] vdd gnd cell_6t
Xbit_r52_c25 bl[25] br[25] wl[52] vdd gnd cell_6t
Xbit_r53_c25 bl[25] br[25] wl[53] vdd gnd cell_6t
Xbit_r54_c25 bl[25] br[25] wl[54] vdd gnd cell_6t
Xbit_r55_c25 bl[25] br[25] wl[55] vdd gnd cell_6t
Xbit_r56_c25 bl[25] br[25] wl[56] vdd gnd cell_6t
Xbit_r57_c25 bl[25] br[25] wl[57] vdd gnd cell_6t
Xbit_r58_c25 bl[25] br[25] wl[58] vdd gnd cell_6t
Xbit_r59_c25 bl[25] br[25] wl[59] vdd gnd cell_6t
Xbit_r60_c25 bl[25] br[25] wl[60] vdd gnd cell_6t
Xbit_r61_c25 bl[25] br[25] wl[61] vdd gnd cell_6t
Xbit_r62_c25 bl[25] br[25] wl[62] vdd gnd cell_6t
Xbit_r63_c25 bl[25] br[25] wl[63] vdd gnd cell_6t
Xbit_r64_c25 bl[25] br[25] wl[64] vdd gnd cell_6t
Xbit_r65_c25 bl[25] br[25] wl[65] vdd gnd cell_6t
Xbit_r66_c25 bl[25] br[25] wl[66] vdd gnd cell_6t
Xbit_r67_c25 bl[25] br[25] wl[67] vdd gnd cell_6t
Xbit_r68_c25 bl[25] br[25] wl[68] vdd gnd cell_6t
Xbit_r69_c25 bl[25] br[25] wl[69] vdd gnd cell_6t
Xbit_r70_c25 bl[25] br[25] wl[70] vdd gnd cell_6t
Xbit_r71_c25 bl[25] br[25] wl[71] vdd gnd cell_6t
Xbit_r72_c25 bl[25] br[25] wl[72] vdd gnd cell_6t
Xbit_r73_c25 bl[25] br[25] wl[73] vdd gnd cell_6t
Xbit_r74_c25 bl[25] br[25] wl[74] vdd gnd cell_6t
Xbit_r75_c25 bl[25] br[25] wl[75] vdd gnd cell_6t
Xbit_r76_c25 bl[25] br[25] wl[76] vdd gnd cell_6t
Xbit_r77_c25 bl[25] br[25] wl[77] vdd gnd cell_6t
Xbit_r78_c25 bl[25] br[25] wl[78] vdd gnd cell_6t
Xbit_r79_c25 bl[25] br[25] wl[79] vdd gnd cell_6t
Xbit_r80_c25 bl[25] br[25] wl[80] vdd gnd cell_6t
Xbit_r81_c25 bl[25] br[25] wl[81] vdd gnd cell_6t
Xbit_r82_c25 bl[25] br[25] wl[82] vdd gnd cell_6t
Xbit_r83_c25 bl[25] br[25] wl[83] vdd gnd cell_6t
Xbit_r84_c25 bl[25] br[25] wl[84] vdd gnd cell_6t
Xbit_r85_c25 bl[25] br[25] wl[85] vdd gnd cell_6t
Xbit_r86_c25 bl[25] br[25] wl[86] vdd gnd cell_6t
Xbit_r87_c25 bl[25] br[25] wl[87] vdd gnd cell_6t
Xbit_r88_c25 bl[25] br[25] wl[88] vdd gnd cell_6t
Xbit_r89_c25 bl[25] br[25] wl[89] vdd gnd cell_6t
Xbit_r90_c25 bl[25] br[25] wl[90] vdd gnd cell_6t
Xbit_r91_c25 bl[25] br[25] wl[91] vdd gnd cell_6t
Xbit_r92_c25 bl[25] br[25] wl[92] vdd gnd cell_6t
Xbit_r93_c25 bl[25] br[25] wl[93] vdd gnd cell_6t
Xbit_r94_c25 bl[25] br[25] wl[94] vdd gnd cell_6t
Xbit_r95_c25 bl[25] br[25] wl[95] vdd gnd cell_6t
Xbit_r96_c25 bl[25] br[25] wl[96] vdd gnd cell_6t
Xbit_r97_c25 bl[25] br[25] wl[97] vdd gnd cell_6t
Xbit_r98_c25 bl[25] br[25] wl[98] vdd gnd cell_6t
Xbit_r99_c25 bl[25] br[25] wl[99] vdd gnd cell_6t
Xbit_r100_c25 bl[25] br[25] wl[100] vdd gnd cell_6t
Xbit_r101_c25 bl[25] br[25] wl[101] vdd gnd cell_6t
Xbit_r102_c25 bl[25] br[25] wl[102] vdd gnd cell_6t
Xbit_r103_c25 bl[25] br[25] wl[103] vdd gnd cell_6t
Xbit_r104_c25 bl[25] br[25] wl[104] vdd gnd cell_6t
Xbit_r105_c25 bl[25] br[25] wl[105] vdd gnd cell_6t
Xbit_r106_c25 bl[25] br[25] wl[106] vdd gnd cell_6t
Xbit_r107_c25 bl[25] br[25] wl[107] vdd gnd cell_6t
Xbit_r108_c25 bl[25] br[25] wl[108] vdd gnd cell_6t
Xbit_r109_c25 bl[25] br[25] wl[109] vdd gnd cell_6t
Xbit_r110_c25 bl[25] br[25] wl[110] vdd gnd cell_6t
Xbit_r111_c25 bl[25] br[25] wl[111] vdd gnd cell_6t
Xbit_r112_c25 bl[25] br[25] wl[112] vdd gnd cell_6t
Xbit_r113_c25 bl[25] br[25] wl[113] vdd gnd cell_6t
Xbit_r114_c25 bl[25] br[25] wl[114] vdd gnd cell_6t
Xbit_r115_c25 bl[25] br[25] wl[115] vdd gnd cell_6t
Xbit_r116_c25 bl[25] br[25] wl[116] vdd gnd cell_6t
Xbit_r117_c25 bl[25] br[25] wl[117] vdd gnd cell_6t
Xbit_r118_c25 bl[25] br[25] wl[118] vdd gnd cell_6t
Xbit_r119_c25 bl[25] br[25] wl[119] vdd gnd cell_6t
Xbit_r120_c25 bl[25] br[25] wl[120] vdd gnd cell_6t
Xbit_r121_c25 bl[25] br[25] wl[121] vdd gnd cell_6t
Xbit_r122_c25 bl[25] br[25] wl[122] vdd gnd cell_6t
Xbit_r123_c25 bl[25] br[25] wl[123] vdd gnd cell_6t
Xbit_r124_c25 bl[25] br[25] wl[124] vdd gnd cell_6t
Xbit_r125_c25 bl[25] br[25] wl[125] vdd gnd cell_6t
Xbit_r126_c25 bl[25] br[25] wl[126] vdd gnd cell_6t
Xbit_r127_c25 bl[25] br[25] wl[127] vdd gnd cell_6t
Xbit_r0_c26 bl[26] br[26] wl[0] vdd gnd cell_6t
Xbit_r1_c26 bl[26] br[26] wl[1] vdd gnd cell_6t
Xbit_r2_c26 bl[26] br[26] wl[2] vdd gnd cell_6t
Xbit_r3_c26 bl[26] br[26] wl[3] vdd gnd cell_6t
Xbit_r4_c26 bl[26] br[26] wl[4] vdd gnd cell_6t
Xbit_r5_c26 bl[26] br[26] wl[5] vdd gnd cell_6t
Xbit_r6_c26 bl[26] br[26] wl[6] vdd gnd cell_6t
Xbit_r7_c26 bl[26] br[26] wl[7] vdd gnd cell_6t
Xbit_r8_c26 bl[26] br[26] wl[8] vdd gnd cell_6t
Xbit_r9_c26 bl[26] br[26] wl[9] vdd gnd cell_6t
Xbit_r10_c26 bl[26] br[26] wl[10] vdd gnd cell_6t
Xbit_r11_c26 bl[26] br[26] wl[11] vdd gnd cell_6t
Xbit_r12_c26 bl[26] br[26] wl[12] vdd gnd cell_6t
Xbit_r13_c26 bl[26] br[26] wl[13] vdd gnd cell_6t
Xbit_r14_c26 bl[26] br[26] wl[14] vdd gnd cell_6t
Xbit_r15_c26 bl[26] br[26] wl[15] vdd gnd cell_6t
Xbit_r16_c26 bl[26] br[26] wl[16] vdd gnd cell_6t
Xbit_r17_c26 bl[26] br[26] wl[17] vdd gnd cell_6t
Xbit_r18_c26 bl[26] br[26] wl[18] vdd gnd cell_6t
Xbit_r19_c26 bl[26] br[26] wl[19] vdd gnd cell_6t
Xbit_r20_c26 bl[26] br[26] wl[20] vdd gnd cell_6t
Xbit_r21_c26 bl[26] br[26] wl[21] vdd gnd cell_6t
Xbit_r22_c26 bl[26] br[26] wl[22] vdd gnd cell_6t
Xbit_r23_c26 bl[26] br[26] wl[23] vdd gnd cell_6t
Xbit_r24_c26 bl[26] br[26] wl[24] vdd gnd cell_6t
Xbit_r25_c26 bl[26] br[26] wl[25] vdd gnd cell_6t
Xbit_r26_c26 bl[26] br[26] wl[26] vdd gnd cell_6t
Xbit_r27_c26 bl[26] br[26] wl[27] vdd gnd cell_6t
Xbit_r28_c26 bl[26] br[26] wl[28] vdd gnd cell_6t
Xbit_r29_c26 bl[26] br[26] wl[29] vdd gnd cell_6t
Xbit_r30_c26 bl[26] br[26] wl[30] vdd gnd cell_6t
Xbit_r31_c26 bl[26] br[26] wl[31] vdd gnd cell_6t
Xbit_r32_c26 bl[26] br[26] wl[32] vdd gnd cell_6t
Xbit_r33_c26 bl[26] br[26] wl[33] vdd gnd cell_6t
Xbit_r34_c26 bl[26] br[26] wl[34] vdd gnd cell_6t
Xbit_r35_c26 bl[26] br[26] wl[35] vdd gnd cell_6t
Xbit_r36_c26 bl[26] br[26] wl[36] vdd gnd cell_6t
Xbit_r37_c26 bl[26] br[26] wl[37] vdd gnd cell_6t
Xbit_r38_c26 bl[26] br[26] wl[38] vdd gnd cell_6t
Xbit_r39_c26 bl[26] br[26] wl[39] vdd gnd cell_6t
Xbit_r40_c26 bl[26] br[26] wl[40] vdd gnd cell_6t
Xbit_r41_c26 bl[26] br[26] wl[41] vdd gnd cell_6t
Xbit_r42_c26 bl[26] br[26] wl[42] vdd gnd cell_6t
Xbit_r43_c26 bl[26] br[26] wl[43] vdd gnd cell_6t
Xbit_r44_c26 bl[26] br[26] wl[44] vdd gnd cell_6t
Xbit_r45_c26 bl[26] br[26] wl[45] vdd gnd cell_6t
Xbit_r46_c26 bl[26] br[26] wl[46] vdd gnd cell_6t
Xbit_r47_c26 bl[26] br[26] wl[47] vdd gnd cell_6t
Xbit_r48_c26 bl[26] br[26] wl[48] vdd gnd cell_6t
Xbit_r49_c26 bl[26] br[26] wl[49] vdd gnd cell_6t
Xbit_r50_c26 bl[26] br[26] wl[50] vdd gnd cell_6t
Xbit_r51_c26 bl[26] br[26] wl[51] vdd gnd cell_6t
Xbit_r52_c26 bl[26] br[26] wl[52] vdd gnd cell_6t
Xbit_r53_c26 bl[26] br[26] wl[53] vdd gnd cell_6t
Xbit_r54_c26 bl[26] br[26] wl[54] vdd gnd cell_6t
Xbit_r55_c26 bl[26] br[26] wl[55] vdd gnd cell_6t
Xbit_r56_c26 bl[26] br[26] wl[56] vdd gnd cell_6t
Xbit_r57_c26 bl[26] br[26] wl[57] vdd gnd cell_6t
Xbit_r58_c26 bl[26] br[26] wl[58] vdd gnd cell_6t
Xbit_r59_c26 bl[26] br[26] wl[59] vdd gnd cell_6t
Xbit_r60_c26 bl[26] br[26] wl[60] vdd gnd cell_6t
Xbit_r61_c26 bl[26] br[26] wl[61] vdd gnd cell_6t
Xbit_r62_c26 bl[26] br[26] wl[62] vdd gnd cell_6t
Xbit_r63_c26 bl[26] br[26] wl[63] vdd gnd cell_6t
Xbit_r64_c26 bl[26] br[26] wl[64] vdd gnd cell_6t
Xbit_r65_c26 bl[26] br[26] wl[65] vdd gnd cell_6t
Xbit_r66_c26 bl[26] br[26] wl[66] vdd gnd cell_6t
Xbit_r67_c26 bl[26] br[26] wl[67] vdd gnd cell_6t
Xbit_r68_c26 bl[26] br[26] wl[68] vdd gnd cell_6t
Xbit_r69_c26 bl[26] br[26] wl[69] vdd gnd cell_6t
Xbit_r70_c26 bl[26] br[26] wl[70] vdd gnd cell_6t
Xbit_r71_c26 bl[26] br[26] wl[71] vdd gnd cell_6t
Xbit_r72_c26 bl[26] br[26] wl[72] vdd gnd cell_6t
Xbit_r73_c26 bl[26] br[26] wl[73] vdd gnd cell_6t
Xbit_r74_c26 bl[26] br[26] wl[74] vdd gnd cell_6t
Xbit_r75_c26 bl[26] br[26] wl[75] vdd gnd cell_6t
Xbit_r76_c26 bl[26] br[26] wl[76] vdd gnd cell_6t
Xbit_r77_c26 bl[26] br[26] wl[77] vdd gnd cell_6t
Xbit_r78_c26 bl[26] br[26] wl[78] vdd gnd cell_6t
Xbit_r79_c26 bl[26] br[26] wl[79] vdd gnd cell_6t
Xbit_r80_c26 bl[26] br[26] wl[80] vdd gnd cell_6t
Xbit_r81_c26 bl[26] br[26] wl[81] vdd gnd cell_6t
Xbit_r82_c26 bl[26] br[26] wl[82] vdd gnd cell_6t
Xbit_r83_c26 bl[26] br[26] wl[83] vdd gnd cell_6t
Xbit_r84_c26 bl[26] br[26] wl[84] vdd gnd cell_6t
Xbit_r85_c26 bl[26] br[26] wl[85] vdd gnd cell_6t
Xbit_r86_c26 bl[26] br[26] wl[86] vdd gnd cell_6t
Xbit_r87_c26 bl[26] br[26] wl[87] vdd gnd cell_6t
Xbit_r88_c26 bl[26] br[26] wl[88] vdd gnd cell_6t
Xbit_r89_c26 bl[26] br[26] wl[89] vdd gnd cell_6t
Xbit_r90_c26 bl[26] br[26] wl[90] vdd gnd cell_6t
Xbit_r91_c26 bl[26] br[26] wl[91] vdd gnd cell_6t
Xbit_r92_c26 bl[26] br[26] wl[92] vdd gnd cell_6t
Xbit_r93_c26 bl[26] br[26] wl[93] vdd gnd cell_6t
Xbit_r94_c26 bl[26] br[26] wl[94] vdd gnd cell_6t
Xbit_r95_c26 bl[26] br[26] wl[95] vdd gnd cell_6t
Xbit_r96_c26 bl[26] br[26] wl[96] vdd gnd cell_6t
Xbit_r97_c26 bl[26] br[26] wl[97] vdd gnd cell_6t
Xbit_r98_c26 bl[26] br[26] wl[98] vdd gnd cell_6t
Xbit_r99_c26 bl[26] br[26] wl[99] vdd gnd cell_6t
Xbit_r100_c26 bl[26] br[26] wl[100] vdd gnd cell_6t
Xbit_r101_c26 bl[26] br[26] wl[101] vdd gnd cell_6t
Xbit_r102_c26 bl[26] br[26] wl[102] vdd gnd cell_6t
Xbit_r103_c26 bl[26] br[26] wl[103] vdd gnd cell_6t
Xbit_r104_c26 bl[26] br[26] wl[104] vdd gnd cell_6t
Xbit_r105_c26 bl[26] br[26] wl[105] vdd gnd cell_6t
Xbit_r106_c26 bl[26] br[26] wl[106] vdd gnd cell_6t
Xbit_r107_c26 bl[26] br[26] wl[107] vdd gnd cell_6t
Xbit_r108_c26 bl[26] br[26] wl[108] vdd gnd cell_6t
Xbit_r109_c26 bl[26] br[26] wl[109] vdd gnd cell_6t
Xbit_r110_c26 bl[26] br[26] wl[110] vdd gnd cell_6t
Xbit_r111_c26 bl[26] br[26] wl[111] vdd gnd cell_6t
Xbit_r112_c26 bl[26] br[26] wl[112] vdd gnd cell_6t
Xbit_r113_c26 bl[26] br[26] wl[113] vdd gnd cell_6t
Xbit_r114_c26 bl[26] br[26] wl[114] vdd gnd cell_6t
Xbit_r115_c26 bl[26] br[26] wl[115] vdd gnd cell_6t
Xbit_r116_c26 bl[26] br[26] wl[116] vdd gnd cell_6t
Xbit_r117_c26 bl[26] br[26] wl[117] vdd gnd cell_6t
Xbit_r118_c26 bl[26] br[26] wl[118] vdd gnd cell_6t
Xbit_r119_c26 bl[26] br[26] wl[119] vdd gnd cell_6t
Xbit_r120_c26 bl[26] br[26] wl[120] vdd gnd cell_6t
Xbit_r121_c26 bl[26] br[26] wl[121] vdd gnd cell_6t
Xbit_r122_c26 bl[26] br[26] wl[122] vdd gnd cell_6t
Xbit_r123_c26 bl[26] br[26] wl[123] vdd gnd cell_6t
Xbit_r124_c26 bl[26] br[26] wl[124] vdd gnd cell_6t
Xbit_r125_c26 bl[26] br[26] wl[125] vdd gnd cell_6t
Xbit_r126_c26 bl[26] br[26] wl[126] vdd gnd cell_6t
Xbit_r127_c26 bl[26] br[26] wl[127] vdd gnd cell_6t
Xbit_r0_c27 bl[27] br[27] wl[0] vdd gnd cell_6t
Xbit_r1_c27 bl[27] br[27] wl[1] vdd gnd cell_6t
Xbit_r2_c27 bl[27] br[27] wl[2] vdd gnd cell_6t
Xbit_r3_c27 bl[27] br[27] wl[3] vdd gnd cell_6t
Xbit_r4_c27 bl[27] br[27] wl[4] vdd gnd cell_6t
Xbit_r5_c27 bl[27] br[27] wl[5] vdd gnd cell_6t
Xbit_r6_c27 bl[27] br[27] wl[6] vdd gnd cell_6t
Xbit_r7_c27 bl[27] br[27] wl[7] vdd gnd cell_6t
Xbit_r8_c27 bl[27] br[27] wl[8] vdd gnd cell_6t
Xbit_r9_c27 bl[27] br[27] wl[9] vdd gnd cell_6t
Xbit_r10_c27 bl[27] br[27] wl[10] vdd gnd cell_6t
Xbit_r11_c27 bl[27] br[27] wl[11] vdd gnd cell_6t
Xbit_r12_c27 bl[27] br[27] wl[12] vdd gnd cell_6t
Xbit_r13_c27 bl[27] br[27] wl[13] vdd gnd cell_6t
Xbit_r14_c27 bl[27] br[27] wl[14] vdd gnd cell_6t
Xbit_r15_c27 bl[27] br[27] wl[15] vdd gnd cell_6t
Xbit_r16_c27 bl[27] br[27] wl[16] vdd gnd cell_6t
Xbit_r17_c27 bl[27] br[27] wl[17] vdd gnd cell_6t
Xbit_r18_c27 bl[27] br[27] wl[18] vdd gnd cell_6t
Xbit_r19_c27 bl[27] br[27] wl[19] vdd gnd cell_6t
Xbit_r20_c27 bl[27] br[27] wl[20] vdd gnd cell_6t
Xbit_r21_c27 bl[27] br[27] wl[21] vdd gnd cell_6t
Xbit_r22_c27 bl[27] br[27] wl[22] vdd gnd cell_6t
Xbit_r23_c27 bl[27] br[27] wl[23] vdd gnd cell_6t
Xbit_r24_c27 bl[27] br[27] wl[24] vdd gnd cell_6t
Xbit_r25_c27 bl[27] br[27] wl[25] vdd gnd cell_6t
Xbit_r26_c27 bl[27] br[27] wl[26] vdd gnd cell_6t
Xbit_r27_c27 bl[27] br[27] wl[27] vdd gnd cell_6t
Xbit_r28_c27 bl[27] br[27] wl[28] vdd gnd cell_6t
Xbit_r29_c27 bl[27] br[27] wl[29] vdd gnd cell_6t
Xbit_r30_c27 bl[27] br[27] wl[30] vdd gnd cell_6t
Xbit_r31_c27 bl[27] br[27] wl[31] vdd gnd cell_6t
Xbit_r32_c27 bl[27] br[27] wl[32] vdd gnd cell_6t
Xbit_r33_c27 bl[27] br[27] wl[33] vdd gnd cell_6t
Xbit_r34_c27 bl[27] br[27] wl[34] vdd gnd cell_6t
Xbit_r35_c27 bl[27] br[27] wl[35] vdd gnd cell_6t
Xbit_r36_c27 bl[27] br[27] wl[36] vdd gnd cell_6t
Xbit_r37_c27 bl[27] br[27] wl[37] vdd gnd cell_6t
Xbit_r38_c27 bl[27] br[27] wl[38] vdd gnd cell_6t
Xbit_r39_c27 bl[27] br[27] wl[39] vdd gnd cell_6t
Xbit_r40_c27 bl[27] br[27] wl[40] vdd gnd cell_6t
Xbit_r41_c27 bl[27] br[27] wl[41] vdd gnd cell_6t
Xbit_r42_c27 bl[27] br[27] wl[42] vdd gnd cell_6t
Xbit_r43_c27 bl[27] br[27] wl[43] vdd gnd cell_6t
Xbit_r44_c27 bl[27] br[27] wl[44] vdd gnd cell_6t
Xbit_r45_c27 bl[27] br[27] wl[45] vdd gnd cell_6t
Xbit_r46_c27 bl[27] br[27] wl[46] vdd gnd cell_6t
Xbit_r47_c27 bl[27] br[27] wl[47] vdd gnd cell_6t
Xbit_r48_c27 bl[27] br[27] wl[48] vdd gnd cell_6t
Xbit_r49_c27 bl[27] br[27] wl[49] vdd gnd cell_6t
Xbit_r50_c27 bl[27] br[27] wl[50] vdd gnd cell_6t
Xbit_r51_c27 bl[27] br[27] wl[51] vdd gnd cell_6t
Xbit_r52_c27 bl[27] br[27] wl[52] vdd gnd cell_6t
Xbit_r53_c27 bl[27] br[27] wl[53] vdd gnd cell_6t
Xbit_r54_c27 bl[27] br[27] wl[54] vdd gnd cell_6t
Xbit_r55_c27 bl[27] br[27] wl[55] vdd gnd cell_6t
Xbit_r56_c27 bl[27] br[27] wl[56] vdd gnd cell_6t
Xbit_r57_c27 bl[27] br[27] wl[57] vdd gnd cell_6t
Xbit_r58_c27 bl[27] br[27] wl[58] vdd gnd cell_6t
Xbit_r59_c27 bl[27] br[27] wl[59] vdd gnd cell_6t
Xbit_r60_c27 bl[27] br[27] wl[60] vdd gnd cell_6t
Xbit_r61_c27 bl[27] br[27] wl[61] vdd gnd cell_6t
Xbit_r62_c27 bl[27] br[27] wl[62] vdd gnd cell_6t
Xbit_r63_c27 bl[27] br[27] wl[63] vdd gnd cell_6t
Xbit_r64_c27 bl[27] br[27] wl[64] vdd gnd cell_6t
Xbit_r65_c27 bl[27] br[27] wl[65] vdd gnd cell_6t
Xbit_r66_c27 bl[27] br[27] wl[66] vdd gnd cell_6t
Xbit_r67_c27 bl[27] br[27] wl[67] vdd gnd cell_6t
Xbit_r68_c27 bl[27] br[27] wl[68] vdd gnd cell_6t
Xbit_r69_c27 bl[27] br[27] wl[69] vdd gnd cell_6t
Xbit_r70_c27 bl[27] br[27] wl[70] vdd gnd cell_6t
Xbit_r71_c27 bl[27] br[27] wl[71] vdd gnd cell_6t
Xbit_r72_c27 bl[27] br[27] wl[72] vdd gnd cell_6t
Xbit_r73_c27 bl[27] br[27] wl[73] vdd gnd cell_6t
Xbit_r74_c27 bl[27] br[27] wl[74] vdd gnd cell_6t
Xbit_r75_c27 bl[27] br[27] wl[75] vdd gnd cell_6t
Xbit_r76_c27 bl[27] br[27] wl[76] vdd gnd cell_6t
Xbit_r77_c27 bl[27] br[27] wl[77] vdd gnd cell_6t
Xbit_r78_c27 bl[27] br[27] wl[78] vdd gnd cell_6t
Xbit_r79_c27 bl[27] br[27] wl[79] vdd gnd cell_6t
Xbit_r80_c27 bl[27] br[27] wl[80] vdd gnd cell_6t
Xbit_r81_c27 bl[27] br[27] wl[81] vdd gnd cell_6t
Xbit_r82_c27 bl[27] br[27] wl[82] vdd gnd cell_6t
Xbit_r83_c27 bl[27] br[27] wl[83] vdd gnd cell_6t
Xbit_r84_c27 bl[27] br[27] wl[84] vdd gnd cell_6t
Xbit_r85_c27 bl[27] br[27] wl[85] vdd gnd cell_6t
Xbit_r86_c27 bl[27] br[27] wl[86] vdd gnd cell_6t
Xbit_r87_c27 bl[27] br[27] wl[87] vdd gnd cell_6t
Xbit_r88_c27 bl[27] br[27] wl[88] vdd gnd cell_6t
Xbit_r89_c27 bl[27] br[27] wl[89] vdd gnd cell_6t
Xbit_r90_c27 bl[27] br[27] wl[90] vdd gnd cell_6t
Xbit_r91_c27 bl[27] br[27] wl[91] vdd gnd cell_6t
Xbit_r92_c27 bl[27] br[27] wl[92] vdd gnd cell_6t
Xbit_r93_c27 bl[27] br[27] wl[93] vdd gnd cell_6t
Xbit_r94_c27 bl[27] br[27] wl[94] vdd gnd cell_6t
Xbit_r95_c27 bl[27] br[27] wl[95] vdd gnd cell_6t
Xbit_r96_c27 bl[27] br[27] wl[96] vdd gnd cell_6t
Xbit_r97_c27 bl[27] br[27] wl[97] vdd gnd cell_6t
Xbit_r98_c27 bl[27] br[27] wl[98] vdd gnd cell_6t
Xbit_r99_c27 bl[27] br[27] wl[99] vdd gnd cell_6t
Xbit_r100_c27 bl[27] br[27] wl[100] vdd gnd cell_6t
Xbit_r101_c27 bl[27] br[27] wl[101] vdd gnd cell_6t
Xbit_r102_c27 bl[27] br[27] wl[102] vdd gnd cell_6t
Xbit_r103_c27 bl[27] br[27] wl[103] vdd gnd cell_6t
Xbit_r104_c27 bl[27] br[27] wl[104] vdd gnd cell_6t
Xbit_r105_c27 bl[27] br[27] wl[105] vdd gnd cell_6t
Xbit_r106_c27 bl[27] br[27] wl[106] vdd gnd cell_6t
Xbit_r107_c27 bl[27] br[27] wl[107] vdd gnd cell_6t
Xbit_r108_c27 bl[27] br[27] wl[108] vdd gnd cell_6t
Xbit_r109_c27 bl[27] br[27] wl[109] vdd gnd cell_6t
Xbit_r110_c27 bl[27] br[27] wl[110] vdd gnd cell_6t
Xbit_r111_c27 bl[27] br[27] wl[111] vdd gnd cell_6t
Xbit_r112_c27 bl[27] br[27] wl[112] vdd gnd cell_6t
Xbit_r113_c27 bl[27] br[27] wl[113] vdd gnd cell_6t
Xbit_r114_c27 bl[27] br[27] wl[114] vdd gnd cell_6t
Xbit_r115_c27 bl[27] br[27] wl[115] vdd gnd cell_6t
Xbit_r116_c27 bl[27] br[27] wl[116] vdd gnd cell_6t
Xbit_r117_c27 bl[27] br[27] wl[117] vdd gnd cell_6t
Xbit_r118_c27 bl[27] br[27] wl[118] vdd gnd cell_6t
Xbit_r119_c27 bl[27] br[27] wl[119] vdd gnd cell_6t
Xbit_r120_c27 bl[27] br[27] wl[120] vdd gnd cell_6t
Xbit_r121_c27 bl[27] br[27] wl[121] vdd gnd cell_6t
Xbit_r122_c27 bl[27] br[27] wl[122] vdd gnd cell_6t
Xbit_r123_c27 bl[27] br[27] wl[123] vdd gnd cell_6t
Xbit_r124_c27 bl[27] br[27] wl[124] vdd gnd cell_6t
Xbit_r125_c27 bl[27] br[27] wl[125] vdd gnd cell_6t
Xbit_r126_c27 bl[27] br[27] wl[126] vdd gnd cell_6t
Xbit_r127_c27 bl[27] br[27] wl[127] vdd gnd cell_6t
Xbit_r0_c28 bl[28] br[28] wl[0] vdd gnd cell_6t
Xbit_r1_c28 bl[28] br[28] wl[1] vdd gnd cell_6t
Xbit_r2_c28 bl[28] br[28] wl[2] vdd gnd cell_6t
Xbit_r3_c28 bl[28] br[28] wl[3] vdd gnd cell_6t
Xbit_r4_c28 bl[28] br[28] wl[4] vdd gnd cell_6t
Xbit_r5_c28 bl[28] br[28] wl[5] vdd gnd cell_6t
Xbit_r6_c28 bl[28] br[28] wl[6] vdd gnd cell_6t
Xbit_r7_c28 bl[28] br[28] wl[7] vdd gnd cell_6t
Xbit_r8_c28 bl[28] br[28] wl[8] vdd gnd cell_6t
Xbit_r9_c28 bl[28] br[28] wl[9] vdd gnd cell_6t
Xbit_r10_c28 bl[28] br[28] wl[10] vdd gnd cell_6t
Xbit_r11_c28 bl[28] br[28] wl[11] vdd gnd cell_6t
Xbit_r12_c28 bl[28] br[28] wl[12] vdd gnd cell_6t
Xbit_r13_c28 bl[28] br[28] wl[13] vdd gnd cell_6t
Xbit_r14_c28 bl[28] br[28] wl[14] vdd gnd cell_6t
Xbit_r15_c28 bl[28] br[28] wl[15] vdd gnd cell_6t
Xbit_r16_c28 bl[28] br[28] wl[16] vdd gnd cell_6t
Xbit_r17_c28 bl[28] br[28] wl[17] vdd gnd cell_6t
Xbit_r18_c28 bl[28] br[28] wl[18] vdd gnd cell_6t
Xbit_r19_c28 bl[28] br[28] wl[19] vdd gnd cell_6t
Xbit_r20_c28 bl[28] br[28] wl[20] vdd gnd cell_6t
Xbit_r21_c28 bl[28] br[28] wl[21] vdd gnd cell_6t
Xbit_r22_c28 bl[28] br[28] wl[22] vdd gnd cell_6t
Xbit_r23_c28 bl[28] br[28] wl[23] vdd gnd cell_6t
Xbit_r24_c28 bl[28] br[28] wl[24] vdd gnd cell_6t
Xbit_r25_c28 bl[28] br[28] wl[25] vdd gnd cell_6t
Xbit_r26_c28 bl[28] br[28] wl[26] vdd gnd cell_6t
Xbit_r27_c28 bl[28] br[28] wl[27] vdd gnd cell_6t
Xbit_r28_c28 bl[28] br[28] wl[28] vdd gnd cell_6t
Xbit_r29_c28 bl[28] br[28] wl[29] vdd gnd cell_6t
Xbit_r30_c28 bl[28] br[28] wl[30] vdd gnd cell_6t
Xbit_r31_c28 bl[28] br[28] wl[31] vdd gnd cell_6t
Xbit_r32_c28 bl[28] br[28] wl[32] vdd gnd cell_6t
Xbit_r33_c28 bl[28] br[28] wl[33] vdd gnd cell_6t
Xbit_r34_c28 bl[28] br[28] wl[34] vdd gnd cell_6t
Xbit_r35_c28 bl[28] br[28] wl[35] vdd gnd cell_6t
Xbit_r36_c28 bl[28] br[28] wl[36] vdd gnd cell_6t
Xbit_r37_c28 bl[28] br[28] wl[37] vdd gnd cell_6t
Xbit_r38_c28 bl[28] br[28] wl[38] vdd gnd cell_6t
Xbit_r39_c28 bl[28] br[28] wl[39] vdd gnd cell_6t
Xbit_r40_c28 bl[28] br[28] wl[40] vdd gnd cell_6t
Xbit_r41_c28 bl[28] br[28] wl[41] vdd gnd cell_6t
Xbit_r42_c28 bl[28] br[28] wl[42] vdd gnd cell_6t
Xbit_r43_c28 bl[28] br[28] wl[43] vdd gnd cell_6t
Xbit_r44_c28 bl[28] br[28] wl[44] vdd gnd cell_6t
Xbit_r45_c28 bl[28] br[28] wl[45] vdd gnd cell_6t
Xbit_r46_c28 bl[28] br[28] wl[46] vdd gnd cell_6t
Xbit_r47_c28 bl[28] br[28] wl[47] vdd gnd cell_6t
Xbit_r48_c28 bl[28] br[28] wl[48] vdd gnd cell_6t
Xbit_r49_c28 bl[28] br[28] wl[49] vdd gnd cell_6t
Xbit_r50_c28 bl[28] br[28] wl[50] vdd gnd cell_6t
Xbit_r51_c28 bl[28] br[28] wl[51] vdd gnd cell_6t
Xbit_r52_c28 bl[28] br[28] wl[52] vdd gnd cell_6t
Xbit_r53_c28 bl[28] br[28] wl[53] vdd gnd cell_6t
Xbit_r54_c28 bl[28] br[28] wl[54] vdd gnd cell_6t
Xbit_r55_c28 bl[28] br[28] wl[55] vdd gnd cell_6t
Xbit_r56_c28 bl[28] br[28] wl[56] vdd gnd cell_6t
Xbit_r57_c28 bl[28] br[28] wl[57] vdd gnd cell_6t
Xbit_r58_c28 bl[28] br[28] wl[58] vdd gnd cell_6t
Xbit_r59_c28 bl[28] br[28] wl[59] vdd gnd cell_6t
Xbit_r60_c28 bl[28] br[28] wl[60] vdd gnd cell_6t
Xbit_r61_c28 bl[28] br[28] wl[61] vdd gnd cell_6t
Xbit_r62_c28 bl[28] br[28] wl[62] vdd gnd cell_6t
Xbit_r63_c28 bl[28] br[28] wl[63] vdd gnd cell_6t
Xbit_r64_c28 bl[28] br[28] wl[64] vdd gnd cell_6t
Xbit_r65_c28 bl[28] br[28] wl[65] vdd gnd cell_6t
Xbit_r66_c28 bl[28] br[28] wl[66] vdd gnd cell_6t
Xbit_r67_c28 bl[28] br[28] wl[67] vdd gnd cell_6t
Xbit_r68_c28 bl[28] br[28] wl[68] vdd gnd cell_6t
Xbit_r69_c28 bl[28] br[28] wl[69] vdd gnd cell_6t
Xbit_r70_c28 bl[28] br[28] wl[70] vdd gnd cell_6t
Xbit_r71_c28 bl[28] br[28] wl[71] vdd gnd cell_6t
Xbit_r72_c28 bl[28] br[28] wl[72] vdd gnd cell_6t
Xbit_r73_c28 bl[28] br[28] wl[73] vdd gnd cell_6t
Xbit_r74_c28 bl[28] br[28] wl[74] vdd gnd cell_6t
Xbit_r75_c28 bl[28] br[28] wl[75] vdd gnd cell_6t
Xbit_r76_c28 bl[28] br[28] wl[76] vdd gnd cell_6t
Xbit_r77_c28 bl[28] br[28] wl[77] vdd gnd cell_6t
Xbit_r78_c28 bl[28] br[28] wl[78] vdd gnd cell_6t
Xbit_r79_c28 bl[28] br[28] wl[79] vdd gnd cell_6t
Xbit_r80_c28 bl[28] br[28] wl[80] vdd gnd cell_6t
Xbit_r81_c28 bl[28] br[28] wl[81] vdd gnd cell_6t
Xbit_r82_c28 bl[28] br[28] wl[82] vdd gnd cell_6t
Xbit_r83_c28 bl[28] br[28] wl[83] vdd gnd cell_6t
Xbit_r84_c28 bl[28] br[28] wl[84] vdd gnd cell_6t
Xbit_r85_c28 bl[28] br[28] wl[85] vdd gnd cell_6t
Xbit_r86_c28 bl[28] br[28] wl[86] vdd gnd cell_6t
Xbit_r87_c28 bl[28] br[28] wl[87] vdd gnd cell_6t
Xbit_r88_c28 bl[28] br[28] wl[88] vdd gnd cell_6t
Xbit_r89_c28 bl[28] br[28] wl[89] vdd gnd cell_6t
Xbit_r90_c28 bl[28] br[28] wl[90] vdd gnd cell_6t
Xbit_r91_c28 bl[28] br[28] wl[91] vdd gnd cell_6t
Xbit_r92_c28 bl[28] br[28] wl[92] vdd gnd cell_6t
Xbit_r93_c28 bl[28] br[28] wl[93] vdd gnd cell_6t
Xbit_r94_c28 bl[28] br[28] wl[94] vdd gnd cell_6t
Xbit_r95_c28 bl[28] br[28] wl[95] vdd gnd cell_6t
Xbit_r96_c28 bl[28] br[28] wl[96] vdd gnd cell_6t
Xbit_r97_c28 bl[28] br[28] wl[97] vdd gnd cell_6t
Xbit_r98_c28 bl[28] br[28] wl[98] vdd gnd cell_6t
Xbit_r99_c28 bl[28] br[28] wl[99] vdd gnd cell_6t
Xbit_r100_c28 bl[28] br[28] wl[100] vdd gnd cell_6t
Xbit_r101_c28 bl[28] br[28] wl[101] vdd gnd cell_6t
Xbit_r102_c28 bl[28] br[28] wl[102] vdd gnd cell_6t
Xbit_r103_c28 bl[28] br[28] wl[103] vdd gnd cell_6t
Xbit_r104_c28 bl[28] br[28] wl[104] vdd gnd cell_6t
Xbit_r105_c28 bl[28] br[28] wl[105] vdd gnd cell_6t
Xbit_r106_c28 bl[28] br[28] wl[106] vdd gnd cell_6t
Xbit_r107_c28 bl[28] br[28] wl[107] vdd gnd cell_6t
Xbit_r108_c28 bl[28] br[28] wl[108] vdd gnd cell_6t
Xbit_r109_c28 bl[28] br[28] wl[109] vdd gnd cell_6t
Xbit_r110_c28 bl[28] br[28] wl[110] vdd gnd cell_6t
Xbit_r111_c28 bl[28] br[28] wl[111] vdd gnd cell_6t
Xbit_r112_c28 bl[28] br[28] wl[112] vdd gnd cell_6t
Xbit_r113_c28 bl[28] br[28] wl[113] vdd gnd cell_6t
Xbit_r114_c28 bl[28] br[28] wl[114] vdd gnd cell_6t
Xbit_r115_c28 bl[28] br[28] wl[115] vdd gnd cell_6t
Xbit_r116_c28 bl[28] br[28] wl[116] vdd gnd cell_6t
Xbit_r117_c28 bl[28] br[28] wl[117] vdd gnd cell_6t
Xbit_r118_c28 bl[28] br[28] wl[118] vdd gnd cell_6t
Xbit_r119_c28 bl[28] br[28] wl[119] vdd gnd cell_6t
Xbit_r120_c28 bl[28] br[28] wl[120] vdd gnd cell_6t
Xbit_r121_c28 bl[28] br[28] wl[121] vdd gnd cell_6t
Xbit_r122_c28 bl[28] br[28] wl[122] vdd gnd cell_6t
Xbit_r123_c28 bl[28] br[28] wl[123] vdd gnd cell_6t
Xbit_r124_c28 bl[28] br[28] wl[124] vdd gnd cell_6t
Xbit_r125_c28 bl[28] br[28] wl[125] vdd gnd cell_6t
Xbit_r126_c28 bl[28] br[28] wl[126] vdd gnd cell_6t
Xbit_r127_c28 bl[28] br[28] wl[127] vdd gnd cell_6t
Xbit_r0_c29 bl[29] br[29] wl[0] vdd gnd cell_6t
Xbit_r1_c29 bl[29] br[29] wl[1] vdd gnd cell_6t
Xbit_r2_c29 bl[29] br[29] wl[2] vdd gnd cell_6t
Xbit_r3_c29 bl[29] br[29] wl[3] vdd gnd cell_6t
Xbit_r4_c29 bl[29] br[29] wl[4] vdd gnd cell_6t
Xbit_r5_c29 bl[29] br[29] wl[5] vdd gnd cell_6t
Xbit_r6_c29 bl[29] br[29] wl[6] vdd gnd cell_6t
Xbit_r7_c29 bl[29] br[29] wl[7] vdd gnd cell_6t
Xbit_r8_c29 bl[29] br[29] wl[8] vdd gnd cell_6t
Xbit_r9_c29 bl[29] br[29] wl[9] vdd gnd cell_6t
Xbit_r10_c29 bl[29] br[29] wl[10] vdd gnd cell_6t
Xbit_r11_c29 bl[29] br[29] wl[11] vdd gnd cell_6t
Xbit_r12_c29 bl[29] br[29] wl[12] vdd gnd cell_6t
Xbit_r13_c29 bl[29] br[29] wl[13] vdd gnd cell_6t
Xbit_r14_c29 bl[29] br[29] wl[14] vdd gnd cell_6t
Xbit_r15_c29 bl[29] br[29] wl[15] vdd gnd cell_6t
Xbit_r16_c29 bl[29] br[29] wl[16] vdd gnd cell_6t
Xbit_r17_c29 bl[29] br[29] wl[17] vdd gnd cell_6t
Xbit_r18_c29 bl[29] br[29] wl[18] vdd gnd cell_6t
Xbit_r19_c29 bl[29] br[29] wl[19] vdd gnd cell_6t
Xbit_r20_c29 bl[29] br[29] wl[20] vdd gnd cell_6t
Xbit_r21_c29 bl[29] br[29] wl[21] vdd gnd cell_6t
Xbit_r22_c29 bl[29] br[29] wl[22] vdd gnd cell_6t
Xbit_r23_c29 bl[29] br[29] wl[23] vdd gnd cell_6t
Xbit_r24_c29 bl[29] br[29] wl[24] vdd gnd cell_6t
Xbit_r25_c29 bl[29] br[29] wl[25] vdd gnd cell_6t
Xbit_r26_c29 bl[29] br[29] wl[26] vdd gnd cell_6t
Xbit_r27_c29 bl[29] br[29] wl[27] vdd gnd cell_6t
Xbit_r28_c29 bl[29] br[29] wl[28] vdd gnd cell_6t
Xbit_r29_c29 bl[29] br[29] wl[29] vdd gnd cell_6t
Xbit_r30_c29 bl[29] br[29] wl[30] vdd gnd cell_6t
Xbit_r31_c29 bl[29] br[29] wl[31] vdd gnd cell_6t
Xbit_r32_c29 bl[29] br[29] wl[32] vdd gnd cell_6t
Xbit_r33_c29 bl[29] br[29] wl[33] vdd gnd cell_6t
Xbit_r34_c29 bl[29] br[29] wl[34] vdd gnd cell_6t
Xbit_r35_c29 bl[29] br[29] wl[35] vdd gnd cell_6t
Xbit_r36_c29 bl[29] br[29] wl[36] vdd gnd cell_6t
Xbit_r37_c29 bl[29] br[29] wl[37] vdd gnd cell_6t
Xbit_r38_c29 bl[29] br[29] wl[38] vdd gnd cell_6t
Xbit_r39_c29 bl[29] br[29] wl[39] vdd gnd cell_6t
Xbit_r40_c29 bl[29] br[29] wl[40] vdd gnd cell_6t
Xbit_r41_c29 bl[29] br[29] wl[41] vdd gnd cell_6t
Xbit_r42_c29 bl[29] br[29] wl[42] vdd gnd cell_6t
Xbit_r43_c29 bl[29] br[29] wl[43] vdd gnd cell_6t
Xbit_r44_c29 bl[29] br[29] wl[44] vdd gnd cell_6t
Xbit_r45_c29 bl[29] br[29] wl[45] vdd gnd cell_6t
Xbit_r46_c29 bl[29] br[29] wl[46] vdd gnd cell_6t
Xbit_r47_c29 bl[29] br[29] wl[47] vdd gnd cell_6t
Xbit_r48_c29 bl[29] br[29] wl[48] vdd gnd cell_6t
Xbit_r49_c29 bl[29] br[29] wl[49] vdd gnd cell_6t
Xbit_r50_c29 bl[29] br[29] wl[50] vdd gnd cell_6t
Xbit_r51_c29 bl[29] br[29] wl[51] vdd gnd cell_6t
Xbit_r52_c29 bl[29] br[29] wl[52] vdd gnd cell_6t
Xbit_r53_c29 bl[29] br[29] wl[53] vdd gnd cell_6t
Xbit_r54_c29 bl[29] br[29] wl[54] vdd gnd cell_6t
Xbit_r55_c29 bl[29] br[29] wl[55] vdd gnd cell_6t
Xbit_r56_c29 bl[29] br[29] wl[56] vdd gnd cell_6t
Xbit_r57_c29 bl[29] br[29] wl[57] vdd gnd cell_6t
Xbit_r58_c29 bl[29] br[29] wl[58] vdd gnd cell_6t
Xbit_r59_c29 bl[29] br[29] wl[59] vdd gnd cell_6t
Xbit_r60_c29 bl[29] br[29] wl[60] vdd gnd cell_6t
Xbit_r61_c29 bl[29] br[29] wl[61] vdd gnd cell_6t
Xbit_r62_c29 bl[29] br[29] wl[62] vdd gnd cell_6t
Xbit_r63_c29 bl[29] br[29] wl[63] vdd gnd cell_6t
Xbit_r64_c29 bl[29] br[29] wl[64] vdd gnd cell_6t
Xbit_r65_c29 bl[29] br[29] wl[65] vdd gnd cell_6t
Xbit_r66_c29 bl[29] br[29] wl[66] vdd gnd cell_6t
Xbit_r67_c29 bl[29] br[29] wl[67] vdd gnd cell_6t
Xbit_r68_c29 bl[29] br[29] wl[68] vdd gnd cell_6t
Xbit_r69_c29 bl[29] br[29] wl[69] vdd gnd cell_6t
Xbit_r70_c29 bl[29] br[29] wl[70] vdd gnd cell_6t
Xbit_r71_c29 bl[29] br[29] wl[71] vdd gnd cell_6t
Xbit_r72_c29 bl[29] br[29] wl[72] vdd gnd cell_6t
Xbit_r73_c29 bl[29] br[29] wl[73] vdd gnd cell_6t
Xbit_r74_c29 bl[29] br[29] wl[74] vdd gnd cell_6t
Xbit_r75_c29 bl[29] br[29] wl[75] vdd gnd cell_6t
Xbit_r76_c29 bl[29] br[29] wl[76] vdd gnd cell_6t
Xbit_r77_c29 bl[29] br[29] wl[77] vdd gnd cell_6t
Xbit_r78_c29 bl[29] br[29] wl[78] vdd gnd cell_6t
Xbit_r79_c29 bl[29] br[29] wl[79] vdd gnd cell_6t
Xbit_r80_c29 bl[29] br[29] wl[80] vdd gnd cell_6t
Xbit_r81_c29 bl[29] br[29] wl[81] vdd gnd cell_6t
Xbit_r82_c29 bl[29] br[29] wl[82] vdd gnd cell_6t
Xbit_r83_c29 bl[29] br[29] wl[83] vdd gnd cell_6t
Xbit_r84_c29 bl[29] br[29] wl[84] vdd gnd cell_6t
Xbit_r85_c29 bl[29] br[29] wl[85] vdd gnd cell_6t
Xbit_r86_c29 bl[29] br[29] wl[86] vdd gnd cell_6t
Xbit_r87_c29 bl[29] br[29] wl[87] vdd gnd cell_6t
Xbit_r88_c29 bl[29] br[29] wl[88] vdd gnd cell_6t
Xbit_r89_c29 bl[29] br[29] wl[89] vdd gnd cell_6t
Xbit_r90_c29 bl[29] br[29] wl[90] vdd gnd cell_6t
Xbit_r91_c29 bl[29] br[29] wl[91] vdd gnd cell_6t
Xbit_r92_c29 bl[29] br[29] wl[92] vdd gnd cell_6t
Xbit_r93_c29 bl[29] br[29] wl[93] vdd gnd cell_6t
Xbit_r94_c29 bl[29] br[29] wl[94] vdd gnd cell_6t
Xbit_r95_c29 bl[29] br[29] wl[95] vdd gnd cell_6t
Xbit_r96_c29 bl[29] br[29] wl[96] vdd gnd cell_6t
Xbit_r97_c29 bl[29] br[29] wl[97] vdd gnd cell_6t
Xbit_r98_c29 bl[29] br[29] wl[98] vdd gnd cell_6t
Xbit_r99_c29 bl[29] br[29] wl[99] vdd gnd cell_6t
Xbit_r100_c29 bl[29] br[29] wl[100] vdd gnd cell_6t
Xbit_r101_c29 bl[29] br[29] wl[101] vdd gnd cell_6t
Xbit_r102_c29 bl[29] br[29] wl[102] vdd gnd cell_6t
Xbit_r103_c29 bl[29] br[29] wl[103] vdd gnd cell_6t
Xbit_r104_c29 bl[29] br[29] wl[104] vdd gnd cell_6t
Xbit_r105_c29 bl[29] br[29] wl[105] vdd gnd cell_6t
Xbit_r106_c29 bl[29] br[29] wl[106] vdd gnd cell_6t
Xbit_r107_c29 bl[29] br[29] wl[107] vdd gnd cell_6t
Xbit_r108_c29 bl[29] br[29] wl[108] vdd gnd cell_6t
Xbit_r109_c29 bl[29] br[29] wl[109] vdd gnd cell_6t
Xbit_r110_c29 bl[29] br[29] wl[110] vdd gnd cell_6t
Xbit_r111_c29 bl[29] br[29] wl[111] vdd gnd cell_6t
Xbit_r112_c29 bl[29] br[29] wl[112] vdd gnd cell_6t
Xbit_r113_c29 bl[29] br[29] wl[113] vdd gnd cell_6t
Xbit_r114_c29 bl[29] br[29] wl[114] vdd gnd cell_6t
Xbit_r115_c29 bl[29] br[29] wl[115] vdd gnd cell_6t
Xbit_r116_c29 bl[29] br[29] wl[116] vdd gnd cell_6t
Xbit_r117_c29 bl[29] br[29] wl[117] vdd gnd cell_6t
Xbit_r118_c29 bl[29] br[29] wl[118] vdd gnd cell_6t
Xbit_r119_c29 bl[29] br[29] wl[119] vdd gnd cell_6t
Xbit_r120_c29 bl[29] br[29] wl[120] vdd gnd cell_6t
Xbit_r121_c29 bl[29] br[29] wl[121] vdd gnd cell_6t
Xbit_r122_c29 bl[29] br[29] wl[122] vdd gnd cell_6t
Xbit_r123_c29 bl[29] br[29] wl[123] vdd gnd cell_6t
Xbit_r124_c29 bl[29] br[29] wl[124] vdd gnd cell_6t
Xbit_r125_c29 bl[29] br[29] wl[125] vdd gnd cell_6t
Xbit_r126_c29 bl[29] br[29] wl[126] vdd gnd cell_6t
Xbit_r127_c29 bl[29] br[29] wl[127] vdd gnd cell_6t
Xbit_r0_c30 bl[30] br[30] wl[0] vdd gnd cell_6t
Xbit_r1_c30 bl[30] br[30] wl[1] vdd gnd cell_6t
Xbit_r2_c30 bl[30] br[30] wl[2] vdd gnd cell_6t
Xbit_r3_c30 bl[30] br[30] wl[3] vdd gnd cell_6t
Xbit_r4_c30 bl[30] br[30] wl[4] vdd gnd cell_6t
Xbit_r5_c30 bl[30] br[30] wl[5] vdd gnd cell_6t
Xbit_r6_c30 bl[30] br[30] wl[6] vdd gnd cell_6t
Xbit_r7_c30 bl[30] br[30] wl[7] vdd gnd cell_6t
Xbit_r8_c30 bl[30] br[30] wl[8] vdd gnd cell_6t
Xbit_r9_c30 bl[30] br[30] wl[9] vdd gnd cell_6t
Xbit_r10_c30 bl[30] br[30] wl[10] vdd gnd cell_6t
Xbit_r11_c30 bl[30] br[30] wl[11] vdd gnd cell_6t
Xbit_r12_c30 bl[30] br[30] wl[12] vdd gnd cell_6t
Xbit_r13_c30 bl[30] br[30] wl[13] vdd gnd cell_6t
Xbit_r14_c30 bl[30] br[30] wl[14] vdd gnd cell_6t
Xbit_r15_c30 bl[30] br[30] wl[15] vdd gnd cell_6t
Xbit_r16_c30 bl[30] br[30] wl[16] vdd gnd cell_6t
Xbit_r17_c30 bl[30] br[30] wl[17] vdd gnd cell_6t
Xbit_r18_c30 bl[30] br[30] wl[18] vdd gnd cell_6t
Xbit_r19_c30 bl[30] br[30] wl[19] vdd gnd cell_6t
Xbit_r20_c30 bl[30] br[30] wl[20] vdd gnd cell_6t
Xbit_r21_c30 bl[30] br[30] wl[21] vdd gnd cell_6t
Xbit_r22_c30 bl[30] br[30] wl[22] vdd gnd cell_6t
Xbit_r23_c30 bl[30] br[30] wl[23] vdd gnd cell_6t
Xbit_r24_c30 bl[30] br[30] wl[24] vdd gnd cell_6t
Xbit_r25_c30 bl[30] br[30] wl[25] vdd gnd cell_6t
Xbit_r26_c30 bl[30] br[30] wl[26] vdd gnd cell_6t
Xbit_r27_c30 bl[30] br[30] wl[27] vdd gnd cell_6t
Xbit_r28_c30 bl[30] br[30] wl[28] vdd gnd cell_6t
Xbit_r29_c30 bl[30] br[30] wl[29] vdd gnd cell_6t
Xbit_r30_c30 bl[30] br[30] wl[30] vdd gnd cell_6t
Xbit_r31_c30 bl[30] br[30] wl[31] vdd gnd cell_6t
Xbit_r32_c30 bl[30] br[30] wl[32] vdd gnd cell_6t
Xbit_r33_c30 bl[30] br[30] wl[33] vdd gnd cell_6t
Xbit_r34_c30 bl[30] br[30] wl[34] vdd gnd cell_6t
Xbit_r35_c30 bl[30] br[30] wl[35] vdd gnd cell_6t
Xbit_r36_c30 bl[30] br[30] wl[36] vdd gnd cell_6t
Xbit_r37_c30 bl[30] br[30] wl[37] vdd gnd cell_6t
Xbit_r38_c30 bl[30] br[30] wl[38] vdd gnd cell_6t
Xbit_r39_c30 bl[30] br[30] wl[39] vdd gnd cell_6t
Xbit_r40_c30 bl[30] br[30] wl[40] vdd gnd cell_6t
Xbit_r41_c30 bl[30] br[30] wl[41] vdd gnd cell_6t
Xbit_r42_c30 bl[30] br[30] wl[42] vdd gnd cell_6t
Xbit_r43_c30 bl[30] br[30] wl[43] vdd gnd cell_6t
Xbit_r44_c30 bl[30] br[30] wl[44] vdd gnd cell_6t
Xbit_r45_c30 bl[30] br[30] wl[45] vdd gnd cell_6t
Xbit_r46_c30 bl[30] br[30] wl[46] vdd gnd cell_6t
Xbit_r47_c30 bl[30] br[30] wl[47] vdd gnd cell_6t
Xbit_r48_c30 bl[30] br[30] wl[48] vdd gnd cell_6t
Xbit_r49_c30 bl[30] br[30] wl[49] vdd gnd cell_6t
Xbit_r50_c30 bl[30] br[30] wl[50] vdd gnd cell_6t
Xbit_r51_c30 bl[30] br[30] wl[51] vdd gnd cell_6t
Xbit_r52_c30 bl[30] br[30] wl[52] vdd gnd cell_6t
Xbit_r53_c30 bl[30] br[30] wl[53] vdd gnd cell_6t
Xbit_r54_c30 bl[30] br[30] wl[54] vdd gnd cell_6t
Xbit_r55_c30 bl[30] br[30] wl[55] vdd gnd cell_6t
Xbit_r56_c30 bl[30] br[30] wl[56] vdd gnd cell_6t
Xbit_r57_c30 bl[30] br[30] wl[57] vdd gnd cell_6t
Xbit_r58_c30 bl[30] br[30] wl[58] vdd gnd cell_6t
Xbit_r59_c30 bl[30] br[30] wl[59] vdd gnd cell_6t
Xbit_r60_c30 bl[30] br[30] wl[60] vdd gnd cell_6t
Xbit_r61_c30 bl[30] br[30] wl[61] vdd gnd cell_6t
Xbit_r62_c30 bl[30] br[30] wl[62] vdd gnd cell_6t
Xbit_r63_c30 bl[30] br[30] wl[63] vdd gnd cell_6t
Xbit_r64_c30 bl[30] br[30] wl[64] vdd gnd cell_6t
Xbit_r65_c30 bl[30] br[30] wl[65] vdd gnd cell_6t
Xbit_r66_c30 bl[30] br[30] wl[66] vdd gnd cell_6t
Xbit_r67_c30 bl[30] br[30] wl[67] vdd gnd cell_6t
Xbit_r68_c30 bl[30] br[30] wl[68] vdd gnd cell_6t
Xbit_r69_c30 bl[30] br[30] wl[69] vdd gnd cell_6t
Xbit_r70_c30 bl[30] br[30] wl[70] vdd gnd cell_6t
Xbit_r71_c30 bl[30] br[30] wl[71] vdd gnd cell_6t
Xbit_r72_c30 bl[30] br[30] wl[72] vdd gnd cell_6t
Xbit_r73_c30 bl[30] br[30] wl[73] vdd gnd cell_6t
Xbit_r74_c30 bl[30] br[30] wl[74] vdd gnd cell_6t
Xbit_r75_c30 bl[30] br[30] wl[75] vdd gnd cell_6t
Xbit_r76_c30 bl[30] br[30] wl[76] vdd gnd cell_6t
Xbit_r77_c30 bl[30] br[30] wl[77] vdd gnd cell_6t
Xbit_r78_c30 bl[30] br[30] wl[78] vdd gnd cell_6t
Xbit_r79_c30 bl[30] br[30] wl[79] vdd gnd cell_6t
Xbit_r80_c30 bl[30] br[30] wl[80] vdd gnd cell_6t
Xbit_r81_c30 bl[30] br[30] wl[81] vdd gnd cell_6t
Xbit_r82_c30 bl[30] br[30] wl[82] vdd gnd cell_6t
Xbit_r83_c30 bl[30] br[30] wl[83] vdd gnd cell_6t
Xbit_r84_c30 bl[30] br[30] wl[84] vdd gnd cell_6t
Xbit_r85_c30 bl[30] br[30] wl[85] vdd gnd cell_6t
Xbit_r86_c30 bl[30] br[30] wl[86] vdd gnd cell_6t
Xbit_r87_c30 bl[30] br[30] wl[87] vdd gnd cell_6t
Xbit_r88_c30 bl[30] br[30] wl[88] vdd gnd cell_6t
Xbit_r89_c30 bl[30] br[30] wl[89] vdd gnd cell_6t
Xbit_r90_c30 bl[30] br[30] wl[90] vdd gnd cell_6t
Xbit_r91_c30 bl[30] br[30] wl[91] vdd gnd cell_6t
Xbit_r92_c30 bl[30] br[30] wl[92] vdd gnd cell_6t
Xbit_r93_c30 bl[30] br[30] wl[93] vdd gnd cell_6t
Xbit_r94_c30 bl[30] br[30] wl[94] vdd gnd cell_6t
Xbit_r95_c30 bl[30] br[30] wl[95] vdd gnd cell_6t
Xbit_r96_c30 bl[30] br[30] wl[96] vdd gnd cell_6t
Xbit_r97_c30 bl[30] br[30] wl[97] vdd gnd cell_6t
Xbit_r98_c30 bl[30] br[30] wl[98] vdd gnd cell_6t
Xbit_r99_c30 bl[30] br[30] wl[99] vdd gnd cell_6t
Xbit_r100_c30 bl[30] br[30] wl[100] vdd gnd cell_6t
Xbit_r101_c30 bl[30] br[30] wl[101] vdd gnd cell_6t
Xbit_r102_c30 bl[30] br[30] wl[102] vdd gnd cell_6t
Xbit_r103_c30 bl[30] br[30] wl[103] vdd gnd cell_6t
Xbit_r104_c30 bl[30] br[30] wl[104] vdd gnd cell_6t
Xbit_r105_c30 bl[30] br[30] wl[105] vdd gnd cell_6t
Xbit_r106_c30 bl[30] br[30] wl[106] vdd gnd cell_6t
Xbit_r107_c30 bl[30] br[30] wl[107] vdd gnd cell_6t
Xbit_r108_c30 bl[30] br[30] wl[108] vdd gnd cell_6t
Xbit_r109_c30 bl[30] br[30] wl[109] vdd gnd cell_6t
Xbit_r110_c30 bl[30] br[30] wl[110] vdd gnd cell_6t
Xbit_r111_c30 bl[30] br[30] wl[111] vdd gnd cell_6t
Xbit_r112_c30 bl[30] br[30] wl[112] vdd gnd cell_6t
Xbit_r113_c30 bl[30] br[30] wl[113] vdd gnd cell_6t
Xbit_r114_c30 bl[30] br[30] wl[114] vdd gnd cell_6t
Xbit_r115_c30 bl[30] br[30] wl[115] vdd gnd cell_6t
Xbit_r116_c30 bl[30] br[30] wl[116] vdd gnd cell_6t
Xbit_r117_c30 bl[30] br[30] wl[117] vdd gnd cell_6t
Xbit_r118_c30 bl[30] br[30] wl[118] vdd gnd cell_6t
Xbit_r119_c30 bl[30] br[30] wl[119] vdd gnd cell_6t
Xbit_r120_c30 bl[30] br[30] wl[120] vdd gnd cell_6t
Xbit_r121_c30 bl[30] br[30] wl[121] vdd gnd cell_6t
Xbit_r122_c30 bl[30] br[30] wl[122] vdd gnd cell_6t
Xbit_r123_c30 bl[30] br[30] wl[123] vdd gnd cell_6t
Xbit_r124_c30 bl[30] br[30] wl[124] vdd gnd cell_6t
Xbit_r125_c30 bl[30] br[30] wl[125] vdd gnd cell_6t
Xbit_r126_c30 bl[30] br[30] wl[126] vdd gnd cell_6t
Xbit_r127_c30 bl[30] br[30] wl[127] vdd gnd cell_6t
Xbit_r0_c31 bl[31] br[31] wl[0] vdd gnd cell_6t
Xbit_r1_c31 bl[31] br[31] wl[1] vdd gnd cell_6t
Xbit_r2_c31 bl[31] br[31] wl[2] vdd gnd cell_6t
Xbit_r3_c31 bl[31] br[31] wl[3] vdd gnd cell_6t
Xbit_r4_c31 bl[31] br[31] wl[4] vdd gnd cell_6t
Xbit_r5_c31 bl[31] br[31] wl[5] vdd gnd cell_6t
Xbit_r6_c31 bl[31] br[31] wl[6] vdd gnd cell_6t
Xbit_r7_c31 bl[31] br[31] wl[7] vdd gnd cell_6t
Xbit_r8_c31 bl[31] br[31] wl[8] vdd gnd cell_6t
Xbit_r9_c31 bl[31] br[31] wl[9] vdd gnd cell_6t
Xbit_r10_c31 bl[31] br[31] wl[10] vdd gnd cell_6t
Xbit_r11_c31 bl[31] br[31] wl[11] vdd gnd cell_6t
Xbit_r12_c31 bl[31] br[31] wl[12] vdd gnd cell_6t
Xbit_r13_c31 bl[31] br[31] wl[13] vdd gnd cell_6t
Xbit_r14_c31 bl[31] br[31] wl[14] vdd gnd cell_6t
Xbit_r15_c31 bl[31] br[31] wl[15] vdd gnd cell_6t
Xbit_r16_c31 bl[31] br[31] wl[16] vdd gnd cell_6t
Xbit_r17_c31 bl[31] br[31] wl[17] vdd gnd cell_6t
Xbit_r18_c31 bl[31] br[31] wl[18] vdd gnd cell_6t
Xbit_r19_c31 bl[31] br[31] wl[19] vdd gnd cell_6t
Xbit_r20_c31 bl[31] br[31] wl[20] vdd gnd cell_6t
Xbit_r21_c31 bl[31] br[31] wl[21] vdd gnd cell_6t
Xbit_r22_c31 bl[31] br[31] wl[22] vdd gnd cell_6t
Xbit_r23_c31 bl[31] br[31] wl[23] vdd gnd cell_6t
Xbit_r24_c31 bl[31] br[31] wl[24] vdd gnd cell_6t
Xbit_r25_c31 bl[31] br[31] wl[25] vdd gnd cell_6t
Xbit_r26_c31 bl[31] br[31] wl[26] vdd gnd cell_6t
Xbit_r27_c31 bl[31] br[31] wl[27] vdd gnd cell_6t
Xbit_r28_c31 bl[31] br[31] wl[28] vdd gnd cell_6t
Xbit_r29_c31 bl[31] br[31] wl[29] vdd gnd cell_6t
Xbit_r30_c31 bl[31] br[31] wl[30] vdd gnd cell_6t
Xbit_r31_c31 bl[31] br[31] wl[31] vdd gnd cell_6t
Xbit_r32_c31 bl[31] br[31] wl[32] vdd gnd cell_6t
Xbit_r33_c31 bl[31] br[31] wl[33] vdd gnd cell_6t
Xbit_r34_c31 bl[31] br[31] wl[34] vdd gnd cell_6t
Xbit_r35_c31 bl[31] br[31] wl[35] vdd gnd cell_6t
Xbit_r36_c31 bl[31] br[31] wl[36] vdd gnd cell_6t
Xbit_r37_c31 bl[31] br[31] wl[37] vdd gnd cell_6t
Xbit_r38_c31 bl[31] br[31] wl[38] vdd gnd cell_6t
Xbit_r39_c31 bl[31] br[31] wl[39] vdd gnd cell_6t
Xbit_r40_c31 bl[31] br[31] wl[40] vdd gnd cell_6t
Xbit_r41_c31 bl[31] br[31] wl[41] vdd gnd cell_6t
Xbit_r42_c31 bl[31] br[31] wl[42] vdd gnd cell_6t
Xbit_r43_c31 bl[31] br[31] wl[43] vdd gnd cell_6t
Xbit_r44_c31 bl[31] br[31] wl[44] vdd gnd cell_6t
Xbit_r45_c31 bl[31] br[31] wl[45] vdd gnd cell_6t
Xbit_r46_c31 bl[31] br[31] wl[46] vdd gnd cell_6t
Xbit_r47_c31 bl[31] br[31] wl[47] vdd gnd cell_6t
Xbit_r48_c31 bl[31] br[31] wl[48] vdd gnd cell_6t
Xbit_r49_c31 bl[31] br[31] wl[49] vdd gnd cell_6t
Xbit_r50_c31 bl[31] br[31] wl[50] vdd gnd cell_6t
Xbit_r51_c31 bl[31] br[31] wl[51] vdd gnd cell_6t
Xbit_r52_c31 bl[31] br[31] wl[52] vdd gnd cell_6t
Xbit_r53_c31 bl[31] br[31] wl[53] vdd gnd cell_6t
Xbit_r54_c31 bl[31] br[31] wl[54] vdd gnd cell_6t
Xbit_r55_c31 bl[31] br[31] wl[55] vdd gnd cell_6t
Xbit_r56_c31 bl[31] br[31] wl[56] vdd gnd cell_6t
Xbit_r57_c31 bl[31] br[31] wl[57] vdd gnd cell_6t
Xbit_r58_c31 bl[31] br[31] wl[58] vdd gnd cell_6t
Xbit_r59_c31 bl[31] br[31] wl[59] vdd gnd cell_6t
Xbit_r60_c31 bl[31] br[31] wl[60] vdd gnd cell_6t
Xbit_r61_c31 bl[31] br[31] wl[61] vdd gnd cell_6t
Xbit_r62_c31 bl[31] br[31] wl[62] vdd gnd cell_6t
Xbit_r63_c31 bl[31] br[31] wl[63] vdd gnd cell_6t
Xbit_r64_c31 bl[31] br[31] wl[64] vdd gnd cell_6t
Xbit_r65_c31 bl[31] br[31] wl[65] vdd gnd cell_6t
Xbit_r66_c31 bl[31] br[31] wl[66] vdd gnd cell_6t
Xbit_r67_c31 bl[31] br[31] wl[67] vdd gnd cell_6t
Xbit_r68_c31 bl[31] br[31] wl[68] vdd gnd cell_6t
Xbit_r69_c31 bl[31] br[31] wl[69] vdd gnd cell_6t
Xbit_r70_c31 bl[31] br[31] wl[70] vdd gnd cell_6t
Xbit_r71_c31 bl[31] br[31] wl[71] vdd gnd cell_6t
Xbit_r72_c31 bl[31] br[31] wl[72] vdd gnd cell_6t
Xbit_r73_c31 bl[31] br[31] wl[73] vdd gnd cell_6t
Xbit_r74_c31 bl[31] br[31] wl[74] vdd gnd cell_6t
Xbit_r75_c31 bl[31] br[31] wl[75] vdd gnd cell_6t
Xbit_r76_c31 bl[31] br[31] wl[76] vdd gnd cell_6t
Xbit_r77_c31 bl[31] br[31] wl[77] vdd gnd cell_6t
Xbit_r78_c31 bl[31] br[31] wl[78] vdd gnd cell_6t
Xbit_r79_c31 bl[31] br[31] wl[79] vdd gnd cell_6t
Xbit_r80_c31 bl[31] br[31] wl[80] vdd gnd cell_6t
Xbit_r81_c31 bl[31] br[31] wl[81] vdd gnd cell_6t
Xbit_r82_c31 bl[31] br[31] wl[82] vdd gnd cell_6t
Xbit_r83_c31 bl[31] br[31] wl[83] vdd gnd cell_6t
Xbit_r84_c31 bl[31] br[31] wl[84] vdd gnd cell_6t
Xbit_r85_c31 bl[31] br[31] wl[85] vdd gnd cell_6t
Xbit_r86_c31 bl[31] br[31] wl[86] vdd gnd cell_6t
Xbit_r87_c31 bl[31] br[31] wl[87] vdd gnd cell_6t
Xbit_r88_c31 bl[31] br[31] wl[88] vdd gnd cell_6t
Xbit_r89_c31 bl[31] br[31] wl[89] vdd gnd cell_6t
Xbit_r90_c31 bl[31] br[31] wl[90] vdd gnd cell_6t
Xbit_r91_c31 bl[31] br[31] wl[91] vdd gnd cell_6t
Xbit_r92_c31 bl[31] br[31] wl[92] vdd gnd cell_6t
Xbit_r93_c31 bl[31] br[31] wl[93] vdd gnd cell_6t
Xbit_r94_c31 bl[31] br[31] wl[94] vdd gnd cell_6t
Xbit_r95_c31 bl[31] br[31] wl[95] vdd gnd cell_6t
Xbit_r96_c31 bl[31] br[31] wl[96] vdd gnd cell_6t
Xbit_r97_c31 bl[31] br[31] wl[97] vdd gnd cell_6t
Xbit_r98_c31 bl[31] br[31] wl[98] vdd gnd cell_6t
Xbit_r99_c31 bl[31] br[31] wl[99] vdd gnd cell_6t
Xbit_r100_c31 bl[31] br[31] wl[100] vdd gnd cell_6t
Xbit_r101_c31 bl[31] br[31] wl[101] vdd gnd cell_6t
Xbit_r102_c31 bl[31] br[31] wl[102] vdd gnd cell_6t
Xbit_r103_c31 bl[31] br[31] wl[103] vdd gnd cell_6t
Xbit_r104_c31 bl[31] br[31] wl[104] vdd gnd cell_6t
Xbit_r105_c31 bl[31] br[31] wl[105] vdd gnd cell_6t
Xbit_r106_c31 bl[31] br[31] wl[106] vdd gnd cell_6t
Xbit_r107_c31 bl[31] br[31] wl[107] vdd gnd cell_6t
Xbit_r108_c31 bl[31] br[31] wl[108] vdd gnd cell_6t
Xbit_r109_c31 bl[31] br[31] wl[109] vdd gnd cell_6t
Xbit_r110_c31 bl[31] br[31] wl[110] vdd gnd cell_6t
Xbit_r111_c31 bl[31] br[31] wl[111] vdd gnd cell_6t
Xbit_r112_c31 bl[31] br[31] wl[112] vdd gnd cell_6t
Xbit_r113_c31 bl[31] br[31] wl[113] vdd gnd cell_6t
Xbit_r114_c31 bl[31] br[31] wl[114] vdd gnd cell_6t
Xbit_r115_c31 bl[31] br[31] wl[115] vdd gnd cell_6t
Xbit_r116_c31 bl[31] br[31] wl[116] vdd gnd cell_6t
Xbit_r117_c31 bl[31] br[31] wl[117] vdd gnd cell_6t
Xbit_r118_c31 bl[31] br[31] wl[118] vdd gnd cell_6t
Xbit_r119_c31 bl[31] br[31] wl[119] vdd gnd cell_6t
Xbit_r120_c31 bl[31] br[31] wl[120] vdd gnd cell_6t
Xbit_r121_c31 bl[31] br[31] wl[121] vdd gnd cell_6t
Xbit_r122_c31 bl[31] br[31] wl[122] vdd gnd cell_6t
Xbit_r123_c31 bl[31] br[31] wl[123] vdd gnd cell_6t
Xbit_r124_c31 bl[31] br[31] wl[124] vdd gnd cell_6t
Xbit_r125_c31 bl[31] br[31] wl[125] vdd gnd cell_6t
Xbit_r126_c31 bl[31] br[31] wl[126] vdd gnd cell_6t
Xbit_r127_c31 bl[31] br[31] wl[127] vdd gnd cell_6t
Xbit_r0_c32 bl[32] br[32] wl[0] vdd gnd cell_6t
Xbit_r1_c32 bl[32] br[32] wl[1] vdd gnd cell_6t
Xbit_r2_c32 bl[32] br[32] wl[2] vdd gnd cell_6t
Xbit_r3_c32 bl[32] br[32] wl[3] vdd gnd cell_6t
Xbit_r4_c32 bl[32] br[32] wl[4] vdd gnd cell_6t
Xbit_r5_c32 bl[32] br[32] wl[5] vdd gnd cell_6t
Xbit_r6_c32 bl[32] br[32] wl[6] vdd gnd cell_6t
Xbit_r7_c32 bl[32] br[32] wl[7] vdd gnd cell_6t
Xbit_r8_c32 bl[32] br[32] wl[8] vdd gnd cell_6t
Xbit_r9_c32 bl[32] br[32] wl[9] vdd gnd cell_6t
Xbit_r10_c32 bl[32] br[32] wl[10] vdd gnd cell_6t
Xbit_r11_c32 bl[32] br[32] wl[11] vdd gnd cell_6t
Xbit_r12_c32 bl[32] br[32] wl[12] vdd gnd cell_6t
Xbit_r13_c32 bl[32] br[32] wl[13] vdd gnd cell_6t
Xbit_r14_c32 bl[32] br[32] wl[14] vdd gnd cell_6t
Xbit_r15_c32 bl[32] br[32] wl[15] vdd gnd cell_6t
Xbit_r16_c32 bl[32] br[32] wl[16] vdd gnd cell_6t
Xbit_r17_c32 bl[32] br[32] wl[17] vdd gnd cell_6t
Xbit_r18_c32 bl[32] br[32] wl[18] vdd gnd cell_6t
Xbit_r19_c32 bl[32] br[32] wl[19] vdd gnd cell_6t
Xbit_r20_c32 bl[32] br[32] wl[20] vdd gnd cell_6t
Xbit_r21_c32 bl[32] br[32] wl[21] vdd gnd cell_6t
Xbit_r22_c32 bl[32] br[32] wl[22] vdd gnd cell_6t
Xbit_r23_c32 bl[32] br[32] wl[23] vdd gnd cell_6t
Xbit_r24_c32 bl[32] br[32] wl[24] vdd gnd cell_6t
Xbit_r25_c32 bl[32] br[32] wl[25] vdd gnd cell_6t
Xbit_r26_c32 bl[32] br[32] wl[26] vdd gnd cell_6t
Xbit_r27_c32 bl[32] br[32] wl[27] vdd gnd cell_6t
Xbit_r28_c32 bl[32] br[32] wl[28] vdd gnd cell_6t
Xbit_r29_c32 bl[32] br[32] wl[29] vdd gnd cell_6t
Xbit_r30_c32 bl[32] br[32] wl[30] vdd gnd cell_6t
Xbit_r31_c32 bl[32] br[32] wl[31] vdd gnd cell_6t
Xbit_r32_c32 bl[32] br[32] wl[32] vdd gnd cell_6t
Xbit_r33_c32 bl[32] br[32] wl[33] vdd gnd cell_6t
Xbit_r34_c32 bl[32] br[32] wl[34] vdd gnd cell_6t
Xbit_r35_c32 bl[32] br[32] wl[35] vdd gnd cell_6t
Xbit_r36_c32 bl[32] br[32] wl[36] vdd gnd cell_6t
Xbit_r37_c32 bl[32] br[32] wl[37] vdd gnd cell_6t
Xbit_r38_c32 bl[32] br[32] wl[38] vdd gnd cell_6t
Xbit_r39_c32 bl[32] br[32] wl[39] vdd gnd cell_6t
Xbit_r40_c32 bl[32] br[32] wl[40] vdd gnd cell_6t
Xbit_r41_c32 bl[32] br[32] wl[41] vdd gnd cell_6t
Xbit_r42_c32 bl[32] br[32] wl[42] vdd gnd cell_6t
Xbit_r43_c32 bl[32] br[32] wl[43] vdd gnd cell_6t
Xbit_r44_c32 bl[32] br[32] wl[44] vdd gnd cell_6t
Xbit_r45_c32 bl[32] br[32] wl[45] vdd gnd cell_6t
Xbit_r46_c32 bl[32] br[32] wl[46] vdd gnd cell_6t
Xbit_r47_c32 bl[32] br[32] wl[47] vdd gnd cell_6t
Xbit_r48_c32 bl[32] br[32] wl[48] vdd gnd cell_6t
Xbit_r49_c32 bl[32] br[32] wl[49] vdd gnd cell_6t
Xbit_r50_c32 bl[32] br[32] wl[50] vdd gnd cell_6t
Xbit_r51_c32 bl[32] br[32] wl[51] vdd gnd cell_6t
Xbit_r52_c32 bl[32] br[32] wl[52] vdd gnd cell_6t
Xbit_r53_c32 bl[32] br[32] wl[53] vdd gnd cell_6t
Xbit_r54_c32 bl[32] br[32] wl[54] vdd gnd cell_6t
Xbit_r55_c32 bl[32] br[32] wl[55] vdd gnd cell_6t
Xbit_r56_c32 bl[32] br[32] wl[56] vdd gnd cell_6t
Xbit_r57_c32 bl[32] br[32] wl[57] vdd gnd cell_6t
Xbit_r58_c32 bl[32] br[32] wl[58] vdd gnd cell_6t
Xbit_r59_c32 bl[32] br[32] wl[59] vdd gnd cell_6t
Xbit_r60_c32 bl[32] br[32] wl[60] vdd gnd cell_6t
Xbit_r61_c32 bl[32] br[32] wl[61] vdd gnd cell_6t
Xbit_r62_c32 bl[32] br[32] wl[62] vdd gnd cell_6t
Xbit_r63_c32 bl[32] br[32] wl[63] vdd gnd cell_6t
Xbit_r64_c32 bl[32] br[32] wl[64] vdd gnd cell_6t
Xbit_r65_c32 bl[32] br[32] wl[65] vdd gnd cell_6t
Xbit_r66_c32 bl[32] br[32] wl[66] vdd gnd cell_6t
Xbit_r67_c32 bl[32] br[32] wl[67] vdd gnd cell_6t
Xbit_r68_c32 bl[32] br[32] wl[68] vdd gnd cell_6t
Xbit_r69_c32 bl[32] br[32] wl[69] vdd gnd cell_6t
Xbit_r70_c32 bl[32] br[32] wl[70] vdd gnd cell_6t
Xbit_r71_c32 bl[32] br[32] wl[71] vdd gnd cell_6t
Xbit_r72_c32 bl[32] br[32] wl[72] vdd gnd cell_6t
Xbit_r73_c32 bl[32] br[32] wl[73] vdd gnd cell_6t
Xbit_r74_c32 bl[32] br[32] wl[74] vdd gnd cell_6t
Xbit_r75_c32 bl[32] br[32] wl[75] vdd gnd cell_6t
Xbit_r76_c32 bl[32] br[32] wl[76] vdd gnd cell_6t
Xbit_r77_c32 bl[32] br[32] wl[77] vdd gnd cell_6t
Xbit_r78_c32 bl[32] br[32] wl[78] vdd gnd cell_6t
Xbit_r79_c32 bl[32] br[32] wl[79] vdd gnd cell_6t
Xbit_r80_c32 bl[32] br[32] wl[80] vdd gnd cell_6t
Xbit_r81_c32 bl[32] br[32] wl[81] vdd gnd cell_6t
Xbit_r82_c32 bl[32] br[32] wl[82] vdd gnd cell_6t
Xbit_r83_c32 bl[32] br[32] wl[83] vdd gnd cell_6t
Xbit_r84_c32 bl[32] br[32] wl[84] vdd gnd cell_6t
Xbit_r85_c32 bl[32] br[32] wl[85] vdd gnd cell_6t
Xbit_r86_c32 bl[32] br[32] wl[86] vdd gnd cell_6t
Xbit_r87_c32 bl[32] br[32] wl[87] vdd gnd cell_6t
Xbit_r88_c32 bl[32] br[32] wl[88] vdd gnd cell_6t
Xbit_r89_c32 bl[32] br[32] wl[89] vdd gnd cell_6t
Xbit_r90_c32 bl[32] br[32] wl[90] vdd gnd cell_6t
Xbit_r91_c32 bl[32] br[32] wl[91] vdd gnd cell_6t
Xbit_r92_c32 bl[32] br[32] wl[92] vdd gnd cell_6t
Xbit_r93_c32 bl[32] br[32] wl[93] vdd gnd cell_6t
Xbit_r94_c32 bl[32] br[32] wl[94] vdd gnd cell_6t
Xbit_r95_c32 bl[32] br[32] wl[95] vdd gnd cell_6t
Xbit_r96_c32 bl[32] br[32] wl[96] vdd gnd cell_6t
Xbit_r97_c32 bl[32] br[32] wl[97] vdd gnd cell_6t
Xbit_r98_c32 bl[32] br[32] wl[98] vdd gnd cell_6t
Xbit_r99_c32 bl[32] br[32] wl[99] vdd gnd cell_6t
Xbit_r100_c32 bl[32] br[32] wl[100] vdd gnd cell_6t
Xbit_r101_c32 bl[32] br[32] wl[101] vdd gnd cell_6t
Xbit_r102_c32 bl[32] br[32] wl[102] vdd gnd cell_6t
Xbit_r103_c32 bl[32] br[32] wl[103] vdd gnd cell_6t
Xbit_r104_c32 bl[32] br[32] wl[104] vdd gnd cell_6t
Xbit_r105_c32 bl[32] br[32] wl[105] vdd gnd cell_6t
Xbit_r106_c32 bl[32] br[32] wl[106] vdd gnd cell_6t
Xbit_r107_c32 bl[32] br[32] wl[107] vdd gnd cell_6t
Xbit_r108_c32 bl[32] br[32] wl[108] vdd gnd cell_6t
Xbit_r109_c32 bl[32] br[32] wl[109] vdd gnd cell_6t
Xbit_r110_c32 bl[32] br[32] wl[110] vdd gnd cell_6t
Xbit_r111_c32 bl[32] br[32] wl[111] vdd gnd cell_6t
Xbit_r112_c32 bl[32] br[32] wl[112] vdd gnd cell_6t
Xbit_r113_c32 bl[32] br[32] wl[113] vdd gnd cell_6t
Xbit_r114_c32 bl[32] br[32] wl[114] vdd gnd cell_6t
Xbit_r115_c32 bl[32] br[32] wl[115] vdd gnd cell_6t
Xbit_r116_c32 bl[32] br[32] wl[116] vdd gnd cell_6t
Xbit_r117_c32 bl[32] br[32] wl[117] vdd gnd cell_6t
Xbit_r118_c32 bl[32] br[32] wl[118] vdd gnd cell_6t
Xbit_r119_c32 bl[32] br[32] wl[119] vdd gnd cell_6t
Xbit_r120_c32 bl[32] br[32] wl[120] vdd gnd cell_6t
Xbit_r121_c32 bl[32] br[32] wl[121] vdd gnd cell_6t
Xbit_r122_c32 bl[32] br[32] wl[122] vdd gnd cell_6t
Xbit_r123_c32 bl[32] br[32] wl[123] vdd gnd cell_6t
Xbit_r124_c32 bl[32] br[32] wl[124] vdd gnd cell_6t
Xbit_r125_c32 bl[32] br[32] wl[125] vdd gnd cell_6t
Xbit_r126_c32 bl[32] br[32] wl[126] vdd gnd cell_6t
Xbit_r127_c32 bl[32] br[32] wl[127] vdd gnd cell_6t
Xbit_r0_c33 bl[33] br[33] wl[0] vdd gnd cell_6t
Xbit_r1_c33 bl[33] br[33] wl[1] vdd gnd cell_6t
Xbit_r2_c33 bl[33] br[33] wl[2] vdd gnd cell_6t
Xbit_r3_c33 bl[33] br[33] wl[3] vdd gnd cell_6t
Xbit_r4_c33 bl[33] br[33] wl[4] vdd gnd cell_6t
Xbit_r5_c33 bl[33] br[33] wl[5] vdd gnd cell_6t
Xbit_r6_c33 bl[33] br[33] wl[6] vdd gnd cell_6t
Xbit_r7_c33 bl[33] br[33] wl[7] vdd gnd cell_6t
Xbit_r8_c33 bl[33] br[33] wl[8] vdd gnd cell_6t
Xbit_r9_c33 bl[33] br[33] wl[9] vdd gnd cell_6t
Xbit_r10_c33 bl[33] br[33] wl[10] vdd gnd cell_6t
Xbit_r11_c33 bl[33] br[33] wl[11] vdd gnd cell_6t
Xbit_r12_c33 bl[33] br[33] wl[12] vdd gnd cell_6t
Xbit_r13_c33 bl[33] br[33] wl[13] vdd gnd cell_6t
Xbit_r14_c33 bl[33] br[33] wl[14] vdd gnd cell_6t
Xbit_r15_c33 bl[33] br[33] wl[15] vdd gnd cell_6t
Xbit_r16_c33 bl[33] br[33] wl[16] vdd gnd cell_6t
Xbit_r17_c33 bl[33] br[33] wl[17] vdd gnd cell_6t
Xbit_r18_c33 bl[33] br[33] wl[18] vdd gnd cell_6t
Xbit_r19_c33 bl[33] br[33] wl[19] vdd gnd cell_6t
Xbit_r20_c33 bl[33] br[33] wl[20] vdd gnd cell_6t
Xbit_r21_c33 bl[33] br[33] wl[21] vdd gnd cell_6t
Xbit_r22_c33 bl[33] br[33] wl[22] vdd gnd cell_6t
Xbit_r23_c33 bl[33] br[33] wl[23] vdd gnd cell_6t
Xbit_r24_c33 bl[33] br[33] wl[24] vdd gnd cell_6t
Xbit_r25_c33 bl[33] br[33] wl[25] vdd gnd cell_6t
Xbit_r26_c33 bl[33] br[33] wl[26] vdd gnd cell_6t
Xbit_r27_c33 bl[33] br[33] wl[27] vdd gnd cell_6t
Xbit_r28_c33 bl[33] br[33] wl[28] vdd gnd cell_6t
Xbit_r29_c33 bl[33] br[33] wl[29] vdd gnd cell_6t
Xbit_r30_c33 bl[33] br[33] wl[30] vdd gnd cell_6t
Xbit_r31_c33 bl[33] br[33] wl[31] vdd gnd cell_6t
Xbit_r32_c33 bl[33] br[33] wl[32] vdd gnd cell_6t
Xbit_r33_c33 bl[33] br[33] wl[33] vdd gnd cell_6t
Xbit_r34_c33 bl[33] br[33] wl[34] vdd gnd cell_6t
Xbit_r35_c33 bl[33] br[33] wl[35] vdd gnd cell_6t
Xbit_r36_c33 bl[33] br[33] wl[36] vdd gnd cell_6t
Xbit_r37_c33 bl[33] br[33] wl[37] vdd gnd cell_6t
Xbit_r38_c33 bl[33] br[33] wl[38] vdd gnd cell_6t
Xbit_r39_c33 bl[33] br[33] wl[39] vdd gnd cell_6t
Xbit_r40_c33 bl[33] br[33] wl[40] vdd gnd cell_6t
Xbit_r41_c33 bl[33] br[33] wl[41] vdd gnd cell_6t
Xbit_r42_c33 bl[33] br[33] wl[42] vdd gnd cell_6t
Xbit_r43_c33 bl[33] br[33] wl[43] vdd gnd cell_6t
Xbit_r44_c33 bl[33] br[33] wl[44] vdd gnd cell_6t
Xbit_r45_c33 bl[33] br[33] wl[45] vdd gnd cell_6t
Xbit_r46_c33 bl[33] br[33] wl[46] vdd gnd cell_6t
Xbit_r47_c33 bl[33] br[33] wl[47] vdd gnd cell_6t
Xbit_r48_c33 bl[33] br[33] wl[48] vdd gnd cell_6t
Xbit_r49_c33 bl[33] br[33] wl[49] vdd gnd cell_6t
Xbit_r50_c33 bl[33] br[33] wl[50] vdd gnd cell_6t
Xbit_r51_c33 bl[33] br[33] wl[51] vdd gnd cell_6t
Xbit_r52_c33 bl[33] br[33] wl[52] vdd gnd cell_6t
Xbit_r53_c33 bl[33] br[33] wl[53] vdd gnd cell_6t
Xbit_r54_c33 bl[33] br[33] wl[54] vdd gnd cell_6t
Xbit_r55_c33 bl[33] br[33] wl[55] vdd gnd cell_6t
Xbit_r56_c33 bl[33] br[33] wl[56] vdd gnd cell_6t
Xbit_r57_c33 bl[33] br[33] wl[57] vdd gnd cell_6t
Xbit_r58_c33 bl[33] br[33] wl[58] vdd gnd cell_6t
Xbit_r59_c33 bl[33] br[33] wl[59] vdd gnd cell_6t
Xbit_r60_c33 bl[33] br[33] wl[60] vdd gnd cell_6t
Xbit_r61_c33 bl[33] br[33] wl[61] vdd gnd cell_6t
Xbit_r62_c33 bl[33] br[33] wl[62] vdd gnd cell_6t
Xbit_r63_c33 bl[33] br[33] wl[63] vdd gnd cell_6t
Xbit_r64_c33 bl[33] br[33] wl[64] vdd gnd cell_6t
Xbit_r65_c33 bl[33] br[33] wl[65] vdd gnd cell_6t
Xbit_r66_c33 bl[33] br[33] wl[66] vdd gnd cell_6t
Xbit_r67_c33 bl[33] br[33] wl[67] vdd gnd cell_6t
Xbit_r68_c33 bl[33] br[33] wl[68] vdd gnd cell_6t
Xbit_r69_c33 bl[33] br[33] wl[69] vdd gnd cell_6t
Xbit_r70_c33 bl[33] br[33] wl[70] vdd gnd cell_6t
Xbit_r71_c33 bl[33] br[33] wl[71] vdd gnd cell_6t
Xbit_r72_c33 bl[33] br[33] wl[72] vdd gnd cell_6t
Xbit_r73_c33 bl[33] br[33] wl[73] vdd gnd cell_6t
Xbit_r74_c33 bl[33] br[33] wl[74] vdd gnd cell_6t
Xbit_r75_c33 bl[33] br[33] wl[75] vdd gnd cell_6t
Xbit_r76_c33 bl[33] br[33] wl[76] vdd gnd cell_6t
Xbit_r77_c33 bl[33] br[33] wl[77] vdd gnd cell_6t
Xbit_r78_c33 bl[33] br[33] wl[78] vdd gnd cell_6t
Xbit_r79_c33 bl[33] br[33] wl[79] vdd gnd cell_6t
Xbit_r80_c33 bl[33] br[33] wl[80] vdd gnd cell_6t
Xbit_r81_c33 bl[33] br[33] wl[81] vdd gnd cell_6t
Xbit_r82_c33 bl[33] br[33] wl[82] vdd gnd cell_6t
Xbit_r83_c33 bl[33] br[33] wl[83] vdd gnd cell_6t
Xbit_r84_c33 bl[33] br[33] wl[84] vdd gnd cell_6t
Xbit_r85_c33 bl[33] br[33] wl[85] vdd gnd cell_6t
Xbit_r86_c33 bl[33] br[33] wl[86] vdd gnd cell_6t
Xbit_r87_c33 bl[33] br[33] wl[87] vdd gnd cell_6t
Xbit_r88_c33 bl[33] br[33] wl[88] vdd gnd cell_6t
Xbit_r89_c33 bl[33] br[33] wl[89] vdd gnd cell_6t
Xbit_r90_c33 bl[33] br[33] wl[90] vdd gnd cell_6t
Xbit_r91_c33 bl[33] br[33] wl[91] vdd gnd cell_6t
Xbit_r92_c33 bl[33] br[33] wl[92] vdd gnd cell_6t
Xbit_r93_c33 bl[33] br[33] wl[93] vdd gnd cell_6t
Xbit_r94_c33 bl[33] br[33] wl[94] vdd gnd cell_6t
Xbit_r95_c33 bl[33] br[33] wl[95] vdd gnd cell_6t
Xbit_r96_c33 bl[33] br[33] wl[96] vdd gnd cell_6t
Xbit_r97_c33 bl[33] br[33] wl[97] vdd gnd cell_6t
Xbit_r98_c33 bl[33] br[33] wl[98] vdd gnd cell_6t
Xbit_r99_c33 bl[33] br[33] wl[99] vdd gnd cell_6t
Xbit_r100_c33 bl[33] br[33] wl[100] vdd gnd cell_6t
Xbit_r101_c33 bl[33] br[33] wl[101] vdd gnd cell_6t
Xbit_r102_c33 bl[33] br[33] wl[102] vdd gnd cell_6t
Xbit_r103_c33 bl[33] br[33] wl[103] vdd gnd cell_6t
Xbit_r104_c33 bl[33] br[33] wl[104] vdd gnd cell_6t
Xbit_r105_c33 bl[33] br[33] wl[105] vdd gnd cell_6t
Xbit_r106_c33 bl[33] br[33] wl[106] vdd gnd cell_6t
Xbit_r107_c33 bl[33] br[33] wl[107] vdd gnd cell_6t
Xbit_r108_c33 bl[33] br[33] wl[108] vdd gnd cell_6t
Xbit_r109_c33 bl[33] br[33] wl[109] vdd gnd cell_6t
Xbit_r110_c33 bl[33] br[33] wl[110] vdd gnd cell_6t
Xbit_r111_c33 bl[33] br[33] wl[111] vdd gnd cell_6t
Xbit_r112_c33 bl[33] br[33] wl[112] vdd gnd cell_6t
Xbit_r113_c33 bl[33] br[33] wl[113] vdd gnd cell_6t
Xbit_r114_c33 bl[33] br[33] wl[114] vdd gnd cell_6t
Xbit_r115_c33 bl[33] br[33] wl[115] vdd gnd cell_6t
Xbit_r116_c33 bl[33] br[33] wl[116] vdd gnd cell_6t
Xbit_r117_c33 bl[33] br[33] wl[117] vdd gnd cell_6t
Xbit_r118_c33 bl[33] br[33] wl[118] vdd gnd cell_6t
Xbit_r119_c33 bl[33] br[33] wl[119] vdd gnd cell_6t
Xbit_r120_c33 bl[33] br[33] wl[120] vdd gnd cell_6t
Xbit_r121_c33 bl[33] br[33] wl[121] vdd gnd cell_6t
Xbit_r122_c33 bl[33] br[33] wl[122] vdd gnd cell_6t
Xbit_r123_c33 bl[33] br[33] wl[123] vdd gnd cell_6t
Xbit_r124_c33 bl[33] br[33] wl[124] vdd gnd cell_6t
Xbit_r125_c33 bl[33] br[33] wl[125] vdd gnd cell_6t
Xbit_r126_c33 bl[33] br[33] wl[126] vdd gnd cell_6t
Xbit_r127_c33 bl[33] br[33] wl[127] vdd gnd cell_6t
Xbit_r0_c34 bl[34] br[34] wl[0] vdd gnd cell_6t
Xbit_r1_c34 bl[34] br[34] wl[1] vdd gnd cell_6t
Xbit_r2_c34 bl[34] br[34] wl[2] vdd gnd cell_6t
Xbit_r3_c34 bl[34] br[34] wl[3] vdd gnd cell_6t
Xbit_r4_c34 bl[34] br[34] wl[4] vdd gnd cell_6t
Xbit_r5_c34 bl[34] br[34] wl[5] vdd gnd cell_6t
Xbit_r6_c34 bl[34] br[34] wl[6] vdd gnd cell_6t
Xbit_r7_c34 bl[34] br[34] wl[7] vdd gnd cell_6t
Xbit_r8_c34 bl[34] br[34] wl[8] vdd gnd cell_6t
Xbit_r9_c34 bl[34] br[34] wl[9] vdd gnd cell_6t
Xbit_r10_c34 bl[34] br[34] wl[10] vdd gnd cell_6t
Xbit_r11_c34 bl[34] br[34] wl[11] vdd gnd cell_6t
Xbit_r12_c34 bl[34] br[34] wl[12] vdd gnd cell_6t
Xbit_r13_c34 bl[34] br[34] wl[13] vdd gnd cell_6t
Xbit_r14_c34 bl[34] br[34] wl[14] vdd gnd cell_6t
Xbit_r15_c34 bl[34] br[34] wl[15] vdd gnd cell_6t
Xbit_r16_c34 bl[34] br[34] wl[16] vdd gnd cell_6t
Xbit_r17_c34 bl[34] br[34] wl[17] vdd gnd cell_6t
Xbit_r18_c34 bl[34] br[34] wl[18] vdd gnd cell_6t
Xbit_r19_c34 bl[34] br[34] wl[19] vdd gnd cell_6t
Xbit_r20_c34 bl[34] br[34] wl[20] vdd gnd cell_6t
Xbit_r21_c34 bl[34] br[34] wl[21] vdd gnd cell_6t
Xbit_r22_c34 bl[34] br[34] wl[22] vdd gnd cell_6t
Xbit_r23_c34 bl[34] br[34] wl[23] vdd gnd cell_6t
Xbit_r24_c34 bl[34] br[34] wl[24] vdd gnd cell_6t
Xbit_r25_c34 bl[34] br[34] wl[25] vdd gnd cell_6t
Xbit_r26_c34 bl[34] br[34] wl[26] vdd gnd cell_6t
Xbit_r27_c34 bl[34] br[34] wl[27] vdd gnd cell_6t
Xbit_r28_c34 bl[34] br[34] wl[28] vdd gnd cell_6t
Xbit_r29_c34 bl[34] br[34] wl[29] vdd gnd cell_6t
Xbit_r30_c34 bl[34] br[34] wl[30] vdd gnd cell_6t
Xbit_r31_c34 bl[34] br[34] wl[31] vdd gnd cell_6t
Xbit_r32_c34 bl[34] br[34] wl[32] vdd gnd cell_6t
Xbit_r33_c34 bl[34] br[34] wl[33] vdd gnd cell_6t
Xbit_r34_c34 bl[34] br[34] wl[34] vdd gnd cell_6t
Xbit_r35_c34 bl[34] br[34] wl[35] vdd gnd cell_6t
Xbit_r36_c34 bl[34] br[34] wl[36] vdd gnd cell_6t
Xbit_r37_c34 bl[34] br[34] wl[37] vdd gnd cell_6t
Xbit_r38_c34 bl[34] br[34] wl[38] vdd gnd cell_6t
Xbit_r39_c34 bl[34] br[34] wl[39] vdd gnd cell_6t
Xbit_r40_c34 bl[34] br[34] wl[40] vdd gnd cell_6t
Xbit_r41_c34 bl[34] br[34] wl[41] vdd gnd cell_6t
Xbit_r42_c34 bl[34] br[34] wl[42] vdd gnd cell_6t
Xbit_r43_c34 bl[34] br[34] wl[43] vdd gnd cell_6t
Xbit_r44_c34 bl[34] br[34] wl[44] vdd gnd cell_6t
Xbit_r45_c34 bl[34] br[34] wl[45] vdd gnd cell_6t
Xbit_r46_c34 bl[34] br[34] wl[46] vdd gnd cell_6t
Xbit_r47_c34 bl[34] br[34] wl[47] vdd gnd cell_6t
Xbit_r48_c34 bl[34] br[34] wl[48] vdd gnd cell_6t
Xbit_r49_c34 bl[34] br[34] wl[49] vdd gnd cell_6t
Xbit_r50_c34 bl[34] br[34] wl[50] vdd gnd cell_6t
Xbit_r51_c34 bl[34] br[34] wl[51] vdd gnd cell_6t
Xbit_r52_c34 bl[34] br[34] wl[52] vdd gnd cell_6t
Xbit_r53_c34 bl[34] br[34] wl[53] vdd gnd cell_6t
Xbit_r54_c34 bl[34] br[34] wl[54] vdd gnd cell_6t
Xbit_r55_c34 bl[34] br[34] wl[55] vdd gnd cell_6t
Xbit_r56_c34 bl[34] br[34] wl[56] vdd gnd cell_6t
Xbit_r57_c34 bl[34] br[34] wl[57] vdd gnd cell_6t
Xbit_r58_c34 bl[34] br[34] wl[58] vdd gnd cell_6t
Xbit_r59_c34 bl[34] br[34] wl[59] vdd gnd cell_6t
Xbit_r60_c34 bl[34] br[34] wl[60] vdd gnd cell_6t
Xbit_r61_c34 bl[34] br[34] wl[61] vdd gnd cell_6t
Xbit_r62_c34 bl[34] br[34] wl[62] vdd gnd cell_6t
Xbit_r63_c34 bl[34] br[34] wl[63] vdd gnd cell_6t
Xbit_r64_c34 bl[34] br[34] wl[64] vdd gnd cell_6t
Xbit_r65_c34 bl[34] br[34] wl[65] vdd gnd cell_6t
Xbit_r66_c34 bl[34] br[34] wl[66] vdd gnd cell_6t
Xbit_r67_c34 bl[34] br[34] wl[67] vdd gnd cell_6t
Xbit_r68_c34 bl[34] br[34] wl[68] vdd gnd cell_6t
Xbit_r69_c34 bl[34] br[34] wl[69] vdd gnd cell_6t
Xbit_r70_c34 bl[34] br[34] wl[70] vdd gnd cell_6t
Xbit_r71_c34 bl[34] br[34] wl[71] vdd gnd cell_6t
Xbit_r72_c34 bl[34] br[34] wl[72] vdd gnd cell_6t
Xbit_r73_c34 bl[34] br[34] wl[73] vdd gnd cell_6t
Xbit_r74_c34 bl[34] br[34] wl[74] vdd gnd cell_6t
Xbit_r75_c34 bl[34] br[34] wl[75] vdd gnd cell_6t
Xbit_r76_c34 bl[34] br[34] wl[76] vdd gnd cell_6t
Xbit_r77_c34 bl[34] br[34] wl[77] vdd gnd cell_6t
Xbit_r78_c34 bl[34] br[34] wl[78] vdd gnd cell_6t
Xbit_r79_c34 bl[34] br[34] wl[79] vdd gnd cell_6t
Xbit_r80_c34 bl[34] br[34] wl[80] vdd gnd cell_6t
Xbit_r81_c34 bl[34] br[34] wl[81] vdd gnd cell_6t
Xbit_r82_c34 bl[34] br[34] wl[82] vdd gnd cell_6t
Xbit_r83_c34 bl[34] br[34] wl[83] vdd gnd cell_6t
Xbit_r84_c34 bl[34] br[34] wl[84] vdd gnd cell_6t
Xbit_r85_c34 bl[34] br[34] wl[85] vdd gnd cell_6t
Xbit_r86_c34 bl[34] br[34] wl[86] vdd gnd cell_6t
Xbit_r87_c34 bl[34] br[34] wl[87] vdd gnd cell_6t
Xbit_r88_c34 bl[34] br[34] wl[88] vdd gnd cell_6t
Xbit_r89_c34 bl[34] br[34] wl[89] vdd gnd cell_6t
Xbit_r90_c34 bl[34] br[34] wl[90] vdd gnd cell_6t
Xbit_r91_c34 bl[34] br[34] wl[91] vdd gnd cell_6t
Xbit_r92_c34 bl[34] br[34] wl[92] vdd gnd cell_6t
Xbit_r93_c34 bl[34] br[34] wl[93] vdd gnd cell_6t
Xbit_r94_c34 bl[34] br[34] wl[94] vdd gnd cell_6t
Xbit_r95_c34 bl[34] br[34] wl[95] vdd gnd cell_6t
Xbit_r96_c34 bl[34] br[34] wl[96] vdd gnd cell_6t
Xbit_r97_c34 bl[34] br[34] wl[97] vdd gnd cell_6t
Xbit_r98_c34 bl[34] br[34] wl[98] vdd gnd cell_6t
Xbit_r99_c34 bl[34] br[34] wl[99] vdd gnd cell_6t
Xbit_r100_c34 bl[34] br[34] wl[100] vdd gnd cell_6t
Xbit_r101_c34 bl[34] br[34] wl[101] vdd gnd cell_6t
Xbit_r102_c34 bl[34] br[34] wl[102] vdd gnd cell_6t
Xbit_r103_c34 bl[34] br[34] wl[103] vdd gnd cell_6t
Xbit_r104_c34 bl[34] br[34] wl[104] vdd gnd cell_6t
Xbit_r105_c34 bl[34] br[34] wl[105] vdd gnd cell_6t
Xbit_r106_c34 bl[34] br[34] wl[106] vdd gnd cell_6t
Xbit_r107_c34 bl[34] br[34] wl[107] vdd gnd cell_6t
Xbit_r108_c34 bl[34] br[34] wl[108] vdd gnd cell_6t
Xbit_r109_c34 bl[34] br[34] wl[109] vdd gnd cell_6t
Xbit_r110_c34 bl[34] br[34] wl[110] vdd gnd cell_6t
Xbit_r111_c34 bl[34] br[34] wl[111] vdd gnd cell_6t
Xbit_r112_c34 bl[34] br[34] wl[112] vdd gnd cell_6t
Xbit_r113_c34 bl[34] br[34] wl[113] vdd gnd cell_6t
Xbit_r114_c34 bl[34] br[34] wl[114] vdd gnd cell_6t
Xbit_r115_c34 bl[34] br[34] wl[115] vdd gnd cell_6t
Xbit_r116_c34 bl[34] br[34] wl[116] vdd gnd cell_6t
Xbit_r117_c34 bl[34] br[34] wl[117] vdd gnd cell_6t
Xbit_r118_c34 bl[34] br[34] wl[118] vdd gnd cell_6t
Xbit_r119_c34 bl[34] br[34] wl[119] vdd gnd cell_6t
Xbit_r120_c34 bl[34] br[34] wl[120] vdd gnd cell_6t
Xbit_r121_c34 bl[34] br[34] wl[121] vdd gnd cell_6t
Xbit_r122_c34 bl[34] br[34] wl[122] vdd gnd cell_6t
Xbit_r123_c34 bl[34] br[34] wl[123] vdd gnd cell_6t
Xbit_r124_c34 bl[34] br[34] wl[124] vdd gnd cell_6t
Xbit_r125_c34 bl[34] br[34] wl[125] vdd gnd cell_6t
Xbit_r126_c34 bl[34] br[34] wl[126] vdd gnd cell_6t
Xbit_r127_c34 bl[34] br[34] wl[127] vdd gnd cell_6t
Xbit_r0_c35 bl[35] br[35] wl[0] vdd gnd cell_6t
Xbit_r1_c35 bl[35] br[35] wl[1] vdd gnd cell_6t
Xbit_r2_c35 bl[35] br[35] wl[2] vdd gnd cell_6t
Xbit_r3_c35 bl[35] br[35] wl[3] vdd gnd cell_6t
Xbit_r4_c35 bl[35] br[35] wl[4] vdd gnd cell_6t
Xbit_r5_c35 bl[35] br[35] wl[5] vdd gnd cell_6t
Xbit_r6_c35 bl[35] br[35] wl[6] vdd gnd cell_6t
Xbit_r7_c35 bl[35] br[35] wl[7] vdd gnd cell_6t
Xbit_r8_c35 bl[35] br[35] wl[8] vdd gnd cell_6t
Xbit_r9_c35 bl[35] br[35] wl[9] vdd gnd cell_6t
Xbit_r10_c35 bl[35] br[35] wl[10] vdd gnd cell_6t
Xbit_r11_c35 bl[35] br[35] wl[11] vdd gnd cell_6t
Xbit_r12_c35 bl[35] br[35] wl[12] vdd gnd cell_6t
Xbit_r13_c35 bl[35] br[35] wl[13] vdd gnd cell_6t
Xbit_r14_c35 bl[35] br[35] wl[14] vdd gnd cell_6t
Xbit_r15_c35 bl[35] br[35] wl[15] vdd gnd cell_6t
Xbit_r16_c35 bl[35] br[35] wl[16] vdd gnd cell_6t
Xbit_r17_c35 bl[35] br[35] wl[17] vdd gnd cell_6t
Xbit_r18_c35 bl[35] br[35] wl[18] vdd gnd cell_6t
Xbit_r19_c35 bl[35] br[35] wl[19] vdd gnd cell_6t
Xbit_r20_c35 bl[35] br[35] wl[20] vdd gnd cell_6t
Xbit_r21_c35 bl[35] br[35] wl[21] vdd gnd cell_6t
Xbit_r22_c35 bl[35] br[35] wl[22] vdd gnd cell_6t
Xbit_r23_c35 bl[35] br[35] wl[23] vdd gnd cell_6t
Xbit_r24_c35 bl[35] br[35] wl[24] vdd gnd cell_6t
Xbit_r25_c35 bl[35] br[35] wl[25] vdd gnd cell_6t
Xbit_r26_c35 bl[35] br[35] wl[26] vdd gnd cell_6t
Xbit_r27_c35 bl[35] br[35] wl[27] vdd gnd cell_6t
Xbit_r28_c35 bl[35] br[35] wl[28] vdd gnd cell_6t
Xbit_r29_c35 bl[35] br[35] wl[29] vdd gnd cell_6t
Xbit_r30_c35 bl[35] br[35] wl[30] vdd gnd cell_6t
Xbit_r31_c35 bl[35] br[35] wl[31] vdd gnd cell_6t
Xbit_r32_c35 bl[35] br[35] wl[32] vdd gnd cell_6t
Xbit_r33_c35 bl[35] br[35] wl[33] vdd gnd cell_6t
Xbit_r34_c35 bl[35] br[35] wl[34] vdd gnd cell_6t
Xbit_r35_c35 bl[35] br[35] wl[35] vdd gnd cell_6t
Xbit_r36_c35 bl[35] br[35] wl[36] vdd gnd cell_6t
Xbit_r37_c35 bl[35] br[35] wl[37] vdd gnd cell_6t
Xbit_r38_c35 bl[35] br[35] wl[38] vdd gnd cell_6t
Xbit_r39_c35 bl[35] br[35] wl[39] vdd gnd cell_6t
Xbit_r40_c35 bl[35] br[35] wl[40] vdd gnd cell_6t
Xbit_r41_c35 bl[35] br[35] wl[41] vdd gnd cell_6t
Xbit_r42_c35 bl[35] br[35] wl[42] vdd gnd cell_6t
Xbit_r43_c35 bl[35] br[35] wl[43] vdd gnd cell_6t
Xbit_r44_c35 bl[35] br[35] wl[44] vdd gnd cell_6t
Xbit_r45_c35 bl[35] br[35] wl[45] vdd gnd cell_6t
Xbit_r46_c35 bl[35] br[35] wl[46] vdd gnd cell_6t
Xbit_r47_c35 bl[35] br[35] wl[47] vdd gnd cell_6t
Xbit_r48_c35 bl[35] br[35] wl[48] vdd gnd cell_6t
Xbit_r49_c35 bl[35] br[35] wl[49] vdd gnd cell_6t
Xbit_r50_c35 bl[35] br[35] wl[50] vdd gnd cell_6t
Xbit_r51_c35 bl[35] br[35] wl[51] vdd gnd cell_6t
Xbit_r52_c35 bl[35] br[35] wl[52] vdd gnd cell_6t
Xbit_r53_c35 bl[35] br[35] wl[53] vdd gnd cell_6t
Xbit_r54_c35 bl[35] br[35] wl[54] vdd gnd cell_6t
Xbit_r55_c35 bl[35] br[35] wl[55] vdd gnd cell_6t
Xbit_r56_c35 bl[35] br[35] wl[56] vdd gnd cell_6t
Xbit_r57_c35 bl[35] br[35] wl[57] vdd gnd cell_6t
Xbit_r58_c35 bl[35] br[35] wl[58] vdd gnd cell_6t
Xbit_r59_c35 bl[35] br[35] wl[59] vdd gnd cell_6t
Xbit_r60_c35 bl[35] br[35] wl[60] vdd gnd cell_6t
Xbit_r61_c35 bl[35] br[35] wl[61] vdd gnd cell_6t
Xbit_r62_c35 bl[35] br[35] wl[62] vdd gnd cell_6t
Xbit_r63_c35 bl[35] br[35] wl[63] vdd gnd cell_6t
Xbit_r64_c35 bl[35] br[35] wl[64] vdd gnd cell_6t
Xbit_r65_c35 bl[35] br[35] wl[65] vdd gnd cell_6t
Xbit_r66_c35 bl[35] br[35] wl[66] vdd gnd cell_6t
Xbit_r67_c35 bl[35] br[35] wl[67] vdd gnd cell_6t
Xbit_r68_c35 bl[35] br[35] wl[68] vdd gnd cell_6t
Xbit_r69_c35 bl[35] br[35] wl[69] vdd gnd cell_6t
Xbit_r70_c35 bl[35] br[35] wl[70] vdd gnd cell_6t
Xbit_r71_c35 bl[35] br[35] wl[71] vdd gnd cell_6t
Xbit_r72_c35 bl[35] br[35] wl[72] vdd gnd cell_6t
Xbit_r73_c35 bl[35] br[35] wl[73] vdd gnd cell_6t
Xbit_r74_c35 bl[35] br[35] wl[74] vdd gnd cell_6t
Xbit_r75_c35 bl[35] br[35] wl[75] vdd gnd cell_6t
Xbit_r76_c35 bl[35] br[35] wl[76] vdd gnd cell_6t
Xbit_r77_c35 bl[35] br[35] wl[77] vdd gnd cell_6t
Xbit_r78_c35 bl[35] br[35] wl[78] vdd gnd cell_6t
Xbit_r79_c35 bl[35] br[35] wl[79] vdd gnd cell_6t
Xbit_r80_c35 bl[35] br[35] wl[80] vdd gnd cell_6t
Xbit_r81_c35 bl[35] br[35] wl[81] vdd gnd cell_6t
Xbit_r82_c35 bl[35] br[35] wl[82] vdd gnd cell_6t
Xbit_r83_c35 bl[35] br[35] wl[83] vdd gnd cell_6t
Xbit_r84_c35 bl[35] br[35] wl[84] vdd gnd cell_6t
Xbit_r85_c35 bl[35] br[35] wl[85] vdd gnd cell_6t
Xbit_r86_c35 bl[35] br[35] wl[86] vdd gnd cell_6t
Xbit_r87_c35 bl[35] br[35] wl[87] vdd gnd cell_6t
Xbit_r88_c35 bl[35] br[35] wl[88] vdd gnd cell_6t
Xbit_r89_c35 bl[35] br[35] wl[89] vdd gnd cell_6t
Xbit_r90_c35 bl[35] br[35] wl[90] vdd gnd cell_6t
Xbit_r91_c35 bl[35] br[35] wl[91] vdd gnd cell_6t
Xbit_r92_c35 bl[35] br[35] wl[92] vdd gnd cell_6t
Xbit_r93_c35 bl[35] br[35] wl[93] vdd gnd cell_6t
Xbit_r94_c35 bl[35] br[35] wl[94] vdd gnd cell_6t
Xbit_r95_c35 bl[35] br[35] wl[95] vdd gnd cell_6t
Xbit_r96_c35 bl[35] br[35] wl[96] vdd gnd cell_6t
Xbit_r97_c35 bl[35] br[35] wl[97] vdd gnd cell_6t
Xbit_r98_c35 bl[35] br[35] wl[98] vdd gnd cell_6t
Xbit_r99_c35 bl[35] br[35] wl[99] vdd gnd cell_6t
Xbit_r100_c35 bl[35] br[35] wl[100] vdd gnd cell_6t
Xbit_r101_c35 bl[35] br[35] wl[101] vdd gnd cell_6t
Xbit_r102_c35 bl[35] br[35] wl[102] vdd gnd cell_6t
Xbit_r103_c35 bl[35] br[35] wl[103] vdd gnd cell_6t
Xbit_r104_c35 bl[35] br[35] wl[104] vdd gnd cell_6t
Xbit_r105_c35 bl[35] br[35] wl[105] vdd gnd cell_6t
Xbit_r106_c35 bl[35] br[35] wl[106] vdd gnd cell_6t
Xbit_r107_c35 bl[35] br[35] wl[107] vdd gnd cell_6t
Xbit_r108_c35 bl[35] br[35] wl[108] vdd gnd cell_6t
Xbit_r109_c35 bl[35] br[35] wl[109] vdd gnd cell_6t
Xbit_r110_c35 bl[35] br[35] wl[110] vdd gnd cell_6t
Xbit_r111_c35 bl[35] br[35] wl[111] vdd gnd cell_6t
Xbit_r112_c35 bl[35] br[35] wl[112] vdd gnd cell_6t
Xbit_r113_c35 bl[35] br[35] wl[113] vdd gnd cell_6t
Xbit_r114_c35 bl[35] br[35] wl[114] vdd gnd cell_6t
Xbit_r115_c35 bl[35] br[35] wl[115] vdd gnd cell_6t
Xbit_r116_c35 bl[35] br[35] wl[116] vdd gnd cell_6t
Xbit_r117_c35 bl[35] br[35] wl[117] vdd gnd cell_6t
Xbit_r118_c35 bl[35] br[35] wl[118] vdd gnd cell_6t
Xbit_r119_c35 bl[35] br[35] wl[119] vdd gnd cell_6t
Xbit_r120_c35 bl[35] br[35] wl[120] vdd gnd cell_6t
Xbit_r121_c35 bl[35] br[35] wl[121] vdd gnd cell_6t
Xbit_r122_c35 bl[35] br[35] wl[122] vdd gnd cell_6t
Xbit_r123_c35 bl[35] br[35] wl[123] vdd gnd cell_6t
Xbit_r124_c35 bl[35] br[35] wl[124] vdd gnd cell_6t
Xbit_r125_c35 bl[35] br[35] wl[125] vdd gnd cell_6t
Xbit_r126_c35 bl[35] br[35] wl[126] vdd gnd cell_6t
Xbit_r127_c35 bl[35] br[35] wl[127] vdd gnd cell_6t
Xbit_r0_c36 bl[36] br[36] wl[0] vdd gnd cell_6t
Xbit_r1_c36 bl[36] br[36] wl[1] vdd gnd cell_6t
Xbit_r2_c36 bl[36] br[36] wl[2] vdd gnd cell_6t
Xbit_r3_c36 bl[36] br[36] wl[3] vdd gnd cell_6t
Xbit_r4_c36 bl[36] br[36] wl[4] vdd gnd cell_6t
Xbit_r5_c36 bl[36] br[36] wl[5] vdd gnd cell_6t
Xbit_r6_c36 bl[36] br[36] wl[6] vdd gnd cell_6t
Xbit_r7_c36 bl[36] br[36] wl[7] vdd gnd cell_6t
Xbit_r8_c36 bl[36] br[36] wl[8] vdd gnd cell_6t
Xbit_r9_c36 bl[36] br[36] wl[9] vdd gnd cell_6t
Xbit_r10_c36 bl[36] br[36] wl[10] vdd gnd cell_6t
Xbit_r11_c36 bl[36] br[36] wl[11] vdd gnd cell_6t
Xbit_r12_c36 bl[36] br[36] wl[12] vdd gnd cell_6t
Xbit_r13_c36 bl[36] br[36] wl[13] vdd gnd cell_6t
Xbit_r14_c36 bl[36] br[36] wl[14] vdd gnd cell_6t
Xbit_r15_c36 bl[36] br[36] wl[15] vdd gnd cell_6t
Xbit_r16_c36 bl[36] br[36] wl[16] vdd gnd cell_6t
Xbit_r17_c36 bl[36] br[36] wl[17] vdd gnd cell_6t
Xbit_r18_c36 bl[36] br[36] wl[18] vdd gnd cell_6t
Xbit_r19_c36 bl[36] br[36] wl[19] vdd gnd cell_6t
Xbit_r20_c36 bl[36] br[36] wl[20] vdd gnd cell_6t
Xbit_r21_c36 bl[36] br[36] wl[21] vdd gnd cell_6t
Xbit_r22_c36 bl[36] br[36] wl[22] vdd gnd cell_6t
Xbit_r23_c36 bl[36] br[36] wl[23] vdd gnd cell_6t
Xbit_r24_c36 bl[36] br[36] wl[24] vdd gnd cell_6t
Xbit_r25_c36 bl[36] br[36] wl[25] vdd gnd cell_6t
Xbit_r26_c36 bl[36] br[36] wl[26] vdd gnd cell_6t
Xbit_r27_c36 bl[36] br[36] wl[27] vdd gnd cell_6t
Xbit_r28_c36 bl[36] br[36] wl[28] vdd gnd cell_6t
Xbit_r29_c36 bl[36] br[36] wl[29] vdd gnd cell_6t
Xbit_r30_c36 bl[36] br[36] wl[30] vdd gnd cell_6t
Xbit_r31_c36 bl[36] br[36] wl[31] vdd gnd cell_6t
Xbit_r32_c36 bl[36] br[36] wl[32] vdd gnd cell_6t
Xbit_r33_c36 bl[36] br[36] wl[33] vdd gnd cell_6t
Xbit_r34_c36 bl[36] br[36] wl[34] vdd gnd cell_6t
Xbit_r35_c36 bl[36] br[36] wl[35] vdd gnd cell_6t
Xbit_r36_c36 bl[36] br[36] wl[36] vdd gnd cell_6t
Xbit_r37_c36 bl[36] br[36] wl[37] vdd gnd cell_6t
Xbit_r38_c36 bl[36] br[36] wl[38] vdd gnd cell_6t
Xbit_r39_c36 bl[36] br[36] wl[39] vdd gnd cell_6t
Xbit_r40_c36 bl[36] br[36] wl[40] vdd gnd cell_6t
Xbit_r41_c36 bl[36] br[36] wl[41] vdd gnd cell_6t
Xbit_r42_c36 bl[36] br[36] wl[42] vdd gnd cell_6t
Xbit_r43_c36 bl[36] br[36] wl[43] vdd gnd cell_6t
Xbit_r44_c36 bl[36] br[36] wl[44] vdd gnd cell_6t
Xbit_r45_c36 bl[36] br[36] wl[45] vdd gnd cell_6t
Xbit_r46_c36 bl[36] br[36] wl[46] vdd gnd cell_6t
Xbit_r47_c36 bl[36] br[36] wl[47] vdd gnd cell_6t
Xbit_r48_c36 bl[36] br[36] wl[48] vdd gnd cell_6t
Xbit_r49_c36 bl[36] br[36] wl[49] vdd gnd cell_6t
Xbit_r50_c36 bl[36] br[36] wl[50] vdd gnd cell_6t
Xbit_r51_c36 bl[36] br[36] wl[51] vdd gnd cell_6t
Xbit_r52_c36 bl[36] br[36] wl[52] vdd gnd cell_6t
Xbit_r53_c36 bl[36] br[36] wl[53] vdd gnd cell_6t
Xbit_r54_c36 bl[36] br[36] wl[54] vdd gnd cell_6t
Xbit_r55_c36 bl[36] br[36] wl[55] vdd gnd cell_6t
Xbit_r56_c36 bl[36] br[36] wl[56] vdd gnd cell_6t
Xbit_r57_c36 bl[36] br[36] wl[57] vdd gnd cell_6t
Xbit_r58_c36 bl[36] br[36] wl[58] vdd gnd cell_6t
Xbit_r59_c36 bl[36] br[36] wl[59] vdd gnd cell_6t
Xbit_r60_c36 bl[36] br[36] wl[60] vdd gnd cell_6t
Xbit_r61_c36 bl[36] br[36] wl[61] vdd gnd cell_6t
Xbit_r62_c36 bl[36] br[36] wl[62] vdd gnd cell_6t
Xbit_r63_c36 bl[36] br[36] wl[63] vdd gnd cell_6t
Xbit_r64_c36 bl[36] br[36] wl[64] vdd gnd cell_6t
Xbit_r65_c36 bl[36] br[36] wl[65] vdd gnd cell_6t
Xbit_r66_c36 bl[36] br[36] wl[66] vdd gnd cell_6t
Xbit_r67_c36 bl[36] br[36] wl[67] vdd gnd cell_6t
Xbit_r68_c36 bl[36] br[36] wl[68] vdd gnd cell_6t
Xbit_r69_c36 bl[36] br[36] wl[69] vdd gnd cell_6t
Xbit_r70_c36 bl[36] br[36] wl[70] vdd gnd cell_6t
Xbit_r71_c36 bl[36] br[36] wl[71] vdd gnd cell_6t
Xbit_r72_c36 bl[36] br[36] wl[72] vdd gnd cell_6t
Xbit_r73_c36 bl[36] br[36] wl[73] vdd gnd cell_6t
Xbit_r74_c36 bl[36] br[36] wl[74] vdd gnd cell_6t
Xbit_r75_c36 bl[36] br[36] wl[75] vdd gnd cell_6t
Xbit_r76_c36 bl[36] br[36] wl[76] vdd gnd cell_6t
Xbit_r77_c36 bl[36] br[36] wl[77] vdd gnd cell_6t
Xbit_r78_c36 bl[36] br[36] wl[78] vdd gnd cell_6t
Xbit_r79_c36 bl[36] br[36] wl[79] vdd gnd cell_6t
Xbit_r80_c36 bl[36] br[36] wl[80] vdd gnd cell_6t
Xbit_r81_c36 bl[36] br[36] wl[81] vdd gnd cell_6t
Xbit_r82_c36 bl[36] br[36] wl[82] vdd gnd cell_6t
Xbit_r83_c36 bl[36] br[36] wl[83] vdd gnd cell_6t
Xbit_r84_c36 bl[36] br[36] wl[84] vdd gnd cell_6t
Xbit_r85_c36 bl[36] br[36] wl[85] vdd gnd cell_6t
Xbit_r86_c36 bl[36] br[36] wl[86] vdd gnd cell_6t
Xbit_r87_c36 bl[36] br[36] wl[87] vdd gnd cell_6t
Xbit_r88_c36 bl[36] br[36] wl[88] vdd gnd cell_6t
Xbit_r89_c36 bl[36] br[36] wl[89] vdd gnd cell_6t
Xbit_r90_c36 bl[36] br[36] wl[90] vdd gnd cell_6t
Xbit_r91_c36 bl[36] br[36] wl[91] vdd gnd cell_6t
Xbit_r92_c36 bl[36] br[36] wl[92] vdd gnd cell_6t
Xbit_r93_c36 bl[36] br[36] wl[93] vdd gnd cell_6t
Xbit_r94_c36 bl[36] br[36] wl[94] vdd gnd cell_6t
Xbit_r95_c36 bl[36] br[36] wl[95] vdd gnd cell_6t
Xbit_r96_c36 bl[36] br[36] wl[96] vdd gnd cell_6t
Xbit_r97_c36 bl[36] br[36] wl[97] vdd gnd cell_6t
Xbit_r98_c36 bl[36] br[36] wl[98] vdd gnd cell_6t
Xbit_r99_c36 bl[36] br[36] wl[99] vdd gnd cell_6t
Xbit_r100_c36 bl[36] br[36] wl[100] vdd gnd cell_6t
Xbit_r101_c36 bl[36] br[36] wl[101] vdd gnd cell_6t
Xbit_r102_c36 bl[36] br[36] wl[102] vdd gnd cell_6t
Xbit_r103_c36 bl[36] br[36] wl[103] vdd gnd cell_6t
Xbit_r104_c36 bl[36] br[36] wl[104] vdd gnd cell_6t
Xbit_r105_c36 bl[36] br[36] wl[105] vdd gnd cell_6t
Xbit_r106_c36 bl[36] br[36] wl[106] vdd gnd cell_6t
Xbit_r107_c36 bl[36] br[36] wl[107] vdd gnd cell_6t
Xbit_r108_c36 bl[36] br[36] wl[108] vdd gnd cell_6t
Xbit_r109_c36 bl[36] br[36] wl[109] vdd gnd cell_6t
Xbit_r110_c36 bl[36] br[36] wl[110] vdd gnd cell_6t
Xbit_r111_c36 bl[36] br[36] wl[111] vdd gnd cell_6t
Xbit_r112_c36 bl[36] br[36] wl[112] vdd gnd cell_6t
Xbit_r113_c36 bl[36] br[36] wl[113] vdd gnd cell_6t
Xbit_r114_c36 bl[36] br[36] wl[114] vdd gnd cell_6t
Xbit_r115_c36 bl[36] br[36] wl[115] vdd gnd cell_6t
Xbit_r116_c36 bl[36] br[36] wl[116] vdd gnd cell_6t
Xbit_r117_c36 bl[36] br[36] wl[117] vdd gnd cell_6t
Xbit_r118_c36 bl[36] br[36] wl[118] vdd gnd cell_6t
Xbit_r119_c36 bl[36] br[36] wl[119] vdd gnd cell_6t
Xbit_r120_c36 bl[36] br[36] wl[120] vdd gnd cell_6t
Xbit_r121_c36 bl[36] br[36] wl[121] vdd gnd cell_6t
Xbit_r122_c36 bl[36] br[36] wl[122] vdd gnd cell_6t
Xbit_r123_c36 bl[36] br[36] wl[123] vdd gnd cell_6t
Xbit_r124_c36 bl[36] br[36] wl[124] vdd gnd cell_6t
Xbit_r125_c36 bl[36] br[36] wl[125] vdd gnd cell_6t
Xbit_r126_c36 bl[36] br[36] wl[126] vdd gnd cell_6t
Xbit_r127_c36 bl[36] br[36] wl[127] vdd gnd cell_6t
Xbit_r0_c37 bl[37] br[37] wl[0] vdd gnd cell_6t
Xbit_r1_c37 bl[37] br[37] wl[1] vdd gnd cell_6t
Xbit_r2_c37 bl[37] br[37] wl[2] vdd gnd cell_6t
Xbit_r3_c37 bl[37] br[37] wl[3] vdd gnd cell_6t
Xbit_r4_c37 bl[37] br[37] wl[4] vdd gnd cell_6t
Xbit_r5_c37 bl[37] br[37] wl[5] vdd gnd cell_6t
Xbit_r6_c37 bl[37] br[37] wl[6] vdd gnd cell_6t
Xbit_r7_c37 bl[37] br[37] wl[7] vdd gnd cell_6t
Xbit_r8_c37 bl[37] br[37] wl[8] vdd gnd cell_6t
Xbit_r9_c37 bl[37] br[37] wl[9] vdd gnd cell_6t
Xbit_r10_c37 bl[37] br[37] wl[10] vdd gnd cell_6t
Xbit_r11_c37 bl[37] br[37] wl[11] vdd gnd cell_6t
Xbit_r12_c37 bl[37] br[37] wl[12] vdd gnd cell_6t
Xbit_r13_c37 bl[37] br[37] wl[13] vdd gnd cell_6t
Xbit_r14_c37 bl[37] br[37] wl[14] vdd gnd cell_6t
Xbit_r15_c37 bl[37] br[37] wl[15] vdd gnd cell_6t
Xbit_r16_c37 bl[37] br[37] wl[16] vdd gnd cell_6t
Xbit_r17_c37 bl[37] br[37] wl[17] vdd gnd cell_6t
Xbit_r18_c37 bl[37] br[37] wl[18] vdd gnd cell_6t
Xbit_r19_c37 bl[37] br[37] wl[19] vdd gnd cell_6t
Xbit_r20_c37 bl[37] br[37] wl[20] vdd gnd cell_6t
Xbit_r21_c37 bl[37] br[37] wl[21] vdd gnd cell_6t
Xbit_r22_c37 bl[37] br[37] wl[22] vdd gnd cell_6t
Xbit_r23_c37 bl[37] br[37] wl[23] vdd gnd cell_6t
Xbit_r24_c37 bl[37] br[37] wl[24] vdd gnd cell_6t
Xbit_r25_c37 bl[37] br[37] wl[25] vdd gnd cell_6t
Xbit_r26_c37 bl[37] br[37] wl[26] vdd gnd cell_6t
Xbit_r27_c37 bl[37] br[37] wl[27] vdd gnd cell_6t
Xbit_r28_c37 bl[37] br[37] wl[28] vdd gnd cell_6t
Xbit_r29_c37 bl[37] br[37] wl[29] vdd gnd cell_6t
Xbit_r30_c37 bl[37] br[37] wl[30] vdd gnd cell_6t
Xbit_r31_c37 bl[37] br[37] wl[31] vdd gnd cell_6t
Xbit_r32_c37 bl[37] br[37] wl[32] vdd gnd cell_6t
Xbit_r33_c37 bl[37] br[37] wl[33] vdd gnd cell_6t
Xbit_r34_c37 bl[37] br[37] wl[34] vdd gnd cell_6t
Xbit_r35_c37 bl[37] br[37] wl[35] vdd gnd cell_6t
Xbit_r36_c37 bl[37] br[37] wl[36] vdd gnd cell_6t
Xbit_r37_c37 bl[37] br[37] wl[37] vdd gnd cell_6t
Xbit_r38_c37 bl[37] br[37] wl[38] vdd gnd cell_6t
Xbit_r39_c37 bl[37] br[37] wl[39] vdd gnd cell_6t
Xbit_r40_c37 bl[37] br[37] wl[40] vdd gnd cell_6t
Xbit_r41_c37 bl[37] br[37] wl[41] vdd gnd cell_6t
Xbit_r42_c37 bl[37] br[37] wl[42] vdd gnd cell_6t
Xbit_r43_c37 bl[37] br[37] wl[43] vdd gnd cell_6t
Xbit_r44_c37 bl[37] br[37] wl[44] vdd gnd cell_6t
Xbit_r45_c37 bl[37] br[37] wl[45] vdd gnd cell_6t
Xbit_r46_c37 bl[37] br[37] wl[46] vdd gnd cell_6t
Xbit_r47_c37 bl[37] br[37] wl[47] vdd gnd cell_6t
Xbit_r48_c37 bl[37] br[37] wl[48] vdd gnd cell_6t
Xbit_r49_c37 bl[37] br[37] wl[49] vdd gnd cell_6t
Xbit_r50_c37 bl[37] br[37] wl[50] vdd gnd cell_6t
Xbit_r51_c37 bl[37] br[37] wl[51] vdd gnd cell_6t
Xbit_r52_c37 bl[37] br[37] wl[52] vdd gnd cell_6t
Xbit_r53_c37 bl[37] br[37] wl[53] vdd gnd cell_6t
Xbit_r54_c37 bl[37] br[37] wl[54] vdd gnd cell_6t
Xbit_r55_c37 bl[37] br[37] wl[55] vdd gnd cell_6t
Xbit_r56_c37 bl[37] br[37] wl[56] vdd gnd cell_6t
Xbit_r57_c37 bl[37] br[37] wl[57] vdd gnd cell_6t
Xbit_r58_c37 bl[37] br[37] wl[58] vdd gnd cell_6t
Xbit_r59_c37 bl[37] br[37] wl[59] vdd gnd cell_6t
Xbit_r60_c37 bl[37] br[37] wl[60] vdd gnd cell_6t
Xbit_r61_c37 bl[37] br[37] wl[61] vdd gnd cell_6t
Xbit_r62_c37 bl[37] br[37] wl[62] vdd gnd cell_6t
Xbit_r63_c37 bl[37] br[37] wl[63] vdd gnd cell_6t
Xbit_r64_c37 bl[37] br[37] wl[64] vdd gnd cell_6t
Xbit_r65_c37 bl[37] br[37] wl[65] vdd gnd cell_6t
Xbit_r66_c37 bl[37] br[37] wl[66] vdd gnd cell_6t
Xbit_r67_c37 bl[37] br[37] wl[67] vdd gnd cell_6t
Xbit_r68_c37 bl[37] br[37] wl[68] vdd gnd cell_6t
Xbit_r69_c37 bl[37] br[37] wl[69] vdd gnd cell_6t
Xbit_r70_c37 bl[37] br[37] wl[70] vdd gnd cell_6t
Xbit_r71_c37 bl[37] br[37] wl[71] vdd gnd cell_6t
Xbit_r72_c37 bl[37] br[37] wl[72] vdd gnd cell_6t
Xbit_r73_c37 bl[37] br[37] wl[73] vdd gnd cell_6t
Xbit_r74_c37 bl[37] br[37] wl[74] vdd gnd cell_6t
Xbit_r75_c37 bl[37] br[37] wl[75] vdd gnd cell_6t
Xbit_r76_c37 bl[37] br[37] wl[76] vdd gnd cell_6t
Xbit_r77_c37 bl[37] br[37] wl[77] vdd gnd cell_6t
Xbit_r78_c37 bl[37] br[37] wl[78] vdd gnd cell_6t
Xbit_r79_c37 bl[37] br[37] wl[79] vdd gnd cell_6t
Xbit_r80_c37 bl[37] br[37] wl[80] vdd gnd cell_6t
Xbit_r81_c37 bl[37] br[37] wl[81] vdd gnd cell_6t
Xbit_r82_c37 bl[37] br[37] wl[82] vdd gnd cell_6t
Xbit_r83_c37 bl[37] br[37] wl[83] vdd gnd cell_6t
Xbit_r84_c37 bl[37] br[37] wl[84] vdd gnd cell_6t
Xbit_r85_c37 bl[37] br[37] wl[85] vdd gnd cell_6t
Xbit_r86_c37 bl[37] br[37] wl[86] vdd gnd cell_6t
Xbit_r87_c37 bl[37] br[37] wl[87] vdd gnd cell_6t
Xbit_r88_c37 bl[37] br[37] wl[88] vdd gnd cell_6t
Xbit_r89_c37 bl[37] br[37] wl[89] vdd gnd cell_6t
Xbit_r90_c37 bl[37] br[37] wl[90] vdd gnd cell_6t
Xbit_r91_c37 bl[37] br[37] wl[91] vdd gnd cell_6t
Xbit_r92_c37 bl[37] br[37] wl[92] vdd gnd cell_6t
Xbit_r93_c37 bl[37] br[37] wl[93] vdd gnd cell_6t
Xbit_r94_c37 bl[37] br[37] wl[94] vdd gnd cell_6t
Xbit_r95_c37 bl[37] br[37] wl[95] vdd gnd cell_6t
Xbit_r96_c37 bl[37] br[37] wl[96] vdd gnd cell_6t
Xbit_r97_c37 bl[37] br[37] wl[97] vdd gnd cell_6t
Xbit_r98_c37 bl[37] br[37] wl[98] vdd gnd cell_6t
Xbit_r99_c37 bl[37] br[37] wl[99] vdd gnd cell_6t
Xbit_r100_c37 bl[37] br[37] wl[100] vdd gnd cell_6t
Xbit_r101_c37 bl[37] br[37] wl[101] vdd gnd cell_6t
Xbit_r102_c37 bl[37] br[37] wl[102] vdd gnd cell_6t
Xbit_r103_c37 bl[37] br[37] wl[103] vdd gnd cell_6t
Xbit_r104_c37 bl[37] br[37] wl[104] vdd gnd cell_6t
Xbit_r105_c37 bl[37] br[37] wl[105] vdd gnd cell_6t
Xbit_r106_c37 bl[37] br[37] wl[106] vdd gnd cell_6t
Xbit_r107_c37 bl[37] br[37] wl[107] vdd gnd cell_6t
Xbit_r108_c37 bl[37] br[37] wl[108] vdd gnd cell_6t
Xbit_r109_c37 bl[37] br[37] wl[109] vdd gnd cell_6t
Xbit_r110_c37 bl[37] br[37] wl[110] vdd gnd cell_6t
Xbit_r111_c37 bl[37] br[37] wl[111] vdd gnd cell_6t
Xbit_r112_c37 bl[37] br[37] wl[112] vdd gnd cell_6t
Xbit_r113_c37 bl[37] br[37] wl[113] vdd gnd cell_6t
Xbit_r114_c37 bl[37] br[37] wl[114] vdd gnd cell_6t
Xbit_r115_c37 bl[37] br[37] wl[115] vdd gnd cell_6t
Xbit_r116_c37 bl[37] br[37] wl[116] vdd gnd cell_6t
Xbit_r117_c37 bl[37] br[37] wl[117] vdd gnd cell_6t
Xbit_r118_c37 bl[37] br[37] wl[118] vdd gnd cell_6t
Xbit_r119_c37 bl[37] br[37] wl[119] vdd gnd cell_6t
Xbit_r120_c37 bl[37] br[37] wl[120] vdd gnd cell_6t
Xbit_r121_c37 bl[37] br[37] wl[121] vdd gnd cell_6t
Xbit_r122_c37 bl[37] br[37] wl[122] vdd gnd cell_6t
Xbit_r123_c37 bl[37] br[37] wl[123] vdd gnd cell_6t
Xbit_r124_c37 bl[37] br[37] wl[124] vdd gnd cell_6t
Xbit_r125_c37 bl[37] br[37] wl[125] vdd gnd cell_6t
Xbit_r126_c37 bl[37] br[37] wl[126] vdd gnd cell_6t
Xbit_r127_c37 bl[37] br[37] wl[127] vdd gnd cell_6t
Xbit_r0_c38 bl[38] br[38] wl[0] vdd gnd cell_6t
Xbit_r1_c38 bl[38] br[38] wl[1] vdd gnd cell_6t
Xbit_r2_c38 bl[38] br[38] wl[2] vdd gnd cell_6t
Xbit_r3_c38 bl[38] br[38] wl[3] vdd gnd cell_6t
Xbit_r4_c38 bl[38] br[38] wl[4] vdd gnd cell_6t
Xbit_r5_c38 bl[38] br[38] wl[5] vdd gnd cell_6t
Xbit_r6_c38 bl[38] br[38] wl[6] vdd gnd cell_6t
Xbit_r7_c38 bl[38] br[38] wl[7] vdd gnd cell_6t
Xbit_r8_c38 bl[38] br[38] wl[8] vdd gnd cell_6t
Xbit_r9_c38 bl[38] br[38] wl[9] vdd gnd cell_6t
Xbit_r10_c38 bl[38] br[38] wl[10] vdd gnd cell_6t
Xbit_r11_c38 bl[38] br[38] wl[11] vdd gnd cell_6t
Xbit_r12_c38 bl[38] br[38] wl[12] vdd gnd cell_6t
Xbit_r13_c38 bl[38] br[38] wl[13] vdd gnd cell_6t
Xbit_r14_c38 bl[38] br[38] wl[14] vdd gnd cell_6t
Xbit_r15_c38 bl[38] br[38] wl[15] vdd gnd cell_6t
Xbit_r16_c38 bl[38] br[38] wl[16] vdd gnd cell_6t
Xbit_r17_c38 bl[38] br[38] wl[17] vdd gnd cell_6t
Xbit_r18_c38 bl[38] br[38] wl[18] vdd gnd cell_6t
Xbit_r19_c38 bl[38] br[38] wl[19] vdd gnd cell_6t
Xbit_r20_c38 bl[38] br[38] wl[20] vdd gnd cell_6t
Xbit_r21_c38 bl[38] br[38] wl[21] vdd gnd cell_6t
Xbit_r22_c38 bl[38] br[38] wl[22] vdd gnd cell_6t
Xbit_r23_c38 bl[38] br[38] wl[23] vdd gnd cell_6t
Xbit_r24_c38 bl[38] br[38] wl[24] vdd gnd cell_6t
Xbit_r25_c38 bl[38] br[38] wl[25] vdd gnd cell_6t
Xbit_r26_c38 bl[38] br[38] wl[26] vdd gnd cell_6t
Xbit_r27_c38 bl[38] br[38] wl[27] vdd gnd cell_6t
Xbit_r28_c38 bl[38] br[38] wl[28] vdd gnd cell_6t
Xbit_r29_c38 bl[38] br[38] wl[29] vdd gnd cell_6t
Xbit_r30_c38 bl[38] br[38] wl[30] vdd gnd cell_6t
Xbit_r31_c38 bl[38] br[38] wl[31] vdd gnd cell_6t
Xbit_r32_c38 bl[38] br[38] wl[32] vdd gnd cell_6t
Xbit_r33_c38 bl[38] br[38] wl[33] vdd gnd cell_6t
Xbit_r34_c38 bl[38] br[38] wl[34] vdd gnd cell_6t
Xbit_r35_c38 bl[38] br[38] wl[35] vdd gnd cell_6t
Xbit_r36_c38 bl[38] br[38] wl[36] vdd gnd cell_6t
Xbit_r37_c38 bl[38] br[38] wl[37] vdd gnd cell_6t
Xbit_r38_c38 bl[38] br[38] wl[38] vdd gnd cell_6t
Xbit_r39_c38 bl[38] br[38] wl[39] vdd gnd cell_6t
Xbit_r40_c38 bl[38] br[38] wl[40] vdd gnd cell_6t
Xbit_r41_c38 bl[38] br[38] wl[41] vdd gnd cell_6t
Xbit_r42_c38 bl[38] br[38] wl[42] vdd gnd cell_6t
Xbit_r43_c38 bl[38] br[38] wl[43] vdd gnd cell_6t
Xbit_r44_c38 bl[38] br[38] wl[44] vdd gnd cell_6t
Xbit_r45_c38 bl[38] br[38] wl[45] vdd gnd cell_6t
Xbit_r46_c38 bl[38] br[38] wl[46] vdd gnd cell_6t
Xbit_r47_c38 bl[38] br[38] wl[47] vdd gnd cell_6t
Xbit_r48_c38 bl[38] br[38] wl[48] vdd gnd cell_6t
Xbit_r49_c38 bl[38] br[38] wl[49] vdd gnd cell_6t
Xbit_r50_c38 bl[38] br[38] wl[50] vdd gnd cell_6t
Xbit_r51_c38 bl[38] br[38] wl[51] vdd gnd cell_6t
Xbit_r52_c38 bl[38] br[38] wl[52] vdd gnd cell_6t
Xbit_r53_c38 bl[38] br[38] wl[53] vdd gnd cell_6t
Xbit_r54_c38 bl[38] br[38] wl[54] vdd gnd cell_6t
Xbit_r55_c38 bl[38] br[38] wl[55] vdd gnd cell_6t
Xbit_r56_c38 bl[38] br[38] wl[56] vdd gnd cell_6t
Xbit_r57_c38 bl[38] br[38] wl[57] vdd gnd cell_6t
Xbit_r58_c38 bl[38] br[38] wl[58] vdd gnd cell_6t
Xbit_r59_c38 bl[38] br[38] wl[59] vdd gnd cell_6t
Xbit_r60_c38 bl[38] br[38] wl[60] vdd gnd cell_6t
Xbit_r61_c38 bl[38] br[38] wl[61] vdd gnd cell_6t
Xbit_r62_c38 bl[38] br[38] wl[62] vdd gnd cell_6t
Xbit_r63_c38 bl[38] br[38] wl[63] vdd gnd cell_6t
Xbit_r64_c38 bl[38] br[38] wl[64] vdd gnd cell_6t
Xbit_r65_c38 bl[38] br[38] wl[65] vdd gnd cell_6t
Xbit_r66_c38 bl[38] br[38] wl[66] vdd gnd cell_6t
Xbit_r67_c38 bl[38] br[38] wl[67] vdd gnd cell_6t
Xbit_r68_c38 bl[38] br[38] wl[68] vdd gnd cell_6t
Xbit_r69_c38 bl[38] br[38] wl[69] vdd gnd cell_6t
Xbit_r70_c38 bl[38] br[38] wl[70] vdd gnd cell_6t
Xbit_r71_c38 bl[38] br[38] wl[71] vdd gnd cell_6t
Xbit_r72_c38 bl[38] br[38] wl[72] vdd gnd cell_6t
Xbit_r73_c38 bl[38] br[38] wl[73] vdd gnd cell_6t
Xbit_r74_c38 bl[38] br[38] wl[74] vdd gnd cell_6t
Xbit_r75_c38 bl[38] br[38] wl[75] vdd gnd cell_6t
Xbit_r76_c38 bl[38] br[38] wl[76] vdd gnd cell_6t
Xbit_r77_c38 bl[38] br[38] wl[77] vdd gnd cell_6t
Xbit_r78_c38 bl[38] br[38] wl[78] vdd gnd cell_6t
Xbit_r79_c38 bl[38] br[38] wl[79] vdd gnd cell_6t
Xbit_r80_c38 bl[38] br[38] wl[80] vdd gnd cell_6t
Xbit_r81_c38 bl[38] br[38] wl[81] vdd gnd cell_6t
Xbit_r82_c38 bl[38] br[38] wl[82] vdd gnd cell_6t
Xbit_r83_c38 bl[38] br[38] wl[83] vdd gnd cell_6t
Xbit_r84_c38 bl[38] br[38] wl[84] vdd gnd cell_6t
Xbit_r85_c38 bl[38] br[38] wl[85] vdd gnd cell_6t
Xbit_r86_c38 bl[38] br[38] wl[86] vdd gnd cell_6t
Xbit_r87_c38 bl[38] br[38] wl[87] vdd gnd cell_6t
Xbit_r88_c38 bl[38] br[38] wl[88] vdd gnd cell_6t
Xbit_r89_c38 bl[38] br[38] wl[89] vdd gnd cell_6t
Xbit_r90_c38 bl[38] br[38] wl[90] vdd gnd cell_6t
Xbit_r91_c38 bl[38] br[38] wl[91] vdd gnd cell_6t
Xbit_r92_c38 bl[38] br[38] wl[92] vdd gnd cell_6t
Xbit_r93_c38 bl[38] br[38] wl[93] vdd gnd cell_6t
Xbit_r94_c38 bl[38] br[38] wl[94] vdd gnd cell_6t
Xbit_r95_c38 bl[38] br[38] wl[95] vdd gnd cell_6t
Xbit_r96_c38 bl[38] br[38] wl[96] vdd gnd cell_6t
Xbit_r97_c38 bl[38] br[38] wl[97] vdd gnd cell_6t
Xbit_r98_c38 bl[38] br[38] wl[98] vdd gnd cell_6t
Xbit_r99_c38 bl[38] br[38] wl[99] vdd gnd cell_6t
Xbit_r100_c38 bl[38] br[38] wl[100] vdd gnd cell_6t
Xbit_r101_c38 bl[38] br[38] wl[101] vdd gnd cell_6t
Xbit_r102_c38 bl[38] br[38] wl[102] vdd gnd cell_6t
Xbit_r103_c38 bl[38] br[38] wl[103] vdd gnd cell_6t
Xbit_r104_c38 bl[38] br[38] wl[104] vdd gnd cell_6t
Xbit_r105_c38 bl[38] br[38] wl[105] vdd gnd cell_6t
Xbit_r106_c38 bl[38] br[38] wl[106] vdd gnd cell_6t
Xbit_r107_c38 bl[38] br[38] wl[107] vdd gnd cell_6t
Xbit_r108_c38 bl[38] br[38] wl[108] vdd gnd cell_6t
Xbit_r109_c38 bl[38] br[38] wl[109] vdd gnd cell_6t
Xbit_r110_c38 bl[38] br[38] wl[110] vdd gnd cell_6t
Xbit_r111_c38 bl[38] br[38] wl[111] vdd gnd cell_6t
Xbit_r112_c38 bl[38] br[38] wl[112] vdd gnd cell_6t
Xbit_r113_c38 bl[38] br[38] wl[113] vdd gnd cell_6t
Xbit_r114_c38 bl[38] br[38] wl[114] vdd gnd cell_6t
Xbit_r115_c38 bl[38] br[38] wl[115] vdd gnd cell_6t
Xbit_r116_c38 bl[38] br[38] wl[116] vdd gnd cell_6t
Xbit_r117_c38 bl[38] br[38] wl[117] vdd gnd cell_6t
Xbit_r118_c38 bl[38] br[38] wl[118] vdd gnd cell_6t
Xbit_r119_c38 bl[38] br[38] wl[119] vdd gnd cell_6t
Xbit_r120_c38 bl[38] br[38] wl[120] vdd gnd cell_6t
Xbit_r121_c38 bl[38] br[38] wl[121] vdd gnd cell_6t
Xbit_r122_c38 bl[38] br[38] wl[122] vdd gnd cell_6t
Xbit_r123_c38 bl[38] br[38] wl[123] vdd gnd cell_6t
Xbit_r124_c38 bl[38] br[38] wl[124] vdd gnd cell_6t
Xbit_r125_c38 bl[38] br[38] wl[125] vdd gnd cell_6t
Xbit_r126_c38 bl[38] br[38] wl[126] vdd gnd cell_6t
Xbit_r127_c38 bl[38] br[38] wl[127] vdd gnd cell_6t
Xbit_r0_c39 bl[39] br[39] wl[0] vdd gnd cell_6t
Xbit_r1_c39 bl[39] br[39] wl[1] vdd gnd cell_6t
Xbit_r2_c39 bl[39] br[39] wl[2] vdd gnd cell_6t
Xbit_r3_c39 bl[39] br[39] wl[3] vdd gnd cell_6t
Xbit_r4_c39 bl[39] br[39] wl[4] vdd gnd cell_6t
Xbit_r5_c39 bl[39] br[39] wl[5] vdd gnd cell_6t
Xbit_r6_c39 bl[39] br[39] wl[6] vdd gnd cell_6t
Xbit_r7_c39 bl[39] br[39] wl[7] vdd gnd cell_6t
Xbit_r8_c39 bl[39] br[39] wl[8] vdd gnd cell_6t
Xbit_r9_c39 bl[39] br[39] wl[9] vdd gnd cell_6t
Xbit_r10_c39 bl[39] br[39] wl[10] vdd gnd cell_6t
Xbit_r11_c39 bl[39] br[39] wl[11] vdd gnd cell_6t
Xbit_r12_c39 bl[39] br[39] wl[12] vdd gnd cell_6t
Xbit_r13_c39 bl[39] br[39] wl[13] vdd gnd cell_6t
Xbit_r14_c39 bl[39] br[39] wl[14] vdd gnd cell_6t
Xbit_r15_c39 bl[39] br[39] wl[15] vdd gnd cell_6t
Xbit_r16_c39 bl[39] br[39] wl[16] vdd gnd cell_6t
Xbit_r17_c39 bl[39] br[39] wl[17] vdd gnd cell_6t
Xbit_r18_c39 bl[39] br[39] wl[18] vdd gnd cell_6t
Xbit_r19_c39 bl[39] br[39] wl[19] vdd gnd cell_6t
Xbit_r20_c39 bl[39] br[39] wl[20] vdd gnd cell_6t
Xbit_r21_c39 bl[39] br[39] wl[21] vdd gnd cell_6t
Xbit_r22_c39 bl[39] br[39] wl[22] vdd gnd cell_6t
Xbit_r23_c39 bl[39] br[39] wl[23] vdd gnd cell_6t
Xbit_r24_c39 bl[39] br[39] wl[24] vdd gnd cell_6t
Xbit_r25_c39 bl[39] br[39] wl[25] vdd gnd cell_6t
Xbit_r26_c39 bl[39] br[39] wl[26] vdd gnd cell_6t
Xbit_r27_c39 bl[39] br[39] wl[27] vdd gnd cell_6t
Xbit_r28_c39 bl[39] br[39] wl[28] vdd gnd cell_6t
Xbit_r29_c39 bl[39] br[39] wl[29] vdd gnd cell_6t
Xbit_r30_c39 bl[39] br[39] wl[30] vdd gnd cell_6t
Xbit_r31_c39 bl[39] br[39] wl[31] vdd gnd cell_6t
Xbit_r32_c39 bl[39] br[39] wl[32] vdd gnd cell_6t
Xbit_r33_c39 bl[39] br[39] wl[33] vdd gnd cell_6t
Xbit_r34_c39 bl[39] br[39] wl[34] vdd gnd cell_6t
Xbit_r35_c39 bl[39] br[39] wl[35] vdd gnd cell_6t
Xbit_r36_c39 bl[39] br[39] wl[36] vdd gnd cell_6t
Xbit_r37_c39 bl[39] br[39] wl[37] vdd gnd cell_6t
Xbit_r38_c39 bl[39] br[39] wl[38] vdd gnd cell_6t
Xbit_r39_c39 bl[39] br[39] wl[39] vdd gnd cell_6t
Xbit_r40_c39 bl[39] br[39] wl[40] vdd gnd cell_6t
Xbit_r41_c39 bl[39] br[39] wl[41] vdd gnd cell_6t
Xbit_r42_c39 bl[39] br[39] wl[42] vdd gnd cell_6t
Xbit_r43_c39 bl[39] br[39] wl[43] vdd gnd cell_6t
Xbit_r44_c39 bl[39] br[39] wl[44] vdd gnd cell_6t
Xbit_r45_c39 bl[39] br[39] wl[45] vdd gnd cell_6t
Xbit_r46_c39 bl[39] br[39] wl[46] vdd gnd cell_6t
Xbit_r47_c39 bl[39] br[39] wl[47] vdd gnd cell_6t
Xbit_r48_c39 bl[39] br[39] wl[48] vdd gnd cell_6t
Xbit_r49_c39 bl[39] br[39] wl[49] vdd gnd cell_6t
Xbit_r50_c39 bl[39] br[39] wl[50] vdd gnd cell_6t
Xbit_r51_c39 bl[39] br[39] wl[51] vdd gnd cell_6t
Xbit_r52_c39 bl[39] br[39] wl[52] vdd gnd cell_6t
Xbit_r53_c39 bl[39] br[39] wl[53] vdd gnd cell_6t
Xbit_r54_c39 bl[39] br[39] wl[54] vdd gnd cell_6t
Xbit_r55_c39 bl[39] br[39] wl[55] vdd gnd cell_6t
Xbit_r56_c39 bl[39] br[39] wl[56] vdd gnd cell_6t
Xbit_r57_c39 bl[39] br[39] wl[57] vdd gnd cell_6t
Xbit_r58_c39 bl[39] br[39] wl[58] vdd gnd cell_6t
Xbit_r59_c39 bl[39] br[39] wl[59] vdd gnd cell_6t
Xbit_r60_c39 bl[39] br[39] wl[60] vdd gnd cell_6t
Xbit_r61_c39 bl[39] br[39] wl[61] vdd gnd cell_6t
Xbit_r62_c39 bl[39] br[39] wl[62] vdd gnd cell_6t
Xbit_r63_c39 bl[39] br[39] wl[63] vdd gnd cell_6t
Xbit_r64_c39 bl[39] br[39] wl[64] vdd gnd cell_6t
Xbit_r65_c39 bl[39] br[39] wl[65] vdd gnd cell_6t
Xbit_r66_c39 bl[39] br[39] wl[66] vdd gnd cell_6t
Xbit_r67_c39 bl[39] br[39] wl[67] vdd gnd cell_6t
Xbit_r68_c39 bl[39] br[39] wl[68] vdd gnd cell_6t
Xbit_r69_c39 bl[39] br[39] wl[69] vdd gnd cell_6t
Xbit_r70_c39 bl[39] br[39] wl[70] vdd gnd cell_6t
Xbit_r71_c39 bl[39] br[39] wl[71] vdd gnd cell_6t
Xbit_r72_c39 bl[39] br[39] wl[72] vdd gnd cell_6t
Xbit_r73_c39 bl[39] br[39] wl[73] vdd gnd cell_6t
Xbit_r74_c39 bl[39] br[39] wl[74] vdd gnd cell_6t
Xbit_r75_c39 bl[39] br[39] wl[75] vdd gnd cell_6t
Xbit_r76_c39 bl[39] br[39] wl[76] vdd gnd cell_6t
Xbit_r77_c39 bl[39] br[39] wl[77] vdd gnd cell_6t
Xbit_r78_c39 bl[39] br[39] wl[78] vdd gnd cell_6t
Xbit_r79_c39 bl[39] br[39] wl[79] vdd gnd cell_6t
Xbit_r80_c39 bl[39] br[39] wl[80] vdd gnd cell_6t
Xbit_r81_c39 bl[39] br[39] wl[81] vdd gnd cell_6t
Xbit_r82_c39 bl[39] br[39] wl[82] vdd gnd cell_6t
Xbit_r83_c39 bl[39] br[39] wl[83] vdd gnd cell_6t
Xbit_r84_c39 bl[39] br[39] wl[84] vdd gnd cell_6t
Xbit_r85_c39 bl[39] br[39] wl[85] vdd gnd cell_6t
Xbit_r86_c39 bl[39] br[39] wl[86] vdd gnd cell_6t
Xbit_r87_c39 bl[39] br[39] wl[87] vdd gnd cell_6t
Xbit_r88_c39 bl[39] br[39] wl[88] vdd gnd cell_6t
Xbit_r89_c39 bl[39] br[39] wl[89] vdd gnd cell_6t
Xbit_r90_c39 bl[39] br[39] wl[90] vdd gnd cell_6t
Xbit_r91_c39 bl[39] br[39] wl[91] vdd gnd cell_6t
Xbit_r92_c39 bl[39] br[39] wl[92] vdd gnd cell_6t
Xbit_r93_c39 bl[39] br[39] wl[93] vdd gnd cell_6t
Xbit_r94_c39 bl[39] br[39] wl[94] vdd gnd cell_6t
Xbit_r95_c39 bl[39] br[39] wl[95] vdd gnd cell_6t
Xbit_r96_c39 bl[39] br[39] wl[96] vdd gnd cell_6t
Xbit_r97_c39 bl[39] br[39] wl[97] vdd gnd cell_6t
Xbit_r98_c39 bl[39] br[39] wl[98] vdd gnd cell_6t
Xbit_r99_c39 bl[39] br[39] wl[99] vdd gnd cell_6t
Xbit_r100_c39 bl[39] br[39] wl[100] vdd gnd cell_6t
Xbit_r101_c39 bl[39] br[39] wl[101] vdd gnd cell_6t
Xbit_r102_c39 bl[39] br[39] wl[102] vdd gnd cell_6t
Xbit_r103_c39 bl[39] br[39] wl[103] vdd gnd cell_6t
Xbit_r104_c39 bl[39] br[39] wl[104] vdd gnd cell_6t
Xbit_r105_c39 bl[39] br[39] wl[105] vdd gnd cell_6t
Xbit_r106_c39 bl[39] br[39] wl[106] vdd gnd cell_6t
Xbit_r107_c39 bl[39] br[39] wl[107] vdd gnd cell_6t
Xbit_r108_c39 bl[39] br[39] wl[108] vdd gnd cell_6t
Xbit_r109_c39 bl[39] br[39] wl[109] vdd gnd cell_6t
Xbit_r110_c39 bl[39] br[39] wl[110] vdd gnd cell_6t
Xbit_r111_c39 bl[39] br[39] wl[111] vdd gnd cell_6t
Xbit_r112_c39 bl[39] br[39] wl[112] vdd gnd cell_6t
Xbit_r113_c39 bl[39] br[39] wl[113] vdd gnd cell_6t
Xbit_r114_c39 bl[39] br[39] wl[114] vdd gnd cell_6t
Xbit_r115_c39 bl[39] br[39] wl[115] vdd gnd cell_6t
Xbit_r116_c39 bl[39] br[39] wl[116] vdd gnd cell_6t
Xbit_r117_c39 bl[39] br[39] wl[117] vdd gnd cell_6t
Xbit_r118_c39 bl[39] br[39] wl[118] vdd gnd cell_6t
Xbit_r119_c39 bl[39] br[39] wl[119] vdd gnd cell_6t
Xbit_r120_c39 bl[39] br[39] wl[120] vdd gnd cell_6t
Xbit_r121_c39 bl[39] br[39] wl[121] vdd gnd cell_6t
Xbit_r122_c39 bl[39] br[39] wl[122] vdd gnd cell_6t
Xbit_r123_c39 bl[39] br[39] wl[123] vdd gnd cell_6t
Xbit_r124_c39 bl[39] br[39] wl[124] vdd gnd cell_6t
Xbit_r125_c39 bl[39] br[39] wl[125] vdd gnd cell_6t
Xbit_r126_c39 bl[39] br[39] wl[126] vdd gnd cell_6t
Xbit_r127_c39 bl[39] br[39] wl[127] vdd gnd cell_6t
Xbit_r0_c40 bl[40] br[40] wl[0] vdd gnd cell_6t
Xbit_r1_c40 bl[40] br[40] wl[1] vdd gnd cell_6t
Xbit_r2_c40 bl[40] br[40] wl[2] vdd gnd cell_6t
Xbit_r3_c40 bl[40] br[40] wl[3] vdd gnd cell_6t
Xbit_r4_c40 bl[40] br[40] wl[4] vdd gnd cell_6t
Xbit_r5_c40 bl[40] br[40] wl[5] vdd gnd cell_6t
Xbit_r6_c40 bl[40] br[40] wl[6] vdd gnd cell_6t
Xbit_r7_c40 bl[40] br[40] wl[7] vdd gnd cell_6t
Xbit_r8_c40 bl[40] br[40] wl[8] vdd gnd cell_6t
Xbit_r9_c40 bl[40] br[40] wl[9] vdd gnd cell_6t
Xbit_r10_c40 bl[40] br[40] wl[10] vdd gnd cell_6t
Xbit_r11_c40 bl[40] br[40] wl[11] vdd gnd cell_6t
Xbit_r12_c40 bl[40] br[40] wl[12] vdd gnd cell_6t
Xbit_r13_c40 bl[40] br[40] wl[13] vdd gnd cell_6t
Xbit_r14_c40 bl[40] br[40] wl[14] vdd gnd cell_6t
Xbit_r15_c40 bl[40] br[40] wl[15] vdd gnd cell_6t
Xbit_r16_c40 bl[40] br[40] wl[16] vdd gnd cell_6t
Xbit_r17_c40 bl[40] br[40] wl[17] vdd gnd cell_6t
Xbit_r18_c40 bl[40] br[40] wl[18] vdd gnd cell_6t
Xbit_r19_c40 bl[40] br[40] wl[19] vdd gnd cell_6t
Xbit_r20_c40 bl[40] br[40] wl[20] vdd gnd cell_6t
Xbit_r21_c40 bl[40] br[40] wl[21] vdd gnd cell_6t
Xbit_r22_c40 bl[40] br[40] wl[22] vdd gnd cell_6t
Xbit_r23_c40 bl[40] br[40] wl[23] vdd gnd cell_6t
Xbit_r24_c40 bl[40] br[40] wl[24] vdd gnd cell_6t
Xbit_r25_c40 bl[40] br[40] wl[25] vdd gnd cell_6t
Xbit_r26_c40 bl[40] br[40] wl[26] vdd gnd cell_6t
Xbit_r27_c40 bl[40] br[40] wl[27] vdd gnd cell_6t
Xbit_r28_c40 bl[40] br[40] wl[28] vdd gnd cell_6t
Xbit_r29_c40 bl[40] br[40] wl[29] vdd gnd cell_6t
Xbit_r30_c40 bl[40] br[40] wl[30] vdd gnd cell_6t
Xbit_r31_c40 bl[40] br[40] wl[31] vdd gnd cell_6t
Xbit_r32_c40 bl[40] br[40] wl[32] vdd gnd cell_6t
Xbit_r33_c40 bl[40] br[40] wl[33] vdd gnd cell_6t
Xbit_r34_c40 bl[40] br[40] wl[34] vdd gnd cell_6t
Xbit_r35_c40 bl[40] br[40] wl[35] vdd gnd cell_6t
Xbit_r36_c40 bl[40] br[40] wl[36] vdd gnd cell_6t
Xbit_r37_c40 bl[40] br[40] wl[37] vdd gnd cell_6t
Xbit_r38_c40 bl[40] br[40] wl[38] vdd gnd cell_6t
Xbit_r39_c40 bl[40] br[40] wl[39] vdd gnd cell_6t
Xbit_r40_c40 bl[40] br[40] wl[40] vdd gnd cell_6t
Xbit_r41_c40 bl[40] br[40] wl[41] vdd gnd cell_6t
Xbit_r42_c40 bl[40] br[40] wl[42] vdd gnd cell_6t
Xbit_r43_c40 bl[40] br[40] wl[43] vdd gnd cell_6t
Xbit_r44_c40 bl[40] br[40] wl[44] vdd gnd cell_6t
Xbit_r45_c40 bl[40] br[40] wl[45] vdd gnd cell_6t
Xbit_r46_c40 bl[40] br[40] wl[46] vdd gnd cell_6t
Xbit_r47_c40 bl[40] br[40] wl[47] vdd gnd cell_6t
Xbit_r48_c40 bl[40] br[40] wl[48] vdd gnd cell_6t
Xbit_r49_c40 bl[40] br[40] wl[49] vdd gnd cell_6t
Xbit_r50_c40 bl[40] br[40] wl[50] vdd gnd cell_6t
Xbit_r51_c40 bl[40] br[40] wl[51] vdd gnd cell_6t
Xbit_r52_c40 bl[40] br[40] wl[52] vdd gnd cell_6t
Xbit_r53_c40 bl[40] br[40] wl[53] vdd gnd cell_6t
Xbit_r54_c40 bl[40] br[40] wl[54] vdd gnd cell_6t
Xbit_r55_c40 bl[40] br[40] wl[55] vdd gnd cell_6t
Xbit_r56_c40 bl[40] br[40] wl[56] vdd gnd cell_6t
Xbit_r57_c40 bl[40] br[40] wl[57] vdd gnd cell_6t
Xbit_r58_c40 bl[40] br[40] wl[58] vdd gnd cell_6t
Xbit_r59_c40 bl[40] br[40] wl[59] vdd gnd cell_6t
Xbit_r60_c40 bl[40] br[40] wl[60] vdd gnd cell_6t
Xbit_r61_c40 bl[40] br[40] wl[61] vdd gnd cell_6t
Xbit_r62_c40 bl[40] br[40] wl[62] vdd gnd cell_6t
Xbit_r63_c40 bl[40] br[40] wl[63] vdd gnd cell_6t
Xbit_r64_c40 bl[40] br[40] wl[64] vdd gnd cell_6t
Xbit_r65_c40 bl[40] br[40] wl[65] vdd gnd cell_6t
Xbit_r66_c40 bl[40] br[40] wl[66] vdd gnd cell_6t
Xbit_r67_c40 bl[40] br[40] wl[67] vdd gnd cell_6t
Xbit_r68_c40 bl[40] br[40] wl[68] vdd gnd cell_6t
Xbit_r69_c40 bl[40] br[40] wl[69] vdd gnd cell_6t
Xbit_r70_c40 bl[40] br[40] wl[70] vdd gnd cell_6t
Xbit_r71_c40 bl[40] br[40] wl[71] vdd gnd cell_6t
Xbit_r72_c40 bl[40] br[40] wl[72] vdd gnd cell_6t
Xbit_r73_c40 bl[40] br[40] wl[73] vdd gnd cell_6t
Xbit_r74_c40 bl[40] br[40] wl[74] vdd gnd cell_6t
Xbit_r75_c40 bl[40] br[40] wl[75] vdd gnd cell_6t
Xbit_r76_c40 bl[40] br[40] wl[76] vdd gnd cell_6t
Xbit_r77_c40 bl[40] br[40] wl[77] vdd gnd cell_6t
Xbit_r78_c40 bl[40] br[40] wl[78] vdd gnd cell_6t
Xbit_r79_c40 bl[40] br[40] wl[79] vdd gnd cell_6t
Xbit_r80_c40 bl[40] br[40] wl[80] vdd gnd cell_6t
Xbit_r81_c40 bl[40] br[40] wl[81] vdd gnd cell_6t
Xbit_r82_c40 bl[40] br[40] wl[82] vdd gnd cell_6t
Xbit_r83_c40 bl[40] br[40] wl[83] vdd gnd cell_6t
Xbit_r84_c40 bl[40] br[40] wl[84] vdd gnd cell_6t
Xbit_r85_c40 bl[40] br[40] wl[85] vdd gnd cell_6t
Xbit_r86_c40 bl[40] br[40] wl[86] vdd gnd cell_6t
Xbit_r87_c40 bl[40] br[40] wl[87] vdd gnd cell_6t
Xbit_r88_c40 bl[40] br[40] wl[88] vdd gnd cell_6t
Xbit_r89_c40 bl[40] br[40] wl[89] vdd gnd cell_6t
Xbit_r90_c40 bl[40] br[40] wl[90] vdd gnd cell_6t
Xbit_r91_c40 bl[40] br[40] wl[91] vdd gnd cell_6t
Xbit_r92_c40 bl[40] br[40] wl[92] vdd gnd cell_6t
Xbit_r93_c40 bl[40] br[40] wl[93] vdd gnd cell_6t
Xbit_r94_c40 bl[40] br[40] wl[94] vdd gnd cell_6t
Xbit_r95_c40 bl[40] br[40] wl[95] vdd gnd cell_6t
Xbit_r96_c40 bl[40] br[40] wl[96] vdd gnd cell_6t
Xbit_r97_c40 bl[40] br[40] wl[97] vdd gnd cell_6t
Xbit_r98_c40 bl[40] br[40] wl[98] vdd gnd cell_6t
Xbit_r99_c40 bl[40] br[40] wl[99] vdd gnd cell_6t
Xbit_r100_c40 bl[40] br[40] wl[100] vdd gnd cell_6t
Xbit_r101_c40 bl[40] br[40] wl[101] vdd gnd cell_6t
Xbit_r102_c40 bl[40] br[40] wl[102] vdd gnd cell_6t
Xbit_r103_c40 bl[40] br[40] wl[103] vdd gnd cell_6t
Xbit_r104_c40 bl[40] br[40] wl[104] vdd gnd cell_6t
Xbit_r105_c40 bl[40] br[40] wl[105] vdd gnd cell_6t
Xbit_r106_c40 bl[40] br[40] wl[106] vdd gnd cell_6t
Xbit_r107_c40 bl[40] br[40] wl[107] vdd gnd cell_6t
Xbit_r108_c40 bl[40] br[40] wl[108] vdd gnd cell_6t
Xbit_r109_c40 bl[40] br[40] wl[109] vdd gnd cell_6t
Xbit_r110_c40 bl[40] br[40] wl[110] vdd gnd cell_6t
Xbit_r111_c40 bl[40] br[40] wl[111] vdd gnd cell_6t
Xbit_r112_c40 bl[40] br[40] wl[112] vdd gnd cell_6t
Xbit_r113_c40 bl[40] br[40] wl[113] vdd gnd cell_6t
Xbit_r114_c40 bl[40] br[40] wl[114] vdd gnd cell_6t
Xbit_r115_c40 bl[40] br[40] wl[115] vdd gnd cell_6t
Xbit_r116_c40 bl[40] br[40] wl[116] vdd gnd cell_6t
Xbit_r117_c40 bl[40] br[40] wl[117] vdd gnd cell_6t
Xbit_r118_c40 bl[40] br[40] wl[118] vdd gnd cell_6t
Xbit_r119_c40 bl[40] br[40] wl[119] vdd gnd cell_6t
Xbit_r120_c40 bl[40] br[40] wl[120] vdd gnd cell_6t
Xbit_r121_c40 bl[40] br[40] wl[121] vdd gnd cell_6t
Xbit_r122_c40 bl[40] br[40] wl[122] vdd gnd cell_6t
Xbit_r123_c40 bl[40] br[40] wl[123] vdd gnd cell_6t
Xbit_r124_c40 bl[40] br[40] wl[124] vdd gnd cell_6t
Xbit_r125_c40 bl[40] br[40] wl[125] vdd gnd cell_6t
Xbit_r126_c40 bl[40] br[40] wl[126] vdd gnd cell_6t
Xbit_r127_c40 bl[40] br[40] wl[127] vdd gnd cell_6t
Xbit_r0_c41 bl[41] br[41] wl[0] vdd gnd cell_6t
Xbit_r1_c41 bl[41] br[41] wl[1] vdd gnd cell_6t
Xbit_r2_c41 bl[41] br[41] wl[2] vdd gnd cell_6t
Xbit_r3_c41 bl[41] br[41] wl[3] vdd gnd cell_6t
Xbit_r4_c41 bl[41] br[41] wl[4] vdd gnd cell_6t
Xbit_r5_c41 bl[41] br[41] wl[5] vdd gnd cell_6t
Xbit_r6_c41 bl[41] br[41] wl[6] vdd gnd cell_6t
Xbit_r7_c41 bl[41] br[41] wl[7] vdd gnd cell_6t
Xbit_r8_c41 bl[41] br[41] wl[8] vdd gnd cell_6t
Xbit_r9_c41 bl[41] br[41] wl[9] vdd gnd cell_6t
Xbit_r10_c41 bl[41] br[41] wl[10] vdd gnd cell_6t
Xbit_r11_c41 bl[41] br[41] wl[11] vdd gnd cell_6t
Xbit_r12_c41 bl[41] br[41] wl[12] vdd gnd cell_6t
Xbit_r13_c41 bl[41] br[41] wl[13] vdd gnd cell_6t
Xbit_r14_c41 bl[41] br[41] wl[14] vdd gnd cell_6t
Xbit_r15_c41 bl[41] br[41] wl[15] vdd gnd cell_6t
Xbit_r16_c41 bl[41] br[41] wl[16] vdd gnd cell_6t
Xbit_r17_c41 bl[41] br[41] wl[17] vdd gnd cell_6t
Xbit_r18_c41 bl[41] br[41] wl[18] vdd gnd cell_6t
Xbit_r19_c41 bl[41] br[41] wl[19] vdd gnd cell_6t
Xbit_r20_c41 bl[41] br[41] wl[20] vdd gnd cell_6t
Xbit_r21_c41 bl[41] br[41] wl[21] vdd gnd cell_6t
Xbit_r22_c41 bl[41] br[41] wl[22] vdd gnd cell_6t
Xbit_r23_c41 bl[41] br[41] wl[23] vdd gnd cell_6t
Xbit_r24_c41 bl[41] br[41] wl[24] vdd gnd cell_6t
Xbit_r25_c41 bl[41] br[41] wl[25] vdd gnd cell_6t
Xbit_r26_c41 bl[41] br[41] wl[26] vdd gnd cell_6t
Xbit_r27_c41 bl[41] br[41] wl[27] vdd gnd cell_6t
Xbit_r28_c41 bl[41] br[41] wl[28] vdd gnd cell_6t
Xbit_r29_c41 bl[41] br[41] wl[29] vdd gnd cell_6t
Xbit_r30_c41 bl[41] br[41] wl[30] vdd gnd cell_6t
Xbit_r31_c41 bl[41] br[41] wl[31] vdd gnd cell_6t
Xbit_r32_c41 bl[41] br[41] wl[32] vdd gnd cell_6t
Xbit_r33_c41 bl[41] br[41] wl[33] vdd gnd cell_6t
Xbit_r34_c41 bl[41] br[41] wl[34] vdd gnd cell_6t
Xbit_r35_c41 bl[41] br[41] wl[35] vdd gnd cell_6t
Xbit_r36_c41 bl[41] br[41] wl[36] vdd gnd cell_6t
Xbit_r37_c41 bl[41] br[41] wl[37] vdd gnd cell_6t
Xbit_r38_c41 bl[41] br[41] wl[38] vdd gnd cell_6t
Xbit_r39_c41 bl[41] br[41] wl[39] vdd gnd cell_6t
Xbit_r40_c41 bl[41] br[41] wl[40] vdd gnd cell_6t
Xbit_r41_c41 bl[41] br[41] wl[41] vdd gnd cell_6t
Xbit_r42_c41 bl[41] br[41] wl[42] vdd gnd cell_6t
Xbit_r43_c41 bl[41] br[41] wl[43] vdd gnd cell_6t
Xbit_r44_c41 bl[41] br[41] wl[44] vdd gnd cell_6t
Xbit_r45_c41 bl[41] br[41] wl[45] vdd gnd cell_6t
Xbit_r46_c41 bl[41] br[41] wl[46] vdd gnd cell_6t
Xbit_r47_c41 bl[41] br[41] wl[47] vdd gnd cell_6t
Xbit_r48_c41 bl[41] br[41] wl[48] vdd gnd cell_6t
Xbit_r49_c41 bl[41] br[41] wl[49] vdd gnd cell_6t
Xbit_r50_c41 bl[41] br[41] wl[50] vdd gnd cell_6t
Xbit_r51_c41 bl[41] br[41] wl[51] vdd gnd cell_6t
Xbit_r52_c41 bl[41] br[41] wl[52] vdd gnd cell_6t
Xbit_r53_c41 bl[41] br[41] wl[53] vdd gnd cell_6t
Xbit_r54_c41 bl[41] br[41] wl[54] vdd gnd cell_6t
Xbit_r55_c41 bl[41] br[41] wl[55] vdd gnd cell_6t
Xbit_r56_c41 bl[41] br[41] wl[56] vdd gnd cell_6t
Xbit_r57_c41 bl[41] br[41] wl[57] vdd gnd cell_6t
Xbit_r58_c41 bl[41] br[41] wl[58] vdd gnd cell_6t
Xbit_r59_c41 bl[41] br[41] wl[59] vdd gnd cell_6t
Xbit_r60_c41 bl[41] br[41] wl[60] vdd gnd cell_6t
Xbit_r61_c41 bl[41] br[41] wl[61] vdd gnd cell_6t
Xbit_r62_c41 bl[41] br[41] wl[62] vdd gnd cell_6t
Xbit_r63_c41 bl[41] br[41] wl[63] vdd gnd cell_6t
Xbit_r64_c41 bl[41] br[41] wl[64] vdd gnd cell_6t
Xbit_r65_c41 bl[41] br[41] wl[65] vdd gnd cell_6t
Xbit_r66_c41 bl[41] br[41] wl[66] vdd gnd cell_6t
Xbit_r67_c41 bl[41] br[41] wl[67] vdd gnd cell_6t
Xbit_r68_c41 bl[41] br[41] wl[68] vdd gnd cell_6t
Xbit_r69_c41 bl[41] br[41] wl[69] vdd gnd cell_6t
Xbit_r70_c41 bl[41] br[41] wl[70] vdd gnd cell_6t
Xbit_r71_c41 bl[41] br[41] wl[71] vdd gnd cell_6t
Xbit_r72_c41 bl[41] br[41] wl[72] vdd gnd cell_6t
Xbit_r73_c41 bl[41] br[41] wl[73] vdd gnd cell_6t
Xbit_r74_c41 bl[41] br[41] wl[74] vdd gnd cell_6t
Xbit_r75_c41 bl[41] br[41] wl[75] vdd gnd cell_6t
Xbit_r76_c41 bl[41] br[41] wl[76] vdd gnd cell_6t
Xbit_r77_c41 bl[41] br[41] wl[77] vdd gnd cell_6t
Xbit_r78_c41 bl[41] br[41] wl[78] vdd gnd cell_6t
Xbit_r79_c41 bl[41] br[41] wl[79] vdd gnd cell_6t
Xbit_r80_c41 bl[41] br[41] wl[80] vdd gnd cell_6t
Xbit_r81_c41 bl[41] br[41] wl[81] vdd gnd cell_6t
Xbit_r82_c41 bl[41] br[41] wl[82] vdd gnd cell_6t
Xbit_r83_c41 bl[41] br[41] wl[83] vdd gnd cell_6t
Xbit_r84_c41 bl[41] br[41] wl[84] vdd gnd cell_6t
Xbit_r85_c41 bl[41] br[41] wl[85] vdd gnd cell_6t
Xbit_r86_c41 bl[41] br[41] wl[86] vdd gnd cell_6t
Xbit_r87_c41 bl[41] br[41] wl[87] vdd gnd cell_6t
Xbit_r88_c41 bl[41] br[41] wl[88] vdd gnd cell_6t
Xbit_r89_c41 bl[41] br[41] wl[89] vdd gnd cell_6t
Xbit_r90_c41 bl[41] br[41] wl[90] vdd gnd cell_6t
Xbit_r91_c41 bl[41] br[41] wl[91] vdd gnd cell_6t
Xbit_r92_c41 bl[41] br[41] wl[92] vdd gnd cell_6t
Xbit_r93_c41 bl[41] br[41] wl[93] vdd gnd cell_6t
Xbit_r94_c41 bl[41] br[41] wl[94] vdd gnd cell_6t
Xbit_r95_c41 bl[41] br[41] wl[95] vdd gnd cell_6t
Xbit_r96_c41 bl[41] br[41] wl[96] vdd gnd cell_6t
Xbit_r97_c41 bl[41] br[41] wl[97] vdd gnd cell_6t
Xbit_r98_c41 bl[41] br[41] wl[98] vdd gnd cell_6t
Xbit_r99_c41 bl[41] br[41] wl[99] vdd gnd cell_6t
Xbit_r100_c41 bl[41] br[41] wl[100] vdd gnd cell_6t
Xbit_r101_c41 bl[41] br[41] wl[101] vdd gnd cell_6t
Xbit_r102_c41 bl[41] br[41] wl[102] vdd gnd cell_6t
Xbit_r103_c41 bl[41] br[41] wl[103] vdd gnd cell_6t
Xbit_r104_c41 bl[41] br[41] wl[104] vdd gnd cell_6t
Xbit_r105_c41 bl[41] br[41] wl[105] vdd gnd cell_6t
Xbit_r106_c41 bl[41] br[41] wl[106] vdd gnd cell_6t
Xbit_r107_c41 bl[41] br[41] wl[107] vdd gnd cell_6t
Xbit_r108_c41 bl[41] br[41] wl[108] vdd gnd cell_6t
Xbit_r109_c41 bl[41] br[41] wl[109] vdd gnd cell_6t
Xbit_r110_c41 bl[41] br[41] wl[110] vdd gnd cell_6t
Xbit_r111_c41 bl[41] br[41] wl[111] vdd gnd cell_6t
Xbit_r112_c41 bl[41] br[41] wl[112] vdd gnd cell_6t
Xbit_r113_c41 bl[41] br[41] wl[113] vdd gnd cell_6t
Xbit_r114_c41 bl[41] br[41] wl[114] vdd gnd cell_6t
Xbit_r115_c41 bl[41] br[41] wl[115] vdd gnd cell_6t
Xbit_r116_c41 bl[41] br[41] wl[116] vdd gnd cell_6t
Xbit_r117_c41 bl[41] br[41] wl[117] vdd gnd cell_6t
Xbit_r118_c41 bl[41] br[41] wl[118] vdd gnd cell_6t
Xbit_r119_c41 bl[41] br[41] wl[119] vdd gnd cell_6t
Xbit_r120_c41 bl[41] br[41] wl[120] vdd gnd cell_6t
Xbit_r121_c41 bl[41] br[41] wl[121] vdd gnd cell_6t
Xbit_r122_c41 bl[41] br[41] wl[122] vdd gnd cell_6t
Xbit_r123_c41 bl[41] br[41] wl[123] vdd gnd cell_6t
Xbit_r124_c41 bl[41] br[41] wl[124] vdd gnd cell_6t
Xbit_r125_c41 bl[41] br[41] wl[125] vdd gnd cell_6t
Xbit_r126_c41 bl[41] br[41] wl[126] vdd gnd cell_6t
Xbit_r127_c41 bl[41] br[41] wl[127] vdd gnd cell_6t
Xbit_r0_c42 bl[42] br[42] wl[0] vdd gnd cell_6t
Xbit_r1_c42 bl[42] br[42] wl[1] vdd gnd cell_6t
Xbit_r2_c42 bl[42] br[42] wl[2] vdd gnd cell_6t
Xbit_r3_c42 bl[42] br[42] wl[3] vdd gnd cell_6t
Xbit_r4_c42 bl[42] br[42] wl[4] vdd gnd cell_6t
Xbit_r5_c42 bl[42] br[42] wl[5] vdd gnd cell_6t
Xbit_r6_c42 bl[42] br[42] wl[6] vdd gnd cell_6t
Xbit_r7_c42 bl[42] br[42] wl[7] vdd gnd cell_6t
Xbit_r8_c42 bl[42] br[42] wl[8] vdd gnd cell_6t
Xbit_r9_c42 bl[42] br[42] wl[9] vdd gnd cell_6t
Xbit_r10_c42 bl[42] br[42] wl[10] vdd gnd cell_6t
Xbit_r11_c42 bl[42] br[42] wl[11] vdd gnd cell_6t
Xbit_r12_c42 bl[42] br[42] wl[12] vdd gnd cell_6t
Xbit_r13_c42 bl[42] br[42] wl[13] vdd gnd cell_6t
Xbit_r14_c42 bl[42] br[42] wl[14] vdd gnd cell_6t
Xbit_r15_c42 bl[42] br[42] wl[15] vdd gnd cell_6t
Xbit_r16_c42 bl[42] br[42] wl[16] vdd gnd cell_6t
Xbit_r17_c42 bl[42] br[42] wl[17] vdd gnd cell_6t
Xbit_r18_c42 bl[42] br[42] wl[18] vdd gnd cell_6t
Xbit_r19_c42 bl[42] br[42] wl[19] vdd gnd cell_6t
Xbit_r20_c42 bl[42] br[42] wl[20] vdd gnd cell_6t
Xbit_r21_c42 bl[42] br[42] wl[21] vdd gnd cell_6t
Xbit_r22_c42 bl[42] br[42] wl[22] vdd gnd cell_6t
Xbit_r23_c42 bl[42] br[42] wl[23] vdd gnd cell_6t
Xbit_r24_c42 bl[42] br[42] wl[24] vdd gnd cell_6t
Xbit_r25_c42 bl[42] br[42] wl[25] vdd gnd cell_6t
Xbit_r26_c42 bl[42] br[42] wl[26] vdd gnd cell_6t
Xbit_r27_c42 bl[42] br[42] wl[27] vdd gnd cell_6t
Xbit_r28_c42 bl[42] br[42] wl[28] vdd gnd cell_6t
Xbit_r29_c42 bl[42] br[42] wl[29] vdd gnd cell_6t
Xbit_r30_c42 bl[42] br[42] wl[30] vdd gnd cell_6t
Xbit_r31_c42 bl[42] br[42] wl[31] vdd gnd cell_6t
Xbit_r32_c42 bl[42] br[42] wl[32] vdd gnd cell_6t
Xbit_r33_c42 bl[42] br[42] wl[33] vdd gnd cell_6t
Xbit_r34_c42 bl[42] br[42] wl[34] vdd gnd cell_6t
Xbit_r35_c42 bl[42] br[42] wl[35] vdd gnd cell_6t
Xbit_r36_c42 bl[42] br[42] wl[36] vdd gnd cell_6t
Xbit_r37_c42 bl[42] br[42] wl[37] vdd gnd cell_6t
Xbit_r38_c42 bl[42] br[42] wl[38] vdd gnd cell_6t
Xbit_r39_c42 bl[42] br[42] wl[39] vdd gnd cell_6t
Xbit_r40_c42 bl[42] br[42] wl[40] vdd gnd cell_6t
Xbit_r41_c42 bl[42] br[42] wl[41] vdd gnd cell_6t
Xbit_r42_c42 bl[42] br[42] wl[42] vdd gnd cell_6t
Xbit_r43_c42 bl[42] br[42] wl[43] vdd gnd cell_6t
Xbit_r44_c42 bl[42] br[42] wl[44] vdd gnd cell_6t
Xbit_r45_c42 bl[42] br[42] wl[45] vdd gnd cell_6t
Xbit_r46_c42 bl[42] br[42] wl[46] vdd gnd cell_6t
Xbit_r47_c42 bl[42] br[42] wl[47] vdd gnd cell_6t
Xbit_r48_c42 bl[42] br[42] wl[48] vdd gnd cell_6t
Xbit_r49_c42 bl[42] br[42] wl[49] vdd gnd cell_6t
Xbit_r50_c42 bl[42] br[42] wl[50] vdd gnd cell_6t
Xbit_r51_c42 bl[42] br[42] wl[51] vdd gnd cell_6t
Xbit_r52_c42 bl[42] br[42] wl[52] vdd gnd cell_6t
Xbit_r53_c42 bl[42] br[42] wl[53] vdd gnd cell_6t
Xbit_r54_c42 bl[42] br[42] wl[54] vdd gnd cell_6t
Xbit_r55_c42 bl[42] br[42] wl[55] vdd gnd cell_6t
Xbit_r56_c42 bl[42] br[42] wl[56] vdd gnd cell_6t
Xbit_r57_c42 bl[42] br[42] wl[57] vdd gnd cell_6t
Xbit_r58_c42 bl[42] br[42] wl[58] vdd gnd cell_6t
Xbit_r59_c42 bl[42] br[42] wl[59] vdd gnd cell_6t
Xbit_r60_c42 bl[42] br[42] wl[60] vdd gnd cell_6t
Xbit_r61_c42 bl[42] br[42] wl[61] vdd gnd cell_6t
Xbit_r62_c42 bl[42] br[42] wl[62] vdd gnd cell_6t
Xbit_r63_c42 bl[42] br[42] wl[63] vdd gnd cell_6t
Xbit_r64_c42 bl[42] br[42] wl[64] vdd gnd cell_6t
Xbit_r65_c42 bl[42] br[42] wl[65] vdd gnd cell_6t
Xbit_r66_c42 bl[42] br[42] wl[66] vdd gnd cell_6t
Xbit_r67_c42 bl[42] br[42] wl[67] vdd gnd cell_6t
Xbit_r68_c42 bl[42] br[42] wl[68] vdd gnd cell_6t
Xbit_r69_c42 bl[42] br[42] wl[69] vdd gnd cell_6t
Xbit_r70_c42 bl[42] br[42] wl[70] vdd gnd cell_6t
Xbit_r71_c42 bl[42] br[42] wl[71] vdd gnd cell_6t
Xbit_r72_c42 bl[42] br[42] wl[72] vdd gnd cell_6t
Xbit_r73_c42 bl[42] br[42] wl[73] vdd gnd cell_6t
Xbit_r74_c42 bl[42] br[42] wl[74] vdd gnd cell_6t
Xbit_r75_c42 bl[42] br[42] wl[75] vdd gnd cell_6t
Xbit_r76_c42 bl[42] br[42] wl[76] vdd gnd cell_6t
Xbit_r77_c42 bl[42] br[42] wl[77] vdd gnd cell_6t
Xbit_r78_c42 bl[42] br[42] wl[78] vdd gnd cell_6t
Xbit_r79_c42 bl[42] br[42] wl[79] vdd gnd cell_6t
Xbit_r80_c42 bl[42] br[42] wl[80] vdd gnd cell_6t
Xbit_r81_c42 bl[42] br[42] wl[81] vdd gnd cell_6t
Xbit_r82_c42 bl[42] br[42] wl[82] vdd gnd cell_6t
Xbit_r83_c42 bl[42] br[42] wl[83] vdd gnd cell_6t
Xbit_r84_c42 bl[42] br[42] wl[84] vdd gnd cell_6t
Xbit_r85_c42 bl[42] br[42] wl[85] vdd gnd cell_6t
Xbit_r86_c42 bl[42] br[42] wl[86] vdd gnd cell_6t
Xbit_r87_c42 bl[42] br[42] wl[87] vdd gnd cell_6t
Xbit_r88_c42 bl[42] br[42] wl[88] vdd gnd cell_6t
Xbit_r89_c42 bl[42] br[42] wl[89] vdd gnd cell_6t
Xbit_r90_c42 bl[42] br[42] wl[90] vdd gnd cell_6t
Xbit_r91_c42 bl[42] br[42] wl[91] vdd gnd cell_6t
Xbit_r92_c42 bl[42] br[42] wl[92] vdd gnd cell_6t
Xbit_r93_c42 bl[42] br[42] wl[93] vdd gnd cell_6t
Xbit_r94_c42 bl[42] br[42] wl[94] vdd gnd cell_6t
Xbit_r95_c42 bl[42] br[42] wl[95] vdd gnd cell_6t
Xbit_r96_c42 bl[42] br[42] wl[96] vdd gnd cell_6t
Xbit_r97_c42 bl[42] br[42] wl[97] vdd gnd cell_6t
Xbit_r98_c42 bl[42] br[42] wl[98] vdd gnd cell_6t
Xbit_r99_c42 bl[42] br[42] wl[99] vdd gnd cell_6t
Xbit_r100_c42 bl[42] br[42] wl[100] vdd gnd cell_6t
Xbit_r101_c42 bl[42] br[42] wl[101] vdd gnd cell_6t
Xbit_r102_c42 bl[42] br[42] wl[102] vdd gnd cell_6t
Xbit_r103_c42 bl[42] br[42] wl[103] vdd gnd cell_6t
Xbit_r104_c42 bl[42] br[42] wl[104] vdd gnd cell_6t
Xbit_r105_c42 bl[42] br[42] wl[105] vdd gnd cell_6t
Xbit_r106_c42 bl[42] br[42] wl[106] vdd gnd cell_6t
Xbit_r107_c42 bl[42] br[42] wl[107] vdd gnd cell_6t
Xbit_r108_c42 bl[42] br[42] wl[108] vdd gnd cell_6t
Xbit_r109_c42 bl[42] br[42] wl[109] vdd gnd cell_6t
Xbit_r110_c42 bl[42] br[42] wl[110] vdd gnd cell_6t
Xbit_r111_c42 bl[42] br[42] wl[111] vdd gnd cell_6t
Xbit_r112_c42 bl[42] br[42] wl[112] vdd gnd cell_6t
Xbit_r113_c42 bl[42] br[42] wl[113] vdd gnd cell_6t
Xbit_r114_c42 bl[42] br[42] wl[114] vdd gnd cell_6t
Xbit_r115_c42 bl[42] br[42] wl[115] vdd gnd cell_6t
Xbit_r116_c42 bl[42] br[42] wl[116] vdd gnd cell_6t
Xbit_r117_c42 bl[42] br[42] wl[117] vdd gnd cell_6t
Xbit_r118_c42 bl[42] br[42] wl[118] vdd gnd cell_6t
Xbit_r119_c42 bl[42] br[42] wl[119] vdd gnd cell_6t
Xbit_r120_c42 bl[42] br[42] wl[120] vdd gnd cell_6t
Xbit_r121_c42 bl[42] br[42] wl[121] vdd gnd cell_6t
Xbit_r122_c42 bl[42] br[42] wl[122] vdd gnd cell_6t
Xbit_r123_c42 bl[42] br[42] wl[123] vdd gnd cell_6t
Xbit_r124_c42 bl[42] br[42] wl[124] vdd gnd cell_6t
Xbit_r125_c42 bl[42] br[42] wl[125] vdd gnd cell_6t
Xbit_r126_c42 bl[42] br[42] wl[126] vdd gnd cell_6t
Xbit_r127_c42 bl[42] br[42] wl[127] vdd gnd cell_6t
Xbit_r0_c43 bl[43] br[43] wl[0] vdd gnd cell_6t
Xbit_r1_c43 bl[43] br[43] wl[1] vdd gnd cell_6t
Xbit_r2_c43 bl[43] br[43] wl[2] vdd gnd cell_6t
Xbit_r3_c43 bl[43] br[43] wl[3] vdd gnd cell_6t
Xbit_r4_c43 bl[43] br[43] wl[4] vdd gnd cell_6t
Xbit_r5_c43 bl[43] br[43] wl[5] vdd gnd cell_6t
Xbit_r6_c43 bl[43] br[43] wl[6] vdd gnd cell_6t
Xbit_r7_c43 bl[43] br[43] wl[7] vdd gnd cell_6t
Xbit_r8_c43 bl[43] br[43] wl[8] vdd gnd cell_6t
Xbit_r9_c43 bl[43] br[43] wl[9] vdd gnd cell_6t
Xbit_r10_c43 bl[43] br[43] wl[10] vdd gnd cell_6t
Xbit_r11_c43 bl[43] br[43] wl[11] vdd gnd cell_6t
Xbit_r12_c43 bl[43] br[43] wl[12] vdd gnd cell_6t
Xbit_r13_c43 bl[43] br[43] wl[13] vdd gnd cell_6t
Xbit_r14_c43 bl[43] br[43] wl[14] vdd gnd cell_6t
Xbit_r15_c43 bl[43] br[43] wl[15] vdd gnd cell_6t
Xbit_r16_c43 bl[43] br[43] wl[16] vdd gnd cell_6t
Xbit_r17_c43 bl[43] br[43] wl[17] vdd gnd cell_6t
Xbit_r18_c43 bl[43] br[43] wl[18] vdd gnd cell_6t
Xbit_r19_c43 bl[43] br[43] wl[19] vdd gnd cell_6t
Xbit_r20_c43 bl[43] br[43] wl[20] vdd gnd cell_6t
Xbit_r21_c43 bl[43] br[43] wl[21] vdd gnd cell_6t
Xbit_r22_c43 bl[43] br[43] wl[22] vdd gnd cell_6t
Xbit_r23_c43 bl[43] br[43] wl[23] vdd gnd cell_6t
Xbit_r24_c43 bl[43] br[43] wl[24] vdd gnd cell_6t
Xbit_r25_c43 bl[43] br[43] wl[25] vdd gnd cell_6t
Xbit_r26_c43 bl[43] br[43] wl[26] vdd gnd cell_6t
Xbit_r27_c43 bl[43] br[43] wl[27] vdd gnd cell_6t
Xbit_r28_c43 bl[43] br[43] wl[28] vdd gnd cell_6t
Xbit_r29_c43 bl[43] br[43] wl[29] vdd gnd cell_6t
Xbit_r30_c43 bl[43] br[43] wl[30] vdd gnd cell_6t
Xbit_r31_c43 bl[43] br[43] wl[31] vdd gnd cell_6t
Xbit_r32_c43 bl[43] br[43] wl[32] vdd gnd cell_6t
Xbit_r33_c43 bl[43] br[43] wl[33] vdd gnd cell_6t
Xbit_r34_c43 bl[43] br[43] wl[34] vdd gnd cell_6t
Xbit_r35_c43 bl[43] br[43] wl[35] vdd gnd cell_6t
Xbit_r36_c43 bl[43] br[43] wl[36] vdd gnd cell_6t
Xbit_r37_c43 bl[43] br[43] wl[37] vdd gnd cell_6t
Xbit_r38_c43 bl[43] br[43] wl[38] vdd gnd cell_6t
Xbit_r39_c43 bl[43] br[43] wl[39] vdd gnd cell_6t
Xbit_r40_c43 bl[43] br[43] wl[40] vdd gnd cell_6t
Xbit_r41_c43 bl[43] br[43] wl[41] vdd gnd cell_6t
Xbit_r42_c43 bl[43] br[43] wl[42] vdd gnd cell_6t
Xbit_r43_c43 bl[43] br[43] wl[43] vdd gnd cell_6t
Xbit_r44_c43 bl[43] br[43] wl[44] vdd gnd cell_6t
Xbit_r45_c43 bl[43] br[43] wl[45] vdd gnd cell_6t
Xbit_r46_c43 bl[43] br[43] wl[46] vdd gnd cell_6t
Xbit_r47_c43 bl[43] br[43] wl[47] vdd gnd cell_6t
Xbit_r48_c43 bl[43] br[43] wl[48] vdd gnd cell_6t
Xbit_r49_c43 bl[43] br[43] wl[49] vdd gnd cell_6t
Xbit_r50_c43 bl[43] br[43] wl[50] vdd gnd cell_6t
Xbit_r51_c43 bl[43] br[43] wl[51] vdd gnd cell_6t
Xbit_r52_c43 bl[43] br[43] wl[52] vdd gnd cell_6t
Xbit_r53_c43 bl[43] br[43] wl[53] vdd gnd cell_6t
Xbit_r54_c43 bl[43] br[43] wl[54] vdd gnd cell_6t
Xbit_r55_c43 bl[43] br[43] wl[55] vdd gnd cell_6t
Xbit_r56_c43 bl[43] br[43] wl[56] vdd gnd cell_6t
Xbit_r57_c43 bl[43] br[43] wl[57] vdd gnd cell_6t
Xbit_r58_c43 bl[43] br[43] wl[58] vdd gnd cell_6t
Xbit_r59_c43 bl[43] br[43] wl[59] vdd gnd cell_6t
Xbit_r60_c43 bl[43] br[43] wl[60] vdd gnd cell_6t
Xbit_r61_c43 bl[43] br[43] wl[61] vdd gnd cell_6t
Xbit_r62_c43 bl[43] br[43] wl[62] vdd gnd cell_6t
Xbit_r63_c43 bl[43] br[43] wl[63] vdd gnd cell_6t
Xbit_r64_c43 bl[43] br[43] wl[64] vdd gnd cell_6t
Xbit_r65_c43 bl[43] br[43] wl[65] vdd gnd cell_6t
Xbit_r66_c43 bl[43] br[43] wl[66] vdd gnd cell_6t
Xbit_r67_c43 bl[43] br[43] wl[67] vdd gnd cell_6t
Xbit_r68_c43 bl[43] br[43] wl[68] vdd gnd cell_6t
Xbit_r69_c43 bl[43] br[43] wl[69] vdd gnd cell_6t
Xbit_r70_c43 bl[43] br[43] wl[70] vdd gnd cell_6t
Xbit_r71_c43 bl[43] br[43] wl[71] vdd gnd cell_6t
Xbit_r72_c43 bl[43] br[43] wl[72] vdd gnd cell_6t
Xbit_r73_c43 bl[43] br[43] wl[73] vdd gnd cell_6t
Xbit_r74_c43 bl[43] br[43] wl[74] vdd gnd cell_6t
Xbit_r75_c43 bl[43] br[43] wl[75] vdd gnd cell_6t
Xbit_r76_c43 bl[43] br[43] wl[76] vdd gnd cell_6t
Xbit_r77_c43 bl[43] br[43] wl[77] vdd gnd cell_6t
Xbit_r78_c43 bl[43] br[43] wl[78] vdd gnd cell_6t
Xbit_r79_c43 bl[43] br[43] wl[79] vdd gnd cell_6t
Xbit_r80_c43 bl[43] br[43] wl[80] vdd gnd cell_6t
Xbit_r81_c43 bl[43] br[43] wl[81] vdd gnd cell_6t
Xbit_r82_c43 bl[43] br[43] wl[82] vdd gnd cell_6t
Xbit_r83_c43 bl[43] br[43] wl[83] vdd gnd cell_6t
Xbit_r84_c43 bl[43] br[43] wl[84] vdd gnd cell_6t
Xbit_r85_c43 bl[43] br[43] wl[85] vdd gnd cell_6t
Xbit_r86_c43 bl[43] br[43] wl[86] vdd gnd cell_6t
Xbit_r87_c43 bl[43] br[43] wl[87] vdd gnd cell_6t
Xbit_r88_c43 bl[43] br[43] wl[88] vdd gnd cell_6t
Xbit_r89_c43 bl[43] br[43] wl[89] vdd gnd cell_6t
Xbit_r90_c43 bl[43] br[43] wl[90] vdd gnd cell_6t
Xbit_r91_c43 bl[43] br[43] wl[91] vdd gnd cell_6t
Xbit_r92_c43 bl[43] br[43] wl[92] vdd gnd cell_6t
Xbit_r93_c43 bl[43] br[43] wl[93] vdd gnd cell_6t
Xbit_r94_c43 bl[43] br[43] wl[94] vdd gnd cell_6t
Xbit_r95_c43 bl[43] br[43] wl[95] vdd gnd cell_6t
Xbit_r96_c43 bl[43] br[43] wl[96] vdd gnd cell_6t
Xbit_r97_c43 bl[43] br[43] wl[97] vdd gnd cell_6t
Xbit_r98_c43 bl[43] br[43] wl[98] vdd gnd cell_6t
Xbit_r99_c43 bl[43] br[43] wl[99] vdd gnd cell_6t
Xbit_r100_c43 bl[43] br[43] wl[100] vdd gnd cell_6t
Xbit_r101_c43 bl[43] br[43] wl[101] vdd gnd cell_6t
Xbit_r102_c43 bl[43] br[43] wl[102] vdd gnd cell_6t
Xbit_r103_c43 bl[43] br[43] wl[103] vdd gnd cell_6t
Xbit_r104_c43 bl[43] br[43] wl[104] vdd gnd cell_6t
Xbit_r105_c43 bl[43] br[43] wl[105] vdd gnd cell_6t
Xbit_r106_c43 bl[43] br[43] wl[106] vdd gnd cell_6t
Xbit_r107_c43 bl[43] br[43] wl[107] vdd gnd cell_6t
Xbit_r108_c43 bl[43] br[43] wl[108] vdd gnd cell_6t
Xbit_r109_c43 bl[43] br[43] wl[109] vdd gnd cell_6t
Xbit_r110_c43 bl[43] br[43] wl[110] vdd gnd cell_6t
Xbit_r111_c43 bl[43] br[43] wl[111] vdd gnd cell_6t
Xbit_r112_c43 bl[43] br[43] wl[112] vdd gnd cell_6t
Xbit_r113_c43 bl[43] br[43] wl[113] vdd gnd cell_6t
Xbit_r114_c43 bl[43] br[43] wl[114] vdd gnd cell_6t
Xbit_r115_c43 bl[43] br[43] wl[115] vdd gnd cell_6t
Xbit_r116_c43 bl[43] br[43] wl[116] vdd gnd cell_6t
Xbit_r117_c43 bl[43] br[43] wl[117] vdd gnd cell_6t
Xbit_r118_c43 bl[43] br[43] wl[118] vdd gnd cell_6t
Xbit_r119_c43 bl[43] br[43] wl[119] vdd gnd cell_6t
Xbit_r120_c43 bl[43] br[43] wl[120] vdd gnd cell_6t
Xbit_r121_c43 bl[43] br[43] wl[121] vdd gnd cell_6t
Xbit_r122_c43 bl[43] br[43] wl[122] vdd gnd cell_6t
Xbit_r123_c43 bl[43] br[43] wl[123] vdd gnd cell_6t
Xbit_r124_c43 bl[43] br[43] wl[124] vdd gnd cell_6t
Xbit_r125_c43 bl[43] br[43] wl[125] vdd gnd cell_6t
Xbit_r126_c43 bl[43] br[43] wl[126] vdd gnd cell_6t
Xbit_r127_c43 bl[43] br[43] wl[127] vdd gnd cell_6t
Xbit_r0_c44 bl[44] br[44] wl[0] vdd gnd cell_6t
Xbit_r1_c44 bl[44] br[44] wl[1] vdd gnd cell_6t
Xbit_r2_c44 bl[44] br[44] wl[2] vdd gnd cell_6t
Xbit_r3_c44 bl[44] br[44] wl[3] vdd gnd cell_6t
Xbit_r4_c44 bl[44] br[44] wl[4] vdd gnd cell_6t
Xbit_r5_c44 bl[44] br[44] wl[5] vdd gnd cell_6t
Xbit_r6_c44 bl[44] br[44] wl[6] vdd gnd cell_6t
Xbit_r7_c44 bl[44] br[44] wl[7] vdd gnd cell_6t
Xbit_r8_c44 bl[44] br[44] wl[8] vdd gnd cell_6t
Xbit_r9_c44 bl[44] br[44] wl[9] vdd gnd cell_6t
Xbit_r10_c44 bl[44] br[44] wl[10] vdd gnd cell_6t
Xbit_r11_c44 bl[44] br[44] wl[11] vdd gnd cell_6t
Xbit_r12_c44 bl[44] br[44] wl[12] vdd gnd cell_6t
Xbit_r13_c44 bl[44] br[44] wl[13] vdd gnd cell_6t
Xbit_r14_c44 bl[44] br[44] wl[14] vdd gnd cell_6t
Xbit_r15_c44 bl[44] br[44] wl[15] vdd gnd cell_6t
Xbit_r16_c44 bl[44] br[44] wl[16] vdd gnd cell_6t
Xbit_r17_c44 bl[44] br[44] wl[17] vdd gnd cell_6t
Xbit_r18_c44 bl[44] br[44] wl[18] vdd gnd cell_6t
Xbit_r19_c44 bl[44] br[44] wl[19] vdd gnd cell_6t
Xbit_r20_c44 bl[44] br[44] wl[20] vdd gnd cell_6t
Xbit_r21_c44 bl[44] br[44] wl[21] vdd gnd cell_6t
Xbit_r22_c44 bl[44] br[44] wl[22] vdd gnd cell_6t
Xbit_r23_c44 bl[44] br[44] wl[23] vdd gnd cell_6t
Xbit_r24_c44 bl[44] br[44] wl[24] vdd gnd cell_6t
Xbit_r25_c44 bl[44] br[44] wl[25] vdd gnd cell_6t
Xbit_r26_c44 bl[44] br[44] wl[26] vdd gnd cell_6t
Xbit_r27_c44 bl[44] br[44] wl[27] vdd gnd cell_6t
Xbit_r28_c44 bl[44] br[44] wl[28] vdd gnd cell_6t
Xbit_r29_c44 bl[44] br[44] wl[29] vdd gnd cell_6t
Xbit_r30_c44 bl[44] br[44] wl[30] vdd gnd cell_6t
Xbit_r31_c44 bl[44] br[44] wl[31] vdd gnd cell_6t
Xbit_r32_c44 bl[44] br[44] wl[32] vdd gnd cell_6t
Xbit_r33_c44 bl[44] br[44] wl[33] vdd gnd cell_6t
Xbit_r34_c44 bl[44] br[44] wl[34] vdd gnd cell_6t
Xbit_r35_c44 bl[44] br[44] wl[35] vdd gnd cell_6t
Xbit_r36_c44 bl[44] br[44] wl[36] vdd gnd cell_6t
Xbit_r37_c44 bl[44] br[44] wl[37] vdd gnd cell_6t
Xbit_r38_c44 bl[44] br[44] wl[38] vdd gnd cell_6t
Xbit_r39_c44 bl[44] br[44] wl[39] vdd gnd cell_6t
Xbit_r40_c44 bl[44] br[44] wl[40] vdd gnd cell_6t
Xbit_r41_c44 bl[44] br[44] wl[41] vdd gnd cell_6t
Xbit_r42_c44 bl[44] br[44] wl[42] vdd gnd cell_6t
Xbit_r43_c44 bl[44] br[44] wl[43] vdd gnd cell_6t
Xbit_r44_c44 bl[44] br[44] wl[44] vdd gnd cell_6t
Xbit_r45_c44 bl[44] br[44] wl[45] vdd gnd cell_6t
Xbit_r46_c44 bl[44] br[44] wl[46] vdd gnd cell_6t
Xbit_r47_c44 bl[44] br[44] wl[47] vdd gnd cell_6t
Xbit_r48_c44 bl[44] br[44] wl[48] vdd gnd cell_6t
Xbit_r49_c44 bl[44] br[44] wl[49] vdd gnd cell_6t
Xbit_r50_c44 bl[44] br[44] wl[50] vdd gnd cell_6t
Xbit_r51_c44 bl[44] br[44] wl[51] vdd gnd cell_6t
Xbit_r52_c44 bl[44] br[44] wl[52] vdd gnd cell_6t
Xbit_r53_c44 bl[44] br[44] wl[53] vdd gnd cell_6t
Xbit_r54_c44 bl[44] br[44] wl[54] vdd gnd cell_6t
Xbit_r55_c44 bl[44] br[44] wl[55] vdd gnd cell_6t
Xbit_r56_c44 bl[44] br[44] wl[56] vdd gnd cell_6t
Xbit_r57_c44 bl[44] br[44] wl[57] vdd gnd cell_6t
Xbit_r58_c44 bl[44] br[44] wl[58] vdd gnd cell_6t
Xbit_r59_c44 bl[44] br[44] wl[59] vdd gnd cell_6t
Xbit_r60_c44 bl[44] br[44] wl[60] vdd gnd cell_6t
Xbit_r61_c44 bl[44] br[44] wl[61] vdd gnd cell_6t
Xbit_r62_c44 bl[44] br[44] wl[62] vdd gnd cell_6t
Xbit_r63_c44 bl[44] br[44] wl[63] vdd gnd cell_6t
Xbit_r64_c44 bl[44] br[44] wl[64] vdd gnd cell_6t
Xbit_r65_c44 bl[44] br[44] wl[65] vdd gnd cell_6t
Xbit_r66_c44 bl[44] br[44] wl[66] vdd gnd cell_6t
Xbit_r67_c44 bl[44] br[44] wl[67] vdd gnd cell_6t
Xbit_r68_c44 bl[44] br[44] wl[68] vdd gnd cell_6t
Xbit_r69_c44 bl[44] br[44] wl[69] vdd gnd cell_6t
Xbit_r70_c44 bl[44] br[44] wl[70] vdd gnd cell_6t
Xbit_r71_c44 bl[44] br[44] wl[71] vdd gnd cell_6t
Xbit_r72_c44 bl[44] br[44] wl[72] vdd gnd cell_6t
Xbit_r73_c44 bl[44] br[44] wl[73] vdd gnd cell_6t
Xbit_r74_c44 bl[44] br[44] wl[74] vdd gnd cell_6t
Xbit_r75_c44 bl[44] br[44] wl[75] vdd gnd cell_6t
Xbit_r76_c44 bl[44] br[44] wl[76] vdd gnd cell_6t
Xbit_r77_c44 bl[44] br[44] wl[77] vdd gnd cell_6t
Xbit_r78_c44 bl[44] br[44] wl[78] vdd gnd cell_6t
Xbit_r79_c44 bl[44] br[44] wl[79] vdd gnd cell_6t
Xbit_r80_c44 bl[44] br[44] wl[80] vdd gnd cell_6t
Xbit_r81_c44 bl[44] br[44] wl[81] vdd gnd cell_6t
Xbit_r82_c44 bl[44] br[44] wl[82] vdd gnd cell_6t
Xbit_r83_c44 bl[44] br[44] wl[83] vdd gnd cell_6t
Xbit_r84_c44 bl[44] br[44] wl[84] vdd gnd cell_6t
Xbit_r85_c44 bl[44] br[44] wl[85] vdd gnd cell_6t
Xbit_r86_c44 bl[44] br[44] wl[86] vdd gnd cell_6t
Xbit_r87_c44 bl[44] br[44] wl[87] vdd gnd cell_6t
Xbit_r88_c44 bl[44] br[44] wl[88] vdd gnd cell_6t
Xbit_r89_c44 bl[44] br[44] wl[89] vdd gnd cell_6t
Xbit_r90_c44 bl[44] br[44] wl[90] vdd gnd cell_6t
Xbit_r91_c44 bl[44] br[44] wl[91] vdd gnd cell_6t
Xbit_r92_c44 bl[44] br[44] wl[92] vdd gnd cell_6t
Xbit_r93_c44 bl[44] br[44] wl[93] vdd gnd cell_6t
Xbit_r94_c44 bl[44] br[44] wl[94] vdd gnd cell_6t
Xbit_r95_c44 bl[44] br[44] wl[95] vdd gnd cell_6t
Xbit_r96_c44 bl[44] br[44] wl[96] vdd gnd cell_6t
Xbit_r97_c44 bl[44] br[44] wl[97] vdd gnd cell_6t
Xbit_r98_c44 bl[44] br[44] wl[98] vdd gnd cell_6t
Xbit_r99_c44 bl[44] br[44] wl[99] vdd gnd cell_6t
Xbit_r100_c44 bl[44] br[44] wl[100] vdd gnd cell_6t
Xbit_r101_c44 bl[44] br[44] wl[101] vdd gnd cell_6t
Xbit_r102_c44 bl[44] br[44] wl[102] vdd gnd cell_6t
Xbit_r103_c44 bl[44] br[44] wl[103] vdd gnd cell_6t
Xbit_r104_c44 bl[44] br[44] wl[104] vdd gnd cell_6t
Xbit_r105_c44 bl[44] br[44] wl[105] vdd gnd cell_6t
Xbit_r106_c44 bl[44] br[44] wl[106] vdd gnd cell_6t
Xbit_r107_c44 bl[44] br[44] wl[107] vdd gnd cell_6t
Xbit_r108_c44 bl[44] br[44] wl[108] vdd gnd cell_6t
Xbit_r109_c44 bl[44] br[44] wl[109] vdd gnd cell_6t
Xbit_r110_c44 bl[44] br[44] wl[110] vdd gnd cell_6t
Xbit_r111_c44 bl[44] br[44] wl[111] vdd gnd cell_6t
Xbit_r112_c44 bl[44] br[44] wl[112] vdd gnd cell_6t
Xbit_r113_c44 bl[44] br[44] wl[113] vdd gnd cell_6t
Xbit_r114_c44 bl[44] br[44] wl[114] vdd gnd cell_6t
Xbit_r115_c44 bl[44] br[44] wl[115] vdd gnd cell_6t
Xbit_r116_c44 bl[44] br[44] wl[116] vdd gnd cell_6t
Xbit_r117_c44 bl[44] br[44] wl[117] vdd gnd cell_6t
Xbit_r118_c44 bl[44] br[44] wl[118] vdd gnd cell_6t
Xbit_r119_c44 bl[44] br[44] wl[119] vdd gnd cell_6t
Xbit_r120_c44 bl[44] br[44] wl[120] vdd gnd cell_6t
Xbit_r121_c44 bl[44] br[44] wl[121] vdd gnd cell_6t
Xbit_r122_c44 bl[44] br[44] wl[122] vdd gnd cell_6t
Xbit_r123_c44 bl[44] br[44] wl[123] vdd gnd cell_6t
Xbit_r124_c44 bl[44] br[44] wl[124] vdd gnd cell_6t
Xbit_r125_c44 bl[44] br[44] wl[125] vdd gnd cell_6t
Xbit_r126_c44 bl[44] br[44] wl[126] vdd gnd cell_6t
Xbit_r127_c44 bl[44] br[44] wl[127] vdd gnd cell_6t
Xbit_r0_c45 bl[45] br[45] wl[0] vdd gnd cell_6t
Xbit_r1_c45 bl[45] br[45] wl[1] vdd gnd cell_6t
Xbit_r2_c45 bl[45] br[45] wl[2] vdd gnd cell_6t
Xbit_r3_c45 bl[45] br[45] wl[3] vdd gnd cell_6t
Xbit_r4_c45 bl[45] br[45] wl[4] vdd gnd cell_6t
Xbit_r5_c45 bl[45] br[45] wl[5] vdd gnd cell_6t
Xbit_r6_c45 bl[45] br[45] wl[6] vdd gnd cell_6t
Xbit_r7_c45 bl[45] br[45] wl[7] vdd gnd cell_6t
Xbit_r8_c45 bl[45] br[45] wl[8] vdd gnd cell_6t
Xbit_r9_c45 bl[45] br[45] wl[9] vdd gnd cell_6t
Xbit_r10_c45 bl[45] br[45] wl[10] vdd gnd cell_6t
Xbit_r11_c45 bl[45] br[45] wl[11] vdd gnd cell_6t
Xbit_r12_c45 bl[45] br[45] wl[12] vdd gnd cell_6t
Xbit_r13_c45 bl[45] br[45] wl[13] vdd gnd cell_6t
Xbit_r14_c45 bl[45] br[45] wl[14] vdd gnd cell_6t
Xbit_r15_c45 bl[45] br[45] wl[15] vdd gnd cell_6t
Xbit_r16_c45 bl[45] br[45] wl[16] vdd gnd cell_6t
Xbit_r17_c45 bl[45] br[45] wl[17] vdd gnd cell_6t
Xbit_r18_c45 bl[45] br[45] wl[18] vdd gnd cell_6t
Xbit_r19_c45 bl[45] br[45] wl[19] vdd gnd cell_6t
Xbit_r20_c45 bl[45] br[45] wl[20] vdd gnd cell_6t
Xbit_r21_c45 bl[45] br[45] wl[21] vdd gnd cell_6t
Xbit_r22_c45 bl[45] br[45] wl[22] vdd gnd cell_6t
Xbit_r23_c45 bl[45] br[45] wl[23] vdd gnd cell_6t
Xbit_r24_c45 bl[45] br[45] wl[24] vdd gnd cell_6t
Xbit_r25_c45 bl[45] br[45] wl[25] vdd gnd cell_6t
Xbit_r26_c45 bl[45] br[45] wl[26] vdd gnd cell_6t
Xbit_r27_c45 bl[45] br[45] wl[27] vdd gnd cell_6t
Xbit_r28_c45 bl[45] br[45] wl[28] vdd gnd cell_6t
Xbit_r29_c45 bl[45] br[45] wl[29] vdd gnd cell_6t
Xbit_r30_c45 bl[45] br[45] wl[30] vdd gnd cell_6t
Xbit_r31_c45 bl[45] br[45] wl[31] vdd gnd cell_6t
Xbit_r32_c45 bl[45] br[45] wl[32] vdd gnd cell_6t
Xbit_r33_c45 bl[45] br[45] wl[33] vdd gnd cell_6t
Xbit_r34_c45 bl[45] br[45] wl[34] vdd gnd cell_6t
Xbit_r35_c45 bl[45] br[45] wl[35] vdd gnd cell_6t
Xbit_r36_c45 bl[45] br[45] wl[36] vdd gnd cell_6t
Xbit_r37_c45 bl[45] br[45] wl[37] vdd gnd cell_6t
Xbit_r38_c45 bl[45] br[45] wl[38] vdd gnd cell_6t
Xbit_r39_c45 bl[45] br[45] wl[39] vdd gnd cell_6t
Xbit_r40_c45 bl[45] br[45] wl[40] vdd gnd cell_6t
Xbit_r41_c45 bl[45] br[45] wl[41] vdd gnd cell_6t
Xbit_r42_c45 bl[45] br[45] wl[42] vdd gnd cell_6t
Xbit_r43_c45 bl[45] br[45] wl[43] vdd gnd cell_6t
Xbit_r44_c45 bl[45] br[45] wl[44] vdd gnd cell_6t
Xbit_r45_c45 bl[45] br[45] wl[45] vdd gnd cell_6t
Xbit_r46_c45 bl[45] br[45] wl[46] vdd gnd cell_6t
Xbit_r47_c45 bl[45] br[45] wl[47] vdd gnd cell_6t
Xbit_r48_c45 bl[45] br[45] wl[48] vdd gnd cell_6t
Xbit_r49_c45 bl[45] br[45] wl[49] vdd gnd cell_6t
Xbit_r50_c45 bl[45] br[45] wl[50] vdd gnd cell_6t
Xbit_r51_c45 bl[45] br[45] wl[51] vdd gnd cell_6t
Xbit_r52_c45 bl[45] br[45] wl[52] vdd gnd cell_6t
Xbit_r53_c45 bl[45] br[45] wl[53] vdd gnd cell_6t
Xbit_r54_c45 bl[45] br[45] wl[54] vdd gnd cell_6t
Xbit_r55_c45 bl[45] br[45] wl[55] vdd gnd cell_6t
Xbit_r56_c45 bl[45] br[45] wl[56] vdd gnd cell_6t
Xbit_r57_c45 bl[45] br[45] wl[57] vdd gnd cell_6t
Xbit_r58_c45 bl[45] br[45] wl[58] vdd gnd cell_6t
Xbit_r59_c45 bl[45] br[45] wl[59] vdd gnd cell_6t
Xbit_r60_c45 bl[45] br[45] wl[60] vdd gnd cell_6t
Xbit_r61_c45 bl[45] br[45] wl[61] vdd gnd cell_6t
Xbit_r62_c45 bl[45] br[45] wl[62] vdd gnd cell_6t
Xbit_r63_c45 bl[45] br[45] wl[63] vdd gnd cell_6t
Xbit_r64_c45 bl[45] br[45] wl[64] vdd gnd cell_6t
Xbit_r65_c45 bl[45] br[45] wl[65] vdd gnd cell_6t
Xbit_r66_c45 bl[45] br[45] wl[66] vdd gnd cell_6t
Xbit_r67_c45 bl[45] br[45] wl[67] vdd gnd cell_6t
Xbit_r68_c45 bl[45] br[45] wl[68] vdd gnd cell_6t
Xbit_r69_c45 bl[45] br[45] wl[69] vdd gnd cell_6t
Xbit_r70_c45 bl[45] br[45] wl[70] vdd gnd cell_6t
Xbit_r71_c45 bl[45] br[45] wl[71] vdd gnd cell_6t
Xbit_r72_c45 bl[45] br[45] wl[72] vdd gnd cell_6t
Xbit_r73_c45 bl[45] br[45] wl[73] vdd gnd cell_6t
Xbit_r74_c45 bl[45] br[45] wl[74] vdd gnd cell_6t
Xbit_r75_c45 bl[45] br[45] wl[75] vdd gnd cell_6t
Xbit_r76_c45 bl[45] br[45] wl[76] vdd gnd cell_6t
Xbit_r77_c45 bl[45] br[45] wl[77] vdd gnd cell_6t
Xbit_r78_c45 bl[45] br[45] wl[78] vdd gnd cell_6t
Xbit_r79_c45 bl[45] br[45] wl[79] vdd gnd cell_6t
Xbit_r80_c45 bl[45] br[45] wl[80] vdd gnd cell_6t
Xbit_r81_c45 bl[45] br[45] wl[81] vdd gnd cell_6t
Xbit_r82_c45 bl[45] br[45] wl[82] vdd gnd cell_6t
Xbit_r83_c45 bl[45] br[45] wl[83] vdd gnd cell_6t
Xbit_r84_c45 bl[45] br[45] wl[84] vdd gnd cell_6t
Xbit_r85_c45 bl[45] br[45] wl[85] vdd gnd cell_6t
Xbit_r86_c45 bl[45] br[45] wl[86] vdd gnd cell_6t
Xbit_r87_c45 bl[45] br[45] wl[87] vdd gnd cell_6t
Xbit_r88_c45 bl[45] br[45] wl[88] vdd gnd cell_6t
Xbit_r89_c45 bl[45] br[45] wl[89] vdd gnd cell_6t
Xbit_r90_c45 bl[45] br[45] wl[90] vdd gnd cell_6t
Xbit_r91_c45 bl[45] br[45] wl[91] vdd gnd cell_6t
Xbit_r92_c45 bl[45] br[45] wl[92] vdd gnd cell_6t
Xbit_r93_c45 bl[45] br[45] wl[93] vdd gnd cell_6t
Xbit_r94_c45 bl[45] br[45] wl[94] vdd gnd cell_6t
Xbit_r95_c45 bl[45] br[45] wl[95] vdd gnd cell_6t
Xbit_r96_c45 bl[45] br[45] wl[96] vdd gnd cell_6t
Xbit_r97_c45 bl[45] br[45] wl[97] vdd gnd cell_6t
Xbit_r98_c45 bl[45] br[45] wl[98] vdd gnd cell_6t
Xbit_r99_c45 bl[45] br[45] wl[99] vdd gnd cell_6t
Xbit_r100_c45 bl[45] br[45] wl[100] vdd gnd cell_6t
Xbit_r101_c45 bl[45] br[45] wl[101] vdd gnd cell_6t
Xbit_r102_c45 bl[45] br[45] wl[102] vdd gnd cell_6t
Xbit_r103_c45 bl[45] br[45] wl[103] vdd gnd cell_6t
Xbit_r104_c45 bl[45] br[45] wl[104] vdd gnd cell_6t
Xbit_r105_c45 bl[45] br[45] wl[105] vdd gnd cell_6t
Xbit_r106_c45 bl[45] br[45] wl[106] vdd gnd cell_6t
Xbit_r107_c45 bl[45] br[45] wl[107] vdd gnd cell_6t
Xbit_r108_c45 bl[45] br[45] wl[108] vdd gnd cell_6t
Xbit_r109_c45 bl[45] br[45] wl[109] vdd gnd cell_6t
Xbit_r110_c45 bl[45] br[45] wl[110] vdd gnd cell_6t
Xbit_r111_c45 bl[45] br[45] wl[111] vdd gnd cell_6t
Xbit_r112_c45 bl[45] br[45] wl[112] vdd gnd cell_6t
Xbit_r113_c45 bl[45] br[45] wl[113] vdd gnd cell_6t
Xbit_r114_c45 bl[45] br[45] wl[114] vdd gnd cell_6t
Xbit_r115_c45 bl[45] br[45] wl[115] vdd gnd cell_6t
Xbit_r116_c45 bl[45] br[45] wl[116] vdd gnd cell_6t
Xbit_r117_c45 bl[45] br[45] wl[117] vdd gnd cell_6t
Xbit_r118_c45 bl[45] br[45] wl[118] vdd gnd cell_6t
Xbit_r119_c45 bl[45] br[45] wl[119] vdd gnd cell_6t
Xbit_r120_c45 bl[45] br[45] wl[120] vdd gnd cell_6t
Xbit_r121_c45 bl[45] br[45] wl[121] vdd gnd cell_6t
Xbit_r122_c45 bl[45] br[45] wl[122] vdd gnd cell_6t
Xbit_r123_c45 bl[45] br[45] wl[123] vdd gnd cell_6t
Xbit_r124_c45 bl[45] br[45] wl[124] vdd gnd cell_6t
Xbit_r125_c45 bl[45] br[45] wl[125] vdd gnd cell_6t
Xbit_r126_c45 bl[45] br[45] wl[126] vdd gnd cell_6t
Xbit_r127_c45 bl[45] br[45] wl[127] vdd gnd cell_6t
Xbit_r0_c46 bl[46] br[46] wl[0] vdd gnd cell_6t
Xbit_r1_c46 bl[46] br[46] wl[1] vdd gnd cell_6t
Xbit_r2_c46 bl[46] br[46] wl[2] vdd gnd cell_6t
Xbit_r3_c46 bl[46] br[46] wl[3] vdd gnd cell_6t
Xbit_r4_c46 bl[46] br[46] wl[4] vdd gnd cell_6t
Xbit_r5_c46 bl[46] br[46] wl[5] vdd gnd cell_6t
Xbit_r6_c46 bl[46] br[46] wl[6] vdd gnd cell_6t
Xbit_r7_c46 bl[46] br[46] wl[7] vdd gnd cell_6t
Xbit_r8_c46 bl[46] br[46] wl[8] vdd gnd cell_6t
Xbit_r9_c46 bl[46] br[46] wl[9] vdd gnd cell_6t
Xbit_r10_c46 bl[46] br[46] wl[10] vdd gnd cell_6t
Xbit_r11_c46 bl[46] br[46] wl[11] vdd gnd cell_6t
Xbit_r12_c46 bl[46] br[46] wl[12] vdd gnd cell_6t
Xbit_r13_c46 bl[46] br[46] wl[13] vdd gnd cell_6t
Xbit_r14_c46 bl[46] br[46] wl[14] vdd gnd cell_6t
Xbit_r15_c46 bl[46] br[46] wl[15] vdd gnd cell_6t
Xbit_r16_c46 bl[46] br[46] wl[16] vdd gnd cell_6t
Xbit_r17_c46 bl[46] br[46] wl[17] vdd gnd cell_6t
Xbit_r18_c46 bl[46] br[46] wl[18] vdd gnd cell_6t
Xbit_r19_c46 bl[46] br[46] wl[19] vdd gnd cell_6t
Xbit_r20_c46 bl[46] br[46] wl[20] vdd gnd cell_6t
Xbit_r21_c46 bl[46] br[46] wl[21] vdd gnd cell_6t
Xbit_r22_c46 bl[46] br[46] wl[22] vdd gnd cell_6t
Xbit_r23_c46 bl[46] br[46] wl[23] vdd gnd cell_6t
Xbit_r24_c46 bl[46] br[46] wl[24] vdd gnd cell_6t
Xbit_r25_c46 bl[46] br[46] wl[25] vdd gnd cell_6t
Xbit_r26_c46 bl[46] br[46] wl[26] vdd gnd cell_6t
Xbit_r27_c46 bl[46] br[46] wl[27] vdd gnd cell_6t
Xbit_r28_c46 bl[46] br[46] wl[28] vdd gnd cell_6t
Xbit_r29_c46 bl[46] br[46] wl[29] vdd gnd cell_6t
Xbit_r30_c46 bl[46] br[46] wl[30] vdd gnd cell_6t
Xbit_r31_c46 bl[46] br[46] wl[31] vdd gnd cell_6t
Xbit_r32_c46 bl[46] br[46] wl[32] vdd gnd cell_6t
Xbit_r33_c46 bl[46] br[46] wl[33] vdd gnd cell_6t
Xbit_r34_c46 bl[46] br[46] wl[34] vdd gnd cell_6t
Xbit_r35_c46 bl[46] br[46] wl[35] vdd gnd cell_6t
Xbit_r36_c46 bl[46] br[46] wl[36] vdd gnd cell_6t
Xbit_r37_c46 bl[46] br[46] wl[37] vdd gnd cell_6t
Xbit_r38_c46 bl[46] br[46] wl[38] vdd gnd cell_6t
Xbit_r39_c46 bl[46] br[46] wl[39] vdd gnd cell_6t
Xbit_r40_c46 bl[46] br[46] wl[40] vdd gnd cell_6t
Xbit_r41_c46 bl[46] br[46] wl[41] vdd gnd cell_6t
Xbit_r42_c46 bl[46] br[46] wl[42] vdd gnd cell_6t
Xbit_r43_c46 bl[46] br[46] wl[43] vdd gnd cell_6t
Xbit_r44_c46 bl[46] br[46] wl[44] vdd gnd cell_6t
Xbit_r45_c46 bl[46] br[46] wl[45] vdd gnd cell_6t
Xbit_r46_c46 bl[46] br[46] wl[46] vdd gnd cell_6t
Xbit_r47_c46 bl[46] br[46] wl[47] vdd gnd cell_6t
Xbit_r48_c46 bl[46] br[46] wl[48] vdd gnd cell_6t
Xbit_r49_c46 bl[46] br[46] wl[49] vdd gnd cell_6t
Xbit_r50_c46 bl[46] br[46] wl[50] vdd gnd cell_6t
Xbit_r51_c46 bl[46] br[46] wl[51] vdd gnd cell_6t
Xbit_r52_c46 bl[46] br[46] wl[52] vdd gnd cell_6t
Xbit_r53_c46 bl[46] br[46] wl[53] vdd gnd cell_6t
Xbit_r54_c46 bl[46] br[46] wl[54] vdd gnd cell_6t
Xbit_r55_c46 bl[46] br[46] wl[55] vdd gnd cell_6t
Xbit_r56_c46 bl[46] br[46] wl[56] vdd gnd cell_6t
Xbit_r57_c46 bl[46] br[46] wl[57] vdd gnd cell_6t
Xbit_r58_c46 bl[46] br[46] wl[58] vdd gnd cell_6t
Xbit_r59_c46 bl[46] br[46] wl[59] vdd gnd cell_6t
Xbit_r60_c46 bl[46] br[46] wl[60] vdd gnd cell_6t
Xbit_r61_c46 bl[46] br[46] wl[61] vdd gnd cell_6t
Xbit_r62_c46 bl[46] br[46] wl[62] vdd gnd cell_6t
Xbit_r63_c46 bl[46] br[46] wl[63] vdd gnd cell_6t
Xbit_r64_c46 bl[46] br[46] wl[64] vdd gnd cell_6t
Xbit_r65_c46 bl[46] br[46] wl[65] vdd gnd cell_6t
Xbit_r66_c46 bl[46] br[46] wl[66] vdd gnd cell_6t
Xbit_r67_c46 bl[46] br[46] wl[67] vdd gnd cell_6t
Xbit_r68_c46 bl[46] br[46] wl[68] vdd gnd cell_6t
Xbit_r69_c46 bl[46] br[46] wl[69] vdd gnd cell_6t
Xbit_r70_c46 bl[46] br[46] wl[70] vdd gnd cell_6t
Xbit_r71_c46 bl[46] br[46] wl[71] vdd gnd cell_6t
Xbit_r72_c46 bl[46] br[46] wl[72] vdd gnd cell_6t
Xbit_r73_c46 bl[46] br[46] wl[73] vdd gnd cell_6t
Xbit_r74_c46 bl[46] br[46] wl[74] vdd gnd cell_6t
Xbit_r75_c46 bl[46] br[46] wl[75] vdd gnd cell_6t
Xbit_r76_c46 bl[46] br[46] wl[76] vdd gnd cell_6t
Xbit_r77_c46 bl[46] br[46] wl[77] vdd gnd cell_6t
Xbit_r78_c46 bl[46] br[46] wl[78] vdd gnd cell_6t
Xbit_r79_c46 bl[46] br[46] wl[79] vdd gnd cell_6t
Xbit_r80_c46 bl[46] br[46] wl[80] vdd gnd cell_6t
Xbit_r81_c46 bl[46] br[46] wl[81] vdd gnd cell_6t
Xbit_r82_c46 bl[46] br[46] wl[82] vdd gnd cell_6t
Xbit_r83_c46 bl[46] br[46] wl[83] vdd gnd cell_6t
Xbit_r84_c46 bl[46] br[46] wl[84] vdd gnd cell_6t
Xbit_r85_c46 bl[46] br[46] wl[85] vdd gnd cell_6t
Xbit_r86_c46 bl[46] br[46] wl[86] vdd gnd cell_6t
Xbit_r87_c46 bl[46] br[46] wl[87] vdd gnd cell_6t
Xbit_r88_c46 bl[46] br[46] wl[88] vdd gnd cell_6t
Xbit_r89_c46 bl[46] br[46] wl[89] vdd gnd cell_6t
Xbit_r90_c46 bl[46] br[46] wl[90] vdd gnd cell_6t
Xbit_r91_c46 bl[46] br[46] wl[91] vdd gnd cell_6t
Xbit_r92_c46 bl[46] br[46] wl[92] vdd gnd cell_6t
Xbit_r93_c46 bl[46] br[46] wl[93] vdd gnd cell_6t
Xbit_r94_c46 bl[46] br[46] wl[94] vdd gnd cell_6t
Xbit_r95_c46 bl[46] br[46] wl[95] vdd gnd cell_6t
Xbit_r96_c46 bl[46] br[46] wl[96] vdd gnd cell_6t
Xbit_r97_c46 bl[46] br[46] wl[97] vdd gnd cell_6t
Xbit_r98_c46 bl[46] br[46] wl[98] vdd gnd cell_6t
Xbit_r99_c46 bl[46] br[46] wl[99] vdd gnd cell_6t
Xbit_r100_c46 bl[46] br[46] wl[100] vdd gnd cell_6t
Xbit_r101_c46 bl[46] br[46] wl[101] vdd gnd cell_6t
Xbit_r102_c46 bl[46] br[46] wl[102] vdd gnd cell_6t
Xbit_r103_c46 bl[46] br[46] wl[103] vdd gnd cell_6t
Xbit_r104_c46 bl[46] br[46] wl[104] vdd gnd cell_6t
Xbit_r105_c46 bl[46] br[46] wl[105] vdd gnd cell_6t
Xbit_r106_c46 bl[46] br[46] wl[106] vdd gnd cell_6t
Xbit_r107_c46 bl[46] br[46] wl[107] vdd gnd cell_6t
Xbit_r108_c46 bl[46] br[46] wl[108] vdd gnd cell_6t
Xbit_r109_c46 bl[46] br[46] wl[109] vdd gnd cell_6t
Xbit_r110_c46 bl[46] br[46] wl[110] vdd gnd cell_6t
Xbit_r111_c46 bl[46] br[46] wl[111] vdd gnd cell_6t
Xbit_r112_c46 bl[46] br[46] wl[112] vdd gnd cell_6t
Xbit_r113_c46 bl[46] br[46] wl[113] vdd gnd cell_6t
Xbit_r114_c46 bl[46] br[46] wl[114] vdd gnd cell_6t
Xbit_r115_c46 bl[46] br[46] wl[115] vdd gnd cell_6t
Xbit_r116_c46 bl[46] br[46] wl[116] vdd gnd cell_6t
Xbit_r117_c46 bl[46] br[46] wl[117] vdd gnd cell_6t
Xbit_r118_c46 bl[46] br[46] wl[118] vdd gnd cell_6t
Xbit_r119_c46 bl[46] br[46] wl[119] vdd gnd cell_6t
Xbit_r120_c46 bl[46] br[46] wl[120] vdd gnd cell_6t
Xbit_r121_c46 bl[46] br[46] wl[121] vdd gnd cell_6t
Xbit_r122_c46 bl[46] br[46] wl[122] vdd gnd cell_6t
Xbit_r123_c46 bl[46] br[46] wl[123] vdd gnd cell_6t
Xbit_r124_c46 bl[46] br[46] wl[124] vdd gnd cell_6t
Xbit_r125_c46 bl[46] br[46] wl[125] vdd gnd cell_6t
Xbit_r126_c46 bl[46] br[46] wl[126] vdd gnd cell_6t
Xbit_r127_c46 bl[46] br[46] wl[127] vdd gnd cell_6t
Xbit_r0_c47 bl[47] br[47] wl[0] vdd gnd cell_6t
Xbit_r1_c47 bl[47] br[47] wl[1] vdd gnd cell_6t
Xbit_r2_c47 bl[47] br[47] wl[2] vdd gnd cell_6t
Xbit_r3_c47 bl[47] br[47] wl[3] vdd gnd cell_6t
Xbit_r4_c47 bl[47] br[47] wl[4] vdd gnd cell_6t
Xbit_r5_c47 bl[47] br[47] wl[5] vdd gnd cell_6t
Xbit_r6_c47 bl[47] br[47] wl[6] vdd gnd cell_6t
Xbit_r7_c47 bl[47] br[47] wl[7] vdd gnd cell_6t
Xbit_r8_c47 bl[47] br[47] wl[8] vdd gnd cell_6t
Xbit_r9_c47 bl[47] br[47] wl[9] vdd gnd cell_6t
Xbit_r10_c47 bl[47] br[47] wl[10] vdd gnd cell_6t
Xbit_r11_c47 bl[47] br[47] wl[11] vdd gnd cell_6t
Xbit_r12_c47 bl[47] br[47] wl[12] vdd gnd cell_6t
Xbit_r13_c47 bl[47] br[47] wl[13] vdd gnd cell_6t
Xbit_r14_c47 bl[47] br[47] wl[14] vdd gnd cell_6t
Xbit_r15_c47 bl[47] br[47] wl[15] vdd gnd cell_6t
Xbit_r16_c47 bl[47] br[47] wl[16] vdd gnd cell_6t
Xbit_r17_c47 bl[47] br[47] wl[17] vdd gnd cell_6t
Xbit_r18_c47 bl[47] br[47] wl[18] vdd gnd cell_6t
Xbit_r19_c47 bl[47] br[47] wl[19] vdd gnd cell_6t
Xbit_r20_c47 bl[47] br[47] wl[20] vdd gnd cell_6t
Xbit_r21_c47 bl[47] br[47] wl[21] vdd gnd cell_6t
Xbit_r22_c47 bl[47] br[47] wl[22] vdd gnd cell_6t
Xbit_r23_c47 bl[47] br[47] wl[23] vdd gnd cell_6t
Xbit_r24_c47 bl[47] br[47] wl[24] vdd gnd cell_6t
Xbit_r25_c47 bl[47] br[47] wl[25] vdd gnd cell_6t
Xbit_r26_c47 bl[47] br[47] wl[26] vdd gnd cell_6t
Xbit_r27_c47 bl[47] br[47] wl[27] vdd gnd cell_6t
Xbit_r28_c47 bl[47] br[47] wl[28] vdd gnd cell_6t
Xbit_r29_c47 bl[47] br[47] wl[29] vdd gnd cell_6t
Xbit_r30_c47 bl[47] br[47] wl[30] vdd gnd cell_6t
Xbit_r31_c47 bl[47] br[47] wl[31] vdd gnd cell_6t
Xbit_r32_c47 bl[47] br[47] wl[32] vdd gnd cell_6t
Xbit_r33_c47 bl[47] br[47] wl[33] vdd gnd cell_6t
Xbit_r34_c47 bl[47] br[47] wl[34] vdd gnd cell_6t
Xbit_r35_c47 bl[47] br[47] wl[35] vdd gnd cell_6t
Xbit_r36_c47 bl[47] br[47] wl[36] vdd gnd cell_6t
Xbit_r37_c47 bl[47] br[47] wl[37] vdd gnd cell_6t
Xbit_r38_c47 bl[47] br[47] wl[38] vdd gnd cell_6t
Xbit_r39_c47 bl[47] br[47] wl[39] vdd gnd cell_6t
Xbit_r40_c47 bl[47] br[47] wl[40] vdd gnd cell_6t
Xbit_r41_c47 bl[47] br[47] wl[41] vdd gnd cell_6t
Xbit_r42_c47 bl[47] br[47] wl[42] vdd gnd cell_6t
Xbit_r43_c47 bl[47] br[47] wl[43] vdd gnd cell_6t
Xbit_r44_c47 bl[47] br[47] wl[44] vdd gnd cell_6t
Xbit_r45_c47 bl[47] br[47] wl[45] vdd gnd cell_6t
Xbit_r46_c47 bl[47] br[47] wl[46] vdd gnd cell_6t
Xbit_r47_c47 bl[47] br[47] wl[47] vdd gnd cell_6t
Xbit_r48_c47 bl[47] br[47] wl[48] vdd gnd cell_6t
Xbit_r49_c47 bl[47] br[47] wl[49] vdd gnd cell_6t
Xbit_r50_c47 bl[47] br[47] wl[50] vdd gnd cell_6t
Xbit_r51_c47 bl[47] br[47] wl[51] vdd gnd cell_6t
Xbit_r52_c47 bl[47] br[47] wl[52] vdd gnd cell_6t
Xbit_r53_c47 bl[47] br[47] wl[53] vdd gnd cell_6t
Xbit_r54_c47 bl[47] br[47] wl[54] vdd gnd cell_6t
Xbit_r55_c47 bl[47] br[47] wl[55] vdd gnd cell_6t
Xbit_r56_c47 bl[47] br[47] wl[56] vdd gnd cell_6t
Xbit_r57_c47 bl[47] br[47] wl[57] vdd gnd cell_6t
Xbit_r58_c47 bl[47] br[47] wl[58] vdd gnd cell_6t
Xbit_r59_c47 bl[47] br[47] wl[59] vdd gnd cell_6t
Xbit_r60_c47 bl[47] br[47] wl[60] vdd gnd cell_6t
Xbit_r61_c47 bl[47] br[47] wl[61] vdd gnd cell_6t
Xbit_r62_c47 bl[47] br[47] wl[62] vdd gnd cell_6t
Xbit_r63_c47 bl[47] br[47] wl[63] vdd gnd cell_6t
Xbit_r64_c47 bl[47] br[47] wl[64] vdd gnd cell_6t
Xbit_r65_c47 bl[47] br[47] wl[65] vdd gnd cell_6t
Xbit_r66_c47 bl[47] br[47] wl[66] vdd gnd cell_6t
Xbit_r67_c47 bl[47] br[47] wl[67] vdd gnd cell_6t
Xbit_r68_c47 bl[47] br[47] wl[68] vdd gnd cell_6t
Xbit_r69_c47 bl[47] br[47] wl[69] vdd gnd cell_6t
Xbit_r70_c47 bl[47] br[47] wl[70] vdd gnd cell_6t
Xbit_r71_c47 bl[47] br[47] wl[71] vdd gnd cell_6t
Xbit_r72_c47 bl[47] br[47] wl[72] vdd gnd cell_6t
Xbit_r73_c47 bl[47] br[47] wl[73] vdd gnd cell_6t
Xbit_r74_c47 bl[47] br[47] wl[74] vdd gnd cell_6t
Xbit_r75_c47 bl[47] br[47] wl[75] vdd gnd cell_6t
Xbit_r76_c47 bl[47] br[47] wl[76] vdd gnd cell_6t
Xbit_r77_c47 bl[47] br[47] wl[77] vdd gnd cell_6t
Xbit_r78_c47 bl[47] br[47] wl[78] vdd gnd cell_6t
Xbit_r79_c47 bl[47] br[47] wl[79] vdd gnd cell_6t
Xbit_r80_c47 bl[47] br[47] wl[80] vdd gnd cell_6t
Xbit_r81_c47 bl[47] br[47] wl[81] vdd gnd cell_6t
Xbit_r82_c47 bl[47] br[47] wl[82] vdd gnd cell_6t
Xbit_r83_c47 bl[47] br[47] wl[83] vdd gnd cell_6t
Xbit_r84_c47 bl[47] br[47] wl[84] vdd gnd cell_6t
Xbit_r85_c47 bl[47] br[47] wl[85] vdd gnd cell_6t
Xbit_r86_c47 bl[47] br[47] wl[86] vdd gnd cell_6t
Xbit_r87_c47 bl[47] br[47] wl[87] vdd gnd cell_6t
Xbit_r88_c47 bl[47] br[47] wl[88] vdd gnd cell_6t
Xbit_r89_c47 bl[47] br[47] wl[89] vdd gnd cell_6t
Xbit_r90_c47 bl[47] br[47] wl[90] vdd gnd cell_6t
Xbit_r91_c47 bl[47] br[47] wl[91] vdd gnd cell_6t
Xbit_r92_c47 bl[47] br[47] wl[92] vdd gnd cell_6t
Xbit_r93_c47 bl[47] br[47] wl[93] vdd gnd cell_6t
Xbit_r94_c47 bl[47] br[47] wl[94] vdd gnd cell_6t
Xbit_r95_c47 bl[47] br[47] wl[95] vdd gnd cell_6t
Xbit_r96_c47 bl[47] br[47] wl[96] vdd gnd cell_6t
Xbit_r97_c47 bl[47] br[47] wl[97] vdd gnd cell_6t
Xbit_r98_c47 bl[47] br[47] wl[98] vdd gnd cell_6t
Xbit_r99_c47 bl[47] br[47] wl[99] vdd gnd cell_6t
Xbit_r100_c47 bl[47] br[47] wl[100] vdd gnd cell_6t
Xbit_r101_c47 bl[47] br[47] wl[101] vdd gnd cell_6t
Xbit_r102_c47 bl[47] br[47] wl[102] vdd gnd cell_6t
Xbit_r103_c47 bl[47] br[47] wl[103] vdd gnd cell_6t
Xbit_r104_c47 bl[47] br[47] wl[104] vdd gnd cell_6t
Xbit_r105_c47 bl[47] br[47] wl[105] vdd gnd cell_6t
Xbit_r106_c47 bl[47] br[47] wl[106] vdd gnd cell_6t
Xbit_r107_c47 bl[47] br[47] wl[107] vdd gnd cell_6t
Xbit_r108_c47 bl[47] br[47] wl[108] vdd gnd cell_6t
Xbit_r109_c47 bl[47] br[47] wl[109] vdd gnd cell_6t
Xbit_r110_c47 bl[47] br[47] wl[110] vdd gnd cell_6t
Xbit_r111_c47 bl[47] br[47] wl[111] vdd gnd cell_6t
Xbit_r112_c47 bl[47] br[47] wl[112] vdd gnd cell_6t
Xbit_r113_c47 bl[47] br[47] wl[113] vdd gnd cell_6t
Xbit_r114_c47 bl[47] br[47] wl[114] vdd gnd cell_6t
Xbit_r115_c47 bl[47] br[47] wl[115] vdd gnd cell_6t
Xbit_r116_c47 bl[47] br[47] wl[116] vdd gnd cell_6t
Xbit_r117_c47 bl[47] br[47] wl[117] vdd gnd cell_6t
Xbit_r118_c47 bl[47] br[47] wl[118] vdd gnd cell_6t
Xbit_r119_c47 bl[47] br[47] wl[119] vdd gnd cell_6t
Xbit_r120_c47 bl[47] br[47] wl[120] vdd gnd cell_6t
Xbit_r121_c47 bl[47] br[47] wl[121] vdd gnd cell_6t
Xbit_r122_c47 bl[47] br[47] wl[122] vdd gnd cell_6t
Xbit_r123_c47 bl[47] br[47] wl[123] vdd gnd cell_6t
Xbit_r124_c47 bl[47] br[47] wl[124] vdd gnd cell_6t
Xbit_r125_c47 bl[47] br[47] wl[125] vdd gnd cell_6t
Xbit_r126_c47 bl[47] br[47] wl[126] vdd gnd cell_6t
Xbit_r127_c47 bl[47] br[47] wl[127] vdd gnd cell_6t
Xbit_r0_c48 bl[48] br[48] wl[0] vdd gnd cell_6t
Xbit_r1_c48 bl[48] br[48] wl[1] vdd gnd cell_6t
Xbit_r2_c48 bl[48] br[48] wl[2] vdd gnd cell_6t
Xbit_r3_c48 bl[48] br[48] wl[3] vdd gnd cell_6t
Xbit_r4_c48 bl[48] br[48] wl[4] vdd gnd cell_6t
Xbit_r5_c48 bl[48] br[48] wl[5] vdd gnd cell_6t
Xbit_r6_c48 bl[48] br[48] wl[6] vdd gnd cell_6t
Xbit_r7_c48 bl[48] br[48] wl[7] vdd gnd cell_6t
Xbit_r8_c48 bl[48] br[48] wl[8] vdd gnd cell_6t
Xbit_r9_c48 bl[48] br[48] wl[9] vdd gnd cell_6t
Xbit_r10_c48 bl[48] br[48] wl[10] vdd gnd cell_6t
Xbit_r11_c48 bl[48] br[48] wl[11] vdd gnd cell_6t
Xbit_r12_c48 bl[48] br[48] wl[12] vdd gnd cell_6t
Xbit_r13_c48 bl[48] br[48] wl[13] vdd gnd cell_6t
Xbit_r14_c48 bl[48] br[48] wl[14] vdd gnd cell_6t
Xbit_r15_c48 bl[48] br[48] wl[15] vdd gnd cell_6t
Xbit_r16_c48 bl[48] br[48] wl[16] vdd gnd cell_6t
Xbit_r17_c48 bl[48] br[48] wl[17] vdd gnd cell_6t
Xbit_r18_c48 bl[48] br[48] wl[18] vdd gnd cell_6t
Xbit_r19_c48 bl[48] br[48] wl[19] vdd gnd cell_6t
Xbit_r20_c48 bl[48] br[48] wl[20] vdd gnd cell_6t
Xbit_r21_c48 bl[48] br[48] wl[21] vdd gnd cell_6t
Xbit_r22_c48 bl[48] br[48] wl[22] vdd gnd cell_6t
Xbit_r23_c48 bl[48] br[48] wl[23] vdd gnd cell_6t
Xbit_r24_c48 bl[48] br[48] wl[24] vdd gnd cell_6t
Xbit_r25_c48 bl[48] br[48] wl[25] vdd gnd cell_6t
Xbit_r26_c48 bl[48] br[48] wl[26] vdd gnd cell_6t
Xbit_r27_c48 bl[48] br[48] wl[27] vdd gnd cell_6t
Xbit_r28_c48 bl[48] br[48] wl[28] vdd gnd cell_6t
Xbit_r29_c48 bl[48] br[48] wl[29] vdd gnd cell_6t
Xbit_r30_c48 bl[48] br[48] wl[30] vdd gnd cell_6t
Xbit_r31_c48 bl[48] br[48] wl[31] vdd gnd cell_6t
Xbit_r32_c48 bl[48] br[48] wl[32] vdd gnd cell_6t
Xbit_r33_c48 bl[48] br[48] wl[33] vdd gnd cell_6t
Xbit_r34_c48 bl[48] br[48] wl[34] vdd gnd cell_6t
Xbit_r35_c48 bl[48] br[48] wl[35] vdd gnd cell_6t
Xbit_r36_c48 bl[48] br[48] wl[36] vdd gnd cell_6t
Xbit_r37_c48 bl[48] br[48] wl[37] vdd gnd cell_6t
Xbit_r38_c48 bl[48] br[48] wl[38] vdd gnd cell_6t
Xbit_r39_c48 bl[48] br[48] wl[39] vdd gnd cell_6t
Xbit_r40_c48 bl[48] br[48] wl[40] vdd gnd cell_6t
Xbit_r41_c48 bl[48] br[48] wl[41] vdd gnd cell_6t
Xbit_r42_c48 bl[48] br[48] wl[42] vdd gnd cell_6t
Xbit_r43_c48 bl[48] br[48] wl[43] vdd gnd cell_6t
Xbit_r44_c48 bl[48] br[48] wl[44] vdd gnd cell_6t
Xbit_r45_c48 bl[48] br[48] wl[45] vdd gnd cell_6t
Xbit_r46_c48 bl[48] br[48] wl[46] vdd gnd cell_6t
Xbit_r47_c48 bl[48] br[48] wl[47] vdd gnd cell_6t
Xbit_r48_c48 bl[48] br[48] wl[48] vdd gnd cell_6t
Xbit_r49_c48 bl[48] br[48] wl[49] vdd gnd cell_6t
Xbit_r50_c48 bl[48] br[48] wl[50] vdd gnd cell_6t
Xbit_r51_c48 bl[48] br[48] wl[51] vdd gnd cell_6t
Xbit_r52_c48 bl[48] br[48] wl[52] vdd gnd cell_6t
Xbit_r53_c48 bl[48] br[48] wl[53] vdd gnd cell_6t
Xbit_r54_c48 bl[48] br[48] wl[54] vdd gnd cell_6t
Xbit_r55_c48 bl[48] br[48] wl[55] vdd gnd cell_6t
Xbit_r56_c48 bl[48] br[48] wl[56] vdd gnd cell_6t
Xbit_r57_c48 bl[48] br[48] wl[57] vdd gnd cell_6t
Xbit_r58_c48 bl[48] br[48] wl[58] vdd gnd cell_6t
Xbit_r59_c48 bl[48] br[48] wl[59] vdd gnd cell_6t
Xbit_r60_c48 bl[48] br[48] wl[60] vdd gnd cell_6t
Xbit_r61_c48 bl[48] br[48] wl[61] vdd gnd cell_6t
Xbit_r62_c48 bl[48] br[48] wl[62] vdd gnd cell_6t
Xbit_r63_c48 bl[48] br[48] wl[63] vdd gnd cell_6t
Xbit_r64_c48 bl[48] br[48] wl[64] vdd gnd cell_6t
Xbit_r65_c48 bl[48] br[48] wl[65] vdd gnd cell_6t
Xbit_r66_c48 bl[48] br[48] wl[66] vdd gnd cell_6t
Xbit_r67_c48 bl[48] br[48] wl[67] vdd gnd cell_6t
Xbit_r68_c48 bl[48] br[48] wl[68] vdd gnd cell_6t
Xbit_r69_c48 bl[48] br[48] wl[69] vdd gnd cell_6t
Xbit_r70_c48 bl[48] br[48] wl[70] vdd gnd cell_6t
Xbit_r71_c48 bl[48] br[48] wl[71] vdd gnd cell_6t
Xbit_r72_c48 bl[48] br[48] wl[72] vdd gnd cell_6t
Xbit_r73_c48 bl[48] br[48] wl[73] vdd gnd cell_6t
Xbit_r74_c48 bl[48] br[48] wl[74] vdd gnd cell_6t
Xbit_r75_c48 bl[48] br[48] wl[75] vdd gnd cell_6t
Xbit_r76_c48 bl[48] br[48] wl[76] vdd gnd cell_6t
Xbit_r77_c48 bl[48] br[48] wl[77] vdd gnd cell_6t
Xbit_r78_c48 bl[48] br[48] wl[78] vdd gnd cell_6t
Xbit_r79_c48 bl[48] br[48] wl[79] vdd gnd cell_6t
Xbit_r80_c48 bl[48] br[48] wl[80] vdd gnd cell_6t
Xbit_r81_c48 bl[48] br[48] wl[81] vdd gnd cell_6t
Xbit_r82_c48 bl[48] br[48] wl[82] vdd gnd cell_6t
Xbit_r83_c48 bl[48] br[48] wl[83] vdd gnd cell_6t
Xbit_r84_c48 bl[48] br[48] wl[84] vdd gnd cell_6t
Xbit_r85_c48 bl[48] br[48] wl[85] vdd gnd cell_6t
Xbit_r86_c48 bl[48] br[48] wl[86] vdd gnd cell_6t
Xbit_r87_c48 bl[48] br[48] wl[87] vdd gnd cell_6t
Xbit_r88_c48 bl[48] br[48] wl[88] vdd gnd cell_6t
Xbit_r89_c48 bl[48] br[48] wl[89] vdd gnd cell_6t
Xbit_r90_c48 bl[48] br[48] wl[90] vdd gnd cell_6t
Xbit_r91_c48 bl[48] br[48] wl[91] vdd gnd cell_6t
Xbit_r92_c48 bl[48] br[48] wl[92] vdd gnd cell_6t
Xbit_r93_c48 bl[48] br[48] wl[93] vdd gnd cell_6t
Xbit_r94_c48 bl[48] br[48] wl[94] vdd gnd cell_6t
Xbit_r95_c48 bl[48] br[48] wl[95] vdd gnd cell_6t
Xbit_r96_c48 bl[48] br[48] wl[96] vdd gnd cell_6t
Xbit_r97_c48 bl[48] br[48] wl[97] vdd gnd cell_6t
Xbit_r98_c48 bl[48] br[48] wl[98] vdd gnd cell_6t
Xbit_r99_c48 bl[48] br[48] wl[99] vdd gnd cell_6t
Xbit_r100_c48 bl[48] br[48] wl[100] vdd gnd cell_6t
Xbit_r101_c48 bl[48] br[48] wl[101] vdd gnd cell_6t
Xbit_r102_c48 bl[48] br[48] wl[102] vdd gnd cell_6t
Xbit_r103_c48 bl[48] br[48] wl[103] vdd gnd cell_6t
Xbit_r104_c48 bl[48] br[48] wl[104] vdd gnd cell_6t
Xbit_r105_c48 bl[48] br[48] wl[105] vdd gnd cell_6t
Xbit_r106_c48 bl[48] br[48] wl[106] vdd gnd cell_6t
Xbit_r107_c48 bl[48] br[48] wl[107] vdd gnd cell_6t
Xbit_r108_c48 bl[48] br[48] wl[108] vdd gnd cell_6t
Xbit_r109_c48 bl[48] br[48] wl[109] vdd gnd cell_6t
Xbit_r110_c48 bl[48] br[48] wl[110] vdd gnd cell_6t
Xbit_r111_c48 bl[48] br[48] wl[111] vdd gnd cell_6t
Xbit_r112_c48 bl[48] br[48] wl[112] vdd gnd cell_6t
Xbit_r113_c48 bl[48] br[48] wl[113] vdd gnd cell_6t
Xbit_r114_c48 bl[48] br[48] wl[114] vdd gnd cell_6t
Xbit_r115_c48 bl[48] br[48] wl[115] vdd gnd cell_6t
Xbit_r116_c48 bl[48] br[48] wl[116] vdd gnd cell_6t
Xbit_r117_c48 bl[48] br[48] wl[117] vdd gnd cell_6t
Xbit_r118_c48 bl[48] br[48] wl[118] vdd gnd cell_6t
Xbit_r119_c48 bl[48] br[48] wl[119] vdd gnd cell_6t
Xbit_r120_c48 bl[48] br[48] wl[120] vdd gnd cell_6t
Xbit_r121_c48 bl[48] br[48] wl[121] vdd gnd cell_6t
Xbit_r122_c48 bl[48] br[48] wl[122] vdd gnd cell_6t
Xbit_r123_c48 bl[48] br[48] wl[123] vdd gnd cell_6t
Xbit_r124_c48 bl[48] br[48] wl[124] vdd gnd cell_6t
Xbit_r125_c48 bl[48] br[48] wl[125] vdd gnd cell_6t
Xbit_r126_c48 bl[48] br[48] wl[126] vdd gnd cell_6t
Xbit_r127_c48 bl[48] br[48] wl[127] vdd gnd cell_6t
Xbit_r0_c49 bl[49] br[49] wl[0] vdd gnd cell_6t
Xbit_r1_c49 bl[49] br[49] wl[1] vdd gnd cell_6t
Xbit_r2_c49 bl[49] br[49] wl[2] vdd gnd cell_6t
Xbit_r3_c49 bl[49] br[49] wl[3] vdd gnd cell_6t
Xbit_r4_c49 bl[49] br[49] wl[4] vdd gnd cell_6t
Xbit_r5_c49 bl[49] br[49] wl[5] vdd gnd cell_6t
Xbit_r6_c49 bl[49] br[49] wl[6] vdd gnd cell_6t
Xbit_r7_c49 bl[49] br[49] wl[7] vdd gnd cell_6t
Xbit_r8_c49 bl[49] br[49] wl[8] vdd gnd cell_6t
Xbit_r9_c49 bl[49] br[49] wl[9] vdd gnd cell_6t
Xbit_r10_c49 bl[49] br[49] wl[10] vdd gnd cell_6t
Xbit_r11_c49 bl[49] br[49] wl[11] vdd gnd cell_6t
Xbit_r12_c49 bl[49] br[49] wl[12] vdd gnd cell_6t
Xbit_r13_c49 bl[49] br[49] wl[13] vdd gnd cell_6t
Xbit_r14_c49 bl[49] br[49] wl[14] vdd gnd cell_6t
Xbit_r15_c49 bl[49] br[49] wl[15] vdd gnd cell_6t
Xbit_r16_c49 bl[49] br[49] wl[16] vdd gnd cell_6t
Xbit_r17_c49 bl[49] br[49] wl[17] vdd gnd cell_6t
Xbit_r18_c49 bl[49] br[49] wl[18] vdd gnd cell_6t
Xbit_r19_c49 bl[49] br[49] wl[19] vdd gnd cell_6t
Xbit_r20_c49 bl[49] br[49] wl[20] vdd gnd cell_6t
Xbit_r21_c49 bl[49] br[49] wl[21] vdd gnd cell_6t
Xbit_r22_c49 bl[49] br[49] wl[22] vdd gnd cell_6t
Xbit_r23_c49 bl[49] br[49] wl[23] vdd gnd cell_6t
Xbit_r24_c49 bl[49] br[49] wl[24] vdd gnd cell_6t
Xbit_r25_c49 bl[49] br[49] wl[25] vdd gnd cell_6t
Xbit_r26_c49 bl[49] br[49] wl[26] vdd gnd cell_6t
Xbit_r27_c49 bl[49] br[49] wl[27] vdd gnd cell_6t
Xbit_r28_c49 bl[49] br[49] wl[28] vdd gnd cell_6t
Xbit_r29_c49 bl[49] br[49] wl[29] vdd gnd cell_6t
Xbit_r30_c49 bl[49] br[49] wl[30] vdd gnd cell_6t
Xbit_r31_c49 bl[49] br[49] wl[31] vdd gnd cell_6t
Xbit_r32_c49 bl[49] br[49] wl[32] vdd gnd cell_6t
Xbit_r33_c49 bl[49] br[49] wl[33] vdd gnd cell_6t
Xbit_r34_c49 bl[49] br[49] wl[34] vdd gnd cell_6t
Xbit_r35_c49 bl[49] br[49] wl[35] vdd gnd cell_6t
Xbit_r36_c49 bl[49] br[49] wl[36] vdd gnd cell_6t
Xbit_r37_c49 bl[49] br[49] wl[37] vdd gnd cell_6t
Xbit_r38_c49 bl[49] br[49] wl[38] vdd gnd cell_6t
Xbit_r39_c49 bl[49] br[49] wl[39] vdd gnd cell_6t
Xbit_r40_c49 bl[49] br[49] wl[40] vdd gnd cell_6t
Xbit_r41_c49 bl[49] br[49] wl[41] vdd gnd cell_6t
Xbit_r42_c49 bl[49] br[49] wl[42] vdd gnd cell_6t
Xbit_r43_c49 bl[49] br[49] wl[43] vdd gnd cell_6t
Xbit_r44_c49 bl[49] br[49] wl[44] vdd gnd cell_6t
Xbit_r45_c49 bl[49] br[49] wl[45] vdd gnd cell_6t
Xbit_r46_c49 bl[49] br[49] wl[46] vdd gnd cell_6t
Xbit_r47_c49 bl[49] br[49] wl[47] vdd gnd cell_6t
Xbit_r48_c49 bl[49] br[49] wl[48] vdd gnd cell_6t
Xbit_r49_c49 bl[49] br[49] wl[49] vdd gnd cell_6t
Xbit_r50_c49 bl[49] br[49] wl[50] vdd gnd cell_6t
Xbit_r51_c49 bl[49] br[49] wl[51] vdd gnd cell_6t
Xbit_r52_c49 bl[49] br[49] wl[52] vdd gnd cell_6t
Xbit_r53_c49 bl[49] br[49] wl[53] vdd gnd cell_6t
Xbit_r54_c49 bl[49] br[49] wl[54] vdd gnd cell_6t
Xbit_r55_c49 bl[49] br[49] wl[55] vdd gnd cell_6t
Xbit_r56_c49 bl[49] br[49] wl[56] vdd gnd cell_6t
Xbit_r57_c49 bl[49] br[49] wl[57] vdd gnd cell_6t
Xbit_r58_c49 bl[49] br[49] wl[58] vdd gnd cell_6t
Xbit_r59_c49 bl[49] br[49] wl[59] vdd gnd cell_6t
Xbit_r60_c49 bl[49] br[49] wl[60] vdd gnd cell_6t
Xbit_r61_c49 bl[49] br[49] wl[61] vdd gnd cell_6t
Xbit_r62_c49 bl[49] br[49] wl[62] vdd gnd cell_6t
Xbit_r63_c49 bl[49] br[49] wl[63] vdd gnd cell_6t
Xbit_r64_c49 bl[49] br[49] wl[64] vdd gnd cell_6t
Xbit_r65_c49 bl[49] br[49] wl[65] vdd gnd cell_6t
Xbit_r66_c49 bl[49] br[49] wl[66] vdd gnd cell_6t
Xbit_r67_c49 bl[49] br[49] wl[67] vdd gnd cell_6t
Xbit_r68_c49 bl[49] br[49] wl[68] vdd gnd cell_6t
Xbit_r69_c49 bl[49] br[49] wl[69] vdd gnd cell_6t
Xbit_r70_c49 bl[49] br[49] wl[70] vdd gnd cell_6t
Xbit_r71_c49 bl[49] br[49] wl[71] vdd gnd cell_6t
Xbit_r72_c49 bl[49] br[49] wl[72] vdd gnd cell_6t
Xbit_r73_c49 bl[49] br[49] wl[73] vdd gnd cell_6t
Xbit_r74_c49 bl[49] br[49] wl[74] vdd gnd cell_6t
Xbit_r75_c49 bl[49] br[49] wl[75] vdd gnd cell_6t
Xbit_r76_c49 bl[49] br[49] wl[76] vdd gnd cell_6t
Xbit_r77_c49 bl[49] br[49] wl[77] vdd gnd cell_6t
Xbit_r78_c49 bl[49] br[49] wl[78] vdd gnd cell_6t
Xbit_r79_c49 bl[49] br[49] wl[79] vdd gnd cell_6t
Xbit_r80_c49 bl[49] br[49] wl[80] vdd gnd cell_6t
Xbit_r81_c49 bl[49] br[49] wl[81] vdd gnd cell_6t
Xbit_r82_c49 bl[49] br[49] wl[82] vdd gnd cell_6t
Xbit_r83_c49 bl[49] br[49] wl[83] vdd gnd cell_6t
Xbit_r84_c49 bl[49] br[49] wl[84] vdd gnd cell_6t
Xbit_r85_c49 bl[49] br[49] wl[85] vdd gnd cell_6t
Xbit_r86_c49 bl[49] br[49] wl[86] vdd gnd cell_6t
Xbit_r87_c49 bl[49] br[49] wl[87] vdd gnd cell_6t
Xbit_r88_c49 bl[49] br[49] wl[88] vdd gnd cell_6t
Xbit_r89_c49 bl[49] br[49] wl[89] vdd gnd cell_6t
Xbit_r90_c49 bl[49] br[49] wl[90] vdd gnd cell_6t
Xbit_r91_c49 bl[49] br[49] wl[91] vdd gnd cell_6t
Xbit_r92_c49 bl[49] br[49] wl[92] vdd gnd cell_6t
Xbit_r93_c49 bl[49] br[49] wl[93] vdd gnd cell_6t
Xbit_r94_c49 bl[49] br[49] wl[94] vdd gnd cell_6t
Xbit_r95_c49 bl[49] br[49] wl[95] vdd gnd cell_6t
Xbit_r96_c49 bl[49] br[49] wl[96] vdd gnd cell_6t
Xbit_r97_c49 bl[49] br[49] wl[97] vdd gnd cell_6t
Xbit_r98_c49 bl[49] br[49] wl[98] vdd gnd cell_6t
Xbit_r99_c49 bl[49] br[49] wl[99] vdd gnd cell_6t
Xbit_r100_c49 bl[49] br[49] wl[100] vdd gnd cell_6t
Xbit_r101_c49 bl[49] br[49] wl[101] vdd gnd cell_6t
Xbit_r102_c49 bl[49] br[49] wl[102] vdd gnd cell_6t
Xbit_r103_c49 bl[49] br[49] wl[103] vdd gnd cell_6t
Xbit_r104_c49 bl[49] br[49] wl[104] vdd gnd cell_6t
Xbit_r105_c49 bl[49] br[49] wl[105] vdd gnd cell_6t
Xbit_r106_c49 bl[49] br[49] wl[106] vdd gnd cell_6t
Xbit_r107_c49 bl[49] br[49] wl[107] vdd gnd cell_6t
Xbit_r108_c49 bl[49] br[49] wl[108] vdd gnd cell_6t
Xbit_r109_c49 bl[49] br[49] wl[109] vdd gnd cell_6t
Xbit_r110_c49 bl[49] br[49] wl[110] vdd gnd cell_6t
Xbit_r111_c49 bl[49] br[49] wl[111] vdd gnd cell_6t
Xbit_r112_c49 bl[49] br[49] wl[112] vdd gnd cell_6t
Xbit_r113_c49 bl[49] br[49] wl[113] vdd gnd cell_6t
Xbit_r114_c49 bl[49] br[49] wl[114] vdd gnd cell_6t
Xbit_r115_c49 bl[49] br[49] wl[115] vdd gnd cell_6t
Xbit_r116_c49 bl[49] br[49] wl[116] vdd gnd cell_6t
Xbit_r117_c49 bl[49] br[49] wl[117] vdd gnd cell_6t
Xbit_r118_c49 bl[49] br[49] wl[118] vdd gnd cell_6t
Xbit_r119_c49 bl[49] br[49] wl[119] vdd gnd cell_6t
Xbit_r120_c49 bl[49] br[49] wl[120] vdd gnd cell_6t
Xbit_r121_c49 bl[49] br[49] wl[121] vdd gnd cell_6t
Xbit_r122_c49 bl[49] br[49] wl[122] vdd gnd cell_6t
Xbit_r123_c49 bl[49] br[49] wl[123] vdd gnd cell_6t
Xbit_r124_c49 bl[49] br[49] wl[124] vdd gnd cell_6t
Xbit_r125_c49 bl[49] br[49] wl[125] vdd gnd cell_6t
Xbit_r126_c49 bl[49] br[49] wl[126] vdd gnd cell_6t
Xbit_r127_c49 bl[49] br[49] wl[127] vdd gnd cell_6t
Xbit_r0_c50 bl[50] br[50] wl[0] vdd gnd cell_6t
Xbit_r1_c50 bl[50] br[50] wl[1] vdd gnd cell_6t
Xbit_r2_c50 bl[50] br[50] wl[2] vdd gnd cell_6t
Xbit_r3_c50 bl[50] br[50] wl[3] vdd gnd cell_6t
Xbit_r4_c50 bl[50] br[50] wl[4] vdd gnd cell_6t
Xbit_r5_c50 bl[50] br[50] wl[5] vdd gnd cell_6t
Xbit_r6_c50 bl[50] br[50] wl[6] vdd gnd cell_6t
Xbit_r7_c50 bl[50] br[50] wl[7] vdd gnd cell_6t
Xbit_r8_c50 bl[50] br[50] wl[8] vdd gnd cell_6t
Xbit_r9_c50 bl[50] br[50] wl[9] vdd gnd cell_6t
Xbit_r10_c50 bl[50] br[50] wl[10] vdd gnd cell_6t
Xbit_r11_c50 bl[50] br[50] wl[11] vdd gnd cell_6t
Xbit_r12_c50 bl[50] br[50] wl[12] vdd gnd cell_6t
Xbit_r13_c50 bl[50] br[50] wl[13] vdd gnd cell_6t
Xbit_r14_c50 bl[50] br[50] wl[14] vdd gnd cell_6t
Xbit_r15_c50 bl[50] br[50] wl[15] vdd gnd cell_6t
Xbit_r16_c50 bl[50] br[50] wl[16] vdd gnd cell_6t
Xbit_r17_c50 bl[50] br[50] wl[17] vdd gnd cell_6t
Xbit_r18_c50 bl[50] br[50] wl[18] vdd gnd cell_6t
Xbit_r19_c50 bl[50] br[50] wl[19] vdd gnd cell_6t
Xbit_r20_c50 bl[50] br[50] wl[20] vdd gnd cell_6t
Xbit_r21_c50 bl[50] br[50] wl[21] vdd gnd cell_6t
Xbit_r22_c50 bl[50] br[50] wl[22] vdd gnd cell_6t
Xbit_r23_c50 bl[50] br[50] wl[23] vdd gnd cell_6t
Xbit_r24_c50 bl[50] br[50] wl[24] vdd gnd cell_6t
Xbit_r25_c50 bl[50] br[50] wl[25] vdd gnd cell_6t
Xbit_r26_c50 bl[50] br[50] wl[26] vdd gnd cell_6t
Xbit_r27_c50 bl[50] br[50] wl[27] vdd gnd cell_6t
Xbit_r28_c50 bl[50] br[50] wl[28] vdd gnd cell_6t
Xbit_r29_c50 bl[50] br[50] wl[29] vdd gnd cell_6t
Xbit_r30_c50 bl[50] br[50] wl[30] vdd gnd cell_6t
Xbit_r31_c50 bl[50] br[50] wl[31] vdd gnd cell_6t
Xbit_r32_c50 bl[50] br[50] wl[32] vdd gnd cell_6t
Xbit_r33_c50 bl[50] br[50] wl[33] vdd gnd cell_6t
Xbit_r34_c50 bl[50] br[50] wl[34] vdd gnd cell_6t
Xbit_r35_c50 bl[50] br[50] wl[35] vdd gnd cell_6t
Xbit_r36_c50 bl[50] br[50] wl[36] vdd gnd cell_6t
Xbit_r37_c50 bl[50] br[50] wl[37] vdd gnd cell_6t
Xbit_r38_c50 bl[50] br[50] wl[38] vdd gnd cell_6t
Xbit_r39_c50 bl[50] br[50] wl[39] vdd gnd cell_6t
Xbit_r40_c50 bl[50] br[50] wl[40] vdd gnd cell_6t
Xbit_r41_c50 bl[50] br[50] wl[41] vdd gnd cell_6t
Xbit_r42_c50 bl[50] br[50] wl[42] vdd gnd cell_6t
Xbit_r43_c50 bl[50] br[50] wl[43] vdd gnd cell_6t
Xbit_r44_c50 bl[50] br[50] wl[44] vdd gnd cell_6t
Xbit_r45_c50 bl[50] br[50] wl[45] vdd gnd cell_6t
Xbit_r46_c50 bl[50] br[50] wl[46] vdd gnd cell_6t
Xbit_r47_c50 bl[50] br[50] wl[47] vdd gnd cell_6t
Xbit_r48_c50 bl[50] br[50] wl[48] vdd gnd cell_6t
Xbit_r49_c50 bl[50] br[50] wl[49] vdd gnd cell_6t
Xbit_r50_c50 bl[50] br[50] wl[50] vdd gnd cell_6t
Xbit_r51_c50 bl[50] br[50] wl[51] vdd gnd cell_6t
Xbit_r52_c50 bl[50] br[50] wl[52] vdd gnd cell_6t
Xbit_r53_c50 bl[50] br[50] wl[53] vdd gnd cell_6t
Xbit_r54_c50 bl[50] br[50] wl[54] vdd gnd cell_6t
Xbit_r55_c50 bl[50] br[50] wl[55] vdd gnd cell_6t
Xbit_r56_c50 bl[50] br[50] wl[56] vdd gnd cell_6t
Xbit_r57_c50 bl[50] br[50] wl[57] vdd gnd cell_6t
Xbit_r58_c50 bl[50] br[50] wl[58] vdd gnd cell_6t
Xbit_r59_c50 bl[50] br[50] wl[59] vdd gnd cell_6t
Xbit_r60_c50 bl[50] br[50] wl[60] vdd gnd cell_6t
Xbit_r61_c50 bl[50] br[50] wl[61] vdd gnd cell_6t
Xbit_r62_c50 bl[50] br[50] wl[62] vdd gnd cell_6t
Xbit_r63_c50 bl[50] br[50] wl[63] vdd gnd cell_6t
Xbit_r64_c50 bl[50] br[50] wl[64] vdd gnd cell_6t
Xbit_r65_c50 bl[50] br[50] wl[65] vdd gnd cell_6t
Xbit_r66_c50 bl[50] br[50] wl[66] vdd gnd cell_6t
Xbit_r67_c50 bl[50] br[50] wl[67] vdd gnd cell_6t
Xbit_r68_c50 bl[50] br[50] wl[68] vdd gnd cell_6t
Xbit_r69_c50 bl[50] br[50] wl[69] vdd gnd cell_6t
Xbit_r70_c50 bl[50] br[50] wl[70] vdd gnd cell_6t
Xbit_r71_c50 bl[50] br[50] wl[71] vdd gnd cell_6t
Xbit_r72_c50 bl[50] br[50] wl[72] vdd gnd cell_6t
Xbit_r73_c50 bl[50] br[50] wl[73] vdd gnd cell_6t
Xbit_r74_c50 bl[50] br[50] wl[74] vdd gnd cell_6t
Xbit_r75_c50 bl[50] br[50] wl[75] vdd gnd cell_6t
Xbit_r76_c50 bl[50] br[50] wl[76] vdd gnd cell_6t
Xbit_r77_c50 bl[50] br[50] wl[77] vdd gnd cell_6t
Xbit_r78_c50 bl[50] br[50] wl[78] vdd gnd cell_6t
Xbit_r79_c50 bl[50] br[50] wl[79] vdd gnd cell_6t
Xbit_r80_c50 bl[50] br[50] wl[80] vdd gnd cell_6t
Xbit_r81_c50 bl[50] br[50] wl[81] vdd gnd cell_6t
Xbit_r82_c50 bl[50] br[50] wl[82] vdd gnd cell_6t
Xbit_r83_c50 bl[50] br[50] wl[83] vdd gnd cell_6t
Xbit_r84_c50 bl[50] br[50] wl[84] vdd gnd cell_6t
Xbit_r85_c50 bl[50] br[50] wl[85] vdd gnd cell_6t
Xbit_r86_c50 bl[50] br[50] wl[86] vdd gnd cell_6t
Xbit_r87_c50 bl[50] br[50] wl[87] vdd gnd cell_6t
Xbit_r88_c50 bl[50] br[50] wl[88] vdd gnd cell_6t
Xbit_r89_c50 bl[50] br[50] wl[89] vdd gnd cell_6t
Xbit_r90_c50 bl[50] br[50] wl[90] vdd gnd cell_6t
Xbit_r91_c50 bl[50] br[50] wl[91] vdd gnd cell_6t
Xbit_r92_c50 bl[50] br[50] wl[92] vdd gnd cell_6t
Xbit_r93_c50 bl[50] br[50] wl[93] vdd gnd cell_6t
Xbit_r94_c50 bl[50] br[50] wl[94] vdd gnd cell_6t
Xbit_r95_c50 bl[50] br[50] wl[95] vdd gnd cell_6t
Xbit_r96_c50 bl[50] br[50] wl[96] vdd gnd cell_6t
Xbit_r97_c50 bl[50] br[50] wl[97] vdd gnd cell_6t
Xbit_r98_c50 bl[50] br[50] wl[98] vdd gnd cell_6t
Xbit_r99_c50 bl[50] br[50] wl[99] vdd gnd cell_6t
Xbit_r100_c50 bl[50] br[50] wl[100] vdd gnd cell_6t
Xbit_r101_c50 bl[50] br[50] wl[101] vdd gnd cell_6t
Xbit_r102_c50 bl[50] br[50] wl[102] vdd gnd cell_6t
Xbit_r103_c50 bl[50] br[50] wl[103] vdd gnd cell_6t
Xbit_r104_c50 bl[50] br[50] wl[104] vdd gnd cell_6t
Xbit_r105_c50 bl[50] br[50] wl[105] vdd gnd cell_6t
Xbit_r106_c50 bl[50] br[50] wl[106] vdd gnd cell_6t
Xbit_r107_c50 bl[50] br[50] wl[107] vdd gnd cell_6t
Xbit_r108_c50 bl[50] br[50] wl[108] vdd gnd cell_6t
Xbit_r109_c50 bl[50] br[50] wl[109] vdd gnd cell_6t
Xbit_r110_c50 bl[50] br[50] wl[110] vdd gnd cell_6t
Xbit_r111_c50 bl[50] br[50] wl[111] vdd gnd cell_6t
Xbit_r112_c50 bl[50] br[50] wl[112] vdd gnd cell_6t
Xbit_r113_c50 bl[50] br[50] wl[113] vdd gnd cell_6t
Xbit_r114_c50 bl[50] br[50] wl[114] vdd gnd cell_6t
Xbit_r115_c50 bl[50] br[50] wl[115] vdd gnd cell_6t
Xbit_r116_c50 bl[50] br[50] wl[116] vdd gnd cell_6t
Xbit_r117_c50 bl[50] br[50] wl[117] vdd gnd cell_6t
Xbit_r118_c50 bl[50] br[50] wl[118] vdd gnd cell_6t
Xbit_r119_c50 bl[50] br[50] wl[119] vdd gnd cell_6t
Xbit_r120_c50 bl[50] br[50] wl[120] vdd gnd cell_6t
Xbit_r121_c50 bl[50] br[50] wl[121] vdd gnd cell_6t
Xbit_r122_c50 bl[50] br[50] wl[122] vdd gnd cell_6t
Xbit_r123_c50 bl[50] br[50] wl[123] vdd gnd cell_6t
Xbit_r124_c50 bl[50] br[50] wl[124] vdd gnd cell_6t
Xbit_r125_c50 bl[50] br[50] wl[125] vdd gnd cell_6t
Xbit_r126_c50 bl[50] br[50] wl[126] vdd gnd cell_6t
Xbit_r127_c50 bl[50] br[50] wl[127] vdd gnd cell_6t
Xbit_r0_c51 bl[51] br[51] wl[0] vdd gnd cell_6t
Xbit_r1_c51 bl[51] br[51] wl[1] vdd gnd cell_6t
Xbit_r2_c51 bl[51] br[51] wl[2] vdd gnd cell_6t
Xbit_r3_c51 bl[51] br[51] wl[3] vdd gnd cell_6t
Xbit_r4_c51 bl[51] br[51] wl[4] vdd gnd cell_6t
Xbit_r5_c51 bl[51] br[51] wl[5] vdd gnd cell_6t
Xbit_r6_c51 bl[51] br[51] wl[6] vdd gnd cell_6t
Xbit_r7_c51 bl[51] br[51] wl[7] vdd gnd cell_6t
Xbit_r8_c51 bl[51] br[51] wl[8] vdd gnd cell_6t
Xbit_r9_c51 bl[51] br[51] wl[9] vdd gnd cell_6t
Xbit_r10_c51 bl[51] br[51] wl[10] vdd gnd cell_6t
Xbit_r11_c51 bl[51] br[51] wl[11] vdd gnd cell_6t
Xbit_r12_c51 bl[51] br[51] wl[12] vdd gnd cell_6t
Xbit_r13_c51 bl[51] br[51] wl[13] vdd gnd cell_6t
Xbit_r14_c51 bl[51] br[51] wl[14] vdd gnd cell_6t
Xbit_r15_c51 bl[51] br[51] wl[15] vdd gnd cell_6t
Xbit_r16_c51 bl[51] br[51] wl[16] vdd gnd cell_6t
Xbit_r17_c51 bl[51] br[51] wl[17] vdd gnd cell_6t
Xbit_r18_c51 bl[51] br[51] wl[18] vdd gnd cell_6t
Xbit_r19_c51 bl[51] br[51] wl[19] vdd gnd cell_6t
Xbit_r20_c51 bl[51] br[51] wl[20] vdd gnd cell_6t
Xbit_r21_c51 bl[51] br[51] wl[21] vdd gnd cell_6t
Xbit_r22_c51 bl[51] br[51] wl[22] vdd gnd cell_6t
Xbit_r23_c51 bl[51] br[51] wl[23] vdd gnd cell_6t
Xbit_r24_c51 bl[51] br[51] wl[24] vdd gnd cell_6t
Xbit_r25_c51 bl[51] br[51] wl[25] vdd gnd cell_6t
Xbit_r26_c51 bl[51] br[51] wl[26] vdd gnd cell_6t
Xbit_r27_c51 bl[51] br[51] wl[27] vdd gnd cell_6t
Xbit_r28_c51 bl[51] br[51] wl[28] vdd gnd cell_6t
Xbit_r29_c51 bl[51] br[51] wl[29] vdd gnd cell_6t
Xbit_r30_c51 bl[51] br[51] wl[30] vdd gnd cell_6t
Xbit_r31_c51 bl[51] br[51] wl[31] vdd gnd cell_6t
Xbit_r32_c51 bl[51] br[51] wl[32] vdd gnd cell_6t
Xbit_r33_c51 bl[51] br[51] wl[33] vdd gnd cell_6t
Xbit_r34_c51 bl[51] br[51] wl[34] vdd gnd cell_6t
Xbit_r35_c51 bl[51] br[51] wl[35] vdd gnd cell_6t
Xbit_r36_c51 bl[51] br[51] wl[36] vdd gnd cell_6t
Xbit_r37_c51 bl[51] br[51] wl[37] vdd gnd cell_6t
Xbit_r38_c51 bl[51] br[51] wl[38] vdd gnd cell_6t
Xbit_r39_c51 bl[51] br[51] wl[39] vdd gnd cell_6t
Xbit_r40_c51 bl[51] br[51] wl[40] vdd gnd cell_6t
Xbit_r41_c51 bl[51] br[51] wl[41] vdd gnd cell_6t
Xbit_r42_c51 bl[51] br[51] wl[42] vdd gnd cell_6t
Xbit_r43_c51 bl[51] br[51] wl[43] vdd gnd cell_6t
Xbit_r44_c51 bl[51] br[51] wl[44] vdd gnd cell_6t
Xbit_r45_c51 bl[51] br[51] wl[45] vdd gnd cell_6t
Xbit_r46_c51 bl[51] br[51] wl[46] vdd gnd cell_6t
Xbit_r47_c51 bl[51] br[51] wl[47] vdd gnd cell_6t
Xbit_r48_c51 bl[51] br[51] wl[48] vdd gnd cell_6t
Xbit_r49_c51 bl[51] br[51] wl[49] vdd gnd cell_6t
Xbit_r50_c51 bl[51] br[51] wl[50] vdd gnd cell_6t
Xbit_r51_c51 bl[51] br[51] wl[51] vdd gnd cell_6t
Xbit_r52_c51 bl[51] br[51] wl[52] vdd gnd cell_6t
Xbit_r53_c51 bl[51] br[51] wl[53] vdd gnd cell_6t
Xbit_r54_c51 bl[51] br[51] wl[54] vdd gnd cell_6t
Xbit_r55_c51 bl[51] br[51] wl[55] vdd gnd cell_6t
Xbit_r56_c51 bl[51] br[51] wl[56] vdd gnd cell_6t
Xbit_r57_c51 bl[51] br[51] wl[57] vdd gnd cell_6t
Xbit_r58_c51 bl[51] br[51] wl[58] vdd gnd cell_6t
Xbit_r59_c51 bl[51] br[51] wl[59] vdd gnd cell_6t
Xbit_r60_c51 bl[51] br[51] wl[60] vdd gnd cell_6t
Xbit_r61_c51 bl[51] br[51] wl[61] vdd gnd cell_6t
Xbit_r62_c51 bl[51] br[51] wl[62] vdd gnd cell_6t
Xbit_r63_c51 bl[51] br[51] wl[63] vdd gnd cell_6t
Xbit_r64_c51 bl[51] br[51] wl[64] vdd gnd cell_6t
Xbit_r65_c51 bl[51] br[51] wl[65] vdd gnd cell_6t
Xbit_r66_c51 bl[51] br[51] wl[66] vdd gnd cell_6t
Xbit_r67_c51 bl[51] br[51] wl[67] vdd gnd cell_6t
Xbit_r68_c51 bl[51] br[51] wl[68] vdd gnd cell_6t
Xbit_r69_c51 bl[51] br[51] wl[69] vdd gnd cell_6t
Xbit_r70_c51 bl[51] br[51] wl[70] vdd gnd cell_6t
Xbit_r71_c51 bl[51] br[51] wl[71] vdd gnd cell_6t
Xbit_r72_c51 bl[51] br[51] wl[72] vdd gnd cell_6t
Xbit_r73_c51 bl[51] br[51] wl[73] vdd gnd cell_6t
Xbit_r74_c51 bl[51] br[51] wl[74] vdd gnd cell_6t
Xbit_r75_c51 bl[51] br[51] wl[75] vdd gnd cell_6t
Xbit_r76_c51 bl[51] br[51] wl[76] vdd gnd cell_6t
Xbit_r77_c51 bl[51] br[51] wl[77] vdd gnd cell_6t
Xbit_r78_c51 bl[51] br[51] wl[78] vdd gnd cell_6t
Xbit_r79_c51 bl[51] br[51] wl[79] vdd gnd cell_6t
Xbit_r80_c51 bl[51] br[51] wl[80] vdd gnd cell_6t
Xbit_r81_c51 bl[51] br[51] wl[81] vdd gnd cell_6t
Xbit_r82_c51 bl[51] br[51] wl[82] vdd gnd cell_6t
Xbit_r83_c51 bl[51] br[51] wl[83] vdd gnd cell_6t
Xbit_r84_c51 bl[51] br[51] wl[84] vdd gnd cell_6t
Xbit_r85_c51 bl[51] br[51] wl[85] vdd gnd cell_6t
Xbit_r86_c51 bl[51] br[51] wl[86] vdd gnd cell_6t
Xbit_r87_c51 bl[51] br[51] wl[87] vdd gnd cell_6t
Xbit_r88_c51 bl[51] br[51] wl[88] vdd gnd cell_6t
Xbit_r89_c51 bl[51] br[51] wl[89] vdd gnd cell_6t
Xbit_r90_c51 bl[51] br[51] wl[90] vdd gnd cell_6t
Xbit_r91_c51 bl[51] br[51] wl[91] vdd gnd cell_6t
Xbit_r92_c51 bl[51] br[51] wl[92] vdd gnd cell_6t
Xbit_r93_c51 bl[51] br[51] wl[93] vdd gnd cell_6t
Xbit_r94_c51 bl[51] br[51] wl[94] vdd gnd cell_6t
Xbit_r95_c51 bl[51] br[51] wl[95] vdd gnd cell_6t
Xbit_r96_c51 bl[51] br[51] wl[96] vdd gnd cell_6t
Xbit_r97_c51 bl[51] br[51] wl[97] vdd gnd cell_6t
Xbit_r98_c51 bl[51] br[51] wl[98] vdd gnd cell_6t
Xbit_r99_c51 bl[51] br[51] wl[99] vdd gnd cell_6t
Xbit_r100_c51 bl[51] br[51] wl[100] vdd gnd cell_6t
Xbit_r101_c51 bl[51] br[51] wl[101] vdd gnd cell_6t
Xbit_r102_c51 bl[51] br[51] wl[102] vdd gnd cell_6t
Xbit_r103_c51 bl[51] br[51] wl[103] vdd gnd cell_6t
Xbit_r104_c51 bl[51] br[51] wl[104] vdd gnd cell_6t
Xbit_r105_c51 bl[51] br[51] wl[105] vdd gnd cell_6t
Xbit_r106_c51 bl[51] br[51] wl[106] vdd gnd cell_6t
Xbit_r107_c51 bl[51] br[51] wl[107] vdd gnd cell_6t
Xbit_r108_c51 bl[51] br[51] wl[108] vdd gnd cell_6t
Xbit_r109_c51 bl[51] br[51] wl[109] vdd gnd cell_6t
Xbit_r110_c51 bl[51] br[51] wl[110] vdd gnd cell_6t
Xbit_r111_c51 bl[51] br[51] wl[111] vdd gnd cell_6t
Xbit_r112_c51 bl[51] br[51] wl[112] vdd gnd cell_6t
Xbit_r113_c51 bl[51] br[51] wl[113] vdd gnd cell_6t
Xbit_r114_c51 bl[51] br[51] wl[114] vdd gnd cell_6t
Xbit_r115_c51 bl[51] br[51] wl[115] vdd gnd cell_6t
Xbit_r116_c51 bl[51] br[51] wl[116] vdd gnd cell_6t
Xbit_r117_c51 bl[51] br[51] wl[117] vdd gnd cell_6t
Xbit_r118_c51 bl[51] br[51] wl[118] vdd gnd cell_6t
Xbit_r119_c51 bl[51] br[51] wl[119] vdd gnd cell_6t
Xbit_r120_c51 bl[51] br[51] wl[120] vdd gnd cell_6t
Xbit_r121_c51 bl[51] br[51] wl[121] vdd gnd cell_6t
Xbit_r122_c51 bl[51] br[51] wl[122] vdd gnd cell_6t
Xbit_r123_c51 bl[51] br[51] wl[123] vdd gnd cell_6t
Xbit_r124_c51 bl[51] br[51] wl[124] vdd gnd cell_6t
Xbit_r125_c51 bl[51] br[51] wl[125] vdd gnd cell_6t
Xbit_r126_c51 bl[51] br[51] wl[126] vdd gnd cell_6t
Xbit_r127_c51 bl[51] br[51] wl[127] vdd gnd cell_6t
Xbit_r0_c52 bl[52] br[52] wl[0] vdd gnd cell_6t
Xbit_r1_c52 bl[52] br[52] wl[1] vdd gnd cell_6t
Xbit_r2_c52 bl[52] br[52] wl[2] vdd gnd cell_6t
Xbit_r3_c52 bl[52] br[52] wl[3] vdd gnd cell_6t
Xbit_r4_c52 bl[52] br[52] wl[4] vdd gnd cell_6t
Xbit_r5_c52 bl[52] br[52] wl[5] vdd gnd cell_6t
Xbit_r6_c52 bl[52] br[52] wl[6] vdd gnd cell_6t
Xbit_r7_c52 bl[52] br[52] wl[7] vdd gnd cell_6t
Xbit_r8_c52 bl[52] br[52] wl[8] vdd gnd cell_6t
Xbit_r9_c52 bl[52] br[52] wl[9] vdd gnd cell_6t
Xbit_r10_c52 bl[52] br[52] wl[10] vdd gnd cell_6t
Xbit_r11_c52 bl[52] br[52] wl[11] vdd gnd cell_6t
Xbit_r12_c52 bl[52] br[52] wl[12] vdd gnd cell_6t
Xbit_r13_c52 bl[52] br[52] wl[13] vdd gnd cell_6t
Xbit_r14_c52 bl[52] br[52] wl[14] vdd gnd cell_6t
Xbit_r15_c52 bl[52] br[52] wl[15] vdd gnd cell_6t
Xbit_r16_c52 bl[52] br[52] wl[16] vdd gnd cell_6t
Xbit_r17_c52 bl[52] br[52] wl[17] vdd gnd cell_6t
Xbit_r18_c52 bl[52] br[52] wl[18] vdd gnd cell_6t
Xbit_r19_c52 bl[52] br[52] wl[19] vdd gnd cell_6t
Xbit_r20_c52 bl[52] br[52] wl[20] vdd gnd cell_6t
Xbit_r21_c52 bl[52] br[52] wl[21] vdd gnd cell_6t
Xbit_r22_c52 bl[52] br[52] wl[22] vdd gnd cell_6t
Xbit_r23_c52 bl[52] br[52] wl[23] vdd gnd cell_6t
Xbit_r24_c52 bl[52] br[52] wl[24] vdd gnd cell_6t
Xbit_r25_c52 bl[52] br[52] wl[25] vdd gnd cell_6t
Xbit_r26_c52 bl[52] br[52] wl[26] vdd gnd cell_6t
Xbit_r27_c52 bl[52] br[52] wl[27] vdd gnd cell_6t
Xbit_r28_c52 bl[52] br[52] wl[28] vdd gnd cell_6t
Xbit_r29_c52 bl[52] br[52] wl[29] vdd gnd cell_6t
Xbit_r30_c52 bl[52] br[52] wl[30] vdd gnd cell_6t
Xbit_r31_c52 bl[52] br[52] wl[31] vdd gnd cell_6t
Xbit_r32_c52 bl[52] br[52] wl[32] vdd gnd cell_6t
Xbit_r33_c52 bl[52] br[52] wl[33] vdd gnd cell_6t
Xbit_r34_c52 bl[52] br[52] wl[34] vdd gnd cell_6t
Xbit_r35_c52 bl[52] br[52] wl[35] vdd gnd cell_6t
Xbit_r36_c52 bl[52] br[52] wl[36] vdd gnd cell_6t
Xbit_r37_c52 bl[52] br[52] wl[37] vdd gnd cell_6t
Xbit_r38_c52 bl[52] br[52] wl[38] vdd gnd cell_6t
Xbit_r39_c52 bl[52] br[52] wl[39] vdd gnd cell_6t
Xbit_r40_c52 bl[52] br[52] wl[40] vdd gnd cell_6t
Xbit_r41_c52 bl[52] br[52] wl[41] vdd gnd cell_6t
Xbit_r42_c52 bl[52] br[52] wl[42] vdd gnd cell_6t
Xbit_r43_c52 bl[52] br[52] wl[43] vdd gnd cell_6t
Xbit_r44_c52 bl[52] br[52] wl[44] vdd gnd cell_6t
Xbit_r45_c52 bl[52] br[52] wl[45] vdd gnd cell_6t
Xbit_r46_c52 bl[52] br[52] wl[46] vdd gnd cell_6t
Xbit_r47_c52 bl[52] br[52] wl[47] vdd gnd cell_6t
Xbit_r48_c52 bl[52] br[52] wl[48] vdd gnd cell_6t
Xbit_r49_c52 bl[52] br[52] wl[49] vdd gnd cell_6t
Xbit_r50_c52 bl[52] br[52] wl[50] vdd gnd cell_6t
Xbit_r51_c52 bl[52] br[52] wl[51] vdd gnd cell_6t
Xbit_r52_c52 bl[52] br[52] wl[52] vdd gnd cell_6t
Xbit_r53_c52 bl[52] br[52] wl[53] vdd gnd cell_6t
Xbit_r54_c52 bl[52] br[52] wl[54] vdd gnd cell_6t
Xbit_r55_c52 bl[52] br[52] wl[55] vdd gnd cell_6t
Xbit_r56_c52 bl[52] br[52] wl[56] vdd gnd cell_6t
Xbit_r57_c52 bl[52] br[52] wl[57] vdd gnd cell_6t
Xbit_r58_c52 bl[52] br[52] wl[58] vdd gnd cell_6t
Xbit_r59_c52 bl[52] br[52] wl[59] vdd gnd cell_6t
Xbit_r60_c52 bl[52] br[52] wl[60] vdd gnd cell_6t
Xbit_r61_c52 bl[52] br[52] wl[61] vdd gnd cell_6t
Xbit_r62_c52 bl[52] br[52] wl[62] vdd gnd cell_6t
Xbit_r63_c52 bl[52] br[52] wl[63] vdd gnd cell_6t
Xbit_r64_c52 bl[52] br[52] wl[64] vdd gnd cell_6t
Xbit_r65_c52 bl[52] br[52] wl[65] vdd gnd cell_6t
Xbit_r66_c52 bl[52] br[52] wl[66] vdd gnd cell_6t
Xbit_r67_c52 bl[52] br[52] wl[67] vdd gnd cell_6t
Xbit_r68_c52 bl[52] br[52] wl[68] vdd gnd cell_6t
Xbit_r69_c52 bl[52] br[52] wl[69] vdd gnd cell_6t
Xbit_r70_c52 bl[52] br[52] wl[70] vdd gnd cell_6t
Xbit_r71_c52 bl[52] br[52] wl[71] vdd gnd cell_6t
Xbit_r72_c52 bl[52] br[52] wl[72] vdd gnd cell_6t
Xbit_r73_c52 bl[52] br[52] wl[73] vdd gnd cell_6t
Xbit_r74_c52 bl[52] br[52] wl[74] vdd gnd cell_6t
Xbit_r75_c52 bl[52] br[52] wl[75] vdd gnd cell_6t
Xbit_r76_c52 bl[52] br[52] wl[76] vdd gnd cell_6t
Xbit_r77_c52 bl[52] br[52] wl[77] vdd gnd cell_6t
Xbit_r78_c52 bl[52] br[52] wl[78] vdd gnd cell_6t
Xbit_r79_c52 bl[52] br[52] wl[79] vdd gnd cell_6t
Xbit_r80_c52 bl[52] br[52] wl[80] vdd gnd cell_6t
Xbit_r81_c52 bl[52] br[52] wl[81] vdd gnd cell_6t
Xbit_r82_c52 bl[52] br[52] wl[82] vdd gnd cell_6t
Xbit_r83_c52 bl[52] br[52] wl[83] vdd gnd cell_6t
Xbit_r84_c52 bl[52] br[52] wl[84] vdd gnd cell_6t
Xbit_r85_c52 bl[52] br[52] wl[85] vdd gnd cell_6t
Xbit_r86_c52 bl[52] br[52] wl[86] vdd gnd cell_6t
Xbit_r87_c52 bl[52] br[52] wl[87] vdd gnd cell_6t
Xbit_r88_c52 bl[52] br[52] wl[88] vdd gnd cell_6t
Xbit_r89_c52 bl[52] br[52] wl[89] vdd gnd cell_6t
Xbit_r90_c52 bl[52] br[52] wl[90] vdd gnd cell_6t
Xbit_r91_c52 bl[52] br[52] wl[91] vdd gnd cell_6t
Xbit_r92_c52 bl[52] br[52] wl[92] vdd gnd cell_6t
Xbit_r93_c52 bl[52] br[52] wl[93] vdd gnd cell_6t
Xbit_r94_c52 bl[52] br[52] wl[94] vdd gnd cell_6t
Xbit_r95_c52 bl[52] br[52] wl[95] vdd gnd cell_6t
Xbit_r96_c52 bl[52] br[52] wl[96] vdd gnd cell_6t
Xbit_r97_c52 bl[52] br[52] wl[97] vdd gnd cell_6t
Xbit_r98_c52 bl[52] br[52] wl[98] vdd gnd cell_6t
Xbit_r99_c52 bl[52] br[52] wl[99] vdd gnd cell_6t
Xbit_r100_c52 bl[52] br[52] wl[100] vdd gnd cell_6t
Xbit_r101_c52 bl[52] br[52] wl[101] vdd gnd cell_6t
Xbit_r102_c52 bl[52] br[52] wl[102] vdd gnd cell_6t
Xbit_r103_c52 bl[52] br[52] wl[103] vdd gnd cell_6t
Xbit_r104_c52 bl[52] br[52] wl[104] vdd gnd cell_6t
Xbit_r105_c52 bl[52] br[52] wl[105] vdd gnd cell_6t
Xbit_r106_c52 bl[52] br[52] wl[106] vdd gnd cell_6t
Xbit_r107_c52 bl[52] br[52] wl[107] vdd gnd cell_6t
Xbit_r108_c52 bl[52] br[52] wl[108] vdd gnd cell_6t
Xbit_r109_c52 bl[52] br[52] wl[109] vdd gnd cell_6t
Xbit_r110_c52 bl[52] br[52] wl[110] vdd gnd cell_6t
Xbit_r111_c52 bl[52] br[52] wl[111] vdd gnd cell_6t
Xbit_r112_c52 bl[52] br[52] wl[112] vdd gnd cell_6t
Xbit_r113_c52 bl[52] br[52] wl[113] vdd gnd cell_6t
Xbit_r114_c52 bl[52] br[52] wl[114] vdd gnd cell_6t
Xbit_r115_c52 bl[52] br[52] wl[115] vdd gnd cell_6t
Xbit_r116_c52 bl[52] br[52] wl[116] vdd gnd cell_6t
Xbit_r117_c52 bl[52] br[52] wl[117] vdd gnd cell_6t
Xbit_r118_c52 bl[52] br[52] wl[118] vdd gnd cell_6t
Xbit_r119_c52 bl[52] br[52] wl[119] vdd gnd cell_6t
Xbit_r120_c52 bl[52] br[52] wl[120] vdd gnd cell_6t
Xbit_r121_c52 bl[52] br[52] wl[121] vdd gnd cell_6t
Xbit_r122_c52 bl[52] br[52] wl[122] vdd gnd cell_6t
Xbit_r123_c52 bl[52] br[52] wl[123] vdd gnd cell_6t
Xbit_r124_c52 bl[52] br[52] wl[124] vdd gnd cell_6t
Xbit_r125_c52 bl[52] br[52] wl[125] vdd gnd cell_6t
Xbit_r126_c52 bl[52] br[52] wl[126] vdd gnd cell_6t
Xbit_r127_c52 bl[52] br[52] wl[127] vdd gnd cell_6t
Xbit_r0_c53 bl[53] br[53] wl[0] vdd gnd cell_6t
Xbit_r1_c53 bl[53] br[53] wl[1] vdd gnd cell_6t
Xbit_r2_c53 bl[53] br[53] wl[2] vdd gnd cell_6t
Xbit_r3_c53 bl[53] br[53] wl[3] vdd gnd cell_6t
Xbit_r4_c53 bl[53] br[53] wl[4] vdd gnd cell_6t
Xbit_r5_c53 bl[53] br[53] wl[5] vdd gnd cell_6t
Xbit_r6_c53 bl[53] br[53] wl[6] vdd gnd cell_6t
Xbit_r7_c53 bl[53] br[53] wl[7] vdd gnd cell_6t
Xbit_r8_c53 bl[53] br[53] wl[8] vdd gnd cell_6t
Xbit_r9_c53 bl[53] br[53] wl[9] vdd gnd cell_6t
Xbit_r10_c53 bl[53] br[53] wl[10] vdd gnd cell_6t
Xbit_r11_c53 bl[53] br[53] wl[11] vdd gnd cell_6t
Xbit_r12_c53 bl[53] br[53] wl[12] vdd gnd cell_6t
Xbit_r13_c53 bl[53] br[53] wl[13] vdd gnd cell_6t
Xbit_r14_c53 bl[53] br[53] wl[14] vdd gnd cell_6t
Xbit_r15_c53 bl[53] br[53] wl[15] vdd gnd cell_6t
Xbit_r16_c53 bl[53] br[53] wl[16] vdd gnd cell_6t
Xbit_r17_c53 bl[53] br[53] wl[17] vdd gnd cell_6t
Xbit_r18_c53 bl[53] br[53] wl[18] vdd gnd cell_6t
Xbit_r19_c53 bl[53] br[53] wl[19] vdd gnd cell_6t
Xbit_r20_c53 bl[53] br[53] wl[20] vdd gnd cell_6t
Xbit_r21_c53 bl[53] br[53] wl[21] vdd gnd cell_6t
Xbit_r22_c53 bl[53] br[53] wl[22] vdd gnd cell_6t
Xbit_r23_c53 bl[53] br[53] wl[23] vdd gnd cell_6t
Xbit_r24_c53 bl[53] br[53] wl[24] vdd gnd cell_6t
Xbit_r25_c53 bl[53] br[53] wl[25] vdd gnd cell_6t
Xbit_r26_c53 bl[53] br[53] wl[26] vdd gnd cell_6t
Xbit_r27_c53 bl[53] br[53] wl[27] vdd gnd cell_6t
Xbit_r28_c53 bl[53] br[53] wl[28] vdd gnd cell_6t
Xbit_r29_c53 bl[53] br[53] wl[29] vdd gnd cell_6t
Xbit_r30_c53 bl[53] br[53] wl[30] vdd gnd cell_6t
Xbit_r31_c53 bl[53] br[53] wl[31] vdd gnd cell_6t
Xbit_r32_c53 bl[53] br[53] wl[32] vdd gnd cell_6t
Xbit_r33_c53 bl[53] br[53] wl[33] vdd gnd cell_6t
Xbit_r34_c53 bl[53] br[53] wl[34] vdd gnd cell_6t
Xbit_r35_c53 bl[53] br[53] wl[35] vdd gnd cell_6t
Xbit_r36_c53 bl[53] br[53] wl[36] vdd gnd cell_6t
Xbit_r37_c53 bl[53] br[53] wl[37] vdd gnd cell_6t
Xbit_r38_c53 bl[53] br[53] wl[38] vdd gnd cell_6t
Xbit_r39_c53 bl[53] br[53] wl[39] vdd gnd cell_6t
Xbit_r40_c53 bl[53] br[53] wl[40] vdd gnd cell_6t
Xbit_r41_c53 bl[53] br[53] wl[41] vdd gnd cell_6t
Xbit_r42_c53 bl[53] br[53] wl[42] vdd gnd cell_6t
Xbit_r43_c53 bl[53] br[53] wl[43] vdd gnd cell_6t
Xbit_r44_c53 bl[53] br[53] wl[44] vdd gnd cell_6t
Xbit_r45_c53 bl[53] br[53] wl[45] vdd gnd cell_6t
Xbit_r46_c53 bl[53] br[53] wl[46] vdd gnd cell_6t
Xbit_r47_c53 bl[53] br[53] wl[47] vdd gnd cell_6t
Xbit_r48_c53 bl[53] br[53] wl[48] vdd gnd cell_6t
Xbit_r49_c53 bl[53] br[53] wl[49] vdd gnd cell_6t
Xbit_r50_c53 bl[53] br[53] wl[50] vdd gnd cell_6t
Xbit_r51_c53 bl[53] br[53] wl[51] vdd gnd cell_6t
Xbit_r52_c53 bl[53] br[53] wl[52] vdd gnd cell_6t
Xbit_r53_c53 bl[53] br[53] wl[53] vdd gnd cell_6t
Xbit_r54_c53 bl[53] br[53] wl[54] vdd gnd cell_6t
Xbit_r55_c53 bl[53] br[53] wl[55] vdd gnd cell_6t
Xbit_r56_c53 bl[53] br[53] wl[56] vdd gnd cell_6t
Xbit_r57_c53 bl[53] br[53] wl[57] vdd gnd cell_6t
Xbit_r58_c53 bl[53] br[53] wl[58] vdd gnd cell_6t
Xbit_r59_c53 bl[53] br[53] wl[59] vdd gnd cell_6t
Xbit_r60_c53 bl[53] br[53] wl[60] vdd gnd cell_6t
Xbit_r61_c53 bl[53] br[53] wl[61] vdd gnd cell_6t
Xbit_r62_c53 bl[53] br[53] wl[62] vdd gnd cell_6t
Xbit_r63_c53 bl[53] br[53] wl[63] vdd gnd cell_6t
Xbit_r64_c53 bl[53] br[53] wl[64] vdd gnd cell_6t
Xbit_r65_c53 bl[53] br[53] wl[65] vdd gnd cell_6t
Xbit_r66_c53 bl[53] br[53] wl[66] vdd gnd cell_6t
Xbit_r67_c53 bl[53] br[53] wl[67] vdd gnd cell_6t
Xbit_r68_c53 bl[53] br[53] wl[68] vdd gnd cell_6t
Xbit_r69_c53 bl[53] br[53] wl[69] vdd gnd cell_6t
Xbit_r70_c53 bl[53] br[53] wl[70] vdd gnd cell_6t
Xbit_r71_c53 bl[53] br[53] wl[71] vdd gnd cell_6t
Xbit_r72_c53 bl[53] br[53] wl[72] vdd gnd cell_6t
Xbit_r73_c53 bl[53] br[53] wl[73] vdd gnd cell_6t
Xbit_r74_c53 bl[53] br[53] wl[74] vdd gnd cell_6t
Xbit_r75_c53 bl[53] br[53] wl[75] vdd gnd cell_6t
Xbit_r76_c53 bl[53] br[53] wl[76] vdd gnd cell_6t
Xbit_r77_c53 bl[53] br[53] wl[77] vdd gnd cell_6t
Xbit_r78_c53 bl[53] br[53] wl[78] vdd gnd cell_6t
Xbit_r79_c53 bl[53] br[53] wl[79] vdd gnd cell_6t
Xbit_r80_c53 bl[53] br[53] wl[80] vdd gnd cell_6t
Xbit_r81_c53 bl[53] br[53] wl[81] vdd gnd cell_6t
Xbit_r82_c53 bl[53] br[53] wl[82] vdd gnd cell_6t
Xbit_r83_c53 bl[53] br[53] wl[83] vdd gnd cell_6t
Xbit_r84_c53 bl[53] br[53] wl[84] vdd gnd cell_6t
Xbit_r85_c53 bl[53] br[53] wl[85] vdd gnd cell_6t
Xbit_r86_c53 bl[53] br[53] wl[86] vdd gnd cell_6t
Xbit_r87_c53 bl[53] br[53] wl[87] vdd gnd cell_6t
Xbit_r88_c53 bl[53] br[53] wl[88] vdd gnd cell_6t
Xbit_r89_c53 bl[53] br[53] wl[89] vdd gnd cell_6t
Xbit_r90_c53 bl[53] br[53] wl[90] vdd gnd cell_6t
Xbit_r91_c53 bl[53] br[53] wl[91] vdd gnd cell_6t
Xbit_r92_c53 bl[53] br[53] wl[92] vdd gnd cell_6t
Xbit_r93_c53 bl[53] br[53] wl[93] vdd gnd cell_6t
Xbit_r94_c53 bl[53] br[53] wl[94] vdd gnd cell_6t
Xbit_r95_c53 bl[53] br[53] wl[95] vdd gnd cell_6t
Xbit_r96_c53 bl[53] br[53] wl[96] vdd gnd cell_6t
Xbit_r97_c53 bl[53] br[53] wl[97] vdd gnd cell_6t
Xbit_r98_c53 bl[53] br[53] wl[98] vdd gnd cell_6t
Xbit_r99_c53 bl[53] br[53] wl[99] vdd gnd cell_6t
Xbit_r100_c53 bl[53] br[53] wl[100] vdd gnd cell_6t
Xbit_r101_c53 bl[53] br[53] wl[101] vdd gnd cell_6t
Xbit_r102_c53 bl[53] br[53] wl[102] vdd gnd cell_6t
Xbit_r103_c53 bl[53] br[53] wl[103] vdd gnd cell_6t
Xbit_r104_c53 bl[53] br[53] wl[104] vdd gnd cell_6t
Xbit_r105_c53 bl[53] br[53] wl[105] vdd gnd cell_6t
Xbit_r106_c53 bl[53] br[53] wl[106] vdd gnd cell_6t
Xbit_r107_c53 bl[53] br[53] wl[107] vdd gnd cell_6t
Xbit_r108_c53 bl[53] br[53] wl[108] vdd gnd cell_6t
Xbit_r109_c53 bl[53] br[53] wl[109] vdd gnd cell_6t
Xbit_r110_c53 bl[53] br[53] wl[110] vdd gnd cell_6t
Xbit_r111_c53 bl[53] br[53] wl[111] vdd gnd cell_6t
Xbit_r112_c53 bl[53] br[53] wl[112] vdd gnd cell_6t
Xbit_r113_c53 bl[53] br[53] wl[113] vdd gnd cell_6t
Xbit_r114_c53 bl[53] br[53] wl[114] vdd gnd cell_6t
Xbit_r115_c53 bl[53] br[53] wl[115] vdd gnd cell_6t
Xbit_r116_c53 bl[53] br[53] wl[116] vdd gnd cell_6t
Xbit_r117_c53 bl[53] br[53] wl[117] vdd gnd cell_6t
Xbit_r118_c53 bl[53] br[53] wl[118] vdd gnd cell_6t
Xbit_r119_c53 bl[53] br[53] wl[119] vdd gnd cell_6t
Xbit_r120_c53 bl[53] br[53] wl[120] vdd gnd cell_6t
Xbit_r121_c53 bl[53] br[53] wl[121] vdd gnd cell_6t
Xbit_r122_c53 bl[53] br[53] wl[122] vdd gnd cell_6t
Xbit_r123_c53 bl[53] br[53] wl[123] vdd gnd cell_6t
Xbit_r124_c53 bl[53] br[53] wl[124] vdd gnd cell_6t
Xbit_r125_c53 bl[53] br[53] wl[125] vdd gnd cell_6t
Xbit_r126_c53 bl[53] br[53] wl[126] vdd gnd cell_6t
Xbit_r127_c53 bl[53] br[53] wl[127] vdd gnd cell_6t
Xbit_r0_c54 bl[54] br[54] wl[0] vdd gnd cell_6t
Xbit_r1_c54 bl[54] br[54] wl[1] vdd gnd cell_6t
Xbit_r2_c54 bl[54] br[54] wl[2] vdd gnd cell_6t
Xbit_r3_c54 bl[54] br[54] wl[3] vdd gnd cell_6t
Xbit_r4_c54 bl[54] br[54] wl[4] vdd gnd cell_6t
Xbit_r5_c54 bl[54] br[54] wl[5] vdd gnd cell_6t
Xbit_r6_c54 bl[54] br[54] wl[6] vdd gnd cell_6t
Xbit_r7_c54 bl[54] br[54] wl[7] vdd gnd cell_6t
Xbit_r8_c54 bl[54] br[54] wl[8] vdd gnd cell_6t
Xbit_r9_c54 bl[54] br[54] wl[9] vdd gnd cell_6t
Xbit_r10_c54 bl[54] br[54] wl[10] vdd gnd cell_6t
Xbit_r11_c54 bl[54] br[54] wl[11] vdd gnd cell_6t
Xbit_r12_c54 bl[54] br[54] wl[12] vdd gnd cell_6t
Xbit_r13_c54 bl[54] br[54] wl[13] vdd gnd cell_6t
Xbit_r14_c54 bl[54] br[54] wl[14] vdd gnd cell_6t
Xbit_r15_c54 bl[54] br[54] wl[15] vdd gnd cell_6t
Xbit_r16_c54 bl[54] br[54] wl[16] vdd gnd cell_6t
Xbit_r17_c54 bl[54] br[54] wl[17] vdd gnd cell_6t
Xbit_r18_c54 bl[54] br[54] wl[18] vdd gnd cell_6t
Xbit_r19_c54 bl[54] br[54] wl[19] vdd gnd cell_6t
Xbit_r20_c54 bl[54] br[54] wl[20] vdd gnd cell_6t
Xbit_r21_c54 bl[54] br[54] wl[21] vdd gnd cell_6t
Xbit_r22_c54 bl[54] br[54] wl[22] vdd gnd cell_6t
Xbit_r23_c54 bl[54] br[54] wl[23] vdd gnd cell_6t
Xbit_r24_c54 bl[54] br[54] wl[24] vdd gnd cell_6t
Xbit_r25_c54 bl[54] br[54] wl[25] vdd gnd cell_6t
Xbit_r26_c54 bl[54] br[54] wl[26] vdd gnd cell_6t
Xbit_r27_c54 bl[54] br[54] wl[27] vdd gnd cell_6t
Xbit_r28_c54 bl[54] br[54] wl[28] vdd gnd cell_6t
Xbit_r29_c54 bl[54] br[54] wl[29] vdd gnd cell_6t
Xbit_r30_c54 bl[54] br[54] wl[30] vdd gnd cell_6t
Xbit_r31_c54 bl[54] br[54] wl[31] vdd gnd cell_6t
Xbit_r32_c54 bl[54] br[54] wl[32] vdd gnd cell_6t
Xbit_r33_c54 bl[54] br[54] wl[33] vdd gnd cell_6t
Xbit_r34_c54 bl[54] br[54] wl[34] vdd gnd cell_6t
Xbit_r35_c54 bl[54] br[54] wl[35] vdd gnd cell_6t
Xbit_r36_c54 bl[54] br[54] wl[36] vdd gnd cell_6t
Xbit_r37_c54 bl[54] br[54] wl[37] vdd gnd cell_6t
Xbit_r38_c54 bl[54] br[54] wl[38] vdd gnd cell_6t
Xbit_r39_c54 bl[54] br[54] wl[39] vdd gnd cell_6t
Xbit_r40_c54 bl[54] br[54] wl[40] vdd gnd cell_6t
Xbit_r41_c54 bl[54] br[54] wl[41] vdd gnd cell_6t
Xbit_r42_c54 bl[54] br[54] wl[42] vdd gnd cell_6t
Xbit_r43_c54 bl[54] br[54] wl[43] vdd gnd cell_6t
Xbit_r44_c54 bl[54] br[54] wl[44] vdd gnd cell_6t
Xbit_r45_c54 bl[54] br[54] wl[45] vdd gnd cell_6t
Xbit_r46_c54 bl[54] br[54] wl[46] vdd gnd cell_6t
Xbit_r47_c54 bl[54] br[54] wl[47] vdd gnd cell_6t
Xbit_r48_c54 bl[54] br[54] wl[48] vdd gnd cell_6t
Xbit_r49_c54 bl[54] br[54] wl[49] vdd gnd cell_6t
Xbit_r50_c54 bl[54] br[54] wl[50] vdd gnd cell_6t
Xbit_r51_c54 bl[54] br[54] wl[51] vdd gnd cell_6t
Xbit_r52_c54 bl[54] br[54] wl[52] vdd gnd cell_6t
Xbit_r53_c54 bl[54] br[54] wl[53] vdd gnd cell_6t
Xbit_r54_c54 bl[54] br[54] wl[54] vdd gnd cell_6t
Xbit_r55_c54 bl[54] br[54] wl[55] vdd gnd cell_6t
Xbit_r56_c54 bl[54] br[54] wl[56] vdd gnd cell_6t
Xbit_r57_c54 bl[54] br[54] wl[57] vdd gnd cell_6t
Xbit_r58_c54 bl[54] br[54] wl[58] vdd gnd cell_6t
Xbit_r59_c54 bl[54] br[54] wl[59] vdd gnd cell_6t
Xbit_r60_c54 bl[54] br[54] wl[60] vdd gnd cell_6t
Xbit_r61_c54 bl[54] br[54] wl[61] vdd gnd cell_6t
Xbit_r62_c54 bl[54] br[54] wl[62] vdd gnd cell_6t
Xbit_r63_c54 bl[54] br[54] wl[63] vdd gnd cell_6t
Xbit_r64_c54 bl[54] br[54] wl[64] vdd gnd cell_6t
Xbit_r65_c54 bl[54] br[54] wl[65] vdd gnd cell_6t
Xbit_r66_c54 bl[54] br[54] wl[66] vdd gnd cell_6t
Xbit_r67_c54 bl[54] br[54] wl[67] vdd gnd cell_6t
Xbit_r68_c54 bl[54] br[54] wl[68] vdd gnd cell_6t
Xbit_r69_c54 bl[54] br[54] wl[69] vdd gnd cell_6t
Xbit_r70_c54 bl[54] br[54] wl[70] vdd gnd cell_6t
Xbit_r71_c54 bl[54] br[54] wl[71] vdd gnd cell_6t
Xbit_r72_c54 bl[54] br[54] wl[72] vdd gnd cell_6t
Xbit_r73_c54 bl[54] br[54] wl[73] vdd gnd cell_6t
Xbit_r74_c54 bl[54] br[54] wl[74] vdd gnd cell_6t
Xbit_r75_c54 bl[54] br[54] wl[75] vdd gnd cell_6t
Xbit_r76_c54 bl[54] br[54] wl[76] vdd gnd cell_6t
Xbit_r77_c54 bl[54] br[54] wl[77] vdd gnd cell_6t
Xbit_r78_c54 bl[54] br[54] wl[78] vdd gnd cell_6t
Xbit_r79_c54 bl[54] br[54] wl[79] vdd gnd cell_6t
Xbit_r80_c54 bl[54] br[54] wl[80] vdd gnd cell_6t
Xbit_r81_c54 bl[54] br[54] wl[81] vdd gnd cell_6t
Xbit_r82_c54 bl[54] br[54] wl[82] vdd gnd cell_6t
Xbit_r83_c54 bl[54] br[54] wl[83] vdd gnd cell_6t
Xbit_r84_c54 bl[54] br[54] wl[84] vdd gnd cell_6t
Xbit_r85_c54 bl[54] br[54] wl[85] vdd gnd cell_6t
Xbit_r86_c54 bl[54] br[54] wl[86] vdd gnd cell_6t
Xbit_r87_c54 bl[54] br[54] wl[87] vdd gnd cell_6t
Xbit_r88_c54 bl[54] br[54] wl[88] vdd gnd cell_6t
Xbit_r89_c54 bl[54] br[54] wl[89] vdd gnd cell_6t
Xbit_r90_c54 bl[54] br[54] wl[90] vdd gnd cell_6t
Xbit_r91_c54 bl[54] br[54] wl[91] vdd gnd cell_6t
Xbit_r92_c54 bl[54] br[54] wl[92] vdd gnd cell_6t
Xbit_r93_c54 bl[54] br[54] wl[93] vdd gnd cell_6t
Xbit_r94_c54 bl[54] br[54] wl[94] vdd gnd cell_6t
Xbit_r95_c54 bl[54] br[54] wl[95] vdd gnd cell_6t
Xbit_r96_c54 bl[54] br[54] wl[96] vdd gnd cell_6t
Xbit_r97_c54 bl[54] br[54] wl[97] vdd gnd cell_6t
Xbit_r98_c54 bl[54] br[54] wl[98] vdd gnd cell_6t
Xbit_r99_c54 bl[54] br[54] wl[99] vdd gnd cell_6t
Xbit_r100_c54 bl[54] br[54] wl[100] vdd gnd cell_6t
Xbit_r101_c54 bl[54] br[54] wl[101] vdd gnd cell_6t
Xbit_r102_c54 bl[54] br[54] wl[102] vdd gnd cell_6t
Xbit_r103_c54 bl[54] br[54] wl[103] vdd gnd cell_6t
Xbit_r104_c54 bl[54] br[54] wl[104] vdd gnd cell_6t
Xbit_r105_c54 bl[54] br[54] wl[105] vdd gnd cell_6t
Xbit_r106_c54 bl[54] br[54] wl[106] vdd gnd cell_6t
Xbit_r107_c54 bl[54] br[54] wl[107] vdd gnd cell_6t
Xbit_r108_c54 bl[54] br[54] wl[108] vdd gnd cell_6t
Xbit_r109_c54 bl[54] br[54] wl[109] vdd gnd cell_6t
Xbit_r110_c54 bl[54] br[54] wl[110] vdd gnd cell_6t
Xbit_r111_c54 bl[54] br[54] wl[111] vdd gnd cell_6t
Xbit_r112_c54 bl[54] br[54] wl[112] vdd gnd cell_6t
Xbit_r113_c54 bl[54] br[54] wl[113] vdd gnd cell_6t
Xbit_r114_c54 bl[54] br[54] wl[114] vdd gnd cell_6t
Xbit_r115_c54 bl[54] br[54] wl[115] vdd gnd cell_6t
Xbit_r116_c54 bl[54] br[54] wl[116] vdd gnd cell_6t
Xbit_r117_c54 bl[54] br[54] wl[117] vdd gnd cell_6t
Xbit_r118_c54 bl[54] br[54] wl[118] vdd gnd cell_6t
Xbit_r119_c54 bl[54] br[54] wl[119] vdd gnd cell_6t
Xbit_r120_c54 bl[54] br[54] wl[120] vdd gnd cell_6t
Xbit_r121_c54 bl[54] br[54] wl[121] vdd gnd cell_6t
Xbit_r122_c54 bl[54] br[54] wl[122] vdd gnd cell_6t
Xbit_r123_c54 bl[54] br[54] wl[123] vdd gnd cell_6t
Xbit_r124_c54 bl[54] br[54] wl[124] vdd gnd cell_6t
Xbit_r125_c54 bl[54] br[54] wl[125] vdd gnd cell_6t
Xbit_r126_c54 bl[54] br[54] wl[126] vdd gnd cell_6t
Xbit_r127_c54 bl[54] br[54] wl[127] vdd gnd cell_6t
Xbit_r0_c55 bl[55] br[55] wl[0] vdd gnd cell_6t
Xbit_r1_c55 bl[55] br[55] wl[1] vdd gnd cell_6t
Xbit_r2_c55 bl[55] br[55] wl[2] vdd gnd cell_6t
Xbit_r3_c55 bl[55] br[55] wl[3] vdd gnd cell_6t
Xbit_r4_c55 bl[55] br[55] wl[4] vdd gnd cell_6t
Xbit_r5_c55 bl[55] br[55] wl[5] vdd gnd cell_6t
Xbit_r6_c55 bl[55] br[55] wl[6] vdd gnd cell_6t
Xbit_r7_c55 bl[55] br[55] wl[7] vdd gnd cell_6t
Xbit_r8_c55 bl[55] br[55] wl[8] vdd gnd cell_6t
Xbit_r9_c55 bl[55] br[55] wl[9] vdd gnd cell_6t
Xbit_r10_c55 bl[55] br[55] wl[10] vdd gnd cell_6t
Xbit_r11_c55 bl[55] br[55] wl[11] vdd gnd cell_6t
Xbit_r12_c55 bl[55] br[55] wl[12] vdd gnd cell_6t
Xbit_r13_c55 bl[55] br[55] wl[13] vdd gnd cell_6t
Xbit_r14_c55 bl[55] br[55] wl[14] vdd gnd cell_6t
Xbit_r15_c55 bl[55] br[55] wl[15] vdd gnd cell_6t
Xbit_r16_c55 bl[55] br[55] wl[16] vdd gnd cell_6t
Xbit_r17_c55 bl[55] br[55] wl[17] vdd gnd cell_6t
Xbit_r18_c55 bl[55] br[55] wl[18] vdd gnd cell_6t
Xbit_r19_c55 bl[55] br[55] wl[19] vdd gnd cell_6t
Xbit_r20_c55 bl[55] br[55] wl[20] vdd gnd cell_6t
Xbit_r21_c55 bl[55] br[55] wl[21] vdd gnd cell_6t
Xbit_r22_c55 bl[55] br[55] wl[22] vdd gnd cell_6t
Xbit_r23_c55 bl[55] br[55] wl[23] vdd gnd cell_6t
Xbit_r24_c55 bl[55] br[55] wl[24] vdd gnd cell_6t
Xbit_r25_c55 bl[55] br[55] wl[25] vdd gnd cell_6t
Xbit_r26_c55 bl[55] br[55] wl[26] vdd gnd cell_6t
Xbit_r27_c55 bl[55] br[55] wl[27] vdd gnd cell_6t
Xbit_r28_c55 bl[55] br[55] wl[28] vdd gnd cell_6t
Xbit_r29_c55 bl[55] br[55] wl[29] vdd gnd cell_6t
Xbit_r30_c55 bl[55] br[55] wl[30] vdd gnd cell_6t
Xbit_r31_c55 bl[55] br[55] wl[31] vdd gnd cell_6t
Xbit_r32_c55 bl[55] br[55] wl[32] vdd gnd cell_6t
Xbit_r33_c55 bl[55] br[55] wl[33] vdd gnd cell_6t
Xbit_r34_c55 bl[55] br[55] wl[34] vdd gnd cell_6t
Xbit_r35_c55 bl[55] br[55] wl[35] vdd gnd cell_6t
Xbit_r36_c55 bl[55] br[55] wl[36] vdd gnd cell_6t
Xbit_r37_c55 bl[55] br[55] wl[37] vdd gnd cell_6t
Xbit_r38_c55 bl[55] br[55] wl[38] vdd gnd cell_6t
Xbit_r39_c55 bl[55] br[55] wl[39] vdd gnd cell_6t
Xbit_r40_c55 bl[55] br[55] wl[40] vdd gnd cell_6t
Xbit_r41_c55 bl[55] br[55] wl[41] vdd gnd cell_6t
Xbit_r42_c55 bl[55] br[55] wl[42] vdd gnd cell_6t
Xbit_r43_c55 bl[55] br[55] wl[43] vdd gnd cell_6t
Xbit_r44_c55 bl[55] br[55] wl[44] vdd gnd cell_6t
Xbit_r45_c55 bl[55] br[55] wl[45] vdd gnd cell_6t
Xbit_r46_c55 bl[55] br[55] wl[46] vdd gnd cell_6t
Xbit_r47_c55 bl[55] br[55] wl[47] vdd gnd cell_6t
Xbit_r48_c55 bl[55] br[55] wl[48] vdd gnd cell_6t
Xbit_r49_c55 bl[55] br[55] wl[49] vdd gnd cell_6t
Xbit_r50_c55 bl[55] br[55] wl[50] vdd gnd cell_6t
Xbit_r51_c55 bl[55] br[55] wl[51] vdd gnd cell_6t
Xbit_r52_c55 bl[55] br[55] wl[52] vdd gnd cell_6t
Xbit_r53_c55 bl[55] br[55] wl[53] vdd gnd cell_6t
Xbit_r54_c55 bl[55] br[55] wl[54] vdd gnd cell_6t
Xbit_r55_c55 bl[55] br[55] wl[55] vdd gnd cell_6t
Xbit_r56_c55 bl[55] br[55] wl[56] vdd gnd cell_6t
Xbit_r57_c55 bl[55] br[55] wl[57] vdd gnd cell_6t
Xbit_r58_c55 bl[55] br[55] wl[58] vdd gnd cell_6t
Xbit_r59_c55 bl[55] br[55] wl[59] vdd gnd cell_6t
Xbit_r60_c55 bl[55] br[55] wl[60] vdd gnd cell_6t
Xbit_r61_c55 bl[55] br[55] wl[61] vdd gnd cell_6t
Xbit_r62_c55 bl[55] br[55] wl[62] vdd gnd cell_6t
Xbit_r63_c55 bl[55] br[55] wl[63] vdd gnd cell_6t
Xbit_r64_c55 bl[55] br[55] wl[64] vdd gnd cell_6t
Xbit_r65_c55 bl[55] br[55] wl[65] vdd gnd cell_6t
Xbit_r66_c55 bl[55] br[55] wl[66] vdd gnd cell_6t
Xbit_r67_c55 bl[55] br[55] wl[67] vdd gnd cell_6t
Xbit_r68_c55 bl[55] br[55] wl[68] vdd gnd cell_6t
Xbit_r69_c55 bl[55] br[55] wl[69] vdd gnd cell_6t
Xbit_r70_c55 bl[55] br[55] wl[70] vdd gnd cell_6t
Xbit_r71_c55 bl[55] br[55] wl[71] vdd gnd cell_6t
Xbit_r72_c55 bl[55] br[55] wl[72] vdd gnd cell_6t
Xbit_r73_c55 bl[55] br[55] wl[73] vdd gnd cell_6t
Xbit_r74_c55 bl[55] br[55] wl[74] vdd gnd cell_6t
Xbit_r75_c55 bl[55] br[55] wl[75] vdd gnd cell_6t
Xbit_r76_c55 bl[55] br[55] wl[76] vdd gnd cell_6t
Xbit_r77_c55 bl[55] br[55] wl[77] vdd gnd cell_6t
Xbit_r78_c55 bl[55] br[55] wl[78] vdd gnd cell_6t
Xbit_r79_c55 bl[55] br[55] wl[79] vdd gnd cell_6t
Xbit_r80_c55 bl[55] br[55] wl[80] vdd gnd cell_6t
Xbit_r81_c55 bl[55] br[55] wl[81] vdd gnd cell_6t
Xbit_r82_c55 bl[55] br[55] wl[82] vdd gnd cell_6t
Xbit_r83_c55 bl[55] br[55] wl[83] vdd gnd cell_6t
Xbit_r84_c55 bl[55] br[55] wl[84] vdd gnd cell_6t
Xbit_r85_c55 bl[55] br[55] wl[85] vdd gnd cell_6t
Xbit_r86_c55 bl[55] br[55] wl[86] vdd gnd cell_6t
Xbit_r87_c55 bl[55] br[55] wl[87] vdd gnd cell_6t
Xbit_r88_c55 bl[55] br[55] wl[88] vdd gnd cell_6t
Xbit_r89_c55 bl[55] br[55] wl[89] vdd gnd cell_6t
Xbit_r90_c55 bl[55] br[55] wl[90] vdd gnd cell_6t
Xbit_r91_c55 bl[55] br[55] wl[91] vdd gnd cell_6t
Xbit_r92_c55 bl[55] br[55] wl[92] vdd gnd cell_6t
Xbit_r93_c55 bl[55] br[55] wl[93] vdd gnd cell_6t
Xbit_r94_c55 bl[55] br[55] wl[94] vdd gnd cell_6t
Xbit_r95_c55 bl[55] br[55] wl[95] vdd gnd cell_6t
Xbit_r96_c55 bl[55] br[55] wl[96] vdd gnd cell_6t
Xbit_r97_c55 bl[55] br[55] wl[97] vdd gnd cell_6t
Xbit_r98_c55 bl[55] br[55] wl[98] vdd gnd cell_6t
Xbit_r99_c55 bl[55] br[55] wl[99] vdd gnd cell_6t
Xbit_r100_c55 bl[55] br[55] wl[100] vdd gnd cell_6t
Xbit_r101_c55 bl[55] br[55] wl[101] vdd gnd cell_6t
Xbit_r102_c55 bl[55] br[55] wl[102] vdd gnd cell_6t
Xbit_r103_c55 bl[55] br[55] wl[103] vdd gnd cell_6t
Xbit_r104_c55 bl[55] br[55] wl[104] vdd gnd cell_6t
Xbit_r105_c55 bl[55] br[55] wl[105] vdd gnd cell_6t
Xbit_r106_c55 bl[55] br[55] wl[106] vdd gnd cell_6t
Xbit_r107_c55 bl[55] br[55] wl[107] vdd gnd cell_6t
Xbit_r108_c55 bl[55] br[55] wl[108] vdd gnd cell_6t
Xbit_r109_c55 bl[55] br[55] wl[109] vdd gnd cell_6t
Xbit_r110_c55 bl[55] br[55] wl[110] vdd gnd cell_6t
Xbit_r111_c55 bl[55] br[55] wl[111] vdd gnd cell_6t
Xbit_r112_c55 bl[55] br[55] wl[112] vdd gnd cell_6t
Xbit_r113_c55 bl[55] br[55] wl[113] vdd gnd cell_6t
Xbit_r114_c55 bl[55] br[55] wl[114] vdd gnd cell_6t
Xbit_r115_c55 bl[55] br[55] wl[115] vdd gnd cell_6t
Xbit_r116_c55 bl[55] br[55] wl[116] vdd gnd cell_6t
Xbit_r117_c55 bl[55] br[55] wl[117] vdd gnd cell_6t
Xbit_r118_c55 bl[55] br[55] wl[118] vdd gnd cell_6t
Xbit_r119_c55 bl[55] br[55] wl[119] vdd gnd cell_6t
Xbit_r120_c55 bl[55] br[55] wl[120] vdd gnd cell_6t
Xbit_r121_c55 bl[55] br[55] wl[121] vdd gnd cell_6t
Xbit_r122_c55 bl[55] br[55] wl[122] vdd gnd cell_6t
Xbit_r123_c55 bl[55] br[55] wl[123] vdd gnd cell_6t
Xbit_r124_c55 bl[55] br[55] wl[124] vdd gnd cell_6t
Xbit_r125_c55 bl[55] br[55] wl[125] vdd gnd cell_6t
Xbit_r126_c55 bl[55] br[55] wl[126] vdd gnd cell_6t
Xbit_r127_c55 bl[55] br[55] wl[127] vdd gnd cell_6t
Xbit_r0_c56 bl[56] br[56] wl[0] vdd gnd cell_6t
Xbit_r1_c56 bl[56] br[56] wl[1] vdd gnd cell_6t
Xbit_r2_c56 bl[56] br[56] wl[2] vdd gnd cell_6t
Xbit_r3_c56 bl[56] br[56] wl[3] vdd gnd cell_6t
Xbit_r4_c56 bl[56] br[56] wl[4] vdd gnd cell_6t
Xbit_r5_c56 bl[56] br[56] wl[5] vdd gnd cell_6t
Xbit_r6_c56 bl[56] br[56] wl[6] vdd gnd cell_6t
Xbit_r7_c56 bl[56] br[56] wl[7] vdd gnd cell_6t
Xbit_r8_c56 bl[56] br[56] wl[8] vdd gnd cell_6t
Xbit_r9_c56 bl[56] br[56] wl[9] vdd gnd cell_6t
Xbit_r10_c56 bl[56] br[56] wl[10] vdd gnd cell_6t
Xbit_r11_c56 bl[56] br[56] wl[11] vdd gnd cell_6t
Xbit_r12_c56 bl[56] br[56] wl[12] vdd gnd cell_6t
Xbit_r13_c56 bl[56] br[56] wl[13] vdd gnd cell_6t
Xbit_r14_c56 bl[56] br[56] wl[14] vdd gnd cell_6t
Xbit_r15_c56 bl[56] br[56] wl[15] vdd gnd cell_6t
Xbit_r16_c56 bl[56] br[56] wl[16] vdd gnd cell_6t
Xbit_r17_c56 bl[56] br[56] wl[17] vdd gnd cell_6t
Xbit_r18_c56 bl[56] br[56] wl[18] vdd gnd cell_6t
Xbit_r19_c56 bl[56] br[56] wl[19] vdd gnd cell_6t
Xbit_r20_c56 bl[56] br[56] wl[20] vdd gnd cell_6t
Xbit_r21_c56 bl[56] br[56] wl[21] vdd gnd cell_6t
Xbit_r22_c56 bl[56] br[56] wl[22] vdd gnd cell_6t
Xbit_r23_c56 bl[56] br[56] wl[23] vdd gnd cell_6t
Xbit_r24_c56 bl[56] br[56] wl[24] vdd gnd cell_6t
Xbit_r25_c56 bl[56] br[56] wl[25] vdd gnd cell_6t
Xbit_r26_c56 bl[56] br[56] wl[26] vdd gnd cell_6t
Xbit_r27_c56 bl[56] br[56] wl[27] vdd gnd cell_6t
Xbit_r28_c56 bl[56] br[56] wl[28] vdd gnd cell_6t
Xbit_r29_c56 bl[56] br[56] wl[29] vdd gnd cell_6t
Xbit_r30_c56 bl[56] br[56] wl[30] vdd gnd cell_6t
Xbit_r31_c56 bl[56] br[56] wl[31] vdd gnd cell_6t
Xbit_r32_c56 bl[56] br[56] wl[32] vdd gnd cell_6t
Xbit_r33_c56 bl[56] br[56] wl[33] vdd gnd cell_6t
Xbit_r34_c56 bl[56] br[56] wl[34] vdd gnd cell_6t
Xbit_r35_c56 bl[56] br[56] wl[35] vdd gnd cell_6t
Xbit_r36_c56 bl[56] br[56] wl[36] vdd gnd cell_6t
Xbit_r37_c56 bl[56] br[56] wl[37] vdd gnd cell_6t
Xbit_r38_c56 bl[56] br[56] wl[38] vdd gnd cell_6t
Xbit_r39_c56 bl[56] br[56] wl[39] vdd gnd cell_6t
Xbit_r40_c56 bl[56] br[56] wl[40] vdd gnd cell_6t
Xbit_r41_c56 bl[56] br[56] wl[41] vdd gnd cell_6t
Xbit_r42_c56 bl[56] br[56] wl[42] vdd gnd cell_6t
Xbit_r43_c56 bl[56] br[56] wl[43] vdd gnd cell_6t
Xbit_r44_c56 bl[56] br[56] wl[44] vdd gnd cell_6t
Xbit_r45_c56 bl[56] br[56] wl[45] vdd gnd cell_6t
Xbit_r46_c56 bl[56] br[56] wl[46] vdd gnd cell_6t
Xbit_r47_c56 bl[56] br[56] wl[47] vdd gnd cell_6t
Xbit_r48_c56 bl[56] br[56] wl[48] vdd gnd cell_6t
Xbit_r49_c56 bl[56] br[56] wl[49] vdd gnd cell_6t
Xbit_r50_c56 bl[56] br[56] wl[50] vdd gnd cell_6t
Xbit_r51_c56 bl[56] br[56] wl[51] vdd gnd cell_6t
Xbit_r52_c56 bl[56] br[56] wl[52] vdd gnd cell_6t
Xbit_r53_c56 bl[56] br[56] wl[53] vdd gnd cell_6t
Xbit_r54_c56 bl[56] br[56] wl[54] vdd gnd cell_6t
Xbit_r55_c56 bl[56] br[56] wl[55] vdd gnd cell_6t
Xbit_r56_c56 bl[56] br[56] wl[56] vdd gnd cell_6t
Xbit_r57_c56 bl[56] br[56] wl[57] vdd gnd cell_6t
Xbit_r58_c56 bl[56] br[56] wl[58] vdd gnd cell_6t
Xbit_r59_c56 bl[56] br[56] wl[59] vdd gnd cell_6t
Xbit_r60_c56 bl[56] br[56] wl[60] vdd gnd cell_6t
Xbit_r61_c56 bl[56] br[56] wl[61] vdd gnd cell_6t
Xbit_r62_c56 bl[56] br[56] wl[62] vdd gnd cell_6t
Xbit_r63_c56 bl[56] br[56] wl[63] vdd gnd cell_6t
Xbit_r64_c56 bl[56] br[56] wl[64] vdd gnd cell_6t
Xbit_r65_c56 bl[56] br[56] wl[65] vdd gnd cell_6t
Xbit_r66_c56 bl[56] br[56] wl[66] vdd gnd cell_6t
Xbit_r67_c56 bl[56] br[56] wl[67] vdd gnd cell_6t
Xbit_r68_c56 bl[56] br[56] wl[68] vdd gnd cell_6t
Xbit_r69_c56 bl[56] br[56] wl[69] vdd gnd cell_6t
Xbit_r70_c56 bl[56] br[56] wl[70] vdd gnd cell_6t
Xbit_r71_c56 bl[56] br[56] wl[71] vdd gnd cell_6t
Xbit_r72_c56 bl[56] br[56] wl[72] vdd gnd cell_6t
Xbit_r73_c56 bl[56] br[56] wl[73] vdd gnd cell_6t
Xbit_r74_c56 bl[56] br[56] wl[74] vdd gnd cell_6t
Xbit_r75_c56 bl[56] br[56] wl[75] vdd gnd cell_6t
Xbit_r76_c56 bl[56] br[56] wl[76] vdd gnd cell_6t
Xbit_r77_c56 bl[56] br[56] wl[77] vdd gnd cell_6t
Xbit_r78_c56 bl[56] br[56] wl[78] vdd gnd cell_6t
Xbit_r79_c56 bl[56] br[56] wl[79] vdd gnd cell_6t
Xbit_r80_c56 bl[56] br[56] wl[80] vdd gnd cell_6t
Xbit_r81_c56 bl[56] br[56] wl[81] vdd gnd cell_6t
Xbit_r82_c56 bl[56] br[56] wl[82] vdd gnd cell_6t
Xbit_r83_c56 bl[56] br[56] wl[83] vdd gnd cell_6t
Xbit_r84_c56 bl[56] br[56] wl[84] vdd gnd cell_6t
Xbit_r85_c56 bl[56] br[56] wl[85] vdd gnd cell_6t
Xbit_r86_c56 bl[56] br[56] wl[86] vdd gnd cell_6t
Xbit_r87_c56 bl[56] br[56] wl[87] vdd gnd cell_6t
Xbit_r88_c56 bl[56] br[56] wl[88] vdd gnd cell_6t
Xbit_r89_c56 bl[56] br[56] wl[89] vdd gnd cell_6t
Xbit_r90_c56 bl[56] br[56] wl[90] vdd gnd cell_6t
Xbit_r91_c56 bl[56] br[56] wl[91] vdd gnd cell_6t
Xbit_r92_c56 bl[56] br[56] wl[92] vdd gnd cell_6t
Xbit_r93_c56 bl[56] br[56] wl[93] vdd gnd cell_6t
Xbit_r94_c56 bl[56] br[56] wl[94] vdd gnd cell_6t
Xbit_r95_c56 bl[56] br[56] wl[95] vdd gnd cell_6t
Xbit_r96_c56 bl[56] br[56] wl[96] vdd gnd cell_6t
Xbit_r97_c56 bl[56] br[56] wl[97] vdd gnd cell_6t
Xbit_r98_c56 bl[56] br[56] wl[98] vdd gnd cell_6t
Xbit_r99_c56 bl[56] br[56] wl[99] vdd gnd cell_6t
Xbit_r100_c56 bl[56] br[56] wl[100] vdd gnd cell_6t
Xbit_r101_c56 bl[56] br[56] wl[101] vdd gnd cell_6t
Xbit_r102_c56 bl[56] br[56] wl[102] vdd gnd cell_6t
Xbit_r103_c56 bl[56] br[56] wl[103] vdd gnd cell_6t
Xbit_r104_c56 bl[56] br[56] wl[104] vdd gnd cell_6t
Xbit_r105_c56 bl[56] br[56] wl[105] vdd gnd cell_6t
Xbit_r106_c56 bl[56] br[56] wl[106] vdd gnd cell_6t
Xbit_r107_c56 bl[56] br[56] wl[107] vdd gnd cell_6t
Xbit_r108_c56 bl[56] br[56] wl[108] vdd gnd cell_6t
Xbit_r109_c56 bl[56] br[56] wl[109] vdd gnd cell_6t
Xbit_r110_c56 bl[56] br[56] wl[110] vdd gnd cell_6t
Xbit_r111_c56 bl[56] br[56] wl[111] vdd gnd cell_6t
Xbit_r112_c56 bl[56] br[56] wl[112] vdd gnd cell_6t
Xbit_r113_c56 bl[56] br[56] wl[113] vdd gnd cell_6t
Xbit_r114_c56 bl[56] br[56] wl[114] vdd gnd cell_6t
Xbit_r115_c56 bl[56] br[56] wl[115] vdd gnd cell_6t
Xbit_r116_c56 bl[56] br[56] wl[116] vdd gnd cell_6t
Xbit_r117_c56 bl[56] br[56] wl[117] vdd gnd cell_6t
Xbit_r118_c56 bl[56] br[56] wl[118] vdd gnd cell_6t
Xbit_r119_c56 bl[56] br[56] wl[119] vdd gnd cell_6t
Xbit_r120_c56 bl[56] br[56] wl[120] vdd gnd cell_6t
Xbit_r121_c56 bl[56] br[56] wl[121] vdd gnd cell_6t
Xbit_r122_c56 bl[56] br[56] wl[122] vdd gnd cell_6t
Xbit_r123_c56 bl[56] br[56] wl[123] vdd gnd cell_6t
Xbit_r124_c56 bl[56] br[56] wl[124] vdd gnd cell_6t
Xbit_r125_c56 bl[56] br[56] wl[125] vdd gnd cell_6t
Xbit_r126_c56 bl[56] br[56] wl[126] vdd gnd cell_6t
Xbit_r127_c56 bl[56] br[56] wl[127] vdd gnd cell_6t
Xbit_r0_c57 bl[57] br[57] wl[0] vdd gnd cell_6t
Xbit_r1_c57 bl[57] br[57] wl[1] vdd gnd cell_6t
Xbit_r2_c57 bl[57] br[57] wl[2] vdd gnd cell_6t
Xbit_r3_c57 bl[57] br[57] wl[3] vdd gnd cell_6t
Xbit_r4_c57 bl[57] br[57] wl[4] vdd gnd cell_6t
Xbit_r5_c57 bl[57] br[57] wl[5] vdd gnd cell_6t
Xbit_r6_c57 bl[57] br[57] wl[6] vdd gnd cell_6t
Xbit_r7_c57 bl[57] br[57] wl[7] vdd gnd cell_6t
Xbit_r8_c57 bl[57] br[57] wl[8] vdd gnd cell_6t
Xbit_r9_c57 bl[57] br[57] wl[9] vdd gnd cell_6t
Xbit_r10_c57 bl[57] br[57] wl[10] vdd gnd cell_6t
Xbit_r11_c57 bl[57] br[57] wl[11] vdd gnd cell_6t
Xbit_r12_c57 bl[57] br[57] wl[12] vdd gnd cell_6t
Xbit_r13_c57 bl[57] br[57] wl[13] vdd gnd cell_6t
Xbit_r14_c57 bl[57] br[57] wl[14] vdd gnd cell_6t
Xbit_r15_c57 bl[57] br[57] wl[15] vdd gnd cell_6t
Xbit_r16_c57 bl[57] br[57] wl[16] vdd gnd cell_6t
Xbit_r17_c57 bl[57] br[57] wl[17] vdd gnd cell_6t
Xbit_r18_c57 bl[57] br[57] wl[18] vdd gnd cell_6t
Xbit_r19_c57 bl[57] br[57] wl[19] vdd gnd cell_6t
Xbit_r20_c57 bl[57] br[57] wl[20] vdd gnd cell_6t
Xbit_r21_c57 bl[57] br[57] wl[21] vdd gnd cell_6t
Xbit_r22_c57 bl[57] br[57] wl[22] vdd gnd cell_6t
Xbit_r23_c57 bl[57] br[57] wl[23] vdd gnd cell_6t
Xbit_r24_c57 bl[57] br[57] wl[24] vdd gnd cell_6t
Xbit_r25_c57 bl[57] br[57] wl[25] vdd gnd cell_6t
Xbit_r26_c57 bl[57] br[57] wl[26] vdd gnd cell_6t
Xbit_r27_c57 bl[57] br[57] wl[27] vdd gnd cell_6t
Xbit_r28_c57 bl[57] br[57] wl[28] vdd gnd cell_6t
Xbit_r29_c57 bl[57] br[57] wl[29] vdd gnd cell_6t
Xbit_r30_c57 bl[57] br[57] wl[30] vdd gnd cell_6t
Xbit_r31_c57 bl[57] br[57] wl[31] vdd gnd cell_6t
Xbit_r32_c57 bl[57] br[57] wl[32] vdd gnd cell_6t
Xbit_r33_c57 bl[57] br[57] wl[33] vdd gnd cell_6t
Xbit_r34_c57 bl[57] br[57] wl[34] vdd gnd cell_6t
Xbit_r35_c57 bl[57] br[57] wl[35] vdd gnd cell_6t
Xbit_r36_c57 bl[57] br[57] wl[36] vdd gnd cell_6t
Xbit_r37_c57 bl[57] br[57] wl[37] vdd gnd cell_6t
Xbit_r38_c57 bl[57] br[57] wl[38] vdd gnd cell_6t
Xbit_r39_c57 bl[57] br[57] wl[39] vdd gnd cell_6t
Xbit_r40_c57 bl[57] br[57] wl[40] vdd gnd cell_6t
Xbit_r41_c57 bl[57] br[57] wl[41] vdd gnd cell_6t
Xbit_r42_c57 bl[57] br[57] wl[42] vdd gnd cell_6t
Xbit_r43_c57 bl[57] br[57] wl[43] vdd gnd cell_6t
Xbit_r44_c57 bl[57] br[57] wl[44] vdd gnd cell_6t
Xbit_r45_c57 bl[57] br[57] wl[45] vdd gnd cell_6t
Xbit_r46_c57 bl[57] br[57] wl[46] vdd gnd cell_6t
Xbit_r47_c57 bl[57] br[57] wl[47] vdd gnd cell_6t
Xbit_r48_c57 bl[57] br[57] wl[48] vdd gnd cell_6t
Xbit_r49_c57 bl[57] br[57] wl[49] vdd gnd cell_6t
Xbit_r50_c57 bl[57] br[57] wl[50] vdd gnd cell_6t
Xbit_r51_c57 bl[57] br[57] wl[51] vdd gnd cell_6t
Xbit_r52_c57 bl[57] br[57] wl[52] vdd gnd cell_6t
Xbit_r53_c57 bl[57] br[57] wl[53] vdd gnd cell_6t
Xbit_r54_c57 bl[57] br[57] wl[54] vdd gnd cell_6t
Xbit_r55_c57 bl[57] br[57] wl[55] vdd gnd cell_6t
Xbit_r56_c57 bl[57] br[57] wl[56] vdd gnd cell_6t
Xbit_r57_c57 bl[57] br[57] wl[57] vdd gnd cell_6t
Xbit_r58_c57 bl[57] br[57] wl[58] vdd gnd cell_6t
Xbit_r59_c57 bl[57] br[57] wl[59] vdd gnd cell_6t
Xbit_r60_c57 bl[57] br[57] wl[60] vdd gnd cell_6t
Xbit_r61_c57 bl[57] br[57] wl[61] vdd gnd cell_6t
Xbit_r62_c57 bl[57] br[57] wl[62] vdd gnd cell_6t
Xbit_r63_c57 bl[57] br[57] wl[63] vdd gnd cell_6t
Xbit_r64_c57 bl[57] br[57] wl[64] vdd gnd cell_6t
Xbit_r65_c57 bl[57] br[57] wl[65] vdd gnd cell_6t
Xbit_r66_c57 bl[57] br[57] wl[66] vdd gnd cell_6t
Xbit_r67_c57 bl[57] br[57] wl[67] vdd gnd cell_6t
Xbit_r68_c57 bl[57] br[57] wl[68] vdd gnd cell_6t
Xbit_r69_c57 bl[57] br[57] wl[69] vdd gnd cell_6t
Xbit_r70_c57 bl[57] br[57] wl[70] vdd gnd cell_6t
Xbit_r71_c57 bl[57] br[57] wl[71] vdd gnd cell_6t
Xbit_r72_c57 bl[57] br[57] wl[72] vdd gnd cell_6t
Xbit_r73_c57 bl[57] br[57] wl[73] vdd gnd cell_6t
Xbit_r74_c57 bl[57] br[57] wl[74] vdd gnd cell_6t
Xbit_r75_c57 bl[57] br[57] wl[75] vdd gnd cell_6t
Xbit_r76_c57 bl[57] br[57] wl[76] vdd gnd cell_6t
Xbit_r77_c57 bl[57] br[57] wl[77] vdd gnd cell_6t
Xbit_r78_c57 bl[57] br[57] wl[78] vdd gnd cell_6t
Xbit_r79_c57 bl[57] br[57] wl[79] vdd gnd cell_6t
Xbit_r80_c57 bl[57] br[57] wl[80] vdd gnd cell_6t
Xbit_r81_c57 bl[57] br[57] wl[81] vdd gnd cell_6t
Xbit_r82_c57 bl[57] br[57] wl[82] vdd gnd cell_6t
Xbit_r83_c57 bl[57] br[57] wl[83] vdd gnd cell_6t
Xbit_r84_c57 bl[57] br[57] wl[84] vdd gnd cell_6t
Xbit_r85_c57 bl[57] br[57] wl[85] vdd gnd cell_6t
Xbit_r86_c57 bl[57] br[57] wl[86] vdd gnd cell_6t
Xbit_r87_c57 bl[57] br[57] wl[87] vdd gnd cell_6t
Xbit_r88_c57 bl[57] br[57] wl[88] vdd gnd cell_6t
Xbit_r89_c57 bl[57] br[57] wl[89] vdd gnd cell_6t
Xbit_r90_c57 bl[57] br[57] wl[90] vdd gnd cell_6t
Xbit_r91_c57 bl[57] br[57] wl[91] vdd gnd cell_6t
Xbit_r92_c57 bl[57] br[57] wl[92] vdd gnd cell_6t
Xbit_r93_c57 bl[57] br[57] wl[93] vdd gnd cell_6t
Xbit_r94_c57 bl[57] br[57] wl[94] vdd gnd cell_6t
Xbit_r95_c57 bl[57] br[57] wl[95] vdd gnd cell_6t
Xbit_r96_c57 bl[57] br[57] wl[96] vdd gnd cell_6t
Xbit_r97_c57 bl[57] br[57] wl[97] vdd gnd cell_6t
Xbit_r98_c57 bl[57] br[57] wl[98] vdd gnd cell_6t
Xbit_r99_c57 bl[57] br[57] wl[99] vdd gnd cell_6t
Xbit_r100_c57 bl[57] br[57] wl[100] vdd gnd cell_6t
Xbit_r101_c57 bl[57] br[57] wl[101] vdd gnd cell_6t
Xbit_r102_c57 bl[57] br[57] wl[102] vdd gnd cell_6t
Xbit_r103_c57 bl[57] br[57] wl[103] vdd gnd cell_6t
Xbit_r104_c57 bl[57] br[57] wl[104] vdd gnd cell_6t
Xbit_r105_c57 bl[57] br[57] wl[105] vdd gnd cell_6t
Xbit_r106_c57 bl[57] br[57] wl[106] vdd gnd cell_6t
Xbit_r107_c57 bl[57] br[57] wl[107] vdd gnd cell_6t
Xbit_r108_c57 bl[57] br[57] wl[108] vdd gnd cell_6t
Xbit_r109_c57 bl[57] br[57] wl[109] vdd gnd cell_6t
Xbit_r110_c57 bl[57] br[57] wl[110] vdd gnd cell_6t
Xbit_r111_c57 bl[57] br[57] wl[111] vdd gnd cell_6t
Xbit_r112_c57 bl[57] br[57] wl[112] vdd gnd cell_6t
Xbit_r113_c57 bl[57] br[57] wl[113] vdd gnd cell_6t
Xbit_r114_c57 bl[57] br[57] wl[114] vdd gnd cell_6t
Xbit_r115_c57 bl[57] br[57] wl[115] vdd gnd cell_6t
Xbit_r116_c57 bl[57] br[57] wl[116] vdd gnd cell_6t
Xbit_r117_c57 bl[57] br[57] wl[117] vdd gnd cell_6t
Xbit_r118_c57 bl[57] br[57] wl[118] vdd gnd cell_6t
Xbit_r119_c57 bl[57] br[57] wl[119] vdd gnd cell_6t
Xbit_r120_c57 bl[57] br[57] wl[120] vdd gnd cell_6t
Xbit_r121_c57 bl[57] br[57] wl[121] vdd gnd cell_6t
Xbit_r122_c57 bl[57] br[57] wl[122] vdd gnd cell_6t
Xbit_r123_c57 bl[57] br[57] wl[123] vdd gnd cell_6t
Xbit_r124_c57 bl[57] br[57] wl[124] vdd gnd cell_6t
Xbit_r125_c57 bl[57] br[57] wl[125] vdd gnd cell_6t
Xbit_r126_c57 bl[57] br[57] wl[126] vdd gnd cell_6t
Xbit_r127_c57 bl[57] br[57] wl[127] vdd gnd cell_6t
Xbit_r0_c58 bl[58] br[58] wl[0] vdd gnd cell_6t
Xbit_r1_c58 bl[58] br[58] wl[1] vdd gnd cell_6t
Xbit_r2_c58 bl[58] br[58] wl[2] vdd gnd cell_6t
Xbit_r3_c58 bl[58] br[58] wl[3] vdd gnd cell_6t
Xbit_r4_c58 bl[58] br[58] wl[4] vdd gnd cell_6t
Xbit_r5_c58 bl[58] br[58] wl[5] vdd gnd cell_6t
Xbit_r6_c58 bl[58] br[58] wl[6] vdd gnd cell_6t
Xbit_r7_c58 bl[58] br[58] wl[7] vdd gnd cell_6t
Xbit_r8_c58 bl[58] br[58] wl[8] vdd gnd cell_6t
Xbit_r9_c58 bl[58] br[58] wl[9] vdd gnd cell_6t
Xbit_r10_c58 bl[58] br[58] wl[10] vdd gnd cell_6t
Xbit_r11_c58 bl[58] br[58] wl[11] vdd gnd cell_6t
Xbit_r12_c58 bl[58] br[58] wl[12] vdd gnd cell_6t
Xbit_r13_c58 bl[58] br[58] wl[13] vdd gnd cell_6t
Xbit_r14_c58 bl[58] br[58] wl[14] vdd gnd cell_6t
Xbit_r15_c58 bl[58] br[58] wl[15] vdd gnd cell_6t
Xbit_r16_c58 bl[58] br[58] wl[16] vdd gnd cell_6t
Xbit_r17_c58 bl[58] br[58] wl[17] vdd gnd cell_6t
Xbit_r18_c58 bl[58] br[58] wl[18] vdd gnd cell_6t
Xbit_r19_c58 bl[58] br[58] wl[19] vdd gnd cell_6t
Xbit_r20_c58 bl[58] br[58] wl[20] vdd gnd cell_6t
Xbit_r21_c58 bl[58] br[58] wl[21] vdd gnd cell_6t
Xbit_r22_c58 bl[58] br[58] wl[22] vdd gnd cell_6t
Xbit_r23_c58 bl[58] br[58] wl[23] vdd gnd cell_6t
Xbit_r24_c58 bl[58] br[58] wl[24] vdd gnd cell_6t
Xbit_r25_c58 bl[58] br[58] wl[25] vdd gnd cell_6t
Xbit_r26_c58 bl[58] br[58] wl[26] vdd gnd cell_6t
Xbit_r27_c58 bl[58] br[58] wl[27] vdd gnd cell_6t
Xbit_r28_c58 bl[58] br[58] wl[28] vdd gnd cell_6t
Xbit_r29_c58 bl[58] br[58] wl[29] vdd gnd cell_6t
Xbit_r30_c58 bl[58] br[58] wl[30] vdd gnd cell_6t
Xbit_r31_c58 bl[58] br[58] wl[31] vdd gnd cell_6t
Xbit_r32_c58 bl[58] br[58] wl[32] vdd gnd cell_6t
Xbit_r33_c58 bl[58] br[58] wl[33] vdd gnd cell_6t
Xbit_r34_c58 bl[58] br[58] wl[34] vdd gnd cell_6t
Xbit_r35_c58 bl[58] br[58] wl[35] vdd gnd cell_6t
Xbit_r36_c58 bl[58] br[58] wl[36] vdd gnd cell_6t
Xbit_r37_c58 bl[58] br[58] wl[37] vdd gnd cell_6t
Xbit_r38_c58 bl[58] br[58] wl[38] vdd gnd cell_6t
Xbit_r39_c58 bl[58] br[58] wl[39] vdd gnd cell_6t
Xbit_r40_c58 bl[58] br[58] wl[40] vdd gnd cell_6t
Xbit_r41_c58 bl[58] br[58] wl[41] vdd gnd cell_6t
Xbit_r42_c58 bl[58] br[58] wl[42] vdd gnd cell_6t
Xbit_r43_c58 bl[58] br[58] wl[43] vdd gnd cell_6t
Xbit_r44_c58 bl[58] br[58] wl[44] vdd gnd cell_6t
Xbit_r45_c58 bl[58] br[58] wl[45] vdd gnd cell_6t
Xbit_r46_c58 bl[58] br[58] wl[46] vdd gnd cell_6t
Xbit_r47_c58 bl[58] br[58] wl[47] vdd gnd cell_6t
Xbit_r48_c58 bl[58] br[58] wl[48] vdd gnd cell_6t
Xbit_r49_c58 bl[58] br[58] wl[49] vdd gnd cell_6t
Xbit_r50_c58 bl[58] br[58] wl[50] vdd gnd cell_6t
Xbit_r51_c58 bl[58] br[58] wl[51] vdd gnd cell_6t
Xbit_r52_c58 bl[58] br[58] wl[52] vdd gnd cell_6t
Xbit_r53_c58 bl[58] br[58] wl[53] vdd gnd cell_6t
Xbit_r54_c58 bl[58] br[58] wl[54] vdd gnd cell_6t
Xbit_r55_c58 bl[58] br[58] wl[55] vdd gnd cell_6t
Xbit_r56_c58 bl[58] br[58] wl[56] vdd gnd cell_6t
Xbit_r57_c58 bl[58] br[58] wl[57] vdd gnd cell_6t
Xbit_r58_c58 bl[58] br[58] wl[58] vdd gnd cell_6t
Xbit_r59_c58 bl[58] br[58] wl[59] vdd gnd cell_6t
Xbit_r60_c58 bl[58] br[58] wl[60] vdd gnd cell_6t
Xbit_r61_c58 bl[58] br[58] wl[61] vdd gnd cell_6t
Xbit_r62_c58 bl[58] br[58] wl[62] vdd gnd cell_6t
Xbit_r63_c58 bl[58] br[58] wl[63] vdd gnd cell_6t
Xbit_r64_c58 bl[58] br[58] wl[64] vdd gnd cell_6t
Xbit_r65_c58 bl[58] br[58] wl[65] vdd gnd cell_6t
Xbit_r66_c58 bl[58] br[58] wl[66] vdd gnd cell_6t
Xbit_r67_c58 bl[58] br[58] wl[67] vdd gnd cell_6t
Xbit_r68_c58 bl[58] br[58] wl[68] vdd gnd cell_6t
Xbit_r69_c58 bl[58] br[58] wl[69] vdd gnd cell_6t
Xbit_r70_c58 bl[58] br[58] wl[70] vdd gnd cell_6t
Xbit_r71_c58 bl[58] br[58] wl[71] vdd gnd cell_6t
Xbit_r72_c58 bl[58] br[58] wl[72] vdd gnd cell_6t
Xbit_r73_c58 bl[58] br[58] wl[73] vdd gnd cell_6t
Xbit_r74_c58 bl[58] br[58] wl[74] vdd gnd cell_6t
Xbit_r75_c58 bl[58] br[58] wl[75] vdd gnd cell_6t
Xbit_r76_c58 bl[58] br[58] wl[76] vdd gnd cell_6t
Xbit_r77_c58 bl[58] br[58] wl[77] vdd gnd cell_6t
Xbit_r78_c58 bl[58] br[58] wl[78] vdd gnd cell_6t
Xbit_r79_c58 bl[58] br[58] wl[79] vdd gnd cell_6t
Xbit_r80_c58 bl[58] br[58] wl[80] vdd gnd cell_6t
Xbit_r81_c58 bl[58] br[58] wl[81] vdd gnd cell_6t
Xbit_r82_c58 bl[58] br[58] wl[82] vdd gnd cell_6t
Xbit_r83_c58 bl[58] br[58] wl[83] vdd gnd cell_6t
Xbit_r84_c58 bl[58] br[58] wl[84] vdd gnd cell_6t
Xbit_r85_c58 bl[58] br[58] wl[85] vdd gnd cell_6t
Xbit_r86_c58 bl[58] br[58] wl[86] vdd gnd cell_6t
Xbit_r87_c58 bl[58] br[58] wl[87] vdd gnd cell_6t
Xbit_r88_c58 bl[58] br[58] wl[88] vdd gnd cell_6t
Xbit_r89_c58 bl[58] br[58] wl[89] vdd gnd cell_6t
Xbit_r90_c58 bl[58] br[58] wl[90] vdd gnd cell_6t
Xbit_r91_c58 bl[58] br[58] wl[91] vdd gnd cell_6t
Xbit_r92_c58 bl[58] br[58] wl[92] vdd gnd cell_6t
Xbit_r93_c58 bl[58] br[58] wl[93] vdd gnd cell_6t
Xbit_r94_c58 bl[58] br[58] wl[94] vdd gnd cell_6t
Xbit_r95_c58 bl[58] br[58] wl[95] vdd gnd cell_6t
Xbit_r96_c58 bl[58] br[58] wl[96] vdd gnd cell_6t
Xbit_r97_c58 bl[58] br[58] wl[97] vdd gnd cell_6t
Xbit_r98_c58 bl[58] br[58] wl[98] vdd gnd cell_6t
Xbit_r99_c58 bl[58] br[58] wl[99] vdd gnd cell_6t
Xbit_r100_c58 bl[58] br[58] wl[100] vdd gnd cell_6t
Xbit_r101_c58 bl[58] br[58] wl[101] vdd gnd cell_6t
Xbit_r102_c58 bl[58] br[58] wl[102] vdd gnd cell_6t
Xbit_r103_c58 bl[58] br[58] wl[103] vdd gnd cell_6t
Xbit_r104_c58 bl[58] br[58] wl[104] vdd gnd cell_6t
Xbit_r105_c58 bl[58] br[58] wl[105] vdd gnd cell_6t
Xbit_r106_c58 bl[58] br[58] wl[106] vdd gnd cell_6t
Xbit_r107_c58 bl[58] br[58] wl[107] vdd gnd cell_6t
Xbit_r108_c58 bl[58] br[58] wl[108] vdd gnd cell_6t
Xbit_r109_c58 bl[58] br[58] wl[109] vdd gnd cell_6t
Xbit_r110_c58 bl[58] br[58] wl[110] vdd gnd cell_6t
Xbit_r111_c58 bl[58] br[58] wl[111] vdd gnd cell_6t
Xbit_r112_c58 bl[58] br[58] wl[112] vdd gnd cell_6t
Xbit_r113_c58 bl[58] br[58] wl[113] vdd gnd cell_6t
Xbit_r114_c58 bl[58] br[58] wl[114] vdd gnd cell_6t
Xbit_r115_c58 bl[58] br[58] wl[115] vdd gnd cell_6t
Xbit_r116_c58 bl[58] br[58] wl[116] vdd gnd cell_6t
Xbit_r117_c58 bl[58] br[58] wl[117] vdd gnd cell_6t
Xbit_r118_c58 bl[58] br[58] wl[118] vdd gnd cell_6t
Xbit_r119_c58 bl[58] br[58] wl[119] vdd gnd cell_6t
Xbit_r120_c58 bl[58] br[58] wl[120] vdd gnd cell_6t
Xbit_r121_c58 bl[58] br[58] wl[121] vdd gnd cell_6t
Xbit_r122_c58 bl[58] br[58] wl[122] vdd gnd cell_6t
Xbit_r123_c58 bl[58] br[58] wl[123] vdd gnd cell_6t
Xbit_r124_c58 bl[58] br[58] wl[124] vdd gnd cell_6t
Xbit_r125_c58 bl[58] br[58] wl[125] vdd gnd cell_6t
Xbit_r126_c58 bl[58] br[58] wl[126] vdd gnd cell_6t
Xbit_r127_c58 bl[58] br[58] wl[127] vdd gnd cell_6t
Xbit_r0_c59 bl[59] br[59] wl[0] vdd gnd cell_6t
Xbit_r1_c59 bl[59] br[59] wl[1] vdd gnd cell_6t
Xbit_r2_c59 bl[59] br[59] wl[2] vdd gnd cell_6t
Xbit_r3_c59 bl[59] br[59] wl[3] vdd gnd cell_6t
Xbit_r4_c59 bl[59] br[59] wl[4] vdd gnd cell_6t
Xbit_r5_c59 bl[59] br[59] wl[5] vdd gnd cell_6t
Xbit_r6_c59 bl[59] br[59] wl[6] vdd gnd cell_6t
Xbit_r7_c59 bl[59] br[59] wl[7] vdd gnd cell_6t
Xbit_r8_c59 bl[59] br[59] wl[8] vdd gnd cell_6t
Xbit_r9_c59 bl[59] br[59] wl[9] vdd gnd cell_6t
Xbit_r10_c59 bl[59] br[59] wl[10] vdd gnd cell_6t
Xbit_r11_c59 bl[59] br[59] wl[11] vdd gnd cell_6t
Xbit_r12_c59 bl[59] br[59] wl[12] vdd gnd cell_6t
Xbit_r13_c59 bl[59] br[59] wl[13] vdd gnd cell_6t
Xbit_r14_c59 bl[59] br[59] wl[14] vdd gnd cell_6t
Xbit_r15_c59 bl[59] br[59] wl[15] vdd gnd cell_6t
Xbit_r16_c59 bl[59] br[59] wl[16] vdd gnd cell_6t
Xbit_r17_c59 bl[59] br[59] wl[17] vdd gnd cell_6t
Xbit_r18_c59 bl[59] br[59] wl[18] vdd gnd cell_6t
Xbit_r19_c59 bl[59] br[59] wl[19] vdd gnd cell_6t
Xbit_r20_c59 bl[59] br[59] wl[20] vdd gnd cell_6t
Xbit_r21_c59 bl[59] br[59] wl[21] vdd gnd cell_6t
Xbit_r22_c59 bl[59] br[59] wl[22] vdd gnd cell_6t
Xbit_r23_c59 bl[59] br[59] wl[23] vdd gnd cell_6t
Xbit_r24_c59 bl[59] br[59] wl[24] vdd gnd cell_6t
Xbit_r25_c59 bl[59] br[59] wl[25] vdd gnd cell_6t
Xbit_r26_c59 bl[59] br[59] wl[26] vdd gnd cell_6t
Xbit_r27_c59 bl[59] br[59] wl[27] vdd gnd cell_6t
Xbit_r28_c59 bl[59] br[59] wl[28] vdd gnd cell_6t
Xbit_r29_c59 bl[59] br[59] wl[29] vdd gnd cell_6t
Xbit_r30_c59 bl[59] br[59] wl[30] vdd gnd cell_6t
Xbit_r31_c59 bl[59] br[59] wl[31] vdd gnd cell_6t
Xbit_r32_c59 bl[59] br[59] wl[32] vdd gnd cell_6t
Xbit_r33_c59 bl[59] br[59] wl[33] vdd gnd cell_6t
Xbit_r34_c59 bl[59] br[59] wl[34] vdd gnd cell_6t
Xbit_r35_c59 bl[59] br[59] wl[35] vdd gnd cell_6t
Xbit_r36_c59 bl[59] br[59] wl[36] vdd gnd cell_6t
Xbit_r37_c59 bl[59] br[59] wl[37] vdd gnd cell_6t
Xbit_r38_c59 bl[59] br[59] wl[38] vdd gnd cell_6t
Xbit_r39_c59 bl[59] br[59] wl[39] vdd gnd cell_6t
Xbit_r40_c59 bl[59] br[59] wl[40] vdd gnd cell_6t
Xbit_r41_c59 bl[59] br[59] wl[41] vdd gnd cell_6t
Xbit_r42_c59 bl[59] br[59] wl[42] vdd gnd cell_6t
Xbit_r43_c59 bl[59] br[59] wl[43] vdd gnd cell_6t
Xbit_r44_c59 bl[59] br[59] wl[44] vdd gnd cell_6t
Xbit_r45_c59 bl[59] br[59] wl[45] vdd gnd cell_6t
Xbit_r46_c59 bl[59] br[59] wl[46] vdd gnd cell_6t
Xbit_r47_c59 bl[59] br[59] wl[47] vdd gnd cell_6t
Xbit_r48_c59 bl[59] br[59] wl[48] vdd gnd cell_6t
Xbit_r49_c59 bl[59] br[59] wl[49] vdd gnd cell_6t
Xbit_r50_c59 bl[59] br[59] wl[50] vdd gnd cell_6t
Xbit_r51_c59 bl[59] br[59] wl[51] vdd gnd cell_6t
Xbit_r52_c59 bl[59] br[59] wl[52] vdd gnd cell_6t
Xbit_r53_c59 bl[59] br[59] wl[53] vdd gnd cell_6t
Xbit_r54_c59 bl[59] br[59] wl[54] vdd gnd cell_6t
Xbit_r55_c59 bl[59] br[59] wl[55] vdd gnd cell_6t
Xbit_r56_c59 bl[59] br[59] wl[56] vdd gnd cell_6t
Xbit_r57_c59 bl[59] br[59] wl[57] vdd gnd cell_6t
Xbit_r58_c59 bl[59] br[59] wl[58] vdd gnd cell_6t
Xbit_r59_c59 bl[59] br[59] wl[59] vdd gnd cell_6t
Xbit_r60_c59 bl[59] br[59] wl[60] vdd gnd cell_6t
Xbit_r61_c59 bl[59] br[59] wl[61] vdd gnd cell_6t
Xbit_r62_c59 bl[59] br[59] wl[62] vdd gnd cell_6t
Xbit_r63_c59 bl[59] br[59] wl[63] vdd gnd cell_6t
Xbit_r64_c59 bl[59] br[59] wl[64] vdd gnd cell_6t
Xbit_r65_c59 bl[59] br[59] wl[65] vdd gnd cell_6t
Xbit_r66_c59 bl[59] br[59] wl[66] vdd gnd cell_6t
Xbit_r67_c59 bl[59] br[59] wl[67] vdd gnd cell_6t
Xbit_r68_c59 bl[59] br[59] wl[68] vdd gnd cell_6t
Xbit_r69_c59 bl[59] br[59] wl[69] vdd gnd cell_6t
Xbit_r70_c59 bl[59] br[59] wl[70] vdd gnd cell_6t
Xbit_r71_c59 bl[59] br[59] wl[71] vdd gnd cell_6t
Xbit_r72_c59 bl[59] br[59] wl[72] vdd gnd cell_6t
Xbit_r73_c59 bl[59] br[59] wl[73] vdd gnd cell_6t
Xbit_r74_c59 bl[59] br[59] wl[74] vdd gnd cell_6t
Xbit_r75_c59 bl[59] br[59] wl[75] vdd gnd cell_6t
Xbit_r76_c59 bl[59] br[59] wl[76] vdd gnd cell_6t
Xbit_r77_c59 bl[59] br[59] wl[77] vdd gnd cell_6t
Xbit_r78_c59 bl[59] br[59] wl[78] vdd gnd cell_6t
Xbit_r79_c59 bl[59] br[59] wl[79] vdd gnd cell_6t
Xbit_r80_c59 bl[59] br[59] wl[80] vdd gnd cell_6t
Xbit_r81_c59 bl[59] br[59] wl[81] vdd gnd cell_6t
Xbit_r82_c59 bl[59] br[59] wl[82] vdd gnd cell_6t
Xbit_r83_c59 bl[59] br[59] wl[83] vdd gnd cell_6t
Xbit_r84_c59 bl[59] br[59] wl[84] vdd gnd cell_6t
Xbit_r85_c59 bl[59] br[59] wl[85] vdd gnd cell_6t
Xbit_r86_c59 bl[59] br[59] wl[86] vdd gnd cell_6t
Xbit_r87_c59 bl[59] br[59] wl[87] vdd gnd cell_6t
Xbit_r88_c59 bl[59] br[59] wl[88] vdd gnd cell_6t
Xbit_r89_c59 bl[59] br[59] wl[89] vdd gnd cell_6t
Xbit_r90_c59 bl[59] br[59] wl[90] vdd gnd cell_6t
Xbit_r91_c59 bl[59] br[59] wl[91] vdd gnd cell_6t
Xbit_r92_c59 bl[59] br[59] wl[92] vdd gnd cell_6t
Xbit_r93_c59 bl[59] br[59] wl[93] vdd gnd cell_6t
Xbit_r94_c59 bl[59] br[59] wl[94] vdd gnd cell_6t
Xbit_r95_c59 bl[59] br[59] wl[95] vdd gnd cell_6t
Xbit_r96_c59 bl[59] br[59] wl[96] vdd gnd cell_6t
Xbit_r97_c59 bl[59] br[59] wl[97] vdd gnd cell_6t
Xbit_r98_c59 bl[59] br[59] wl[98] vdd gnd cell_6t
Xbit_r99_c59 bl[59] br[59] wl[99] vdd gnd cell_6t
Xbit_r100_c59 bl[59] br[59] wl[100] vdd gnd cell_6t
Xbit_r101_c59 bl[59] br[59] wl[101] vdd gnd cell_6t
Xbit_r102_c59 bl[59] br[59] wl[102] vdd gnd cell_6t
Xbit_r103_c59 bl[59] br[59] wl[103] vdd gnd cell_6t
Xbit_r104_c59 bl[59] br[59] wl[104] vdd gnd cell_6t
Xbit_r105_c59 bl[59] br[59] wl[105] vdd gnd cell_6t
Xbit_r106_c59 bl[59] br[59] wl[106] vdd gnd cell_6t
Xbit_r107_c59 bl[59] br[59] wl[107] vdd gnd cell_6t
Xbit_r108_c59 bl[59] br[59] wl[108] vdd gnd cell_6t
Xbit_r109_c59 bl[59] br[59] wl[109] vdd gnd cell_6t
Xbit_r110_c59 bl[59] br[59] wl[110] vdd gnd cell_6t
Xbit_r111_c59 bl[59] br[59] wl[111] vdd gnd cell_6t
Xbit_r112_c59 bl[59] br[59] wl[112] vdd gnd cell_6t
Xbit_r113_c59 bl[59] br[59] wl[113] vdd gnd cell_6t
Xbit_r114_c59 bl[59] br[59] wl[114] vdd gnd cell_6t
Xbit_r115_c59 bl[59] br[59] wl[115] vdd gnd cell_6t
Xbit_r116_c59 bl[59] br[59] wl[116] vdd gnd cell_6t
Xbit_r117_c59 bl[59] br[59] wl[117] vdd gnd cell_6t
Xbit_r118_c59 bl[59] br[59] wl[118] vdd gnd cell_6t
Xbit_r119_c59 bl[59] br[59] wl[119] vdd gnd cell_6t
Xbit_r120_c59 bl[59] br[59] wl[120] vdd gnd cell_6t
Xbit_r121_c59 bl[59] br[59] wl[121] vdd gnd cell_6t
Xbit_r122_c59 bl[59] br[59] wl[122] vdd gnd cell_6t
Xbit_r123_c59 bl[59] br[59] wl[123] vdd gnd cell_6t
Xbit_r124_c59 bl[59] br[59] wl[124] vdd gnd cell_6t
Xbit_r125_c59 bl[59] br[59] wl[125] vdd gnd cell_6t
Xbit_r126_c59 bl[59] br[59] wl[126] vdd gnd cell_6t
Xbit_r127_c59 bl[59] br[59] wl[127] vdd gnd cell_6t
Xbit_r0_c60 bl[60] br[60] wl[0] vdd gnd cell_6t
Xbit_r1_c60 bl[60] br[60] wl[1] vdd gnd cell_6t
Xbit_r2_c60 bl[60] br[60] wl[2] vdd gnd cell_6t
Xbit_r3_c60 bl[60] br[60] wl[3] vdd gnd cell_6t
Xbit_r4_c60 bl[60] br[60] wl[4] vdd gnd cell_6t
Xbit_r5_c60 bl[60] br[60] wl[5] vdd gnd cell_6t
Xbit_r6_c60 bl[60] br[60] wl[6] vdd gnd cell_6t
Xbit_r7_c60 bl[60] br[60] wl[7] vdd gnd cell_6t
Xbit_r8_c60 bl[60] br[60] wl[8] vdd gnd cell_6t
Xbit_r9_c60 bl[60] br[60] wl[9] vdd gnd cell_6t
Xbit_r10_c60 bl[60] br[60] wl[10] vdd gnd cell_6t
Xbit_r11_c60 bl[60] br[60] wl[11] vdd gnd cell_6t
Xbit_r12_c60 bl[60] br[60] wl[12] vdd gnd cell_6t
Xbit_r13_c60 bl[60] br[60] wl[13] vdd gnd cell_6t
Xbit_r14_c60 bl[60] br[60] wl[14] vdd gnd cell_6t
Xbit_r15_c60 bl[60] br[60] wl[15] vdd gnd cell_6t
Xbit_r16_c60 bl[60] br[60] wl[16] vdd gnd cell_6t
Xbit_r17_c60 bl[60] br[60] wl[17] vdd gnd cell_6t
Xbit_r18_c60 bl[60] br[60] wl[18] vdd gnd cell_6t
Xbit_r19_c60 bl[60] br[60] wl[19] vdd gnd cell_6t
Xbit_r20_c60 bl[60] br[60] wl[20] vdd gnd cell_6t
Xbit_r21_c60 bl[60] br[60] wl[21] vdd gnd cell_6t
Xbit_r22_c60 bl[60] br[60] wl[22] vdd gnd cell_6t
Xbit_r23_c60 bl[60] br[60] wl[23] vdd gnd cell_6t
Xbit_r24_c60 bl[60] br[60] wl[24] vdd gnd cell_6t
Xbit_r25_c60 bl[60] br[60] wl[25] vdd gnd cell_6t
Xbit_r26_c60 bl[60] br[60] wl[26] vdd gnd cell_6t
Xbit_r27_c60 bl[60] br[60] wl[27] vdd gnd cell_6t
Xbit_r28_c60 bl[60] br[60] wl[28] vdd gnd cell_6t
Xbit_r29_c60 bl[60] br[60] wl[29] vdd gnd cell_6t
Xbit_r30_c60 bl[60] br[60] wl[30] vdd gnd cell_6t
Xbit_r31_c60 bl[60] br[60] wl[31] vdd gnd cell_6t
Xbit_r32_c60 bl[60] br[60] wl[32] vdd gnd cell_6t
Xbit_r33_c60 bl[60] br[60] wl[33] vdd gnd cell_6t
Xbit_r34_c60 bl[60] br[60] wl[34] vdd gnd cell_6t
Xbit_r35_c60 bl[60] br[60] wl[35] vdd gnd cell_6t
Xbit_r36_c60 bl[60] br[60] wl[36] vdd gnd cell_6t
Xbit_r37_c60 bl[60] br[60] wl[37] vdd gnd cell_6t
Xbit_r38_c60 bl[60] br[60] wl[38] vdd gnd cell_6t
Xbit_r39_c60 bl[60] br[60] wl[39] vdd gnd cell_6t
Xbit_r40_c60 bl[60] br[60] wl[40] vdd gnd cell_6t
Xbit_r41_c60 bl[60] br[60] wl[41] vdd gnd cell_6t
Xbit_r42_c60 bl[60] br[60] wl[42] vdd gnd cell_6t
Xbit_r43_c60 bl[60] br[60] wl[43] vdd gnd cell_6t
Xbit_r44_c60 bl[60] br[60] wl[44] vdd gnd cell_6t
Xbit_r45_c60 bl[60] br[60] wl[45] vdd gnd cell_6t
Xbit_r46_c60 bl[60] br[60] wl[46] vdd gnd cell_6t
Xbit_r47_c60 bl[60] br[60] wl[47] vdd gnd cell_6t
Xbit_r48_c60 bl[60] br[60] wl[48] vdd gnd cell_6t
Xbit_r49_c60 bl[60] br[60] wl[49] vdd gnd cell_6t
Xbit_r50_c60 bl[60] br[60] wl[50] vdd gnd cell_6t
Xbit_r51_c60 bl[60] br[60] wl[51] vdd gnd cell_6t
Xbit_r52_c60 bl[60] br[60] wl[52] vdd gnd cell_6t
Xbit_r53_c60 bl[60] br[60] wl[53] vdd gnd cell_6t
Xbit_r54_c60 bl[60] br[60] wl[54] vdd gnd cell_6t
Xbit_r55_c60 bl[60] br[60] wl[55] vdd gnd cell_6t
Xbit_r56_c60 bl[60] br[60] wl[56] vdd gnd cell_6t
Xbit_r57_c60 bl[60] br[60] wl[57] vdd gnd cell_6t
Xbit_r58_c60 bl[60] br[60] wl[58] vdd gnd cell_6t
Xbit_r59_c60 bl[60] br[60] wl[59] vdd gnd cell_6t
Xbit_r60_c60 bl[60] br[60] wl[60] vdd gnd cell_6t
Xbit_r61_c60 bl[60] br[60] wl[61] vdd gnd cell_6t
Xbit_r62_c60 bl[60] br[60] wl[62] vdd gnd cell_6t
Xbit_r63_c60 bl[60] br[60] wl[63] vdd gnd cell_6t
Xbit_r64_c60 bl[60] br[60] wl[64] vdd gnd cell_6t
Xbit_r65_c60 bl[60] br[60] wl[65] vdd gnd cell_6t
Xbit_r66_c60 bl[60] br[60] wl[66] vdd gnd cell_6t
Xbit_r67_c60 bl[60] br[60] wl[67] vdd gnd cell_6t
Xbit_r68_c60 bl[60] br[60] wl[68] vdd gnd cell_6t
Xbit_r69_c60 bl[60] br[60] wl[69] vdd gnd cell_6t
Xbit_r70_c60 bl[60] br[60] wl[70] vdd gnd cell_6t
Xbit_r71_c60 bl[60] br[60] wl[71] vdd gnd cell_6t
Xbit_r72_c60 bl[60] br[60] wl[72] vdd gnd cell_6t
Xbit_r73_c60 bl[60] br[60] wl[73] vdd gnd cell_6t
Xbit_r74_c60 bl[60] br[60] wl[74] vdd gnd cell_6t
Xbit_r75_c60 bl[60] br[60] wl[75] vdd gnd cell_6t
Xbit_r76_c60 bl[60] br[60] wl[76] vdd gnd cell_6t
Xbit_r77_c60 bl[60] br[60] wl[77] vdd gnd cell_6t
Xbit_r78_c60 bl[60] br[60] wl[78] vdd gnd cell_6t
Xbit_r79_c60 bl[60] br[60] wl[79] vdd gnd cell_6t
Xbit_r80_c60 bl[60] br[60] wl[80] vdd gnd cell_6t
Xbit_r81_c60 bl[60] br[60] wl[81] vdd gnd cell_6t
Xbit_r82_c60 bl[60] br[60] wl[82] vdd gnd cell_6t
Xbit_r83_c60 bl[60] br[60] wl[83] vdd gnd cell_6t
Xbit_r84_c60 bl[60] br[60] wl[84] vdd gnd cell_6t
Xbit_r85_c60 bl[60] br[60] wl[85] vdd gnd cell_6t
Xbit_r86_c60 bl[60] br[60] wl[86] vdd gnd cell_6t
Xbit_r87_c60 bl[60] br[60] wl[87] vdd gnd cell_6t
Xbit_r88_c60 bl[60] br[60] wl[88] vdd gnd cell_6t
Xbit_r89_c60 bl[60] br[60] wl[89] vdd gnd cell_6t
Xbit_r90_c60 bl[60] br[60] wl[90] vdd gnd cell_6t
Xbit_r91_c60 bl[60] br[60] wl[91] vdd gnd cell_6t
Xbit_r92_c60 bl[60] br[60] wl[92] vdd gnd cell_6t
Xbit_r93_c60 bl[60] br[60] wl[93] vdd gnd cell_6t
Xbit_r94_c60 bl[60] br[60] wl[94] vdd gnd cell_6t
Xbit_r95_c60 bl[60] br[60] wl[95] vdd gnd cell_6t
Xbit_r96_c60 bl[60] br[60] wl[96] vdd gnd cell_6t
Xbit_r97_c60 bl[60] br[60] wl[97] vdd gnd cell_6t
Xbit_r98_c60 bl[60] br[60] wl[98] vdd gnd cell_6t
Xbit_r99_c60 bl[60] br[60] wl[99] vdd gnd cell_6t
Xbit_r100_c60 bl[60] br[60] wl[100] vdd gnd cell_6t
Xbit_r101_c60 bl[60] br[60] wl[101] vdd gnd cell_6t
Xbit_r102_c60 bl[60] br[60] wl[102] vdd gnd cell_6t
Xbit_r103_c60 bl[60] br[60] wl[103] vdd gnd cell_6t
Xbit_r104_c60 bl[60] br[60] wl[104] vdd gnd cell_6t
Xbit_r105_c60 bl[60] br[60] wl[105] vdd gnd cell_6t
Xbit_r106_c60 bl[60] br[60] wl[106] vdd gnd cell_6t
Xbit_r107_c60 bl[60] br[60] wl[107] vdd gnd cell_6t
Xbit_r108_c60 bl[60] br[60] wl[108] vdd gnd cell_6t
Xbit_r109_c60 bl[60] br[60] wl[109] vdd gnd cell_6t
Xbit_r110_c60 bl[60] br[60] wl[110] vdd gnd cell_6t
Xbit_r111_c60 bl[60] br[60] wl[111] vdd gnd cell_6t
Xbit_r112_c60 bl[60] br[60] wl[112] vdd gnd cell_6t
Xbit_r113_c60 bl[60] br[60] wl[113] vdd gnd cell_6t
Xbit_r114_c60 bl[60] br[60] wl[114] vdd gnd cell_6t
Xbit_r115_c60 bl[60] br[60] wl[115] vdd gnd cell_6t
Xbit_r116_c60 bl[60] br[60] wl[116] vdd gnd cell_6t
Xbit_r117_c60 bl[60] br[60] wl[117] vdd gnd cell_6t
Xbit_r118_c60 bl[60] br[60] wl[118] vdd gnd cell_6t
Xbit_r119_c60 bl[60] br[60] wl[119] vdd gnd cell_6t
Xbit_r120_c60 bl[60] br[60] wl[120] vdd gnd cell_6t
Xbit_r121_c60 bl[60] br[60] wl[121] vdd gnd cell_6t
Xbit_r122_c60 bl[60] br[60] wl[122] vdd gnd cell_6t
Xbit_r123_c60 bl[60] br[60] wl[123] vdd gnd cell_6t
Xbit_r124_c60 bl[60] br[60] wl[124] vdd gnd cell_6t
Xbit_r125_c60 bl[60] br[60] wl[125] vdd gnd cell_6t
Xbit_r126_c60 bl[60] br[60] wl[126] vdd gnd cell_6t
Xbit_r127_c60 bl[60] br[60] wl[127] vdd gnd cell_6t
Xbit_r0_c61 bl[61] br[61] wl[0] vdd gnd cell_6t
Xbit_r1_c61 bl[61] br[61] wl[1] vdd gnd cell_6t
Xbit_r2_c61 bl[61] br[61] wl[2] vdd gnd cell_6t
Xbit_r3_c61 bl[61] br[61] wl[3] vdd gnd cell_6t
Xbit_r4_c61 bl[61] br[61] wl[4] vdd gnd cell_6t
Xbit_r5_c61 bl[61] br[61] wl[5] vdd gnd cell_6t
Xbit_r6_c61 bl[61] br[61] wl[6] vdd gnd cell_6t
Xbit_r7_c61 bl[61] br[61] wl[7] vdd gnd cell_6t
Xbit_r8_c61 bl[61] br[61] wl[8] vdd gnd cell_6t
Xbit_r9_c61 bl[61] br[61] wl[9] vdd gnd cell_6t
Xbit_r10_c61 bl[61] br[61] wl[10] vdd gnd cell_6t
Xbit_r11_c61 bl[61] br[61] wl[11] vdd gnd cell_6t
Xbit_r12_c61 bl[61] br[61] wl[12] vdd gnd cell_6t
Xbit_r13_c61 bl[61] br[61] wl[13] vdd gnd cell_6t
Xbit_r14_c61 bl[61] br[61] wl[14] vdd gnd cell_6t
Xbit_r15_c61 bl[61] br[61] wl[15] vdd gnd cell_6t
Xbit_r16_c61 bl[61] br[61] wl[16] vdd gnd cell_6t
Xbit_r17_c61 bl[61] br[61] wl[17] vdd gnd cell_6t
Xbit_r18_c61 bl[61] br[61] wl[18] vdd gnd cell_6t
Xbit_r19_c61 bl[61] br[61] wl[19] vdd gnd cell_6t
Xbit_r20_c61 bl[61] br[61] wl[20] vdd gnd cell_6t
Xbit_r21_c61 bl[61] br[61] wl[21] vdd gnd cell_6t
Xbit_r22_c61 bl[61] br[61] wl[22] vdd gnd cell_6t
Xbit_r23_c61 bl[61] br[61] wl[23] vdd gnd cell_6t
Xbit_r24_c61 bl[61] br[61] wl[24] vdd gnd cell_6t
Xbit_r25_c61 bl[61] br[61] wl[25] vdd gnd cell_6t
Xbit_r26_c61 bl[61] br[61] wl[26] vdd gnd cell_6t
Xbit_r27_c61 bl[61] br[61] wl[27] vdd gnd cell_6t
Xbit_r28_c61 bl[61] br[61] wl[28] vdd gnd cell_6t
Xbit_r29_c61 bl[61] br[61] wl[29] vdd gnd cell_6t
Xbit_r30_c61 bl[61] br[61] wl[30] vdd gnd cell_6t
Xbit_r31_c61 bl[61] br[61] wl[31] vdd gnd cell_6t
Xbit_r32_c61 bl[61] br[61] wl[32] vdd gnd cell_6t
Xbit_r33_c61 bl[61] br[61] wl[33] vdd gnd cell_6t
Xbit_r34_c61 bl[61] br[61] wl[34] vdd gnd cell_6t
Xbit_r35_c61 bl[61] br[61] wl[35] vdd gnd cell_6t
Xbit_r36_c61 bl[61] br[61] wl[36] vdd gnd cell_6t
Xbit_r37_c61 bl[61] br[61] wl[37] vdd gnd cell_6t
Xbit_r38_c61 bl[61] br[61] wl[38] vdd gnd cell_6t
Xbit_r39_c61 bl[61] br[61] wl[39] vdd gnd cell_6t
Xbit_r40_c61 bl[61] br[61] wl[40] vdd gnd cell_6t
Xbit_r41_c61 bl[61] br[61] wl[41] vdd gnd cell_6t
Xbit_r42_c61 bl[61] br[61] wl[42] vdd gnd cell_6t
Xbit_r43_c61 bl[61] br[61] wl[43] vdd gnd cell_6t
Xbit_r44_c61 bl[61] br[61] wl[44] vdd gnd cell_6t
Xbit_r45_c61 bl[61] br[61] wl[45] vdd gnd cell_6t
Xbit_r46_c61 bl[61] br[61] wl[46] vdd gnd cell_6t
Xbit_r47_c61 bl[61] br[61] wl[47] vdd gnd cell_6t
Xbit_r48_c61 bl[61] br[61] wl[48] vdd gnd cell_6t
Xbit_r49_c61 bl[61] br[61] wl[49] vdd gnd cell_6t
Xbit_r50_c61 bl[61] br[61] wl[50] vdd gnd cell_6t
Xbit_r51_c61 bl[61] br[61] wl[51] vdd gnd cell_6t
Xbit_r52_c61 bl[61] br[61] wl[52] vdd gnd cell_6t
Xbit_r53_c61 bl[61] br[61] wl[53] vdd gnd cell_6t
Xbit_r54_c61 bl[61] br[61] wl[54] vdd gnd cell_6t
Xbit_r55_c61 bl[61] br[61] wl[55] vdd gnd cell_6t
Xbit_r56_c61 bl[61] br[61] wl[56] vdd gnd cell_6t
Xbit_r57_c61 bl[61] br[61] wl[57] vdd gnd cell_6t
Xbit_r58_c61 bl[61] br[61] wl[58] vdd gnd cell_6t
Xbit_r59_c61 bl[61] br[61] wl[59] vdd gnd cell_6t
Xbit_r60_c61 bl[61] br[61] wl[60] vdd gnd cell_6t
Xbit_r61_c61 bl[61] br[61] wl[61] vdd gnd cell_6t
Xbit_r62_c61 bl[61] br[61] wl[62] vdd gnd cell_6t
Xbit_r63_c61 bl[61] br[61] wl[63] vdd gnd cell_6t
Xbit_r64_c61 bl[61] br[61] wl[64] vdd gnd cell_6t
Xbit_r65_c61 bl[61] br[61] wl[65] vdd gnd cell_6t
Xbit_r66_c61 bl[61] br[61] wl[66] vdd gnd cell_6t
Xbit_r67_c61 bl[61] br[61] wl[67] vdd gnd cell_6t
Xbit_r68_c61 bl[61] br[61] wl[68] vdd gnd cell_6t
Xbit_r69_c61 bl[61] br[61] wl[69] vdd gnd cell_6t
Xbit_r70_c61 bl[61] br[61] wl[70] vdd gnd cell_6t
Xbit_r71_c61 bl[61] br[61] wl[71] vdd gnd cell_6t
Xbit_r72_c61 bl[61] br[61] wl[72] vdd gnd cell_6t
Xbit_r73_c61 bl[61] br[61] wl[73] vdd gnd cell_6t
Xbit_r74_c61 bl[61] br[61] wl[74] vdd gnd cell_6t
Xbit_r75_c61 bl[61] br[61] wl[75] vdd gnd cell_6t
Xbit_r76_c61 bl[61] br[61] wl[76] vdd gnd cell_6t
Xbit_r77_c61 bl[61] br[61] wl[77] vdd gnd cell_6t
Xbit_r78_c61 bl[61] br[61] wl[78] vdd gnd cell_6t
Xbit_r79_c61 bl[61] br[61] wl[79] vdd gnd cell_6t
Xbit_r80_c61 bl[61] br[61] wl[80] vdd gnd cell_6t
Xbit_r81_c61 bl[61] br[61] wl[81] vdd gnd cell_6t
Xbit_r82_c61 bl[61] br[61] wl[82] vdd gnd cell_6t
Xbit_r83_c61 bl[61] br[61] wl[83] vdd gnd cell_6t
Xbit_r84_c61 bl[61] br[61] wl[84] vdd gnd cell_6t
Xbit_r85_c61 bl[61] br[61] wl[85] vdd gnd cell_6t
Xbit_r86_c61 bl[61] br[61] wl[86] vdd gnd cell_6t
Xbit_r87_c61 bl[61] br[61] wl[87] vdd gnd cell_6t
Xbit_r88_c61 bl[61] br[61] wl[88] vdd gnd cell_6t
Xbit_r89_c61 bl[61] br[61] wl[89] vdd gnd cell_6t
Xbit_r90_c61 bl[61] br[61] wl[90] vdd gnd cell_6t
Xbit_r91_c61 bl[61] br[61] wl[91] vdd gnd cell_6t
Xbit_r92_c61 bl[61] br[61] wl[92] vdd gnd cell_6t
Xbit_r93_c61 bl[61] br[61] wl[93] vdd gnd cell_6t
Xbit_r94_c61 bl[61] br[61] wl[94] vdd gnd cell_6t
Xbit_r95_c61 bl[61] br[61] wl[95] vdd gnd cell_6t
Xbit_r96_c61 bl[61] br[61] wl[96] vdd gnd cell_6t
Xbit_r97_c61 bl[61] br[61] wl[97] vdd gnd cell_6t
Xbit_r98_c61 bl[61] br[61] wl[98] vdd gnd cell_6t
Xbit_r99_c61 bl[61] br[61] wl[99] vdd gnd cell_6t
Xbit_r100_c61 bl[61] br[61] wl[100] vdd gnd cell_6t
Xbit_r101_c61 bl[61] br[61] wl[101] vdd gnd cell_6t
Xbit_r102_c61 bl[61] br[61] wl[102] vdd gnd cell_6t
Xbit_r103_c61 bl[61] br[61] wl[103] vdd gnd cell_6t
Xbit_r104_c61 bl[61] br[61] wl[104] vdd gnd cell_6t
Xbit_r105_c61 bl[61] br[61] wl[105] vdd gnd cell_6t
Xbit_r106_c61 bl[61] br[61] wl[106] vdd gnd cell_6t
Xbit_r107_c61 bl[61] br[61] wl[107] vdd gnd cell_6t
Xbit_r108_c61 bl[61] br[61] wl[108] vdd gnd cell_6t
Xbit_r109_c61 bl[61] br[61] wl[109] vdd gnd cell_6t
Xbit_r110_c61 bl[61] br[61] wl[110] vdd gnd cell_6t
Xbit_r111_c61 bl[61] br[61] wl[111] vdd gnd cell_6t
Xbit_r112_c61 bl[61] br[61] wl[112] vdd gnd cell_6t
Xbit_r113_c61 bl[61] br[61] wl[113] vdd gnd cell_6t
Xbit_r114_c61 bl[61] br[61] wl[114] vdd gnd cell_6t
Xbit_r115_c61 bl[61] br[61] wl[115] vdd gnd cell_6t
Xbit_r116_c61 bl[61] br[61] wl[116] vdd gnd cell_6t
Xbit_r117_c61 bl[61] br[61] wl[117] vdd gnd cell_6t
Xbit_r118_c61 bl[61] br[61] wl[118] vdd gnd cell_6t
Xbit_r119_c61 bl[61] br[61] wl[119] vdd gnd cell_6t
Xbit_r120_c61 bl[61] br[61] wl[120] vdd gnd cell_6t
Xbit_r121_c61 bl[61] br[61] wl[121] vdd gnd cell_6t
Xbit_r122_c61 bl[61] br[61] wl[122] vdd gnd cell_6t
Xbit_r123_c61 bl[61] br[61] wl[123] vdd gnd cell_6t
Xbit_r124_c61 bl[61] br[61] wl[124] vdd gnd cell_6t
Xbit_r125_c61 bl[61] br[61] wl[125] vdd gnd cell_6t
Xbit_r126_c61 bl[61] br[61] wl[126] vdd gnd cell_6t
Xbit_r127_c61 bl[61] br[61] wl[127] vdd gnd cell_6t
Xbit_r0_c62 bl[62] br[62] wl[0] vdd gnd cell_6t
Xbit_r1_c62 bl[62] br[62] wl[1] vdd gnd cell_6t
Xbit_r2_c62 bl[62] br[62] wl[2] vdd gnd cell_6t
Xbit_r3_c62 bl[62] br[62] wl[3] vdd gnd cell_6t
Xbit_r4_c62 bl[62] br[62] wl[4] vdd gnd cell_6t
Xbit_r5_c62 bl[62] br[62] wl[5] vdd gnd cell_6t
Xbit_r6_c62 bl[62] br[62] wl[6] vdd gnd cell_6t
Xbit_r7_c62 bl[62] br[62] wl[7] vdd gnd cell_6t
Xbit_r8_c62 bl[62] br[62] wl[8] vdd gnd cell_6t
Xbit_r9_c62 bl[62] br[62] wl[9] vdd gnd cell_6t
Xbit_r10_c62 bl[62] br[62] wl[10] vdd gnd cell_6t
Xbit_r11_c62 bl[62] br[62] wl[11] vdd gnd cell_6t
Xbit_r12_c62 bl[62] br[62] wl[12] vdd gnd cell_6t
Xbit_r13_c62 bl[62] br[62] wl[13] vdd gnd cell_6t
Xbit_r14_c62 bl[62] br[62] wl[14] vdd gnd cell_6t
Xbit_r15_c62 bl[62] br[62] wl[15] vdd gnd cell_6t
Xbit_r16_c62 bl[62] br[62] wl[16] vdd gnd cell_6t
Xbit_r17_c62 bl[62] br[62] wl[17] vdd gnd cell_6t
Xbit_r18_c62 bl[62] br[62] wl[18] vdd gnd cell_6t
Xbit_r19_c62 bl[62] br[62] wl[19] vdd gnd cell_6t
Xbit_r20_c62 bl[62] br[62] wl[20] vdd gnd cell_6t
Xbit_r21_c62 bl[62] br[62] wl[21] vdd gnd cell_6t
Xbit_r22_c62 bl[62] br[62] wl[22] vdd gnd cell_6t
Xbit_r23_c62 bl[62] br[62] wl[23] vdd gnd cell_6t
Xbit_r24_c62 bl[62] br[62] wl[24] vdd gnd cell_6t
Xbit_r25_c62 bl[62] br[62] wl[25] vdd gnd cell_6t
Xbit_r26_c62 bl[62] br[62] wl[26] vdd gnd cell_6t
Xbit_r27_c62 bl[62] br[62] wl[27] vdd gnd cell_6t
Xbit_r28_c62 bl[62] br[62] wl[28] vdd gnd cell_6t
Xbit_r29_c62 bl[62] br[62] wl[29] vdd gnd cell_6t
Xbit_r30_c62 bl[62] br[62] wl[30] vdd gnd cell_6t
Xbit_r31_c62 bl[62] br[62] wl[31] vdd gnd cell_6t
Xbit_r32_c62 bl[62] br[62] wl[32] vdd gnd cell_6t
Xbit_r33_c62 bl[62] br[62] wl[33] vdd gnd cell_6t
Xbit_r34_c62 bl[62] br[62] wl[34] vdd gnd cell_6t
Xbit_r35_c62 bl[62] br[62] wl[35] vdd gnd cell_6t
Xbit_r36_c62 bl[62] br[62] wl[36] vdd gnd cell_6t
Xbit_r37_c62 bl[62] br[62] wl[37] vdd gnd cell_6t
Xbit_r38_c62 bl[62] br[62] wl[38] vdd gnd cell_6t
Xbit_r39_c62 bl[62] br[62] wl[39] vdd gnd cell_6t
Xbit_r40_c62 bl[62] br[62] wl[40] vdd gnd cell_6t
Xbit_r41_c62 bl[62] br[62] wl[41] vdd gnd cell_6t
Xbit_r42_c62 bl[62] br[62] wl[42] vdd gnd cell_6t
Xbit_r43_c62 bl[62] br[62] wl[43] vdd gnd cell_6t
Xbit_r44_c62 bl[62] br[62] wl[44] vdd gnd cell_6t
Xbit_r45_c62 bl[62] br[62] wl[45] vdd gnd cell_6t
Xbit_r46_c62 bl[62] br[62] wl[46] vdd gnd cell_6t
Xbit_r47_c62 bl[62] br[62] wl[47] vdd gnd cell_6t
Xbit_r48_c62 bl[62] br[62] wl[48] vdd gnd cell_6t
Xbit_r49_c62 bl[62] br[62] wl[49] vdd gnd cell_6t
Xbit_r50_c62 bl[62] br[62] wl[50] vdd gnd cell_6t
Xbit_r51_c62 bl[62] br[62] wl[51] vdd gnd cell_6t
Xbit_r52_c62 bl[62] br[62] wl[52] vdd gnd cell_6t
Xbit_r53_c62 bl[62] br[62] wl[53] vdd gnd cell_6t
Xbit_r54_c62 bl[62] br[62] wl[54] vdd gnd cell_6t
Xbit_r55_c62 bl[62] br[62] wl[55] vdd gnd cell_6t
Xbit_r56_c62 bl[62] br[62] wl[56] vdd gnd cell_6t
Xbit_r57_c62 bl[62] br[62] wl[57] vdd gnd cell_6t
Xbit_r58_c62 bl[62] br[62] wl[58] vdd gnd cell_6t
Xbit_r59_c62 bl[62] br[62] wl[59] vdd gnd cell_6t
Xbit_r60_c62 bl[62] br[62] wl[60] vdd gnd cell_6t
Xbit_r61_c62 bl[62] br[62] wl[61] vdd gnd cell_6t
Xbit_r62_c62 bl[62] br[62] wl[62] vdd gnd cell_6t
Xbit_r63_c62 bl[62] br[62] wl[63] vdd gnd cell_6t
Xbit_r64_c62 bl[62] br[62] wl[64] vdd gnd cell_6t
Xbit_r65_c62 bl[62] br[62] wl[65] vdd gnd cell_6t
Xbit_r66_c62 bl[62] br[62] wl[66] vdd gnd cell_6t
Xbit_r67_c62 bl[62] br[62] wl[67] vdd gnd cell_6t
Xbit_r68_c62 bl[62] br[62] wl[68] vdd gnd cell_6t
Xbit_r69_c62 bl[62] br[62] wl[69] vdd gnd cell_6t
Xbit_r70_c62 bl[62] br[62] wl[70] vdd gnd cell_6t
Xbit_r71_c62 bl[62] br[62] wl[71] vdd gnd cell_6t
Xbit_r72_c62 bl[62] br[62] wl[72] vdd gnd cell_6t
Xbit_r73_c62 bl[62] br[62] wl[73] vdd gnd cell_6t
Xbit_r74_c62 bl[62] br[62] wl[74] vdd gnd cell_6t
Xbit_r75_c62 bl[62] br[62] wl[75] vdd gnd cell_6t
Xbit_r76_c62 bl[62] br[62] wl[76] vdd gnd cell_6t
Xbit_r77_c62 bl[62] br[62] wl[77] vdd gnd cell_6t
Xbit_r78_c62 bl[62] br[62] wl[78] vdd gnd cell_6t
Xbit_r79_c62 bl[62] br[62] wl[79] vdd gnd cell_6t
Xbit_r80_c62 bl[62] br[62] wl[80] vdd gnd cell_6t
Xbit_r81_c62 bl[62] br[62] wl[81] vdd gnd cell_6t
Xbit_r82_c62 bl[62] br[62] wl[82] vdd gnd cell_6t
Xbit_r83_c62 bl[62] br[62] wl[83] vdd gnd cell_6t
Xbit_r84_c62 bl[62] br[62] wl[84] vdd gnd cell_6t
Xbit_r85_c62 bl[62] br[62] wl[85] vdd gnd cell_6t
Xbit_r86_c62 bl[62] br[62] wl[86] vdd gnd cell_6t
Xbit_r87_c62 bl[62] br[62] wl[87] vdd gnd cell_6t
Xbit_r88_c62 bl[62] br[62] wl[88] vdd gnd cell_6t
Xbit_r89_c62 bl[62] br[62] wl[89] vdd gnd cell_6t
Xbit_r90_c62 bl[62] br[62] wl[90] vdd gnd cell_6t
Xbit_r91_c62 bl[62] br[62] wl[91] vdd gnd cell_6t
Xbit_r92_c62 bl[62] br[62] wl[92] vdd gnd cell_6t
Xbit_r93_c62 bl[62] br[62] wl[93] vdd gnd cell_6t
Xbit_r94_c62 bl[62] br[62] wl[94] vdd gnd cell_6t
Xbit_r95_c62 bl[62] br[62] wl[95] vdd gnd cell_6t
Xbit_r96_c62 bl[62] br[62] wl[96] vdd gnd cell_6t
Xbit_r97_c62 bl[62] br[62] wl[97] vdd gnd cell_6t
Xbit_r98_c62 bl[62] br[62] wl[98] vdd gnd cell_6t
Xbit_r99_c62 bl[62] br[62] wl[99] vdd gnd cell_6t
Xbit_r100_c62 bl[62] br[62] wl[100] vdd gnd cell_6t
Xbit_r101_c62 bl[62] br[62] wl[101] vdd gnd cell_6t
Xbit_r102_c62 bl[62] br[62] wl[102] vdd gnd cell_6t
Xbit_r103_c62 bl[62] br[62] wl[103] vdd gnd cell_6t
Xbit_r104_c62 bl[62] br[62] wl[104] vdd gnd cell_6t
Xbit_r105_c62 bl[62] br[62] wl[105] vdd gnd cell_6t
Xbit_r106_c62 bl[62] br[62] wl[106] vdd gnd cell_6t
Xbit_r107_c62 bl[62] br[62] wl[107] vdd gnd cell_6t
Xbit_r108_c62 bl[62] br[62] wl[108] vdd gnd cell_6t
Xbit_r109_c62 bl[62] br[62] wl[109] vdd gnd cell_6t
Xbit_r110_c62 bl[62] br[62] wl[110] vdd gnd cell_6t
Xbit_r111_c62 bl[62] br[62] wl[111] vdd gnd cell_6t
Xbit_r112_c62 bl[62] br[62] wl[112] vdd gnd cell_6t
Xbit_r113_c62 bl[62] br[62] wl[113] vdd gnd cell_6t
Xbit_r114_c62 bl[62] br[62] wl[114] vdd gnd cell_6t
Xbit_r115_c62 bl[62] br[62] wl[115] vdd gnd cell_6t
Xbit_r116_c62 bl[62] br[62] wl[116] vdd gnd cell_6t
Xbit_r117_c62 bl[62] br[62] wl[117] vdd gnd cell_6t
Xbit_r118_c62 bl[62] br[62] wl[118] vdd gnd cell_6t
Xbit_r119_c62 bl[62] br[62] wl[119] vdd gnd cell_6t
Xbit_r120_c62 bl[62] br[62] wl[120] vdd gnd cell_6t
Xbit_r121_c62 bl[62] br[62] wl[121] vdd gnd cell_6t
Xbit_r122_c62 bl[62] br[62] wl[122] vdd gnd cell_6t
Xbit_r123_c62 bl[62] br[62] wl[123] vdd gnd cell_6t
Xbit_r124_c62 bl[62] br[62] wl[124] vdd gnd cell_6t
Xbit_r125_c62 bl[62] br[62] wl[125] vdd gnd cell_6t
Xbit_r126_c62 bl[62] br[62] wl[126] vdd gnd cell_6t
Xbit_r127_c62 bl[62] br[62] wl[127] vdd gnd cell_6t
Xbit_r0_c63 bl[63] br[63] wl[0] vdd gnd cell_6t
Xbit_r1_c63 bl[63] br[63] wl[1] vdd gnd cell_6t
Xbit_r2_c63 bl[63] br[63] wl[2] vdd gnd cell_6t
Xbit_r3_c63 bl[63] br[63] wl[3] vdd gnd cell_6t
Xbit_r4_c63 bl[63] br[63] wl[4] vdd gnd cell_6t
Xbit_r5_c63 bl[63] br[63] wl[5] vdd gnd cell_6t
Xbit_r6_c63 bl[63] br[63] wl[6] vdd gnd cell_6t
Xbit_r7_c63 bl[63] br[63] wl[7] vdd gnd cell_6t
Xbit_r8_c63 bl[63] br[63] wl[8] vdd gnd cell_6t
Xbit_r9_c63 bl[63] br[63] wl[9] vdd gnd cell_6t
Xbit_r10_c63 bl[63] br[63] wl[10] vdd gnd cell_6t
Xbit_r11_c63 bl[63] br[63] wl[11] vdd gnd cell_6t
Xbit_r12_c63 bl[63] br[63] wl[12] vdd gnd cell_6t
Xbit_r13_c63 bl[63] br[63] wl[13] vdd gnd cell_6t
Xbit_r14_c63 bl[63] br[63] wl[14] vdd gnd cell_6t
Xbit_r15_c63 bl[63] br[63] wl[15] vdd gnd cell_6t
Xbit_r16_c63 bl[63] br[63] wl[16] vdd gnd cell_6t
Xbit_r17_c63 bl[63] br[63] wl[17] vdd gnd cell_6t
Xbit_r18_c63 bl[63] br[63] wl[18] vdd gnd cell_6t
Xbit_r19_c63 bl[63] br[63] wl[19] vdd gnd cell_6t
Xbit_r20_c63 bl[63] br[63] wl[20] vdd gnd cell_6t
Xbit_r21_c63 bl[63] br[63] wl[21] vdd gnd cell_6t
Xbit_r22_c63 bl[63] br[63] wl[22] vdd gnd cell_6t
Xbit_r23_c63 bl[63] br[63] wl[23] vdd gnd cell_6t
Xbit_r24_c63 bl[63] br[63] wl[24] vdd gnd cell_6t
Xbit_r25_c63 bl[63] br[63] wl[25] vdd gnd cell_6t
Xbit_r26_c63 bl[63] br[63] wl[26] vdd gnd cell_6t
Xbit_r27_c63 bl[63] br[63] wl[27] vdd gnd cell_6t
Xbit_r28_c63 bl[63] br[63] wl[28] vdd gnd cell_6t
Xbit_r29_c63 bl[63] br[63] wl[29] vdd gnd cell_6t
Xbit_r30_c63 bl[63] br[63] wl[30] vdd gnd cell_6t
Xbit_r31_c63 bl[63] br[63] wl[31] vdd gnd cell_6t
Xbit_r32_c63 bl[63] br[63] wl[32] vdd gnd cell_6t
Xbit_r33_c63 bl[63] br[63] wl[33] vdd gnd cell_6t
Xbit_r34_c63 bl[63] br[63] wl[34] vdd gnd cell_6t
Xbit_r35_c63 bl[63] br[63] wl[35] vdd gnd cell_6t
Xbit_r36_c63 bl[63] br[63] wl[36] vdd gnd cell_6t
Xbit_r37_c63 bl[63] br[63] wl[37] vdd gnd cell_6t
Xbit_r38_c63 bl[63] br[63] wl[38] vdd gnd cell_6t
Xbit_r39_c63 bl[63] br[63] wl[39] vdd gnd cell_6t
Xbit_r40_c63 bl[63] br[63] wl[40] vdd gnd cell_6t
Xbit_r41_c63 bl[63] br[63] wl[41] vdd gnd cell_6t
Xbit_r42_c63 bl[63] br[63] wl[42] vdd gnd cell_6t
Xbit_r43_c63 bl[63] br[63] wl[43] vdd gnd cell_6t
Xbit_r44_c63 bl[63] br[63] wl[44] vdd gnd cell_6t
Xbit_r45_c63 bl[63] br[63] wl[45] vdd gnd cell_6t
Xbit_r46_c63 bl[63] br[63] wl[46] vdd gnd cell_6t
Xbit_r47_c63 bl[63] br[63] wl[47] vdd gnd cell_6t
Xbit_r48_c63 bl[63] br[63] wl[48] vdd gnd cell_6t
Xbit_r49_c63 bl[63] br[63] wl[49] vdd gnd cell_6t
Xbit_r50_c63 bl[63] br[63] wl[50] vdd gnd cell_6t
Xbit_r51_c63 bl[63] br[63] wl[51] vdd gnd cell_6t
Xbit_r52_c63 bl[63] br[63] wl[52] vdd gnd cell_6t
Xbit_r53_c63 bl[63] br[63] wl[53] vdd gnd cell_6t
Xbit_r54_c63 bl[63] br[63] wl[54] vdd gnd cell_6t
Xbit_r55_c63 bl[63] br[63] wl[55] vdd gnd cell_6t
Xbit_r56_c63 bl[63] br[63] wl[56] vdd gnd cell_6t
Xbit_r57_c63 bl[63] br[63] wl[57] vdd gnd cell_6t
Xbit_r58_c63 bl[63] br[63] wl[58] vdd gnd cell_6t
Xbit_r59_c63 bl[63] br[63] wl[59] vdd gnd cell_6t
Xbit_r60_c63 bl[63] br[63] wl[60] vdd gnd cell_6t
Xbit_r61_c63 bl[63] br[63] wl[61] vdd gnd cell_6t
Xbit_r62_c63 bl[63] br[63] wl[62] vdd gnd cell_6t
Xbit_r63_c63 bl[63] br[63] wl[63] vdd gnd cell_6t
Xbit_r64_c63 bl[63] br[63] wl[64] vdd gnd cell_6t
Xbit_r65_c63 bl[63] br[63] wl[65] vdd gnd cell_6t
Xbit_r66_c63 bl[63] br[63] wl[66] vdd gnd cell_6t
Xbit_r67_c63 bl[63] br[63] wl[67] vdd gnd cell_6t
Xbit_r68_c63 bl[63] br[63] wl[68] vdd gnd cell_6t
Xbit_r69_c63 bl[63] br[63] wl[69] vdd gnd cell_6t
Xbit_r70_c63 bl[63] br[63] wl[70] vdd gnd cell_6t
Xbit_r71_c63 bl[63] br[63] wl[71] vdd gnd cell_6t
Xbit_r72_c63 bl[63] br[63] wl[72] vdd gnd cell_6t
Xbit_r73_c63 bl[63] br[63] wl[73] vdd gnd cell_6t
Xbit_r74_c63 bl[63] br[63] wl[74] vdd gnd cell_6t
Xbit_r75_c63 bl[63] br[63] wl[75] vdd gnd cell_6t
Xbit_r76_c63 bl[63] br[63] wl[76] vdd gnd cell_6t
Xbit_r77_c63 bl[63] br[63] wl[77] vdd gnd cell_6t
Xbit_r78_c63 bl[63] br[63] wl[78] vdd gnd cell_6t
Xbit_r79_c63 bl[63] br[63] wl[79] vdd gnd cell_6t
Xbit_r80_c63 bl[63] br[63] wl[80] vdd gnd cell_6t
Xbit_r81_c63 bl[63] br[63] wl[81] vdd gnd cell_6t
Xbit_r82_c63 bl[63] br[63] wl[82] vdd gnd cell_6t
Xbit_r83_c63 bl[63] br[63] wl[83] vdd gnd cell_6t
Xbit_r84_c63 bl[63] br[63] wl[84] vdd gnd cell_6t
Xbit_r85_c63 bl[63] br[63] wl[85] vdd gnd cell_6t
Xbit_r86_c63 bl[63] br[63] wl[86] vdd gnd cell_6t
Xbit_r87_c63 bl[63] br[63] wl[87] vdd gnd cell_6t
Xbit_r88_c63 bl[63] br[63] wl[88] vdd gnd cell_6t
Xbit_r89_c63 bl[63] br[63] wl[89] vdd gnd cell_6t
Xbit_r90_c63 bl[63] br[63] wl[90] vdd gnd cell_6t
Xbit_r91_c63 bl[63] br[63] wl[91] vdd gnd cell_6t
Xbit_r92_c63 bl[63] br[63] wl[92] vdd gnd cell_6t
Xbit_r93_c63 bl[63] br[63] wl[93] vdd gnd cell_6t
Xbit_r94_c63 bl[63] br[63] wl[94] vdd gnd cell_6t
Xbit_r95_c63 bl[63] br[63] wl[95] vdd gnd cell_6t
Xbit_r96_c63 bl[63] br[63] wl[96] vdd gnd cell_6t
Xbit_r97_c63 bl[63] br[63] wl[97] vdd gnd cell_6t
Xbit_r98_c63 bl[63] br[63] wl[98] vdd gnd cell_6t
Xbit_r99_c63 bl[63] br[63] wl[99] vdd gnd cell_6t
Xbit_r100_c63 bl[63] br[63] wl[100] vdd gnd cell_6t
Xbit_r101_c63 bl[63] br[63] wl[101] vdd gnd cell_6t
Xbit_r102_c63 bl[63] br[63] wl[102] vdd gnd cell_6t
Xbit_r103_c63 bl[63] br[63] wl[103] vdd gnd cell_6t
Xbit_r104_c63 bl[63] br[63] wl[104] vdd gnd cell_6t
Xbit_r105_c63 bl[63] br[63] wl[105] vdd gnd cell_6t
Xbit_r106_c63 bl[63] br[63] wl[106] vdd gnd cell_6t
Xbit_r107_c63 bl[63] br[63] wl[107] vdd gnd cell_6t
Xbit_r108_c63 bl[63] br[63] wl[108] vdd gnd cell_6t
Xbit_r109_c63 bl[63] br[63] wl[109] vdd gnd cell_6t
Xbit_r110_c63 bl[63] br[63] wl[110] vdd gnd cell_6t
Xbit_r111_c63 bl[63] br[63] wl[111] vdd gnd cell_6t
Xbit_r112_c63 bl[63] br[63] wl[112] vdd gnd cell_6t
Xbit_r113_c63 bl[63] br[63] wl[113] vdd gnd cell_6t
Xbit_r114_c63 bl[63] br[63] wl[114] vdd gnd cell_6t
Xbit_r115_c63 bl[63] br[63] wl[115] vdd gnd cell_6t
Xbit_r116_c63 bl[63] br[63] wl[116] vdd gnd cell_6t
Xbit_r117_c63 bl[63] br[63] wl[117] vdd gnd cell_6t
Xbit_r118_c63 bl[63] br[63] wl[118] vdd gnd cell_6t
Xbit_r119_c63 bl[63] br[63] wl[119] vdd gnd cell_6t
Xbit_r120_c63 bl[63] br[63] wl[120] vdd gnd cell_6t
Xbit_r121_c63 bl[63] br[63] wl[121] vdd gnd cell_6t
Xbit_r122_c63 bl[63] br[63] wl[122] vdd gnd cell_6t
Xbit_r123_c63 bl[63] br[63] wl[123] vdd gnd cell_6t
Xbit_r124_c63 bl[63] br[63] wl[124] vdd gnd cell_6t
Xbit_r125_c63 bl[63] br[63] wl[125] vdd gnd cell_6t
Xbit_r126_c63 bl[63] br[63] wl[126] vdd gnd cell_6t
Xbit_r127_c63 bl[63] br[63] wl[127] vdd gnd cell_6t
Xbit_r0_c64 bl[64] br[64] wl[0] vdd gnd cell_6t
Xbit_r1_c64 bl[64] br[64] wl[1] vdd gnd cell_6t
Xbit_r2_c64 bl[64] br[64] wl[2] vdd gnd cell_6t
Xbit_r3_c64 bl[64] br[64] wl[3] vdd gnd cell_6t
Xbit_r4_c64 bl[64] br[64] wl[4] vdd gnd cell_6t
Xbit_r5_c64 bl[64] br[64] wl[5] vdd gnd cell_6t
Xbit_r6_c64 bl[64] br[64] wl[6] vdd gnd cell_6t
Xbit_r7_c64 bl[64] br[64] wl[7] vdd gnd cell_6t
Xbit_r8_c64 bl[64] br[64] wl[8] vdd gnd cell_6t
Xbit_r9_c64 bl[64] br[64] wl[9] vdd gnd cell_6t
Xbit_r10_c64 bl[64] br[64] wl[10] vdd gnd cell_6t
Xbit_r11_c64 bl[64] br[64] wl[11] vdd gnd cell_6t
Xbit_r12_c64 bl[64] br[64] wl[12] vdd gnd cell_6t
Xbit_r13_c64 bl[64] br[64] wl[13] vdd gnd cell_6t
Xbit_r14_c64 bl[64] br[64] wl[14] vdd gnd cell_6t
Xbit_r15_c64 bl[64] br[64] wl[15] vdd gnd cell_6t
Xbit_r16_c64 bl[64] br[64] wl[16] vdd gnd cell_6t
Xbit_r17_c64 bl[64] br[64] wl[17] vdd gnd cell_6t
Xbit_r18_c64 bl[64] br[64] wl[18] vdd gnd cell_6t
Xbit_r19_c64 bl[64] br[64] wl[19] vdd gnd cell_6t
Xbit_r20_c64 bl[64] br[64] wl[20] vdd gnd cell_6t
Xbit_r21_c64 bl[64] br[64] wl[21] vdd gnd cell_6t
Xbit_r22_c64 bl[64] br[64] wl[22] vdd gnd cell_6t
Xbit_r23_c64 bl[64] br[64] wl[23] vdd gnd cell_6t
Xbit_r24_c64 bl[64] br[64] wl[24] vdd gnd cell_6t
Xbit_r25_c64 bl[64] br[64] wl[25] vdd gnd cell_6t
Xbit_r26_c64 bl[64] br[64] wl[26] vdd gnd cell_6t
Xbit_r27_c64 bl[64] br[64] wl[27] vdd gnd cell_6t
Xbit_r28_c64 bl[64] br[64] wl[28] vdd gnd cell_6t
Xbit_r29_c64 bl[64] br[64] wl[29] vdd gnd cell_6t
Xbit_r30_c64 bl[64] br[64] wl[30] vdd gnd cell_6t
Xbit_r31_c64 bl[64] br[64] wl[31] vdd gnd cell_6t
Xbit_r32_c64 bl[64] br[64] wl[32] vdd gnd cell_6t
Xbit_r33_c64 bl[64] br[64] wl[33] vdd gnd cell_6t
Xbit_r34_c64 bl[64] br[64] wl[34] vdd gnd cell_6t
Xbit_r35_c64 bl[64] br[64] wl[35] vdd gnd cell_6t
Xbit_r36_c64 bl[64] br[64] wl[36] vdd gnd cell_6t
Xbit_r37_c64 bl[64] br[64] wl[37] vdd gnd cell_6t
Xbit_r38_c64 bl[64] br[64] wl[38] vdd gnd cell_6t
Xbit_r39_c64 bl[64] br[64] wl[39] vdd gnd cell_6t
Xbit_r40_c64 bl[64] br[64] wl[40] vdd gnd cell_6t
Xbit_r41_c64 bl[64] br[64] wl[41] vdd gnd cell_6t
Xbit_r42_c64 bl[64] br[64] wl[42] vdd gnd cell_6t
Xbit_r43_c64 bl[64] br[64] wl[43] vdd gnd cell_6t
Xbit_r44_c64 bl[64] br[64] wl[44] vdd gnd cell_6t
Xbit_r45_c64 bl[64] br[64] wl[45] vdd gnd cell_6t
Xbit_r46_c64 bl[64] br[64] wl[46] vdd gnd cell_6t
Xbit_r47_c64 bl[64] br[64] wl[47] vdd gnd cell_6t
Xbit_r48_c64 bl[64] br[64] wl[48] vdd gnd cell_6t
Xbit_r49_c64 bl[64] br[64] wl[49] vdd gnd cell_6t
Xbit_r50_c64 bl[64] br[64] wl[50] vdd gnd cell_6t
Xbit_r51_c64 bl[64] br[64] wl[51] vdd gnd cell_6t
Xbit_r52_c64 bl[64] br[64] wl[52] vdd gnd cell_6t
Xbit_r53_c64 bl[64] br[64] wl[53] vdd gnd cell_6t
Xbit_r54_c64 bl[64] br[64] wl[54] vdd gnd cell_6t
Xbit_r55_c64 bl[64] br[64] wl[55] vdd gnd cell_6t
Xbit_r56_c64 bl[64] br[64] wl[56] vdd gnd cell_6t
Xbit_r57_c64 bl[64] br[64] wl[57] vdd gnd cell_6t
Xbit_r58_c64 bl[64] br[64] wl[58] vdd gnd cell_6t
Xbit_r59_c64 bl[64] br[64] wl[59] vdd gnd cell_6t
Xbit_r60_c64 bl[64] br[64] wl[60] vdd gnd cell_6t
Xbit_r61_c64 bl[64] br[64] wl[61] vdd gnd cell_6t
Xbit_r62_c64 bl[64] br[64] wl[62] vdd gnd cell_6t
Xbit_r63_c64 bl[64] br[64] wl[63] vdd gnd cell_6t
Xbit_r64_c64 bl[64] br[64] wl[64] vdd gnd cell_6t
Xbit_r65_c64 bl[64] br[64] wl[65] vdd gnd cell_6t
Xbit_r66_c64 bl[64] br[64] wl[66] vdd gnd cell_6t
Xbit_r67_c64 bl[64] br[64] wl[67] vdd gnd cell_6t
Xbit_r68_c64 bl[64] br[64] wl[68] vdd gnd cell_6t
Xbit_r69_c64 bl[64] br[64] wl[69] vdd gnd cell_6t
Xbit_r70_c64 bl[64] br[64] wl[70] vdd gnd cell_6t
Xbit_r71_c64 bl[64] br[64] wl[71] vdd gnd cell_6t
Xbit_r72_c64 bl[64] br[64] wl[72] vdd gnd cell_6t
Xbit_r73_c64 bl[64] br[64] wl[73] vdd gnd cell_6t
Xbit_r74_c64 bl[64] br[64] wl[74] vdd gnd cell_6t
Xbit_r75_c64 bl[64] br[64] wl[75] vdd gnd cell_6t
Xbit_r76_c64 bl[64] br[64] wl[76] vdd gnd cell_6t
Xbit_r77_c64 bl[64] br[64] wl[77] vdd gnd cell_6t
Xbit_r78_c64 bl[64] br[64] wl[78] vdd gnd cell_6t
Xbit_r79_c64 bl[64] br[64] wl[79] vdd gnd cell_6t
Xbit_r80_c64 bl[64] br[64] wl[80] vdd gnd cell_6t
Xbit_r81_c64 bl[64] br[64] wl[81] vdd gnd cell_6t
Xbit_r82_c64 bl[64] br[64] wl[82] vdd gnd cell_6t
Xbit_r83_c64 bl[64] br[64] wl[83] vdd gnd cell_6t
Xbit_r84_c64 bl[64] br[64] wl[84] vdd gnd cell_6t
Xbit_r85_c64 bl[64] br[64] wl[85] vdd gnd cell_6t
Xbit_r86_c64 bl[64] br[64] wl[86] vdd gnd cell_6t
Xbit_r87_c64 bl[64] br[64] wl[87] vdd gnd cell_6t
Xbit_r88_c64 bl[64] br[64] wl[88] vdd gnd cell_6t
Xbit_r89_c64 bl[64] br[64] wl[89] vdd gnd cell_6t
Xbit_r90_c64 bl[64] br[64] wl[90] vdd gnd cell_6t
Xbit_r91_c64 bl[64] br[64] wl[91] vdd gnd cell_6t
Xbit_r92_c64 bl[64] br[64] wl[92] vdd gnd cell_6t
Xbit_r93_c64 bl[64] br[64] wl[93] vdd gnd cell_6t
Xbit_r94_c64 bl[64] br[64] wl[94] vdd gnd cell_6t
Xbit_r95_c64 bl[64] br[64] wl[95] vdd gnd cell_6t
Xbit_r96_c64 bl[64] br[64] wl[96] vdd gnd cell_6t
Xbit_r97_c64 bl[64] br[64] wl[97] vdd gnd cell_6t
Xbit_r98_c64 bl[64] br[64] wl[98] vdd gnd cell_6t
Xbit_r99_c64 bl[64] br[64] wl[99] vdd gnd cell_6t
Xbit_r100_c64 bl[64] br[64] wl[100] vdd gnd cell_6t
Xbit_r101_c64 bl[64] br[64] wl[101] vdd gnd cell_6t
Xbit_r102_c64 bl[64] br[64] wl[102] vdd gnd cell_6t
Xbit_r103_c64 bl[64] br[64] wl[103] vdd gnd cell_6t
Xbit_r104_c64 bl[64] br[64] wl[104] vdd gnd cell_6t
Xbit_r105_c64 bl[64] br[64] wl[105] vdd gnd cell_6t
Xbit_r106_c64 bl[64] br[64] wl[106] vdd gnd cell_6t
Xbit_r107_c64 bl[64] br[64] wl[107] vdd gnd cell_6t
Xbit_r108_c64 bl[64] br[64] wl[108] vdd gnd cell_6t
Xbit_r109_c64 bl[64] br[64] wl[109] vdd gnd cell_6t
Xbit_r110_c64 bl[64] br[64] wl[110] vdd gnd cell_6t
Xbit_r111_c64 bl[64] br[64] wl[111] vdd gnd cell_6t
Xbit_r112_c64 bl[64] br[64] wl[112] vdd gnd cell_6t
Xbit_r113_c64 bl[64] br[64] wl[113] vdd gnd cell_6t
Xbit_r114_c64 bl[64] br[64] wl[114] vdd gnd cell_6t
Xbit_r115_c64 bl[64] br[64] wl[115] vdd gnd cell_6t
Xbit_r116_c64 bl[64] br[64] wl[116] vdd gnd cell_6t
Xbit_r117_c64 bl[64] br[64] wl[117] vdd gnd cell_6t
Xbit_r118_c64 bl[64] br[64] wl[118] vdd gnd cell_6t
Xbit_r119_c64 bl[64] br[64] wl[119] vdd gnd cell_6t
Xbit_r120_c64 bl[64] br[64] wl[120] vdd gnd cell_6t
Xbit_r121_c64 bl[64] br[64] wl[121] vdd gnd cell_6t
Xbit_r122_c64 bl[64] br[64] wl[122] vdd gnd cell_6t
Xbit_r123_c64 bl[64] br[64] wl[123] vdd gnd cell_6t
Xbit_r124_c64 bl[64] br[64] wl[124] vdd gnd cell_6t
Xbit_r125_c64 bl[64] br[64] wl[125] vdd gnd cell_6t
Xbit_r126_c64 bl[64] br[64] wl[126] vdd gnd cell_6t
Xbit_r127_c64 bl[64] br[64] wl[127] vdd gnd cell_6t
Xbit_r0_c65 bl[65] br[65] wl[0] vdd gnd cell_6t
Xbit_r1_c65 bl[65] br[65] wl[1] vdd gnd cell_6t
Xbit_r2_c65 bl[65] br[65] wl[2] vdd gnd cell_6t
Xbit_r3_c65 bl[65] br[65] wl[3] vdd gnd cell_6t
Xbit_r4_c65 bl[65] br[65] wl[4] vdd gnd cell_6t
Xbit_r5_c65 bl[65] br[65] wl[5] vdd gnd cell_6t
Xbit_r6_c65 bl[65] br[65] wl[6] vdd gnd cell_6t
Xbit_r7_c65 bl[65] br[65] wl[7] vdd gnd cell_6t
Xbit_r8_c65 bl[65] br[65] wl[8] vdd gnd cell_6t
Xbit_r9_c65 bl[65] br[65] wl[9] vdd gnd cell_6t
Xbit_r10_c65 bl[65] br[65] wl[10] vdd gnd cell_6t
Xbit_r11_c65 bl[65] br[65] wl[11] vdd gnd cell_6t
Xbit_r12_c65 bl[65] br[65] wl[12] vdd gnd cell_6t
Xbit_r13_c65 bl[65] br[65] wl[13] vdd gnd cell_6t
Xbit_r14_c65 bl[65] br[65] wl[14] vdd gnd cell_6t
Xbit_r15_c65 bl[65] br[65] wl[15] vdd gnd cell_6t
Xbit_r16_c65 bl[65] br[65] wl[16] vdd gnd cell_6t
Xbit_r17_c65 bl[65] br[65] wl[17] vdd gnd cell_6t
Xbit_r18_c65 bl[65] br[65] wl[18] vdd gnd cell_6t
Xbit_r19_c65 bl[65] br[65] wl[19] vdd gnd cell_6t
Xbit_r20_c65 bl[65] br[65] wl[20] vdd gnd cell_6t
Xbit_r21_c65 bl[65] br[65] wl[21] vdd gnd cell_6t
Xbit_r22_c65 bl[65] br[65] wl[22] vdd gnd cell_6t
Xbit_r23_c65 bl[65] br[65] wl[23] vdd gnd cell_6t
Xbit_r24_c65 bl[65] br[65] wl[24] vdd gnd cell_6t
Xbit_r25_c65 bl[65] br[65] wl[25] vdd gnd cell_6t
Xbit_r26_c65 bl[65] br[65] wl[26] vdd gnd cell_6t
Xbit_r27_c65 bl[65] br[65] wl[27] vdd gnd cell_6t
Xbit_r28_c65 bl[65] br[65] wl[28] vdd gnd cell_6t
Xbit_r29_c65 bl[65] br[65] wl[29] vdd gnd cell_6t
Xbit_r30_c65 bl[65] br[65] wl[30] vdd gnd cell_6t
Xbit_r31_c65 bl[65] br[65] wl[31] vdd gnd cell_6t
Xbit_r32_c65 bl[65] br[65] wl[32] vdd gnd cell_6t
Xbit_r33_c65 bl[65] br[65] wl[33] vdd gnd cell_6t
Xbit_r34_c65 bl[65] br[65] wl[34] vdd gnd cell_6t
Xbit_r35_c65 bl[65] br[65] wl[35] vdd gnd cell_6t
Xbit_r36_c65 bl[65] br[65] wl[36] vdd gnd cell_6t
Xbit_r37_c65 bl[65] br[65] wl[37] vdd gnd cell_6t
Xbit_r38_c65 bl[65] br[65] wl[38] vdd gnd cell_6t
Xbit_r39_c65 bl[65] br[65] wl[39] vdd gnd cell_6t
Xbit_r40_c65 bl[65] br[65] wl[40] vdd gnd cell_6t
Xbit_r41_c65 bl[65] br[65] wl[41] vdd gnd cell_6t
Xbit_r42_c65 bl[65] br[65] wl[42] vdd gnd cell_6t
Xbit_r43_c65 bl[65] br[65] wl[43] vdd gnd cell_6t
Xbit_r44_c65 bl[65] br[65] wl[44] vdd gnd cell_6t
Xbit_r45_c65 bl[65] br[65] wl[45] vdd gnd cell_6t
Xbit_r46_c65 bl[65] br[65] wl[46] vdd gnd cell_6t
Xbit_r47_c65 bl[65] br[65] wl[47] vdd gnd cell_6t
Xbit_r48_c65 bl[65] br[65] wl[48] vdd gnd cell_6t
Xbit_r49_c65 bl[65] br[65] wl[49] vdd gnd cell_6t
Xbit_r50_c65 bl[65] br[65] wl[50] vdd gnd cell_6t
Xbit_r51_c65 bl[65] br[65] wl[51] vdd gnd cell_6t
Xbit_r52_c65 bl[65] br[65] wl[52] vdd gnd cell_6t
Xbit_r53_c65 bl[65] br[65] wl[53] vdd gnd cell_6t
Xbit_r54_c65 bl[65] br[65] wl[54] vdd gnd cell_6t
Xbit_r55_c65 bl[65] br[65] wl[55] vdd gnd cell_6t
Xbit_r56_c65 bl[65] br[65] wl[56] vdd gnd cell_6t
Xbit_r57_c65 bl[65] br[65] wl[57] vdd gnd cell_6t
Xbit_r58_c65 bl[65] br[65] wl[58] vdd gnd cell_6t
Xbit_r59_c65 bl[65] br[65] wl[59] vdd gnd cell_6t
Xbit_r60_c65 bl[65] br[65] wl[60] vdd gnd cell_6t
Xbit_r61_c65 bl[65] br[65] wl[61] vdd gnd cell_6t
Xbit_r62_c65 bl[65] br[65] wl[62] vdd gnd cell_6t
Xbit_r63_c65 bl[65] br[65] wl[63] vdd gnd cell_6t
Xbit_r64_c65 bl[65] br[65] wl[64] vdd gnd cell_6t
Xbit_r65_c65 bl[65] br[65] wl[65] vdd gnd cell_6t
Xbit_r66_c65 bl[65] br[65] wl[66] vdd gnd cell_6t
Xbit_r67_c65 bl[65] br[65] wl[67] vdd gnd cell_6t
Xbit_r68_c65 bl[65] br[65] wl[68] vdd gnd cell_6t
Xbit_r69_c65 bl[65] br[65] wl[69] vdd gnd cell_6t
Xbit_r70_c65 bl[65] br[65] wl[70] vdd gnd cell_6t
Xbit_r71_c65 bl[65] br[65] wl[71] vdd gnd cell_6t
Xbit_r72_c65 bl[65] br[65] wl[72] vdd gnd cell_6t
Xbit_r73_c65 bl[65] br[65] wl[73] vdd gnd cell_6t
Xbit_r74_c65 bl[65] br[65] wl[74] vdd gnd cell_6t
Xbit_r75_c65 bl[65] br[65] wl[75] vdd gnd cell_6t
Xbit_r76_c65 bl[65] br[65] wl[76] vdd gnd cell_6t
Xbit_r77_c65 bl[65] br[65] wl[77] vdd gnd cell_6t
Xbit_r78_c65 bl[65] br[65] wl[78] vdd gnd cell_6t
Xbit_r79_c65 bl[65] br[65] wl[79] vdd gnd cell_6t
Xbit_r80_c65 bl[65] br[65] wl[80] vdd gnd cell_6t
Xbit_r81_c65 bl[65] br[65] wl[81] vdd gnd cell_6t
Xbit_r82_c65 bl[65] br[65] wl[82] vdd gnd cell_6t
Xbit_r83_c65 bl[65] br[65] wl[83] vdd gnd cell_6t
Xbit_r84_c65 bl[65] br[65] wl[84] vdd gnd cell_6t
Xbit_r85_c65 bl[65] br[65] wl[85] vdd gnd cell_6t
Xbit_r86_c65 bl[65] br[65] wl[86] vdd gnd cell_6t
Xbit_r87_c65 bl[65] br[65] wl[87] vdd gnd cell_6t
Xbit_r88_c65 bl[65] br[65] wl[88] vdd gnd cell_6t
Xbit_r89_c65 bl[65] br[65] wl[89] vdd gnd cell_6t
Xbit_r90_c65 bl[65] br[65] wl[90] vdd gnd cell_6t
Xbit_r91_c65 bl[65] br[65] wl[91] vdd gnd cell_6t
Xbit_r92_c65 bl[65] br[65] wl[92] vdd gnd cell_6t
Xbit_r93_c65 bl[65] br[65] wl[93] vdd gnd cell_6t
Xbit_r94_c65 bl[65] br[65] wl[94] vdd gnd cell_6t
Xbit_r95_c65 bl[65] br[65] wl[95] vdd gnd cell_6t
Xbit_r96_c65 bl[65] br[65] wl[96] vdd gnd cell_6t
Xbit_r97_c65 bl[65] br[65] wl[97] vdd gnd cell_6t
Xbit_r98_c65 bl[65] br[65] wl[98] vdd gnd cell_6t
Xbit_r99_c65 bl[65] br[65] wl[99] vdd gnd cell_6t
Xbit_r100_c65 bl[65] br[65] wl[100] vdd gnd cell_6t
Xbit_r101_c65 bl[65] br[65] wl[101] vdd gnd cell_6t
Xbit_r102_c65 bl[65] br[65] wl[102] vdd gnd cell_6t
Xbit_r103_c65 bl[65] br[65] wl[103] vdd gnd cell_6t
Xbit_r104_c65 bl[65] br[65] wl[104] vdd gnd cell_6t
Xbit_r105_c65 bl[65] br[65] wl[105] vdd gnd cell_6t
Xbit_r106_c65 bl[65] br[65] wl[106] vdd gnd cell_6t
Xbit_r107_c65 bl[65] br[65] wl[107] vdd gnd cell_6t
Xbit_r108_c65 bl[65] br[65] wl[108] vdd gnd cell_6t
Xbit_r109_c65 bl[65] br[65] wl[109] vdd gnd cell_6t
Xbit_r110_c65 bl[65] br[65] wl[110] vdd gnd cell_6t
Xbit_r111_c65 bl[65] br[65] wl[111] vdd gnd cell_6t
Xbit_r112_c65 bl[65] br[65] wl[112] vdd gnd cell_6t
Xbit_r113_c65 bl[65] br[65] wl[113] vdd gnd cell_6t
Xbit_r114_c65 bl[65] br[65] wl[114] vdd gnd cell_6t
Xbit_r115_c65 bl[65] br[65] wl[115] vdd gnd cell_6t
Xbit_r116_c65 bl[65] br[65] wl[116] vdd gnd cell_6t
Xbit_r117_c65 bl[65] br[65] wl[117] vdd gnd cell_6t
Xbit_r118_c65 bl[65] br[65] wl[118] vdd gnd cell_6t
Xbit_r119_c65 bl[65] br[65] wl[119] vdd gnd cell_6t
Xbit_r120_c65 bl[65] br[65] wl[120] vdd gnd cell_6t
Xbit_r121_c65 bl[65] br[65] wl[121] vdd gnd cell_6t
Xbit_r122_c65 bl[65] br[65] wl[122] vdd gnd cell_6t
Xbit_r123_c65 bl[65] br[65] wl[123] vdd gnd cell_6t
Xbit_r124_c65 bl[65] br[65] wl[124] vdd gnd cell_6t
Xbit_r125_c65 bl[65] br[65] wl[125] vdd gnd cell_6t
Xbit_r126_c65 bl[65] br[65] wl[126] vdd gnd cell_6t
Xbit_r127_c65 bl[65] br[65] wl[127] vdd gnd cell_6t
Xbit_r0_c66 bl[66] br[66] wl[0] vdd gnd cell_6t
Xbit_r1_c66 bl[66] br[66] wl[1] vdd gnd cell_6t
Xbit_r2_c66 bl[66] br[66] wl[2] vdd gnd cell_6t
Xbit_r3_c66 bl[66] br[66] wl[3] vdd gnd cell_6t
Xbit_r4_c66 bl[66] br[66] wl[4] vdd gnd cell_6t
Xbit_r5_c66 bl[66] br[66] wl[5] vdd gnd cell_6t
Xbit_r6_c66 bl[66] br[66] wl[6] vdd gnd cell_6t
Xbit_r7_c66 bl[66] br[66] wl[7] vdd gnd cell_6t
Xbit_r8_c66 bl[66] br[66] wl[8] vdd gnd cell_6t
Xbit_r9_c66 bl[66] br[66] wl[9] vdd gnd cell_6t
Xbit_r10_c66 bl[66] br[66] wl[10] vdd gnd cell_6t
Xbit_r11_c66 bl[66] br[66] wl[11] vdd gnd cell_6t
Xbit_r12_c66 bl[66] br[66] wl[12] vdd gnd cell_6t
Xbit_r13_c66 bl[66] br[66] wl[13] vdd gnd cell_6t
Xbit_r14_c66 bl[66] br[66] wl[14] vdd gnd cell_6t
Xbit_r15_c66 bl[66] br[66] wl[15] vdd gnd cell_6t
Xbit_r16_c66 bl[66] br[66] wl[16] vdd gnd cell_6t
Xbit_r17_c66 bl[66] br[66] wl[17] vdd gnd cell_6t
Xbit_r18_c66 bl[66] br[66] wl[18] vdd gnd cell_6t
Xbit_r19_c66 bl[66] br[66] wl[19] vdd gnd cell_6t
Xbit_r20_c66 bl[66] br[66] wl[20] vdd gnd cell_6t
Xbit_r21_c66 bl[66] br[66] wl[21] vdd gnd cell_6t
Xbit_r22_c66 bl[66] br[66] wl[22] vdd gnd cell_6t
Xbit_r23_c66 bl[66] br[66] wl[23] vdd gnd cell_6t
Xbit_r24_c66 bl[66] br[66] wl[24] vdd gnd cell_6t
Xbit_r25_c66 bl[66] br[66] wl[25] vdd gnd cell_6t
Xbit_r26_c66 bl[66] br[66] wl[26] vdd gnd cell_6t
Xbit_r27_c66 bl[66] br[66] wl[27] vdd gnd cell_6t
Xbit_r28_c66 bl[66] br[66] wl[28] vdd gnd cell_6t
Xbit_r29_c66 bl[66] br[66] wl[29] vdd gnd cell_6t
Xbit_r30_c66 bl[66] br[66] wl[30] vdd gnd cell_6t
Xbit_r31_c66 bl[66] br[66] wl[31] vdd gnd cell_6t
Xbit_r32_c66 bl[66] br[66] wl[32] vdd gnd cell_6t
Xbit_r33_c66 bl[66] br[66] wl[33] vdd gnd cell_6t
Xbit_r34_c66 bl[66] br[66] wl[34] vdd gnd cell_6t
Xbit_r35_c66 bl[66] br[66] wl[35] vdd gnd cell_6t
Xbit_r36_c66 bl[66] br[66] wl[36] vdd gnd cell_6t
Xbit_r37_c66 bl[66] br[66] wl[37] vdd gnd cell_6t
Xbit_r38_c66 bl[66] br[66] wl[38] vdd gnd cell_6t
Xbit_r39_c66 bl[66] br[66] wl[39] vdd gnd cell_6t
Xbit_r40_c66 bl[66] br[66] wl[40] vdd gnd cell_6t
Xbit_r41_c66 bl[66] br[66] wl[41] vdd gnd cell_6t
Xbit_r42_c66 bl[66] br[66] wl[42] vdd gnd cell_6t
Xbit_r43_c66 bl[66] br[66] wl[43] vdd gnd cell_6t
Xbit_r44_c66 bl[66] br[66] wl[44] vdd gnd cell_6t
Xbit_r45_c66 bl[66] br[66] wl[45] vdd gnd cell_6t
Xbit_r46_c66 bl[66] br[66] wl[46] vdd gnd cell_6t
Xbit_r47_c66 bl[66] br[66] wl[47] vdd gnd cell_6t
Xbit_r48_c66 bl[66] br[66] wl[48] vdd gnd cell_6t
Xbit_r49_c66 bl[66] br[66] wl[49] vdd gnd cell_6t
Xbit_r50_c66 bl[66] br[66] wl[50] vdd gnd cell_6t
Xbit_r51_c66 bl[66] br[66] wl[51] vdd gnd cell_6t
Xbit_r52_c66 bl[66] br[66] wl[52] vdd gnd cell_6t
Xbit_r53_c66 bl[66] br[66] wl[53] vdd gnd cell_6t
Xbit_r54_c66 bl[66] br[66] wl[54] vdd gnd cell_6t
Xbit_r55_c66 bl[66] br[66] wl[55] vdd gnd cell_6t
Xbit_r56_c66 bl[66] br[66] wl[56] vdd gnd cell_6t
Xbit_r57_c66 bl[66] br[66] wl[57] vdd gnd cell_6t
Xbit_r58_c66 bl[66] br[66] wl[58] vdd gnd cell_6t
Xbit_r59_c66 bl[66] br[66] wl[59] vdd gnd cell_6t
Xbit_r60_c66 bl[66] br[66] wl[60] vdd gnd cell_6t
Xbit_r61_c66 bl[66] br[66] wl[61] vdd gnd cell_6t
Xbit_r62_c66 bl[66] br[66] wl[62] vdd gnd cell_6t
Xbit_r63_c66 bl[66] br[66] wl[63] vdd gnd cell_6t
Xbit_r64_c66 bl[66] br[66] wl[64] vdd gnd cell_6t
Xbit_r65_c66 bl[66] br[66] wl[65] vdd gnd cell_6t
Xbit_r66_c66 bl[66] br[66] wl[66] vdd gnd cell_6t
Xbit_r67_c66 bl[66] br[66] wl[67] vdd gnd cell_6t
Xbit_r68_c66 bl[66] br[66] wl[68] vdd gnd cell_6t
Xbit_r69_c66 bl[66] br[66] wl[69] vdd gnd cell_6t
Xbit_r70_c66 bl[66] br[66] wl[70] vdd gnd cell_6t
Xbit_r71_c66 bl[66] br[66] wl[71] vdd gnd cell_6t
Xbit_r72_c66 bl[66] br[66] wl[72] vdd gnd cell_6t
Xbit_r73_c66 bl[66] br[66] wl[73] vdd gnd cell_6t
Xbit_r74_c66 bl[66] br[66] wl[74] vdd gnd cell_6t
Xbit_r75_c66 bl[66] br[66] wl[75] vdd gnd cell_6t
Xbit_r76_c66 bl[66] br[66] wl[76] vdd gnd cell_6t
Xbit_r77_c66 bl[66] br[66] wl[77] vdd gnd cell_6t
Xbit_r78_c66 bl[66] br[66] wl[78] vdd gnd cell_6t
Xbit_r79_c66 bl[66] br[66] wl[79] vdd gnd cell_6t
Xbit_r80_c66 bl[66] br[66] wl[80] vdd gnd cell_6t
Xbit_r81_c66 bl[66] br[66] wl[81] vdd gnd cell_6t
Xbit_r82_c66 bl[66] br[66] wl[82] vdd gnd cell_6t
Xbit_r83_c66 bl[66] br[66] wl[83] vdd gnd cell_6t
Xbit_r84_c66 bl[66] br[66] wl[84] vdd gnd cell_6t
Xbit_r85_c66 bl[66] br[66] wl[85] vdd gnd cell_6t
Xbit_r86_c66 bl[66] br[66] wl[86] vdd gnd cell_6t
Xbit_r87_c66 bl[66] br[66] wl[87] vdd gnd cell_6t
Xbit_r88_c66 bl[66] br[66] wl[88] vdd gnd cell_6t
Xbit_r89_c66 bl[66] br[66] wl[89] vdd gnd cell_6t
Xbit_r90_c66 bl[66] br[66] wl[90] vdd gnd cell_6t
Xbit_r91_c66 bl[66] br[66] wl[91] vdd gnd cell_6t
Xbit_r92_c66 bl[66] br[66] wl[92] vdd gnd cell_6t
Xbit_r93_c66 bl[66] br[66] wl[93] vdd gnd cell_6t
Xbit_r94_c66 bl[66] br[66] wl[94] vdd gnd cell_6t
Xbit_r95_c66 bl[66] br[66] wl[95] vdd gnd cell_6t
Xbit_r96_c66 bl[66] br[66] wl[96] vdd gnd cell_6t
Xbit_r97_c66 bl[66] br[66] wl[97] vdd gnd cell_6t
Xbit_r98_c66 bl[66] br[66] wl[98] vdd gnd cell_6t
Xbit_r99_c66 bl[66] br[66] wl[99] vdd gnd cell_6t
Xbit_r100_c66 bl[66] br[66] wl[100] vdd gnd cell_6t
Xbit_r101_c66 bl[66] br[66] wl[101] vdd gnd cell_6t
Xbit_r102_c66 bl[66] br[66] wl[102] vdd gnd cell_6t
Xbit_r103_c66 bl[66] br[66] wl[103] vdd gnd cell_6t
Xbit_r104_c66 bl[66] br[66] wl[104] vdd gnd cell_6t
Xbit_r105_c66 bl[66] br[66] wl[105] vdd gnd cell_6t
Xbit_r106_c66 bl[66] br[66] wl[106] vdd gnd cell_6t
Xbit_r107_c66 bl[66] br[66] wl[107] vdd gnd cell_6t
Xbit_r108_c66 bl[66] br[66] wl[108] vdd gnd cell_6t
Xbit_r109_c66 bl[66] br[66] wl[109] vdd gnd cell_6t
Xbit_r110_c66 bl[66] br[66] wl[110] vdd gnd cell_6t
Xbit_r111_c66 bl[66] br[66] wl[111] vdd gnd cell_6t
Xbit_r112_c66 bl[66] br[66] wl[112] vdd gnd cell_6t
Xbit_r113_c66 bl[66] br[66] wl[113] vdd gnd cell_6t
Xbit_r114_c66 bl[66] br[66] wl[114] vdd gnd cell_6t
Xbit_r115_c66 bl[66] br[66] wl[115] vdd gnd cell_6t
Xbit_r116_c66 bl[66] br[66] wl[116] vdd gnd cell_6t
Xbit_r117_c66 bl[66] br[66] wl[117] vdd gnd cell_6t
Xbit_r118_c66 bl[66] br[66] wl[118] vdd gnd cell_6t
Xbit_r119_c66 bl[66] br[66] wl[119] vdd gnd cell_6t
Xbit_r120_c66 bl[66] br[66] wl[120] vdd gnd cell_6t
Xbit_r121_c66 bl[66] br[66] wl[121] vdd gnd cell_6t
Xbit_r122_c66 bl[66] br[66] wl[122] vdd gnd cell_6t
Xbit_r123_c66 bl[66] br[66] wl[123] vdd gnd cell_6t
Xbit_r124_c66 bl[66] br[66] wl[124] vdd gnd cell_6t
Xbit_r125_c66 bl[66] br[66] wl[125] vdd gnd cell_6t
Xbit_r126_c66 bl[66] br[66] wl[126] vdd gnd cell_6t
Xbit_r127_c66 bl[66] br[66] wl[127] vdd gnd cell_6t
Xbit_r0_c67 bl[67] br[67] wl[0] vdd gnd cell_6t
Xbit_r1_c67 bl[67] br[67] wl[1] vdd gnd cell_6t
Xbit_r2_c67 bl[67] br[67] wl[2] vdd gnd cell_6t
Xbit_r3_c67 bl[67] br[67] wl[3] vdd gnd cell_6t
Xbit_r4_c67 bl[67] br[67] wl[4] vdd gnd cell_6t
Xbit_r5_c67 bl[67] br[67] wl[5] vdd gnd cell_6t
Xbit_r6_c67 bl[67] br[67] wl[6] vdd gnd cell_6t
Xbit_r7_c67 bl[67] br[67] wl[7] vdd gnd cell_6t
Xbit_r8_c67 bl[67] br[67] wl[8] vdd gnd cell_6t
Xbit_r9_c67 bl[67] br[67] wl[9] vdd gnd cell_6t
Xbit_r10_c67 bl[67] br[67] wl[10] vdd gnd cell_6t
Xbit_r11_c67 bl[67] br[67] wl[11] vdd gnd cell_6t
Xbit_r12_c67 bl[67] br[67] wl[12] vdd gnd cell_6t
Xbit_r13_c67 bl[67] br[67] wl[13] vdd gnd cell_6t
Xbit_r14_c67 bl[67] br[67] wl[14] vdd gnd cell_6t
Xbit_r15_c67 bl[67] br[67] wl[15] vdd gnd cell_6t
Xbit_r16_c67 bl[67] br[67] wl[16] vdd gnd cell_6t
Xbit_r17_c67 bl[67] br[67] wl[17] vdd gnd cell_6t
Xbit_r18_c67 bl[67] br[67] wl[18] vdd gnd cell_6t
Xbit_r19_c67 bl[67] br[67] wl[19] vdd gnd cell_6t
Xbit_r20_c67 bl[67] br[67] wl[20] vdd gnd cell_6t
Xbit_r21_c67 bl[67] br[67] wl[21] vdd gnd cell_6t
Xbit_r22_c67 bl[67] br[67] wl[22] vdd gnd cell_6t
Xbit_r23_c67 bl[67] br[67] wl[23] vdd gnd cell_6t
Xbit_r24_c67 bl[67] br[67] wl[24] vdd gnd cell_6t
Xbit_r25_c67 bl[67] br[67] wl[25] vdd gnd cell_6t
Xbit_r26_c67 bl[67] br[67] wl[26] vdd gnd cell_6t
Xbit_r27_c67 bl[67] br[67] wl[27] vdd gnd cell_6t
Xbit_r28_c67 bl[67] br[67] wl[28] vdd gnd cell_6t
Xbit_r29_c67 bl[67] br[67] wl[29] vdd gnd cell_6t
Xbit_r30_c67 bl[67] br[67] wl[30] vdd gnd cell_6t
Xbit_r31_c67 bl[67] br[67] wl[31] vdd gnd cell_6t
Xbit_r32_c67 bl[67] br[67] wl[32] vdd gnd cell_6t
Xbit_r33_c67 bl[67] br[67] wl[33] vdd gnd cell_6t
Xbit_r34_c67 bl[67] br[67] wl[34] vdd gnd cell_6t
Xbit_r35_c67 bl[67] br[67] wl[35] vdd gnd cell_6t
Xbit_r36_c67 bl[67] br[67] wl[36] vdd gnd cell_6t
Xbit_r37_c67 bl[67] br[67] wl[37] vdd gnd cell_6t
Xbit_r38_c67 bl[67] br[67] wl[38] vdd gnd cell_6t
Xbit_r39_c67 bl[67] br[67] wl[39] vdd gnd cell_6t
Xbit_r40_c67 bl[67] br[67] wl[40] vdd gnd cell_6t
Xbit_r41_c67 bl[67] br[67] wl[41] vdd gnd cell_6t
Xbit_r42_c67 bl[67] br[67] wl[42] vdd gnd cell_6t
Xbit_r43_c67 bl[67] br[67] wl[43] vdd gnd cell_6t
Xbit_r44_c67 bl[67] br[67] wl[44] vdd gnd cell_6t
Xbit_r45_c67 bl[67] br[67] wl[45] vdd gnd cell_6t
Xbit_r46_c67 bl[67] br[67] wl[46] vdd gnd cell_6t
Xbit_r47_c67 bl[67] br[67] wl[47] vdd gnd cell_6t
Xbit_r48_c67 bl[67] br[67] wl[48] vdd gnd cell_6t
Xbit_r49_c67 bl[67] br[67] wl[49] vdd gnd cell_6t
Xbit_r50_c67 bl[67] br[67] wl[50] vdd gnd cell_6t
Xbit_r51_c67 bl[67] br[67] wl[51] vdd gnd cell_6t
Xbit_r52_c67 bl[67] br[67] wl[52] vdd gnd cell_6t
Xbit_r53_c67 bl[67] br[67] wl[53] vdd gnd cell_6t
Xbit_r54_c67 bl[67] br[67] wl[54] vdd gnd cell_6t
Xbit_r55_c67 bl[67] br[67] wl[55] vdd gnd cell_6t
Xbit_r56_c67 bl[67] br[67] wl[56] vdd gnd cell_6t
Xbit_r57_c67 bl[67] br[67] wl[57] vdd gnd cell_6t
Xbit_r58_c67 bl[67] br[67] wl[58] vdd gnd cell_6t
Xbit_r59_c67 bl[67] br[67] wl[59] vdd gnd cell_6t
Xbit_r60_c67 bl[67] br[67] wl[60] vdd gnd cell_6t
Xbit_r61_c67 bl[67] br[67] wl[61] vdd gnd cell_6t
Xbit_r62_c67 bl[67] br[67] wl[62] vdd gnd cell_6t
Xbit_r63_c67 bl[67] br[67] wl[63] vdd gnd cell_6t
Xbit_r64_c67 bl[67] br[67] wl[64] vdd gnd cell_6t
Xbit_r65_c67 bl[67] br[67] wl[65] vdd gnd cell_6t
Xbit_r66_c67 bl[67] br[67] wl[66] vdd gnd cell_6t
Xbit_r67_c67 bl[67] br[67] wl[67] vdd gnd cell_6t
Xbit_r68_c67 bl[67] br[67] wl[68] vdd gnd cell_6t
Xbit_r69_c67 bl[67] br[67] wl[69] vdd gnd cell_6t
Xbit_r70_c67 bl[67] br[67] wl[70] vdd gnd cell_6t
Xbit_r71_c67 bl[67] br[67] wl[71] vdd gnd cell_6t
Xbit_r72_c67 bl[67] br[67] wl[72] vdd gnd cell_6t
Xbit_r73_c67 bl[67] br[67] wl[73] vdd gnd cell_6t
Xbit_r74_c67 bl[67] br[67] wl[74] vdd gnd cell_6t
Xbit_r75_c67 bl[67] br[67] wl[75] vdd gnd cell_6t
Xbit_r76_c67 bl[67] br[67] wl[76] vdd gnd cell_6t
Xbit_r77_c67 bl[67] br[67] wl[77] vdd gnd cell_6t
Xbit_r78_c67 bl[67] br[67] wl[78] vdd gnd cell_6t
Xbit_r79_c67 bl[67] br[67] wl[79] vdd gnd cell_6t
Xbit_r80_c67 bl[67] br[67] wl[80] vdd gnd cell_6t
Xbit_r81_c67 bl[67] br[67] wl[81] vdd gnd cell_6t
Xbit_r82_c67 bl[67] br[67] wl[82] vdd gnd cell_6t
Xbit_r83_c67 bl[67] br[67] wl[83] vdd gnd cell_6t
Xbit_r84_c67 bl[67] br[67] wl[84] vdd gnd cell_6t
Xbit_r85_c67 bl[67] br[67] wl[85] vdd gnd cell_6t
Xbit_r86_c67 bl[67] br[67] wl[86] vdd gnd cell_6t
Xbit_r87_c67 bl[67] br[67] wl[87] vdd gnd cell_6t
Xbit_r88_c67 bl[67] br[67] wl[88] vdd gnd cell_6t
Xbit_r89_c67 bl[67] br[67] wl[89] vdd gnd cell_6t
Xbit_r90_c67 bl[67] br[67] wl[90] vdd gnd cell_6t
Xbit_r91_c67 bl[67] br[67] wl[91] vdd gnd cell_6t
Xbit_r92_c67 bl[67] br[67] wl[92] vdd gnd cell_6t
Xbit_r93_c67 bl[67] br[67] wl[93] vdd gnd cell_6t
Xbit_r94_c67 bl[67] br[67] wl[94] vdd gnd cell_6t
Xbit_r95_c67 bl[67] br[67] wl[95] vdd gnd cell_6t
Xbit_r96_c67 bl[67] br[67] wl[96] vdd gnd cell_6t
Xbit_r97_c67 bl[67] br[67] wl[97] vdd gnd cell_6t
Xbit_r98_c67 bl[67] br[67] wl[98] vdd gnd cell_6t
Xbit_r99_c67 bl[67] br[67] wl[99] vdd gnd cell_6t
Xbit_r100_c67 bl[67] br[67] wl[100] vdd gnd cell_6t
Xbit_r101_c67 bl[67] br[67] wl[101] vdd gnd cell_6t
Xbit_r102_c67 bl[67] br[67] wl[102] vdd gnd cell_6t
Xbit_r103_c67 bl[67] br[67] wl[103] vdd gnd cell_6t
Xbit_r104_c67 bl[67] br[67] wl[104] vdd gnd cell_6t
Xbit_r105_c67 bl[67] br[67] wl[105] vdd gnd cell_6t
Xbit_r106_c67 bl[67] br[67] wl[106] vdd gnd cell_6t
Xbit_r107_c67 bl[67] br[67] wl[107] vdd gnd cell_6t
Xbit_r108_c67 bl[67] br[67] wl[108] vdd gnd cell_6t
Xbit_r109_c67 bl[67] br[67] wl[109] vdd gnd cell_6t
Xbit_r110_c67 bl[67] br[67] wl[110] vdd gnd cell_6t
Xbit_r111_c67 bl[67] br[67] wl[111] vdd gnd cell_6t
Xbit_r112_c67 bl[67] br[67] wl[112] vdd gnd cell_6t
Xbit_r113_c67 bl[67] br[67] wl[113] vdd gnd cell_6t
Xbit_r114_c67 bl[67] br[67] wl[114] vdd gnd cell_6t
Xbit_r115_c67 bl[67] br[67] wl[115] vdd gnd cell_6t
Xbit_r116_c67 bl[67] br[67] wl[116] vdd gnd cell_6t
Xbit_r117_c67 bl[67] br[67] wl[117] vdd gnd cell_6t
Xbit_r118_c67 bl[67] br[67] wl[118] vdd gnd cell_6t
Xbit_r119_c67 bl[67] br[67] wl[119] vdd gnd cell_6t
Xbit_r120_c67 bl[67] br[67] wl[120] vdd gnd cell_6t
Xbit_r121_c67 bl[67] br[67] wl[121] vdd gnd cell_6t
Xbit_r122_c67 bl[67] br[67] wl[122] vdd gnd cell_6t
Xbit_r123_c67 bl[67] br[67] wl[123] vdd gnd cell_6t
Xbit_r124_c67 bl[67] br[67] wl[124] vdd gnd cell_6t
Xbit_r125_c67 bl[67] br[67] wl[125] vdd gnd cell_6t
Xbit_r126_c67 bl[67] br[67] wl[126] vdd gnd cell_6t
Xbit_r127_c67 bl[67] br[67] wl[127] vdd gnd cell_6t
Xbit_r0_c68 bl[68] br[68] wl[0] vdd gnd cell_6t
Xbit_r1_c68 bl[68] br[68] wl[1] vdd gnd cell_6t
Xbit_r2_c68 bl[68] br[68] wl[2] vdd gnd cell_6t
Xbit_r3_c68 bl[68] br[68] wl[3] vdd gnd cell_6t
Xbit_r4_c68 bl[68] br[68] wl[4] vdd gnd cell_6t
Xbit_r5_c68 bl[68] br[68] wl[5] vdd gnd cell_6t
Xbit_r6_c68 bl[68] br[68] wl[6] vdd gnd cell_6t
Xbit_r7_c68 bl[68] br[68] wl[7] vdd gnd cell_6t
Xbit_r8_c68 bl[68] br[68] wl[8] vdd gnd cell_6t
Xbit_r9_c68 bl[68] br[68] wl[9] vdd gnd cell_6t
Xbit_r10_c68 bl[68] br[68] wl[10] vdd gnd cell_6t
Xbit_r11_c68 bl[68] br[68] wl[11] vdd gnd cell_6t
Xbit_r12_c68 bl[68] br[68] wl[12] vdd gnd cell_6t
Xbit_r13_c68 bl[68] br[68] wl[13] vdd gnd cell_6t
Xbit_r14_c68 bl[68] br[68] wl[14] vdd gnd cell_6t
Xbit_r15_c68 bl[68] br[68] wl[15] vdd gnd cell_6t
Xbit_r16_c68 bl[68] br[68] wl[16] vdd gnd cell_6t
Xbit_r17_c68 bl[68] br[68] wl[17] vdd gnd cell_6t
Xbit_r18_c68 bl[68] br[68] wl[18] vdd gnd cell_6t
Xbit_r19_c68 bl[68] br[68] wl[19] vdd gnd cell_6t
Xbit_r20_c68 bl[68] br[68] wl[20] vdd gnd cell_6t
Xbit_r21_c68 bl[68] br[68] wl[21] vdd gnd cell_6t
Xbit_r22_c68 bl[68] br[68] wl[22] vdd gnd cell_6t
Xbit_r23_c68 bl[68] br[68] wl[23] vdd gnd cell_6t
Xbit_r24_c68 bl[68] br[68] wl[24] vdd gnd cell_6t
Xbit_r25_c68 bl[68] br[68] wl[25] vdd gnd cell_6t
Xbit_r26_c68 bl[68] br[68] wl[26] vdd gnd cell_6t
Xbit_r27_c68 bl[68] br[68] wl[27] vdd gnd cell_6t
Xbit_r28_c68 bl[68] br[68] wl[28] vdd gnd cell_6t
Xbit_r29_c68 bl[68] br[68] wl[29] vdd gnd cell_6t
Xbit_r30_c68 bl[68] br[68] wl[30] vdd gnd cell_6t
Xbit_r31_c68 bl[68] br[68] wl[31] vdd gnd cell_6t
Xbit_r32_c68 bl[68] br[68] wl[32] vdd gnd cell_6t
Xbit_r33_c68 bl[68] br[68] wl[33] vdd gnd cell_6t
Xbit_r34_c68 bl[68] br[68] wl[34] vdd gnd cell_6t
Xbit_r35_c68 bl[68] br[68] wl[35] vdd gnd cell_6t
Xbit_r36_c68 bl[68] br[68] wl[36] vdd gnd cell_6t
Xbit_r37_c68 bl[68] br[68] wl[37] vdd gnd cell_6t
Xbit_r38_c68 bl[68] br[68] wl[38] vdd gnd cell_6t
Xbit_r39_c68 bl[68] br[68] wl[39] vdd gnd cell_6t
Xbit_r40_c68 bl[68] br[68] wl[40] vdd gnd cell_6t
Xbit_r41_c68 bl[68] br[68] wl[41] vdd gnd cell_6t
Xbit_r42_c68 bl[68] br[68] wl[42] vdd gnd cell_6t
Xbit_r43_c68 bl[68] br[68] wl[43] vdd gnd cell_6t
Xbit_r44_c68 bl[68] br[68] wl[44] vdd gnd cell_6t
Xbit_r45_c68 bl[68] br[68] wl[45] vdd gnd cell_6t
Xbit_r46_c68 bl[68] br[68] wl[46] vdd gnd cell_6t
Xbit_r47_c68 bl[68] br[68] wl[47] vdd gnd cell_6t
Xbit_r48_c68 bl[68] br[68] wl[48] vdd gnd cell_6t
Xbit_r49_c68 bl[68] br[68] wl[49] vdd gnd cell_6t
Xbit_r50_c68 bl[68] br[68] wl[50] vdd gnd cell_6t
Xbit_r51_c68 bl[68] br[68] wl[51] vdd gnd cell_6t
Xbit_r52_c68 bl[68] br[68] wl[52] vdd gnd cell_6t
Xbit_r53_c68 bl[68] br[68] wl[53] vdd gnd cell_6t
Xbit_r54_c68 bl[68] br[68] wl[54] vdd gnd cell_6t
Xbit_r55_c68 bl[68] br[68] wl[55] vdd gnd cell_6t
Xbit_r56_c68 bl[68] br[68] wl[56] vdd gnd cell_6t
Xbit_r57_c68 bl[68] br[68] wl[57] vdd gnd cell_6t
Xbit_r58_c68 bl[68] br[68] wl[58] vdd gnd cell_6t
Xbit_r59_c68 bl[68] br[68] wl[59] vdd gnd cell_6t
Xbit_r60_c68 bl[68] br[68] wl[60] vdd gnd cell_6t
Xbit_r61_c68 bl[68] br[68] wl[61] vdd gnd cell_6t
Xbit_r62_c68 bl[68] br[68] wl[62] vdd gnd cell_6t
Xbit_r63_c68 bl[68] br[68] wl[63] vdd gnd cell_6t
Xbit_r64_c68 bl[68] br[68] wl[64] vdd gnd cell_6t
Xbit_r65_c68 bl[68] br[68] wl[65] vdd gnd cell_6t
Xbit_r66_c68 bl[68] br[68] wl[66] vdd gnd cell_6t
Xbit_r67_c68 bl[68] br[68] wl[67] vdd gnd cell_6t
Xbit_r68_c68 bl[68] br[68] wl[68] vdd gnd cell_6t
Xbit_r69_c68 bl[68] br[68] wl[69] vdd gnd cell_6t
Xbit_r70_c68 bl[68] br[68] wl[70] vdd gnd cell_6t
Xbit_r71_c68 bl[68] br[68] wl[71] vdd gnd cell_6t
Xbit_r72_c68 bl[68] br[68] wl[72] vdd gnd cell_6t
Xbit_r73_c68 bl[68] br[68] wl[73] vdd gnd cell_6t
Xbit_r74_c68 bl[68] br[68] wl[74] vdd gnd cell_6t
Xbit_r75_c68 bl[68] br[68] wl[75] vdd gnd cell_6t
Xbit_r76_c68 bl[68] br[68] wl[76] vdd gnd cell_6t
Xbit_r77_c68 bl[68] br[68] wl[77] vdd gnd cell_6t
Xbit_r78_c68 bl[68] br[68] wl[78] vdd gnd cell_6t
Xbit_r79_c68 bl[68] br[68] wl[79] vdd gnd cell_6t
Xbit_r80_c68 bl[68] br[68] wl[80] vdd gnd cell_6t
Xbit_r81_c68 bl[68] br[68] wl[81] vdd gnd cell_6t
Xbit_r82_c68 bl[68] br[68] wl[82] vdd gnd cell_6t
Xbit_r83_c68 bl[68] br[68] wl[83] vdd gnd cell_6t
Xbit_r84_c68 bl[68] br[68] wl[84] vdd gnd cell_6t
Xbit_r85_c68 bl[68] br[68] wl[85] vdd gnd cell_6t
Xbit_r86_c68 bl[68] br[68] wl[86] vdd gnd cell_6t
Xbit_r87_c68 bl[68] br[68] wl[87] vdd gnd cell_6t
Xbit_r88_c68 bl[68] br[68] wl[88] vdd gnd cell_6t
Xbit_r89_c68 bl[68] br[68] wl[89] vdd gnd cell_6t
Xbit_r90_c68 bl[68] br[68] wl[90] vdd gnd cell_6t
Xbit_r91_c68 bl[68] br[68] wl[91] vdd gnd cell_6t
Xbit_r92_c68 bl[68] br[68] wl[92] vdd gnd cell_6t
Xbit_r93_c68 bl[68] br[68] wl[93] vdd gnd cell_6t
Xbit_r94_c68 bl[68] br[68] wl[94] vdd gnd cell_6t
Xbit_r95_c68 bl[68] br[68] wl[95] vdd gnd cell_6t
Xbit_r96_c68 bl[68] br[68] wl[96] vdd gnd cell_6t
Xbit_r97_c68 bl[68] br[68] wl[97] vdd gnd cell_6t
Xbit_r98_c68 bl[68] br[68] wl[98] vdd gnd cell_6t
Xbit_r99_c68 bl[68] br[68] wl[99] vdd gnd cell_6t
Xbit_r100_c68 bl[68] br[68] wl[100] vdd gnd cell_6t
Xbit_r101_c68 bl[68] br[68] wl[101] vdd gnd cell_6t
Xbit_r102_c68 bl[68] br[68] wl[102] vdd gnd cell_6t
Xbit_r103_c68 bl[68] br[68] wl[103] vdd gnd cell_6t
Xbit_r104_c68 bl[68] br[68] wl[104] vdd gnd cell_6t
Xbit_r105_c68 bl[68] br[68] wl[105] vdd gnd cell_6t
Xbit_r106_c68 bl[68] br[68] wl[106] vdd gnd cell_6t
Xbit_r107_c68 bl[68] br[68] wl[107] vdd gnd cell_6t
Xbit_r108_c68 bl[68] br[68] wl[108] vdd gnd cell_6t
Xbit_r109_c68 bl[68] br[68] wl[109] vdd gnd cell_6t
Xbit_r110_c68 bl[68] br[68] wl[110] vdd gnd cell_6t
Xbit_r111_c68 bl[68] br[68] wl[111] vdd gnd cell_6t
Xbit_r112_c68 bl[68] br[68] wl[112] vdd gnd cell_6t
Xbit_r113_c68 bl[68] br[68] wl[113] vdd gnd cell_6t
Xbit_r114_c68 bl[68] br[68] wl[114] vdd gnd cell_6t
Xbit_r115_c68 bl[68] br[68] wl[115] vdd gnd cell_6t
Xbit_r116_c68 bl[68] br[68] wl[116] vdd gnd cell_6t
Xbit_r117_c68 bl[68] br[68] wl[117] vdd gnd cell_6t
Xbit_r118_c68 bl[68] br[68] wl[118] vdd gnd cell_6t
Xbit_r119_c68 bl[68] br[68] wl[119] vdd gnd cell_6t
Xbit_r120_c68 bl[68] br[68] wl[120] vdd gnd cell_6t
Xbit_r121_c68 bl[68] br[68] wl[121] vdd gnd cell_6t
Xbit_r122_c68 bl[68] br[68] wl[122] vdd gnd cell_6t
Xbit_r123_c68 bl[68] br[68] wl[123] vdd gnd cell_6t
Xbit_r124_c68 bl[68] br[68] wl[124] vdd gnd cell_6t
Xbit_r125_c68 bl[68] br[68] wl[125] vdd gnd cell_6t
Xbit_r126_c68 bl[68] br[68] wl[126] vdd gnd cell_6t
Xbit_r127_c68 bl[68] br[68] wl[127] vdd gnd cell_6t
Xbit_r0_c69 bl[69] br[69] wl[0] vdd gnd cell_6t
Xbit_r1_c69 bl[69] br[69] wl[1] vdd gnd cell_6t
Xbit_r2_c69 bl[69] br[69] wl[2] vdd gnd cell_6t
Xbit_r3_c69 bl[69] br[69] wl[3] vdd gnd cell_6t
Xbit_r4_c69 bl[69] br[69] wl[4] vdd gnd cell_6t
Xbit_r5_c69 bl[69] br[69] wl[5] vdd gnd cell_6t
Xbit_r6_c69 bl[69] br[69] wl[6] vdd gnd cell_6t
Xbit_r7_c69 bl[69] br[69] wl[7] vdd gnd cell_6t
Xbit_r8_c69 bl[69] br[69] wl[8] vdd gnd cell_6t
Xbit_r9_c69 bl[69] br[69] wl[9] vdd gnd cell_6t
Xbit_r10_c69 bl[69] br[69] wl[10] vdd gnd cell_6t
Xbit_r11_c69 bl[69] br[69] wl[11] vdd gnd cell_6t
Xbit_r12_c69 bl[69] br[69] wl[12] vdd gnd cell_6t
Xbit_r13_c69 bl[69] br[69] wl[13] vdd gnd cell_6t
Xbit_r14_c69 bl[69] br[69] wl[14] vdd gnd cell_6t
Xbit_r15_c69 bl[69] br[69] wl[15] vdd gnd cell_6t
Xbit_r16_c69 bl[69] br[69] wl[16] vdd gnd cell_6t
Xbit_r17_c69 bl[69] br[69] wl[17] vdd gnd cell_6t
Xbit_r18_c69 bl[69] br[69] wl[18] vdd gnd cell_6t
Xbit_r19_c69 bl[69] br[69] wl[19] vdd gnd cell_6t
Xbit_r20_c69 bl[69] br[69] wl[20] vdd gnd cell_6t
Xbit_r21_c69 bl[69] br[69] wl[21] vdd gnd cell_6t
Xbit_r22_c69 bl[69] br[69] wl[22] vdd gnd cell_6t
Xbit_r23_c69 bl[69] br[69] wl[23] vdd gnd cell_6t
Xbit_r24_c69 bl[69] br[69] wl[24] vdd gnd cell_6t
Xbit_r25_c69 bl[69] br[69] wl[25] vdd gnd cell_6t
Xbit_r26_c69 bl[69] br[69] wl[26] vdd gnd cell_6t
Xbit_r27_c69 bl[69] br[69] wl[27] vdd gnd cell_6t
Xbit_r28_c69 bl[69] br[69] wl[28] vdd gnd cell_6t
Xbit_r29_c69 bl[69] br[69] wl[29] vdd gnd cell_6t
Xbit_r30_c69 bl[69] br[69] wl[30] vdd gnd cell_6t
Xbit_r31_c69 bl[69] br[69] wl[31] vdd gnd cell_6t
Xbit_r32_c69 bl[69] br[69] wl[32] vdd gnd cell_6t
Xbit_r33_c69 bl[69] br[69] wl[33] vdd gnd cell_6t
Xbit_r34_c69 bl[69] br[69] wl[34] vdd gnd cell_6t
Xbit_r35_c69 bl[69] br[69] wl[35] vdd gnd cell_6t
Xbit_r36_c69 bl[69] br[69] wl[36] vdd gnd cell_6t
Xbit_r37_c69 bl[69] br[69] wl[37] vdd gnd cell_6t
Xbit_r38_c69 bl[69] br[69] wl[38] vdd gnd cell_6t
Xbit_r39_c69 bl[69] br[69] wl[39] vdd gnd cell_6t
Xbit_r40_c69 bl[69] br[69] wl[40] vdd gnd cell_6t
Xbit_r41_c69 bl[69] br[69] wl[41] vdd gnd cell_6t
Xbit_r42_c69 bl[69] br[69] wl[42] vdd gnd cell_6t
Xbit_r43_c69 bl[69] br[69] wl[43] vdd gnd cell_6t
Xbit_r44_c69 bl[69] br[69] wl[44] vdd gnd cell_6t
Xbit_r45_c69 bl[69] br[69] wl[45] vdd gnd cell_6t
Xbit_r46_c69 bl[69] br[69] wl[46] vdd gnd cell_6t
Xbit_r47_c69 bl[69] br[69] wl[47] vdd gnd cell_6t
Xbit_r48_c69 bl[69] br[69] wl[48] vdd gnd cell_6t
Xbit_r49_c69 bl[69] br[69] wl[49] vdd gnd cell_6t
Xbit_r50_c69 bl[69] br[69] wl[50] vdd gnd cell_6t
Xbit_r51_c69 bl[69] br[69] wl[51] vdd gnd cell_6t
Xbit_r52_c69 bl[69] br[69] wl[52] vdd gnd cell_6t
Xbit_r53_c69 bl[69] br[69] wl[53] vdd gnd cell_6t
Xbit_r54_c69 bl[69] br[69] wl[54] vdd gnd cell_6t
Xbit_r55_c69 bl[69] br[69] wl[55] vdd gnd cell_6t
Xbit_r56_c69 bl[69] br[69] wl[56] vdd gnd cell_6t
Xbit_r57_c69 bl[69] br[69] wl[57] vdd gnd cell_6t
Xbit_r58_c69 bl[69] br[69] wl[58] vdd gnd cell_6t
Xbit_r59_c69 bl[69] br[69] wl[59] vdd gnd cell_6t
Xbit_r60_c69 bl[69] br[69] wl[60] vdd gnd cell_6t
Xbit_r61_c69 bl[69] br[69] wl[61] vdd gnd cell_6t
Xbit_r62_c69 bl[69] br[69] wl[62] vdd gnd cell_6t
Xbit_r63_c69 bl[69] br[69] wl[63] vdd gnd cell_6t
Xbit_r64_c69 bl[69] br[69] wl[64] vdd gnd cell_6t
Xbit_r65_c69 bl[69] br[69] wl[65] vdd gnd cell_6t
Xbit_r66_c69 bl[69] br[69] wl[66] vdd gnd cell_6t
Xbit_r67_c69 bl[69] br[69] wl[67] vdd gnd cell_6t
Xbit_r68_c69 bl[69] br[69] wl[68] vdd gnd cell_6t
Xbit_r69_c69 bl[69] br[69] wl[69] vdd gnd cell_6t
Xbit_r70_c69 bl[69] br[69] wl[70] vdd gnd cell_6t
Xbit_r71_c69 bl[69] br[69] wl[71] vdd gnd cell_6t
Xbit_r72_c69 bl[69] br[69] wl[72] vdd gnd cell_6t
Xbit_r73_c69 bl[69] br[69] wl[73] vdd gnd cell_6t
Xbit_r74_c69 bl[69] br[69] wl[74] vdd gnd cell_6t
Xbit_r75_c69 bl[69] br[69] wl[75] vdd gnd cell_6t
Xbit_r76_c69 bl[69] br[69] wl[76] vdd gnd cell_6t
Xbit_r77_c69 bl[69] br[69] wl[77] vdd gnd cell_6t
Xbit_r78_c69 bl[69] br[69] wl[78] vdd gnd cell_6t
Xbit_r79_c69 bl[69] br[69] wl[79] vdd gnd cell_6t
Xbit_r80_c69 bl[69] br[69] wl[80] vdd gnd cell_6t
Xbit_r81_c69 bl[69] br[69] wl[81] vdd gnd cell_6t
Xbit_r82_c69 bl[69] br[69] wl[82] vdd gnd cell_6t
Xbit_r83_c69 bl[69] br[69] wl[83] vdd gnd cell_6t
Xbit_r84_c69 bl[69] br[69] wl[84] vdd gnd cell_6t
Xbit_r85_c69 bl[69] br[69] wl[85] vdd gnd cell_6t
Xbit_r86_c69 bl[69] br[69] wl[86] vdd gnd cell_6t
Xbit_r87_c69 bl[69] br[69] wl[87] vdd gnd cell_6t
Xbit_r88_c69 bl[69] br[69] wl[88] vdd gnd cell_6t
Xbit_r89_c69 bl[69] br[69] wl[89] vdd gnd cell_6t
Xbit_r90_c69 bl[69] br[69] wl[90] vdd gnd cell_6t
Xbit_r91_c69 bl[69] br[69] wl[91] vdd gnd cell_6t
Xbit_r92_c69 bl[69] br[69] wl[92] vdd gnd cell_6t
Xbit_r93_c69 bl[69] br[69] wl[93] vdd gnd cell_6t
Xbit_r94_c69 bl[69] br[69] wl[94] vdd gnd cell_6t
Xbit_r95_c69 bl[69] br[69] wl[95] vdd gnd cell_6t
Xbit_r96_c69 bl[69] br[69] wl[96] vdd gnd cell_6t
Xbit_r97_c69 bl[69] br[69] wl[97] vdd gnd cell_6t
Xbit_r98_c69 bl[69] br[69] wl[98] vdd gnd cell_6t
Xbit_r99_c69 bl[69] br[69] wl[99] vdd gnd cell_6t
Xbit_r100_c69 bl[69] br[69] wl[100] vdd gnd cell_6t
Xbit_r101_c69 bl[69] br[69] wl[101] vdd gnd cell_6t
Xbit_r102_c69 bl[69] br[69] wl[102] vdd gnd cell_6t
Xbit_r103_c69 bl[69] br[69] wl[103] vdd gnd cell_6t
Xbit_r104_c69 bl[69] br[69] wl[104] vdd gnd cell_6t
Xbit_r105_c69 bl[69] br[69] wl[105] vdd gnd cell_6t
Xbit_r106_c69 bl[69] br[69] wl[106] vdd gnd cell_6t
Xbit_r107_c69 bl[69] br[69] wl[107] vdd gnd cell_6t
Xbit_r108_c69 bl[69] br[69] wl[108] vdd gnd cell_6t
Xbit_r109_c69 bl[69] br[69] wl[109] vdd gnd cell_6t
Xbit_r110_c69 bl[69] br[69] wl[110] vdd gnd cell_6t
Xbit_r111_c69 bl[69] br[69] wl[111] vdd gnd cell_6t
Xbit_r112_c69 bl[69] br[69] wl[112] vdd gnd cell_6t
Xbit_r113_c69 bl[69] br[69] wl[113] vdd gnd cell_6t
Xbit_r114_c69 bl[69] br[69] wl[114] vdd gnd cell_6t
Xbit_r115_c69 bl[69] br[69] wl[115] vdd gnd cell_6t
Xbit_r116_c69 bl[69] br[69] wl[116] vdd gnd cell_6t
Xbit_r117_c69 bl[69] br[69] wl[117] vdd gnd cell_6t
Xbit_r118_c69 bl[69] br[69] wl[118] vdd gnd cell_6t
Xbit_r119_c69 bl[69] br[69] wl[119] vdd gnd cell_6t
Xbit_r120_c69 bl[69] br[69] wl[120] vdd gnd cell_6t
Xbit_r121_c69 bl[69] br[69] wl[121] vdd gnd cell_6t
Xbit_r122_c69 bl[69] br[69] wl[122] vdd gnd cell_6t
Xbit_r123_c69 bl[69] br[69] wl[123] vdd gnd cell_6t
Xbit_r124_c69 bl[69] br[69] wl[124] vdd gnd cell_6t
Xbit_r125_c69 bl[69] br[69] wl[125] vdd gnd cell_6t
Xbit_r126_c69 bl[69] br[69] wl[126] vdd gnd cell_6t
Xbit_r127_c69 bl[69] br[69] wl[127] vdd gnd cell_6t
Xbit_r0_c70 bl[70] br[70] wl[0] vdd gnd cell_6t
Xbit_r1_c70 bl[70] br[70] wl[1] vdd gnd cell_6t
Xbit_r2_c70 bl[70] br[70] wl[2] vdd gnd cell_6t
Xbit_r3_c70 bl[70] br[70] wl[3] vdd gnd cell_6t
Xbit_r4_c70 bl[70] br[70] wl[4] vdd gnd cell_6t
Xbit_r5_c70 bl[70] br[70] wl[5] vdd gnd cell_6t
Xbit_r6_c70 bl[70] br[70] wl[6] vdd gnd cell_6t
Xbit_r7_c70 bl[70] br[70] wl[7] vdd gnd cell_6t
Xbit_r8_c70 bl[70] br[70] wl[8] vdd gnd cell_6t
Xbit_r9_c70 bl[70] br[70] wl[9] vdd gnd cell_6t
Xbit_r10_c70 bl[70] br[70] wl[10] vdd gnd cell_6t
Xbit_r11_c70 bl[70] br[70] wl[11] vdd gnd cell_6t
Xbit_r12_c70 bl[70] br[70] wl[12] vdd gnd cell_6t
Xbit_r13_c70 bl[70] br[70] wl[13] vdd gnd cell_6t
Xbit_r14_c70 bl[70] br[70] wl[14] vdd gnd cell_6t
Xbit_r15_c70 bl[70] br[70] wl[15] vdd gnd cell_6t
Xbit_r16_c70 bl[70] br[70] wl[16] vdd gnd cell_6t
Xbit_r17_c70 bl[70] br[70] wl[17] vdd gnd cell_6t
Xbit_r18_c70 bl[70] br[70] wl[18] vdd gnd cell_6t
Xbit_r19_c70 bl[70] br[70] wl[19] vdd gnd cell_6t
Xbit_r20_c70 bl[70] br[70] wl[20] vdd gnd cell_6t
Xbit_r21_c70 bl[70] br[70] wl[21] vdd gnd cell_6t
Xbit_r22_c70 bl[70] br[70] wl[22] vdd gnd cell_6t
Xbit_r23_c70 bl[70] br[70] wl[23] vdd gnd cell_6t
Xbit_r24_c70 bl[70] br[70] wl[24] vdd gnd cell_6t
Xbit_r25_c70 bl[70] br[70] wl[25] vdd gnd cell_6t
Xbit_r26_c70 bl[70] br[70] wl[26] vdd gnd cell_6t
Xbit_r27_c70 bl[70] br[70] wl[27] vdd gnd cell_6t
Xbit_r28_c70 bl[70] br[70] wl[28] vdd gnd cell_6t
Xbit_r29_c70 bl[70] br[70] wl[29] vdd gnd cell_6t
Xbit_r30_c70 bl[70] br[70] wl[30] vdd gnd cell_6t
Xbit_r31_c70 bl[70] br[70] wl[31] vdd gnd cell_6t
Xbit_r32_c70 bl[70] br[70] wl[32] vdd gnd cell_6t
Xbit_r33_c70 bl[70] br[70] wl[33] vdd gnd cell_6t
Xbit_r34_c70 bl[70] br[70] wl[34] vdd gnd cell_6t
Xbit_r35_c70 bl[70] br[70] wl[35] vdd gnd cell_6t
Xbit_r36_c70 bl[70] br[70] wl[36] vdd gnd cell_6t
Xbit_r37_c70 bl[70] br[70] wl[37] vdd gnd cell_6t
Xbit_r38_c70 bl[70] br[70] wl[38] vdd gnd cell_6t
Xbit_r39_c70 bl[70] br[70] wl[39] vdd gnd cell_6t
Xbit_r40_c70 bl[70] br[70] wl[40] vdd gnd cell_6t
Xbit_r41_c70 bl[70] br[70] wl[41] vdd gnd cell_6t
Xbit_r42_c70 bl[70] br[70] wl[42] vdd gnd cell_6t
Xbit_r43_c70 bl[70] br[70] wl[43] vdd gnd cell_6t
Xbit_r44_c70 bl[70] br[70] wl[44] vdd gnd cell_6t
Xbit_r45_c70 bl[70] br[70] wl[45] vdd gnd cell_6t
Xbit_r46_c70 bl[70] br[70] wl[46] vdd gnd cell_6t
Xbit_r47_c70 bl[70] br[70] wl[47] vdd gnd cell_6t
Xbit_r48_c70 bl[70] br[70] wl[48] vdd gnd cell_6t
Xbit_r49_c70 bl[70] br[70] wl[49] vdd gnd cell_6t
Xbit_r50_c70 bl[70] br[70] wl[50] vdd gnd cell_6t
Xbit_r51_c70 bl[70] br[70] wl[51] vdd gnd cell_6t
Xbit_r52_c70 bl[70] br[70] wl[52] vdd gnd cell_6t
Xbit_r53_c70 bl[70] br[70] wl[53] vdd gnd cell_6t
Xbit_r54_c70 bl[70] br[70] wl[54] vdd gnd cell_6t
Xbit_r55_c70 bl[70] br[70] wl[55] vdd gnd cell_6t
Xbit_r56_c70 bl[70] br[70] wl[56] vdd gnd cell_6t
Xbit_r57_c70 bl[70] br[70] wl[57] vdd gnd cell_6t
Xbit_r58_c70 bl[70] br[70] wl[58] vdd gnd cell_6t
Xbit_r59_c70 bl[70] br[70] wl[59] vdd gnd cell_6t
Xbit_r60_c70 bl[70] br[70] wl[60] vdd gnd cell_6t
Xbit_r61_c70 bl[70] br[70] wl[61] vdd gnd cell_6t
Xbit_r62_c70 bl[70] br[70] wl[62] vdd gnd cell_6t
Xbit_r63_c70 bl[70] br[70] wl[63] vdd gnd cell_6t
Xbit_r64_c70 bl[70] br[70] wl[64] vdd gnd cell_6t
Xbit_r65_c70 bl[70] br[70] wl[65] vdd gnd cell_6t
Xbit_r66_c70 bl[70] br[70] wl[66] vdd gnd cell_6t
Xbit_r67_c70 bl[70] br[70] wl[67] vdd gnd cell_6t
Xbit_r68_c70 bl[70] br[70] wl[68] vdd gnd cell_6t
Xbit_r69_c70 bl[70] br[70] wl[69] vdd gnd cell_6t
Xbit_r70_c70 bl[70] br[70] wl[70] vdd gnd cell_6t
Xbit_r71_c70 bl[70] br[70] wl[71] vdd gnd cell_6t
Xbit_r72_c70 bl[70] br[70] wl[72] vdd gnd cell_6t
Xbit_r73_c70 bl[70] br[70] wl[73] vdd gnd cell_6t
Xbit_r74_c70 bl[70] br[70] wl[74] vdd gnd cell_6t
Xbit_r75_c70 bl[70] br[70] wl[75] vdd gnd cell_6t
Xbit_r76_c70 bl[70] br[70] wl[76] vdd gnd cell_6t
Xbit_r77_c70 bl[70] br[70] wl[77] vdd gnd cell_6t
Xbit_r78_c70 bl[70] br[70] wl[78] vdd gnd cell_6t
Xbit_r79_c70 bl[70] br[70] wl[79] vdd gnd cell_6t
Xbit_r80_c70 bl[70] br[70] wl[80] vdd gnd cell_6t
Xbit_r81_c70 bl[70] br[70] wl[81] vdd gnd cell_6t
Xbit_r82_c70 bl[70] br[70] wl[82] vdd gnd cell_6t
Xbit_r83_c70 bl[70] br[70] wl[83] vdd gnd cell_6t
Xbit_r84_c70 bl[70] br[70] wl[84] vdd gnd cell_6t
Xbit_r85_c70 bl[70] br[70] wl[85] vdd gnd cell_6t
Xbit_r86_c70 bl[70] br[70] wl[86] vdd gnd cell_6t
Xbit_r87_c70 bl[70] br[70] wl[87] vdd gnd cell_6t
Xbit_r88_c70 bl[70] br[70] wl[88] vdd gnd cell_6t
Xbit_r89_c70 bl[70] br[70] wl[89] vdd gnd cell_6t
Xbit_r90_c70 bl[70] br[70] wl[90] vdd gnd cell_6t
Xbit_r91_c70 bl[70] br[70] wl[91] vdd gnd cell_6t
Xbit_r92_c70 bl[70] br[70] wl[92] vdd gnd cell_6t
Xbit_r93_c70 bl[70] br[70] wl[93] vdd gnd cell_6t
Xbit_r94_c70 bl[70] br[70] wl[94] vdd gnd cell_6t
Xbit_r95_c70 bl[70] br[70] wl[95] vdd gnd cell_6t
Xbit_r96_c70 bl[70] br[70] wl[96] vdd gnd cell_6t
Xbit_r97_c70 bl[70] br[70] wl[97] vdd gnd cell_6t
Xbit_r98_c70 bl[70] br[70] wl[98] vdd gnd cell_6t
Xbit_r99_c70 bl[70] br[70] wl[99] vdd gnd cell_6t
Xbit_r100_c70 bl[70] br[70] wl[100] vdd gnd cell_6t
Xbit_r101_c70 bl[70] br[70] wl[101] vdd gnd cell_6t
Xbit_r102_c70 bl[70] br[70] wl[102] vdd gnd cell_6t
Xbit_r103_c70 bl[70] br[70] wl[103] vdd gnd cell_6t
Xbit_r104_c70 bl[70] br[70] wl[104] vdd gnd cell_6t
Xbit_r105_c70 bl[70] br[70] wl[105] vdd gnd cell_6t
Xbit_r106_c70 bl[70] br[70] wl[106] vdd gnd cell_6t
Xbit_r107_c70 bl[70] br[70] wl[107] vdd gnd cell_6t
Xbit_r108_c70 bl[70] br[70] wl[108] vdd gnd cell_6t
Xbit_r109_c70 bl[70] br[70] wl[109] vdd gnd cell_6t
Xbit_r110_c70 bl[70] br[70] wl[110] vdd gnd cell_6t
Xbit_r111_c70 bl[70] br[70] wl[111] vdd gnd cell_6t
Xbit_r112_c70 bl[70] br[70] wl[112] vdd gnd cell_6t
Xbit_r113_c70 bl[70] br[70] wl[113] vdd gnd cell_6t
Xbit_r114_c70 bl[70] br[70] wl[114] vdd gnd cell_6t
Xbit_r115_c70 bl[70] br[70] wl[115] vdd gnd cell_6t
Xbit_r116_c70 bl[70] br[70] wl[116] vdd gnd cell_6t
Xbit_r117_c70 bl[70] br[70] wl[117] vdd gnd cell_6t
Xbit_r118_c70 bl[70] br[70] wl[118] vdd gnd cell_6t
Xbit_r119_c70 bl[70] br[70] wl[119] vdd gnd cell_6t
Xbit_r120_c70 bl[70] br[70] wl[120] vdd gnd cell_6t
Xbit_r121_c70 bl[70] br[70] wl[121] vdd gnd cell_6t
Xbit_r122_c70 bl[70] br[70] wl[122] vdd gnd cell_6t
Xbit_r123_c70 bl[70] br[70] wl[123] vdd gnd cell_6t
Xbit_r124_c70 bl[70] br[70] wl[124] vdd gnd cell_6t
Xbit_r125_c70 bl[70] br[70] wl[125] vdd gnd cell_6t
Xbit_r126_c70 bl[70] br[70] wl[126] vdd gnd cell_6t
Xbit_r127_c70 bl[70] br[70] wl[127] vdd gnd cell_6t
Xbit_r0_c71 bl[71] br[71] wl[0] vdd gnd cell_6t
Xbit_r1_c71 bl[71] br[71] wl[1] vdd gnd cell_6t
Xbit_r2_c71 bl[71] br[71] wl[2] vdd gnd cell_6t
Xbit_r3_c71 bl[71] br[71] wl[3] vdd gnd cell_6t
Xbit_r4_c71 bl[71] br[71] wl[4] vdd gnd cell_6t
Xbit_r5_c71 bl[71] br[71] wl[5] vdd gnd cell_6t
Xbit_r6_c71 bl[71] br[71] wl[6] vdd gnd cell_6t
Xbit_r7_c71 bl[71] br[71] wl[7] vdd gnd cell_6t
Xbit_r8_c71 bl[71] br[71] wl[8] vdd gnd cell_6t
Xbit_r9_c71 bl[71] br[71] wl[9] vdd gnd cell_6t
Xbit_r10_c71 bl[71] br[71] wl[10] vdd gnd cell_6t
Xbit_r11_c71 bl[71] br[71] wl[11] vdd gnd cell_6t
Xbit_r12_c71 bl[71] br[71] wl[12] vdd gnd cell_6t
Xbit_r13_c71 bl[71] br[71] wl[13] vdd gnd cell_6t
Xbit_r14_c71 bl[71] br[71] wl[14] vdd gnd cell_6t
Xbit_r15_c71 bl[71] br[71] wl[15] vdd gnd cell_6t
Xbit_r16_c71 bl[71] br[71] wl[16] vdd gnd cell_6t
Xbit_r17_c71 bl[71] br[71] wl[17] vdd gnd cell_6t
Xbit_r18_c71 bl[71] br[71] wl[18] vdd gnd cell_6t
Xbit_r19_c71 bl[71] br[71] wl[19] vdd gnd cell_6t
Xbit_r20_c71 bl[71] br[71] wl[20] vdd gnd cell_6t
Xbit_r21_c71 bl[71] br[71] wl[21] vdd gnd cell_6t
Xbit_r22_c71 bl[71] br[71] wl[22] vdd gnd cell_6t
Xbit_r23_c71 bl[71] br[71] wl[23] vdd gnd cell_6t
Xbit_r24_c71 bl[71] br[71] wl[24] vdd gnd cell_6t
Xbit_r25_c71 bl[71] br[71] wl[25] vdd gnd cell_6t
Xbit_r26_c71 bl[71] br[71] wl[26] vdd gnd cell_6t
Xbit_r27_c71 bl[71] br[71] wl[27] vdd gnd cell_6t
Xbit_r28_c71 bl[71] br[71] wl[28] vdd gnd cell_6t
Xbit_r29_c71 bl[71] br[71] wl[29] vdd gnd cell_6t
Xbit_r30_c71 bl[71] br[71] wl[30] vdd gnd cell_6t
Xbit_r31_c71 bl[71] br[71] wl[31] vdd gnd cell_6t
Xbit_r32_c71 bl[71] br[71] wl[32] vdd gnd cell_6t
Xbit_r33_c71 bl[71] br[71] wl[33] vdd gnd cell_6t
Xbit_r34_c71 bl[71] br[71] wl[34] vdd gnd cell_6t
Xbit_r35_c71 bl[71] br[71] wl[35] vdd gnd cell_6t
Xbit_r36_c71 bl[71] br[71] wl[36] vdd gnd cell_6t
Xbit_r37_c71 bl[71] br[71] wl[37] vdd gnd cell_6t
Xbit_r38_c71 bl[71] br[71] wl[38] vdd gnd cell_6t
Xbit_r39_c71 bl[71] br[71] wl[39] vdd gnd cell_6t
Xbit_r40_c71 bl[71] br[71] wl[40] vdd gnd cell_6t
Xbit_r41_c71 bl[71] br[71] wl[41] vdd gnd cell_6t
Xbit_r42_c71 bl[71] br[71] wl[42] vdd gnd cell_6t
Xbit_r43_c71 bl[71] br[71] wl[43] vdd gnd cell_6t
Xbit_r44_c71 bl[71] br[71] wl[44] vdd gnd cell_6t
Xbit_r45_c71 bl[71] br[71] wl[45] vdd gnd cell_6t
Xbit_r46_c71 bl[71] br[71] wl[46] vdd gnd cell_6t
Xbit_r47_c71 bl[71] br[71] wl[47] vdd gnd cell_6t
Xbit_r48_c71 bl[71] br[71] wl[48] vdd gnd cell_6t
Xbit_r49_c71 bl[71] br[71] wl[49] vdd gnd cell_6t
Xbit_r50_c71 bl[71] br[71] wl[50] vdd gnd cell_6t
Xbit_r51_c71 bl[71] br[71] wl[51] vdd gnd cell_6t
Xbit_r52_c71 bl[71] br[71] wl[52] vdd gnd cell_6t
Xbit_r53_c71 bl[71] br[71] wl[53] vdd gnd cell_6t
Xbit_r54_c71 bl[71] br[71] wl[54] vdd gnd cell_6t
Xbit_r55_c71 bl[71] br[71] wl[55] vdd gnd cell_6t
Xbit_r56_c71 bl[71] br[71] wl[56] vdd gnd cell_6t
Xbit_r57_c71 bl[71] br[71] wl[57] vdd gnd cell_6t
Xbit_r58_c71 bl[71] br[71] wl[58] vdd gnd cell_6t
Xbit_r59_c71 bl[71] br[71] wl[59] vdd gnd cell_6t
Xbit_r60_c71 bl[71] br[71] wl[60] vdd gnd cell_6t
Xbit_r61_c71 bl[71] br[71] wl[61] vdd gnd cell_6t
Xbit_r62_c71 bl[71] br[71] wl[62] vdd gnd cell_6t
Xbit_r63_c71 bl[71] br[71] wl[63] vdd gnd cell_6t
Xbit_r64_c71 bl[71] br[71] wl[64] vdd gnd cell_6t
Xbit_r65_c71 bl[71] br[71] wl[65] vdd gnd cell_6t
Xbit_r66_c71 bl[71] br[71] wl[66] vdd gnd cell_6t
Xbit_r67_c71 bl[71] br[71] wl[67] vdd gnd cell_6t
Xbit_r68_c71 bl[71] br[71] wl[68] vdd gnd cell_6t
Xbit_r69_c71 bl[71] br[71] wl[69] vdd gnd cell_6t
Xbit_r70_c71 bl[71] br[71] wl[70] vdd gnd cell_6t
Xbit_r71_c71 bl[71] br[71] wl[71] vdd gnd cell_6t
Xbit_r72_c71 bl[71] br[71] wl[72] vdd gnd cell_6t
Xbit_r73_c71 bl[71] br[71] wl[73] vdd gnd cell_6t
Xbit_r74_c71 bl[71] br[71] wl[74] vdd gnd cell_6t
Xbit_r75_c71 bl[71] br[71] wl[75] vdd gnd cell_6t
Xbit_r76_c71 bl[71] br[71] wl[76] vdd gnd cell_6t
Xbit_r77_c71 bl[71] br[71] wl[77] vdd gnd cell_6t
Xbit_r78_c71 bl[71] br[71] wl[78] vdd gnd cell_6t
Xbit_r79_c71 bl[71] br[71] wl[79] vdd gnd cell_6t
Xbit_r80_c71 bl[71] br[71] wl[80] vdd gnd cell_6t
Xbit_r81_c71 bl[71] br[71] wl[81] vdd gnd cell_6t
Xbit_r82_c71 bl[71] br[71] wl[82] vdd gnd cell_6t
Xbit_r83_c71 bl[71] br[71] wl[83] vdd gnd cell_6t
Xbit_r84_c71 bl[71] br[71] wl[84] vdd gnd cell_6t
Xbit_r85_c71 bl[71] br[71] wl[85] vdd gnd cell_6t
Xbit_r86_c71 bl[71] br[71] wl[86] vdd gnd cell_6t
Xbit_r87_c71 bl[71] br[71] wl[87] vdd gnd cell_6t
Xbit_r88_c71 bl[71] br[71] wl[88] vdd gnd cell_6t
Xbit_r89_c71 bl[71] br[71] wl[89] vdd gnd cell_6t
Xbit_r90_c71 bl[71] br[71] wl[90] vdd gnd cell_6t
Xbit_r91_c71 bl[71] br[71] wl[91] vdd gnd cell_6t
Xbit_r92_c71 bl[71] br[71] wl[92] vdd gnd cell_6t
Xbit_r93_c71 bl[71] br[71] wl[93] vdd gnd cell_6t
Xbit_r94_c71 bl[71] br[71] wl[94] vdd gnd cell_6t
Xbit_r95_c71 bl[71] br[71] wl[95] vdd gnd cell_6t
Xbit_r96_c71 bl[71] br[71] wl[96] vdd gnd cell_6t
Xbit_r97_c71 bl[71] br[71] wl[97] vdd gnd cell_6t
Xbit_r98_c71 bl[71] br[71] wl[98] vdd gnd cell_6t
Xbit_r99_c71 bl[71] br[71] wl[99] vdd gnd cell_6t
Xbit_r100_c71 bl[71] br[71] wl[100] vdd gnd cell_6t
Xbit_r101_c71 bl[71] br[71] wl[101] vdd gnd cell_6t
Xbit_r102_c71 bl[71] br[71] wl[102] vdd gnd cell_6t
Xbit_r103_c71 bl[71] br[71] wl[103] vdd gnd cell_6t
Xbit_r104_c71 bl[71] br[71] wl[104] vdd gnd cell_6t
Xbit_r105_c71 bl[71] br[71] wl[105] vdd gnd cell_6t
Xbit_r106_c71 bl[71] br[71] wl[106] vdd gnd cell_6t
Xbit_r107_c71 bl[71] br[71] wl[107] vdd gnd cell_6t
Xbit_r108_c71 bl[71] br[71] wl[108] vdd gnd cell_6t
Xbit_r109_c71 bl[71] br[71] wl[109] vdd gnd cell_6t
Xbit_r110_c71 bl[71] br[71] wl[110] vdd gnd cell_6t
Xbit_r111_c71 bl[71] br[71] wl[111] vdd gnd cell_6t
Xbit_r112_c71 bl[71] br[71] wl[112] vdd gnd cell_6t
Xbit_r113_c71 bl[71] br[71] wl[113] vdd gnd cell_6t
Xbit_r114_c71 bl[71] br[71] wl[114] vdd gnd cell_6t
Xbit_r115_c71 bl[71] br[71] wl[115] vdd gnd cell_6t
Xbit_r116_c71 bl[71] br[71] wl[116] vdd gnd cell_6t
Xbit_r117_c71 bl[71] br[71] wl[117] vdd gnd cell_6t
Xbit_r118_c71 bl[71] br[71] wl[118] vdd gnd cell_6t
Xbit_r119_c71 bl[71] br[71] wl[119] vdd gnd cell_6t
Xbit_r120_c71 bl[71] br[71] wl[120] vdd gnd cell_6t
Xbit_r121_c71 bl[71] br[71] wl[121] vdd gnd cell_6t
Xbit_r122_c71 bl[71] br[71] wl[122] vdd gnd cell_6t
Xbit_r123_c71 bl[71] br[71] wl[123] vdd gnd cell_6t
Xbit_r124_c71 bl[71] br[71] wl[124] vdd gnd cell_6t
Xbit_r125_c71 bl[71] br[71] wl[125] vdd gnd cell_6t
Xbit_r126_c71 bl[71] br[71] wl[126] vdd gnd cell_6t
Xbit_r127_c71 bl[71] br[71] wl[127] vdd gnd cell_6t
Xbit_r0_c72 bl[72] br[72] wl[0] vdd gnd cell_6t
Xbit_r1_c72 bl[72] br[72] wl[1] vdd gnd cell_6t
Xbit_r2_c72 bl[72] br[72] wl[2] vdd gnd cell_6t
Xbit_r3_c72 bl[72] br[72] wl[3] vdd gnd cell_6t
Xbit_r4_c72 bl[72] br[72] wl[4] vdd gnd cell_6t
Xbit_r5_c72 bl[72] br[72] wl[5] vdd gnd cell_6t
Xbit_r6_c72 bl[72] br[72] wl[6] vdd gnd cell_6t
Xbit_r7_c72 bl[72] br[72] wl[7] vdd gnd cell_6t
Xbit_r8_c72 bl[72] br[72] wl[8] vdd gnd cell_6t
Xbit_r9_c72 bl[72] br[72] wl[9] vdd gnd cell_6t
Xbit_r10_c72 bl[72] br[72] wl[10] vdd gnd cell_6t
Xbit_r11_c72 bl[72] br[72] wl[11] vdd gnd cell_6t
Xbit_r12_c72 bl[72] br[72] wl[12] vdd gnd cell_6t
Xbit_r13_c72 bl[72] br[72] wl[13] vdd gnd cell_6t
Xbit_r14_c72 bl[72] br[72] wl[14] vdd gnd cell_6t
Xbit_r15_c72 bl[72] br[72] wl[15] vdd gnd cell_6t
Xbit_r16_c72 bl[72] br[72] wl[16] vdd gnd cell_6t
Xbit_r17_c72 bl[72] br[72] wl[17] vdd gnd cell_6t
Xbit_r18_c72 bl[72] br[72] wl[18] vdd gnd cell_6t
Xbit_r19_c72 bl[72] br[72] wl[19] vdd gnd cell_6t
Xbit_r20_c72 bl[72] br[72] wl[20] vdd gnd cell_6t
Xbit_r21_c72 bl[72] br[72] wl[21] vdd gnd cell_6t
Xbit_r22_c72 bl[72] br[72] wl[22] vdd gnd cell_6t
Xbit_r23_c72 bl[72] br[72] wl[23] vdd gnd cell_6t
Xbit_r24_c72 bl[72] br[72] wl[24] vdd gnd cell_6t
Xbit_r25_c72 bl[72] br[72] wl[25] vdd gnd cell_6t
Xbit_r26_c72 bl[72] br[72] wl[26] vdd gnd cell_6t
Xbit_r27_c72 bl[72] br[72] wl[27] vdd gnd cell_6t
Xbit_r28_c72 bl[72] br[72] wl[28] vdd gnd cell_6t
Xbit_r29_c72 bl[72] br[72] wl[29] vdd gnd cell_6t
Xbit_r30_c72 bl[72] br[72] wl[30] vdd gnd cell_6t
Xbit_r31_c72 bl[72] br[72] wl[31] vdd gnd cell_6t
Xbit_r32_c72 bl[72] br[72] wl[32] vdd gnd cell_6t
Xbit_r33_c72 bl[72] br[72] wl[33] vdd gnd cell_6t
Xbit_r34_c72 bl[72] br[72] wl[34] vdd gnd cell_6t
Xbit_r35_c72 bl[72] br[72] wl[35] vdd gnd cell_6t
Xbit_r36_c72 bl[72] br[72] wl[36] vdd gnd cell_6t
Xbit_r37_c72 bl[72] br[72] wl[37] vdd gnd cell_6t
Xbit_r38_c72 bl[72] br[72] wl[38] vdd gnd cell_6t
Xbit_r39_c72 bl[72] br[72] wl[39] vdd gnd cell_6t
Xbit_r40_c72 bl[72] br[72] wl[40] vdd gnd cell_6t
Xbit_r41_c72 bl[72] br[72] wl[41] vdd gnd cell_6t
Xbit_r42_c72 bl[72] br[72] wl[42] vdd gnd cell_6t
Xbit_r43_c72 bl[72] br[72] wl[43] vdd gnd cell_6t
Xbit_r44_c72 bl[72] br[72] wl[44] vdd gnd cell_6t
Xbit_r45_c72 bl[72] br[72] wl[45] vdd gnd cell_6t
Xbit_r46_c72 bl[72] br[72] wl[46] vdd gnd cell_6t
Xbit_r47_c72 bl[72] br[72] wl[47] vdd gnd cell_6t
Xbit_r48_c72 bl[72] br[72] wl[48] vdd gnd cell_6t
Xbit_r49_c72 bl[72] br[72] wl[49] vdd gnd cell_6t
Xbit_r50_c72 bl[72] br[72] wl[50] vdd gnd cell_6t
Xbit_r51_c72 bl[72] br[72] wl[51] vdd gnd cell_6t
Xbit_r52_c72 bl[72] br[72] wl[52] vdd gnd cell_6t
Xbit_r53_c72 bl[72] br[72] wl[53] vdd gnd cell_6t
Xbit_r54_c72 bl[72] br[72] wl[54] vdd gnd cell_6t
Xbit_r55_c72 bl[72] br[72] wl[55] vdd gnd cell_6t
Xbit_r56_c72 bl[72] br[72] wl[56] vdd gnd cell_6t
Xbit_r57_c72 bl[72] br[72] wl[57] vdd gnd cell_6t
Xbit_r58_c72 bl[72] br[72] wl[58] vdd gnd cell_6t
Xbit_r59_c72 bl[72] br[72] wl[59] vdd gnd cell_6t
Xbit_r60_c72 bl[72] br[72] wl[60] vdd gnd cell_6t
Xbit_r61_c72 bl[72] br[72] wl[61] vdd gnd cell_6t
Xbit_r62_c72 bl[72] br[72] wl[62] vdd gnd cell_6t
Xbit_r63_c72 bl[72] br[72] wl[63] vdd gnd cell_6t
Xbit_r64_c72 bl[72] br[72] wl[64] vdd gnd cell_6t
Xbit_r65_c72 bl[72] br[72] wl[65] vdd gnd cell_6t
Xbit_r66_c72 bl[72] br[72] wl[66] vdd gnd cell_6t
Xbit_r67_c72 bl[72] br[72] wl[67] vdd gnd cell_6t
Xbit_r68_c72 bl[72] br[72] wl[68] vdd gnd cell_6t
Xbit_r69_c72 bl[72] br[72] wl[69] vdd gnd cell_6t
Xbit_r70_c72 bl[72] br[72] wl[70] vdd gnd cell_6t
Xbit_r71_c72 bl[72] br[72] wl[71] vdd gnd cell_6t
Xbit_r72_c72 bl[72] br[72] wl[72] vdd gnd cell_6t
Xbit_r73_c72 bl[72] br[72] wl[73] vdd gnd cell_6t
Xbit_r74_c72 bl[72] br[72] wl[74] vdd gnd cell_6t
Xbit_r75_c72 bl[72] br[72] wl[75] vdd gnd cell_6t
Xbit_r76_c72 bl[72] br[72] wl[76] vdd gnd cell_6t
Xbit_r77_c72 bl[72] br[72] wl[77] vdd gnd cell_6t
Xbit_r78_c72 bl[72] br[72] wl[78] vdd gnd cell_6t
Xbit_r79_c72 bl[72] br[72] wl[79] vdd gnd cell_6t
Xbit_r80_c72 bl[72] br[72] wl[80] vdd gnd cell_6t
Xbit_r81_c72 bl[72] br[72] wl[81] vdd gnd cell_6t
Xbit_r82_c72 bl[72] br[72] wl[82] vdd gnd cell_6t
Xbit_r83_c72 bl[72] br[72] wl[83] vdd gnd cell_6t
Xbit_r84_c72 bl[72] br[72] wl[84] vdd gnd cell_6t
Xbit_r85_c72 bl[72] br[72] wl[85] vdd gnd cell_6t
Xbit_r86_c72 bl[72] br[72] wl[86] vdd gnd cell_6t
Xbit_r87_c72 bl[72] br[72] wl[87] vdd gnd cell_6t
Xbit_r88_c72 bl[72] br[72] wl[88] vdd gnd cell_6t
Xbit_r89_c72 bl[72] br[72] wl[89] vdd gnd cell_6t
Xbit_r90_c72 bl[72] br[72] wl[90] vdd gnd cell_6t
Xbit_r91_c72 bl[72] br[72] wl[91] vdd gnd cell_6t
Xbit_r92_c72 bl[72] br[72] wl[92] vdd gnd cell_6t
Xbit_r93_c72 bl[72] br[72] wl[93] vdd gnd cell_6t
Xbit_r94_c72 bl[72] br[72] wl[94] vdd gnd cell_6t
Xbit_r95_c72 bl[72] br[72] wl[95] vdd gnd cell_6t
Xbit_r96_c72 bl[72] br[72] wl[96] vdd gnd cell_6t
Xbit_r97_c72 bl[72] br[72] wl[97] vdd gnd cell_6t
Xbit_r98_c72 bl[72] br[72] wl[98] vdd gnd cell_6t
Xbit_r99_c72 bl[72] br[72] wl[99] vdd gnd cell_6t
Xbit_r100_c72 bl[72] br[72] wl[100] vdd gnd cell_6t
Xbit_r101_c72 bl[72] br[72] wl[101] vdd gnd cell_6t
Xbit_r102_c72 bl[72] br[72] wl[102] vdd gnd cell_6t
Xbit_r103_c72 bl[72] br[72] wl[103] vdd gnd cell_6t
Xbit_r104_c72 bl[72] br[72] wl[104] vdd gnd cell_6t
Xbit_r105_c72 bl[72] br[72] wl[105] vdd gnd cell_6t
Xbit_r106_c72 bl[72] br[72] wl[106] vdd gnd cell_6t
Xbit_r107_c72 bl[72] br[72] wl[107] vdd gnd cell_6t
Xbit_r108_c72 bl[72] br[72] wl[108] vdd gnd cell_6t
Xbit_r109_c72 bl[72] br[72] wl[109] vdd gnd cell_6t
Xbit_r110_c72 bl[72] br[72] wl[110] vdd gnd cell_6t
Xbit_r111_c72 bl[72] br[72] wl[111] vdd gnd cell_6t
Xbit_r112_c72 bl[72] br[72] wl[112] vdd gnd cell_6t
Xbit_r113_c72 bl[72] br[72] wl[113] vdd gnd cell_6t
Xbit_r114_c72 bl[72] br[72] wl[114] vdd gnd cell_6t
Xbit_r115_c72 bl[72] br[72] wl[115] vdd gnd cell_6t
Xbit_r116_c72 bl[72] br[72] wl[116] vdd gnd cell_6t
Xbit_r117_c72 bl[72] br[72] wl[117] vdd gnd cell_6t
Xbit_r118_c72 bl[72] br[72] wl[118] vdd gnd cell_6t
Xbit_r119_c72 bl[72] br[72] wl[119] vdd gnd cell_6t
Xbit_r120_c72 bl[72] br[72] wl[120] vdd gnd cell_6t
Xbit_r121_c72 bl[72] br[72] wl[121] vdd gnd cell_6t
Xbit_r122_c72 bl[72] br[72] wl[122] vdd gnd cell_6t
Xbit_r123_c72 bl[72] br[72] wl[123] vdd gnd cell_6t
Xbit_r124_c72 bl[72] br[72] wl[124] vdd gnd cell_6t
Xbit_r125_c72 bl[72] br[72] wl[125] vdd gnd cell_6t
Xbit_r126_c72 bl[72] br[72] wl[126] vdd gnd cell_6t
Xbit_r127_c72 bl[72] br[72] wl[127] vdd gnd cell_6t
Xbit_r0_c73 bl[73] br[73] wl[0] vdd gnd cell_6t
Xbit_r1_c73 bl[73] br[73] wl[1] vdd gnd cell_6t
Xbit_r2_c73 bl[73] br[73] wl[2] vdd gnd cell_6t
Xbit_r3_c73 bl[73] br[73] wl[3] vdd gnd cell_6t
Xbit_r4_c73 bl[73] br[73] wl[4] vdd gnd cell_6t
Xbit_r5_c73 bl[73] br[73] wl[5] vdd gnd cell_6t
Xbit_r6_c73 bl[73] br[73] wl[6] vdd gnd cell_6t
Xbit_r7_c73 bl[73] br[73] wl[7] vdd gnd cell_6t
Xbit_r8_c73 bl[73] br[73] wl[8] vdd gnd cell_6t
Xbit_r9_c73 bl[73] br[73] wl[9] vdd gnd cell_6t
Xbit_r10_c73 bl[73] br[73] wl[10] vdd gnd cell_6t
Xbit_r11_c73 bl[73] br[73] wl[11] vdd gnd cell_6t
Xbit_r12_c73 bl[73] br[73] wl[12] vdd gnd cell_6t
Xbit_r13_c73 bl[73] br[73] wl[13] vdd gnd cell_6t
Xbit_r14_c73 bl[73] br[73] wl[14] vdd gnd cell_6t
Xbit_r15_c73 bl[73] br[73] wl[15] vdd gnd cell_6t
Xbit_r16_c73 bl[73] br[73] wl[16] vdd gnd cell_6t
Xbit_r17_c73 bl[73] br[73] wl[17] vdd gnd cell_6t
Xbit_r18_c73 bl[73] br[73] wl[18] vdd gnd cell_6t
Xbit_r19_c73 bl[73] br[73] wl[19] vdd gnd cell_6t
Xbit_r20_c73 bl[73] br[73] wl[20] vdd gnd cell_6t
Xbit_r21_c73 bl[73] br[73] wl[21] vdd gnd cell_6t
Xbit_r22_c73 bl[73] br[73] wl[22] vdd gnd cell_6t
Xbit_r23_c73 bl[73] br[73] wl[23] vdd gnd cell_6t
Xbit_r24_c73 bl[73] br[73] wl[24] vdd gnd cell_6t
Xbit_r25_c73 bl[73] br[73] wl[25] vdd gnd cell_6t
Xbit_r26_c73 bl[73] br[73] wl[26] vdd gnd cell_6t
Xbit_r27_c73 bl[73] br[73] wl[27] vdd gnd cell_6t
Xbit_r28_c73 bl[73] br[73] wl[28] vdd gnd cell_6t
Xbit_r29_c73 bl[73] br[73] wl[29] vdd gnd cell_6t
Xbit_r30_c73 bl[73] br[73] wl[30] vdd gnd cell_6t
Xbit_r31_c73 bl[73] br[73] wl[31] vdd gnd cell_6t
Xbit_r32_c73 bl[73] br[73] wl[32] vdd gnd cell_6t
Xbit_r33_c73 bl[73] br[73] wl[33] vdd gnd cell_6t
Xbit_r34_c73 bl[73] br[73] wl[34] vdd gnd cell_6t
Xbit_r35_c73 bl[73] br[73] wl[35] vdd gnd cell_6t
Xbit_r36_c73 bl[73] br[73] wl[36] vdd gnd cell_6t
Xbit_r37_c73 bl[73] br[73] wl[37] vdd gnd cell_6t
Xbit_r38_c73 bl[73] br[73] wl[38] vdd gnd cell_6t
Xbit_r39_c73 bl[73] br[73] wl[39] vdd gnd cell_6t
Xbit_r40_c73 bl[73] br[73] wl[40] vdd gnd cell_6t
Xbit_r41_c73 bl[73] br[73] wl[41] vdd gnd cell_6t
Xbit_r42_c73 bl[73] br[73] wl[42] vdd gnd cell_6t
Xbit_r43_c73 bl[73] br[73] wl[43] vdd gnd cell_6t
Xbit_r44_c73 bl[73] br[73] wl[44] vdd gnd cell_6t
Xbit_r45_c73 bl[73] br[73] wl[45] vdd gnd cell_6t
Xbit_r46_c73 bl[73] br[73] wl[46] vdd gnd cell_6t
Xbit_r47_c73 bl[73] br[73] wl[47] vdd gnd cell_6t
Xbit_r48_c73 bl[73] br[73] wl[48] vdd gnd cell_6t
Xbit_r49_c73 bl[73] br[73] wl[49] vdd gnd cell_6t
Xbit_r50_c73 bl[73] br[73] wl[50] vdd gnd cell_6t
Xbit_r51_c73 bl[73] br[73] wl[51] vdd gnd cell_6t
Xbit_r52_c73 bl[73] br[73] wl[52] vdd gnd cell_6t
Xbit_r53_c73 bl[73] br[73] wl[53] vdd gnd cell_6t
Xbit_r54_c73 bl[73] br[73] wl[54] vdd gnd cell_6t
Xbit_r55_c73 bl[73] br[73] wl[55] vdd gnd cell_6t
Xbit_r56_c73 bl[73] br[73] wl[56] vdd gnd cell_6t
Xbit_r57_c73 bl[73] br[73] wl[57] vdd gnd cell_6t
Xbit_r58_c73 bl[73] br[73] wl[58] vdd gnd cell_6t
Xbit_r59_c73 bl[73] br[73] wl[59] vdd gnd cell_6t
Xbit_r60_c73 bl[73] br[73] wl[60] vdd gnd cell_6t
Xbit_r61_c73 bl[73] br[73] wl[61] vdd gnd cell_6t
Xbit_r62_c73 bl[73] br[73] wl[62] vdd gnd cell_6t
Xbit_r63_c73 bl[73] br[73] wl[63] vdd gnd cell_6t
Xbit_r64_c73 bl[73] br[73] wl[64] vdd gnd cell_6t
Xbit_r65_c73 bl[73] br[73] wl[65] vdd gnd cell_6t
Xbit_r66_c73 bl[73] br[73] wl[66] vdd gnd cell_6t
Xbit_r67_c73 bl[73] br[73] wl[67] vdd gnd cell_6t
Xbit_r68_c73 bl[73] br[73] wl[68] vdd gnd cell_6t
Xbit_r69_c73 bl[73] br[73] wl[69] vdd gnd cell_6t
Xbit_r70_c73 bl[73] br[73] wl[70] vdd gnd cell_6t
Xbit_r71_c73 bl[73] br[73] wl[71] vdd gnd cell_6t
Xbit_r72_c73 bl[73] br[73] wl[72] vdd gnd cell_6t
Xbit_r73_c73 bl[73] br[73] wl[73] vdd gnd cell_6t
Xbit_r74_c73 bl[73] br[73] wl[74] vdd gnd cell_6t
Xbit_r75_c73 bl[73] br[73] wl[75] vdd gnd cell_6t
Xbit_r76_c73 bl[73] br[73] wl[76] vdd gnd cell_6t
Xbit_r77_c73 bl[73] br[73] wl[77] vdd gnd cell_6t
Xbit_r78_c73 bl[73] br[73] wl[78] vdd gnd cell_6t
Xbit_r79_c73 bl[73] br[73] wl[79] vdd gnd cell_6t
Xbit_r80_c73 bl[73] br[73] wl[80] vdd gnd cell_6t
Xbit_r81_c73 bl[73] br[73] wl[81] vdd gnd cell_6t
Xbit_r82_c73 bl[73] br[73] wl[82] vdd gnd cell_6t
Xbit_r83_c73 bl[73] br[73] wl[83] vdd gnd cell_6t
Xbit_r84_c73 bl[73] br[73] wl[84] vdd gnd cell_6t
Xbit_r85_c73 bl[73] br[73] wl[85] vdd gnd cell_6t
Xbit_r86_c73 bl[73] br[73] wl[86] vdd gnd cell_6t
Xbit_r87_c73 bl[73] br[73] wl[87] vdd gnd cell_6t
Xbit_r88_c73 bl[73] br[73] wl[88] vdd gnd cell_6t
Xbit_r89_c73 bl[73] br[73] wl[89] vdd gnd cell_6t
Xbit_r90_c73 bl[73] br[73] wl[90] vdd gnd cell_6t
Xbit_r91_c73 bl[73] br[73] wl[91] vdd gnd cell_6t
Xbit_r92_c73 bl[73] br[73] wl[92] vdd gnd cell_6t
Xbit_r93_c73 bl[73] br[73] wl[93] vdd gnd cell_6t
Xbit_r94_c73 bl[73] br[73] wl[94] vdd gnd cell_6t
Xbit_r95_c73 bl[73] br[73] wl[95] vdd gnd cell_6t
Xbit_r96_c73 bl[73] br[73] wl[96] vdd gnd cell_6t
Xbit_r97_c73 bl[73] br[73] wl[97] vdd gnd cell_6t
Xbit_r98_c73 bl[73] br[73] wl[98] vdd gnd cell_6t
Xbit_r99_c73 bl[73] br[73] wl[99] vdd gnd cell_6t
Xbit_r100_c73 bl[73] br[73] wl[100] vdd gnd cell_6t
Xbit_r101_c73 bl[73] br[73] wl[101] vdd gnd cell_6t
Xbit_r102_c73 bl[73] br[73] wl[102] vdd gnd cell_6t
Xbit_r103_c73 bl[73] br[73] wl[103] vdd gnd cell_6t
Xbit_r104_c73 bl[73] br[73] wl[104] vdd gnd cell_6t
Xbit_r105_c73 bl[73] br[73] wl[105] vdd gnd cell_6t
Xbit_r106_c73 bl[73] br[73] wl[106] vdd gnd cell_6t
Xbit_r107_c73 bl[73] br[73] wl[107] vdd gnd cell_6t
Xbit_r108_c73 bl[73] br[73] wl[108] vdd gnd cell_6t
Xbit_r109_c73 bl[73] br[73] wl[109] vdd gnd cell_6t
Xbit_r110_c73 bl[73] br[73] wl[110] vdd gnd cell_6t
Xbit_r111_c73 bl[73] br[73] wl[111] vdd gnd cell_6t
Xbit_r112_c73 bl[73] br[73] wl[112] vdd gnd cell_6t
Xbit_r113_c73 bl[73] br[73] wl[113] vdd gnd cell_6t
Xbit_r114_c73 bl[73] br[73] wl[114] vdd gnd cell_6t
Xbit_r115_c73 bl[73] br[73] wl[115] vdd gnd cell_6t
Xbit_r116_c73 bl[73] br[73] wl[116] vdd gnd cell_6t
Xbit_r117_c73 bl[73] br[73] wl[117] vdd gnd cell_6t
Xbit_r118_c73 bl[73] br[73] wl[118] vdd gnd cell_6t
Xbit_r119_c73 bl[73] br[73] wl[119] vdd gnd cell_6t
Xbit_r120_c73 bl[73] br[73] wl[120] vdd gnd cell_6t
Xbit_r121_c73 bl[73] br[73] wl[121] vdd gnd cell_6t
Xbit_r122_c73 bl[73] br[73] wl[122] vdd gnd cell_6t
Xbit_r123_c73 bl[73] br[73] wl[123] vdd gnd cell_6t
Xbit_r124_c73 bl[73] br[73] wl[124] vdd gnd cell_6t
Xbit_r125_c73 bl[73] br[73] wl[125] vdd gnd cell_6t
Xbit_r126_c73 bl[73] br[73] wl[126] vdd gnd cell_6t
Xbit_r127_c73 bl[73] br[73] wl[127] vdd gnd cell_6t
Xbit_r0_c74 bl[74] br[74] wl[0] vdd gnd cell_6t
Xbit_r1_c74 bl[74] br[74] wl[1] vdd gnd cell_6t
Xbit_r2_c74 bl[74] br[74] wl[2] vdd gnd cell_6t
Xbit_r3_c74 bl[74] br[74] wl[3] vdd gnd cell_6t
Xbit_r4_c74 bl[74] br[74] wl[4] vdd gnd cell_6t
Xbit_r5_c74 bl[74] br[74] wl[5] vdd gnd cell_6t
Xbit_r6_c74 bl[74] br[74] wl[6] vdd gnd cell_6t
Xbit_r7_c74 bl[74] br[74] wl[7] vdd gnd cell_6t
Xbit_r8_c74 bl[74] br[74] wl[8] vdd gnd cell_6t
Xbit_r9_c74 bl[74] br[74] wl[9] vdd gnd cell_6t
Xbit_r10_c74 bl[74] br[74] wl[10] vdd gnd cell_6t
Xbit_r11_c74 bl[74] br[74] wl[11] vdd gnd cell_6t
Xbit_r12_c74 bl[74] br[74] wl[12] vdd gnd cell_6t
Xbit_r13_c74 bl[74] br[74] wl[13] vdd gnd cell_6t
Xbit_r14_c74 bl[74] br[74] wl[14] vdd gnd cell_6t
Xbit_r15_c74 bl[74] br[74] wl[15] vdd gnd cell_6t
Xbit_r16_c74 bl[74] br[74] wl[16] vdd gnd cell_6t
Xbit_r17_c74 bl[74] br[74] wl[17] vdd gnd cell_6t
Xbit_r18_c74 bl[74] br[74] wl[18] vdd gnd cell_6t
Xbit_r19_c74 bl[74] br[74] wl[19] vdd gnd cell_6t
Xbit_r20_c74 bl[74] br[74] wl[20] vdd gnd cell_6t
Xbit_r21_c74 bl[74] br[74] wl[21] vdd gnd cell_6t
Xbit_r22_c74 bl[74] br[74] wl[22] vdd gnd cell_6t
Xbit_r23_c74 bl[74] br[74] wl[23] vdd gnd cell_6t
Xbit_r24_c74 bl[74] br[74] wl[24] vdd gnd cell_6t
Xbit_r25_c74 bl[74] br[74] wl[25] vdd gnd cell_6t
Xbit_r26_c74 bl[74] br[74] wl[26] vdd gnd cell_6t
Xbit_r27_c74 bl[74] br[74] wl[27] vdd gnd cell_6t
Xbit_r28_c74 bl[74] br[74] wl[28] vdd gnd cell_6t
Xbit_r29_c74 bl[74] br[74] wl[29] vdd gnd cell_6t
Xbit_r30_c74 bl[74] br[74] wl[30] vdd gnd cell_6t
Xbit_r31_c74 bl[74] br[74] wl[31] vdd gnd cell_6t
Xbit_r32_c74 bl[74] br[74] wl[32] vdd gnd cell_6t
Xbit_r33_c74 bl[74] br[74] wl[33] vdd gnd cell_6t
Xbit_r34_c74 bl[74] br[74] wl[34] vdd gnd cell_6t
Xbit_r35_c74 bl[74] br[74] wl[35] vdd gnd cell_6t
Xbit_r36_c74 bl[74] br[74] wl[36] vdd gnd cell_6t
Xbit_r37_c74 bl[74] br[74] wl[37] vdd gnd cell_6t
Xbit_r38_c74 bl[74] br[74] wl[38] vdd gnd cell_6t
Xbit_r39_c74 bl[74] br[74] wl[39] vdd gnd cell_6t
Xbit_r40_c74 bl[74] br[74] wl[40] vdd gnd cell_6t
Xbit_r41_c74 bl[74] br[74] wl[41] vdd gnd cell_6t
Xbit_r42_c74 bl[74] br[74] wl[42] vdd gnd cell_6t
Xbit_r43_c74 bl[74] br[74] wl[43] vdd gnd cell_6t
Xbit_r44_c74 bl[74] br[74] wl[44] vdd gnd cell_6t
Xbit_r45_c74 bl[74] br[74] wl[45] vdd gnd cell_6t
Xbit_r46_c74 bl[74] br[74] wl[46] vdd gnd cell_6t
Xbit_r47_c74 bl[74] br[74] wl[47] vdd gnd cell_6t
Xbit_r48_c74 bl[74] br[74] wl[48] vdd gnd cell_6t
Xbit_r49_c74 bl[74] br[74] wl[49] vdd gnd cell_6t
Xbit_r50_c74 bl[74] br[74] wl[50] vdd gnd cell_6t
Xbit_r51_c74 bl[74] br[74] wl[51] vdd gnd cell_6t
Xbit_r52_c74 bl[74] br[74] wl[52] vdd gnd cell_6t
Xbit_r53_c74 bl[74] br[74] wl[53] vdd gnd cell_6t
Xbit_r54_c74 bl[74] br[74] wl[54] vdd gnd cell_6t
Xbit_r55_c74 bl[74] br[74] wl[55] vdd gnd cell_6t
Xbit_r56_c74 bl[74] br[74] wl[56] vdd gnd cell_6t
Xbit_r57_c74 bl[74] br[74] wl[57] vdd gnd cell_6t
Xbit_r58_c74 bl[74] br[74] wl[58] vdd gnd cell_6t
Xbit_r59_c74 bl[74] br[74] wl[59] vdd gnd cell_6t
Xbit_r60_c74 bl[74] br[74] wl[60] vdd gnd cell_6t
Xbit_r61_c74 bl[74] br[74] wl[61] vdd gnd cell_6t
Xbit_r62_c74 bl[74] br[74] wl[62] vdd gnd cell_6t
Xbit_r63_c74 bl[74] br[74] wl[63] vdd gnd cell_6t
Xbit_r64_c74 bl[74] br[74] wl[64] vdd gnd cell_6t
Xbit_r65_c74 bl[74] br[74] wl[65] vdd gnd cell_6t
Xbit_r66_c74 bl[74] br[74] wl[66] vdd gnd cell_6t
Xbit_r67_c74 bl[74] br[74] wl[67] vdd gnd cell_6t
Xbit_r68_c74 bl[74] br[74] wl[68] vdd gnd cell_6t
Xbit_r69_c74 bl[74] br[74] wl[69] vdd gnd cell_6t
Xbit_r70_c74 bl[74] br[74] wl[70] vdd gnd cell_6t
Xbit_r71_c74 bl[74] br[74] wl[71] vdd gnd cell_6t
Xbit_r72_c74 bl[74] br[74] wl[72] vdd gnd cell_6t
Xbit_r73_c74 bl[74] br[74] wl[73] vdd gnd cell_6t
Xbit_r74_c74 bl[74] br[74] wl[74] vdd gnd cell_6t
Xbit_r75_c74 bl[74] br[74] wl[75] vdd gnd cell_6t
Xbit_r76_c74 bl[74] br[74] wl[76] vdd gnd cell_6t
Xbit_r77_c74 bl[74] br[74] wl[77] vdd gnd cell_6t
Xbit_r78_c74 bl[74] br[74] wl[78] vdd gnd cell_6t
Xbit_r79_c74 bl[74] br[74] wl[79] vdd gnd cell_6t
Xbit_r80_c74 bl[74] br[74] wl[80] vdd gnd cell_6t
Xbit_r81_c74 bl[74] br[74] wl[81] vdd gnd cell_6t
Xbit_r82_c74 bl[74] br[74] wl[82] vdd gnd cell_6t
Xbit_r83_c74 bl[74] br[74] wl[83] vdd gnd cell_6t
Xbit_r84_c74 bl[74] br[74] wl[84] vdd gnd cell_6t
Xbit_r85_c74 bl[74] br[74] wl[85] vdd gnd cell_6t
Xbit_r86_c74 bl[74] br[74] wl[86] vdd gnd cell_6t
Xbit_r87_c74 bl[74] br[74] wl[87] vdd gnd cell_6t
Xbit_r88_c74 bl[74] br[74] wl[88] vdd gnd cell_6t
Xbit_r89_c74 bl[74] br[74] wl[89] vdd gnd cell_6t
Xbit_r90_c74 bl[74] br[74] wl[90] vdd gnd cell_6t
Xbit_r91_c74 bl[74] br[74] wl[91] vdd gnd cell_6t
Xbit_r92_c74 bl[74] br[74] wl[92] vdd gnd cell_6t
Xbit_r93_c74 bl[74] br[74] wl[93] vdd gnd cell_6t
Xbit_r94_c74 bl[74] br[74] wl[94] vdd gnd cell_6t
Xbit_r95_c74 bl[74] br[74] wl[95] vdd gnd cell_6t
Xbit_r96_c74 bl[74] br[74] wl[96] vdd gnd cell_6t
Xbit_r97_c74 bl[74] br[74] wl[97] vdd gnd cell_6t
Xbit_r98_c74 bl[74] br[74] wl[98] vdd gnd cell_6t
Xbit_r99_c74 bl[74] br[74] wl[99] vdd gnd cell_6t
Xbit_r100_c74 bl[74] br[74] wl[100] vdd gnd cell_6t
Xbit_r101_c74 bl[74] br[74] wl[101] vdd gnd cell_6t
Xbit_r102_c74 bl[74] br[74] wl[102] vdd gnd cell_6t
Xbit_r103_c74 bl[74] br[74] wl[103] vdd gnd cell_6t
Xbit_r104_c74 bl[74] br[74] wl[104] vdd gnd cell_6t
Xbit_r105_c74 bl[74] br[74] wl[105] vdd gnd cell_6t
Xbit_r106_c74 bl[74] br[74] wl[106] vdd gnd cell_6t
Xbit_r107_c74 bl[74] br[74] wl[107] vdd gnd cell_6t
Xbit_r108_c74 bl[74] br[74] wl[108] vdd gnd cell_6t
Xbit_r109_c74 bl[74] br[74] wl[109] vdd gnd cell_6t
Xbit_r110_c74 bl[74] br[74] wl[110] vdd gnd cell_6t
Xbit_r111_c74 bl[74] br[74] wl[111] vdd gnd cell_6t
Xbit_r112_c74 bl[74] br[74] wl[112] vdd gnd cell_6t
Xbit_r113_c74 bl[74] br[74] wl[113] vdd gnd cell_6t
Xbit_r114_c74 bl[74] br[74] wl[114] vdd gnd cell_6t
Xbit_r115_c74 bl[74] br[74] wl[115] vdd gnd cell_6t
Xbit_r116_c74 bl[74] br[74] wl[116] vdd gnd cell_6t
Xbit_r117_c74 bl[74] br[74] wl[117] vdd gnd cell_6t
Xbit_r118_c74 bl[74] br[74] wl[118] vdd gnd cell_6t
Xbit_r119_c74 bl[74] br[74] wl[119] vdd gnd cell_6t
Xbit_r120_c74 bl[74] br[74] wl[120] vdd gnd cell_6t
Xbit_r121_c74 bl[74] br[74] wl[121] vdd gnd cell_6t
Xbit_r122_c74 bl[74] br[74] wl[122] vdd gnd cell_6t
Xbit_r123_c74 bl[74] br[74] wl[123] vdd gnd cell_6t
Xbit_r124_c74 bl[74] br[74] wl[124] vdd gnd cell_6t
Xbit_r125_c74 bl[74] br[74] wl[125] vdd gnd cell_6t
Xbit_r126_c74 bl[74] br[74] wl[126] vdd gnd cell_6t
Xbit_r127_c74 bl[74] br[74] wl[127] vdd gnd cell_6t
Xbit_r0_c75 bl[75] br[75] wl[0] vdd gnd cell_6t
Xbit_r1_c75 bl[75] br[75] wl[1] vdd gnd cell_6t
Xbit_r2_c75 bl[75] br[75] wl[2] vdd gnd cell_6t
Xbit_r3_c75 bl[75] br[75] wl[3] vdd gnd cell_6t
Xbit_r4_c75 bl[75] br[75] wl[4] vdd gnd cell_6t
Xbit_r5_c75 bl[75] br[75] wl[5] vdd gnd cell_6t
Xbit_r6_c75 bl[75] br[75] wl[6] vdd gnd cell_6t
Xbit_r7_c75 bl[75] br[75] wl[7] vdd gnd cell_6t
Xbit_r8_c75 bl[75] br[75] wl[8] vdd gnd cell_6t
Xbit_r9_c75 bl[75] br[75] wl[9] vdd gnd cell_6t
Xbit_r10_c75 bl[75] br[75] wl[10] vdd gnd cell_6t
Xbit_r11_c75 bl[75] br[75] wl[11] vdd gnd cell_6t
Xbit_r12_c75 bl[75] br[75] wl[12] vdd gnd cell_6t
Xbit_r13_c75 bl[75] br[75] wl[13] vdd gnd cell_6t
Xbit_r14_c75 bl[75] br[75] wl[14] vdd gnd cell_6t
Xbit_r15_c75 bl[75] br[75] wl[15] vdd gnd cell_6t
Xbit_r16_c75 bl[75] br[75] wl[16] vdd gnd cell_6t
Xbit_r17_c75 bl[75] br[75] wl[17] vdd gnd cell_6t
Xbit_r18_c75 bl[75] br[75] wl[18] vdd gnd cell_6t
Xbit_r19_c75 bl[75] br[75] wl[19] vdd gnd cell_6t
Xbit_r20_c75 bl[75] br[75] wl[20] vdd gnd cell_6t
Xbit_r21_c75 bl[75] br[75] wl[21] vdd gnd cell_6t
Xbit_r22_c75 bl[75] br[75] wl[22] vdd gnd cell_6t
Xbit_r23_c75 bl[75] br[75] wl[23] vdd gnd cell_6t
Xbit_r24_c75 bl[75] br[75] wl[24] vdd gnd cell_6t
Xbit_r25_c75 bl[75] br[75] wl[25] vdd gnd cell_6t
Xbit_r26_c75 bl[75] br[75] wl[26] vdd gnd cell_6t
Xbit_r27_c75 bl[75] br[75] wl[27] vdd gnd cell_6t
Xbit_r28_c75 bl[75] br[75] wl[28] vdd gnd cell_6t
Xbit_r29_c75 bl[75] br[75] wl[29] vdd gnd cell_6t
Xbit_r30_c75 bl[75] br[75] wl[30] vdd gnd cell_6t
Xbit_r31_c75 bl[75] br[75] wl[31] vdd gnd cell_6t
Xbit_r32_c75 bl[75] br[75] wl[32] vdd gnd cell_6t
Xbit_r33_c75 bl[75] br[75] wl[33] vdd gnd cell_6t
Xbit_r34_c75 bl[75] br[75] wl[34] vdd gnd cell_6t
Xbit_r35_c75 bl[75] br[75] wl[35] vdd gnd cell_6t
Xbit_r36_c75 bl[75] br[75] wl[36] vdd gnd cell_6t
Xbit_r37_c75 bl[75] br[75] wl[37] vdd gnd cell_6t
Xbit_r38_c75 bl[75] br[75] wl[38] vdd gnd cell_6t
Xbit_r39_c75 bl[75] br[75] wl[39] vdd gnd cell_6t
Xbit_r40_c75 bl[75] br[75] wl[40] vdd gnd cell_6t
Xbit_r41_c75 bl[75] br[75] wl[41] vdd gnd cell_6t
Xbit_r42_c75 bl[75] br[75] wl[42] vdd gnd cell_6t
Xbit_r43_c75 bl[75] br[75] wl[43] vdd gnd cell_6t
Xbit_r44_c75 bl[75] br[75] wl[44] vdd gnd cell_6t
Xbit_r45_c75 bl[75] br[75] wl[45] vdd gnd cell_6t
Xbit_r46_c75 bl[75] br[75] wl[46] vdd gnd cell_6t
Xbit_r47_c75 bl[75] br[75] wl[47] vdd gnd cell_6t
Xbit_r48_c75 bl[75] br[75] wl[48] vdd gnd cell_6t
Xbit_r49_c75 bl[75] br[75] wl[49] vdd gnd cell_6t
Xbit_r50_c75 bl[75] br[75] wl[50] vdd gnd cell_6t
Xbit_r51_c75 bl[75] br[75] wl[51] vdd gnd cell_6t
Xbit_r52_c75 bl[75] br[75] wl[52] vdd gnd cell_6t
Xbit_r53_c75 bl[75] br[75] wl[53] vdd gnd cell_6t
Xbit_r54_c75 bl[75] br[75] wl[54] vdd gnd cell_6t
Xbit_r55_c75 bl[75] br[75] wl[55] vdd gnd cell_6t
Xbit_r56_c75 bl[75] br[75] wl[56] vdd gnd cell_6t
Xbit_r57_c75 bl[75] br[75] wl[57] vdd gnd cell_6t
Xbit_r58_c75 bl[75] br[75] wl[58] vdd gnd cell_6t
Xbit_r59_c75 bl[75] br[75] wl[59] vdd gnd cell_6t
Xbit_r60_c75 bl[75] br[75] wl[60] vdd gnd cell_6t
Xbit_r61_c75 bl[75] br[75] wl[61] vdd gnd cell_6t
Xbit_r62_c75 bl[75] br[75] wl[62] vdd gnd cell_6t
Xbit_r63_c75 bl[75] br[75] wl[63] vdd gnd cell_6t
Xbit_r64_c75 bl[75] br[75] wl[64] vdd gnd cell_6t
Xbit_r65_c75 bl[75] br[75] wl[65] vdd gnd cell_6t
Xbit_r66_c75 bl[75] br[75] wl[66] vdd gnd cell_6t
Xbit_r67_c75 bl[75] br[75] wl[67] vdd gnd cell_6t
Xbit_r68_c75 bl[75] br[75] wl[68] vdd gnd cell_6t
Xbit_r69_c75 bl[75] br[75] wl[69] vdd gnd cell_6t
Xbit_r70_c75 bl[75] br[75] wl[70] vdd gnd cell_6t
Xbit_r71_c75 bl[75] br[75] wl[71] vdd gnd cell_6t
Xbit_r72_c75 bl[75] br[75] wl[72] vdd gnd cell_6t
Xbit_r73_c75 bl[75] br[75] wl[73] vdd gnd cell_6t
Xbit_r74_c75 bl[75] br[75] wl[74] vdd gnd cell_6t
Xbit_r75_c75 bl[75] br[75] wl[75] vdd gnd cell_6t
Xbit_r76_c75 bl[75] br[75] wl[76] vdd gnd cell_6t
Xbit_r77_c75 bl[75] br[75] wl[77] vdd gnd cell_6t
Xbit_r78_c75 bl[75] br[75] wl[78] vdd gnd cell_6t
Xbit_r79_c75 bl[75] br[75] wl[79] vdd gnd cell_6t
Xbit_r80_c75 bl[75] br[75] wl[80] vdd gnd cell_6t
Xbit_r81_c75 bl[75] br[75] wl[81] vdd gnd cell_6t
Xbit_r82_c75 bl[75] br[75] wl[82] vdd gnd cell_6t
Xbit_r83_c75 bl[75] br[75] wl[83] vdd gnd cell_6t
Xbit_r84_c75 bl[75] br[75] wl[84] vdd gnd cell_6t
Xbit_r85_c75 bl[75] br[75] wl[85] vdd gnd cell_6t
Xbit_r86_c75 bl[75] br[75] wl[86] vdd gnd cell_6t
Xbit_r87_c75 bl[75] br[75] wl[87] vdd gnd cell_6t
Xbit_r88_c75 bl[75] br[75] wl[88] vdd gnd cell_6t
Xbit_r89_c75 bl[75] br[75] wl[89] vdd gnd cell_6t
Xbit_r90_c75 bl[75] br[75] wl[90] vdd gnd cell_6t
Xbit_r91_c75 bl[75] br[75] wl[91] vdd gnd cell_6t
Xbit_r92_c75 bl[75] br[75] wl[92] vdd gnd cell_6t
Xbit_r93_c75 bl[75] br[75] wl[93] vdd gnd cell_6t
Xbit_r94_c75 bl[75] br[75] wl[94] vdd gnd cell_6t
Xbit_r95_c75 bl[75] br[75] wl[95] vdd gnd cell_6t
Xbit_r96_c75 bl[75] br[75] wl[96] vdd gnd cell_6t
Xbit_r97_c75 bl[75] br[75] wl[97] vdd gnd cell_6t
Xbit_r98_c75 bl[75] br[75] wl[98] vdd gnd cell_6t
Xbit_r99_c75 bl[75] br[75] wl[99] vdd gnd cell_6t
Xbit_r100_c75 bl[75] br[75] wl[100] vdd gnd cell_6t
Xbit_r101_c75 bl[75] br[75] wl[101] vdd gnd cell_6t
Xbit_r102_c75 bl[75] br[75] wl[102] vdd gnd cell_6t
Xbit_r103_c75 bl[75] br[75] wl[103] vdd gnd cell_6t
Xbit_r104_c75 bl[75] br[75] wl[104] vdd gnd cell_6t
Xbit_r105_c75 bl[75] br[75] wl[105] vdd gnd cell_6t
Xbit_r106_c75 bl[75] br[75] wl[106] vdd gnd cell_6t
Xbit_r107_c75 bl[75] br[75] wl[107] vdd gnd cell_6t
Xbit_r108_c75 bl[75] br[75] wl[108] vdd gnd cell_6t
Xbit_r109_c75 bl[75] br[75] wl[109] vdd gnd cell_6t
Xbit_r110_c75 bl[75] br[75] wl[110] vdd gnd cell_6t
Xbit_r111_c75 bl[75] br[75] wl[111] vdd gnd cell_6t
Xbit_r112_c75 bl[75] br[75] wl[112] vdd gnd cell_6t
Xbit_r113_c75 bl[75] br[75] wl[113] vdd gnd cell_6t
Xbit_r114_c75 bl[75] br[75] wl[114] vdd gnd cell_6t
Xbit_r115_c75 bl[75] br[75] wl[115] vdd gnd cell_6t
Xbit_r116_c75 bl[75] br[75] wl[116] vdd gnd cell_6t
Xbit_r117_c75 bl[75] br[75] wl[117] vdd gnd cell_6t
Xbit_r118_c75 bl[75] br[75] wl[118] vdd gnd cell_6t
Xbit_r119_c75 bl[75] br[75] wl[119] vdd gnd cell_6t
Xbit_r120_c75 bl[75] br[75] wl[120] vdd gnd cell_6t
Xbit_r121_c75 bl[75] br[75] wl[121] vdd gnd cell_6t
Xbit_r122_c75 bl[75] br[75] wl[122] vdd gnd cell_6t
Xbit_r123_c75 bl[75] br[75] wl[123] vdd gnd cell_6t
Xbit_r124_c75 bl[75] br[75] wl[124] vdd gnd cell_6t
Xbit_r125_c75 bl[75] br[75] wl[125] vdd gnd cell_6t
Xbit_r126_c75 bl[75] br[75] wl[126] vdd gnd cell_6t
Xbit_r127_c75 bl[75] br[75] wl[127] vdd gnd cell_6t
Xbit_r0_c76 bl[76] br[76] wl[0] vdd gnd cell_6t
Xbit_r1_c76 bl[76] br[76] wl[1] vdd gnd cell_6t
Xbit_r2_c76 bl[76] br[76] wl[2] vdd gnd cell_6t
Xbit_r3_c76 bl[76] br[76] wl[3] vdd gnd cell_6t
Xbit_r4_c76 bl[76] br[76] wl[4] vdd gnd cell_6t
Xbit_r5_c76 bl[76] br[76] wl[5] vdd gnd cell_6t
Xbit_r6_c76 bl[76] br[76] wl[6] vdd gnd cell_6t
Xbit_r7_c76 bl[76] br[76] wl[7] vdd gnd cell_6t
Xbit_r8_c76 bl[76] br[76] wl[8] vdd gnd cell_6t
Xbit_r9_c76 bl[76] br[76] wl[9] vdd gnd cell_6t
Xbit_r10_c76 bl[76] br[76] wl[10] vdd gnd cell_6t
Xbit_r11_c76 bl[76] br[76] wl[11] vdd gnd cell_6t
Xbit_r12_c76 bl[76] br[76] wl[12] vdd gnd cell_6t
Xbit_r13_c76 bl[76] br[76] wl[13] vdd gnd cell_6t
Xbit_r14_c76 bl[76] br[76] wl[14] vdd gnd cell_6t
Xbit_r15_c76 bl[76] br[76] wl[15] vdd gnd cell_6t
Xbit_r16_c76 bl[76] br[76] wl[16] vdd gnd cell_6t
Xbit_r17_c76 bl[76] br[76] wl[17] vdd gnd cell_6t
Xbit_r18_c76 bl[76] br[76] wl[18] vdd gnd cell_6t
Xbit_r19_c76 bl[76] br[76] wl[19] vdd gnd cell_6t
Xbit_r20_c76 bl[76] br[76] wl[20] vdd gnd cell_6t
Xbit_r21_c76 bl[76] br[76] wl[21] vdd gnd cell_6t
Xbit_r22_c76 bl[76] br[76] wl[22] vdd gnd cell_6t
Xbit_r23_c76 bl[76] br[76] wl[23] vdd gnd cell_6t
Xbit_r24_c76 bl[76] br[76] wl[24] vdd gnd cell_6t
Xbit_r25_c76 bl[76] br[76] wl[25] vdd gnd cell_6t
Xbit_r26_c76 bl[76] br[76] wl[26] vdd gnd cell_6t
Xbit_r27_c76 bl[76] br[76] wl[27] vdd gnd cell_6t
Xbit_r28_c76 bl[76] br[76] wl[28] vdd gnd cell_6t
Xbit_r29_c76 bl[76] br[76] wl[29] vdd gnd cell_6t
Xbit_r30_c76 bl[76] br[76] wl[30] vdd gnd cell_6t
Xbit_r31_c76 bl[76] br[76] wl[31] vdd gnd cell_6t
Xbit_r32_c76 bl[76] br[76] wl[32] vdd gnd cell_6t
Xbit_r33_c76 bl[76] br[76] wl[33] vdd gnd cell_6t
Xbit_r34_c76 bl[76] br[76] wl[34] vdd gnd cell_6t
Xbit_r35_c76 bl[76] br[76] wl[35] vdd gnd cell_6t
Xbit_r36_c76 bl[76] br[76] wl[36] vdd gnd cell_6t
Xbit_r37_c76 bl[76] br[76] wl[37] vdd gnd cell_6t
Xbit_r38_c76 bl[76] br[76] wl[38] vdd gnd cell_6t
Xbit_r39_c76 bl[76] br[76] wl[39] vdd gnd cell_6t
Xbit_r40_c76 bl[76] br[76] wl[40] vdd gnd cell_6t
Xbit_r41_c76 bl[76] br[76] wl[41] vdd gnd cell_6t
Xbit_r42_c76 bl[76] br[76] wl[42] vdd gnd cell_6t
Xbit_r43_c76 bl[76] br[76] wl[43] vdd gnd cell_6t
Xbit_r44_c76 bl[76] br[76] wl[44] vdd gnd cell_6t
Xbit_r45_c76 bl[76] br[76] wl[45] vdd gnd cell_6t
Xbit_r46_c76 bl[76] br[76] wl[46] vdd gnd cell_6t
Xbit_r47_c76 bl[76] br[76] wl[47] vdd gnd cell_6t
Xbit_r48_c76 bl[76] br[76] wl[48] vdd gnd cell_6t
Xbit_r49_c76 bl[76] br[76] wl[49] vdd gnd cell_6t
Xbit_r50_c76 bl[76] br[76] wl[50] vdd gnd cell_6t
Xbit_r51_c76 bl[76] br[76] wl[51] vdd gnd cell_6t
Xbit_r52_c76 bl[76] br[76] wl[52] vdd gnd cell_6t
Xbit_r53_c76 bl[76] br[76] wl[53] vdd gnd cell_6t
Xbit_r54_c76 bl[76] br[76] wl[54] vdd gnd cell_6t
Xbit_r55_c76 bl[76] br[76] wl[55] vdd gnd cell_6t
Xbit_r56_c76 bl[76] br[76] wl[56] vdd gnd cell_6t
Xbit_r57_c76 bl[76] br[76] wl[57] vdd gnd cell_6t
Xbit_r58_c76 bl[76] br[76] wl[58] vdd gnd cell_6t
Xbit_r59_c76 bl[76] br[76] wl[59] vdd gnd cell_6t
Xbit_r60_c76 bl[76] br[76] wl[60] vdd gnd cell_6t
Xbit_r61_c76 bl[76] br[76] wl[61] vdd gnd cell_6t
Xbit_r62_c76 bl[76] br[76] wl[62] vdd gnd cell_6t
Xbit_r63_c76 bl[76] br[76] wl[63] vdd gnd cell_6t
Xbit_r64_c76 bl[76] br[76] wl[64] vdd gnd cell_6t
Xbit_r65_c76 bl[76] br[76] wl[65] vdd gnd cell_6t
Xbit_r66_c76 bl[76] br[76] wl[66] vdd gnd cell_6t
Xbit_r67_c76 bl[76] br[76] wl[67] vdd gnd cell_6t
Xbit_r68_c76 bl[76] br[76] wl[68] vdd gnd cell_6t
Xbit_r69_c76 bl[76] br[76] wl[69] vdd gnd cell_6t
Xbit_r70_c76 bl[76] br[76] wl[70] vdd gnd cell_6t
Xbit_r71_c76 bl[76] br[76] wl[71] vdd gnd cell_6t
Xbit_r72_c76 bl[76] br[76] wl[72] vdd gnd cell_6t
Xbit_r73_c76 bl[76] br[76] wl[73] vdd gnd cell_6t
Xbit_r74_c76 bl[76] br[76] wl[74] vdd gnd cell_6t
Xbit_r75_c76 bl[76] br[76] wl[75] vdd gnd cell_6t
Xbit_r76_c76 bl[76] br[76] wl[76] vdd gnd cell_6t
Xbit_r77_c76 bl[76] br[76] wl[77] vdd gnd cell_6t
Xbit_r78_c76 bl[76] br[76] wl[78] vdd gnd cell_6t
Xbit_r79_c76 bl[76] br[76] wl[79] vdd gnd cell_6t
Xbit_r80_c76 bl[76] br[76] wl[80] vdd gnd cell_6t
Xbit_r81_c76 bl[76] br[76] wl[81] vdd gnd cell_6t
Xbit_r82_c76 bl[76] br[76] wl[82] vdd gnd cell_6t
Xbit_r83_c76 bl[76] br[76] wl[83] vdd gnd cell_6t
Xbit_r84_c76 bl[76] br[76] wl[84] vdd gnd cell_6t
Xbit_r85_c76 bl[76] br[76] wl[85] vdd gnd cell_6t
Xbit_r86_c76 bl[76] br[76] wl[86] vdd gnd cell_6t
Xbit_r87_c76 bl[76] br[76] wl[87] vdd gnd cell_6t
Xbit_r88_c76 bl[76] br[76] wl[88] vdd gnd cell_6t
Xbit_r89_c76 bl[76] br[76] wl[89] vdd gnd cell_6t
Xbit_r90_c76 bl[76] br[76] wl[90] vdd gnd cell_6t
Xbit_r91_c76 bl[76] br[76] wl[91] vdd gnd cell_6t
Xbit_r92_c76 bl[76] br[76] wl[92] vdd gnd cell_6t
Xbit_r93_c76 bl[76] br[76] wl[93] vdd gnd cell_6t
Xbit_r94_c76 bl[76] br[76] wl[94] vdd gnd cell_6t
Xbit_r95_c76 bl[76] br[76] wl[95] vdd gnd cell_6t
Xbit_r96_c76 bl[76] br[76] wl[96] vdd gnd cell_6t
Xbit_r97_c76 bl[76] br[76] wl[97] vdd gnd cell_6t
Xbit_r98_c76 bl[76] br[76] wl[98] vdd gnd cell_6t
Xbit_r99_c76 bl[76] br[76] wl[99] vdd gnd cell_6t
Xbit_r100_c76 bl[76] br[76] wl[100] vdd gnd cell_6t
Xbit_r101_c76 bl[76] br[76] wl[101] vdd gnd cell_6t
Xbit_r102_c76 bl[76] br[76] wl[102] vdd gnd cell_6t
Xbit_r103_c76 bl[76] br[76] wl[103] vdd gnd cell_6t
Xbit_r104_c76 bl[76] br[76] wl[104] vdd gnd cell_6t
Xbit_r105_c76 bl[76] br[76] wl[105] vdd gnd cell_6t
Xbit_r106_c76 bl[76] br[76] wl[106] vdd gnd cell_6t
Xbit_r107_c76 bl[76] br[76] wl[107] vdd gnd cell_6t
Xbit_r108_c76 bl[76] br[76] wl[108] vdd gnd cell_6t
Xbit_r109_c76 bl[76] br[76] wl[109] vdd gnd cell_6t
Xbit_r110_c76 bl[76] br[76] wl[110] vdd gnd cell_6t
Xbit_r111_c76 bl[76] br[76] wl[111] vdd gnd cell_6t
Xbit_r112_c76 bl[76] br[76] wl[112] vdd gnd cell_6t
Xbit_r113_c76 bl[76] br[76] wl[113] vdd gnd cell_6t
Xbit_r114_c76 bl[76] br[76] wl[114] vdd gnd cell_6t
Xbit_r115_c76 bl[76] br[76] wl[115] vdd gnd cell_6t
Xbit_r116_c76 bl[76] br[76] wl[116] vdd gnd cell_6t
Xbit_r117_c76 bl[76] br[76] wl[117] vdd gnd cell_6t
Xbit_r118_c76 bl[76] br[76] wl[118] vdd gnd cell_6t
Xbit_r119_c76 bl[76] br[76] wl[119] vdd gnd cell_6t
Xbit_r120_c76 bl[76] br[76] wl[120] vdd gnd cell_6t
Xbit_r121_c76 bl[76] br[76] wl[121] vdd gnd cell_6t
Xbit_r122_c76 bl[76] br[76] wl[122] vdd gnd cell_6t
Xbit_r123_c76 bl[76] br[76] wl[123] vdd gnd cell_6t
Xbit_r124_c76 bl[76] br[76] wl[124] vdd gnd cell_6t
Xbit_r125_c76 bl[76] br[76] wl[125] vdd gnd cell_6t
Xbit_r126_c76 bl[76] br[76] wl[126] vdd gnd cell_6t
Xbit_r127_c76 bl[76] br[76] wl[127] vdd gnd cell_6t
Xbit_r0_c77 bl[77] br[77] wl[0] vdd gnd cell_6t
Xbit_r1_c77 bl[77] br[77] wl[1] vdd gnd cell_6t
Xbit_r2_c77 bl[77] br[77] wl[2] vdd gnd cell_6t
Xbit_r3_c77 bl[77] br[77] wl[3] vdd gnd cell_6t
Xbit_r4_c77 bl[77] br[77] wl[4] vdd gnd cell_6t
Xbit_r5_c77 bl[77] br[77] wl[5] vdd gnd cell_6t
Xbit_r6_c77 bl[77] br[77] wl[6] vdd gnd cell_6t
Xbit_r7_c77 bl[77] br[77] wl[7] vdd gnd cell_6t
Xbit_r8_c77 bl[77] br[77] wl[8] vdd gnd cell_6t
Xbit_r9_c77 bl[77] br[77] wl[9] vdd gnd cell_6t
Xbit_r10_c77 bl[77] br[77] wl[10] vdd gnd cell_6t
Xbit_r11_c77 bl[77] br[77] wl[11] vdd gnd cell_6t
Xbit_r12_c77 bl[77] br[77] wl[12] vdd gnd cell_6t
Xbit_r13_c77 bl[77] br[77] wl[13] vdd gnd cell_6t
Xbit_r14_c77 bl[77] br[77] wl[14] vdd gnd cell_6t
Xbit_r15_c77 bl[77] br[77] wl[15] vdd gnd cell_6t
Xbit_r16_c77 bl[77] br[77] wl[16] vdd gnd cell_6t
Xbit_r17_c77 bl[77] br[77] wl[17] vdd gnd cell_6t
Xbit_r18_c77 bl[77] br[77] wl[18] vdd gnd cell_6t
Xbit_r19_c77 bl[77] br[77] wl[19] vdd gnd cell_6t
Xbit_r20_c77 bl[77] br[77] wl[20] vdd gnd cell_6t
Xbit_r21_c77 bl[77] br[77] wl[21] vdd gnd cell_6t
Xbit_r22_c77 bl[77] br[77] wl[22] vdd gnd cell_6t
Xbit_r23_c77 bl[77] br[77] wl[23] vdd gnd cell_6t
Xbit_r24_c77 bl[77] br[77] wl[24] vdd gnd cell_6t
Xbit_r25_c77 bl[77] br[77] wl[25] vdd gnd cell_6t
Xbit_r26_c77 bl[77] br[77] wl[26] vdd gnd cell_6t
Xbit_r27_c77 bl[77] br[77] wl[27] vdd gnd cell_6t
Xbit_r28_c77 bl[77] br[77] wl[28] vdd gnd cell_6t
Xbit_r29_c77 bl[77] br[77] wl[29] vdd gnd cell_6t
Xbit_r30_c77 bl[77] br[77] wl[30] vdd gnd cell_6t
Xbit_r31_c77 bl[77] br[77] wl[31] vdd gnd cell_6t
Xbit_r32_c77 bl[77] br[77] wl[32] vdd gnd cell_6t
Xbit_r33_c77 bl[77] br[77] wl[33] vdd gnd cell_6t
Xbit_r34_c77 bl[77] br[77] wl[34] vdd gnd cell_6t
Xbit_r35_c77 bl[77] br[77] wl[35] vdd gnd cell_6t
Xbit_r36_c77 bl[77] br[77] wl[36] vdd gnd cell_6t
Xbit_r37_c77 bl[77] br[77] wl[37] vdd gnd cell_6t
Xbit_r38_c77 bl[77] br[77] wl[38] vdd gnd cell_6t
Xbit_r39_c77 bl[77] br[77] wl[39] vdd gnd cell_6t
Xbit_r40_c77 bl[77] br[77] wl[40] vdd gnd cell_6t
Xbit_r41_c77 bl[77] br[77] wl[41] vdd gnd cell_6t
Xbit_r42_c77 bl[77] br[77] wl[42] vdd gnd cell_6t
Xbit_r43_c77 bl[77] br[77] wl[43] vdd gnd cell_6t
Xbit_r44_c77 bl[77] br[77] wl[44] vdd gnd cell_6t
Xbit_r45_c77 bl[77] br[77] wl[45] vdd gnd cell_6t
Xbit_r46_c77 bl[77] br[77] wl[46] vdd gnd cell_6t
Xbit_r47_c77 bl[77] br[77] wl[47] vdd gnd cell_6t
Xbit_r48_c77 bl[77] br[77] wl[48] vdd gnd cell_6t
Xbit_r49_c77 bl[77] br[77] wl[49] vdd gnd cell_6t
Xbit_r50_c77 bl[77] br[77] wl[50] vdd gnd cell_6t
Xbit_r51_c77 bl[77] br[77] wl[51] vdd gnd cell_6t
Xbit_r52_c77 bl[77] br[77] wl[52] vdd gnd cell_6t
Xbit_r53_c77 bl[77] br[77] wl[53] vdd gnd cell_6t
Xbit_r54_c77 bl[77] br[77] wl[54] vdd gnd cell_6t
Xbit_r55_c77 bl[77] br[77] wl[55] vdd gnd cell_6t
Xbit_r56_c77 bl[77] br[77] wl[56] vdd gnd cell_6t
Xbit_r57_c77 bl[77] br[77] wl[57] vdd gnd cell_6t
Xbit_r58_c77 bl[77] br[77] wl[58] vdd gnd cell_6t
Xbit_r59_c77 bl[77] br[77] wl[59] vdd gnd cell_6t
Xbit_r60_c77 bl[77] br[77] wl[60] vdd gnd cell_6t
Xbit_r61_c77 bl[77] br[77] wl[61] vdd gnd cell_6t
Xbit_r62_c77 bl[77] br[77] wl[62] vdd gnd cell_6t
Xbit_r63_c77 bl[77] br[77] wl[63] vdd gnd cell_6t
Xbit_r64_c77 bl[77] br[77] wl[64] vdd gnd cell_6t
Xbit_r65_c77 bl[77] br[77] wl[65] vdd gnd cell_6t
Xbit_r66_c77 bl[77] br[77] wl[66] vdd gnd cell_6t
Xbit_r67_c77 bl[77] br[77] wl[67] vdd gnd cell_6t
Xbit_r68_c77 bl[77] br[77] wl[68] vdd gnd cell_6t
Xbit_r69_c77 bl[77] br[77] wl[69] vdd gnd cell_6t
Xbit_r70_c77 bl[77] br[77] wl[70] vdd gnd cell_6t
Xbit_r71_c77 bl[77] br[77] wl[71] vdd gnd cell_6t
Xbit_r72_c77 bl[77] br[77] wl[72] vdd gnd cell_6t
Xbit_r73_c77 bl[77] br[77] wl[73] vdd gnd cell_6t
Xbit_r74_c77 bl[77] br[77] wl[74] vdd gnd cell_6t
Xbit_r75_c77 bl[77] br[77] wl[75] vdd gnd cell_6t
Xbit_r76_c77 bl[77] br[77] wl[76] vdd gnd cell_6t
Xbit_r77_c77 bl[77] br[77] wl[77] vdd gnd cell_6t
Xbit_r78_c77 bl[77] br[77] wl[78] vdd gnd cell_6t
Xbit_r79_c77 bl[77] br[77] wl[79] vdd gnd cell_6t
Xbit_r80_c77 bl[77] br[77] wl[80] vdd gnd cell_6t
Xbit_r81_c77 bl[77] br[77] wl[81] vdd gnd cell_6t
Xbit_r82_c77 bl[77] br[77] wl[82] vdd gnd cell_6t
Xbit_r83_c77 bl[77] br[77] wl[83] vdd gnd cell_6t
Xbit_r84_c77 bl[77] br[77] wl[84] vdd gnd cell_6t
Xbit_r85_c77 bl[77] br[77] wl[85] vdd gnd cell_6t
Xbit_r86_c77 bl[77] br[77] wl[86] vdd gnd cell_6t
Xbit_r87_c77 bl[77] br[77] wl[87] vdd gnd cell_6t
Xbit_r88_c77 bl[77] br[77] wl[88] vdd gnd cell_6t
Xbit_r89_c77 bl[77] br[77] wl[89] vdd gnd cell_6t
Xbit_r90_c77 bl[77] br[77] wl[90] vdd gnd cell_6t
Xbit_r91_c77 bl[77] br[77] wl[91] vdd gnd cell_6t
Xbit_r92_c77 bl[77] br[77] wl[92] vdd gnd cell_6t
Xbit_r93_c77 bl[77] br[77] wl[93] vdd gnd cell_6t
Xbit_r94_c77 bl[77] br[77] wl[94] vdd gnd cell_6t
Xbit_r95_c77 bl[77] br[77] wl[95] vdd gnd cell_6t
Xbit_r96_c77 bl[77] br[77] wl[96] vdd gnd cell_6t
Xbit_r97_c77 bl[77] br[77] wl[97] vdd gnd cell_6t
Xbit_r98_c77 bl[77] br[77] wl[98] vdd gnd cell_6t
Xbit_r99_c77 bl[77] br[77] wl[99] vdd gnd cell_6t
Xbit_r100_c77 bl[77] br[77] wl[100] vdd gnd cell_6t
Xbit_r101_c77 bl[77] br[77] wl[101] vdd gnd cell_6t
Xbit_r102_c77 bl[77] br[77] wl[102] vdd gnd cell_6t
Xbit_r103_c77 bl[77] br[77] wl[103] vdd gnd cell_6t
Xbit_r104_c77 bl[77] br[77] wl[104] vdd gnd cell_6t
Xbit_r105_c77 bl[77] br[77] wl[105] vdd gnd cell_6t
Xbit_r106_c77 bl[77] br[77] wl[106] vdd gnd cell_6t
Xbit_r107_c77 bl[77] br[77] wl[107] vdd gnd cell_6t
Xbit_r108_c77 bl[77] br[77] wl[108] vdd gnd cell_6t
Xbit_r109_c77 bl[77] br[77] wl[109] vdd gnd cell_6t
Xbit_r110_c77 bl[77] br[77] wl[110] vdd gnd cell_6t
Xbit_r111_c77 bl[77] br[77] wl[111] vdd gnd cell_6t
Xbit_r112_c77 bl[77] br[77] wl[112] vdd gnd cell_6t
Xbit_r113_c77 bl[77] br[77] wl[113] vdd gnd cell_6t
Xbit_r114_c77 bl[77] br[77] wl[114] vdd gnd cell_6t
Xbit_r115_c77 bl[77] br[77] wl[115] vdd gnd cell_6t
Xbit_r116_c77 bl[77] br[77] wl[116] vdd gnd cell_6t
Xbit_r117_c77 bl[77] br[77] wl[117] vdd gnd cell_6t
Xbit_r118_c77 bl[77] br[77] wl[118] vdd gnd cell_6t
Xbit_r119_c77 bl[77] br[77] wl[119] vdd gnd cell_6t
Xbit_r120_c77 bl[77] br[77] wl[120] vdd gnd cell_6t
Xbit_r121_c77 bl[77] br[77] wl[121] vdd gnd cell_6t
Xbit_r122_c77 bl[77] br[77] wl[122] vdd gnd cell_6t
Xbit_r123_c77 bl[77] br[77] wl[123] vdd gnd cell_6t
Xbit_r124_c77 bl[77] br[77] wl[124] vdd gnd cell_6t
Xbit_r125_c77 bl[77] br[77] wl[125] vdd gnd cell_6t
Xbit_r126_c77 bl[77] br[77] wl[126] vdd gnd cell_6t
Xbit_r127_c77 bl[77] br[77] wl[127] vdd gnd cell_6t
Xbit_r0_c78 bl[78] br[78] wl[0] vdd gnd cell_6t
Xbit_r1_c78 bl[78] br[78] wl[1] vdd gnd cell_6t
Xbit_r2_c78 bl[78] br[78] wl[2] vdd gnd cell_6t
Xbit_r3_c78 bl[78] br[78] wl[3] vdd gnd cell_6t
Xbit_r4_c78 bl[78] br[78] wl[4] vdd gnd cell_6t
Xbit_r5_c78 bl[78] br[78] wl[5] vdd gnd cell_6t
Xbit_r6_c78 bl[78] br[78] wl[6] vdd gnd cell_6t
Xbit_r7_c78 bl[78] br[78] wl[7] vdd gnd cell_6t
Xbit_r8_c78 bl[78] br[78] wl[8] vdd gnd cell_6t
Xbit_r9_c78 bl[78] br[78] wl[9] vdd gnd cell_6t
Xbit_r10_c78 bl[78] br[78] wl[10] vdd gnd cell_6t
Xbit_r11_c78 bl[78] br[78] wl[11] vdd gnd cell_6t
Xbit_r12_c78 bl[78] br[78] wl[12] vdd gnd cell_6t
Xbit_r13_c78 bl[78] br[78] wl[13] vdd gnd cell_6t
Xbit_r14_c78 bl[78] br[78] wl[14] vdd gnd cell_6t
Xbit_r15_c78 bl[78] br[78] wl[15] vdd gnd cell_6t
Xbit_r16_c78 bl[78] br[78] wl[16] vdd gnd cell_6t
Xbit_r17_c78 bl[78] br[78] wl[17] vdd gnd cell_6t
Xbit_r18_c78 bl[78] br[78] wl[18] vdd gnd cell_6t
Xbit_r19_c78 bl[78] br[78] wl[19] vdd gnd cell_6t
Xbit_r20_c78 bl[78] br[78] wl[20] vdd gnd cell_6t
Xbit_r21_c78 bl[78] br[78] wl[21] vdd gnd cell_6t
Xbit_r22_c78 bl[78] br[78] wl[22] vdd gnd cell_6t
Xbit_r23_c78 bl[78] br[78] wl[23] vdd gnd cell_6t
Xbit_r24_c78 bl[78] br[78] wl[24] vdd gnd cell_6t
Xbit_r25_c78 bl[78] br[78] wl[25] vdd gnd cell_6t
Xbit_r26_c78 bl[78] br[78] wl[26] vdd gnd cell_6t
Xbit_r27_c78 bl[78] br[78] wl[27] vdd gnd cell_6t
Xbit_r28_c78 bl[78] br[78] wl[28] vdd gnd cell_6t
Xbit_r29_c78 bl[78] br[78] wl[29] vdd gnd cell_6t
Xbit_r30_c78 bl[78] br[78] wl[30] vdd gnd cell_6t
Xbit_r31_c78 bl[78] br[78] wl[31] vdd gnd cell_6t
Xbit_r32_c78 bl[78] br[78] wl[32] vdd gnd cell_6t
Xbit_r33_c78 bl[78] br[78] wl[33] vdd gnd cell_6t
Xbit_r34_c78 bl[78] br[78] wl[34] vdd gnd cell_6t
Xbit_r35_c78 bl[78] br[78] wl[35] vdd gnd cell_6t
Xbit_r36_c78 bl[78] br[78] wl[36] vdd gnd cell_6t
Xbit_r37_c78 bl[78] br[78] wl[37] vdd gnd cell_6t
Xbit_r38_c78 bl[78] br[78] wl[38] vdd gnd cell_6t
Xbit_r39_c78 bl[78] br[78] wl[39] vdd gnd cell_6t
Xbit_r40_c78 bl[78] br[78] wl[40] vdd gnd cell_6t
Xbit_r41_c78 bl[78] br[78] wl[41] vdd gnd cell_6t
Xbit_r42_c78 bl[78] br[78] wl[42] vdd gnd cell_6t
Xbit_r43_c78 bl[78] br[78] wl[43] vdd gnd cell_6t
Xbit_r44_c78 bl[78] br[78] wl[44] vdd gnd cell_6t
Xbit_r45_c78 bl[78] br[78] wl[45] vdd gnd cell_6t
Xbit_r46_c78 bl[78] br[78] wl[46] vdd gnd cell_6t
Xbit_r47_c78 bl[78] br[78] wl[47] vdd gnd cell_6t
Xbit_r48_c78 bl[78] br[78] wl[48] vdd gnd cell_6t
Xbit_r49_c78 bl[78] br[78] wl[49] vdd gnd cell_6t
Xbit_r50_c78 bl[78] br[78] wl[50] vdd gnd cell_6t
Xbit_r51_c78 bl[78] br[78] wl[51] vdd gnd cell_6t
Xbit_r52_c78 bl[78] br[78] wl[52] vdd gnd cell_6t
Xbit_r53_c78 bl[78] br[78] wl[53] vdd gnd cell_6t
Xbit_r54_c78 bl[78] br[78] wl[54] vdd gnd cell_6t
Xbit_r55_c78 bl[78] br[78] wl[55] vdd gnd cell_6t
Xbit_r56_c78 bl[78] br[78] wl[56] vdd gnd cell_6t
Xbit_r57_c78 bl[78] br[78] wl[57] vdd gnd cell_6t
Xbit_r58_c78 bl[78] br[78] wl[58] vdd gnd cell_6t
Xbit_r59_c78 bl[78] br[78] wl[59] vdd gnd cell_6t
Xbit_r60_c78 bl[78] br[78] wl[60] vdd gnd cell_6t
Xbit_r61_c78 bl[78] br[78] wl[61] vdd gnd cell_6t
Xbit_r62_c78 bl[78] br[78] wl[62] vdd gnd cell_6t
Xbit_r63_c78 bl[78] br[78] wl[63] vdd gnd cell_6t
Xbit_r64_c78 bl[78] br[78] wl[64] vdd gnd cell_6t
Xbit_r65_c78 bl[78] br[78] wl[65] vdd gnd cell_6t
Xbit_r66_c78 bl[78] br[78] wl[66] vdd gnd cell_6t
Xbit_r67_c78 bl[78] br[78] wl[67] vdd gnd cell_6t
Xbit_r68_c78 bl[78] br[78] wl[68] vdd gnd cell_6t
Xbit_r69_c78 bl[78] br[78] wl[69] vdd gnd cell_6t
Xbit_r70_c78 bl[78] br[78] wl[70] vdd gnd cell_6t
Xbit_r71_c78 bl[78] br[78] wl[71] vdd gnd cell_6t
Xbit_r72_c78 bl[78] br[78] wl[72] vdd gnd cell_6t
Xbit_r73_c78 bl[78] br[78] wl[73] vdd gnd cell_6t
Xbit_r74_c78 bl[78] br[78] wl[74] vdd gnd cell_6t
Xbit_r75_c78 bl[78] br[78] wl[75] vdd gnd cell_6t
Xbit_r76_c78 bl[78] br[78] wl[76] vdd gnd cell_6t
Xbit_r77_c78 bl[78] br[78] wl[77] vdd gnd cell_6t
Xbit_r78_c78 bl[78] br[78] wl[78] vdd gnd cell_6t
Xbit_r79_c78 bl[78] br[78] wl[79] vdd gnd cell_6t
Xbit_r80_c78 bl[78] br[78] wl[80] vdd gnd cell_6t
Xbit_r81_c78 bl[78] br[78] wl[81] vdd gnd cell_6t
Xbit_r82_c78 bl[78] br[78] wl[82] vdd gnd cell_6t
Xbit_r83_c78 bl[78] br[78] wl[83] vdd gnd cell_6t
Xbit_r84_c78 bl[78] br[78] wl[84] vdd gnd cell_6t
Xbit_r85_c78 bl[78] br[78] wl[85] vdd gnd cell_6t
Xbit_r86_c78 bl[78] br[78] wl[86] vdd gnd cell_6t
Xbit_r87_c78 bl[78] br[78] wl[87] vdd gnd cell_6t
Xbit_r88_c78 bl[78] br[78] wl[88] vdd gnd cell_6t
Xbit_r89_c78 bl[78] br[78] wl[89] vdd gnd cell_6t
Xbit_r90_c78 bl[78] br[78] wl[90] vdd gnd cell_6t
Xbit_r91_c78 bl[78] br[78] wl[91] vdd gnd cell_6t
Xbit_r92_c78 bl[78] br[78] wl[92] vdd gnd cell_6t
Xbit_r93_c78 bl[78] br[78] wl[93] vdd gnd cell_6t
Xbit_r94_c78 bl[78] br[78] wl[94] vdd gnd cell_6t
Xbit_r95_c78 bl[78] br[78] wl[95] vdd gnd cell_6t
Xbit_r96_c78 bl[78] br[78] wl[96] vdd gnd cell_6t
Xbit_r97_c78 bl[78] br[78] wl[97] vdd gnd cell_6t
Xbit_r98_c78 bl[78] br[78] wl[98] vdd gnd cell_6t
Xbit_r99_c78 bl[78] br[78] wl[99] vdd gnd cell_6t
Xbit_r100_c78 bl[78] br[78] wl[100] vdd gnd cell_6t
Xbit_r101_c78 bl[78] br[78] wl[101] vdd gnd cell_6t
Xbit_r102_c78 bl[78] br[78] wl[102] vdd gnd cell_6t
Xbit_r103_c78 bl[78] br[78] wl[103] vdd gnd cell_6t
Xbit_r104_c78 bl[78] br[78] wl[104] vdd gnd cell_6t
Xbit_r105_c78 bl[78] br[78] wl[105] vdd gnd cell_6t
Xbit_r106_c78 bl[78] br[78] wl[106] vdd gnd cell_6t
Xbit_r107_c78 bl[78] br[78] wl[107] vdd gnd cell_6t
Xbit_r108_c78 bl[78] br[78] wl[108] vdd gnd cell_6t
Xbit_r109_c78 bl[78] br[78] wl[109] vdd gnd cell_6t
Xbit_r110_c78 bl[78] br[78] wl[110] vdd gnd cell_6t
Xbit_r111_c78 bl[78] br[78] wl[111] vdd gnd cell_6t
Xbit_r112_c78 bl[78] br[78] wl[112] vdd gnd cell_6t
Xbit_r113_c78 bl[78] br[78] wl[113] vdd gnd cell_6t
Xbit_r114_c78 bl[78] br[78] wl[114] vdd gnd cell_6t
Xbit_r115_c78 bl[78] br[78] wl[115] vdd gnd cell_6t
Xbit_r116_c78 bl[78] br[78] wl[116] vdd gnd cell_6t
Xbit_r117_c78 bl[78] br[78] wl[117] vdd gnd cell_6t
Xbit_r118_c78 bl[78] br[78] wl[118] vdd gnd cell_6t
Xbit_r119_c78 bl[78] br[78] wl[119] vdd gnd cell_6t
Xbit_r120_c78 bl[78] br[78] wl[120] vdd gnd cell_6t
Xbit_r121_c78 bl[78] br[78] wl[121] vdd gnd cell_6t
Xbit_r122_c78 bl[78] br[78] wl[122] vdd gnd cell_6t
Xbit_r123_c78 bl[78] br[78] wl[123] vdd gnd cell_6t
Xbit_r124_c78 bl[78] br[78] wl[124] vdd gnd cell_6t
Xbit_r125_c78 bl[78] br[78] wl[125] vdd gnd cell_6t
Xbit_r126_c78 bl[78] br[78] wl[126] vdd gnd cell_6t
Xbit_r127_c78 bl[78] br[78] wl[127] vdd gnd cell_6t
Xbit_r0_c79 bl[79] br[79] wl[0] vdd gnd cell_6t
Xbit_r1_c79 bl[79] br[79] wl[1] vdd gnd cell_6t
Xbit_r2_c79 bl[79] br[79] wl[2] vdd gnd cell_6t
Xbit_r3_c79 bl[79] br[79] wl[3] vdd gnd cell_6t
Xbit_r4_c79 bl[79] br[79] wl[4] vdd gnd cell_6t
Xbit_r5_c79 bl[79] br[79] wl[5] vdd gnd cell_6t
Xbit_r6_c79 bl[79] br[79] wl[6] vdd gnd cell_6t
Xbit_r7_c79 bl[79] br[79] wl[7] vdd gnd cell_6t
Xbit_r8_c79 bl[79] br[79] wl[8] vdd gnd cell_6t
Xbit_r9_c79 bl[79] br[79] wl[9] vdd gnd cell_6t
Xbit_r10_c79 bl[79] br[79] wl[10] vdd gnd cell_6t
Xbit_r11_c79 bl[79] br[79] wl[11] vdd gnd cell_6t
Xbit_r12_c79 bl[79] br[79] wl[12] vdd gnd cell_6t
Xbit_r13_c79 bl[79] br[79] wl[13] vdd gnd cell_6t
Xbit_r14_c79 bl[79] br[79] wl[14] vdd gnd cell_6t
Xbit_r15_c79 bl[79] br[79] wl[15] vdd gnd cell_6t
Xbit_r16_c79 bl[79] br[79] wl[16] vdd gnd cell_6t
Xbit_r17_c79 bl[79] br[79] wl[17] vdd gnd cell_6t
Xbit_r18_c79 bl[79] br[79] wl[18] vdd gnd cell_6t
Xbit_r19_c79 bl[79] br[79] wl[19] vdd gnd cell_6t
Xbit_r20_c79 bl[79] br[79] wl[20] vdd gnd cell_6t
Xbit_r21_c79 bl[79] br[79] wl[21] vdd gnd cell_6t
Xbit_r22_c79 bl[79] br[79] wl[22] vdd gnd cell_6t
Xbit_r23_c79 bl[79] br[79] wl[23] vdd gnd cell_6t
Xbit_r24_c79 bl[79] br[79] wl[24] vdd gnd cell_6t
Xbit_r25_c79 bl[79] br[79] wl[25] vdd gnd cell_6t
Xbit_r26_c79 bl[79] br[79] wl[26] vdd gnd cell_6t
Xbit_r27_c79 bl[79] br[79] wl[27] vdd gnd cell_6t
Xbit_r28_c79 bl[79] br[79] wl[28] vdd gnd cell_6t
Xbit_r29_c79 bl[79] br[79] wl[29] vdd gnd cell_6t
Xbit_r30_c79 bl[79] br[79] wl[30] vdd gnd cell_6t
Xbit_r31_c79 bl[79] br[79] wl[31] vdd gnd cell_6t
Xbit_r32_c79 bl[79] br[79] wl[32] vdd gnd cell_6t
Xbit_r33_c79 bl[79] br[79] wl[33] vdd gnd cell_6t
Xbit_r34_c79 bl[79] br[79] wl[34] vdd gnd cell_6t
Xbit_r35_c79 bl[79] br[79] wl[35] vdd gnd cell_6t
Xbit_r36_c79 bl[79] br[79] wl[36] vdd gnd cell_6t
Xbit_r37_c79 bl[79] br[79] wl[37] vdd gnd cell_6t
Xbit_r38_c79 bl[79] br[79] wl[38] vdd gnd cell_6t
Xbit_r39_c79 bl[79] br[79] wl[39] vdd gnd cell_6t
Xbit_r40_c79 bl[79] br[79] wl[40] vdd gnd cell_6t
Xbit_r41_c79 bl[79] br[79] wl[41] vdd gnd cell_6t
Xbit_r42_c79 bl[79] br[79] wl[42] vdd gnd cell_6t
Xbit_r43_c79 bl[79] br[79] wl[43] vdd gnd cell_6t
Xbit_r44_c79 bl[79] br[79] wl[44] vdd gnd cell_6t
Xbit_r45_c79 bl[79] br[79] wl[45] vdd gnd cell_6t
Xbit_r46_c79 bl[79] br[79] wl[46] vdd gnd cell_6t
Xbit_r47_c79 bl[79] br[79] wl[47] vdd gnd cell_6t
Xbit_r48_c79 bl[79] br[79] wl[48] vdd gnd cell_6t
Xbit_r49_c79 bl[79] br[79] wl[49] vdd gnd cell_6t
Xbit_r50_c79 bl[79] br[79] wl[50] vdd gnd cell_6t
Xbit_r51_c79 bl[79] br[79] wl[51] vdd gnd cell_6t
Xbit_r52_c79 bl[79] br[79] wl[52] vdd gnd cell_6t
Xbit_r53_c79 bl[79] br[79] wl[53] vdd gnd cell_6t
Xbit_r54_c79 bl[79] br[79] wl[54] vdd gnd cell_6t
Xbit_r55_c79 bl[79] br[79] wl[55] vdd gnd cell_6t
Xbit_r56_c79 bl[79] br[79] wl[56] vdd gnd cell_6t
Xbit_r57_c79 bl[79] br[79] wl[57] vdd gnd cell_6t
Xbit_r58_c79 bl[79] br[79] wl[58] vdd gnd cell_6t
Xbit_r59_c79 bl[79] br[79] wl[59] vdd gnd cell_6t
Xbit_r60_c79 bl[79] br[79] wl[60] vdd gnd cell_6t
Xbit_r61_c79 bl[79] br[79] wl[61] vdd gnd cell_6t
Xbit_r62_c79 bl[79] br[79] wl[62] vdd gnd cell_6t
Xbit_r63_c79 bl[79] br[79] wl[63] vdd gnd cell_6t
Xbit_r64_c79 bl[79] br[79] wl[64] vdd gnd cell_6t
Xbit_r65_c79 bl[79] br[79] wl[65] vdd gnd cell_6t
Xbit_r66_c79 bl[79] br[79] wl[66] vdd gnd cell_6t
Xbit_r67_c79 bl[79] br[79] wl[67] vdd gnd cell_6t
Xbit_r68_c79 bl[79] br[79] wl[68] vdd gnd cell_6t
Xbit_r69_c79 bl[79] br[79] wl[69] vdd gnd cell_6t
Xbit_r70_c79 bl[79] br[79] wl[70] vdd gnd cell_6t
Xbit_r71_c79 bl[79] br[79] wl[71] vdd gnd cell_6t
Xbit_r72_c79 bl[79] br[79] wl[72] vdd gnd cell_6t
Xbit_r73_c79 bl[79] br[79] wl[73] vdd gnd cell_6t
Xbit_r74_c79 bl[79] br[79] wl[74] vdd gnd cell_6t
Xbit_r75_c79 bl[79] br[79] wl[75] vdd gnd cell_6t
Xbit_r76_c79 bl[79] br[79] wl[76] vdd gnd cell_6t
Xbit_r77_c79 bl[79] br[79] wl[77] vdd gnd cell_6t
Xbit_r78_c79 bl[79] br[79] wl[78] vdd gnd cell_6t
Xbit_r79_c79 bl[79] br[79] wl[79] vdd gnd cell_6t
Xbit_r80_c79 bl[79] br[79] wl[80] vdd gnd cell_6t
Xbit_r81_c79 bl[79] br[79] wl[81] vdd gnd cell_6t
Xbit_r82_c79 bl[79] br[79] wl[82] vdd gnd cell_6t
Xbit_r83_c79 bl[79] br[79] wl[83] vdd gnd cell_6t
Xbit_r84_c79 bl[79] br[79] wl[84] vdd gnd cell_6t
Xbit_r85_c79 bl[79] br[79] wl[85] vdd gnd cell_6t
Xbit_r86_c79 bl[79] br[79] wl[86] vdd gnd cell_6t
Xbit_r87_c79 bl[79] br[79] wl[87] vdd gnd cell_6t
Xbit_r88_c79 bl[79] br[79] wl[88] vdd gnd cell_6t
Xbit_r89_c79 bl[79] br[79] wl[89] vdd gnd cell_6t
Xbit_r90_c79 bl[79] br[79] wl[90] vdd gnd cell_6t
Xbit_r91_c79 bl[79] br[79] wl[91] vdd gnd cell_6t
Xbit_r92_c79 bl[79] br[79] wl[92] vdd gnd cell_6t
Xbit_r93_c79 bl[79] br[79] wl[93] vdd gnd cell_6t
Xbit_r94_c79 bl[79] br[79] wl[94] vdd gnd cell_6t
Xbit_r95_c79 bl[79] br[79] wl[95] vdd gnd cell_6t
Xbit_r96_c79 bl[79] br[79] wl[96] vdd gnd cell_6t
Xbit_r97_c79 bl[79] br[79] wl[97] vdd gnd cell_6t
Xbit_r98_c79 bl[79] br[79] wl[98] vdd gnd cell_6t
Xbit_r99_c79 bl[79] br[79] wl[99] vdd gnd cell_6t
Xbit_r100_c79 bl[79] br[79] wl[100] vdd gnd cell_6t
Xbit_r101_c79 bl[79] br[79] wl[101] vdd gnd cell_6t
Xbit_r102_c79 bl[79] br[79] wl[102] vdd gnd cell_6t
Xbit_r103_c79 bl[79] br[79] wl[103] vdd gnd cell_6t
Xbit_r104_c79 bl[79] br[79] wl[104] vdd gnd cell_6t
Xbit_r105_c79 bl[79] br[79] wl[105] vdd gnd cell_6t
Xbit_r106_c79 bl[79] br[79] wl[106] vdd gnd cell_6t
Xbit_r107_c79 bl[79] br[79] wl[107] vdd gnd cell_6t
Xbit_r108_c79 bl[79] br[79] wl[108] vdd gnd cell_6t
Xbit_r109_c79 bl[79] br[79] wl[109] vdd gnd cell_6t
Xbit_r110_c79 bl[79] br[79] wl[110] vdd gnd cell_6t
Xbit_r111_c79 bl[79] br[79] wl[111] vdd gnd cell_6t
Xbit_r112_c79 bl[79] br[79] wl[112] vdd gnd cell_6t
Xbit_r113_c79 bl[79] br[79] wl[113] vdd gnd cell_6t
Xbit_r114_c79 bl[79] br[79] wl[114] vdd gnd cell_6t
Xbit_r115_c79 bl[79] br[79] wl[115] vdd gnd cell_6t
Xbit_r116_c79 bl[79] br[79] wl[116] vdd gnd cell_6t
Xbit_r117_c79 bl[79] br[79] wl[117] vdd gnd cell_6t
Xbit_r118_c79 bl[79] br[79] wl[118] vdd gnd cell_6t
Xbit_r119_c79 bl[79] br[79] wl[119] vdd gnd cell_6t
Xbit_r120_c79 bl[79] br[79] wl[120] vdd gnd cell_6t
Xbit_r121_c79 bl[79] br[79] wl[121] vdd gnd cell_6t
Xbit_r122_c79 bl[79] br[79] wl[122] vdd gnd cell_6t
Xbit_r123_c79 bl[79] br[79] wl[123] vdd gnd cell_6t
Xbit_r124_c79 bl[79] br[79] wl[124] vdd gnd cell_6t
Xbit_r125_c79 bl[79] br[79] wl[125] vdd gnd cell_6t
Xbit_r126_c79 bl[79] br[79] wl[126] vdd gnd cell_6t
Xbit_r127_c79 bl[79] br[79] wl[127] vdd gnd cell_6t
Xbit_r0_c80 bl[80] br[80] wl[0] vdd gnd cell_6t
Xbit_r1_c80 bl[80] br[80] wl[1] vdd gnd cell_6t
Xbit_r2_c80 bl[80] br[80] wl[2] vdd gnd cell_6t
Xbit_r3_c80 bl[80] br[80] wl[3] vdd gnd cell_6t
Xbit_r4_c80 bl[80] br[80] wl[4] vdd gnd cell_6t
Xbit_r5_c80 bl[80] br[80] wl[5] vdd gnd cell_6t
Xbit_r6_c80 bl[80] br[80] wl[6] vdd gnd cell_6t
Xbit_r7_c80 bl[80] br[80] wl[7] vdd gnd cell_6t
Xbit_r8_c80 bl[80] br[80] wl[8] vdd gnd cell_6t
Xbit_r9_c80 bl[80] br[80] wl[9] vdd gnd cell_6t
Xbit_r10_c80 bl[80] br[80] wl[10] vdd gnd cell_6t
Xbit_r11_c80 bl[80] br[80] wl[11] vdd gnd cell_6t
Xbit_r12_c80 bl[80] br[80] wl[12] vdd gnd cell_6t
Xbit_r13_c80 bl[80] br[80] wl[13] vdd gnd cell_6t
Xbit_r14_c80 bl[80] br[80] wl[14] vdd gnd cell_6t
Xbit_r15_c80 bl[80] br[80] wl[15] vdd gnd cell_6t
Xbit_r16_c80 bl[80] br[80] wl[16] vdd gnd cell_6t
Xbit_r17_c80 bl[80] br[80] wl[17] vdd gnd cell_6t
Xbit_r18_c80 bl[80] br[80] wl[18] vdd gnd cell_6t
Xbit_r19_c80 bl[80] br[80] wl[19] vdd gnd cell_6t
Xbit_r20_c80 bl[80] br[80] wl[20] vdd gnd cell_6t
Xbit_r21_c80 bl[80] br[80] wl[21] vdd gnd cell_6t
Xbit_r22_c80 bl[80] br[80] wl[22] vdd gnd cell_6t
Xbit_r23_c80 bl[80] br[80] wl[23] vdd gnd cell_6t
Xbit_r24_c80 bl[80] br[80] wl[24] vdd gnd cell_6t
Xbit_r25_c80 bl[80] br[80] wl[25] vdd gnd cell_6t
Xbit_r26_c80 bl[80] br[80] wl[26] vdd gnd cell_6t
Xbit_r27_c80 bl[80] br[80] wl[27] vdd gnd cell_6t
Xbit_r28_c80 bl[80] br[80] wl[28] vdd gnd cell_6t
Xbit_r29_c80 bl[80] br[80] wl[29] vdd gnd cell_6t
Xbit_r30_c80 bl[80] br[80] wl[30] vdd gnd cell_6t
Xbit_r31_c80 bl[80] br[80] wl[31] vdd gnd cell_6t
Xbit_r32_c80 bl[80] br[80] wl[32] vdd gnd cell_6t
Xbit_r33_c80 bl[80] br[80] wl[33] vdd gnd cell_6t
Xbit_r34_c80 bl[80] br[80] wl[34] vdd gnd cell_6t
Xbit_r35_c80 bl[80] br[80] wl[35] vdd gnd cell_6t
Xbit_r36_c80 bl[80] br[80] wl[36] vdd gnd cell_6t
Xbit_r37_c80 bl[80] br[80] wl[37] vdd gnd cell_6t
Xbit_r38_c80 bl[80] br[80] wl[38] vdd gnd cell_6t
Xbit_r39_c80 bl[80] br[80] wl[39] vdd gnd cell_6t
Xbit_r40_c80 bl[80] br[80] wl[40] vdd gnd cell_6t
Xbit_r41_c80 bl[80] br[80] wl[41] vdd gnd cell_6t
Xbit_r42_c80 bl[80] br[80] wl[42] vdd gnd cell_6t
Xbit_r43_c80 bl[80] br[80] wl[43] vdd gnd cell_6t
Xbit_r44_c80 bl[80] br[80] wl[44] vdd gnd cell_6t
Xbit_r45_c80 bl[80] br[80] wl[45] vdd gnd cell_6t
Xbit_r46_c80 bl[80] br[80] wl[46] vdd gnd cell_6t
Xbit_r47_c80 bl[80] br[80] wl[47] vdd gnd cell_6t
Xbit_r48_c80 bl[80] br[80] wl[48] vdd gnd cell_6t
Xbit_r49_c80 bl[80] br[80] wl[49] vdd gnd cell_6t
Xbit_r50_c80 bl[80] br[80] wl[50] vdd gnd cell_6t
Xbit_r51_c80 bl[80] br[80] wl[51] vdd gnd cell_6t
Xbit_r52_c80 bl[80] br[80] wl[52] vdd gnd cell_6t
Xbit_r53_c80 bl[80] br[80] wl[53] vdd gnd cell_6t
Xbit_r54_c80 bl[80] br[80] wl[54] vdd gnd cell_6t
Xbit_r55_c80 bl[80] br[80] wl[55] vdd gnd cell_6t
Xbit_r56_c80 bl[80] br[80] wl[56] vdd gnd cell_6t
Xbit_r57_c80 bl[80] br[80] wl[57] vdd gnd cell_6t
Xbit_r58_c80 bl[80] br[80] wl[58] vdd gnd cell_6t
Xbit_r59_c80 bl[80] br[80] wl[59] vdd gnd cell_6t
Xbit_r60_c80 bl[80] br[80] wl[60] vdd gnd cell_6t
Xbit_r61_c80 bl[80] br[80] wl[61] vdd gnd cell_6t
Xbit_r62_c80 bl[80] br[80] wl[62] vdd gnd cell_6t
Xbit_r63_c80 bl[80] br[80] wl[63] vdd gnd cell_6t
Xbit_r64_c80 bl[80] br[80] wl[64] vdd gnd cell_6t
Xbit_r65_c80 bl[80] br[80] wl[65] vdd gnd cell_6t
Xbit_r66_c80 bl[80] br[80] wl[66] vdd gnd cell_6t
Xbit_r67_c80 bl[80] br[80] wl[67] vdd gnd cell_6t
Xbit_r68_c80 bl[80] br[80] wl[68] vdd gnd cell_6t
Xbit_r69_c80 bl[80] br[80] wl[69] vdd gnd cell_6t
Xbit_r70_c80 bl[80] br[80] wl[70] vdd gnd cell_6t
Xbit_r71_c80 bl[80] br[80] wl[71] vdd gnd cell_6t
Xbit_r72_c80 bl[80] br[80] wl[72] vdd gnd cell_6t
Xbit_r73_c80 bl[80] br[80] wl[73] vdd gnd cell_6t
Xbit_r74_c80 bl[80] br[80] wl[74] vdd gnd cell_6t
Xbit_r75_c80 bl[80] br[80] wl[75] vdd gnd cell_6t
Xbit_r76_c80 bl[80] br[80] wl[76] vdd gnd cell_6t
Xbit_r77_c80 bl[80] br[80] wl[77] vdd gnd cell_6t
Xbit_r78_c80 bl[80] br[80] wl[78] vdd gnd cell_6t
Xbit_r79_c80 bl[80] br[80] wl[79] vdd gnd cell_6t
Xbit_r80_c80 bl[80] br[80] wl[80] vdd gnd cell_6t
Xbit_r81_c80 bl[80] br[80] wl[81] vdd gnd cell_6t
Xbit_r82_c80 bl[80] br[80] wl[82] vdd gnd cell_6t
Xbit_r83_c80 bl[80] br[80] wl[83] vdd gnd cell_6t
Xbit_r84_c80 bl[80] br[80] wl[84] vdd gnd cell_6t
Xbit_r85_c80 bl[80] br[80] wl[85] vdd gnd cell_6t
Xbit_r86_c80 bl[80] br[80] wl[86] vdd gnd cell_6t
Xbit_r87_c80 bl[80] br[80] wl[87] vdd gnd cell_6t
Xbit_r88_c80 bl[80] br[80] wl[88] vdd gnd cell_6t
Xbit_r89_c80 bl[80] br[80] wl[89] vdd gnd cell_6t
Xbit_r90_c80 bl[80] br[80] wl[90] vdd gnd cell_6t
Xbit_r91_c80 bl[80] br[80] wl[91] vdd gnd cell_6t
Xbit_r92_c80 bl[80] br[80] wl[92] vdd gnd cell_6t
Xbit_r93_c80 bl[80] br[80] wl[93] vdd gnd cell_6t
Xbit_r94_c80 bl[80] br[80] wl[94] vdd gnd cell_6t
Xbit_r95_c80 bl[80] br[80] wl[95] vdd gnd cell_6t
Xbit_r96_c80 bl[80] br[80] wl[96] vdd gnd cell_6t
Xbit_r97_c80 bl[80] br[80] wl[97] vdd gnd cell_6t
Xbit_r98_c80 bl[80] br[80] wl[98] vdd gnd cell_6t
Xbit_r99_c80 bl[80] br[80] wl[99] vdd gnd cell_6t
Xbit_r100_c80 bl[80] br[80] wl[100] vdd gnd cell_6t
Xbit_r101_c80 bl[80] br[80] wl[101] vdd gnd cell_6t
Xbit_r102_c80 bl[80] br[80] wl[102] vdd gnd cell_6t
Xbit_r103_c80 bl[80] br[80] wl[103] vdd gnd cell_6t
Xbit_r104_c80 bl[80] br[80] wl[104] vdd gnd cell_6t
Xbit_r105_c80 bl[80] br[80] wl[105] vdd gnd cell_6t
Xbit_r106_c80 bl[80] br[80] wl[106] vdd gnd cell_6t
Xbit_r107_c80 bl[80] br[80] wl[107] vdd gnd cell_6t
Xbit_r108_c80 bl[80] br[80] wl[108] vdd gnd cell_6t
Xbit_r109_c80 bl[80] br[80] wl[109] vdd gnd cell_6t
Xbit_r110_c80 bl[80] br[80] wl[110] vdd gnd cell_6t
Xbit_r111_c80 bl[80] br[80] wl[111] vdd gnd cell_6t
Xbit_r112_c80 bl[80] br[80] wl[112] vdd gnd cell_6t
Xbit_r113_c80 bl[80] br[80] wl[113] vdd gnd cell_6t
Xbit_r114_c80 bl[80] br[80] wl[114] vdd gnd cell_6t
Xbit_r115_c80 bl[80] br[80] wl[115] vdd gnd cell_6t
Xbit_r116_c80 bl[80] br[80] wl[116] vdd gnd cell_6t
Xbit_r117_c80 bl[80] br[80] wl[117] vdd gnd cell_6t
Xbit_r118_c80 bl[80] br[80] wl[118] vdd gnd cell_6t
Xbit_r119_c80 bl[80] br[80] wl[119] vdd gnd cell_6t
Xbit_r120_c80 bl[80] br[80] wl[120] vdd gnd cell_6t
Xbit_r121_c80 bl[80] br[80] wl[121] vdd gnd cell_6t
Xbit_r122_c80 bl[80] br[80] wl[122] vdd gnd cell_6t
Xbit_r123_c80 bl[80] br[80] wl[123] vdd gnd cell_6t
Xbit_r124_c80 bl[80] br[80] wl[124] vdd gnd cell_6t
Xbit_r125_c80 bl[80] br[80] wl[125] vdd gnd cell_6t
Xbit_r126_c80 bl[80] br[80] wl[126] vdd gnd cell_6t
Xbit_r127_c80 bl[80] br[80] wl[127] vdd gnd cell_6t
Xbit_r0_c81 bl[81] br[81] wl[0] vdd gnd cell_6t
Xbit_r1_c81 bl[81] br[81] wl[1] vdd gnd cell_6t
Xbit_r2_c81 bl[81] br[81] wl[2] vdd gnd cell_6t
Xbit_r3_c81 bl[81] br[81] wl[3] vdd gnd cell_6t
Xbit_r4_c81 bl[81] br[81] wl[4] vdd gnd cell_6t
Xbit_r5_c81 bl[81] br[81] wl[5] vdd gnd cell_6t
Xbit_r6_c81 bl[81] br[81] wl[6] vdd gnd cell_6t
Xbit_r7_c81 bl[81] br[81] wl[7] vdd gnd cell_6t
Xbit_r8_c81 bl[81] br[81] wl[8] vdd gnd cell_6t
Xbit_r9_c81 bl[81] br[81] wl[9] vdd gnd cell_6t
Xbit_r10_c81 bl[81] br[81] wl[10] vdd gnd cell_6t
Xbit_r11_c81 bl[81] br[81] wl[11] vdd gnd cell_6t
Xbit_r12_c81 bl[81] br[81] wl[12] vdd gnd cell_6t
Xbit_r13_c81 bl[81] br[81] wl[13] vdd gnd cell_6t
Xbit_r14_c81 bl[81] br[81] wl[14] vdd gnd cell_6t
Xbit_r15_c81 bl[81] br[81] wl[15] vdd gnd cell_6t
Xbit_r16_c81 bl[81] br[81] wl[16] vdd gnd cell_6t
Xbit_r17_c81 bl[81] br[81] wl[17] vdd gnd cell_6t
Xbit_r18_c81 bl[81] br[81] wl[18] vdd gnd cell_6t
Xbit_r19_c81 bl[81] br[81] wl[19] vdd gnd cell_6t
Xbit_r20_c81 bl[81] br[81] wl[20] vdd gnd cell_6t
Xbit_r21_c81 bl[81] br[81] wl[21] vdd gnd cell_6t
Xbit_r22_c81 bl[81] br[81] wl[22] vdd gnd cell_6t
Xbit_r23_c81 bl[81] br[81] wl[23] vdd gnd cell_6t
Xbit_r24_c81 bl[81] br[81] wl[24] vdd gnd cell_6t
Xbit_r25_c81 bl[81] br[81] wl[25] vdd gnd cell_6t
Xbit_r26_c81 bl[81] br[81] wl[26] vdd gnd cell_6t
Xbit_r27_c81 bl[81] br[81] wl[27] vdd gnd cell_6t
Xbit_r28_c81 bl[81] br[81] wl[28] vdd gnd cell_6t
Xbit_r29_c81 bl[81] br[81] wl[29] vdd gnd cell_6t
Xbit_r30_c81 bl[81] br[81] wl[30] vdd gnd cell_6t
Xbit_r31_c81 bl[81] br[81] wl[31] vdd gnd cell_6t
Xbit_r32_c81 bl[81] br[81] wl[32] vdd gnd cell_6t
Xbit_r33_c81 bl[81] br[81] wl[33] vdd gnd cell_6t
Xbit_r34_c81 bl[81] br[81] wl[34] vdd gnd cell_6t
Xbit_r35_c81 bl[81] br[81] wl[35] vdd gnd cell_6t
Xbit_r36_c81 bl[81] br[81] wl[36] vdd gnd cell_6t
Xbit_r37_c81 bl[81] br[81] wl[37] vdd gnd cell_6t
Xbit_r38_c81 bl[81] br[81] wl[38] vdd gnd cell_6t
Xbit_r39_c81 bl[81] br[81] wl[39] vdd gnd cell_6t
Xbit_r40_c81 bl[81] br[81] wl[40] vdd gnd cell_6t
Xbit_r41_c81 bl[81] br[81] wl[41] vdd gnd cell_6t
Xbit_r42_c81 bl[81] br[81] wl[42] vdd gnd cell_6t
Xbit_r43_c81 bl[81] br[81] wl[43] vdd gnd cell_6t
Xbit_r44_c81 bl[81] br[81] wl[44] vdd gnd cell_6t
Xbit_r45_c81 bl[81] br[81] wl[45] vdd gnd cell_6t
Xbit_r46_c81 bl[81] br[81] wl[46] vdd gnd cell_6t
Xbit_r47_c81 bl[81] br[81] wl[47] vdd gnd cell_6t
Xbit_r48_c81 bl[81] br[81] wl[48] vdd gnd cell_6t
Xbit_r49_c81 bl[81] br[81] wl[49] vdd gnd cell_6t
Xbit_r50_c81 bl[81] br[81] wl[50] vdd gnd cell_6t
Xbit_r51_c81 bl[81] br[81] wl[51] vdd gnd cell_6t
Xbit_r52_c81 bl[81] br[81] wl[52] vdd gnd cell_6t
Xbit_r53_c81 bl[81] br[81] wl[53] vdd gnd cell_6t
Xbit_r54_c81 bl[81] br[81] wl[54] vdd gnd cell_6t
Xbit_r55_c81 bl[81] br[81] wl[55] vdd gnd cell_6t
Xbit_r56_c81 bl[81] br[81] wl[56] vdd gnd cell_6t
Xbit_r57_c81 bl[81] br[81] wl[57] vdd gnd cell_6t
Xbit_r58_c81 bl[81] br[81] wl[58] vdd gnd cell_6t
Xbit_r59_c81 bl[81] br[81] wl[59] vdd gnd cell_6t
Xbit_r60_c81 bl[81] br[81] wl[60] vdd gnd cell_6t
Xbit_r61_c81 bl[81] br[81] wl[61] vdd gnd cell_6t
Xbit_r62_c81 bl[81] br[81] wl[62] vdd gnd cell_6t
Xbit_r63_c81 bl[81] br[81] wl[63] vdd gnd cell_6t
Xbit_r64_c81 bl[81] br[81] wl[64] vdd gnd cell_6t
Xbit_r65_c81 bl[81] br[81] wl[65] vdd gnd cell_6t
Xbit_r66_c81 bl[81] br[81] wl[66] vdd gnd cell_6t
Xbit_r67_c81 bl[81] br[81] wl[67] vdd gnd cell_6t
Xbit_r68_c81 bl[81] br[81] wl[68] vdd gnd cell_6t
Xbit_r69_c81 bl[81] br[81] wl[69] vdd gnd cell_6t
Xbit_r70_c81 bl[81] br[81] wl[70] vdd gnd cell_6t
Xbit_r71_c81 bl[81] br[81] wl[71] vdd gnd cell_6t
Xbit_r72_c81 bl[81] br[81] wl[72] vdd gnd cell_6t
Xbit_r73_c81 bl[81] br[81] wl[73] vdd gnd cell_6t
Xbit_r74_c81 bl[81] br[81] wl[74] vdd gnd cell_6t
Xbit_r75_c81 bl[81] br[81] wl[75] vdd gnd cell_6t
Xbit_r76_c81 bl[81] br[81] wl[76] vdd gnd cell_6t
Xbit_r77_c81 bl[81] br[81] wl[77] vdd gnd cell_6t
Xbit_r78_c81 bl[81] br[81] wl[78] vdd gnd cell_6t
Xbit_r79_c81 bl[81] br[81] wl[79] vdd gnd cell_6t
Xbit_r80_c81 bl[81] br[81] wl[80] vdd gnd cell_6t
Xbit_r81_c81 bl[81] br[81] wl[81] vdd gnd cell_6t
Xbit_r82_c81 bl[81] br[81] wl[82] vdd gnd cell_6t
Xbit_r83_c81 bl[81] br[81] wl[83] vdd gnd cell_6t
Xbit_r84_c81 bl[81] br[81] wl[84] vdd gnd cell_6t
Xbit_r85_c81 bl[81] br[81] wl[85] vdd gnd cell_6t
Xbit_r86_c81 bl[81] br[81] wl[86] vdd gnd cell_6t
Xbit_r87_c81 bl[81] br[81] wl[87] vdd gnd cell_6t
Xbit_r88_c81 bl[81] br[81] wl[88] vdd gnd cell_6t
Xbit_r89_c81 bl[81] br[81] wl[89] vdd gnd cell_6t
Xbit_r90_c81 bl[81] br[81] wl[90] vdd gnd cell_6t
Xbit_r91_c81 bl[81] br[81] wl[91] vdd gnd cell_6t
Xbit_r92_c81 bl[81] br[81] wl[92] vdd gnd cell_6t
Xbit_r93_c81 bl[81] br[81] wl[93] vdd gnd cell_6t
Xbit_r94_c81 bl[81] br[81] wl[94] vdd gnd cell_6t
Xbit_r95_c81 bl[81] br[81] wl[95] vdd gnd cell_6t
Xbit_r96_c81 bl[81] br[81] wl[96] vdd gnd cell_6t
Xbit_r97_c81 bl[81] br[81] wl[97] vdd gnd cell_6t
Xbit_r98_c81 bl[81] br[81] wl[98] vdd gnd cell_6t
Xbit_r99_c81 bl[81] br[81] wl[99] vdd gnd cell_6t
Xbit_r100_c81 bl[81] br[81] wl[100] vdd gnd cell_6t
Xbit_r101_c81 bl[81] br[81] wl[101] vdd gnd cell_6t
Xbit_r102_c81 bl[81] br[81] wl[102] vdd gnd cell_6t
Xbit_r103_c81 bl[81] br[81] wl[103] vdd gnd cell_6t
Xbit_r104_c81 bl[81] br[81] wl[104] vdd gnd cell_6t
Xbit_r105_c81 bl[81] br[81] wl[105] vdd gnd cell_6t
Xbit_r106_c81 bl[81] br[81] wl[106] vdd gnd cell_6t
Xbit_r107_c81 bl[81] br[81] wl[107] vdd gnd cell_6t
Xbit_r108_c81 bl[81] br[81] wl[108] vdd gnd cell_6t
Xbit_r109_c81 bl[81] br[81] wl[109] vdd gnd cell_6t
Xbit_r110_c81 bl[81] br[81] wl[110] vdd gnd cell_6t
Xbit_r111_c81 bl[81] br[81] wl[111] vdd gnd cell_6t
Xbit_r112_c81 bl[81] br[81] wl[112] vdd gnd cell_6t
Xbit_r113_c81 bl[81] br[81] wl[113] vdd gnd cell_6t
Xbit_r114_c81 bl[81] br[81] wl[114] vdd gnd cell_6t
Xbit_r115_c81 bl[81] br[81] wl[115] vdd gnd cell_6t
Xbit_r116_c81 bl[81] br[81] wl[116] vdd gnd cell_6t
Xbit_r117_c81 bl[81] br[81] wl[117] vdd gnd cell_6t
Xbit_r118_c81 bl[81] br[81] wl[118] vdd gnd cell_6t
Xbit_r119_c81 bl[81] br[81] wl[119] vdd gnd cell_6t
Xbit_r120_c81 bl[81] br[81] wl[120] vdd gnd cell_6t
Xbit_r121_c81 bl[81] br[81] wl[121] vdd gnd cell_6t
Xbit_r122_c81 bl[81] br[81] wl[122] vdd gnd cell_6t
Xbit_r123_c81 bl[81] br[81] wl[123] vdd gnd cell_6t
Xbit_r124_c81 bl[81] br[81] wl[124] vdd gnd cell_6t
Xbit_r125_c81 bl[81] br[81] wl[125] vdd gnd cell_6t
Xbit_r126_c81 bl[81] br[81] wl[126] vdd gnd cell_6t
Xbit_r127_c81 bl[81] br[81] wl[127] vdd gnd cell_6t
Xbit_r0_c82 bl[82] br[82] wl[0] vdd gnd cell_6t
Xbit_r1_c82 bl[82] br[82] wl[1] vdd gnd cell_6t
Xbit_r2_c82 bl[82] br[82] wl[2] vdd gnd cell_6t
Xbit_r3_c82 bl[82] br[82] wl[3] vdd gnd cell_6t
Xbit_r4_c82 bl[82] br[82] wl[4] vdd gnd cell_6t
Xbit_r5_c82 bl[82] br[82] wl[5] vdd gnd cell_6t
Xbit_r6_c82 bl[82] br[82] wl[6] vdd gnd cell_6t
Xbit_r7_c82 bl[82] br[82] wl[7] vdd gnd cell_6t
Xbit_r8_c82 bl[82] br[82] wl[8] vdd gnd cell_6t
Xbit_r9_c82 bl[82] br[82] wl[9] vdd gnd cell_6t
Xbit_r10_c82 bl[82] br[82] wl[10] vdd gnd cell_6t
Xbit_r11_c82 bl[82] br[82] wl[11] vdd gnd cell_6t
Xbit_r12_c82 bl[82] br[82] wl[12] vdd gnd cell_6t
Xbit_r13_c82 bl[82] br[82] wl[13] vdd gnd cell_6t
Xbit_r14_c82 bl[82] br[82] wl[14] vdd gnd cell_6t
Xbit_r15_c82 bl[82] br[82] wl[15] vdd gnd cell_6t
Xbit_r16_c82 bl[82] br[82] wl[16] vdd gnd cell_6t
Xbit_r17_c82 bl[82] br[82] wl[17] vdd gnd cell_6t
Xbit_r18_c82 bl[82] br[82] wl[18] vdd gnd cell_6t
Xbit_r19_c82 bl[82] br[82] wl[19] vdd gnd cell_6t
Xbit_r20_c82 bl[82] br[82] wl[20] vdd gnd cell_6t
Xbit_r21_c82 bl[82] br[82] wl[21] vdd gnd cell_6t
Xbit_r22_c82 bl[82] br[82] wl[22] vdd gnd cell_6t
Xbit_r23_c82 bl[82] br[82] wl[23] vdd gnd cell_6t
Xbit_r24_c82 bl[82] br[82] wl[24] vdd gnd cell_6t
Xbit_r25_c82 bl[82] br[82] wl[25] vdd gnd cell_6t
Xbit_r26_c82 bl[82] br[82] wl[26] vdd gnd cell_6t
Xbit_r27_c82 bl[82] br[82] wl[27] vdd gnd cell_6t
Xbit_r28_c82 bl[82] br[82] wl[28] vdd gnd cell_6t
Xbit_r29_c82 bl[82] br[82] wl[29] vdd gnd cell_6t
Xbit_r30_c82 bl[82] br[82] wl[30] vdd gnd cell_6t
Xbit_r31_c82 bl[82] br[82] wl[31] vdd gnd cell_6t
Xbit_r32_c82 bl[82] br[82] wl[32] vdd gnd cell_6t
Xbit_r33_c82 bl[82] br[82] wl[33] vdd gnd cell_6t
Xbit_r34_c82 bl[82] br[82] wl[34] vdd gnd cell_6t
Xbit_r35_c82 bl[82] br[82] wl[35] vdd gnd cell_6t
Xbit_r36_c82 bl[82] br[82] wl[36] vdd gnd cell_6t
Xbit_r37_c82 bl[82] br[82] wl[37] vdd gnd cell_6t
Xbit_r38_c82 bl[82] br[82] wl[38] vdd gnd cell_6t
Xbit_r39_c82 bl[82] br[82] wl[39] vdd gnd cell_6t
Xbit_r40_c82 bl[82] br[82] wl[40] vdd gnd cell_6t
Xbit_r41_c82 bl[82] br[82] wl[41] vdd gnd cell_6t
Xbit_r42_c82 bl[82] br[82] wl[42] vdd gnd cell_6t
Xbit_r43_c82 bl[82] br[82] wl[43] vdd gnd cell_6t
Xbit_r44_c82 bl[82] br[82] wl[44] vdd gnd cell_6t
Xbit_r45_c82 bl[82] br[82] wl[45] vdd gnd cell_6t
Xbit_r46_c82 bl[82] br[82] wl[46] vdd gnd cell_6t
Xbit_r47_c82 bl[82] br[82] wl[47] vdd gnd cell_6t
Xbit_r48_c82 bl[82] br[82] wl[48] vdd gnd cell_6t
Xbit_r49_c82 bl[82] br[82] wl[49] vdd gnd cell_6t
Xbit_r50_c82 bl[82] br[82] wl[50] vdd gnd cell_6t
Xbit_r51_c82 bl[82] br[82] wl[51] vdd gnd cell_6t
Xbit_r52_c82 bl[82] br[82] wl[52] vdd gnd cell_6t
Xbit_r53_c82 bl[82] br[82] wl[53] vdd gnd cell_6t
Xbit_r54_c82 bl[82] br[82] wl[54] vdd gnd cell_6t
Xbit_r55_c82 bl[82] br[82] wl[55] vdd gnd cell_6t
Xbit_r56_c82 bl[82] br[82] wl[56] vdd gnd cell_6t
Xbit_r57_c82 bl[82] br[82] wl[57] vdd gnd cell_6t
Xbit_r58_c82 bl[82] br[82] wl[58] vdd gnd cell_6t
Xbit_r59_c82 bl[82] br[82] wl[59] vdd gnd cell_6t
Xbit_r60_c82 bl[82] br[82] wl[60] vdd gnd cell_6t
Xbit_r61_c82 bl[82] br[82] wl[61] vdd gnd cell_6t
Xbit_r62_c82 bl[82] br[82] wl[62] vdd gnd cell_6t
Xbit_r63_c82 bl[82] br[82] wl[63] vdd gnd cell_6t
Xbit_r64_c82 bl[82] br[82] wl[64] vdd gnd cell_6t
Xbit_r65_c82 bl[82] br[82] wl[65] vdd gnd cell_6t
Xbit_r66_c82 bl[82] br[82] wl[66] vdd gnd cell_6t
Xbit_r67_c82 bl[82] br[82] wl[67] vdd gnd cell_6t
Xbit_r68_c82 bl[82] br[82] wl[68] vdd gnd cell_6t
Xbit_r69_c82 bl[82] br[82] wl[69] vdd gnd cell_6t
Xbit_r70_c82 bl[82] br[82] wl[70] vdd gnd cell_6t
Xbit_r71_c82 bl[82] br[82] wl[71] vdd gnd cell_6t
Xbit_r72_c82 bl[82] br[82] wl[72] vdd gnd cell_6t
Xbit_r73_c82 bl[82] br[82] wl[73] vdd gnd cell_6t
Xbit_r74_c82 bl[82] br[82] wl[74] vdd gnd cell_6t
Xbit_r75_c82 bl[82] br[82] wl[75] vdd gnd cell_6t
Xbit_r76_c82 bl[82] br[82] wl[76] vdd gnd cell_6t
Xbit_r77_c82 bl[82] br[82] wl[77] vdd gnd cell_6t
Xbit_r78_c82 bl[82] br[82] wl[78] vdd gnd cell_6t
Xbit_r79_c82 bl[82] br[82] wl[79] vdd gnd cell_6t
Xbit_r80_c82 bl[82] br[82] wl[80] vdd gnd cell_6t
Xbit_r81_c82 bl[82] br[82] wl[81] vdd gnd cell_6t
Xbit_r82_c82 bl[82] br[82] wl[82] vdd gnd cell_6t
Xbit_r83_c82 bl[82] br[82] wl[83] vdd gnd cell_6t
Xbit_r84_c82 bl[82] br[82] wl[84] vdd gnd cell_6t
Xbit_r85_c82 bl[82] br[82] wl[85] vdd gnd cell_6t
Xbit_r86_c82 bl[82] br[82] wl[86] vdd gnd cell_6t
Xbit_r87_c82 bl[82] br[82] wl[87] vdd gnd cell_6t
Xbit_r88_c82 bl[82] br[82] wl[88] vdd gnd cell_6t
Xbit_r89_c82 bl[82] br[82] wl[89] vdd gnd cell_6t
Xbit_r90_c82 bl[82] br[82] wl[90] vdd gnd cell_6t
Xbit_r91_c82 bl[82] br[82] wl[91] vdd gnd cell_6t
Xbit_r92_c82 bl[82] br[82] wl[92] vdd gnd cell_6t
Xbit_r93_c82 bl[82] br[82] wl[93] vdd gnd cell_6t
Xbit_r94_c82 bl[82] br[82] wl[94] vdd gnd cell_6t
Xbit_r95_c82 bl[82] br[82] wl[95] vdd gnd cell_6t
Xbit_r96_c82 bl[82] br[82] wl[96] vdd gnd cell_6t
Xbit_r97_c82 bl[82] br[82] wl[97] vdd gnd cell_6t
Xbit_r98_c82 bl[82] br[82] wl[98] vdd gnd cell_6t
Xbit_r99_c82 bl[82] br[82] wl[99] vdd gnd cell_6t
Xbit_r100_c82 bl[82] br[82] wl[100] vdd gnd cell_6t
Xbit_r101_c82 bl[82] br[82] wl[101] vdd gnd cell_6t
Xbit_r102_c82 bl[82] br[82] wl[102] vdd gnd cell_6t
Xbit_r103_c82 bl[82] br[82] wl[103] vdd gnd cell_6t
Xbit_r104_c82 bl[82] br[82] wl[104] vdd gnd cell_6t
Xbit_r105_c82 bl[82] br[82] wl[105] vdd gnd cell_6t
Xbit_r106_c82 bl[82] br[82] wl[106] vdd gnd cell_6t
Xbit_r107_c82 bl[82] br[82] wl[107] vdd gnd cell_6t
Xbit_r108_c82 bl[82] br[82] wl[108] vdd gnd cell_6t
Xbit_r109_c82 bl[82] br[82] wl[109] vdd gnd cell_6t
Xbit_r110_c82 bl[82] br[82] wl[110] vdd gnd cell_6t
Xbit_r111_c82 bl[82] br[82] wl[111] vdd gnd cell_6t
Xbit_r112_c82 bl[82] br[82] wl[112] vdd gnd cell_6t
Xbit_r113_c82 bl[82] br[82] wl[113] vdd gnd cell_6t
Xbit_r114_c82 bl[82] br[82] wl[114] vdd gnd cell_6t
Xbit_r115_c82 bl[82] br[82] wl[115] vdd gnd cell_6t
Xbit_r116_c82 bl[82] br[82] wl[116] vdd gnd cell_6t
Xbit_r117_c82 bl[82] br[82] wl[117] vdd gnd cell_6t
Xbit_r118_c82 bl[82] br[82] wl[118] vdd gnd cell_6t
Xbit_r119_c82 bl[82] br[82] wl[119] vdd gnd cell_6t
Xbit_r120_c82 bl[82] br[82] wl[120] vdd gnd cell_6t
Xbit_r121_c82 bl[82] br[82] wl[121] vdd gnd cell_6t
Xbit_r122_c82 bl[82] br[82] wl[122] vdd gnd cell_6t
Xbit_r123_c82 bl[82] br[82] wl[123] vdd gnd cell_6t
Xbit_r124_c82 bl[82] br[82] wl[124] vdd gnd cell_6t
Xbit_r125_c82 bl[82] br[82] wl[125] vdd gnd cell_6t
Xbit_r126_c82 bl[82] br[82] wl[126] vdd gnd cell_6t
Xbit_r127_c82 bl[82] br[82] wl[127] vdd gnd cell_6t
Xbit_r0_c83 bl[83] br[83] wl[0] vdd gnd cell_6t
Xbit_r1_c83 bl[83] br[83] wl[1] vdd gnd cell_6t
Xbit_r2_c83 bl[83] br[83] wl[2] vdd gnd cell_6t
Xbit_r3_c83 bl[83] br[83] wl[3] vdd gnd cell_6t
Xbit_r4_c83 bl[83] br[83] wl[4] vdd gnd cell_6t
Xbit_r5_c83 bl[83] br[83] wl[5] vdd gnd cell_6t
Xbit_r6_c83 bl[83] br[83] wl[6] vdd gnd cell_6t
Xbit_r7_c83 bl[83] br[83] wl[7] vdd gnd cell_6t
Xbit_r8_c83 bl[83] br[83] wl[8] vdd gnd cell_6t
Xbit_r9_c83 bl[83] br[83] wl[9] vdd gnd cell_6t
Xbit_r10_c83 bl[83] br[83] wl[10] vdd gnd cell_6t
Xbit_r11_c83 bl[83] br[83] wl[11] vdd gnd cell_6t
Xbit_r12_c83 bl[83] br[83] wl[12] vdd gnd cell_6t
Xbit_r13_c83 bl[83] br[83] wl[13] vdd gnd cell_6t
Xbit_r14_c83 bl[83] br[83] wl[14] vdd gnd cell_6t
Xbit_r15_c83 bl[83] br[83] wl[15] vdd gnd cell_6t
Xbit_r16_c83 bl[83] br[83] wl[16] vdd gnd cell_6t
Xbit_r17_c83 bl[83] br[83] wl[17] vdd gnd cell_6t
Xbit_r18_c83 bl[83] br[83] wl[18] vdd gnd cell_6t
Xbit_r19_c83 bl[83] br[83] wl[19] vdd gnd cell_6t
Xbit_r20_c83 bl[83] br[83] wl[20] vdd gnd cell_6t
Xbit_r21_c83 bl[83] br[83] wl[21] vdd gnd cell_6t
Xbit_r22_c83 bl[83] br[83] wl[22] vdd gnd cell_6t
Xbit_r23_c83 bl[83] br[83] wl[23] vdd gnd cell_6t
Xbit_r24_c83 bl[83] br[83] wl[24] vdd gnd cell_6t
Xbit_r25_c83 bl[83] br[83] wl[25] vdd gnd cell_6t
Xbit_r26_c83 bl[83] br[83] wl[26] vdd gnd cell_6t
Xbit_r27_c83 bl[83] br[83] wl[27] vdd gnd cell_6t
Xbit_r28_c83 bl[83] br[83] wl[28] vdd gnd cell_6t
Xbit_r29_c83 bl[83] br[83] wl[29] vdd gnd cell_6t
Xbit_r30_c83 bl[83] br[83] wl[30] vdd gnd cell_6t
Xbit_r31_c83 bl[83] br[83] wl[31] vdd gnd cell_6t
Xbit_r32_c83 bl[83] br[83] wl[32] vdd gnd cell_6t
Xbit_r33_c83 bl[83] br[83] wl[33] vdd gnd cell_6t
Xbit_r34_c83 bl[83] br[83] wl[34] vdd gnd cell_6t
Xbit_r35_c83 bl[83] br[83] wl[35] vdd gnd cell_6t
Xbit_r36_c83 bl[83] br[83] wl[36] vdd gnd cell_6t
Xbit_r37_c83 bl[83] br[83] wl[37] vdd gnd cell_6t
Xbit_r38_c83 bl[83] br[83] wl[38] vdd gnd cell_6t
Xbit_r39_c83 bl[83] br[83] wl[39] vdd gnd cell_6t
Xbit_r40_c83 bl[83] br[83] wl[40] vdd gnd cell_6t
Xbit_r41_c83 bl[83] br[83] wl[41] vdd gnd cell_6t
Xbit_r42_c83 bl[83] br[83] wl[42] vdd gnd cell_6t
Xbit_r43_c83 bl[83] br[83] wl[43] vdd gnd cell_6t
Xbit_r44_c83 bl[83] br[83] wl[44] vdd gnd cell_6t
Xbit_r45_c83 bl[83] br[83] wl[45] vdd gnd cell_6t
Xbit_r46_c83 bl[83] br[83] wl[46] vdd gnd cell_6t
Xbit_r47_c83 bl[83] br[83] wl[47] vdd gnd cell_6t
Xbit_r48_c83 bl[83] br[83] wl[48] vdd gnd cell_6t
Xbit_r49_c83 bl[83] br[83] wl[49] vdd gnd cell_6t
Xbit_r50_c83 bl[83] br[83] wl[50] vdd gnd cell_6t
Xbit_r51_c83 bl[83] br[83] wl[51] vdd gnd cell_6t
Xbit_r52_c83 bl[83] br[83] wl[52] vdd gnd cell_6t
Xbit_r53_c83 bl[83] br[83] wl[53] vdd gnd cell_6t
Xbit_r54_c83 bl[83] br[83] wl[54] vdd gnd cell_6t
Xbit_r55_c83 bl[83] br[83] wl[55] vdd gnd cell_6t
Xbit_r56_c83 bl[83] br[83] wl[56] vdd gnd cell_6t
Xbit_r57_c83 bl[83] br[83] wl[57] vdd gnd cell_6t
Xbit_r58_c83 bl[83] br[83] wl[58] vdd gnd cell_6t
Xbit_r59_c83 bl[83] br[83] wl[59] vdd gnd cell_6t
Xbit_r60_c83 bl[83] br[83] wl[60] vdd gnd cell_6t
Xbit_r61_c83 bl[83] br[83] wl[61] vdd gnd cell_6t
Xbit_r62_c83 bl[83] br[83] wl[62] vdd gnd cell_6t
Xbit_r63_c83 bl[83] br[83] wl[63] vdd gnd cell_6t
Xbit_r64_c83 bl[83] br[83] wl[64] vdd gnd cell_6t
Xbit_r65_c83 bl[83] br[83] wl[65] vdd gnd cell_6t
Xbit_r66_c83 bl[83] br[83] wl[66] vdd gnd cell_6t
Xbit_r67_c83 bl[83] br[83] wl[67] vdd gnd cell_6t
Xbit_r68_c83 bl[83] br[83] wl[68] vdd gnd cell_6t
Xbit_r69_c83 bl[83] br[83] wl[69] vdd gnd cell_6t
Xbit_r70_c83 bl[83] br[83] wl[70] vdd gnd cell_6t
Xbit_r71_c83 bl[83] br[83] wl[71] vdd gnd cell_6t
Xbit_r72_c83 bl[83] br[83] wl[72] vdd gnd cell_6t
Xbit_r73_c83 bl[83] br[83] wl[73] vdd gnd cell_6t
Xbit_r74_c83 bl[83] br[83] wl[74] vdd gnd cell_6t
Xbit_r75_c83 bl[83] br[83] wl[75] vdd gnd cell_6t
Xbit_r76_c83 bl[83] br[83] wl[76] vdd gnd cell_6t
Xbit_r77_c83 bl[83] br[83] wl[77] vdd gnd cell_6t
Xbit_r78_c83 bl[83] br[83] wl[78] vdd gnd cell_6t
Xbit_r79_c83 bl[83] br[83] wl[79] vdd gnd cell_6t
Xbit_r80_c83 bl[83] br[83] wl[80] vdd gnd cell_6t
Xbit_r81_c83 bl[83] br[83] wl[81] vdd gnd cell_6t
Xbit_r82_c83 bl[83] br[83] wl[82] vdd gnd cell_6t
Xbit_r83_c83 bl[83] br[83] wl[83] vdd gnd cell_6t
Xbit_r84_c83 bl[83] br[83] wl[84] vdd gnd cell_6t
Xbit_r85_c83 bl[83] br[83] wl[85] vdd gnd cell_6t
Xbit_r86_c83 bl[83] br[83] wl[86] vdd gnd cell_6t
Xbit_r87_c83 bl[83] br[83] wl[87] vdd gnd cell_6t
Xbit_r88_c83 bl[83] br[83] wl[88] vdd gnd cell_6t
Xbit_r89_c83 bl[83] br[83] wl[89] vdd gnd cell_6t
Xbit_r90_c83 bl[83] br[83] wl[90] vdd gnd cell_6t
Xbit_r91_c83 bl[83] br[83] wl[91] vdd gnd cell_6t
Xbit_r92_c83 bl[83] br[83] wl[92] vdd gnd cell_6t
Xbit_r93_c83 bl[83] br[83] wl[93] vdd gnd cell_6t
Xbit_r94_c83 bl[83] br[83] wl[94] vdd gnd cell_6t
Xbit_r95_c83 bl[83] br[83] wl[95] vdd gnd cell_6t
Xbit_r96_c83 bl[83] br[83] wl[96] vdd gnd cell_6t
Xbit_r97_c83 bl[83] br[83] wl[97] vdd gnd cell_6t
Xbit_r98_c83 bl[83] br[83] wl[98] vdd gnd cell_6t
Xbit_r99_c83 bl[83] br[83] wl[99] vdd gnd cell_6t
Xbit_r100_c83 bl[83] br[83] wl[100] vdd gnd cell_6t
Xbit_r101_c83 bl[83] br[83] wl[101] vdd gnd cell_6t
Xbit_r102_c83 bl[83] br[83] wl[102] vdd gnd cell_6t
Xbit_r103_c83 bl[83] br[83] wl[103] vdd gnd cell_6t
Xbit_r104_c83 bl[83] br[83] wl[104] vdd gnd cell_6t
Xbit_r105_c83 bl[83] br[83] wl[105] vdd gnd cell_6t
Xbit_r106_c83 bl[83] br[83] wl[106] vdd gnd cell_6t
Xbit_r107_c83 bl[83] br[83] wl[107] vdd gnd cell_6t
Xbit_r108_c83 bl[83] br[83] wl[108] vdd gnd cell_6t
Xbit_r109_c83 bl[83] br[83] wl[109] vdd gnd cell_6t
Xbit_r110_c83 bl[83] br[83] wl[110] vdd gnd cell_6t
Xbit_r111_c83 bl[83] br[83] wl[111] vdd gnd cell_6t
Xbit_r112_c83 bl[83] br[83] wl[112] vdd gnd cell_6t
Xbit_r113_c83 bl[83] br[83] wl[113] vdd gnd cell_6t
Xbit_r114_c83 bl[83] br[83] wl[114] vdd gnd cell_6t
Xbit_r115_c83 bl[83] br[83] wl[115] vdd gnd cell_6t
Xbit_r116_c83 bl[83] br[83] wl[116] vdd gnd cell_6t
Xbit_r117_c83 bl[83] br[83] wl[117] vdd gnd cell_6t
Xbit_r118_c83 bl[83] br[83] wl[118] vdd gnd cell_6t
Xbit_r119_c83 bl[83] br[83] wl[119] vdd gnd cell_6t
Xbit_r120_c83 bl[83] br[83] wl[120] vdd gnd cell_6t
Xbit_r121_c83 bl[83] br[83] wl[121] vdd gnd cell_6t
Xbit_r122_c83 bl[83] br[83] wl[122] vdd gnd cell_6t
Xbit_r123_c83 bl[83] br[83] wl[123] vdd gnd cell_6t
Xbit_r124_c83 bl[83] br[83] wl[124] vdd gnd cell_6t
Xbit_r125_c83 bl[83] br[83] wl[125] vdd gnd cell_6t
Xbit_r126_c83 bl[83] br[83] wl[126] vdd gnd cell_6t
Xbit_r127_c83 bl[83] br[83] wl[127] vdd gnd cell_6t
Xbit_r0_c84 bl[84] br[84] wl[0] vdd gnd cell_6t
Xbit_r1_c84 bl[84] br[84] wl[1] vdd gnd cell_6t
Xbit_r2_c84 bl[84] br[84] wl[2] vdd gnd cell_6t
Xbit_r3_c84 bl[84] br[84] wl[3] vdd gnd cell_6t
Xbit_r4_c84 bl[84] br[84] wl[4] vdd gnd cell_6t
Xbit_r5_c84 bl[84] br[84] wl[5] vdd gnd cell_6t
Xbit_r6_c84 bl[84] br[84] wl[6] vdd gnd cell_6t
Xbit_r7_c84 bl[84] br[84] wl[7] vdd gnd cell_6t
Xbit_r8_c84 bl[84] br[84] wl[8] vdd gnd cell_6t
Xbit_r9_c84 bl[84] br[84] wl[9] vdd gnd cell_6t
Xbit_r10_c84 bl[84] br[84] wl[10] vdd gnd cell_6t
Xbit_r11_c84 bl[84] br[84] wl[11] vdd gnd cell_6t
Xbit_r12_c84 bl[84] br[84] wl[12] vdd gnd cell_6t
Xbit_r13_c84 bl[84] br[84] wl[13] vdd gnd cell_6t
Xbit_r14_c84 bl[84] br[84] wl[14] vdd gnd cell_6t
Xbit_r15_c84 bl[84] br[84] wl[15] vdd gnd cell_6t
Xbit_r16_c84 bl[84] br[84] wl[16] vdd gnd cell_6t
Xbit_r17_c84 bl[84] br[84] wl[17] vdd gnd cell_6t
Xbit_r18_c84 bl[84] br[84] wl[18] vdd gnd cell_6t
Xbit_r19_c84 bl[84] br[84] wl[19] vdd gnd cell_6t
Xbit_r20_c84 bl[84] br[84] wl[20] vdd gnd cell_6t
Xbit_r21_c84 bl[84] br[84] wl[21] vdd gnd cell_6t
Xbit_r22_c84 bl[84] br[84] wl[22] vdd gnd cell_6t
Xbit_r23_c84 bl[84] br[84] wl[23] vdd gnd cell_6t
Xbit_r24_c84 bl[84] br[84] wl[24] vdd gnd cell_6t
Xbit_r25_c84 bl[84] br[84] wl[25] vdd gnd cell_6t
Xbit_r26_c84 bl[84] br[84] wl[26] vdd gnd cell_6t
Xbit_r27_c84 bl[84] br[84] wl[27] vdd gnd cell_6t
Xbit_r28_c84 bl[84] br[84] wl[28] vdd gnd cell_6t
Xbit_r29_c84 bl[84] br[84] wl[29] vdd gnd cell_6t
Xbit_r30_c84 bl[84] br[84] wl[30] vdd gnd cell_6t
Xbit_r31_c84 bl[84] br[84] wl[31] vdd gnd cell_6t
Xbit_r32_c84 bl[84] br[84] wl[32] vdd gnd cell_6t
Xbit_r33_c84 bl[84] br[84] wl[33] vdd gnd cell_6t
Xbit_r34_c84 bl[84] br[84] wl[34] vdd gnd cell_6t
Xbit_r35_c84 bl[84] br[84] wl[35] vdd gnd cell_6t
Xbit_r36_c84 bl[84] br[84] wl[36] vdd gnd cell_6t
Xbit_r37_c84 bl[84] br[84] wl[37] vdd gnd cell_6t
Xbit_r38_c84 bl[84] br[84] wl[38] vdd gnd cell_6t
Xbit_r39_c84 bl[84] br[84] wl[39] vdd gnd cell_6t
Xbit_r40_c84 bl[84] br[84] wl[40] vdd gnd cell_6t
Xbit_r41_c84 bl[84] br[84] wl[41] vdd gnd cell_6t
Xbit_r42_c84 bl[84] br[84] wl[42] vdd gnd cell_6t
Xbit_r43_c84 bl[84] br[84] wl[43] vdd gnd cell_6t
Xbit_r44_c84 bl[84] br[84] wl[44] vdd gnd cell_6t
Xbit_r45_c84 bl[84] br[84] wl[45] vdd gnd cell_6t
Xbit_r46_c84 bl[84] br[84] wl[46] vdd gnd cell_6t
Xbit_r47_c84 bl[84] br[84] wl[47] vdd gnd cell_6t
Xbit_r48_c84 bl[84] br[84] wl[48] vdd gnd cell_6t
Xbit_r49_c84 bl[84] br[84] wl[49] vdd gnd cell_6t
Xbit_r50_c84 bl[84] br[84] wl[50] vdd gnd cell_6t
Xbit_r51_c84 bl[84] br[84] wl[51] vdd gnd cell_6t
Xbit_r52_c84 bl[84] br[84] wl[52] vdd gnd cell_6t
Xbit_r53_c84 bl[84] br[84] wl[53] vdd gnd cell_6t
Xbit_r54_c84 bl[84] br[84] wl[54] vdd gnd cell_6t
Xbit_r55_c84 bl[84] br[84] wl[55] vdd gnd cell_6t
Xbit_r56_c84 bl[84] br[84] wl[56] vdd gnd cell_6t
Xbit_r57_c84 bl[84] br[84] wl[57] vdd gnd cell_6t
Xbit_r58_c84 bl[84] br[84] wl[58] vdd gnd cell_6t
Xbit_r59_c84 bl[84] br[84] wl[59] vdd gnd cell_6t
Xbit_r60_c84 bl[84] br[84] wl[60] vdd gnd cell_6t
Xbit_r61_c84 bl[84] br[84] wl[61] vdd gnd cell_6t
Xbit_r62_c84 bl[84] br[84] wl[62] vdd gnd cell_6t
Xbit_r63_c84 bl[84] br[84] wl[63] vdd gnd cell_6t
Xbit_r64_c84 bl[84] br[84] wl[64] vdd gnd cell_6t
Xbit_r65_c84 bl[84] br[84] wl[65] vdd gnd cell_6t
Xbit_r66_c84 bl[84] br[84] wl[66] vdd gnd cell_6t
Xbit_r67_c84 bl[84] br[84] wl[67] vdd gnd cell_6t
Xbit_r68_c84 bl[84] br[84] wl[68] vdd gnd cell_6t
Xbit_r69_c84 bl[84] br[84] wl[69] vdd gnd cell_6t
Xbit_r70_c84 bl[84] br[84] wl[70] vdd gnd cell_6t
Xbit_r71_c84 bl[84] br[84] wl[71] vdd gnd cell_6t
Xbit_r72_c84 bl[84] br[84] wl[72] vdd gnd cell_6t
Xbit_r73_c84 bl[84] br[84] wl[73] vdd gnd cell_6t
Xbit_r74_c84 bl[84] br[84] wl[74] vdd gnd cell_6t
Xbit_r75_c84 bl[84] br[84] wl[75] vdd gnd cell_6t
Xbit_r76_c84 bl[84] br[84] wl[76] vdd gnd cell_6t
Xbit_r77_c84 bl[84] br[84] wl[77] vdd gnd cell_6t
Xbit_r78_c84 bl[84] br[84] wl[78] vdd gnd cell_6t
Xbit_r79_c84 bl[84] br[84] wl[79] vdd gnd cell_6t
Xbit_r80_c84 bl[84] br[84] wl[80] vdd gnd cell_6t
Xbit_r81_c84 bl[84] br[84] wl[81] vdd gnd cell_6t
Xbit_r82_c84 bl[84] br[84] wl[82] vdd gnd cell_6t
Xbit_r83_c84 bl[84] br[84] wl[83] vdd gnd cell_6t
Xbit_r84_c84 bl[84] br[84] wl[84] vdd gnd cell_6t
Xbit_r85_c84 bl[84] br[84] wl[85] vdd gnd cell_6t
Xbit_r86_c84 bl[84] br[84] wl[86] vdd gnd cell_6t
Xbit_r87_c84 bl[84] br[84] wl[87] vdd gnd cell_6t
Xbit_r88_c84 bl[84] br[84] wl[88] vdd gnd cell_6t
Xbit_r89_c84 bl[84] br[84] wl[89] vdd gnd cell_6t
Xbit_r90_c84 bl[84] br[84] wl[90] vdd gnd cell_6t
Xbit_r91_c84 bl[84] br[84] wl[91] vdd gnd cell_6t
Xbit_r92_c84 bl[84] br[84] wl[92] vdd gnd cell_6t
Xbit_r93_c84 bl[84] br[84] wl[93] vdd gnd cell_6t
Xbit_r94_c84 bl[84] br[84] wl[94] vdd gnd cell_6t
Xbit_r95_c84 bl[84] br[84] wl[95] vdd gnd cell_6t
Xbit_r96_c84 bl[84] br[84] wl[96] vdd gnd cell_6t
Xbit_r97_c84 bl[84] br[84] wl[97] vdd gnd cell_6t
Xbit_r98_c84 bl[84] br[84] wl[98] vdd gnd cell_6t
Xbit_r99_c84 bl[84] br[84] wl[99] vdd gnd cell_6t
Xbit_r100_c84 bl[84] br[84] wl[100] vdd gnd cell_6t
Xbit_r101_c84 bl[84] br[84] wl[101] vdd gnd cell_6t
Xbit_r102_c84 bl[84] br[84] wl[102] vdd gnd cell_6t
Xbit_r103_c84 bl[84] br[84] wl[103] vdd gnd cell_6t
Xbit_r104_c84 bl[84] br[84] wl[104] vdd gnd cell_6t
Xbit_r105_c84 bl[84] br[84] wl[105] vdd gnd cell_6t
Xbit_r106_c84 bl[84] br[84] wl[106] vdd gnd cell_6t
Xbit_r107_c84 bl[84] br[84] wl[107] vdd gnd cell_6t
Xbit_r108_c84 bl[84] br[84] wl[108] vdd gnd cell_6t
Xbit_r109_c84 bl[84] br[84] wl[109] vdd gnd cell_6t
Xbit_r110_c84 bl[84] br[84] wl[110] vdd gnd cell_6t
Xbit_r111_c84 bl[84] br[84] wl[111] vdd gnd cell_6t
Xbit_r112_c84 bl[84] br[84] wl[112] vdd gnd cell_6t
Xbit_r113_c84 bl[84] br[84] wl[113] vdd gnd cell_6t
Xbit_r114_c84 bl[84] br[84] wl[114] vdd gnd cell_6t
Xbit_r115_c84 bl[84] br[84] wl[115] vdd gnd cell_6t
Xbit_r116_c84 bl[84] br[84] wl[116] vdd gnd cell_6t
Xbit_r117_c84 bl[84] br[84] wl[117] vdd gnd cell_6t
Xbit_r118_c84 bl[84] br[84] wl[118] vdd gnd cell_6t
Xbit_r119_c84 bl[84] br[84] wl[119] vdd gnd cell_6t
Xbit_r120_c84 bl[84] br[84] wl[120] vdd gnd cell_6t
Xbit_r121_c84 bl[84] br[84] wl[121] vdd gnd cell_6t
Xbit_r122_c84 bl[84] br[84] wl[122] vdd gnd cell_6t
Xbit_r123_c84 bl[84] br[84] wl[123] vdd gnd cell_6t
Xbit_r124_c84 bl[84] br[84] wl[124] vdd gnd cell_6t
Xbit_r125_c84 bl[84] br[84] wl[125] vdd gnd cell_6t
Xbit_r126_c84 bl[84] br[84] wl[126] vdd gnd cell_6t
Xbit_r127_c84 bl[84] br[84] wl[127] vdd gnd cell_6t
Xbit_r0_c85 bl[85] br[85] wl[0] vdd gnd cell_6t
Xbit_r1_c85 bl[85] br[85] wl[1] vdd gnd cell_6t
Xbit_r2_c85 bl[85] br[85] wl[2] vdd gnd cell_6t
Xbit_r3_c85 bl[85] br[85] wl[3] vdd gnd cell_6t
Xbit_r4_c85 bl[85] br[85] wl[4] vdd gnd cell_6t
Xbit_r5_c85 bl[85] br[85] wl[5] vdd gnd cell_6t
Xbit_r6_c85 bl[85] br[85] wl[6] vdd gnd cell_6t
Xbit_r7_c85 bl[85] br[85] wl[7] vdd gnd cell_6t
Xbit_r8_c85 bl[85] br[85] wl[8] vdd gnd cell_6t
Xbit_r9_c85 bl[85] br[85] wl[9] vdd gnd cell_6t
Xbit_r10_c85 bl[85] br[85] wl[10] vdd gnd cell_6t
Xbit_r11_c85 bl[85] br[85] wl[11] vdd gnd cell_6t
Xbit_r12_c85 bl[85] br[85] wl[12] vdd gnd cell_6t
Xbit_r13_c85 bl[85] br[85] wl[13] vdd gnd cell_6t
Xbit_r14_c85 bl[85] br[85] wl[14] vdd gnd cell_6t
Xbit_r15_c85 bl[85] br[85] wl[15] vdd gnd cell_6t
Xbit_r16_c85 bl[85] br[85] wl[16] vdd gnd cell_6t
Xbit_r17_c85 bl[85] br[85] wl[17] vdd gnd cell_6t
Xbit_r18_c85 bl[85] br[85] wl[18] vdd gnd cell_6t
Xbit_r19_c85 bl[85] br[85] wl[19] vdd gnd cell_6t
Xbit_r20_c85 bl[85] br[85] wl[20] vdd gnd cell_6t
Xbit_r21_c85 bl[85] br[85] wl[21] vdd gnd cell_6t
Xbit_r22_c85 bl[85] br[85] wl[22] vdd gnd cell_6t
Xbit_r23_c85 bl[85] br[85] wl[23] vdd gnd cell_6t
Xbit_r24_c85 bl[85] br[85] wl[24] vdd gnd cell_6t
Xbit_r25_c85 bl[85] br[85] wl[25] vdd gnd cell_6t
Xbit_r26_c85 bl[85] br[85] wl[26] vdd gnd cell_6t
Xbit_r27_c85 bl[85] br[85] wl[27] vdd gnd cell_6t
Xbit_r28_c85 bl[85] br[85] wl[28] vdd gnd cell_6t
Xbit_r29_c85 bl[85] br[85] wl[29] vdd gnd cell_6t
Xbit_r30_c85 bl[85] br[85] wl[30] vdd gnd cell_6t
Xbit_r31_c85 bl[85] br[85] wl[31] vdd gnd cell_6t
Xbit_r32_c85 bl[85] br[85] wl[32] vdd gnd cell_6t
Xbit_r33_c85 bl[85] br[85] wl[33] vdd gnd cell_6t
Xbit_r34_c85 bl[85] br[85] wl[34] vdd gnd cell_6t
Xbit_r35_c85 bl[85] br[85] wl[35] vdd gnd cell_6t
Xbit_r36_c85 bl[85] br[85] wl[36] vdd gnd cell_6t
Xbit_r37_c85 bl[85] br[85] wl[37] vdd gnd cell_6t
Xbit_r38_c85 bl[85] br[85] wl[38] vdd gnd cell_6t
Xbit_r39_c85 bl[85] br[85] wl[39] vdd gnd cell_6t
Xbit_r40_c85 bl[85] br[85] wl[40] vdd gnd cell_6t
Xbit_r41_c85 bl[85] br[85] wl[41] vdd gnd cell_6t
Xbit_r42_c85 bl[85] br[85] wl[42] vdd gnd cell_6t
Xbit_r43_c85 bl[85] br[85] wl[43] vdd gnd cell_6t
Xbit_r44_c85 bl[85] br[85] wl[44] vdd gnd cell_6t
Xbit_r45_c85 bl[85] br[85] wl[45] vdd gnd cell_6t
Xbit_r46_c85 bl[85] br[85] wl[46] vdd gnd cell_6t
Xbit_r47_c85 bl[85] br[85] wl[47] vdd gnd cell_6t
Xbit_r48_c85 bl[85] br[85] wl[48] vdd gnd cell_6t
Xbit_r49_c85 bl[85] br[85] wl[49] vdd gnd cell_6t
Xbit_r50_c85 bl[85] br[85] wl[50] vdd gnd cell_6t
Xbit_r51_c85 bl[85] br[85] wl[51] vdd gnd cell_6t
Xbit_r52_c85 bl[85] br[85] wl[52] vdd gnd cell_6t
Xbit_r53_c85 bl[85] br[85] wl[53] vdd gnd cell_6t
Xbit_r54_c85 bl[85] br[85] wl[54] vdd gnd cell_6t
Xbit_r55_c85 bl[85] br[85] wl[55] vdd gnd cell_6t
Xbit_r56_c85 bl[85] br[85] wl[56] vdd gnd cell_6t
Xbit_r57_c85 bl[85] br[85] wl[57] vdd gnd cell_6t
Xbit_r58_c85 bl[85] br[85] wl[58] vdd gnd cell_6t
Xbit_r59_c85 bl[85] br[85] wl[59] vdd gnd cell_6t
Xbit_r60_c85 bl[85] br[85] wl[60] vdd gnd cell_6t
Xbit_r61_c85 bl[85] br[85] wl[61] vdd gnd cell_6t
Xbit_r62_c85 bl[85] br[85] wl[62] vdd gnd cell_6t
Xbit_r63_c85 bl[85] br[85] wl[63] vdd gnd cell_6t
Xbit_r64_c85 bl[85] br[85] wl[64] vdd gnd cell_6t
Xbit_r65_c85 bl[85] br[85] wl[65] vdd gnd cell_6t
Xbit_r66_c85 bl[85] br[85] wl[66] vdd gnd cell_6t
Xbit_r67_c85 bl[85] br[85] wl[67] vdd gnd cell_6t
Xbit_r68_c85 bl[85] br[85] wl[68] vdd gnd cell_6t
Xbit_r69_c85 bl[85] br[85] wl[69] vdd gnd cell_6t
Xbit_r70_c85 bl[85] br[85] wl[70] vdd gnd cell_6t
Xbit_r71_c85 bl[85] br[85] wl[71] vdd gnd cell_6t
Xbit_r72_c85 bl[85] br[85] wl[72] vdd gnd cell_6t
Xbit_r73_c85 bl[85] br[85] wl[73] vdd gnd cell_6t
Xbit_r74_c85 bl[85] br[85] wl[74] vdd gnd cell_6t
Xbit_r75_c85 bl[85] br[85] wl[75] vdd gnd cell_6t
Xbit_r76_c85 bl[85] br[85] wl[76] vdd gnd cell_6t
Xbit_r77_c85 bl[85] br[85] wl[77] vdd gnd cell_6t
Xbit_r78_c85 bl[85] br[85] wl[78] vdd gnd cell_6t
Xbit_r79_c85 bl[85] br[85] wl[79] vdd gnd cell_6t
Xbit_r80_c85 bl[85] br[85] wl[80] vdd gnd cell_6t
Xbit_r81_c85 bl[85] br[85] wl[81] vdd gnd cell_6t
Xbit_r82_c85 bl[85] br[85] wl[82] vdd gnd cell_6t
Xbit_r83_c85 bl[85] br[85] wl[83] vdd gnd cell_6t
Xbit_r84_c85 bl[85] br[85] wl[84] vdd gnd cell_6t
Xbit_r85_c85 bl[85] br[85] wl[85] vdd gnd cell_6t
Xbit_r86_c85 bl[85] br[85] wl[86] vdd gnd cell_6t
Xbit_r87_c85 bl[85] br[85] wl[87] vdd gnd cell_6t
Xbit_r88_c85 bl[85] br[85] wl[88] vdd gnd cell_6t
Xbit_r89_c85 bl[85] br[85] wl[89] vdd gnd cell_6t
Xbit_r90_c85 bl[85] br[85] wl[90] vdd gnd cell_6t
Xbit_r91_c85 bl[85] br[85] wl[91] vdd gnd cell_6t
Xbit_r92_c85 bl[85] br[85] wl[92] vdd gnd cell_6t
Xbit_r93_c85 bl[85] br[85] wl[93] vdd gnd cell_6t
Xbit_r94_c85 bl[85] br[85] wl[94] vdd gnd cell_6t
Xbit_r95_c85 bl[85] br[85] wl[95] vdd gnd cell_6t
Xbit_r96_c85 bl[85] br[85] wl[96] vdd gnd cell_6t
Xbit_r97_c85 bl[85] br[85] wl[97] vdd gnd cell_6t
Xbit_r98_c85 bl[85] br[85] wl[98] vdd gnd cell_6t
Xbit_r99_c85 bl[85] br[85] wl[99] vdd gnd cell_6t
Xbit_r100_c85 bl[85] br[85] wl[100] vdd gnd cell_6t
Xbit_r101_c85 bl[85] br[85] wl[101] vdd gnd cell_6t
Xbit_r102_c85 bl[85] br[85] wl[102] vdd gnd cell_6t
Xbit_r103_c85 bl[85] br[85] wl[103] vdd gnd cell_6t
Xbit_r104_c85 bl[85] br[85] wl[104] vdd gnd cell_6t
Xbit_r105_c85 bl[85] br[85] wl[105] vdd gnd cell_6t
Xbit_r106_c85 bl[85] br[85] wl[106] vdd gnd cell_6t
Xbit_r107_c85 bl[85] br[85] wl[107] vdd gnd cell_6t
Xbit_r108_c85 bl[85] br[85] wl[108] vdd gnd cell_6t
Xbit_r109_c85 bl[85] br[85] wl[109] vdd gnd cell_6t
Xbit_r110_c85 bl[85] br[85] wl[110] vdd gnd cell_6t
Xbit_r111_c85 bl[85] br[85] wl[111] vdd gnd cell_6t
Xbit_r112_c85 bl[85] br[85] wl[112] vdd gnd cell_6t
Xbit_r113_c85 bl[85] br[85] wl[113] vdd gnd cell_6t
Xbit_r114_c85 bl[85] br[85] wl[114] vdd gnd cell_6t
Xbit_r115_c85 bl[85] br[85] wl[115] vdd gnd cell_6t
Xbit_r116_c85 bl[85] br[85] wl[116] vdd gnd cell_6t
Xbit_r117_c85 bl[85] br[85] wl[117] vdd gnd cell_6t
Xbit_r118_c85 bl[85] br[85] wl[118] vdd gnd cell_6t
Xbit_r119_c85 bl[85] br[85] wl[119] vdd gnd cell_6t
Xbit_r120_c85 bl[85] br[85] wl[120] vdd gnd cell_6t
Xbit_r121_c85 bl[85] br[85] wl[121] vdd gnd cell_6t
Xbit_r122_c85 bl[85] br[85] wl[122] vdd gnd cell_6t
Xbit_r123_c85 bl[85] br[85] wl[123] vdd gnd cell_6t
Xbit_r124_c85 bl[85] br[85] wl[124] vdd gnd cell_6t
Xbit_r125_c85 bl[85] br[85] wl[125] vdd gnd cell_6t
Xbit_r126_c85 bl[85] br[85] wl[126] vdd gnd cell_6t
Xbit_r127_c85 bl[85] br[85] wl[127] vdd gnd cell_6t
Xbit_r0_c86 bl[86] br[86] wl[0] vdd gnd cell_6t
Xbit_r1_c86 bl[86] br[86] wl[1] vdd gnd cell_6t
Xbit_r2_c86 bl[86] br[86] wl[2] vdd gnd cell_6t
Xbit_r3_c86 bl[86] br[86] wl[3] vdd gnd cell_6t
Xbit_r4_c86 bl[86] br[86] wl[4] vdd gnd cell_6t
Xbit_r5_c86 bl[86] br[86] wl[5] vdd gnd cell_6t
Xbit_r6_c86 bl[86] br[86] wl[6] vdd gnd cell_6t
Xbit_r7_c86 bl[86] br[86] wl[7] vdd gnd cell_6t
Xbit_r8_c86 bl[86] br[86] wl[8] vdd gnd cell_6t
Xbit_r9_c86 bl[86] br[86] wl[9] vdd gnd cell_6t
Xbit_r10_c86 bl[86] br[86] wl[10] vdd gnd cell_6t
Xbit_r11_c86 bl[86] br[86] wl[11] vdd gnd cell_6t
Xbit_r12_c86 bl[86] br[86] wl[12] vdd gnd cell_6t
Xbit_r13_c86 bl[86] br[86] wl[13] vdd gnd cell_6t
Xbit_r14_c86 bl[86] br[86] wl[14] vdd gnd cell_6t
Xbit_r15_c86 bl[86] br[86] wl[15] vdd gnd cell_6t
Xbit_r16_c86 bl[86] br[86] wl[16] vdd gnd cell_6t
Xbit_r17_c86 bl[86] br[86] wl[17] vdd gnd cell_6t
Xbit_r18_c86 bl[86] br[86] wl[18] vdd gnd cell_6t
Xbit_r19_c86 bl[86] br[86] wl[19] vdd gnd cell_6t
Xbit_r20_c86 bl[86] br[86] wl[20] vdd gnd cell_6t
Xbit_r21_c86 bl[86] br[86] wl[21] vdd gnd cell_6t
Xbit_r22_c86 bl[86] br[86] wl[22] vdd gnd cell_6t
Xbit_r23_c86 bl[86] br[86] wl[23] vdd gnd cell_6t
Xbit_r24_c86 bl[86] br[86] wl[24] vdd gnd cell_6t
Xbit_r25_c86 bl[86] br[86] wl[25] vdd gnd cell_6t
Xbit_r26_c86 bl[86] br[86] wl[26] vdd gnd cell_6t
Xbit_r27_c86 bl[86] br[86] wl[27] vdd gnd cell_6t
Xbit_r28_c86 bl[86] br[86] wl[28] vdd gnd cell_6t
Xbit_r29_c86 bl[86] br[86] wl[29] vdd gnd cell_6t
Xbit_r30_c86 bl[86] br[86] wl[30] vdd gnd cell_6t
Xbit_r31_c86 bl[86] br[86] wl[31] vdd gnd cell_6t
Xbit_r32_c86 bl[86] br[86] wl[32] vdd gnd cell_6t
Xbit_r33_c86 bl[86] br[86] wl[33] vdd gnd cell_6t
Xbit_r34_c86 bl[86] br[86] wl[34] vdd gnd cell_6t
Xbit_r35_c86 bl[86] br[86] wl[35] vdd gnd cell_6t
Xbit_r36_c86 bl[86] br[86] wl[36] vdd gnd cell_6t
Xbit_r37_c86 bl[86] br[86] wl[37] vdd gnd cell_6t
Xbit_r38_c86 bl[86] br[86] wl[38] vdd gnd cell_6t
Xbit_r39_c86 bl[86] br[86] wl[39] vdd gnd cell_6t
Xbit_r40_c86 bl[86] br[86] wl[40] vdd gnd cell_6t
Xbit_r41_c86 bl[86] br[86] wl[41] vdd gnd cell_6t
Xbit_r42_c86 bl[86] br[86] wl[42] vdd gnd cell_6t
Xbit_r43_c86 bl[86] br[86] wl[43] vdd gnd cell_6t
Xbit_r44_c86 bl[86] br[86] wl[44] vdd gnd cell_6t
Xbit_r45_c86 bl[86] br[86] wl[45] vdd gnd cell_6t
Xbit_r46_c86 bl[86] br[86] wl[46] vdd gnd cell_6t
Xbit_r47_c86 bl[86] br[86] wl[47] vdd gnd cell_6t
Xbit_r48_c86 bl[86] br[86] wl[48] vdd gnd cell_6t
Xbit_r49_c86 bl[86] br[86] wl[49] vdd gnd cell_6t
Xbit_r50_c86 bl[86] br[86] wl[50] vdd gnd cell_6t
Xbit_r51_c86 bl[86] br[86] wl[51] vdd gnd cell_6t
Xbit_r52_c86 bl[86] br[86] wl[52] vdd gnd cell_6t
Xbit_r53_c86 bl[86] br[86] wl[53] vdd gnd cell_6t
Xbit_r54_c86 bl[86] br[86] wl[54] vdd gnd cell_6t
Xbit_r55_c86 bl[86] br[86] wl[55] vdd gnd cell_6t
Xbit_r56_c86 bl[86] br[86] wl[56] vdd gnd cell_6t
Xbit_r57_c86 bl[86] br[86] wl[57] vdd gnd cell_6t
Xbit_r58_c86 bl[86] br[86] wl[58] vdd gnd cell_6t
Xbit_r59_c86 bl[86] br[86] wl[59] vdd gnd cell_6t
Xbit_r60_c86 bl[86] br[86] wl[60] vdd gnd cell_6t
Xbit_r61_c86 bl[86] br[86] wl[61] vdd gnd cell_6t
Xbit_r62_c86 bl[86] br[86] wl[62] vdd gnd cell_6t
Xbit_r63_c86 bl[86] br[86] wl[63] vdd gnd cell_6t
Xbit_r64_c86 bl[86] br[86] wl[64] vdd gnd cell_6t
Xbit_r65_c86 bl[86] br[86] wl[65] vdd gnd cell_6t
Xbit_r66_c86 bl[86] br[86] wl[66] vdd gnd cell_6t
Xbit_r67_c86 bl[86] br[86] wl[67] vdd gnd cell_6t
Xbit_r68_c86 bl[86] br[86] wl[68] vdd gnd cell_6t
Xbit_r69_c86 bl[86] br[86] wl[69] vdd gnd cell_6t
Xbit_r70_c86 bl[86] br[86] wl[70] vdd gnd cell_6t
Xbit_r71_c86 bl[86] br[86] wl[71] vdd gnd cell_6t
Xbit_r72_c86 bl[86] br[86] wl[72] vdd gnd cell_6t
Xbit_r73_c86 bl[86] br[86] wl[73] vdd gnd cell_6t
Xbit_r74_c86 bl[86] br[86] wl[74] vdd gnd cell_6t
Xbit_r75_c86 bl[86] br[86] wl[75] vdd gnd cell_6t
Xbit_r76_c86 bl[86] br[86] wl[76] vdd gnd cell_6t
Xbit_r77_c86 bl[86] br[86] wl[77] vdd gnd cell_6t
Xbit_r78_c86 bl[86] br[86] wl[78] vdd gnd cell_6t
Xbit_r79_c86 bl[86] br[86] wl[79] vdd gnd cell_6t
Xbit_r80_c86 bl[86] br[86] wl[80] vdd gnd cell_6t
Xbit_r81_c86 bl[86] br[86] wl[81] vdd gnd cell_6t
Xbit_r82_c86 bl[86] br[86] wl[82] vdd gnd cell_6t
Xbit_r83_c86 bl[86] br[86] wl[83] vdd gnd cell_6t
Xbit_r84_c86 bl[86] br[86] wl[84] vdd gnd cell_6t
Xbit_r85_c86 bl[86] br[86] wl[85] vdd gnd cell_6t
Xbit_r86_c86 bl[86] br[86] wl[86] vdd gnd cell_6t
Xbit_r87_c86 bl[86] br[86] wl[87] vdd gnd cell_6t
Xbit_r88_c86 bl[86] br[86] wl[88] vdd gnd cell_6t
Xbit_r89_c86 bl[86] br[86] wl[89] vdd gnd cell_6t
Xbit_r90_c86 bl[86] br[86] wl[90] vdd gnd cell_6t
Xbit_r91_c86 bl[86] br[86] wl[91] vdd gnd cell_6t
Xbit_r92_c86 bl[86] br[86] wl[92] vdd gnd cell_6t
Xbit_r93_c86 bl[86] br[86] wl[93] vdd gnd cell_6t
Xbit_r94_c86 bl[86] br[86] wl[94] vdd gnd cell_6t
Xbit_r95_c86 bl[86] br[86] wl[95] vdd gnd cell_6t
Xbit_r96_c86 bl[86] br[86] wl[96] vdd gnd cell_6t
Xbit_r97_c86 bl[86] br[86] wl[97] vdd gnd cell_6t
Xbit_r98_c86 bl[86] br[86] wl[98] vdd gnd cell_6t
Xbit_r99_c86 bl[86] br[86] wl[99] vdd gnd cell_6t
Xbit_r100_c86 bl[86] br[86] wl[100] vdd gnd cell_6t
Xbit_r101_c86 bl[86] br[86] wl[101] vdd gnd cell_6t
Xbit_r102_c86 bl[86] br[86] wl[102] vdd gnd cell_6t
Xbit_r103_c86 bl[86] br[86] wl[103] vdd gnd cell_6t
Xbit_r104_c86 bl[86] br[86] wl[104] vdd gnd cell_6t
Xbit_r105_c86 bl[86] br[86] wl[105] vdd gnd cell_6t
Xbit_r106_c86 bl[86] br[86] wl[106] vdd gnd cell_6t
Xbit_r107_c86 bl[86] br[86] wl[107] vdd gnd cell_6t
Xbit_r108_c86 bl[86] br[86] wl[108] vdd gnd cell_6t
Xbit_r109_c86 bl[86] br[86] wl[109] vdd gnd cell_6t
Xbit_r110_c86 bl[86] br[86] wl[110] vdd gnd cell_6t
Xbit_r111_c86 bl[86] br[86] wl[111] vdd gnd cell_6t
Xbit_r112_c86 bl[86] br[86] wl[112] vdd gnd cell_6t
Xbit_r113_c86 bl[86] br[86] wl[113] vdd gnd cell_6t
Xbit_r114_c86 bl[86] br[86] wl[114] vdd gnd cell_6t
Xbit_r115_c86 bl[86] br[86] wl[115] vdd gnd cell_6t
Xbit_r116_c86 bl[86] br[86] wl[116] vdd gnd cell_6t
Xbit_r117_c86 bl[86] br[86] wl[117] vdd gnd cell_6t
Xbit_r118_c86 bl[86] br[86] wl[118] vdd gnd cell_6t
Xbit_r119_c86 bl[86] br[86] wl[119] vdd gnd cell_6t
Xbit_r120_c86 bl[86] br[86] wl[120] vdd gnd cell_6t
Xbit_r121_c86 bl[86] br[86] wl[121] vdd gnd cell_6t
Xbit_r122_c86 bl[86] br[86] wl[122] vdd gnd cell_6t
Xbit_r123_c86 bl[86] br[86] wl[123] vdd gnd cell_6t
Xbit_r124_c86 bl[86] br[86] wl[124] vdd gnd cell_6t
Xbit_r125_c86 bl[86] br[86] wl[125] vdd gnd cell_6t
Xbit_r126_c86 bl[86] br[86] wl[126] vdd gnd cell_6t
Xbit_r127_c86 bl[86] br[86] wl[127] vdd gnd cell_6t
Xbit_r0_c87 bl[87] br[87] wl[0] vdd gnd cell_6t
Xbit_r1_c87 bl[87] br[87] wl[1] vdd gnd cell_6t
Xbit_r2_c87 bl[87] br[87] wl[2] vdd gnd cell_6t
Xbit_r3_c87 bl[87] br[87] wl[3] vdd gnd cell_6t
Xbit_r4_c87 bl[87] br[87] wl[4] vdd gnd cell_6t
Xbit_r5_c87 bl[87] br[87] wl[5] vdd gnd cell_6t
Xbit_r6_c87 bl[87] br[87] wl[6] vdd gnd cell_6t
Xbit_r7_c87 bl[87] br[87] wl[7] vdd gnd cell_6t
Xbit_r8_c87 bl[87] br[87] wl[8] vdd gnd cell_6t
Xbit_r9_c87 bl[87] br[87] wl[9] vdd gnd cell_6t
Xbit_r10_c87 bl[87] br[87] wl[10] vdd gnd cell_6t
Xbit_r11_c87 bl[87] br[87] wl[11] vdd gnd cell_6t
Xbit_r12_c87 bl[87] br[87] wl[12] vdd gnd cell_6t
Xbit_r13_c87 bl[87] br[87] wl[13] vdd gnd cell_6t
Xbit_r14_c87 bl[87] br[87] wl[14] vdd gnd cell_6t
Xbit_r15_c87 bl[87] br[87] wl[15] vdd gnd cell_6t
Xbit_r16_c87 bl[87] br[87] wl[16] vdd gnd cell_6t
Xbit_r17_c87 bl[87] br[87] wl[17] vdd gnd cell_6t
Xbit_r18_c87 bl[87] br[87] wl[18] vdd gnd cell_6t
Xbit_r19_c87 bl[87] br[87] wl[19] vdd gnd cell_6t
Xbit_r20_c87 bl[87] br[87] wl[20] vdd gnd cell_6t
Xbit_r21_c87 bl[87] br[87] wl[21] vdd gnd cell_6t
Xbit_r22_c87 bl[87] br[87] wl[22] vdd gnd cell_6t
Xbit_r23_c87 bl[87] br[87] wl[23] vdd gnd cell_6t
Xbit_r24_c87 bl[87] br[87] wl[24] vdd gnd cell_6t
Xbit_r25_c87 bl[87] br[87] wl[25] vdd gnd cell_6t
Xbit_r26_c87 bl[87] br[87] wl[26] vdd gnd cell_6t
Xbit_r27_c87 bl[87] br[87] wl[27] vdd gnd cell_6t
Xbit_r28_c87 bl[87] br[87] wl[28] vdd gnd cell_6t
Xbit_r29_c87 bl[87] br[87] wl[29] vdd gnd cell_6t
Xbit_r30_c87 bl[87] br[87] wl[30] vdd gnd cell_6t
Xbit_r31_c87 bl[87] br[87] wl[31] vdd gnd cell_6t
Xbit_r32_c87 bl[87] br[87] wl[32] vdd gnd cell_6t
Xbit_r33_c87 bl[87] br[87] wl[33] vdd gnd cell_6t
Xbit_r34_c87 bl[87] br[87] wl[34] vdd gnd cell_6t
Xbit_r35_c87 bl[87] br[87] wl[35] vdd gnd cell_6t
Xbit_r36_c87 bl[87] br[87] wl[36] vdd gnd cell_6t
Xbit_r37_c87 bl[87] br[87] wl[37] vdd gnd cell_6t
Xbit_r38_c87 bl[87] br[87] wl[38] vdd gnd cell_6t
Xbit_r39_c87 bl[87] br[87] wl[39] vdd gnd cell_6t
Xbit_r40_c87 bl[87] br[87] wl[40] vdd gnd cell_6t
Xbit_r41_c87 bl[87] br[87] wl[41] vdd gnd cell_6t
Xbit_r42_c87 bl[87] br[87] wl[42] vdd gnd cell_6t
Xbit_r43_c87 bl[87] br[87] wl[43] vdd gnd cell_6t
Xbit_r44_c87 bl[87] br[87] wl[44] vdd gnd cell_6t
Xbit_r45_c87 bl[87] br[87] wl[45] vdd gnd cell_6t
Xbit_r46_c87 bl[87] br[87] wl[46] vdd gnd cell_6t
Xbit_r47_c87 bl[87] br[87] wl[47] vdd gnd cell_6t
Xbit_r48_c87 bl[87] br[87] wl[48] vdd gnd cell_6t
Xbit_r49_c87 bl[87] br[87] wl[49] vdd gnd cell_6t
Xbit_r50_c87 bl[87] br[87] wl[50] vdd gnd cell_6t
Xbit_r51_c87 bl[87] br[87] wl[51] vdd gnd cell_6t
Xbit_r52_c87 bl[87] br[87] wl[52] vdd gnd cell_6t
Xbit_r53_c87 bl[87] br[87] wl[53] vdd gnd cell_6t
Xbit_r54_c87 bl[87] br[87] wl[54] vdd gnd cell_6t
Xbit_r55_c87 bl[87] br[87] wl[55] vdd gnd cell_6t
Xbit_r56_c87 bl[87] br[87] wl[56] vdd gnd cell_6t
Xbit_r57_c87 bl[87] br[87] wl[57] vdd gnd cell_6t
Xbit_r58_c87 bl[87] br[87] wl[58] vdd gnd cell_6t
Xbit_r59_c87 bl[87] br[87] wl[59] vdd gnd cell_6t
Xbit_r60_c87 bl[87] br[87] wl[60] vdd gnd cell_6t
Xbit_r61_c87 bl[87] br[87] wl[61] vdd gnd cell_6t
Xbit_r62_c87 bl[87] br[87] wl[62] vdd gnd cell_6t
Xbit_r63_c87 bl[87] br[87] wl[63] vdd gnd cell_6t
Xbit_r64_c87 bl[87] br[87] wl[64] vdd gnd cell_6t
Xbit_r65_c87 bl[87] br[87] wl[65] vdd gnd cell_6t
Xbit_r66_c87 bl[87] br[87] wl[66] vdd gnd cell_6t
Xbit_r67_c87 bl[87] br[87] wl[67] vdd gnd cell_6t
Xbit_r68_c87 bl[87] br[87] wl[68] vdd gnd cell_6t
Xbit_r69_c87 bl[87] br[87] wl[69] vdd gnd cell_6t
Xbit_r70_c87 bl[87] br[87] wl[70] vdd gnd cell_6t
Xbit_r71_c87 bl[87] br[87] wl[71] vdd gnd cell_6t
Xbit_r72_c87 bl[87] br[87] wl[72] vdd gnd cell_6t
Xbit_r73_c87 bl[87] br[87] wl[73] vdd gnd cell_6t
Xbit_r74_c87 bl[87] br[87] wl[74] vdd gnd cell_6t
Xbit_r75_c87 bl[87] br[87] wl[75] vdd gnd cell_6t
Xbit_r76_c87 bl[87] br[87] wl[76] vdd gnd cell_6t
Xbit_r77_c87 bl[87] br[87] wl[77] vdd gnd cell_6t
Xbit_r78_c87 bl[87] br[87] wl[78] vdd gnd cell_6t
Xbit_r79_c87 bl[87] br[87] wl[79] vdd gnd cell_6t
Xbit_r80_c87 bl[87] br[87] wl[80] vdd gnd cell_6t
Xbit_r81_c87 bl[87] br[87] wl[81] vdd gnd cell_6t
Xbit_r82_c87 bl[87] br[87] wl[82] vdd gnd cell_6t
Xbit_r83_c87 bl[87] br[87] wl[83] vdd gnd cell_6t
Xbit_r84_c87 bl[87] br[87] wl[84] vdd gnd cell_6t
Xbit_r85_c87 bl[87] br[87] wl[85] vdd gnd cell_6t
Xbit_r86_c87 bl[87] br[87] wl[86] vdd gnd cell_6t
Xbit_r87_c87 bl[87] br[87] wl[87] vdd gnd cell_6t
Xbit_r88_c87 bl[87] br[87] wl[88] vdd gnd cell_6t
Xbit_r89_c87 bl[87] br[87] wl[89] vdd gnd cell_6t
Xbit_r90_c87 bl[87] br[87] wl[90] vdd gnd cell_6t
Xbit_r91_c87 bl[87] br[87] wl[91] vdd gnd cell_6t
Xbit_r92_c87 bl[87] br[87] wl[92] vdd gnd cell_6t
Xbit_r93_c87 bl[87] br[87] wl[93] vdd gnd cell_6t
Xbit_r94_c87 bl[87] br[87] wl[94] vdd gnd cell_6t
Xbit_r95_c87 bl[87] br[87] wl[95] vdd gnd cell_6t
Xbit_r96_c87 bl[87] br[87] wl[96] vdd gnd cell_6t
Xbit_r97_c87 bl[87] br[87] wl[97] vdd gnd cell_6t
Xbit_r98_c87 bl[87] br[87] wl[98] vdd gnd cell_6t
Xbit_r99_c87 bl[87] br[87] wl[99] vdd gnd cell_6t
Xbit_r100_c87 bl[87] br[87] wl[100] vdd gnd cell_6t
Xbit_r101_c87 bl[87] br[87] wl[101] vdd gnd cell_6t
Xbit_r102_c87 bl[87] br[87] wl[102] vdd gnd cell_6t
Xbit_r103_c87 bl[87] br[87] wl[103] vdd gnd cell_6t
Xbit_r104_c87 bl[87] br[87] wl[104] vdd gnd cell_6t
Xbit_r105_c87 bl[87] br[87] wl[105] vdd gnd cell_6t
Xbit_r106_c87 bl[87] br[87] wl[106] vdd gnd cell_6t
Xbit_r107_c87 bl[87] br[87] wl[107] vdd gnd cell_6t
Xbit_r108_c87 bl[87] br[87] wl[108] vdd gnd cell_6t
Xbit_r109_c87 bl[87] br[87] wl[109] vdd gnd cell_6t
Xbit_r110_c87 bl[87] br[87] wl[110] vdd gnd cell_6t
Xbit_r111_c87 bl[87] br[87] wl[111] vdd gnd cell_6t
Xbit_r112_c87 bl[87] br[87] wl[112] vdd gnd cell_6t
Xbit_r113_c87 bl[87] br[87] wl[113] vdd gnd cell_6t
Xbit_r114_c87 bl[87] br[87] wl[114] vdd gnd cell_6t
Xbit_r115_c87 bl[87] br[87] wl[115] vdd gnd cell_6t
Xbit_r116_c87 bl[87] br[87] wl[116] vdd gnd cell_6t
Xbit_r117_c87 bl[87] br[87] wl[117] vdd gnd cell_6t
Xbit_r118_c87 bl[87] br[87] wl[118] vdd gnd cell_6t
Xbit_r119_c87 bl[87] br[87] wl[119] vdd gnd cell_6t
Xbit_r120_c87 bl[87] br[87] wl[120] vdd gnd cell_6t
Xbit_r121_c87 bl[87] br[87] wl[121] vdd gnd cell_6t
Xbit_r122_c87 bl[87] br[87] wl[122] vdd gnd cell_6t
Xbit_r123_c87 bl[87] br[87] wl[123] vdd gnd cell_6t
Xbit_r124_c87 bl[87] br[87] wl[124] vdd gnd cell_6t
Xbit_r125_c87 bl[87] br[87] wl[125] vdd gnd cell_6t
Xbit_r126_c87 bl[87] br[87] wl[126] vdd gnd cell_6t
Xbit_r127_c87 bl[87] br[87] wl[127] vdd gnd cell_6t
Xbit_r0_c88 bl[88] br[88] wl[0] vdd gnd cell_6t
Xbit_r1_c88 bl[88] br[88] wl[1] vdd gnd cell_6t
Xbit_r2_c88 bl[88] br[88] wl[2] vdd gnd cell_6t
Xbit_r3_c88 bl[88] br[88] wl[3] vdd gnd cell_6t
Xbit_r4_c88 bl[88] br[88] wl[4] vdd gnd cell_6t
Xbit_r5_c88 bl[88] br[88] wl[5] vdd gnd cell_6t
Xbit_r6_c88 bl[88] br[88] wl[6] vdd gnd cell_6t
Xbit_r7_c88 bl[88] br[88] wl[7] vdd gnd cell_6t
Xbit_r8_c88 bl[88] br[88] wl[8] vdd gnd cell_6t
Xbit_r9_c88 bl[88] br[88] wl[9] vdd gnd cell_6t
Xbit_r10_c88 bl[88] br[88] wl[10] vdd gnd cell_6t
Xbit_r11_c88 bl[88] br[88] wl[11] vdd gnd cell_6t
Xbit_r12_c88 bl[88] br[88] wl[12] vdd gnd cell_6t
Xbit_r13_c88 bl[88] br[88] wl[13] vdd gnd cell_6t
Xbit_r14_c88 bl[88] br[88] wl[14] vdd gnd cell_6t
Xbit_r15_c88 bl[88] br[88] wl[15] vdd gnd cell_6t
Xbit_r16_c88 bl[88] br[88] wl[16] vdd gnd cell_6t
Xbit_r17_c88 bl[88] br[88] wl[17] vdd gnd cell_6t
Xbit_r18_c88 bl[88] br[88] wl[18] vdd gnd cell_6t
Xbit_r19_c88 bl[88] br[88] wl[19] vdd gnd cell_6t
Xbit_r20_c88 bl[88] br[88] wl[20] vdd gnd cell_6t
Xbit_r21_c88 bl[88] br[88] wl[21] vdd gnd cell_6t
Xbit_r22_c88 bl[88] br[88] wl[22] vdd gnd cell_6t
Xbit_r23_c88 bl[88] br[88] wl[23] vdd gnd cell_6t
Xbit_r24_c88 bl[88] br[88] wl[24] vdd gnd cell_6t
Xbit_r25_c88 bl[88] br[88] wl[25] vdd gnd cell_6t
Xbit_r26_c88 bl[88] br[88] wl[26] vdd gnd cell_6t
Xbit_r27_c88 bl[88] br[88] wl[27] vdd gnd cell_6t
Xbit_r28_c88 bl[88] br[88] wl[28] vdd gnd cell_6t
Xbit_r29_c88 bl[88] br[88] wl[29] vdd gnd cell_6t
Xbit_r30_c88 bl[88] br[88] wl[30] vdd gnd cell_6t
Xbit_r31_c88 bl[88] br[88] wl[31] vdd gnd cell_6t
Xbit_r32_c88 bl[88] br[88] wl[32] vdd gnd cell_6t
Xbit_r33_c88 bl[88] br[88] wl[33] vdd gnd cell_6t
Xbit_r34_c88 bl[88] br[88] wl[34] vdd gnd cell_6t
Xbit_r35_c88 bl[88] br[88] wl[35] vdd gnd cell_6t
Xbit_r36_c88 bl[88] br[88] wl[36] vdd gnd cell_6t
Xbit_r37_c88 bl[88] br[88] wl[37] vdd gnd cell_6t
Xbit_r38_c88 bl[88] br[88] wl[38] vdd gnd cell_6t
Xbit_r39_c88 bl[88] br[88] wl[39] vdd gnd cell_6t
Xbit_r40_c88 bl[88] br[88] wl[40] vdd gnd cell_6t
Xbit_r41_c88 bl[88] br[88] wl[41] vdd gnd cell_6t
Xbit_r42_c88 bl[88] br[88] wl[42] vdd gnd cell_6t
Xbit_r43_c88 bl[88] br[88] wl[43] vdd gnd cell_6t
Xbit_r44_c88 bl[88] br[88] wl[44] vdd gnd cell_6t
Xbit_r45_c88 bl[88] br[88] wl[45] vdd gnd cell_6t
Xbit_r46_c88 bl[88] br[88] wl[46] vdd gnd cell_6t
Xbit_r47_c88 bl[88] br[88] wl[47] vdd gnd cell_6t
Xbit_r48_c88 bl[88] br[88] wl[48] vdd gnd cell_6t
Xbit_r49_c88 bl[88] br[88] wl[49] vdd gnd cell_6t
Xbit_r50_c88 bl[88] br[88] wl[50] vdd gnd cell_6t
Xbit_r51_c88 bl[88] br[88] wl[51] vdd gnd cell_6t
Xbit_r52_c88 bl[88] br[88] wl[52] vdd gnd cell_6t
Xbit_r53_c88 bl[88] br[88] wl[53] vdd gnd cell_6t
Xbit_r54_c88 bl[88] br[88] wl[54] vdd gnd cell_6t
Xbit_r55_c88 bl[88] br[88] wl[55] vdd gnd cell_6t
Xbit_r56_c88 bl[88] br[88] wl[56] vdd gnd cell_6t
Xbit_r57_c88 bl[88] br[88] wl[57] vdd gnd cell_6t
Xbit_r58_c88 bl[88] br[88] wl[58] vdd gnd cell_6t
Xbit_r59_c88 bl[88] br[88] wl[59] vdd gnd cell_6t
Xbit_r60_c88 bl[88] br[88] wl[60] vdd gnd cell_6t
Xbit_r61_c88 bl[88] br[88] wl[61] vdd gnd cell_6t
Xbit_r62_c88 bl[88] br[88] wl[62] vdd gnd cell_6t
Xbit_r63_c88 bl[88] br[88] wl[63] vdd gnd cell_6t
Xbit_r64_c88 bl[88] br[88] wl[64] vdd gnd cell_6t
Xbit_r65_c88 bl[88] br[88] wl[65] vdd gnd cell_6t
Xbit_r66_c88 bl[88] br[88] wl[66] vdd gnd cell_6t
Xbit_r67_c88 bl[88] br[88] wl[67] vdd gnd cell_6t
Xbit_r68_c88 bl[88] br[88] wl[68] vdd gnd cell_6t
Xbit_r69_c88 bl[88] br[88] wl[69] vdd gnd cell_6t
Xbit_r70_c88 bl[88] br[88] wl[70] vdd gnd cell_6t
Xbit_r71_c88 bl[88] br[88] wl[71] vdd gnd cell_6t
Xbit_r72_c88 bl[88] br[88] wl[72] vdd gnd cell_6t
Xbit_r73_c88 bl[88] br[88] wl[73] vdd gnd cell_6t
Xbit_r74_c88 bl[88] br[88] wl[74] vdd gnd cell_6t
Xbit_r75_c88 bl[88] br[88] wl[75] vdd gnd cell_6t
Xbit_r76_c88 bl[88] br[88] wl[76] vdd gnd cell_6t
Xbit_r77_c88 bl[88] br[88] wl[77] vdd gnd cell_6t
Xbit_r78_c88 bl[88] br[88] wl[78] vdd gnd cell_6t
Xbit_r79_c88 bl[88] br[88] wl[79] vdd gnd cell_6t
Xbit_r80_c88 bl[88] br[88] wl[80] vdd gnd cell_6t
Xbit_r81_c88 bl[88] br[88] wl[81] vdd gnd cell_6t
Xbit_r82_c88 bl[88] br[88] wl[82] vdd gnd cell_6t
Xbit_r83_c88 bl[88] br[88] wl[83] vdd gnd cell_6t
Xbit_r84_c88 bl[88] br[88] wl[84] vdd gnd cell_6t
Xbit_r85_c88 bl[88] br[88] wl[85] vdd gnd cell_6t
Xbit_r86_c88 bl[88] br[88] wl[86] vdd gnd cell_6t
Xbit_r87_c88 bl[88] br[88] wl[87] vdd gnd cell_6t
Xbit_r88_c88 bl[88] br[88] wl[88] vdd gnd cell_6t
Xbit_r89_c88 bl[88] br[88] wl[89] vdd gnd cell_6t
Xbit_r90_c88 bl[88] br[88] wl[90] vdd gnd cell_6t
Xbit_r91_c88 bl[88] br[88] wl[91] vdd gnd cell_6t
Xbit_r92_c88 bl[88] br[88] wl[92] vdd gnd cell_6t
Xbit_r93_c88 bl[88] br[88] wl[93] vdd gnd cell_6t
Xbit_r94_c88 bl[88] br[88] wl[94] vdd gnd cell_6t
Xbit_r95_c88 bl[88] br[88] wl[95] vdd gnd cell_6t
Xbit_r96_c88 bl[88] br[88] wl[96] vdd gnd cell_6t
Xbit_r97_c88 bl[88] br[88] wl[97] vdd gnd cell_6t
Xbit_r98_c88 bl[88] br[88] wl[98] vdd gnd cell_6t
Xbit_r99_c88 bl[88] br[88] wl[99] vdd gnd cell_6t
Xbit_r100_c88 bl[88] br[88] wl[100] vdd gnd cell_6t
Xbit_r101_c88 bl[88] br[88] wl[101] vdd gnd cell_6t
Xbit_r102_c88 bl[88] br[88] wl[102] vdd gnd cell_6t
Xbit_r103_c88 bl[88] br[88] wl[103] vdd gnd cell_6t
Xbit_r104_c88 bl[88] br[88] wl[104] vdd gnd cell_6t
Xbit_r105_c88 bl[88] br[88] wl[105] vdd gnd cell_6t
Xbit_r106_c88 bl[88] br[88] wl[106] vdd gnd cell_6t
Xbit_r107_c88 bl[88] br[88] wl[107] vdd gnd cell_6t
Xbit_r108_c88 bl[88] br[88] wl[108] vdd gnd cell_6t
Xbit_r109_c88 bl[88] br[88] wl[109] vdd gnd cell_6t
Xbit_r110_c88 bl[88] br[88] wl[110] vdd gnd cell_6t
Xbit_r111_c88 bl[88] br[88] wl[111] vdd gnd cell_6t
Xbit_r112_c88 bl[88] br[88] wl[112] vdd gnd cell_6t
Xbit_r113_c88 bl[88] br[88] wl[113] vdd gnd cell_6t
Xbit_r114_c88 bl[88] br[88] wl[114] vdd gnd cell_6t
Xbit_r115_c88 bl[88] br[88] wl[115] vdd gnd cell_6t
Xbit_r116_c88 bl[88] br[88] wl[116] vdd gnd cell_6t
Xbit_r117_c88 bl[88] br[88] wl[117] vdd gnd cell_6t
Xbit_r118_c88 bl[88] br[88] wl[118] vdd gnd cell_6t
Xbit_r119_c88 bl[88] br[88] wl[119] vdd gnd cell_6t
Xbit_r120_c88 bl[88] br[88] wl[120] vdd gnd cell_6t
Xbit_r121_c88 bl[88] br[88] wl[121] vdd gnd cell_6t
Xbit_r122_c88 bl[88] br[88] wl[122] vdd gnd cell_6t
Xbit_r123_c88 bl[88] br[88] wl[123] vdd gnd cell_6t
Xbit_r124_c88 bl[88] br[88] wl[124] vdd gnd cell_6t
Xbit_r125_c88 bl[88] br[88] wl[125] vdd gnd cell_6t
Xbit_r126_c88 bl[88] br[88] wl[126] vdd gnd cell_6t
Xbit_r127_c88 bl[88] br[88] wl[127] vdd gnd cell_6t
Xbit_r0_c89 bl[89] br[89] wl[0] vdd gnd cell_6t
Xbit_r1_c89 bl[89] br[89] wl[1] vdd gnd cell_6t
Xbit_r2_c89 bl[89] br[89] wl[2] vdd gnd cell_6t
Xbit_r3_c89 bl[89] br[89] wl[3] vdd gnd cell_6t
Xbit_r4_c89 bl[89] br[89] wl[4] vdd gnd cell_6t
Xbit_r5_c89 bl[89] br[89] wl[5] vdd gnd cell_6t
Xbit_r6_c89 bl[89] br[89] wl[6] vdd gnd cell_6t
Xbit_r7_c89 bl[89] br[89] wl[7] vdd gnd cell_6t
Xbit_r8_c89 bl[89] br[89] wl[8] vdd gnd cell_6t
Xbit_r9_c89 bl[89] br[89] wl[9] vdd gnd cell_6t
Xbit_r10_c89 bl[89] br[89] wl[10] vdd gnd cell_6t
Xbit_r11_c89 bl[89] br[89] wl[11] vdd gnd cell_6t
Xbit_r12_c89 bl[89] br[89] wl[12] vdd gnd cell_6t
Xbit_r13_c89 bl[89] br[89] wl[13] vdd gnd cell_6t
Xbit_r14_c89 bl[89] br[89] wl[14] vdd gnd cell_6t
Xbit_r15_c89 bl[89] br[89] wl[15] vdd gnd cell_6t
Xbit_r16_c89 bl[89] br[89] wl[16] vdd gnd cell_6t
Xbit_r17_c89 bl[89] br[89] wl[17] vdd gnd cell_6t
Xbit_r18_c89 bl[89] br[89] wl[18] vdd gnd cell_6t
Xbit_r19_c89 bl[89] br[89] wl[19] vdd gnd cell_6t
Xbit_r20_c89 bl[89] br[89] wl[20] vdd gnd cell_6t
Xbit_r21_c89 bl[89] br[89] wl[21] vdd gnd cell_6t
Xbit_r22_c89 bl[89] br[89] wl[22] vdd gnd cell_6t
Xbit_r23_c89 bl[89] br[89] wl[23] vdd gnd cell_6t
Xbit_r24_c89 bl[89] br[89] wl[24] vdd gnd cell_6t
Xbit_r25_c89 bl[89] br[89] wl[25] vdd gnd cell_6t
Xbit_r26_c89 bl[89] br[89] wl[26] vdd gnd cell_6t
Xbit_r27_c89 bl[89] br[89] wl[27] vdd gnd cell_6t
Xbit_r28_c89 bl[89] br[89] wl[28] vdd gnd cell_6t
Xbit_r29_c89 bl[89] br[89] wl[29] vdd gnd cell_6t
Xbit_r30_c89 bl[89] br[89] wl[30] vdd gnd cell_6t
Xbit_r31_c89 bl[89] br[89] wl[31] vdd gnd cell_6t
Xbit_r32_c89 bl[89] br[89] wl[32] vdd gnd cell_6t
Xbit_r33_c89 bl[89] br[89] wl[33] vdd gnd cell_6t
Xbit_r34_c89 bl[89] br[89] wl[34] vdd gnd cell_6t
Xbit_r35_c89 bl[89] br[89] wl[35] vdd gnd cell_6t
Xbit_r36_c89 bl[89] br[89] wl[36] vdd gnd cell_6t
Xbit_r37_c89 bl[89] br[89] wl[37] vdd gnd cell_6t
Xbit_r38_c89 bl[89] br[89] wl[38] vdd gnd cell_6t
Xbit_r39_c89 bl[89] br[89] wl[39] vdd gnd cell_6t
Xbit_r40_c89 bl[89] br[89] wl[40] vdd gnd cell_6t
Xbit_r41_c89 bl[89] br[89] wl[41] vdd gnd cell_6t
Xbit_r42_c89 bl[89] br[89] wl[42] vdd gnd cell_6t
Xbit_r43_c89 bl[89] br[89] wl[43] vdd gnd cell_6t
Xbit_r44_c89 bl[89] br[89] wl[44] vdd gnd cell_6t
Xbit_r45_c89 bl[89] br[89] wl[45] vdd gnd cell_6t
Xbit_r46_c89 bl[89] br[89] wl[46] vdd gnd cell_6t
Xbit_r47_c89 bl[89] br[89] wl[47] vdd gnd cell_6t
Xbit_r48_c89 bl[89] br[89] wl[48] vdd gnd cell_6t
Xbit_r49_c89 bl[89] br[89] wl[49] vdd gnd cell_6t
Xbit_r50_c89 bl[89] br[89] wl[50] vdd gnd cell_6t
Xbit_r51_c89 bl[89] br[89] wl[51] vdd gnd cell_6t
Xbit_r52_c89 bl[89] br[89] wl[52] vdd gnd cell_6t
Xbit_r53_c89 bl[89] br[89] wl[53] vdd gnd cell_6t
Xbit_r54_c89 bl[89] br[89] wl[54] vdd gnd cell_6t
Xbit_r55_c89 bl[89] br[89] wl[55] vdd gnd cell_6t
Xbit_r56_c89 bl[89] br[89] wl[56] vdd gnd cell_6t
Xbit_r57_c89 bl[89] br[89] wl[57] vdd gnd cell_6t
Xbit_r58_c89 bl[89] br[89] wl[58] vdd gnd cell_6t
Xbit_r59_c89 bl[89] br[89] wl[59] vdd gnd cell_6t
Xbit_r60_c89 bl[89] br[89] wl[60] vdd gnd cell_6t
Xbit_r61_c89 bl[89] br[89] wl[61] vdd gnd cell_6t
Xbit_r62_c89 bl[89] br[89] wl[62] vdd gnd cell_6t
Xbit_r63_c89 bl[89] br[89] wl[63] vdd gnd cell_6t
Xbit_r64_c89 bl[89] br[89] wl[64] vdd gnd cell_6t
Xbit_r65_c89 bl[89] br[89] wl[65] vdd gnd cell_6t
Xbit_r66_c89 bl[89] br[89] wl[66] vdd gnd cell_6t
Xbit_r67_c89 bl[89] br[89] wl[67] vdd gnd cell_6t
Xbit_r68_c89 bl[89] br[89] wl[68] vdd gnd cell_6t
Xbit_r69_c89 bl[89] br[89] wl[69] vdd gnd cell_6t
Xbit_r70_c89 bl[89] br[89] wl[70] vdd gnd cell_6t
Xbit_r71_c89 bl[89] br[89] wl[71] vdd gnd cell_6t
Xbit_r72_c89 bl[89] br[89] wl[72] vdd gnd cell_6t
Xbit_r73_c89 bl[89] br[89] wl[73] vdd gnd cell_6t
Xbit_r74_c89 bl[89] br[89] wl[74] vdd gnd cell_6t
Xbit_r75_c89 bl[89] br[89] wl[75] vdd gnd cell_6t
Xbit_r76_c89 bl[89] br[89] wl[76] vdd gnd cell_6t
Xbit_r77_c89 bl[89] br[89] wl[77] vdd gnd cell_6t
Xbit_r78_c89 bl[89] br[89] wl[78] vdd gnd cell_6t
Xbit_r79_c89 bl[89] br[89] wl[79] vdd gnd cell_6t
Xbit_r80_c89 bl[89] br[89] wl[80] vdd gnd cell_6t
Xbit_r81_c89 bl[89] br[89] wl[81] vdd gnd cell_6t
Xbit_r82_c89 bl[89] br[89] wl[82] vdd gnd cell_6t
Xbit_r83_c89 bl[89] br[89] wl[83] vdd gnd cell_6t
Xbit_r84_c89 bl[89] br[89] wl[84] vdd gnd cell_6t
Xbit_r85_c89 bl[89] br[89] wl[85] vdd gnd cell_6t
Xbit_r86_c89 bl[89] br[89] wl[86] vdd gnd cell_6t
Xbit_r87_c89 bl[89] br[89] wl[87] vdd gnd cell_6t
Xbit_r88_c89 bl[89] br[89] wl[88] vdd gnd cell_6t
Xbit_r89_c89 bl[89] br[89] wl[89] vdd gnd cell_6t
Xbit_r90_c89 bl[89] br[89] wl[90] vdd gnd cell_6t
Xbit_r91_c89 bl[89] br[89] wl[91] vdd gnd cell_6t
Xbit_r92_c89 bl[89] br[89] wl[92] vdd gnd cell_6t
Xbit_r93_c89 bl[89] br[89] wl[93] vdd gnd cell_6t
Xbit_r94_c89 bl[89] br[89] wl[94] vdd gnd cell_6t
Xbit_r95_c89 bl[89] br[89] wl[95] vdd gnd cell_6t
Xbit_r96_c89 bl[89] br[89] wl[96] vdd gnd cell_6t
Xbit_r97_c89 bl[89] br[89] wl[97] vdd gnd cell_6t
Xbit_r98_c89 bl[89] br[89] wl[98] vdd gnd cell_6t
Xbit_r99_c89 bl[89] br[89] wl[99] vdd gnd cell_6t
Xbit_r100_c89 bl[89] br[89] wl[100] vdd gnd cell_6t
Xbit_r101_c89 bl[89] br[89] wl[101] vdd gnd cell_6t
Xbit_r102_c89 bl[89] br[89] wl[102] vdd gnd cell_6t
Xbit_r103_c89 bl[89] br[89] wl[103] vdd gnd cell_6t
Xbit_r104_c89 bl[89] br[89] wl[104] vdd gnd cell_6t
Xbit_r105_c89 bl[89] br[89] wl[105] vdd gnd cell_6t
Xbit_r106_c89 bl[89] br[89] wl[106] vdd gnd cell_6t
Xbit_r107_c89 bl[89] br[89] wl[107] vdd gnd cell_6t
Xbit_r108_c89 bl[89] br[89] wl[108] vdd gnd cell_6t
Xbit_r109_c89 bl[89] br[89] wl[109] vdd gnd cell_6t
Xbit_r110_c89 bl[89] br[89] wl[110] vdd gnd cell_6t
Xbit_r111_c89 bl[89] br[89] wl[111] vdd gnd cell_6t
Xbit_r112_c89 bl[89] br[89] wl[112] vdd gnd cell_6t
Xbit_r113_c89 bl[89] br[89] wl[113] vdd gnd cell_6t
Xbit_r114_c89 bl[89] br[89] wl[114] vdd gnd cell_6t
Xbit_r115_c89 bl[89] br[89] wl[115] vdd gnd cell_6t
Xbit_r116_c89 bl[89] br[89] wl[116] vdd gnd cell_6t
Xbit_r117_c89 bl[89] br[89] wl[117] vdd gnd cell_6t
Xbit_r118_c89 bl[89] br[89] wl[118] vdd gnd cell_6t
Xbit_r119_c89 bl[89] br[89] wl[119] vdd gnd cell_6t
Xbit_r120_c89 bl[89] br[89] wl[120] vdd gnd cell_6t
Xbit_r121_c89 bl[89] br[89] wl[121] vdd gnd cell_6t
Xbit_r122_c89 bl[89] br[89] wl[122] vdd gnd cell_6t
Xbit_r123_c89 bl[89] br[89] wl[123] vdd gnd cell_6t
Xbit_r124_c89 bl[89] br[89] wl[124] vdd gnd cell_6t
Xbit_r125_c89 bl[89] br[89] wl[125] vdd gnd cell_6t
Xbit_r126_c89 bl[89] br[89] wl[126] vdd gnd cell_6t
Xbit_r127_c89 bl[89] br[89] wl[127] vdd gnd cell_6t
Xbit_r0_c90 bl[90] br[90] wl[0] vdd gnd cell_6t
Xbit_r1_c90 bl[90] br[90] wl[1] vdd gnd cell_6t
Xbit_r2_c90 bl[90] br[90] wl[2] vdd gnd cell_6t
Xbit_r3_c90 bl[90] br[90] wl[3] vdd gnd cell_6t
Xbit_r4_c90 bl[90] br[90] wl[4] vdd gnd cell_6t
Xbit_r5_c90 bl[90] br[90] wl[5] vdd gnd cell_6t
Xbit_r6_c90 bl[90] br[90] wl[6] vdd gnd cell_6t
Xbit_r7_c90 bl[90] br[90] wl[7] vdd gnd cell_6t
Xbit_r8_c90 bl[90] br[90] wl[8] vdd gnd cell_6t
Xbit_r9_c90 bl[90] br[90] wl[9] vdd gnd cell_6t
Xbit_r10_c90 bl[90] br[90] wl[10] vdd gnd cell_6t
Xbit_r11_c90 bl[90] br[90] wl[11] vdd gnd cell_6t
Xbit_r12_c90 bl[90] br[90] wl[12] vdd gnd cell_6t
Xbit_r13_c90 bl[90] br[90] wl[13] vdd gnd cell_6t
Xbit_r14_c90 bl[90] br[90] wl[14] vdd gnd cell_6t
Xbit_r15_c90 bl[90] br[90] wl[15] vdd gnd cell_6t
Xbit_r16_c90 bl[90] br[90] wl[16] vdd gnd cell_6t
Xbit_r17_c90 bl[90] br[90] wl[17] vdd gnd cell_6t
Xbit_r18_c90 bl[90] br[90] wl[18] vdd gnd cell_6t
Xbit_r19_c90 bl[90] br[90] wl[19] vdd gnd cell_6t
Xbit_r20_c90 bl[90] br[90] wl[20] vdd gnd cell_6t
Xbit_r21_c90 bl[90] br[90] wl[21] vdd gnd cell_6t
Xbit_r22_c90 bl[90] br[90] wl[22] vdd gnd cell_6t
Xbit_r23_c90 bl[90] br[90] wl[23] vdd gnd cell_6t
Xbit_r24_c90 bl[90] br[90] wl[24] vdd gnd cell_6t
Xbit_r25_c90 bl[90] br[90] wl[25] vdd gnd cell_6t
Xbit_r26_c90 bl[90] br[90] wl[26] vdd gnd cell_6t
Xbit_r27_c90 bl[90] br[90] wl[27] vdd gnd cell_6t
Xbit_r28_c90 bl[90] br[90] wl[28] vdd gnd cell_6t
Xbit_r29_c90 bl[90] br[90] wl[29] vdd gnd cell_6t
Xbit_r30_c90 bl[90] br[90] wl[30] vdd gnd cell_6t
Xbit_r31_c90 bl[90] br[90] wl[31] vdd gnd cell_6t
Xbit_r32_c90 bl[90] br[90] wl[32] vdd gnd cell_6t
Xbit_r33_c90 bl[90] br[90] wl[33] vdd gnd cell_6t
Xbit_r34_c90 bl[90] br[90] wl[34] vdd gnd cell_6t
Xbit_r35_c90 bl[90] br[90] wl[35] vdd gnd cell_6t
Xbit_r36_c90 bl[90] br[90] wl[36] vdd gnd cell_6t
Xbit_r37_c90 bl[90] br[90] wl[37] vdd gnd cell_6t
Xbit_r38_c90 bl[90] br[90] wl[38] vdd gnd cell_6t
Xbit_r39_c90 bl[90] br[90] wl[39] vdd gnd cell_6t
Xbit_r40_c90 bl[90] br[90] wl[40] vdd gnd cell_6t
Xbit_r41_c90 bl[90] br[90] wl[41] vdd gnd cell_6t
Xbit_r42_c90 bl[90] br[90] wl[42] vdd gnd cell_6t
Xbit_r43_c90 bl[90] br[90] wl[43] vdd gnd cell_6t
Xbit_r44_c90 bl[90] br[90] wl[44] vdd gnd cell_6t
Xbit_r45_c90 bl[90] br[90] wl[45] vdd gnd cell_6t
Xbit_r46_c90 bl[90] br[90] wl[46] vdd gnd cell_6t
Xbit_r47_c90 bl[90] br[90] wl[47] vdd gnd cell_6t
Xbit_r48_c90 bl[90] br[90] wl[48] vdd gnd cell_6t
Xbit_r49_c90 bl[90] br[90] wl[49] vdd gnd cell_6t
Xbit_r50_c90 bl[90] br[90] wl[50] vdd gnd cell_6t
Xbit_r51_c90 bl[90] br[90] wl[51] vdd gnd cell_6t
Xbit_r52_c90 bl[90] br[90] wl[52] vdd gnd cell_6t
Xbit_r53_c90 bl[90] br[90] wl[53] vdd gnd cell_6t
Xbit_r54_c90 bl[90] br[90] wl[54] vdd gnd cell_6t
Xbit_r55_c90 bl[90] br[90] wl[55] vdd gnd cell_6t
Xbit_r56_c90 bl[90] br[90] wl[56] vdd gnd cell_6t
Xbit_r57_c90 bl[90] br[90] wl[57] vdd gnd cell_6t
Xbit_r58_c90 bl[90] br[90] wl[58] vdd gnd cell_6t
Xbit_r59_c90 bl[90] br[90] wl[59] vdd gnd cell_6t
Xbit_r60_c90 bl[90] br[90] wl[60] vdd gnd cell_6t
Xbit_r61_c90 bl[90] br[90] wl[61] vdd gnd cell_6t
Xbit_r62_c90 bl[90] br[90] wl[62] vdd gnd cell_6t
Xbit_r63_c90 bl[90] br[90] wl[63] vdd gnd cell_6t
Xbit_r64_c90 bl[90] br[90] wl[64] vdd gnd cell_6t
Xbit_r65_c90 bl[90] br[90] wl[65] vdd gnd cell_6t
Xbit_r66_c90 bl[90] br[90] wl[66] vdd gnd cell_6t
Xbit_r67_c90 bl[90] br[90] wl[67] vdd gnd cell_6t
Xbit_r68_c90 bl[90] br[90] wl[68] vdd gnd cell_6t
Xbit_r69_c90 bl[90] br[90] wl[69] vdd gnd cell_6t
Xbit_r70_c90 bl[90] br[90] wl[70] vdd gnd cell_6t
Xbit_r71_c90 bl[90] br[90] wl[71] vdd gnd cell_6t
Xbit_r72_c90 bl[90] br[90] wl[72] vdd gnd cell_6t
Xbit_r73_c90 bl[90] br[90] wl[73] vdd gnd cell_6t
Xbit_r74_c90 bl[90] br[90] wl[74] vdd gnd cell_6t
Xbit_r75_c90 bl[90] br[90] wl[75] vdd gnd cell_6t
Xbit_r76_c90 bl[90] br[90] wl[76] vdd gnd cell_6t
Xbit_r77_c90 bl[90] br[90] wl[77] vdd gnd cell_6t
Xbit_r78_c90 bl[90] br[90] wl[78] vdd gnd cell_6t
Xbit_r79_c90 bl[90] br[90] wl[79] vdd gnd cell_6t
Xbit_r80_c90 bl[90] br[90] wl[80] vdd gnd cell_6t
Xbit_r81_c90 bl[90] br[90] wl[81] vdd gnd cell_6t
Xbit_r82_c90 bl[90] br[90] wl[82] vdd gnd cell_6t
Xbit_r83_c90 bl[90] br[90] wl[83] vdd gnd cell_6t
Xbit_r84_c90 bl[90] br[90] wl[84] vdd gnd cell_6t
Xbit_r85_c90 bl[90] br[90] wl[85] vdd gnd cell_6t
Xbit_r86_c90 bl[90] br[90] wl[86] vdd gnd cell_6t
Xbit_r87_c90 bl[90] br[90] wl[87] vdd gnd cell_6t
Xbit_r88_c90 bl[90] br[90] wl[88] vdd gnd cell_6t
Xbit_r89_c90 bl[90] br[90] wl[89] vdd gnd cell_6t
Xbit_r90_c90 bl[90] br[90] wl[90] vdd gnd cell_6t
Xbit_r91_c90 bl[90] br[90] wl[91] vdd gnd cell_6t
Xbit_r92_c90 bl[90] br[90] wl[92] vdd gnd cell_6t
Xbit_r93_c90 bl[90] br[90] wl[93] vdd gnd cell_6t
Xbit_r94_c90 bl[90] br[90] wl[94] vdd gnd cell_6t
Xbit_r95_c90 bl[90] br[90] wl[95] vdd gnd cell_6t
Xbit_r96_c90 bl[90] br[90] wl[96] vdd gnd cell_6t
Xbit_r97_c90 bl[90] br[90] wl[97] vdd gnd cell_6t
Xbit_r98_c90 bl[90] br[90] wl[98] vdd gnd cell_6t
Xbit_r99_c90 bl[90] br[90] wl[99] vdd gnd cell_6t
Xbit_r100_c90 bl[90] br[90] wl[100] vdd gnd cell_6t
Xbit_r101_c90 bl[90] br[90] wl[101] vdd gnd cell_6t
Xbit_r102_c90 bl[90] br[90] wl[102] vdd gnd cell_6t
Xbit_r103_c90 bl[90] br[90] wl[103] vdd gnd cell_6t
Xbit_r104_c90 bl[90] br[90] wl[104] vdd gnd cell_6t
Xbit_r105_c90 bl[90] br[90] wl[105] vdd gnd cell_6t
Xbit_r106_c90 bl[90] br[90] wl[106] vdd gnd cell_6t
Xbit_r107_c90 bl[90] br[90] wl[107] vdd gnd cell_6t
Xbit_r108_c90 bl[90] br[90] wl[108] vdd gnd cell_6t
Xbit_r109_c90 bl[90] br[90] wl[109] vdd gnd cell_6t
Xbit_r110_c90 bl[90] br[90] wl[110] vdd gnd cell_6t
Xbit_r111_c90 bl[90] br[90] wl[111] vdd gnd cell_6t
Xbit_r112_c90 bl[90] br[90] wl[112] vdd gnd cell_6t
Xbit_r113_c90 bl[90] br[90] wl[113] vdd gnd cell_6t
Xbit_r114_c90 bl[90] br[90] wl[114] vdd gnd cell_6t
Xbit_r115_c90 bl[90] br[90] wl[115] vdd gnd cell_6t
Xbit_r116_c90 bl[90] br[90] wl[116] vdd gnd cell_6t
Xbit_r117_c90 bl[90] br[90] wl[117] vdd gnd cell_6t
Xbit_r118_c90 bl[90] br[90] wl[118] vdd gnd cell_6t
Xbit_r119_c90 bl[90] br[90] wl[119] vdd gnd cell_6t
Xbit_r120_c90 bl[90] br[90] wl[120] vdd gnd cell_6t
Xbit_r121_c90 bl[90] br[90] wl[121] vdd gnd cell_6t
Xbit_r122_c90 bl[90] br[90] wl[122] vdd gnd cell_6t
Xbit_r123_c90 bl[90] br[90] wl[123] vdd gnd cell_6t
Xbit_r124_c90 bl[90] br[90] wl[124] vdd gnd cell_6t
Xbit_r125_c90 bl[90] br[90] wl[125] vdd gnd cell_6t
Xbit_r126_c90 bl[90] br[90] wl[126] vdd gnd cell_6t
Xbit_r127_c90 bl[90] br[90] wl[127] vdd gnd cell_6t
Xbit_r0_c91 bl[91] br[91] wl[0] vdd gnd cell_6t
Xbit_r1_c91 bl[91] br[91] wl[1] vdd gnd cell_6t
Xbit_r2_c91 bl[91] br[91] wl[2] vdd gnd cell_6t
Xbit_r3_c91 bl[91] br[91] wl[3] vdd gnd cell_6t
Xbit_r4_c91 bl[91] br[91] wl[4] vdd gnd cell_6t
Xbit_r5_c91 bl[91] br[91] wl[5] vdd gnd cell_6t
Xbit_r6_c91 bl[91] br[91] wl[6] vdd gnd cell_6t
Xbit_r7_c91 bl[91] br[91] wl[7] vdd gnd cell_6t
Xbit_r8_c91 bl[91] br[91] wl[8] vdd gnd cell_6t
Xbit_r9_c91 bl[91] br[91] wl[9] vdd gnd cell_6t
Xbit_r10_c91 bl[91] br[91] wl[10] vdd gnd cell_6t
Xbit_r11_c91 bl[91] br[91] wl[11] vdd gnd cell_6t
Xbit_r12_c91 bl[91] br[91] wl[12] vdd gnd cell_6t
Xbit_r13_c91 bl[91] br[91] wl[13] vdd gnd cell_6t
Xbit_r14_c91 bl[91] br[91] wl[14] vdd gnd cell_6t
Xbit_r15_c91 bl[91] br[91] wl[15] vdd gnd cell_6t
Xbit_r16_c91 bl[91] br[91] wl[16] vdd gnd cell_6t
Xbit_r17_c91 bl[91] br[91] wl[17] vdd gnd cell_6t
Xbit_r18_c91 bl[91] br[91] wl[18] vdd gnd cell_6t
Xbit_r19_c91 bl[91] br[91] wl[19] vdd gnd cell_6t
Xbit_r20_c91 bl[91] br[91] wl[20] vdd gnd cell_6t
Xbit_r21_c91 bl[91] br[91] wl[21] vdd gnd cell_6t
Xbit_r22_c91 bl[91] br[91] wl[22] vdd gnd cell_6t
Xbit_r23_c91 bl[91] br[91] wl[23] vdd gnd cell_6t
Xbit_r24_c91 bl[91] br[91] wl[24] vdd gnd cell_6t
Xbit_r25_c91 bl[91] br[91] wl[25] vdd gnd cell_6t
Xbit_r26_c91 bl[91] br[91] wl[26] vdd gnd cell_6t
Xbit_r27_c91 bl[91] br[91] wl[27] vdd gnd cell_6t
Xbit_r28_c91 bl[91] br[91] wl[28] vdd gnd cell_6t
Xbit_r29_c91 bl[91] br[91] wl[29] vdd gnd cell_6t
Xbit_r30_c91 bl[91] br[91] wl[30] vdd gnd cell_6t
Xbit_r31_c91 bl[91] br[91] wl[31] vdd gnd cell_6t
Xbit_r32_c91 bl[91] br[91] wl[32] vdd gnd cell_6t
Xbit_r33_c91 bl[91] br[91] wl[33] vdd gnd cell_6t
Xbit_r34_c91 bl[91] br[91] wl[34] vdd gnd cell_6t
Xbit_r35_c91 bl[91] br[91] wl[35] vdd gnd cell_6t
Xbit_r36_c91 bl[91] br[91] wl[36] vdd gnd cell_6t
Xbit_r37_c91 bl[91] br[91] wl[37] vdd gnd cell_6t
Xbit_r38_c91 bl[91] br[91] wl[38] vdd gnd cell_6t
Xbit_r39_c91 bl[91] br[91] wl[39] vdd gnd cell_6t
Xbit_r40_c91 bl[91] br[91] wl[40] vdd gnd cell_6t
Xbit_r41_c91 bl[91] br[91] wl[41] vdd gnd cell_6t
Xbit_r42_c91 bl[91] br[91] wl[42] vdd gnd cell_6t
Xbit_r43_c91 bl[91] br[91] wl[43] vdd gnd cell_6t
Xbit_r44_c91 bl[91] br[91] wl[44] vdd gnd cell_6t
Xbit_r45_c91 bl[91] br[91] wl[45] vdd gnd cell_6t
Xbit_r46_c91 bl[91] br[91] wl[46] vdd gnd cell_6t
Xbit_r47_c91 bl[91] br[91] wl[47] vdd gnd cell_6t
Xbit_r48_c91 bl[91] br[91] wl[48] vdd gnd cell_6t
Xbit_r49_c91 bl[91] br[91] wl[49] vdd gnd cell_6t
Xbit_r50_c91 bl[91] br[91] wl[50] vdd gnd cell_6t
Xbit_r51_c91 bl[91] br[91] wl[51] vdd gnd cell_6t
Xbit_r52_c91 bl[91] br[91] wl[52] vdd gnd cell_6t
Xbit_r53_c91 bl[91] br[91] wl[53] vdd gnd cell_6t
Xbit_r54_c91 bl[91] br[91] wl[54] vdd gnd cell_6t
Xbit_r55_c91 bl[91] br[91] wl[55] vdd gnd cell_6t
Xbit_r56_c91 bl[91] br[91] wl[56] vdd gnd cell_6t
Xbit_r57_c91 bl[91] br[91] wl[57] vdd gnd cell_6t
Xbit_r58_c91 bl[91] br[91] wl[58] vdd gnd cell_6t
Xbit_r59_c91 bl[91] br[91] wl[59] vdd gnd cell_6t
Xbit_r60_c91 bl[91] br[91] wl[60] vdd gnd cell_6t
Xbit_r61_c91 bl[91] br[91] wl[61] vdd gnd cell_6t
Xbit_r62_c91 bl[91] br[91] wl[62] vdd gnd cell_6t
Xbit_r63_c91 bl[91] br[91] wl[63] vdd gnd cell_6t
Xbit_r64_c91 bl[91] br[91] wl[64] vdd gnd cell_6t
Xbit_r65_c91 bl[91] br[91] wl[65] vdd gnd cell_6t
Xbit_r66_c91 bl[91] br[91] wl[66] vdd gnd cell_6t
Xbit_r67_c91 bl[91] br[91] wl[67] vdd gnd cell_6t
Xbit_r68_c91 bl[91] br[91] wl[68] vdd gnd cell_6t
Xbit_r69_c91 bl[91] br[91] wl[69] vdd gnd cell_6t
Xbit_r70_c91 bl[91] br[91] wl[70] vdd gnd cell_6t
Xbit_r71_c91 bl[91] br[91] wl[71] vdd gnd cell_6t
Xbit_r72_c91 bl[91] br[91] wl[72] vdd gnd cell_6t
Xbit_r73_c91 bl[91] br[91] wl[73] vdd gnd cell_6t
Xbit_r74_c91 bl[91] br[91] wl[74] vdd gnd cell_6t
Xbit_r75_c91 bl[91] br[91] wl[75] vdd gnd cell_6t
Xbit_r76_c91 bl[91] br[91] wl[76] vdd gnd cell_6t
Xbit_r77_c91 bl[91] br[91] wl[77] vdd gnd cell_6t
Xbit_r78_c91 bl[91] br[91] wl[78] vdd gnd cell_6t
Xbit_r79_c91 bl[91] br[91] wl[79] vdd gnd cell_6t
Xbit_r80_c91 bl[91] br[91] wl[80] vdd gnd cell_6t
Xbit_r81_c91 bl[91] br[91] wl[81] vdd gnd cell_6t
Xbit_r82_c91 bl[91] br[91] wl[82] vdd gnd cell_6t
Xbit_r83_c91 bl[91] br[91] wl[83] vdd gnd cell_6t
Xbit_r84_c91 bl[91] br[91] wl[84] vdd gnd cell_6t
Xbit_r85_c91 bl[91] br[91] wl[85] vdd gnd cell_6t
Xbit_r86_c91 bl[91] br[91] wl[86] vdd gnd cell_6t
Xbit_r87_c91 bl[91] br[91] wl[87] vdd gnd cell_6t
Xbit_r88_c91 bl[91] br[91] wl[88] vdd gnd cell_6t
Xbit_r89_c91 bl[91] br[91] wl[89] vdd gnd cell_6t
Xbit_r90_c91 bl[91] br[91] wl[90] vdd gnd cell_6t
Xbit_r91_c91 bl[91] br[91] wl[91] vdd gnd cell_6t
Xbit_r92_c91 bl[91] br[91] wl[92] vdd gnd cell_6t
Xbit_r93_c91 bl[91] br[91] wl[93] vdd gnd cell_6t
Xbit_r94_c91 bl[91] br[91] wl[94] vdd gnd cell_6t
Xbit_r95_c91 bl[91] br[91] wl[95] vdd gnd cell_6t
Xbit_r96_c91 bl[91] br[91] wl[96] vdd gnd cell_6t
Xbit_r97_c91 bl[91] br[91] wl[97] vdd gnd cell_6t
Xbit_r98_c91 bl[91] br[91] wl[98] vdd gnd cell_6t
Xbit_r99_c91 bl[91] br[91] wl[99] vdd gnd cell_6t
Xbit_r100_c91 bl[91] br[91] wl[100] vdd gnd cell_6t
Xbit_r101_c91 bl[91] br[91] wl[101] vdd gnd cell_6t
Xbit_r102_c91 bl[91] br[91] wl[102] vdd gnd cell_6t
Xbit_r103_c91 bl[91] br[91] wl[103] vdd gnd cell_6t
Xbit_r104_c91 bl[91] br[91] wl[104] vdd gnd cell_6t
Xbit_r105_c91 bl[91] br[91] wl[105] vdd gnd cell_6t
Xbit_r106_c91 bl[91] br[91] wl[106] vdd gnd cell_6t
Xbit_r107_c91 bl[91] br[91] wl[107] vdd gnd cell_6t
Xbit_r108_c91 bl[91] br[91] wl[108] vdd gnd cell_6t
Xbit_r109_c91 bl[91] br[91] wl[109] vdd gnd cell_6t
Xbit_r110_c91 bl[91] br[91] wl[110] vdd gnd cell_6t
Xbit_r111_c91 bl[91] br[91] wl[111] vdd gnd cell_6t
Xbit_r112_c91 bl[91] br[91] wl[112] vdd gnd cell_6t
Xbit_r113_c91 bl[91] br[91] wl[113] vdd gnd cell_6t
Xbit_r114_c91 bl[91] br[91] wl[114] vdd gnd cell_6t
Xbit_r115_c91 bl[91] br[91] wl[115] vdd gnd cell_6t
Xbit_r116_c91 bl[91] br[91] wl[116] vdd gnd cell_6t
Xbit_r117_c91 bl[91] br[91] wl[117] vdd gnd cell_6t
Xbit_r118_c91 bl[91] br[91] wl[118] vdd gnd cell_6t
Xbit_r119_c91 bl[91] br[91] wl[119] vdd gnd cell_6t
Xbit_r120_c91 bl[91] br[91] wl[120] vdd gnd cell_6t
Xbit_r121_c91 bl[91] br[91] wl[121] vdd gnd cell_6t
Xbit_r122_c91 bl[91] br[91] wl[122] vdd gnd cell_6t
Xbit_r123_c91 bl[91] br[91] wl[123] vdd gnd cell_6t
Xbit_r124_c91 bl[91] br[91] wl[124] vdd gnd cell_6t
Xbit_r125_c91 bl[91] br[91] wl[125] vdd gnd cell_6t
Xbit_r126_c91 bl[91] br[91] wl[126] vdd gnd cell_6t
Xbit_r127_c91 bl[91] br[91] wl[127] vdd gnd cell_6t
Xbit_r0_c92 bl[92] br[92] wl[0] vdd gnd cell_6t
Xbit_r1_c92 bl[92] br[92] wl[1] vdd gnd cell_6t
Xbit_r2_c92 bl[92] br[92] wl[2] vdd gnd cell_6t
Xbit_r3_c92 bl[92] br[92] wl[3] vdd gnd cell_6t
Xbit_r4_c92 bl[92] br[92] wl[4] vdd gnd cell_6t
Xbit_r5_c92 bl[92] br[92] wl[5] vdd gnd cell_6t
Xbit_r6_c92 bl[92] br[92] wl[6] vdd gnd cell_6t
Xbit_r7_c92 bl[92] br[92] wl[7] vdd gnd cell_6t
Xbit_r8_c92 bl[92] br[92] wl[8] vdd gnd cell_6t
Xbit_r9_c92 bl[92] br[92] wl[9] vdd gnd cell_6t
Xbit_r10_c92 bl[92] br[92] wl[10] vdd gnd cell_6t
Xbit_r11_c92 bl[92] br[92] wl[11] vdd gnd cell_6t
Xbit_r12_c92 bl[92] br[92] wl[12] vdd gnd cell_6t
Xbit_r13_c92 bl[92] br[92] wl[13] vdd gnd cell_6t
Xbit_r14_c92 bl[92] br[92] wl[14] vdd gnd cell_6t
Xbit_r15_c92 bl[92] br[92] wl[15] vdd gnd cell_6t
Xbit_r16_c92 bl[92] br[92] wl[16] vdd gnd cell_6t
Xbit_r17_c92 bl[92] br[92] wl[17] vdd gnd cell_6t
Xbit_r18_c92 bl[92] br[92] wl[18] vdd gnd cell_6t
Xbit_r19_c92 bl[92] br[92] wl[19] vdd gnd cell_6t
Xbit_r20_c92 bl[92] br[92] wl[20] vdd gnd cell_6t
Xbit_r21_c92 bl[92] br[92] wl[21] vdd gnd cell_6t
Xbit_r22_c92 bl[92] br[92] wl[22] vdd gnd cell_6t
Xbit_r23_c92 bl[92] br[92] wl[23] vdd gnd cell_6t
Xbit_r24_c92 bl[92] br[92] wl[24] vdd gnd cell_6t
Xbit_r25_c92 bl[92] br[92] wl[25] vdd gnd cell_6t
Xbit_r26_c92 bl[92] br[92] wl[26] vdd gnd cell_6t
Xbit_r27_c92 bl[92] br[92] wl[27] vdd gnd cell_6t
Xbit_r28_c92 bl[92] br[92] wl[28] vdd gnd cell_6t
Xbit_r29_c92 bl[92] br[92] wl[29] vdd gnd cell_6t
Xbit_r30_c92 bl[92] br[92] wl[30] vdd gnd cell_6t
Xbit_r31_c92 bl[92] br[92] wl[31] vdd gnd cell_6t
Xbit_r32_c92 bl[92] br[92] wl[32] vdd gnd cell_6t
Xbit_r33_c92 bl[92] br[92] wl[33] vdd gnd cell_6t
Xbit_r34_c92 bl[92] br[92] wl[34] vdd gnd cell_6t
Xbit_r35_c92 bl[92] br[92] wl[35] vdd gnd cell_6t
Xbit_r36_c92 bl[92] br[92] wl[36] vdd gnd cell_6t
Xbit_r37_c92 bl[92] br[92] wl[37] vdd gnd cell_6t
Xbit_r38_c92 bl[92] br[92] wl[38] vdd gnd cell_6t
Xbit_r39_c92 bl[92] br[92] wl[39] vdd gnd cell_6t
Xbit_r40_c92 bl[92] br[92] wl[40] vdd gnd cell_6t
Xbit_r41_c92 bl[92] br[92] wl[41] vdd gnd cell_6t
Xbit_r42_c92 bl[92] br[92] wl[42] vdd gnd cell_6t
Xbit_r43_c92 bl[92] br[92] wl[43] vdd gnd cell_6t
Xbit_r44_c92 bl[92] br[92] wl[44] vdd gnd cell_6t
Xbit_r45_c92 bl[92] br[92] wl[45] vdd gnd cell_6t
Xbit_r46_c92 bl[92] br[92] wl[46] vdd gnd cell_6t
Xbit_r47_c92 bl[92] br[92] wl[47] vdd gnd cell_6t
Xbit_r48_c92 bl[92] br[92] wl[48] vdd gnd cell_6t
Xbit_r49_c92 bl[92] br[92] wl[49] vdd gnd cell_6t
Xbit_r50_c92 bl[92] br[92] wl[50] vdd gnd cell_6t
Xbit_r51_c92 bl[92] br[92] wl[51] vdd gnd cell_6t
Xbit_r52_c92 bl[92] br[92] wl[52] vdd gnd cell_6t
Xbit_r53_c92 bl[92] br[92] wl[53] vdd gnd cell_6t
Xbit_r54_c92 bl[92] br[92] wl[54] vdd gnd cell_6t
Xbit_r55_c92 bl[92] br[92] wl[55] vdd gnd cell_6t
Xbit_r56_c92 bl[92] br[92] wl[56] vdd gnd cell_6t
Xbit_r57_c92 bl[92] br[92] wl[57] vdd gnd cell_6t
Xbit_r58_c92 bl[92] br[92] wl[58] vdd gnd cell_6t
Xbit_r59_c92 bl[92] br[92] wl[59] vdd gnd cell_6t
Xbit_r60_c92 bl[92] br[92] wl[60] vdd gnd cell_6t
Xbit_r61_c92 bl[92] br[92] wl[61] vdd gnd cell_6t
Xbit_r62_c92 bl[92] br[92] wl[62] vdd gnd cell_6t
Xbit_r63_c92 bl[92] br[92] wl[63] vdd gnd cell_6t
Xbit_r64_c92 bl[92] br[92] wl[64] vdd gnd cell_6t
Xbit_r65_c92 bl[92] br[92] wl[65] vdd gnd cell_6t
Xbit_r66_c92 bl[92] br[92] wl[66] vdd gnd cell_6t
Xbit_r67_c92 bl[92] br[92] wl[67] vdd gnd cell_6t
Xbit_r68_c92 bl[92] br[92] wl[68] vdd gnd cell_6t
Xbit_r69_c92 bl[92] br[92] wl[69] vdd gnd cell_6t
Xbit_r70_c92 bl[92] br[92] wl[70] vdd gnd cell_6t
Xbit_r71_c92 bl[92] br[92] wl[71] vdd gnd cell_6t
Xbit_r72_c92 bl[92] br[92] wl[72] vdd gnd cell_6t
Xbit_r73_c92 bl[92] br[92] wl[73] vdd gnd cell_6t
Xbit_r74_c92 bl[92] br[92] wl[74] vdd gnd cell_6t
Xbit_r75_c92 bl[92] br[92] wl[75] vdd gnd cell_6t
Xbit_r76_c92 bl[92] br[92] wl[76] vdd gnd cell_6t
Xbit_r77_c92 bl[92] br[92] wl[77] vdd gnd cell_6t
Xbit_r78_c92 bl[92] br[92] wl[78] vdd gnd cell_6t
Xbit_r79_c92 bl[92] br[92] wl[79] vdd gnd cell_6t
Xbit_r80_c92 bl[92] br[92] wl[80] vdd gnd cell_6t
Xbit_r81_c92 bl[92] br[92] wl[81] vdd gnd cell_6t
Xbit_r82_c92 bl[92] br[92] wl[82] vdd gnd cell_6t
Xbit_r83_c92 bl[92] br[92] wl[83] vdd gnd cell_6t
Xbit_r84_c92 bl[92] br[92] wl[84] vdd gnd cell_6t
Xbit_r85_c92 bl[92] br[92] wl[85] vdd gnd cell_6t
Xbit_r86_c92 bl[92] br[92] wl[86] vdd gnd cell_6t
Xbit_r87_c92 bl[92] br[92] wl[87] vdd gnd cell_6t
Xbit_r88_c92 bl[92] br[92] wl[88] vdd gnd cell_6t
Xbit_r89_c92 bl[92] br[92] wl[89] vdd gnd cell_6t
Xbit_r90_c92 bl[92] br[92] wl[90] vdd gnd cell_6t
Xbit_r91_c92 bl[92] br[92] wl[91] vdd gnd cell_6t
Xbit_r92_c92 bl[92] br[92] wl[92] vdd gnd cell_6t
Xbit_r93_c92 bl[92] br[92] wl[93] vdd gnd cell_6t
Xbit_r94_c92 bl[92] br[92] wl[94] vdd gnd cell_6t
Xbit_r95_c92 bl[92] br[92] wl[95] vdd gnd cell_6t
Xbit_r96_c92 bl[92] br[92] wl[96] vdd gnd cell_6t
Xbit_r97_c92 bl[92] br[92] wl[97] vdd gnd cell_6t
Xbit_r98_c92 bl[92] br[92] wl[98] vdd gnd cell_6t
Xbit_r99_c92 bl[92] br[92] wl[99] vdd gnd cell_6t
Xbit_r100_c92 bl[92] br[92] wl[100] vdd gnd cell_6t
Xbit_r101_c92 bl[92] br[92] wl[101] vdd gnd cell_6t
Xbit_r102_c92 bl[92] br[92] wl[102] vdd gnd cell_6t
Xbit_r103_c92 bl[92] br[92] wl[103] vdd gnd cell_6t
Xbit_r104_c92 bl[92] br[92] wl[104] vdd gnd cell_6t
Xbit_r105_c92 bl[92] br[92] wl[105] vdd gnd cell_6t
Xbit_r106_c92 bl[92] br[92] wl[106] vdd gnd cell_6t
Xbit_r107_c92 bl[92] br[92] wl[107] vdd gnd cell_6t
Xbit_r108_c92 bl[92] br[92] wl[108] vdd gnd cell_6t
Xbit_r109_c92 bl[92] br[92] wl[109] vdd gnd cell_6t
Xbit_r110_c92 bl[92] br[92] wl[110] vdd gnd cell_6t
Xbit_r111_c92 bl[92] br[92] wl[111] vdd gnd cell_6t
Xbit_r112_c92 bl[92] br[92] wl[112] vdd gnd cell_6t
Xbit_r113_c92 bl[92] br[92] wl[113] vdd gnd cell_6t
Xbit_r114_c92 bl[92] br[92] wl[114] vdd gnd cell_6t
Xbit_r115_c92 bl[92] br[92] wl[115] vdd gnd cell_6t
Xbit_r116_c92 bl[92] br[92] wl[116] vdd gnd cell_6t
Xbit_r117_c92 bl[92] br[92] wl[117] vdd gnd cell_6t
Xbit_r118_c92 bl[92] br[92] wl[118] vdd gnd cell_6t
Xbit_r119_c92 bl[92] br[92] wl[119] vdd gnd cell_6t
Xbit_r120_c92 bl[92] br[92] wl[120] vdd gnd cell_6t
Xbit_r121_c92 bl[92] br[92] wl[121] vdd gnd cell_6t
Xbit_r122_c92 bl[92] br[92] wl[122] vdd gnd cell_6t
Xbit_r123_c92 bl[92] br[92] wl[123] vdd gnd cell_6t
Xbit_r124_c92 bl[92] br[92] wl[124] vdd gnd cell_6t
Xbit_r125_c92 bl[92] br[92] wl[125] vdd gnd cell_6t
Xbit_r126_c92 bl[92] br[92] wl[126] vdd gnd cell_6t
Xbit_r127_c92 bl[92] br[92] wl[127] vdd gnd cell_6t
Xbit_r0_c93 bl[93] br[93] wl[0] vdd gnd cell_6t
Xbit_r1_c93 bl[93] br[93] wl[1] vdd gnd cell_6t
Xbit_r2_c93 bl[93] br[93] wl[2] vdd gnd cell_6t
Xbit_r3_c93 bl[93] br[93] wl[3] vdd gnd cell_6t
Xbit_r4_c93 bl[93] br[93] wl[4] vdd gnd cell_6t
Xbit_r5_c93 bl[93] br[93] wl[5] vdd gnd cell_6t
Xbit_r6_c93 bl[93] br[93] wl[6] vdd gnd cell_6t
Xbit_r7_c93 bl[93] br[93] wl[7] vdd gnd cell_6t
Xbit_r8_c93 bl[93] br[93] wl[8] vdd gnd cell_6t
Xbit_r9_c93 bl[93] br[93] wl[9] vdd gnd cell_6t
Xbit_r10_c93 bl[93] br[93] wl[10] vdd gnd cell_6t
Xbit_r11_c93 bl[93] br[93] wl[11] vdd gnd cell_6t
Xbit_r12_c93 bl[93] br[93] wl[12] vdd gnd cell_6t
Xbit_r13_c93 bl[93] br[93] wl[13] vdd gnd cell_6t
Xbit_r14_c93 bl[93] br[93] wl[14] vdd gnd cell_6t
Xbit_r15_c93 bl[93] br[93] wl[15] vdd gnd cell_6t
Xbit_r16_c93 bl[93] br[93] wl[16] vdd gnd cell_6t
Xbit_r17_c93 bl[93] br[93] wl[17] vdd gnd cell_6t
Xbit_r18_c93 bl[93] br[93] wl[18] vdd gnd cell_6t
Xbit_r19_c93 bl[93] br[93] wl[19] vdd gnd cell_6t
Xbit_r20_c93 bl[93] br[93] wl[20] vdd gnd cell_6t
Xbit_r21_c93 bl[93] br[93] wl[21] vdd gnd cell_6t
Xbit_r22_c93 bl[93] br[93] wl[22] vdd gnd cell_6t
Xbit_r23_c93 bl[93] br[93] wl[23] vdd gnd cell_6t
Xbit_r24_c93 bl[93] br[93] wl[24] vdd gnd cell_6t
Xbit_r25_c93 bl[93] br[93] wl[25] vdd gnd cell_6t
Xbit_r26_c93 bl[93] br[93] wl[26] vdd gnd cell_6t
Xbit_r27_c93 bl[93] br[93] wl[27] vdd gnd cell_6t
Xbit_r28_c93 bl[93] br[93] wl[28] vdd gnd cell_6t
Xbit_r29_c93 bl[93] br[93] wl[29] vdd gnd cell_6t
Xbit_r30_c93 bl[93] br[93] wl[30] vdd gnd cell_6t
Xbit_r31_c93 bl[93] br[93] wl[31] vdd gnd cell_6t
Xbit_r32_c93 bl[93] br[93] wl[32] vdd gnd cell_6t
Xbit_r33_c93 bl[93] br[93] wl[33] vdd gnd cell_6t
Xbit_r34_c93 bl[93] br[93] wl[34] vdd gnd cell_6t
Xbit_r35_c93 bl[93] br[93] wl[35] vdd gnd cell_6t
Xbit_r36_c93 bl[93] br[93] wl[36] vdd gnd cell_6t
Xbit_r37_c93 bl[93] br[93] wl[37] vdd gnd cell_6t
Xbit_r38_c93 bl[93] br[93] wl[38] vdd gnd cell_6t
Xbit_r39_c93 bl[93] br[93] wl[39] vdd gnd cell_6t
Xbit_r40_c93 bl[93] br[93] wl[40] vdd gnd cell_6t
Xbit_r41_c93 bl[93] br[93] wl[41] vdd gnd cell_6t
Xbit_r42_c93 bl[93] br[93] wl[42] vdd gnd cell_6t
Xbit_r43_c93 bl[93] br[93] wl[43] vdd gnd cell_6t
Xbit_r44_c93 bl[93] br[93] wl[44] vdd gnd cell_6t
Xbit_r45_c93 bl[93] br[93] wl[45] vdd gnd cell_6t
Xbit_r46_c93 bl[93] br[93] wl[46] vdd gnd cell_6t
Xbit_r47_c93 bl[93] br[93] wl[47] vdd gnd cell_6t
Xbit_r48_c93 bl[93] br[93] wl[48] vdd gnd cell_6t
Xbit_r49_c93 bl[93] br[93] wl[49] vdd gnd cell_6t
Xbit_r50_c93 bl[93] br[93] wl[50] vdd gnd cell_6t
Xbit_r51_c93 bl[93] br[93] wl[51] vdd gnd cell_6t
Xbit_r52_c93 bl[93] br[93] wl[52] vdd gnd cell_6t
Xbit_r53_c93 bl[93] br[93] wl[53] vdd gnd cell_6t
Xbit_r54_c93 bl[93] br[93] wl[54] vdd gnd cell_6t
Xbit_r55_c93 bl[93] br[93] wl[55] vdd gnd cell_6t
Xbit_r56_c93 bl[93] br[93] wl[56] vdd gnd cell_6t
Xbit_r57_c93 bl[93] br[93] wl[57] vdd gnd cell_6t
Xbit_r58_c93 bl[93] br[93] wl[58] vdd gnd cell_6t
Xbit_r59_c93 bl[93] br[93] wl[59] vdd gnd cell_6t
Xbit_r60_c93 bl[93] br[93] wl[60] vdd gnd cell_6t
Xbit_r61_c93 bl[93] br[93] wl[61] vdd gnd cell_6t
Xbit_r62_c93 bl[93] br[93] wl[62] vdd gnd cell_6t
Xbit_r63_c93 bl[93] br[93] wl[63] vdd gnd cell_6t
Xbit_r64_c93 bl[93] br[93] wl[64] vdd gnd cell_6t
Xbit_r65_c93 bl[93] br[93] wl[65] vdd gnd cell_6t
Xbit_r66_c93 bl[93] br[93] wl[66] vdd gnd cell_6t
Xbit_r67_c93 bl[93] br[93] wl[67] vdd gnd cell_6t
Xbit_r68_c93 bl[93] br[93] wl[68] vdd gnd cell_6t
Xbit_r69_c93 bl[93] br[93] wl[69] vdd gnd cell_6t
Xbit_r70_c93 bl[93] br[93] wl[70] vdd gnd cell_6t
Xbit_r71_c93 bl[93] br[93] wl[71] vdd gnd cell_6t
Xbit_r72_c93 bl[93] br[93] wl[72] vdd gnd cell_6t
Xbit_r73_c93 bl[93] br[93] wl[73] vdd gnd cell_6t
Xbit_r74_c93 bl[93] br[93] wl[74] vdd gnd cell_6t
Xbit_r75_c93 bl[93] br[93] wl[75] vdd gnd cell_6t
Xbit_r76_c93 bl[93] br[93] wl[76] vdd gnd cell_6t
Xbit_r77_c93 bl[93] br[93] wl[77] vdd gnd cell_6t
Xbit_r78_c93 bl[93] br[93] wl[78] vdd gnd cell_6t
Xbit_r79_c93 bl[93] br[93] wl[79] vdd gnd cell_6t
Xbit_r80_c93 bl[93] br[93] wl[80] vdd gnd cell_6t
Xbit_r81_c93 bl[93] br[93] wl[81] vdd gnd cell_6t
Xbit_r82_c93 bl[93] br[93] wl[82] vdd gnd cell_6t
Xbit_r83_c93 bl[93] br[93] wl[83] vdd gnd cell_6t
Xbit_r84_c93 bl[93] br[93] wl[84] vdd gnd cell_6t
Xbit_r85_c93 bl[93] br[93] wl[85] vdd gnd cell_6t
Xbit_r86_c93 bl[93] br[93] wl[86] vdd gnd cell_6t
Xbit_r87_c93 bl[93] br[93] wl[87] vdd gnd cell_6t
Xbit_r88_c93 bl[93] br[93] wl[88] vdd gnd cell_6t
Xbit_r89_c93 bl[93] br[93] wl[89] vdd gnd cell_6t
Xbit_r90_c93 bl[93] br[93] wl[90] vdd gnd cell_6t
Xbit_r91_c93 bl[93] br[93] wl[91] vdd gnd cell_6t
Xbit_r92_c93 bl[93] br[93] wl[92] vdd gnd cell_6t
Xbit_r93_c93 bl[93] br[93] wl[93] vdd gnd cell_6t
Xbit_r94_c93 bl[93] br[93] wl[94] vdd gnd cell_6t
Xbit_r95_c93 bl[93] br[93] wl[95] vdd gnd cell_6t
Xbit_r96_c93 bl[93] br[93] wl[96] vdd gnd cell_6t
Xbit_r97_c93 bl[93] br[93] wl[97] vdd gnd cell_6t
Xbit_r98_c93 bl[93] br[93] wl[98] vdd gnd cell_6t
Xbit_r99_c93 bl[93] br[93] wl[99] vdd gnd cell_6t
Xbit_r100_c93 bl[93] br[93] wl[100] vdd gnd cell_6t
Xbit_r101_c93 bl[93] br[93] wl[101] vdd gnd cell_6t
Xbit_r102_c93 bl[93] br[93] wl[102] vdd gnd cell_6t
Xbit_r103_c93 bl[93] br[93] wl[103] vdd gnd cell_6t
Xbit_r104_c93 bl[93] br[93] wl[104] vdd gnd cell_6t
Xbit_r105_c93 bl[93] br[93] wl[105] vdd gnd cell_6t
Xbit_r106_c93 bl[93] br[93] wl[106] vdd gnd cell_6t
Xbit_r107_c93 bl[93] br[93] wl[107] vdd gnd cell_6t
Xbit_r108_c93 bl[93] br[93] wl[108] vdd gnd cell_6t
Xbit_r109_c93 bl[93] br[93] wl[109] vdd gnd cell_6t
Xbit_r110_c93 bl[93] br[93] wl[110] vdd gnd cell_6t
Xbit_r111_c93 bl[93] br[93] wl[111] vdd gnd cell_6t
Xbit_r112_c93 bl[93] br[93] wl[112] vdd gnd cell_6t
Xbit_r113_c93 bl[93] br[93] wl[113] vdd gnd cell_6t
Xbit_r114_c93 bl[93] br[93] wl[114] vdd gnd cell_6t
Xbit_r115_c93 bl[93] br[93] wl[115] vdd gnd cell_6t
Xbit_r116_c93 bl[93] br[93] wl[116] vdd gnd cell_6t
Xbit_r117_c93 bl[93] br[93] wl[117] vdd gnd cell_6t
Xbit_r118_c93 bl[93] br[93] wl[118] vdd gnd cell_6t
Xbit_r119_c93 bl[93] br[93] wl[119] vdd gnd cell_6t
Xbit_r120_c93 bl[93] br[93] wl[120] vdd gnd cell_6t
Xbit_r121_c93 bl[93] br[93] wl[121] vdd gnd cell_6t
Xbit_r122_c93 bl[93] br[93] wl[122] vdd gnd cell_6t
Xbit_r123_c93 bl[93] br[93] wl[123] vdd gnd cell_6t
Xbit_r124_c93 bl[93] br[93] wl[124] vdd gnd cell_6t
Xbit_r125_c93 bl[93] br[93] wl[125] vdd gnd cell_6t
Xbit_r126_c93 bl[93] br[93] wl[126] vdd gnd cell_6t
Xbit_r127_c93 bl[93] br[93] wl[127] vdd gnd cell_6t
Xbit_r0_c94 bl[94] br[94] wl[0] vdd gnd cell_6t
Xbit_r1_c94 bl[94] br[94] wl[1] vdd gnd cell_6t
Xbit_r2_c94 bl[94] br[94] wl[2] vdd gnd cell_6t
Xbit_r3_c94 bl[94] br[94] wl[3] vdd gnd cell_6t
Xbit_r4_c94 bl[94] br[94] wl[4] vdd gnd cell_6t
Xbit_r5_c94 bl[94] br[94] wl[5] vdd gnd cell_6t
Xbit_r6_c94 bl[94] br[94] wl[6] vdd gnd cell_6t
Xbit_r7_c94 bl[94] br[94] wl[7] vdd gnd cell_6t
Xbit_r8_c94 bl[94] br[94] wl[8] vdd gnd cell_6t
Xbit_r9_c94 bl[94] br[94] wl[9] vdd gnd cell_6t
Xbit_r10_c94 bl[94] br[94] wl[10] vdd gnd cell_6t
Xbit_r11_c94 bl[94] br[94] wl[11] vdd gnd cell_6t
Xbit_r12_c94 bl[94] br[94] wl[12] vdd gnd cell_6t
Xbit_r13_c94 bl[94] br[94] wl[13] vdd gnd cell_6t
Xbit_r14_c94 bl[94] br[94] wl[14] vdd gnd cell_6t
Xbit_r15_c94 bl[94] br[94] wl[15] vdd gnd cell_6t
Xbit_r16_c94 bl[94] br[94] wl[16] vdd gnd cell_6t
Xbit_r17_c94 bl[94] br[94] wl[17] vdd gnd cell_6t
Xbit_r18_c94 bl[94] br[94] wl[18] vdd gnd cell_6t
Xbit_r19_c94 bl[94] br[94] wl[19] vdd gnd cell_6t
Xbit_r20_c94 bl[94] br[94] wl[20] vdd gnd cell_6t
Xbit_r21_c94 bl[94] br[94] wl[21] vdd gnd cell_6t
Xbit_r22_c94 bl[94] br[94] wl[22] vdd gnd cell_6t
Xbit_r23_c94 bl[94] br[94] wl[23] vdd gnd cell_6t
Xbit_r24_c94 bl[94] br[94] wl[24] vdd gnd cell_6t
Xbit_r25_c94 bl[94] br[94] wl[25] vdd gnd cell_6t
Xbit_r26_c94 bl[94] br[94] wl[26] vdd gnd cell_6t
Xbit_r27_c94 bl[94] br[94] wl[27] vdd gnd cell_6t
Xbit_r28_c94 bl[94] br[94] wl[28] vdd gnd cell_6t
Xbit_r29_c94 bl[94] br[94] wl[29] vdd gnd cell_6t
Xbit_r30_c94 bl[94] br[94] wl[30] vdd gnd cell_6t
Xbit_r31_c94 bl[94] br[94] wl[31] vdd gnd cell_6t
Xbit_r32_c94 bl[94] br[94] wl[32] vdd gnd cell_6t
Xbit_r33_c94 bl[94] br[94] wl[33] vdd gnd cell_6t
Xbit_r34_c94 bl[94] br[94] wl[34] vdd gnd cell_6t
Xbit_r35_c94 bl[94] br[94] wl[35] vdd gnd cell_6t
Xbit_r36_c94 bl[94] br[94] wl[36] vdd gnd cell_6t
Xbit_r37_c94 bl[94] br[94] wl[37] vdd gnd cell_6t
Xbit_r38_c94 bl[94] br[94] wl[38] vdd gnd cell_6t
Xbit_r39_c94 bl[94] br[94] wl[39] vdd gnd cell_6t
Xbit_r40_c94 bl[94] br[94] wl[40] vdd gnd cell_6t
Xbit_r41_c94 bl[94] br[94] wl[41] vdd gnd cell_6t
Xbit_r42_c94 bl[94] br[94] wl[42] vdd gnd cell_6t
Xbit_r43_c94 bl[94] br[94] wl[43] vdd gnd cell_6t
Xbit_r44_c94 bl[94] br[94] wl[44] vdd gnd cell_6t
Xbit_r45_c94 bl[94] br[94] wl[45] vdd gnd cell_6t
Xbit_r46_c94 bl[94] br[94] wl[46] vdd gnd cell_6t
Xbit_r47_c94 bl[94] br[94] wl[47] vdd gnd cell_6t
Xbit_r48_c94 bl[94] br[94] wl[48] vdd gnd cell_6t
Xbit_r49_c94 bl[94] br[94] wl[49] vdd gnd cell_6t
Xbit_r50_c94 bl[94] br[94] wl[50] vdd gnd cell_6t
Xbit_r51_c94 bl[94] br[94] wl[51] vdd gnd cell_6t
Xbit_r52_c94 bl[94] br[94] wl[52] vdd gnd cell_6t
Xbit_r53_c94 bl[94] br[94] wl[53] vdd gnd cell_6t
Xbit_r54_c94 bl[94] br[94] wl[54] vdd gnd cell_6t
Xbit_r55_c94 bl[94] br[94] wl[55] vdd gnd cell_6t
Xbit_r56_c94 bl[94] br[94] wl[56] vdd gnd cell_6t
Xbit_r57_c94 bl[94] br[94] wl[57] vdd gnd cell_6t
Xbit_r58_c94 bl[94] br[94] wl[58] vdd gnd cell_6t
Xbit_r59_c94 bl[94] br[94] wl[59] vdd gnd cell_6t
Xbit_r60_c94 bl[94] br[94] wl[60] vdd gnd cell_6t
Xbit_r61_c94 bl[94] br[94] wl[61] vdd gnd cell_6t
Xbit_r62_c94 bl[94] br[94] wl[62] vdd gnd cell_6t
Xbit_r63_c94 bl[94] br[94] wl[63] vdd gnd cell_6t
Xbit_r64_c94 bl[94] br[94] wl[64] vdd gnd cell_6t
Xbit_r65_c94 bl[94] br[94] wl[65] vdd gnd cell_6t
Xbit_r66_c94 bl[94] br[94] wl[66] vdd gnd cell_6t
Xbit_r67_c94 bl[94] br[94] wl[67] vdd gnd cell_6t
Xbit_r68_c94 bl[94] br[94] wl[68] vdd gnd cell_6t
Xbit_r69_c94 bl[94] br[94] wl[69] vdd gnd cell_6t
Xbit_r70_c94 bl[94] br[94] wl[70] vdd gnd cell_6t
Xbit_r71_c94 bl[94] br[94] wl[71] vdd gnd cell_6t
Xbit_r72_c94 bl[94] br[94] wl[72] vdd gnd cell_6t
Xbit_r73_c94 bl[94] br[94] wl[73] vdd gnd cell_6t
Xbit_r74_c94 bl[94] br[94] wl[74] vdd gnd cell_6t
Xbit_r75_c94 bl[94] br[94] wl[75] vdd gnd cell_6t
Xbit_r76_c94 bl[94] br[94] wl[76] vdd gnd cell_6t
Xbit_r77_c94 bl[94] br[94] wl[77] vdd gnd cell_6t
Xbit_r78_c94 bl[94] br[94] wl[78] vdd gnd cell_6t
Xbit_r79_c94 bl[94] br[94] wl[79] vdd gnd cell_6t
Xbit_r80_c94 bl[94] br[94] wl[80] vdd gnd cell_6t
Xbit_r81_c94 bl[94] br[94] wl[81] vdd gnd cell_6t
Xbit_r82_c94 bl[94] br[94] wl[82] vdd gnd cell_6t
Xbit_r83_c94 bl[94] br[94] wl[83] vdd gnd cell_6t
Xbit_r84_c94 bl[94] br[94] wl[84] vdd gnd cell_6t
Xbit_r85_c94 bl[94] br[94] wl[85] vdd gnd cell_6t
Xbit_r86_c94 bl[94] br[94] wl[86] vdd gnd cell_6t
Xbit_r87_c94 bl[94] br[94] wl[87] vdd gnd cell_6t
Xbit_r88_c94 bl[94] br[94] wl[88] vdd gnd cell_6t
Xbit_r89_c94 bl[94] br[94] wl[89] vdd gnd cell_6t
Xbit_r90_c94 bl[94] br[94] wl[90] vdd gnd cell_6t
Xbit_r91_c94 bl[94] br[94] wl[91] vdd gnd cell_6t
Xbit_r92_c94 bl[94] br[94] wl[92] vdd gnd cell_6t
Xbit_r93_c94 bl[94] br[94] wl[93] vdd gnd cell_6t
Xbit_r94_c94 bl[94] br[94] wl[94] vdd gnd cell_6t
Xbit_r95_c94 bl[94] br[94] wl[95] vdd gnd cell_6t
Xbit_r96_c94 bl[94] br[94] wl[96] vdd gnd cell_6t
Xbit_r97_c94 bl[94] br[94] wl[97] vdd gnd cell_6t
Xbit_r98_c94 bl[94] br[94] wl[98] vdd gnd cell_6t
Xbit_r99_c94 bl[94] br[94] wl[99] vdd gnd cell_6t
Xbit_r100_c94 bl[94] br[94] wl[100] vdd gnd cell_6t
Xbit_r101_c94 bl[94] br[94] wl[101] vdd gnd cell_6t
Xbit_r102_c94 bl[94] br[94] wl[102] vdd gnd cell_6t
Xbit_r103_c94 bl[94] br[94] wl[103] vdd gnd cell_6t
Xbit_r104_c94 bl[94] br[94] wl[104] vdd gnd cell_6t
Xbit_r105_c94 bl[94] br[94] wl[105] vdd gnd cell_6t
Xbit_r106_c94 bl[94] br[94] wl[106] vdd gnd cell_6t
Xbit_r107_c94 bl[94] br[94] wl[107] vdd gnd cell_6t
Xbit_r108_c94 bl[94] br[94] wl[108] vdd gnd cell_6t
Xbit_r109_c94 bl[94] br[94] wl[109] vdd gnd cell_6t
Xbit_r110_c94 bl[94] br[94] wl[110] vdd gnd cell_6t
Xbit_r111_c94 bl[94] br[94] wl[111] vdd gnd cell_6t
Xbit_r112_c94 bl[94] br[94] wl[112] vdd gnd cell_6t
Xbit_r113_c94 bl[94] br[94] wl[113] vdd gnd cell_6t
Xbit_r114_c94 bl[94] br[94] wl[114] vdd gnd cell_6t
Xbit_r115_c94 bl[94] br[94] wl[115] vdd gnd cell_6t
Xbit_r116_c94 bl[94] br[94] wl[116] vdd gnd cell_6t
Xbit_r117_c94 bl[94] br[94] wl[117] vdd gnd cell_6t
Xbit_r118_c94 bl[94] br[94] wl[118] vdd gnd cell_6t
Xbit_r119_c94 bl[94] br[94] wl[119] vdd gnd cell_6t
Xbit_r120_c94 bl[94] br[94] wl[120] vdd gnd cell_6t
Xbit_r121_c94 bl[94] br[94] wl[121] vdd gnd cell_6t
Xbit_r122_c94 bl[94] br[94] wl[122] vdd gnd cell_6t
Xbit_r123_c94 bl[94] br[94] wl[123] vdd gnd cell_6t
Xbit_r124_c94 bl[94] br[94] wl[124] vdd gnd cell_6t
Xbit_r125_c94 bl[94] br[94] wl[125] vdd gnd cell_6t
Xbit_r126_c94 bl[94] br[94] wl[126] vdd gnd cell_6t
Xbit_r127_c94 bl[94] br[94] wl[127] vdd gnd cell_6t
Xbit_r0_c95 bl[95] br[95] wl[0] vdd gnd cell_6t
Xbit_r1_c95 bl[95] br[95] wl[1] vdd gnd cell_6t
Xbit_r2_c95 bl[95] br[95] wl[2] vdd gnd cell_6t
Xbit_r3_c95 bl[95] br[95] wl[3] vdd gnd cell_6t
Xbit_r4_c95 bl[95] br[95] wl[4] vdd gnd cell_6t
Xbit_r5_c95 bl[95] br[95] wl[5] vdd gnd cell_6t
Xbit_r6_c95 bl[95] br[95] wl[6] vdd gnd cell_6t
Xbit_r7_c95 bl[95] br[95] wl[7] vdd gnd cell_6t
Xbit_r8_c95 bl[95] br[95] wl[8] vdd gnd cell_6t
Xbit_r9_c95 bl[95] br[95] wl[9] vdd gnd cell_6t
Xbit_r10_c95 bl[95] br[95] wl[10] vdd gnd cell_6t
Xbit_r11_c95 bl[95] br[95] wl[11] vdd gnd cell_6t
Xbit_r12_c95 bl[95] br[95] wl[12] vdd gnd cell_6t
Xbit_r13_c95 bl[95] br[95] wl[13] vdd gnd cell_6t
Xbit_r14_c95 bl[95] br[95] wl[14] vdd gnd cell_6t
Xbit_r15_c95 bl[95] br[95] wl[15] vdd gnd cell_6t
Xbit_r16_c95 bl[95] br[95] wl[16] vdd gnd cell_6t
Xbit_r17_c95 bl[95] br[95] wl[17] vdd gnd cell_6t
Xbit_r18_c95 bl[95] br[95] wl[18] vdd gnd cell_6t
Xbit_r19_c95 bl[95] br[95] wl[19] vdd gnd cell_6t
Xbit_r20_c95 bl[95] br[95] wl[20] vdd gnd cell_6t
Xbit_r21_c95 bl[95] br[95] wl[21] vdd gnd cell_6t
Xbit_r22_c95 bl[95] br[95] wl[22] vdd gnd cell_6t
Xbit_r23_c95 bl[95] br[95] wl[23] vdd gnd cell_6t
Xbit_r24_c95 bl[95] br[95] wl[24] vdd gnd cell_6t
Xbit_r25_c95 bl[95] br[95] wl[25] vdd gnd cell_6t
Xbit_r26_c95 bl[95] br[95] wl[26] vdd gnd cell_6t
Xbit_r27_c95 bl[95] br[95] wl[27] vdd gnd cell_6t
Xbit_r28_c95 bl[95] br[95] wl[28] vdd gnd cell_6t
Xbit_r29_c95 bl[95] br[95] wl[29] vdd gnd cell_6t
Xbit_r30_c95 bl[95] br[95] wl[30] vdd gnd cell_6t
Xbit_r31_c95 bl[95] br[95] wl[31] vdd gnd cell_6t
Xbit_r32_c95 bl[95] br[95] wl[32] vdd gnd cell_6t
Xbit_r33_c95 bl[95] br[95] wl[33] vdd gnd cell_6t
Xbit_r34_c95 bl[95] br[95] wl[34] vdd gnd cell_6t
Xbit_r35_c95 bl[95] br[95] wl[35] vdd gnd cell_6t
Xbit_r36_c95 bl[95] br[95] wl[36] vdd gnd cell_6t
Xbit_r37_c95 bl[95] br[95] wl[37] vdd gnd cell_6t
Xbit_r38_c95 bl[95] br[95] wl[38] vdd gnd cell_6t
Xbit_r39_c95 bl[95] br[95] wl[39] vdd gnd cell_6t
Xbit_r40_c95 bl[95] br[95] wl[40] vdd gnd cell_6t
Xbit_r41_c95 bl[95] br[95] wl[41] vdd gnd cell_6t
Xbit_r42_c95 bl[95] br[95] wl[42] vdd gnd cell_6t
Xbit_r43_c95 bl[95] br[95] wl[43] vdd gnd cell_6t
Xbit_r44_c95 bl[95] br[95] wl[44] vdd gnd cell_6t
Xbit_r45_c95 bl[95] br[95] wl[45] vdd gnd cell_6t
Xbit_r46_c95 bl[95] br[95] wl[46] vdd gnd cell_6t
Xbit_r47_c95 bl[95] br[95] wl[47] vdd gnd cell_6t
Xbit_r48_c95 bl[95] br[95] wl[48] vdd gnd cell_6t
Xbit_r49_c95 bl[95] br[95] wl[49] vdd gnd cell_6t
Xbit_r50_c95 bl[95] br[95] wl[50] vdd gnd cell_6t
Xbit_r51_c95 bl[95] br[95] wl[51] vdd gnd cell_6t
Xbit_r52_c95 bl[95] br[95] wl[52] vdd gnd cell_6t
Xbit_r53_c95 bl[95] br[95] wl[53] vdd gnd cell_6t
Xbit_r54_c95 bl[95] br[95] wl[54] vdd gnd cell_6t
Xbit_r55_c95 bl[95] br[95] wl[55] vdd gnd cell_6t
Xbit_r56_c95 bl[95] br[95] wl[56] vdd gnd cell_6t
Xbit_r57_c95 bl[95] br[95] wl[57] vdd gnd cell_6t
Xbit_r58_c95 bl[95] br[95] wl[58] vdd gnd cell_6t
Xbit_r59_c95 bl[95] br[95] wl[59] vdd gnd cell_6t
Xbit_r60_c95 bl[95] br[95] wl[60] vdd gnd cell_6t
Xbit_r61_c95 bl[95] br[95] wl[61] vdd gnd cell_6t
Xbit_r62_c95 bl[95] br[95] wl[62] vdd gnd cell_6t
Xbit_r63_c95 bl[95] br[95] wl[63] vdd gnd cell_6t
Xbit_r64_c95 bl[95] br[95] wl[64] vdd gnd cell_6t
Xbit_r65_c95 bl[95] br[95] wl[65] vdd gnd cell_6t
Xbit_r66_c95 bl[95] br[95] wl[66] vdd gnd cell_6t
Xbit_r67_c95 bl[95] br[95] wl[67] vdd gnd cell_6t
Xbit_r68_c95 bl[95] br[95] wl[68] vdd gnd cell_6t
Xbit_r69_c95 bl[95] br[95] wl[69] vdd gnd cell_6t
Xbit_r70_c95 bl[95] br[95] wl[70] vdd gnd cell_6t
Xbit_r71_c95 bl[95] br[95] wl[71] vdd gnd cell_6t
Xbit_r72_c95 bl[95] br[95] wl[72] vdd gnd cell_6t
Xbit_r73_c95 bl[95] br[95] wl[73] vdd gnd cell_6t
Xbit_r74_c95 bl[95] br[95] wl[74] vdd gnd cell_6t
Xbit_r75_c95 bl[95] br[95] wl[75] vdd gnd cell_6t
Xbit_r76_c95 bl[95] br[95] wl[76] vdd gnd cell_6t
Xbit_r77_c95 bl[95] br[95] wl[77] vdd gnd cell_6t
Xbit_r78_c95 bl[95] br[95] wl[78] vdd gnd cell_6t
Xbit_r79_c95 bl[95] br[95] wl[79] vdd gnd cell_6t
Xbit_r80_c95 bl[95] br[95] wl[80] vdd gnd cell_6t
Xbit_r81_c95 bl[95] br[95] wl[81] vdd gnd cell_6t
Xbit_r82_c95 bl[95] br[95] wl[82] vdd gnd cell_6t
Xbit_r83_c95 bl[95] br[95] wl[83] vdd gnd cell_6t
Xbit_r84_c95 bl[95] br[95] wl[84] vdd gnd cell_6t
Xbit_r85_c95 bl[95] br[95] wl[85] vdd gnd cell_6t
Xbit_r86_c95 bl[95] br[95] wl[86] vdd gnd cell_6t
Xbit_r87_c95 bl[95] br[95] wl[87] vdd gnd cell_6t
Xbit_r88_c95 bl[95] br[95] wl[88] vdd gnd cell_6t
Xbit_r89_c95 bl[95] br[95] wl[89] vdd gnd cell_6t
Xbit_r90_c95 bl[95] br[95] wl[90] vdd gnd cell_6t
Xbit_r91_c95 bl[95] br[95] wl[91] vdd gnd cell_6t
Xbit_r92_c95 bl[95] br[95] wl[92] vdd gnd cell_6t
Xbit_r93_c95 bl[95] br[95] wl[93] vdd gnd cell_6t
Xbit_r94_c95 bl[95] br[95] wl[94] vdd gnd cell_6t
Xbit_r95_c95 bl[95] br[95] wl[95] vdd gnd cell_6t
Xbit_r96_c95 bl[95] br[95] wl[96] vdd gnd cell_6t
Xbit_r97_c95 bl[95] br[95] wl[97] vdd gnd cell_6t
Xbit_r98_c95 bl[95] br[95] wl[98] vdd gnd cell_6t
Xbit_r99_c95 bl[95] br[95] wl[99] vdd gnd cell_6t
Xbit_r100_c95 bl[95] br[95] wl[100] vdd gnd cell_6t
Xbit_r101_c95 bl[95] br[95] wl[101] vdd gnd cell_6t
Xbit_r102_c95 bl[95] br[95] wl[102] vdd gnd cell_6t
Xbit_r103_c95 bl[95] br[95] wl[103] vdd gnd cell_6t
Xbit_r104_c95 bl[95] br[95] wl[104] vdd gnd cell_6t
Xbit_r105_c95 bl[95] br[95] wl[105] vdd gnd cell_6t
Xbit_r106_c95 bl[95] br[95] wl[106] vdd gnd cell_6t
Xbit_r107_c95 bl[95] br[95] wl[107] vdd gnd cell_6t
Xbit_r108_c95 bl[95] br[95] wl[108] vdd gnd cell_6t
Xbit_r109_c95 bl[95] br[95] wl[109] vdd gnd cell_6t
Xbit_r110_c95 bl[95] br[95] wl[110] vdd gnd cell_6t
Xbit_r111_c95 bl[95] br[95] wl[111] vdd gnd cell_6t
Xbit_r112_c95 bl[95] br[95] wl[112] vdd gnd cell_6t
Xbit_r113_c95 bl[95] br[95] wl[113] vdd gnd cell_6t
Xbit_r114_c95 bl[95] br[95] wl[114] vdd gnd cell_6t
Xbit_r115_c95 bl[95] br[95] wl[115] vdd gnd cell_6t
Xbit_r116_c95 bl[95] br[95] wl[116] vdd gnd cell_6t
Xbit_r117_c95 bl[95] br[95] wl[117] vdd gnd cell_6t
Xbit_r118_c95 bl[95] br[95] wl[118] vdd gnd cell_6t
Xbit_r119_c95 bl[95] br[95] wl[119] vdd gnd cell_6t
Xbit_r120_c95 bl[95] br[95] wl[120] vdd gnd cell_6t
Xbit_r121_c95 bl[95] br[95] wl[121] vdd gnd cell_6t
Xbit_r122_c95 bl[95] br[95] wl[122] vdd gnd cell_6t
Xbit_r123_c95 bl[95] br[95] wl[123] vdd gnd cell_6t
Xbit_r124_c95 bl[95] br[95] wl[124] vdd gnd cell_6t
Xbit_r125_c95 bl[95] br[95] wl[125] vdd gnd cell_6t
Xbit_r126_c95 bl[95] br[95] wl[126] vdd gnd cell_6t
Xbit_r127_c95 bl[95] br[95] wl[127] vdd gnd cell_6t
Xbit_r0_c96 bl[96] br[96] wl[0] vdd gnd cell_6t
Xbit_r1_c96 bl[96] br[96] wl[1] vdd gnd cell_6t
Xbit_r2_c96 bl[96] br[96] wl[2] vdd gnd cell_6t
Xbit_r3_c96 bl[96] br[96] wl[3] vdd gnd cell_6t
Xbit_r4_c96 bl[96] br[96] wl[4] vdd gnd cell_6t
Xbit_r5_c96 bl[96] br[96] wl[5] vdd gnd cell_6t
Xbit_r6_c96 bl[96] br[96] wl[6] vdd gnd cell_6t
Xbit_r7_c96 bl[96] br[96] wl[7] vdd gnd cell_6t
Xbit_r8_c96 bl[96] br[96] wl[8] vdd gnd cell_6t
Xbit_r9_c96 bl[96] br[96] wl[9] vdd gnd cell_6t
Xbit_r10_c96 bl[96] br[96] wl[10] vdd gnd cell_6t
Xbit_r11_c96 bl[96] br[96] wl[11] vdd gnd cell_6t
Xbit_r12_c96 bl[96] br[96] wl[12] vdd gnd cell_6t
Xbit_r13_c96 bl[96] br[96] wl[13] vdd gnd cell_6t
Xbit_r14_c96 bl[96] br[96] wl[14] vdd gnd cell_6t
Xbit_r15_c96 bl[96] br[96] wl[15] vdd gnd cell_6t
Xbit_r16_c96 bl[96] br[96] wl[16] vdd gnd cell_6t
Xbit_r17_c96 bl[96] br[96] wl[17] vdd gnd cell_6t
Xbit_r18_c96 bl[96] br[96] wl[18] vdd gnd cell_6t
Xbit_r19_c96 bl[96] br[96] wl[19] vdd gnd cell_6t
Xbit_r20_c96 bl[96] br[96] wl[20] vdd gnd cell_6t
Xbit_r21_c96 bl[96] br[96] wl[21] vdd gnd cell_6t
Xbit_r22_c96 bl[96] br[96] wl[22] vdd gnd cell_6t
Xbit_r23_c96 bl[96] br[96] wl[23] vdd gnd cell_6t
Xbit_r24_c96 bl[96] br[96] wl[24] vdd gnd cell_6t
Xbit_r25_c96 bl[96] br[96] wl[25] vdd gnd cell_6t
Xbit_r26_c96 bl[96] br[96] wl[26] vdd gnd cell_6t
Xbit_r27_c96 bl[96] br[96] wl[27] vdd gnd cell_6t
Xbit_r28_c96 bl[96] br[96] wl[28] vdd gnd cell_6t
Xbit_r29_c96 bl[96] br[96] wl[29] vdd gnd cell_6t
Xbit_r30_c96 bl[96] br[96] wl[30] vdd gnd cell_6t
Xbit_r31_c96 bl[96] br[96] wl[31] vdd gnd cell_6t
Xbit_r32_c96 bl[96] br[96] wl[32] vdd gnd cell_6t
Xbit_r33_c96 bl[96] br[96] wl[33] vdd gnd cell_6t
Xbit_r34_c96 bl[96] br[96] wl[34] vdd gnd cell_6t
Xbit_r35_c96 bl[96] br[96] wl[35] vdd gnd cell_6t
Xbit_r36_c96 bl[96] br[96] wl[36] vdd gnd cell_6t
Xbit_r37_c96 bl[96] br[96] wl[37] vdd gnd cell_6t
Xbit_r38_c96 bl[96] br[96] wl[38] vdd gnd cell_6t
Xbit_r39_c96 bl[96] br[96] wl[39] vdd gnd cell_6t
Xbit_r40_c96 bl[96] br[96] wl[40] vdd gnd cell_6t
Xbit_r41_c96 bl[96] br[96] wl[41] vdd gnd cell_6t
Xbit_r42_c96 bl[96] br[96] wl[42] vdd gnd cell_6t
Xbit_r43_c96 bl[96] br[96] wl[43] vdd gnd cell_6t
Xbit_r44_c96 bl[96] br[96] wl[44] vdd gnd cell_6t
Xbit_r45_c96 bl[96] br[96] wl[45] vdd gnd cell_6t
Xbit_r46_c96 bl[96] br[96] wl[46] vdd gnd cell_6t
Xbit_r47_c96 bl[96] br[96] wl[47] vdd gnd cell_6t
Xbit_r48_c96 bl[96] br[96] wl[48] vdd gnd cell_6t
Xbit_r49_c96 bl[96] br[96] wl[49] vdd gnd cell_6t
Xbit_r50_c96 bl[96] br[96] wl[50] vdd gnd cell_6t
Xbit_r51_c96 bl[96] br[96] wl[51] vdd gnd cell_6t
Xbit_r52_c96 bl[96] br[96] wl[52] vdd gnd cell_6t
Xbit_r53_c96 bl[96] br[96] wl[53] vdd gnd cell_6t
Xbit_r54_c96 bl[96] br[96] wl[54] vdd gnd cell_6t
Xbit_r55_c96 bl[96] br[96] wl[55] vdd gnd cell_6t
Xbit_r56_c96 bl[96] br[96] wl[56] vdd gnd cell_6t
Xbit_r57_c96 bl[96] br[96] wl[57] vdd gnd cell_6t
Xbit_r58_c96 bl[96] br[96] wl[58] vdd gnd cell_6t
Xbit_r59_c96 bl[96] br[96] wl[59] vdd gnd cell_6t
Xbit_r60_c96 bl[96] br[96] wl[60] vdd gnd cell_6t
Xbit_r61_c96 bl[96] br[96] wl[61] vdd gnd cell_6t
Xbit_r62_c96 bl[96] br[96] wl[62] vdd gnd cell_6t
Xbit_r63_c96 bl[96] br[96] wl[63] vdd gnd cell_6t
Xbit_r64_c96 bl[96] br[96] wl[64] vdd gnd cell_6t
Xbit_r65_c96 bl[96] br[96] wl[65] vdd gnd cell_6t
Xbit_r66_c96 bl[96] br[96] wl[66] vdd gnd cell_6t
Xbit_r67_c96 bl[96] br[96] wl[67] vdd gnd cell_6t
Xbit_r68_c96 bl[96] br[96] wl[68] vdd gnd cell_6t
Xbit_r69_c96 bl[96] br[96] wl[69] vdd gnd cell_6t
Xbit_r70_c96 bl[96] br[96] wl[70] vdd gnd cell_6t
Xbit_r71_c96 bl[96] br[96] wl[71] vdd gnd cell_6t
Xbit_r72_c96 bl[96] br[96] wl[72] vdd gnd cell_6t
Xbit_r73_c96 bl[96] br[96] wl[73] vdd gnd cell_6t
Xbit_r74_c96 bl[96] br[96] wl[74] vdd gnd cell_6t
Xbit_r75_c96 bl[96] br[96] wl[75] vdd gnd cell_6t
Xbit_r76_c96 bl[96] br[96] wl[76] vdd gnd cell_6t
Xbit_r77_c96 bl[96] br[96] wl[77] vdd gnd cell_6t
Xbit_r78_c96 bl[96] br[96] wl[78] vdd gnd cell_6t
Xbit_r79_c96 bl[96] br[96] wl[79] vdd gnd cell_6t
Xbit_r80_c96 bl[96] br[96] wl[80] vdd gnd cell_6t
Xbit_r81_c96 bl[96] br[96] wl[81] vdd gnd cell_6t
Xbit_r82_c96 bl[96] br[96] wl[82] vdd gnd cell_6t
Xbit_r83_c96 bl[96] br[96] wl[83] vdd gnd cell_6t
Xbit_r84_c96 bl[96] br[96] wl[84] vdd gnd cell_6t
Xbit_r85_c96 bl[96] br[96] wl[85] vdd gnd cell_6t
Xbit_r86_c96 bl[96] br[96] wl[86] vdd gnd cell_6t
Xbit_r87_c96 bl[96] br[96] wl[87] vdd gnd cell_6t
Xbit_r88_c96 bl[96] br[96] wl[88] vdd gnd cell_6t
Xbit_r89_c96 bl[96] br[96] wl[89] vdd gnd cell_6t
Xbit_r90_c96 bl[96] br[96] wl[90] vdd gnd cell_6t
Xbit_r91_c96 bl[96] br[96] wl[91] vdd gnd cell_6t
Xbit_r92_c96 bl[96] br[96] wl[92] vdd gnd cell_6t
Xbit_r93_c96 bl[96] br[96] wl[93] vdd gnd cell_6t
Xbit_r94_c96 bl[96] br[96] wl[94] vdd gnd cell_6t
Xbit_r95_c96 bl[96] br[96] wl[95] vdd gnd cell_6t
Xbit_r96_c96 bl[96] br[96] wl[96] vdd gnd cell_6t
Xbit_r97_c96 bl[96] br[96] wl[97] vdd gnd cell_6t
Xbit_r98_c96 bl[96] br[96] wl[98] vdd gnd cell_6t
Xbit_r99_c96 bl[96] br[96] wl[99] vdd gnd cell_6t
Xbit_r100_c96 bl[96] br[96] wl[100] vdd gnd cell_6t
Xbit_r101_c96 bl[96] br[96] wl[101] vdd gnd cell_6t
Xbit_r102_c96 bl[96] br[96] wl[102] vdd gnd cell_6t
Xbit_r103_c96 bl[96] br[96] wl[103] vdd gnd cell_6t
Xbit_r104_c96 bl[96] br[96] wl[104] vdd gnd cell_6t
Xbit_r105_c96 bl[96] br[96] wl[105] vdd gnd cell_6t
Xbit_r106_c96 bl[96] br[96] wl[106] vdd gnd cell_6t
Xbit_r107_c96 bl[96] br[96] wl[107] vdd gnd cell_6t
Xbit_r108_c96 bl[96] br[96] wl[108] vdd gnd cell_6t
Xbit_r109_c96 bl[96] br[96] wl[109] vdd gnd cell_6t
Xbit_r110_c96 bl[96] br[96] wl[110] vdd gnd cell_6t
Xbit_r111_c96 bl[96] br[96] wl[111] vdd gnd cell_6t
Xbit_r112_c96 bl[96] br[96] wl[112] vdd gnd cell_6t
Xbit_r113_c96 bl[96] br[96] wl[113] vdd gnd cell_6t
Xbit_r114_c96 bl[96] br[96] wl[114] vdd gnd cell_6t
Xbit_r115_c96 bl[96] br[96] wl[115] vdd gnd cell_6t
Xbit_r116_c96 bl[96] br[96] wl[116] vdd gnd cell_6t
Xbit_r117_c96 bl[96] br[96] wl[117] vdd gnd cell_6t
Xbit_r118_c96 bl[96] br[96] wl[118] vdd gnd cell_6t
Xbit_r119_c96 bl[96] br[96] wl[119] vdd gnd cell_6t
Xbit_r120_c96 bl[96] br[96] wl[120] vdd gnd cell_6t
Xbit_r121_c96 bl[96] br[96] wl[121] vdd gnd cell_6t
Xbit_r122_c96 bl[96] br[96] wl[122] vdd gnd cell_6t
Xbit_r123_c96 bl[96] br[96] wl[123] vdd gnd cell_6t
Xbit_r124_c96 bl[96] br[96] wl[124] vdd gnd cell_6t
Xbit_r125_c96 bl[96] br[96] wl[125] vdd gnd cell_6t
Xbit_r126_c96 bl[96] br[96] wl[126] vdd gnd cell_6t
Xbit_r127_c96 bl[96] br[96] wl[127] vdd gnd cell_6t
Xbit_r0_c97 bl[97] br[97] wl[0] vdd gnd cell_6t
Xbit_r1_c97 bl[97] br[97] wl[1] vdd gnd cell_6t
Xbit_r2_c97 bl[97] br[97] wl[2] vdd gnd cell_6t
Xbit_r3_c97 bl[97] br[97] wl[3] vdd gnd cell_6t
Xbit_r4_c97 bl[97] br[97] wl[4] vdd gnd cell_6t
Xbit_r5_c97 bl[97] br[97] wl[5] vdd gnd cell_6t
Xbit_r6_c97 bl[97] br[97] wl[6] vdd gnd cell_6t
Xbit_r7_c97 bl[97] br[97] wl[7] vdd gnd cell_6t
Xbit_r8_c97 bl[97] br[97] wl[8] vdd gnd cell_6t
Xbit_r9_c97 bl[97] br[97] wl[9] vdd gnd cell_6t
Xbit_r10_c97 bl[97] br[97] wl[10] vdd gnd cell_6t
Xbit_r11_c97 bl[97] br[97] wl[11] vdd gnd cell_6t
Xbit_r12_c97 bl[97] br[97] wl[12] vdd gnd cell_6t
Xbit_r13_c97 bl[97] br[97] wl[13] vdd gnd cell_6t
Xbit_r14_c97 bl[97] br[97] wl[14] vdd gnd cell_6t
Xbit_r15_c97 bl[97] br[97] wl[15] vdd gnd cell_6t
Xbit_r16_c97 bl[97] br[97] wl[16] vdd gnd cell_6t
Xbit_r17_c97 bl[97] br[97] wl[17] vdd gnd cell_6t
Xbit_r18_c97 bl[97] br[97] wl[18] vdd gnd cell_6t
Xbit_r19_c97 bl[97] br[97] wl[19] vdd gnd cell_6t
Xbit_r20_c97 bl[97] br[97] wl[20] vdd gnd cell_6t
Xbit_r21_c97 bl[97] br[97] wl[21] vdd gnd cell_6t
Xbit_r22_c97 bl[97] br[97] wl[22] vdd gnd cell_6t
Xbit_r23_c97 bl[97] br[97] wl[23] vdd gnd cell_6t
Xbit_r24_c97 bl[97] br[97] wl[24] vdd gnd cell_6t
Xbit_r25_c97 bl[97] br[97] wl[25] vdd gnd cell_6t
Xbit_r26_c97 bl[97] br[97] wl[26] vdd gnd cell_6t
Xbit_r27_c97 bl[97] br[97] wl[27] vdd gnd cell_6t
Xbit_r28_c97 bl[97] br[97] wl[28] vdd gnd cell_6t
Xbit_r29_c97 bl[97] br[97] wl[29] vdd gnd cell_6t
Xbit_r30_c97 bl[97] br[97] wl[30] vdd gnd cell_6t
Xbit_r31_c97 bl[97] br[97] wl[31] vdd gnd cell_6t
Xbit_r32_c97 bl[97] br[97] wl[32] vdd gnd cell_6t
Xbit_r33_c97 bl[97] br[97] wl[33] vdd gnd cell_6t
Xbit_r34_c97 bl[97] br[97] wl[34] vdd gnd cell_6t
Xbit_r35_c97 bl[97] br[97] wl[35] vdd gnd cell_6t
Xbit_r36_c97 bl[97] br[97] wl[36] vdd gnd cell_6t
Xbit_r37_c97 bl[97] br[97] wl[37] vdd gnd cell_6t
Xbit_r38_c97 bl[97] br[97] wl[38] vdd gnd cell_6t
Xbit_r39_c97 bl[97] br[97] wl[39] vdd gnd cell_6t
Xbit_r40_c97 bl[97] br[97] wl[40] vdd gnd cell_6t
Xbit_r41_c97 bl[97] br[97] wl[41] vdd gnd cell_6t
Xbit_r42_c97 bl[97] br[97] wl[42] vdd gnd cell_6t
Xbit_r43_c97 bl[97] br[97] wl[43] vdd gnd cell_6t
Xbit_r44_c97 bl[97] br[97] wl[44] vdd gnd cell_6t
Xbit_r45_c97 bl[97] br[97] wl[45] vdd gnd cell_6t
Xbit_r46_c97 bl[97] br[97] wl[46] vdd gnd cell_6t
Xbit_r47_c97 bl[97] br[97] wl[47] vdd gnd cell_6t
Xbit_r48_c97 bl[97] br[97] wl[48] vdd gnd cell_6t
Xbit_r49_c97 bl[97] br[97] wl[49] vdd gnd cell_6t
Xbit_r50_c97 bl[97] br[97] wl[50] vdd gnd cell_6t
Xbit_r51_c97 bl[97] br[97] wl[51] vdd gnd cell_6t
Xbit_r52_c97 bl[97] br[97] wl[52] vdd gnd cell_6t
Xbit_r53_c97 bl[97] br[97] wl[53] vdd gnd cell_6t
Xbit_r54_c97 bl[97] br[97] wl[54] vdd gnd cell_6t
Xbit_r55_c97 bl[97] br[97] wl[55] vdd gnd cell_6t
Xbit_r56_c97 bl[97] br[97] wl[56] vdd gnd cell_6t
Xbit_r57_c97 bl[97] br[97] wl[57] vdd gnd cell_6t
Xbit_r58_c97 bl[97] br[97] wl[58] vdd gnd cell_6t
Xbit_r59_c97 bl[97] br[97] wl[59] vdd gnd cell_6t
Xbit_r60_c97 bl[97] br[97] wl[60] vdd gnd cell_6t
Xbit_r61_c97 bl[97] br[97] wl[61] vdd gnd cell_6t
Xbit_r62_c97 bl[97] br[97] wl[62] vdd gnd cell_6t
Xbit_r63_c97 bl[97] br[97] wl[63] vdd gnd cell_6t
Xbit_r64_c97 bl[97] br[97] wl[64] vdd gnd cell_6t
Xbit_r65_c97 bl[97] br[97] wl[65] vdd gnd cell_6t
Xbit_r66_c97 bl[97] br[97] wl[66] vdd gnd cell_6t
Xbit_r67_c97 bl[97] br[97] wl[67] vdd gnd cell_6t
Xbit_r68_c97 bl[97] br[97] wl[68] vdd gnd cell_6t
Xbit_r69_c97 bl[97] br[97] wl[69] vdd gnd cell_6t
Xbit_r70_c97 bl[97] br[97] wl[70] vdd gnd cell_6t
Xbit_r71_c97 bl[97] br[97] wl[71] vdd gnd cell_6t
Xbit_r72_c97 bl[97] br[97] wl[72] vdd gnd cell_6t
Xbit_r73_c97 bl[97] br[97] wl[73] vdd gnd cell_6t
Xbit_r74_c97 bl[97] br[97] wl[74] vdd gnd cell_6t
Xbit_r75_c97 bl[97] br[97] wl[75] vdd gnd cell_6t
Xbit_r76_c97 bl[97] br[97] wl[76] vdd gnd cell_6t
Xbit_r77_c97 bl[97] br[97] wl[77] vdd gnd cell_6t
Xbit_r78_c97 bl[97] br[97] wl[78] vdd gnd cell_6t
Xbit_r79_c97 bl[97] br[97] wl[79] vdd gnd cell_6t
Xbit_r80_c97 bl[97] br[97] wl[80] vdd gnd cell_6t
Xbit_r81_c97 bl[97] br[97] wl[81] vdd gnd cell_6t
Xbit_r82_c97 bl[97] br[97] wl[82] vdd gnd cell_6t
Xbit_r83_c97 bl[97] br[97] wl[83] vdd gnd cell_6t
Xbit_r84_c97 bl[97] br[97] wl[84] vdd gnd cell_6t
Xbit_r85_c97 bl[97] br[97] wl[85] vdd gnd cell_6t
Xbit_r86_c97 bl[97] br[97] wl[86] vdd gnd cell_6t
Xbit_r87_c97 bl[97] br[97] wl[87] vdd gnd cell_6t
Xbit_r88_c97 bl[97] br[97] wl[88] vdd gnd cell_6t
Xbit_r89_c97 bl[97] br[97] wl[89] vdd gnd cell_6t
Xbit_r90_c97 bl[97] br[97] wl[90] vdd gnd cell_6t
Xbit_r91_c97 bl[97] br[97] wl[91] vdd gnd cell_6t
Xbit_r92_c97 bl[97] br[97] wl[92] vdd gnd cell_6t
Xbit_r93_c97 bl[97] br[97] wl[93] vdd gnd cell_6t
Xbit_r94_c97 bl[97] br[97] wl[94] vdd gnd cell_6t
Xbit_r95_c97 bl[97] br[97] wl[95] vdd gnd cell_6t
Xbit_r96_c97 bl[97] br[97] wl[96] vdd gnd cell_6t
Xbit_r97_c97 bl[97] br[97] wl[97] vdd gnd cell_6t
Xbit_r98_c97 bl[97] br[97] wl[98] vdd gnd cell_6t
Xbit_r99_c97 bl[97] br[97] wl[99] vdd gnd cell_6t
Xbit_r100_c97 bl[97] br[97] wl[100] vdd gnd cell_6t
Xbit_r101_c97 bl[97] br[97] wl[101] vdd gnd cell_6t
Xbit_r102_c97 bl[97] br[97] wl[102] vdd gnd cell_6t
Xbit_r103_c97 bl[97] br[97] wl[103] vdd gnd cell_6t
Xbit_r104_c97 bl[97] br[97] wl[104] vdd gnd cell_6t
Xbit_r105_c97 bl[97] br[97] wl[105] vdd gnd cell_6t
Xbit_r106_c97 bl[97] br[97] wl[106] vdd gnd cell_6t
Xbit_r107_c97 bl[97] br[97] wl[107] vdd gnd cell_6t
Xbit_r108_c97 bl[97] br[97] wl[108] vdd gnd cell_6t
Xbit_r109_c97 bl[97] br[97] wl[109] vdd gnd cell_6t
Xbit_r110_c97 bl[97] br[97] wl[110] vdd gnd cell_6t
Xbit_r111_c97 bl[97] br[97] wl[111] vdd gnd cell_6t
Xbit_r112_c97 bl[97] br[97] wl[112] vdd gnd cell_6t
Xbit_r113_c97 bl[97] br[97] wl[113] vdd gnd cell_6t
Xbit_r114_c97 bl[97] br[97] wl[114] vdd gnd cell_6t
Xbit_r115_c97 bl[97] br[97] wl[115] vdd gnd cell_6t
Xbit_r116_c97 bl[97] br[97] wl[116] vdd gnd cell_6t
Xbit_r117_c97 bl[97] br[97] wl[117] vdd gnd cell_6t
Xbit_r118_c97 bl[97] br[97] wl[118] vdd gnd cell_6t
Xbit_r119_c97 bl[97] br[97] wl[119] vdd gnd cell_6t
Xbit_r120_c97 bl[97] br[97] wl[120] vdd gnd cell_6t
Xbit_r121_c97 bl[97] br[97] wl[121] vdd gnd cell_6t
Xbit_r122_c97 bl[97] br[97] wl[122] vdd gnd cell_6t
Xbit_r123_c97 bl[97] br[97] wl[123] vdd gnd cell_6t
Xbit_r124_c97 bl[97] br[97] wl[124] vdd gnd cell_6t
Xbit_r125_c97 bl[97] br[97] wl[125] vdd gnd cell_6t
Xbit_r126_c97 bl[97] br[97] wl[126] vdd gnd cell_6t
Xbit_r127_c97 bl[97] br[97] wl[127] vdd gnd cell_6t
Xbit_r0_c98 bl[98] br[98] wl[0] vdd gnd cell_6t
Xbit_r1_c98 bl[98] br[98] wl[1] vdd gnd cell_6t
Xbit_r2_c98 bl[98] br[98] wl[2] vdd gnd cell_6t
Xbit_r3_c98 bl[98] br[98] wl[3] vdd gnd cell_6t
Xbit_r4_c98 bl[98] br[98] wl[4] vdd gnd cell_6t
Xbit_r5_c98 bl[98] br[98] wl[5] vdd gnd cell_6t
Xbit_r6_c98 bl[98] br[98] wl[6] vdd gnd cell_6t
Xbit_r7_c98 bl[98] br[98] wl[7] vdd gnd cell_6t
Xbit_r8_c98 bl[98] br[98] wl[8] vdd gnd cell_6t
Xbit_r9_c98 bl[98] br[98] wl[9] vdd gnd cell_6t
Xbit_r10_c98 bl[98] br[98] wl[10] vdd gnd cell_6t
Xbit_r11_c98 bl[98] br[98] wl[11] vdd gnd cell_6t
Xbit_r12_c98 bl[98] br[98] wl[12] vdd gnd cell_6t
Xbit_r13_c98 bl[98] br[98] wl[13] vdd gnd cell_6t
Xbit_r14_c98 bl[98] br[98] wl[14] vdd gnd cell_6t
Xbit_r15_c98 bl[98] br[98] wl[15] vdd gnd cell_6t
Xbit_r16_c98 bl[98] br[98] wl[16] vdd gnd cell_6t
Xbit_r17_c98 bl[98] br[98] wl[17] vdd gnd cell_6t
Xbit_r18_c98 bl[98] br[98] wl[18] vdd gnd cell_6t
Xbit_r19_c98 bl[98] br[98] wl[19] vdd gnd cell_6t
Xbit_r20_c98 bl[98] br[98] wl[20] vdd gnd cell_6t
Xbit_r21_c98 bl[98] br[98] wl[21] vdd gnd cell_6t
Xbit_r22_c98 bl[98] br[98] wl[22] vdd gnd cell_6t
Xbit_r23_c98 bl[98] br[98] wl[23] vdd gnd cell_6t
Xbit_r24_c98 bl[98] br[98] wl[24] vdd gnd cell_6t
Xbit_r25_c98 bl[98] br[98] wl[25] vdd gnd cell_6t
Xbit_r26_c98 bl[98] br[98] wl[26] vdd gnd cell_6t
Xbit_r27_c98 bl[98] br[98] wl[27] vdd gnd cell_6t
Xbit_r28_c98 bl[98] br[98] wl[28] vdd gnd cell_6t
Xbit_r29_c98 bl[98] br[98] wl[29] vdd gnd cell_6t
Xbit_r30_c98 bl[98] br[98] wl[30] vdd gnd cell_6t
Xbit_r31_c98 bl[98] br[98] wl[31] vdd gnd cell_6t
Xbit_r32_c98 bl[98] br[98] wl[32] vdd gnd cell_6t
Xbit_r33_c98 bl[98] br[98] wl[33] vdd gnd cell_6t
Xbit_r34_c98 bl[98] br[98] wl[34] vdd gnd cell_6t
Xbit_r35_c98 bl[98] br[98] wl[35] vdd gnd cell_6t
Xbit_r36_c98 bl[98] br[98] wl[36] vdd gnd cell_6t
Xbit_r37_c98 bl[98] br[98] wl[37] vdd gnd cell_6t
Xbit_r38_c98 bl[98] br[98] wl[38] vdd gnd cell_6t
Xbit_r39_c98 bl[98] br[98] wl[39] vdd gnd cell_6t
Xbit_r40_c98 bl[98] br[98] wl[40] vdd gnd cell_6t
Xbit_r41_c98 bl[98] br[98] wl[41] vdd gnd cell_6t
Xbit_r42_c98 bl[98] br[98] wl[42] vdd gnd cell_6t
Xbit_r43_c98 bl[98] br[98] wl[43] vdd gnd cell_6t
Xbit_r44_c98 bl[98] br[98] wl[44] vdd gnd cell_6t
Xbit_r45_c98 bl[98] br[98] wl[45] vdd gnd cell_6t
Xbit_r46_c98 bl[98] br[98] wl[46] vdd gnd cell_6t
Xbit_r47_c98 bl[98] br[98] wl[47] vdd gnd cell_6t
Xbit_r48_c98 bl[98] br[98] wl[48] vdd gnd cell_6t
Xbit_r49_c98 bl[98] br[98] wl[49] vdd gnd cell_6t
Xbit_r50_c98 bl[98] br[98] wl[50] vdd gnd cell_6t
Xbit_r51_c98 bl[98] br[98] wl[51] vdd gnd cell_6t
Xbit_r52_c98 bl[98] br[98] wl[52] vdd gnd cell_6t
Xbit_r53_c98 bl[98] br[98] wl[53] vdd gnd cell_6t
Xbit_r54_c98 bl[98] br[98] wl[54] vdd gnd cell_6t
Xbit_r55_c98 bl[98] br[98] wl[55] vdd gnd cell_6t
Xbit_r56_c98 bl[98] br[98] wl[56] vdd gnd cell_6t
Xbit_r57_c98 bl[98] br[98] wl[57] vdd gnd cell_6t
Xbit_r58_c98 bl[98] br[98] wl[58] vdd gnd cell_6t
Xbit_r59_c98 bl[98] br[98] wl[59] vdd gnd cell_6t
Xbit_r60_c98 bl[98] br[98] wl[60] vdd gnd cell_6t
Xbit_r61_c98 bl[98] br[98] wl[61] vdd gnd cell_6t
Xbit_r62_c98 bl[98] br[98] wl[62] vdd gnd cell_6t
Xbit_r63_c98 bl[98] br[98] wl[63] vdd gnd cell_6t
Xbit_r64_c98 bl[98] br[98] wl[64] vdd gnd cell_6t
Xbit_r65_c98 bl[98] br[98] wl[65] vdd gnd cell_6t
Xbit_r66_c98 bl[98] br[98] wl[66] vdd gnd cell_6t
Xbit_r67_c98 bl[98] br[98] wl[67] vdd gnd cell_6t
Xbit_r68_c98 bl[98] br[98] wl[68] vdd gnd cell_6t
Xbit_r69_c98 bl[98] br[98] wl[69] vdd gnd cell_6t
Xbit_r70_c98 bl[98] br[98] wl[70] vdd gnd cell_6t
Xbit_r71_c98 bl[98] br[98] wl[71] vdd gnd cell_6t
Xbit_r72_c98 bl[98] br[98] wl[72] vdd gnd cell_6t
Xbit_r73_c98 bl[98] br[98] wl[73] vdd gnd cell_6t
Xbit_r74_c98 bl[98] br[98] wl[74] vdd gnd cell_6t
Xbit_r75_c98 bl[98] br[98] wl[75] vdd gnd cell_6t
Xbit_r76_c98 bl[98] br[98] wl[76] vdd gnd cell_6t
Xbit_r77_c98 bl[98] br[98] wl[77] vdd gnd cell_6t
Xbit_r78_c98 bl[98] br[98] wl[78] vdd gnd cell_6t
Xbit_r79_c98 bl[98] br[98] wl[79] vdd gnd cell_6t
Xbit_r80_c98 bl[98] br[98] wl[80] vdd gnd cell_6t
Xbit_r81_c98 bl[98] br[98] wl[81] vdd gnd cell_6t
Xbit_r82_c98 bl[98] br[98] wl[82] vdd gnd cell_6t
Xbit_r83_c98 bl[98] br[98] wl[83] vdd gnd cell_6t
Xbit_r84_c98 bl[98] br[98] wl[84] vdd gnd cell_6t
Xbit_r85_c98 bl[98] br[98] wl[85] vdd gnd cell_6t
Xbit_r86_c98 bl[98] br[98] wl[86] vdd gnd cell_6t
Xbit_r87_c98 bl[98] br[98] wl[87] vdd gnd cell_6t
Xbit_r88_c98 bl[98] br[98] wl[88] vdd gnd cell_6t
Xbit_r89_c98 bl[98] br[98] wl[89] vdd gnd cell_6t
Xbit_r90_c98 bl[98] br[98] wl[90] vdd gnd cell_6t
Xbit_r91_c98 bl[98] br[98] wl[91] vdd gnd cell_6t
Xbit_r92_c98 bl[98] br[98] wl[92] vdd gnd cell_6t
Xbit_r93_c98 bl[98] br[98] wl[93] vdd gnd cell_6t
Xbit_r94_c98 bl[98] br[98] wl[94] vdd gnd cell_6t
Xbit_r95_c98 bl[98] br[98] wl[95] vdd gnd cell_6t
Xbit_r96_c98 bl[98] br[98] wl[96] vdd gnd cell_6t
Xbit_r97_c98 bl[98] br[98] wl[97] vdd gnd cell_6t
Xbit_r98_c98 bl[98] br[98] wl[98] vdd gnd cell_6t
Xbit_r99_c98 bl[98] br[98] wl[99] vdd gnd cell_6t
Xbit_r100_c98 bl[98] br[98] wl[100] vdd gnd cell_6t
Xbit_r101_c98 bl[98] br[98] wl[101] vdd gnd cell_6t
Xbit_r102_c98 bl[98] br[98] wl[102] vdd gnd cell_6t
Xbit_r103_c98 bl[98] br[98] wl[103] vdd gnd cell_6t
Xbit_r104_c98 bl[98] br[98] wl[104] vdd gnd cell_6t
Xbit_r105_c98 bl[98] br[98] wl[105] vdd gnd cell_6t
Xbit_r106_c98 bl[98] br[98] wl[106] vdd gnd cell_6t
Xbit_r107_c98 bl[98] br[98] wl[107] vdd gnd cell_6t
Xbit_r108_c98 bl[98] br[98] wl[108] vdd gnd cell_6t
Xbit_r109_c98 bl[98] br[98] wl[109] vdd gnd cell_6t
Xbit_r110_c98 bl[98] br[98] wl[110] vdd gnd cell_6t
Xbit_r111_c98 bl[98] br[98] wl[111] vdd gnd cell_6t
Xbit_r112_c98 bl[98] br[98] wl[112] vdd gnd cell_6t
Xbit_r113_c98 bl[98] br[98] wl[113] vdd gnd cell_6t
Xbit_r114_c98 bl[98] br[98] wl[114] vdd gnd cell_6t
Xbit_r115_c98 bl[98] br[98] wl[115] vdd gnd cell_6t
Xbit_r116_c98 bl[98] br[98] wl[116] vdd gnd cell_6t
Xbit_r117_c98 bl[98] br[98] wl[117] vdd gnd cell_6t
Xbit_r118_c98 bl[98] br[98] wl[118] vdd gnd cell_6t
Xbit_r119_c98 bl[98] br[98] wl[119] vdd gnd cell_6t
Xbit_r120_c98 bl[98] br[98] wl[120] vdd gnd cell_6t
Xbit_r121_c98 bl[98] br[98] wl[121] vdd gnd cell_6t
Xbit_r122_c98 bl[98] br[98] wl[122] vdd gnd cell_6t
Xbit_r123_c98 bl[98] br[98] wl[123] vdd gnd cell_6t
Xbit_r124_c98 bl[98] br[98] wl[124] vdd gnd cell_6t
Xbit_r125_c98 bl[98] br[98] wl[125] vdd gnd cell_6t
Xbit_r126_c98 bl[98] br[98] wl[126] vdd gnd cell_6t
Xbit_r127_c98 bl[98] br[98] wl[127] vdd gnd cell_6t
Xbit_r0_c99 bl[99] br[99] wl[0] vdd gnd cell_6t
Xbit_r1_c99 bl[99] br[99] wl[1] vdd gnd cell_6t
Xbit_r2_c99 bl[99] br[99] wl[2] vdd gnd cell_6t
Xbit_r3_c99 bl[99] br[99] wl[3] vdd gnd cell_6t
Xbit_r4_c99 bl[99] br[99] wl[4] vdd gnd cell_6t
Xbit_r5_c99 bl[99] br[99] wl[5] vdd gnd cell_6t
Xbit_r6_c99 bl[99] br[99] wl[6] vdd gnd cell_6t
Xbit_r7_c99 bl[99] br[99] wl[7] vdd gnd cell_6t
Xbit_r8_c99 bl[99] br[99] wl[8] vdd gnd cell_6t
Xbit_r9_c99 bl[99] br[99] wl[9] vdd gnd cell_6t
Xbit_r10_c99 bl[99] br[99] wl[10] vdd gnd cell_6t
Xbit_r11_c99 bl[99] br[99] wl[11] vdd gnd cell_6t
Xbit_r12_c99 bl[99] br[99] wl[12] vdd gnd cell_6t
Xbit_r13_c99 bl[99] br[99] wl[13] vdd gnd cell_6t
Xbit_r14_c99 bl[99] br[99] wl[14] vdd gnd cell_6t
Xbit_r15_c99 bl[99] br[99] wl[15] vdd gnd cell_6t
Xbit_r16_c99 bl[99] br[99] wl[16] vdd gnd cell_6t
Xbit_r17_c99 bl[99] br[99] wl[17] vdd gnd cell_6t
Xbit_r18_c99 bl[99] br[99] wl[18] vdd gnd cell_6t
Xbit_r19_c99 bl[99] br[99] wl[19] vdd gnd cell_6t
Xbit_r20_c99 bl[99] br[99] wl[20] vdd gnd cell_6t
Xbit_r21_c99 bl[99] br[99] wl[21] vdd gnd cell_6t
Xbit_r22_c99 bl[99] br[99] wl[22] vdd gnd cell_6t
Xbit_r23_c99 bl[99] br[99] wl[23] vdd gnd cell_6t
Xbit_r24_c99 bl[99] br[99] wl[24] vdd gnd cell_6t
Xbit_r25_c99 bl[99] br[99] wl[25] vdd gnd cell_6t
Xbit_r26_c99 bl[99] br[99] wl[26] vdd gnd cell_6t
Xbit_r27_c99 bl[99] br[99] wl[27] vdd gnd cell_6t
Xbit_r28_c99 bl[99] br[99] wl[28] vdd gnd cell_6t
Xbit_r29_c99 bl[99] br[99] wl[29] vdd gnd cell_6t
Xbit_r30_c99 bl[99] br[99] wl[30] vdd gnd cell_6t
Xbit_r31_c99 bl[99] br[99] wl[31] vdd gnd cell_6t
Xbit_r32_c99 bl[99] br[99] wl[32] vdd gnd cell_6t
Xbit_r33_c99 bl[99] br[99] wl[33] vdd gnd cell_6t
Xbit_r34_c99 bl[99] br[99] wl[34] vdd gnd cell_6t
Xbit_r35_c99 bl[99] br[99] wl[35] vdd gnd cell_6t
Xbit_r36_c99 bl[99] br[99] wl[36] vdd gnd cell_6t
Xbit_r37_c99 bl[99] br[99] wl[37] vdd gnd cell_6t
Xbit_r38_c99 bl[99] br[99] wl[38] vdd gnd cell_6t
Xbit_r39_c99 bl[99] br[99] wl[39] vdd gnd cell_6t
Xbit_r40_c99 bl[99] br[99] wl[40] vdd gnd cell_6t
Xbit_r41_c99 bl[99] br[99] wl[41] vdd gnd cell_6t
Xbit_r42_c99 bl[99] br[99] wl[42] vdd gnd cell_6t
Xbit_r43_c99 bl[99] br[99] wl[43] vdd gnd cell_6t
Xbit_r44_c99 bl[99] br[99] wl[44] vdd gnd cell_6t
Xbit_r45_c99 bl[99] br[99] wl[45] vdd gnd cell_6t
Xbit_r46_c99 bl[99] br[99] wl[46] vdd gnd cell_6t
Xbit_r47_c99 bl[99] br[99] wl[47] vdd gnd cell_6t
Xbit_r48_c99 bl[99] br[99] wl[48] vdd gnd cell_6t
Xbit_r49_c99 bl[99] br[99] wl[49] vdd gnd cell_6t
Xbit_r50_c99 bl[99] br[99] wl[50] vdd gnd cell_6t
Xbit_r51_c99 bl[99] br[99] wl[51] vdd gnd cell_6t
Xbit_r52_c99 bl[99] br[99] wl[52] vdd gnd cell_6t
Xbit_r53_c99 bl[99] br[99] wl[53] vdd gnd cell_6t
Xbit_r54_c99 bl[99] br[99] wl[54] vdd gnd cell_6t
Xbit_r55_c99 bl[99] br[99] wl[55] vdd gnd cell_6t
Xbit_r56_c99 bl[99] br[99] wl[56] vdd gnd cell_6t
Xbit_r57_c99 bl[99] br[99] wl[57] vdd gnd cell_6t
Xbit_r58_c99 bl[99] br[99] wl[58] vdd gnd cell_6t
Xbit_r59_c99 bl[99] br[99] wl[59] vdd gnd cell_6t
Xbit_r60_c99 bl[99] br[99] wl[60] vdd gnd cell_6t
Xbit_r61_c99 bl[99] br[99] wl[61] vdd gnd cell_6t
Xbit_r62_c99 bl[99] br[99] wl[62] vdd gnd cell_6t
Xbit_r63_c99 bl[99] br[99] wl[63] vdd gnd cell_6t
Xbit_r64_c99 bl[99] br[99] wl[64] vdd gnd cell_6t
Xbit_r65_c99 bl[99] br[99] wl[65] vdd gnd cell_6t
Xbit_r66_c99 bl[99] br[99] wl[66] vdd gnd cell_6t
Xbit_r67_c99 bl[99] br[99] wl[67] vdd gnd cell_6t
Xbit_r68_c99 bl[99] br[99] wl[68] vdd gnd cell_6t
Xbit_r69_c99 bl[99] br[99] wl[69] vdd gnd cell_6t
Xbit_r70_c99 bl[99] br[99] wl[70] vdd gnd cell_6t
Xbit_r71_c99 bl[99] br[99] wl[71] vdd gnd cell_6t
Xbit_r72_c99 bl[99] br[99] wl[72] vdd gnd cell_6t
Xbit_r73_c99 bl[99] br[99] wl[73] vdd gnd cell_6t
Xbit_r74_c99 bl[99] br[99] wl[74] vdd gnd cell_6t
Xbit_r75_c99 bl[99] br[99] wl[75] vdd gnd cell_6t
Xbit_r76_c99 bl[99] br[99] wl[76] vdd gnd cell_6t
Xbit_r77_c99 bl[99] br[99] wl[77] vdd gnd cell_6t
Xbit_r78_c99 bl[99] br[99] wl[78] vdd gnd cell_6t
Xbit_r79_c99 bl[99] br[99] wl[79] vdd gnd cell_6t
Xbit_r80_c99 bl[99] br[99] wl[80] vdd gnd cell_6t
Xbit_r81_c99 bl[99] br[99] wl[81] vdd gnd cell_6t
Xbit_r82_c99 bl[99] br[99] wl[82] vdd gnd cell_6t
Xbit_r83_c99 bl[99] br[99] wl[83] vdd gnd cell_6t
Xbit_r84_c99 bl[99] br[99] wl[84] vdd gnd cell_6t
Xbit_r85_c99 bl[99] br[99] wl[85] vdd gnd cell_6t
Xbit_r86_c99 bl[99] br[99] wl[86] vdd gnd cell_6t
Xbit_r87_c99 bl[99] br[99] wl[87] vdd gnd cell_6t
Xbit_r88_c99 bl[99] br[99] wl[88] vdd gnd cell_6t
Xbit_r89_c99 bl[99] br[99] wl[89] vdd gnd cell_6t
Xbit_r90_c99 bl[99] br[99] wl[90] vdd gnd cell_6t
Xbit_r91_c99 bl[99] br[99] wl[91] vdd gnd cell_6t
Xbit_r92_c99 bl[99] br[99] wl[92] vdd gnd cell_6t
Xbit_r93_c99 bl[99] br[99] wl[93] vdd gnd cell_6t
Xbit_r94_c99 bl[99] br[99] wl[94] vdd gnd cell_6t
Xbit_r95_c99 bl[99] br[99] wl[95] vdd gnd cell_6t
Xbit_r96_c99 bl[99] br[99] wl[96] vdd gnd cell_6t
Xbit_r97_c99 bl[99] br[99] wl[97] vdd gnd cell_6t
Xbit_r98_c99 bl[99] br[99] wl[98] vdd gnd cell_6t
Xbit_r99_c99 bl[99] br[99] wl[99] vdd gnd cell_6t
Xbit_r100_c99 bl[99] br[99] wl[100] vdd gnd cell_6t
Xbit_r101_c99 bl[99] br[99] wl[101] vdd gnd cell_6t
Xbit_r102_c99 bl[99] br[99] wl[102] vdd gnd cell_6t
Xbit_r103_c99 bl[99] br[99] wl[103] vdd gnd cell_6t
Xbit_r104_c99 bl[99] br[99] wl[104] vdd gnd cell_6t
Xbit_r105_c99 bl[99] br[99] wl[105] vdd gnd cell_6t
Xbit_r106_c99 bl[99] br[99] wl[106] vdd gnd cell_6t
Xbit_r107_c99 bl[99] br[99] wl[107] vdd gnd cell_6t
Xbit_r108_c99 bl[99] br[99] wl[108] vdd gnd cell_6t
Xbit_r109_c99 bl[99] br[99] wl[109] vdd gnd cell_6t
Xbit_r110_c99 bl[99] br[99] wl[110] vdd gnd cell_6t
Xbit_r111_c99 bl[99] br[99] wl[111] vdd gnd cell_6t
Xbit_r112_c99 bl[99] br[99] wl[112] vdd gnd cell_6t
Xbit_r113_c99 bl[99] br[99] wl[113] vdd gnd cell_6t
Xbit_r114_c99 bl[99] br[99] wl[114] vdd gnd cell_6t
Xbit_r115_c99 bl[99] br[99] wl[115] vdd gnd cell_6t
Xbit_r116_c99 bl[99] br[99] wl[116] vdd gnd cell_6t
Xbit_r117_c99 bl[99] br[99] wl[117] vdd gnd cell_6t
Xbit_r118_c99 bl[99] br[99] wl[118] vdd gnd cell_6t
Xbit_r119_c99 bl[99] br[99] wl[119] vdd gnd cell_6t
Xbit_r120_c99 bl[99] br[99] wl[120] vdd gnd cell_6t
Xbit_r121_c99 bl[99] br[99] wl[121] vdd gnd cell_6t
Xbit_r122_c99 bl[99] br[99] wl[122] vdd gnd cell_6t
Xbit_r123_c99 bl[99] br[99] wl[123] vdd gnd cell_6t
Xbit_r124_c99 bl[99] br[99] wl[124] vdd gnd cell_6t
Xbit_r125_c99 bl[99] br[99] wl[125] vdd gnd cell_6t
Xbit_r126_c99 bl[99] br[99] wl[126] vdd gnd cell_6t
Xbit_r127_c99 bl[99] br[99] wl[127] vdd gnd cell_6t
Xbit_r0_c100 bl[100] br[100] wl[0] vdd gnd cell_6t
Xbit_r1_c100 bl[100] br[100] wl[1] vdd gnd cell_6t
Xbit_r2_c100 bl[100] br[100] wl[2] vdd gnd cell_6t
Xbit_r3_c100 bl[100] br[100] wl[3] vdd gnd cell_6t
Xbit_r4_c100 bl[100] br[100] wl[4] vdd gnd cell_6t
Xbit_r5_c100 bl[100] br[100] wl[5] vdd gnd cell_6t
Xbit_r6_c100 bl[100] br[100] wl[6] vdd gnd cell_6t
Xbit_r7_c100 bl[100] br[100] wl[7] vdd gnd cell_6t
Xbit_r8_c100 bl[100] br[100] wl[8] vdd gnd cell_6t
Xbit_r9_c100 bl[100] br[100] wl[9] vdd gnd cell_6t
Xbit_r10_c100 bl[100] br[100] wl[10] vdd gnd cell_6t
Xbit_r11_c100 bl[100] br[100] wl[11] vdd gnd cell_6t
Xbit_r12_c100 bl[100] br[100] wl[12] vdd gnd cell_6t
Xbit_r13_c100 bl[100] br[100] wl[13] vdd gnd cell_6t
Xbit_r14_c100 bl[100] br[100] wl[14] vdd gnd cell_6t
Xbit_r15_c100 bl[100] br[100] wl[15] vdd gnd cell_6t
Xbit_r16_c100 bl[100] br[100] wl[16] vdd gnd cell_6t
Xbit_r17_c100 bl[100] br[100] wl[17] vdd gnd cell_6t
Xbit_r18_c100 bl[100] br[100] wl[18] vdd gnd cell_6t
Xbit_r19_c100 bl[100] br[100] wl[19] vdd gnd cell_6t
Xbit_r20_c100 bl[100] br[100] wl[20] vdd gnd cell_6t
Xbit_r21_c100 bl[100] br[100] wl[21] vdd gnd cell_6t
Xbit_r22_c100 bl[100] br[100] wl[22] vdd gnd cell_6t
Xbit_r23_c100 bl[100] br[100] wl[23] vdd gnd cell_6t
Xbit_r24_c100 bl[100] br[100] wl[24] vdd gnd cell_6t
Xbit_r25_c100 bl[100] br[100] wl[25] vdd gnd cell_6t
Xbit_r26_c100 bl[100] br[100] wl[26] vdd gnd cell_6t
Xbit_r27_c100 bl[100] br[100] wl[27] vdd gnd cell_6t
Xbit_r28_c100 bl[100] br[100] wl[28] vdd gnd cell_6t
Xbit_r29_c100 bl[100] br[100] wl[29] vdd gnd cell_6t
Xbit_r30_c100 bl[100] br[100] wl[30] vdd gnd cell_6t
Xbit_r31_c100 bl[100] br[100] wl[31] vdd gnd cell_6t
Xbit_r32_c100 bl[100] br[100] wl[32] vdd gnd cell_6t
Xbit_r33_c100 bl[100] br[100] wl[33] vdd gnd cell_6t
Xbit_r34_c100 bl[100] br[100] wl[34] vdd gnd cell_6t
Xbit_r35_c100 bl[100] br[100] wl[35] vdd gnd cell_6t
Xbit_r36_c100 bl[100] br[100] wl[36] vdd gnd cell_6t
Xbit_r37_c100 bl[100] br[100] wl[37] vdd gnd cell_6t
Xbit_r38_c100 bl[100] br[100] wl[38] vdd gnd cell_6t
Xbit_r39_c100 bl[100] br[100] wl[39] vdd gnd cell_6t
Xbit_r40_c100 bl[100] br[100] wl[40] vdd gnd cell_6t
Xbit_r41_c100 bl[100] br[100] wl[41] vdd gnd cell_6t
Xbit_r42_c100 bl[100] br[100] wl[42] vdd gnd cell_6t
Xbit_r43_c100 bl[100] br[100] wl[43] vdd gnd cell_6t
Xbit_r44_c100 bl[100] br[100] wl[44] vdd gnd cell_6t
Xbit_r45_c100 bl[100] br[100] wl[45] vdd gnd cell_6t
Xbit_r46_c100 bl[100] br[100] wl[46] vdd gnd cell_6t
Xbit_r47_c100 bl[100] br[100] wl[47] vdd gnd cell_6t
Xbit_r48_c100 bl[100] br[100] wl[48] vdd gnd cell_6t
Xbit_r49_c100 bl[100] br[100] wl[49] vdd gnd cell_6t
Xbit_r50_c100 bl[100] br[100] wl[50] vdd gnd cell_6t
Xbit_r51_c100 bl[100] br[100] wl[51] vdd gnd cell_6t
Xbit_r52_c100 bl[100] br[100] wl[52] vdd gnd cell_6t
Xbit_r53_c100 bl[100] br[100] wl[53] vdd gnd cell_6t
Xbit_r54_c100 bl[100] br[100] wl[54] vdd gnd cell_6t
Xbit_r55_c100 bl[100] br[100] wl[55] vdd gnd cell_6t
Xbit_r56_c100 bl[100] br[100] wl[56] vdd gnd cell_6t
Xbit_r57_c100 bl[100] br[100] wl[57] vdd gnd cell_6t
Xbit_r58_c100 bl[100] br[100] wl[58] vdd gnd cell_6t
Xbit_r59_c100 bl[100] br[100] wl[59] vdd gnd cell_6t
Xbit_r60_c100 bl[100] br[100] wl[60] vdd gnd cell_6t
Xbit_r61_c100 bl[100] br[100] wl[61] vdd gnd cell_6t
Xbit_r62_c100 bl[100] br[100] wl[62] vdd gnd cell_6t
Xbit_r63_c100 bl[100] br[100] wl[63] vdd gnd cell_6t
Xbit_r64_c100 bl[100] br[100] wl[64] vdd gnd cell_6t
Xbit_r65_c100 bl[100] br[100] wl[65] vdd gnd cell_6t
Xbit_r66_c100 bl[100] br[100] wl[66] vdd gnd cell_6t
Xbit_r67_c100 bl[100] br[100] wl[67] vdd gnd cell_6t
Xbit_r68_c100 bl[100] br[100] wl[68] vdd gnd cell_6t
Xbit_r69_c100 bl[100] br[100] wl[69] vdd gnd cell_6t
Xbit_r70_c100 bl[100] br[100] wl[70] vdd gnd cell_6t
Xbit_r71_c100 bl[100] br[100] wl[71] vdd gnd cell_6t
Xbit_r72_c100 bl[100] br[100] wl[72] vdd gnd cell_6t
Xbit_r73_c100 bl[100] br[100] wl[73] vdd gnd cell_6t
Xbit_r74_c100 bl[100] br[100] wl[74] vdd gnd cell_6t
Xbit_r75_c100 bl[100] br[100] wl[75] vdd gnd cell_6t
Xbit_r76_c100 bl[100] br[100] wl[76] vdd gnd cell_6t
Xbit_r77_c100 bl[100] br[100] wl[77] vdd gnd cell_6t
Xbit_r78_c100 bl[100] br[100] wl[78] vdd gnd cell_6t
Xbit_r79_c100 bl[100] br[100] wl[79] vdd gnd cell_6t
Xbit_r80_c100 bl[100] br[100] wl[80] vdd gnd cell_6t
Xbit_r81_c100 bl[100] br[100] wl[81] vdd gnd cell_6t
Xbit_r82_c100 bl[100] br[100] wl[82] vdd gnd cell_6t
Xbit_r83_c100 bl[100] br[100] wl[83] vdd gnd cell_6t
Xbit_r84_c100 bl[100] br[100] wl[84] vdd gnd cell_6t
Xbit_r85_c100 bl[100] br[100] wl[85] vdd gnd cell_6t
Xbit_r86_c100 bl[100] br[100] wl[86] vdd gnd cell_6t
Xbit_r87_c100 bl[100] br[100] wl[87] vdd gnd cell_6t
Xbit_r88_c100 bl[100] br[100] wl[88] vdd gnd cell_6t
Xbit_r89_c100 bl[100] br[100] wl[89] vdd gnd cell_6t
Xbit_r90_c100 bl[100] br[100] wl[90] vdd gnd cell_6t
Xbit_r91_c100 bl[100] br[100] wl[91] vdd gnd cell_6t
Xbit_r92_c100 bl[100] br[100] wl[92] vdd gnd cell_6t
Xbit_r93_c100 bl[100] br[100] wl[93] vdd gnd cell_6t
Xbit_r94_c100 bl[100] br[100] wl[94] vdd gnd cell_6t
Xbit_r95_c100 bl[100] br[100] wl[95] vdd gnd cell_6t
Xbit_r96_c100 bl[100] br[100] wl[96] vdd gnd cell_6t
Xbit_r97_c100 bl[100] br[100] wl[97] vdd gnd cell_6t
Xbit_r98_c100 bl[100] br[100] wl[98] vdd gnd cell_6t
Xbit_r99_c100 bl[100] br[100] wl[99] vdd gnd cell_6t
Xbit_r100_c100 bl[100] br[100] wl[100] vdd gnd cell_6t
Xbit_r101_c100 bl[100] br[100] wl[101] vdd gnd cell_6t
Xbit_r102_c100 bl[100] br[100] wl[102] vdd gnd cell_6t
Xbit_r103_c100 bl[100] br[100] wl[103] vdd gnd cell_6t
Xbit_r104_c100 bl[100] br[100] wl[104] vdd gnd cell_6t
Xbit_r105_c100 bl[100] br[100] wl[105] vdd gnd cell_6t
Xbit_r106_c100 bl[100] br[100] wl[106] vdd gnd cell_6t
Xbit_r107_c100 bl[100] br[100] wl[107] vdd gnd cell_6t
Xbit_r108_c100 bl[100] br[100] wl[108] vdd gnd cell_6t
Xbit_r109_c100 bl[100] br[100] wl[109] vdd gnd cell_6t
Xbit_r110_c100 bl[100] br[100] wl[110] vdd gnd cell_6t
Xbit_r111_c100 bl[100] br[100] wl[111] vdd gnd cell_6t
Xbit_r112_c100 bl[100] br[100] wl[112] vdd gnd cell_6t
Xbit_r113_c100 bl[100] br[100] wl[113] vdd gnd cell_6t
Xbit_r114_c100 bl[100] br[100] wl[114] vdd gnd cell_6t
Xbit_r115_c100 bl[100] br[100] wl[115] vdd gnd cell_6t
Xbit_r116_c100 bl[100] br[100] wl[116] vdd gnd cell_6t
Xbit_r117_c100 bl[100] br[100] wl[117] vdd gnd cell_6t
Xbit_r118_c100 bl[100] br[100] wl[118] vdd gnd cell_6t
Xbit_r119_c100 bl[100] br[100] wl[119] vdd gnd cell_6t
Xbit_r120_c100 bl[100] br[100] wl[120] vdd gnd cell_6t
Xbit_r121_c100 bl[100] br[100] wl[121] vdd gnd cell_6t
Xbit_r122_c100 bl[100] br[100] wl[122] vdd gnd cell_6t
Xbit_r123_c100 bl[100] br[100] wl[123] vdd gnd cell_6t
Xbit_r124_c100 bl[100] br[100] wl[124] vdd gnd cell_6t
Xbit_r125_c100 bl[100] br[100] wl[125] vdd gnd cell_6t
Xbit_r126_c100 bl[100] br[100] wl[126] vdd gnd cell_6t
Xbit_r127_c100 bl[100] br[100] wl[127] vdd gnd cell_6t
Xbit_r0_c101 bl[101] br[101] wl[0] vdd gnd cell_6t
Xbit_r1_c101 bl[101] br[101] wl[1] vdd gnd cell_6t
Xbit_r2_c101 bl[101] br[101] wl[2] vdd gnd cell_6t
Xbit_r3_c101 bl[101] br[101] wl[3] vdd gnd cell_6t
Xbit_r4_c101 bl[101] br[101] wl[4] vdd gnd cell_6t
Xbit_r5_c101 bl[101] br[101] wl[5] vdd gnd cell_6t
Xbit_r6_c101 bl[101] br[101] wl[6] vdd gnd cell_6t
Xbit_r7_c101 bl[101] br[101] wl[7] vdd gnd cell_6t
Xbit_r8_c101 bl[101] br[101] wl[8] vdd gnd cell_6t
Xbit_r9_c101 bl[101] br[101] wl[9] vdd gnd cell_6t
Xbit_r10_c101 bl[101] br[101] wl[10] vdd gnd cell_6t
Xbit_r11_c101 bl[101] br[101] wl[11] vdd gnd cell_6t
Xbit_r12_c101 bl[101] br[101] wl[12] vdd gnd cell_6t
Xbit_r13_c101 bl[101] br[101] wl[13] vdd gnd cell_6t
Xbit_r14_c101 bl[101] br[101] wl[14] vdd gnd cell_6t
Xbit_r15_c101 bl[101] br[101] wl[15] vdd gnd cell_6t
Xbit_r16_c101 bl[101] br[101] wl[16] vdd gnd cell_6t
Xbit_r17_c101 bl[101] br[101] wl[17] vdd gnd cell_6t
Xbit_r18_c101 bl[101] br[101] wl[18] vdd gnd cell_6t
Xbit_r19_c101 bl[101] br[101] wl[19] vdd gnd cell_6t
Xbit_r20_c101 bl[101] br[101] wl[20] vdd gnd cell_6t
Xbit_r21_c101 bl[101] br[101] wl[21] vdd gnd cell_6t
Xbit_r22_c101 bl[101] br[101] wl[22] vdd gnd cell_6t
Xbit_r23_c101 bl[101] br[101] wl[23] vdd gnd cell_6t
Xbit_r24_c101 bl[101] br[101] wl[24] vdd gnd cell_6t
Xbit_r25_c101 bl[101] br[101] wl[25] vdd gnd cell_6t
Xbit_r26_c101 bl[101] br[101] wl[26] vdd gnd cell_6t
Xbit_r27_c101 bl[101] br[101] wl[27] vdd gnd cell_6t
Xbit_r28_c101 bl[101] br[101] wl[28] vdd gnd cell_6t
Xbit_r29_c101 bl[101] br[101] wl[29] vdd gnd cell_6t
Xbit_r30_c101 bl[101] br[101] wl[30] vdd gnd cell_6t
Xbit_r31_c101 bl[101] br[101] wl[31] vdd gnd cell_6t
Xbit_r32_c101 bl[101] br[101] wl[32] vdd gnd cell_6t
Xbit_r33_c101 bl[101] br[101] wl[33] vdd gnd cell_6t
Xbit_r34_c101 bl[101] br[101] wl[34] vdd gnd cell_6t
Xbit_r35_c101 bl[101] br[101] wl[35] vdd gnd cell_6t
Xbit_r36_c101 bl[101] br[101] wl[36] vdd gnd cell_6t
Xbit_r37_c101 bl[101] br[101] wl[37] vdd gnd cell_6t
Xbit_r38_c101 bl[101] br[101] wl[38] vdd gnd cell_6t
Xbit_r39_c101 bl[101] br[101] wl[39] vdd gnd cell_6t
Xbit_r40_c101 bl[101] br[101] wl[40] vdd gnd cell_6t
Xbit_r41_c101 bl[101] br[101] wl[41] vdd gnd cell_6t
Xbit_r42_c101 bl[101] br[101] wl[42] vdd gnd cell_6t
Xbit_r43_c101 bl[101] br[101] wl[43] vdd gnd cell_6t
Xbit_r44_c101 bl[101] br[101] wl[44] vdd gnd cell_6t
Xbit_r45_c101 bl[101] br[101] wl[45] vdd gnd cell_6t
Xbit_r46_c101 bl[101] br[101] wl[46] vdd gnd cell_6t
Xbit_r47_c101 bl[101] br[101] wl[47] vdd gnd cell_6t
Xbit_r48_c101 bl[101] br[101] wl[48] vdd gnd cell_6t
Xbit_r49_c101 bl[101] br[101] wl[49] vdd gnd cell_6t
Xbit_r50_c101 bl[101] br[101] wl[50] vdd gnd cell_6t
Xbit_r51_c101 bl[101] br[101] wl[51] vdd gnd cell_6t
Xbit_r52_c101 bl[101] br[101] wl[52] vdd gnd cell_6t
Xbit_r53_c101 bl[101] br[101] wl[53] vdd gnd cell_6t
Xbit_r54_c101 bl[101] br[101] wl[54] vdd gnd cell_6t
Xbit_r55_c101 bl[101] br[101] wl[55] vdd gnd cell_6t
Xbit_r56_c101 bl[101] br[101] wl[56] vdd gnd cell_6t
Xbit_r57_c101 bl[101] br[101] wl[57] vdd gnd cell_6t
Xbit_r58_c101 bl[101] br[101] wl[58] vdd gnd cell_6t
Xbit_r59_c101 bl[101] br[101] wl[59] vdd gnd cell_6t
Xbit_r60_c101 bl[101] br[101] wl[60] vdd gnd cell_6t
Xbit_r61_c101 bl[101] br[101] wl[61] vdd gnd cell_6t
Xbit_r62_c101 bl[101] br[101] wl[62] vdd gnd cell_6t
Xbit_r63_c101 bl[101] br[101] wl[63] vdd gnd cell_6t
Xbit_r64_c101 bl[101] br[101] wl[64] vdd gnd cell_6t
Xbit_r65_c101 bl[101] br[101] wl[65] vdd gnd cell_6t
Xbit_r66_c101 bl[101] br[101] wl[66] vdd gnd cell_6t
Xbit_r67_c101 bl[101] br[101] wl[67] vdd gnd cell_6t
Xbit_r68_c101 bl[101] br[101] wl[68] vdd gnd cell_6t
Xbit_r69_c101 bl[101] br[101] wl[69] vdd gnd cell_6t
Xbit_r70_c101 bl[101] br[101] wl[70] vdd gnd cell_6t
Xbit_r71_c101 bl[101] br[101] wl[71] vdd gnd cell_6t
Xbit_r72_c101 bl[101] br[101] wl[72] vdd gnd cell_6t
Xbit_r73_c101 bl[101] br[101] wl[73] vdd gnd cell_6t
Xbit_r74_c101 bl[101] br[101] wl[74] vdd gnd cell_6t
Xbit_r75_c101 bl[101] br[101] wl[75] vdd gnd cell_6t
Xbit_r76_c101 bl[101] br[101] wl[76] vdd gnd cell_6t
Xbit_r77_c101 bl[101] br[101] wl[77] vdd gnd cell_6t
Xbit_r78_c101 bl[101] br[101] wl[78] vdd gnd cell_6t
Xbit_r79_c101 bl[101] br[101] wl[79] vdd gnd cell_6t
Xbit_r80_c101 bl[101] br[101] wl[80] vdd gnd cell_6t
Xbit_r81_c101 bl[101] br[101] wl[81] vdd gnd cell_6t
Xbit_r82_c101 bl[101] br[101] wl[82] vdd gnd cell_6t
Xbit_r83_c101 bl[101] br[101] wl[83] vdd gnd cell_6t
Xbit_r84_c101 bl[101] br[101] wl[84] vdd gnd cell_6t
Xbit_r85_c101 bl[101] br[101] wl[85] vdd gnd cell_6t
Xbit_r86_c101 bl[101] br[101] wl[86] vdd gnd cell_6t
Xbit_r87_c101 bl[101] br[101] wl[87] vdd gnd cell_6t
Xbit_r88_c101 bl[101] br[101] wl[88] vdd gnd cell_6t
Xbit_r89_c101 bl[101] br[101] wl[89] vdd gnd cell_6t
Xbit_r90_c101 bl[101] br[101] wl[90] vdd gnd cell_6t
Xbit_r91_c101 bl[101] br[101] wl[91] vdd gnd cell_6t
Xbit_r92_c101 bl[101] br[101] wl[92] vdd gnd cell_6t
Xbit_r93_c101 bl[101] br[101] wl[93] vdd gnd cell_6t
Xbit_r94_c101 bl[101] br[101] wl[94] vdd gnd cell_6t
Xbit_r95_c101 bl[101] br[101] wl[95] vdd gnd cell_6t
Xbit_r96_c101 bl[101] br[101] wl[96] vdd gnd cell_6t
Xbit_r97_c101 bl[101] br[101] wl[97] vdd gnd cell_6t
Xbit_r98_c101 bl[101] br[101] wl[98] vdd gnd cell_6t
Xbit_r99_c101 bl[101] br[101] wl[99] vdd gnd cell_6t
Xbit_r100_c101 bl[101] br[101] wl[100] vdd gnd cell_6t
Xbit_r101_c101 bl[101] br[101] wl[101] vdd gnd cell_6t
Xbit_r102_c101 bl[101] br[101] wl[102] vdd gnd cell_6t
Xbit_r103_c101 bl[101] br[101] wl[103] vdd gnd cell_6t
Xbit_r104_c101 bl[101] br[101] wl[104] vdd gnd cell_6t
Xbit_r105_c101 bl[101] br[101] wl[105] vdd gnd cell_6t
Xbit_r106_c101 bl[101] br[101] wl[106] vdd gnd cell_6t
Xbit_r107_c101 bl[101] br[101] wl[107] vdd gnd cell_6t
Xbit_r108_c101 bl[101] br[101] wl[108] vdd gnd cell_6t
Xbit_r109_c101 bl[101] br[101] wl[109] vdd gnd cell_6t
Xbit_r110_c101 bl[101] br[101] wl[110] vdd gnd cell_6t
Xbit_r111_c101 bl[101] br[101] wl[111] vdd gnd cell_6t
Xbit_r112_c101 bl[101] br[101] wl[112] vdd gnd cell_6t
Xbit_r113_c101 bl[101] br[101] wl[113] vdd gnd cell_6t
Xbit_r114_c101 bl[101] br[101] wl[114] vdd gnd cell_6t
Xbit_r115_c101 bl[101] br[101] wl[115] vdd gnd cell_6t
Xbit_r116_c101 bl[101] br[101] wl[116] vdd gnd cell_6t
Xbit_r117_c101 bl[101] br[101] wl[117] vdd gnd cell_6t
Xbit_r118_c101 bl[101] br[101] wl[118] vdd gnd cell_6t
Xbit_r119_c101 bl[101] br[101] wl[119] vdd gnd cell_6t
Xbit_r120_c101 bl[101] br[101] wl[120] vdd gnd cell_6t
Xbit_r121_c101 bl[101] br[101] wl[121] vdd gnd cell_6t
Xbit_r122_c101 bl[101] br[101] wl[122] vdd gnd cell_6t
Xbit_r123_c101 bl[101] br[101] wl[123] vdd gnd cell_6t
Xbit_r124_c101 bl[101] br[101] wl[124] vdd gnd cell_6t
Xbit_r125_c101 bl[101] br[101] wl[125] vdd gnd cell_6t
Xbit_r126_c101 bl[101] br[101] wl[126] vdd gnd cell_6t
Xbit_r127_c101 bl[101] br[101] wl[127] vdd gnd cell_6t
Xbit_r0_c102 bl[102] br[102] wl[0] vdd gnd cell_6t
Xbit_r1_c102 bl[102] br[102] wl[1] vdd gnd cell_6t
Xbit_r2_c102 bl[102] br[102] wl[2] vdd gnd cell_6t
Xbit_r3_c102 bl[102] br[102] wl[3] vdd gnd cell_6t
Xbit_r4_c102 bl[102] br[102] wl[4] vdd gnd cell_6t
Xbit_r5_c102 bl[102] br[102] wl[5] vdd gnd cell_6t
Xbit_r6_c102 bl[102] br[102] wl[6] vdd gnd cell_6t
Xbit_r7_c102 bl[102] br[102] wl[7] vdd gnd cell_6t
Xbit_r8_c102 bl[102] br[102] wl[8] vdd gnd cell_6t
Xbit_r9_c102 bl[102] br[102] wl[9] vdd gnd cell_6t
Xbit_r10_c102 bl[102] br[102] wl[10] vdd gnd cell_6t
Xbit_r11_c102 bl[102] br[102] wl[11] vdd gnd cell_6t
Xbit_r12_c102 bl[102] br[102] wl[12] vdd gnd cell_6t
Xbit_r13_c102 bl[102] br[102] wl[13] vdd gnd cell_6t
Xbit_r14_c102 bl[102] br[102] wl[14] vdd gnd cell_6t
Xbit_r15_c102 bl[102] br[102] wl[15] vdd gnd cell_6t
Xbit_r16_c102 bl[102] br[102] wl[16] vdd gnd cell_6t
Xbit_r17_c102 bl[102] br[102] wl[17] vdd gnd cell_6t
Xbit_r18_c102 bl[102] br[102] wl[18] vdd gnd cell_6t
Xbit_r19_c102 bl[102] br[102] wl[19] vdd gnd cell_6t
Xbit_r20_c102 bl[102] br[102] wl[20] vdd gnd cell_6t
Xbit_r21_c102 bl[102] br[102] wl[21] vdd gnd cell_6t
Xbit_r22_c102 bl[102] br[102] wl[22] vdd gnd cell_6t
Xbit_r23_c102 bl[102] br[102] wl[23] vdd gnd cell_6t
Xbit_r24_c102 bl[102] br[102] wl[24] vdd gnd cell_6t
Xbit_r25_c102 bl[102] br[102] wl[25] vdd gnd cell_6t
Xbit_r26_c102 bl[102] br[102] wl[26] vdd gnd cell_6t
Xbit_r27_c102 bl[102] br[102] wl[27] vdd gnd cell_6t
Xbit_r28_c102 bl[102] br[102] wl[28] vdd gnd cell_6t
Xbit_r29_c102 bl[102] br[102] wl[29] vdd gnd cell_6t
Xbit_r30_c102 bl[102] br[102] wl[30] vdd gnd cell_6t
Xbit_r31_c102 bl[102] br[102] wl[31] vdd gnd cell_6t
Xbit_r32_c102 bl[102] br[102] wl[32] vdd gnd cell_6t
Xbit_r33_c102 bl[102] br[102] wl[33] vdd gnd cell_6t
Xbit_r34_c102 bl[102] br[102] wl[34] vdd gnd cell_6t
Xbit_r35_c102 bl[102] br[102] wl[35] vdd gnd cell_6t
Xbit_r36_c102 bl[102] br[102] wl[36] vdd gnd cell_6t
Xbit_r37_c102 bl[102] br[102] wl[37] vdd gnd cell_6t
Xbit_r38_c102 bl[102] br[102] wl[38] vdd gnd cell_6t
Xbit_r39_c102 bl[102] br[102] wl[39] vdd gnd cell_6t
Xbit_r40_c102 bl[102] br[102] wl[40] vdd gnd cell_6t
Xbit_r41_c102 bl[102] br[102] wl[41] vdd gnd cell_6t
Xbit_r42_c102 bl[102] br[102] wl[42] vdd gnd cell_6t
Xbit_r43_c102 bl[102] br[102] wl[43] vdd gnd cell_6t
Xbit_r44_c102 bl[102] br[102] wl[44] vdd gnd cell_6t
Xbit_r45_c102 bl[102] br[102] wl[45] vdd gnd cell_6t
Xbit_r46_c102 bl[102] br[102] wl[46] vdd gnd cell_6t
Xbit_r47_c102 bl[102] br[102] wl[47] vdd gnd cell_6t
Xbit_r48_c102 bl[102] br[102] wl[48] vdd gnd cell_6t
Xbit_r49_c102 bl[102] br[102] wl[49] vdd gnd cell_6t
Xbit_r50_c102 bl[102] br[102] wl[50] vdd gnd cell_6t
Xbit_r51_c102 bl[102] br[102] wl[51] vdd gnd cell_6t
Xbit_r52_c102 bl[102] br[102] wl[52] vdd gnd cell_6t
Xbit_r53_c102 bl[102] br[102] wl[53] vdd gnd cell_6t
Xbit_r54_c102 bl[102] br[102] wl[54] vdd gnd cell_6t
Xbit_r55_c102 bl[102] br[102] wl[55] vdd gnd cell_6t
Xbit_r56_c102 bl[102] br[102] wl[56] vdd gnd cell_6t
Xbit_r57_c102 bl[102] br[102] wl[57] vdd gnd cell_6t
Xbit_r58_c102 bl[102] br[102] wl[58] vdd gnd cell_6t
Xbit_r59_c102 bl[102] br[102] wl[59] vdd gnd cell_6t
Xbit_r60_c102 bl[102] br[102] wl[60] vdd gnd cell_6t
Xbit_r61_c102 bl[102] br[102] wl[61] vdd gnd cell_6t
Xbit_r62_c102 bl[102] br[102] wl[62] vdd gnd cell_6t
Xbit_r63_c102 bl[102] br[102] wl[63] vdd gnd cell_6t
Xbit_r64_c102 bl[102] br[102] wl[64] vdd gnd cell_6t
Xbit_r65_c102 bl[102] br[102] wl[65] vdd gnd cell_6t
Xbit_r66_c102 bl[102] br[102] wl[66] vdd gnd cell_6t
Xbit_r67_c102 bl[102] br[102] wl[67] vdd gnd cell_6t
Xbit_r68_c102 bl[102] br[102] wl[68] vdd gnd cell_6t
Xbit_r69_c102 bl[102] br[102] wl[69] vdd gnd cell_6t
Xbit_r70_c102 bl[102] br[102] wl[70] vdd gnd cell_6t
Xbit_r71_c102 bl[102] br[102] wl[71] vdd gnd cell_6t
Xbit_r72_c102 bl[102] br[102] wl[72] vdd gnd cell_6t
Xbit_r73_c102 bl[102] br[102] wl[73] vdd gnd cell_6t
Xbit_r74_c102 bl[102] br[102] wl[74] vdd gnd cell_6t
Xbit_r75_c102 bl[102] br[102] wl[75] vdd gnd cell_6t
Xbit_r76_c102 bl[102] br[102] wl[76] vdd gnd cell_6t
Xbit_r77_c102 bl[102] br[102] wl[77] vdd gnd cell_6t
Xbit_r78_c102 bl[102] br[102] wl[78] vdd gnd cell_6t
Xbit_r79_c102 bl[102] br[102] wl[79] vdd gnd cell_6t
Xbit_r80_c102 bl[102] br[102] wl[80] vdd gnd cell_6t
Xbit_r81_c102 bl[102] br[102] wl[81] vdd gnd cell_6t
Xbit_r82_c102 bl[102] br[102] wl[82] vdd gnd cell_6t
Xbit_r83_c102 bl[102] br[102] wl[83] vdd gnd cell_6t
Xbit_r84_c102 bl[102] br[102] wl[84] vdd gnd cell_6t
Xbit_r85_c102 bl[102] br[102] wl[85] vdd gnd cell_6t
Xbit_r86_c102 bl[102] br[102] wl[86] vdd gnd cell_6t
Xbit_r87_c102 bl[102] br[102] wl[87] vdd gnd cell_6t
Xbit_r88_c102 bl[102] br[102] wl[88] vdd gnd cell_6t
Xbit_r89_c102 bl[102] br[102] wl[89] vdd gnd cell_6t
Xbit_r90_c102 bl[102] br[102] wl[90] vdd gnd cell_6t
Xbit_r91_c102 bl[102] br[102] wl[91] vdd gnd cell_6t
Xbit_r92_c102 bl[102] br[102] wl[92] vdd gnd cell_6t
Xbit_r93_c102 bl[102] br[102] wl[93] vdd gnd cell_6t
Xbit_r94_c102 bl[102] br[102] wl[94] vdd gnd cell_6t
Xbit_r95_c102 bl[102] br[102] wl[95] vdd gnd cell_6t
Xbit_r96_c102 bl[102] br[102] wl[96] vdd gnd cell_6t
Xbit_r97_c102 bl[102] br[102] wl[97] vdd gnd cell_6t
Xbit_r98_c102 bl[102] br[102] wl[98] vdd gnd cell_6t
Xbit_r99_c102 bl[102] br[102] wl[99] vdd gnd cell_6t
Xbit_r100_c102 bl[102] br[102] wl[100] vdd gnd cell_6t
Xbit_r101_c102 bl[102] br[102] wl[101] vdd gnd cell_6t
Xbit_r102_c102 bl[102] br[102] wl[102] vdd gnd cell_6t
Xbit_r103_c102 bl[102] br[102] wl[103] vdd gnd cell_6t
Xbit_r104_c102 bl[102] br[102] wl[104] vdd gnd cell_6t
Xbit_r105_c102 bl[102] br[102] wl[105] vdd gnd cell_6t
Xbit_r106_c102 bl[102] br[102] wl[106] vdd gnd cell_6t
Xbit_r107_c102 bl[102] br[102] wl[107] vdd gnd cell_6t
Xbit_r108_c102 bl[102] br[102] wl[108] vdd gnd cell_6t
Xbit_r109_c102 bl[102] br[102] wl[109] vdd gnd cell_6t
Xbit_r110_c102 bl[102] br[102] wl[110] vdd gnd cell_6t
Xbit_r111_c102 bl[102] br[102] wl[111] vdd gnd cell_6t
Xbit_r112_c102 bl[102] br[102] wl[112] vdd gnd cell_6t
Xbit_r113_c102 bl[102] br[102] wl[113] vdd gnd cell_6t
Xbit_r114_c102 bl[102] br[102] wl[114] vdd gnd cell_6t
Xbit_r115_c102 bl[102] br[102] wl[115] vdd gnd cell_6t
Xbit_r116_c102 bl[102] br[102] wl[116] vdd gnd cell_6t
Xbit_r117_c102 bl[102] br[102] wl[117] vdd gnd cell_6t
Xbit_r118_c102 bl[102] br[102] wl[118] vdd gnd cell_6t
Xbit_r119_c102 bl[102] br[102] wl[119] vdd gnd cell_6t
Xbit_r120_c102 bl[102] br[102] wl[120] vdd gnd cell_6t
Xbit_r121_c102 bl[102] br[102] wl[121] vdd gnd cell_6t
Xbit_r122_c102 bl[102] br[102] wl[122] vdd gnd cell_6t
Xbit_r123_c102 bl[102] br[102] wl[123] vdd gnd cell_6t
Xbit_r124_c102 bl[102] br[102] wl[124] vdd gnd cell_6t
Xbit_r125_c102 bl[102] br[102] wl[125] vdd gnd cell_6t
Xbit_r126_c102 bl[102] br[102] wl[126] vdd gnd cell_6t
Xbit_r127_c102 bl[102] br[102] wl[127] vdd gnd cell_6t
Xbit_r0_c103 bl[103] br[103] wl[0] vdd gnd cell_6t
Xbit_r1_c103 bl[103] br[103] wl[1] vdd gnd cell_6t
Xbit_r2_c103 bl[103] br[103] wl[2] vdd gnd cell_6t
Xbit_r3_c103 bl[103] br[103] wl[3] vdd gnd cell_6t
Xbit_r4_c103 bl[103] br[103] wl[4] vdd gnd cell_6t
Xbit_r5_c103 bl[103] br[103] wl[5] vdd gnd cell_6t
Xbit_r6_c103 bl[103] br[103] wl[6] vdd gnd cell_6t
Xbit_r7_c103 bl[103] br[103] wl[7] vdd gnd cell_6t
Xbit_r8_c103 bl[103] br[103] wl[8] vdd gnd cell_6t
Xbit_r9_c103 bl[103] br[103] wl[9] vdd gnd cell_6t
Xbit_r10_c103 bl[103] br[103] wl[10] vdd gnd cell_6t
Xbit_r11_c103 bl[103] br[103] wl[11] vdd gnd cell_6t
Xbit_r12_c103 bl[103] br[103] wl[12] vdd gnd cell_6t
Xbit_r13_c103 bl[103] br[103] wl[13] vdd gnd cell_6t
Xbit_r14_c103 bl[103] br[103] wl[14] vdd gnd cell_6t
Xbit_r15_c103 bl[103] br[103] wl[15] vdd gnd cell_6t
Xbit_r16_c103 bl[103] br[103] wl[16] vdd gnd cell_6t
Xbit_r17_c103 bl[103] br[103] wl[17] vdd gnd cell_6t
Xbit_r18_c103 bl[103] br[103] wl[18] vdd gnd cell_6t
Xbit_r19_c103 bl[103] br[103] wl[19] vdd gnd cell_6t
Xbit_r20_c103 bl[103] br[103] wl[20] vdd gnd cell_6t
Xbit_r21_c103 bl[103] br[103] wl[21] vdd gnd cell_6t
Xbit_r22_c103 bl[103] br[103] wl[22] vdd gnd cell_6t
Xbit_r23_c103 bl[103] br[103] wl[23] vdd gnd cell_6t
Xbit_r24_c103 bl[103] br[103] wl[24] vdd gnd cell_6t
Xbit_r25_c103 bl[103] br[103] wl[25] vdd gnd cell_6t
Xbit_r26_c103 bl[103] br[103] wl[26] vdd gnd cell_6t
Xbit_r27_c103 bl[103] br[103] wl[27] vdd gnd cell_6t
Xbit_r28_c103 bl[103] br[103] wl[28] vdd gnd cell_6t
Xbit_r29_c103 bl[103] br[103] wl[29] vdd gnd cell_6t
Xbit_r30_c103 bl[103] br[103] wl[30] vdd gnd cell_6t
Xbit_r31_c103 bl[103] br[103] wl[31] vdd gnd cell_6t
Xbit_r32_c103 bl[103] br[103] wl[32] vdd gnd cell_6t
Xbit_r33_c103 bl[103] br[103] wl[33] vdd gnd cell_6t
Xbit_r34_c103 bl[103] br[103] wl[34] vdd gnd cell_6t
Xbit_r35_c103 bl[103] br[103] wl[35] vdd gnd cell_6t
Xbit_r36_c103 bl[103] br[103] wl[36] vdd gnd cell_6t
Xbit_r37_c103 bl[103] br[103] wl[37] vdd gnd cell_6t
Xbit_r38_c103 bl[103] br[103] wl[38] vdd gnd cell_6t
Xbit_r39_c103 bl[103] br[103] wl[39] vdd gnd cell_6t
Xbit_r40_c103 bl[103] br[103] wl[40] vdd gnd cell_6t
Xbit_r41_c103 bl[103] br[103] wl[41] vdd gnd cell_6t
Xbit_r42_c103 bl[103] br[103] wl[42] vdd gnd cell_6t
Xbit_r43_c103 bl[103] br[103] wl[43] vdd gnd cell_6t
Xbit_r44_c103 bl[103] br[103] wl[44] vdd gnd cell_6t
Xbit_r45_c103 bl[103] br[103] wl[45] vdd gnd cell_6t
Xbit_r46_c103 bl[103] br[103] wl[46] vdd gnd cell_6t
Xbit_r47_c103 bl[103] br[103] wl[47] vdd gnd cell_6t
Xbit_r48_c103 bl[103] br[103] wl[48] vdd gnd cell_6t
Xbit_r49_c103 bl[103] br[103] wl[49] vdd gnd cell_6t
Xbit_r50_c103 bl[103] br[103] wl[50] vdd gnd cell_6t
Xbit_r51_c103 bl[103] br[103] wl[51] vdd gnd cell_6t
Xbit_r52_c103 bl[103] br[103] wl[52] vdd gnd cell_6t
Xbit_r53_c103 bl[103] br[103] wl[53] vdd gnd cell_6t
Xbit_r54_c103 bl[103] br[103] wl[54] vdd gnd cell_6t
Xbit_r55_c103 bl[103] br[103] wl[55] vdd gnd cell_6t
Xbit_r56_c103 bl[103] br[103] wl[56] vdd gnd cell_6t
Xbit_r57_c103 bl[103] br[103] wl[57] vdd gnd cell_6t
Xbit_r58_c103 bl[103] br[103] wl[58] vdd gnd cell_6t
Xbit_r59_c103 bl[103] br[103] wl[59] vdd gnd cell_6t
Xbit_r60_c103 bl[103] br[103] wl[60] vdd gnd cell_6t
Xbit_r61_c103 bl[103] br[103] wl[61] vdd gnd cell_6t
Xbit_r62_c103 bl[103] br[103] wl[62] vdd gnd cell_6t
Xbit_r63_c103 bl[103] br[103] wl[63] vdd gnd cell_6t
Xbit_r64_c103 bl[103] br[103] wl[64] vdd gnd cell_6t
Xbit_r65_c103 bl[103] br[103] wl[65] vdd gnd cell_6t
Xbit_r66_c103 bl[103] br[103] wl[66] vdd gnd cell_6t
Xbit_r67_c103 bl[103] br[103] wl[67] vdd gnd cell_6t
Xbit_r68_c103 bl[103] br[103] wl[68] vdd gnd cell_6t
Xbit_r69_c103 bl[103] br[103] wl[69] vdd gnd cell_6t
Xbit_r70_c103 bl[103] br[103] wl[70] vdd gnd cell_6t
Xbit_r71_c103 bl[103] br[103] wl[71] vdd gnd cell_6t
Xbit_r72_c103 bl[103] br[103] wl[72] vdd gnd cell_6t
Xbit_r73_c103 bl[103] br[103] wl[73] vdd gnd cell_6t
Xbit_r74_c103 bl[103] br[103] wl[74] vdd gnd cell_6t
Xbit_r75_c103 bl[103] br[103] wl[75] vdd gnd cell_6t
Xbit_r76_c103 bl[103] br[103] wl[76] vdd gnd cell_6t
Xbit_r77_c103 bl[103] br[103] wl[77] vdd gnd cell_6t
Xbit_r78_c103 bl[103] br[103] wl[78] vdd gnd cell_6t
Xbit_r79_c103 bl[103] br[103] wl[79] vdd gnd cell_6t
Xbit_r80_c103 bl[103] br[103] wl[80] vdd gnd cell_6t
Xbit_r81_c103 bl[103] br[103] wl[81] vdd gnd cell_6t
Xbit_r82_c103 bl[103] br[103] wl[82] vdd gnd cell_6t
Xbit_r83_c103 bl[103] br[103] wl[83] vdd gnd cell_6t
Xbit_r84_c103 bl[103] br[103] wl[84] vdd gnd cell_6t
Xbit_r85_c103 bl[103] br[103] wl[85] vdd gnd cell_6t
Xbit_r86_c103 bl[103] br[103] wl[86] vdd gnd cell_6t
Xbit_r87_c103 bl[103] br[103] wl[87] vdd gnd cell_6t
Xbit_r88_c103 bl[103] br[103] wl[88] vdd gnd cell_6t
Xbit_r89_c103 bl[103] br[103] wl[89] vdd gnd cell_6t
Xbit_r90_c103 bl[103] br[103] wl[90] vdd gnd cell_6t
Xbit_r91_c103 bl[103] br[103] wl[91] vdd gnd cell_6t
Xbit_r92_c103 bl[103] br[103] wl[92] vdd gnd cell_6t
Xbit_r93_c103 bl[103] br[103] wl[93] vdd gnd cell_6t
Xbit_r94_c103 bl[103] br[103] wl[94] vdd gnd cell_6t
Xbit_r95_c103 bl[103] br[103] wl[95] vdd gnd cell_6t
Xbit_r96_c103 bl[103] br[103] wl[96] vdd gnd cell_6t
Xbit_r97_c103 bl[103] br[103] wl[97] vdd gnd cell_6t
Xbit_r98_c103 bl[103] br[103] wl[98] vdd gnd cell_6t
Xbit_r99_c103 bl[103] br[103] wl[99] vdd gnd cell_6t
Xbit_r100_c103 bl[103] br[103] wl[100] vdd gnd cell_6t
Xbit_r101_c103 bl[103] br[103] wl[101] vdd gnd cell_6t
Xbit_r102_c103 bl[103] br[103] wl[102] vdd gnd cell_6t
Xbit_r103_c103 bl[103] br[103] wl[103] vdd gnd cell_6t
Xbit_r104_c103 bl[103] br[103] wl[104] vdd gnd cell_6t
Xbit_r105_c103 bl[103] br[103] wl[105] vdd gnd cell_6t
Xbit_r106_c103 bl[103] br[103] wl[106] vdd gnd cell_6t
Xbit_r107_c103 bl[103] br[103] wl[107] vdd gnd cell_6t
Xbit_r108_c103 bl[103] br[103] wl[108] vdd gnd cell_6t
Xbit_r109_c103 bl[103] br[103] wl[109] vdd gnd cell_6t
Xbit_r110_c103 bl[103] br[103] wl[110] vdd gnd cell_6t
Xbit_r111_c103 bl[103] br[103] wl[111] vdd gnd cell_6t
Xbit_r112_c103 bl[103] br[103] wl[112] vdd gnd cell_6t
Xbit_r113_c103 bl[103] br[103] wl[113] vdd gnd cell_6t
Xbit_r114_c103 bl[103] br[103] wl[114] vdd gnd cell_6t
Xbit_r115_c103 bl[103] br[103] wl[115] vdd gnd cell_6t
Xbit_r116_c103 bl[103] br[103] wl[116] vdd gnd cell_6t
Xbit_r117_c103 bl[103] br[103] wl[117] vdd gnd cell_6t
Xbit_r118_c103 bl[103] br[103] wl[118] vdd gnd cell_6t
Xbit_r119_c103 bl[103] br[103] wl[119] vdd gnd cell_6t
Xbit_r120_c103 bl[103] br[103] wl[120] vdd gnd cell_6t
Xbit_r121_c103 bl[103] br[103] wl[121] vdd gnd cell_6t
Xbit_r122_c103 bl[103] br[103] wl[122] vdd gnd cell_6t
Xbit_r123_c103 bl[103] br[103] wl[123] vdd gnd cell_6t
Xbit_r124_c103 bl[103] br[103] wl[124] vdd gnd cell_6t
Xbit_r125_c103 bl[103] br[103] wl[125] vdd gnd cell_6t
Xbit_r126_c103 bl[103] br[103] wl[126] vdd gnd cell_6t
Xbit_r127_c103 bl[103] br[103] wl[127] vdd gnd cell_6t
Xbit_r0_c104 bl[104] br[104] wl[0] vdd gnd cell_6t
Xbit_r1_c104 bl[104] br[104] wl[1] vdd gnd cell_6t
Xbit_r2_c104 bl[104] br[104] wl[2] vdd gnd cell_6t
Xbit_r3_c104 bl[104] br[104] wl[3] vdd gnd cell_6t
Xbit_r4_c104 bl[104] br[104] wl[4] vdd gnd cell_6t
Xbit_r5_c104 bl[104] br[104] wl[5] vdd gnd cell_6t
Xbit_r6_c104 bl[104] br[104] wl[6] vdd gnd cell_6t
Xbit_r7_c104 bl[104] br[104] wl[7] vdd gnd cell_6t
Xbit_r8_c104 bl[104] br[104] wl[8] vdd gnd cell_6t
Xbit_r9_c104 bl[104] br[104] wl[9] vdd gnd cell_6t
Xbit_r10_c104 bl[104] br[104] wl[10] vdd gnd cell_6t
Xbit_r11_c104 bl[104] br[104] wl[11] vdd gnd cell_6t
Xbit_r12_c104 bl[104] br[104] wl[12] vdd gnd cell_6t
Xbit_r13_c104 bl[104] br[104] wl[13] vdd gnd cell_6t
Xbit_r14_c104 bl[104] br[104] wl[14] vdd gnd cell_6t
Xbit_r15_c104 bl[104] br[104] wl[15] vdd gnd cell_6t
Xbit_r16_c104 bl[104] br[104] wl[16] vdd gnd cell_6t
Xbit_r17_c104 bl[104] br[104] wl[17] vdd gnd cell_6t
Xbit_r18_c104 bl[104] br[104] wl[18] vdd gnd cell_6t
Xbit_r19_c104 bl[104] br[104] wl[19] vdd gnd cell_6t
Xbit_r20_c104 bl[104] br[104] wl[20] vdd gnd cell_6t
Xbit_r21_c104 bl[104] br[104] wl[21] vdd gnd cell_6t
Xbit_r22_c104 bl[104] br[104] wl[22] vdd gnd cell_6t
Xbit_r23_c104 bl[104] br[104] wl[23] vdd gnd cell_6t
Xbit_r24_c104 bl[104] br[104] wl[24] vdd gnd cell_6t
Xbit_r25_c104 bl[104] br[104] wl[25] vdd gnd cell_6t
Xbit_r26_c104 bl[104] br[104] wl[26] vdd gnd cell_6t
Xbit_r27_c104 bl[104] br[104] wl[27] vdd gnd cell_6t
Xbit_r28_c104 bl[104] br[104] wl[28] vdd gnd cell_6t
Xbit_r29_c104 bl[104] br[104] wl[29] vdd gnd cell_6t
Xbit_r30_c104 bl[104] br[104] wl[30] vdd gnd cell_6t
Xbit_r31_c104 bl[104] br[104] wl[31] vdd gnd cell_6t
Xbit_r32_c104 bl[104] br[104] wl[32] vdd gnd cell_6t
Xbit_r33_c104 bl[104] br[104] wl[33] vdd gnd cell_6t
Xbit_r34_c104 bl[104] br[104] wl[34] vdd gnd cell_6t
Xbit_r35_c104 bl[104] br[104] wl[35] vdd gnd cell_6t
Xbit_r36_c104 bl[104] br[104] wl[36] vdd gnd cell_6t
Xbit_r37_c104 bl[104] br[104] wl[37] vdd gnd cell_6t
Xbit_r38_c104 bl[104] br[104] wl[38] vdd gnd cell_6t
Xbit_r39_c104 bl[104] br[104] wl[39] vdd gnd cell_6t
Xbit_r40_c104 bl[104] br[104] wl[40] vdd gnd cell_6t
Xbit_r41_c104 bl[104] br[104] wl[41] vdd gnd cell_6t
Xbit_r42_c104 bl[104] br[104] wl[42] vdd gnd cell_6t
Xbit_r43_c104 bl[104] br[104] wl[43] vdd gnd cell_6t
Xbit_r44_c104 bl[104] br[104] wl[44] vdd gnd cell_6t
Xbit_r45_c104 bl[104] br[104] wl[45] vdd gnd cell_6t
Xbit_r46_c104 bl[104] br[104] wl[46] vdd gnd cell_6t
Xbit_r47_c104 bl[104] br[104] wl[47] vdd gnd cell_6t
Xbit_r48_c104 bl[104] br[104] wl[48] vdd gnd cell_6t
Xbit_r49_c104 bl[104] br[104] wl[49] vdd gnd cell_6t
Xbit_r50_c104 bl[104] br[104] wl[50] vdd gnd cell_6t
Xbit_r51_c104 bl[104] br[104] wl[51] vdd gnd cell_6t
Xbit_r52_c104 bl[104] br[104] wl[52] vdd gnd cell_6t
Xbit_r53_c104 bl[104] br[104] wl[53] vdd gnd cell_6t
Xbit_r54_c104 bl[104] br[104] wl[54] vdd gnd cell_6t
Xbit_r55_c104 bl[104] br[104] wl[55] vdd gnd cell_6t
Xbit_r56_c104 bl[104] br[104] wl[56] vdd gnd cell_6t
Xbit_r57_c104 bl[104] br[104] wl[57] vdd gnd cell_6t
Xbit_r58_c104 bl[104] br[104] wl[58] vdd gnd cell_6t
Xbit_r59_c104 bl[104] br[104] wl[59] vdd gnd cell_6t
Xbit_r60_c104 bl[104] br[104] wl[60] vdd gnd cell_6t
Xbit_r61_c104 bl[104] br[104] wl[61] vdd gnd cell_6t
Xbit_r62_c104 bl[104] br[104] wl[62] vdd gnd cell_6t
Xbit_r63_c104 bl[104] br[104] wl[63] vdd gnd cell_6t
Xbit_r64_c104 bl[104] br[104] wl[64] vdd gnd cell_6t
Xbit_r65_c104 bl[104] br[104] wl[65] vdd gnd cell_6t
Xbit_r66_c104 bl[104] br[104] wl[66] vdd gnd cell_6t
Xbit_r67_c104 bl[104] br[104] wl[67] vdd gnd cell_6t
Xbit_r68_c104 bl[104] br[104] wl[68] vdd gnd cell_6t
Xbit_r69_c104 bl[104] br[104] wl[69] vdd gnd cell_6t
Xbit_r70_c104 bl[104] br[104] wl[70] vdd gnd cell_6t
Xbit_r71_c104 bl[104] br[104] wl[71] vdd gnd cell_6t
Xbit_r72_c104 bl[104] br[104] wl[72] vdd gnd cell_6t
Xbit_r73_c104 bl[104] br[104] wl[73] vdd gnd cell_6t
Xbit_r74_c104 bl[104] br[104] wl[74] vdd gnd cell_6t
Xbit_r75_c104 bl[104] br[104] wl[75] vdd gnd cell_6t
Xbit_r76_c104 bl[104] br[104] wl[76] vdd gnd cell_6t
Xbit_r77_c104 bl[104] br[104] wl[77] vdd gnd cell_6t
Xbit_r78_c104 bl[104] br[104] wl[78] vdd gnd cell_6t
Xbit_r79_c104 bl[104] br[104] wl[79] vdd gnd cell_6t
Xbit_r80_c104 bl[104] br[104] wl[80] vdd gnd cell_6t
Xbit_r81_c104 bl[104] br[104] wl[81] vdd gnd cell_6t
Xbit_r82_c104 bl[104] br[104] wl[82] vdd gnd cell_6t
Xbit_r83_c104 bl[104] br[104] wl[83] vdd gnd cell_6t
Xbit_r84_c104 bl[104] br[104] wl[84] vdd gnd cell_6t
Xbit_r85_c104 bl[104] br[104] wl[85] vdd gnd cell_6t
Xbit_r86_c104 bl[104] br[104] wl[86] vdd gnd cell_6t
Xbit_r87_c104 bl[104] br[104] wl[87] vdd gnd cell_6t
Xbit_r88_c104 bl[104] br[104] wl[88] vdd gnd cell_6t
Xbit_r89_c104 bl[104] br[104] wl[89] vdd gnd cell_6t
Xbit_r90_c104 bl[104] br[104] wl[90] vdd gnd cell_6t
Xbit_r91_c104 bl[104] br[104] wl[91] vdd gnd cell_6t
Xbit_r92_c104 bl[104] br[104] wl[92] vdd gnd cell_6t
Xbit_r93_c104 bl[104] br[104] wl[93] vdd gnd cell_6t
Xbit_r94_c104 bl[104] br[104] wl[94] vdd gnd cell_6t
Xbit_r95_c104 bl[104] br[104] wl[95] vdd gnd cell_6t
Xbit_r96_c104 bl[104] br[104] wl[96] vdd gnd cell_6t
Xbit_r97_c104 bl[104] br[104] wl[97] vdd gnd cell_6t
Xbit_r98_c104 bl[104] br[104] wl[98] vdd gnd cell_6t
Xbit_r99_c104 bl[104] br[104] wl[99] vdd gnd cell_6t
Xbit_r100_c104 bl[104] br[104] wl[100] vdd gnd cell_6t
Xbit_r101_c104 bl[104] br[104] wl[101] vdd gnd cell_6t
Xbit_r102_c104 bl[104] br[104] wl[102] vdd gnd cell_6t
Xbit_r103_c104 bl[104] br[104] wl[103] vdd gnd cell_6t
Xbit_r104_c104 bl[104] br[104] wl[104] vdd gnd cell_6t
Xbit_r105_c104 bl[104] br[104] wl[105] vdd gnd cell_6t
Xbit_r106_c104 bl[104] br[104] wl[106] vdd gnd cell_6t
Xbit_r107_c104 bl[104] br[104] wl[107] vdd gnd cell_6t
Xbit_r108_c104 bl[104] br[104] wl[108] vdd gnd cell_6t
Xbit_r109_c104 bl[104] br[104] wl[109] vdd gnd cell_6t
Xbit_r110_c104 bl[104] br[104] wl[110] vdd gnd cell_6t
Xbit_r111_c104 bl[104] br[104] wl[111] vdd gnd cell_6t
Xbit_r112_c104 bl[104] br[104] wl[112] vdd gnd cell_6t
Xbit_r113_c104 bl[104] br[104] wl[113] vdd gnd cell_6t
Xbit_r114_c104 bl[104] br[104] wl[114] vdd gnd cell_6t
Xbit_r115_c104 bl[104] br[104] wl[115] vdd gnd cell_6t
Xbit_r116_c104 bl[104] br[104] wl[116] vdd gnd cell_6t
Xbit_r117_c104 bl[104] br[104] wl[117] vdd gnd cell_6t
Xbit_r118_c104 bl[104] br[104] wl[118] vdd gnd cell_6t
Xbit_r119_c104 bl[104] br[104] wl[119] vdd gnd cell_6t
Xbit_r120_c104 bl[104] br[104] wl[120] vdd gnd cell_6t
Xbit_r121_c104 bl[104] br[104] wl[121] vdd gnd cell_6t
Xbit_r122_c104 bl[104] br[104] wl[122] vdd gnd cell_6t
Xbit_r123_c104 bl[104] br[104] wl[123] vdd gnd cell_6t
Xbit_r124_c104 bl[104] br[104] wl[124] vdd gnd cell_6t
Xbit_r125_c104 bl[104] br[104] wl[125] vdd gnd cell_6t
Xbit_r126_c104 bl[104] br[104] wl[126] vdd gnd cell_6t
Xbit_r127_c104 bl[104] br[104] wl[127] vdd gnd cell_6t
Xbit_r0_c105 bl[105] br[105] wl[0] vdd gnd cell_6t
Xbit_r1_c105 bl[105] br[105] wl[1] vdd gnd cell_6t
Xbit_r2_c105 bl[105] br[105] wl[2] vdd gnd cell_6t
Xbit_r3_c105 bl[105] br[105] wl[3] vdd gnd cell_6t
Xbit_r4_c105 bl[105] br[105] wl[4] vdd gnd cell_6t
Xbit_r5_c105 bl[105] br[105] wl[5] vdd gnd cell_6t
Xbit_r6_c105 bl[105] br[105] wl[6] vdd gnd cell_6t
Xbit_r7_c105 bl[105] br[105] wl[7] vdd gnd cell_6t
Xbit_r8_c105 bl[105] br[105] wl[8] vdd gnd cell_6t
Xbit_r9_c105 bl[105] br[105] wl[9] vdd gnd cell_6t
Xbit_r10_c105 bl[105] br[105] wl[10] vdd gnd cell_6t
Xbit_r11_c105 bl[105] br[105] wl[11] vdd gnd cell_6t
Xbit_r12_c105 bl[105] br[105] wl[12] vdd gnd cell_6t
Xbit_r13_c105 bl[105] br[105] wl[13] vdd gnd cell_6t
Xbit_r14_c105 bl[105] br[105] wl[14] vdd gnd cell_6t
Xbit_r15_c105 bl[105] br[105] wl[15] vdd gnd cell_6t
Xbit_r16_c105 bl[105] br[105] wl[16] vdd gnd cell_6t
Xbit_r17_c105 bl[105] br[105] wl[17] vdd gnd cell_6t
Xbit_r18_c105 bl[105] br[105] wl[18] vdd gnd cell_6t
Xbit_r19_c105 bl[105] br[105] wl[19] vdd gnd cell_6t
Xbit_r20_c105 bl[105] br[105] wl[20] vdd gnd cell_6t
Xbit_r21_c105 bl[105] br[105] wl[21] vdd gnd cell_6t
Xbit_r22_c105 bl[105] br[105] wl[22] vdd gnd cell_6t
Xbit_r23_c105 bl[105] br[105] wl[23] vdd gnd cell_6t
Xbit_r24_c105 bl[105] br[105] wl[24] vdd gnd cell_6t
Xbit_r25_c105 bl[105] br[105] wl[25] vdd gnd cell_6t
Xbit_r26_c105 bl[105] br[105] wl[26] vdd gnd cell_6t
Xbit_r27_c105 bl[105] br[105] wl[27] vdd gnd cell_6t
Xbit_r28_c105 bl[105] br[105] wl[28] vdd gnd cell_6t
Xbit_r29_c105 bl[105] br[105] wl[29] vdd gnd cell_6t
Xbit_r30_c105 bl[105] br[105] wl[30] vdd gnd cell_6t
Xbit_r31_c105 bl[105] br[105] wl[31] vdd gnd cell_6t
Xbit_r32_c105 bl[105] br[105] wl[32] vdd gnd cell_6t
Xbit_r33_c105 bl[105] br[105] wl[33] vdd gnd cell_6t
Xbit_r34_c105 bl[105] br[105] wl[34] vdd gnd cell_6t
Xbit_r35_c105 bl[105] br[105] wl[35] vdd gnd cell_6t
Xbit_r36_c105 bl[105] br[105] wl[36] vdd gnd cell_6t
Xbit_r37_c105 bl[105] br[105] wl[37] vdd gnd cell_6t
Xbit_r38_c105 bl[105] br[105] wl[38] vdd gnd cell_6t
Xbit_r39_c105 bl[105] br[105] wl[39] vdd gnd cell_6t
Xbit_r40_c105 bl[105] br[105] wl[40] vdd gnd cell_6t
Xbit_r41_c105 bl[105] br[105] wl[41] vdd gnd cell_6t
Xbit_r42_c105 bl[105] br[105] wl[42] vdd gnd cell_6t
Xbit_r43_c105 bl[105] br[105] wl[43] vdd gnd cell_6t
Xbit_r44_c105 bl[105] br[105] wl[44] vdd gnd cell_6t
Xbit_r45_c105 bl[105] br[105] wl[45] vdd gnd cell_6t
Xbit_r46_c105 bl[105] br[105] wl[46] vdd gnd cell_6t
Xbit_r47_c105 bl[105] br[105] wl[47] vdd gnd cell_6t
Xbit_r48_c105 bl[105] br[105] wl[48] vdd gnd cell_6t
Xbit_r49_c105 bl[105] br[105] wl[49] vdd gnd cell_6t
Xbit_r50_c105 bl[105] br[105] wl[50] vdd gnd cell_6t
Xbit_r51_c105 bl[105] br[105] wl[51] vdd gnd cell_6t
Xbit_r52_c105 bl[105] br[105] wl[52] vdd gnd cell_6t
Xbit_r53_c105 bl[105] br[105] wl[53] vdd gnd cell_6t
Xbit_r54_c105 bl[105] br[105] wl[54] vdd gnd cell_6t
Xbit_r55_c105 bl[105] br[105] wl[55] vdd gnd cell_6t
Xbit_r56_c105 bl[105] br[105] wl[56] vdd gnd cell_6t
Xbit_r57_c105 bl[105] br[105] wl[57] vdd gnd cell_6t
Xbit_r58_c105 bl[105] br[105] wl[58] vdd gnd cell_6t
Xbit_r59_c105 bl[105] br[105] wl[59] vdd gnd cell_6t
Xbit_r60_c105 bl[105] br[105] wl[60] vdd gnd cell_6t
Xbit_r61_c105 bl[105] br[105] wl[61] vdd gnd cell_6t
Xbit_r62_c105 bl[105] br[105] wl[62] vdd gnd cell_6t
Xbit_r63_c105 bl[105] br[105] wl[63] vdd gnd cell_6t
Xbit_r64_c105 bl[105] br[105] wl[64] vdd gnd cell_6t
Xbit_r65_c105 bl[105] br[105] wl[65] vdd gnd cell_6t
Xbit_r66_c105 bl[105] br[105] wl[66] vdd gnd cell_6t
Xbit_r67_c105 bl[105] br[105] wl[67] vdd gnd cell_6t
Xbit_r68_c105 bl[105] br[105] wl[68] vdd gnd cell_6t
Xbit_r69_c105 bl[105] br[105] wl[69] vdd gnd cell_6t
Xbit_r70_c105 bl[105] br[105] wl[70] vdd gnd cell_6t
Xbit_r71_c105 bl[105] br[105] wl[71] vdd gnd cell_6t
Xbit_r72_c105 bl[105] br[105] wl[72] vdd gnd cell_6t
Xbit_r73_c105 bl[105] br[105] wl[73] vdd gnd cell_6t
Xbit_r74_c105 bl[105] br[105] wl[74] vdd gnd cell_6t
Xbit_r75_c105 bl[105] br[105] wl[75] vdd gnd cell_6t
Xbit_r76_c105 bl[105] br[105] wl[76] vdd gnd cell_6t
Xbit_r77_c105 bl[105] br[105] wl[77] vdd gnd cell_6t
Xbit_r78_c105 bl[105] br[105] wl[78] vdd gnd cell_6t
Xbit_r79_c105 bl[105] br[105] wl[79] vdd gnd cell_6t
Xbit_r80_c105 bl[105] br[105] wl[80] vdd gnd cell_6t
Xbit_r81_c105 bl[105] br[105] wl[81] vdd gnd cell_6t
Xbit_r82_c105 bl[105] br[105] wl[82] vdd gnd cell_6t
Xbit_r83_c105 bl[105] br[105] wl[83] vdd gnd cell_6t
Xbit_r84_c105 bl[105] br[105] wl[84] vdd gnd cell_6t
Xbit_r85_c105 bl[105] br[105] wl[85] vdd gnd cell_6t
Xbit_r86_c105 bl[105] br[105] wl[86] vdd gnd cell_6t
Xbit_r87_c105 bl[105] br[105] wl[87] vdd gnd cell_6t
Xbit_r88_c105 bl[105] br[105] wl[88] vdd gnd cell_6t
Xbit_r89_c105 bl[105] br[105] wl[89] vdd gnd cell_6t
Xbit_r90_c105 bl[105] br[105] wl[90] vdd gnd cell_6t
Xbit_r91_c105 bl[105] br[105] wl[91] vdd gnd cell_6t
Xbit_r92_c105 bl[105] br[105] wl[92] vdd gnd cell_6t
Xbit_r93_c105 bl[105] br[105] wl[93] vdd gnd cell_6t
Xbit_r94_c105 bl[105] br[105] wl[94] vdd gnd cell_6t
Xbit_r95_c105 bl[105] br[105] wl[95] vdd gnd cell_6t
Xbit_r96_c105 bl[105] br[105] wl[96] vdd gnd cell_6t
Xbit_r97_c105 bl[105] br[105] wl[97] vdd gnd cell_6t
Xbit_r98_c105 bl[105] br[105] wl[98] vdd gnd cell_6t
Xbit_r99_c105 bl[105] br[105] wl[99] vdd gnd cell_6t
Xbit_r100_c105 bl[105] br[105] wl[100] vdd gnd cell_6t
Xbit_r101_c105 bl[105] br[105] wl[101] vdd gnd cell_6t
Xbit_r102_c105 bl[105] br[105] wl[102] vdd gnd cell_6t
Xbit_r103_c105 bl[105] br[105] wl[103] vdd gnd cell_6t
Xbit_r104_c105 bl[105] br[105] wl[104] vdd gnd cell_6t
Xbit_r105_c105 bl[105] br[105] wl[105] vdd gnd cell_6t
Xbit_r106_c105 bl[105] br[105] wl[106] vdd gnd cell_6t
Xbit_r107_c105 bl[105] br[105] wl[107] vdd gnd cell_6t
Xbit_r108_c105 bl[105] br[105] wl[108] vdd gnd cell_6t
Xbit_r109_c105 bl[105] br[105] wl[109] vdd gnd cell_6t
Xbit_r110_c105 bl[105] br[105] wl[110] vdd gnd cell_6t
Xbit_r111_c105 bl[105] br[105] wl[111] vdd gnd cell_6t
Xbit_r112_c105 bl[105] br[105] wl[112] vdd gnd cell_6t
Xbit_r113_c105 bl[105] br[105] wl[113] vdd gnd cell_6t
Xbit_r114_c105 bl[105] br[105] wl[114] vdd gnd cell_6t
Xbit_r115_c105 bl[105] br[105] wl[115] vdd gnd cell_6t
Xbit_r116_c105 bl[105] br[105] wl[116] vdd gnd cell_6t
Xbit_r117_c105 bl[105] br[105] wl[117] vdd gnd cell_6t
Xbit_r118_c105 bl[105] br[105] wl[118] vdd gnd cell_6t
Xbit_r119_c105 bl[105] br[105] wl[119] vdd gnd cell_6t
Xbit_r120_c105 bl[105] br[105] wl[120] vdd gnd cell_6t
Xbit_r121_c105 bl[105] br[105] wl[121] vdd gnd cell_6t
Xbit_r122_c105 bl[105] br[105] wl[122] vdd gnd cell_6t
Xbit_r123_c105 bl[105] br[105] wl[123] vdd gnd cell_6t
Xbit_r124_c105 bl[105] br[105] wl[124] vdd gnd cell_6t
Xbit_r125_c105 bl[105] br[105] wl[125] vdd gnd cell_6t
Xbit_r126_c105 bl[105] br[105] wl[126] vdd gnd cell_6t
Xbit_r127_c105 bl[105] br[105] wl[127] vdd gnd cell_6t
Xbit_r0_c106 bl[106] br[106] wl[0] vdd gnd cell_6t
Xbit_r1_c106 bl[106] br[106] wl[1] vdd gnd cell_6t
Xbit_r2_c106 bl[106] br[106] wl[2] vdd gnd cell_6t
Xbit_r3_c106 bl[106] br[106] wl[3] vdd gnd cell_6t
Xbit_r4_c106 bl[106] br[106] wl[4] vdd gnd cell_6t
Xbit_r5_c106 bl[106] br[106] wl[5] vdd gnd cell_6t
Xbit_r6_c106 bl[106] br[106] wl[6] vdd gnd cell_6t
Xbit_r7_c106 bl[106] br[106] wl[7] vdd gnd cell_6t
Xbit_r8_c106 bl[106] br[106] wl[8] vdd gnd cell_6t
Xbit_r9_c106 bl[106] br[106] wl[9] vdd gnd cell_6t
Xbit_r10_c106 bl[106] br[106] wl[10] vdd gnd cell_6t
Xbit_r11_c106 bl[106] br[106] wl[11] vdd gnd cell_6t
Xbit_r12_c106 bl[106] br[106] wl[12] vdd gnd cell_6t
Xbit_r13_c106 bl[106] br[106] wl[13] vdd gnd cell_6t
Xbit_r14_c106 bl[106] br[106] wl[14] vdd gnd cell_6t
Xbit_r15_c106 bl[106] br[106] wl[15] vdd gnd cell_6t
Xbit_r16_c106 bl[106] br[106] wl[16] vdd gnd cell_6t
Xbit_r17_c106 bl[106] br[106] wl[17] vdd gnd cell_6t
Xbit_r18_c106 bl[106] br[106] wl[18] vdd gnd cell_6t
Xbit_r19_c106 bl[106] br[106] wl[19] vdd gnd cell_6t
Xbit_r20_c106 bl[106] br[106] wl[20] vdd gnd cell_6t
Xbit_r21_c106 bl[106] br[106] wl[21] vdd gnd cell_6t
Xbit_r22_c106 bl[106] br[106] wl[22] vdd gnd cell_6t
Xbit_r23_c106 bl[106] br[106] wl[23] vdd gnd cell_6t
Xbit_r24_c106 bl[106] br[106] wl[24] vdd gnd cell_6t
Xbit_r25_c106 bl[106] br[106] wl[25] vdd gnd cell_6t
Xbit_r26_c106 bl[106] br[106] wl[26] vdd gnd cell_6t
Xbit_r27_c106 bl[106] br[106] wl[27] vdd gnd cell_6t
Xbit_r28_c106 bl[106] br[106] wl[28] vdd gnd cell_6t
Xbit_r29_c106 bl[106] br[106] wl[29] vdd gnd cell_6t
Xbit_r30_c106 bl[106] br[106] wl[30] vdd gnd cell_6t
Xbit_r31_c106 bl[106] br[106] wl[31] vdd gnd cell_6t
Xbit_r32_c106 bl[106] br[106] wl[32] vdd gnd cell_6t
Xbit_r33_c106 bl[106] br[106] wl[33] vdd gnd cell_6t
Xbit_r34_c106 bl[106] br[106] wl[34] vdd gnd cell_6t
Xbit_r35_c106 bl[106] br[106] wl[35] vdd gnd cell_6t
Xbit_r36_c106 bl[106] br[106] wl[36] vdd gnd cell_6t
Xbit_r37_c106 bl[106] br[106] wl[37] vdd gnd cell_6t
Xbit_r38_c106 bl[106] br[106] wl[38] vdd gnd cell_6t
Xbit_r39_c106 bl[106] br[106] wl[39] vdd gnd cell_6t
Xbit_r40_c106 bl[106] br[106] wl[40] vdd gnd cell_6t
Xbit_r41_c106 bl[106] br[106] wl[41] vdd gnd cell_6t
Xbit_r42_c106 bl[106] br[106] wl[42] vdd gnd cell_6t
Xbit_r43_c106 bl[106] br[106] wl[43] vdd gnd cell_6t
Xbit_r44_c106 bl[106] br[106] wl[44] vdd gnd cell_6t
Xbit_r45_c106 bl[106] br[106] wl[45] vdd gnd cell_6t
Xbit_r46_c106 bl[106] br[106] wl[46] vdd gnd cell_6t
Xbit_r47_c106 bl[106] br[106] wl[47] vdd gnd cell_6t
Xbit_r48_c106 bl[106] br[106] wl[48] vdd gnd cell_6t
Xbit_r49_c106 bl[106] br[106] wl[49] vdd gnd cell_6t
Xbit_r50_c106 bl[106] br[106] wl[50] vdd gnd cell_6t
Xbit_r51_c106 bl[106] br[106] wl[51] vdd gnd cell_6t
Xbit_r52_c106 bl[106] br[106] wl[52] vdd gnd cell_6t
Xbit_r53_c106 bl[106] br[106] wl[53] vdd gnd cell_6t
Xbit_r54_c106 bl[106] br[106] wl[54] vdd gnd cell_6t
Xbit_r55_c106 bl[106] br[106] wl[55] vdd gnd cell_6t
Xbit_r56_c106 bl[106] br[106] wl[56] vdd gnd cell_6t
Xbit_r57_c106 bl[106] br[106] wl[57] vdd gnd cell_6t
Xbit_r58_c106 bl[106] br[106] wl[58] vdd gnd cell_6t
Xbit_r59_c106 bl[106] br[106] wl[59] vdd gnd cell_6t
Xbit_r60_c106 bl[106] br[106] wl[60] vdd gnd cell_6t
Xbit_r61_c106 bl[106] br[106] wl[61] vdd gnd cell_6t
Xbit_r62_c106 bl[106] br[106] wl[62] vdd gnd cell_6t
Xbit_r63_c106 bl[106] br[106] wl[63] vdd gnd cell_6t
Xbit_r64_c106 bl[106] br[106] wl[64] vdd gnd cell_6t
Xbit_r65_c106 bl[106] br[106] wl[65] vdd gnd cell_6t
Xbit_r66_c106 bl[106] br[106] wl[66] vdd gnd cell_6t
Xbit_r67_c106 bl[106] br[106] wl[67] vdd gnd cell_6t
Xbit_r68_c106 bl[106] br[106] wl[68] vdd gnd cell_6t
Xbit_r69_c106 bl[106] br[106] wl[69] vdd gnd cell_6t
Xbit_r70_c106 bl[106] br[106] wl[70] vdd gnd cell_6t
Xbit_r71_c106 bl[106] br[106] wl[71] vdd gnd cell_6t
Xbit_r72_c106 bl[106] br[106] wl[72] vdd gnd cell_6t
Xbit_r73_c106 bl[106] br[106] wl[73] vdd gnd cell_6t
Xbit_r74_c106 bl[106] br[106] wl[74] vdd gnd cell_6t
Xbit_r75_c106 bl[106] br[106] wl[75] vdd gnd cell_6t
Xbit_r76_c106 bl[106] br[106] wl[76] vdd gnd cell_6t
Xbit_r77_c106 bl[106] br[106] wl[77] vdd gnd cell_6t
Xbit_r78_c106 bl[106] br[106] wl[78] vdd gnd cell_6t
Xbit_r79_c106 bl[106] br[106] wl[79] vdd gnd cell_6t
Xbit_r80_c106 bl[106] br[106] wl[80] vdd gnd cell_6t
Xbit_r81_c106 bl[106] br[106] wl[81] vdd gnd cell_6t
Xbit_r82_c106 bl[106] br[106] wl[82] vdd gnd cell_6t
Xbit_r83_c106 bl[106] br[106] wl[83] vdd gnd cell_6t
Xbit_r84_c106 bl[106] br[106] wl[84] vdd gnd cell_6t
Xbit_r85_c106 bl[106] br[106] wl[85] vdd gnd cell_6t
Xbit_r86_c106 bl[106] br[106] wl[86] vdd gnd cell_6t
Xbit_r87_c106 bl[106] br[106] wl[87] vdd gnd cell_6t
Xbit_r88_c106 bl[106] br[106] wl[88] vdd gnd cell_6t
Xbit_r89_c106 bl[106] br[106] wl[89] vdd gnd cell_6t
Xbit_r90_c106 bl[106] br[106] wl[90] vdd gnd cell_6t
Xbit_r91_c106 bl[106] br[106] wl[91] vdd gnd cell_6t
Xbit_r92_c106 bl[106] br[106] wl[92] vdd gnd cell_6t
Xbit_r93_c106 bl[106] br[106] wl[93] vdd gnd cell_6t
Xbit_r94_c106 bl[106] br[106] wl[94] vdd gnd cell_6t
Xbit_r95_c106 bl[106] br[106] wl[95] vdd gnd cell_6t
Xbit_r96_c106 bl[106] br[106] wl[96] vdd gnd cell_6t
Xbit_r97_c106 bl[106] br[106] wl[97] vdd gnd cell_6t
Xbit_r98_c106 bl[106] br[106] wl[98] vdd gnd cell_6t
Xbit_r99_c106 bl[106] br[106] wl[99] vdd gnd cell_6t
Xbit_r100_c106 bl[106] br[106] wl[100] vdd gnd cell_6t
Xbit_r101_c106 bl[106] br[106] wl[101] vdd gnd cell_6t
Xbit_r102_c106 bl[106] br[106] wl[102] vdd gnd cell_6t
Xbit_r103_c106 bl[106] br[106] wl[103] vdd gnd cell_6t
Xbit_r104_c106 bl[106] br[106] wl[104] vdd gnd cell_6t
Xbit_r105_c106 bl[106] br[106] wl[105] vdd gnd cell_6t
Xbit_r106_c106 bl[106] br[106] wl[106] vdd gnd cell_6t
Xbit_r107_c106 bl[106] br[106] wl[107] vdd gnd cell_6t
Xbit_r108_c106 bl[106] br[106] wl[108] vdd gnd cell_6t
Xbit_r109_c106 bl[106] br[106] wl[109] vdd gnd cell_6t
Xbit_r110_c106 bl[106] br[106] wl[110] vdd gnd cell_6t
Xbit_r111_c106 bl[106] br[106] wl[111] vdd gnd cell_6t
Xbit_r112_c106 bl[106] br[106] wl[112] vdd gnd cell_6t
Xbit_r113_c106 bl[106] br[106] wl[113] vdd gnd cell_6t
Xbit_r114_c106 bl[106] br[106] wl[114] vdd gnd cell_6t
Xbit_r115_c106 bl[106] br[106] wl[115] vdd gnd cell_6t
Xbit_r116_c106 bl[106] br[106] wl[116] vdd gnd cell_6t
Xbit_r117_c106 bl[106] br[106] wl[117] vdd gnd cell_6t
Xbit_r118_c106 bl[106] br[106] wl[118] vdd gnd cell_6t
Xbit_r119_c106 bl[106] br[106] wl[119] vdd gnd cell_6t
Xbit_r120_c106 bl[106] br[106] wl[120] vdd gnd cell_6t
Xbit_r121_c106 bl[106] br[106] wl[121] vdd gnd cell_6t
Xbit_r122_c106 bl[106] br[106] wl[122] vdd gnd cell_6t
Xbit_r123_c106 bl[106] br[106] wl[123] vdd gnd cell_6t
Xbit_r124_c106 bl[106] br[106] wl[124] vdd gnd cell_6t
Xbit_r125_c106 bl[106] br[106] wl[125] vdd gnd cell_6t
Xbit_r126_c106 bl[106] br[106] wl[126] vdd gnd cell_6t
Xbit_r127_c106 bl[106] br[106] wl[127] vdd gnd cell_6t
Xbit_r0_c107 bl[107] br[107] wl[0] vdd gnd cell_6t
Xbit_r1_c107 bl[107] br[107] wl[1] vdd gnd cell_6t
Xbit_r2_c107 bl[107] br[107] wl[2] vdd gnd cell_6t
Xbit_r3_c107 bl[107] br[107] wl[3] vdd gnd cell_6t
Xbit_r4_c107 bl[107] br[107] wl[4] vdd gnd cell_6t
Xbit_r5_c107 bl[107] br[107] wl[5] vdd gnd cell_6t
Xbit_r6_c107 bl[107] br[107] wl[6] vdd gnd cell_6t
Xbit_r7_c107 bl[107] br[107] wl[7] vdd gnd cell_6t
Xbit_r8_c107 bl[107] br[107] wl[8] vdd gnd cell_6t
Xbit_r9_c107 bl[107] br[107] wl[9] vdd gnd cell_6t
Xbit_r10_c107 bl[107] br[107] wl[10] vdd gnd cell_6t
Xbit_r11_c107 bl[107] br[107] wl[11] vdd gnd cell_6t
Xbit_r12_c107 bl[107] br[107] wl[12] vdd gnd cell_6t
Xbit_r13_c107 bl[107] br[107] wl[13] vdd gnd cell_6t
Xbit_r14_c107 bl[107] br[107] wl[14] vdd gnd cell_6t
Xbit_r15_c107 bl[107] br[107] wl[15] vdd gnd cell_6t
Xbit_r16_c107 bl[107] br[107] wl[16] vdd gnd cell_6t
Xbit_r17_c107 bl[107] br[107] wl[17] vdd gnd cell_6t
Xbit_r18_c107 bl[107] br[107] wl[18] vdd gnd cell_6t
Xbit_r19_c107 bl[107] br[107] wl[19] vdd gnd cell_6t
Xbit_r20_c107 bl[107] br[107] wl[20] vdd gnd cell_6t
Xbit_r21_c107 bl[107] br[107] wl[21] vdd gnd cell_6t
Xbit_r22_c107 bl[107] br[107] wl[22] vdd gnd cell_6t
Xbit_r23_c107 bl[107] br[107] wl[23] vdd gnd cell_6t
Xbit_r24_c107 bl[107] br[107] wl[24] vdd gnd cell_6t
Xbit_r25_c107 bl[107] br[107] wl[25] vdd gnd cell_6t
Xbit_r26_c107 bl[107] br[107] wl[26] vdd gnd cell_6t
Xbit_r27_c107 bl[107] br[107] wl[27] vdd gnd cell_6t
Xbit_r28_c107 bl[107] br[107] wl[28] vdd gnd cell_6t
Xbit_r29_c107 bl[107] br[107] wl[29] vdd gnd cell_6t
Xbit_r30_c107 bl[107] br[107] wl[30] vdd gnd cell_6t
Xbit_r31_c107 bl[107] br[107] wl[31] vdd gnd cell_6t
Xbit_r32_c107 bl[107] br[107] wl[32] vdd gnd cell_6t
Xbit_r33_c107 bl[107] br[107] wl[33] vdd gnd cell_6t
Xbit_r34_c107 bl[107] br[107] wl[34] vdd gnd cell_6t
Xbit_r35_c107 bl[107] br[107] wl[35] vdd gnd cell_6t
Xbit_r36_c107 bl[107] br[107] wl[36] vdd gnd cell_6t
Xbit_r37_c107 bl[107] br[107] wl[37] vdd gnd cell_6t
Xbit_r38_c107 bl[107] br[107] wl[38] vdd gnd cell_6t
Xbit_r39_c107 bl[107] br[107] wl[39] vdd gnd cell_6t
Xbit_r40_c107 bl[107] br[107] wl[40] vdd gnd cell_6t
Xbit_r41_c107 bl[107] br[107] wl[41] vdd gnd cell_6t
Xbit_r42_c107 bl[107] br[107] wl[42] vdd gnd cell_6t
Xbit_r43_c107 bl[107] br[107] wl[43] vdd gnd cell_6t
Xbit_r44_c107 bl[107] br[107] wl[44] vdd gnd cell_6t
Xbit_r45_c107 bl[107] br[107] wl[45] vdd gnd cell_6t
Xbit_r46_c107 bl[107] br[107] wl[46] vdd gnd cell_6t
Xbit_r47_c107 bl[107] br[107] wl[47] vdd gnd cell_6t
Xbit_r48_c107 bl[107] br[107] wl[48] vdd gnd cell_6t
Xbit_r49_c107 bl[107] br[107] wl[49] vdd gnd cell_6t
Xbit_r50_c107 bl[107] br[107] wl[50] vdd gnd cell_6t
Xbit_r51_c107 bl[107] br[107] wl[51] vdd gnd cell_6t
Xbit_r52_c107 bl[107] br[107] wl[52] vdd gnd cell_6t
Xbit_r53_c107 bl[107] br[107] wl[53] vdd gnd cell_6t
Xbit_r54_c107 bl[107] br[107] wl[54] vdd gnd cell_6t
Xbit_r55_c107 bl[107] br[107] wl[55] vdd gnd cell_6t
Xbit_r56_c107 bl[107] br[107] wl[56] vdd gnd cell_6t
Xbit_r57_c107 bl[107] br[107] wl[57] vdd gnd cell_6t
Xbit_r58_c107 bl[107] br[107] wl[58] vdd gnd cell_6t
Xbit_r59_c107 bl[107] br[107] wl[59] vdd gnd cell_6t
Xbit_r60_c107 bl[107] br[107] wl[60] vdd gnd cell_6t
Xbit_r61_c107 bl[107] br[107] wl[61] vdd gnd cell_6t
Xbit_r62_c107 bl[107] br[107] wl[62] vdd gnd cell_6t
Xbit_r63_c107 bl[107] br[107] wl[63] vdd gnd cell_6t
Xbit_r64_c107 bl[107] br[107] wl[64] vdd gnd cell_6t
Xbit_r65_c107 bl[107] br[107] wl[65] vdd gnd cell_6t
Xbit_r66_c107 bl[107] br[107] wl[66] vdd gnd cell_6t
Xbit_r67_c107 bl[107] br[107] wl[67] vdd gnd cell_6t
Xbit_r68_c107 bl[107] br[107] wl[68] vdd gnd cell_6t
Xbit_r69_c107 bl[107] br[107] wl[69] vdd gnd cell_6t
Xbit_r70_c107 bl[107] br[107] wl[70] vdd gnd cell_6t
Xbit_r71_c107 bl[107] br[107] wl[71] vdd gnd cell_6t
Xbit_r72_c107 bl[107] br[107] wl[72] vdd gnd cell_6t
Xbit_r73_c107 bl[107] br[107] wl[73] vdd gnd cell_6t
Xbit_r74_c107 bl[107] br[107] wl[74] vdd gnd cell_6t
Xbit_r75_c107 bl[107] br[107] wl[75] vdd gnd cell_6t
Xbit_r76_c107 bl[107] br[107] wl[76] vdd gnd cell_6t
Xbit_r77_c107 bl[107] br[107] wl[77] vdd gnd cell_6t
Xbit_r78_c107 bl[107] br[107] wl[78] vdd gnd cell_6t
Xbit_r79_c107 bl[107] br[107] wl[79] vdd gnd cell_6t
Xbit_r80_c107 bl[107] br[107] wl[80] vdd gnd cell_6t
Xbit_r81_c107 bl[107] br[107] wl[81] vdd gnd cell_6t
Xbit_r82_c107 bl[107] br[107] wl[82] vdd gnd cell_6t
Xbit_r83_c107 bl[107] br[107] wl[83] vdd gnd cell_6t
Xbit_r84_c107 bl[107] br[107] wl[84] vdd gnd cell_6t
Xbit_r85_c107 bl[107] br[107] wl[85] vdd gnd cell_6t
Xbit_r86_c107 bl[107] br[107] wl[86] vdd gnd cell_6t
Xbit_r87_c107 bl[107] br[107] wl[87] vdd gnd cell_6t
Xbit_r88_c107 bl[107] br[107] wl[88] vdd gnd cell_6t
Xbit_r89_c107 bl[107] br[107] wl[89] vdd gnd cell_6t
Xbit_r90_c107 bl[107] br[107] wl[90] vdd gnd cell_6t
Xbit_r91_c107 bl[107] br[107] wl[91] vdd gnd cell_6t
Xbit_r92_c107 bl[107] br[107] wl[92] vdd gnd cell_6t
Xbit_r93_c107 bl[107] br[107] wl[93] vdd gnd cell_6t
Xbit_r94_c107 bl[107] br[107] wl[94] vdd gnd cell_6t
Xbit_r95_c107 bl[107] br[107] wl[95] vdd gnd cell_6t
Xbit_r96_c107 bl[107] br[107] wl[96] vdd gnd cell_6t
Xbit_r97_c107 bl[107] br[107] wl[97] vdd gnd cell_6t
Xbit_r98_c107 bl[107] br[107] wl[98] vdd gnd cell_6t
Xbit_r99_c107 bl[107] br[107] wl[99] vdd gnd cell_6t
Xbit_r100_c107 bl[107] br[107] wl[100] vdd gnd cell_6t
Xbit_r101_c107 bl[107] br[107] wl[101] vdd gnd cell_6t
Xbit_r102_c107 bl[107] br[107] wl[102] vdd gnd cell_6t
Xbit_r103_c107 bl[107] br[107] wl[103] vdd gnd cell_6t
Xbit_r104_c107 bl[107] br[107] wl[104] vdd gnd cell_6t
Xbit_r105_c107 bl[107] br[107] wl[105] vdd gnd cell_6t
Xbit_r106_c107 bl[107] br[107] wl[106] vdd gnd cell_6t
Xbit_r107_c107 bl[107] br[107] wl[107] vdd gnd cell_6t
Xbit_r108_c107 bl[107] br[107] wl[108] vdd gnd cell_6t
Xbit_r109_c107 bl[107] br[107] wl[109] vdd gnd cell_6t
Xbit_r110_c107 bl[107] br[107] wl[110] vdd gnd cell_6t
Xbit_r111_c107 bl[107] br[107] wl[111] vdd gnd cell_6t
Xbit_r112_c107 bl[107] br[107] wl[112] vdd gnd cell_6t
Xbit_r113_c107 bl[107] br[107] wl[113] vdd gnd cell_6t
Xbit_r114_c107 bl[107] br[107] wl[114] vdd gnd cell_6t
Xbit_r115_c107 bl[107] br[107] wl[115] vdd gnd cell_6t
Xbit_r116_c107 bl[107] br[107] wl[116] vdd gnd cell_6t
Xbit_r117_c107 bl[107] br[107] wl[117] vdd gnd cell_6t
Xbit_r118_c107 bl[107] br[107] wl[118] vdd gnd cell_6t
Xbit_r119_c107 bl[107] br[107] wl[119] vdd gnd cell_6t
Xbit_r120_c107 bl[107] br[107] wl[120] vdd gnd cell_6t
Xbit_r121_c107 bl[107] br[107] wl[121] vdd gnd cell_6t
Xbit_r122_c107 bl[107] br[107] wl[122] vdd gnd cell_6t
Xbit_r123_c107 bl[107] br[107] wl[123] vdd gnd cell_6t
Xbit_r124_c107 bl[107] br[107] wl[124] vdd gnd cell_6t
Xbit_r125_c107 bl[107] br[107] wl[125] vdd gnd cell_6t
Xbit_r126_c107 bl[107] br[107] wl[126] vdd gnd cell_6t
Xbit_r127_c107 bl[107] br[107] wl[127] vdd gnd cell_6t
Xbit_r0_c108 bl[108] br[108] wl[0] vdd gnd cell_6t
Xbit_r1_c108 bl[108] br[108] wl[1] vdd gnd cell_6t
Xbit_r2_c108 bl[108] br[108] wl[2] vdd gnd cell_6t
Xbit_r3_c108 bl[108] br[108] wl[3] vdd gnd cell_6t
Xbit_r4_c108 bl[108] br[108] wl[4] vdd gnd cell_6t
Xbit_r5_c108 bl[108] br[108] wl[5] vdd gnd cell_6t
Xbit_r6_c108 bl[108] br[108] wl[6] vdd gnd cell_6t
Xbit_r7_c108 bl[108] br[108] wl[7] vdd gnd cell_6t
Xbit_r8_c108 bl[108] br[108] wl[8] vdd gnd cell_6t
Xbit_r9_c108 bl[108] br[108] wl[9] vdd gnd cell_6t
Xbit_r10_c108 bl[108] br[108] wl[10] vdd gnd cell_6t
Xbit_r11_c108 bl[108] br[108] wl[11] vdd gnd cell_6t
Xbit_r12_c108 bl[108] br[108] wl[12] vdd gnd cell_6t
Xbit_r13_c108 bl[108] br[108] wl[13] vdd gnd cell_6t
Xbit_r14_c108 bl[108] br[108] wl[14] vdd gnd cell_6t
Xbit_r15_c108 bl[108] br[108] wl[15] vdd gnd cell_6t
Xbit_r16_c108 bl[108] br[108] wl[16] vdd gnd cell_6t
Xbit_r17_c108 bl[108] br[108] wl[17] vdd gnd cell_6t
Xbit_r18_c108 bl[108] br[108] wl[18] vdd gnd cell_6t
Xbit_r19_c108 bl[108] br[108] wl[19] vdd gnd cell_6t
Xbit_r20_c108 bl[108] br[108] wl[20] vdd gnd cell_6t
Xbit_r21_c108 bl[108] br[108] wl[21] vdd gnd cell_6t
Xbit_r22_c108 bl[108] br[108] wl[22] vdd gnd cell_6t
Xbit_r23_c108 bl[108] br[108] wl[23] vdd gnd cell_6t
Xbit_r24_c108 bl[108] br[108] wl[24] vdd gnd cell_6t
Xbit_r25_c108 bl[108] br[108] wl[25] vdd gnd cell_6t
Xbit_r26_c108 bl[108] br[108] wl[26] vdd gnd cell_6t
Xbit_r27_c108 bl[108] br[108] wl[27] vdd gnd cell_6t
Xbit_r28_c108 bl[108] br[108] wl[28] vdd gnd cell_6t
Xbit_r29_c108 bl[108] br[108] wl[29] vdd gnd cell_6t
Xbit_r30_c108 bl[108] br[108] wl[30] vdd gnd cell_6t
Xbit_r31_c108 bl[108] br[108] wl[31] vdd gnd cell_6t
Xbit_r32_c108 bl[108] br[108] wl[32] vdd gnd cell_6t
Xbit_r33_c108 bl[108] br[108] wl[33] vdd gnd cell_6t
Xbit_r34_c108 bl[108] br[108] wl[34] vdd gnd cell_6t
Xbit_r35_c108 bl[108] br[108] wl[35] vdd gnd cell_6t
Xbit_r36_c108 bl[108] br[108] wl[36] vdd gnd cell_6t
Xbit_r37_c108 bl[108] br[108] wl[37] vdd gnd cell_6t
Xbit_r38_c108 bl[108] br[108] wl[38] vdd gnd cell_6t
Xbit_r39_c108 bl[108] br[108] wl[39] vdd gnd cell_6t
Xbit_r40_c108 bl[108] br[108] wl[40] vdd gnd cell_6t
Xbit_r41_c108 bl[108] br[108] wl[41] vdd gnd cell_6t
Xbit_r42_c108 bl[108] br[108] wl[42] vdd gnd cell_6t
Xbit_r43_c108 bl[108] br[108] wl[43] vdd gnd cell_6t
Xbit_r44_c108 bl[108] br[108] wl[44] vdd gnd cell_6t
Xbit_r45_c108 bl[108] br[108] wl[45] vdd gnd cell_6t
Xbit_r46_c108 bl[108] br[108] wl[46] vdd gnd cell_6t
Xbit_r47_c108 bl[108] br[108] wl[47] vdd gnd cell_6t
Xbit_r48_c108 bl[108] br[108] wl[48] vdd gnd cell_6t
Xbit_r49_c108 bl[108] br[108] wl[49] vdd gnd cell_6t
Xbit_r50_c108 bl[108] br[108] wl[50] vdd gnd cell_6t
Xbit_r51_c108 bl[108] br[108] wl[51] vdd gnd cell_6t
Xbit_r52_c108 bl[108] br[108] wl[52] vdd gnd cell_6t
Xbit_r53_c108 bl[108] br[108] wl[53] vdd gnd cell_6t
Xbit_r54_c108 bl[108] br[108] wl[54] vdd gnd cell_6t
Xbit_r55_c108 bl[108] br[108] wl[55] vdd gnd cell_6t
Xbit_r56_c108 bl[108] br[108] wl[56] vdd gnd cell_6t
Xbit_r57_c108 bl[108] br[108] wl[57] vdd gnd cell_6t
Xbit_r58_c108 bl[108] br[108] wl[58] vdd gnd cell_6t
Xbit_r59_c108 bl[108] br[108] wl[59] vdd gnd cell_6t
Xbit_r60_c108 bl[108] br[108] wl[60] vdd gnd cell_6t
Xbit_r61_c108 bl[108] br[108] wl[61] vdd gnd cell_6t
Xbit_r62_c108 bl[108] br[108] wl[62] vdd gnd cell_6t
Xbit_r63_c108 bl[108] br[108] wl[63] vdd gnd cell_6t
Xbit_r64_c108 bl[108] br[108] wl[64] vdd gnd cell_6t
Xbit_r65_c108 bl[108] br[108] wl[65] vdd gnd cell_6t
Xbit_r66_c108 bl[108] br[108] wl[66] vdd gnd cell_6t
Xbit_r67_c108 bl[108] br[108] wl[67] vdd gnd cell_6t
Xbit_r68_c108 bl[108] br[108] wl[68] vdd gnd cell_6t
Xbit_r69_c108 bl[108] br[108] wl[69] vdd gnd cell_6t
Xbit_r70_c108 bl[108] br[108] wl[70] vdd gnd cell_6t
Xbit_r71_c108 bl[108] br[108] wl[71] vdd gnd cell_6t
Xbit_r72_c108 bl[108] br[108] wl[72] vdd gnd cell_6t
Xbit_r73_c108 bl[108] br[108] wl[73] vdd gnd cell_6t
Xbit_r74_c108 bl[108] br[108] wl[74] vdd gnd cell_6t
Xbit_r75_c108 bl[108] br[108] wl[75] vdd gnd cell_6t
Xbit_r76_c108 bl[108] br[108] wl[76] vdd gnd cell_6t
Xbit_r77_c108 bl[108] br[108] wl[77] vdd gnd cell_6t
Xbit_r78_c108 bl[108] br[108] wl[78] vdd gnd cell_6t
Xbit_r79_c108 bl[108] br[108] wl[79] vdd gnd cell_6t
Xbit_r80_c108 bl[108] br[108] wl[80] vdd gnd cell_6t
Xbit_r81_c108 bl[108] br[108] wl[81] vdd gnd cell_6t
Xbit_r82_c108 bl[108] br[108] wl[82] vdd gnd cell_6t
Xbit_r83_c108 bl[108] br[108] wl[83] vdd gnd cell_6t
Xbit_r84_c108 bl[108] br[108] wl[84] vdd gnd cell_6t
Xbit_r85_c108 bl[108] br[108] wl[85] vdd gnd cell_6t
Xbit_r86_c108 bl[108] br[108] wl[86] vdd gnd cell_6t
Xbit_r87_c108 bl[108] br[108] wl[87] vdd gnd cell_6t
Xbit_r88_c108 bl[108] br[108] wl[88] vdd gnd cell_6t
Xbit_r89_c108 bl[108] br[108] wl[89] vdd gnd cell_6t
Xbit_r90_c108 bl[108] br[108] wl[90] vdd gnd cell_6t
Xbit_r91_c108 bl[108] br[108] wl[91] vdd gnd cell_6t
Xbit_r92_c108 bl[108] br[108] wl[92] vdd gnd cell_6t
Xbit_r93_c108 bl[108] br[108] wl[93] vdd gnd cell_6t
Xbit_r94_c108 bl[108] br[108] wl[94] vdd gnd cell_6t
Xbit_r95_c108 bl[108] br[108] wl[95] vdd gnd cell_6t
Xbit_r96_c108 bl[108] br[108] wl[96] vdd gnd cell_6t
Xbit_r97_c108 bl[108] br[108] wl[97] vdd gnd cell_6t
Xbit_r98_c108 bl[108] br[108] wl[98] vdd gnd cell_6t
Xbit_r99_c108 bl[108] br[108] wl[99] vdd gnd cell_6t
Xbit_r100_c108 bl[108] br[108] wl[100] vdd gnd cell_6t
Xbit_r101_c108 bl[108] br[108] wl[101] vdd gnd cell_6t
Xbit_r102_c108 bl[108] br[108] wl[102] vdd gnd cell_6t
Xbit_r103_c108 bl[108] br[108] wl[103] vdd gnd cell_6t
Xbit_r104_c108 bl[108] br[108] wl[104] vdd gnd cell_6t
Xbit_r105_c108 bl[108] br[108] wl[105] vdd gnd cell_6t
Xbit_r106_c108 bl[108] br[108] wl[106] vdd gnd cell_6t
Xbit_r107_c108 bl[108] br[108] wl[107] vdd gnd cell_6t
Xbit_r108_c108 bl[108] br[108] wl[108] vdd gnd cell_6t
Xbit_r109_c108 bl[108] br[108] wl[109] vdd gnd cell_6t
Xbit_r110_c108 bl[108] br[108] wl[110] vdd gnd cell_6t
Xbit_r111_c108 bl[108] br[108] wl[111] vdd gnd cell_6t
Xbit_r112_c108 bl[108] br[108] wl[112] vdd gnd cell_6t
Xbit_r113_c108 bl[108] br[108] wl[113] vdd gnd cell_6t
Xbit_r114_c108 bl[108] br[108] wl[114] vdd gnd cell_6t
Xbit_r115_c108 bl[108] br[108] wl[115] vdd gnd cell_6t
Xbit_r116_c108 bl[108] br[108] wl[116] vdd gnd cell_6t
Xbit_r117_c108 bl[108] br[108] wl[117] vdd gnd cell_6t
Xbit_r118_c108 bl[108] br[108] wl[118] vdd gnd cell_6t
Xbit_r119_c108 bl[108] br[108] wl[119] vdd gnd cell_6t
Xbit_r120_c108 bl[108] br[108] wl[120] vdd gnd cell_6t
Xbit_r121_c108 bl[108] br[108] wl[121] vdd gnd cell_6t
Xbit_r122_c108 bl[108] br[108] wl[122] vdd gnd cell_6t
Xbit_r123_c108 bl[108] br[108] wl[123] vdd gnd cell_6t
Xbit_r124_c108 bl[108] br[108] wl[124] vdd gnd cell_6t
Xbit_r125_c108 bl[108] br[108] wl[125] vdd gnd cell_6t
Xbit_r126_c108 bl[108] br[108] wl[126] vdd gnd cell_6t
Xbit_r127_c108 bl[108] br[108] wl[127] vdd gnd cell_6t
Xbit_r0_c109 bl[109] br[109] wl[0] vdd gnd cell_6t
Xbit_r1_c109 bl[109] br[109] wl[1] vdd gnd cell_6t
Xbit_r2_c109 bl[109] br[109] wl[2] vdd gnd cell_6t
Xbit_r3_c109 bl[109] br[109] wl[3] vdd gnd cell_6t
Xbit_r4_c109 bl[109] br[109] wl[4] vdd gnd cell_6t
Xbit_r5_c109 bl[109] br[109] wl[5] vdd gnd cell_6t
Xbit_r6_c109 bl[109] br[109] wl[6] vdd gnd cell_6t
Xbit_r7_c109 bl[109] br[109] wl[7] vdd gnd cell_6t
Xbit_r8_c109 bl[109] br[109] wl[8] vdd gnd cell_6t
Xbit_r9_c109 bl[109] br[109] wl[9] vdd gnd cell_6t
Xbit_r10_c109 bl[109] br[109] wl[10] vdd gnd cell_6t
Xbit_r11_c109 bl[109] br[109] wl[11] vdd gnd cell_6t
Xbit_r12_c109 bl[109] br[109] wl[12] vdd gnd cell_6t
Xbit_r13_c109 bl[109] br[109] wl[13] vdd gnd cell_6t
Xbit_r14_c109 bl[109] br[109] wl[14] vdd gnd cell_6t
Xbit_r15_c109 bl[109] br[109] wl[15] vdd gnd cell_6t
Xbit_r16_c109 bl[109] br[109] wl[16] vdd gnd cell_6t
Xbit_r17_c109 bl[109] br[109] wl[17] vdd gnd cell_6t
Xbit_r18_c109 bl[109] br[109] wl[18] vdd gnd cell_6t
Xbit_r19_c109 bl[109] br[109] wl[19] vdd gnd cell_6t
Xbit_r20_c109 bl[109] br[109] wl[20] vdd gnd cell_6t
Xbit_r21_c109 bl[109] br[109] wl[21] vdd gnd cell_6t
Xbit_r22_c109 bl[109] br[109] wl[22] vdd gnd cell_6t
Xbit_r23_c109 bl[109] br[109] wl[23] vdd gnd cell_6t
Xbit_r24_c109 bl[109] br[109] wl[24] vdd gnd cell_6t
Xbit_r25_c109 bl[109] br[109] wl[25] vdd gnd cell_6t
Xbit_r26_c109 bl[109] br[109] wl[26] vdd gnd cell_6t
Xbit_r27_c109 bl[109] br[109] wl[27] vdd gnd cell_6t
Xbit_r28_c109 bl[109] br[109] wl[28] vdd gnd cell_6t
Xbit_r29_c109 bl[109] br[109] wl[29] vdd gnd cell_6t
Xbit_r30_c109 bl[109] br[109] wl[30] vdd gnd cell_6t
Xbit_r31_c109 bl[109] br[109] wl[31] vdd gnd cell_6t
Xbit_r32_c109 bl[109] br[109] wl[32] vdd gnd cell_6t
Xbit_r33_c109 bl[109] br[109] wl[33] vdd gnd cell_6t
Xbit_r34_c109 bl[109] br[109] wl[34] vdd gnd cell_6t
Xbit_r35_c109 bl[109] br[109] wl[35] vdd gnd cell_6t
Xbit_r36_c109 bl[109] br[109] wl[36] vdd gnd cell_6t
Xbit_r37_c109 bl[109] br[109] wl[37] vdd gnd cell_6t
Xbit_r38_c109 bl[109] br[109] wl[38] vdd gnd cell_6t
Xbit_r39_c109 bl[109] br[109] wl[39] vdd gnd cell_6t
Xbit_r40_c109 bl[109] br[109] wl[40] vdd gnd cell_6t
Xbit_r41_c109 bl[109] br[109] wl[41] vdd gnd cell_6t
Xbit_r42_c109 bl[109] br[109] wl[42] vdd gnd cell_6t
Xbit_r43_c109 bl[109] br[109] wl[43] vdd gnd cell_6t
Xbit_r44_c109 bl[109] br[109] wl[44] vdd gnd cell_6t
Xbit_r45_c109 bl[109] br[109] wl[45] vdd gnd cell_6t
Xbit_r46_c109 bl[109] br[109] wl[46] vdd gnd cell_6t
Xbit_r47_c109 bl[109] br[109] wl[47] vdd gnd cell_6t
Xbit_r48_c109 bl[109] br[109] wl[48] vdd gnd cell_6t
Xbit_r49_c109 bl[109] br[109] wl[49] vdd gnd cell_6t
Xbit_r50_c109 bl[109] br[109] wl[50] vdd gnd cell_6t
Xbit_r51_c109 bl[109] br[109] wl[51] vdd gnd cell_6t
Xbit_r52_c109 bl[109] br[109] wl[52] vdd gnd cell_6t
Xbit_r53_c109 bl[109] br[109] wl[53] vdd gnd cell_6t
Xbit_r54_c109 bl[109] br[109] wl[54] vdd gnd cell_6t
Xbit_r55_c109 bl[109] br[109] wl[55] vdd gnd cell_6t
Xbit_r56_c109 bl[109] br[109] wl[56] vdd gnd cell_6t
Xbit_r57_c109 bl[109] br[109] wl[57] vdd gnd cell_6t
Xbit_r58_c109 bl[109] br[109] wl[58] vdd gnd cell_6t
Xbit_r59_c109 bl[109] br[109] wl[59] vdd gnd cell_6t
Xbit_r60_c109 bl[109] br[109] wl[60] vdd gnd cell_6t
Xbit_r61_c109 bl[109] br[109] wl[61] vdd gnd cell_6t
Xbit_r62_c109 bl[109] br[109] wl[62] vdd gnd cell_6t
Xbit_r63_c109 bl[109] br[109] wl[63] vdd gnd cell_6t
Xbit_r64_c109 bl[109] br[109] wl[64] vdd gnd cell_6t
Xbit_r65_c109 bl[109] br[109] wl[65] vdd gnd cell_6t
Xbit_r66_c109 bl[109] br[109] wl[66] vdd gnd cell_6t
Xbit_r67_c109 bl[109] br[109] wl[67] vdd gnd cell_6t
Xbit_r68_c109 bl[109] br[109] wl[68] vdd gnd cell_6t
Xbit_r69_c109 bl[109] br[109] wl[69] vdd gnd cell_6t
Xbit_r70_c109 bl[109] br[109] wl[70] vdd gnd cell_6t
Xbit_r71_c109 bl[109] br[109] wl[71] vdd gnd cell_6t
Xbit_r72_c109 bl[109] br[109] wl[72] vdd gnd cell_6t
Xbit_r73_c109 bl[109] br[109] wl[73] vdd gnd cell_6t
Xbit_r74_c109 bl[109] br[109] wl[74] vdd gnd cell_6t
Xbit_r75_c109 bl[109] br[109] wl[75] vdd gnd cell_6t
Xbit_r76_c109 bl[109] br[109] wl[76] vdd gnd cell_6t
Xbit_r77_c109 bl[109] br[109] wl[77] vdd gnd cell_6t
Xbit_r78_c109 bl[109] br[109] wl[78] vdd gnd cell_6t
Xbit_r79_c109 bl[109] br[109] wl[79] vdd gnd cell_6t
Xbit_r80_c109 bl[109] br[109] wl[80] vdd gnd cell_6t
Xbit_r81_c109 bl[109] br[109] wl[81] vdd gnd cell_6t
Xbit_r82_c109 bl[109] br[109] wl[82] vdd gnd cell_6t
Xbit_r83_c109 bl[109] br[109] wl[83] vdd gnd cell_6t
Xbit_r84_c109 bl[109] br[109] wl[84] vdd gnd cell_6t
Xbit_r85_c109 bl[109] br[109] wl[85] vdd gnd cell_6t
Xbit_r86_c109 bl[109] br[109] wl[86] vdd gnd cell_6t
Xbit_r87_c109 bl[109] br[109] wl[87] vdd gnd cell_6t
Xbit_r88_c109 bl[109] br[109] wl[88] vdd gnd cell_6t
Xbit_r89_c109 bl[109] br[109] wl[89] vdd gnd cell_6t
Xbit_r90_c109 bl[109] br[109] wl[90] vdd gnd cell_6t
Xbit_r91_c109 bl[109] br[109] wl[91] vdd gnd cell_6t
Xbit_r92_c109 bl[109] br[109] wl[92] vdd gnd cell_6t
Xbit_r93_c109 bl[109] br[109] wl[93] vdd gnd cell_6t
Xbit_r94_c109 bl[109] br[109] wl[94] vdd gnd cell_6t
Xbit_r95_c109 bl[109] br[109] wl[95] vdd gnd cell_6t
Xbit_r96_c109 bl[109] br[109] wl[96] vdd gnd cell_6t
Xbit_r97_c109 bl[109] br[109] wl[97] vdd gnd cell_6t
Xbit_r98_c109 bl[109] br[109] wl[98] vdd gnd cell_6t
Xbit_r99_c109 bl[109] br[109] wl[99] vdd gnd cell_6t
Xbit_r100_c109 bl[109] br[109] wl[100] vdd gnd cell_6t
Xbit_r101_c109 bl[109] br[109] wl[101] vdd gnd cell_6t
Xbit_r102_c109 bl[109] br[109] wl[102] vdd gnd cell_6t
Xbit_r103_c109 bl[109] br[109] wl[103] vdd gnd cell_6t
Xbit_r104_c109 bl[109] br[109] wl[104] vdd gnd cell_6t
Xbit_r105_c109 bl[109] br[109] wl[105] vdd gnd cell_6t
Xbit_r106_c109 bl[109] br[109] wl[106] vdd gnd cell_6t
Xbit_r107_c109 bl[109] br[109] wl[107] vdd gnd cell_6t
Xbit_r108_c109 bl[109] br[109] wl[108] vdd gnd cell_6t
Xbit_r109_c109 bl[109] br[109] wl[109] vdd gnd cell_6t
Xbit_r110_c109 bl[109] br[109] wl[110] vdd gnd cell_6t
Xbit_r111_c109 bl[109] br[109] wl[111] vdd gnd cell_6t
Xbit_r112_c109 bl[109] br[109] wl[112] vdd gnd cell_6t
Xbit_r113_c109 bl[109] br[109] wl[113] vdd gnd cell_6t
Xbit_r114_c109 bl[109] br[109] wl[114] vdd gnd cell_6t
Xbit_r115_c109 bl[109] br[109] wl[115] vdd gnd cell_6t
Xbit_r116_c109 bl[109] br[109] wl[116] vdd gnd cell_6t
Xbit_r117_c109 bl[109] br[109] wl[117] vdd gnd cell_6t
Xbit_r118_c109 bl[109] br[109] wl[118] vdd gnd cell_6t
Xbit_r119_c109 bl[109] br[109] wl[119] vdd gnd cell_6t
Xbit_r120_c109 bl[109] br[109] wl[120] vdd gnd cell_6t
Xbit_r121_c109 bl[109] br[109] wl[121] vdd gnd cell_6t
Xbit_r122_c109 bl[109] br[109] wl[122] vdd gnd cell_6t
Xbit_r123_c109 bl[109] br[109] wl[123] vdd gnd cell_6t
Xbit_r124_c109 bl[109] br[109] wl[124] vdd gnd cell_6t
Xbit_r125_c109 bl[109] br[109] wl[125] vdd gnd cell_6t
Xbit_r126_c109 bl[109] br[109] wl[126] vdd gnd cell_6t
Xbit_r127_c109 bl[109] br[109] wl[127] vdd gnd cell_6t
Xbit_r0_c110 bl[110] br[110] wl[0] vdd gnd cell_6t
Xbit_r1_c110 bl[110] br[110] wl[1] vdd gnd cell_6t
Xbit_r2_c110 bl[110] br[110] wl[2] vdd gnd cell_6t
Xbit_r3_c110 bl[110] br[110] wl[3] vdd gnd cell_6t
Xbit_r4_c110 bl[110] br[110] wl[4] vdd gnd cell_6t
Xbit_r5_c110 bl[110] br[110] wl[5] vdd gnd cell_6t
Xbit_r6_c110 bl[110] br[110] wl[6] vdd gnd cell_6t
Xbit_r7_c110 bl[110] br[110] wl[7] vdd gnd cell_6t
Xbit_r8_c110 bl[110] br[110] wl[8] vdd gnd cell_6t
Xbit_r9_c110 bl[110] br[110] wl[9] vdd gnd cell_6t
Xbit_r10_c110 bl[110] br[110] wl[10] vdd gnd cell_6t
Xbit_r11_c110 bl[110] br[110] wl[11] vdd gnd cell_6t
Xbit_r12_c110 bl[110] br[110] wl[12] vdd gnd cell_6t
Xbit_r13_c110 bl[110] br[110] wl[13] vdd gnd cell_6t
Xbit_r14_c110 bl[110] br[110] wl[14] vdd gnd cell_6t
Xbit_r15_c110 bl[110] br[110] wl[15] vdd gnd cell_6t
Xbit_r16_c110 bl[110] br[110] wl[16] vdd gnd cell_6t
Xbit_r17_c110 bl[110] br[110] wl[17] vdd gnd cell_6t
Xbit_r18_c110 bl[110] br[110] wl[18] vdd gnd cell_6t
Xbit_r19_c110 bl[110] br[110] wl[19] vdd gnd cell_6t
Xbit_r20_c110 bl[110] br[110] wl[20] vdd gnd cell_6t
Xbit_r21_c110 bl[110] br[110] wl[21] vdd gnd cell_6t
Xbit_r22_c110 bl[110] br[110] wl[22] vdd gnd cell_6t
Xbit_r23_c110 bl[110] br[110] wl[23] vdd gnd cell_6t
Xbit_r24_c110 bl[110] br[110] wl[24] vdd gnd cell_6t
Xbit_r25_c110 bl[110] br[110] wl[25] vdd gnd cell_6t
Xbit_r26_c110 bl[110] br[110] wl[26] vdd gnd cell_6t
Xbit_r27_c110 bl[110] br[110] wl[27] vdd gnd cell_6t
Xbit_r28_c110 bl[110] br[110] wl[28] vdd gnd cell_6t
Xbit_r29_c110 bl[110] br[110] wl[29] vdd gnd cell_6t
Xbit_r30_c110 bl[110] br[110] wl[30] vdd gnd cell_6t
Xbit_r31_c110 bl[110] br[110] wl[31] vdd gnd cell_6t
Xbit_r32_c110 bl[110] br[110] wl[32] vdd gnd cell_6t
Xbit_r33_c110 bl[110] br[110] wl[33] vdd gnd cell_6t
Xbit_r34_c110 bl[110] br[110] wl[34] vdd gnd cell_6t
Xbit_r35_c110 bl[110] br[110] wl[35] vdd gnd cell_6t
Xbit_r36_c110 bl[110] br[110] wl[36] vdd gnd cell_6t
Xbit_r37_c110 bl[110] br[110] wl[37] vdd gnd cell_6t
Xbit_r38_c110 bl[110] br[110] wl[38] vdd gnd cell_6t
Xbit_r39_c110 bl[110] br[110] wl[39] vdd gnd cell_6t
Xbit_r40_c110 bl[110] br[110] wl[40] vdd gnd cell_6t
Xbit_r41_c110 bl[110] br[110] wl[41] vdd gnd cell_6t
Xbit_r42_c110 bl[110] br[110] wl[42] vdd gnd cell_6t
Xbit_r43_c110 bl[110] br[110] wl[43] vdd gnd cell_6t
Xbit_r44_c110 bl[110] br[110] wl[44] vdd gnd cell_6t
Xbit_r45_c110 bl[110] br[110] wl[45] vdd gnd cell_6t
Xbit_r46_c110 bl[110] br[110] wl[46] vdd gnd cell_6t
Xbit_r47_c110 bl[110] br[110] wl[47] vdd gnd cell_6t
Xbit_r48_c110 bl[110] br[110] wl[48] vdd gnd cell_6t
Xbit_r49_c110 bl[110] br[110] wl[49] vdd gnd cell_6t
Xbit_r50_c110 bl[110] br[110] wl[50] vdd gnd cell_6t
Xbit_r51_c110 bl[110] br[110] wl[51] vdd gnd cell_6t
Xbit_r52_c110 bl[110] br[110] wl[52] vdd gnd cell_6t
Xbit_r53_c110 bl[110] br[110] wl[53] vdd gnd cell_6t
Xbit_r54_c110 bl[110] br[110] wl[54] vdd gnd cell_6t
Xbit_r55_c110 bl[110] br[110] wl[55] vdd gnd cell_6t
Xbit_r56_c110 bl[110] br[110] wl[56] vdd gnd cell_6t
Xbit_r57_c110 bl[110] br[110] wl[57] vdd gnd cell_6t
Xbit_r58_c110 bl[110] br[110] wl[58] vdd gnd cell_6t
Xbit_r59_c110 bl[110] br[110] wl[59] vdd gnd cell_6t
Xbit_r60_c110 bl[110] br[110] wl[60] vdd gnd cell_6t
Xbit_r61_c110 bl[110] br[110] wl[61] vdd gnd cell_6t
Xbit_r62_c110 bl[110] br[110] wl[62] vdd gnd cell_6t
Xbit_r63_c110 bl[110] br[110] wl[63] vdd gnd cell_6t
Xbit_r64_c110 bl[110] br[110] wl[64] vdd gnd cell_6t
Xbit_r65_c110 bl[110] br[110] wl[65] vdd gnd cell_6t
Xbit_r66_c110 bl[110] br[110] wl[66] vdd gnd cell_6t
Xbit_r67_c110 bl[110] br[110] wl[67] vdd gnd cell_6t
Xbit_r68_c110 bl[110] br[110] wl[68] vdd gnd cell_6t
Xbit_r69_c110 bl[110] br[110] wl[69] vdd gnd cell_6t
Xbit_r70_c110 bl[110] br[110] wl[70] vdd gnd cell_6t
Xbit_r71_c110 bl[110] br[110] wl[71] vdd gnd cell_6t
Xbit_r72_c110 bl[110] br[110] wl[72] vdd gnd cell_6t
Xbit_r73_c110 bl[110] br[110] wl[73] vdd gnd cell_6t
Xbit_r74_c110 bl[110] br[110] wl[74] vdd gnd cell_6t
Xbit_r75_c110 bl[110] br[110] wl[75] vdd gnd cell_6t
Xbit_r76_c110 bl[110] br[110] wl[76] vdd gnd cell_6t
Xbit_r77_c110 bl[110] br[110] wl[77] vdd gnd cell_6t
Xbit_r78_c110 bl[110] br[110] wl[78] vdd gnd cell_6t
Xbit_r79_c110 bl[110] br[110] wl[79] vdd gnd cell_6t
Xbit_r80_c110 bl[110] br[110] wl[80] vdd gnd cell_6t
Xbit_r81_c110 bl[110] br[110] wl[81] vdd gnd cell_6t
Xbit_r82_c110 bl[110] br[110] wl[82] vdd gnd cell_6t
Xbit_r83_c110 bl[110] br[110] wl[83] vdd gnd cell_6t
Xbit_r84_c110 bl[110] br[110] wl[84] vdd gnd cell_6t
Xbit_r85_c110 bl[110] br[110] wl[85] vdd gnd cell_6t
Xbit_r86_c110 bl[110] br[110] wl[86] vdd gnd cell_6t
Xbit_r87_c110 bl[110] br[110] wl[87] vdd gnd cell_6t
Xbit_r88_c110 bl[110] br[110] wl[88] vdd gnd cell_6t
Xbit_r89_c110 bl[110] br[110] wl[89] vdd gnd cell_6t
Xbit_r90_c110 bl[110] br[110] wl[90] vdd gnd cell_6t
Xbit_r91_c110 bl[110] br[110] wl[91] vdd gnd cell_6t
Xbit_r92_c110 bl[110] br[110] wl[92] vdd gnd cell_6t
Xbit_r93_c110 bl[110] br[110] wl[93] vdd gnd cell_6t
Xbit_r94_c110 bl[110] br[110] wl[94] vdd gnd cell_6t
Xbit_r95_c110 bl[110] br[110] wl[95] vdd gnd cell_6t
Xbit_r96_c110 bl[110] br[110] wl[96] vdd gnd cell_6t
Xbit_r97_c110 bl[110] br[110] wl[97] vdd gnd cell_6t
Xbit_r98_c110 bl[110] br[110] wl[98] vdd gnd cell_6t
Xbit_r99_c110 bl[110] br[110] wl[99] vdd gnd cell_6t
Xbit_r100_c110 bl[110] br[110] wl[100] vdd gnd cell_6t
Xbit_r101_c110 bl[110] br[110] wl[101] vdd gnd cell_6t
Xbit_r102_c110 bl[110] br[110] wl[102] vdd gnd cell_6t
Xbit_r103_c110 bl[110] br[110] wl[103] vdd gnd cell_6t
Xbit_r104_c110 bl[110] br[110] wl[104] vdd gnd cell_6t
Xbit_r105_c110 bl[110] br[110] wl[105] vdd gnd cell_6t
Xbit_r106_c110 bl[110] br[110] wl[106] vdd gnd cell_6t
Xbit_r107_c110 bl[110] br[110] wl[107] vdd gnd cell_6t
Xbit_r108_c110 bl[110] br[110] wl[108] vdd gnd cell_6t
Xbit_r109_c110 bl[110] br[110] wl[109] vdd gnd cell_6t
Xbit_r110_c110 bl[110] br[110] wl[110] vdd gnd cell_6t
Xbit_r111_c110 bl[110] br[110] wl[111] vdd gnd cell_6t
Xbit_r112_c110 bl[110] br[110] wl[112] vdd gnd cell_6t
Xbit_r113_c110 bl[110] br[110] wl[113] vdd gnd cell_6t
Xbit_r114_c110 bl[110] br[110] wl[114] vdd gnd cell_6t
Xbit_r115_c110 bl[110] br[110] wl[115] vdd gnd cell_6t
Xbit_r116_c110 bl[110] br[110] wl[116] vdd gnd cell_6t
Xbit_r117_c110 bl[110] br[110] wl[117] vdd gnd cell_6t
Xbit_r118_c110 bl[110] br[110] wl[118] vdd gnd cell_6t
Xbit_r119_c110 bl[110] br[110] wl[119] vdd gnd cell_6t
Xbit_r120_c110 bl[110] br[110] wl[120] vdd gnd cell_6t
Xbit_r121_c110 bl[110] br[110] wl[121] vdd gnd cell_6t
Xbit_r122_c110 bl[110] br[110] wl[122] vdd gnd cell_6t
Xbit_r123_c110 bl[110] br[110] wl[123] vdd gnd cell_6t
Xbit_r124_c110 bl[110] br[110] wl[124] vdd gnd cell_6t
Xbit_r125_c110 bl[110] br[110] wl[125] vdd gnd cell_6t
Xbit_r126_c110 bl[110] br[110] wl[126] vdd gnd cell_6t
Xbit_r127_c110 bl[110] br[110] wl[127] vdd gnd cell_6t
Xbit_r0_c111 bl[111] br[111] wl[0] vdd gnd cell_6t
Xbit_r1_c111 bl[111] br[111] wl[1] vdd gnd cell_6t
Xbit_r2_c111 bl[111] br[111] wl[2] vdd gnd cell_6t
Xbit_r3_c111 bl[111] br[111] wl[3] vdd gnd cell_6t
Xbit_r4_c111 bl[111] br[111] wl[4] vdd gnd cell_6t
Xbit_r5_c111 bl[111] br[111] wl[5] vdd gnd cell_6t
Xbit_r6_c111 bl[111] br[111] wl[6] vdd gnd cell_6t
Xbit_r7_c111 bl[111] br[111] wl[7] vdd gnd cell_6t
Xbit_r8_c111 bl[111] br[111] wl[8] vdd gnd cell_6t
Xbit_r9_c111 bl[111] br[111] wl[9] vdd gnd cell_6t
Xbit_r10_c111 bl[111] br[111] wl[10] vdd gnd cell_6t
Xbit_r11_c111 bl[111] br[111] wl[11] vdd gnd cell_6t
Xbit_r12_c111 bl[111] br[111] wl[12] vdd gnd cell_6t
Xbit_r13_c111 bl[111] br[111] wl[13] vdd gnd cell_6t
Xbit_r14_c111 bl[111] br[111] wl[14] vdd gnd cell_6t
Xbit_r15_c111 bl[111] br[111] wl[15] vdd gnd cell_6t
Xbit_r16_c111 bl[111] br[111] wl[16] vdd gnd cell_6t
Xbit_r17_c111 bl[111] br[111] wl[17] vdd gnd cell_6t
Xbit_r18_c111 bl[111] br[111] wl[18] vdd gnd cell_6t
Xbit_r19_c111 bl[111] br[111] wl[19] vdd gnd cell_6t
Xbit_r20_c111 bl[111] br[111] wl[20] vdd gnd cell_6t
Xbit_r21_c111 bl[111] br[111] wl[21] vdd gnd cell_6t
Xbit_r22_c111 bl[111] br[111] wl[22] vdd gnd cell_6t
Xbit_r23_c111 bl[111] br[111] wl[23] vdd gnd cell_6t
Xbit_r24_c111 bl[111] br[111] wl[24] vdd gnd cell_6t
Xbit_r25_c111 bl[111] br[111] wl[25] vdd gnd cell_6t
Xbit_r26_c111 bl[111] br[111] wl[26] vdd gnd cell_6t
Xbit_r27_c111 bl[111] br[111] wl[27] vdd gnd cell_6t
Xbit_r28_c111 bl[111] br[111] wl[28] vdd gnd cell_6t
Xbit_r29_c111 bl[111] br[111] wl[29] vdd gnd cell_6t
Xbit_r30_c111 bl[111] br[111] wl[30] vdd gnd cell_6t
Xbit_r31_c111 bl[111] br[111] wl[31] vdd gnd cell_6t
Xbit_r32_c111 bl[111] br[111] wl[32] vdd gnd cell_6t
Xbit_r33_c111 bl[111] br[111] wl[33] vdd gnd cell_6t
Xbit_r34_c111 bl[111] br[111] wl[34] vdd gnd cell_6t
Xbit_r35_c111 bl[111] br[111] wl[35] vdd gnd cell_6t
Xbit_r36_c111 bl[111] br[111] wl[36] vdd gnd cell_6t
Xbit_r37_c111 bl[111] br[111] wl[37] vdd gnd cell_6t
Xbit_r38_c111 bl[111] br[111] wl[38] vdd gnd cell_6t
Xbit_r39_c111 bl[111] br[111] wl[39] vdd gnd cell_6t
Xbit_r40_c111 bl[111] br[111] wl[40] vdd gnd cell_6t
Xbit_r41_c111 bl[111] br[111] wl[41] vdd gnd cell_6t
Xbit_r42_c111 bl[111] br[111] wl[42] vdd gnd cell_6t
Xbit_r43_c111 bl[111] br[111] wl[43] vdd gnd cell_6t
Xbit_r44_c111 bl[111] br[111] wl[44] vdd gnd cell_6t
Xbit_r45_c111 bl[111] br[111] wl[45] vdd gnd cell_6t
Xbit_r46_c111 bl[111] br[111] wl[46] vdd gnd cell_6t
Xbit_r47_c111 bl[111] br[111] wl[47] vdd gnd cell_6t
Xbit_r48_c111 bl[111] br[111] wl[48] vdd gnd cell_6t
Xbit_r49_c111 bl[111] br[111] wl[49] vdd gnd cell_6t
Xbit_r50_c111 bl[111] br[111] wl[50] vdd gnd cell_6t
Xbit_r51_c111 bl[111] br[111] wl[51] vdd gnd cell_6t
Xbit_r52_c111 bl[111] br[111] wl[52] vdd gnd cell_6t
Xbit_r53_c111 bl[111] br[111] wl[53] vdd gnd cell_6t
Xbit_r54_c111 bl[111] br[111] wl[54] vdd gnd cell_6t
Xbit_r55_c111 bl[111] br[111] wl[55] vdd gnd cell_6t
Xbit_r56_c111 bl[111] br[111] wl[56] vdd gnd cell_6t
Xbit_r57_c111 bl[111] br[111] wl[57] vdd gnd cell_6t
Xbit_r58_c111 bl[111] br[111] wl[58] vdd gnd cell_6t
Xbit_r59_c111 bl[111] br[111] wl[59] vdd gnd cell_6t
Xbit_r60_c111 bl[111] br[111] wl[60] vdd gnd cell_6t
Xbit_r61_c111 bl[111] br[111] wl[61] vdd gnd cell_6t
Xbit_r62_c111 bl[111] br[111] wl[62] vdd gnd cell_6t
Xbit_r63_c111 bl[111] br[111] wl[63] vdd gnd cell_6t
Xbit_r64_c111 bl[111] br[111] wl[64] vdd gnd cell_6t
Xbit_r65_c111 bl[111] br[111] wl[65] vdd gnd cell_6t
Xbit_r66_c111 bl[111] br[111] wl[66] vdd gnd cell_6t
Xbit_r67_c111 bl[111] br[111] wl[67] vdd gnd cell_6t
Xbit_r68_c111 bl[111] br[111] wl[68] vdd gnd cell_6t
Xbit_r69_c111 bl[111] br[111] wl[69] vdd gnd cell_6t
Xbit_r70_c111 bl[111] br[111] wl[70] vdd gnd cell_6t
Xbit_r71_c111 bl[111] br[111] wl[71] vdd gnd cell_6t
Xbit_r72_c111 bl[111] br[111] wl[72] vdd gnd cell_6t
Xbit_r73_c111 bl[111] br[111] wl[73] vdd gnd cell_6t
Xbit_r74_c111 bl[111] br[111] wl[74] vdd gnd cell_6t
Xbit_r75_c111 bl[111] br[111] wl[75] vdd gnd cell_6t
Xbit_r76_c111 bl[111] br[111] wl[76] vdd gnd cell_6t
Xbit_r77_c111 bl[111] br[111] wl[77] vdd gnd cell_6t
Xbit_r78_c111 bl[111] br[111] wl[78] vdd gnd cell_6t
Xbit_r79_c111 bl[111] br[111] wl[79] vdd gnd cell_6t
Xbit_r80_c111 bl[111] br[111] wl[80] vdd gnd cell_6t
Xbit_r81_c111 bl[111] br[111] wl[81] vdd gnd cell_6t
Xbit_r82_c111 bl[111] br[111] wl[82] vdd gnd cell_6t
Xbit_r83_c111 bl[111] br[111] wl[83] vdd gnd cell_6t
Xbit_r84_c111 bl[111] br[111] wl[84] vdd gnd cell_6t
Xbit_r85_c111 bl[111] br[111] wl[85] vdd gnd cell_6t
Xbit_r86_c111 bl[111] br[111] wl[86] vdd gnd cell_6t
Xbit_r87_c111 bl[111] br[111] wl[87] vdd gnd cell_6t
Xbit_r88_c111 bl[111] br[111] wl[88] vdd gnd cell_6t
Xbit_r89_c111 bl[111] br[111] wl[89] vdd gnd cell_6t
Xbit_r90_c111 bl[111] br[111] wl[90] vdd gnd cell_6t
Xbit_r91_c111 bl[111] br[111] wl[91] vdd gnd cell_6t
Xbit_r92_c111 bl[111] br[111] wl[92] vdd gnd cell_6t
Xbit_r93_c111 bl[111] br[111] wl[93] vdd gnd cell_6t
Xbit_r94_c111 bl[111] br[111] wl[94] vdd gnd cell_6t
Xbit_r95_c111 bl[111] br[111] wl[95] vdd gnd cell_6t
Xbit_r96_c111 bl[111] br[111] wl[96] vdd gnd cell_6t
Xbit_r97_c111 bl[111] br[111] wl[97] vdd gnd cell_6t
Xbit_r98_c111 bl[111] br[111] wl[98] vdd gnd cell_6t
Xbit_r99_c111 bl[111] br[111] wl[99] vdd gnd cell_6t
Xbit_r100_c111 bl[111] br[111] wl[100] vdd gnd cell_6t
Xbit_r101_c111 bl[111] br[111] wl[101] vdd gnd cell_6t
Xbit_r102_c111 bl[111] br[111] wl[102] vdd gnd cell_6t
Xbit_r103_c111 bl[111] br[111] wl[103] vdd gnd cell_6t
Xbit_r104_c111 bl[111] br[111] wl[104] vdd gnd cell_6t
Xbit_r105_c111 bl[111] br[111] wl[105] vdd gnd cell_6t
Xbit_r106_c111 bl[111] br[111] wl[106] vdd gnd cell_6t
Xbit_r107_c111 bl[111] br[111] wl[107] vdd gnd cell_6t
Xbit_r108_c111 bl[111] br[111] wl[108] vdd gnd cell_6t
Xbit_r109_c111 bl[111] br[111] wl[109] vdd gnd cell_6t
Xbit_r110_c111 bl[111] br[111] wl[110] vdd gnd cell_6t
Xbit_r111_c111 bl[111] br[111] wl[111] vdd gnd cell_6t
Xbit_r112_c111 bl[111] br[111] wl[112] vdd gnd cell_6t
Xbit_r113_c111 bl[111] br[111] wl[113] vdd gnd cell_6t
Xbit_r114_c111 bl[111] br[111] wl[114] vdd gnd cell_6t
Xbit_r115_c111 bl[111] br[111] wl[115] vdd gnd cell_6t
Xbit_r116_c111 bl[111] br[111] wl[116] vdd gnd cell_6t
Xbit_r117_c111 bl[111] br[111] wl[117] vdd gnd cell_6t
Xbit_r118_c111 bl[111] br[111] wl[118] vdd gnd cell_6t
Xbit_r119_c111 bl[111] br[111] wl[119] vdd gnd cell_6t
Xbit_r120_c111 bl[111] br[111] wl[120] vdd gnd cell_6t
Xbit_r121_c111 bl[111] br[111] wl[121] vdd gnd cell_6t
Xbit_r122_c111 bl[111] br[111] wl[122] vdd gnd cell_6t
Xbit_r123_c111 bl[111] br[111] wl[123] vdd gnd cell_6t
Xbit_r124_c111 bl[111] br[111] wl[124] vdd gnd cell_6t
Xbit_r125_c111 bl[111] br[111] wl[125] vdd gnd cell_6t
Xbit_r126_c111 bl[111] br[111] wl[126] vdd gnd cell_6t
Xbit_r127_c111 bl[111] br[111] wl[127] vdd gnd cell_6t
Xbit_r0_c112 bl[112] br[112] wl[0] vdd gnd cell_6t
Xbit_r1_c112 bl[112] br[112] wl[1] vdd gnd cell_6t
Xbit_r2_c112 bl[112] br[112] wl[2] vdd gnd cell_6t
Xbit_r3_c112 bl[112] br[112] wl[3] vdd gnd cell_6t
Xbit_r4_c112 bl[112] br[112] wl[4] vdd gnd cell_6t
Xbit_r5_c112 bl[112] br[112] wl[5] vdd gnd cell_6t
Xbit_r6_c112 bl[112] br[112] wl[6] vdd gnd cell_6t
Xbit_r7_c112 bl[112] br[112] wl[7] vdd gnd cell_6t
Xbit_r8_c112 bl[112] br[112] wl[8] vdd gnd cell_6t
Xbit_r9_c112 bl[112] br[112] wl[9] vdd gnd cell_6t
Xbit_r10_c112 bl[112] br[112] wl[10] vdd gnd cell_6t
Xbit_r11_c112 bl[112] br[112] wl[11] vdd gnd cell_6t
Xbit_r12_c112 bl[112] br[112] wl[12] vdd gnd cell_6t
Xbit_r13_c112 bl[112] br[112] wl[13] vdd gnd cell_6t
Xbit_r14_c112 bl[112] br[112] wl[14] vdd gnd cell_6t
Xbit_r15_c112 bl[112] br[112] wl[15] vdd gnd cell_6t
Xbit_r16_c112 bl[112] br[112] wl[16] vdd gnd cell_6t
Xbit_r17_c112 bl[112] br[112] wl[17] vdd gnd cell_6t
Xbit_r18_c112 bl[112] br[112] wl[18] vdd gnd cell_6t
Xbit_r19_c112 bl[112] br[112] wl[19] vdd gnd cell_6t
Xbit_r20_c112 bl[112] br[112] wl[20] vdd gnd cell_6t
Xbit_r21_c112 bl[112] br[112] wl[21] vdd gnd cell_6t
Xbit_r22_c112 bl[112] br[112] wl[22] vdd gnd cell_6t
Xbit_r23_c112 bl[112] br[112] wl[23] vdd gnd cell_6t
Xbit_r24_c112 bl[112] br[112] wl[24] vdd gnd cell_6t
Xbit_r25_c112 bl[112] br[112] wl[25] vdd gnd cell_6t
Xbit_r26_c112 bl[112] br[112] wl[26] vdd gnd cell_6t
Xbit_r27_c112 bl[112] br[112] wl[27] vdd gnd cell_6t
Xbit_r28_c112 bl[112] br[112] wl[28] vdd gnd cell_6t
Xbit_r29_c112 bl[112] br[112] wl[29] vdd gnd cell_6t
Xbit_r30_c112 bl[112] br[112] wl[30] vdd gnd cell_6t
Xbit_r31_c112 bl[112] br[112] wl[31] vdd gnd cell_6t
Xbit_r32_c112 bl[112] br[112] wl[32] vdd gnd cell_6t
Xbit_r33_c112 bl[112] br[112] wl[33] vdd gnd cell_6t
Xbit_r34_c112 bl[112] br[112] wl[34] vdd gnd cell_6t
Xbit_r35_c112 bl[112] br[112] wl[35] vdd gnd cell_6t
Xbit_r36_c112 bl[112] br[112] wl[36] vdd gnd cell_6t
Xbit_r37_c112 bl[112] br[112] wl[37] vdd gnd cell_6t
Xbit_r38_c112 bl[112] br[112] wl[38] vdd gnd cell_6t
Xbit_r39_c112 bl[112] br[112] wl[39] vdd gnd cell_6t
Xbit_r40_c112 bl[112] br[112] wl[40] vdd gnd cell_6t
Xbit_r41_c112 bl[112] br[112] wl[41] vdd gnd cell_6t
Xbit_r42_c112 bl[112] br[112] wl[42] vdd gnd cell_6t
Xbit_r43_c112 bl[112] br[112] wl[43] vdd gnd cell_6t
Xbit_r44_c112 bl[112] br[112] wl[44] vdd gnd cell_6t
Xbit_r45_c112 bl[112] br[112] wl[45] vdd gnd cell_6t
Xbit_r46_c112 bl[112] br[112] wl[46] vdd gnd cell_6t
Xbit_r47_c112 bl[112] br[112] wl[47] vdd gnd cell_6t
Xbit_r48_c112 bl[112] br[112] wl[48] vdd gnd cell_6t
Xbit_r49_c112 bl[112] br[112] wl[49] vdd gnd cell_6t
Xbit_r50_c112 bl[112] br[112] wl[50] vdd gnd cell_6t
Xbit_r51_c112 bl[112] br[112] wl[51] vdd gnd cell_6t
Xbit_r52_c112 bl[112] br[112] wl[52] vdd gnd cell_6t
Xbit_r53_c112 bl[112] br[112] wl[53] vdd gnd cell_6t
Xbit_r54_c112 bl[112] br[112] wl[54] vdd gnd cell_6t
Xbit_r55_c112 bl[112] br[112] wl[55] vdd gnd cell_6t
Xbit_r56_c112 bl[112] br[112] wl[56] vdd gnd cell_6t
Xbit_r57_c112 bl[112] br[112] wl[57] vdd gnd cell_6t
Xbit_r58_c112 bl[112] br[112] wl[58] vdd gnd cell_6t
Xbit_r59_c112 bl[112] br[112] wl[59] vdd gnd cell_6t
Xbit_r60_c112 bl[112] br[112] wl[60] vdd gnd cell_6t
Xbit_r61_c112 bl[112] br[112] wl[61] vdd gnd cell_6t
Xbit_r62_c112 bl[112] br[112] wl[62] vdd gnd cell_6t
Xbit_r63_c112 bl[112] br[112] wl[63] vdd gnd cell_6t
Xbit_r64_c112 bl[112] br[112] wl[64] vdd gnd cell_6t
Xbit_r65_c112 bl[112] br[112] wl[65] vdd gnd cell_6t
Xbit_r66_c112 bl[112] br[112] wl[66] vdd gnd cell_6t
Xbit_r67_c112 bl[112] br[112] wl[67] vdd gnd cell_6t
Xbit_r68_c112 bl[112] br[112] wl[68] vdd gnd cell_6t
Xbit_r69_c112 bl[112] br[112] wl[69] vdd gnd cell_6t
Xbit_r70_c112 bl[112] br[112] wl[70] vdd gnd cell_6t
Xbit_r71_c112 bl[112] br[112] wl[71] vdd gnd cell_6t
Xbit_r72_c112 bl[112] br[112] wl[72] vdd gnd cell_6t
Xbit_r73_c112 bl[112] br[112] wl[73] vdd gnd cell_6t
Xbit_r74_c112 bl[112] br[112] wl[74] vdd gnd cell_6t
Xbit_r75_c112 bl[112] br[112] wl[75] vdd gnd cell_6t
Xbit_r76_c112 bl[112] br[112] wl[76] vdd gnd cell_6t
Xbit_r77_c112 bl[112] br[112] wl[77] vdd gnd cell_6t
Xbit_r78_c112 bl[112] br[112] wl[78] vdd gnd cell_6t
Xbit_r79_c112 bl[112] br[112] wl[79] vdd gnd cell_6t
Xbit_r80_c112 bl[112] br[112] wl[80] vdd gnd cell_6t
Xbit_r81_c112 bl[112] br[112] wl[81] vdd gnd cell_6t
Xbit_r82_c112 bl[112] br[112] wl[82] vdd gnd cell_6t
Xbit_r83_c112 bl[112] br[112] wl[83] vdd gnd cell_6t
Xbit_r84_c112 bl[112] br[112] wl[84] vdd gnd cell_6t
Xbit_r85_c112 bl[112] br[112] wl[85] vdd gnd cell_6t
Xbit_r86_c112 bl[112] br[112] wl[86] vdd gnd cell_6t
Xbit_r87_c112 bl[112] br[112] wl[87] vdd gnd cell_6t
Xbit_r88_c112 bl[112] br[112] wl[88] vdd gnd cell_6t
Xbit_r89_c112 bl[112] br[112] wl[89] vdd gnd cell_6t
Xbit_r90_c112 bl[112] br[112] wl[90] vdd gnd cell_6t
Xbit_r91_c112 bl[112] br[112] wl[91] vdd gnd cell_6t
Xbit_r92_c112 bl[112] br[112] wl[92] vdd gnd cell_6t
Xbit_r93_c112 bl[112] br[112] wl[93] vdd gnd cell_6t
Xbit_r94_c112 bl[112] br[112] wl[94] vdd gnd cell_6t
Xbit_r95_c112 bl[112] br[112] wl[95] vdd gnd cell_6t
Xbit_r96_c112 bl[112] br[112] wl[96] vdd gnd cell_6t
Xbit_r97_c112 bl[112] br[112] wl[97] vdd gnd cell_6t
Xbit_r98_c112 bl[112] br[112] wl[98] vdd gnd cell_6t
Xbit_r99_c112 bl[112] br[112] wl[99] vdd gnd cell_6t
Xbit_r100_c112 bl[112] br[112] wl[100] vdd gnd cell_6t
Xbit_r101_c112 bl[112] br[112] wl[101] vdd gnd cell_6t
Xbit_r102_c112 bl[112] br[112] wl[102] vdd gnd cell_6t
Xbit_r103_c112 bl[112] br[112] wl[103] vdd gnd cell_6t
Xbit_r104_c112 bl[112] br[112] wl[104] vdd gnd cell_6t
Xbit_r105_c112 bl[112] br[112] wl[105] vdd gnd cell_6t
Xbit_r106_c112 bl[112] br[112] wl[106] vdd gnd cell_6t
Xbit_r107_c112 bl[112] br[112] wl[107] vdd gnd cell_6t
Xbit_r108_c112 bl[112] br[112] wl[108] vdd gnd cell_6t
Xbit_r109_c112 bl[112] br[112] wl[109] vdd gnd cell_6t
Xbit_r110_c112 bl[112] br[112] wl[110] vdd gnd cell_6t
Xbit_r111_c112 bl[112] br[112] wl[111] vdd gnd cell_6t
Xbit_r112_c112 bl[112] br[112] wl[112] vdd gnd cell_6t
Xbit_r113_c112 bl[112] br[112] wl[113] vdd gnd cell_6t
Xbit_r114_c112 bl[112] br[112] wl[114] vdd gnd cell_6t
Xbit_r115_c112 bl[112] br[112] wl[115] vdd gnd cell_6t
Xbit_r116_c112 bl[112] br[112] wl[116] vdd gnd cell_6t
Xbit_r117_c112 bl[112] br[112] wl[117] vdd gnd cell_6t
Xbit_r118_c112 bl[112] br[112] wl[118] vdd gnd cell_6t
Xbit_r119_c112 bl[112] br[112] wl[119] vdd gnd cell_6t
Xbit_r120_c112 bl[112] br[112] wl[120] vdd gnd cell_6t
Xbit_r121_c112 bl[112] br[112] wl[121] vdd gnd cell_6t
Xbit_r122_c112 bl[112] br[112] wl[122] vdd gnd cell_6t
Xbit_r123_c112 bl[112] br[112] wl[123] vdd gnd cell_6t
Xbit_r124_c112 bl[112] br[112] wl[124] vdd gnd cell_6t
Xbit_r125_c112 bl[112] br[112] wl[125] vdd gnd cell_6t
Xbit_r126_c112 bl[112] br[112] wl[126] vdd gnd cell_6t
Xbit_r127_c112 bl[112] br[112] wl[127] vdd gnd cell_6t
Xbit_r0_c113 bl[113] br[113] wl[0] vdd gnd cell_6t
Xbit_r1_c113 bl[113] br[113] wl[1] vdd gnd cell_6t
Xbit_r2_c113 bl[113] br[113] wl[2] vdd gnd cell_6t
Xbit_r3_c113 bl[113] br[113] wl[3] vdd gnd cell_6t
Xbit_r4_c113 bl[113] br[113] wl[4] vdd gnd cell_6t
Xbit_r5_c113 bl[113] br[113] wl[5] vdd gnd cell_6t
Xbit_r6_c113 bl[113] br[113] wl[6] vdd gnd cell_6t
Xbit_r7_c113 bl[113] br[113] wl[7] vdd gnd cell_6t
Xbit_r8_c113 bl[113] br[113] wl[8] vdd gnd cell_6t
Xbit_r9_c113 bl[113] br[113] wl[9] vdd gnd cell_6t
Xbit_r10_c113 bl[113] br[113] wl[10] vdd gnd cell_6t
Xbit_r11_c113 bl[113] br[113] wl[11] vdd gnd cell_6t
Xbit_r12_c113 bl[113] br[113] wl[12] vdd gnd cell_6t
Xbit_r13_c113 bl[113] br[113] wl[13] vdd gnd cell_6t
Xbit_r14_c113 bl[113] br[113] wl[14] vdd gnd cell_6t
Xbit_r15_c113 bl[113] br[113] wl[15] vdd gnd cell_6t
Xbit_r16_c113 bl[113] br[113] wl[16] vdd gnd cell_6t
Xbit_r17_c113 bl[113] br[113] wl[17] vdd gnd cell_6t
Xbit_r18_c113 bl[113] br[113] wl[18] vdd gnd cell_6t
Xbit_r19_c113 bl[113] br[113] wl[19] vdd gnd cell_6t
Xbit_r20_c113 bl[113] br[113] wl[20] vdd gnd cell_6t
Xbit_r21_c113 bl[113] br[113] wl[21] vdd gnd cell_6t
Xbit_r22_c113 bl[113] br[113] wl[22] vdd gnd cell_6t
Xbit_r23_c113 bl[113] br[113] wl[23] vdd gnd cell_6t
Xbit_r24_c113 bl[113] br[113] wl[24] vdd gnd cell_6t
Xbit_r25_c113 bl[113] br[113] wl[25] vdd gnd cell_6t
Xbit_r26_c113 bl[113] br[113] wl[26] vdd gnd cell_6t
Xbit_r27_c113 bl[113] br[113] wl[27] vdd gnd cell_6t
Xbit_r28_c113 bl[113] br[113] wl[28] vdd gnd cell_6t
Xbit_r29_c113 bl[113] br[113] wl[29] vdd gnd cell_6t
Xbit_r30_c113 bl[113] br[113] wl[30] vdd gnd cell_6t
Xbit_r31_c113 bl[113] br[113] wl[31] vdd gnd cell_6t
Xbit_r32_c113 bl[113] br[113] wl[32] vdd gnd cell_6t
Xbit_r33_c113 bl[113] br[113] wl[33] vdd gnd cell_6t
Xbit_r34_c113 bl[113] br[113] wl[34] vdd gnd cell_6t
Xbit_r35_c113 bl[113] br[113] wl[35] vdd gnd cell_6t
Xbit_r36_c113 bl[113] br[113] wl[36] vdd gnd cell_6t
Xbit_r37_c113 bl[113] br[113] wl[37] vdd gnd cell_6t
Xbit_r38_c113 bl[113] br[113] wl[38] vdd gnd cell_6t
Xbit_r39_c113 bl[113] br[113] wl[39] vdd gnd cell_6t
Xbit_r40_c113 bl[113] br[113] wl[40] vdd gnd cell_6t
Xbit_r41_c113 bl[113] br[113] wl[41] vdd gnd cell_6t
Xbit_r42_c113 bl[113] br[113] wl[42] vdd gnd cell_6t
Xbit_r43_c113 bl[113] br[113] wl[43] vdd gnd cell_6t
Xbit_r44_c113 bl[113] br[113] wl[44] vdd gnd cell_6t
Xbit_r45_c113 bl[113] br[113] wl[45] vdd gnd cell_6t
Xbit_r46_c113 bl[113] br[113] wl[46] vdd gnd cell_6t
Xbit_r47_c113 bl[113] br[113] wl[47] vdd gnd cell_6t
Xbit_r48_c113 bl[113] br[113] wl[48] vdd gnd cell_6t
Xbit_r49_c113 bl[113] br[113] wl[49] vdd gnd cell_6t
Xbit_r50_c113 bl[113] br[113] wl[50] vdd gnd cell_6t
Xbit_r51_c113 bl[113] br[113] wl[51] vdd gnd cell_6t
Xbit_r52_c113 bl[113] br[113] wl[52] vdd gnd cell_6t
Xbit_r53_c113 bl[113] br[113] wl[53] vdd gnd cell_6t
Xbit_r54_c113 bl[113] br[113] wl[54] vdd gnd cell_6t
Xbit_r55_c113 bl[113] br[113] wl[55] vdd gnd cell_6t
Xbit_r56_c113 bl[113] br[113] wl[56] vdd gnd cell_6t
Xbit_r57_c113 bl[113] br[113] wl[57] vdd gnd cell_6t
Xbit_r58_c113 bl[113] br[113] wl[58] vdd gnd cell_6t
Xbit_r59_c113 bl[113] br[113] wl[59] vdd gnd cell_6t
Xbit_r60_c113 bl[113] br[113] wl[60] vdd gnd cell_6t
Xbit_r61_c113 bl[113] br[113] wl[61] vdd gnd cell_6t
Xbit_r62_c113 bl[113] br[113] wl[62] vdd gnd cell_6t
Xbit_r63_c113 bl[113] br[113] wl[63] vdd gnd cell_6t
Xbit_r64_c113 bl[113] br[113] wl[64] vdd gnd cell_6t
Xbit_r65_c113 bl[113] br[113] wl[65] vdd gnd cell_6t
Xbit_r66_c113 bl[113] br[113] wl[66] vdd gnd cell_6t
Xbit_r67_c113 bl[113] br[113] wl[67] vdd gnd cell_6t
Xbit_r68_c113 bl[113] br[113] wl[68] vdd gnd cell_6t
Xbit_r69_c113 bl[113] br[113] wl[69] vdd gnd cell_6t
Xbit_r70_c113 bl[113] br[113] wl[70] vdd gnd cell_6t
Xbit_r71_c113 bl[113] br[113] wl[71] vdd gnd cell_6t
Xbit_r72_c113 bl[113] br[113] wl[72] vdd gnd cell_6t
Xbit_r73_c113 bl[113] br[113] wl[73] vdd gnd cell_6t
Xbit_r74_c113 bl[113] br[113] wl[74] vdd gnd cell_6t
Xbit_r75_c113 bl[113] br[113] wl[75] vdd gnd cell_6t
Xbit_r76_c113 bl[113] br[113] wl[76] vdd gnd cell_6t
Xbit_r77_c113 bl[113] br[113] wl[77] vdd gnd cell_6t
Xbit_r78_c113 bl[113] br[113] wl[78] vdd gnd cell_6t
Xbit_r79_c113 bl[113] br[113] wl[79] vdd gnd cell_6t
Xbit_r80_c113 bl[113] br[113] wl[80] vdd gnd cell_6t
Xbit_r81_c113 bl[113] br[113] wl[81] vdd gnd cell_6t
Xbit_r82_c113 bl[113] br[113] wl[82] vdd gnd cell_6t
Xbit_r83_c113 bl[113] br[113] wl[83] vdd gnd cell_6t
Xbit_r84_c113 bl[113] br[113] wl[84] vdd gnd cell_6t
Xbit_r85_c113 bl[113] br[113] wl[85] vdd gnd cell_6t
Xbit_r86_c113 bl[113] br[113] wl[86] vdd gnd cell_6t
Xbit_r87_c113 bl[113] br[113] wl[87] vdd gnd cell_6t
Xbit_r88_c113 bl[113] br[113] wl[88] vdd gnd cell_6t
Xbit_r89_c113 bl[113] br[113] wl[89] vdd gnd cell_6t
Xbit_r90_c113 bl[113] br[113] wl[90] vdd gnd cell_6t
Xbit_r91_c113 bl[113] br[113] wl[91] vdd gnd cell_6t
Xbit_r92_c113 bl[113] br[113] wl[92] vdd gnd cell_6t
Xbit_r93_c113 bl[113] br[113] wl[93] vdd gnd cell_6t
Xbit_r94_c113 bl[113] br[113] wl[94] vdd gnd cell_6t
Xbit_r95_c113 bl[113] br[113] wl[95] vdd gnd cell_6t
Xbit_r96_c113 bl[113] br[113] wl[96] vdd gnd cell_6t
Xbit_r97_c113 bl[113] br[113] wl[97] vdd gnd cell_6t
Xbit_r98_c113 bl[113] br[113] wl[98] vdd gnd cell_6t
Xbit_r99_c113 bl[113] br[113] wl[99] vdd gnd cell_6t
Xbit_r100_c113 bl[113] br[113] wl[100] vdd gnd cell_6t
Xbit_r101_c113 bl[113] br[113] wl[101] vdd gnd cell_6t
Xbit_r102_c113 bl[113] br[113] wl[102] vdd gnd cell_6t
Xbit_r103_c113 bl[113] br[113] wl[103] vdd gnd cell_6t
Xbit_r104_c113 bl[113] br[113] wl[104] vdd gnd cell_6t
Xbit_r105_c113 bl[113] br[113] wl[105] vdd gnd cell_6t
Xbit_r106_c113 bl[113] br[113] wl[106] vdd gnd cell_6t
Xbit_r107_c113 bl[113] br[113] wl[107] vdd gnd cell_6t
Xbit_r108_c113 bl[113] br[113] wl[108] vdd gnd cell_6t
Xbit_r109_c113 bl[113] br[113] wl[109] vdd gnd cell_6t
Xbit_r110_c113 bl[113] br[113] wl[110] vdd gnd cell_6t
Xbit_r111_c113 bl[113] br[113] wl[111] vdd gnd cell_6t
Xbit_r112_c113 bl[113] br[113] wl[112] vdd gnd cell_6t
Xbit_r113_c113 bl[113] br[113] wl[113] vdd gnd cell_6t
Xbit_r114_c113 bl[113] br[113] wl[114] vdd gnd cell_6t
Xbit_r115_c113 bl[113] br[113] wl[115] vdd gnd cell_6t
Xbit_r116_c113 bl[113] br[113] wl[116] vdd gnd cell_6t
Xbit_r117_c113 bl[113] br[113] wl[117] vdd gnd cell_6t
Xbit_r118_c113 bl[113] br[113] wl[118] vdd gnd cell_6t
Xbit_r119_c113 bl[113] br[113] wl[119] vdd gnd cell_6t
Xbit_r120_c113 bl[113] br[113] wl[120] vdd gnd cell_6t
Xbit_r121_c113 bl[113] br[113] wl[121] vdd gnd cell_6t
Xbit_r122_c113 bl[113] br[113] wl[122] vdd gnd cell_6t
Xbit_r123_c113 bl[113] br[113] wl[123] vdd gnd cell_6t
Xbit_r124_c113 bl[113] br[113] wl[124] vdd gnd cell_6t
Xbit_r125_c113 bl[113] br[113] wl[125] vdd gnd cell_6t
Xbit_r126_c113 bl[113] br[113] wl[126] vdd gnd cell_6t
Xbit_r127_c113 bl[113] br[113] wl[127] vdd gnd cell_6t
Xbit_r0_c114 bl[114] br[114] wl[0] vdd gnd cell_6t
Xbit_r1_c114 bl[114] br[114] wl[1] vdd gnd cell_6t
Xbit_r2_c114 bl[114] br[114] wl[2] vdd gnd cell_6t
Xbit_r3_c114 bl[114] br[114] wl[3] vdd gnd cell_6t
Xbit_r4_c114 bl[114] br[114] wl[4] vdd gnd cell_6t
Xbit_r5_c114 bl[114] br[114] wl[5] vdd gnd cell_6t
Xbit_r6_c114 bl[114] br[114] wl[6] vdd gnd cell_6t
Xbit_r7_c114 bl[114] br[114] wl[7] vdd gnd cell_6t
Xbit_r8_c114 bl[114] br[114] wl[8] vdd gnd cell_6t
Xbit_r9_c114 bl[114] br[114] wl[9] vdd gnd cell_6t
Xbit_r10_c114 bl[114] br[114] wl[10] vdd gnd cell_6t
Xbit_r11_c114 bl[114] br[114] wl[11] vdd gnd cell_6t
Xbit_r12_c114 bl[114] br[114] wl[12] vdd gnd cell_6t
Xbit_r13_c114 bl[114] br[114] wl[13] vdd gnd cell_6t
Xbit_r14_c114 bl[114] br[114] wl[14] vdd gnd cell_6t
Xbit_r15_c114 bl[114] br[114] wl[15] vdd gnd cell_6t
Xbit_r16_c114 bl[114] br[114] wl[16] vdd gnd cell_6t
Xbit_r17_c114 bl[114] br[114] wl[17] vdd gnd cell_6t
Xbit_r18_c114 bl[114] br[114] wl[18] vdd gnd cell_6t
Xbit_r19_c114 bl[114] br[114] wl[19] vdd gnd cell_6t
Xbit_r20_c114 bl[114] br[114] wl[20] vdd gnd cell_6t
Xbit_r21_c114 bl[114] br[114] wl[21] vdd gnd cell_6t
Xbit_r22_c114 bl[114] br[114] wl[22] vdd gnd cell_6t
Xbit_r23_c114 bl[114] br[114] wl[23] vdd gnd cell_6t
Xbit_r24_c114 bl[114] br[114] wl[24] vdd gnd cell_6t
Xbit_r25_c114 bl[114] br[114] wl[25] vdd gnd cell_6t
Xbit_r26_c114 bl[114] br[114] wl[26] vdd gnd cell_6t
Xbit_r27_c114 bl[114] br[114] wl[27] vdd gnd cell_6t
Xbit_r28_c114 bl[114] br[114] wl[28] vdd gnd cell_6t
Xbit_r29_c114 bl[114] br[114] wl[29] vdd gnd cell_6t
Xbit_r30_c114 bl[114] br[114] wl[30] vdd gnd cell_6t
Xbit_r31_c114 bl[114] br[114] wl[31] vdd gnd cell_6t
Xbit_r32_c114 bl[114] br[114] wl[32] vdd gnd cell_6t
Xbit_r33_c114 bl[114] br[114] wl[33] vdd gnd cell_6t
Xbit_r34_c114 bl[114] br[114] wl[34] vdd gnd cell_6t
Xbit_r35_c114 bl[114] br[114] wl[35] vdd gnd cell_6t
Xbit_r36_c114 bl[114] br[114] wl[36] vdd gnd cell_6t
Xbit_r37_c114 bl[114] br[114] wl[37] vdd gnd cell_6t
Xbit_r38_c114 bl[114] br[114] wl[38] vdd gnd cell_6t
Xbit_r39_c114 bl[114] br[114] wl[39] vdd gnd cell_6t
Xbit_r40_c114 bl[114] br[114] wl[40] vdd gnd cell_6t
Xbit_r41_c114 bl[114] br[114] wl[41] vdd gnd cell_6t
Xbit_r42_c114 bl[114] br[114] wl[42] vdd gnd cell_6t
Xbit_r43_c114 bl[114] br[114] wl[43] vdd gnd cell_6t
Xbit_r44_c114 bl[114] br[114] wl[44] vdd gnd cell_6t
Xbit_r45_c114 bl[114] br[114] wl[45] vdd gnd cell_6t
Xbit_r46_c114 bl[114] br[114] wl[46] vdd gnd cell_6t
Xbit_r47_c114 bl[114] br[114] wl[47] vdd gnd cell_6t
Xbit_r48_c114 bl[114] br[114] wl[48] vdd gnd cell_6t
Xbit_r49_c114 bl[114] br[114] wl[49] vdd gnd cell_6t
Xbit_r50_c114 bl[114] br[114] wl[50] vdd gnd cell_6t
Xbit_r51_c114 bl[114] br[114] wl[51] vdd gnd cell_6t
Xbit_r52_c114 bl[114] br[114] wl[52] vdd gnd cell_6t
Xbit_r53_c114 bl[114] br[114] wl[53] vdd gnd cell_6t
Xbit_r54_c114 bl[114] br[114] wl[54] vdd gnd cell_6t
Xbit_r55_c114 bl[114] br[114] wl[55] vdd gnd cell_6t
Xbit_r56_c114 bl[114] br[114] wl[56] vdd gnd cell_6t
Xbit_r57_c114 bl[114] br[114] wl[57] vdd gnd cell_6t
Xbit_r58_c114 bl[114] br[114] wl[58] vdd gnd cell_6t
Xbit_r59_c114 bl[114] br[114] wl[59] vdd gnd cell_6t
Xbit_r60_c114 bl[114] br[114] wl[60] vdd gnd cell_6t
Xbit_r61_c114 bl[114] br[114] wl[61] vdd gnd cell_6t
Xbit_r62_c114 bl[114] br[114] wl[62] vdd gnd cell_6t
Xbit_r63_c114 bl[114] br[114] wl[63] vdd gnd cell_6t
Xbit_r64_c114 bl[114] br[114] wl[64] vdd gnd cell_6t
Xbit_r65_c114 bl[114] br[114] wl[65] vdd gnd cell_6t
Xbit_r66_c114 bl[114] br[114] wl[66] vdd gnd cell_6t
Xbit_r67_c114 bl[114] br[114] wl[67] vdd gnd cell_6t
Xbit_r68_c114 bl[114] br[114] wl[68] vdd gnd cell_6t
Xbit_r69_c114 bl[114] br[114] wl[69] vdd gnd cell_6t
Xbit_r70_c114 bl[114] br[114] wl[70] vdd gnd cell_6t
Xbit_r71_c114 bl[114] br[114] wl[71] vdd gnd cell_6t
Xbit_r72_c114 bl[114] br[114] wl[72] vdd gnd cell_6t
Xbit_r73_c114 bl[114] br[114] wl[73] vdd gnd cell_6t
Xbit_r74_c114 bl[114] br[114] wl[74] vdd gnd cell_6t
Xbit_r75_c114 bl[114] br[114] wl[75] vdd gnd cell_6t
Xbit_r76_c114 bl[114] br[114] wl[76] vdd gnd cell_6t
Xbit_r77_c114 bl[114] br[114] wl[77] vdd gnd cell_6t
Xbit_r78_c114 bl[114] br[114] wl[78] vdd gnd cell_6t
Xbit_r79_c114 bl[114] br[114] wl[79] vdd gnd cell_6t
Xbit_r80_c114 bl[114] br[114] wl[80] vdd gnd cell_6t
Xbit_r81_c114 bl[114] br[114] wl[81] vdd gnd cell_6t
Xbit_r82_c114 bl[114] br[114] wl[82] vdd gnd cell_6t
Xbit_r83_c114 bl[114] br[114] wl[83] vdd gnd cell_6t
Xbit_r84_c114 bl[114] br[114] wl[84] vdd gnd cell_6t
Xbit_r85_c114 bl[114] br[114] wl[85] vdd gnd cell_6t
Xbit_r86_c114 bl[114] br[114] wl[86] vdd gnd cell_6t
Xbit_r87_c114 bl[114] br[114] wl[87] vdd gnd cell_6t
Xbit_r88_c114 bl[114] br[114] wl[88] vdd gnd cell_6t
Xbit_r89_c114 bl[114] br[114] wl[89] vdd gnd cell_6t
Xbit_r90_c114 bl[114] br[114] wl[90] vdd gnd cell_6t
Xbit_r91_c114 bl[114] br[114] wl[91] vdd gnd cell_6t
Xbit_r92_c114 bl[114] br[114] wl[92] vdd gnd cell_6t
Xbit_r93_c114 bl[114] br[114] wl[93] vdd gnd cell_6t
Xbit_r94_c114 bl[114] br[114] wl[94] vdd gnd cell_6t
Xbit_r95_c114 bl[114] br[114] wl[95] vdd gnd cell_6t
Xbit_r96_c114 bl[114] br[114] wl[96] vdd gnd cell_6t
Xbit_r97_c114 bl[114] br[114] wl[97] vdd gnd cell_6t
Xbit_r98_c114 bl[114] br[114] wl[98] vdd gnd cell_6t
Xbit_r99_c114 bl[114] br[114] wl[99] vdd gnd cell_6t
Xbit_r100_c114 bl[114] br[114] wl[100] vdd gnd cell_6t
Xbit_r101_c114 bl[114] br[114] wl[101] vdd gnd cell_6t
Xbit_r102_c114 bl[114] br[114] wl[102] vdd gnd cell_6t
Xbit_r103_c114 bl[114] br[114] wl[103] vdd gnd cell_6t
Xbit_r104_c114 bl[114] br[114] wl[104] vdd gnd cell_6t
Xbit_r105_c114 bl[114] br[114] wl[105] vdd gnd cell_6t
Xbit_r106_c114 bl[114] br[114] wl[106] vdd gnd cell_6t
Xbit_r107_c114 bl[114] br[114] wl[107] vdd gnd cell_6t
Xbit_r108_c114 bl[114] br[114] wl[108] vdd gnd cell_6t
Xbit_r109_c114 bl[114] br[114] wl[109] vdd gnd cell_6t
Xbit_r110_c114 bl[114] br[114] wl[110] vdd gnd cell_6t
Xbit_r111_c114 bl[114] br[114] wl[111] vdd gnd cell_6t
Xbit_r112_c114 bl[114] br[114] wl[112] vdd gnd cell_6t
Xbit_r113_c114 bl[114] br[114] wl[113] vdd gnd cell_6t
Xbit_r114_c114 bl[114] br[114] wl[114] vdd gnd cell_6t
Xbit_r115_c114 bl[114] br[114] wl[115] vdd gnd cell_6t
Xbit_r116_c114 bl[114] br[114] wl[116] vdd gnd cell_6t
Xbit_r117_c114 bl[114] br[114] wl[117] vdd gnd cell_6t
Xbit_r118_c114 bl[114] br[114] wl[118] vdd gnd cell_6t
Xbit_r119_c114 bl[114] br[114] wl[119] vdd gnd cell_6t
Xbit_r120_c114 bl[114] br[114] wl[120] vdd gnd cell_6t
Xbit_r121_c114 bl[114] br[114] wl[121] vdd gnd cell_6t
Xbit_r122_c114 bl[114] br[114] wl[122] vdd gnd cell_6t
Xbit_r123_c114 bl[114] br[114] wl[123] vdd gnd cell_6t
Xbit_r124_c114 bl[114] br[114] wl[124] vdd gnd cell_6t
Xbit_r125_c114 bl[114] br[114] wl[125] vdd gnd cell_6t
Xbit_r126_c114 bl[114] br[114] wl[126] vdd gnd cell_6t
Xbit_r127_c114 bl[114] br[114] wl[127] vdd gnd cell_6t
Xbit_r0_c115 bl[115] br[115] wl[0] vdd gnd cell_6t
Xbit_r1_c115 bl[115] br[115] wl[1] vdd gnd cell_6t
Xbit_r2_c115 bl[115] br[115] wl[2] vdd gnd cell_6t
Xbit_r3_c115 bl[115] br[115] wl[3] vdd gnd cell_6t
Xbit_r4_c115 bl[115] br[115] wl[4] vdd gnd cell_6t
Xbit_r5_c115 bl[115] br[115] wl[5] vdd gnd cell_6t
Xbit_r6_c115 bl[115] br[115] wl[6] vdd gnd cell_6t
Xbit_r7_c115 bl[115] br[115] wl[7] vdd gnd cell_6t
Xbit_r8_c115 bl[115] br[115] wl[8] vdd gnd cell_6t
Xbit_r9_c115 bl[115] br[115] wl[9] vdd gnd cell_6t
Xbit_r10_c115 bl[115] br[115] wl[10] vdd gnd cell_6t
Xbit_r11_c115 bl[115] br[115] wl[11] vdd gnd cell_6t
Xbit_r12_c115 bl[115] br[115] wl[12] vdd gnd cell_6t
Xbit_r13_c115 bl[115] br[115] wl[13] vdd gnd cell_6t
Xbit_r14_c115 bl[115] br[115] wl[14] vdd gnd cell_6t
Xbit_r15_c115 bl[115] br[115] wl[15] vdd gnd cell_6t
Xbit_r16_c115 bl[115] br[115] wl[16] vdd gnd cell_6t
Xbit_r17_c115 bl[115] br[115] wl[17] vdd gnd cell_6t
Xbit_r18_c115 bl[115] br[115] wl[18] vdd gnd cell_6t
Xbit_r19_c115 bl[115] br[115] wl[19] vdd gnd cell_6t
Xbit_r20_c115 bl[115] br[115] wl[20] vdd gnd cell_6t
Xbit_r21_c115 bl[115] br[115] wl[21] vdd gnd cell_6t
Xbit_r22_c115 bl[115] br[115] wl[22] vdd gnd cell_6t
Xbit_r23_c115 bl[115] br[115] wl[23] vdd gnd cell_6t
Xbit_r24_c115 bl[115] br[115] wl[24] vdd gnd cell_6t
Xbit_r25_c115 bl[115] br[115] wl[25] vdd gnd cell_6t
Xbit_r26_c115 bl[115] br[115] wl[26] vdd gnd cell_6t
Xbit_r27_c115 bl[115] br[115] wl[27] vdd gnd cell_6t
Xbit_r28_c115 bl[115] br[115] wl[28] vdd gnd cell_6t
Xbit_r29_c115 bl[115] br[115] wl[29] vdd gnd cell_6t
Xbit_r30_c115 bl[115] br[115] wl[30] vdd gnd cell_6t
Xbit_r31_c115 bl[115] br[115] wl[31] vdd gnd cell_6t
Xbit_r32_c115 bl[115] br[115] wl[32] vdd gnd cell_6t
Xbit_r33_c115 bl[115] br[115] wl[33] vdd gnd cell_6t
Xbit_r34_c115 bl[115] br[115] wl[34] vdd gnd cell_6t
Xbit_r35_c115 bl[115] br[115] wl[35] vdd gnd cell_6t
Xbit_r36_c115 bl[115] br[115] wl[36] vdd gnd cell_6t
Xbit_r37_c115 bl[115] br[115] wl[37] vdd gnd cell_6t
Xbit_r38_c115 bl[115] br[115] wl[38] vdd gnd cell_6t
Xbit_r39_c115 bl[115] br[115] wl[39] vdd gnd cell_6t
Xbit_r40_c115 bl[115] br[115] wl[40] vdd gnd cell_6t
Xbit_r41_c115 bl[115] br[115] wl[41] vdd gnd cell_6t
Xbit_r42_c115 bl[115] br[115] wl[42] vdd gnd cell_6t
Xbit_r43_c115 bl[115] br[115] wl[43] vdd gnd cell_6t
Xbit_r44_c115 bl[115] br[115] wl[44] vdd gnd cell_6t
Xbit_r45_c115 bl[115] br[115] wl[45] vdd gnd cell_6t
Xbit_r46_c115 bl[115] br[115] wl[46] vdd gnd cell_6t
Xbit_r47_c115 bl[115] br[115] wl[47] vdd gnd cell_6t
Xbit_r48_c115 bl[115] br[115] wl[48] vdd gnd cell_6t
Xbit_r49_c115 bl[115] br[115] wl[49] vdd gnd cell_6t
Xbit_r50_c115 bl[115] br[115] wl[50] vdd gnd cell_6t
Xbit_r51_c115 bl[115] br[115] wl[51] vdd gnd cell_6t
Xbit_r52_c115 bl[115] br[115] wl[52] vdd gnd cell_6t
Xbit_r53_c115 bl[115] br[115] wl[53] vdd gnd cell_6t
Xbit_r54_c115 bl[115] br[115] wl[54] vdd gnd cell_6t
Xbit_r55_c115 bl[115] br[115] wl[55] vdd gnd cell_6t
Xbit_r56_c115 bl[115] br[115] wl[56] vdd gnd cell_6t
Xbit_r57_c115 bl[115] br[115] wl[57] vdd gnd cell_6t
Xbit_r58_c115 bl[115] br[115] wl[58] vdd gnd cell_6t
Xbit_r59_c115 bl[115] br[115] wl[59] vdd gnd cell_6t
Xbit_r60_c115 bl[115] br[115] wl[60] vdd gnd cell_6t
Xbit_r61_c115 bl[115] br[115] wl[61] vdd gnd cell_6t
Xbit_r62_c115 bl[115] br[115] wl[62] vdd gnd cell_6t
Xbit_r63_c115 bl[115] br[115] wl[63] vdd gnd cell_6t
Xbit_r64_c115 bl[115] br[115] wl[64] vdd gnd cell_6t
Xbit_r65_c115 bl[115] br[115] wl[65] vdd gnd cell_6t
Xbit_r66_c115 bl[115] br[115] wl[66] vdd gnd cell_6t
Xbit_r67_c115 bl[115] br[115] wl[67] vdd gnd cell_6t
Xbit_r68_c115 bl[115] br[115] wl[68] vdd gnd cell_6t
Xbit_r69_c115 bl[115] br[115] wl[69] vdd gnd cell_6t
Xbit_r70_c115 bl[115] br[115] wl[70] vdd gnd cell_6t
Xbit_r71_c115 bl[115] br[115] wl[71] vdd gnd cell_6t
Xbit_r72_c115 bl[115] br[115] wl[72] vdd gnd cell_6t
Xbit_r73_c115 bl[115] br[115] wl[73] vdd gnd cell_6t
Xbit_r74_c115 bl[115] br[115] wl[74] vdd gnd cell_6t
Xbit_r75_c115 bl[115] br[115] wl[75] vdd gnd cell_6t
Xbit_r76_c115 bl[115] br[115] wl[76] vdd gnd cell_6t
Xbit_r77_c115 bl[115] br[115] wl[77] vdd gnd cell_6t
Xbit_r78_c115 bl[115] br[115] wl[78] vdd gnd cell_6t
Xbit_r79_c115 bl[115] br[115] wl[79] vdd gnd cell_6t
Xbit_r80_c115 bl[115] br[115] wl[80] vdd gnd cell_6t
Xbit_r81_c115 bl[115] br[115] wl[81] vdd gnd cell_6t
Xbit_r82_c115 bl[115] br[115] wl[82] vdd gnd cell_6t
Xbit_r83_c115 bl[115] br[115] wl[83] vdd gnd cell_6t
Xbit_r84_c115 bl[115] br[115] wl[84] vdd gnd cell_6t
Xbit_r85_c115 bl[115] br[115] wl[85] vdd gnd cell_6t
Xbit_r86_c115 bl[115] br[115] wl[86] vdd gnd cell_6t
Xbit_r87_c115 bl[115] br[115] wl[87] vdd gnd cell_6t
Xbit_r88_c115 bl[115] br[115] wl[88] vdd gnd cell_6t
Xbit_r89_c115 bl[115] br[115] wl[89] vdd gnd cell_6t
Xbit_r90_c115 bl[115] br[115] wl[90] vdd gnd cell_6t
Xbit_r91_c115 bl[115] br[115] wl[91] vdd gnd cell_6t
Xbit_r92_c115 bl[115] br[115] wl[92] vdd gnd cell_6t
Xbit_r93_c115 bl[115] br[115] wl[93] vdd gnd cell_6t
Xbit_r94_c115 bl[115] br[115] wl[94] vdd gnd cell_6t
Xbit_r95_c115 bl[115] br[115] wl[95] vdd gnd cell_6t
Xbit_r96_c115 bl[115] br[115] wl[96] vdd gnd cell_6t
Xbit_r97_c115 bl[115] br[115] wl[97] vdd gnd cell_6t
Xbit_r98_c115 bl[115] br[115] wl[98] vdd gnd cell_6t
Xbit_r99_c115 bl[115] br[115] wl[99] vdd gnd cell_6t
Xbit_r100_c115 bl[115] br[115] wl[100] vdd gnd cell_6t
Xbit_r101_c115 bl[115] br[115] wl[101] vdd gnd cell_6t
Xbit_r102_c115 bl[115] br[115] wl[102] vdd gnd cell_6t
Xbit_r103_c115 bl[115] br[115] wl[103] vdd gnd cell_6t
Xbit_r104_c115 bl[115] br[115] wl[104] vdd gnd cell_6t
Xbit_r105_c115 bl[115] br[115] wl[105] vdd gnd cell_6t
Xbit_r106_c115 bl[115] br[115] wl[106] vdd gnd cell_6t
Xbit_r107_c115 bl[115] br[115] wl[107] vdd gnd cell_6t
Xbit_r108_c115 bl[115] br[115] wl[108] vdd gnd cell_6t
Xbit_r109_c115 bl[115] br[115] wl[109] vdd gnd cell_6t
Xbit_r110_c115 bl[115] br[115] wl[110] vdd gnd cell_6t
Xbit_r111_c115 bl[115] br[115] wl[111] vdd gnd cell_6t
Xbit_r112_c115 bl[115] br[115] wl[112] vdd gnd cell_6t
Xbit_r113_c115 bl[115] br[115] wl[113] vdd gnd cell_6t
Xbit_r114_c115 bl[115] br[115] wl[114] vdd gnd cell_6t
Xbit_r115_c115 bl[115] br[115] wl[115] vdd gnd cell_6t
Xbit_r116_c115 bl[115] br[115] wl[116] vdd gnd cell_6t
Xbit_r117_c115 bl[115] br[115] wl[117] vdd gnd cell_6t
Xbit_r118_c115 bl[115] br[115] wl[118] vdd gnd cell_6t
Xbit_r119_c115 bl[115] br[115] wl[119] vdd gnd cell_6t
Xbit_r120_c115 bl[115] br[115] wl[120] vdd gnd cell_6t
Xbit_r121_c115 bl[115] br[115] wl[121] vdd gnd cell_6t
Xbit_r122_c115 bl[115] br[115] wl[122] vdd gnd cell_6t
Xbit_r123_c115 bl[115] br[115] wl[123] vdd gnd cell_6t
Xbit_r124_c115 bl[115] br[115] wl[124] vdd gnd cell_6t
Xbit_r125_c115 bl[115] br[115] wl[125] vdd gnd cell_6t
Xbit_r126_c115 bl[115] br[115] wl[126] vdd gnd cell_6t
Xbit_r127_c115 bl[115] br[115] wl[127] vdd gnd cell_6t
Xbit_r0_c116 bl[116] br[116] wl[0] vdd gnd cell_6t
Xbit_r1_c116 bl[116] br[116] wl[1] vdd gnd cell_6t
Xbit_r2_c116 bl[116] br[116] wl[2] vdd gnd cell_6t
Xbit_r3_c116 bl[116] br[116] wl[3] vdd gnd cell_6t
Xbit_r4_c116 bl[116] br[116] wl[4] vdd gnd cell_6t
Xbit_r5_c116 bl[116] br[116] wl[5] vdd gnd cell_6t
Xbit_r6_c116 bl[116] br[116] wl[6] vdd gnd cell_6t
Xbit_r7_c116 bl[116] br[116] wl[7] vdd gnd cell_6t
Xbit_r8_c116 bl[116] br[116] wl[8] vdd gnd cell_6t
Xbit_r9_c116 bl[116] br[116] wl[9] vdd gnd cell_6t
Xbit_r10_c116 bl[116] br[116] wl[10] vdd gnd cell_6t
Xbit_r11_c116 bl[116] br[116] wl[11] vdd gnd cell_6t
Xbit_r12_c116 bl[116] br[116] wl[12] vdd gnd cell_6t
Xbit_r13_c116 bl[116] br[116] wl[13] vdd gnd cell_6t
Xbit_r14_c116 bl[116] br[116] wl[14] vdd gnd cell_6t
Xbit_r15_c116 bl[116] br[116] wl[15] vdd gnd cell_6t
Xbit_r16_c116 bl[116] br[116] wl[16] vdd gnd cell_6t
Xbit_r17_c116 bl[116] br[116] wl[17] vdd gnd cell_6t
Xbit_r18_c116 bl[116] br[116] wl[18] vdd gnd cell_6t
Xbit_r19_c116 bl[116] br[116] wl[19] vdd gnd cell_6t
Xbit_r20_c116 bl[116] br[116] wl[20] vdd gnd cell_6t
Xbit_r21_c116 bl[116] br[116] wl[21] vdd gnd cell_6t
Xbit_r22_c116 bl[116] br[116] wl[22] vdd gnd cell_6t
Xbit_r23_c116 bl[116] br[116] wl[23] vdd gnd cell_6t
Xbit_r24_c116 bl[116] br[116] wl[24] vdd gnd cell_6t
Xbit_r25_c116 bl[116] br[116] wl[25] vdd gnd cell_6t
Xbit_r26_c116 bl[116] br[116] wl[26] vdd gnd cell_6t
Xbit_r27_c116 bl[116] br[116] wl[27] vdd gnd cell_6t
Xbit_r28_c116 bl[116] br[116] wl[28] vdd gnd cell_6t
Xbit_r29_c116 bl[116] br[116] wl[29] vdd gnd cell_6t
Xbit_r30_c116 bl[116] br[116] wl[30] vdd gnd cell_6t
Xbit_r31_c116 bl[116] br[116] wl[31] vdd gnd cell_6t
Xbit_r32_c116 bl[116] br[116] wl[32] vdd gnd cell_6t
Xbit_r33_c116 bl[116] br[116] wl[33] vdd gnd cell_6t
Xbit_r34_c116 bl[116] br[116] wl[34] vdd gnd cell_6t
Xbit_r35_c116 bl[116] br[116] wl[35] vdd gnd cell_6t
Xbit_r36_c116 bl[116] br[116] wl[36] vdd gnd cell_6t
Xbit_r37_c116 bl[116] br[116] wl[37] vdd gnd cell_6t
Xbit_r38_c116 bl[116] br[116] wl[38] vdd gnd cell_6t
Xbit_r39_c116 bl[116] br[116] wl[39] vdd gnd cell_6t
Xbit_r40_c116 bl[116] br[116] wl[40] vdd gnd cell_6t
Xbit_r41_c116 bl[116] br[116] wl[41] vdd gnd cell_6t
Xbit_r42_c116 bl[116] br[116] wl[42] vdd gnd cell_6t
Xbit_r43_c116 bl[116] br[116] wl[43] vdd gnd cell_6t
Xbit_r44_c116 bl[116] br[116] wl[44] vdd gnd cell_6t
Xbit_r45_c116 bl[116] br[116] wl[45] vdd gnd cell_6t
Xbit_r46_c116 bl[116] br[116] wl[46] vdd gnd cell_6t
Xbit_r47_c116 bl[116] br[116] wl[47] vdd gnd cell_6t
Xbit_r48_c116 bl[116] br[116] wl[48] vdd gnd cell_6t
Xbit_r49_c116 bl[116] br[116] wl[49] vdd gnd cell_6t
Xbit_r50_c116 bl[116] br[116] wl[50] vdd gnd cell_6t
Xbit_r51_c116 bl[116] br[116] wl[51] vdd gnd cell_6t
Xbit_r52_c116 bl[116] br[116] wl[52] vdd gnd cell_6t
Xbit_r53_c116 bl[116] br[116] wl[53] vdd gnd cell_6t
Xbit_r54_c116 bl[116] br[116] wl[54] vdd gnd cell_6t
Xbit_r55_c116 bl[116] br[116] wl[55] vdd gnd cell_6t
Xbit_r56_c116 bl[116] br[116] wl[56] vdd gnd cell_6t
Xbit_r57_c116 bl[116] br[116] wl[57] vdd gnd cell_6t
Xbit_r58_c116 bl[116] br[116] wl[58] vdd gnd cell_6t
Xbit_r59_c116 bl[116] br[116] wl[59] vdd gnd cell_6t
Xbit_r60_c116 bl[116] br[116] wl[60] vdd gnd cell_6t
Xbit_r61_c116 bl[116] br[116] wl[61] vdd gnd cell_6t
Xbit_r62_c116 bl[116] br[116] wl[62] vdd gnd cell_6t
Xbit_r63_c116 bl[116] br[116] wl[63] vdd gnd cell_6t
Xbit_r64_c116 bl[116] br[116] wl[64] vdd gnd cell_6t
Xbit_r65_c116 bl[116] br[116] wl[65] vdd gnd cell_6t
Xbit_r66_c116 bl[116] br[116] wl[66] vdd gnd cell_6t
Xbit_r67_c116 bl[116] br[116] wl[67] vdd gnd cell_6t
Xbit_r68_c116 bl[116] br[116] wl[68] vdd gnd cell_6t
Xbit_r69_c116 bl[116] br[116] wl[69] vdd gnd cell_6t
Xbit_r70_c116 bl[116] br[116] wl[70] vdd gnd cell_6t
Xbit_r71_c116 bl[116] br[116] wl[71] vdd gnd cell_6t
Xbit_r72_c116 bl[116] br[116] wl[72] vdd gnd cell_6t
Xbit_r73_c116 bl[116] br[116] wl[73] vdd gnd cell_6t
Xbit_r74_c116 bl[116] br[116] wl[74] vdd gnd cell_6t
Xbit_r75_c116 bl[116] br[116] wl[75] vdd gnd cell_6t
Xbit_r76_c116 bl[116] br[116] wl[76] vdd gnd cell_6t
Xbit_r77_c116 bl[116] br[116] wl[77] vdd gnd cell_6t
Xbit_r78_c116 bl[116] br[116] wl[78] vdd gnd cell_6t
Xbit_r79_c116 bl[116] br[116] wl[79] vdd gnd cell_6t
Xbit_r80_c116 bl[116] br[116] wl[80] vdd gnd cell_6t
Xbit_r81_c116 bl[116] br[116] wl[81] vdd gnd cell_6t
Xbit_r82_c116 bl[116] br[116] wl[82] vdd gnd cell_6t
Xbit_r83_c116 bl[116] br[116] wl[83] vdd gnd cell_6t
Xbit_r84_c116 bl[116] br[116] wl[84] vdd gnd cell_6t
Xbit_r85_c116 bl[116] br[116] wl[85] vdd gnd cell_6t
Xbit_r86_c116 bl[116] br[116] wl[86] vdd gnd cell_6t
Xbit_r87_c116 bl[116] br[116] wl[87] vdd gnd cell_6t
Xbit_r88_c116 bl[116] br[116] wl[88] vdd gnd cell_6t
Xbit_r89_c116 bl[116] br[116] wl[89] vdd gnd cell_6t
Xbit_r90_c116 bl[116] br[116] wl[90] vdd gnd cell_6t
Xbit_r91_c116 bl[116] br[116] wl[91] vdd gnd cell_6t
Xbit_r92_c116 bl[116] br[116] wl[92] vdd gnd cell_6t
Xbit_r93_c116 bl[116] br[116] wl[93] vdd gnd cell_6t
Xbit_r94_c116 bl[116] br[116] wl[94] vdd gnd cell_6t
Xbit_r95_c116 bl[116] br[116] wl[95] vdd gnd cell_6t
Xbit_r96_c116 bl[116] br[116] wl[96] vdd gnd cell_6t
Xbit_r97_c116 bl[116] br[116] wl[97] vdd gnd cell_6t
Xbit_r98_c116 bl[116] br[116] wl[98] vdd gnd cell_6t
Xbit_r99_c116 bl[116] br[116] wl[99] vdd gnd cell_6t
Xbit_r100_c116 bl[116] br[116] wl[100] vdd gnd cell_6t
Xbit_r101_c116 bl[116] br[116] wl[101] vdd gnd cell_6t
Xbit_r102_c116 bl[116] br[116] wl[102] vdd gnd cell_6t
Xbit_r103_c116 bl[116] br[116] wl[103] vdd gnd cell_6t
Xbit_r104_c116 bl[116] br[116] wl[104] vdd gnd cell_6t
Xbit_r105_c116 bl[116] br[116] wl[105] vdd gnd cell_6t
Xbit_r106_c116 bl[116] br[116] wl[106] vdd gnd cell_6t
Xbit_r107_c116 bl[116] br[116] wl[107] vdd gnd cell_6t
Xbit_r108_c116 bl[116] br[116] wl[108] vdd gnd cell_6t
Xbit_r109_c116 bl[116] br[116] wl[109] vdd gnd cell_6t
Xbit_r110_c116 bl[116] br[116] wl[110] vdd gnd cell_6t
Xbit_r111_c116 bl[116] br[116] wl[111] vdd gnd cell_6t
Xbit_r112_c116 bl[116] br[116] wl[112] vdd gnd cell_6t
Xbit_r113_c116 bl[116] br[116] wl[113] vdd gnd cell_6t
Xbit_r114_c116 bl[116] br[116] wl[114] vdd gnd cell_6t
Xbit_r115_c116 bl[116] br[116] wl[115] vdd gnd cell_6t
Xbit_r116_c116 bl[116] br[116] wl[116] vdd gnd cell_6t
Xbit_r117_c116 bl[116] br[116] wl[117] vdd gnd cell_6t
Xbit_r118_c116 bl[116] br[116] wl[118] vdd gnd cell_6t
Xbit_r119_c116 bl[116] br[116] wl[119] vdd gnd cell_6t
Xbit_r120_c116 bl[116] br[116] wl[120] vdd gnd cell_6t
Xbit_r121_c116 bl[116] br[116] wl[121] vdd gnd cell_6t
Xbit_r122_c116 bl[116] br[116] wl[122] vdd gnd cell_6t
Xbit_r123_c116 bl[116] br[116] wl[123] vdd gnd cell_6t
Xbit_r124_c116 bl[116] br[116] wl[124] vdd gnd cell_6t
Xbit_r125_c116 bl[116] br[116] wl[125] vdd gnd cell_6t
Xbit_r126_c116 bl[116] br[116] wl[126] vdd gnd cell_6t
Xbit_r127_c116 bl[116] br[116] wl[127] vdd gnd cell_6t
Xbit_r0_c117 bl[117] br[117] wl[0] vdd gnd cell_6t
Xbit_r1_c117 bl[117] br[117] wl[1] vdd gnd cell_6t
Xbit_r2_c117 bl[117] br[117] wl[2] vdd gnd cell_6t
Xbit_r3_c117 bl[117] br[117] wl[3] vdd gnd cell_6t
Xbit_r4_c117 bl[117] br[117] wl[4] vdd gnd cell_6t
Xbit_r5_c117 bl[117] br[117] wl[5] vdd gnd cell_6t
Xbit_r6_c117 bl[117] br[117] wl[6] vdd gnd cell_6t
Xbit_r7_c117 bl[117] br[117] wl[7] vdd gnd cell_6t
Xbit_r8_c117 bl[117] br[117] wl[8] vdd gnd cell_6t
Xbit_r9_c117 bl[117] br[117] wl[9] vdd gnd cell_6t
Xbit_r10_c117 bl[117] br[117] wl[10] vdd gnd cell_6t
Xbit_r11_c117 bl[117] br[117] wl[11] vdd gnd cell_6t
Xbit_r12_c117 bl[117] br[117] wl[12] vdd gnd cell_6t
Xbit_r13_c117 bl[117] br[117] wl[13] vdd gnd cell_6t
Xbit_r14_c117 bl[117] br[117] wl[14] vdd gnd cell_6t
Xbit_r15_c117 bl[117] br[117] wl[15] vdd gnd cell_6t
Xbit_r16_c117 bl[117] br[117] wl[16] vdd gnd cell_6t
Xbit_r17_c117 bl[117] br[117] wl[17] vdd gnd cell_6t
Xbit_r18_c117 bl[117] br[117] wl[18] vdd gnd cell_6t
Xbit_r19_c117 bl[117] br[117] wl[19] vdd gnd cell_6t
Xbit_r20_c117 bl[117] br[117] wl[20] vdd gnd cell_6t
Xbit_r21_c117 bl[117] br[117] wl[21] vdd gnd cell_6t
Xbit_r22_c117 bl[117] br[117] wl[22] vdd gnd cell_6t
Xbit_r23_c117 bl[117] br[117] wl[23] vdd gnd cell_6t
Xbit_r24_c117 bl[117] br[117] wl[24] vdd gnd cell_6t
Xbit_r25_c117 bl[117] br[117] wl[25] vdd gnd cell_6t
Xbit_r26_c117 bl[117] br[117] wl[26] vdd gnd cell_6t
Xbit_r27_c117 bl[117] br[117] wl[27] vdd gnd cell_6t
Xbit_r28_c117 bl[117] br[117] wl[28] vdd gnd cell_6t
Xbit_r29_c117 bl[117] br[117] wl[29] vdd gnd cell_6t
Xbit_r30_c117 bl[117] br[117] wl[30] vdd gnd cell_6t
Xbit_r31_c117 bl[117] br[117] wl[31] vdd gnd cell_6t
Xbit_r32_c117 bl[117] br[117] wl[32] vdd gnd cell_6t
Xbit_r33_c117 bl[117] br[117] wl[33] vdd gnd cell_6t
Xbit_r34_c117 bl[117] br[117] wl[34] vdd gnd cell_6t
Xbit_r35_c117 bl[117] br[117] wl[35] vdd gnd cell_6t
Xbit_r36_c117 bl[117] br[117] wl[36] vdd gnd cell_6t
Xbit_r37_c117 bl[117] br[117] wl[37] vdd gnd cell_6t
Xbit_r38_c117 bl[117] br[117] wl[38] vdd gnd cell_6t
Xbit_r39_c117 bl[117] br[117] wl[39] vdd gnd cell_6t
Xbit_r40_c117 bl[117] br[117] wl[40] vdd gnd cell_6t
Xbit_r41_c117 bl[117] br[117] wl[41] vdd gnd cell_6t
Xbit_r42_c117 bl[117] br[117] wl[42] vdd gnd cell_6t
Xbit_r43_c117 bl[117] br[117] wl[43] vdd gnd cell_6t
Xbit_r44_c117 bl[117] br[117] wl[44] vdd gnd cell_6t
Xbit_r45_c117 bl[117] br[117] wl[45] vdd gnd cell_6t
Xbit_r46_c117 bl[117] br[117] wl[46] vdd gnd cell_6t
Xbit_r47_c117 bl[117] br[117] wl[47] vdd gnd cell_6t
Xbit_r48_c117 bl[117] br[117] wl[48] vdd gnd cell_6t
Xbit_r49_c117 bl[117] br[117] wl[49] vdd gnd cell_6t
Xbit_r50_c117 bl[117] br[117] wl[50] vdd gnd cell_6t
Xbit_r51_c117 bl[117] br[117] wl[51] vdd gnd cell_6t
Xbit_r52_c117 bl[117] br[117] wl[52] vdd gnd cell_6t
Xbit_r53_c117 bl[117] br[117] wl[53] vdd gnd cell_6t
Xbit_r54_c117 bl[117] br[117] wl[54] vdd gnd cell_6t
Xbit_r55_c117 bl[117] br[117] wl[55] vdd gnd cell_6t
Xbit_r56_c117 bl[117] br[117] wl[56] vdd gnd cell_6t
Xbit_r57_c117 bl[117] br[117] wl[57] vdd gnd cell_6t
Xbit_r58_c117 bl[117] br[117] wl[58] vdd gnd cell_6t
Xbit_r59_c117 bl[117] br[117] wl[59] vdd gnd cell_6t
Xbit_r60_c117 bl[117] br[117] wl[60] vdd gnd cell_6t
Xbit_r61_c117 bl[117] br[117] wl[61] vdd gnd cell_6t
Xbit_r62_c117 bl[117] br[117] wl[62] vdd gnd cell_6t
Xbit_r63_c117 bl[117] br[117] wl[63] vdd gnd cell_6t
Xbit_r64_c117 bl[117] br[117] wl[64] vdd gnd cell_6t
Xbit_r65_c117 bl[117] br[117] wl[65] vdd gnd cell_6t
Xbit_r66_c117 bl[117] br[117] wl[66] vdd gnd cell_6t
Xbit_r67_c117 bl[117] br[117] wl[67] vdd gnd cell_6t
Xbit_r68_c117 bl[117] br[117] wl[68] vdd gnd cell_6t
Xbit_r69_c117 bl[117] br[117] wl[69] vdd gnd cell_6t
Xbit_r70_c117 bl[117] br[117] wl[70] vdd gnd cell_6t
Xbit_r71_c117 bl[117] br[117] wl[71] vdd gnd cell_6t
Xbit_r72_c117 bl[117] br[117] wl[72] vdd gnd cell_6t
Xbit_r73_c117 bl[117] br[117] wl[73] vdd gnd cell_6t
Xbit_r74_c117 bl[117] br[117] wl[74] vdd gnd cell_6t
Xbit_r75_c117 bl[117] br[117] wl[75] vdd gnd cell_6t
Xbit_r76_c117 bl[117] br[117] wl[76] vdd gnd cell_6t
Xbit_r77_c117 bl[117] br[117] wl[77] vdd gnd cell_6t
Xbit_r78_c117 bl[117] br[117] wl[78] vdd gnd cell_6t
Xbit_r79_c117 bl[117] br[117] wl[79] vdd gnd cell_6t
Xbit_r80_c117 bl[117] br[117] wl[80] vdd gnd cell_6t
Xbit_r81_c117 bl[117] br[117] wl[81] vdd gnd cell_6t
Xbit_r82_c117 bl[117] br[117] wl[82] vdd gnd cell_6t
Xbit_r83_c117 bl[117] br[117] wl[83] vdd gnd cell_6t
Xbit_r84_c117 bl[117] br[117] wl[84] vdd gnd cell_6t
Xbit_r85_c117 bl[117] br[117] wl[85] vdd gnd cell_6t
Xbit_r86_c117 bl[117] br[117] wl[86] vdd gnd cell_6t
Xbit_r87_c117 bl[117] br[117] wl[87] vdd gnd cell_6t
Xbit_r88_c117 bl[117] br[117] wl[88] vdd gnd cell_6t
Xbit_r89_c117 bl[117] br[117] wl[89] vdd gnd cell_6t
Xbit_r90_c117 bl[117] br[117] wl[90] vdd gnd cell_6t
Xbit_r91_c117 bl[117] br[117] wl[91] vdd gnd cell_6t
Xbit_r92_c117 bl[117] br[117] wl[92] vdd gnd cell_6t
Xbit_r93_c117 bl[117] br[117] wl[93] vdd gnd cell_6t
Xbit_r94_c117 bl[117] br[117] wl[94] vdd gnd cell_6t
Xbit_r95_c117 bl[117] br[117] wl[95] vdd gnd cell_6t
Xbit_r96_c117 bl[117] br[117] wl[96] vdd gnd cell_6t
Xbit_r97_c117 bl[117] br[117] wl[97] vdd gnd cell_6t
Xbit_r98_c117 bl[117] br[117] wl[98] vdd gnd cell_6t
Xbit_r99_c117 bl[117] br[117] wl[99] vdd gnd cell_6t
Xbit_r100_c117 bl[117] br[117] wl[100] vdd gnd cell_6t
Xbit_r101_c117 bl[117] br[117] wl[101] vdd gnd cell_6t
Xbit_r102_c117 bl[117] br[117] wl[102] vdd gnd cell_6t
Xbit_r103_c117 bl[117] br[117] wl[103] vdd gnd cell_6t
Xbit_r104_c117 bl[117] br[117] wl[104] vdd gnd cell_6t
Xbit_r105_c117 bl[117] br[117] wl[105] vdd gnd cell_6t
Xbit_r106_c117 bl[117] br[117] wl[106] vdd gnd cell_6t
Xbit_r107_c117 bl[117] br[117] wl[107] vdd gnd cell_6t
Xbit_r108_c117 bl[117] br[117] wl[108] vdd gnd cell_6t
Xbit_r109_c117 bl[117] br[117] wl[109] vdd gnd cell_6t
Xbit_r110_c117 bl[117] br[117] wl[110] vdd gnd cell_6t
Xbit_r111_c117 bl[117] br[117] wl[111] vdd gnd cell_6t
Xbit_r112_c117 bl[117] br[117] wl[112] vdd gnd cell_6t
Xbit_r113_c117 bl[117] br[117] wl[113] vdd gnd cell_6t
Xbit_r114_c117 bl[117] br[117] wl[114] vdd gnd cell_6t
Xbit_r115_c117 bl[117] br[117] wl[115] vdd gnd cell_6t
Xbit_r116_c117 bl[117] br[117] wl[116] vdd gnd cell_6t
Xbit_r117_c117 bl[117] br[117] wl[117] vdd gnd cell_6t
Xbit_r118_c117 bl[117] br[117] wl[118] vdd gnd cell_6t
Xbit_r119_c117 bl[117] br[117] wl[119] vdd gnd cell_6t
Xbit_r120_c117 bl[117] br[117] wl[120] vdd gnd cell_6t
Xbit_r121_c117 bl[117] br[117] wl[121] vdd gnd cell_6t
Xbit_r122_c117 bl[117] br[117] wl[122] vdd gnd cell_6t
Xbit_r123_c117 bl[117] br[117] wl[123] vdd gnd cell_6t
Xbit_r124_c117 bl[117] br[117] wl[124] vdd gnd cell_6t
Xbit_r125_c117 bl[117] br[117] wl[125] vdd gnd cell_6t
Xbit_r126_c117 bl[117] br[117] wl[126] vdd gnd cell_6t
Xbit_r127_c117 bl[117] br[117] wl[127] vdd gnd cell_6t
Xbit_r0_c118 bl[118] br[118] wl[0] vdd gnd cell_6t
Xbit_r1_c118 bl[118] br[118] wl[1] vdd gnd cell_6t
Xbit_r2_c118 bl[118] br[118] wl[2] vdd gnd cell_6t
Xbit_r3_c118 bl[118] br[118] wl[3] vdd gnd cell_6t
Xbit_r4_c118 bl[118] br[118] wl[4] vdd gnd cell_6t
Xbit_r5_c118 bl[118] br[118] wl[5] vdd gnd cell_6t
Xbit_r6_c118 bl[118] br[118] wl[6] vdd gnd cell_6t
Xbit_r7_c118 bl[118] br[118] wl[7] vdd gnd cell_6t
Xbit_r8_c118 bl[118] br[118] wl[8] vdd gnd cell_6t
Xbit_r9_c118 bl[118] br[118] wl[9] vdd gnd cell_6t
Xbit_r10_c118 bl[118] br[118] wl[10] vdd gnd cell_6t
Xbit_r11_c118 bl[118] br[118] wl[11] vdd gnd cell_6t
Xbit_r12_c118 bl[118] br[118] wl[12] vdd gnd cell_6t
Xbit_r13_c118 bl[118] br[118] wl[13] vdd gnd cell_6t
Xbit_r14_c118 bl[118] br[118] wl[14] vdd gnd cell_6t
Xbit_r15_c118 bl[118] br[118] wl[15] vdd gnd cell_6t
Xbit_r16_c118 bl[118] br[118] wl[16] vdd gnd cell_6t
Xbit_r17_c118 bl[118] br[118] wl[17] vdd gnd cell_6t
Xbit_r18_c118 bl[118] br[118] wl[18] vdd gnd cell_6t
Xbit_r19_c118 bl[118] br[118] wl[19] vdd gnd cell_6t
Xbit_r20_c118 bl[118] br[118] wl[20] vdd gnd cell_6t
Xbit_r21_c118 bl[118] br[118] wl[21] vdd gnd cell_6t
Xbit_r22_c118 bl[118] br[118] wl[22] vdd gnd cell_6t
Xbit_r23_c118 bl[118] br[118] wl[23] vdd gnd cell_6t
Xbit_r24_c118 bl[118] br[118] wl[24] vdd gnd cell_6t
Xbit_r25_c118 bl[118] br[118] wl[25] vdd gnd cell_6t
Xbit_r26_c118 bl[118] br[118] wl[26] vdd gnd cell_6t
Xbit_r27_c118 bl[118] br[118] wl[27] vdd gnd cell_6t
Xbit_r28_c118 bl[118] br[118] wl[28] vdd gnd cell_6t
Xbit_r29_c118 bl[118] br[118] wl[29] vdd gnd cell_6t
Xbit_r30_c118 bl[118] br[118] wl[30] vdd gnd cell_6t
Xbit_r31_c118 bl[118] br[118] wl[31] vdd gnd cell_6t
Xbit_r32_c118 bl[118] br[118] wl[32] vdd gnd cell_6t
Xbit_r33_c118 bl[118] br[118] wl[33] vdd gnd cell_6t
Xbit_r34_c118 bl[118] br[118] wl[34] vdd gnd cell_6t
Xbit_r35_c118 bl[118] br[118] wl[35] vdd gnd cell_6t
Xbit_r36_c118 bl[118] br[118] wl[36] vdd gnd cell_6t
Xbit_r37_c118 bl[118] br[118] wl[37] vdd gnd cell_6t
Xbit_r38_c118 bl[118] br[118] wl[38] vdd gnd cell_6t
Xbit_r39_c118 bl[118] br[118] wl[39] vdd gnd cell_6t
Xbit_r40_c118 bl[118] br[118] wl[40] vdd gnd cell_6t
Xbit_r41_c118 bl[118] br[118] wl[41] vdd gnd cell_6t
Xbit_r42_c118 bl[118] br[118] wl[42] vdd gnd cell_6t
Xbit_r43_c118 bl[118] br[118] wl[43] vdd gnd cell_6t
Xbit_r44_c118 bl[118] br[118] wl[44] vdd gnd cell_6t
Xbit_r45_c118 bl[118] br[118] wl[45] vdd gnd cell_6t
Xbit_r46_c118 bl[118] br[118] wl[46] vdd gnd cell_6t
Xbit_r47_c118 bl[118] br[118] wl[47] vdd gnd cell_6t
Xbit_r48_c118 bl[118] br[118] wl[48] vdd gnd cell_6t
Xbit_r49_c118 bl[118] br[118] wl[49] vdd gnd cell_6t
Xbit_r50_c118 bl[118] br[118] wl[50] vdd gnd cell_6t
Xbit_r51_c118 bl[118] br[118] wl[51] vdd gnd cell_6t
Xbit_r52_c118 bl[118] br[118] wl[52] vdd gnd cell_6t
Xbit_r53_c118 bl[118] br[118] wl[53] vdd gnd cell_6t
Xbit_r54_c118 bl[118] br[118] wl[54] vdd gnd cell_6t
Xbit_r55_c118 bl[118] br[118] wl[55] vdd gnd cell_6t
Xbit_r56_c118 bl[118] br[118] wl[56] vdd gnd cell_6t
Xbit_r57_c118 bl[118] br[118] wl[57] vdd gnd cell_6t
Xbit_r58_c118 bl[118] br[118] wl[58] vdd gnd cell_6t
Xbit_r59_c118 bl[118] br[118] wl[59] vdd gnd cell_6t
Xbit_r60_c118 bl[118] br[118] wl[60] vdd gnd cell_6t
Xbit_r61_c118 bl[118] br[118] wl[61] vdd gnd cell_6t
Xbit_r62_c118 bl[118] br[118] wl[62] vdd gnd cell_6t
Xbit_r63_c118 bl[118] br[118] wl[63] vdd gnd cell_6t
Xbit_r64_c118 bl[118] br[118] wl[64] vdd gnd cell_6t
Xbit_r65_c118 bl[118] br[118] wl[65] vdd gnd cell_6t
Xbit_r66_c118 bl[118] br[118] wl[66] vdd gnd cell_6t
Xbit_r67_c118 bl[118] br[118] wl[67] vdd gnd cell_6t
Xbit_r68_c118 bl[118] br[118] wl[68] vdd gnd cell_6t
Xbit_r69_c118 bl[118] br[118] wl[69] vdd gnd cell_6t
Xbit_r70_c118 bl[118] br[118] wl[70] vdd gnd cell_6t
Xbit_r71_c118 bl[118] br[118] wl[71] vdd gnd cell_6t
Xbit_r72_c118 bl[118] br[118] wl[72] vdd gnd cell_6t
Xbit_r73_c118 bl[118] br[118] wl[73] vdd gnd cell_6t
Xbit_r74_c118 bl[118] br[118] wl[74] vdd gnd cell_6t
Xbit_r75_c118 bl[118] br[118] wl[75] vdd gnd cell_6t
Xbit_r76_c118 bl[118] br[118] wl[76] vdd gnd cell_6t
Xbit_r77_c118 bl[118] br[118] wl[77] vdd gnd cell_6t
Xbit_r78_c118 bl[118] br[118] wl[78] vdd gnd cell_6t
Xbit_r79_c118 bl[118] br[118] wl[79] vdd gnd cell_6t
Xbit_r80_c118 bl[118] br[118] wl[80] vdd gnd cell_6t
Xbit_r81_c118 bl[118] br[118] wl[81] vdd gnd cell_6t
Xbit_r82_c118 bl[118] br[118] wl[82] vdd gnd cell_6t
Xbit_r83_c118 bl[118] br[118] wl[83] vdd gnd cell_6t
Xbit_r84_c118 bl[118] br[118] wl[84] vdd gnd cell_6t
Xbit_r85_c118 bl[118] br[118] wl[85] vdd gnd cell_6t
Xbit_r86_c118 bl[118] br[118] wl[86] vdd gnd cell_6t
Xbit_r87_c118 bl[118] br[118] wl[87] vdd gnd cell_6t
Xbit_r88_c118 bl[118] br[118] wl[88] vdd gnd cell_6t
Xbit_r89_c118 bl[118] br[118] wl[89] vdd gnd cell_6t
Xbit_r90_c118 bl[118] br[118] wl[90] vdd gnd cell_6t
Xbit_r91_c118 bl[118] br[118] wl[91] vdd gnd cell_6t
Xbit_r92_c118 bl[118] br[118] wl[92] vdd gnd cell_6t
Xbit_r93_c118 bl[118] br[118] wl[93] vdd gnd cell_6t
Xbit_r94_c118 bl[118] br[118] wl[94] vdd gnd cell_6t
Xbit_r95_c118 bl[118] br[118] wl[95] vdd gnd cell_6t
Xbit_r96_c118 bl[118] br[118] wl[96] vdd gnd cell_6t
Xbit_r97_c118 bl[118] br[118] wl[97] vdd gnd cell_6t
Xbit_r98_c118 bl[118] br[118] wl[98] vdd gnd cell_6t
Xbit_r99_c118 bl[118] br[118] wl[99] vdd gnd cell_6t
Xbit_r100_c118 bl[118] br[118] wl[100] vdd gnd cell_6t
Xbit_r101_c118 bl[118] br[118] wl[101] vdd gnd cell_6t
Xbit_r102_c118 bl[118] br[118] wl[102] vdd gnd cell_6t
Xbit_r103_c118 bl[118] br[118] wl[103] vdd gnd cell_6t
Xbit_r104_c118 bl[118] br[118] wl[104] vdd gnd cell_6t
Xbit_r105_c118 bl[118] br[118] wl[105] vdd gnd cell_6t
Xbit_r106_c118 bl[118] br[118] wl[106] vdd gnd cell_6t
Xbit_r107_c118 bl[118] br[118] wl[107] vdd gnd cell_6t
Xbit_r108_c118 bl[118] br[118] wl[108] vdd gnd cell_6t
Xbit_r109_c118 bl[118] br[118] wl[109] vdd gnd cell_6t
Xbit_r110_c118 bl[118] br[118] wl[110] vdd gnd cell_6t
Xbit_r111_c118 bl[118] br[118] wl[111] vdd gnd cell_6t
Xbit_r112_c118 bl[118] br[118] wl[112] vdd gnd cell_6t
Xbit_r113_c118 bl[118] br[118] wl[113] vdd gnd cell_6t
Xbit_r114_c118 bl[118] br[118] wl[114] vdd gnd cell_6t
Xbit_r115_c118 bl[118] br[118] wl[115] vdd gnd cell_6t
Xbit_r116_c118 bl[118] br[118] wl[116] vdd gnd cell_6t
Xbit_r117_c118 bl[118] br[118] wl[117] vdd gnd cell_6t
Xbit_r118_c118 bl[118] br[118] wl[118] vdd gnd cell_6t
Xbit_r119_c118 bl[118] br[118] wl[119] vdd gnd cell_6t
Xbit_r120_c118 bl[118] br[118] wl[120] vdd gnd cell_6t
Xbit_r121_c118 bl[118] br[118] wl[121] vdd gnd cell_6t
Xbit_r122_c118 bl[118] br[118] wl[122] vdd gnd cell_6t
Xbit_r123_c118 bl[118] br[118] wl[123] vdd gnd cell_6t
Xbit_r124_c118 bl[118] br[118] wl[124] vdd gnd cell_6t
Xbit_r125_c118 bl[118] br[118] wl[125] vdd gnd cell_6t
Xbit_r126_c118 bl[118] br[118] wl[126] vdd gnd cell_6t
Xbit_r127_c118 bl[118] br[118] wl[127] vdd gnd cell_6t
Xbit_r0_c119 bl[119] br[119] wl[0] vdd gnd cell_6t
Xbit_r1_c119 bl[119] br[119] wl[1] vdd gnd cell_6t
Xbit_r2_c119 bl[119] br[119] wl[2] vdd gnd cell_6t
Xbit_r3_c119 bl[119] br[119] wl[3] vdd gnd cell_6t
Xbit_r4_c119 bl[119] br[119] wl[4] vdd gnd cell_6t
Xbit_r5_c119 bl[119] br[119] wl[5] vdd gnd cell_6t
Xbit_r6_c119 bl[119] br[119] wl[6] vdd gnd cell_6t
Xbit_r7_c119 bl[119] br[119] wl[7] vdd gnd cell_6t
Xbit_r8_c119 bl[119] br[119] wl[8] vdd gnd cell_6t
Xbit_r9_c119 bl[119] br[119] wl[9] vdd gnd cell_6t
Xbit_r10_c119 bl[119] br[119] wl[10] vdd gnd cell_6t
Xbit_r11_c119 bl[119] br[119] wl[11] vdd gnd cell_6t
Xbit_r12_c119 bl[119] br[119] wl[12] vdd gnd cell_6t
Xbit_r13_c119 bl[119] br[119] wl[13] vdd gnd cell_6t
Xbit_r14_c119 bl[119] br[119] wl[14] vdd gnd cell_6t
Xbit_r15_c119 bl[119] br[119] wl[15] vdd gnd cell_6t
Xbit_r16_c119 bl[119] br[119] wl[16] vdd gnd cell_6t
Xbit_r17_c119 bl[119] br[119] wl[17] vdd gnd cell_6t
Xbit_r18_c119 bl[119] br[119] wl[18] vdd gnd cell_6t
Xbit_r19_c119 bl[119] br[119] wl[19] vdd gnd cell_6t
Xbit_r20_c119 bl[119] br[119] wl[20] vdd gnd cell_6t
Xbit_r21_c119 bl[119] br[119] wl[21] vdd gnd cell_6t
Xbit_r22_c119 bl[119] br[119] wl[22] vdd gnd cell_6t
Xbit_r23_c119 bl[119] br[119] wl[23] vdd gnd cell_6t
Xbit_r24_c119 bl[119] br[119] wl[24] vdd gnd cell_6t
Xbit_r25_c119 bl[119] br[119] wl[25] vdd gnd cell_6t
Xbit_r26_c119 bl[119] br[119] wl[26] vdd gnd cell_6t
Xbit_r27_c119 bl[119] br[119] wl[27] vdd gnd cell_6t
Xbit_r28_c119 bl[119] br[119] wl[28] vdd gnd cell_6t
Xbit_r29_c119 bl[119] br[119] wl[29] vdd gnd cell_6t
Xbit_r30_c119 bl[119] br[119] wl[30] vdd gnd cell_6t
Xbit_r31_c119 bl[119] br[119] wl[31] vdd gnd cell_6t
Xbit_r32_c119 bl[119] br[119] wl[32] vdd gnd cell_6t
Xbit_r33_c119 bl[119] br[119] wl[33] vdd gnd cell_6t
Xbit_r34_c119 bl[119] br[119] wl[34] vdd gnd cell_6t
Xbit_r35_c119 bl[119] br[119] wl[35] vdd gnd cell_6t
Xbit_r36_c119 bl[119] br[119] wl[36] vdd gnd cell_6t
Xbit_r37_c119 bl[119] br[119] wl[37] vdd gnd cell_6t
Xbit_r38_c119 bl[119] br[119] wl[38] vdd gnd cell_6t
Xbit_r39_c119 bl[119] br[119] wl[39] vdd gnd cell_6t
Xbit_r40_c119 bl[119] br[119] wl[40] vdd gnd cell_6t
Xbit_r41_c119 bl[119] br[119] wl[41] vdd gnd cell_6t
Xbit_r42_c119 bl[119] br[119] wl[42] vdd gnd cell_6t
Xbit_r43_c119 bl[119] br[119] wl[43] vdd gnd cell_6t
Xbit_r44_c119 bl[119] br[119] wl[44] vdd gnd cell_6t
Xbit_r45_c119 bl[119] br[119] wl[45] vdd gnd cell_6t
Xbit_r46_c119 bl[119] br[119] wl[46] vdd gnd cell_6t
Xbit_r47_c119 bl[119] br[119] wl[47] vdd gnd cell_6t
Xbit_r48_c119 bl[119] br[119] wl[48] vdd gnd cell_6t
Xbit_r49_c119 bl[119] br[119] wl[49] vdd gnd cell_6t
Xbit_r50_c119 bl[119] br[119] wl[50] vdd gnd cell_6t
Xbit_r51_c119 bl[119] br[119] wl[51] vdd gnd cell_6t
Xbit_r52_c119 bl[119] br[119] wl[52] vdd gnd cell_6t
Xbit_r53_c119 bl[119] br[119] wl[53] vdd gnd cell_6t
Xbit_r54_c119 bl[119] br[119] wl[54] vdd gnd cell_6t
Xbit_r55_c119 bl[119] br[119] wl[55] vdd gnd cell_6t
Xbit_r56_c119 bl[119] br[119] wl[56] vdd gnd cell_6t
Xbit_r57_c119 bl[119] br[119] wl[57] vdd gnd cell_6t
Xbit_r58_c119 bl[119] br[119] wl[58] vdd gnd cell_6t
Xbit_r59_c119 bl[119] br[119] wl[59] vdd gnd cell_6t
Xbit_r60_c119 bl[119] br[119] wl[60] vdd gnd cell_6t
Xbit_r61_c119 bl[119] br[119] wl[61] vdd gnd cell_6t
Xbit_r62_c119 bl[119] br[119] wl[62] vdd gnd cell_6t
Xbit_r63_c119 bl[119] br[119] wl[63] vdd gnd cell_6t
Xbit_r64_c119 bl[119] br[119] wl[64] vdd gnd cell_6t
Xbit_r65_c119 bl[119] br[119] wl[65] vdd gnd cell_6t
Xbit_r66_c119 bl[119] br[119] wl[66] vdd gnd cell_6t
Xbit_r67_c119 bl[119] br[119] wl[67] vdd gnd cell_6t
Xbit_r68_c119 bl[119] br[119] wl[68] vdd gnd cell_6t
Xbit_r69_c119 bl[119] br[119] wl[69] vdd gnd cell_6t
Xbit_r70_c119 bl[119] br[119] wl[70] vdd gnd cell_6t
Xbit_r71_c119 bl[119] br[119] wl[71] vdd gnd cell_6t
Xbit_r72_c119 bl[119] br[119] wl[72] vdd gnd cell_6t
Xbit_r73_c119 bl[119] br[119] wl[73] vdd gnd cell_6t
Xbit_r74_c119 bl[119] br[119] wl[74] vdd gnd cell_6t
Xbit_r75_c119 bl[119] br[119] wl[75] vdd gnd cell_6t
Xbit_r76_c119 bl[119] br[119] wl[76] vdd gnd cell_6t
Xbit_r77_c119 bl[119] br[119] wl[77] vdd gnd cell_6t
Xbit_r78_c119 bl[119] br[119] wl[78] vdd gnd cell_6t
Xbit_r79_c119 bl[119] br[119] wl[79] vdd gnd cell_6t
Xbit_r80_c119 bl[119] br[119] wl[80] vdd gnd cell_6t
Xbit_r81_c119 bl[119] br[119] wl[81] vdd gnd cell_6t
Xbit_r82_c119 bl[119] br[119] wl[82] vdd gnd cell_6t
Xbit_r83_c119 bl[119] br[119] wl[83] vdd gnd cell_6t
Xbit_r84_c119 bl[119] br[119] wl[84] vdd gnd cell_6t
Xbit_r85_c119 bl[119] br[119] wl[85] vdd gnd cell_6t
Xbit_r86_c119 bl[119] br[119] wl[86] vdd gnd cell_6t
Xbit_r87_c119 bl[119] br[119] wl[87] vdd gnd cell_6t
Xbit_r88_c119 bl[119] br[119] wl[88] vdd gnd cell_6t
Xbit_r89_c119 bl[119] br[119] wl[89] vdd gnd cell_6t
Xbit_r90_c119 bl[119] br[119] wl[90] vdd gnd cell_6t
Xbit_r91_c119 bl[119] br[119] wl[91] vdd gnd cell_6t
Xbit_r92_c119 bl[119] br[119] wl[92] vdd gnd cell_6t
Xbit_r93_c119 bl[119] br[119] wl[93] vdd gnd cell_6t
Xbit_r94_c119 bl[119] br[119] wl[94] vdd gnd cell_6t
Xbit_r95_c119 bl[119] br[119] wl[95] vdd gnd cell_6t
Xbit_r96_c119 bl[119] br[119] wl[96] vdd gnd cell_6t
Xbit_r97_c119 bl[119] br[119] wl[97] vdd gnd cell_6t
Xbit_r98_c119 bl[119] br[119] wl[98] vdd gnd cell_6t
Xbit_r99_c119 bl[119] br[119] wl[99] vdd gnd cell_6t
Xbit_r100_c119 bl[119] br[119] wl[100] vdd gnd cell_6t
Xbit_r101_c119 bl[119] br[119] wl[101] vdd gnd cell_6t
Xbit_r102_c119 bl[119] br[119] wl[102] vdd gnd cell_6t
Xbit_r103_c119 bl[119] br[119] wl[103] vdd gnd cell_6t
Xbit_r104_c119 bl[119] br[119] wl[104] vdd gnd cell_6t
Xbit_r105_c119 bl[119] br[119] wl[105] vdd gnd cell_6t
Xbit_r106_c119 bl[119] br[119] wl[106] vdd gnd cell_6t
Xbit_r107_c119 bl[119] br[119] wl[107] vdd gnd cell_6t
Xbit_r108_c119 bl[119] br[119] wl[108] vdd gnd cell_6t
Xbit_r109_c119 bl[119] br[119] wl[109] vdd gnd cell_6t
Xbit_r110_c119 bl[119] br[119] wl[110] vdd gnd cell_6t
Xbit_r111_c119 bl[119] br[119] wl[111] vdd gnd cell_6t
Xbit_r112_c119 bl[119] br[119] wl[112] vdd gnd cell_6t
Xbit_r113_c119 bl[119] br[119] wl[113] vdd gnd cell_6t
Xbit_r114_c119 bl[119] br[119] wl[114] vdd gnd cell_6t
Xbit_r115_c119 bl[119] br[119] wl[115] vdd gnd cell_6t
Xbit_r116_c119 bl[119] br[119] wl[116] vdd gnd cell_6t
Xbit_r117_c119 bl[119] br[119] wl[117] vdd gnd cell_6t
Xbit_r118_c119 bl[119] br[119] wl[118] vdd gnd cell_6t
Xbit_r119_c119 bl[119] br[119] wl[119] vdd gnd cell_6t
Xbit_r120_c119 bl[119] br[119] wl[120] vdd gnd cell_6t
Xbit_r121_c119 bl[119] br[119] wl[121] vdd gnd cell_6t
Xbit_r122_c119 bl[119] br[119] wl[122] vdd gnd cell_6t
Xbit_r123_c119 bl[119] br[119] wl[123] vdd gnd cell_6t
Xbit_r124_c119 bl[119] br[119] wl[124] vdd gnd cell_6t
Xbit_r125_c119 bl[119] br[119] wl[125] vdd gnd cell_6t
Xbit_r126_c119 bl[119] br[119] wl[126] vdd gnd cell_6t
Xbit_r127_c119 bl[119] br[119] wl[127] vdd gnd cell_6t
Xbit_r0_c120 bl[120] br[120] wl[0] vdd gnd cell_6t
Xbit_r1_c120 bl[120] br[120] wl[1] vdd gnd cell_6t
Xbit_r2_c120 bl[120] br[120] wl[2] vdd gnd cell_6t
Xbit_r3_c120 bl[120] br[120] wl[3] vdd gnd cell_6t
Xbit_r4_c120 bl[120] br[120] wl[4] vdd gnd cell_6t
Xbit_r5_c120 bl[120] br[120] wl[5] vdd gnd cell_6t
Xbit_r6_c120 bl[120] br[120] wl[6] vdd gnd cell_6t
Xbit_r7_c120 bl[120] br[120] wl[7] vdd gnd cell_6t
Xbit_r8_c120 bl[120] br[120] wl[8] vdd gnd cell_6t
Xbit_r9_c120 bl[120] br[120] wl[9] vdd gnd cell_6t
Xbit_r10_c120 bl[120] br[120] wl[10] vdd gnd cell_6t
Xbit_r11_c120 bl[120] br[120] wl[11] vdd gnd cell_6t
Xbit_r12_c120 bl[120] br[120] wl[12] vdd gnd cell_6t
Xbit_r13_c120 bl[120] br[120] wl[13] vdd gnd cell_6t
Xbit_r14_c120 bl[120] br[120] wl[14] vdd gnd cell_6t
Xbit_r15_c120 bl[120] br[120] wl[15] vdd gnd cell_6t
Xbit_r16_c120 bl[120] br[120] wl[16] vdd gnd cell_6t
Xbit_r17_c120 bl[120] br[120] wl[17] vdd gnd cell_6t
Xbit_r18_c120 bl[120] br[120] wl[18] vdd gnd cell_6t
Xbit_r19_c120 bl[120] br[120] wl[19] vdd gnd cell_6t
Xbit_r20_c120 bl[120] br[120] wl[20] vdd gnd cell_6t
Xbit_r21_c120 bl[120] br[120] wl[21] vdd gnd cell_6t
Xbit_r22_c120 bl[120] br[120] wl[22] vdd gnd cell_6t
Xbit_r23_c120 bl[120] br[120] wl[23] vdd gnd cell_6t
Xbit_r24_c120 bl[120] br[120] wl[24] vdd gnd cell_6t
Xbit_r25_c120 bl[120] br[120] wl[25] vdd gnd cell_6t
Xbit_r26_c120 bl[120] br[120] wl[26] vdd gnd cell_6t
Xbit_r27_c120 bl[120] br[120] wl[27] vdd gnd cell_6t
Xbit_r28_c120 bl[120] br[120] wl[28] vdd gnd cell_6t
Xbit_r29_c120 bl[120] br[120] wl[29] vdd gnd cell_6t
Xbit_r30_c120 bl[120] br[120] wl[30] vdd gnd cell_6t
Xbit_r31_c120 bl[120] br[120] wl[31] vdd gnd cell_6t
Xbit_r32_c120 bl[120] br[120] wl[32] vdd gnd cell_6t
Xbit_r33_c120 bl[120] br[120] wl[33] vdd gnd cell_6t
Xbit_r34_c120 bl[120] br[120] wl[34] vdd gnd cell_6t
Xbit_r35_c120 bl[120] br[120] wl[35] vdd gnd cell_6t
Xbit_r36_c120 bl[120] br[120] wl[36] vdd gnd cell_6t
Xbit_r37_c120 bl[120] br[120] wl[37] vdd gnd cell_6t
Xbit_r38_c120 bl[120] br[120] wl[38] vdd gnd cell_6t
Xbit_r39_c120 bl[120] br[120] wl[39] vdd gnd cell_6t
Xbit_r40_c120 bl[120] br[120] wl[40] vdd gnd cell_6t
Xbit_r41_c120 bl[120] br[120] wl[41] vdd gnd cell_6t
Xbit_r42_c120 bl[120] br[120] wl[42] vdd gnd cell_6t
Xbit_r43_c120 bl[120] br[120] wl[43] vdd gnd cell_6t
Xbit_r44_c120 bl[120] br[120] wl[44] vdd gnd cell_6t
Xbit_r45_c120 bl[120] br[120] wl[45] vdd gnd cell_6t
Xbit_r46_c120 bl[120] br[120] wl[46] vdd gnd cell_6t
Xbit_r47_c120 bl[120] br[120] wl[47] vdd gnd cell_6t
Xbit_r48_c120 bl[120] br[120] wl[48] vdd gnd cell_6t
Xbit_r49_c120 bl[120] br[120] wl[49] vdd gnd cell_6t
Xbit_r50_c120 bl[120] br[120] wl[50] vdd gnd cell_6t
Xbit_r51_c120 bl[120] br[120] wl[51] vdd gnd cell_6t
Xbit_r52_c120 bl[120] br[120] wl[52] vdd gnd cell_6t
Xbit_r53_c120 bl[120] br[120] wl[53] vdd gnd cell_6t
Xbit_r54_c120 bl[120] br[120] wl[54] vdd gnd cell_6t
Xbit_r55_c120 bl[120] br[120] wl[55] vdd gnd cell_6t
Xbit_r56_c120 bl[120] br[120] wl[56] vdd gnd cell_6t
Xbit_r57_c120 bl[120] br[120] wl[57] vdd gnd cell_6t
Xbit_r58_c120 bl[120] br[120] wl[58] vdd gnd cell_6t
Xbit_r59_c120 bl[120] br[120] wl[59] vdd gnd cell_6t
Xbit_r60_c120 bl[120] br[120] wl[60] vdd gnd cell_6t
Xbit_r61_c120 bl[120] br[120] wl[61] vdd gnd cell_6t
Xbit_r62_c120 bl[120] br[120] wl[62] vdd gnd cell_6t
Xbit_r63_c120 bl[120] br[120] wl[63] vdd gnd cell_6t
Xbit_r64_c120 bl[120] br[120] wl[64] vdd gnd cell_6t
Xbit_r65_c120 bl[120] br[120] wl[65] vdd gnd cell_6t
Xbit_r66_c120 bl[120] br[120] wl[66] vdd gnd cell_6t
Xbit_r67_c120 bl[120] br[120] wl[67] vdd gnd cell_6t
Xbit_r68_c120 bl[120] br[120] wl[68] vdd gnd cell_6t
Xbit_r69_c120 bl[120] br[120] wl[69] vdd gnd cell_6t
Xbit_r70_c120 bl[120] br[120] wl[70] vdd gnd cell_6t
Xbit_r71_c120 bl[120] br[120] wl[71] vdd gnd cell_6t
Xbit_r72_c120 bl[120] br[120] wl[72] vdd gnd cell_6t
Xbit_r73_c120 bl[120] br[120] wl[73] vdd gnd cell_6t
Xbit_r74_c120 bl[120] br[120] wl[74] vdd gnd cell_6t
Xbit_r75_c120 bl[120] br[120] wl[75] vdd gnd cell_6t
Xbit_r76_c120 bl[120] br[120] wl[76] vdd gnd cell_6t
Xbit_r77_c120 bl[120] br[120] wl[77] vdd gnd cell_6t
Xbit_r78_c120 bl[120] br[120] wl[78] vdd gnd cell_6t
Xbit_r79_c120 bl[120] br[120] wl[79] vdd gnd cell_6t
Xbit_r80_c120 bl[120] br[120] wl[80] vdd gnd cell_6t
Xbit_r81_c120 bl[120] br[120] wl[81] vdd gnd cell_6t
Xbit_r82_c120 bl[120] br[120] wl[82] vdd gnd cell_6t
Xbit_r83_c120 bl[120] br[120] wl[83] vdd gnd cell_6t
Xbit_r84_c120 bl[120] br[120] wl[84] vdd gnd cell_6t
Xbit_r85_c120 bl[120] br[120] wl[85] vdd gnd cell_6t
Xbit_r86_c120 bl[120] br[120] wl[86] vdd gnd cell_6t
Xbit_r87_c120 bl[120] br[120] wl[87] vdd gnd cell_6t
Xbit_r88_c120 bl[120] br[120] wl[88] vdd gnd cell_6t
Xbit_r89_c120 bl[120] br[120] wl[89] vdd gnd cell_6t
Xbit_r90_c120 bl[120] br[120] wl[90] vdd gnd cell_6t
Xbit_r91_c120 bl[120] br[120] wl[91] vdd gnd cell_6t
Xbit_r92_c120 bl[120] br[120] wl[92] vdd gnd cell_6t
Xbit_r93_c120 bl[120] br[120] wl[93] vdd gnd cell_6t
Xbit_r94_c120 bl[120] br[120] wl[94] vdd gnd cell_6t
Xbit_r95_c120 bl[120] br[120] wl[95] vdd gnd cell_6t
Xbit_r96_c120 bl[120] br[120] wl[96] vdd gnd cell_6t
Xbit_r97_c120 bl[120] br[120] wl[97] vdd gnd cell_6t
Xbit_r98_c120 bl[120] br[120] wl[98] vdd gnd cell_6t
Xbit_r99_c120 bl[120] br[120] wl[99] vdd gnd cell_6t
Xbit_r100_c120 bl[120] br[120] wl[100] vdd gnd cell_6t
Xbit_r101_c120 bl[120] br[120] wl[101] vdd gnd cell_6t
Xbit_r102_c120 bl[120] br[120] wl[102] vdd gnd cell_6t
Xbit_r103_c120 bl[120] br[120] wl[103] vdd gnd cell_6t
Xbit_r104_c120 bl[120] br[120] wl[104] vdd gnd cell_6t
Xbit_r105_c120 bl[120] br[120] wl[105] vdd gnd cell_6t
Xbit_r106_c120 bl[120] br[120] wl[106] vdd gnd cell_6t
Xbit_r107_c120 bl[120] br[120] wl[107] vdd gnd cell_6t
Xbit_r108_c120 bl[120] br[120] wl[108] vdd gnd cell_6t
Xbit_r109_c120 bl[120] br[120] wl[109] vdd gnd cell_6t
Xbit_r110_c120 bl[120] br[120] wl[110] vdd gnd cell_6t
Xbit_r111_c120 bl[120] br[120] wl[111] vdd gnd cell_6t
Xbit_r112_c120 bl[120] br[120] wl[112] vdd gnd cell_6t
Xbit_r113_c120 bl[120] br[120] wl[113] vdd gnd cell_6t
Xbit_r114_c120 bl[120] br[120] wl[114] vdd gnd cell_6t
Xbit_r115_c120 bl[120] br[120] wl[115] vdd gnd cell_6t
Xbit_r116_c120 bl[120] br[120] wl[116] vdd gnd cell_6t
Xbit_r117_c120 bl[120] br[120] wl[117] vdd gnd cell_6t
Xbit_r118_c120 bl[120] br[120] wl[118] vdd gnd cell_6t
Xbit_r119_c120 bl[120] br[120] wl[119] vdd gnd cell_6t
Xbit_r120_c120 bl[120] br[120] wl[120] vdd gnd cell_6t
Xbit_r121_c120 bl[120] br[120] wl[121] vdd gnd cell_6t
Xbit_r122_c120 bl[120] br[120] wl[122] vdd gnd cell_6t
Xbit_r123_c120 bl[120] br[120] wl[123] vdd gnd cell_6t
Xbit_r124_c120 bl[120] br[120] wl[124] vdd gnd cell_6t
Xbit_r125_c120 bl[120] br[120] wl[125] vdd gnd cell_6t
Xbit_r126_c120 bl[120] br[120] wl[126] vdd gnd cell_6t
Xbit_r127_c120 bl[120] br[120] wl[127] vdd gnd cell_6t
Xbit_r0_c121 bl[121] br[121] wl[0] vdd gnd cell_6t
Xbit_r1_c121 bl[121] br[121] wl[1] vdd gnd cell_6t
Xbit_r2_c121 bl[121] br[121] wl[2] vdd gnd cell_6t
Xbit_r3_c121 bl[121] br[121] wl[3] vdd gnd cell_6t
Xbit_r4_c121 bl[121] br[121] wl[4] vdd gnd cell_6t
Xbit_r5_c121 bl[121] br[121] wl[5] vdd gnd cell_6t
Xbit_r6_c121 bl[121] br[121] wl[6] vdd gnd cell_6t
Xbit_r7_c121 bl[121] br[121] wl[7] vdd gnd cell_6t
Xbit_r8_c121 bl[121] br[121] wl[8] vdd gnd cell_6t
Xbit_r9_c121 bl[121] br[121] wl[9] vdd gnd cell_6t
Xbit_r10_c121 bl[121] br[121] wl[10] vdd gnd cell_6t
Xbit_r11_c121 bl[121] br[121] wl[11] vdd gnd cell_6t
Xbit_r12_c121 bl[121] br[121] wl[12] vdd gnd cell_6t
Xbit_r13_c121 bl[121] br[121] wl[13] vdd gnd cell_6t
Xbit_r14_c121 bl[121] br[121] wl[14] vdd gnd cell_6t
Xbit_r15_c121 bl[121] br[121] wl[15] vdd gnd cell_6t
Xbit_r16_c121 bl[121] br[121] wl[16] vdd gnd cell_6t
Xbit_r17_c121 bl[121] br[121] wl[17] vdd gnd cell_6t
Xbit_r18_c121 bl[121] br[121] wl[18] vdd gnd cell_6t
Xbit_r19_c121 bl[121] br[121] wl[19] vdd gnd cell_6t
Xbit_r20_c121 bl[121] br[121] wl[20] vdd gnd cell_6t
Xbit_r21_c121 bl[121] br[121] wl[21] vdd gnd cell_6t
Xbit_r22_c121 bl[121] br[121] wl[22] vdd gnd cell_6t
Xbit_r23_c121 bl[121] br[121] wl[23] vdd gnd cell_6t
Xbit_r24_c121 bl[121] br[121] wl[24] vdd gnd cell_6t
Xbit_r25_c121 bl[121] br[121] wl[25] vdd gnd cell_6t
Xbit_r26_c121 bl[121] br[121] wl[26] vdd gnd cell_6t
Xbit_r27_c121 bl[121] br[121] wl[27] vdd gnd cell_6t
Xbit_r28_c121 bl[121] br[121] wl[28] vdd gnd cell_6t
Xbit_r29_c121 bl[121] br[121] wl[29] vdd gnd cell_6t
Xbit_r30_c121 bl[121] br[121] wl[30] vdd gnd cell_6t
Xbit_r31_c121 bl[121] br[121] wl[31] vdd gnd cell_6t
Xbit_r32_c121 bl[121] br[121] wl[32] vdd gnd cell_6t
Xbit_r33_c121 bl[121] br[121] wl[33] vdd gnd cell_6t
Xbit_r34_c121 bl[121] br[121] wl[34] vdd gnd cell_6t
Xbit_r35_c121 bl[121] br[121] wl[35] vdd gnd cell_6t
Xbit_r36_c121 bl[121] br[121] wl[36] vdd gnd cell_6t
Xbit_r37_c121 bl[121] br[121] wl[37] vdd gnd cell_6t
Xbit_r38_c121 bl[121] br[121] wl[38] vdd gnd cell_6t
Xbit_r39_c121 bl[121] br[121] wl[39] vdd gnd cell_6t
Xbit_r40_c121 bl[121] br[121] wl[40] vdd gnd cell_6t
Xbit_r41_c121 bl[121] br[121] wl[41] vdd gnd cell_6t
Xbit_r42_c121 bl[121] br[121] wl[42] vdd gnd cell_6t
Xbit_r43_c121 bl[121] br[121] wl[43] vdd gnd cell_6t
Xbit_r44_c121 bl[121] br[121] wl[44] vdd gnd cell_6t
Xbit_r45_c121 bl[121] br[121] wl[45] vdd gnd cell_6t
Xbit_r46_c121 bl[121] br[121] wl[46] vdd gnd cell_6t
Xbit_r47_c121 bl[121] br[121] wl[47] vdd gnd cell_6t
Xbit_r48_c121 bl[121] br[121] wl[48] vdd gnd cell_6t
Xbit_r49_c121 bl[121] br[121] wl[49] vdd gnd cell_6t
Xbit_r50_c121 bl[121] br[121] wl[50] vdd gnd cell_6t
Xbit_r51_c121 bl[121] br[121] wl[51] vdd gnd cell_6t
Xbit_r52_c121 bl[121] br[121] wl[52] vdd gnd cell_6t
Xbit_r53_c121 bl[121] br[121] wl[53] vdd gnd cell_6t
Xbit_r54_c121 bl[121] br[121] wl[54] vdd gnd cell_6t
Xbit_r55_c121 bl[121] br[121] wl[55] vdd gnd cell_6t
Xbit_r56_c121 bl[121] br[121] wl[56] vdd gnd cell_6t
Xbit_r57_c121 bl[121] br[121] wl[57] vdd gnd cell_6t
Xbit_r58_c121 bl[121] br[121] wl[58] vdd gnd cell_6t
Xbit_r59_c121 bl[121] br[121] wl[59] vdd gnd cell_6t
Xbit_r60_c121 bl[121] br[121] wl[60] vdd gnd cell_6t
Xbit_r61_c121 bl[121] br[121] wl[61] vdd gnd cell_6t
Xbit_r62_c121 bl[121] br[121] wl[62] vdd gnd cell_6t
Xbit_r63_c121 bl[121] br[121] wl[63] vdd gnd cell_6t
Xbit_r64_c121 bl[121] br[121] wl[64] vdd gnd cell_6t
Xbit_r65_c121 bl[121] br[121] wl[65] vdd gnd cell_6t
Xbit_r66_c121 bl[121] br[121] wl[66] vdd gnd cell_6t
Xbit_r67_c121 bl[121] br[121] wl[67] vdd gnd cell_6t
Xbit_r68_c121 bl[121] br[121] wl[68] vdd gnd cell_6t
Xbit_r69_c121 bl[121] br[121] wl[69] vdd gnd cell_6t
Xbit_r70_c121 bl[121] br[121] wl[70] vdd gnd cell_6t
Xbit_r71_c121 bl[121] br[121] wl[71] vdd gnd cell_6t
Xbit_r72_c121 bl[121] br[121] wl[72] vdd gnd cell_6t
Xbit_r73_c121 bl[121] br[121] wl[73] vdd gnd cell_6t
Xbit_r74_c121 bl[121] br[121] wl[74] vdd gnd cell_6t
Xbit_r75_c121 bl[121] br[121] wl[75] vdd gnd cell_6t
Xbit_r76_c121 bl[121] br[121] wl[76] vdd gnd cell_6t
Xbit_r77_c121 bl[121] br[121] wl[77] vdd gnd cell_6t
Xbit_r78_c121 bl[121] br[121] wl[78] vdd gnd cell_6t
Xbit_r79_c121 bl[121] br[121] wl[79] vdd gnd cell_6t
Xbit_r80_c121 bl[121] br[121] wl[80] vdd gnd cell_6t
Xbit_r81_c121 bl[121] br[121] wl[81] vdd gnd cell_6t
Xbit_r82_c121 bl[121] br[121] wl[82] vdd gnd cell_6t
Xbit_r83_c121 bl[121] br[121] wl[83] vdd gnd cell_6t
Xbit_r84_c121 bl[121] br[121] wl[84] vdd gnd cell_6t
Xbit_r85_c121 bl[121] br[121] wl[85] vdd gnd cell_6t
Xbit_r86_c121 bl[121] br[121] wl[86] vdd gnd cell_6t
Xbit_r87_c121 bl[121] br[121] wl[87] vdd gnd cell_6t
Xbit_r88_c121 bl[121] br[121] wl[88] vdd gnd cell_6t
Xbit_r89_c121 bl[121] br[121] wl[89] vdd gnd cell_6t
Xbit_r90_c121 bl[121] br[121] wl[90] vdd gnd cell_6t
Xbit_r91_c121 bl[121] br[121] wl[91] vdd gnd cell_6t
Xbit_r92_c121 bl[121] br[121] wl[92] vdd gnd cell_6t
Xbit_r93_c121 bl[121] br[121] wl[93] vdd gnd cell_6t
Xbit_r94_c121 bl[121] br[121] wl[94] vdd gnd cell_6t
Xbit_r95_c121 bl[121] br[121] wl[95] vdd gnd cell_6t
Xbit_r96_c121 bl[121] br[121] wl[96] vdd gnd cell_6t
Xbit_r97_c121 bl[121] br[121] wl[97] vdd gnd cell_6t
Xbit_r98_c121 bl[121] br[121] wl[98] vdd gnd cell_6t
Xbit_r99_c121 bl[121] br[121] wl[99] vdd gnd cell_6t
Xbit_r100_c121 bl[121] br[121] wl[100] vdd gnd cell_6t
Xbit_r101_c121 bl[121] br[121] wl[101] vdd gnd cell_6t
Xbit_r102_c121 bl[121] br[121] wl[102] vdd gnd cell_6t
Xbit_r103_c121 bl[121] br[121] wl[103] vdd gnd cell_6t
Xbit_r104_c121 bl[121] br[121] wl[104] vdd gnd cell_6t
Xbit_r105_c121 bl[121] br[121] wl[105] vdd gnd cell_6t
Xbit_r106_c121 bl[121] br[121] wl[106] vdd gnd cell_6t
Xbit_r107_c121 bl[121] br[121] wl[107] vdd gnd cell_6t
Xbit_r108_c121 bl[121] br[121] wl[108] vdd gnd cell_6t
Xbit_r109_c121 bl[121] br[121] wl[109] vdd gnd cell_6t
Xbit_r110_c121 bl[121] br[121] wl[110] vdd gnd cell_6t
Xbit_r111_c121 bl[121] br[121] wl[111] vdd gnd cell_6t
Xbit_r112_c121 bl[121] br[121] wl[112] vdd gnd cell_6t
Xbit_r113_c121 bl[121] br[121] wl[113] vdd gnd cell_6t
Xbit_r114_c121 bl[121] br[121] wl[114] vdd gnd cell_6t
Xbit_r115_c121 bl[121] br[121] wl[115] vdd gnd cell_6t
Xbit_r116_c121 bl[121] br[121] wl[116] vdd gnd cell_6t
Xbit_r117_c121 bl[121] br[121] wl[117] vdd gnd cell_6t
Xbit_r118_c121 bl[121] br[121] wl[118] vdd gnd cell_6t
Xbit_r119_c121 bl[121] br[121] wl[119] vdd gnd cell_6t
Xbit_r120_c121 bl[121] br[121] wl[120] vdd gnd cell_6t
Xbit_r121_c121 bl[121] br[121] wl[121] vdd gnd cell_6t
Xbit_r122_c121 bl[121] br[121] wl[122] vdd gnd cell_6t
Xbit_r123_c121 bl[121] br[121] wl[123] vdd gnd cell_6t
Xbit_r124_c121 bl[121] br[121] wl[124] vdd gnd cell_6t
Xbit_r125_c121 bl[121] br[121] wl[125] vdd gnd cell_6t
Xbit_r126_c121 bl[121] br[121] wl[126] vdd gnd cell_6t
Xbit_r127_c121 bl[121] br[121] wl[127] vdd gnd cell_6t
Xbit_r0_c122 bl[122] br[122] wl[0] vdd gnd cell_6t
Xbit_r1_c122 bl[122] br[122] wl[1] vdd gnd cell_6t
Xbit_r2_c122 bl[122] br[122] wl[2] vdd gnd cell_6t
Xbit_r3_c122 bl[122] br[122] wl[3] vdd gnd cell_6t
Xbit_r4_c122 bl[122] br[122] wl[4] vdd gnd cell_6t
Xbit_r5_c122 bl[122] br[122] wl[5] vdd gnd cell_6t
Xbit_r6_c122 bl[122] br[122] wl[6] vdd gnd cell_6t
Xbit_r7_c122 bl[122] br[122] wl[7] vdd gnd cell_6t
Xbit_r8_c122 bl[122] br[122] wl[8] vdd gnd cell_6t
Xbit_r9_c122 bl[122] br[122] wl[9] vdd gnd cell_6t
Xbit_r10_c122 bl[122] br[122] wl[10] vdd gnd cell_6t
Xbit_r11_c122 bl[122] br[122] wl[11] vdd gnd cell_6t
Xbit_r12_c122 bl[122] br[122] wl[12] vdd gnd cell_6t
Xbit_r13_c122 bl[122] br[122] wl[13] vdd gnd cell_6t
Xbit_r14_c122 bl[122] br[122] wl[14] vdd gnd cell_6t
Xbit_r15_c122 bl[122] br[122] wl[15] vdd gnd cell_6t
Xbit_r16_c122 bl[122] br[122] wl[16] vdd gnd cell_6t
Xbit_r17_c122 bl[122] br[122] wl[17] vdd gnd cell_6t
Xbit_r18_c122 bl[122] br[122] wl[18] vdd gnd cell_6t
Xbit_r19_c122 bl[122] br[122] wl[19] vdd gnd cell_6t
Xbit_r20_c122 bl[122] br[122] wl[20] vdd gnd cell_6t
Xbit_r21_c122 bl[122] br[122] wl[21] vdd gnd cell_6t
Xbit_r22_c122 bl[122] br[122] wl[22] vdd gnd cell_6t
Xbit_r23_c122 bl[122] br[122] wl[23] vdd gnd cell_6t
Xbit_r24_c122 bl[122] br[122] wl[24] vdd gnd cell_6t
Xbit_r25_c122 bl[122] br[122] wl[25] vdd gnd cell_6t
Xbit_r26_c122 bl[122] br[122] wl[26] vdd gnd cell_6t
Xbit_r27_c122 bl[122] br[122] wl[27] vdd gnd cell_6t
Xbit_r28_c122 bl[122] br[122] wl[28] vdd gnd cell_6t
Xbit_r29_c122 bl[122] br[122] wl[29] vdd gnd cell_6t
Xbit_r30_c122 bl[122] br[122] wl[30] vdd gnd cell_6t
Xbit_r31_c122 bl[122] br[122] wl[31] vdd gnd cell_6t
Xbit_r32_c122 bl[122] br[122] wl[32] vdd gnd cell_6t
Xbit_r33_c122 bl[122] br[122] wl[33] vdd gnd cell_6t
Xbit_r34_c122 bl[122] br[122] wl[34] vdd gnd cell_6t
Xbit_r35_c122 bl[122] br[122] wl[35] vdd gnd cell_6t
Xbit_r36_c122 bl[122] br[122] wl[36] vdd gnd cell_6t
Xbit_r37_c122 bl[122] br[122] wl[37] vdd gnd cell_6t
Xbit_r38_c122 bl[122] br[122] wl[38] vdd gnd cell_6t
Xbit_r39_c122 bl[122] br[122] wl[39] vdd gnd cell_6t
Xbit_r40_c122 bl[122] br[122] wl[40] vdd gnd cell_6t
Xbit_r41_c122 bl[122] br[122] wl[41] vdd gnd cell_6t
Xbit_r42_c122 bl[122] br[122] wl[42] vdd gnd cell_6t
Xbit_r43_c122 bl[122] br[122] wl[43] vdd gnd cell_6t
Xbit_r44_c122 bl[122] br[122] wl[44] vdd gnd cell_6t
Xbit_r45_c122 bl[122] br[122] wl[45] vdd gnd cell_6t
Xbit_r46_c122 bl[122] br[122] wl[46] vdd gnd cell_6t
Xbit_r47_c122 bl[122] br[122] wl[47] vdd gnd cell_6t
Xbit_r48_c122 bl[122] br[122] wl[48] vdd gnd cell_6t
Xbit_r49_c122 bl[122] br[122] wl[49] vdd gnd cell_6t
Xbit_r50_c122 bl[122] br[122] wl[50] vdd gnd cell_6t
Xbit_r51_c122 bl[122] br[122] wl[51] vdd gnd cell_6t
Xbit_r52_c122 bl[122] br[122] wl[52] vdd gnd cell_6t
Xbit_r53_c122 bl[122] br[122] wl[53] vdd gnd cell_6t
Xbit_r54_c122 bl[122] br[122] wl[54] vdd gnd cell_6t
Xbit_r55_c122 bl[122] br[122] wl[55] vdd gnd cell_6t
Xbit_r56_c122 bl[122] br[122] wl[56] vdd gnd cell_6t
Xbit_r57_c122 bl[122] br[122] wl[57] vdd gnd cell_6t
Xbit_r58_c122 bl[122] br[122] wl[58] vdd gnd cell_6t
Xbit_r59_c122 bl[122] br[122] wl[59] vdd gnd cell_6t
Xbit_r60_c122 bl[122] br[122] wl[60] vdd gnd cell_6t
Xbit_r61_c122 bl[122] br[122] wl[61] vdd gnd cell_6t
Xbit_r62_c122 bl[122] br[122] wl[62] vdd gnd cell_6t
Xbit_r63_c122 bl[122] br[122] wl[63] vdd gnd cell_6t
Xbit_r64_c122 bl[122] br[122] wl[64] vdd gnd cell_6t
Xbit_r65_c122 bl[122] br[122] wl[65] vdd gnd cell_6t
Xbit_r66_c122 bl[122] br[122] wl[66] vdd gnd cell_6t
Xbit_r67_c122 bl[122] br[122] wl[67] vdd gnd cell_6t
Xbit_r68_c122 bl[122] br[122] wl[68] vdd gnd cell_6t
Xbit_r69_c122 bl[122] br[122] wl[69] vdd gnd cell_6t
Xbit_r70_c122 bl[122] br[122] wl[70] vdd gnd cell_6t
Xbit_r71_c122 bl[122] br[122] wl[71] vdd gnd cell_6t
Xbit_r72_c122 bl[122] br[122] wl[72] vdd gnd cell_6t
Xbit_r73_c122 bl[122] br[122] wl[73] vdd gnd cell_6t
Xbit_r74_c122 bl[122] br[122] wl[74] vdd gnd cell_6t
Xbit_r75_c122 bl[122] br[122] wl[75] vdd gnd cell_6t
Xbit_r76_c122 bl[122] br[122] wl[76] vdd gnd cell_6t
Xbit_r77_c122 bl[122] br[122] wl[77] vdd gnd cell_6t
Xbit_r78_c122 bl[122] br[122] wl[78] vdd gnd cell_6t
Xbit_r79_c122 bl[122] br[122] wl[79] vdd gnd cell_6t
Xbit_r80_c122 bl[122] br[122] wl[80] vdd gnd cell_6t
Xbit_r81_c122 bl[122] br[122] wl[81] vdd gnd cell_6t
Xbit_r82_c122 bl[122] br[122] wl[82] vdd gnd cell_6t
Xbit_r83_c122 bl[122] br[122] wl[83] vdd gnd cell_6t
Xbit_r84_c122 bl[122] br[122] wl[84] vdd gnd cell_6t
Xbit_r85_c122 bl[122] br[122] wl[85] vdd gnd cell_6t
Xbit_r86_c122 bl[122] br[122] wl[86] vdd gnd cell_6t
Xbit_r87_c122 bl[122] br[122] wl[87] vdd gnd cell_6t
Xbit_r88_c122 bl[122] br[122] wl[88] vdd gnd cell_6t
Xbit_r89_c122 bl[122] br[122] wl[89] vdd gnd cell_6t
Xbit_r90_c122 bl[122] br[122] wl[90] vdd gnd cell_6t
Xbit_r91_c122 bl[122] br[122] wl[91] vdd gnd cell_6t
Xbit_r92_c122 bl[122] br[122] wl[92] vdd gnd cell_6t
Xbit_r93_c122 bl[122] br[122] wl[93] vdd gnd cell_6t
Xbit_r94_c122 bl[122] br[122] wl[94] vdd gnd cell_6t
Xbit_r95_c122 bl[122] br[122] wl[95] vdd gnd cell_6t
Xbit_r96_c122 bl[122] br[122] wl[96] vdd gnd cell_6t
Xbit_r97_c122 bl[122] br[122] wl[97] vdd gnd cell_6t
Xbit_r98_c122 bl[122] br[122] wl[98] vdd gnd cell_6t
Xbit_r99_c122 bl[122] br[122] wl[99] vdd gnd cell_6t
Xbit_r100_c122 bl[122] br[122] wl[100] vdd gnd cell_6t
Xbit_r101_c122 bl[122] br[122] wl[101] vdd gnd cell_6t
Xbit_r102_c122 bl[122] br[122] wl[102] vdd gnd cell_6t
Xbit_r103_c122 bl[122] br[122] wl[103] vdd gnd cell_6t
Xbit_r104_c122 bl[122] br[122] wl[104] vdd gnd cell_6t
Xbit_r105_c122 bl[122] br[122] wl[105] vdd gnd cell_6t
Xbit_r106_c122 bl[122] br[122] wl[106] vdd gnd cell_6t
Xbit_r107_c122 bl[122] br[122] wl[107] vdd gnd cell_6t
Xbit_r108_c122 bl[122] br[122] wl[108] vdd gnd cell_6t
Xbit_r109_c122 bl[122] br[122] wl[109] vdd gnd cell_6t
Xbit_r110_c122 bl[122] br[122] wl[110] vdd gnd cell_6t
Xbit_r111_c122 bl[122] br[122] wl[111] vdd gnd cell_6t
Xbit_r112_c122 bl[122] br[122] wl[112] vdd gnd cell_6t
Xbit_r113_c122 bl[122] br[122] wl[113] vdd gnd cell_6t
Xbit_r114_c122 bl[122] br[122] wl[114] vdd gnd cell_6t
Xbit_r115_c122 bl[122] br[122] wl[115] vdd gnd cell_6t
Xbit_r116_c122 bl[122] br[122] wl[116] vdd gnd cell_6t
Xbit_r117_c122 bl[122] br[122] wl[117] vdd gnd cell_6t
Xbit_r118_c122 bl[122] br[122] wl[118] vdd gnd cell_6t
Xbit_r119_c122 bl[122] br[122] wl[119] vdd gnd cell_6t
Xbit_r120_c122 bl[122] br[122] wl[120] vdd gnd cell_6t
Xbit_r121_c122 bl[122] br[122] wl[121] vdd gnd cell_6t
Xbit_r122_c122 bl[122] br[122] wl[122] vdd gnd cell_6t
Xbit_r123_c122 bl[122] br[122] wl[123] vdd gnd cell_6t
Xbit_r124_c122 bl[122] br[122] wl[124] vdd gnd cell_6t
Xbit_r125_c122 bl[122] br[122] wl[125] vdd gnd cell_6t
Xbit_r126_c122 bl[122] br[122] wl[126] vdd gnd cell_6t
Xbit_r127_c122 bl[122] br[122] wl[127] vdd gnd cell_6t
Xbit_r0_c123 bl[123] br[123] wl[0] vdd gnd cell_6t
Xbit_r1_c123 bl[123] br[123] wl[1] vdd gnd cell_6t
Xbit_r2_c123 bl[123] br[123] wl[2] vdd gnd cell_6t
Xbit_r3_c123 bl[123] br[123] wl[3] vdd gnd cell_6t
Xbit_r4_c123 bl[123] br[123] wl[4] vdd gnd cell_6t
Xbit_r5_c123 bl[123] br[123] wl[5] vdd gnd cell_6t
Xbit_r6_c123 bl[123] br[123] wl[6] vdd gnd cell_6t
Xbit_r7_c123 bl[123] br[123] wl[7] vdd gnd cell_6t
Xbit_r8_c123 bl[123] br[123] wl[8] vdd gnd cell_6t
Xbit_r9_c123 bl[123] br[123] wl[9] vdd gnd cell_6t
Xbit_r10_c123 bl[123] br[123] wl[10] vdd gnd cell_6t
Xbit_r11_c123 bl[123] br[123] wl[11] vdd gnd cell_6t
Xbit_r12_c123 bl[123] br[123] wl[12] vdd gnd cell_6t
Xbit_r13_c123 bl[123] br[123] wl[13] vdd gnd cell_6t
Xbit_r14_c123 bl[123] br[123] wl[14] vdd gnd cell_6t
Xbit_r15_c123 bl[123] br[123] wl[15] vdd gnd cell_6t
Xbit_r16_c123 bl[123] br[123] wl[16] vdd gnd cell_6t
Xbit_r17_c123 bl[123] br[123] wl[17] vdd gnd cell_6t
Xbit_r18_c123 bl[123] br[123] wl[18] vdd gnd cell_6t
Xbit_r19_c123 bl[123] br[123] wl[19] vdd gnd cell_6t
Xbit_r20_c123 bl[123] br[123] wl[20] vdd gnd cell_6t
Xbit_r21_c123 bl[123] br[123] wl[21] vdd gnd cell_6t
Xbit_r22_c123 bl[123] br[123] wl[22] vdd gnd cell_6t
Xbit_r23_c123 bl[123] br[123] wl[23] vdd gnd cell_6t
Xbit_r24_c123 bl[123] br[123] wl[24] vdd gnd cell_6t
Xbit_r25_c123 bl[123] br[123] wl[25] vdd gnd cell_6t
Xbit_r26_c123 bl[123] br[123] wl[26] vdd gnd cell_6t
Xbit_r27_c123 bl[123] br[123] wl[27] vdd gnd cell_6t
Xbit_r28_c123 bl[123] br[123] wl[28] vdd gnd cell_6t
Xbit_r29_c123 bl[123] br[123] wl[29] vdd gnd cell_6t
Xbit_r30_c123 bl[123] br[123] wl[30] vdd gnd cell_6t
Xbit_r31_c123 bl[123] br[123] wl[31] vdd gnd cell_6t
Xbit_r32_c123 bl[123] br[123] wl[32] vdd gnd cell_6t
Xbit_r33_c123 bl[123] br[123] wl[33] vdd gnd cell_6t
Xbit_r34_c123 bl[123] br[123] wl[34] vdd gnd cell_6t
Xbit_r35_c123 bl[123] br[123] wl[35] vdd gnd cell_6t
Xbit_r36_c123 bl[123] br[123] wl[36] vdd gnd cell_6t
Xbit_r37_c123 bl[123] br[123] wl[37] vdd gnd cell_6t
Xbit_r38_c123 bl[123] br[123] wl[38] vdd gnd cell_6t
Xbit_r39_c123 bl[123] br[123] wl[39] vdd gnd cell_6t
Xbit_r40_c123 bl[123] br[123] wl[40] vdd gnd cell_6t
Xbit_r41_c123 bl[123] br[123] wl[41] vdd gnd cell_6t
Xbit_r42_c123 bl[123] br[123] wl[42] vdd gnd cell_6t
Xbit_r43_c123 bl[123] br[123] wl[43] vdd gnd cell_6t
Xbit_r44_c123 bl[123] br[123] wl[44] vdd gnd cell_6t
Xbit_r45_c123 bl[123] br[123] wl[45] vdd gnd cell_6t
Xbit_r46_c123 bl[123] br[123] wl[46] vdd gnd cell_6t
Xbit_r47_c123 bl[123] br[123] wl[47] vdd gnd cell_6t
Xbit_r48_c123 bl[123] br[123] wl[48] vdd gnd cell_6t
Xbit_r49_c123 bl[123] br[123] wl[49] vdd gnd cell_6t
Xbit_r50_c123 bl[123] br[123] wl[50] vdd gnd cell_6t
Xbit_r51_c123 bl[123] br[123] wl[51] vdd gnd cell_6t
Xbit_r52_c123 bl[123] br[123] wl[52] vdd gnd cell_6t
Xbit_r53_c123 bl[123] br[123] wl[53] vdd gnd cell_6t
Xbit_r54_c123 bl[123] br[123] wl[54] vdd gnd cell_6t
Xbit_r55_c123 bl[123] br[123] wl[55] vdd gnd cell_6t
Xbit_r56_c123 bl[123] br[123] wl[56] vdd gnd cell_6t
Xbit_r57_c123 bl[123] br[123] wl[57] vdd gnd cell_6t
Xbit_r58_c123 bl[123] br[123] wl[58] vdd gnd cell_6t
Xbit_r59_c123 bl[123] br[123] wl[59] vdd gnd cell_6t
Xbit_r60_c123 bl[123] br[123] wl[60] vdd gnd cell_6t
Xbit_r61_c123 bl[123] br[123] wl[61] vdd gnd cell_6t
Xbit_r62_c123 bl[123] br[123] wl[62] vdd gnd cell_6t
Xbit_r63_c123 bl[123] br[123] wl[63] vdd gnd cell_6t
Xbit_r64_c123 bl[123] br[123] wl[64] vdd gnd cell_6t
Xbit_r65_c123 bl[123] br[123] wl[65] vdd gnd cell_6t
Xbit_r66_c123 bl[123] br[123] wl[66] vdd gnd cell_6t
Xbit_r67_c123 bl[123] br[123] wl[67] vdd gnd cell_6t
Xbit_r68_c123 bl[123] br[123] wl[68] vdd gnd cell_6t
Xbit_r69_c123 bl[123] br[123] wl[69] vdd gnd cell_6t
Xbit_r70_c123 bl[123] br[123] wl[70] vdd gnd cell_6t
Xbit_r71_c123 bl[123] br[123] wl[71] vdd gnd cell_6t
Xbit_r72_c123 bl[123] br[123] wl[72] vdd gnd cell_6t
Xbit_r73_c123 bl[123] br[123] wl[73] vdd gnd cell_6t
Xbit_r74_c123 bl[123] br[123] wl[74] vdd gnd cell_6t
Xbit_r75_c123 bl[123] br[123] wl[75] vdd gnd cell_6t
Xbit_r76_c123 bl[123] br[123] wl[76] vdd gnd cell_6t
Xbit_r77_c123 bl[123] br[123] wl[77] vdd gnd cell_6t
Xbit_r78_c123 bl[123] br[123] wl[78] vdd gnd cell_6t
Xbit_r79_c123 bl[123] br[123] wl[79] vdd gnd cell_6t
Xbit_r80_c123 bl[123] br[123] wl[80] vdd gnd cell_6t
Xbit_r81_c123 bl[123] br[123] wl[81] vdd gnd cell_6t
Xbit_r82_c123 bl[123] br[123] wl[82] vdd gnd cell_6t
Xbit_r83_c123 bl[123] br[123] wl[83] vdd gnd cell_6t
Xbit_r84_c123 bl[123] br[123] wl[84] vdd gnd cell_6t
Xbit_r85_c123 bl[123] br[123] wl[85] vdd gnd cell_6t
Xbit_r86_c123 bl[123] br[123] wl[86] vdd gnd cell_6t
Xbit_r87_c123 bl[123] br[123] wl[87] vdd gnd cell_6t
Xbit_r88_c123 bl[123] br[123] wl[88] vdd gnd cell_6t
Xbit_r89_c123 bl[123] br[123] wl[89] vdd gnd cell_6t
Xbit_r90_c123 bl[123] br[123] wl[90] vdd gnd cell_6t
Xbit_r91_c123 bl[123] br[123] wl[91] vdd gnd cell_6t
Xbit_r92_c123 bl[123] br[123] wl[92] vdd gnd cell_6t
Xbit_r93_c123 bl[123] br[123] wl[93] vdd gnd cell_6t
Xbit_r94_c123 bl[123] br[123] wl[94] vdd gnd cell_6t
Xbit_r95_c123 bl[123] br[123] wl[95] vdd gnd cell_6t
Xbit_r96_c123 bl[123] br[123] wl[96] vdd gnd cell_6t
Xbit_r97_c123 bl[123] br[123] wl[97] vdd gnd cell_6t
Xbit_r98_c123 bl[123] br[123] wl[98] vdd gnd cell_6t
Xbit_r99_c123 bl[123] br[123] wl[99] vdd gnd cell_6t
Xbit_r100_c123 bl[123] br[123] wl[100] vdd gnd cell_6t
Xbit_r101_c123 bl[123] br[123] wl[101] vdd gnd cell_6t
Xbit_r102_c123 bl[123] br[123] wl[102] vdd gnd cell_6t
Xbit_r103_c123 bl[123] br[123] wl[103] vdd gnd cell_6t
Xbit_r104_c123 bl[123] br[123] wl[104] vdd gnd cell_6t
Xbit_r105_c123 bl[123] br[123] wl[105] vdd gnd cell_6t
Xbit_r106_c123 bl[123] br[123] wl[106] vdd gnd cell_6t
Xbit_r107_c123 bl[123] br[123] wl[107] vdd gnd cell_6t
Xbit_r108_c123 bl[123] br[123] wl[108] vdd gnd cell_6t
Xbit_r109_c123 bl[123] br[123] wl[109] vdd gnd cell_6t
Xbit_r110_c123 bl[123] br[123] wl[110] vdd gnd cell_6t
Xbit_r111_c123 bl[123] br[123] wl[111] vdd gnd cell_6t
Xbit_r112_c123 bl[123] br[123] wl[112] vdd gnd cell_6t
Xbit_r113_c123 bl[123] br[123] wl[113] vdd gnd cell_6t
Xbit_r114_c123 bl[123] br[123] wl[114] vdd gnd cell_6t
Xbit_r115_c123 bl[123] br[123] wl[115] vdd gnd cell_6t
Xbit_r116_c123 bl[123] br[123] wl[116] vdd gnd cell_6t
Xbit_r117_c123 bl[123] br[123] wl[117] vdd gnd cell_6t
Xbit_r118_c123 bl[123] br[123] wl[118] vdd gnd cell_6t
Xbit_r119_c123 bl[123] br[123] wl[119] vdd gnd cell_6t
Xbit_r120_c123 bl[123] br[123] wl[120] vdd gnd cell_6t
Xbit_r121_c123 bl[123] br[123] wl[121] vdd gnd cell_6t
Xbit_r122_c123 bl[123] br[123] wl[122] vdd gnd cell_6t
Xbit_r123_c123 bl[123] br[123] wl[123] vdd gnd cell_6t
Xbit_r124_c123 bl[123] br[123] wl[124] vdd gnd cell_6t
Xbit_r125_c123 bl[123] br[123] wl[125] vdd gnd cell_6t
Xbit_r126_c123 bl[123] br[123] wl[126] vdd gnd cell_6t
Xbit_r127_c123 bl[123] br[123] wl[127] vdd gnd cell_6t
Xbit_r0_c124 bl[124] br[124] wl[0] vdd gnd cell_6t
Xbit_r1_c124 bl[124] br[124] wl[1] vdd gnd cell_6t
Xbit_r2_c124 bl[124] br[124] wl[2] vdd gnd cell_6t
Xbit_r3_c124 bl[124] br[124] wl[3] vdd gnd cell_6t
Xbit_r4_c124 bl[124] br[124] wl[4] vdd gnd cell_6t
Xbit_r5_c124 bl[124] br[124] wl[5] vdd gnd cell_6t
Xbit_r6_c124 bl[124] br[124] wl[6] vdd gnd cell_6t
Xbit_r7_c124 bl[124] br[124] wl[7] vdd gnd cell_6t
Xbit_r8_c124 bl[124] br[124] wl[8] vdd gnd cell_6t
Xbit_r9_c124 bl[124] br[124] wl[9] vdd gnd cell_6t
Xbit_r10_c124 bl[124] br[124] wl[10] vdd gnd cell_6t
Xbit_r11_c124 bl[124] br[124] wl[11] vdd gnd cell_6t
Xbit_r12_c124 bl[124] br[124] wl[12] vdd gnd cell_6t
Xbit_r13_c124 bl[124] br[124] wl[13] vdd gnd cell_6t
Xbit_r14_c124 bl[124] br[124] wl[14] vdd gnd cell_6t
Xbit_r15_c124 bl[124] br[124] wl[15] vdd gnd cell_6t
Xbit_r16_c124 bl[124] br[124] wl[16] vdd gnd cell_6t
Xbit_r17_c124 bl[124] br[124] wl[17] vdd gnd cell_6t
Xbit_r18_c124 bl[124] br[124] wl[18] vdd gnd cell_6t
Xbit_r19_c124 bl[124] br[124] wl[19] vdd gnd cell_6t
Xbit_r20_c124 bl[124] br[124] wl[20] vdd gnd cell_6t
Xbit_r21_c124 bl[124] br[124] wl[21] vdd gnd cell_6t
Xbit_r22_c124 bl[124] br[124] wl[22] vdd gnd cell_6t
Xbit_r23_c124 bl[124] br[124] wl[23] vdd gnd cell_6t
Xbit_r24_c124 bl[124] br[124] wl[24] vdd gnd cell_6t
Xbit_r25_c124 bl[124] br[124] wl[25] vdd gnd cell_6t
Xbit_r26_c124 bl[124] br[124] wl[26] vdd gnd cell_6t
Xbit_r27_c124 bl[124] br[124] wl[27] vdd gnd cell_6t
Xbit_r28_c124 bl[124] br[124] wl[28] vdd gnd cell_6t
Xbit_r29_c124 bl[124] br[124] wl[29] vdd gnd cell_6t
Xbit_r30_c124 bl[124] br[124] wl[30] vdd gnd cell_6t
Xbit_r31_c124 bl[124] br[124] wl[31] vdd gnd cell_6t
Xbit_r32_c124 bl[124] br[124] wl[32] vdd gnd cell_6t
Xbit_r33_c124 bl[124] br[124] wl[33] vdd gnd cell_6t
Xbit_r34_c124 bl[124] br[124] wl[34] vdd gnd cell_6t
Xbit_r35_c124 bl[124] br[124] wl[35] vdd gnd cell_6t
Xbit_r36_c124 bl[124] br[124] wl[36] vdd gnd cell_6t
Xbit_r37_c124 bl[124] br[124] wl[37] vdd gnd cell_6t
Xbit_r38_c124 bl[124] br[124] wl[38] vdd gnd cell_6t
Xbit_r39_c124 bl[124] br[124] wl[39] vdd gnd cell_6t
Xbit_r40_c124 bl[124] br[124] wl[40] vdd gnd cell_6t
Xbit_r41_c124 bl[124] br[124] wl[41] vdd gnd cell_6t
Xbit_r42_c124 bl[124] br[124] wl[42] vdd gnd cell_6t
Xbit_r43_c124 bl[124] br[124] wl[43] vdd gnd cell_6t
Xbit_r44_c124 bl[124] br[124] wl[44] vdd gnd cell_6t
Xbit_r45_c124 bl[124] br[124] wl[45] vdd gnd cell_6t
Xbit_r46_c124 bl[124] br[124] wl[46] vdd gnd cell_6t
Xbit_r47_c124 bl[124] br[124] wl[47] vdd gnd cell_6t
Xbit_r48_c124 bl[124] br[124] wl[48] vdd gnd cell_6t
Xbit_r49_c124 bl[124] br[124] wl[49] vdd gnd cell_6t
Xbit_r50_c124 bl[124] br[124] wl[50] vdd gnd cell_6t
Xbit_r51_c124 bl[124] br[124] wl[51] vdd gnd cell_6t
Xbit_r52_c124 bl[124] br[124] wl[52] vdd gnd cell_6t
Xbit_r53_c124 bl[124] br[124] wl[53] vdd gnd cell_6t
Xbit_r54_c124 bl[124] br[124] wl[54] vdd gnd cell_6t
Xbit_r55_c124 bl[124] br[124] wl[55] vdd gnd cell_6t
Xbit_r56_c124 bl[124] br[124] wl[56] vdd gnd cell_6t
Xbit_r57_c124 bl[124] br[124] wl[57] vdd gnd cell_6t
Xbit_r58_c124 bl[124] br[124] wl[58] vdd gnd cell_6t
Xbit_r59_c124 bl[124] br[124] wl[59] vdd gnd cell_6t
Xbit_r60_c124 bl[124] br[124] wl[60] vdd gnd cell_6t
Xbit_r61_c124 bl[124] br[124] wl[61] vdd gnd cell_6t
Xbit_r62_c124 bl[124] br[124] wl[62] vdd gnd cell_6t
Xbit_r63_c124 bl[124] br[124] wl[63] vdd gnd cell_6t
Xbit_r64_c124 bl[124] br[124] wl[64] vdd gnd cell_6t
Xbit_r65_c124 bl[124] br[124] wl[65] vdd gnd cell_6t
Xbit_r66_c124 bl[124] br[124] wl[66] vdd gnd cell_6t
Xbit_r67_c124 bl[124] br[124] wl[67] vdd gnd cell_6t
Xbit_r68_c124 bl[124] br[124] wl[68] vdd gnd cell_6t
Xbit_r69_c124 bl[124] br[124] wl[69] vdd gnd cell_6t
Xbit_r70_c124 bl[124] br[124] wl[70] vdd gnd cell_6t
Xbit_r71_c124 bl[124] br[124] wl[71] vdd gnd cell_6t
Xbit_r72_c124 bl[124] br[124] wl[72] vdd gnd cell_6t
Xbit_r73_c124 bl[124] br[124] wl[73] vdd gnd cell_6t
Xbit_r74_c124 bl[124] br[124] wl[74] vdd gnd cell_6t
Xbit_r75_c124 bl[124] br[124] wl[75] vdd gnd cell_6t
Xbit_r76_c124 bl[124] br[124] wl[76] vdd gnd cell_6t
Xbit_r77_c124 bl[124] br[124] wl[77] vdd gnd cell_6t
Xbit_r78_c124 bl[124] br[124] wl[78] vdd gnd cell_6t
Xbit_r79_c124 bl[124] br[124] wl[79] vdd gnd cell_6t
Xbit_r80_c124 bl[124] br[124] wl[80] vdd gnd cell_6t
Xbit_r81_c124 bl[124] br[124] wl[81] vdd gnd cell_6t
Xbit_r82_c124 bl[124] br[124] wl[82] vdd gnd cell_6t
Xbit_r83_c124 bl[124] br[124] wl[83] vdd gnd cell_6t
Xbit_r84_c124 bl[124] br[124] wl[84] vdd gnd cell_6t
Xbit_r85_c124 bl[124] br[124] wl[85] vdd gnd cell_6t
Xbit_r86_c124 bl[124] br[124] wl[86] vdd gnd cell_6t
Xbit_r87_c124 bl[124] br[124] wl[87] vdd gnd cell_6t
Xbit_r88_c124 bl[124] br[124] wl[88] vdd gnd cell_6t
Xbit_r89_c124 bl[124] br[124] wl[89] vdd gnd cell_6t
Xbit_r90_c124 bl[124] br[124] wl[90] vdd gnd cell_6t
Xbit_r91_c124 bl[124] br[124] wl[91] vdd gnd cell_6t
Xbit_r92_c124 bl[124] br[124] wl[92] vdd gnd cell_6t
Xbit_r93_c124 bl[124] br[124] wl[93] vdd gnd cell_6t
Xbit_r94_c124 bl[124] br[124] wl[94] vdd gnd cell_6t
Xbit_r95_c124 bl[124] br[124] wl[95] vdd gnd cell_6t
Xbit_r96_c124 bl[124] br[124] wl[96] vdd gnd cell_6t
Xbit_r97_c124 bl[124] br[124] wl[97] vdd gnd cell_6t
Xbit_r98_c124 bl[124] br[124] wl[98] vdd gnd cell_6t
Xbit_r99_c124 bl[124] br[124] wl[99] vdd gnd cell_6t
Xbit_r100_c124 bl[124] br[124] wl[100] vdd gnd cell_6t
Xbit_r101_c124 bl[124] br[124] wl[101] vdd gnd cell_6t
Xbit_r102_c124 bl[124] br[124] wl[102] vdd gnd cell_6t
Xbit_r103_c124 bl[124] br[124] wl[103] vdd gnd cell_6t
Xbit_r104_c124 bl[124] br[124] wl[104] vdd gnd cell_6t
Xbit_r105_c124 bl[124] br[124] wl[105] vdd gnd cell_6t
Xbit_r106_c124 bl[124] br[124] wl[106] vdd gnd cell_6t
Xbit_r107_c124 bl[124] br[124] wl[107] vdd gnd cell_6t
Xbit_r108_c124 bl[124] br[124] wl[108] vdd gnd cell_6t
Xbit_r109_c124 bl[124] br[124] wl[109] vdd gnd cell_6t
Xbit_r110_c124 bl[124] br[124] wl[110] vdd gnd cell_6t
Xbit_r111_c124 bl[124] br[124] wl[111] vdd gnd cell_6t
Xbit_r112_c124 bl[124] br[124] wl[112] vdd gnd cell_6t
Xbit_r113_c124 bl[124] br[124] wl[113] vdd gnd cell_6t
Xbit_r114_c124 bl[124] br[124] wl[114] vdd gnd cell_6t
Xbit_r115_c124 bl[124] br[124] wl[115] vdd gnd cell_6t
Xbit_r116_c124 bl[124] br[124] wl[116] vdd gnd cell_6t
Xbit_r117_c124 bl[124] br[124] wl[117] vdd gnd cell_6t
Xbit_r118_c124 bl[124] br[124] wl[118] vdd gnd cell_6t
Xbit_r119_c124 bl[124] br[124] wl[119] vdd gnd cell_6t
Xbit_r120_c124 bl[124] br[124] wl[120] vdd gnd cell_6t
Xbit_r121_c124 bl[124] br[124] wl[121] vdd gnd cell_6t
Xbit_r122_c124 bl[124] br[124] wl[122] vdd gnd cell_6t
Xbit_r123_c124 bl[124] br[124] wl[123] vdd gnd cell_6t
Xbit_r124_c124 bl[124] br[124] wl[124] vdd gnd cell_6t
Xbit_r125_c124 bl[124] br[124] wl[125] vdd gnd cell_6t
Xbit_r126_c124 bl[124] br[124] wl[126] vdd gnd cell_6t
Xbit_r127_c124 bl[124] br[124] wl[127] vdd gnd cell_6t
Xbit_r0_c125 bl[125] br[125] wl[0] vdd gnd cell_6t
Xbit_r1_c125 bl[125] br[125] wl[1] vdd gnd cell_6t
Xbit_r2_c125 bl[125] br[125] wl[2] vdd gnd cell_6t
Xbit_r3_c125 bl[125] br[125] wl[3] vdd gnd cell_6t
Xbit_r4_c125 bl[125] br[125] wl[4] vdd gnd cell_6t
Xbit_r5_c125 bl[125] br[125] wl[5] vdd gnd cell_6t
Xbit_r6_c125 bl[125] br[125] wl[6] vdd gnd cell_6t
Xbit_r7_c125 bl[125] br[125] wl[7] vdd gnd cell_6t
Xbit_r8_c125 bl[125] br[125] wl[8] vdd gnd cell_6t
Xbit_r9_c125 bl[125] br[125] wl[9] vdd gnd cell_6t
Xbit_r10_c125 bl[125] br[125] wl[10] vdd gnd cell_6t
Xbit_r11_c125 bl[125] br[125] wl[11] vdd gnd cell_6t
Xbit_r12_c125 bl[125] br[125] wl[12] vdd gnd cell_6t
Xbit_r13_c125 bl[125] br[125] wl[13] vdd gnd cell_6t
Xbit_r14_c125 bl[125] br[125] wl[14] vdd gnd cell_6t
Xbit_r15_c125 bl[125] br[125] wl[15] vdd gnd cell_6t
Xbit_r16_c125 bl[125] br[125] wl[16] vdd gnd cell_6t
Xbit_r17_c125 bl[125] br[125] wl[17] vdd gnd cell_6t
Xbit_r18_c125 bl[125] br[125] wl[18] vdd gnd cell_6t
Xbit_r19_c125 bl[125] br[125] wl[19] vdd gnd cell_6t
Xbit_r20_c125 bl[125] br[125] wl[20] vdd gnd cell_6t
Xbit_r21_c125 bl[125] br[125] wl[21] vdd gnd cell_6t
Xbit_r22_c125 bl[125] br[125] wl[22] vdd gnd cell_6t
Xbit_r23_c125 bl[125] br[125] wl[23] vdd gnd cell_6t
Xbit_r24_c125 bl[125] br[125] wl[24] vdd gnd cell_6t
Xbit_r25_c125 bl[125] br[125] wl[25] vdd gnd cell_6t
Xbit_r26_c125 bl[125] br[125] wl[26] vdd gnd cell_6t
Xbit_r27_c125 bl[125] br[125] wl[27] vdd gnd cell_6t
Xbit_r28_c125 bl[125] br[125] wl[28] vdd gnd cell_6t
Xbit_r29_c125 bl[125] br[125] wl[29] vdd gnd cell_6t
Xbit_r30_c125 bl[125] br[125] wl[30] vdd gnd cell_6t
Xbit_r31_c125 bl[125] br[125] wl[31] vdd gnd cell_6t
Xbit_r32_c125 bl[125] br[125] wl[32] vdd gnd cell_6t
Xbit_r33_c125 bl[125] br[125] wl[33] vdd gnd cell_6t
Xbit_r34_c125 bl[125] br[125] wl[34] vdd gnd cell_6t
Xbit_r35_c125 bl[125] br[125] wl[35] vdd gnd cell_6t
Xbit_r36_c125 bl[125] br[125] wl[36] vdd gnd cell_6t
Xbit_r37_c125 bl[125] br[125] wl[37] vdd gnd cell_6t
Xbit_r38_c125 bl[125] br[125] wl[38] vdd gnd cell_6t
Xbit_r39_c125 bl[125] br[125] wl[39] vdd gnd cell_6t
Xbit_r40_c125 bl[125] br[125] wl[40] vdd gnd cell_6t
Xbit_r41_c125 bl[125] br[125] wl[41] vdd gnd cell_6t
Xbit_r42_c125 bl[125] br[125] wl[42] vdd gnd cell_6t
Xbit_r43_c125 bl[125] br[125] wl[43] vdd gnd cell_6t
Xbit_r44_c125 bl[125] br[125] wl[44] vdd gnd cell_6t
Xbit_r45_c125 bl[125] br[125] wl[45] vdd gnd cell_6t
Xbit_r46_c125 bl[125] br[125] wl[46] vdd gnd cell_6t
Xbit_r47_c125 bl[125] br[125] wl[47] vdd gnd cell_6t
Xbit_r48_c125 bl[125] br[125] wl[48] vdd gnd cell_6t
Xbit_r49_c125 bl[125] br[125] wl[49] vdd gnd cell_6t
Xbit_r50_c125 bl[125] br[125] wl[50] vdd gnd cell_6t
Xbit_r51_c125 bl[125] br[125] wl[51] vdd gnd cell_6t
Xbit_r52_c125 bl[125] br[125] wl[52] vdd gnd cell_6t
Xbit_r53_c125 bl[125] br[125] wl[53] vdd gnd cell_6t
Xbit_r54_c125 bl[125] br[125] wl[54] vdd gnd cell_6t
Xbit_r55_c125 bl[125] br[125] wl[55] vdd gnd cell_6t
Xbit_r56_c125 bl[125] br[125] wl[56] vdd gnd cell_6t
Xbit_r57_c125 bl[125] br[125] wl[57] vdd gnd cell_6t
Xbit_r58_c125 bl[125] br[125] wl[58] vdd gnd cell_6t
Xbit_r59_c125 bl[125] br[125] wl[59] vdd gnd cell_6t
Xbit_r60_c125 bl[125] br[125] wl[60] vdd gnd cell_6t
Xbit_r61_c125 bl[125] br[125] wl[61] vdd gnd cell_6t
Xbit_r62_c125 bl[125] br[125] wl[62] vdd gnd cell_6t
Xbit_r63_c125 bl[125] br[125] wl[63] vdd gnd cell_6t
Xbit_r64_c125 bl[125] br[125] wl[64] vdd gnd cell_6t
Xbit_r65_c125 bl[125] br[125] wl[65] vdd gnd cell_6t
Xbit_r66_c125 bl[125] br[125] wl[66] vdd gnd cell_6t
Xbit_r67_c125 bl[125] br[125] wl[67] vdd gnd cell_6t
Xbit_r68_c125 bl[125] br[125] wl[68] vdd gnd cell_6t
Xbit_r69_c125 bl[125] br[125] wl[69] vdd gnd cell_6t
Xbit_r70_c125 bl[125] br[125] wl[70] vdd gnd cell_6t
Xbit_r71_c125 bl[125] br[125] wl[71] vdd gnd cell_6t
Xbit_r72_c125 bl[125] br[125] wl[72] vdd gnd cell_6t
Xbit_r73_c125 bl[125] br[125] wl[73] vdd gnd cell_6t
Xbit_r74_c125 bl[125] br[125] wl[74] vdd gnd cell_6t
Xbit_r75_c125 bl[125] br[125] wl[75] vdd gnd cell_6t
Xbit_r76_c125 bl[125] br[125] wl[76] vdd gnd cell_6t
Xbit_r77_c125 bl[125] br[125] wl[77] vdd gnd cell_6t
Xbit_r78_c125 bl[125] br[125] wl[78] vdd gnd cell_6t
Xbit_r79_c125 bl[125] br[125] wl[79] vdd gnd cell_6t
Xbit_r80_c125 bl[125] br[125] wl[80] vdd gnd cell_6t
Xbit_r81_c125 bl[125] br[125] wl[81] vdd gnd cell_6t
Xbit_r82_c125 bl[125] br[125] wl[82] vdd gnd cell_6t
Xbit_r83_c125 bl[125] br[125] wl[83] vdd gnd cell_6t
Xbit_r84_c125 bl[125] br[125] wl[84] vdd gnd cell_6t
Xbit_r85_c125 bl[125] br[125] wl[85] vdd gnd cell_6t
Xbit_r86_c125 bl[125] br[125] wl[86] vdd gnd cell_6t
Xbit_r87_c125 bl[125] br[125] wl[87] vdd gnd cell_6t
Xbit_r88_c125 bl[125] br[125] wl[88] vdd gnd cell_6t
Xbit_r89_c125 bl[125] br[125] wl[89] vdd gnd cell_6t
Xbit_r90_c125 bl[125] br[125] wl[90] vdd gnd cell_6t
Xbit_r91_c125 bl[125] br[125] wl[91] vdd gnd cell_6t
Xbit_r92_c125 bl[125] br[125] wl[92] vdd gnd cell_6t
Xbit_r93_c125 bl[125] br[125] wl[93] vdd gnd cell_6t
Xbit_r94_c125 bl[125] br[125] wl[94] vdd gnd cell_6t
Xbit_r95_c125 bl[125] br[125] wl[95] vdd gnd cell_6t
Xbit_r96_c125 bl[125] br[125] wl[96] vdd gnd cell_6t
Xbit_r97_c125 bl[125] br[125] wl[97] vdd gnd cell_6t
Xbit_r98_c125 bl[125] br[125] wl[98] vdd gnd cell_6t
Xbit_r99_c125 bl[125] br[125] wl[99] vdd gnd cell_6t
Xbit_r100_c125 bl[125] br[125] wl[100] vdd gnd cell_6t
Xbit_r101_c125 bl[125] br[125] wl[101] vdd gnd cell_6t
Xbit_r102_c125 bl[125] br[125] wl[102] vdd gnd cell_6t
Xbit_r103_c125 bl[125] br[125] wl[103] vdd gnd cell_6t
Xbit_r104_c125 bl[125] br[125] wl[104] vdd gnd cell_6t
Xbit_r105_c125 bl[125] br[125] wl[105] vdd gnd cell_6t
Xbit_r106_c125 bl[125] br[125] wl[106] vdd gnd cell_6t
Xbit_r107_c125 bl[125] br[125] wl[107] vdd gnd cell_6t
Xbit_r108_c125 bl[125] br[125] wl[108] vdd gnd cell_6t
Xbit_r109_c125 bl[125] br[125] wl[109] vdd gnd cell_6t
Xbit_r110_c125 bl[125] br[125] wl[110] vdd gnd cell_6t
Xbit_r111_c125 bl[125] br[125] wl[111] vdd gnd cell_6t
Xbit_r112_c125 bl[125] br[125] wl[112] vdd gnd cell_6t
Xbit_r113_c125 bl[125] br[125] wl[113] vdd gnd cell_6t
Xbit_r114_c125 bl[125] br[125] wl[114] vdd gnd cell_6t
Xbit_r115_c125 bl[125] br[125] wl[115] vdd gnd cell_6t
Xbit_r116_c125 bl[125] br[125] wl[116] vdd gnd cell_6t
Xbit_r117_c125 bl[125] br[125] wl[117] vdd gnd cell_6t
Xbit_r118_c125 bl[125] br[125] wl[118] vdd gnd cell_6t
Xbit_r119_c125 bl[125] br[125] wl[119] vdd gnd cell_6t
Xbit_r120_c125 bl[125] br[125] wl[120] vdd gnd cell_6t
Xbit_r121_c125 bl[125] br[125] wl[121] vdd gnd cell_6t
Xbit_r122_c125 bl[125] br[125] wl[122] vdd gnd cell_6t
Xbit_r123_c125 bl[125] br[125] wl[123] vdd gnd cell_6t
Xbit_r124_c125 bl[125] br[125] wl[124] vdd gnd cell_6t
Xbit_r125_c125 bl[125] br[125] wl[125] vdd gnd cell_6t
Xbit_r126_c125 bl[125] br[125] wl[126] vdd gnd cell_6t
Xbit_r127_c125 bl[125] br[125] wl[127] vdd gnd cell_6t
Xbit_r0_c126 bl[126] br[126] wl[0] vdd gnd cell_6t
Xbit_r1_c126 bl[126] br[126] wl[1] vdd gnd cell_6t
Xbit_r2_c126 bl[126] br[126] wl[2] vdd gnd cell_6t
Xbit_r3_c126 bl[126] br[126] wl[3] vdd gnd cell_6t
Xbit_r4_c126 bl[126] br[126] wl[4] vdd gnd cell_6t
Xbit_r5_c126 bl[126] br[126] wl[5] vdd gnd cell_6t
Xbit_r6_c126 bl[126] br[126] wl[6] vdd gnd cell_6t
Xbit_r7_c126 bl[126] br[126] wl[7] vdd gnd cell_6t
Xbit_r8_c126 bl[126] br[126] wl[8] vdd gnd cell_6t
Xbit_r9_c126 bl[126] br[126] wl[9] vdd gnd cell_6t
Xbit_r10_c126 bl[126] br[126] wl[10] vdd gnd cell_6t
Xbit_r11_c126 bl[126] br[126] wl[11] vdd gnd cell_6t
Xbit_r12_c126 bl[126] br[126] wl[12] vdd gnd cell_6t
Xbit_r13_c126 bl[126] br[126] wl[13] vdd gnd cell_6t
Xbit_r14_c126 bl[126] br[126] wl[14] vdd gnd cell_6t
Xbit_r15_c126 bl[126] br[126] wl[15] vdd gnd cell_6t
Xbit_r16_c126 bl[126] br[126] wl[16] vdd gnd cell_6t
Xbit_r17_c126 bl[126] br[126] wl[17] vdd gnd cell_6t
Xbit_r18_c126 bl[126] br[126] wl[18] vdd gnd cell_6t
Xbit_r19_c126 bl[126] br[126] wl[19] vdd gnd cell_6t
Xbit_r20_c126 bl[126] br[126] wl[20] vdd gnd cell_6t
Xbit_r21_c126 bl[126] br[126] wl[21] vdd gnd cell_6t
Xbit_r22_c126 bl[126] br[126] wl[22] vdd gnd cell_6t
Xbit_r23_c126 bl[126] br[126] wl[23] vdd gnd cell_6t
Xbit_r24_c126 bl[126] br[126] wl[24] vdd gnd cell_6t
Xbit_r25_c126 bl[126] br[126] wl[25] vdd gnd cell_6t
Xbit_r26_c126 bl[126] br[126] wl[26] vdd gnd cell_6t
Xbit_r27_c126 bl[126] br[126] wl[27] vdd gnd cell_6t
Xbit_r28_c126 bl[126] br[126] wl[28] vdd gnd cell_6t
Xbit_r29_c126 bl[126] br[126] wl[29] vdd gnd cell_6t
Xbit_r30_c126 bl[126] br[126] wl[30] vdd gnd cell_6t
Xbit_r31_c126 bl[126] br[126] wl[31] vdd gnd cell_6t
Xbit_r32_c126 bl[126] br[126] wl[32] vdd gnd cell_6t
Xbit_r33_c126 bl[126] br[126] wl[33] vdd gnd cell_6t
Xbit_r34_c126 bl[126] br[126] wl[34] vdd gnd cell_6t
Xbit_r35_c126 bl[126] br[126] wl[35] vdd gnd cell_6t
Xbit_r36_c126 bl[126] br[126] wl[36] vdd gnd cell_6t
Xbit_r37_c126 bl[126] br[126] wl[37] vdd gnd cell_6t
Xbit_r38_c126 bl[126] br[126] wl[38] vdd gnd cell_6t
Xbit_r39_c126 bl[126] br[126] wl[39] vdd gnd cell_6t
Xbit_r40_c126 bl[126] br[126] wl[40] vdd gnd cell_6t
Xbit_r41_c126 bl[126] br[126] wl[41] vdd gnd cell_6t
Xbit_r42_c126 bl[126] br[126] wl[42] vdd gnd cell_6t
Xbit_r43_c126 bl[126] br[126] wl[43] vdd gnd cell_6t
Xbit_r44_c126 bl[126] br[126] wl[44] vdd gnd cell_6t
Xbit_r45_c126 bl[126] br[126] wl[45] vdd gnd cell_6t
Xbit_r46_c126 bl[126] br[126] wl[46] vdd gnd cell_6t
Xbit_r47_c126 bl[126] br[126] wl[47] vdd gnd cell_6t
Xbit_r48_c126 bl[126] br[126] wl[48] vdd gnd cell_6t
Xbit_r49_c126 bl[126] br[126] wl[49] vdd gnd cell_6t
Xbit_r50_c126 bl[126] br[126] wl[50] vdd gnd cell_6t
Xbit_r51_c126 bl[126] br[126] wl[51] vdd gnd cell_6t
Xbit_r52_c126 bl[126] br[126] wl[52] vdd gnd cell_6t
Xbit_r53_c126 bl[126] br[126] wl[53] vdd gnd cell_6t
Xbit_r54_c126 bl[126] br[126] wl[54] vdd gnd cell_6t
Xbit_r55_c126 bl[126] br[126] wl[55] vdd gnd cell_6t
Xbit_r56_c126 bl[126] br[126] wl[56] vdd gnd cell_6t
Xbit_r57_c126 bl[126] br[126] wl[57] vdd gnd cell_6t
Xbit_r58_c126 bl[126] br[126] wl[58] vdd gnd cell_6t
Xbit_r59_c126 bl[126] br[126] wl[59] vdd gnd cell_6t
Xbit_r60_c126 bl[126] br[126] wl[60] vdd gnd cell_6t
Xbit_r61_c126 bl[126] br[126] wl[61] vdd gnd cell_6t
Xbit_r62_c126 bl[126] br[126] wl[62] vdd gnd cell_6t
Xbit_r63_c126 bl[126] br[126] wl[63] vdd gnd cell_6t
Xbit_r64_c126 bl[126] br[126] wl[64] vdd gnd cell_6t
Xbit_r65_c126 bl[126] br[126] wl[65] vdd gnd cell_6t
Xbit_r66_c126 bl[126] br[126] wl[66] vdd gnd cell_6t
Xbit_r67_c126 bl[126] br[126] wl[67] vdd gnd cell_6t
Xbit_r68_c126 bl[126] br[126] wl[68] vdd gnd cell_6t
Xbit_r69_c126 bl[126] br[126] wl[69] vdd gnd cell_6t
Xbit_r70_c126 bl[126] br[126] wl[70] vdd gnd cell_6t
Xbit_r71_c126 bl[126] br[126] wl[71] vdd gnd cell_6t
Xbit_r72_c126 bl[126] br[126] wl[72] vdd gnd cell_6t
Xbit_r73_c126 bl[126] br[126] wl[73] vdd gnd cell_6t
Xbit_r74_c126 bl[126] br[126] wl[74] vdd gnd cell_6t
Xbit_r75_c126 bl[126] br[126] wl[75] vdd gnd cell_6t
Xbit_r76_c126 bl[126] br[126] wl[76] vdd gnd cell_6t
Xbit_r77_c126 bl[126] br[126] wl[77] vdd gnd cell_6t
Xbit_r78_c126 bl[126] br[126] wl[78] vdd gnd cell_6t
Xbit_r79_c126 bl[126] br[126] wl[79] vdd gnd cell_6t
Xbit_r80_c126 bl[126] br[126] wl[80] vdd gnd cell_6t
Xbit_r81_c126 bl[126] br[126] wl[81] vdd gnd cell_6t
Xbit_r82_c126 bl[126] br[126] wl[82] vdd gnd cell_6t
Xbit_r83_c126 bl[126] br[126] wl[83] vdd gnd cell_6t
Xbit_r84_c126 bl[126] br[126] wl[84] vdd gnd cell_6t
Xbit_r85_c126 bl[126] br[126] wl[85] vdd gnd cell_6t
Xbit_r86_c126 bl[126] br[126] wl[86] vdd gnd cell_6t
Xbit_r87_c126 bl[126] br[126] wl[87] vdd gnd cell_6t
Xbit_r88_c126 bl[126] br[126] wl[88] vdd gnd cell_6t
Xbit_r89_c126 bl[126] br[126] wl[89] vdd gnd cell_6t
Xbit_r90_c126 bl[126] br[126] wl[90] vdd gnd cell_6t
Xbit_r91_c126 bl[126] br[126] wl[91] vdd gnd cell_6t
Xbit_r92_c126 bl[126] br[126] wl[92] vdd gnd cell_6t
Xbit_r93_c126 bl[126] br[126] wl[93] vdd gnd cell_6t
Xbit_r94_c126 bl[126] br[126] wl[94] vdd gnd cell_6t
Xbit_r95_c126 bl[126] br[126] wl[95] vdd gnd cell_6t
Xbit_r96_c126 bl[126] br[126] wl[96] vdd gnd cell_6t
Xbit_r97_c126 bl[126] br[126] wl[97] vdd gnd cell_6t
Xbit_r98_c126 bl[126] br[126] wl[98] vdd gnd cell_6t
Xbit_r99_c126 bl[126] br[126] wl[99] vdd gnd cell_6t
Xbit_r100_c126 bl[126] br[126] wl[100] vdd gnd cell_6t
Xbit_r101_c126 bl[126] br[126] wl[101] vdd gnd cell_6t
Xbit_r102_c126 bl[126] br[126] wl[102] vdd gnd cell_6t
Xbit_r103_c126 bl[126] br[126] wl[103] vdd gnd cell_6t
Xbit_r104_c126 bl[126] br[126] wl[104] vdd gnd cell_6t
Xbit_r105_c126 bl[126] br[126] wl[105] vdd gnd cell_6t
Xbit_r106_c126 bl[126] br[126] wl[106] vdd gnd cell_6t
Xbit_r107_c126 bl[126] br[126] wl[107] vdd gnd cell_6t
Xbit_r108_c126 bl[126] br[126] wl[108] vdd gnd cell_6t
Xbit_r109_c126 bl[126] br[126] wl[109] vdd gnd cell_6t
Xbit_r110_c126 bl[126] br[126] wl[110] vdd gnd cell_6t
Xbit_r111_c126 bl[126] br[126] wl[111] vdd gnd cell_6t
Xbit_r112_c126 bl[126] br[126] wl[112] vdd gnd cell_6t
Xbit_r113_c126 bl[126] br[126] wl[113] vdd gnd cell_6t
Xbit_r114_c126 bl[126] br[126] wl[114] vdd gnd cell_6t
Xbit_r115_c126 bl[126] br[126] wl[115] vdd gnd cell_6t
Xbit_r116_c126 bl[126] br[126] wl[116] vdd gnd cell_6t
Xbit_r117_c126 bl[126] br[126] wl[117] vdd gnd cell_6t
Xbit_r118_c126 bl[126] br[126] wl[118] vdd gnd cell_6t
Xbit_r119_c126 bl[126] br[126] wl[119] vdd gnd cell_6t
Xbit_r120_c126 bl[126] br[126] wl[120] vdd gnd cell_6t
Xbit_r121_c126 bl[126] br[126] wl[121] vdd gnd cell_6t
Xbit_r122_c126 bl[126] br[126] wl[122] vdd gnd cell_6t
Xbit_r123_c126 bl[126] br[126] wl[123] vdd gnd cell_6t
Xbit_r124_c126 bl[126] br[126] wl[124] vdd gnd cell_6t
Xbit_r125_c126 bl[126] br[126] wl[125] vdd gnd cell_6t
Xbit_r126_c126 bl[126] br[126] wl[126] vdd gnd cell_6t
Xbit_r127_c126 bl[126] br[126] wl[127] vdd gnd cell_6t
Xbit_r0_c127 bl[127] br[127] wl[0] vdd gnd cell_6t
Xbit_r1_c127 bl[127] br[127] wl[1] vdd gnd cell_6t
Xbit_r2_c127 bl[127] br[127] wl[2] vdd gnd cell_6t
Xbit_r3_c127 bl[127] br[127] wl[3] vdd gnd cell_6t
Xbit_r4_c127 bl[127] br[127] wl[4] vdd gnd cell_6t
Xbit_r5_c127 bl[127] br[127] wl[5] vdd gnd cell_6t
Xbit_r6_c127 bl[127] br[127] wl[6] vdd gnd cell_6t
Xbit_r7_c127 bl[127] br[127] wl[7] vdd gnd cell_6t
Xbit_r8_c127 bl[127] br[127] wl[8] vdd gnd cell_6t
Xbit_r9_c127 bl[127] br[127] wl[9] vdd gnd cell_6t
Xbit_r10_c127 bl[127] br[127] wl[10] vdd gnd cell_6t
Xbit_r11_c127 bl[127] br[127] wl[11] vdd gnd cell_6t
Xbit_r12_c127 bl[127] br[127] wl[12] vdd gnd cell_6t
Xbit_r13_c127 bl[127] br[127] wl[13] vdd gnd cell_6t
Xbit_r14_c127 bl[127] br[127] wl[14] vdd gnd cell_6t
Xbit_r15_c127 bl[127] br[127] wl[15] vdd gnd cell_6t
Xbit_r16_c127 bl[127] br[127] wl[16] vdd gnd cell_6t
Xbit_r17_c127 bl[127] br[127] wl[17] vdd gnd cell_6t
Xbit_r18_c127 bl[127] br[127] wl[18] vdd gnd cell_6t
Xbit_r19_c127 bl[127] br[127] wl[19] vdd gnd cell_6t
Xbit_r20_c127 bl[127] br[127] wl[20] vdd gnd cell_6t
Xbit_r21_c127 bl[127] br[127] wl[21] vdd gnd cell_6t
Xbit_r22_c127 bl[127] br[127] wl[22] vdd gnd cell_6t
Xbit_r23_c127 bl[127] br[127] wl[23] vdd gnd cell_6t
Xbit_r24_c127 bl[127] br[127] wl[24] vdd gnd cell_6t
Xbit_r25_c127 bl[127] br[127] wl[25] vdd gnd cell_6t
Xbit_r26_c127 bl[127] br[127] wl[26] vdd gnd cell_6t
Xbit_r27_c127 bl[127] br[127] wl[27] vdd gnd cell_6t
Xbit_r28_c127 bl[127] br[127] wl[28] vdd gnd cell_6t
Xbit_r29_c127 bl[127] br[127] wl[29] vdd gnd cell_6t
Xbit_r30_c127 bl[127] br[127] wl[30] vdd gnd cell_6t
Xbit_r31_c127 bl[127] br[127] wl[31] vdd gnd cell_6t
Xbit_r32_c127 bl[127] br[127] wl[32] vdd gnd cell_6t
Xbit_r33_c127 bl[127] br[127] wl[33] vdd gnd cell_6t
Xbit_r34_c127 bl[127] br[127] wl[34] vdd gnd cell_6t
Xbit_r35_c127 bl[127] br[127] wl[35] vdd gnd cell_6t
Xbit_r36_c127 bl[127] br[127] wl[36] vdd gnd cell_6t
Xbit_r37_c127 bl[127] br[127] wl[37] vdd gnd cell_6t
Xbit_r38_c127 bl[127] br[127] wl[38] vdd gnd cell_6t
Xbit_r39_c127 bl[127] br[127] wl[39] vdd gnd cell_6t
Xbit_r40_c127 bl[127] br[127] wl[40] vdd gnd cell_6t
Xbit_r41_c127 bl[127] br[127] wl[41] vdd gnd cell_6t
Xbit_r42_c127 bl[127] br[127] wl[42] vdd gnd cell_6t
Xbit_r43_c127 bl[127] br[127] wl[43] vdd gnd cell_6t
Xbit_r44_c127 bl[127] br[127] wl[44] vdd gnd cell_6t
Xbit_r45_c127 bl[127] br[127] wl[45] vdd gnd cell_6t
Xbit_r46_c127 bl[127] br[127] wl[46] vdd gnd cell_6t
Xbit_r47_c127 bl[127] br[127] wl[47] vdd gnd cell_6t
Xbit_r48_c127 bl[127] br[127] wl[48] vdd gnd cell_6t
Xbit_r49_c127 bl[127] br[127] wl[49] vdd gnd cell_6t
Xbit_r50_c127 bl[127] br[127] wl[50] vdd gnd cell_6t
Xbit_r51_c127 bl[127] br[127] wl[51] vdd gnd cell_6t
Xbit_r52_c127 bl[127] br[127] wl[52] vdd gnd cell_6t
Xbit_r53_c127 bl[127] br[127] wl[53] vdd gnd cell_6t
Xbit_r54_c127 bl[127] br[127] wl[54] vdd gnd cell_6t
Xbit_r55_c127 bl[127] br[127] wl[55] vdd gnd cell_6t
Xbit_r56_c127 bl[127] br[127] wl[56] vdd gnd cell_6t
Xbit_r57_c127 bl[127] br[127] wl[57] vdd gnd cell_6t
Xbit_r58_c127 bl[127] br[127] wl[58] vdd gnd cell_6t
Xbit_r59_c127 bl[127] br[127] wl[59] vdd gnd cell_6t
Xbit_r60_c127 bl[127] br[127] wl[60] vdd gnd cell_6t
Xbit_r61_c127 bl[127] br[127] wl[61] vdd gnd cell_6t
Xbit_r62_c127 bl[127] br[127] wl[62] vdd gnd cell_6t
Xbit_r63_c127 bl[127] br[127] wl[63] vdd gnd cell_6t
Xbit_r64_c127 bl[127] br[127] wl[64] vdd gnd cell_6t
Xbit_r65_c127 bl[127] br[127] wl[65] vdd gnd cell_6t
Xbit_r66_c127 bl[127] br[127] wl[66] vdd gnd cell_6t
Xbit_r67_c127 bl[127] br[127] wl[67] vdd gnd cell_6t
Xbit_r68_c127 bl[127] br[127] wl[68] vdd gnd cell_6t
Xbit_r69_c127 bl[127] br[127] wl[69] vdd gnd cell_6t
Xbit_r70_c127 bl[127] br[127] wl[70] vdd gnd cell_6t
Xbit_r71_c127 bl[127] br[127] wl[71] vdd gnd cell_6t
Xbit_r72_c127 bl[127] br[127] wl[72] vdd gnd cell_6t
Xbit_r73_c127 bl[127] br[127] wl[73] vdd gnd cell_6t
Xbit_r74_c127 bl[127] br[127] wl[74] vdd gnd cell_6t
Xbit_r75_c127 bl[127] br[127] wl[75] vdd gnd cell_6t
Xbit_r76_c127 bl[127] br[127] wl[76] vdd gnd cell_6t
Xbit_r77_c127 bl[127] br[127] wl[77] vdd gnd cell_6t
Xbit_r78_c127 bl[127] br[127] wl[78] vdd gnd cell_6t
Xbit_r79_c127 bl[127] br[127] wl[79] vdd gnd cell_6t
Xbit_r80_c127 bl[127] br[127] wl[80] vdd gnd cell_6t
Xbit_r81_c127 bl[127] br[127] wl[81] vdd gnd cell_6t
Xbit_r82_c127 bl[127] br[127] wl[82] vdd gnd cell_6t
Xbit_r83_c127 bl[127] br[127] wl[83] vdd gnd cell_6t
Xbit_r84_c127 bl[127] br[127] wl[84] vdd gnd cell_6t
Xbit_r85_c127 bl[127] br[127] wl[85] vdd gnd cell_6t
Xbit_r86_c127 bl[127] br[127] wl[86] vdd gnd cell_6t
Xbit_r87_c127 bl[127] br[127] wl[87] vdd gnd cell_6t
Xbit_r88_c127 bl[127] br[127] wl[88] vdd gnd cell_6t
Xbit_r89_c127 bl[127] br[127] wl[89] vdd gnd cell_6t
Xbit_r90_c127 bl[127] br[127] wl[90] vdd gnd cell_6t
Xbit_r91_c127 bl[127] br[127] wl[91] vdd gnd cell_6t
Xbit_r92_c127 bl[127] br[127] wl[92] vdd gnd cell_6t
Xbit_r93_c127 bl[127] br[127] wl[93] vdd gnd cell_6t
Xbit_r94_c127 bl[127] br[127] wl[94] vdd gnd cell_6t
Xbit_r95_c127 bl[127] br[127] wl[95] vdd gnd cell_6t
Xbit_r96_c127 bl[127] br[127] wl[96] vdd gnd cell_6t
Xbit_r97_c127 bl[127] br[127] wl[97] vdd gnd cell_6t
Xbit_r98_c127 bl[127] br[127] wl[98] vdd gnd cell_6t
Xbit_r99_c127 bl[127] br[127] wl[99] vdd gnd cell_6t
Xbit_r100_c127 bl[127] br[127] wl[100] vdd gnd cell_6t
Xbit_r101_c127 bl[127] br[127] wl[101] vdd gnd cell_6t
Xbit_r102_c127 bl[127] br[127] wl[102] vdd gnd cell_6t
Xbit_r103_c127 bl[127] br[127] wl[103] vdd gnd cell_6t
Xbit_r104_c127 bl[127] br[127] wl[104] vdd gnd cell_6t
Xbit_r105_c127 bl[127] br[127] wl[105] vdd gnd cell_6t
Xbit_r106_c127 bl[127] br[127] wl[106] vdd gnd cell_6t
Xbit_r107_c127 bl[127] br[127] wl[107] vdd gnd cell_6t
Xbit_r108_c127 bl[127] br[127] wl[108] vdd gnd cell_6t
Xbit_r109_c127 bl[127] br[127] wl[109] vdd gnd cell_6t
Xbit_r110_c127 bl[127] br[127] wl[110] vdd gnd cell_6t
Xbit_r111_c127 bl[127] br[127] wl[111] vdd gnd cell_6t
Xbit_r112_c127 bl[127] br[127] wl[112] vdd gnd cell_6t
Xbit_r113_c127 bl[127] br[127] wl[113] vdd gnd cell_6t
Xbit_r114_c127 bl[127] br[127] wl[114] vdd gnd cell_6t
Xbit_r115_c127 bl[127] br[127] wl[115] vdd gnd cell_6t
Xbit_r116_c127 bl[127] br[127] wl[116] vdd gnd cell_6t
Xbit_r117_c127 bl[127] br[127] wl[117] vdd gnd cell_6t
Xbit_r118_c127 bl[127] br[127] wl[118] vdd gnd cell_6t
Xbit_r119_c127 bl[127] br[127] wl[119] vdd gnd cell_6t
Xbit_r120_c127 bl[127] br[127] wl[120] vdd gnd cell_6t
Xbit_r121_c127 bl[127] br[127] wl[121] vdd gnd cell_6t
Xbit_r122_c127 bl[127] br[127] wl[122] vdd gnd cell_6t
Xbit_r123_c127 bl[127] br[127] wl[123] vdd gnd cell_6t
Xbit_r124_c127 bl[127] br[127] wl[124] vdd gnd cell_6t
Xbit_r125_c127 bl[127] br[127] wl[125] vdd gnd cell_6t
Xbit_r126_c127 bl[127] br[127] wl[126] vdd gnd cell_6t
Xbit_r127_c127 bl[127] br[127] wl[127] vdd gnd cell_6t
Xbit_r0_c128 bl[128] br[128] wl[0] vdd gnd cell_6t
Xbit_r1_c128 bl[128] br[128] wl[1] vdd gnd cell_6t
Xbit_r2_c128 bl[128] br[128] wl[2] vdd gnd cell_6t
Xbit_r3_c128 bl[128] br[128] wl[3] vdd gnd cell_6t
Xbit_r4_c128 bl[128] br[128] wl[4] vdd gnd cell_6t
Xbit_r5_c128 bl[128] br[128] wl[5] vdd gnd cell_6t
Xbit_r6_c128 bl[128] br[128] wl[6] vdd gnd cell_6t
Xbit_r7_c128 bl[128] br[128] wl[7] vdd gnd cell_6t
Xbit_r8_c128 bl[128] br[128] wl[8] vdd gnd cell_6t
Xbit_r9_c128 bl[128] br[128] wl[9] vdd gnd cell_6t
Xbit_r10_c128 bl[128] br[128] wl[10] vdd gnd cell_6t
Xbit_r11_c128 bl[128] br[128] wl[11] vdd gnd cell_6t
Xbit_r12_c128 bl[128] br[128] wl[12] vdd gnd cell_6t
Xbit_r13_c128 bl[128] br[128] wl[13] vdd gnd cell_6t
Xbit_r14_c128 bl[128] br[128] wl[14] vdd gnd cell_6t
Xbit_r15_c128 bl[128] br[128] wl[15] vdd gnd cell_6t
Xbit_r16_c128 bl[128] br[128] wl[16] vdd gnd cell_6t
Xbit_r17_c128 bl[128] br[128] wl[17] vdd gnd cell_6t
Xbit_r18_c128 bl[128] br[128] wl[18] vdd gnd cell_6t
Xbit_r19_c128 bl[128] br[128] wl[19] vdd gnd cell_6t
Xbit_r20_c128 bl[128] br[128] wl[20] vdd gnd cell_6t
Xbit_r21_c128 bl[128] br[128] wl[21] vdd gnd cell_6t
Xbit_r22_c128 bl[128] br[128] wl[22] vdd gnd cell_6t
Xbit_r23_c128 bl[128] br[128] wl[23] vdd gnd cell_6t
Xbit_r24_c128 bl[128] br[128] wl[24] vdd gnd cell_6t
Xbit_r25_c128 bl[128] br[128] wl[25] vdd gnd cell_6t
Xbit_r26_c128 bl[128] br[128] wl[26] vdd gnd cell_6t
Xbit_r27_c128 bl[128] br[128] wl[27] vdd gnd cell_6t
Xbit_r28_c128 bl[128] br[128] wl[28] vdd gnd cell_6t
Xbit_r29_c128 bl[128] br[128] wl[29] vdd gnd cell_6t
Xbit_r30_c128 bl[128] br[128] wl[30] vdd gnd cell_6t
Xbit_r31_c128 bl[128] br[128] wl[31] vdd gnd cell_6t
Xbit_r32_c128 bl[128] br[128] wl[32] vdd gnd cell_6t
Xbit_r33_c128 bl[128] br[128] wl[33] vdd gnd cell_6t
Xbit_r34_c128 bl[128] br[128] wl[34] vdd gnd cell_6t
Xbit_r35_c128 bl[128] br[128] wl[35] vdd gnd cell_6t
Xbit_r36_c128 bl[128] br[128] wl[36] vdd gnd cell_6t
Xbit_r37_c128 bl[128] br[128] wl[37] vdd gnd cell_6t
Xbit_r38_c128 bl[128] br[128] wl[38] vdd gnd cell_6t
Xbit_r39_c128 bl[128] br[128] wl[39] vdd gnd cell_6t
Xbit_r40_c128 bl[128] br[128] wl[40] vdd gnd cell_6t
Xbit_r41_c128 bl[128] br[128] wl[41] vdd gnd cell_6t
Xbit_r42_c128 bl[128] br[128] wl[42] vdd gnd cell_6t
Xbit_r43_c128 bl[128] br[128] wl[43] vdd gnd cell_6t
Xbit_r44_c128 bl[128] br[128] wl[44] vdd gnd cell_6t
Xbit_r45_c128 bl[128] br[128] wl[45] vdd gnd cell_6t
Xbit_r46_c128 bl[128] br[128] wl[46] vdd gnd cell_6t
Xbit_r47_c128 bl[128] br[128] wl[47] vdd gnd cell_6t
Xbit_r48_c128 bl[128] br[128] wl[48] vdd gnd cell_6t
Xbit_r49_c128 bl[128] br[128] wl[49] vdd gnd cell_6t
Xbit_r50_c128 bl[128] br[128] wl[50] vdd gnd cell_6t
Xbit_r51_c128 bl[128] br[128] wl[51] vdd gnd cell_6t
Xbit_r52_c128 bl[128] br[128] wl[52] vdd gnd cell_6t
Xbit_r53_c128 bl[128] br[128] wl[53] vdd gnd cell_6t
Xbit_r54_c128 bl[128] br[128] wl[54] vdd gnd cell_6t
Xbit_r55_c128 bl[128] br[128] wl[55] vdd gnd cell_6t
Xbit_r56_c128 bl[128] br[128] wl[56] vdd gnd cell_6t
Xbit_r57_c128 bl[128] br[128] wl[57] vdd gnd cell_6t
Xbit_r58_c128 bl[128] br[128] wl[58] vdd gnd cell_6t
Xbit_r59_c128 bl[128] br[128] wl[59] vdd gnd cell_6t
Xbit_r60_c128 bl[128] br[128] wl[60] vdd gnd cell_6t
Xbit_r61_c128 bl[128] br[128] wl[61] vdd gnd cell_6t
Xbit_r62_c128 bl[128] br[128] wl[62] vdd gnd cell_6t
Xbit_r63_c128 bl[128] br[128] wl[63] vdd gnd cell_6t
Xbit_r64_c128 bl[128] br[128] wl[64] vdd gnd cell_6t
Xbit_r65_c128 bl[128] br[128] wl[65] vdd gnd cell_6t
Xbit_r66_c128 bl[128] br[128] wl[66] vdd gnd cell_6t
Xbit_r67_c128 bl[128] br[128] wl[67] vdd gnd cell_6t
Xbit_r68_c128 bl[128] br[128] wl[68] vdd gnd cell_6t
Xbit_r69_c128 bl[128] br[128] wl[69] vdd gnd cell_6t
Xbit_r70_c128 bl[128] br[128] wl[70] vdd gnd cell_6t
Xbit_r71_c128 bl[128] br[128] wl[71] vdd gnd cell_6t
Xbit_r72_c128 bl[128] br[128] wl[72] vdd gnd cell_6t
Xbit_r73_c128 bl[128] br[128] wl[73] vdd gnd cell_6t
Xbit_r74_c128 bl[128] br[128] wl[74] vdd gnd cell_6t
Xbit_r75_c128 bl[128] br[128] wl[75] vdd gnd cell_6t
Xbit_r76_c128 bl[128] br[128] wl[76] vdd gnd cell_6t
Xbit_r77_c128 bl[128] br[128] wl[77] vdd gnd cell_6t
Xbit_r78_c128 bl[128] br[128] wl[78] vdd gnd cell_6t
Xbit_r79_c128 bl[128] br[128] wl[79] vdd gnd cell_6t
Xbit_r80_c128 bl[128] br[128] wl[80] vdd gnd cell_6t
Xbit_r81_c128 bl[128] br[128] wl[81] vdd gnd cell_6t
Xbit_r82_c128 bl[128] br[128] wl[82] vdd gnd cell_6t
Xbit_r83_c128 bl[128] br[128] wl[83] vdd gnd cell_6t
Xbit_r84_c128 bl[128] br[128] wl[84] vdd gnd cell_6t
Xbit_r85_c128 bl[128] br[128] wl[85] vdd gnd cell_6t
Xbit_r86_c128 bl[128] br[128] wl[86] vdd gnd cell_6t
Xbit_r87_c128 bl[128] br[128] wl[87] vdd gnd cell_6t
Xbit_r88_c128 bl[128] br[128] wl[88] vdd gnd cell_6t
Xbit_r89_c128 bl[128] br[128] wl[89] vdd gnd cell_6t
Xbit_r90_c128 bl[128] br[128] wl[90] vdd gnd cell_6t
Xbit_r91_c128 bl[128] br[128] wl[91] vdd gnd cell_6t
Xbit_r92_c128 bl[128] br[128] wl[92] vdd gnd cell_6t
Xbit_r93_c128 bl[128] br[128] wl[93] vdd gnd cell_6t
Xbit_r94_c128 bl[128] br[128] wl[94] vdd gnd cell_6t
Xbit_r95_c128 bl[128] br[128] wl[95] vdd gnd cell_6t
Xbit_r96_c128 bl[128] br[128] wl[96] vdd gnd cell_6t
Xbit_r97_c128 bl[128] br[128] wl[97] vdd gnd cell_6t
Xbit_r98_c128 bl[128] br[128] wl[98] vdd gnd cell_6t
Xbit_r99_c128 bl[128] br[128] wl[99] vdd gnd cell_6t
Xbit_r100_c128 bl[128] br[128] wl[100] vdd gnd cell_6t
Xbit_r101_c128 bl[128] br[128] wl[101] vdd gnd cell_6t
Xbit_r102_c128 bl[128] br[128] wl[102] vdd gnd cell_6t
Xbit_r103_c128 bl[128] br[128] wl[103] vdd gnd cell_6t
Xbit_r104_c128 bl[128] br[128] wl[104] vdd gnd cell_6t
Xbit_r105_c128 bl[128] br[128] wl[105] vdd gnd cell_6t
Xbit_r106_c128 bl[128] br[128] wl[106] vdd gnd cell_6t
Xbit_r107_c128 bl[128] br[128] wl[107] vdd gnd cell_6t
Xbit_r108_c128 bl[128] br[128] wl[108] vdd gnd cell_6t
Xbit_r109_c128 bl[128] br[128] wl[109] vdd gnd cell_6t
Xbit_r110_c128 bl[128] br[128] wl[110] vdd gnd cell_6t
Xbit_r111_c128 bl[128] br[128] wl[111] vdd gnd cell_6t
Xbit_r112_c128 bl[128] br[128] wl[112] vdd gnd cell_6t
Xbit_r113_c128 bl[128] br[128] wl[113] vdd gnd cell_6t
Xbit_r114_c128 bl[128] br[128] wl[114] vdd gnd cell_6t
Xbit_r115_c128 bl[128] br[128] wl[115] vdd gnd cell_6t
Xbit_r116_c128 bl[128] br[128] wl[116] vdd gnd cell_6t
Xbit_r117_c128 bl[128] br[128] wl[117] vdd gnd cell_6t
Xbit_r118_c128 bl[128] br[128] wl[118] vdd gnd cell_6t
Xbit_r119_c128 bl[128] br[128] wl[119] vdd gnd cell_6t
Xbit_r120_c128 bl[128] br[128] wl[120] vdd gnd cell_6t
Xbit_r121_c128 bl[128] br[128] wl[121] vdd gnd cell_6t
Xbit_r122_c128 bl[128] br[128] wl[122] vdd gnd cell_6t
Xbit_r123_c128 bl[128] br[128] wl[123] vdd gnd cell_6t
Xbit_r124_c128 bl[128] br[128] wl[124] vdd gnd cell_6t
Xbit_r125_c128 bl[128] br[128] wl[125] vdd gnd cell_6t
Xbit_r126_c128 bl[128] br[128] wl[126] vdd gnd cell_6t
Xbit_r127_c128 bl[128] br[128] wl[127] vdd gnd cell_6t
Xbit_r0_c129 bl[129] br[129] wl[0] vdd gnd cell_6t
Xbit_r1_c129 bl[129] br[129] wl[1] vdd gnd cell_6t
Xbit_r2_c129 bl[129] br[129] wl[2] vdd gnd cell_6t
Xbit_r3_c129 bl[129] br[129] wl[3] vdd gnd cell_6t
Xbit_r4_c129 bl[129] br[129] wl[4] vdd gnd cell_6t
Xbit_r5_c129 bl[129] br[129] wl[5] vdd gnd cell_6t
Xbit_r6_c129 bl[129] br[129] wl[6] vdd gnd cell_6t
Xbit_r7_c129 bl[129] br[129] wl[7] vdd gnd cell_6t
Xbit_r8_c129 bl[129] br[129] wl[8] vdd gnd cell_6t
Xbit_r9_c129 bl[129] br[129] wl[9] vdd gnd cell_6t
Xbit_r10_c129 bl[129] br[129] wl[10] vdd gnd cell_6t
Xbit_r11_c129 bl[129] br[129] wl[11] vdd gnd cell_6t
Xbit_r12_c129 bl[129] br[129] wl[12] vdd gnd cell_6t
Xbit_r13_c129 bl[129] br[129] wl[13] vdd gnd cell_6t
Xbit_r14_c129 bl[129] br[129] wl[14] vdd gnd cell_6t
Xbit_r15_c129 bl[129] br[129] wl[15] vdd gnd cell_6t
Xbit_r16_c129 bl[129] br[129] wl[16] vdd gnd cell_6t
Xbit_r17_c129 bl[129] br[129] wl[17] vdd gnd cell_6t
Xbit_r18_c129 bl[129] br[129] wl[18] vdd gnd cell_6t
Xbit_r19_c129 bl[129] br[129] wl[19] vdd gnd cell_6t
Xbit_r20_c129 bl[129] br[129] wl[20] vdd gnd cell_6t
Xbit_r21_c129 bl[129] br[129] wl[21] vdd gnd cell_6t
Xbit_r22_c129 bl[129] br[129] wl[22] vdd gnd cell_6t
Xbit_r23_c129 bl[129] br[129] wl[23] vdd gnd cell_6t
Xbit_r24_c129 bl[129] br[129] wl[24] vdd gnd cell_6t
Xbit_r25_c129 bl[129] br[129] wl[25] vdd gnd cell_6t
Xbit_r26_c129 bl[129] br[129] wl[26] vdd gnd cell_6t
Xbit_r27_c129 bl[129] br[129] wl[27] vdd gnd cell_6t
Xbit_r28_c129 bl[129] br[129] wl[28] vdd gnd cell_6t
Xbit_r29_c129 bl[129] br[129] wl[29] vdd gnd cell_6t
Xbit_r30_c129 bl[129] br[129] wl[30] vdd gnd cell_6t
Xbit_r31_c129 bl[129] br[129] wl[31] vdd gnd cell_6t
Xbit_r32_c129 bl[129] br[129] wl[32] vdd gnd cell_6t
Xbit_r33_c129 bl[129] br[129] wl[33] vdd gnd cell_6t
Xbit_r34_c129 bl[129] br[129] wl[34] vdd gnd cell_6t
Xbit_r35_c129 bl[129] br[129] wl[35] vdd gnd cell_6t
Xbit_r36_c129 bl[129] br[129] wl[36] vdd gnd cell_6t
Xbit_r37_c129 bl[129] br[129] wl[37] vdd gnd cell_6t
Xbit_r38_c129 bl[129] br[129] wl[38] vdd gnd cell_6t
Xbit_r39_c129 bl[129] br[129] wl[39] vdd gnd cell_6t
Xbit_r40_c129 bl[129] br[129] wl[40] vdd gnd cell_6t
Xbit_r41_c129 bl[129] br[129] wl[41] vdd gnd cell_6t
Xbit_r42_c129 bl[129] br[129] wl[42] vdd gnd cell_6t
Xbit_r43_c129 bl[129] br[129] wl[43] vdd gnd cell_6t
Xbit_r44_c129 bl[129] br[129] wl[44] vdd gnd cell_6t
Xbit_r45_c129 bl[129] br[129] wl[45] vdd gnd cell_6t
Xbit_r46_c129 bl[129] br[129] wl[46] vdd gnd cell_6t
Xbit_r47_c129 bl[129] br[129] wl[47] vdd gnd cell_6t
Xbit_r48_c129 bl[129] br[129] wl[48] vdd gnd cell_6t
Xbit_r49_c129 bl[129] br[129] wl[49] vdd gnd cell_6t
Xbit_r50_c129 bl[129] br[129] wl[50] vdd gnd cell_6t
Xbit_r51_c129 bl[129] br[129] wl[51] vdd gnd cell_6t
Xbit_r52_c129 bl[129] br[129] wl[52] vdd gnd cell_6t
Xbit_r53_c129 bl[129] br[129] wl[53] vdd gnd cell_6t
Xbit_r54_c129 bl[129] br[129] wl[54] vdd gnd cell_6t
Xbit_r55_c129 bl[129] br[129] wl[55] vdd gnd cell_6t
Xbit_r56_c129 bl[129] br[129] wl[56] vdd gnd cell_6t
Xbit_r57_c129 bl[129] br[129] wl[57] vdd gnd cell_6t
Xbit_r58_c129 bl[129] br[129] wl[58] vdd gnd cell_6t
Xbit_r59_c129 bl[129] br[129] wl[59] vdd gnd cell_6t
Xbit_r60_c129 bl[129] br[129] wl[60] vdd gnd cell_6t
Xbit_r61_c129 bl[129] br[129] wl[61] vdd gnd cell_6t
Xbit_r62_c129 bl[129] br[129] wl[62] vdd gnd cell_6t
Xbit_r63_c129 bl[129] br[129] wl[63] vdd gnd cell_6t
Xbit_r64_c129 bl[129] br[129] wl[64] vdd gnd cell_6t
Xbit_r65_c129 bl[129] br[129] wl[65] vdd gnd cell_6t
Xbit_r66_c129 bl[129] br[129] wl[66] vdd gnd cell_6t
Xbit_r67_c129 bl[129] br[129] wl[67] vdd gnd cell_6t
Xbit_r68_c129 bl[129] br[129] wl[68] vdd gnd cell_6t
Xbit_r69_c129 bl[129] br[129] wl[69] vdd gnd cell_6t
Xbit_r70_c129 bl[129] br[129] wl[70] vdd gnd cell_6t
Xbit_r71_c129 bl[129] br[129] wl[71] vdd gnd cell_6t
Xbit_r72_c129 bl[129] br[129] wl[72] vdd gnd cell_6t
Xbit_r73_c129 bl[129] br[129] wl[73] vdd gnd cell_6t
Xbit_r74_c129 bl[129] br[129] wl[74] vdd gnd cell_6t
Xbit_r75_c129 bl[129] br[129] wl[75] vdd gnd cell_6t
Xbit_r76_c129 bl[129] br[129] wl[76] vdd gnd cell_6t
Xbit_r77_c129 bl[129] br[129] wl[77] vdd gnd cell_6t
Xbit_r78_c129 bl[129] br[129] wl[78] vdd gnd cell_6t
Xbit_r79_c129 bl[129] br[129] wl[79] vdd gnd cell_6t
Xbit_r80_c129 bl[129] br[129] wl[80] vdd gnd cell_6t
Xbit_r81_c129 bl[129] br[129] wl[81] vdd gnd cell_6t
Xbit_r82_c129 bl[129] br[129] wl[82] vdd gnd cell_6t
Xbit_r83_c129 bl[129] br[129] wl[83] vdd gnd cell_6t
Xbit_r84_c129 bl[129] br[129] wl[84] vdd gnd cell_6t
Xbit_r85_c129 bl[129] br[129] wl[85] vdd gnd cell_6t
Xbit_r86_c129 bl[129] br[129] wl[86] vdd gnd cell_6t
Xbit_r87_c129 bl[129] br[129] wl[87] vdd gnd cell_6t
Xbit_r88_c129 bl[129] br[129] wl[88] vdd gnd cell_6t
Xbit_r89_c129 bl[129] br[129] wl[89] vdd gnd cell_6t
Xbit_r90_c129 bl[129] br[129] wl[90] vdd gnd cell_6t
Xbit_r91_c129 bl[129] br[129] wl[91] vdd gnd cell_6t
Xbit_r92_c129 bl[129] br[129] wl[92] vdd gnd cell_6t
Xbit_r93_c129 bl[129] br[129] wl[93] vdd gnd cell_6t
Xbit_r94_c129 bl[129] br[129] wl[94] vdd gnd cell_6t
Xbit_r95_c129 bl[129] br[129] wl[95] vdd gnd cell_6t
Xbit_r96_c129 bl[129] br[129] wl[96] vdd gnd cell_6t
Xbit_r97_c129 bl[129] br[129] wl[97] vdd gnd cell_6t
Xbit_r98_c129 bl[129] br[129] wl[98] vdd gnd cell_6t
Xbit_r99_c129 bl[129] br[129] wl[99] vdd gnd cell_6t
Xbit_r100_c129 bl[129] br[129] wl[100] vdd gnd cell_6t
Xbit_r101_c129 bl[129] br[129] wl[101] vdd gnd cell_6t
Xbit_r102_c129 bl[129] br[129] wl[102] vdd gnd cell_6t
Xbit_r103_c129 bl[129] br[129] wl[103] vdd gnd cell_6t
Xbit_r104_c129 bl[129] br[129] wl[104] vdd gnd cell_6t
Xbit_r105_c129 bl[129] br[129] wl[105] vdd gnd cell_6t
Xbit_r106_c129 bl[129] br[129] wl[106] vdd gnd cell_6t
Xbit_r107_c129 bl[129] br[129] wl[107] vdd gnd cell_6t
Xbit_r108_c129 bl[129] br[129] wl[108] vdd gnd cell_6t
Xbit_r109_c129 bl[129] br[129] wl[109] vdd gnd cell_6t
Xbit_r110_c129 bl[129] br[129] wl[110] vdd gnd cell_6t
Xbit_r111_c129 bl[129] br[129] wl[111] vdd gnd cell_6t
Xbit_r112_c129 bl[129] br[129] wl[112] vdd gnd cell_6t
Xbit_r113_c129 bl[129] br[129] wl[113] vdd gnd cell_6t
Xbit_r114_c129 bl[129] br[129] wl[114] vdd gnd cell_6t
Xbit_r115_c129 bl[129] br[129] wl[115] vdd gnd cell_6t
Xbit_r116_c129 bl[129] br[129] wl[116] vdd gnd cell_6t
Xbit_r117_c129 bl[129] br[129] wl[117] vdd gnd cell_6t
Xbit_r118_c129 bl[129] br[129] wl[118] vdd gnd cell_6t
Xbit_r119_c129 bl[129] br[129] wl[119] vdd gnd cell_6t
Xbit_r120_c129 bl[129] br[129] wl[120] vdd gnd cell_6t
Xbit_r121_c129 bl[129] br[129] wl[121] vdd gnd cell_6t
Xbit_r122_c129 bl[129] br[129] wl[122] vdd gnd cell_6t
Xbit_r123_c129 bl[129] br[129] wl[123] vdd gnd cell_6t
Xbit_r124_c129 bl[129] br[129] wl[124] vdd gnd cell_6t
Xbit_r125_c129 bl[129] br[129] wl[125] vdd gnd cell_6t
Xbit_r126_c129 bl[129] br[129] wl[126] vdd gnd cell_6t
Xbit_r127_c129 bl[129] br[129] wl[127] vdd gnd cell_6t
Xbit_r0_c130 bl[130] br[130] wl[0] vdd gnd cell_6t
Xbit_r1_c130 bl[130] br[130] wl[1] vdd gnd cell_6t
Xbit_r2_c130 bl[130] br[130] wl[2] vdd gnd cell_6t
Xbit_r3_c130 bl[130] br[130] wl[3] vdd gnd cell_6t
Xbit_r4_c130 bl[130] br[130] wl[4] vdd gnd cell_6t
Xbit_r5_c130 bl[130] br[130] wl[5] vdd gnd cell_6t
Xbit_r6_c130 bl[130] br[130] wl[6] vdd gnd cell_6t
Xbit_r7_c130 bl[130] br[130] wl[7] vdd gnd cell_6t
Xbit_r8_c130 bl[130] br[130] wl[8] vdd gnd cell_6t
Xbit_r9_c130 bl[130] br[130] wl[9] vdd gnd cell_6t
Xbit_r10_c130 bl[130] br[130] wl[10] vdd gnd cell_6t
Xbit_r11_c130 bl[130] br[130] wl[11] vdd gnd cell_6t
Xbit_r12_c130 bl[130] br[130] wl[12] vdd gnd cell_6t
Xbit_r13_c130 bl[130] br[130] wl[13] vdd gnd cell_6t
Xbit_r14_c130 bl[130] br[130] wl[14] vdd gnd cell_6t
Xbit_r15_c130 bl[130] br[130] wl[15] vdd gnd cell_6t
Xbit_r16_c130 bl[130] br[130] wl[16] vdd gnd cell_6t
Xbit_r17_c130 bl[130] br[130] wl[17] vdd gnd cell_6t
Xbit_r18_c130 bl[130] br[130] wl[18] vdd gnd cell_6t
Xbit_r19_c130 bl[130] br[130] wl[19] vdd gnd cell_6t
Xbit_r20_c130 bl[130] br[130] wl[20] vdd gnd cell_6t
Xbit_r21_c130 bl[130] br[130] wl[21] vdd gnd cell_6t
Xbit_r22_c130 bl[130] br[130] wl[22] vdd gnd cell_6t
Xbit_r23_c130 bl[130] br[130] wl[23] vdd gnd cell_6t
Xbit_r24_c130 bl[130] br[130] wl[24] vdd gnd cell_6t
Xbit_r25_c130 bl[130] br[130] wl[25] vdd gnd cell_6t
Xbit_r26_c130 bl[130] br[130] wl[26] vdd gnd cell_6t
Xbit_r27_c130 bl[130] br[130] wl[27] vdd gnd cell_6t
Xbit_r28_c130 bl[130] br[130] wl[28] vdd gnd cell_6t
Xbit_r29_c130 bl[130] br[130] wl[29] vdd gnd cell_6t
Xbit_r30_c130 bl[130] br[130] wl[30] vdd gnd cell_6t
Xbit_r31_c130 bl[130] br[130] wl[31] vdd gnd cell_6t
Xbit_r32_c130 bl[130] br[130] wl[32] vdd gnd cell_6t
Xbit_r33_c130 bl[130] br[130] wl[33] vdd gnd cell_6t
Xbit_r34_c130 bl[130] br[130] wl[34] vdd gnd cell_6t
Xbit_r35_c130 bl[130] br[130] wl[35] vdd gnd cell_6t
Xbit_r36_c130 bl[130] br[130] wl[36] vdd gnd cell_6t
Xbit_r37_c130 bl[130] br[130] wl[37] vdd gnd cell_6t
Xbit_r38_c130 bl[130] br[130] wl[38] vdd gnd cell_6t
Xbit_r39_c130 bl[130] br[130] wl[39] vdd gnd cell_6t
Xbit_r40_c130 bl[130] br[130] wl[40] vdd gnd cell_6t
Xbit_r41_c130 bl[130] br[130] wl[41] vdd gnd cell_6t
Xbit_r42_c130 bl[130] br[130] wl[42] vdd gnd cell_6t
Xbit_r43_c130 bl[130] br[130] wl[43] vdd gnd cell_6t
Xbit_r44_c130 bl[130] br[130] wl[44] vdd gnd cell_6t
Xbit_r45_c130 bl[130] br[130] wl[45] vdd gnd cell_6t
Xbit_r46_c130 bl[130] br[130] wl[46] vdd gnd cell_6t
Xbit_r47_c130 bl[130] br[130] wl[47] vdd gnd cell_6t
Xbit_r48_c130 bl[130] br[130] wl[48] vdd gnd cell_6t
Xbit_r49_c130 bl[130] br[130] wl[49] vdd gnd cell_6t
Xbit_r50_c130 bl[130] br[130] wl[50] vdd gnd cell_6t
Xbit_r51_c130 bl[130] br[130] wl[51] vdd gnd cell_6t
Xbit_r52_c130 bl[130] br[130] wl[52] vdd gnd cell_6t
Xbit_r53_c130 bl[130] br[130] wl[53] vdd gnd cell_6t
Xbit_r54_c130 bl[130] br[130] wl[54] vdd gnd cell_6t
Xbit_r55_c130 bl[130] br[130] wl[55] vdd gnd cell_6t
Xbit_r56_c130 bl[130] br[130] wl[56] vdd gnd cell_6t
Xbit_r57_c130 bl[130] br[130] wl[57] vdd gnd cell_6t
Xbit_r58_c130 bl[130] br[130] wl[58] vdd gnd cell_6t
Xbit_r59_c130 bl[130] br[130] wl[59] vdd gnd cell_6t
Xbit_r60_c130 bl[130] br[130] wl[60] vdd gnd cell_6t
Xbit_r61_c130 bl[130] br[130] wl[61] vdd gnd cell_6t
Xbit_r62_c130 bl[130] br[130] wl[62] vdd gnd cell_6t
Xbit_r63_c130 bl[130] br[130] wl[63] vdd gnd cell_6t
Xbit_r64_c130 bl[130] br[130] wl[64] vdd gnd cell_6t
Xbit_r65_c130 bl[130] br[130] wl[65] vdd gnd cell_6t
Xbit_r66_c130 bl[130] br[130] wl[66] vdd gnd cell_6t
Xbit_r67_c130 bl[130] br[130] wl[67] vdd gnd cell_6t
Xbit_r68_c130 bl[130] br[130] wl[68] vdd gnd cell_6t
Xbit_r69_c130 bl[130] br[130] wl[69] vdd gnd cell_6t
Xbit_r70_c130 bl[130] br[130] wl[70] vdd gnd cell_6t
Xbit_r71_c130 bl[130] br[130] wl[71] vdd gnd cell_6t
Xbit_r72_c130 bl[130] br[130] wl[72] vdd gnd cell_6t
Xbit_r73_c130 bl[130] br[130] wl[73] vdd gnd cell_6t
Xbit_r74_c130 bl[130] br[130] wl[74] vdd gnd cell_6t
Xbit_r75_c130 bl[130] br[130] wl[75] vdd gnd cell_6t
Xbit_r76_c130 bl[130] br[130] wl[76] vdd gnd cell_6t
Xbit_r77_c130 bl[130] br[130] wl[77] vdd gnd cell_6t
Xbit_r78_c130 bl[130] br[130] wl[78] vdd gnd cell_6t
Xbit_r79_c130 bl[130] br[130] wl[79] vdd gnd cell_6t
Xbit_r80_c130 bl[130] br[130] wl[80] vdd gnd cell_6t
Xbit_r81_c130 bl[130] br[130] wl[81] vdd gnd cell_6t
Xbit_r82_c130 bl[130] br[130] wl[82] vdd gnd cell_6t
Xbit_r83_c130 bl[130] br[130] wl[83] vdd gnd cell_6t
Xbit_r84_c130 bl[130] br[130] wl[84] vdd gnd cell_6t
Xbit_r85_c130 bl[130] br[130] wl[85] vdd gnd cell_6t
Xbit_r86_c130 bl[130] br[130] wl[86] vdd gnd cell_6t
Xbit_r87_c130 bl[130] br[130] wl[87] vdd gnd cell_6t
Xbit_r88_c130 bl[130] br[130] wl[88] vdd gnd cell_6t
Xbit_r89_c130 bl[130] br[130] wl[89] vdd gnd cell_6t
Xbit_r90_c130 bl[130] br[130] wl[90] vdd gnd cell_6t
Xbit_r91_c130 bl[130] br[130] wl[91] vdd gnd cell_6t
Xbit_r92_c130 bl[130] br[130] wl[92] vdd gnd cell_6t
Xbit_r93_c130 bl[130] br[130] wl[93] vdd gnd cell_6t
Xbit_r94_c130 bl[130] br[130] wl[94] vdd gnd cell_6t
Xbit_r95_c130 bl[130] br[130] wl[95] vdd gnd cell_6t
Xbit_r96_c130 bl[130] br[130] wl[96] vdd gnd cell_6t
Xbit_r97_c130 bl[130] br[130] wl[97] vdd gnd cell_6t
Xbit_r98_c130 bl[130] br[130] wl[98] vdd gnd cell_6t
Xbit_r99_c130 bl[130] br[130] wl[99] vdd gnd cell_6t
Xbit_r100_c130 bl[130] br[130] wl[100] vdd gnd cell_6t
Xbit_r101_c130 bl[130] br[130] wl[101] vdd gnd cell_6t
Xbit_r102_c130 bl[130] br[130] wl[102] vdd gnd cell_6t
Xbit_r103_c130 bl[130] br[130] wl[103] vdd gnd cell_6t
Xbit_r104_c130 bl[130] br[130] wl[104] vdd gnd cell_6t
Xbit_r105_c130 bl[130] br[130] wl[105] vdd gnd cell_6t
Xbit_r106_c130 bl[130] br[130] wl[106] vdd gnd cell_6t
Xbit_r107_c130 bl[130] br[130] wl[107] vdd gnd cell_6t
Xbit_r108_c130 bl[130] br[130] wl[108] vdd gnd cell_6t
Xbit_r109_c130 bl[130] br[130] wl[109] vdd gnd cell_6t
Xbit_r110_c130 bl[130] br[130] wl[110] vdd gnd cell_6t
Xbit_r111_c130 bl[130] br[130] wl[111] vdd gnd cell_6t
Xbit_r112_c130 bl[130] br[130] wl[112] vdd gnd cell_6t
Xbit_r113_c130 bl[130] br[130] wl[113] vdd gnd cell_6t
Xbit_r114_c130 bl[130] br[130] wl[114] vdd gnd cell_6t
Xbit_r115_c130 bl[130] br[130] wl[115] vdd gnd cell_6t
Xbit_r116_c130 bl[130] br[130] wl[116] vdd gnd cell_6t
Xbit_r117_c130 bl[130] br[130] wl[117] vdd gnd cell_6t
Xbit_r118_c130 bl[130] br[130] wl[118] vdd gnd cell_6t
Xbit_r119_c130 bl[130] br[130] wl[119] vdd gnd cell_6t
Xbit_r120_c130 bl[130] br[130] wl[120] vdd gnd cell_6t
Xbit_r121_c130 bl[130] br[130] wl[121] vdd gnd cell_6t
Xbit_r122_c130 bl[130] br[130] wl[122] vdd gnd cell_6t
Xbit_r123_c130 bl[130] br[130] wl[123] vdd gnd cell_6t
Xbit_r124_c130 bl[130] br[130] wl[124] vdd gnd cell_6t
Xbit_r125_c130 bl[130] br[130] wl[125] vdd gnd cell_6t
Xbit_r126_c130 bl[130] br[130] wl[126] vdd gnd cell_6t
Xbit_r127_c130 bl[130] br[130] wl[127] vdd gnd cell_6t
Xbit_r0_c131 bl[131] br[131] wl[0] vdd gnd cell_6t
Xbit_r1_c131 bl[131] br[131] wl[1] vdd gnd cell_6t
Xbit_r2_c131 bl[131] br[131] wl[2] vdd gnd cell_6t
Xbit_r3_c131 bl[131] br[131] wl[3] vdd gnd cell_6t
Xbit_r4_c131 bl[131] br[131] wl[4] vdd gnd cell_6t
Xbit_r5_c131 bl[131] br[131] wl[5] vdd gnd cell_6t
Xbit_r6_c131 bl[131] br[131] wl[6] vdd gnd cell_6t
Xbit_r7_c131 bl[131] br[131] wl[7] vdd gnd cell_6t
Xbit_r8_c131 bl[131] br[131] wl[8] vdd gnd cell_6t
Xbit_r9_c131 bl[131] br[131] wl[9] vdd gnd cell_6t
Xbit_r10_c131 bl[131] br[131] wl[10] vdd gnd cell_6t
Xbit_r11_c131 bl[131] br[131] wl[11] vdd gnd cell_6t
Xbit_r12_c131 bl[131] br[131] wl[12] vdd gnd cell_6t
Xbit_r13_c131 bl[131] br[131] wl[13] vdd gnd cell_6t
Xbit_r14_c131 bl[131] br[131] wl[14] vdd gnd cell_6t
Xbit_r15_c131 bl[131] br[131] wl[15] vdd gnd cell_6t
Xbit_r16_c131 bl[131] br[131] wl[16] vdd gnd cell_6t
Xbit_r17_c131 bl[131] br[131] wl[17] vdd gnd cell_6t
Xbit_r18_c131 bl[131] br[131] wl[18] vdd gnd cell_6t
Xbit_r19_c131 bl[131] br[131] wl[19] vdd gnd cell_6t
Xbit_r20_c131 bl[131] br[131] wl[20] vdd gnd cell_6t
Xbit_r21_c131 bl[131] br[131] wl[21] vdd gnd cell_6t
Xbit_r22_c131 bl[131] br[131] wl[22] vdd gnd cell_6t
Xbit_r23_c131 bl[131] br[131] wl[23] vdd gnd cell_6t
Xbit_r24_c131 bl[131] br[131] wl[24] vdd gnd cell_6t
Xbit_r25_c131 bl[131] br[131] wl[25] vdd gnd cell_6t
Xbit_r26_c131 bl[131] br[131] wl[26] vdd gnd cell_6t
Xbit_r27_c131 bl[131] br[131] wl[27] vdd gnd cell_6t
Xbit_r28_c131 bl[131] br[131] wl[28] vdd gnd cell_6t
Xbit_r29_c131 bl[131] br[131] wl[29] vdd gnd cell_6t
Xbit_r30_c131 bl[131] br[131] wl[30] vdd gnd cell_6t
Xbit_r31_c131 bl[131] br[131] wl[31] vdd gnd cell_6t
Xbit_r32_c131 bl[131] br[131] wl[32] vdd gnd cell_6t
Xbit_r33_c131 bl[131] br[131] wl[33] vdd gnd cell_6t
Xbit_r34_c131 bl[131] br[131] wl[34] vdd gnd cell_6t
Xbit_r35_c131 bl[131] br[131] wl[35] vdd gnd cell_6t
Xbit_r36_c131 bl[131] br[131] wl[36] vdd gnd cell_6t
Xbit_r37_c131 bl[131] br[131] wl[37] vdd gnd cell_6t
Xbit_r38_c131 bl[131] br[131] wl[38] vdd gnd cell_6t
Xbit_r39_c131 bl[131] br[131] wl[39] vdd gnd cell_6t
Xbit_r40_c131 bl[131] br[131] wl[40] vdd gnd cell_6t
Xbit_r41_c131 bl[131] br[131] wl[41] vdd gnd cell_6t
Xbit_r42_c131 bl[131] br[131] wl[42] vdd gnd cell_6t
Xbit_r43_c131 bl[131] br[131] wl[43] vdd gnd cell_6t
Xbit_r44_c131 bl[131] br[131] wl[44] vdd gnd cell_6t
Xbit_r45_c131 bl[131] br[131] wl[45] vdd gnd cell_6t
Xbit_r46_c131 bl[131] br[131] wl[46] vdd gnd cell_6t
Xbit_r47_c131 bl[131] br[131] wl[47] vdd gnd cell_6t
Xbit_r48_c131 bl[131] br[131] wl[48] vdd gnd cell_6t
Xbit_r49_c131 bl[131] br[131] wl[49] vdd gnd cell_6t
Xbit_r50_c131 bl[131] br[131] wl[50] vdd gnd cell_6t
Xbit_r51_c131 bl[131] br[131] wl[51] vdd gnd cell_6t
Xbit_r52_c131 bl[131] br[131] wl[52] vdd gnd cell_6t
Xbit_r53_c131 bl[131] br[131] wl[53] vdd gnd cell_6t
Xbit_r54_c131 bl[131] br[131] wl[54] vdd gnd cell_6t
Xbit_r55_c131 bl[131] br[131] wl[55] vdd gnd cell_6t
Xbit_r56_c131 bl[131] br[131] wl[56] vdd gnd cell_6t
Xbit_r57_c131 bl[131] br[131] wl[57] vdd gnd cell_6t
Xbit_r58_c131 bl[131] br[131] wl[58] vdd gnd cell_6t
Xbit_r59_c131 bl[131] br[131] wl[59] vdd gnd cell_6t
Xbit_r60_c131 bl[131] br[131] wl[60] vdd gnd cell_6t
Xbit_r61_c131 bl[131] br[131] wl[61] vdd gnd cell_6t
Xbit_r62_c131 bl[131] br[131] wl[62] vdd gnd cell_6t
Xbit_r63_c131 bl[131] br[131] wl[63] vdd gnd cell_6t
Xbit_r64_c131 bl[131] br[131] wl[64] vdd gnd cell_6t
Xbit_r65_c131 bl[131] br[131] wl[65] vdd gnd cell_6t
Xbit_r66_c131 bl[131] br[131] wl[66] vdd gnd cell_6t
Xbit_r67_c131 bl[131] br[131] wl[67] vdd gnd cell_6t
Xbit_r68_c131 bl[131] br[131] wl[68] vdd gnd cell_6t
Xbit_r69_c131 bl[131] br[131] wl[69] vdd gnd cell_6t
Xbit_r70_c131 bl[131] br[131] wl[70] vdd gnd cell_6t
Xbit_r71_c131 bl[131] br[131] wl[71] vdd gnd cell_6t
Xbit_r72_c131 bl[131] br[131] wl[72] vdd gnd cell_6t
Xbit_r73_c131 bl[131] br[131] wl[73] vdd gnd cell_6t
Xbit_r74_c131 bl[131] br[131] wl[74] vdd gnd cell_6t
Xbit_r75_c131 bl[131] br[131] wl[75] vdd gnd cell_6t
Xbit_r76_c131 bl[131] br[131] wl[76] vdd gnd cell_6t
Xbit_r77_c131 bl[131] br[131] wl[77] vdd gnd cell_6t
Xbit_r78_c131 bl[131] br[131] wl[78] vdd gnd cell_6t
Xbit_r79_c131 bl[131] br[131] wl[79] vdd gnd cell_6t
Xbit_r80_c131 bl[131] br[131] wl[80] vdd gnd cell_6t
Xbit_r81_c131 bl[131] br[131] wl[81] vdd gnd cell_6t
Xbit_r82_c131 bl[131] br[131] wl[82] vdd gnd cell_6t
Xbit_r83_c131 bl[131] br[131] wl[83] vdd gnd cell_6t
Xbit_r84_c131 bl[131] br[131] wl[84] vdd gnd cell_6t
Xbit_r85_c131 bl[131] br[131] wl[85] vdd gnd cell_6t
Xbit_r86_c131 bl[131] br[131] wl[86] vdd gnd cell_6t
Xbit_r87_c131 bl[131] br[131] wl[87] vdd gnd cell_6t
Xbit_r88_c131 bl[131] br[131] wl[88] vdd gnd cell_6t
Xbit_r89_c131 bl[131] br[131] wl[89] vdd gnd cell_6t
Xbit_r90_c131 bl[131] br[131] wl[90] vdd gnd cell_6t
Xbit_r91_c131 bl[131] br[131] wl[91] vdd gnd cell_6t
Xbit_r92_c131 bl[131] br[131] wl[92] vdd gnd cell_6t
Xbit_r93_c131 bl[131] br[131] wl[93] vdd gnd cell_6t
Xbit_r94_c131 bl[131] br[131] wl[94] vdd gnd cell_6t
Xbit_r95_c131 bl[131] br[131] wl[95] vdd gnd cell_6t
Xbit_r96_c131 bl[131] br[131] wl[96] vdd gnd cell_6t
Xbit_r97_c131 bl[131] br[131] wl[97] vdd gnd cell_6t
Xbit_r98_c131 bl[131] br[131] wl[98] vdd gnd cell_6t
Xbit_r99_c131 bl[131] br[131] wl[99] vdd gnd cell_6t
Xbit_r100_c131 bl[131] br[131] wl[100] vdd gnd cell_6t
Xbit_r101_c131 bl[131] br[131] wl[101] vdd gnd cell_6t
Xbit_r102_c131 bl[131] br[131] wl[102] vdd gnd cell_6t
Xbit_r103_c131 bl[131] br[131] wl[103] vdd gnd cell_6t
Xbit_r104_c131 bl[131] br[131] wl[104] vdd gnd cell_6t
Xbit_r105_c131 bl[131] br[131] wl[105] vdd gnd cell_6t
Xbit_r106_c131 bl[131] br[131] wl[106] vdd gnd cell_6t
Xbit_r107_c131 bl[131] br[131] wl[107] vdd gnd cell_6t
Xbit_r108_c131 bl[131] br[131] wl[108] vdd gnd cell_6t
Xbit_r109_c131 bl[131] br[131] wl[109] vdd gnd cell_6t
Xbit_r110_c131 bl[131] br[131] wl[110] vdd gnd cell_6t
Xbit_r111_c131 bl[131] br[131] wl[111] vdd gnd cell_6t
Xbit_r112_c131 bl[131] br[131] wl[112] vdd gnd cell_6t
Xbit_r113_c131 bl[131] br[131] wl[113] vdd gnd cell_6t
Xbit_r114_c131 bl[131] br[131] wl[114] vdd gnd cell_6t
Xbit_r115_c131 bl[131] br[131] wl[115] vdd gnd cell_6t
Xbit_r116_c131 bl[131] br[131] wl[116] vdd gnd cell_6t
Xbit_r117_c131 bl[131] br[131] wl[117] vdd gnd cell_6t
Xbit_r118_c131 bl[131] br[131] wl[118] vdd gnd cell_6t
Xbit_r119_c131 bl[131] br[131] wl[119] vdd gnd cell_6t
Xbit_r120_c131 bl[131] br[131] wl[120] vdd gnd cell_6t
Xbit_r121_c131 bl[131] br[131] wl[121] vdd gnd cell_6t
Xbit_r122_c131 bl[131] br[131] wl[122] vdd gnd cell_6t
Xbit_r123_c131 bl[131] br[131] wl[123] vdd gnd cell_6t
Xbit_r124_c131 bl[131] br[131] wl[124] vdd gnd cell_6t
Xbit_r125_c131 bl[131] br[131] wl[125] vdd gnd cell_6t
Xbit_r126_c131 bl[131] br[131] wl[126] vdd gnd cell_6t
Xbit_r127_c131 bl[131] br[131] wl[127] vdd gnd cell_6t
Xbit_r0_c132 bl[132] br[132] wl[0] vdd gnd cell_6t
Xbit_r1_c132 bl[132] br[132] wl[1] vdd gnd cell_6t
Xbit_r2_c132 bl[132] br[132] wl[2] vdd gnd cell_6t
Xbit_r3_c132 bl[132] br[132] wl[3] vdd gnd cell_6t
Xbit_r4_c132 bl[132] br[132] wl[4] vdd gnd cell_6t
Xbit_r5_c132 bl[132] br[132] wl[5] vdd gnd cell_6t
Xbit_r6_c132 bl[132] br[132] wl[6] vdd gnd cell_6t
Xbit_r7_c132 bl[132] br[132] wl[7] vdd gnd cell_6t
Xbit_r8_c132 bl[132] br[132] wl[8] vdd gnd cell_6t
Xbit_r9_c132 bl[132] br[132] wl[9] vdd gnd cell_6t
Xbit_r10_c132 bl[132] br[132] wl[10] vdd gnd cell_6t
Xbit_r11_c132 bl[132] br[132] wl[11] vdd gnd cell_6t
Xbit_r12_c132 bl[132] br[132] wl[12] vdd gnd cell_6t
Xbit_r13_c132 bl[132] br[132] wl[13] vdd gnd cell_6t
Xbit_r14_c132 bl[132] br[132] wl[14] vdd gnd cell_6t
Xbit_r15_c132 bl[132] br[132] wl[15] vdd gnd cell_6t
Xbit_r16_c132 bl[132] br[132] wl[16] vdd gnd cell_6t
Xbit_r17_c132 bl[132] br[132] wl[17] vdd gnd cell_6t
Xbit_r18_c132 bl[132] br[132] wl[18] vdd gnd cell_6t
Xbit_r19_c132 bl[132] br[132] wl[19] vdd gnd cell_6t
Xbit_r20_c132 bl[132] br[132] wl[20] vdd gnd cell_6t
Xbit_r21_c132 bl[132] br[132] wl[21] vdd gnd cell_6t
Xbit_r22_c132 bl[132] br[132] wl[22] vdd gnd cell_6t
Xbit_r23_c132 bl[132] br[132] wl[23] vdd gnd cell_6t
Xbit_r24_c132 bl[132] br[132] wl[24] vdd gnd cell_6t
Xbit_r25_c132 bl[132] br[132] wl[25] vdd gnd cell_6t
Xbit_r26_c132 bl[132] br[132] wl[26] vdd gnd cell_6t
Xbit_r27_c132 bl[132] br[132] wl[27] vdd gnd cell_6t
Xbit_r28_c132 bl[132] br[132] wl[28] vdd gnd cell_6t
Xbit_r29_c132 bl[132] br[132] wl[29] vdd gnd cell_6t
Xbit_r30_c132 bl[132] br[132] wl[30] vdd gnd cell_6t
Xbit_r31_c132 bl[132] br[132] wl[31] vdd gnd cell_6t
Xbit_r32_c132 bl[132] br[132] wl[32] vdd gnd cell_6t
Xbit_r33_c132 bl[132] br[132] wl[33] vdd gnd cell_6t
Xbit_r34_c132 bl[132] br[132] wl[34] vdd gnd cell_6t
Xbit_r35_c132 bl[132] br[132] wl[35] vdd gnd cell_6t
Xbit_r36_c132 bl[132] br[132] wl[36] vdd gnd cell_6t
Xbit_r37_c132 bl[132] br[132] wl[37] vdd gnd cell_6t
Xbit_r38_c132 bl[132] br[132] wl[38] vdd gnd cell_6t
Xbit_r39_c132 bl[132] br[132] wl[39] vdd gnd cell_6t
Xbit_r40_c132 bl[132] br[132] wl[40] vdd gnd cell_6t
Xbit_r41_c132 bl[132] br[132] wl[41] vdd gnd cell_6t
Xbit_r42_c132 bl[132] br[132] wl[42] vdd gnd cell_6t
Xbit_r43_c132 bl[132] br[132] wl[43] vdd gnd cell_6t
Xbit_r44_c132 bl[132] br[132] wl[44] vdd gnd cell_6t
Xbit_r45_c132 bl[132] br[132] wl[45] vdd gnd cell_6t
Xbit_r46_c132 bl[132] br[132] wl[46] vdd gnd cell_6t
Xbit_r47_c132 bl[132] br[132] wl[47] vdd gnd cell_6t
Xbit_r48_c132 bl[132] br[132] wl[48] vdd gnd cell_6t
Xbit_r49_c132 bl[132] br[132] wl[49] vdd gnd cell_6t
Xbit_r50_c132 bl[132] br[132] wl[50] vdd gnd cell_6t
Xbit_r51_c132 bl[132] br[132] wl[51] vdd gnd cell_6t
Xbit_r52_c132 bl[132] br[132] wl[52] vdd gnd cell_6t
Xbit_r53_c132 bl[132] br[132] wl[53] vdd gnd cell_6t
Xbit_r54_c132 bl[132] br[132] wl[54] vdd gnd cell_6t
Xbit_r55_c132 bl[132] br[132] wl[55] vdd gnd cell_6t
Xbit_r56_c132 bl[132] br[132] wl[56] vdd gnd cell_6t
Xbit_r57_c132 bl[132] br[132] wl[57] vdd gnd cell_6t
Xbit_r58_c132 bl[132] br[132] wl[58] vdd gnd cell_6t
Xbit_r59_c132 bl[132] br[132] wl[59] vdd gnd cell_6t
Xbit_r60_c132 bl[132] br[132] wl[60] vdd gnd cell_6t
Xbit_r61_c132 bl[132] br[132] wl[61] vdd gnd cell_6t
Xbit_r62_c132 bl[132] br[132] wl[62] vdd gnd cell_6t
Xbit_r63_c132 bl[132] br[132] wl[63] vdd gnd cell_6t
Xbit_r64_c132 bl[132] br[132] wl[64] vdd gnd cell_6t
Xbit_r65_c132 bl[132] br[132] wl[65] vdd gnd cell_6t
Xbit_r66_c132 bl[132] br[132] wl[66] vdd gnd cell_6t
Xbit_r67_c132 bl[132] br[132] wl[67] vdd gnd cell_6t
Xbit_r68_c132 bl[132] br[132] wl[68] vdd gnd cell_6t
Xbit_r69_c132 bl[132] br[132] wl[69] vdd gnd cell_6t
Xbit_r70_c132 bl[132] br[132] wl[70] vdd gnd cell_6t
Xbit_r71_c132 bl[132] br[132] wl[71] vdd gnd cell_6t
Xbit_r72_c132 bl[132] br[132] wl[72] vdd gnd cell_6t
Xbit_r73_c132 bl[132] br[132] wl[73] vdd gnd cell_6t
Xbit_r74_c132 bl[132] br[132] wl[74] vdd gnd cell_6t
Xbit_r75_c132 bl[132] br[132] wl[75] vdd gnd cell_6t
Xbit_r76_c132 bl[132] br[132] wl[76] vdd gnd cell_6t
Xbit_r77_c132 bl[132] br[132] wl[77] vdd gnd cell_6t
Xbit_r78_c132 bl[132] br[132] wl[78] vdd gnd cell_6t
Xbit_r79_c132 bl[132] br[132] wl[79] vdd gnd cell_6t
Xbit_r80_c132 bl[132] br[132] wl[80] vdd gnd cell_6t
Xbit_r81_c132 bl[132] br[132] wl[81] vdd gnd cell_6t
Xbit_r82_c132 bl[132] br[132] wl[82] vdd gnd cell_6t
Xbit_r83_c132 bl[132] br[132] wl[83] vdd gnd cell_6t
Xbit_r84_c132 bl[132] br[132] wl[84] vdd gnd cell_6t
Xbit_r85_c132 bl[132] br[132] wl[85] vdd gnd cell_6t
Xbit_r86_c132 bl[132] br[132] wl[86] vdd gnd cell_6t
Xbit_r87_c132 bl[132] br[132] wl[87] vdd gnd cell_6t
Xbit_r88_c132 bl[132] br[132] wl[88] vdd gnd cell_6t
Xbit_r89_c132 bl[132] br[132] wl[89] vdd gnd cell_6t
Xbit_r90_c132 bl[132] br[132] wl[90] vdd gnd cell_6t
Xbit_r91_c132 bl[132] br[132] wl[91] vdd gnd cell_6t
Xbit_r92_c132 bl[132] br[132] wl[92] vdd gnd cell_6t
Xbit_r93_c132 bl[132] br[132] wl[93] vdd gnd cell_6t
Xbit_r94_c132 bl[132] br[132] wl[94] vdd gnd cell_6t
Xbit_r95_c132 bl[132] br[132] wl[95] vdd gnd cell_6t
Xbit_r96_c132 bl[132] br[132] wl[96] vdd gnd cell_6t
Xbit_r97_c132 bl[132] br[132] wl[97] vdd gnd cell_6t
Xbit_r98_c132 bl[132] br[132] wl[98] vdd gnd cell_6t
Xbit_r99_c132 bl[132] br[132] wl[99] vdd gnd cell_6t
Xbit_r100_c132 bl[132] br[132] wl[100] vdd gnd cell_6t
Xbit_r101_c132 bl[132] br[132] wl[101] vdd gnd cell_6t
Xbit_r102_c132 bl[132] br[132] wl[102] vdd gnd cell_6t
Xbit_r103_c132 bl[132] br[132] wl[103] vdd gnd cell_6t
Xbit_r104_c132 bl[132] br[132] wl[104] vdd gnd cell_6t
Xbit_r105_c132 bl[132] br[132] wl[105] vdd gnd cell_6t
Xbit_r106_c132 bl[132] br[132] wl[106] vdd gnd cell_6t
Xbit_r107_c132 bl[132] br[132] wl[107] vdd gnd cell_6t
Xbit_r108_c132 bl[132] br[132] wl[108] vdd gnd cell_6t
Xbit_r109_c132 bl[132] br[132] wl[109] vdd gnd cell_6t
Xbit_r110_c132 bl[132] br[132] wl[110] vdd gnd cell_6t
Xbit_r111_c132 bl[132] br[132] wl[111] vdd gnd cell_6t
Xbit_r112_c132 bl[132] br[132] wl[112] vdd gnd cell_6t
Xbit_r113_c132 bl[132] br[132] wl[113] vdd gnd cell_6t
Xbit_r114_c132 bl[132] br[132] wl[114] vdd gnd cell_6t
Xbit_r115_c132 bl[132] br[132] wl[115] vdd gnd cell_6t
Xbit_r116_c132 bl[132] br[132] wl[116] vdd gnd cell_6t
Xbit_r117_c132 bl[132] br[132] wl[117] vdd gnd cell_6t
Xbit_r118_c132 bl[132] br[132] wl[118] vdd gnd cell_6t
Xbit_r119_c132 bl[132] br[132] wl[119] vdd gnd cell_6t
Xbit_r120_c132 bl[132] br[132] wl[120] vdd gnd cell_6t
Xbit_r121_c132 bl[132] br[132] wl[121] vdd gnd cell_6t
Xbit_r122_c132 bl[132] br[132] wl[122] vdd gnd cell_6t
Xbit_r123_c132 bl[132] br[132] wl[123] vdd gnd cell_6t
Xbit_r124_c132 bl[132] br[132] wl[124] vdd gnd cell_6t
Xbit_r125_c132 bl[132] br[132] wl[125] vdd gnd cell_6t
Xbit_r126_c132 bl[132] br[132] wl[126] vdd gnd cell_6t
Xbit_r127_c132 bl[132] br[132] wl[127] vdd gnd cell_6t
Xbit_r0_c133 bl[133] br[133] wl[0] vdd gnd cell_6t
Xbit_r1_c133 bl[133] br[133] wl[1] vdd gnd cell_6t
Xbit_r2_c133 bl[133] br[133] wl[2] vdd gnd cell_6t
Xbit_r3_c133 bl[133] br[133] wl[3] vdd gnd cell_6t
Xbit_r4_c133 bl[133] br[133] wl[4] vdd gnd cell_6t
Xbit_r5_c133 bl[133] br[133] wl[5] vdd gnd cell_6t
Xbit_r6_c133 bl[133] br[133] wl[6] vdd gnd cell_6t
Xbit_r7_c133 bl[133] br[133] wl[7] vdd gnd cell_6t
Xbit_r8_c133 bl[133] br[133] wl[8] vdd gnd cell_6t
Xbit_r9_c133 bl[133] br[133] wl[9] vdd gnd cell_6t
Xbit_r10_c133 bl[133] br[133] wl[10] vdd gnd cell_6t
Xbit_r11_c133 bl[133] br[133] wl[11] vdd gnd cell_6t
Xbit_r12_c133 bl[133] br[133] wl[12] vdd gnd cell_6t
Xbit_r13_c133 bl[133] br[133] wl[13] vdd gnd cell_6t
Xbit_r14_c133 bl[133] br[133] wl[14] vdd gnd cell_6t
Xbit_r15_c133 bl[133] br[133] wl[15] vdd gnd cell_6t
Xbit_r16_c133 bl[133] br[133] wl[16] vdd gnd cell_6t
Xbit_r17_c133 bl[133] br[133] wl[17] vdd gnd cell_6t
Xbit_r18_c133 bl[133] br[133] wl[18] vdd gnd cell_6t
Xbit_r19_c133 bl[133] br[133] wl[19] vdd gnd cell_6t
Xbit_r20_c133 bl[133] br[133] wl[20] vdd gnd cell_6t
Xbit_r21_c133 bl[133] br[133] wl[21] vdd gnd cell_6t
Xbit_r22_c133 bl[133] br[133] wl[22] vdd gnd cell_6t
Xbit_r23_c133 bl[133] br[133] wl[23] vdd gnd cell_6t
Xbit_r24_c133 bl[133] br[133] wl[24] vdd gnd cell_6t
Xbit_r25_c133 bl[133] br[133] wl[25] vdd gnd cell_6t
Xbit_r26_c133 bl[133] br[133] wl[26] vdd gnd cell_6t
Xbit_r27_c133 bl[133] br[133] wl[27] vdd gnd cell_6t
Xbit_r28_c133 bl[133] br[133] wl[28] vdd gnd cell_6t
Xbit_r29_c133 bl[133] br[133] wl[29] vdd gnd cell_6t
Xbit_r30_c133 bl[133] br[133] wl[30] vdd gnd cell_6t
Xbit_r31_c133 bl[133] br[133] wl[31] vdd gnd cell_6t
Xbit_r32_c133 bl[133] br[133] wl[32] vdd gnd cell_6t
Xbit_r33_c133 bl[133] br[133] wl[33] vdd gnd cell_6t
Xbit_r34_c133 bl[133] br[133] wl[34] vdd gnd cell_6t
Xbit_r35_c133 bl[133] br[133] wl[35] vdd gnd cell_6t
Xbit_r36_c133 bl[133] br[133] wl[36] vdd gnd cell_6t
Xbit_r37_c133 bl[133] br[133] wl[37] vdd gnd cell_6t
Xbit_r38_c133 bl[133] br[133] wl[38] vdd gnd cell_6t
Xbit_r39_c133 bl[133] br[133] wl[39] vdd gnd cell_6t
Xbit_r40_c133 bl[133] br[133] wl[40] vdd gnd cell_6t
Xbit_r41_c133 bl[133] br[133] wl[41] vdd gnd cell_6t
Xbit_r42_c133 bl[133] br[133] wl[42] vdd gnd cell_6t
Xbit_r43_c133 bl[133] br[133] wl[43] vdd gnd cell_6t
Xbit_r44_c133 bl[133] br[133] wl[44] vdd gnd cell_6t
Xbit_r45_c133 bl[133] br[133] wl[45] vdd gnd cell_6t
Xbit_r46_c133 bl[133] br[133] wl[46] vdd gnd cell_6t
Xbit_r47_c133 bl[133] br[133] wl[47] vdd gnd cell_6t
Xbit_r48_c133 bl[133] br[133] wl[48] vdd gnd cell_6t
Xbit_r49_c133 bl[133] br[133] wl[49] vdd gnd cell_6t
Xbit_r50_c133 bl[133] br[133] wl[50] vdd gnd cell_6t
Xbit_r51_c133 bl[133] br[133] wl[51] vdd gnd cell_6t
Xbit_r52_c133 bl[133] br[133] wl[52] vdd gnd cell_6t
Xbit_r53_c133 bl[133] br[133] wl[53] vdd gnd cell_6t
Xbit_r54_c133 bl[133] br[133] wl[54] vdd gnd cell_6t
Xbit_r55_c133 bl[133] br[133] wl[55] vdd gnd cell_6t
Xbit_r56_c133 bl[133] br[133] wl[56] vdd gnd cell_6t
Xbit_r57_c133 bl[133] br[133] wl[57] vdd gnd cell_6t
Xbit_r58_c133 bl[133] br[133] wl[58] vdd gnd cell_6t
Xbit_r59_c133 bl[133] br[133] wl[59] vdd gnd cell_6t
Xbit_r60_c133 bl[133] br[133] wl[60] vdd gnd cell_6t
Xbit_r61_c133 bl[133] br[133] wl[61] vdd gnd cell_6t
Xbit_r62_c133 bl[133] br[133] wl[62] vdd gnd cell_6t
Xbit_r63_c133 bl[133] br[133] wl[63] vdd gnd cell_6t
Xbit_r64_c133 bl[133] br[133] wl[64] vdd gnd cell_6t
Xbit_r65_c133 bl[133] br[133] wl[65] vdd gnd cell_6t
Xbit_r66_c133 bl[133] br[133] wl[66] vdd gnd cell_6t
Xbit_r67_c133 bl[133] br[133] wl[67] vdd gnd cell_6t
Xbit_r68_c133 bl[133] br[133] wl[68] vdd gnd cell_6t
Xbit_r69_c133 bl[133] br[133] wl[69] vdd gnd cell_6t
Xbit_r70_c133 bl[133] br[133] wl[70] vdd gnd cell_6t
Xbit_r71_c133 bl[133] br[133] wl[71] vdd gnd cell_6t
Xbit_r72_c133 bl[133] br[133] wl[72] vdd gnd cell_6t
Xbit_r73_c133 bl[133] br[133] wl[73] vdd gnd cell_6t
Xbit_r74_c133 bl[133] br[133] wl[74] vdd gnd cell_6t
Xbit_r75_c133 bl[133] br[133] wl[75] vdd gnd cell_6t
Xbit_r76_c133 bl[133] br[133] wl[76] vdd gnd cell_6t
Xbit_r77_c133 bl[133] br[133] wl[77] vdd gnd cell_6t
Xbit_r78_c133 bl[133] br[133] wl[78] vdd gnd cell_6t
Xbit_r79_c133 bl[133] br[133] wl[79] vdd gnd cell_6t
Xbit_r80_c133 bl[133] br[133] wl[80] vdd gnd cell_6t
Xbit_r81_c133 bl[133] br[133] wl[81] vdd gnd cell_6t
Xbit_r82_c133 bl[133] br[133] wl[82] vdd gnd cell_6t
Xbit_r83_c133 bl[133] br[133] wl[83] vdd gnd cell_6t
Xbit_r84_c133 bl[133] br[133] wl[84] vdd gnd cell_6t
Xbit_r85_c133 bl[133] br[133] wl[85] vdd gnd cell_6t
Xbit_r86_c133 bl[133] br[133] wl[86] vdd gnd cell_6t
Xbit_r87_c133 bl[133] br[133] wl[87] vdd gnd cell_6t
Xbit_r88_c133 bl[133] br[133] wl[88] vdd gnd cell_6t
Xbit_r89_c133 bl[133] br[133] wl[89] vdd gnd cell_6t
Xbit_r90_c133 bl[133] br[133] wl[90] vdd gnd cell_6t
Xbit_r91_c133 bl[133] br[133] wl[91] vdd gnd cell_6t
Xbit_r92_c133 bl[133] br[133] wl[92] vdd gnd cell_6t
Xbit_r93_c133 bl[133] br[133] wl[93] vdd gnd cell_6t
Xbit_r94_c133 bl[133] br[133] wl[94] vdd gnd cell_6t
Xbit_r95_c133 bl[133] br[133] wl[95] vdd gnd cell_6t
Xbit_r96_c133 bl[133] br[133] wl[96] vdd gnd cell_6t
Xbit_r97_c133 bl[133] br[133] wl[97] vdd gnd cell_6t
Xbit_r98_c133 bl[133] br[133] wl[98] vdd gnd cell_6t
Xbit_r99_c133 bl[133] br[133] wl[99] vdd gnd cell_6t
Xbit_r100_c133 bl[133] br[133] wl[100] vdd gnd cell_6t
Xbit_r101_c133 bl[133] br[133] wl[101] vdd gnd cell_6t
Xbit_r102_c133 bl[133] br[133] wl[102] vdd gnd cell_6t
Xbit_r103_c133 bl[133] br[133] wl[103] vdd gnd cell_6t
Xbit_r104_c133 bl[133] br[133] wl[104] vdd gnd cell_6t
Xbit_r105_c133 bl[133] br[133] wl[105] vdd gnd cell_6t
Xbit_r106_c133 bl[133] br[133] wl[106] vdd gnd cell_6t
Xbit_r107_c133 bl[133] br[133] wl[107] vdd gnd cell_6t
Xbit_r108_c133 bl[133] br[133] wl[108] vdd gnd cell_6t
Xbit_r109_c133 bl[133] br[133] wl[109] vdd gnd cell_6t
Xbit_r110_c133 bl[133] br[133] wl[110] vdd gnd cell_6t
Xbit_r111_c133 bl[133] br[133] wl[111] vdd gnd cell_6t
Xbit_r112_c133 bl[133] br[133] wl[112] vdd gnd cell_6t
Xbit_r113_c133 bl[133] br[133] wl[113] vdd gnd cell_6t
Xbit_r114_c133 bl[133] br[133] wl[114] vdd gnd cell_6t
Xbit_r115_c133 bl[133] br[133] wl[115] vdd gnd cell_6t
Xbit_r116_c133 bl[133] br[133] wl[116] vdd gnd cell_6t
Xbit_r117_c133 bl[133] br[133] wl[117] vdd gnd cell_6t
Xbit_r118_c133 bl[133] br[133] wl[118] vdd gnd cell_6t
Xbit_r119_c133 bl[133] br[133] wl[119] vdd gnd cell_6t
Xbit_r120_c133 bl[133] br[133] wl[120] vdd gnd cell_6t
Xbit_r121_c133 bl[133] br[133] wl[121] vdd gnd cell_6t
Xbit_r122_c133 bl[133] br[133] wl[122] vdd gnd cell_6t
Xbit_r123_c133 bl[133] br[133] wl[123] vdd gnd cell_6t
Xbit_r124_c133 bl[133] br[133] wl[124] vdd gnd cell_6t
Xbit_r125_c133 bl[133] br[133] wl[125] vdd gnd cell_6t
Xbit_r126_c133 bl[133] br[133] wl[126] vdd gnd cell_6t
Xbit_r127_c133 bl[133] br[133] wl[127] vdd gnd cell_6t
Xbit_r0_c134 bl[134] br[134] wl[0] vdd gnd cell_6t
Xbit_r1_c134 bl[134] br[134] wl[1] vdd gnd cell_6t
Xbit_r2_c134 bl[134] br[134] wl[2] vdd gnd cell_6t
Xbit_r3_c134 bl[134] br[134] wl[3] vdd gnd cell_6t
Xbit_r4_c134 bl[134] br[134] wl[4] vdd gnd cell_6t
Xbit_r5_c134 bl[134] br[134] wl[5] vdd gnd cell_6t
Xbit_r6_c134 bl[134] br[134] wl[6] vdd gnd cell_6t
Xbit_r7_c134 bl[134] br[134] wl[7] vdd gnd cell_6t
Xbit_r8_c134 bl[134] br[134] wl[8] vdd gnd cell_6t
Xbit_r9_c134 bl[134] br[134] wl[9] vdd gnd cell_6t
Xbit_r10_c134 bl[134] br[134] wl[10] vdd gnd cell_6t
Xbit_r11_c134 bl[134] br[134] wl[11] vdd gnd cell_6t
Xbit_r12_c134 bl[134] br[134] wl[12] vdd gnd cell_6t
Xbit_r13_c134 bl[134] br[134] wl[13] vdd gnd cell_6t
Xbit_r14_c134 bl[134] br[134] wl[14] vdd gnd cell_6t
Xbit_r15_c134 bl[134] br[134] wl[15] vdd gnd cell_6t
Xbit_r16_c134 bl[134] br[134] wl[16] vdd gnd cell_6t
Xbit_r17_c134 bl[134] br[134] wl[17] vdd gnd cell_6t
Xbit_r18_c134 bl[134] br[134] wl[18] vdd gnd cell_6t
Xbit_r19_c134 bl[134] br[134] wl[19] vdd gnd cell_6t
Xbit_r20_c134 bl[134] br[134] wl[20] vdd gnd cell_6t
Xbit_r21_c134 bl[134] br[134] wl[21] vdd gnd cell_6t
Xbit_r22_c134 bl[134] br[134] wl[22] vdd gnd cell_6t
Xbit_r23_c134 bl[134] br[134] wl[23] vdd gnd cell_6t
Xbit_r24_c134 bl[134] br[134] wl[24] vdd gnd cell_6t
Xbit_r25_c134 bl[134] br[134] wl[25] vdd gnd cell_6t
Xbit_r26_c134 bl[134] br[134] wl[26] vdd gnd cell_6t
Xbit_r27_c134 bl[134] br[134] wl[27] vdd gnd cell_6t
Xbit_r28_c134 bl[134] br[134] wl[28] vdd gnd cell_6t
Xbit_r29_c134 bl[134] br[134] wl[29] vdd gnd cell_6t
Xbit_r30_c134 bl[134] br[134] wl[30] vdd gnd cell_6t
Xbit_r31_c134 bl[134] br[134] wl[31] vdd gnd cell_6t
Xbit_r32_c134 bl[134] br[134] wl[32] vdd gnd cell_6t
Xbit_r33_c134 bl[134] br[134] wl[33] vdd gnd cell_6t
Xbit_r34_c134 bl[134] br[134] wl[34] vdd gnd cell_6t
Xbit_r35_c134 bl[134] br[134] wl[35] vdd gnd cell_6t
Xbit_r36_c134 bl[134] br[134] wl[36] vdd gnd cell_6t
Xbit_r37_c134 bl[134] br[134] wl[37] vdd gnd cell_6t
Xbit_r38_c134 bl[134] br[134] wl[38] vdd gnd cell_6t
Xbit_r39_c134 bl[134] br[134] wl[39] vdd gnd cell_6t
Xbit_r40_c134 bl[134] br[134] wl[40] vdd gnd cell_6t
Xbit_r41_c134 bl[134] br[134] wl[41] vdd gnd cell_6t
Xbit_r42_c134 bl[134] br[134] wl[42] vdd gnd cell_6t
Xbit_r43_c134 bl[134] br[134] wl[43] vdd gnd cell_6t
Xbit_r44_c134 bl[134] br[134] wl[44] vdd gnd cell_6t
Xbit_r45_c134 bl[134] br[134] wl[45] vdd gnd cell_6t
Xbit_r46_c134 bl[134] br[134] wl[46] vdd gnd cell_6t
Xbit_r47_c134 bl[134] br[134] wl[47] vdd gnd cell_6t
Xbit_r48_c134 bl[134] br[134] wl[48] vdd gnd cell_6t
Xbit_r49_c134 bl[134] br[134] wl[49] vdd gnd cell_6t
Xbit_r50_c134 bl[134] br[134] wl[50] vdd gnd cell_6t
Xbit_r51_c134 bl[134] br[134] wl[51] vdd gnd cell_6t
Xbit_r52_c134 bl[134] br[134] wl[52] vdd gnd cell_6t
Xbit_r53_c134 bl[134] br[134] wl[53] vdd gnd cell_6t
Xbit_r54_c134 bl[134] br[134] wl[54] vdd gnd cell_6t
Xbit_r55_c134 bl[134] br[134] wl[55] vdd gnd cell_6t
Xbit_r56_c134 bl[134] br[134] wl[56] vdd gnd cell_6t
Xbit_r57_c134 bl[134] br[134] wl[57] vdd gnd cell_6t
Xbit_r58_c134 bl[134] br[134] wl[58] vdd gnd cell_6t
Xbit_r59_c134 bl[134] br[134] wl[59] vdd gnd cell_6t
Xbit_r60_c134 bl[134] br[134] wl[60] vdd gnd cell_6t
Xbit_r61_c134 bl[134] br[134] wl[61] vdd gnd cell_6t
Xbit_r62_c134 bl[134] br[134] wl[62] vdd gnd cell_6t
Xbit_r63_c134 bl[134] br[134] wl[63] vdd gnd cell_6t
Xbit_r64_c134 bl[134] br[134] wl[64] vdd gnd cell_6t
Xbit_r65_c134 bl[134] br[134] wl[65] vdd gnd cell_6t
Xbit_r66_c134 bl[134] br[134] wl[66] vdd gnd cell_6t
Xbit_r67_c134 bl[134] br[134] wl[67] vdd gnd cell_6t
Xbit_r68_c134 bl[134] br[134] wl[68] vdd gnd cell_6t
Xbit_r69_c134 bl[134] br[134] wl[69] vdd gnd cell_6t
Xbit_r70_c134 bl[134] br[134] wl[70] vdd gnd cell_6t
Xbit_r71_c134 bl[134] br[134] wl[71] vdd gnd cell_6t
Xbit_r72_c134 bl[134] br[134] wl[72] vdd gnd cell_6t
Xbit_r73_c134 bl[134] br[134] wl[73] vdd gnd cell_6t
Xbit_r74_c134 bl[134] br[134] wl[74] vdd gnd cell_6t
Xbit_r75_c134 bl[134] br[134] wl[75] vdd gnd cell_6t
Xbit_r76_c134 bl[134] br[134] wl[76] vdd gnd cell_6t
Xbit_r77_c134 bl[134] br[134] wl[77] vdd gnd cell_6t
Xbit_r78_c134 bl[134] br[134] wl[78] vdd gnd cell_6t
Xbit_r79_c134 bl[134] br[134] wl[79] vdd gnd cell_6t
Xbit_r80_c134 bl[134] br[134] wl[80] vdd gnd cell_6t
Xbit_r81_c134 bl[134] br[134] wl[81] vdd gnd cell_6t
Xbit_r82_c134 bl[134] br[134] wl[82] vdd gnd cell_6t
Xbit_r83_c134 bl[134] br[134] wl[83] vdd gnd cell_6t
Xbit_r84_c134 bl[134] br[134] wl[84] vdd gnd cell_6t
Xbit_r85_c134 bl[134] br[134] wl[85] vdd gnd cell_6t
Xbit_r86_c134 bl[134] br[134] wl[86] vdd gnd cell_6t
Xbit_r87_c134 bl[134] br[134] wl[87] vdd gnd cell_6t
Xbit_r88_c134 bl[134] br[134] wl[88] vdd gnd cell_6t
Xbit_r89_c134 bl[134] br[134] wl[89] vdd gnd cell_6t
Xbit_r90_c134 bl[134] br[134] wl[90] vdd gnd cell_6t
Xbit_r91_c134 bl[134] br[134] wl[91] vdd gnd cell_6t
Xbit_r92_c134 bl[134] br[134] wl[92] vdd gnd cell_6t
Xbit_r93_c134 bl[134] br[134] wl[93] vdd gnd cell_6t
Xbit_r94_c134 bl[134] br[134] wl[94] vdd gnd cell_6t
Xbit_r95_c134 bl[134] br[134] wl[95] vdd gnd cell_6t
Xbit_r96_c134 bl[134] br[134] wl[96] vdd gnd cell_6t
Xbit_r97_c134 bl[134] br[134] wl[97] vdd gnd cell_6t
Xbit_r98_c134 bl[134] br[134] wl[98] vdd gnd cell_6t
Xbit_r99_c134 bl[134] br[134] wl[99] vdd gnd cell_6t
Xbit_r100_c134 bl[134] br[134] wl[100] vdd gnd cell_6t
Xbit_r101_c134 bl[134] br[134] wl[101] vdd gnd cell_6t
Xbit_r102_c134 bl[134] br[134] wl[102] vdd gnd cell_6t
Xbit_r103_c134 bl[134] br[134] wl[103] vdd gnd cell_6t
Xbit_r104_c134 bl[134] br[134] wl[104] vdd gnd cell_6t
Xbit_r105_c134 bl[134] br[134] wl[105] vdd gnd cell_6t
Xbit_r106_c134 bl[134] br[134] wl[106] vdd gnd cell_6t
Xbit_r107_c134 bl[134] br[134] wl[107] vdd gnd cell_6t
Xbit_r108_c134 bl[134] br[134] wl[108] vdd gnd cell_6t
Xbit_r109_c134 bl[134] br[134] wl[109] vdd gnd cell_6t
Xbit_r110_c134 bl[134] br[134] wl[110] vdd gnd cell_6t
Xbit_r111_c134 bl[134] br[134] wl[111] vdd gnd cell_6t
Xbit_r112_c134 bl[134] br[134] wl[112] vdd gnd cell_6t
Xbit_r113_c134 bl[134] br[134] wl[113] vdd gnd cell_6t
Xbit_r114_c134 bl[134] br[134] wl[114] vdd gnd cell_6t
Xbit_r115_c134 bl[134] br[134] wl[115] vdd gnd cell_6t
Xbit_r116_c134 bl[134] br[134] wl[116] vdd gnd cell_6t
Xbit_r117_c134 bl[134] br[134] wl[117] vdd gnd cell_6t
Xbit_r118_c134 bl[134] br[134] wl[118] vdd gnd cell_6t
Xbit_r119_c134 bl[134] br[134] wl[119] vdd gnd cell_6t
Xbit_r120_c134 bl[134] br[134] wl[120] vdd gnd cell_6t
Xbit_r121_c134 bl[134] br[134] wl[121] vdd gnd cell_6t
Xbit_r122_c134 bl[134] br[134] wl[122] vdd gnd cell_6t
Xbit_r123_c134 bl[134] br[134] wl[123] vdd gnd cell_6t
Xbit_r124_c134 bl[134] br[134] wl[124] vdd gnd cell_6t
Xbit_r125_c134 bl[134] br[134] wl[125] vdd gnd cell_6t
Xbit_r126_c134 bl[134] br[134] wl[126] vdd gnd cell_6t
Xbit_r127_c134 bl[134] br[134] wl[127] vdd gnd cell_6t
Xbit_r0_c135 bl[135] br[135] wl[0] vdd gnd cell_6t
Xbit_r1_c135 bl[135] br[135] wl[1] vdd gnd cell_6t
Xbit_r2_c135 bl[135] br[135] wl[2] vdd gnd cell_6t
Xbit_r3_c135 bl[135] br[135] wl[3] vdd gnd cell_6t
Xbit_r4_c135 bl[135] br[135] wl[4] vdd gnd cell_6t
Xbit_r5_c135 bl[135] br[135] wl[5] vdd gnd cell_6t
Xbit_r6_c135 bl[135] br[135] wl[6] vdd gnd cell_6t
Xbit_r7_c135 bl[135] br[135] wl[7] vdd gnd cell_6t
Xbit_r8_c135 bl[135] br[135] wl[8] vdd gnd cell_6t
Xbit_r9_c135 bl[135] br[135] wl[9] vdd gnd cell_6t
Xbit_r10_c135 bl[135] br[135] wl[10] vdd gnd cell_6t
Xbit_r11_c135 bl[135] br[135] wl[11] vdd gnd cell_6t
Xbit_r12_c135 bl[135] br[135] wl[12] vdd gnd cell_6t
Xbit_r13_c135 bl[135] br[135] wl[13] vdd gnd cell_6t
Xbit_r14_c135 bl[135] br[135] wl[14] vdd gnd cell_6t
Xbit_r15_c135 bl[135] br[135] wl[15] vdd gnd cell_6t
Xbit_r16_c135 bl[135] br[135] wl[16] vdd gnd cell_6t
Xbit_r17_c135 bl[135] br[135] wl[17] vdd gnd cell_6t
Xbit_r18_c135 bl[135] br[135] wl[18] vdd gnd cell_6t
Xbit_r19_c135 bl[135] br[135] wl[19] vdd gnd cell_6t
Xbit_r20_c135 bl[135] br[135] wl[20] vdd gnd cell_6t
Xbit_r21_c135 bl[135] br[135] wl[21] vdd gnd cell_6t
Xbit_r22_c135 bl[135] br[135] wl[22] vdd gnd cell_6t
Xbit_r23_c135 bl[135] br[135] wl[23] vdd gnd cell_6t
Xbit_r24_c135 bl[135] br[135] wl[24] vdd gnd cell_6t
Xbit_r25_c135 bl[135] br[135] wl[25] vdd gnd cell_6t
Xbit_r26_c135 bl[135] br[135] wl[26] vdd gnd cell_6t
Xbit_r27_c135 bl[135] br[135] wl[27] vdd gnd cell_6t
Xbit_r28_c135 bl[135] br[135] wl[28] vdd gnd cell_6t
Xbit_r29_c135 bl[135] br[135] wl[29] vdd gnd cell_6t
Xbit_r30_c135 bl[135] br[135] wl[30] vdd gnd cell_6t
Xbit_r31_c135 bl[135] br[135] wl[31] vdd gnd cell_6t
Xbit_r32_c135 bl[135] br[135] wl[32] vdd gnd cell_6t
Xbit_r33_c135 bl[135] br[135] wl[33] vdd gnd cell_6t
Xbit_r34_c135 bl[135] br[135] wl[34] vdd gnd cell_6t
Xbit_r35_c135 bl[135] br[135] wl[35] vdd gnd cell_6t
Xbit_r36_c135 bl[135] br[135] wl[36] vdd gnd cell_6t
Xbit_r37_c135 bl[135] br[135] wl[37] vdd gnd cell_6t
Xbit_r38_c135 bl[135] br[135] wl[38] vdd gnd cell_6t
Xbit_r39_c135 bl[135] br[135] wl[39] vdd gnd cell_6t
Xbit_r40_c135 bl[135] br[135] wl[40] vdd gnd cell_6t
Xbit_r41_c135 bl[135] br[135] wl[41] vdd gnd cell_6t
Xbit_r42_c135 bl[135] br[135] wl[42] vdd gnd cell_6t
Xbit_r43_c135 bl[135] br[135] wl[43] vdd gnd cell_6t
Xbit_r44_c135 bl[135] br[135] wl[44] vdd gnd cell_6t
Xbit_r45_c135 bl[135] br[135] wl[45] vdd gnd cell_6t
Xbit_r46_c135 bl[135] br[135] wl[46] vdd gnd cell_6t
Xbit_r47_c135 bl[135] br[135] wl[47] vdd gnd cell_6t
Xbit_r48_c135 bl[135] br[135] wl[48] vdd gnd cell_6t
Xbit_r49_c135 bl[135] br[135] wl[49] vdd gnd cell_6t
Xbit_r50_c135 bl[135] br[135] wl[50] vdd gnd cell_6t
Xbit_r51_c135 bl[135] br[135] wl[51] vdd gnd cell_6t
Xbit_r52_c135 bl[135] br[135] wl[52] vdd gnd cell_6t
Xbit_r53_c135 bl[135] br[135] wl[53] vdd gnd cell_6t
Xbit_r54_c135 bl[135] br[135] wl[54] vdd gnd cell_6t
Xbit_r55_c135 bl[135] br[135] wl[55] vdd gnd cell_6t
Xbit_r56_c135 bl[135] br[135] wl[56] vdd gnd cell_6t
Xbit_r57_c135 bl[135] br[135] wl[57] vdd gnd cell_6t
Xbit_r58_c135 bl[135] br[135] wl[58] vdd gnd cell_6t
Xbit_r59_c135 bl[135] br[135] wl[59] vdd gnd cell_6t
Xbit_r60_c135 bl[135] br[135] wl[60] vdd gnd cell_6t
Xbit_r61_c135 bl[135] br[135] wl[61] vdd gnd cell_6t
Xbit_r62_c135 bl[135] br[135] wl[62] vdd gnd cell_6t
Xbit_r63_c135 bl[135] br[135] wl[63] vdd gnd cell_6t
Xbit_r64_c135 bl[135] br[135] wl[64] vdd gnd cell_6t
Xbit_r65_c135 bl[135] br[135] wl[65] vdd gnd cell_6t
Xbit_r66_c135 bl[135] br[135] wl[66] vdd gnd cell_6t
Xbit_r67_c135 bl[135] br[135] wl[67] vdd gnd cell_6t
Xbit_r68_c135 bl[135] br[135] wl[68] vdd gnd cell_6t
Xbit_r69_c135 bl[135] br[135] wl[69] vdd gnd cell_6t
Xbit_r70_c135 bl[135] br[135] wl[70] vdd gnd cell_6t
Xbit_r71_c135 bl[135] br[135] wl[71] vdd gnd cell_6t
Xbit_r72_c135 bl[135] br[135] wl[72] vdd gnd cell_6t
Xbit_r73_c135 bl[135] br[135] wl[73] vdd gnd cell_6t
Xbit_r74_c135 bl[135] br[135] wl[74] vdd gnd cell_6t
Xbit_r75_c135 bl[135] br[135] wl[75] vdd gnd cell_6t
Xbit_r76_c135 bl[135] br[135] wl[76] vdd gnd cell_6t
Xbit_r77_c135 bl[135] br[135] wl[77] vdd gnd cell_6t
Xbit_r78_c135 bl[135] br[135] wl[78] vdd gnd cell_6t
Xbit_r79_c135 bl[135] br[135] wl[79] vdd gnd cell_6t
Xbit_r80_c135 bl[135] br[135] wl[80] vdd gnd cell_6t
Xbit_r81_c135 bl[135] br[135] wl[81] vdd gnd cell_6t
Xbit_r82_c135 bl[135] br[135] wl[82] vdd gnd cell_6t
Xbit_r83_c135 bl[135] br[135] wl[83] vdd gnd cell_6t
Xbit_r84_c135 bl[135] br[135] wl[84] vdd gnd cell_6t
Xbit_r85_c135 bl[135] br[135] wl[85] vdd gnd cell_6t
Xbit_r86_c135 bl[135] br[135] wl[86] vdd gnd cell_6t
Xbit_r87_c135 bl[135] br[135] wl[87] vdd gnd cell_6t
Xbit_r88_c135 bl[135] br[135] wl[88] vdd gnd cell_6t
Xbit_r89_c135 bl[135] br[135] wl[89] vdd gnd cell_6t
Xbit_r90_c135 bl[135] br[135] wl[90] vdd gnd cell_6t
Xbit_r91_c135 bl[135] br[135] wl[91] vdd gnd cell_6t
Xbit_r92_c135 bl[135] br[135] wl[92] vdd gnd cell_6t
Xbit_r93_c135 bl[135] br[135] wl[93] vdd gnd cell_6t
Xbit_r94_c135 bl[135] br[135] wl[94] vdd gnd cell_6t
Xbit_r95_c135 bl[135] br[135] wl[95] vdd gnd cell_6t
Xbit_r96_c135 bl[135] br[135] wl[96] vdd gnd cell_6t
Xbit_r97_c135 bl[135] br[135] wl[97] vdd gnd cell_6t
Xbit_r98_c135 bl[135] br[135] wl[98] vdd gnd cell_6t
Xbit_r99_c135 bl[135] br[135] wl[99] vdd gnd cell_6t
Xbit_r100_c135 bl[135] br[135] wl[100] vdd gnd cell_6t
Xbit_r101_c135 bl[135] br[135] wl[101] vdd gnd cell_6t
Xbit_r102_c135 bl[135] br[135] wl[102] vdd gnd cell_6t
Xbit_r103_c135 bl[135] br[135] wl[103] vdd gnd cell_6t
Xbit_r104_c135 bl[135] br[135] wl[104] vdd gnd cell_6t
Xbit_r105_c135 bl[135] br[135] wl[105] vdd gnd cell_6t
Xbit_r106_c135 bl[135] br[135] wl[106] vdd gnd cell_6t
Xbit_r107_c135 bl[135] br[135] wl[107] vdd gnd cell_6t
Xbit_r108_c135 bl[135] br[135] wl[108] vdd gnd cell_6t
Xbit_r109_c135 bl[135] br[135] wl[109] vdd gnd cell_6t
Xbit_r110_c135 bl[135] br[135] wl[110] vdd gnd cell_6t
Xbit_r111_c135 bl[135] br[135] wl[111] vdd gnd cell_6t
Xbit_r112_c135 bl[135] br[135] wl[112] vdd gnd cell_6t
Xbit_r113_c135 bl[135] br[135] wl[113] vdd gnd cell_6t
Xbit_r114_c135 bl[135] br[135] wl[114] vdd gnd cell_6t
Xbit_r115_c135 bl[135] br[135] wl[115] vdd gnd cell_6t
Xbit_r116_c135 bl[135] br[135] wl[116] vdd gnd cell_6t
Xbit_r117_c135 bl[135] br[135] wl[117] vdd gnd cell_6t
Xbit_r118_c135 bl[135] br[135] wl[118] vdd gnd cell_6t
Xbit_r119_c135 bl[135] br[135] wl[119] vdd gnd cell_6t
Xbit_r120_c135 bl[135] br[135] wl[120] vdd gnd cell_6t
Xbit_r121_c135 bl[135] br[135] wl[121] vdd gnd cell_6t
Xbit_r122_c135 bl[135] br[135] wl[122] vdd gnd cell_6t
Xbit_r123_c135 bl[135] br[135] wl[123] vdd gnd cell_6t
Xbit_r124_c135 bl[135] br[135] wl[124] vdd gnd cell_6t
Xbit_r125_c135 bl[135] br[135] wl[125] vdd gnd cell_6t
Xbit_r126_c135 bl[135] br[135] wl[126] vdd gnd cell_6t
Xbit_r127_c135 bl[135] br[135] wl[127] vdd gnd cell_6t
Xbit_r0_c136 bl[136] br[136] wl[0] vdd gnd cell_6t
Xbit_r1_c136 bl[136] br[136] wl[1] vdd gnd cell_6t
Xbit_r2_c136 bl[136] br[136] wl[2] vdd gnd cell_6t
Xbit_r3_c136 bl[136] br[136] wl[3] vdd gnd cell_6t
Xbit_r4_c136 bl[136] br[136] wl[4] vdd gnd cell_6t
Xbit_r5_c136 bl[136] br[136] wl[5] vdd gnd cell_6t
Xbit_r6_c136 bl[136] br[136] wl[6] vdd gnd cell_6t
Xbit_r7_c136 bl[136] br[136] wl[7] vdd gnd cell_6t
Xbit_r8_c136 bl[136] br[136] wl[8] vdd gnd cell_6t
Xbit_r9_c136 bl[136] br[136] wl[9] vdd gnd cell_6t
Xbit_r10_c136 bl[136] br[136] wl[10] vdd gnd cell_6t
Xbit_r11_c136 bl[136] br[136] wl[11] vdd gnd cell_6t
Xbit_r12_c136 bl[136] br[136] wl[12] vdd gnd cell_6t
Xbit_r13_c136 bl[136] br[136] wl[13] vdd gnd cell_6t
Xbit_r14_c136 bl[136] br[136] wl[14] vdd gnd cell_6t
Xbit_r15_c136 bl[136] br[136] wl[15] vdd gnd cell_6t
Xbit_r16_c136 bl[136] br[136] wl[16] vdd gnd cell_6t
Xbit_r17_c136 bl[136] br[136] wl[17] vdd gnd cell_6t
Xbit_r18_c136 bl[136] br[136] wl[18] vdd gnd cell_6t
Xbit_r19_c136 bl[136] br[136] wl[19] vdd gnd cell_6t
Xbit_r20_c136 bl[136] br[136] wl[20] vdd gnd cell_6t
Xbit_r21_c136 bl[136] br[136] wl[21] vdd gnd cell_6t
Xbit_r22_c136 bl[136] br[136] wl[22] vdd gnd cell_6t
Xbit_r23_c136 bl[136] br[136] wl[23] vdd gnd cell_6t
Xbit_r24_c136 bl[136] br[136] wl[24] vdd gnd cell_6t
Xbit_r25_c136 bl[136] br[136] wl[25] vdd gnd cell_6t
Xbit_r26_c136 bl[136] br[136] wl[26] vdd gnd cell_6t
Xbit_r27_c136 bl[136] br[136] wl[27] vdd gnd cell_6t
Xbit_r28_c136 bl[136] br[136] wl[28] vdd gnd cell_6t
Xbit_r29_c136 bl[136] br[136] wl[29] vdd gnd cell_6t
Xbit_r30_c136 bl[136] br[136] wl[30] vdd gnd cell_6t
Xbit_r31_c136 bl[136] br[136] wl[31] vdd gnd cell_6t
Xbit_r32_c136 bl[136] br[136] wl[32] vdd gnd cell_6t
Xbit_r33_c136 bl[136] br[136] wl[33] vdd gnd cell_6t
Xbit_r34_c136 bl[136] br[136] wl[34] vdd gnd cell_6t
Xbit_r35_c136 bl[136] br[136] wl[35] vdd gnd cell_6t
Xbit_r36_c136 bl[136] br[136] wl[36] vdd gnd cell_6t
Xbit_r37_c136 bl[136] br[136] wl[37] vdd gnd cell_6t
Xbit_r38_c136 bl[136] br[136] wl[38] vdd gnd cell_6t
Xbit_r39_c136 bl[136] br[136] wl[39] vdd gnd cell_6t
Xbit_r40_c136 bl[136] br[136] wl[40] vdd gnd cell_6t
Xbit_r41_c136 bl[136] br[136] wl[41] vdd gnd cell_6t
Xbit_r42_c136 bl[136] br[136] wl[42] vdd gnd cell_6t
Xbit_r43_c136 bl[136] br[136] wl[43] vdd gnd cell_6t
Xbit_r44_c136 bl[136] br[136] wl[44] vdd gnd cell_6t
Xbit_r45_c136 bl[136] br[136] wl[45] vdd gnd cell_6t
Xbit_r46_c136 bl[136] br[136] wl[46] vdd gnd cell_6t
Xbit_r47_c136 bl[136] br[136] wl[47] vdd gnd cell_6t
Xbit_r48_c136 bl[136] br[136] wl[48] vdd gnd cell_6t
Xbit_r49_c136 bl[136] br[136] wl[49] vdd gnd cell_6t
Xbit_r50_c136 bl[136] br[136] wl[50] vdd gnd cell_6t
Xbit_r51_c136 bl[136] br[136] wl[51] vdd gnd cell_6t
Xbit_r52_c136 bl[136] br[136] wl[52] vdd gnd cell_6t
Xbit_r53_c136 bl[136] br[136] wl[53] vdd gnd cell_6t
Xbit_r54_c136 bl[136] br[136] wl[54] vdd gnd cell_6t
Xbit_r55_c136 bl[136] br[136] wl[55] vdd gnd cell_6t
Xbit_r56_c136 bl[136] br[136] wl[56] vdd gnd cell_6t
Xbit_r57_c136 bl[136] br[136] wl[57] vdd gnd cell_6t
Xbit_r58_c136 bl[136] br[136] wl[58] vdd gnd cell_6t
Xbit_r59_c136 bl[136] br[136] wl[59] vdd gnd cell_6t
Xbit_r60_c136 bl[136] br[136] wl[60] vdd gnd cell_6t
Xbit_r61_c136 bl[136] br[136] wl[61] vdd gnd cell_6t
Xbit_r62_c136 bl[136] br[136] wl[62] vdd gnd cell_6t
Xbit_r63_c136 bl[136] br[136] wl[63] vdd gnd cell_6t
Xbit_r64_c136 bl[136] br[136] wl[64] vdd gnd cell_6t
Xbit_r65_c136 bl[136] br[136] wl[65] vdd gnd cell_6t
Xbit_r66_c136 bl[136] br[136] wl[66] vdd gnd cell_6t
Xbit_r67_c136 bl[136] br[136] wl[67] vdd gnd cell_6t
Xbit_r68_c136 bl[136] br[136] wl[68] vdd gnd cell_6t
Xbit_r69_c136 bl[136] br[136] wl[69] vdd gnd cell_6t
Xbit_r70_c136 bl[136] br[136] wl[70] vdd gnd cell_6t
Xbit_r71_c136 bl[136] br[136] wl[71] vdd gnd cell_6t
Xbit_r72_c136 bl[136] br[136] wl[72] vdd gnd cell_6t
Xbit_r73_c136 bl[136] br[136] wl[73] vdd gnd cell_6t
Xbit_r74_c136 bl[136] br[136] wl[74] vdd gnd cell_6t
Xbit_r75_c136 bl[136] br[136] wl[75] vdd gnd cell_6t
Xbit_r76_c136 bl[136] br[136] wl[76] vdd gnd cell_6t
Xbit_r77_c136 bl[136] br[136] wl[77] vdd gnd cell_6t
Xbit_r78_c136 bl[136] br[136] wl[78] vdd gnd cell_6t
Xbit_r79_c136 bl[136] br[136] wl[79] vdd gnd cell_6t
Xbit_r80_c136 bl[136] br[136] wl[80] vdd gnd cell_6t
Xbit_r81_c136 bl[136] br[136] wl[81] vdd gnd cell_6t
Xbit_r82_c136 bl[136] br[136] wl[82] vdd gnd cell_6t
Xbit_r83_c136 bl[136] br[136] wl[83] vdd gnd cell_6t
Xbit_r84_c136 bl[136] br[136] wl[84] vdd gnd cell_6t
Xbit_r85_c136 bl[136] br[136] wl[85] vdd gnd cell_6t
Xbit_r86_c136 bl[136] br[136] wl[86] vdd gnd cell_6t
Xbit_r87_c136 bl[136] br[136] wl[87] vdd gnd cell_6t
Xbit_r88_c136 bl[136] br[136] wl[88] vdd gnd cell_6t
Xbit_r89_c136 bl[136] br[136] wl[89] vdd gnd cell_6t
Xbit_r90_c136 bl[136] br[136] wl[90] vdd gnd cell_6t
Xbit_r91_c136 bl[136] br[136] wl[91] vdd gnd cell_6t
Xbit_r92_c136 bl[136] br[136] wl[92] vdd gnd cell_6t
Xbit_r93_c136 bl[136] br[136] wl[93] vdd gnd cell_6t
Xbit_r94_c136 bl[136] br[136] wl[94] vdd gnd cell_6t
Xbit_r95_c136 bl[136] br[136] wl[95] vdd gnd cell_6t
Xbit_r96_c136 bl[136] br[136] wl[96] vdd gnd cell_6t
Xbit_r97_c136 bl[136] br[136] wl[97] vdd gnd cell_6t
Xbit_r98_c136 bl[136] br[136] wl[98] vdd gnd cell_6t
Xbit_r99_c136 bl[136] br[136] wl[99] vdd gnd cell_6t
Xbit_r100_c136 bl[136] br[136] wl[100] vdd gnd cell_6t
Xbit_r101_c136 bl[136] br[136] wl[101] vdd gnd cell_6t
Xbit_r102_c136 bl[136] br[136] wl[102] vdd gnd cell_6t
Xbit_r103_c136 bl[136] br[136] wl[103] vdd gnd cell_6t
Xbit_r104_c136 bl[136] br[136] wl[104] vdd gnd cell_6t
Xbit_r105_c136 bl[136] br[136] wl[105] vdd gnd cell_6t
Xbit_r106_c136 bl[136] br[136] wl[106] vdd gnd cell_6t
Xbit_r107_c136 bl[136] br[136] wl[107] vdd gnd cell_6t
Xbit_r108_c136 bl[136] br[136] wl[108] vdd gnd cell_6t
Xbit_r109_c136 bl[136] br[136] wl[109] vdd gnd cell_6t
Xbit_r110_c136 bl[136] br[136] wl[110] vdd gnd cell_6t
Xbit_r111_c136 bl[136] br[136] wl[111] vdd gnd cell_6t
Xbit_r112_c136 bl[136] br[136] wl[112] vdd gnd cell_6t
Xbit_r113_c136 bl[136] br[136] wl[113] vdd gnd cell_6t
Xbit_r114_c136 bl[136] br[136] wl[114] vdd gnd cell_6t
Xbit_r115_c136 bl[136] br[136] wl[115] vdd gnd cell_6t
Xbit_r116_c136 bl[136] br[136] wl[116] vdd gnd cell_6t
Xbit_r117_c136 bl[136] br[136] wl[117] vdd gnd cell_6t
Xbit_r118_c136 bl[136] br[136] wl[118] vdd gnd cell_6t
Xbit_r119_c136 bl[136] br[136] wl[119] vdd gnd cell_6t
Xbit_r120_c136 bl[136] br[136] wl[120] vdd gnd cell_6t
Xbit_r121_c136 bl[136] br[136] wl[121] vdd gnd cell_6t
Xbit_r122_c136 bl[136] br[136] wl[122] vdd gnd cell_6t
Xbit_r123_c136 bl[136] br[136] wl[123] vdd gnd cell_6t
Xbit_r124_c136 bl[136] br[136] wl[124] vdd gnd cell_6t
Xbit_r125_c136 bl[136] br[136] wl[125] vdd gnd cell_6t
Xbit_r126_c136 bl[136] br[136] wl[126] vdd gnd cell_6t
Xbit_r127_c136 bl[136] br[136] wl[127] vdd gnd cell_6t
Xbit_r0_c137 bl[137] br[137] wl[0] vdd gnd cell_6t
Xbit_r1_c137 bl[137] br[137] wl[1] vdd gnd cell_6t
Xbit_r2_c137 bl[137] br[137] wl[2] vdd gnd cell_6t
Xbit_r3_c137 bl[137] br[137] wl[3] vdd gnd cell_6t
Xbit_r4_c137 bl[137] br[137] wl[4] vdd gnd cell_6t
Xbit_r5_c137 bl[137] br[137] wl[5] vdd gnd cell_6t
Xbit_r6_c137 bl[137] br[137] wl[6] vdd gnd cell_6t
Xbit_r7_c137 bl[137] br[137] wl[7] vdd gnd cell_6t
Xbit_r8_c137 bl[137] br[137] wl[8] vdd gnd cell_6t
Xbit_r9_c137 bl[137] br[137] wl[9] vdd gnd cell_6t
Xbit_r10_c137 bl[137] br[137] wl[10] vdd gnd cell_6t
Xbit_r11_c137 bl[137] br[137] wl[11] vdd gnd cell_6t
Xbit_r12_c137 bl[137] br[137] wl[12] vdd gnd cell_6t
Xbit_r13_c137 bl[137] br[137] wl[13] vdd gnd cell_6t
Xbit_r14_c137 bl[137] br[137] wl[14] vdd gnd cell_6t
Xbit_r15_c137 bl[137] br[137] wl[15] vdd gnd cell_6t
Xbit_r16_c137 bl[137] br[137] wl[16] vdd gnd cell_6t
Xbit_r17_c137 bl[137] br[137] wl[17] vdd gnd cell_6t
Xbit_r18_c137 bl[137] br[137] wl[18] vdd gnd cell_6t
Xbit_r19_c137 bl[137] br[137] wl[19] vdd gnd cell_6t
Xbit_r20_c137 bl[137] br[137] wl[20] vdd gnd cell_6t
Xbit_r21_c137 bl[137] br[137] wl[21] vdd gnd cell_6t
Xbit_r22_c137 bl[137] br[137] wl[22] vdd gnd cell_6t
Xbit_r23_c137 bl[137] br[137] wl[23] vdd gnd cell_6t
Xbit_r24_c137 bl[137] br[137] wl[24] vdd gnd cell_6t
Xbit_r25_c137 bl[137] br[137] wl[25] vdd gnd cell_6t
Xbit_r26_c137 bl[137] br[137] wl[26] vdd gnd cell_6t
Xbit_r27_c137 bl[137] br[137] wl[27] vdd gnd cell_6t
Xbit_r28_c137 bl[137] br[137] wl[28] vdd gnd cell_6t
Xbit_r29_c137 bl[137] br[137] wl[29] vdd gnd cell_6t
Xbit_r30_c137 bl[137] br[137] wl[30] vdd gnd cell_6t
Xbit_r31_c137 bl[137] br[137] wl[31] vdd gnd cell_6t
Xbit_r32_c137 bl[137] br[137] wl[32] vdd gnd cell_6t
Xbit_r33_c137 bl[137] br[137] wl[33] vdd gnd cell_6t
Xbit_r34_c137 bl[137] br[137] wl[34] vdd gnd cell_6t
Xbit_r35_c137 bl[137] br[137] wl[35] vdd gnd cell_6t
Xbit_r36_c137 bl[137] br[137] wl[36] vdd gnd cell_6t
Xbit_r37_c137 bl[137] br[137] wl[37] vdd gnd cell_6t
Xbit_r38_c137 bl[137] br[137] wl[38] vdd gnd cell_6t
Xbit_r39_c137 bl[137] br[137] wl[39] vdd gnd cell_6t
Xbit_r40_c137 bl[137] br[137] wl[40] vdd gnd cell_6t
Xbit_r41_c137 bl[137] br[137] wl[41] vdd gnd cell_6t
Xbit_r42_c137 bl[137] br[137] wl[42] vdd gnd cell_6t
Xbit_r43_c137 bl[137] br[137] wl[43] vdd gnd cell_6t
Xbit_r44_c137 bl[137] br[137] wl[44] vdd gnd cell_6t
Xbit_r45_c137 bl[137] br[137] wl[45] vdd gnd cell_6t
Xbit_r46_c137 bl[137] br[137] wl[46] vdd gnd cell_6t
Xbit_r47_c137 bl[137] br[137] wl[47] vdd gnd cell_6t
Xbit_r48_c137 bl[137] br[137] wl[48] vdd gnd cell_6t
Xbit_r49_c137 bl[137] br[137] wl[49] vdd gnd cell_6t
Xbit_r50_c137 bl[137] br[137] wl[50] vdd gnd cell_6t
Xbit_r51_c137 bl[137] br[137] wl[51] vdd gnd cell_6t
Xbit_r52_c137 bl[137] br[137] wl[52] vdd gnd cell_6t
Xbit_r53_c137 bl[137] br[137] wl[53] vdd gnd cell_6t
Xbit_r54_c137 bl[137] br[137] wl[54] vdd gnd cell_6t
Xbit_r55_c137 bl[137] br[137] wl[55] vdd gnd cell_6t
Xbit_r56_c137 bl[137] br[137] wl[56] vdd gnd cell_6t
Xbit_r57_c137 bl[137] br[137] wl[57] vdd gnd cell_6t
Xbit_r58_c137 bl[137] br[137] wl[58] vdd gnd cell_6t
Xbit_r59_c137 bl[137] br[137] wl[59] vdd gnd cell_6t
Xbit_r60_c137 bl[137] br[137] wl[60] vdd gnd cell_6t
Xbit_r61_c137 bl[137] br[137] wl[61] vdd gnd cell_6t
Xbit_r62_c137 bl[137] br[137] wl[62] vdd gnd cell_6t
Xbit_r63_c137 bl[137] br[137] wl[63] vdd gnd cell_6t
Xbit_r64_c137 bl[137] br[137] wl[64] vdd gnd cell_6t
Xbit_r65_c137 bl[137] br[137] wl[65] vdd gnd cell_6t
Xbit_r66_c137 bl[137] br[137] wl[66] vdd gnd cell_6t
Xbit_r67_c137 bl[137] br[137] wl[67] vdd gnd cell_6t
Xbit_r68_c137 bl[137] br[137] wl[68] vdd gnd cell_6t
Xbit_r69_c137 bl[137] br[137] wl[69] vdd gnd cell_6t
Xbit_r70_c137 bl[137] br[137] wl[70] vdd gnd cell_6t
Xbit_r71_c137 bl[137] br[137] wl[71] vdd gnd cell_6t
Xbit_r72_c137 bl[137] br[137] wl[72] vdd gnd cell_6t
Xbit_r73_c137 bl[137] br[137] wl[73] vdd gnd cell_6t
Xbit_r74_c137 bl[137] br[137] wl[74] vdd gnd cell_6t
Xbit_r75_c137 bl[137] br[137] wl[75] vdd gnd cell_6t
Xbit_r76_c137 bl[137] br[137] wl[76] vdd gnd cell_6t
Xbit_r77_c137 bl[137] br[137] wl[77] vdd gnd cell_6t
Xbit_r78_c137 bl[137] br[137] wl[78] vdd gnd cell_6t
Xbit_r79_c137 bl[137] br[137] wl[79] vdd gnd cell_6t
Xbit_r80_c137 bl[137] br[137] wl[80] vdd gnd cell_6t
Xbit_r81_c137 bl[137] br[137] wl[81] vdd gnd cell_6t
Xbit_r82_c137 bl[137] br[137] wl[82] vdd gnd cell_6t
Xbit_r83_c137 bl[137] br[137] wl[83] vdd gnd cell_6t
Xbit_r84_c137 bl[137] br[137] wl[84] vdd gnd cell_6t
Xbit_r85_c137 bl[137] br[137] wl[85] vdd gnd cell_6t
Xbit_r86_c137 bl[137] br[137] wl[86] vdd gnd cell_6t
Xbit_r87_c137 bl[137] br[137] wl[87] vdd gnd cell_6t
Xbit_r88_c137 bl[137] br[137] wl[88] vdd gnd cell_6t
Xbit_r89_c137 bl[137] br[137] wl[89] vdd gnd cell_6t
Xbit_r90_c137 bl[137] br[137] wl[90] vdd gnd cell_6t
Xbit_r91_c137 bl[137] br[137] wl[91] vdd gnd cell_6t
Xbit_r92_c137 bl[137] br[137] wl[92] vdd gnd cell_6t
Xbit_r93_c137 bl[137] br[137] wl[93] vdd gnd cell_6t
Xbit_r94_c137 bl[137] br[137] wl[94] vdd gnd cell_6t
Xbit_r95_c137 bl[137] br[137] wl[95] vdd gnd cell_6t
Xbit_r96_c137 bl[137] br[137] wl[96] vdd gnd cell_6t
Xbit_r97_c137 bl[137] br[137] wl[97] vdd gnd cell_6t
Xbit_r98_c137 bl[137] br[137] wl[98] vdd gnd cell_6t
Xbit_r99_c137 bl[137] br[137] wl[99] vdd gnd cell_6t
Xbit_r100_c137 bl[137] br[137] wl[100] vdd gnd cell_6t
Xbit_r101_c137 bl[137] br[137] wl[101] vdd gnd cell_6t
Xbit_r102_c137 bl[137] br[137] wl[102] vdd gnd cell_6t
Xbit_r103_c137 bl[137] br[137] wl[103] vdd gnd cell_6t
Xbit_r104_c137 bl[137] br[137] wl[104] vdd gnd cell_6t
Xbit_r105_c137 bl[137] br[137] wl[105] vdd gnd cell_6t
Xbit_r106_c137 bl[137] br[137] wl[106] vdd gnd cell_6t
Xbit_r107_c137 bl[137] br[137] wl[107] vdd gnd cell_6t
Xbit_r108_c137 bl[137] br[137] wl[108] vdd gnd cell_6t
Xbit_r109_c137 bl[137] br[137] wl[109] vdd gnd cell_6t
Xbit_r110_c137 bl[137] br[137] wl[110] vdd gnd cell_6t
Xbit_r111_c137 bl[137] br[137] wl[111] vdd gnd cell_6t
Xbit_r112_c137 bl[137] br[137] wl[112] vdd gnd cell_6t
Xbit_r113_c137 bl[137] br[137] wl[113] vdd gnd cell_6t
Xbit_r114_c137 bl[137] br[137] wl[114] vdd gnd cell_6t
Xbit_r115_c137 bl[137] br[137] wl[115] vdd gnd cell_6t
Xbit_r116_c137 bl[137] br[137] wl[116] vdd gnd cell_6t
Xbit_r117_c137 bl[137] br[137] wl[117] vdd gnd cell_6t
Xbit_r118_c137 bl[137] br[137] wl[118] vdd gnd cell_6t
Xbit_r119_c137 bl[137] br[137] wl[119] vdd gnd cell_6t
Xbit_r120_c137 bl[137] br[137] wl[120] vdd gnd cell_6t
Xbit_r121_c137 bl[137] br[137] wl[121] vdd gnd cell_6t
Xbit_r122_c137 bl[137] br[137] wl[122] vdd gnd cell_6t
Xbit_r123_c137 bl[137] br[137] wl[123] vdd gnd cell_6t
Xbit_r124_c137 bl[137] br[137] wl[124] vdd gnd cell_6t
Xbit_r125_c137 bl[137] br[137] wl[125] vdd gnd cell_6t
Xbit_r126_c137 bl[137] br[137] wl[126] vdd gnd cell_6t
Xbit_r127_c137 bl[137] br[137] wl[127] vdd gnd cell_6t
Xbit_r0_c138 bl[138] br[138] wl[0] vdd gnd cell_6t
Xbit_r1_c138 bl[138] br[138] wl[1] vdd gnd cell_6t
Xbit_r2_c138 bl[138] br[138] wl[2] vdd gnd cell_6t
Xbit_r3_c138 bl[138] br[138] wl[3] vdd gnd cell_6t
Xbit_r4_c138 bl[138] br[138] wl[4] vdd gnd cell_6t
Xbit_r5_c138 bl[138] br[138] wl[5] vdd gnd cell_6t
Xbit_r6_c138 bl[138] br[138] wl[6] vdd gnd cell_6t
Xbit_r7_c138 bl[138] br[138] wl[7] vdd gnd cell_6t
Xbit_r8_c138 bl[138] br[138] wl[8] vdd gnd cell_6t
Xbit_r9_c138 bl[138] br[138] wl[9] vdd gnd cell_6t
Xbit_r10_c138 bl[138] br[138] wl[10] vdd gnd cell_6t
Xbit_r11_c138 bl[138] br[138] wl[11] vdd gnd cell_6t
Xbit_r12_c138 bl[138] br[138] wl[12] vdd gnd cell_6t
Xbit_r13_c138 bl[138] br[138] wl[13] vdd gnd cell_6t
Xbit_r14_c138 bl[138] br[138] wl[14] vdd gnd cell_6t
Xbit_r15_c138 bl[138] br[138] wl[15] vdd gnd cell_6t
Xbit_r16_c138 bl[138] br[138] wl[16] vdd gnd cell_6t
Xbit_r17_c138 bl[138] br[138] wl[17] vdd gnd cell_6t
Xbit_r18_c138 bl[138] br[138] wl[18] vdd gnd cell_6t
Xbit_r19_c138 bl[138] br[138] wl[19] vdd gnd cell_6t
Xbit_r20_c138 bl[138] br[138] wl[20] vdd gnd cell_6t
Xbit_r21_c138 bl[138] br[138] wl[21] vdd gnd cell_6t
Xbit_r22_c138 bl[138] br[138] wl[22] vdd gnd cell_6t
Xbit_r23_c138 bl[138] br[138] wl[23] vdd gnd cell_6t
Xbit_r24_c138 bl[138] br[138] wl[24] vdd gnd cell_6t
Xbit_r25_c138 bl[138] br[138] wl[25] vdd gnd cell_6t
Xbit_r26_c138 bl[138] br[138] wl[26] vdd gnd cell_6t
Xbit_r27_c138 bl[138] br[138] wl[27] vdd gnd cell_6t
Xbit_r28_c138 bl[138] br[138] wl[28] vdd gnd cell_6t
Xbit_r29_c138 bl[138] br[138] wl[29] vdd gnd cell_6t
Xbit_r30_c138 bl[138] br[138] wl[30] vdd gnd cell_6t
Xbit_r31_c138 bl[138] br[138] wl[31] vdd gnd cell_6t
Xbit_r32_c138 bl[138] br[138] wl[32] vdd gnd cell_6t
Xbit_r33_c138 bl[138] br[138] wl[33] vdd gnd cell_6t
Xbit_r34_c138 bl[138] br[138] wl[34] vdd gnd cell_6t
Xbit_r35_c138 bl[138] br[138] wl[35] vdd gnd cell_6t
Xbit_r36_c138 bl[138] br[138] wl[36] vdd gnd cell_6t
Xbit_r37_c138 bl[138] br[138] wl[37] vdd gnd cell_6t
Xbit_r38_c138 bl[138] br[138] wl[38] vdd gnd cell_6t
Xbit_r39_c138 bl[138] br[138] wl[39] vdd gnd cell_6t
Xbit_r40_c138 bl[138] br[138] wl[40] vdd gnd cell_6t
Xbit_r41_c138 bl[138] br[138] wl[41] vdd gnd cell_6t
Xbit_r42_c138 bl[138] br[138] wl[42] vdd gnd cell_6t
Xbit_r43_c138 bl[138] br[138] wl[43] vdd gnd cell_6t
Xbit_r44_c138 bl[138] br[138] wl[44] vdd gnd cell_6t
Xbit_r45_c138 bl[138] br[138] wl[45] vdd gnd cell_6t
Xbit_r46_c138 bl[138] br[138] wl[46] vdd gnd cell_6t
Xbit_r47_c138 bl[138] br[138] wl[47] vdd gnd cell_6t
Xbit_r48_c138 bl[138] br[138] wl[48] vdd gnd cell_6t
Xbit_r49_c138 bl[138] br[138] wl[49] vdd gnd cell_6t
Xbit_r50_c138 bl[138] br[138] wl[50] vdd gnd cell_6t
Xbit_r51_c138 bl[138] br[138] wl[51] vdd gnd cell_6t
Xbit_r52_c138 bl[138] br[138] wl[52] vdd gnd cell_6t
Xbit_r53_c138 bl[138] br[138] wl[53] vdd gnd cell_6t
Xbit_r54_c138 bl[138] br[138] wl[54] vdd gnd cell_6t
Xbit_r55_c138 bl[138] br[138] wl[55] vdd gnd cell_6t
Xbit_r56_c138 bl[138] br[138] wl[56] vdd gnd cell_6t
Xbit_r57_c138 bl[138] br[138] wl[57] vdd gnd cell_6t
Xbit_r58_c138 bl[138] br[138] wl[58] vdd gnd cell_6t
Xbit_r59_c138 bl[138] br[138] wl[59] vdd gnd cell_6t
Xbit_r60_c138 bl[138] br[138] wl[60] vdd gnd cell_6t
Xbit_r61_c138 bl[138] br[138] wl[61] vdd gnd cell_6t
Xbit_r62_c138 bl[138] br[138] wl[62] vdd gnd cell_6t
Xbit_r63_c138 bl[138] br[138] wl[63] vdd gnd cell_6t
Xbit_r64_c138 bl[138] br[138] wl[64] vdd gnd cell_6t
Xbit_r65_c138 bl[138] br[138] wl[65] vdd gnd cell_6t
Xbit_r66_c138 bl[138] br[138] wl[66] vdd gnd cell_6t
Xbit_r67_c138 bl[138] br[138] wl[67] vdd gnd cell_6t
Xbit_r68_c138 bl[138] br[138] wl[68] vdd gnd cell_6t
Xbit_r69_c138 bl[138] br[138] wl[69] vdd gnd cell_6t
Xbit_r70_c138 bl[138] br[138] wl[70] vdd gnd cell_6t
Xbit_r71_c138 bl[138] br[138] wl[71] vdd gnd cell_6t
Xbit_r72_c138 bl[138] br[138] wl[72] vdd gnd cell_6t
Xbit_r73_c138 bl[138] br[138] wl[73] vdd gnd cell_6t
Xbit_r74_c138 bl[138] br[138] wl[74] vdd gnd cell_6t
Xbit_r75_c138 bl[138] br[138] wl[75] vdd gnd cell_6t
Xbit_r76_c138 bl[138] br[138] wl[76] vdd gnd cell_6t
Xbit_r77_c138 bl[138] br[138] wl[77] vdd gnd cell_6t
Xbit_r78_c138 bl[138] br[138] wl[78] vdd gnd cell_6t
Xbit_r79_c138 bl[138] br[138] wl[79] vdd gnd cell_6t
Xbit_r80_c138 bl[138] br[138] wl[80] vdd gnd cell_6t
Xbit_r81_c138 bl[138] br[138] wl[81] vdd gnd cell_6t
Xbit_r82_c138 bl[138] br[138] wl[82] vdd gnd cell_6t
Xbit_r83_c138 bl[138] br[138] wl[83] vdd gnd cell_6t
Xbit_r84_c138 bl[138] br[138] wl[84] vdd gnd cell_6t
Xbit_r85_c138 bl[138] br[138] wl[85] vdd gnd cell_6t
Xbit_r86_c138 bl[138] br[138] wl[86] vdd gnd cell_6t
Xbit_r87_c138 bl[138] br[138] wl[87] vdd gnd cell_6t
Xbit_r88_c138 bl[138] br[138] wl[88] vdd gnd cell_6t
Xbit_r89_c138 bl[138] br[138] wl[89] vdd gnd cell_6t
Xbit_r90_c138 bl[138] br[138] wl[90] vdd gnd cell_6t
Xbit_r91_c138 bl[138] br[138] wl[91] vdd gnd cell_6t
Xbit_r92_c138 bl[138] br[138] wl[92] vdd gnd cell_6t
Xbit_r93_c138 bl[138] br[138] wl[93] vdd gnd cell_6t
Xbit_r94_c138 bl[138] br[138] wl[94] vdd gnd cell_6t
Xbit_r95_c138 bl[138] br[138] wl[95] vdd gnd cell_6t
Xbit_r96_c138 bl[138] br[138] wl[96] vdd gnd cell_6t
Xbit_r97_c138 bl[138] br[138] wl[97] vdd gnd cell_6t
Xbit_r98_c138 bl[138] br[138] wl[98] vdd gnd cell_6t
Xbit_r99_c138 bl[138] br[138] wl[99] vdd gnd cell_6t
Xbit_r100_c138 bl[138] br[138] wl[100] vdd gnd cell_6t
Xbit_r101_c138 bl[138] br[138] wl[101] vdd gnd cell_6t
Xbit_r102_c138 bl[138] br[138] wl[102] vdd gnd cell_6t
Xbit_r103_c138 bl[138] br[138] wl[103] vdd gnd cell_6t
Xbit_r104_c138 bl[138] br[138] wl[104] vdd gnd cell_6t
Xbit_r105_c138 bl[138] br[138] wl[105] vdd gnd cell_6t
Xbit_r106_c138 bl[138] br[138] wl[106] vdd gnd cell_6t
Xbit_r107_c138 bl[138] br[138] wl[107] vdd gnd cell_6t
Xbit_r108_c138 bl[138] br[138] wl[108] vdd gnd cell_6t
Xbit_r109_c138 bl[138] br[138] wl[109] vdd gnd cell_6t
Xbit_r110_c138 bl[138] br[138] wl[110] vdd gnd cell_6t
Xbit_r111_c138 bl[138] br[138] wl[111] vdd gnd cell_6t
Xbit_r112_c138 bl[138] br[138] wl[112] vdd gnd cell_6t
Xbit_r113_c138 bl[138] br[138] wl[113] vdd gnd cell_6t
Xbit_r114_c138 bl[138] br[138] wl[114] vdd gnd cell_6t
Xbit_r115_c138 bl[138] br[138] wl[115] vdd gnd cell_6t
Xbit_r116_c138 bl[138] br[138] wl[116] vdd gnd cell_6t
Xbit_r117_c138 bl[138] br[138] wl[117] vdd gnd cell_6t
Xbit_r118_c138 bl[138] br[138] wl[118] vdd gnd cell_6t
Xbit_r119_c138 bl[138] br[138] wl[119] vdd gnd cell_6t
Xbit_r120_c138 bl[138] br[138] wl[120] vdd gnd cell_6t
Xbit_r121_c138 bl[138] br[138] wl[121] vdd gnd cell_6t
Xbit_r122_c138 bl[138] br[138] wl[122] vdd gnd cell_6t
Xbit_r123_c138 bl[138] br[138] wl[123] vdd gnd cell_6t
Xbit_r124_c138 bl[138] br[138] wl[124] vdd gnd cell_6t
Xbit_r125_c138 bl[138] br[138] wl[125] vdd gnd cell_6t
Xbit_r126_c138 bl[138] br[138] wl[126] vdd gnd cell_6t
Xbit_r127_c138 bl[138] br[138] wl[127] vdd gnd cell_6t
Xbit_r0_c139 bl[139] br[139] wl[0] vdd gnd cell_6t
Xbit_r1_c139 bl[139] br[139] wl[1] vdd gnd cell_6t
Xbit_r2_c139 bl[139] br[139] wl[2] vdd gnd cell_6t
Xbit_r3_c139 bl[139] br[139] wl[3] vdd gnd cell_6t
Xbit_r4_c139 bl[139] br[139] wl[4] vdd gnd cell_6t
Xbit_r5_c139 bl[139] br[139] wl[5] vdd gnd cell_6t
Xbit_r6_c139 bl[139] br[139] wl[6] vdd gnd cell_6t
Xbit_r7_c139 bl[139] br[139] wl[7] vdd gnd cell_6t
Xbit_r8_c139 bl[139] br[139] wl[8] vdd gnd cell_6t
Xbit_r9_c139 bl[139] br[139] wl[9] vdd gnd cell_6t
Xbit_r10_c139 bl[139] br[139] wl[10] vdd gnd cell_6t
Xbit_r11_c139 bl[139] br[139] wl[11] vdd gnd cell_6t
Xbit_r12_c139 bl[139] br[139] wl[12] vdd gnd cell_6t
Xbit_r13_c139 bl[139] br[139] wl[13] vdd gnd cell_6t
Xbit_r14_c139 bl[139] br[139] wl[14] vdd gnd cell_6t
Xbit_r15_c139 bl[139] br[139] wl[15] vdd gnd cell_6t
Xbit_r16_c139 bl[139] br[139] wl[16] vdd gnd cell_6t
Xbit_r17_c139 bl[139] br[139] wl[17] vdd gnd cell_6t
Xbit_r18_c139 bl[139] br[139] wl[18] vdd gnd cell_6t
Xbit_r19_c139 bl[139] br[139] wl[19] vdd gnd cell_6t
Xbit_r20_c139 bl[139] br[139] wl[20] vdd gnd cell_6t
Xbit_r21_c139 bl[139] br[139] wl[21] vdd gnd cell_6t
Xbit_r22_c139 bl[139] br[139] wl[22] vdd gnd cell_6t
Xbit_r23_c139 bl[139] br[139] wl[23] vdd gnd cell_6t
Xbit_r24_c139 bl[139] br[139] wl[24] vdd gnd cell_6t
Xbit_r25_c139 bl[139] br[139] wl[25] vdd gnd cell_6t
Xbit_r26_c139 bl[139] br[139] wl[26] vdd gnd cell_6t
Xbit_r27_c139 bl[139] br[139] wl[27] vdd gnd cell_6t
Xbit_r28_c139 bl[139] br[139] wl[28] vdd gnd cell_6t
Xbit_r29_c139 bl[139] br[139] wl[29] vdd gnd cell_6t
Xbit_r30_c139 bl[139] br[139] wl[30] vdd gnd cell_6t
Xbit_r31_c139 bl[139] br[139] wl[31] vdd gnd cell_6t
Xbit_r32_c139 bl[139] br[139] wl[32] vdd gnd cell_6t
Xbit_r33_c139 bl[139] br[139] wl[33] vdd gnd cell_6t
Xbit_r34_c139 bl[139] br[139] wl[34] vdd gnd cell_6t
Xbit_r35_c139 bl[139] br[139] wl[35] vdd gnd cell_6t
Xbit_r36_c139 bl[139] br[139] wl[36] vdd gnd cell_6t
Xbit_r37_c139 bl[139] br[139] wl[37] vdd gnd cell_6t
Xbit_r38_c139 bl[139] br[139] wl[38] vdd gnd cell_6t
Xbit_r39_c139 bl[139] br[139] wl[39] vdd gnd cell_6t
Xbit_r40_c139 bl[139] br[139] wl[40] vdd gnd cell_6t
Xbit_r41_c139 bl[139] br[139] wl[41] vdd gnd cell_6t
Xbit_r42_c139 bl[139] br[139] wl[42] vdd gnd cell_6t
Xbit_r43_c139 bl[139] br[139] wl[43] vdd gnd cell_6t
Xbit_r44_c139 bl[139] br[139] wl[44] vdd gnd cell_6t
Xbit_r45_c139 bl[139] br[139] wl[45] vdd gnd cell_6t
Xbit_r46_c139 bl[139] br[139] wl[46] vdd gnd cell_6t
Xbit_r47_c139 bl[139] br[139] wl[47] vdd gnd cell_6t
Xbit_r48_c139 bl[139] br[139] wl[48] vdd gnd cell_6t
Xbit_r49_c139 bl[139] br[139] wl[49] vdd gnd cell_6t
Xbit_r50_c139 bl[139] br[139] wl[50] vdd gnd cell_6t
Xbit_r51_c139 bl[139] br[139] wl[51] vdd gnd cell_6t
Xbit_r52_c139 bl[139] br[139] wl[52] vdd gnd cell_6t
Xbit_r53_c139 bl[139] br[139] wl[53] vdd gnd cell_6t
Xbit_r54_c139 bl[139] br[139] wl[54] vdd gnd cell_6t
Xbit_r55_c139 bl[139] br[139] wl[55] vdd gnd cell_6t
Xbit_r56_c139 bl[139] br[139] wl[56] vdd gnd cell_6t
Xbit_r57_c139 bl[139] br[139] wl[57] vdd gnd cell_6t
Xbit_r58_c139 bl[139] br[139] wl[58] vdd gnd cell_6t
Xbit_r59_c139 bl[139] br[139] wl[59] vdd gnd cell_6t
Xbit_r60_c139 bl[139] br[139] wl[60] vdd gnd cell_6t
Xbit_r61_c139 bl[139] br[139] wl[61] vdd gnd cell_6t
Xbit_r62_c139 bl[139] br[139] wl[62] vdd gnd cell_6t
Xbit_r63_c139 bl[139] br[139] wl[63] vdd gnd cell_6t
Xbit_r64_c139 bl[139] br[139] wl[64] vdd gnd cell_6t
Xbit_r65_c139 bl[139] br[139] wl[65] vdd gnd cell_6t
Xbit_r66_c139 bl[139] br[139] wl[66] vdd gnd cell_6t
Xbit_r67_c139 bl[139] br[139] wl[67] vdd gnd cell_6t
Xbit_r68_c139 bl[139] br[139] wl[68] vdd gnd cell_6t
Xbit_r69_c139 bl[139] br[139] wl[69] vdd gnd cell_6t
Xbit_r70_c139 bl[139] br[139] wl[70] vdd gnd cell_6t
Xbit_r71_c139 bl[139] br[139] wl[71] vdd gnd cell_6t
Xbit_r72_c139 bl[139] br[139] wl[72] vdd gnd cell_6t
Xbit_r73_c139 bl[139] br[139] wl[73] vdd gnd cell_6t
Xbit_r74_c139 bl[139] br[139] wl[74] vdd gnd cell_6t
Xbit_r75_c139 bl[139] br[139] wl[75] vdd gnd cell_6t
Xbit_r76_c139 bl[139] br[139] wl[76] vdd gnd cell_6t
Xbit_r77_c139 bl[139] br[139] wl[77] vdd gnd cell_6t
Xbit_r78_c139 bl[139] br[139] wl[78] vdd gnd cell_6t
Xbit_r79_c139 bl[139] br[139] wl[79] vdd gnd cell_6t
Xbit_r80_c139 bl[139] br[139] wl[80] vdd gnd cell_6t
Xbit_r81_c139 bl[139] br[139] wl[81] vdd gnd cell_6t
Xbit_r82_c139 bl[139] br[139] wl[82] vdd gnd cell_6t
Xbit_r83_c139 bl[139] br[139] wl[83] vdd gnd cell_6t
Xbit_r84_c139 bl[139] br[139] wl[84] vdd gnd cell_6t
Xbit_r85_c139 bl[139] br[139] wl[85] vdd gnd cell_6t
Xbit_r86_c139 bl[139] br[139] wl[86] vdd gnd cell_6t
Xbit_r87_c139 bl[139] br[139] wl[87] vdd gnd cell_6t
Xbit_r88_c139 bl[139] br[139] wl[88] vdd gnd cell_6t
Xbit_r89_c139 bl[139] br[139] wl[89] vdd gnd cell_6t
Xbit_r90_c139 bl[139] br[139] wl[90] vdd gnd cell_6t
Xbit_r91_c139 bl[139] br[139] wl[91] vdd gnd cell_6t
Xbit_r92_c139 bl[139] br[139] wl[92] vdd gnd cell_6t
Xbit_r93_c139 bl[139] br[139] wl[93] vdd gnd cell_6t
Xbit_r94_c139 bl[139] br[139] wl[94] vdd gnd cell_6t
Xbit_r95_c139 bl[139] br[139] wl[95] vdd gnd cell_6t
Xbit_r96_c139 bl[139] br[139] wl[96] vdd gnd cell_6t
Xbit_r97_c139 bl[139] br[139] wl[97] vdd gnd cell_6t
Xbit_r98_c139 bl[139] br[139] wl[98] vdd gnd cell_6t
Xbit_r99_c139 bl[139] br[139] wl[99] vdd gnd cell_6t
Xbit_r100_c139 bl[139] br[139] wl[100] vdd gnd cell_6t
Xbit_r101_c139 bl[139] br[139] wl[101] vdd gnd cell_6t
Xbit_r102_c139 bl[139] br[139] wl[102] vdd gnd cell_6t
Xbit_r103_c139 bl[139] br[139] wl[103] vdd gnd cell_6t
Xbit_r104_c139 bl[139] br[139] wl[104] vdd gnd cell_6t
Xbit_r105_c139 bl[139] br[139] wl[105] vdd gnd cell_6t
Xbit_r106_c139 bl[139] br[139] wl[106] vdd gnd cell_6t
Xbit_r107_c139 bl[139] br[139] wl[107] vdd gnd cell_6t
Xbit_r108_c139 bl[139] br[139] wl[108] vdd gnd cell_6t
Xbit_r109_c139 bl[139] br[139] wl[109] vdd gnd cell_6t
Xbit_r110_c139 bl[139] br[139] wl[110] vdd gnd cell_6t
Xbit_r111_c139 bl[139] br[139] wl[111] vdd gnd cell_6t
Xbit_r112_c139 bl[139] br[139] wl[112] vdd gnd cell_6t
Xbit_r113_c139 bl[139] br[139] wl[113] vdd gnd cell_6t
Xbit_r114_c139 bl[139] br[139] wl[114] vdd gnd cell_6t
Xbit_r115_c139 bl[139] br[139] wl[115] vdd gnd cell_6t
Xbit_r116_c139 bl[139] br[139] wl[116] vdd gnd cell_6t
Xbit_r117_c139 bl[139] br[139] wl[117] vdd gnd cell_6t
Xbit_r118_c139 bl[139] br[139] wl[118] vdd gnd cell_6t
Xbit_r119_c139 bl[139] br[139] wl[119] vdd gnd cell_6t
Xbit_r120_c139 bl[139] br[139] wl[120] vdd gnd cell_6t
Xbit_r121_c139 bl[139] br[139] wl[121] vdd gnd cell_6t
Xbit_r122_c139 bl[139] br[139] wl[122] vdd gnd cell_6t
Xbit_r123_c139 bl[139] br[139] wl[123] vdd gnd cell_6t
Xbit_r124_c139 bl[139] br[139] wl[124] vdd gnd cell_6t
Xbit_r125_c139 bl[139] br[139] wl[125] vdd gnd cell_6t
Xbit_r126_c139 bl[139] br[139] wl[126] vdd gnd cell_6t
Xbit_r127_c139 bl[139] br[139] wl[127] vdd gnd cell_6t
Xbit_r0_c140 bl[140] br[140] wl[0] vdd gnd cell_6t
Xbit_r1_c140 bl[140] br[140] wl[1] vdd gnd cell_6t
Xbit_r2_c140 bl[140] br[140] wl[2] vdd gnd cell_6t
Xbit_r3_c140 bl[140] br[140] wl[3] vdd gnd cell_6t
Xbit_r4_c140 bl[140] br[140] wl[4] vdd gnd cell_6t
Xbit_r5_c140 bl[140] br[140] wl[5] vdd gnd cell_6t
Xbit_r6_c140 bl[140] br[140] wl[6] vdd gnd cell_6t
Xbit_r7_c140 bl[140] br[140] wl[7] vdd gnd cell_6t
Xbit_r8_c140 bl[140] br[140] wl[8] vdd gnd cell_6t
Xbit_r9_c140 bl[140] br[140] wl[9] vdd gnd cell_6t
Xbit_r10_c140 bl[140] br[140] wl[10] vdd gnd cell_6t
Xbit_r11_c140 bl[140] br[140] wl[11] vdd gnd cell_6t
Xbit_r12_c140 bl[140] br[140] wl[12] vdd gnd cell_6t
Xbit_r13_c140 bl[140] br[140] wl[13] vdd gnd cell_6t
Xbit_r14_c140 bl[140] br[140] wl[14] vdd gnd cell_6t
Xbit_r15_c140 bl[140] br[140] wl[15] vdd gnd cell_6t
Xbit_r16_c140 bl[140] br[140] wl[16] vdd gnd cell_6t
Xbit_r17_c140 bl[140] br[140] wl[17] vdd gnd cell_6t
Xbit_r18_c140 bl[140] br[140] wl[18] vdd gnd cell_6t
Xbit_r19_c140 bl[140] br[140] wl[19] vdd gnd cell_6t
Xbit_r20_c140 bl[140] br[140] wl[20] vdd gnd cell_6t
Xbit_r21_c140 bl[140] br[140] wl[21] vdd gnd cell_6t
Xbit_r22_c140 bl[140] br[140] wl[22] vdd gnd cell_6t
Xbit_r23_c140 bl[140] br[140] wl[23] vdd gnd cell_6t
Xbit_r24_c140 bl[140] br[140] wl[24] vdd gnd cell_6t
Xbit_r25_c140 bl[140] br[140] wl[25] vdd gnd cell_6t
Xbit_r26_c140 bl[140] br[140] wl[26] vdd gnd cell_6t
Xbit_r27_c140 bl[140] br[140] wl[27] vdd gnd cell_6t
Xbit_r28_c140 bl[140] br[140] wl[28] vdd gnd cell_6t
Xbit_r29_c140 bl[140] br[140] wl[29] vdd gnd cell_6t
Xbit_r30_c140 bl[140] br[140] wl[30] vdd gnd cell_6t
Xbit_r31_c140 bl[140] br[140] wl[31] vdd gnd cell_6t
Xbit_r32_c140 bl[140] br[140] wl[32] vdd gnd cell_6t
Xbit_r33_c140 bl[140] br[140] wl[33] vdd gnd cell_6t
Xbit_r34_c140 bl[140] br[140] wl[34] vdd gnd cell_6t
Xbit_r35_c140 bl[140] br[140] wl[35] vdd gnd cell_6t
Xbit_r36_c140 bl[140] br[140] wl[36] vdd gnd cell_6t
Xbit_r37_c140 bl[140] br[140] wl[37] vdd gnd cell_6t
Xbit_r38_c140 bl[140] br[140] wl[38] vdd gnd cell_6t
Xbit_r39_c140 bl[140] br[140] wl[39] vdd gnd cell_6t
Xbit_r40_c140 bl[140] br[140] wl[40] vdd gnd cell_6t
Xbit_r41_c140 bl[140] br[140] wl[41] vdd gnd cell_6t
Xbit_r42_c140 bl[140] br[140] wl[42] vdd gnd cell_6t
Xbit_r43_c140 bl[140] br[140] wl[43] vdd gnd cell_6t
Xbit_r44_c140 bl[140] br[140] wl[44] vdd gnd cell_6t
Xbit_r45_c140 bl[140] br[140] wl[45] vdd gnd cell_6t
Xbit_r46_c140 bl[140] br[140] wl[46] vdd gnd cell_6t
Xbit_r47_c140 bl[140] br[140] wl[47] vdd gnd cell_6t
Xbit_r48_c140 bl[140] br[140] wl[48] vdd gnd cell_6t
Xbit_r49_c140 bl[140] br[140] wl[49] vdd gnd cell_6t
Xbit_r50_c140 bl[140] br[140] wl[50] vdd gnd cell_6t
Xbit_r51_c140 bl[140] br[140] wl[51] vdd gnd cell_6t
Xbit_r52_c140 bl[140] br[140] wl[52] vdd gnd cell_6t
Xbit_r53_c140 bl[140] br[140] wl[53] vdd gnd cell_6t
Xbit_r54_c140 bl[140] br[140] wl[54] vdd gnd cell_6t
Xbit_r55_c140 bl[140] br[140] wl[55] vdd gnd cell_6t
Xbit_r56_c140 bl[140] br[140] wl[56] vdd gnd cell_6t
Xbit_r57_c140 bl[140] br[140] wl[57] vdd gnd cell_6t
Xbit_r58_c140 bl[140] br[140] wl[58] vdd gnd cell_6t
Xbit_r59_c140 bl[140] br[140] wl[59] vdd gnd cell_6t
Xbit_r60_c140 bl[140] br[140] wl[60] vdd gnd cell_6t
Xbit_r61_c140 bl[140] br[140] wl[61] vdd gnd cell_6t
Xbit_r62_c140 bl[140] br[140] wl[62] vdd gnd cell_6t
Xbit_r63_c140 bl[140] br[140] wl[63] vdd gnd cell_6t
Xbit_r64_c140 bl[140] br[140] wl[64] vdd gnd cell_6t
Xbit_r65_c140 bl[140] br[140] wl[65] vdd gnd cell_6t
Xbit_r66_c140 bl[140] br[140] wl[66] vdd gnd cell_6t
Xbit_r67_c140 bl[140] br[140] wl[67] vdd gnd cell_6t
Xbit_r68_c140 bl[140] br[140] wl[68] vdd gnd cell_6t
Xbit_r69_c140 bl[140] br[140] wl[69] vdd gnd cell_6t
Xbit_r70_c140 bl[140] br[140] wl[70] vdd gnd cell_6t
Xbit_r71_c140 bl[140] br[140] wl[71] vdd gnd cell_6t
Xbit_r72_c140 bl[140] br[140] wl[72] vdd gnd cell_6t
Xbit_r73_c140 bl[140] br[140] wl[73] vdd gnd cell_6t
Xbit_r74_c140 bl[140] br[140] wl[74] vdd gnd cell_6t
Xbit_r75_c140 bl[140] br[140] wl[75] vdd gnd cell_6t
Xbit_r76_c140 bl[140] br[140] wl[76] vdd gnd cell_6t
Xbit_r77_c140 bl[140] br[140] wl[77] vdd gnd cell_6t
Xbit_r78_c140 bl[140] br[140] wl[78] vdd gnd cell_6t
Xbit_r79_c140 bl[140] br[140] wl[79] vdd gnd cell_6t
Xbit_r80_c140 bl[140] br[140] wl[80] vdd gnd cell_6t
Xbit_r81_c140 bl[140] br[140] wl[81] vdd gnd cell_6t
Xbit_r82_c140 bl[140] br[140] wl[82] vdd gnd cell_6t
Xbit_r83_c140 bl[140] br[140] wl[83] vdd gnd cell_6t
Xbit_r84_c140 bl[140] br[140] wl[84] vdd gnd cell_6t
Xbit_r85_c140 bl[140] br[140] wl[85] vdd gnd cell_6t
Xbit_r86_c140 bl[140] br[140] wl[86] vdd gnd cell_6t
Xbit_r87_c140 bl[140] br[140] wl[87] vdd gnd cell_6t
Xbit_r88_c140 bl[140] br[140] wl[88] vdd gnd cell_6t
Xbit_r89_c140 bl[140] br[140] wl[89] vdd gnd cell_6t
Xbit_r90_c140 bl[140] br[140] wl[90] vdd gnd cell_6t
Xbit_r91_c140 bl[140] br[140] wl[91] vdd gnd cell_6t
Xbit_r92_c140 bl[140] br[140] wl[92] vdd gnd cell_6t
Xbit_r93_c140 bl[140] br[140] wl[93] vdd gnd cell_6t
Xbit_r94_c140 bl[140] br[140] wl[94] vdd gnd cell_6t
Xbit_r95_c140 bl[140] br[140] wl[95] vdd gnd cell_6t
Xbit_r96_c140 bl[140] br[140] wl[96] vdd gnd cell_6t
Xbit_r97_c140 bl[140] br[140] wl[97] vdd gnd cell_6t
Xbit_r98_c140 bl[140] br[140] wl[98] vdd gnd cell_6t
Xbit_r99_c140 bl[140] br[140] wl[99] vdd gnd cell_6t
Xbit_r100_c140 bl[140] br[140] wl[100] vdd gnd cell_6t
Xbit_r101_c140 bl[140] br[140] wl[101] vdd gnd cell_6t
Xbit_r102_c140 bl[140] br[140] wl[102] vdd gnd cell_6t
Xbit_r103_c140 bl[140] br[140] wl[103] vdd gnd cell_6t
Xbit_r104_c140 bl[140] br[140] wl[104] vdd gnd cell_6t
Xbit_r105_c140 bl[140] br[140] wl[105] vdd gnd cell_6t
Xbit_r106_c140 bl[140] br[140] wl[106] vdd gnd cell_6t
Xbit_r107_c140 bl[140] br[140] wl[107] vdd gnd cell_6t
Xbit_r108_c140 bl[140] br[140] wl[108] vdd gnd cell_6t
Xbit_r109_c140 bl[140] br[140] wl[109] vdd gnd cell_6t
Xbit_r110_c140 bl[140] br[140] wl[110] vdd gnd cell_6t
Xbit_r111_c140 bl[140] br[140] wl[111] vdd gnd cell_6t
Xbit_r112_c140 bl[140] br[140] wl[112] vdd gnd cell_6t
Xbit_r113_c140 bl[140] br[140] wl[113] vdd gnd cell_6t
Xbit_r114_c140 bl[140] br[140] wl[114] vdd gnd cell_6t
Xbit_r115_c140 bl[140] br[140] wl[115] vdd gnd cell_6t
Xbit_r116_c140 bl[140] br[140] wl[116] vdd gnd cell_6t
Xbit_r117_c140 bl[140] br[140] wl[117] vdd gnd cell_6t
Xbit_r118_c140 bl[140] br[140] wl[118] vdd gnd cell_6t
Xbit_r119_c140 bl[140] br[140] wl[119] vdd gnd cell_6t
Xbit_r120_c140 bl[140] br[140] wl[120] vdd gnd cell_6t
Xbit_r121_c140 bl[140] br[140] wl[121] vdd gnd cell_6t
Xbit_r122_c140 bl[140] br[140] wl[122] vdd gnd cell_6t
Xbit_r123_c140 bl[140] br[140] wl[123] vdd gnd cell_6t
Xbit_r124_c140 bl[140] br[140] wl[124] vdd gnd cell_6t
Xbit_r125_c140 bl[140] br[140] wl[125] vdd gnd cell_6t
Xbit_r126_c140 bl[140] br[140] wl[126] vdd gnd cell_6t
Xbit_r127_c140 bl[140] br[140] wl[127] vdd gnd cell_6t
Xbit_r0_c141 bl[141] br[141] wl[0] vdd gnd cell_6t
Xbit_r1_c141 bl[141] br[141] wl[1] vdd gnd cell_6t
Xbit_r2_c141 bl[141] br[141] wl[2] vdd gnd cell_6t
Xbit_r3_c141 bl[141] br[141] wl[3] vdd gnd cell_6t
Xbit_r4_c141 bl[141] br[141] wl[4] vdd gnd cell_6t
Xbit_r5_c141 bl[141] br[141] wl[5] vdd gnd cell_6t
Xbit_r6_c141 bl[141] br[141] wl[6] vdd gnd cell_6t
Xbit_r7_c141 bl[141] br[141] wl[7] vdd gnd cell_6t
Xbit_r8_c141 bl[141] br[141] wl[8] vdd gnd cell_6t
Xbit_r9_c141 bl[141] br[141] wl[9] vdd gnd cell_6t
Xbit_r10_c141 bl[141] br[141] wl[10] vdd gnd cell_6t
Xbit_r11_c141 bl[141] br[141] wl[11] vdd gnd cell_6t
Xbit_r12_c141 bl[141] br[141] wl[12] vdd gnd cell_6t
Xbit_r13_c141 bl[141] br[141] wl[13] vdd gnd cell_6t
Xbit_r14_c141 bl[141] br[141] wl[14] vdd gnd cell_6t
Xbit_r15_c141 bl[141] br[141] wl[15] vdd gnd cell_6t
Xbit_r16_c141 bl[141] br[141] wl[16] vdd gnd cell_6t
Xbit_r17_c141 bl[141] br[141] wl[17] vdd gnd cell_6t
Xbit_r18_c141 bl[141] br[141] wl[18] vdd gnd cell_6t
Xbit_r19_c141 bl[141] br[141] wl[19] vdd gnd cell_6t
Xbit_r20_c141 bl[141] br[141] wl[20] vdd gnd cell_6t
Xbit_r21_c141 bl[141] br[141] wl[21] vdd gnd cell_6t
Xbit_r22_c141 bl[141] br[141] wl[22] vdd gnd cell_6t
Xbit_r23_c141 bl[141] br[141] wl[23] vdd gnd cell_6t
Xbit_r24_c141 bl[141] br[141] wl[24] vdd gnd cell_6t
Xbit_r25_c141 bl[141] br[141] wl[25] vdd gnd cell_6t
Xbit_r26_c141 bl[141] br[141] wl[26] vdd gnd cell_6t
Xbit_r27_c141 bl[141] br[141] wl[27] vdd gnd cell_6t
Xbit_r28_c141 bl[141] br[141] wl[28] vdd gnd cell_6t
Xbit_r29_c141 bl[141] br[141] wl[29] vdd gnd cell_6t
Xbit_r30_c141 bl[141] br[141] wl[30] vdd gnd cell_6t
Xbit_r31_c141 bl[141] br[141] wl[31] vdd gnd cell_6t
Xbit_r32_c141 bl[141] br[141] wl[32] vdd gnd cell_6t
Xbit_r33_c141 bl[141] br[141] wl[33] vdd gnd cell_6t
Xbit_r34_c141 bl[141] br[141] wl[34] vdd gnd cell_6t
Xbit_r35_c141 bl[141] br[141] wl[35] vdd gnd cell_6t
Xbit_r36_c141 bl[141] br[141] wl[36] vdd gnd cell_6t
Xbit_r37_c141 bl[141] br[141] wl[37] vdd gnd cell_6t
Xbit_r38_c141 bl[141] br[141] wl[38] vdd gnd cell_6t
Xbit_r39_c141 bl[141] br[141] wl[39] vdd gnd cell_6t
Xbit_r40_c141 bl[141] br[141] wl[40] vdd gnd cell_6t
Xbit_r41_c141 bl[141] br[141] wl[41] vdd gnd cell_6t
Xbit_r42_c141 bl[141] br[141] wl[42] vdd gnd cell_6t
Xbit_r43_c141 bl[141] br[141] wl[43] vdd gnd cell_6t
Xbit_r44_c141 bl[141] br[141] wl[44] vdd gnd cell_6t
Xbit_r45_c141 bl[141] br[141] wl[45] vdd gnd cell_6t
Xbit_r46_c141 bl[141] br[141] wl[46] vdd gnd cell_6t
Xbit_r47_c141 bl[141] br[141] wl[47] vdd gnd cell_6t
Xbit_r48_c141 bl[141] br[141] wl[48] vdd gnd cell_6t
Xbit_r49_c141 bl[141] br[141] wl[49] vdd gnd cell_6t
Xbit_r50_c141 bl[141] br[141] wl[50] vdd gnd cell_6t
Xbit_r51_c141 bl[141] br[141] wl[51] vdd gnd cell_6t
Xbit_r52_c141 bl[141] br[141] wl[52] vdd gnd cell_6t
Xbit_r53_c141 bl[141] br[141] wl[53] vdd gnd cell_6t
Xbit_r54_c141 bl[141] br[141] wl[54] vdd gnd cell_6t
Xbit_r55_c141 bl[141] br[141] wl[55] vdd gnd cell_6t
Xbit_r56_c141 bl[141] br[141] wl[56] vdd gnd cell_6t
Xbit_r57_c141 bl[141] br[141] wl[57] vdd gnd cell_6t
Xbit_r58_c141 bl[141] br[141] wl[58] vdd gnd cell_6t
Xbit_r59_c141 bl[141] br[141] wl[59] vdd gnd cell_6t
Xbit_r60_c141 bl[141] br[141] wl[60] vdd gnd cell_6t
Xbit_r61_c141 bl[141] br[141] wl[61] vdd gnd cell_6t
Xbit_r62_c141 bl[141] br[141] wl[62] vdd gnd cell_6t
Xbit_r63_c141 bl[141] br[141] wl[63] vdd gnd cell_6t
Xbit_r64_c141 bl[141] br[141] wl[64] vdd gnd cell_6t
Xbit_r65_c141 bl[141] br[141] wl[65] vdd gnd cell_6t
Xbit_r66_c141 bl[141] br[141] wl[66] vdd gnd cell_6t
Xbit_r67_c141 bl[141] br[141] wl[67] vdd gnd cell_6t
Xbit_r68_c141 bl[141] br[141] wl[68] vdd gnd cell_6t
Xbit_r69_c141 bl[141] br[141] wl[69] vdd gnd cell_6t
Xbit_r70_c141 bl[141] br[141] wl[70] vdd gnd cell_6t
Xbit_r71_c141 bl[141] br[141] wl[71] vdd gnd cell_6t
Xbit_r72_c141 bl[141] br[141] wl[72] vdd gnd cell_6t
Xbit_r73_c141 bl[141] br[141] wl[73] vdd gnd cell_6t
Xbit_r74_c141 bl[141] br[141] wl[74] vdd gnd cell_6t
Xbit_r75_c141 bl[141] br[141] wl[75] vdd gnd cell_6t
Xbit_r76_c141 bl[141] br[141] wl[76] vdd gnd cell_6t
Xbit_r77_c141 bl[141] br[141] wl[77] vdd gnd cell_6t
Xbit_r78_c141 bl[141] br[141] wl[78] vdd gnd cell_6t
Xbit_r79_c141 bl[141] br[141] wl[79] vdd gnd cell_6t
Xbit_r80_c141 bl[141] br[141] wl[80] vdd gnd cell_6t
Xbit_r81_c141 bl[141] br[141] wl[81] vdd gnd cell_6t
Xbit_r82_c141 bl[141] br[141] wl[82] vdd gnd cell_6t
Xbit_r83_c141 bl[141] br[141] wl[83] vdd gnd cell_6t
Xbit_r84_c141 bl[141] br[141] wl[84] vdd gnd cell_6t
Xbit_r85_c141 bl[141] br[141] wl[85] vdd gnd cell_6t
Xbit_r86_c141 bl[141] br[141] wl[86] vdd gnd cell_6t
Xbit_r87_c141 bl[141] br[141] wl[87] vdd gnd cell_6t
Xbit_r88_c141 bl[141] br[141] wl[88] vdd gnd cell_6t
Xbit_r89_c141 bl[141] br[141] wl[89] vdd gnd cell_6t
Xbit_r90_c141 bl[141] br[141] wl[90] vdd gnd cell_6t
Xbit_r91_c141 bl[141] br[141] wl[91] vdd gnd cell_6t
Xbit_r92_c141 bl[141] br[141] wl[92] vdd gnd cell_6t
Xbit_r93_c141 bl[141] br[141] wl[93] vdd gnd cell_6t
Xbit_r94_c141 bl[141] br[141] wl[94] vdd gnd cell_6t
Xbit_r95_c141 bl[141] br[141] wl[95] vdd gnd cell_6t
Xbit_r96_c141 bl[141] br[141] wl[96] vdd gnd cell_6t
Xbit_r97_c141 bl[141] br[141] wl[97] vdd gnd cell_6t
Xbit_r98_c141 bl[141] br[141] wl[98] vdd gnd cell_6t
Xbit_r99_c141 bl[141] br[141] wl[99] vdd gnd cell_6t
Xbit_r100_c141 bl[141] br[141] wl[100] vdd gnd cell_6t
Xbit_r101_c141 bl[141] br[141] wl[101] vdd gnd cell_6t
Xbit_r102_c141 bl[141] br[141] wl[102] vdd gnd cell_6t
Xbit_r103_c141 bl[141] br[141] wl[103] vdd gnd cell_6t
Xbit_r104_c141 bl[141] br[141] wl[104] vdd gnd cell_6t
Xbit_r105_c141 bl[141] br[141] wl[105] vdd gnd cell_6t
Xbit_r106_c141 bl[141] br[141] wl[106] vdd gnd cell_6t
Xbit_r107_c141 bl[141] br[141] wl[107] vdd gnd cell_6t
Xbit_r108_c141 bl[141] br[141] wl[108] vdd gnd cell_6t
Xbit_r109_c141 bl[141] br[141] wl[109] vdd gnd cell_6t
Xbit_r110_c141 bl[141] br[141] wl[110] vdd gnd cell_6t
Xbit_r111_c141 bl[141] br[141] wl[111] vdd gnd cell_6t
Xbit_r112_c141 bl[141] br[141] wl[112] vdd gnd cell_6t
Xbit_r113_c141 bl[141] br[141] wl[113] vdd gnd cell_6t
Xbit_r114_c141 bl[141] br[141] wl[114] vdd gnd cell_6t
Xbit_r115_c141 bl[141] br[141] wl[115] vdd gnd cell_6t
Xbit_r116_c141 bl[141] br[141] wl[116] vdd gnd cell_6t
Xbit_r117_c141 bl[141] br[141] wl[117] vdd gnd cell_6t
Xbit_r118_c141 bl[141] br[141] wl[118] vdd gnd cell_6t
Xbit_r119_c141 bl[141] br[141] wl[119] vdd gnd cell_6t
Xbit_r120_c141 bl[141] br[141] wl[120] vdd gnd cell_6t
Xbit_r121_c141 bl[141] br[141] wl[121] vdd gnd cell_6t
Xbit_r122_c141 bl[141] br[141] wl[122] vdd gnd cell_6t
Xbit_r123_c141 bl[141] br[141] wl[123] vdd gnd cell_6t
Xbit_r124_c141 bl[141] br[141] wl[124] vdd gnd cell_6t
Xbit_r125_c141 bl[141] br[141] wl[125] vdd gnd cell_6t
Xbit_r126_c141 bl[141] br[141] wl[126] vdd gnd cell_6t
Xbit_r127_c141 bl[141] br[141] wl[127] vdd gnd cell_6t
Xbit_r0_c142 bl[142] br[142] wl[0] vdd gnd cell_6t
Xbit_r1_c142 bl[142] br[142] wl[1] vdd gnd cell_6t
Xbit_r2_c142 bl[142] br[142] wl[2] vdd gnd cell_6t
Xbit_r3_c142 bl[142] br[142] wl[3] vdd gnd cell_6t
Xbit_r4_c142 bl[142] br[142] wl[4] vdd gnd cell_6t
Xbit_r5_c142 bl[142] br[142] wl[5] vdd gnd cell_6t
Xbit_r6_c142 bl[142] br[142] wl[6] vdd gnd cell_6t
Xbit_r7_c142 bl[142] br[142] wl[7] vdd gnd cell_6t
Xbit_r8_c142 bl[142] br[142] wl[8] vdd gnd cell_6t
Xbit_r9_c142 bl[142] br[142] wl[9] vdd gnd cell_6t
Xbit_r10_c142 bl[142] br[142] wl[10] vdd gnd cell_6t
Xbit_r11_c142 bl[142] br[142] wl[11] vdd gnd cell_6t
Xbit_r12_c142 bl[142] br[142] wl[12] vdd gnd cell_6t
Xbit_r13_c142 bl[142] br[142] wl[13] vdd gnd cell_6t
Xbit_r14_c142 bl[142] br[142] wl[14] vdd gnd cell_6t
Xbit_r15_c142 bl[142] br[142] wl[15] vdd gnd cell_6t
Xbit_r16_c142 bl[142] br[142] wl[16] vdd gnd cell_6t
Xbit_r17_c142 bl[142] br[142] wl[17] vdd gnd cell_6t
Xbit_r18_c142 bl[142] br[142] wl[18] vdd gnd cell_6t
Xbit_r19_c142 bl[142] br[142] wl[19] vdd gnd cell_6t
Xbit_r20_c142 bl[142] br[142] wl[20] vdd gnd cell_6t
Xbit_r21_c142 bl[142] br[142] wl[21] vdd gnd cell_6t
Xbit_r22_c142 bl[142] br[142] wl[22] vdd gnd cell_6t
Xbit_r23_c142 bl[142] br[142] wl[23] vdd gnd cell_6t
Xbit_r24_c142 bl[142] br[142] wl[24] vdd gnd cell_6t
Xbit_r25_c142 bl[142] br[142] wl[25] vdd gnd cell_6t
Xbit_r26_c142 bl[142] br[142] wl[26] vdd gnd cell_6t
Xbit_r27_c142 bl[142] br[142] wl[27] vdd gnd cell_6t
Xbit_r28_c142 bl[142] br[142] wl[28] vdd gnd cell_6t
Xbit_r29_c142 bl[142] br[142] wl[29] vdd gnd cell_6t
Xbit_r30_c142 bl[142] br[142] wl[30] vdd gnd cell_6t
Xbit_r31_c142 bl[142] br[142] wl[31] vdd gnd cell_6t
Xbit_r32_c142 bl[142] br[142] wl[32] vdd gnd cell_6t
Xbit_r33_c142 bl[142] br[142] wl[33] vdd gnd cell_6t
Xbit_r34_c142 bl[142] br[142] wl[34] vdd gnd cell_6t
Xbit_r35_c142 bl[142] br[142] wl[35] vdd gnd cell_6t
Xbit_r36_c142 bl[142] br[142] wl[36] vdd gnd cell_6t
Xbit_r37_c142 bl[142] br[142] wl[37] vdd gnd cell_6t
Xbit_r38_c142 bl[142] br[142] wl[38] vdd gnd cell_6t
Xbit_r39_c142 bl[142] br[142] wl[39] vdd gnd cell_6t
Xbit_r40_c142 bl[142] br[142] wl[40] vdd gnd cell_6t
Xbit_r41_c142 bl[142] br[142] wl[41] vdd gnd cell_6t
Xbit_r42_c142 bl[142] br[142] wl[42] vdd gnd cell_6t
Xbit_r43_c142 bl[142] br[142] wl[43] vdd gnd cell_6t
Xbit_r44_c142 bl[142] br[142] wl[44] vdd gnd cell_6t
Xbit_r45_c142 bl[142] br[142] wl[45] vdd gnd cell_6t
Xbit_r46_c142 bl[142] br[142] wl[46] vdd gnd cell_6t
Xbit_r47_c142 bl[142] br[142] wl[47] vdd gnd cell_6t
Xbit_r48_c142 bl[142] br[142] wl[48] vdd gnd cell_6t
Xbit_r49_c142 bl[142] br[142] wl[49] vdd gnd cell_6t
Xbit_r50_c142 bl[142] br[142] wl[50] vdd gnd cell_6t
Xbit_r51_c142 bl[142] br[142] wl[51] vdd gnd cell_6t
Xbit_r52_c142 bl[142] br[142] wl[52] vdd gnd cell_6t
Xbit_r53_c142 bl[142] br[142] wl[53] vdd gnd cell_6t
Xbit_r54_c142 bl[142] br[142] wl[54] vdd gnd cell_6t
Xbit_r55_c142 bl[142] br[142] wl[55] vdd gnd cell_6t
Xbit_r56_c142 bl[142] br[142] wl[56] vdd gnd cell_6t
Xbit_r57_c142 bl[142] br[142] wl[57] vdd gnd cell_6t
Xbit_r58_c142 bl[142] br[142] wl[58] vdd gnd cell_6t
Xbit_r59_c142 bl[142] br[142] wl[59] vdd gnd cell_6t
Xbit_r60_c142 bl[142] br[142] wl[60] vdd gnd cell_6t
Xbit_r61_c142 bl[142] br[142] wl[61] vdd gnd cell_6t
Xbit_r62_c142 bl[142] br[142] wl[62] vdd gnd cell_6t
Xbit_r63_c142 bl[142] br[142] wl[63] vdd gnd cell_6t
Xbit_r64_c142 bl[142] br[142] wl[64] vdd gnd cell_6t
Xbit_r65_c142 bl[142] br[142] wl[65] vdd gnd cell_6t
Xbit_r66_c142 bl[142] br[142] wl[66] vdd gnd cell_6t
Xbit_r67_c142 bl[142] br[142] wl[67] vdd gnd cell_6t
Xbit_r68_c142 bl[142] br[142] wl[68] vdd gnd cell_6t
Xbit_r69_c142 bl[142] br[142] wl[69] vdd gnd cell_6t
Xbit_r70_c142 bl[142] br[142] wl[70] vdd gnd cell_6t
Xbit_r71_c142 bl[142] br[142] wl[71] vdd gnd cell_6t
Xbit_r72_c142 bl[142] br[142] wl[72] vdd gnd cell_6t
Xbit_r73_c142 bl[142] br[142] wl[73] vdd gnd cell_6t
Xbit_r74_c142 bl[142] br[142] wl[74] vdd gnd cell_6t
Xbit_r75_c142 bl[142] br[142] wl[75] vdd gnd cell_6t
Xbit_r76_c142 bl[142] br[142] wl[76] vdd gnd cell_6t
Xbit_r77_c142 bl[142] br[142] wl[77] vdd gnd cell_6t
Xbit_r78_c142 bl[142] br[142] wl[78] vdd gnd cell_6t
Xbit_r79_c142 bl[142] br[142] wl[79] vdd gnd cell_6t
Xbit_r80_c142 bl[142] br[142] wl[80] vdd gnd cell_6t
Xbit_r81_c142 bl[142] br[142] wl[81] vdd gnd cell_6t
Xbit_r82_c142 bl[142] br[142] wl[82] vdd gnd cell_6t
Xbit_r83_c142 bl[142] br[142] wl[83] vdd gnd cell_6t
Xbit_r84_c142 bl[142] br[142] wl[84] vdd gnd cell_6t
Xbit_r85_c142 bl[142] br[142] wl[85] vdd gnd cell_6t
Xbit_r86_c142 bl[142] br[142] wl[86] vdd gnd cell_6t
Xbit_r87_c142 bl[142] br[142] wl[87] vdd gnd cell_6t
Xbit_r88_c142 bl[142] br[142] wl[88] vdd gnd cell_6t
Xbit_r89_c142 bl[142] br[142] wl[89] vdd gnd cell_6t
Xbit_r90_c142 bl[142] br[142] wl[90] vdd gnd cell_6t
Xbit_r91_c142 bl[142] br[142] wl[91] vdd gnd cell_6t
Xbit_r92_c142 bl[142] br[142] wl[92] vdd gnd cell_6t
Xbit_r93_c142 bl[142] br[142] wl[93] vdd gnd cell_6t
Xbit_r94_c142 bl[142] br[142] wl[94] vdd gnd cell_6t
Xbit_r95_c142 bl[142] br[142] wl[95] vdd gnd cell_6t
Xbit_r96_c142 bl[142] br[142] wl[96] vdd gnd cell_6t
Xbit_r97_c142 bl[142] br[142] wl[97] vdd gnd cell_6t
Xbit_r98_c142 bl[142] br[142] wl[98] vdd gnd cell_6t
Xbit_r99_c142 bl[142] br[142] wl[99] vdd gnd cell_6t
Xbit_r100_c142 bl[142] br[142] wl[100] vdd gnd cell_6t
Xbit_r101_c142 bl[142] br[142] wl[101] vdd gnd cell_6t
Xbit_r102_c142 bl[142] br[142] wl[102] vdd gnd cell_6t
Xbit_r103_c142 bl[142] br[142] wl[103] vdd gnd cell_6t
Xbit_r104_c142 bl[142] br[142] wl[104] vdd gnd cell_6t
Xbit_r105_c142 bl[142] br[142] wl[105] vdd gnd cell_6t
Xbit_r106_c142 bl[142] br[142] wl[106] vdd gnd cell_6t
Xbit_r107_c142 bl[142] br[142] wl[107] vdd gnd cell_6t
Xbit_r108_c142 bl[142] br[142] wl[108] vdd gnd cell_6t
Xbit_r109_c142 bl[142] br[142] wl[109] vdd gnd cell_6t
Xbit_r110_c142 bl[142] br[142] wl[110] vdd gnd cell_6t
Xbit_r111_c142 bl[142] br[142] wl[111] vdd gnd cell_6t
Xbit_r112_c142 bl[142] br[142] wl[112] vdd gnd cell_6t
Xbit_r113_c142 bl[142] br[142] wl[113] vdd gnd cell_6t
Xbit_r114_c142 bl[142] br[142] wl[114] vdd gnd cell_6t
Xbit_r115_c142 bl[142] br[142] wl[115] vdd gnd cell_6t
Xbit_r116_c142 bl[142] br[142] wl[116] vdd gnd cell_6t
Xbit_r117_c142 bl[142] br[142] wl[117] vdd gnd cell_6t
Xbit_r118_c142 bl[142] br[142] wl[118] vdd gnd cell_6t
Xbit_r119_c142 bl[142] br[142] wl[119] vdd gnd cell_6t
Xbit_r120_c142 bl[142] br[142] wl[120] vdd gnd cell_6t
Xbit_r121_c142 bl[142] br[142] wl[121] vdd gnd cell_6t
Xbit_r122_c142 bl[142] br[142] wl[122] vdd gnd cell_6t
Xbit_r123_c142 bl[142] br[142] wl[123] vdd gnd cell_6t
Xbit_r124_c142 bl[142] br[142] wl[124] vdd gnd cell_6t
Xbit_r125_c142 bl[142] br[142] wl[125] vdd gnd cell_6t
Xbit_r126_c142 bl[142] br[142] wl[126] vdd gnd cell_6t
Xbit_r127_c142 bl[142] br[142] wl[127] vdd gnd cell_6t
Xbit_r0_c143 bl[143] br[143] wl[0] vdd gnd cell_6t
Xbit_r1_c143 bl[143] br[143] wl[1] vdd gnd cell_6t
Xbit_r2_c143 bl[143] br[143] wl[2] vdd gnd cell_6t
Xbit_r3_c143 bl[143] br[143] wl[3] vdd gnd cell_6t
Xbit_r4_c143 bl[143] br[143] wl[4] vdd gnd cell_6t
Xbit_r5_c143 bl[143] br[143] wl[5] vdd gnd cell_6t
Xbit_r6_c143 bl[143] br[143] wl[6] vdd gnd cell_6t
Xbit_r7_c143 bl[143] br[143] wl[7] vdd gnd cell_6t
Xbit_r8_c143 bl[143] br[143] wl[8] vdd gnd cell_6t
Xbit_r9_c143 bl[143] br[143] wl[9] vdd gnd cell_6t
Xbit_r10_c143 bl[143] br[143] wl[10] vdd gnd cell_6t
Xbit_r11_c143 bl[143] br[143] wl[11] vdd gnd cell_6t
Xbit_r12_c143 bl[143] br[143] wl[12] vdd gnd cell_6t
Xbit_r13_c143 bl[143] br[143] wl[13] vdd gnd cell_6t
Xbit_r14_c143 bl[143] br[143] wl[14] vdd gnd cell_6t
Xbit_r15_c143 bl[143] br[143] wl[15] vdd gnd cell_6t
Xbit_r16_c143 bl[143] br[143] wl[16] vdd gnd cell_6t
Xbit_r17_c143 bl[143] br[143] wl[17] vdd gnd cell_6t
Xbit_r18_c143 bl[143] br[143] wl[18] vdd gnd cell_6t
Xbit_r19_c143 bl[143] br[143] wl[19] vdd gnd cell_6t
Xbit_r20_c143 bl[143] br[143] wl[20] vdd gnd cell_6t
Xbit_r21_c143 bl[143] br[143] wl[21] vdd gnd cell_6t
Xbit_r22_c143 bl[143] br[143] wl[22] vdd gnd cell_6t
Xbit_r23_c143 bl[143] br[143] wl[23] vdd gnd cell_6t
Xbit_r24_c143 bl[143] br[143] wl[24] vdd gnd cell_6t
Xbit_r25_c143 bl[143] br[143] wl[25] vdd gnd cell_6t
Xbit_r26_c143 bl[143] br[143] wl[26] vdd gnd cell_6t
Xbit_r27_c143 bl[143] br[143] wl[27] vdd gnd cell_6t
Xbit_r28_c143 bl[143] br[143] wl[28] vdd gnd cell_6t
Xbit_r29_c143 bl[143] br[143] wl[29] vdd gnd cell_6t
Xbit_r30_c143 bl[143] br[143] wl[30] vdd gnd cell_6t
Xbit_r31_c143 bl[143] br[143] wl[31] vdd gnd cell_6t
Xbit_r32_c143 bl[143] br[143] wl[32] vdd gnd cell_6t
Xbit_r33_c143 bl[143] br[143] wl[33] vdd gnd cell_6t
Xbit_r34_c143 bl[143] br[143] wl[34] vdd gnd cell_6t
Xbit_r35_c143 bl[143] br[143] wl[35] vdd gnd cell_6t
Xbit_r36_c143 bl[143] br[143] wl[36] vdd gnd cell_6t
Xbit_r37_c143 bl[143] br[143] wl[37] vdd gnd cell_6t
Xbit_r38_c143 bl[143] br[143] wl[38] vdd gnd cell_6t
Xbit_r39_c143 bl[143] br[143] wl[39] vdd gnd cell_6t
Xbit_r40_c143 bl[143] br[143] wl[40] vdd gnd cell_6t
Xbit_r41_c143 bl[143] br[143] wl[41] vdd gnd cell_6t
Xbit_r42_c143 bl[143] br[143] wl[42] vdd gnd cell_6t
Xbit_r43_c143 bl[143] br[143] wl[43] vdd gnd cell_6t
Xbit_r44_c143 bl[143] br[143] wl[44] vdd gnd cell_6t
Xbit_r45_c143 bl[143] br[143] wl[45] vdd gnd cell_6t
Xbit_r46_c143 bl[143] br[143] wl[46] vdd gnd cell_6t
Xbit_r47_c143 bl[143] br[143] wl[47] vdd gnd cell_6t
Xbit_r48_c143 bl[143] br[143] wl[48] vdd gnd cell_6t
Xbit_r49_c143 bl[143] br[143] wl[49] vdd gnd cell_6t
Xbit_r50_c143 bl[143] br[143] wl[50] vdd gnd cell_6t
Xbit_r51_c143 bl[143] br[143] wl[51] vdd gnd cell_6t
Xbit_r52_c143 bl[143] br[143] wl[52] vdd gnd cell_6t
Xbit_r53_c143 bl[143] br[143] wl[53] vdd gnd cell_6t
Xbit_r54_c143 bl[143] br[143] wl[54] vdd gnd cell_6t
Xbit_r55_c143 bl[143] br[143] wl[55] vdd gnd cell_6t
Xbit_r56_c143 bl[143] br[143] wl[56] vdd gnd cell_6t
Xbit_r57_c143 bl[143] br[143] wl[57] vdd gnd cell_6t
Xbit_r58_c143 bl[143] br[143] wl[58] vdd gnd cell_6t
Xbit_r59_c143 bl[143] br[143] wl[59] vdd gnd cell_6t
Xbit_r60_c143 bl[143] br[143] wl[60] vdd gnd cell_6t
Xbit_r61_c143 bl[143] br[143] wl[61] vdd gnd cell_6t
Xbit_r62_c143 bl[143] br[143] wl[62] vdd gnd cell_6t
Xbit_r63_c143 bl[143] br[143] wl[63] vdd gnd cell_6t
Xbit_r64_c143 bl[143] br[143] wl[64] vdd gnd cell_6t
Xbit_r65_c143 bl[143] br[143] wl[65] vdd gnd cell_6t
Xbit_r66_c143 bl[143] br[143] wl[66] vdd gnd cell_6t
Xbit_r67_c143 bl[143] br[143] wl[67] vdd gnd cell_6t
Xbit_r68_c143 bl[143] br[143] wl[68] vdd gnd cell_6t
Xbit_r69_c143 bl[143] br[143] wl[69] vdd gnd cell_6t
Xbit_r70_c143 bl[143] br[143] wl[70] vdd gnd cell_6t
Xbit_r71_c143 bl[143] br[143] wl[71] vdd gnd cell_6t
Xbit_r72_c143 bl[143] br[143] wl[72] vdd gnd cell_6t
Xbit_r73_c143 bl[143] br[143] wl[73] vdd gnd cell_6t
Xbit_r74_c143 bl[143] br[143] wl[74] vdd gnd cell_6t
Xbit_r75_c143 bl[143] br[143] wl[75] vdd gnd cell_6t
Xbit_r76_c143 bl[143] br[143] wl[76] vdd gnd cell_6t
Xbit_r77_c143 bl[143] br[143] wl[77] vdd gnd cell_6t
Xbit_r78_c143 bl[143] br[143] wl[78] vdd gnd cell_6t
Xbit_r79_c143 bl[143] br[143] wl[79] vdd gnd cell_6t
Xbit_r80_c143 bl[143] br[143] wl[80] vdd gnd cell_6t
Xbit_r81_c143 bl[143] br[143] wl[81] vdd gnd cell_6t
Xbit_r82_c143 bl[143] br[143] wl[82] vdd gnd cell_6t
Xbit_r83_c143 bl[143] br[143] wl[83] vdd gnd cell_6t
Xbit_r84_c143 bl[143] br[143] wl[84] vdd gnd cell_6t
Xbit_r85_c143 bl[143] br[143] wl[85] vdd gnd cell_6t
Xbit_r86_c143 bl[143] br[143] wl[86] vdd gnd cell_6t
Xbit_r87_c143 bl[143] br[143] wl[87] vdd gnd cell_6t
Xbit_r88_c143 bl[143] br[143] wl[88] vdd gnd cell_6t
Xbit_r89_c143 bl[143] br[143] wl[89] vdd gnd cell_6t
Xbit_r90_c143 bl[143] br[143] wl[90] vdd gnd cell_6t
Xbit_r91_c143 bl[143] br[143] wl[91] vdd gnd cell_6t
Xbit_r92_c143 bl[143] br[143] wl[92] vdd gnd cell_6t
Xbit_r93_c143 bl[143] br[143] wl[93] vdd gnd cell_6t
Xbit_r94_c143 bl[143] br[143] wl[94] vdd gnd cell_6t
Xbit_r95_c143 bl[143] br[143] wl[95] vdd gnd cell_6t
Xbit_r96_c143 bl[143] br[143] wl[96] vdd gnd cell_6t
Xbit_r97_c143 bl[143] br[143] wl[97] vdd gnd cell_6t
Xbit_r98_c143 bl[143] br[143] wl[98] vdd gnd cell_6t
Xbit_r99_c143 bl[143] br[143] wl[99] vdd gnd cell_6t
Xbit_r100_c143 bl[143] br[143] wl[100] vdd gnd cell_6t
Xbit_r101_c143 bl[143] br[143] wl[101] vdd gnd cell_6t
Xbit_r102_c143 bl[143] br[143] wl[102] vdd gnd cell_6t
Xbit_r103_c143 bl[143] br[143] wl[103] vdd gnd cell_6t
Xbit_r104_c143 bl[143] br[143] wl[104] vdd gnd cell_6t
Xbit_r105_c143 bl[143] br[143] wl[105] vdd gnd cell_6t
Xbit_r106_c143 bl[143] br[143] wl[106] vdd gnd cell_6t
Xbit_r107_c143 bl[143] br[143] wl[107] vdd gnd cell_6t
Xbit_r108_c143 bl[143] br[143] wl[108] vdd gnd cell_6t
Xbit_r109_c143 bl[143] br[143] wl[109] vdd gnd cell_6t
Xbit_r110_c143 bl[143] br[143] wl[110] vdd gnd cell_6t
Xbit_r111_c143 bl[143] br[143] wl[111] vdd gnd cell_6t
Xbit_r112_c143 bl[143] br[143] wl[112] vdd gnd cell_6t
Xbit_r113_c143 bl[143] br[143] wl[113] vdd gnd cell_6t
Xbit_r114_c143 bl[143] br[143] wl[114] vdd gnd cell_6t
Xbit_r115_c143 bl[143] br[143] wl[115] vdd gnd cell_6t
Xbit_r116_c143 bl[143] br[143] wl[116] vdd gnd cell_6t
Xbit_r117_c143 bl[143] br[143] wl[117] vdd gnd cell_6t
Xbit_r118_c143 bl[143] br[143] wl[118] vdd gnd cell_6t
Xbit_r119_c143 bl[143] br[143] wl[119] vdd gnd cell_6t
Xbit_r120_c143 bl[143] br[143] wl[120] vdd gnd cell_6t
Xbit_r121_c143 bl[143] br[143] wl[121] vdd gnd cell_6t
Xbit_r122_c143 bl[143] br[143] wl[122] vdd gnd cell_6t
Xbit_r123_c143 bl[143] br[143] wl[123] vdd gnd cell_6t
Xbit_r124_c143 bl[143] br[143] wl[124] vdd gnd cell_6t
Xbit_r125_c143 bl[143] br[143] wl[125] vdd gnd cell_6t
Xbit_r126_c143 bl[143] br[143] wl[126] vdd gnd cell_6t
Xbit_r127_c143 bl[143] br[143] wl[127] vdd gnd cell_6t
Xbit_r0_c144 bl[144] br[144] wl[0] vdd gnd cell_6t
Xbit_r1_c144 bl[144] br[144] wl[1] vdd gnd cell_6t
Xbit_r2_c144 bl[144] br[144] wl[2] vdd gnd cell_6t
Xbit_r3_c144 bl[144] br[144] wl[3] vdd gnd cell_6t
Xbit_r4_c144 bl[144] br[144] wl[4] vdd gnd cell_6t
Xbit_r5_c144 bl[144] br[144] wl[5] vdd gnd cell_6t
Xbit_r6_c144 bl[144] br[144] wl[6] vdd gnd cell_6t
Xbit_r7_c144 bl[144] br[144] wl[7] vdd gnd cell_6t
Xbit_r8_c144 bl[144] br[144] wl[8] vdd gnd cell_6t
Xbit_r9_c144 bl[144] br[144] wl[9] vdd gnd cell_6t
Xbit_r10_c144 bl[144] br[144] wl[10] vdd gnd cell_6t
Xbit_r11_c144 bl[144] br[144] wl[11] vdd gnd cell_6t
Xbit_r12_c144 bl[144] br[144] wl[12] vdd gnd cell_6t
Xbit_r13_c144 bl[144] br[144] wl[13] vdd gnd cell_6t
Xbit_r14_c144 bl[144] br[144] wl[14] vdd gnd cell_6t
Xbit_r15_c144 bl[144] br[144] wl[15] vdd gnd cell_6t
Xbit_r16_c144 bl[144] br[144] wl[16] vdd gnd cell_6t
Xbit_r17_c144 bl[144] br[144] wl[17] vdd gnd cell_6t
Xbit_r18_c144 bl[144] br[144] wl[18] vdd gnd cell_6t
Xbit_r19_c144 bl[144] br[144] wl[19] vdd gnd cell_6t
Xbit_r20_c144 bl[144] br[144] wl[20] vdd gnd cell_6t
Xbit_r21_c144 bl[144] br[144] wl[21] vdd gnd cell_6t
Xbit_r22_c144 bl[144] br[144] wl[22] vdd gnd cell_6t
Xbit_r23_c144 bl[144] br[144] wl[23] vdd gnd cell_6t
Xbit_r24_c144 bl[144] br[144] wl[24] vdd gnd cell_6t
Xbit_r25_c144 bl[144] br[144] wl[25] vdd gnd cell_6t
Xbit_r26_c144 bl[144] br[144] wl[26] vdd gnd cell_6t
Xbit_r27_c144 bl[144] br[144] wl[27] vdd gnd cell_6t
Xbit_r28_c144 bl[144] br[144] wl[28] vdd gnd cell_6t
Xbit_r29_c144 bl[144] br[144] wl[29] vdd gnd cell_6t
Xbit_r30_c144 bl[144] br[144] wl[30] vdd gnd cell_6t
Xbit_r31_c144 bl[144] br[144] wl[31] vdd gnd cell_6t
Xbit_r32_c144 bl[144] br[144] wl[32] vdd gnd cell_6t
Xbit_r33_c144 bl[144] br[144] wl[33] vdd gnd cell_6t
Xbit_r34_c144 bl[144] br[144] wl[34] vdd gnd cell_6t
Xbit_r35_c144 bl[144] br[144] wl[35] vdd gnd cell_6t
Xbit_r36_c144 bl[144] br[144] wl[36] vdd gnd cell_6t
Xbit_r37_c144 bl[144] br[144] wl[37] vdd gnd cell_6t
Xbit_r38_c144 bl[144] br[144] wl[38] vdd gnd cell_6t
Xbit_r39_c144 bl[144] br[144] wl[39] vdd gnd cell_6t
Xbit_r40_c144 bl[144] br[144] wl[40] vdd gnd cell_6t
Xbit_r41_c144 bl[144] br[144] wl[41] vdd gnd cell_6t
Xbit_r42_c144 bl[144] br[144] wl[42] vdd gnd cell_6t
Xbit_r43_c144 bl[144] br[144] wl[43] vdd gnd cell_6t
Xbit_r44_c144 bl[144] br[144] wl[44] vdd gnd cell_6t
Xbit_r45_c144 bl[144] br[144] wl[45] vdd gnd cell_6t
Xbit_r46_c144 bl[144] br[144] wl[46] vdd gnd cell_6t
Xbit_r47_c144 bl[144] br[144] wl[47] vdd gnd cell_6t
Xbit_r48_c144 bl[144] br[144] wl[48] vdd gnd cell_6t
Xbit_r49_c144 bl[144] br[144] wl[49] vdd gnd cell_6t
Xbit_r50_c144 bl[144] br[144] wl[50] vdd gnd cell_6t
Xbit_r51_c144 bl[144] br[144] wl[51] vdd gnd cell_6t
Xbit_r52_c144 bl[144] br[144] wl[52] vdd gnd cell_6t
Xbit_r53_c144 bl[144] br[144] wl[53] vdd gnd cell_6t
Xbit_r54_c144 bl[144] br[144] wl[54] vdd gnd cell_6t
Xbit_r55_c144 bl[144] br[144] wl[55] vdd gnd cell_6t
Xbit_r56_c144 bl[144] br[144] wl[56] vdd gnd cell_6t
Xbit_r57_c144 bl[144] br[144] wl[57] vdd gnd cell_6t
Xbit_r58_c144 bl[144] br[144] wl[58] vdd gnd cell_6t
Xbit_r59_c144 bl[144] br[144] wl[59] vdd gnd cell_6t
Xbit_r60_c144 bl[144] br[144] wl[60] vdd gnd cell_6t
Xbit_r61_c144 bl[144] br[144] wl[61] vdd gnd cell_6t
Xbit_r62_c144 bl[144] br[144] wl[62] vdd gnd cell_6t
Xbit_r63_c144 bl[144] br[144] wl[63] vdd gnd cell_6t
Xbit_r64_c144 bl[144] br[144] wl[64] vdd gnd cell_6t
Xbit_r65_c144 bl[144] br[144] wl[65] vdd gnd cell_6t
Xbit_r66_c144 bl[144] br[144] wl[66] vdd gnd cell_6t
Xbit_r67_c144 bl[144] br[144] wl[67] vdd gnd cell_6t
Xbit_r68_c144 bl[144] br[144] wl[68] vdd gnd cell_6t
Xbit_r69_c144 bl[144] br[144] wl[69] vdd gnd cell_6t
Xbit_r70_c144 bl[144] br[144] wl[70] vdd gnd cell_6t
Xbit_r71_c144 bl[144] br[144] wl[71] vdd gnd cell_6t
Xbit_r72_c144 bl[144] br[144] wl[72] vdd gnd cell_6t
Xbit_r73_c144 bl[144] br[144] wl[73] vdd gnd cell_6t
Xbit_r74_c144 bl[144] br[144] wl[74] vdd gnd cell_6t
Xbit_r75_c144 bl[144] br[144] wl[75] vdd gnd cell_6t
Xbit_r76_c144 bl[144] br[144] wl[76] vdd gnd cell_6t
Xbit_r77_c144 bl[144] br[144] wl[77] vdd gnd cell_6t
Xbit_r78_c144 bl[144] br[144] wl[78] vdd gnd cell_6t
Xbit_r79_c144 bl[144] br[144] wl[79] vdd gnd cell_6t
Xbit_r80_c144 bl[144] br[144] wl[80] vdd gnd cell_6t
Xbit_r81_c144 bl[144] br[144] wl[81] vdd gnd cell_6t
Xbit_r82_c144 bl[144] br[144] wl[82] vdd gnd cell_6t
Xbit_r83_c144 bl[144] br[144] wl[83] vdd gnd cell_6t
Xbit_r84_c144 bl[144] br[144] wl[84] vdd gnd cell_6t
Xbit_r85_c144 bl[144] br[144] wl[85] vdd gnd cell_6t
Xbit_r86_c144 bl[144] br[144] wl[86] vdd gnd cell_6t
Xbit_r87_c144 bl[144] br[144] wl[87] vdd gnd cell_6t
Xbit_r88_c144 bl[144] br[144] wl[88] vdd gnd cell_6t
Xbit_r89_c144 bl[144] br[144] wl[89] vdd gnd cell_6t
Xbit_r90_c144 bl[144] br[144] wl[90] vdd gnd cell_6t
Xbit_r91_c144 bl[144] br[144] wl[91] vdd gnd cell_6t
Xbit_r92_c144 bl[144] br[144] wl[92] vdd gnd cell_6t
Xbit_r93_c144 bl[144] br[144] wl[93] vdd gnd cell_6t
Xbit_r94_c144 bl[144] br[144] wl[94] vdd gnd cell_6t
Xbit_r95_c144 bl[144] br[144] wl[95] vdd gnd cell_6t
Xbit_r96_c144 bl[144] br[144] wl[96] vdd gnd cell_6t
Xbit_r97_c144 bl[144] br[144] wl[97] vdd gnd cell_6t
Xbit_r98_c144 bl[144] br[144] wl[98] vdd gnd cell_6t
Xbit_r99_c144 bl[144] br[144] wl[99] vdd gnd cell_6t
Xbit_r100_c144 bl[144] br[144] wl[100] vdd gnd cell_6t
Xbit_r101_c144 bl[144] br[144] wl[101] vdd gnd cell_6t
Xbit_r102_c144 bl[144] br[144] wl[102] vdd gnd cell_6t
Xbit_r103_c144 bl[144] br[144] wl[103] vdd gnd cell_6t
Xbit_r104_c144 bl[144] br[144] wl[104] vdd gnd cell_6t
Xbit_r105_c144 bl[144] br[144] wl[105] vdd gnd cell_6t
Xbit_r106_c144 bl[144] br[144] wl[106] vdd gnd cell_6t
Xbit_r107_c144 bl[144] br[144] wl[107] vdd gnd cell_6t
Xbit_r108_c144 bl[144] br[144] wl[108] vdd gnd cell_6t
Xbit_r109_c144 bl[144] br[144] wl[109] vdd gnd cell_6t
Xbit_r110_c144 bl[144] br[144] wl[110] vdd gnd cell_6t
Xbit_r111_c144 bl[144] br[144] wl[111] vdd gnd cell_6t
Xbit_r112_c144 bl[144] br[144] wl[112] vdd gnd cell_6t
Xbit_r113_c144 bl[144] br[144] wl[113] vdd gnd cell_6t
Xbit_r114_c144 bl[144] br[144] wl[114] vdd gnd cell_6t
Xbit_r115_c144 bl[144] br[144] wl[115] vdd gnd cell_6t
Xbit_r116_c144 bl[144] br[144] wl[116] vdd gnd cell_6t
Xbit_r117_c144 bl[144] br[144] wl[117] vdd gnd cell_6t
Xbit_r118_c144 bl[144] br[144] wl[118] vdd gnd cell_6t
Xbit_r119_c144 bl[144] br[144] wl[119] vdd gnd cell_6t
Xbit_r120_c144 bl[144] br[144] wl[120] vdd gnd cell_6t
Xbit_r121_c144 bl[144] br[144] wl[121] vdd gnd cell_6t
Xbit_r122_c144 bl[144] br[144] wl[122] vdd gnd cell_6t
Xbit_r123_c144 bl[144] br[144] wl[123] vdd gnd cell_6t
Xbit_r124_c144 bl[144] br[144] wl[124] vdd gnd cell_6t
Xbit_r125_c144 bl[144] br[144] wl[125] vdd gnd cell_6t
Xbit_r126_c144 bl[144] br[144] wl[126] vdd gnd cell_6t
Xbit_r127_c144 bl[144] br[144] wl[127] vdd gnd cell_6t
Xbit_r0_c145 bl[145] br[145] wl[0] vdd gnd cell_6t
Xbit_r1_c145 bl[145] br[145] wl[1] vdd gnd cell_6t
Xbit_r2_c145 bl[145] br[145] wl[2] vdd gnd cell_6t
Xbit_r3_c145 bl[145] br[145] wl[3] vdd gnd cell_6t
Xbit_r4_c145 bl[145] br[145] wl[4] vdd gnd cell_6t
Xbit_r5_c145 bl[145] br[145] wl[5] vdd gnd cell_6t
Xbit_r6_c145 bl[145] br[145] wl[6] vdd gnd cell_6t
Xbit_r7_c145 bl[145] br[145] wl[7] vdd gnd cell_6t
Xbit_r8_c145 bl[145] br[145] wl[8] vdd gnd cell_6t
Xbit_r9_c145 bl[145] br[145] wl[9] vdd gnd cell_6t
Xbit_r10_c145 bl[145] br[145] wl[10] vdd gnd cell_6t
Xbit_r11_c145 bl[145] br[145] wl[11] vdd gnd cell_6t
Xbit_r12_c145 bl[145] br[145] wl[12] vdd gnd cell_6t
Xbit_r13_c145 bl[145] br[145] wl[13] vdd gnd cell_6t
Xbit_r14_c145 bl[145] br[145] wl[14] vdd gnd cell_6t
Xbit_r15_c145 bl[145] br[145] wl[15] vdd gnd cell_6t
Xbit_r16_c145 bl[145] br[145] wl[16] vdd gnd cell_6t
Xbit_r17_c145 bl[145] br[145] wl[17] vdd gnd cell_6t
Xbit_r18_c145 bl[145] br[145] wl[18] vdd gnd cell_6t
Xbit_r19_c145 bl[145] br[145] wl[19] vdd gnd cell_6t
Xbit_r20_c145 bl[145] br[145] wl[20] vdd gnd cell_6t
Xbit_r21_c145 bl[145] br[145] wl[21] vdd gnd cell_6t
Xbit_r22_c145 bl[145] br[145] wl[22] vdd gnd cell_6t
Xbit_r23_c145 bl[145] br[145] wl[23] vdd gnd cell_6t
Xbit_r24_c145 bl[145] br[145] wl[24] vdd gnd cell_6t
Xbit_r25_c145 bl[145] br[145] wl[25] vdd gnd cell_6t
Xbit_r26_c145 bl[145] br[145] wl[26] vdd gnd cell_6t
Xbit_r27_c145 bl[145] br[145] wl[27] vdd gnd cell_6t
Xbit_r28_c145 bl[145] br[145] wl[28] vdd gnd cell_6t
Xbit_r29_c145 bl[145] br[145] wl[29] vdd gnd cell_6t
Xbit_r30_c145 bl[145] br[145] wl[30] vdd gnd cell_6t
Xbit_r31_c145 bl[145] br[145] wl[31] vdd gnd cell_6t
Xbit_r32_c145 bl[145] br[145] wl[32] vdd gnd cell_6t
Xbit_r33_c145 bl[145] br[145] wl[33] vdd gnd cell_6t
Xbit_r34_c145 bl[145] br[145] wl[34] vdd gnd cell_6t
Xbit_r35_c145 bl[145] br[145] wl[35] vdd gnd cell_6t
Xbit_r36_c145 bl[145] br[145] wl[36] vdd gnd cell_6t
Xbit_r37_c145 bl[145] br[145] wl[37] vdd gnd cell_6t
Xbit_r38_c145 bl[145] br[145] wl[38] vdd gnd cell_6t
Xbit_r39_c145 bl[145] br[145] wl[39] vdd gnd cell_6t
Xbit_r40_c145 bl[145] br[145] wl[40] vdd gnd cell_6t
Xbit_r41_c145 bl[145] br[145] wl[41] vdd gnd cell_6t
Xbit_r42_c145 bl[145] br[145] wl[42] vdd gnd cell_6t
Xbit_r43_c145 bl[145] br[145] wl[43] vdd gnd cell_6t
Xbit_r44_c145 bl[145] br[145] wl[44] vdd gnd cell_6t
Xbit_r45_c145 bl[145] br[145] wl[45] vdd gnd cell_6t
Xbit_r46_c145 bl[145] br[145] wl[46] vdd gnd cell_6t
Xbit_r47_c145 bl[145] br[145] wl[47] vdd gnd cell_6t
Xbit_r48_c145 bl[145] br[145] wl[48] vdd gnd cell_6t
Xbit_r49_c145 bl[145] br[145] wl[49] vdd gnd cell_6t
Xbit_r50_c145 bl[145] br[145] wl[50] vdd gnd cell_6t
Xbit_r51_c145 bl[145] br[145] wl[51] vdd gnd cell_6t
Xbit_r52_c145 bl[145] br[145] wl[52] vdd gnd cell_6t
Xbit_r53_c145 bl[145] br[145] wl[53] vdd gnd cell_6t
Xbit_r54_c145 bl[145] br[145] wl[54] vdd gnd cell_6t
Xbit_r55_c145 bl[145] br[145] wl[55] vdd gnd cell_6t
Xbit_r56_c145 bl[145] br[145] wl[56] vdd gnd cell_6t
Xbit_r57_c145 bl[145] br[145] wl[57] vdd gnd cell_6t
Xbit_r58_c145 bl[145] br[145] wl[58] vdd gnd cell_6t
Xbit_r59_c145 bl[145] br[145] wl[59] vdd gnd cell_6t
Xbit_r60_c145 bl[145] br[145] wl[60] vdd gnd cell_6t
Xbit_r61_c145 bl[145] br[145] wl[61] vdd gnd cell_6t
Xbit_r62_c145 bl[145] br[145] wl[62] vdd gnd cell_6t
Xbit_r63_c145 bl[145] br[145] wl[63] vdd gnd cell_6t
Xbit_r64_c145 bl[145] br[145] wl[64] vdd gnd cell_6t
Xbit_r65_c145 bl[145] br[145] wl[65] vdd gnd cell_6t
Xbit_r66_c145 bl[145] br[145] wl[66] vdd gnd cell_6t
Xbit_r67_c145 bl[145] br[145] wl[67] vdd gnd cell_6t
Xbit_r68_c145 bl[145] br[145] wl[68] vdd gnd cell_6t
Xbit_r69_c145 bl[145] br[145] wl[69] vdd gnd cell_6t
Xbit_r70_c145 bl[145] br[145] wl[70] vdd gnd cell_6t
Xbit_r71_c145 bl[145] br[145] wl[71] vdd gnd cell_6t
Xbit_r72_c145 bl[145] br[145] wl[72] vdd gnd cell_6t
Xbit_r73_c145 bl[145] br[145] wl[73] vdd gnd cell_6t
Xbit_r74_c145 bl[145] br[145] wl[74] vdd gnd cell_6t
Xbit_r75_c145 bl[145] br[145] wl[75] vdd gnd cell_6t
Xbit_r76_c145 bl[145] br[145] wl[76] vdd gnd cell_6t
Xbit_r77_c145 bl[145] br[145] wl[77] vdd gnd cell_6t
Xbit_r78_c145 bl[145] br[145] wl[78] vdd gnd cell_6t
Xbit_r79_c145 bl[145] br[145] wl[79] vdd gnd cell_6t
Xbit_r80_c145 bl[145] br[145] wl[80] vdd gnd cell_6t
Xbit_r81_c145 bl[145] br[145] wl[81] vdd gnd cell_6t
Xbit_r82_c145 bl[145] br[145] wl[82] vdd gnd cell_6t
Xbit_r83_c145 bl[145] br[145] wl[83] vdd gnd cell_6t
Xbit_r84_c145 bl[145] br[145] wl[84] vdd gnd cell_6t
Xbit_r85_c145 bl[145] br[145] wl[85] vdd gnd cell_6t
Xbit_r86_c145 bl[145] br[145] wl[86] vdd gnd cell_6t
Xbit_r87_c145 bl[145] br[145] wl[87] vdd gnd cell_6t
Xbit_r88_c145 bl[145] br[145] wl[88] vdd gnd cell_6t
Xbit_r89_c145 bl[145] br[145] wl[89] vdd gnd cell_6t
Xbit_r90_c145 bl[145] br[145] wl[90] vdd gnd cell_6t
Xbit_r91_c145 bl[145] br[145] wl[91] vdd gnd cell_6t
Xbit_r92_c145 bl[145] br[145] wl[92] vdd gnd cell_6t
Xbit_r93_c145 bl[145] br[145] wl[93] vdd gnd cell_6t
Xbit_r94_c145 bl[145] br[145] wl[94] vdd gnd cell_6t
Xbit_r95_c145 bl[145] br[145] wl[95] vdd gnd cell_6t
Xbit_r96_c145 bl[145] br[145] wl[96] vdd gnd cell_6t
Xbit_r97_c145 bl[145] br[145] wl[97] vdd gnd cell_6t
Xbit_r98_c145 bl[145] br[145] wl[98] vdd gnd cell_6t
Xbit_r99_c145 bl[145] br[145] wl[99] vdd gnd cell_6t
Xbit_r100_c145 bl[145] br[145] wl[100] vdd gnd cell_6t
Xbit_r101_c145 bl[145] br[145] wl[101] vdd gnd cell_6t
Xbit_r102_c145 bl[145] br[145] wl[102] vdd gnd cell_6t
Xbit_r103_c145 bl[145] br[145] wl[103] vdd gnd cell_6t
Xbit_r104_c145 bl[145] br[145] wl[104] vdd gnd cell_6t
Xbit_r105_c145 bl[145] br[145] wl[105] vdd gnd cell_6t
Xbit_r106_c145 bl[145] br[145] wl[106] vdd gnd cell_6t
Xbit_r107_c145 bl[145] br[145] wl[107] vdd gnd cell_6t
Xbit_r108_c145 bl[145] br[145] wl[108] vdd gnd cell_6t
Xbit_r109_c145 bl[145] br[145] wl[109] vdd gnd cell_6t
Xbit_r110_c145 bl[145] br[145] wl[110] vdd gnd cell_6t
Xbit_r111_c145 bl[145] br[145] wl[111] vdd gnd cell_6t
Xbit_r112_c145 bl[145] br[145] wl[112] vdd gnd cell_6t
Xbit_r113_c145 bl[145] br[145] wl[113] vdd gnd cell_6t
Xbit_r114_c145 bl[145] br[145] wl[114] vdd gnd cell_6t
Xbit_r115_c145 bl[145] br[145] wl[115] vdd gnd cell_6t
Xbit_r116_c145 bl[145] br[145] wl[116] vdd gnd cell_6t
Xbit_r117_c145 bl[145] br[145] wl[117] vdd gnd cell_6t
Xbit_r118_c145 bl[145] br[145] wl[118] vdd gnd cell_6t
Xbit_r119_c145 bl[145] br[145] wl[119] vdd gnd cell_6t
Xbit_r120_c145 bl[145] br[145] wl[120] vdd gnd cell_6t
Xbit_r121_c145 bl[145] br[145] wl[121] vdd gnd cell_6t
Xbit_r122_c145 bl[145] br[145] wl[122] vdd gnd cell_6t
Xbit_r123_c145 bl[145] br[145] wl[123] vdd gnd cell_6t
Xbit_r124_c145 bl[145] br[145] wl[124] vdd gnd cell_6t
Xbit_r125_c145 bl[145] br[145] wl[125] vdd gnd cell_6t
Xbit_r126_c145 bl[145] br[145] wl[126] vdd gnd cell_6t
Xbit_r127_c145 bl[145] br[145] wl[127] vdd gnd cell_6t
Xbit_r0_c146 bl[146] br[146] wl[0] vdd gnd cell_6t
Xbit_r1_c146 bl[146] br[146] wl[1] vdd gnd cell_6t
Xbit_r2_c146 bl[146] br[146] wl[2] vdd gnd cell_6t
Xbit_r3_c146 bl[146] br[146] wl[3] vdd gnd cell_6t
Xbit_r4_c146 bl[146] br[146] wl[4] vdd gnd cell_6t
Xbit_r5_c146 bl[146] br[146] wl[5] vdd gnd cell_6t
Xbit_r6_c146 bl[146] br[146] wl[6] vdd gnd cell_6t
Xbit_r7_c146 bl[146] br[146] wl[7] vdd gnd cell_6t
Xbit_r8_c146 bl[146] br[146] wl[8] vdd gnd cell_6t
Xbit_r9_c146 bl[146] br[146] wl[9] vdd gnd cell_6t
Xbit_r10_c146 bl[146] br[146] wl[10] vdd gnd cell_6t
Xbit_r11_c146 bl[146] br[146] wl[11] vdd gnd cell_6t
Xbit_r12_c146 bl[146] br[146] wl[12] vdd gnd cell_6t
Xbit_r13_c146 bl[146] br[146] wl[13] vdd gnd cell_6t
Xbit_r14_c146 bl[146] br[146] wl[14] vdd gnd cell_6t
Xbit_r15_c146 bl[146] br[146] wl[15] vdd gnd cell_6t
Xbit_r16_c146 bl[146] br[146] wl[16] vdd gnd cell_6t
Xbit_r17_c146 bl[146] br[146] wl[17] vdd gnd cell_6t
Xbit_r18_c146 bl[146] br[146] wl[18] vdd gnd cell_6t
Xbit_r19_c146 bl[146] br[146] wl[19] vdd gnd cell_6t
Xbit_r20_c146 bl[146] br[146] wl[20] vdd gnd cell_6t
Xbit_r21_c146 bl[146] br[146] wl[21] vdd gnd cell_6t
Xbit_r22_c146 bl[146] br[146] wl[22] vdd gnd cell_6t
Xbit_r23_c146 bl[146] br[146] wl[23] vdd gnd cell_6t
Xbit_r24_c146 bl[146] br[146] wl[24] vdd gnd cell_6t
Xbit_r25_c146 bl[146] br[146] wl[25] vdd gnd cell_6t
Xbit_r26_c146 bl[146] br[146] wl[26] vdd gnd cell_6t
Xbit_r27_c146 bl[146] br[146] wl[27] vdd gnd cell_6t
Xbit_r28_c146 bl[146] br[146] wl[28] vdd gnd cell_6t
Xbit_r29_c146 bl[146] br[146] wl[29] vdd gnd cell_6t
Xbit_r30_c146 bl[146] br[146] wl[30] vdd gnd cell_6t
Xbit_r31_c146 bl[146] br[146] wl[31] vdd gnd cell_6t
Xbit_r32_c146 bl[146] br[146] wl[32] vdd gnd cell_6t
Xbit_r33_c146 bl[146] br[146] wl[33] vdd gnd cell_6t
Xbit_r34_c146 bl[146] br[146] wl[34] vdd gnd cell_6t
Xbit_r35_c146 bl[146] br[146] wl[35] vdd gnd cell_6t
Xbit_r36_c146 bl[146] br[146] wl[36] vdd gnd cell_6t
Xbit_r37_c146 bl[146] br[146] wl[37] vdd gnd cell_6t
Xbit_r38_c146 bl[146] br[146] wl[38] vdd gnd cell_6t
Xbit_r39_c146 bl[146] br[146] wl[39] vdd gnd cell_6t
Xbit_r40_c146 bl[146] br[146] wl[40] vdd gnd cell_6t
Xbit_r41_c146 bl[146] br[146] wl[41] vdd gnd cell_6t
Xbit_r42_c146 bl[146] br[146] wl[42] vdd gnd cell_6t
Xbit_r43_c146 bl[146] br[146] wl[43] vdd gnd cell_6t
Xbit_r44_c146 bl[146] br[146] wl[44] vdd gnd cell_6t
Xbit_r45_c146 bl[146] br[146] wl[45] vdd gnd cell_6t
Xbit_r46_c146 bl[146] br[146] wl[46] vdd gnd cell_6t
Xbit_r47_c146 bl[146] br[146] wl[47] vdd gnd cell_6t
Xbit_r48_c146 bl[146] br[146] wl[48] vdd gnd cell_6t
Xbit_r49_c146 bl[146] br[146] wl[49] vdd gnd cell_6t
Xbit_r50_c146 bl[146] br[146] wl[50] vdd gnd cell_6t
Xbit_r51_c146 bl[146] br[146] wl[51] vdd gnd cell_6t
Xbit_r52_c146 bl[146] br[146] wl[52] vdd gnd cell_6t
Xbit_r53_c146 bl[146] br[146] wl[53] vdd gnd cell_6t
Xbit_r54_c146 bl[146] br[146] wl[54] vdd gnd cell_6t
Xbit_r55_c146 bl[146] br[146] wl[55] vdd gnd cell_6t
Xbit_r56_c146 bl[146] br[146] wl[56] vdd gnd cell_6t
Xbit_r57_c146 bl[146] br[146] wl[57] vdd gnd cell_6t
Xbit_r58_c146 bl[146] br[146] wl[58] vdd gnd cell_6t
Xbit_r59_c146 bl[146] br[146] wl[59] vdd gnd cell_6t
Xbit_r60_c146 bl[146] br[146] wl[60] vdd gnd cell_6t
Xbit_r61_c146 bl[146] br[146] wl[61] vdd gnd cell_6t
Xbit_r62_c146 bl[146] br[146] wl[62] vdd gnd cell_6t
Xbit_r63_c146 bl[146] br[146] wl[63] vdd gnd cell_6t
Xbit_r64_c146 bl[146] br[146] wl[64] vdd gnd cell_6t
Xbit_r65_c146 bl[146] br[146] wl[65] vdd gnd cell_6t
Xbit_r66_c146 bl[146] br[146] wl[66] vdd gnd cell_6t
Xbit_r67_c146 bl[146] br[146] wl[67] vdd gnd cell_6t
Xbit_r68_c146 bl[146] br[146] wl[68] vdd gnd cell_6t
Xbit_r69_c146 bl[146] br[146] wl[69] vdd gnd cell_6t
Xbit_r70_c146 bl[146] br[146] wl[70] vdd gnd cell_6t
Xbit_r71_c146 bl[146] br[146] wl[71] vdd gnd cell_6t
Xbit_r72_c146 bl[146] br[146] wl[72] vdd gnd cell_6t
Xbit_r73_c146 bl[146] br[146] wl[73] vdd gnd cell_6t
Xbit_r74_c146 bl[146] br[146] wl[74] vdd gnd cell_6t
Xbit_r75_c146 bl[146] br[146] wl[75] vdd gnd cell_6t
Xbit_r76_c146 bl[146] br[146] wl[76] vdd gnd cell_6t
Xbit_r77_c146 bl[146] br[146] wl[77] vdd gnd cell_6t
Xbit_r78_c146 bl[146] br[146] wl[78] vdd gnd cell_6t
Xbit_r79_c146 bl[146] br[146] wl[79] vdd gnd cell_6t
Xbit_r80_c146 bl[146] br[146] wl[80] vdd gnd cell_6t
Xbit_r81_c146 bl[146] br[146] wl[81] vdd gnd cell_6t
Xbit_r82_c146 bl[146] br[146] wl[82] vdd gnd cell_6t
Xbit_r83_c146 bl[146] br[146] wl[83] vdd gnd cell_6t
Xbit_r84_c146 bl[146] br[146] wl[84] vdd gnd cell_6t
Xbit_r85_c146 bl[146] br[146] wl[85] vdd gnd cell_6t
Xbit_r86_c146 bl[146] br[146] wl[86] vdd gnd cell_6t
Xbit_r87_c146 bl[146] br[146] wl[87] vdd gnd cell_6t
Xbit_r88_c146 bl[146] br[146] wl[88] vdd gnd cell_6t
Xbit_r89_c146 bl[146] br[146] wl[89] vdd gnd cell_6t
Xbit_r90_c146 bl[146] br[146] wl[90] vdd gnd cell_6t
Xbit_r91_c146 bl[146] br[146] wl[91] vdd gnd cell_6t
Xbit_r92_c146 bl[146] br[146] wl[92] vdd gnd cell_6t
Xbit_r93_c146 bl[146] br[146] wl[93] vdd gnd cell_6t
Xbit_r94_c146 bl[146] br[146] wl[94] vdd gnd cell_6t
Xbit_r95_c146 bl[146] br[146] wl[95] vdd gnd cell_6t
Xbit_r96_c146 bl[146] br[146] wl[96] vdd gnd cell_6t
Xbit_r97_c146 bl[146] br[146] wl[97] vdd gnd cell_6t
Xbit_r98_c146 bl[146] br[146] wl[98] vdd gnd cell_6t
Xbit_r99_c146 bl[146] br[146] wl[99] vdd gnd cell_6t
Xbit_r100_c146 bl[146] br[146] wl[100] vdd gnd cell_6t
Xbit_r101_c146 bl[146] br[146] wl[101] vdd gnd cell_6t
Xbit_r102_c146 bl[146] br[146] wl[102] vdd gnd cell_6t
Xbit_r103_c146 bl[146] br[146] wl[103] vdd gnd cell_6t
Xbit_r104_c146 bl[146] br[146] wl[104] vdd gnd cell_6t
Xbit_r105_c146 bl[146] br[146] wl[105] vdd gnd cell_6t
Xbit_r106_c146 bl[146] br[146] wl[106] vdd gnd cell_6t
Xbit_r107_c146 bl[146] br[146] wl[107] vdd gnd cell_6t
Xbit_r108_c146 bl[146] br[146] wl[108] vdd gnd cell_6t
Xbit_r109_c146 bl[146] br[146] wl[109] vdd gnd cell_6t
Xbit_r110_c146 bl[146] br[146] wl[110] vdd gnd cell_6t
Xbit_r111_c146 bl[146] br[146] wl[111] vdd gnd cell_6t
Xbit_r112_c146 bl[146] br[146] wl[112] vdd gnd cell_6t
Xbit_r113_c146 bl[146] br[146] wl[113] vdd gnd cell_6t
Xbit_r114_c146 bl[146] br[146] wl[114] vdd gnd cell_6t
Xbit_r115_c146 bl[146] br[146] wl[115] vdd gnd cell_6t
Xbit_r116_c146 bl[146] br[146] wl[116] vdd gnd cell_6t
Xbit_r117_c146 bl[146] br[146] wl[117] vdd gnd cell_6t
Xbit_r118_c146 bl[146] br[146] wl[118] vdd gnd cell_6t
Xbit_r119_c146 bl[146] br[146] wl[119] vdd gnd cell_6t
Xbit_r120_c146 bl[146] br[146] wl[120] vdd gnd cell_6t
Xbit_r121_c146 bl[146] br[146] wl[121] vdd gnd cell_6t
Xbit_r122_c146 bl[146] br[146] wl[122] vdd gnd cell_6t
Xbit_r123_c146 bl[146] br[146] wl[123] vdd gnd cell_6t
Xbit_r124_c146 bl[146] br[146] wl[124] vdd gnd cell_6t
Xbit_r125_c146 bl[146] br[146] wl[125] vdd gnd cell_6t
Xbit_r126_c146 bl[146] br[146] wl[126] vdd gnd cell_6t
Xbit_r127_c146 bl[146] br[146] wl[127] vdd gnd cell_6t
Xbit_r0_c147 bl[147] br[147] wl[0] vdd gnd cell_6t
Xbit_r1_c147 bl[147] br[147] wl[1] vdd gnd cell_6t
Xbit_r2_c147 bl[147] br[147] wl[2] vdd gnd cell_6t
Xbit_r3_c147 bl[147] br[147] wl[3] vdd gnd cell_6t
Xbit_r4_c147 bl[147] br[147] wl[4] vdd gnd cell_6t
Xbit_r5_c147 bl[147] br[147] wl[5] vdd gnd cell_6t
Xbit_r6_c147 bl[147] br[147] wl[6] vdd gnd cell_6t
Xbit_r7_c147 bl[147] br[147] wl[7] vdd gnd cell_6t
Xbit_r8_c147 bl[147] br[147] wl[8] vdd gnd cell_6t
Xbit_r9_c147 bl[147] br[147] wl[9] vdd gnd cell_6t
Xbit_r10_c147 bl[147] br[147] wl[10] vdd gnd cell_6t
Xbit_r11_c147 bl[147] br[147] wl[11] vdd gnd cell_6t
Xbit_r12_c147 bl[147] br[147] wl[12] vdd gnd cell_6t
Xbit_r13_c147 bl[147] br[147] wl[13] vdd gnd cell_6t
Xbit_r14_c147 bl[147] br[147] wl[14] vdd gnd cell_6t
Xbit_r15_c147 bl[147] br[147] wl[15] vdd gnd cell_6t
Xbit_r16_c147 bl[147] br[147] wl[16] vdd gnd cell_6t
Xbit_r17_c147 bl[147] br[147] wl[17] vdd gnd cell_6t
Xbit_r18_c147 bl[147] br[147] wl[18] vdd gnd cell_6t
Xbit_r19_c147 bl[147] br[147] wl[19] vdd gnd cell_6t
Xbit_r20_c147 bl[147] br[147] wl[20] vdd gnd cell_6t
Xbit_r21_c147 bl[147] br[147] wl[21] vdd gnd cell_6t
Xbit_r22_c147 bl[147] br[147] wl[22] vdd gnd cell_6t
Xbit_r23_c147 bl[147] br[147] wl[23] vdd gnd cell_6t
Xbit_r24_c147 bl[147] br[147] wl[24] vdd gnd cell_6t
Xbit_r25_c147 bl[147] br[147] wl[25] vdd gnd cell_6t
Xbit_r26_c147 bl[147] br[147] wl[26] vdd gnd cell_6t
Xbit_r27_c147 bl[147] br[147] wl[27] vdd gnd cell_6t
Xbit_r28_c147 bl[147] br[147] wl[28] vdd gnd cell_6t
Xbit_r29_c147 bl[147] br[147] wl[29] vdd gnd cell_6t
Xbit_r30_c147 bl[147] br[147] wl[30] vdd gnd cell_6t
Xbit_r31_c147 bl[147] br[147] wl[31] vdd gnd cell_6t
Xbit_r32_c147 bl[147] br[147] wl[32] vdd gnd cell_6t
Xbit_r33_c147 bl[147] br[147] wl[33] vdd gnd cell_6t
Xbit_r34_c147 bl[147] br[147] wl[34] vdd gnd cell_6t
Xbit_r35_c147 bl[147] br[147] wl[35] vdd gnd cell_6t
Xbit_r36_c147 bl[147] br[147] wl[36] vdd gnd cell_6t
Xbit_r37_c147 bl[147] br[147] wl[37] vdd gnd cell_6t
Xbit_r38_c147 bl[147] br[147] wl[38] vdd gnd cell_6t
Xbit_r39_c147 bl[147] br[147] wl[39] vdd gnd cell_6t
Xbit_r40_c147 bl[147] br[147] wl[40] vdd gnd cell_6t
Xbit_r41_c147 bl[147] br[147] wl[41] vdd gnd cell_6t
Xbit_r42_c147 bl[147] br[147] wl[42] vdd gnd cell_6t
Xbit_r43_c147 bl[147] br[147] wl[43] vdd gnd cell_6t
Xbit_r44_c147 bl[147] br[147] wl[44] vdd gnd cell_6t
Xbit_r45_c147 bl[147] br[147] wl[45] vdd gnd cell_6t
Xbit_r46_c147 bl[147] br[147] wl[46] vdd gnd cell_6t
Xbit_r47_c147 bl[147] br[147] wl[47] vdd gnd cell_6t
Xbit_r48_c147 bl[147] br[147] wl[48] vdd gnd cell_6t
Xbit_r49_c147 bl[147] br[147] wl[49] vdd gnd cell_6t
Xbit_r50_c147 bl[147] br[147] wl[50] vdd gnd cell_6t
Xbit_r51_c147 bl[147] br[147] wl[51] vdd gnd cell_6t
Xbit_r52_c147 bl[147] br[147] wl[52] vdd gnd cell_6t
Xbit_r53_c147 bl[147] br[147] wl[53] vdd gnd cell_6t
Xbit_r54_c147 bl[147] br[147] wl[54] vdd gnd cell_6t
Xbit_r55_c147 bl[147] br[147] wl[55] vdd gnd cell_6t
Xbit_r56_c147 bl[147] br[147] wl[56] vdd gnd cell_6t
Xbit_r57_c147 bl[147] br[147] wl[57] vdd gnd cell_6t
Xbit_r58_c147 bl[147] br[147] wl[58] vdd gnd cell_6t
Xbit_r59_c147 bl[147] br[147] wl[59] vdd gnd cell_6t
Xbit_r60_c147 bl[147] br[147] wl[60] vdd gnd cell_6t
Xbit_r61_c147 bl[147] br[147] wl[61] vdd gnd cell_6t
Xbit_r62_c147 bl[147] br[147] wl[62] vdd gnd cell_6t
Xbit_r63_c147 bl[147] br[147] wl[63] vdd gnd cell_6t
Xbit_r64_c147 bl[147] br[147] wl[64] vdd gnd cell_6t
Xbit_r65_c147 bl[147] br[147] wl[65] vdd gnd cell_6t
Xbit_r66_c147 bl[147] br[147] wl[66] vdd gnd cell_6t
Xbit_r67_c147 bl[147] br[147] wl[67] vdd gnd cell_6t
Xbit_r68_c147 bl[147] br[147] wl[68] vdd gnd cell_6t
Xbit_r69_c147 bl[147] br[147] wl[69] vdd gnd cell_6t
Xbit_r70_c147 bl[147] br[147] wl[70] vdd gnd cell_6t
Xbit_r71_c147 bl[147] br[147] wl[71] vdd gnd cell_6t
Xbit_r72_c147 bl[147] br[147] wl[72] vdd gnd cell_6t
Xbit_r73_c147 bl[147] br[147] wl[73] vdd gnd cell_6t
Xbit_r74_c147 bl[147] br[147] wl[74] vdd gnd cell_6t
Xbit_r75_c147 bl[147] br[147] wl[75] vdd gnd cell_6t
Xbit_r76_c147 bl[147] br[147] wl[76] vdd gnd cell_6t
Xbit_r77_c147 bl[147] br[147] wl[77] vdd gnd cell_6t
Xbit_r78_c147 bl[147] br[147] wl[78] vdd gnd cell_6t
Xbit_r79_c147 bl[147] br[147] wl[79] vdd gnd cell_6t
Xbit_r80_c147 bl[147] br[147] wl[80] vdd gnd cell_6t
Xbit_r81_c147 bl[147] br[147] wl[81] vdd gnd cell_6t
Xbit_r82_c147 bl[147] br[147] wl[82] vdd gnd cell_6t
Xbit_r83_c147 bl[147] br[147] wl[83] vdd gnd cell_6t
Xbit_r84_c147 bl[147] br[147] wl[84] vdd gnd cell_6t
Xbit_r85_c147 bl[147] br[147] wl[85] vdd gnd cell_6t
Xbit_r86_c147 bl[147] br[147] wl[86] vdd gnd cell_6t
Xbit_r87_c147 bl[147] br[147] wl[87] vdd gnd cell_6t
Xbit_r88_c147 bl[147] br[147] wl[88] vdd gnd cell_6t
Xbit_r89_c147 bl[147] br[147] wl[89] vdd gnd cell_6t
Xbit_r90_c147 bl[147] br[147] wl[90] vdd gnd cell_6t
Xbit_r91_c147 bl[147] br[147] wl[91] vdd gnd cell_6t
Xbit_r92_c147 bl[147] br[147] wl[92] vdd gnd cell_6t
Xbit_r93_c147 bl[147] br[147] wl[93] vdd gnd cell_6t
Xbit_r94_c147 bl[147] br[147] wl[94] vdd gnd cell_6t
Xbit_r95_c147 bl[147] br[147] wl[95] vdd gnd cell_6t
Xbit_r96_c147 bl[147] br[147] wl[96] vdd gnd cell_6t
Xbit_r97_c147 bl[147] br[147] wl[97] vdd gnd cell_6t
Xbit_r98_c147 bl[147] br[147] wl[98] vdd gnd cell_6t
Xbit_r99_c147 bl[147] br[147] wl[99] vdd gnd cell_6t
Xbit_r100_c147 bl[147] br[147] wl[100] vdd gnd cell_6t
Xbit_r101_c147 bl[147] br[147] wl[101] vdd gnd cell_6t
Xbit_r102_c147 bl[147] br[147] wl[102] vdd gnd cell_6t
Xbit_r103_c147 bl[147] br[147] wl[103] vdd gnd cell_6t
Xbit_r104_c147 bl[147] br[147] wl[104] vdd gnd cell_6t
Xbit_r105_c147 bl[147] br[147] wl[105] vdd gnd cell_6t
Xbit_r106_c147 bl[147] br[147] wl[106] vdd gnd cell_6t
Xbit_r107_c147 bl[147] br[147] wl[107] vdd gnd cell_6t
Xbit_r108_c147 bl[147] br[147] wl[108] vdd gnd cell_6t
Xbit_r109_c147 bl[147] br[147] wl[109] vdd gnd cell_6t
Xbit_r110_c147 bl[147] br[147] wl[110] vdd gnd cell_6t
Xbit_r111_c147 bl[147] br[147] wl[111] vdd gnd cell_6t
Xbit_r112_c147 bl[147] br[147] wl[112] vdd gnd cell_6t
Xbit_r113_c147 bl[147] br[147] wl[113] vdd gnd cell_6t
Xbit_r114_c147 bl[147] br[147] wl[114] vdd gnd cell_6t
Xbit_r115_c147 bl[147] br[147] wl[115] vdd gnd cell_6t
Xbit_r116_c147 bl[147] br[147] wl[116] vdd gnd cell_6t
Xbit_r117_c147 bl[147] br[147] wl[117] vdd gnd cell_6t
Xbit_r118_c147 bl[147] br[147] wl[118] vdd gnd cell_6t
Xbit_r119_c147 bl[147] br[147] wl[119] vdd gnd cell_6t
Xbit_r120_c147 bl[147] br[147] wl[120] vdd gnd cell_6t
Xbit_r121_c147 bl[147] br[147] wl[121] vdd gnd cell_6t
Xbit_r122_c147 bl[147] br[147] wl[122] vdd gnd cell_6t
Xbit_r123_c147 bl[147] br[147] wl[123] vdd gnd cell_6t
Xbit_r124_c147 bl[147] br[147] wl[124] vdd gnd cell_6t
Xbit_r125_c147 bl[147] br[147] wl[125] vdd gnd cell_6t
Xbit_r126_c147 bl[147] br[147] wl[126] vdd gnd cell_6t
Xbit_r127_c147 bl[147] br[147] wl[127] vdd gnd cell_6t
Xbit_r0_c148 bl[148] br[148] wl[0] vdd gnd cell_6t
Xbit_r1_c148 bl[148] br[148] wl[1] vdd gnd cell_6t
Xbit_r2_c148 bl[148] br[148] wl[2] vdd gnd cell_6t
Xbit_r3_c148 bl[148] br[148] wl[3] vdd gnd cell_6t
Xbit_r4_c148 bl[148] br[148] wl[4] vdd gnd cell_6t
Xbit_r5_c148 bl[148] br[148] wl[5] vdd gnd cell_6t
Xbit_r6_c148 bl[148] br[148] wl[6] vdd gnd cell_6t
Xbit_r7_c148 bl[148] br[148] wl[7] vdd gnd cell_6t
Xbit_r8_c148 bl[148] br[148] wl[8] vdd gnd cell_6t
Xbit_r9_c148 bl[148] br[148] wl[9] vdd gnd cell_6t
Xbit_r10_c148 bl[148] br[148] wl[10] vdd gnd cell_6t
Xbit_r11_c148 bl[148] br[148] wl[11] vdd gnd cell_6t
Xbit_r12_c148 bl[148] br[148] wl[12] vdd gnd cell_6t
Xbit_r13_c148 bl[148] br[148] wl[13] vdd gnd cell_6t
Xbit_r14_c148 bl[148] br[148] wl[14] vdd gnd cell_6t
Xbit_r15_c148 bl[148] br[148] wl[15] vdd gnd cell_6t
Xbit_r16_c148 bl[148] br[148] wl[16] vdd gnd cell_6t
Xbit_r17_c148 bl[148] br[148] wl[17] vdd gnd cell_6t
Xbit_r18_c148 bl[148] br[148] wl[18] vdd gnd cell_6t
Xbit_r19_c148 bl[148] br[148] wl[19] vdd gnd cell_6t
Xbit_r20_c148 bl[148] br[148] wl[20] vdd gnd cell_6t
Xbit_r21_c148 bl[148] br[148] wl[21] vdd gnd cell_6t
Xbit_r22_c148 bl[148] br[148] wl[22] vdd gnd cell_6t
Xbit_r23_c148 bl[148] br[148] wl[23] vdd gnd cell_6t
Xbit_r24_c148 bl[148] br[148] wl[24] vdd gnd cell_6t
Xbit_r25_c148 bl[148] br[148] wl[25] vdd gnd cell_6t
Xbit_r26_c148 bl[148] br[148] wl[26] vdd gnd cell_6t
Xbit_r27_c148 bl[148] br[148] wl[27] vdd gnd cell_6t
Xbit_r28_c148 bl[148] br[148] wl[28] vdd gnd cell_6t
Xbit_r29_c148 bl[148] br[148] wl[29] vdd gnd cell_6t
Xbit_r30_c148 bl[148] br[148] wl[30] vdd gnd cell_6t
Xbit_r31_c148 bl[148] br[148] wl[31] vdd gnd cell_6t
Xbit_r32_c148 bl[148] br[148] wl[32] vdd gnd cell_6t
Xbit_r33_c148 bl[148] br[148] wl[33] vdd gnd cell_6t
Xbit_r34_c148 bl[148] br[148] wl[34] vdd gnd cell_6t
Xbit_r35_c148 bl[148] br[148] wl[35] vdd gnd cell_6t
Xbit_r36_c148 bl[148] br[148] wl[36] vdd gnd cell_6t
Xbit_r37_c148 bl[148] br[148] wl[37] vdd gnd cell_6t
Xbit_r38_c148 bl[148] br[148] wl[38] vdd gnd cell_6t
Xbit_r39_c148 bl[148] br[148] wl[39] vdd gnd cell_6t
Xbit_r40_c148 bl[148] br[148] wl[40] vdd gnd cell_6t
Xbit_r41_c148 bl[148] br[148] wl[41] vdd gnd cell_6t
Xbit_r42_c148 bl[148] br[148] wl[42] vdd gnd cell_6t
Xbit_r43_c148 bl[148] br[148] wl[43] vdd gnd cell_6t
Xbit_r44_c148 bl[148] br[148] wl[44] vdd gnd cell_6t
Xbit_r45_c148 bl[148] br[148] wl[45] vdd gnd cell_6t
Xbit_r46_c148 bl[148] br[148] wl[46] vdd gnd cell_6t
Xbit_r47_c148 bl[148] br[148] wl[47] vdd gnd cell_6t
Xbit_r48_c148 bl[148] br[148] wl[48] vdd gnd cell_6t
Xbit_r49_c148 bl[148] br[148] wl[49] vdd gnd cell_6t
Xbit_r50_c148 bl[148] br[148] wl[50] vdd gnd cell_6t
Xbit_r51_c148 bl[148] br[148] wl[51] vdd gnd cell_6t
Xbit_r52_c148 bl[148] br[148] wl[52] vdd gnd cell_6t
Xbit_r53_c148 bl[148] br[148] wl[53] vdd gnd cell_6t
Xbit_r54_c148 bl[148] br[148] wl[54] vdd gnd cell_6t
Xbit_r55_c148 bl[148] br[148] wl[55] vdd gnd cell_6t
Xbit_r56_c148 bl[148] br[148] wl[56] vdd gnd cell_6t
Xbit_r57_c148 bl[148] br[148] wl[57] vdd gnd cell_6t
Xbit_r58_c148 bl[148] br[148] wl[58] vdd gnd cell_6t
Xbit_r59_c148 bl[148] br[148] wl[59] vdd gnd cell_6t
Xbit_r60_c148 bl[148] br[148] wl[60] vdd gnd cell_6t
Xbit_r61_c148 bl[148] br[148] wl[61] vdd gnd cell_6t
Xbit_r62_c148 bl[148] br[148] wl[62] vdd gnd cell_6t
Xbit_r63_c148 bl[148] br[148] wl[63] vdd gnd cell_6t
Xbit_r64_c148 bl[148] br[148] wl[64] vdd gnd cell_6t
Xbit_r65_c148 bl[148] br[148] wl[65] vdd gnd cell_6t
Xbit_r66_c148 bl[148] br[148] wl[66] vdd gnd cell_6t
Xbit_r67_c148 bl[148] br[148] wl[67] vdd gnd cell_6t
Xbit_r68_c148 bl[148] br[148] wl[68] vdd gnd cell_6t
Xbit_r69_c148 bl[148] br[148] wl[69] vdd gnd cell_6t
Xbit_r70_c148 bl[148] br[148] wl[70] vdd gnd cell_6t
Xbit_r71_c148 bl[148] br[148] wl[71] vdd gnd cell_6t
Xbit_r72_c148 bl[148] br[148] wl[72] vdd gnd cell_6t
Xbit_r73_c148 bl[148] br[148] wl[73] vdd gnd cell_6t
Xbit_r74_c148 bl[148] br[148] wl[74] vdd gnd cell_6t
Xbit_r75_c148 bl[148] br[148] wl[75] vdd gnd cell_6t
Xbit_r76_c148 bl[148] br[148] wl[76] vdd gnd cell_6t
Xbit_r77_c148 bl[148] br[148] wl[77] vdd gnd cell_6t
Xbit_r78_c148 bl[148] br[148] wl[78] vdd gnd cell_6t
Xbit_r79_c148 bl[148] br[148] wl[79] vdd gnd cell_6t
Xbit_r80_c148 bl[148] br[148] wl[80] vdd gnd cell_6t
Xbit_r81_c148 bl[148] br[148] wl[81] vdd gnd cell_6t
Xbit_r82_c148 bl[148] br[148] wl[82] vdd gnd cell_6t
Xbit_r83_c148 bl[148] br[148] wl[83] vdd gnd cell_6t
Xbit_r84_c148 bl[148] br[148] wl[84] vdd gnd cell_6t
Xbit_r85_c148 bl[148] br[148] wl[85] vdd gnd cell_6t
Xbit_r86_c148 bl[148] br[148] wl[86] vdd gnd cell_6t
Xbit_r87_c148 bl[148] br[148] wl[87] vdd gnd cell_6t
Xbit_r88_c148 bl[148] br[148] wl[88] vdd gnd cell_6t
Xbit_r89_c148 bl[148] br[148] wl[89] vdd gnd cell_6t
Xbit_r90_c148 bl[148] br[148] wl[90] vdd gnd cell_6t
Xbit_r91_c148 bl[148] br[148] wl[91] vdd gnd cell_6t
Xbit_r92_c148 bl[148] br[148] wl[92] vdd gnd cell_6t
Xbit_r93_c148 bl[148] br[148] wl[93] vdd gnd cell_6t
Xbit_r94_c148 bl[148] br[148] wl[94] vdd gnd cell_6t
Xbit_r95_c148 bl[148] br[148] wl[95] vdd gnd cell_6t
Xbit_r96_c148 bl[148] br[148] wl[96] vdd gnd cell_6t
Xbit_r97_c148 bl[148] br[148] wl[97] vdd gnd cell_6t
Xbit_r98_c148 bl[148] br[148] wl[98] vdd gnd cell_6t
Xbit_r99_c148 bl[148] br[148] wl[99] vdd gnd cell_6t
Xbit_r100_c148 bl[148] br[148] wl[100] vdd gnd cell_6t
Xbit_r101_c148 bl[148] br[148] wl[101] vdd gnd cell_6t
Xbit_r102_c148 bl[148] br[148] wl[102] vdd gnd cell_6t
Xbit_r103_c148 bl[148] br[148] wl[103] vdd gnd cell_6t
Xbit_r104_c148 bl[148] br[148] wl[104] vdd gnd cell_6t
Xbit_r105_c148 bl[148] br[148] wl[105] vdd gnd cell_6t
Xbit_r106_c148 bl[148] br[148] wl[106] vdd gnd cell_6t
Xbit_r107_c148 bl[148] br[148] wl[107] vdd gnd cell_6t
Xbit_r108_c148 bl[148] br[148] wl[108] vdd gnd cell_6t
Xbit_r109_c148 bl[148] br[148] wl[109] vdd gnd cell_6t
Xbit_r110_c148 bl[148] br[148] wl[110] vdd gnd cell_6t
Xbit_r111_c148 bl[148] br[148] wl[111] vdd gnd cell_6t
Xbit_r112_c148 bl[148] br[148] wl[112] vdd gnd cell_6t
Xbit_r113_c148 bl[148] br[148] wl[113] vdd gnd cell_6t
Xbit_r114_c148 bl[148] br[148] wl[114] vdd gnd cell_6t
Xbit_r115_c148 bl[148] br[148] wl[115] vdd gnd cell_6t
Xbit_r116_c148 bl[148] br[148] wl[116] vdd gnd cell_6t
Xbit_r117_c148 bl[148] br[148] wl[117] vdd gnd cell_6t
Xbit_r118_c148 bl[148] br[148] wl[118] vdd gnd cell_6t
Xbit_r119_c148 bl[148] br[148] wl[119] vdd gnd cell_6t
Xbit_r120_c148 bl[148] br[148] wl[120] vdd gnd cell_6t
Xbit_r121_c148 bl[148] br[148] wl[121] vdd gnd cell_6t
Xbit_r122_c148 bl[148] br[148] wl[122] vdd gnd cell_6t
Xbit_r123_c148 bl[148] br[148] wl[123] vdd gnd cell_6t
Xbit_r124_c148 bl[148] br[148] wl[124] vdd gnd cell_6t
Xbit_r125_c148 bl[148] br[148] wl[125] vdd gnd cell_6t
Xbit_r126_c148 bl[148] br[148] wl[126] vdd gnd cell_6t
Xbit_r127_c148 bl[148] br[148] wl[127] vdd gnd cell_6t
Xbit_r0_c149 bl[149] br[149] wl[0] vdd gnd cell_6t
Xbit_r1_c149 bl[149] br[149] wl[1] vdd gnd cell_6t
Xbit_r2_c149 bl[149] br[149] wl[2] vdd gnd cell_6t
Xbit_r3_c149 bl[149] br[149] wl[3] vdd gnd cell_6t
Xbit_r4_c149 bl[149] br[149] wl[4] vdd gnd cell_6t
Xbit_r5_c149 bl[149] br[149] wl[5] vdd gnd cell_6t
Xbit_r6_c149 bl[149] br[149] wl[6] vdd gnd cell_6t
Xbit_r7_c149 bl[149] br[149] wl[7] vdd gnd cell_6t
Xbit_r8_c149 bl[149] br[149] wl[8] vdd gnd cell_6t
Xbit_r9_c149 bl[149] br[149] wl[9] vdd gnd cell_6t
Xbit_r10_c149 bl[149] br[149] wl[10] vdd gnd cell_6t
Xbit_r11_c149 bl[149] br[149] wl[11] vdd gnd cell_6t
Xbit_r12_c149 bl[149] br[149] wl[12] vdd gnd cell_6t
Xbit_r13_c149 bl[149] br[149] wl[13] vdd gnd cell_6t
Xbit_r14_c149 bl[149] br[149] wl[14] vdd gnd cell_6t
Xbit_r15_c149 bl[149] br[149] wl[15] vdd gnd cell_6t
Xbit_r16_c149 bl[149] br[149] wl[16] vdd gnd cell_6t
Xbit_r17_c149 bl[149] br[149] wl[17] vdd gnd cell_6t
Xbit_r18_c149 bl[149] br[149] wl[18] vdd gnd cell_6t
Xbit_r19_c149 bl[149] br[149] wl[19] vdd gnd cell_6t
Xbit_r20_c149 bl[149] br[149] wl[20] vdd gnd cell_6t
Xbit_r21_c149 bl[149] br[149] wl[21] vdd gnd cell_6t
Xbit_r22_c149 bl[149] br[149] wl[22] vdd gnd cell_6t
Xbit_r23_c149 bl[149] br[149] wl[23] vdd gnd cell_6t
Xbit_r24_c149 bl[149] br[149] wl[24] vdd gnd cell_6t
Xbit_r25_c149 bl[149] br[149] wl[25] vdd gnd cell_6t
Xbit_r26_c149 bl[149] br[149] wl[26] vdd gnd cell_6t
Xbit_r27_c149 bl[149] br[149] wl[27] vdd gnd cell_6t
Xbit_r28_c149 bl[149] br[149] wl[28] vdd gnd cell_6t
Xbit_r29_c149 bl[149] br[149] wl[29] vdd gnd cell_6t
Xbit_r30_c149 bl[149] br[149] wl[30] vdd gnd cell_6t
Xbit_r31_c149 bl[149] br[149] wl[31] vdd gnd cell_6t
Xbit_r32_c149 bl[149] br[149] wl[32] vdd gnd cell_6t
Xbit_r33_c149 bl[149] br[149] wl[33] vdd gnd cell_6t
Xbit_r34_c149 bl[149] br[149] wl[34] vdd gnd cell_6t
Xbit_r35_c149 bl[149] br[149] wl[35] vdd gnd cell_6t
Xbit_r36_c149 bl[149] br[149] wl[36] vdd gnd cell_6t
Xbit_r37_c149 bl[149] br[149] wl[37] vdd gnd cell_6t
Xbit_r38_c149 bl[149] br[149] wl[38] vdd gnd cell_6t
Xbit_r39_c149 bl[149] br[149] wl[39] vdd gnd cell_6t
Xbit_r40_c149 bl[149] br[149] wl[40] vdd gnd cell_6t
Xbit_r41_c149 bl[149] br[149] wl[41] vdd gnd cell_6t
Xbit_r42_c149 bl[149] br[149] wl[42] vdd gnd cell_6t
Xbit_r43_c149 bl[149] br[149] wl[43] vdd gnd cell_6t
Xbit_r44_c149 bl[149] br[149] wl[44] vdd gnd cell_6t
Xbit_r45_c149 bl[149] br[149] wl[45] vdd gnd cell_6t
Xbit_r46_c149 bl[149] br[149] wl[46] vdd gnd cell_6t
Xbit_r47_c149 bl[149] br[149] wl[47] vdd gnd cell_6t
Xbit_r48_c149 bl[149] br[149] wl[48] vdd gnd cell_6t
Xbit_r49_c149 bl[149] br[149] wl[49] vdd gnd cell_6t
Xbit_r50_c149 bl[149] br[149] wl[50] vdd gnd cell_6t
Xbit_r51_c149 bl[149] br[149] wl[51] vdd gnd cell_6t
Xbit_r52_c149 bl[149] br[149] wl[52] vdd gnd cell_6t
Xbit_r53_c149 bl[149] br[149] wl[53] vdd gnd cell_6t
Xbit_r54_c149 bl[149] br[149] wl[54] vdd gnd cell_6t
Xbit_r55_c149 bl[149] br[149] wl[55] vdd gnd cell_6t
Xbit_r56_c149 bl[149] br[149] wl[56] vdd gnd cell_6t
Xbit_r57_c149 bl[149] br[149] wl[57] vdd gnd cell_6t
Xbit_r58_c149 bl[149] br[149] wl[58] vdd gnd cell_6t
Xbit_r59_c149 bl[149] br[149] wl[59] vdd gnd cell_6t
Xbit_r60_c149 bl[149] br[149] wl[60] vdd gnd cell_6t
Xbit_r61_c149 bl[149] br[149] wl[61] vdd gnd cell_6t
Xbit_r62_c149 bl[149] br[149] wl[62] vdd gnd cell_6t
Xbit_r63_c149 bl[149] br[149] wl[63] vdd gnd cell_6t
Xbit_r64_c149 bl[149] br[149] wl[64] vdd gnd cell_6t
Xbit_r65_c149 bl[149] br[149] wl[65] vdd gnd cell_6t
Xbit_r66_c149 bl[149] br[149] wl[66] vdd gnd cell_6t
Xbit_r67_c149 bl[149] br[149] wl[67] vdd gnd cell_6t
Xbit_r68_c149 bl[149] br[149] wl[68] vdd gnd cell_6t
Xbit_r69_c149 bl[149] br[149] wl[69] vdd gnd cell_6t
Xbit_r70_c149 bl[149] br[149] wl[70] vdd gnd cell_6t
Xbit_r71_c149 bl[149] br[149] wl[71] vdd gnd cell_6t
Xbit_r72_c149 bl[149] br[149] wl[72] vdd gnd cell_6t
Xbit_r73_c149 bl[149] br[149] wl[73] vdd gnd cell_6t
Xbit_r74_c149 bl[149] br[149] wl[74] vdd gnd cell_6t
Xbit_r75_c149 bl[149] br[149] wl[75] vdd gnd cell_6t
Xbit_r76_c149 bl[149] br[149] wl[76] vdd gnd cell_6t
Xbit_r77_c149 bl[149] br[149] wl[77] vdd gnd cell_6t
Xbit_r78_c149 bl[149] br[149] wl[78] vdd gnd cell_6t
Xbit_r79_c149 bl[149] br[149] wl[79] vdd gnd cell_6t
Xbit_r80_c149 bl[149] br[149] wl[80] vdd gnd cell_6t
Xbit_r81_c149 bl[149] br[149] wl[81] vdd gnd cell_6t
Xbit_r82_c149 bl[149] br[149] wl[82] vdd gnd cell_6t
Xbit_r83_c149 bl[149] br[149] wl[83] vdd gnd cell_6t
Xbit_r84_c149 bl[149] br[149] wl[84] vdd gnd cell_6t
Xbit_r85_c149 bl[149] br[149] wl[85] vdd gnd cell_6t
Xbit_r86_c149 bl[149] br[149] wl[86] vdd gnd cell_6t
Xbit_r87_c149 bl[149] br[149] wl[87] vdd gnd cell_6t
Xbit_r88_c149 bl[149] br[149] wl[88] vdd gnd cell_6t
Xbit_r89_c149 bl[149] br[149] wl[89] vdd gnd cell_6t
Xbit_r90_c149 bl[149] br[149] wl[90] vdd gnd cell_6t
Xbit_r91_c149 bl[149] br[149] wl[91] vdd gnd cell_6t
Xbit_r92_c149 bl[149] br[149] wl[92] vdd gnd cell_6t
Xbit_r93_c149 bl[149] br[149] wl[93] vdd gnd cell_6t
Xbit_r94_c149 bl[149] br[149] wl[94] vdd gnd cell_6t
Xbit_r95_c149 bl[149] br[149] wl[95] vdd gnd cell_6t
Xbit_r96_c149 bl[149] br[149] wl[96] vdd gnd cell_6t
Xbit_r97_c149 bl[149] br[149] wl[97] vdd gnd cell_6t
Xbit_r98_c149 bl[149] br[149] wl[98] vdd gnd cell_6t
Xbit_r99_c149 bl[149] br[149] wl[99] vdd gnd cell_6t
Xbit_r100_c149 bl[149] br[149] wl[100] vdd gnd cell_6t
Xbit_r101_c149 bl[149] br[149] wl[101] vdd gnd cell_6t
Xbit_r102_c149 bl[149] br[149] wl[102] vdd gnd cell_6t
Xbit_r103_c149 bl[149] br[149] wl[103] vdd gnd cell_6t
Xbit_r104_c149 bl[149] br[149] wl[104] vdd gnd cell_6t
Xbit_r105_c149 bl[149] br[149] wl[105] vdd gnd cell_6t
Xbit_r106_c149 bl[149] br[149] wl[106] vdd gnd cell_6t
Xbit_r107_c149 bl[149] br[149] wl[107] vdd gnd cell_6t
Xbit_r108_c149 bl[149] br[149] wl[108] vdd gnd cell_6t
Xbit_r109_c149 bl[149] br[149] wl[109] vdd gnd cell_6t
Xbit_r110_c149 bl[149] br[149] wl[110] vdd gnd cell_6t
Xbit_r111_c149 bl[149] br[149] wl[111] vdd gnd cell_6t
Xbit_r112_c149 bl[149] br[149] wl[112] vdd gnd cell_6t
Xbit_r113_c149 bl[149] br[149] wl[113] vdd gnd cell_6t
Xbit_r114_c149 bl[149] br[149] wl[114] vdd gnd cell_6t
Xbit_r115_c149 bl[149] br[149] wl[115] vdd gnd cell_6t
Xbit_r116_c149 bl[149] br[149] wl[116] vdd gnd cell_6t
Xbit_r117_c149 bl[149] br[149] wl[117] vdd gnd cell_6t
Xbit_r118_c149 bl[149] br[149] wl[118] vdd gnd cell_6t
Xbit_r119_c149 bl[149] br[149] wl[119] vdd gnd cell_6t
Xbit_r120_c149 bl[149] br[149] wl[120] vdd gnd cell_6t
Xbit_r121_c149 bl[149] br[149] wl[121] vdd gnd cell_6t
Xbit_r122_c149 bl[149] br[149] wl[122] vdd gnd cell_6t
Xbit_r123_c149 bl[149] br[149] wl[123] vdd gnd cell_6t
Xbit_r124_c149 bl[149] br[149] wl[124] vdd gnd cell_6t
Xbit_r125_c149 bl[149] br[149] wl[125] vdd gnd cell_6t
Xbit_r126_c149 bl[149] br[149] wl[126] vdd gnd cell_6t
Xbit_r127_c149 bl[149] br[149] wl[127] vdd gnd cell_6t
Xbit_r0_c150 bl[150] br[150] wl[0] vdd gnd cell_6t
Xbit_r1_c150 bl[150] br[150] wl[1] vdd gnd cell_6t
Xbit_r2_c150 bl[150] br[150] wl[2] vdd gnd cell_6t
Xbit_r3_c150 bl[150] br[150] wl[3] vdd gnd cell_6t
Xbit_r4_c150 bl[150] br[150] wl[4] vdd gnd cell_6t
Xbit_r5_c150 bl[150] br[150] wl[5] vdd gnd cell_6t
Xbit_r6_c150 bl[150] br[150] wl[6] vdd gnd cell_6t
Xbit_r7_c150 bl[150] br[150] wl[7] vdd gnd cell_6t
Xbit_r8_c150 bl[150] br[150] wl[8] vdd gnd cell_6t
Xbit_r9_c150 bl[150] br[150] wl[9] vdd gnd cell_6t
Xbit_r10_c150 bl[150] br[150] wl[10] vdd gnd cell_6t
Xbit_r11_c150 bl[150] br[150] wl[11] vdd gnd cell_6t
Xbit_r12_c150 bl[150] br[150] wl[12] vdd gnd cell_6t
Xbit_r13_c150 bl[150] br[150] wl[13] vdd gnd cell_6t
Xbit_r14_c150 bl[150] br[150] wl[14] vdd gnd cell_6t
Xbit_r15_c150 bl[150] br[150] wl[15] vdd gnd cell_6t
Xbit_r16_c150 bl[150] br[150] wl[16] vdd gnd cell_6t
Xbit_r17_c150 bl[150] br[150] wl[17] vdd gnd cell_6t
Xbit_r18_c150 bl[150] br[150] wl[18] vdd gnd cell_6t
Xbit_r19_c150 bl[150] br[150] wl[19] vdd gnd cell_6t
Xbit_r20_c150 bl[150] br[150] wl[20] vdd gnd cell_6t
Xbit_r21_c150 bl[150] br[150] wl[21] vdd gnd cell_6t
Xbit_r22_c150 bl[150] br[150] wl[22] vdd gnd cell_6t
Xbit_r23_c150 bl[150] br[150] wl[23] vdd gnd cell_6t
Xbit_r24_c150 bl[150] br[150] wl[24] vdd gnd cell_6t
Xbit_r25_c150 bl[150] br[150] wl[25] vdd gnd cell_6t
Xbit_r26_c150 bl[150] br[150] wl[26] vdd gnd cell_6t
Xbit_r27_c150 bl[150] br[150] wl[27] vdd gnd cell_6t
Xbit_r28_c150 bl[150] br[150] wl[28] vdd gnd cell_6t
Xbit_r29_c150 bl[150] br[150] wl[29] vdd gnd cell_6t
Xbit_r30_c150 bl[150] br[150] wl[30] vdd gnd cell_6t
Xbit_r31_c150 bl[150] br[150] wl[31] vdd gnd cell_6t
Xbit_r32_c150 bl[150] br[150] wl[32] vdd gnd cell_6t
Xbit_r33_c150 bl[150] br[150] wl[33] vdd gnd cell_6t
Xbit_r34_c150 bl[150] br[150] wl[34] vdd gnd cell_6t
Xbit_r35_c150 bl[150] br[150] wl[35] vdd gnd cell_6t
Xbit_r36_c150 bl[150] br[150] wl[36] vdd gnd cell_6t
Xbit_r37_c150 bl[150] br[150] wl[37] vdd gnd cell_6t
Xbit_r38_c150 bl[150] br[150] wl[38] vdd gnd cell_6t
Xbit_r39_c150 bl[150] br[150] wl[39] vdd gnd cell_6t
Xbit_r40_c150 bl[150] br[150] wl[40] vdd gnd cell_6t
Xbit_r41_c150 bl[150] br[150] wl[41] vdd gnd cell_6t
Xbit_r42_c150 bl[150] br[150] wl[42] vdd gnd cell_6t
Xbit_r43_c150 bl[150] br[150] wl[43] vdd gnd cell_6t
Xbit_r44_c150 bl[150] br[150] wl[44] vdd gnd cell_6t
Xbit_r45_c150 bl[150] br[150] wl[45] vdd gnd cell_6t
Xbit_r46_c150 bl[150] br[150] wl[46] vdd gnd cell_6t
Xbit_r47_c150 bl[150] br[150] wl[47] vdd gnd cell_6t
Xbit_r48_c150 bl[150] br[150] wl[48] vdd gnd cell_6t
Xbit_r49_c150 bl[150] br[150] wl[49] vdd gnd cell_6t
Xbit_r50_c150 bl[150] br[150] wl[50] vdd gnd cell_6t
Xbit_r51_c150 bl[150] br[150] wl[51] vdd gnd cell_6t
Xbit_r52_c150 bl[150] br[150] wl[52] vdd gnd cell_6t
Xbit_r53_c150 bl[150] br[150] wl[53] vdd gnd cell_6t
Xbit_r54_c150 bl[150] br[150] wl[54] vdd gnd cell_6t
Xbit_r55_c150 bl[150] br[150] wl[55] vdd gnd cell_6t
Xbit_r56_c150 bl[150] br[150] wl[56] vdd gnd cell_6t
Xbit_r57_c150 bl[150] br[150] wl[57] vdd gnd cell_6t
Xbit_r58_c150 bl[150] br[150] wl[58] vdd gnd cell_6t
Xbit_r59_c150 bl[150] br[150] wl[59] vdd gnd cell_6t
Xbit_r60_c150 bl[150] br[150] wl[60] vdd gnd cell_6t
Xbit_r61_c150 bl[150] br[150] wl[61] vdd gnd cell_6t
Xbit_r62_c150 bl[150] br[150] wl[62] vdd gnd cell_6t
Xbit_r63_c150 bl[150] br[150] wl[63] vdd gnd cell_6t
Xbit_r64_c150 bl[150] br[150] wl[64] vdd gnd cell_6t
Xbit_r65_c150 bl[150] br[150] wl[65] vdd gnd cell_6t
Xbit_r66_c150 bl[150] br[150] wl[66] vdd gnd cell_6t
Xbit_r67_c150 bl[150] br[150] wl[67] vdd gnd cell_6t
Xbit_r68_c150 bl[150] br[150] wl[68] vdd gnd cell_6t
Xbit_r69_c150 bl[150] br[150] wl[69] vdd gnd cell_6t
Xbit_r70_c150 bl[150] br[150] wl[70] vdd gnd cell_6t
Xbit_r71_c150 bl[150] br[150] wl[71] vdd gnd cell_6t
Xbit_r72_c150 bl[150] br[150] wl[72] vdd gnd cell_6t
Xbit_r73_c150 bl[150] br[150] wl[73] vdd gnd cell_6t
Xbit_r74_c150 bl[150] br[150] wl[74] vdd gnd cell_6t
Xbit_r75_c150 bl[150] br[150] wl[75] vdd gnd cell_6t
Xbit_r76_c150 bl[150] br[150] wl[76] vdd gnd cell_6t
Xbit_r77_c150 bl[150] br[150] wl[77] vdd gnd cell_6t
Xbit_r78_c150 bl[150] br[150] wl[78] vdd gnd cell_6t
Xbit_r79_c150 bl[150] br[150] wl[79] vdd gnd cell_6t
Xbit_r80_c150 bl[150] br[150] wl[80] vdd gnd cell_6t
Xbit_r81_c150 bl[150] br[150] wl[81] vdd gnd cell_6t
Xbit_r82_c150 bl[150] br[150] wl[82] vdd gnd cell_6t
Xbit_r83_c150 bl[150] br[150] wl[83] vdd gnd cell_6t
Xbit_r84_c150 bl[150] br[150] wl[84] vdd gnd cell_6t
Xbit_r85_c150 bl[150] br[150] wl[85] vdd gnd cell_6t
Xbit_r86_c150 bl[150] br[150] wl[86] vdd gnd cell_6t
Xbit_r87_c150 bl[150] br[150] wl[87] vdd gnd cell_6t
Xbit_r88_c150 bl[150] br[150] wl[88] vdd gnd cell_6t
Xbit_r89_c150 bl[150] br[150] wl[89] vdd gnd cell_6t
Xbit_r90_c150 bl[150] br[150] wl[90] vdd gnd cell_6t
Xbit_r91_c150 bl[150] br[150] wl[91] vdd gnd cell_6t
Xbit_r92_c150 bl[150] br[150] wl[92] vdd gnd cell_6t
Xbit_r93_c150 bl[150] br[150] wl[93] vdd gnd cell_6t
Xbit_r94_c150 bl[150] br[150] wl[94] vdd gnd cell_6t
Xbit_r95_c150 bl[150] br[150] wl[95] vdd gnd cell_6t
Xbit_r96_c150 bl[150] br[150] wl[96] vdd gnd cell_6t
Xbit_r97_c150 bl[150] br[150] wl[97] vdd gnd cell_6t
Xbit_r98_c150 bl[150] br[150] wl[98] vdd gnd cell_6t
Xbit_r99_c150 bl[150] br[150] wl[99] vdd gnd cell_6t
Xbit_r100_c150 bl[150] br[150] wl[100] vdd gnd cell_6t
Xbit_r101_c150 bl[150] br[150] wl[101] vdd gnd cell_6t
Xbit_r102_c150 bl[150] br[150] wl[102] vdd gnd cell_6t
Xbit_r103_c150 bl[150] br[150] wl[103] vdd gnd cell_6t
Xbit_r104_c150 bl[150] br[150] wl[104] vdd gnd cell_6t
Xbit_r105_c150 bl[150] br[150] wl[105] vdd gnd cell_6t
Xbit_r106_c150 bl[150] br[150] wl[106] vdd gnd cell_6t
Xbit_r107_c150 bl[150] br[150] wl[107] vdd gnd cell_6t
Xbit_r108_c150 bl[150] br[150] wl[108] vdd gnd cell_6t
Xbit_r109_c150 bl[150] br[150] wl[109] vdd gnd cell_6t
Xbit_r110_c150 bl[150] br[150] wl[110] vdd gnd cell_6t
Xbit_r111_c150 bl[150] br[150] wl[111] vdd gnd cell_6t
Xbit_r112_c150 bl[150] br[150] wl[112] vdd gnd cell_6t
Xbit_r113_c150 bl[150] br[150] wl[113] vdd gnd cell_6t
Xbit_r114_c150 bl[150] br[150] wl[114] vdd gnd cell_6t
Xbit_r115_c150 bl[150] br[150] wl[115] vdd gnd cell_6t
Xbit_r116_c150 bl[150] br[150] wl[116] vdd gnd cell_6t
Xbit_r117_c150 bl[150] br[150] wl[117] vdd gnd cell_6t
Xbit_r118_c150 bl[150] br[150] wl[118] vdd gnd cell_6t
Xbit_r119_c150 bl[150] br[150] wl[119] vdd gnd cell_6t
Xbit_r120_c150 bl[150] br[150] wl[120] vdd gnd cell_6t
Xbit_r121_c150 bl[150] br[150] wl[121] vdd gnd cell_6t
Xbit_r122_c150 bl[150] br[150] wl[122] vdd gnd cell_6t
Xbit_r123_c150 bl[150] br[150] wl[123] vdd gnd cell_6t
Xbit_r124_c150 bl[150] br[150] wl[124] vdd gnd cell_6t
Xbit_r125_c150 bl[150] br[150] wl[125] vdd gnd cell_6t
Xbit_r126_c150 bl[150] br[150] wl[126] vdd gnd cell_6t
Xbit_r127_c150 bl[150] br[150] wl[127] vdd gnd cell_6t
Xbit_r0_c151 bl[151] br[151] wl[0] vdd gnd cell_6t
Xbit_r1_c151 bl[151] br[151] wl[1] vdd gnd cell_6t
Xbit_r2_c151 bl[151] br[151] wl[2] vdd gnd cell_6t
Xbit_r3_c151 bl[151] br[151] wl[3] vdd gnd cell_6t
Xbit_r4_c151 bl[151] br[151] wl[4] vdd gnd cell_6t
Xbit_r5_c151 bl[151] br[151] wl[5] vdd gnd cell_6t
Xbit_r6_c151 bl[151] br[151] wl[6] vdd gnd cell_6t
Xbit_r7_c151 bl[151] br[151] wl[7] vdd gnd cell_6t
Xbit_r8_c151 bl[151] br[151] wl[8] vdd gnd cell_6t
Xbit_r9_c151 bl[151] br[151] wl[9] vdd gnd cell_6t
Xbit_r10_c151 bl[151] br[151] wl[10] vdd gnd cell_6t
Xbit_r11_c151 bl[151] br[151] wl[11] vdd gnd cell_6t
Xbit_r12_c151 bl[151] br[151] wl[12] vdd gnd cell_6t
Xbit_r13_c151 bl[151] br[151] wl[13] vdd gnd cell_6t
Xbit_r14_c151 bl[151] br[151] wl[14] vdd gnd cell_6t
Xbit_r15_c151 bl[151] br[151] wl[15] vdd gnd cell_6t
Xbit_r16_c151 bl[151] br[151] wl[16] vdd gnd cell_6t
Xbit_r17_c151 bl[151] br[151] wl[17] vdd gnd cell_6t
Xbit_r18_c151 bl[151] br[151] wl[18] vdd gnd cell_6t
Xbit_r19_c151 bl[151] br[151] wl[19] vdd gnd cell_6t
Xbit_r20_c151 bl[151] br[151] wl[20] vdd gnd cell_6t
Xbit_r21_c151 bl[151] br[151] wl[21] vdd gnd cell_6t
Xbit_r22_c151 bl[151] br[151] wl[22] vdd gnd cell_6t
Xbit_r23_c151 bl[151] br[151] wl[23] vdd gnd cell_6t
Xbit_r24_c151 bl[151] br[151] wl[24] vdd gnd cell_6t
Xbit_r25_c151 bl[151] br[151] wl[25] vdd gnd cell_6t
Xbit_r26_c151 bl[151] br[151] wl[26] vdd gnd cell_6t
Xbit_r27_c151 bl[151] br[151] wl[27] vdd gnd cell_6t
Xbit_r28_c151 bl[151] br[151] wl[28] vdd gnd cell_6t
Xbit_r29_c151 bl[151] br[151] wl[29] vdd gnd cell_6t
Xbit_r30_c151 bl[151] br[151] wl[30] vdd gnd cell_6t
Xbit_r31_c151 bl[151] br[151] wl[31] vdd gnd cell_6t
Xbit_r32_c151 bl[151] br[151] wl[32] vdd gnd cell_6t
Xbit_r33_c151 bl[151] br[151] wl[33] vdd gnd cell_6t
Xbit_r34_c151 bl[151] br[151] wl[34] vdd gnd cell_6t
Xbit_r35_c151 bl[151] br[151] wl[35] vdd gnd cell_6t
Xbit_r36_c151 bl[151] br[151] wl[36] vdd gnd cell_6t
Xbit_r37_c151 bl[151] br[151] wl[37] vdd gnd cell_6t
Xbit_r38_c151 bl[151] br[151] wl[38] vdd gnd cell_6t
Xbit_r39_c151 bl[151] br[151] wl[39] vdd gnd cell_6t
Xbit_r40_c151 bl[151] br[151] wl[40] vdd gnd cell_6t
Xbit_r41_c151 bl[151] br[151] wl[41] vdd gnd cell_6t
Xbit_r42_c151 bl[151] br[151] wl[42] vdd gnd cell_6t
Xbit_r43_c151 bl[151] br[151] wl[43] vdd gnd cell_6t
Xbit_r44_c151 bl[151] br[151] wl[44] vdd gnd cell_6t
Xbit_r45_c151 bl[151] br[151] wl[45] vdd gnd cell_6t
Xbit_r46_c151 bl[151] br[151] wl[46] vdd gnd cell_6t
Xbit_r47_c151 bl[151] br[151] wl[47] vdd gnd cell_6t
Xbit_r48_c151 bl[151] br[151] wl[48] vdd gnd cell_6t
Xbit_r49_c151 bl[151] br[151] wl[49] vdd gnd cell_6t
Xbit_r50_c151 bl[151] br[151] wl[50] vdd gnd cell_6t
Xbit_r51_c151 bl[151] br[151] wl[51] vdd gnd cell_6t
Xbit_r52_c151 bl[151] br[151] wl[52] vdd gnd cell_6t
Xbit_r53_c151 bl[151] br[151] wl[53] vdd gnd cell_6t
Xbit_r54_c151 bl[151] br[151] wl[54] vdd gnd cell_6t
Xbit_r55_c151 bl[151] br[151] wl[55] vdd gnd cell_6t
Xbit_r56_c151 bl[151] br[151] wl[56] vdd gnd cell_6t
Xbit_r57_c151 bl[151] br[151] wl[57] vdd gnd cell_6t
Xbit_r58_c151 bl[151] br[151] wl[58] vdd gnd cell_6t
Xbit_r59_c151 bl[151] br[151] wl[59] vdd gnd cell_6t
Xbit_r60_c151 bl[151] br[151] wl[60] vdd gnd cell_6t
Xbit_r61_c151 bl[151] br[151] wl[61] vdd gnd cell_6t
Xbit_r62_c151 bl[151] br[151] wl[62] vdd gnd cell_6t
Xbit_r63_c151 bl[151] br[151] wl[63] vdd gnd cell_6t
Xbit_r64_c151 bl[151] br[151] wl[64] vdd gnd cell_6t
Xbit_r65_c151 bl[151] br[151] wl[65] vdd gnd cell_6t
Xbit_r66_c151 bl[151] br[151] wl[66] vdd gnd cell_6t
Xbit_r67_c151 bl[151] br[151] wl[67] vdd gnd cell_6t
Xbit_r68_c151 bl[151] br[151] wl[68] vdd gnd cell_6t
Xbit_r69_c151 bl[151] br[151] wl[69] vdd gnd cell_6t
Xbit_r70_c151 bl[151] br[151] wl[70] vdd gnd cell_6t
Xbit_r71_c151 bl[151] br[151] wl[71] vdd gnd cell_6t
Xbit_r72_c151 bl[151] br[151] wl[72] vdd gnd cell_6t
Xbit_r73_c151 bl[151] br[151] wl[73] vdd gnd cell_6t
Xbit_r74_c151 bl[151] br[151] wl[74] vdd gnd cell_6t
Xbit_r75_c151 bl[151] br[151] wl[75] vdd gnd cell_6t
Xbit_r76_c151 bl[151] br[151] wl[76] vdd gnd cell_6t
Xbit_r77_c151 bl[151] br[151] wl[77] vdd gnd cell_6t
Xbit_r78_c151 bl[151] br[151] wl[78] vdd gnd cell_6t
Xbit_r79_c151 bl[151] br[151] wl[79] vdd gnd cell_6t
Xbit_r80_c151 bl[151] br[151] wl[80] vdd gnd cell_6t
Xbit_r81_c151 bl[151] br[151] wl[81] vdd gnd cell_6t
Xbit_r82_c151 bl[151] br[151] wl[82] vdd gnd cell_6t
Xbit_r83_c151 bl[151] br[151] wl[83] vdd gnd cell_6t
Xbit_r84_c151 bl[151] br[151] wl[84] vdd gnd cell_6t
Xbit_r85_c151 bl[151] br[151] wl[85] vdd gnd cell_6t
Xbit_r86_c151 bl[151] br[151] wl[86] vdd gnd cell_6t
Xbit_r87_c151 bl[151] br[151] wl[87] vdd gnd cell_6t
Xbit_r88_c151 bl[151] br[151] wl[88] vdd gnd cell_6t
Xbit_r89_c151 bl[151] br[151] wl[89] vdd gnd cell_6t
Xbit_r90_c151 bl[151] br[151] wl[90] vdd gnd cell_6t
Xbit_r91_c151 bl[151] br[151] wl[91] vdd gnd cell_6t
Xbit_r92_c151 bl[151] br[151] wl[92] vdd gnd cell_6t
Xbit_r93_c151 bl[151] br[151] wl[93] vdd gnd cell_6t
Xbit_r94_c151 bl[151] br[151] wl[94] vdd gnd cell_6t
Xbit_r95_c151 bl[151] br[151] wl[95] vdd gnd cell_6t
Xbit_r96_c151 bl[151] br[151] wl[96] vdd gnd cell_6t
Xbit_r97_c151 bl[151] br[151] wl[97] vdd gnd cell_6t
Xbit_r98_c151 bl[151] br[151] wl[98] vdd gnd cell_6t
Xbit_r99_c151 bl[151] br[151] wl[99] vdd gnd cell_6t
Xbit_r100_c151 bl[151] br[151] wl[100] vdd gnd cell_6t
Xbit_r101_c151 bl[151] br[151] wl[101] vdd gnd cell_6t
Xbit_r102_c151 bl[151] br[151] wl[102] vdd gnd cell_6t
Xbit_r103_c151 bl[151] br[151] wl[103] vdd gnd cell_6t
Xbit_r104_c151 bl[151] br[151] wl[104] vdd gnd cell_6t
Xbit_r105_c151 bl[151] br[151] wl[105] vdd gnd cell_6t
Xbit_r106_c151 bl[151] br[151] wl[106] vdd gnd cell_6t
Xbit_r107_c151 bl[151] br[151] wl[107] vdd gnd cell_6t
Xbit_r108_c151 bl[151] br[151] wl[108] vdd gnd cell_6t
Xbit_r109_c151 bl[151] br[151] wl[109] vdd gnd cell_6t
Xbit_r110_c151 bl[151] br[151] wl[110] vdd gnd cell_6t
Xbit_r111_c151 bl[151] br[151] wl[111] vdd gnd cell_6t
Xbit_r112_c151 bl[151] br[151] wl[112] vdd gnd cell_6t
Xbit_r113_c151 bl[151] br[151] wl[113] vdd gnd cell_6t
Xbit_r114_c151 bl[151] br[151] wl[114] vdd gnd cell_6t
Xbit_r115_c151 bl[151] br[151] wl[115] vdd gnd cell_6t
Xbit_r116_c151 bl[151] br[151] wl[116] vdd gnd cell_6t
Xbit_r117_c151 bl[151] br[151] wl[117] vdd gnd cell_6t
Xbit_r118_c151 bl[151] br[151] wl[118] vdd gnd cell_6t
Xbit_r119_c151 bl[151] br[151] wl[119] vdd gnd cell_6t
Xbit_r120_c151 bl[151] br[151] wl[120] vdd gnd cell_6t
Xbit_r121_c151 bl[151] br[151] wl[121] vdd gnd cell_6t
Xbit_r122_c151 bl[151] br[151] wl[122] vdd gnd cell_6t
Xbit_r123_c151 bl[151] br[151] wl[123] vdd gnd cell_6t
Xbit_r124_c151 bl[151] br[151] wl[124] vdd gnd cell_6t
Xbit_r125_c151 bl[151] br[151] wl[125] vdd gnd cell_6t
Xbit_r126_c151 bl[151] br[151] wl[126] vdd gnd cell_6t
Xbit_r127_c151 bl[151] br[151] wl[127] vdd gnd cell_6t
Xbit_r0_c152 bl[152] br[152] wl[0] vdd gnd cell_6t
Xbit_r1_c152 bl[152] br[152] wl[1] vdd gnd cell_6t
Xbit_r2_c152 bl[152] br[152] wl[2] vdd gnd cell_6t
Xbit_r3_c152 bl[152] br[152] wl[3] vdd gnd cell_6t
Xbit_r4_c152 bl[152] br[152] wl[4] vdd gnd cell_6t
Xbit_r5_c152 bl[152] br[152] wl[5] vdd gnd cell_6t
Xbit_r6_c152 bl[152] br[152] wl[6] vdd gnd cell_6t
Xbit_r7_c152 bl[152] br[152] wl[7] vdd gnd cell_6t
Xbit_r8_c152 bl[152] br[152] wl[8] vdd gnd cell_6t
Xbit_r9_c152 bl[152] br[152] wl[9] vdd gnd cell_6t
Xbit_r10_c152 bl[152] br[152] wl[10] vdd gnd cell_6t
Xbit_r11_c152 bl[152] br[152] wl[11] vdd gnd cell_6t
Xbit_r12_c152 bl[152] br[152] wl[12] vdd gnd cell_6t
Xbit_r13_c152 bl[152] br[152] wl[13] vdd gnd cell_6t
Xbit_r14_c152 bl[152] br[152] wl[14] vdd gnd cell_6t
Xbit_r15_c152 bl[152] br[152] wl[15] vdd gnd cell_6t
Xbit_r16_c152 bl[152] br[152] wl[16] vdd gnd cell_6t
Xbit_r17_c152 bl[152] br[152] wl[17] vdd gnd cell_6t
Xbit_r18_c152 bl[152] br[152] wl[18] vdd gnd cell_6t
Xbit_r19_c152 bl[152] br[152] wl[19] vdd gnd cell_6t
Xbit_r20_c152 bl[152] br[152] wl[20] vdd gnd cell_6t
Xbit_r21_c152 bl[152] br[152] wl[21] vdd gnd cell_6t
Xbit_r22_c152 bl[152] br[152] wl[22] vdd gnd cell_6t
Xbit_r23_c152 bl[152] br[152] wl[23] vdd gnd cell_6t
Xbit_r24_c152 bl[152] br[152] wl[24] vdd gnd cell_6t
Xbit_r25_c152 bl[152] br[152] wl[25] vdd gnd cell_6t
Xbit_r26_c152 bl[152] br[152] wl[26] vdd gnd cell_6t
Xbit_r27_c152 bl[152] br[152] wl[27] vdd gnd cell_6t
Xbit_r28_c152 bl[152] br[152] wl[28] vdd gnd cell_6t
Xbit_r29_c152 bl[152] br[152] wl[29] vdd gnd cell_6t
Xbit_r30_c152 bl[152] br[152] wl[30] vdd gnd cell_6t
Xbit_r31_c152 bl[152] br[152] wl[31] vdd gnd cell_6t
Xbit_r32_c152 bl[152] br[152] wl[32] vdd gnd cell_6t
Xbit_r33_c152 bl[152] br[152] wl[33] vdd gnd cell_6t
Xbit_r34_c152 bl[152] br[152] wl[34] vdd gnd cell_6t
Xbit_r35_c152 bl[152] br[152] wl[35] vdd gnd cell_6t
Xbit_r36_c152 bl[152] br[152] wl[36] vdd gnd cell_6t
Xbit_r37_c152 bl[152] br[152] wl[37] vdd gnd cell_6t
Xbit_r38_c152 bl[152] br[152] wl[38] vdd gnd cell_6t
Xbit_r39_c152 bl[152] br[152] wl[39] vdd gnd cell_6t
Xbit_r40_c152 bl[152] br[152] wl[40] vdd gnd cell_6t
Xbit_r41_c152 bl[152] br[152] wl[41] vdd gnd cell_6t
Xbit_r42_c152 bl[152] br[152] wl[42] vdd gnd cell_6t
Xbit_r43_c152 bl[152] br[152] wl[43] vdd gnd cell_6t
Xbit_r44_c152 bl[152] br[152] wl[44] vdd gnd cell_6t
Xbit_r45_c152 bl[152] br[152] wl[45] vdd gnd cell_6t
Xbit_r46_c152 bl[152] br[152] wl[46] vdd gnd cell_6t
Xbit_r47_c152 bl[152] br[152] wl[47] vdd gnd cell_6t
Xbit_r48_c152 bl[152] br[152] wl[48] vdd gnd cell_6t
Xbit_r49_c152 bl[152] br[152] wl[49] vdd gnd cell_6t
Xbit_r50_c152 bl[152] br[152] wl[50] vdd gnd cell_6t
Xbit_r51_c152 bl[152] br[152] wl[51] vdd gnd cell_6t
Xbit_r52_c152 bl[152] br[152] wl[52] vdd gnd cell_6t
Xbit_r53_c152 bl[152] br[152] wl[53] vdd gnd cell_6t
Xbit_r54_c152 bl[152] br[152] wl[54] vdd gnd cell_6t
Xbit_r55_c152 bl[152] br[152] wl[55] vdd gnd cell_6t
Xbit_r56_c152 bl[152] br[152] wl[56] vdd gnd cell_6t
Xbit_r57_c152 bl[152] br[152] wl[57] vdd gnd cell_6t
Xbit_r58_c152 bl[152] br[152] wl[58] vdd gnd cell_6t
Xbit_r59_c152 bl[152] br[152] wl[59] vdd gnd cell_6t
Xbit_r60_c152 bl[152] br[152] wl[60] vdd gnd cell_6t
Xbit_r61_c152 bl[152] br[152] wl[61] vdd gnd cell_6t
Xbit_r62_c152 bl[152] br[152] wl[62] vdd gnd cell_6t
Xbit_r63_c152 bl[152] br[152] wl[63] vdd gnd cell_6t
Xbit_r64_c152 bl[152] br[152] wl[64] vdd gnd cell_6t
Xbit_r65_c152 bl[152] br[152] wl[65] vdd gnd cell_6t
Xbit_r66_c152 bl[152] br[152] wl[66] vdd gnd cell_6t
Xbit_r67_c152 bl[152] br[152] wl[67] vdd gnd cell_6t
Xbit_r68_c152 bl[152] br[152] wl[68] vdd gnd cell_6t
Xbit_r69_c152 bl[152] br[152] wl[69] vdd gnd cell_6t
Xbit_r70_c152 bl[152] br[152] wl[70] vdd gnd cell_6t
Xbit_r71_c152 bl[152] br[152] wl[71] vdd gnd cell_6t
Xbit_r72_c152 bl[152] br[152] wl[72] vdd gnd cell_6t
Xbit_r73_c152 bl[152] br[152] wl[73] vdd gnd cell_6t
Xbit_r74_c152 bl[152] br[152] wl[74] vdd gnd cell_6t
Xbit_r75_c152 bl[152] br[152] wl[75] vdd gnd cell_6t
Xbit_r76_c152 bl[152] br[152] wl[76] vdd gnd cell_6t
Xbit_r77_c152 bl[152] br[152] wl[77] vdd gnd cell_6t
Xbit_r78_c152 bl[152] br[152] wl[78] vdd gnd cell_6t
Xbit_r79_c152 bl[152] br[152] wl[79] vdd gnd cell_6t
Xbit_r80_c152 bl[152] br[152] wl[80] vdd gnd cell_6t
Xbit_r81_c152 bl[152] br[152] wl[81] vdd gnd cell_6t
Xbit_r82_c152 bl[152] br[152] wl[82] vdd gnd cell_6t
Xbit_r83_c152 bl[152] br[152] wl[83] vdd gnd cell_6t
Xbit_r84_c152 bl[152] br[152] wl[84] vdd gnd cell_6t
Xbit_r85_c152 bl[152] br[152] wl[85] vdd gnd cell_6t
Xbit_r86_c152 bl[152] br[152] wl[86] vdd gnd cell_6t
Xbit_r87_c152 bl[152] br[152] wl[87] vdd gnd cell_6t
Xbit_r88_c152 bl[152] br[152] wl[88] vdd gnd cell_6t
Xbit_r89_c152 bl[152] br[152] wl[89] vdd gnd cell_6t
Xbit_r90_c152 bl[152] br[152] wl[90] vdd gnd cell_6t
Xbit_r91_c152 bl[152] br[152] wl[91] vdd gnd cell_6t
Xbit_r92_c152 bl[152] br[152] wl[92] vdd gnd cell_6t
Xbit_r93_c152 bl[152] br[152] wl[93] vdd gnd cell_6t
Xbit_r94_c152 bl[152] br[152] wl[94] vdd gnd cell_6t
Xbit_r95_c152 bl[152] br[152] wl[95] vdd gnd cell_6t
Xbit_r96_c152 bl[152] br[152] wl[96] vdd gnd cell_6t
Xbit_r97_c152 bl[152] br[152] wl[97] vdd gnd cell_6t
Xbit_r98_c152 bl[152] br[152] wl[98] vdd gnd cell_6t
Xbit_r99_c152 bl[152] br[152] wl[99] vdd gnd cell_6t
Xbit_r100_c152 bl[152] br[152] wl[100] vdd gnd cell_6t
Xbit_r101_c152 bl[152] br[152] wl[101] vdd gnd cell_6t
Xbit_r102_c152 bl[152] br[152] wl[102] vdd gnd cell_6t
Xbit_r103_c152 bl[152] br[152] wl[103] vdd gnd cell_6t
Xbit_r104_c152 bl[152] br[152] wl[104] vdd gnd cell_6t
Xbit_r105_c152 bl[152] br[152] wl[105] vdd gnd cell_6t
Xbit_r106_c152 bl[152] br[152] wl[106] vdd gnd cell_6t
Xbit_r107_c152 bl[152] br[152] wl[107] vdd gnd cell_6t
Xbit_r108_c152 bl[152] br[152] wl[108] vdd gnd cell_6t
Xbit_r109_c152 bl[152] br[152] wl[109] vdd gnd cell_6t
Xbit_r110_c152 bl[152] br[152] wl[110] vdd gnd cell_6t
Xbit_r111_c152 bl[152] br[152] wl[111] vdd gnd cell_6t
Xbit_r112_c152 bl[152] br[152] wl[112] vdd gnd cell_6t
Xbit_r113_c152 bl[152] br[152] wl[113] vdd gnd cell_6t
Xbit_r114_c152 bl[152] br[152] wl[114] vdd gnd cell_6t
Xbit_r115_c152 bl[152] br[152] wl[115] vdd gnd cell_6t
Xbit_r116_c152 bl[152] br[152] wl[116] vdd gnd cell_6t
Xbit_r117_c152 bl[152] br[152] wl[117] vdd gnd cell_6t
Xbit_r118_c152 bl[152] br[152] wl[118] vdd gnd cell_6t
Xbit_r119_c152 bl[152] br[152] wl[119] vdd gnd cell_6t
Xbit_r120_c152 bl[152] br[152] wl[120] vdd gnd cell_6t
Xbit_r121_c152 bl[152] br[152] wl[121] vdd gnd cell_6t
Xbit_r122_c152 bl[152] br[152] wl[122] vdd gnd cell_6t
Xbit_r123_c152 bl[152] br[152] wl[123] vdd gnd cell_6t
Xbit_r124_c152 bl[152] br[152] wl[124] vdd gnd cell_6t
Xbit_r125_c152 bl[152] br[152] wl[125] vdd gnd cell_6t
Xbit_r126_c152 bl[152] br[152] wl[126] vdd gnd cell_6t
Xbit_r127_c152 bl[152] br[152] wl[127] vdd gnd cell_6t
Xbit_r0_c153 bl[153] br[153] wl[0] vdd gnd cell_6t
Xbit_r1_c153 bl[153] br[153] wl[1] vdd gnd cell_6t
Xbit_r2_c153 bl[153] br[153] wl[2] vdd gnd cell_6t
Xbit_r3_c153 bl[153] br[153] wl[3] vdd gnd cell_6t
Xbit_r4_c153 bl[153] br[153] wl[4] vdd gnd cell_6t
Xbit_r5_c153 bl[153] br[153] wl[5] vdd gnd cell_6t
Xbit_r6_c153 bl[153] br[153] wl[6] vdd gnd cell_6t
Xbit_r7_c153 bl[153] br[153] wl[7] vdd gnd cell_6t
Xbit_r8_c153 bl[153] br[153] wl[8] vdd gnd cell_6t
Xbit_r9_c153 bl[153] br[153] wl[9] vdd gnd cell_6t
Xbit_r10_c153 bl[153] br[153] wl[10] vdd gnd cell_6t
Xbit_r11_c153 bl[153] br[153] wl[11] vdd gnd cell_6t
Xbit_r12_c153 bl[153] br[153] wl[12] vdd gnd cell_6t
Xbit_r13_c153 bl[153] br[153] wl[13] vdd gnd cell_6t
Xbit_r14_c153 bl[153] br[153] wl[14] vdd gnd cell_6t
Xbit_r15_c153 bl[153] br[153] wl[15] vdd gnd cell_6t
Xbit_r16_c153 bl[153] br[153] wl[16] vdd gnd cell_6t
Xbit_r17_c153 bl[153] br[153] wl[17] vdd gnd cell_6t
Xbit_r18_c153 bl[153] br[153] wl[18] vdd gnd cell_6t
Xbit_r19_c153 bl[153] br[153] wl[19] vdd gnd cell_6t
Xbit_r20_c153 bl[153] br[153] wl[20] vdd gnd cell_6t
Xbit_r21_c153 bl[153] br[153] wl[21] vdd gnd cell_6t
Xbit_r22_c153 bl[153] br[153] wl[22] vdd gnd cell_6t
Xbit_r23_c153 bl[153] br[153] wl[23] vdd gnd cell_6t
Xbit_r24_c153 bl[153] br[153] wl[24] vdd gnd cell_6t
Xbit_r25_c153 bl[153] br[153] wl[25] vdd gnd cell_6t
Xbit_r26_c153 bl[153] br[153] wl[26] vdd gnd cell_6t
Xbit_r27_c153 bl[153] br[153] wl[27] vdd gnd cell_6t
Xbit_r28_c153 bl[153] br[153] wl[28] vdd gnd cell_6t
Xbit_r29_c153 bl[153] br[153] wl[29] vdd gnd cell_6t
Xbit_r30_c153 bl[153] br[153] wl[30] vdd gnd cell_6t
Xbit_r31_c153 bl[153] br[153] wl[31] vdd gnd cell_6t
Xbit_r32_c153 bl[153] br[153] wl[32] vdd gnd cell_6t
Xbit_r33_c153 bl[153] br[153] wl[33] vdd gnd cell_6t
Xbit_r34_c153 bl[153] br[153] wl[34] vdd gnd cell_6t
Xbit_r35_c153 bl[153] br[153] wl[35] vdd gnd cell_6t
Xbit_r36_c153 bl[153] br[153] wl[36] vdd gnd cell_6t
Xbit_r37_c153 bl[153] br[153] wl[37] vdd gnd cell_6t
Xbit_r38_c153 bl[153] br[153] wl[38] vdd gnd cell_6t
Xbit_r39_c153 bl[153] br[153] wl[39] vdd gnd cell_6t
Xbit_r40_c153 bl[153] br[153] wl[40] vdd gnd cell_6t
Xbit_r41_c153 bl[153] br[153] wl[41] vdd gnd cell_6t
Xbit_r42_c153 bl[153] br[153] wl[42] vdd gnd cell_6t
Xbit_r43_c153 bl[153] br[153] wl[43] vdd gnd cell_6t
Xbit_r44_c153 bl[153] br[153] wl[44] vdd gnd cell_6t
Xbit_r45_c153 bl[153] br[153] wl[45] vdd gnd cell_6t
Xbit_r46_c153 bl[153] br[153] wl[46] vdd gnd cell_6t
Xbit_r47_c153 bl[153] br[153] wl[47] vdd gnd cell_6t
Xbit_r48_c153 bl[153] br[153] wl[48] vdd gnd cell_6t
Xbit_r49_c153 bl[153] br[153] wl[49] vdd gnd cell_6t
Xbit_r50_c153 bl[153] br[153] wl[50] vdd gnd cell_6t
Xbit_r51_c153 bl[153] br[153] wl[51] vdd gnd cell_6t
Xbit_r52_c153 bl[153] br[153] wl[52] vdd gnd cell_6t
Xbit_r53_c153 bl[153] br[153] wl[53] vdd gnd cell_6t
Xbit_r54_c153 bl[153] br[153] wl[54] vdd gnd cell_6t
Xbit_r55_c153 bl[153] br[153] wl[55] vdd gnd cell_6t
Xbit_r56_c153 bl[153] br[153] wl[56] vdd gnd cell_6t
Xbit_r57_c153 bl[153] br[153] wl[57] vdd gnd cell_6t
Xbit_r58_c153 bl[153] br[153] wl[58] vdd gnd cell_6t
Xbit_r59_c153 bl[153] br[153] wl[59] vdd gnd cell_6t
Xbit_r60_c153 bl[153] br[153] wl[60] vdd gnd cell_6t
Xbit_r61_c153 bl[153] br[153] wl[61] vdd gnd cell_6t
Xbit_r62_c153 bl[153] br[153] wl[62] vdd gnd cell_6t
Xbit_r63_c153 bl[153] br[153] wl[63] vdd gnd cell_6t
Xbit_r64_c153 bl[153] br[153] wl[64] vdd gnd cell_6t
Xbit_r65_c153 bl[153] br[153] wl[65] vdd gnd cell_6t
Xbit_r66_c153 bl[153] br[153] wl[66] vdd gnd cell_6t
Xbit_r67_c153 bl[153] br[153] wl[67] vdd gnd cell_6t
Xbit_r68_c153 bl[153] br[153] wl[68] vdd gnd cell_6t
Xbit_r69_c153 bl[153] br[153] wl[69] vdd gnd cell_6t
Xbit_r70_c153 bl[153] br[153] wl[70] vdd gnd cell_6t
Xbit_r71_c153 bl[153] br[153] wl[71] vdd gnd cell_6t
Xbit_r72_c153 bl[153] br[153] wl[72] vdd gnd cell_6t
Xbit_r73_c153 bl[153] br[153] wl[73] vdd gnd cell_6t
Xbit_r74_c153 bl[153] br[153] wl[74] vdd gnd cell_6t
Xbit_r75_c153 bl[153] br[153] wl[75] vdd gnd cell_6t
Xbit_r76_c153 bl[153] br[153] wl[76] vdd gnd cell_6t
Xbit_r77_c153 bl[153] br[153] wl[77] vdd gnd cell_6t
Xbit_r78_c153 bl[153] br[153] wl[78] vdd gnd cell_6t
Xbit_r79_c153 bl[153] br[153] wl[79] vdd gnd cell_6t
Xbit_r80_c153 bl[153] br[153] wl[80] vdd gnd cell_6t
Xbit_r81_c153 bl[153] br[153] wl[81] vdd gnd cell_6t
Xbit_r82_c153 bl[153] br[153] wl[82] vdd gnd cell_6t
Xbit_r83_c153 bl[153] br[153] wl[83] vdd gnd cell_6t
Xbit_r84_c153 bl[153] br[153] wl[84] vdd gnd cell_6t
Xbit_r85_c153 bl[153] br[153] wl[85] vdd gnd cell_6t
Xbit_r86_c153 bl[153] br[153] wl[86] vdd gnd cell_6t
Xbit_r87_c153 bl[153] br[153] wl[87] vdd gnd cell_6t
Xbit_r88_c153 bl[153] br[153] wl[88] vdd gnd cell_6t
Xbit_r89_c153 bl[153] br[153] wl[89] vdd gnd cell_6t
Xbit_r90_c153 bl[153] br[153] wl[90] vdd gnd cell_6t
Xbit_r91_c153 bl[153] br[153] wl[91] vdd gnd cell_6t
Xbit_r92_c153 bl[153] br[153] wl[92] vdd gnd cell_6t
Xbit_r93_c153 bl[153] br[153] wl[93] vdd gnd cell_6t
Xbit_r94_c153 bl[153] br[153] wl[94] vdd gnd cell_6t
Xbit_r95_c153 bl[153] br[153] wl[95] vdd gnd cell_6t
Xbit_r96_c153 bl[153] br[153] wl[96] vdd gnd cell_6t
Xbit_r97_c153 bl[153] br[153] wl[97] vdd gnd cell_6t
Xbit_r98_c153 bl[153] br[153] wl[98] vdd gnd cell_6t
Xbit_r99_c153 bl[153] br[153] wl[99] vdd gnd cell_6t
Xbit_r100_c153 bl[153] br[153] wl[100] vdd gnd cell_6t
Xbit_r101_c153 bl[153] br[153] wl[101] vdd gnd cell_6t
Xbit_r102_c153 bl[153] br[153] wl[102] vdd gnd cell_6t
Xbit_r103_c153 bl[153] br[153] wl[103] vdd gnd cell_6t
Xbit_r104_c153 bl[153] br[153] wl[104] vdd gnd cell_6t
Xbit_r105_c153 bl[153] br[153] wl[105] vdd gnd cell_6t
Xbit_r106_c153 bl[153] br[153] wl[106] vdd gnd cell_6t
Xbit_r107_c153 bl[153] br[153] wl[107] vdd gnd cell_6t
Xbit_r108_c153 bl[153] br[153] wl[108] vdd gnd cell_6t
Xbit_r109_c153 bl[153] br[153] wl[109] vdd gnd cell_6t
Xbit_r110_c153 bl[153] br[153] wl[110] vdd gnd cell_6t
Xbit_r111_c153 bl[153] br[153] wl[111] vdd gnd cell_6t
Xbit_r112_c153 bl[153] br[153] wl[112] vdd gnd cell_6t
Xbit_r113_c153 bl[153] br[153] wl[113] vdd gnd cell_6t
Xbit_r114_c153 bl[153] br[153] wl[114] vdd gnd cell_6t
Xbit_r115_c153 bl[153] br[153] wl[115] vdd gnd cell_6t
Xbit_r116_c153 bl[153] br[153] wl[116] vdd gnd cell_6t
Xbit_r117_c153 bl[153] br[153] wl[117] vdd gnd cell_6t
Xbit_r118_c153 bl[153] br[153] wl[118] vdd gnd cell_6t
Xbit_r119_c153 bl[153] br[153] wl[119] vdd gnd cell_6t
Xbit_r120_c153 bl[153] br[153] wl[120] vdd gnd cell_6t
Xbit_r121_c153 bl[153] br[153] wl[121] vdd gnd cell_6t
Xbit_r122_c153 bl[153] br[153] wl[122] vdd gnd cell_6t
Xbit_r123_c153 bl[153] br[153] wl[123] vdd gnd cell_6t
Xbit_r124_c153 bl[153] br[153] wl[124] vdd gnd cell_6t
Xbit_r125_c153 bl[153] br[153] wl[125] vdd gnd cell_6t
Xbit_r126_c153 bl[153] br[153] wl[126] vdd gnd cell_6t
Xbit_r127_c153 bl[153] br[153] wl[127] vdd gnd cell_6t
Xbit_r0_c154 bl[154] br[154] wl[0] vdd gnd cell_6t
Xbit_r1_c154 bl[154] br[154] wl[1] vdd gnd cell_6t
Xbit_r2_c154 bl[154] br[154] wl[2] vdd gnd cell_6t
Xbit_r3_c154 bl[154] br[154] wl[3] vdd gnd cell_6t
Xbit_r4_c154 bl[154] br[154] wl[4] vdd gnd cell_6t
Xbit_r5_c154 bl[154] br[154] wl[5] vdd gnd cell_6t
Xbit_r6_c154 bl[154] br[154] wl[6] vdd gnd cell_6t
Xbit_r7_c154 bl[154] br[154] wl[7] vdd gnd cell_6t
Xbit_r8_c154 bl[154] br[154] wl[8] vdd gnd cell_6t
Xbit_r9_c154 bl[154] br[154] wl[9] vdd gnd cell_6t
Xbit_r10_c154 bl[154] br[154] wl[10] vdd gnd cell_6t
Xbit_r11_c154 bl[154] br[154] wl[11] vdd gnd cell_6t
Xbit_r12_c154 bl[154] br[154] wl[12] vdd gnd cell_6t
Xbit_r13_c154 bl[154] br[154] wl[13] vdd gnd cell_6t
Xbit_r14_c154 bl[154] br[154] wl[14] vdd gnd cell_6t
Xbit_r15_c154 bl[154] br[154] wl[15] vdd gnd cell_6t
Xbit_r16_c154 bl[154] br[154] wl[16] vdd gnd cell_6t
Xbit_r17_c154 bl[154] br[154] wl[17] vdd gnd cell_6t
Xbit_r18_c154 bl[154] br[154] wl[18] vdd gnd cell_6t
Xbit_r19_c154 bl[154] br[154] wl[19] vdd gnd cell_6t
Xbit_r20_c154 bl[154] br[154] wl[20] vdd gnd cell_6t
Xbit_r21_c154 bl[154] br[154] wl[21] vdd gnd cell_6t
Xbit_r22_c154 bl[154] br[154] wl[22] vdd gnd cell_6t
Xbit_r23_c154 bl[154] br[154] wl[23] vdd gnd cell_6t
Xbit_r24_c154 bl[154] br[154] wl[24] vdd gnd cell_6t
Xbit_r25_c154 bl[154] br[154] wl[25] vdd gnd cell_6t
Xbit_r26_c154 bl[154] br[154] wl[26] vdd gnd cell_6t
Xbit_r27_c154 bl[154] br[154] wl[27] vdd gnd cell_6t
Xbit_r28_c154 bl[154] br[154] wl[28] vdd gnd cell_6t
Xbit_r29_c154 bl[154] br[154] wl[29] vdd gnd cell_6t
Xbit_r30_c154 bl[154] br[154] wl[30] vdd gnd cell_6t
Xbit_r31_c154 bl[154] br[154] wl[31] vdd gnd cell_6t
Xbit_r32_c154 bl[154] br[154] wl[32] vdd gnd cell_6t
Xbit_r33_c154 bl[154] br[154] wl[33] vdd gnd cell_6t
Xbit_r34_c154 bl[154] br[154] wl[34] vdd gnd cell_6t
Xbit_r35_c154 bl[154] br[154] wl[35] vdd gnd cell_6t
Xbit_r36_c154 bl[154] br[154] wl[36] vdd gnd cell_6t
Xbit_r37_c154 bl[154] br[154] wl[37] vdd gnd cell_6t
Xbit_r38_c154 bl[154] br[154] wl[38] vdd gnd cell_6t
Xbit_r39_c154 bl[154] br[154] wl[39] vdd gnd cell_6t
Xbit_r40_c154 bl[154] br[154] wl[40] vdd gnd cell_6t
Xbit_r41_c154 bl[154] br[154] wl[41] vdd gnd cell_6t
Xbit_r42_c154 bl[154] br[154] wl[42] vdd gnd cell_6t
Xbit_r43_c154 bl[154] br[154] wl[43] vdd gnd cell_6t
Xbit_r44_c154 bl[154] br[154] wl[44] vdd gnd cell_6t
Xbit_r45_c154 bl[154] br[154] wl[45] vdd gnd cell_6t
Xbit_r46_c154 bl[154] br[154] wl[46] vdd gnd cell_6t
Xbit_r47_c154 bl[154] br[154] wl[47] vdd gnd cell_6t
Xbit_r48_c154 bl[154] br[154] wl[48] vdd gnd cell_6t
Xbit_r49_c154 bl[154] br[154] wl[49] vdd gnd cell_6t
Xbit_r50_c154 bl[154] br[154] wl[50] vdd gnd cell_6t
Xbit_r51_c154 bl[154] br[154] wl[51] vdd gnd cell_6t
Xbit_r52_c154 bl[154] br[154] wl[52] vdd gnd cell_6t
Xbit_r53_c154 bl[154] br[154] wl[53] vdd gnd cell_6t
Xbit_r54_c154 bl[154] br[154] wl[54] vdd gnd cell_6t
Xbit_r55_c154 bl[154] br[154] wl[55] vdd gnd cell_6t
Xbit_r56_c154 bl[154] br[154] wl[56] vdd gnd cell_6t
Xbit_r57_c154 bl[154] br[154] wl[57] vdd gnd cell_6t
Xbit_r58_c154 bl[154] br[154] wl[58] vdd gnd cell_6t
Xbit_r59_c154 bl[154] br[154] wl[59] vdd gnd cell_6t
Xbit_r60_c154 bl[154] br[154] wl[60] vdd gnd cell_6t
Xbit_r61_c154 bl[154] br[154] wl[61] vdd gnd cell_6t
Xbit_r62_c154 bl[154] br[154] wl[62] vdd gnd cell_6t
Xbit_r63_c154 bl[154] br[154] wl[63] vdd gnd cell_6t
Xbit_r64_c154 bl[154] br[154] wl[64] vdd gnd cell_6t
Xbit_r65_c154 bl[154] br[154] wl[65] vdd gnd cell_6t
Xbit_r66_c154 bl[154] br[154] wl[66] vdd gnd cell_6t
Xbit_r67_c154 bl[154] br[154] wl[67] vdd gnd cell_6t
Xbit_r68_c154 bl[154] br[154] wl[68] vdd gnd cell_6t
Xbit_r69_c154 bl[154] br[154] wl[69] vdd gnd cell_6t
Xbit_r70_c154 bl[154] br[154] wl[70] vdd gnd cell_6t
Xbit_r71_c154 bl[154] br[154] wl[71] vdd gnd cell_6t
Xbit_r72_c154 bl[154] br[154] wl[72] vdd gnd cell_6t
Xbit_r73_c154 bl[154] br[154] wl[73] vdd gnd cell_6t
Xbit_r74_c154 bl[154] br[154] wl[74] vdd gnd cell_6t
Xbit_r75_c154 bl[154] br[154] wl[75] vdd gnd cell_6t
Xbit_r76_c154 bl[154] br[154] wl[76] vdd gnd cell_6t
Xbit_r77_c154 bl[154] br[154] wl[77] vdd gnd cell_6t
Xbit_r78_c154 bl[154] br[154] wl[78] vdd gnd cell_6t
Xbit_r79_c154 bl[154] br[154] wl[79] vdd gnd cell_6t
Xbit_r80_c154 bl[154] br[154] wl[80] vdd gnd cell_6t
Xbit_r81_c154 bl[154] br[154] wl[81] vdd gnd cell_6t
Xbit_r82_c154 bl[154] br[154] wl[82] vdd gnd cell_6t
Xbit_r83_c154 bl[154] br[154] wl[83] vdd gnd cell_6t
Xbit_r84_c154 bl[154] br[154] wl[84] vdd gnd cell_6t
Xbit_r85_c154 bl[154] br[154] wl[85] vdd gnd cell_6t
Xbit_r86_c154 bl[154] br[154] wl[86] vdd gnd cell_6t
Xbit_r87_c154 bl[154] br[154] wl[87] vdd gnd cell_6t
Xbit_r88_c154 bl[154] br[154] wl[88] vdd gnd cell_6t
Xbit_r89_c154 bl[154] br[154] wl[89] vdd gnd cell_6t
Xbit_r90_c154 bl[154] br[154] wl[90] vdd gnd cell_6t
Xbit_r91_c154 bl[154] br[154] wl[91] vdd gnd cell_6t
Xbit_r92_c154 bl[154] br[154] wl[92] vdd gnd cell_6t
Xbit_r93_c154 bl[154] br[154] wl[93] vdd gnd cell_6t
Xbit_r94_c154 bl[154] br[154] wl[94] vdd gnd cell_6t
Xbit_r95_c154 bl[154] br[154] wl[95] vdd gnd cell_6t
Xbit_r96_c154 bl[154] br[154] wl[96] vdd gnd cell_6t
Xbit_r97_c154 bl[154] br[154] wl[97] vdd gnd cell_6t
Xbit_r98_c154 bl[154] br[154] wl[98] vdd gnd cell_6t
Xbit_r99_c154 bl[154] br[154] wl[99] vdd gnd cell_6t
Xbit_r100_c154 bl[154] br[154] wl[100] vdd gnd cell_6t
Xbit_r101_c154 bl[154] br[154] wl[101] vdd gnd cell_6t
Xbit_r102_c154 bl[154] br[154] wl[102] vdd gnd cell_6t
Xbit_r103_c154 bl[154] br[154] wl[103] vdd gnd cell_6t
Xbit_r104_c154 bl[154] br[154] wl[104] vdd gnd cell_6t
Xbit_r105_c154 bl[154] br[154] wl[105] vdd gnd cell_6t
Xbit_r106_c154 bl[154] br[154] wl[106] vdd gnd cell_6t
Xbit_r107_c154 bl[154] br[154] wl[107] vdd gnd cell_6t
Xbit_r108_c154 bl[154] br[154] wl[108] vdd gnd cell_6t
Xbit_r109_c154 bl[154] br[154] wl[109] vdd gnd cell_6t
Xbit_r110_c154 bl[154] br[154] wl[110] vdd gnd cell_6t
Xbit_r111_c154 bl[154] br[154] wl[111] vdd gnd cell_6t
Xbit_r112_c154 bl[154] br[154] wl[112] vdd gnd cell_6t
Xbit_r113_c154 bl[154] br[154] wl[113] vdd gnd cell_6t
Xbit_r114_c154 bl[154] br[154] wl[114] vdd gnd cell_6t
Xbit_r115_c154 bl[154] br[154] wl[115] vdd gnd cell_6t
Xbit_r116_c154 bl[154] br[154] wl[116] vdd gnd cell_6t
Xbit_r117_c154 bl[154] br[154] wl[117] vdd gnd cell_6t
Xbit_r118_c154 bl[154] br[154] wl[118] vdd gnd cell_6t
Xbit_r119_c154 bl[154] br[154] wl[119] vdd gnd cell_6t
Xbit_r120_c154 bl[154] br[154] wl[120] vdd gnd cell_6t
Xbit_r121_c154 bl[154] br[154] wl[121] vdd gnd cell_6t
Xbit_r122_c154 bl[154] br[154] wl[122] vdd gnd cell_6t
Xbit_r123_c154 bl[154] br[154] wl[123] vdd gnd cell_6t
Xbit_r124_c154 bl[154] br[154] wl[124] vdd gnd cell_6t
Xbit_r125_c154 bl[154] br[154] wl[125] vdd gnd cell_6t
Xbit_r126_c154 bl[154] br[154] wl[126] vdd gnd cell_6t
Xbit_r127_c154 bl[154] br[154] wl[127] vdd gnd cell_6t
Xbit_r0_c155 bl[155] br[155] wl[0] vdd gnd cell_6t
Xbit_r1_c155 bl[155] br[155] wl[1] vdd gnd cell_6t
Xbit_r2_c155 bl[155] br[155] wl[2] vdd gnd cell_6t
Xbit_r3_c155 bl[155] br[155] wl[3] vdd gnd cell_6t
Xbit_r4_c155 bl[155] br[155] wl[4] vdd gnd cell_6t
Xbit_r5_c155 bl[155] br[155] wl[5] vdd gnd cell_6t
Xbit_r6_c155 bl[155] br[155] wl[6] vdd gnd cell_6t
Xbit_r7_c155 bl[155] br[155] wl[7] vdd gnd cell_6t
Xbit_r8_c155 bl[155] br[155] wl[8] vdd gnd cell_6t
Xbit_r9_c155 bl[155] br[155] wl[9] vdd gnd cell_6t
Xbit_r10_c155 bl[155] br[155] wl[10] vdd gnd cell_6t
Xbit_r11_c155 bl[155] br[155] wl[11] vdd gnd cell_6t
Xbit_r12_c155 bl[155] br[155] wl[12] vdd gnd cell_6t
Xbit_r13_c155 bl[155] br[155] wl[13] vdd gnd cell_6t
Xbit_r14_c155 bl[155] br[155] wl[14] vdd gnd cell_6t
Xbit_r15_c155 bl[155] br[155] wl[15] vdd gnd cell_6t
Xbit_r16_c155 bl[155] br[155] wl[16] vdd gnd cell_6t
Xbit_r17_c155 bl[155] br[155] wl[17] vdd gnd cell_6t
Xbit_r18_c155 bl[155] br[155] wl[18] vdd gnd cell_6t
Xbit_r19_c155 bl[155] br[155] wl[19] vdd gnd cell_6t
Xbit_r20_c155 bl[155] br[155] wl[20] vdd gnd cell_6t
Xbit_r21_c155 bl[155] br[155] wl[21] vdd gnd cell_6t
Xbit_r22_c155 bl[155] br[155] wl[22] vdd gnd cell_6t
Xbit_r23_c155 bl[155] br[155] wl[23] vdd gnd cell_6t
Xbit_r24_c155 bl[155] br[155] wl[24] vdd gnd cell_6t
Xbit_r25_c155 bl[155] br[155] wl[25] vdd gnd cell_6t
Xbit_r26_c155 bl[155] br[155] wl[26] vdd gnd cell_6t
Xbit_r27_c155 bl[155] br[155] wl[27] vdd gnd cell_6t
Xbit_r28_c155 bl[155] br[155] wl[28] vdd gnd cell_6t
Xbit_r29_c155 bl[155] br[155] wl[29] vdd gnd cell_6t
Xbit_r30_c155 bl[155] br[155] wl[30] vdd gnd cell_6t
Xbit_r31_c155 bl[155] br[155] wl[31] vdd gnd cell_6t
Xbit_r32_c155 bl[155] br[155] wl[32] vdd gnd cell_6t
Xbit_r33_c155 bl[155] br[155] wl[33] vdd gnd cell_6t
Xbit_r34_c155 bl[155] br[155] wl[34] vdd gnd cell_6t
Xbit_r35_c155 bl[155] br[155] wl[35] vdd gnd cell_6t
Xbit_r36_c155 bl[155] br[155] wl[36] vdd gnd cell_6t
Xbit_r37_c155 bl[155] br[155] wl[37] vdd gnd cell_6t
Xbit_r38_c155 bl[155] br[155] wl[38] vdd gnd cell_6t
Xbit_r39_c155 bl[155] br[155] wl[39] vdd gnd cell_6t
Xbit_r40_c155 bl[155] br[155] wl[40] vdd gnd cell_6t
Xbit_r41_c155 bl[155] br[155] wl[41] vdd gnd cell_6t
Xbit_r42_c155 bl[155] br[155] wl[42] vdd gnd cell_6t
Xbit_r43_c155 bl[155] br[155] wl[43] vdd gnd cell_6t
Xbit_r44_c155 bl[155] br[155] wl[44] vdd gnd cell_6t
Xbit_r45_c155 bl[155] br[155] wl[45] vdd gnd cell_6t
Xbit_r46_c155 bl[155] br[155] wl[46] vdd gnd cell_6t
Xbit_r47_c155 bl[155] br[155] wl[47] vdd gnd cell_6t
Xbit_r48_c155 bl[155] br[155] wl[48] vdd gnd cell_6t
Xbit_r49_c155 bl[155] br[155] wl[49] vdd gnd cell_6t
Xbit_r50_c155 bl[155] br[155] wl[50] vdd gnd cell_6t
Xbit_r51_c155 bl[155] br[155] wl[51] vdd gnd cell_6t
Xbit_r52_c155 bl[155] br[155] wl[52] vdd gnd cell_6t
Xbit_r53_c155 bl[155] br[155] wl[53] vdd gnd cell_6t
Xbit_r54_c155 bl[155] br[155] wl[54] vdd gnd cell_6t
Xbit_r55_c155 bl[155] br[155] wl[55] vdd gnd cell_6t
Xbit_r56_c155 bl[155] br[155] wl[56] vdd gnd cell_6t
Xbit_r57_c155 bl[155] br[155] wl[57] vdd gnd cell_6t
Xbit_r58_c155 bl[155] br[155] wl[58] vdd gnd cell_6t
Xbit_r59_c155 bl[155] br[155] wl[59] vdd gnd cell_6t
Xbit_r60_c155 bl[155] br[155] wl[60] vdd gnd cell_6t
Xbit_r61_c155 bl[155] br[155] wl[61] vdd gnd cell_6t
Xbit_r62_c155 bl[155] br[155] wl[62] vdd gnd cell_6t
Xbit_r63_c155 bl[155] br[155] wl[63] vdd gnd cell_6t
Xbit_r64_c155 bl[155] br[155] wl[64] vdd gnd cell_6t
Xbit_r65_c155 bl[155] br[155] wl[65] vdd gnd cell_6t
Xbit_r66_c155 bl[155] br[155] wl[66] vdd gnd cell_6t
Xbit_r67_c155 bl[155] br[155] wl[67] vdd gnd cell_6t
Xbit_r68_c155 bl[155] br[155] wl[68] vdd gnd cell_6t
Xbit_r69_c155 bl[155] br[155] wl[69] vdd gnd cell_6t
Xbit_r70_c155 bl[155] br[155] wl[70] vdd gnd cell_6t
Xbit_r71_c155 bl[155] br[155] wl[71] vdd gnd cell_6t
Xbit_r72_c155 bl[155] br[155] wl[72] vdd gnd cell_6t
Xbit_r73_c155 bl[155] br[155] wl[73] vdd gnd cell_6t
Xbit_r74_c155 bl[155] br[155] wl[74] vdd gnd cell_6t
Xbit_r75_c155 bl[155] br[155] wl[75] vdd gnd cell_6t
Xbit_r76_c155 bl[155] br[155] wl[76] vdd gnd cell_6t
Xbit_r77_c155 bl[155] br[155] wl[77] vdd gnd cell_6t
Xbit_r78_c155 bl[155] br[155] wl[78] vdd gnd cell_6t
Xbit_r79_c155 bl[155] br[155] wl[79] vdd gnd cell_6t
Xbit_r80_c155 bl[155] br[155] wl[80] vdd gnd cell_6t
Xbit_r81_c155 bl[155] br[155] wl[81] vdd gnd cell_6t
Xbit_r82_c155 bl[155] br[155] wl[82] vdd gnd cell_6t
Xbit_r83_c155 bl[155] br[155] wl[83] vdd gnd cell_6t
Xbit_r84_c155 bl[155] br[155] wl[84] vdd gnd cell_6t
Xbit_r85_c155 bl[155] br[155] wl[85] vdd gnd cell_6t
Xbit_r86_c155 bl[155] br[155] wl[86] vdd gnd cell_6t
Xbit_r87_c155 bl[155] br[155] wl[87] vdd gnd cell_6t
Xbit_r88_c155 bl[155] br[155] wl[88] vdd gnd cell_6t
Xbit_r89_c155 bl[155] br[155] wl[89] vdd gnd cell_6t
Xbit_r90_c155 bl[155] br[155] wl[90] vdd gnd cell_6t
Xbit_r91_c155 bl[155] br[155] wl[91] vdd gnd cell_6t
Xbit_r92_c155 bl[155] br[155] wl[92] vdd gnd cell_6t
Xbit_r93_c155 bl[155] br[155] wl[93] vdd gnd cell_6t
Xbit_r94_c155 bl[155] br[155] wl[94] vdd gnd cell_6t
Xbit_r95_c155 bl[155] br[155] wl[95] vdd gnd cell_6t
Xbit_r96_c155 bl[155] br[155] wl[96] vdd gnd cell_6t
Xbit_r97_c155 bl[155] br[155] wl[97] vdd gnd cell_6t
Xbit_r98_c155 bl[155] br[155] wl[98] vdd gnd cell_6t
Xbit_r99_c155 bl[155] br[155] wl[99] vdd gnd cell_6t
Xbit_r100_c155 bl[155] br[155] wl[100] vdd gnd cell_6t
Xbit_r101_c155 bl[155] br[155] wl[101] vdd gnd cell_6t
Xbit_r102_c155 bl[155] br[155] wl[102] vdd gnd cell_6t
Xbit_r103_c155 bl[155] br[155] wl[103] vdd gnd cell_6t
Xbit_r104_c155 bl[155] br[155] wl[104] vdd gnd cell_6t
Xbit_r105_c155 bl[155] br[155] wl[105] vdd gnd cell_6t
Xbit_r106_c155 bl[155] br[155] wl[106] vdd gnd cell_6t
Xbit_r107_c155 bl[155] br[155] wl[107] vdd gnd cell_6t
Xbit_r108_c155 bl[155] br[155] wl[108] vdd gnd cell_6t
Xbit_r109_c155 bl[155] br[155] wl[109] vdd gnd cell_6t
Xbit_r110_c155 bl[155] br[155] wl[110] vdd gnd cell_6t
Xbit_r111_c155 bl[155] br[155] wl[111] vdd gnd cell_6t
Xbit_r112_c155 bl[155] br[155] wl[112] vdd gnd cell_6t
Xbit_r113_c155 bl[155] br[155] wl[113] vdd gnd cell_6t
Xbit_r114_c155 bl[155] br[155] wl[114] vdd gnd cell_6t
Xbit_r115_c155 bl[155] br[155] wl[115] vdd gnd cell_6t
Xbit_r116_c155 bl[155] br[155] wl[116] vdd gnd cell_6t
Xbit_r117_c155 bl[155] br[155] wl[117] vdd gnd cell_6t
Xbit_r118_c155 bl[155] br[155] wl[118] vdd gnd cell_6t
Xbit_r119_c155 bl[155] br[155] wl[119] vdd gnd cell_6t
Xbit_r120_c155 bl[155] br[155] wl[120] vdd gnd cell_6t
Xbit_r121_c155 bl[155] br[155] wl[121] vdd gnd cell_6t
Xbit_r122_c155 bl[155] br[155] wl[122] vdd gnd cell_6t
Xbit_r123_c155 bl[155] br[155] wl[123] vdd gnd cell_6t
Xbit_r124_c155 bl[155] br[155] wl[124] vdd gnd cell_6t
Xbit_r125_c155 bl[155] br[155] wl[125] vdd gnd cell_6t
Xbit_r126_c155 bl[155] br[155] wl[126] vdd gnd cell_6t
Xbit_r127_c155 bl[155] br[155] wl[127] vdd gnd cell_6t
Xbit_r0_c156 bl[156] br[156] wl[0] vdd gnd cell_6t
Xbit_r1_c156 bl[156] br[156] wl[1] vdd gnd cell_6t
Xbit_r2_c156 bl[156] br[156] wl[2] vdd gnd cell_6t
Xbit_r3_c156 bl[156] br[156] wl[3] vdd gnd cell_6t
Xbit_r4_c156 bl[156] br[156] wl[4] vdd gnd cell_6t
Xbit_r5_c156 bl[156] br[156] wl[5] vdd gnd cell_6t
Xbit_r6_c156 bl[156] br[156] wl[6] vdd gnd cell_6t
Xbit_r7_c156 bl[156] br[156] wl[7] vdd gnd cell_6t
Xbit_r8_c156 bl[156] br[156] wl[8] vdd gnd cell_6t
Xbit_r9_c156 bl[156] br[156] wl[9] vdd gnd cell_6t
Xbit_r10_c156 bl[156] br[156] wl[10] vdd gnd cell_6t
Xbit_r11_c156 bl[156] br[156] wl[11] vdd gnd cell_6t
Xbit_r12_c156 bl[156] br[156] wl[12] vdd gnd cell_6t
Xbit_r13_c156 bl[156] br[156] wl[13] vdd gnd cell_6t
Xbit_r14_c156 bl[156] br[156] wl[14] vdd gnd cell_6t
Xbit_r15_c156 bl[156] br[156] wl[15] vdd gnd cell_6t
Xbit_r16_c156 bl[156] br[156] wl[16] vdd gnd cell_6t
Xbit_r17_c156 bl[156] br[156] wl[17] vdd gnd cell_6t
Xbit_r18_c156 bl[156] br[156] wl[18] vdd gnd cell_6t
Xbit_r19_c156 bl[156] br[156] wl[19] vdd gnd cell_6t
Xbit_r20_c156 bl[156] br[156] wl[20] vdd gnd cell_6t
Xbit_r21_c156 bl[156] br[156] wl[21] vdd gnd cell_6t
Xbit_r22_c156 bl[156] br[156] wl[22] vdd gnd cell_6t
Xbit_r23_c156 bl[156] br[156] wl[23] vdd gnd cell_6t
Xbit_r24_c156 bl[156] br[156] wl[24] vdd gnd cell_6t
Xbit_r25_c156 bl[156] br[156] wl[25] vdd gnd cell_6t
Xbit_r26_c156 bl[156] br[156] wl[26] vdd gnd cell_6t
Xbit_r27_c156 bl[156] br[156] wl[27] vdd gnd cell_6t
Xbit_r28_c156 bl[156] br[156] wl[28] vdd gnd cell_6t
Xbit_r29_c156 bl[156] br[156] wl[29] vdd gnd cell_6t
Xbit_r30_c156 bl[156] br[156] wl[30] vdd gnd cell_6t
Xbit_r31_c156 bl[156] br[156] wl[31] vdd gnd cell_6t
Xbit_r32_c156 bl[156] br[156] wl[32] vdd gnd cell_6t
Xbit_r33_c156 bl[156] br[156] wl[33] vdd gnd cell_6t
Xbit_r34_c156 bl[156] br[156] wl[34] vdd gnd cell_6t
Xbit_r35_c156 bl[156] br[156] wl[35] vdd gnd cell_6t
Xbit_r36_c156 bl[156] br[156] wl[36] vdd gnd cell_6t
Xbit_r37_c156 bl[156] br[156] wl[37] vdd gnd cell_6t
Xbit_r38_c156 bl[156] br[156] wl[38] vdd gnd cell_6t
Xbit_r39_c156 bl[156] br[156] wl[39] vdd gnd cell_6t
Xbit_r40_c156 bl[156] br[156] wl[40] vdd gnd cell_6t
Xbit_r41_c156 bl[156] br[156] wl[41] vdd gnd cell_6t
Xbit_r42_c156 bl[156] br[156] wl[42] vdd gnd cell_6t
Xbit_r43_c156 bl[156] br[156] wl[43] vdd gnd cell_6t
Xbit_r44_c156 bl[156] br[156] wl[44] vdd gnd cell_6t
Xbit_r45_c156 bl[156] br[156] wl[45] vdd gnd cell_6t
Xbit_r46_c156 bl[156] br[156] wl[46] vdd gnd cell_6t
Xbit_r47_c156 bl[156] br[156] wl[47] vdd gnd cell_6t
Xbit_r48_c156 bl[156] br[156] wl[48] vdd gnd cell_6t
Xbit_r49_c156 bl[156] br[156] wl[49] vdd gnd cell_6t
Xbit_r50_c156 bl[156] br[156] wl[50] vdd gnd cell_6t
Xbit_r51_c156 bl[156] br[156] wl[51] vdd gnd cell_6t
Xbit_r52_c156 bl[156] br[156] wl[52] vdd gnd cell_6t
Xbit_r53_c156 bl[156] br[156] wl[53] vdd gnd cell_6t
Xbit_r54_c156 bl[156] br[156] wl[54] vdd gnd cell_6t
Xbit_r55_c156 bl[156] br[156] wl[55] vdd gnd cell_6t
Xbit_r56_c156 bl[156] br[156] wl[56] vdd gnd cell_6t
Xbit_r57_c156 bl[156] br[156] wl[57] vdd gnd cell_6t
Xbit_r58_c156 bl[156] br[156] wl[58] vdd gnd cell_6t
Xbit_r59_c156 bl[156] br[156] wl[59] vdd gnd cell_6t
Xbit_r60_c156 bl[156] br[156] wl[60] vdd gnd cell_6t
Xbit_r61_c156 bl[156] br[156] wl[61] vdd gnd cell_6t
Xbit_r62_c156 bl[156] br[156] wl[62] vdd gnd cell_6t
Xbit_r63_c156 bl[156] br[156] wl[63] vdd gnd cell_6t
Xbit_r64_c156 bl[156] br[156] wl[64] vdd gnd cell_6t
Xbit_r65_c156 bl[156] br[156] wl[65] vdd gnd cell_6t
Xbit_r66_c156 bl[156] br[156] wl[66] vdd gnd cell_6t
Xbit_r67_c156 bl[156] br[156] wl[67] vdd gnd cell_6t
Xbit_r68_c156 bl[156] br[156] wl[68] vdd gnd cell_6t
Xbit_r69_c156 bl[156] br[156] wl[69] vdd gnd cell_6t
Xbit_r70_c156 bl[156] br[156] wl[70] vdd gnd cell_6t
Xbit_r71_c156 bl[156] br[156] wl[71] vdd gnd cell_6t
Xbit_r72_c156 bl[156] br[156] wl[72] vdd gnd cell_6t
Xbit_r73_c156 bl[156] br[156] wl[73] vdd gnd cell_6t
Xbit_r74_c156 bl[156] br[156] wl[74] vdd gnd cell_6t
Xbit_r75_c156 bl[156] br[156] wl[75] vdd gnd cell_6t
Xbit_r76_c156 bl[156] br[156] wl[76] vdd gnd cell_6t
Xbit_r77_c156 bl[156] br[156] wl[77] vdd gnd cell_6t
Xbit_r78_c156 bl[156] br[156] wl[78] vdd gnd cell_6t
Xbit_r79_c156 bl[156] br[156] wl[79] vdd gnd cell_6t
Xbit_r80_c156 bl[156] br[156] wl[80] vdd gnd cell_6t
Xbit_r81_c156 bl[156] br[156] wl[81] vdd gnd cell_6t
Xbit_r82_c156 bl[156] br[156] wl[82] vdd gnd cell_6t
Xbit_r83_c156 bl[156] br[156] wl[83] vdd gnd cell_6t
Xbit_r84_c156 bl[156] br[156] wl[84] vdd gnd cell_6t
Xbit_r85_c156 bl[156] br[156] wl[85] vdd gnd cell_6t
Xbit_r86_c156 bl[156] br[156] wl[86] vdd gnd cell_6t
Xbit_r87_c156 bl[156] br[156] wl[87] vdd gnd cell_6t
Xbit_r88_c156 bl[156] br[156] wl[88] vdd gnd cell_6t
Xbit_r89_c156 bl[156] br[156] wl[89] vdd gnd cell_6t
Xbit_r90_c156 bl[156] br[156] wl[90] vdd gnd cell_6t
Xbit_r91_c156 bl[156] br[156] wl[91] vdd gnd cell_6t
Xbit_r92_c156 bl[156] br[156] wl[92] vdd gnd cell_6t
Xbit_r93_c156 bl[156] br[156] wl[93] vdd gnd cell_6t
Xbit_r94_c156 bl[156] br[156] wl[94] vdd gnd cell_6t
Xbit_r95_c156 bl[156] br[156] wl[95] vdd gnd cell_6t
Xbit_r96_c156 bl[156] br[156] wl[96] vdd gnd cell_6t
Xbit_r97_c156 bl[156] br[156] wl[97] vdd gnd cell_6t
Xbit_r98_c156 bl[156] br[156] wl[98] vdd gnd cell_6t
Xbit_r99_c156 bl[156] br[156] wl[99] vdd gnd cell_6t
Xbit_r100_c156 bl[156] br[156] wl[100] vdd gnd cell_6t
Xbit_r101_c156 bl[156] br[156] wl[101] vdd gnd cell_6t
Xbit_r102_c156 bl[156] br[156] wl[102] vdd gnd cell_6t
Xbit_r103_c156 bl[156] br[156] wl[103] vdd gnd cell_6t
Xbit_r104_c156 bl[156] br[156] wl[104] vdd gnd cell_6t
Xbit_r105_c156 bl[156] br[156] wl[105] vdd gnd cell_6t
Xbit_r106_c156 bl[156] br[156] wl[106] vdd gnd cell_6t
Xbit_r107_c156 bl[156] br[156] wl[107] vdd gnd cell_6t
Xbit_r108_c156 bl[156] br[156] wl[108] vdd gnd cell_6t
Xbit_r109_c156 bl[156] br[156] wl[109] vdd gnd cell_6t
Xbit_r110_c156 bl[156] br[156] wl[110] vdd gnd cell_6t
Xbit_r111_c156 bl[156] br[156] wl[111] vdd gnd cell_6t
Xbit_r112_c156 bl[156] br[156] wl[112] vdd gnd cell_6t
Xbit_r113_c156 bl[156] br[156] wl[113] vdd gnd cell_6t
Xbit_r114_c156 bl[156] br[156] wl[114] vdd gnd cell_6t
Xbit_r115_c156 bl[156] br[156] wl[115] vdd gnd cell_6t
Xbit_r116_c156 bl[156] br[156] wl[116] vdd gnd cell_6t
Xbit_r117_c156 bl[156] br[156] wl[117] vdd gnd cell_6t
Xbit_r118_c156 bl[156] br[156] wl[118] vdd gnd cell_6t
Xbit_r119_c156 bl[156] br[156] wl[119] vdd gnd cell_6t
Xbit_r120_c156 bl[156] br[156] wl[120] vdd gnd cell_6t
Xbit_r121_c156 bl[156] br[156] wl[121] vdd gnd cell_6t
Xbit_r122_c156 bl[156] br[156] wl[122] vdd gnd cell_6t
Xbit_r123_c156 bl[156] br[156] wl[123] vdd gnd cell_6t
Xbit_r124_c156 bl[156] br[156] wl[124] vdd gnd cell_6t
Xbit_r125_c156 bl[156] br[156] wl[125] vdd gnd cell_6t
Xbit_r126_c156 bl[156] br[156] wl[126] vdd gnd cell_6t
Xbit_r127_c156 bl[156] br[156] wl[127] vdd gnd cell_6t
Xbit_r0_c157 bl[157] br[157] wl[0] vdd gnd cell_6t
Xbit_r1_c157 bl[157] br[157] wl[1] vdd gnd cell_6t
Xbit_r2_c157 bl[157] br[157] wl[2] vdd gnd cell_6t
Xbit_r3_c157 bl[157] br[157] wl[3] vdd gnd cell_6t
Xbit_r4_c157 bl[157] br[157] wl[4] vdd gnd cell_6t
Xbit_r5_c157 bl[157] br[157] wl[5] vdd gnd cell_6t
Xbit_r6_c157 bl[157] br[157] wl[6] vdd gnd cell_6t
Xbit_r7_c157 bl[157] br[157] wl[7] vdd gnd cell_6t
Xbit_r8_c157 bl[157] br[157] wl[8] vdd gnd cell_6t
Xbit_r9_c157 bl[157] br[157] wl[9] vdd gnd cell_6t
Xbit_r10_c157 bl[157] br[157] wl[10] vdd gnd cell_6t
Xbit_r11_c157 bl[157] br[157] wl[11] vdd gnd cell_6t
Xbit_r12_c157 bl[157] br[157] wl[12] vdd gnd cell_6t
Xbit_r13_c157 bl[157] br[157] wl[13] vdd gnd cell_6t
Xbit_r14_c157 bl[157] br[157] wl[14] vdd gnd cell_6t
Xbit_r15_c157 bl[157] br[157] wl[15] vdd gnd cell_6t
Xbit_r16_c157 bl[157] br[157] wl[16] vdd gnd cell_6t
Xbit_r17_c157 bl[157] br[157] wl[17] vdd gnd cell_6t
Xbit_r18_c157 bl[157] br[157] wl[18] vdd gnd cell_6t
Xbit_r19_c157 bl[157] br[157] wl[19] vdd gnd cell_6t
Xbit_r20_c157 bl[157] br[157] wl[20] vdd gnd cell_6t
Xbit_r21_c157 bl[157] br[157] wl[21] vdd gnd cell_6t
Xbit_r22_c157 bl[157] br[157] wl[22] vdd gnd cell_6t
Xbit_r23_c157 bl[157] br[157] wl[23] vdd gnd cell_6t
Xbit_r24_c157 bl[157] br[157] wl[24] vdd gnd cell_6t
Xbit_r25_c157 bl[157] br[157] wl[25] vdd gnd cell_6t
Xbit_r26_c157 bl[157] br[157] wl[26] vdd gnd cell_6t
Xbit_r27_c157 bl[157] br[157] wl[27] vdd gnd cell_6t
Xbit_r28_c157 bl[157] br[157] wl[28] vdd gnd cell_6t
Xbit_r29_c157 bl[157] br[157] wl[29] vdd gnd cell_6t
Xbit_r30_c157 bl[157] br[157] wl[30] vdd gnd cell_6t
Xbit_r31_c157 bl[157] br[157] wl[31] vdd gnd cell_6t
Xbit_r32_c157 bl[157] br[157] wl[32] vdd gnd cell_6t
Xbit_r33_c157 bl[157] br[157] wl[33] vdd gnd cell_6t
Xbit_r34_c157 bl[157] br[157] wl[34] vdd gnd cell_6t
Xbit_r35_c157 bl[157] br[157] wl[35] vdd gnd cell_6t
Xbit_r36_c157 bl[157] br[157] wl[36] vdd gnd cell_6t
Xbit_r37_c157 bl[157] br[157] wl[37] vdd gnd cell_6t
Xbit_r38_c157 bl[157] br[157] wl[38] vdd gnd cell_6t
Xbit_r39_c157 bl[157] br[157] wl[39] vdd gnd cell_6t
Xbit_r40_c157 bl[157] br[157] wl[40] vdd gnd cell_6t
Xbit_r41_c157 bl[157] br[157] wl[41] vdd gnd cell_6t
Xbit_r42_c157 bl[157] br[157] wl[42] vdd gnd cell_6t
Xbit_r43_c157 bl[157] br[157] wl[43] vdd gnd cell_6t
Xbit_r44_c157 bl[157] br[157] wl[44] vdd gnd cell_6t
Xbit_r45_c157 bl[157] br[157] wl[45] vdd gnd cell_6t
Xbit_r46_c157 bl[157] br[157] wl[46] vdd gnd cell_6t
Xbit_r47_c157 bl[157] br[157] wl[47] vdd gnd cell_6t
Xbit_r48_c157 bl[157] br[157] wl[48] vdd gnd cell_6t
Xbit_r49_c157 bl[157] br[157] wl[49] vdd gnd cell_6t
Xbit_r50_c157 bl[157] br[157] wl[50] vdd gnd cell_6t
Xbit_r51_c157 bl[157] br[157] wl[51] vdd gnd cell_6t
Xbit_r52_c157 bl[157] br[157] wl[52] vdd gnd cell_6t
Xbit_r53_c157 bl[157] br[157] wl[53] vdd gnd cell_6t
Xbit_r54_c157 bl[157] br[157] wl[54] vdd gnd cell_6t
Xbit_r55_c157 bl[157] br[157] wl[55] vdd gnd cell_6t
Xbit_r56_c157 bl[157] br[157] wl[56] vdd gnd cell_6t
Xbit_r57_c157 bl[157] br[157] wl[57] vdd gnd cell_6t
Xbit_r58_c157 bl[157] br[157] wl[58] vdd gnd cell_6t
Xbit_r59_c157 bl[157] br[157] wl[59] vdd gnd cell_6t
Xbit_r60_c157 bl[157] br[157] wl[60] vdd gnd cell_6t
Xbit_r61_c157 bl[157] br[157] wl[61] vdd gnd cell_6t
Xbit_r62_c157 bl[157] br[157] wl[62] vdd gnd cell_6t
Xbit_r63_c157 bl[157] br[157] wl[63] vdd gnd cell_6t
Xbit_r64_c157 bl[157] br[157] wl[64] vdd gnd cell_6t
Xbit_r65_c157 bl[157] br[157] wl[65] vdd gnd cell_6t
Xbit_r66_c157 bl[157] br[157] wl[66] vdd gnd cell_6t
Xbit_r67_c157 bl[157] br[157] wl[67] vdd gnd cell_6t
Xbit_r68_c157 bl[157] br[157] wl[68] vdd gnd cell_6t
Xbit_r69_c157 bl[157] br[157] wl[69] vdd gnd cell_6t
Xbit_r70_c157 bl[157] br[157] wl[70] vdd gnd cell_6t
Xbit_r71_c157 bl[157] br[157] wl[71] vdd gnd cell_6t
Xbit_r72_c157 bl[157] br[157] wl[72] vdd gnd cell_6t
Xbit_r73_c157 bl[157] br[157] wl[73] vdd gnd cell_6t
Xbit_r74_c157 bl[157] br[157] wl[74] vdd gnd cell_6t
Xbit_r75_c157 bl[157] br[157] wl[75] vdd gnd cell_6t
Xbit_r76_c157 bl[157] br[157] wl[76] vdd gnd cell_6t
Xbit_r77_c157 bl[157] br[157] wl[77] vdd gnd cell_6t
Xbit_r78_c157 bl[157] br[157] wl[78] vdd gnd cell_6t
Xbit_r79_c157 bl[157] br[157] wl[79] vdd gnd cell_6t
Xbit_r80_c157 bl[157] br[157] wl[80] vdd gnd cell_6t
Xbit_r81_c157 bl[157] br[157] wl[81] vdd gnd cell_6t
Xbit_r82_c157 bl[157] br[157] wl[82] vdd gnd cell_6t
Xbit_r83_c157 bl[157] br[157] wl[83] vdd gnd cell_6t
Xbit_r84_c157 bl[157] br[157] wl[84] vdd gnd cell_6t
Xbit_r85_c157 bl[157] br[157] wl[85] vdd gnd cell_6t
Xbit_r86_c157 bl[157] br[157] wl[86] vdd gnd cell_6t
Xbit_r87_c157 bl[157] br[157] wl[87] vdd gnd cell_6t
Xbit_r88_c157 bl[157] br[157] wl[88] vdd gnd cell_6t
Xbit_r89_c157 bl[157] br[157] wl[89] vdd gnd cell_6t
Xbit_r90_c157 bl[157] br[157] wl[90] vdd gnd cell_6t
Xbit_r91_c157 bl[157] br[157] wl[91] vdd gnd cell_6t
Xbit_r92_c157 bl[157] br[157] wl[92] vdd gnd cell_6t
Xbit_r93_c157 bl[157] br[157] wl[93] vdd gnd cell_6t
Xbit_r94_c157 bl[157] br[157] wl[94] vdd gnd cell_6t
Xbit_r95_c157 bl[157] br[157] wl[95] vdd gnd cell_6t
Xbit_r96_c157 bl[157] br[157] wl[96] vdd gnd cell_6t
Xbit_r97_c157 bl[157] br[157] wl[97] vdd gnd cell_6t
Xbit_r98_c157 bl[157] br[157] wl[98] vdd gnd cell_6t
Xbit_r99_c157 bl[157] br[157] wl[99] vdd gnd cell_6t
Xbit_r100_c157 bl[157] br[157] wl[100] vdd gnd cell_6t
Xbit_r101_c157 bl[157] br[157] wl[101] vdd gnd cell_6t
Xbit_r102_c157 bl[157] br[157] wl[102] vdd gnd cell_6t
Xbit_r103_c157 bl[157] br[157] wl[103] vdd gnd cell_6t
Xbit_r104_c157 bl[157] br[157] wl[104] vdd gnd cell_6t
Xbit_r105_c157 bl[157] br[157] wl[105] vdd gnd cell_6t
Xbit_r106_c157 bl[157] br[157] wl[106] vdd gnd cell_6t
Xbit_r107_c157 bl[157] br[157] wl[107] vdd gnd cell_6t
Xbit_r108_c157 bl[157] br[157] wl[108] vdd gnd cell_6t
Xbit_r109_c157 bl[157] br[157] wl[109] vdd gnd cell_6t
Xbit_r110_c157 bl[157] br[157] wl[110] vdd gnd cell_6t
Xbit_r111_c157 bl[157] br[157] wl[111] vdd gnd cell_6t
Xbit_r112_c157 bl[157] br[157] wl[112] vdd gnd cell_6t
Xbit_r113_c157 bl[157] br[157] wl[113] vdd gnd cell_6t
Xbit_r114_c157 bl[157] br[157] wl[114] vdd gnd cell_6t
Xbit_r115_c157 bl[157] br[157] wl[115] vdd gnd cell_6t
Xbit_r116_c157 bl[157] br[157] wl[116] vdd gnd cell_6t
Xbit_r117_c157 bl[157] br[157] wl[117] vdd gnd cell_6t
Xbit_r118_c157 bl[157] br[157] wl[118] vdd gnd cell_6t
Xbit_r119_c157 bl[157] br[157] wl[119] vdd gnd cell_6t
Xbit_r120_c157 bl[157] br[157] wl[120] vdd gnd cell_6t
Xbit_r121_c157 bl[157] br[157] wl[121] vdd gnd cell_6t
Xbit_r122_c157 bl[157] br[157] wl[122] vdd gnd cell_6t
Xbit_r123_c157 bl[157] br[157] wl[123] vdd gnd cell_6t
Xbit_r124_c157 bl[157] br[157] wl[124] vdd gnd cell_6t
Xbit_r125_c157 bl[157] br[157] wl[125] vdd gnd cell_6t
Xbit_r126_c157 bl[157] br[157] wl[126] vdd gnd cell_6t
Xbit_r127_c157 bl[157] br[157] wl[127] vdd gnd cell_6t
Xbit_r0_c158 bl[158] br[158] wl[0] vdd gnd cell_6t
Xbit_r1_c158 bl[158] br[158] wl[1] vdd gnd cell_6t
Xbit_r2_c158 bl[158] br[158] wl[2] vdd gnd cell_6t
Xbit_r3_c158 bl[158] br[158] wl[3] vdd gnd cell_6t
Xbit_r4_c158 bl[158] br[158] wl[4] vdd gnd cell_6t
Xbit_r5_c158 bl[158] br[158] wl[5] vdd gnd cell_6t
Xbit_r6_c158 bl[158] br[158] wl[6] vdd gnd cell_6t
Xbit_r7_c158 bl[158] br[158] wl[7] vdd gnd cell_6t
Xbit_r8_c158 bl[158] br[158] wl[8] vdd gnd cell_6t
Xbit_r9_c158 bl[158] br[158] wl[9] vdd gnd cell_6t
Xbit_r10_c158 bl[158] br[158] wl[10] vdd gnd cell_6t
Xbit_r11_c158 bl[158] br[158] wl[11] vdd gnd cell_6t
Xbit_r12_c158 bl[158] br[158] wl[12] vdd gnd cell_6t
Xbit_r13_c158 bl[158] br[158] wl[13] vdd gnd cell_6t
Xbit_r14_c158 bl[158] br[158] wl[14] vdd gnd cell_6t
Xbit_r15_c158 bl[158] br[158] wl[15] vdd gnd cell_6t
Xbit_r16_c158 bl[158] br[158] wl[16] vdd gnd cell_6t
Xbit_r17_c158 bl[158] br[158] wl[17] vdd gnd cell_6t
Xbit_r18_c158 bl[158] br[158] wl[18] vdd gnd cell_6t
Xbit_r19_c158 bl[158] br[158] wl[19] vdd gnd cell_6t
Xbit_r20_c158 bl[158] br[158] wl[20] vdd gnd cell_6t
Xbit_r21_c158 bl[158] br[158] wl[21] vdd gnd cell_6t
Xbit_r22_c158 bl[158] br[158] wl[22] vdd gnd cell_6t
Xbit_r23_c158 bl[158] br[158] wl[23] vdd gnd cell_6t
Xbit_r24_c158 bl[158] br[158] wl[24] vdd gnd cell_6t
Xbit_r25_c158 bl[158] br[158] wl[25] vdd gnd cell_6t
Xbit_r26_c158 bl[158] br[158] wl[26] vdd gnd cell_6t
Xbit_r27_c158 bl[158] br[158] wl[27] vdd gnd cell_6t
Xbit_r28_c158 bl[158] br[158] wl[28] vdd gnd cell_6t
Xbit_r29_c158 bl[158] br[158] wl[29] vdd gnd cell_6t
Xbit_r30_c158 bl[158] br[158] wl[30] vdd gnd cell_6t
Xbit_r31_c158 bl[158] br[158] wl[31] vdd gnd cell_6t
Xbit_r32_c158 bl[158] br[158] wl[32] vdd gnd cell_6t
Xbit_r33_c158 bl[158] br[158] wl[33] vdd gnd cell_6t
Xbit_r34_c158 bl[158] br[158] wl[34] vdd gnd cell_6t
Xbit_r35_c158 bl[158] br[158] wl[35] vdd gnd cell_6t
Xbit_r36_c158 bl[158] br[158] wl[36] vdd gnd cell_6t
Xbit_r37_c158 bl[158] br[158] wl[37] vdd gnd cell_6t
Xbit_r38_c158 bl[158] br[158] wl[38] vdd gnd cell_6t
Xbit_r39_c158 bl[158] br[158] wl[39] vdd gnd cell_6t
Xbit_r40_c158 bl[158] br[158] wl[40] vdd gnd cell_6t
Xbit_r41_c158 bl[158] br[158] wl[41] vdd gnd cell_6t
Xbit_r42_c158 bl[158] br[158] wl[42] vdd gnd cell_6t
Xbit_r43_c158 bl[158] br[158] wl[43] vdd gnd cell_6t
Xbit_r44_c158 bl[158] br[158] wl[44] vdd gnd cell_6t
Xbit_r45_c158 bl[158] br[158] wl[45] vdd gnd cell_6t
Xbit_r46_c158 bl[158] br[158] wl[46] vdd gnd cell_6t
Xbit_r47_c158 bl[158] br[158] wl[47] vdd gnd cell_6t
Xbit_r48_c158 bl[158] br[158] wl[48] vdd gnd cell_6t
Xbit_r49_c158 bl[158] br[158] wl[49] vdd gnd cell_6t
Xbit_r50_c158 bl[158] br[158] wl[50] vdd gnd cell_6t
Xbit_r51_c158 bl[158] br[158] wl[51] vdd gnd cell_6t
Xbit_r52_c158 bl[158] br[158] wl[52] vdd gnd cell_6t
Xbit_r53_c158 bl[158] br[158] wl[53] vdd gnd cell_6t
Xbit_r54_c158 bl[158] br[158] wl[54] vdd gnd cell_6t
Xbit_r55_c158 bl[158] br[158] wl[55] vdd gnd cell_6t
Xbit_r56_c158 bl[158] br[158] wl[56] vdd gnd cell_6t
Xbit_r57_c158 bl[158] br[158] wl[57] vdd gnd cell_6t
Xbit_r58_c158 bl[158] br[158] wl[58] vdd gnd cell_6t
Xbit_r59_c158 bl[158] br[158] wl[59] vdd gnd cell_6t
Xbit_r60_c158 bl[158] br[158] wl[60] vdd gnd cell_6t
Xbit_r61_c158 bl[158] br[158] wl[61] vdd gnd cell_6t
Xbit_r62_c158 bl[158] br[158] wl[62] vdd gnd cell_6t
Xbit_r63_c158 bl[158] br[158] wl[63] vdd gnd cell_6t
Xbit_r64_c158 bl[158] br[158] wl[64] vdd gnd cell_6t
Xbit_r65_c158 bl[158] br[158] wl[65] vdd gnd cell_6t
Xbit_r66_c158 bl[158] br[158] wl[66] vdd gnd cell_6t
Xbit_r67_c158 bl[158] br[158] wl[67] vdd gnd cell_6t
Xbit_r68_c158 bl[158] br[158] wl[68] vdd gnd cell_6t
Xbit_r69_c158 bl[158] br[158] wl[69] vdd gnd cell_6t
Xbit_r70_c158 bl[158] br[158] wl[70] vdd gnd cell_6t
Xbit_r71_c158 bl[158] br[158] wl[71] vdd gnd cell_6t
Xbit_r72_c158 bl[158] br[158] wl[72] vdd gnd cell_6t
Xbit_r73_c158 bl[158] br[158] wl[73] vdd gnd cell_6t
Xbit_r74_c158 bl[158] br[158] wl[74] vdd gnd cell_6t
Xbit_r75_c158 bl[158] br[158] wl[75] vdd gnd cell_6t
Xbit_r76_c158 bl[158] br[158] wl[76] vdd gnd cell_6t
Xbit_r77_c158 bl[158] br[158] wl[77] vdd gnd cell_6t
Xbit_r78_c158 bl[158] br[158] wl[78] vdd gnd cell_6t
Xbit_r79_c158 bl[158] br[158] wl[79] vdd gnd cell_6t
Xbit_r80_c158 bl[158] br[158] wl[80] vdd gnd cell_6t
Xbit_r81_c158 bl[158] br[158] wl[81] vdd gnd cell_6t
Xbit_r82_c158 bl[158] br[158] wl[82] vdd gnd cell_6t
Xbit_r83_c158 bl[158] br[158] wl[83] vdd gnd cell_6t
Xbit_r84_c158 bl[158] br[158] wl[84] vdd gnd cell_6t
Xbit_r85_c158 bl[158] br[158] wl[85] vdd gnd cell_6t
Xbit_r86_c158 bl[158] br[158] wl[86] vdd gnd cell_6t
Xbit_r87_c158 bl[158] br[158] wl[87] vdd gnd cell_6t
Xbit_r88_c158 bl[158] br[158] wl[88] vdd gnd cell_6t
Xbit_r89_c158 bl[158] br[158] wl[89] vdd gnd cell_6t
Xbit_r90_c158 bl[158] br[158] wl[90] vdd gnd cell_6t
Xbit_r91_c158 bl[158] br[158] wl[91] vdd gnd cell_6t
Xbit_r92_c158 bl[158] br[158] wl[92] vdd gnd cell_6t
Xbit_r93_c158 bl[158] br[158] wl[93] vdd gnd cell_6t
Xbit_r94_c158 bl[158] br[158] wl[94] vdd gnd cell_6t
Xbit_r95_c158 bl[158] br[158] wl[95] vdd gnd cell_6t
Xbit_r96_c158 bl[158] br[158] wl[96] vdd gnd cell_6t
Xbit_r97_c158 bl[158] br[158] wl[97] vdd gnd cell_6t
Xbit_r98_c158 bl[158] br[158] wl[98] vdd gnd cell_6t
Xbit_r99_c158 bl[158] br[158] wl[99] vdd gnd cell_6t
Xbit_r100_c158 bl[158] br[158] wl[100] vdd gnd cell_6t
Xbit_r101_c158 bl[158] br[158] wl[101] vdd gnd cell_6t
Xbit_r102_c158 bl[158] br[158] wl[102] vdd gnd cell_6t
Xbit_r103_c158 bl[158] br[158] wl[103] vdd gnd cell_6t
Xbit_r104_c158 bl[158] br[158] wl[104] vdd gnd cell_6t
Xbit_r105_c158 bl[158] br[158] wl[105] vdd gnd cell_6t
Xbit_r106_c158 bl[158] br[158] wl[106] vdd gnd cell_6t
Xbit_r107_c158 bl[158] br[158] wl[107] vdd gnd cell_6t
Xbit_r108_c158 bl[158] br[158] wl[108] vdd gnd cell_6t
Xbit_r109_c158 bl[158] br[158] wl[109] vdd gnd cell_6t
Xbit_r110_c158 bl[158] br[158] wl[110] vdd gnd cell_6t
Xbit_r111_c158 bl[158] br[158] wl[111] vdd gnd cell_6t
Xbit_r112_c158 bl[158] br[158] wl[112] vdd gnd cell_6t
Xbit_r113_c158 bl[158] br[158] wl[113] vdd gnd cell_6t
Xbit_r114_c158 bl[158] br[158] wl[114] vdd gnd cell_6t
Xbit_r115_c158 bl[158] br[158] wl[115] vdd gnd cell_6t
Xbit_r116_c158 bl[158] br[158] wl[116] vdd gnd cell_6t
Xbit_r117_c158 bl[158] br[158] wl[117] vdd gnd cell_6t
Xbit_r118_c158 bl[158] br[158] wl[118] vdd gnd cell_6t
Xbit_r119_c158 bl[158] br[158] wl[119] vdd gnd cell_6t
Xbit_r120_c158 bl[158] br[158] wl[120] vdd gnd cell_6t
Xbit_r121_c158 bl[158] br[158] wl[121] vdd gnd cell_6t
Xbit_r122_c158 bl[158] br[158] wl[122] vdd gnd cell_6t
Xbit_r123_c158 bl[158] br[158] wl[123] vdd gnd cell_6t
Xbit_r124_c158 bl[158] br[158] wl[124] vdd gnd cell_6t
Xbit_r125_c158 bl[158] br[158] wl[125] vdd gnd cell_6t
Xbit_r126_c158 bl[158] br[158] wl[126] vdd gnd cell_6t
Xbit_r127_c158 bl[158] br[158] wl[127] vdd gnd cell_6t
Xbit_r0_c159 bl[159] br[159] wl[0] vdd gnd cell_6t
Xbit_r1_c159 bl[159] br[159] wl[1] vdd gnd cell_6t
Xbit_r2_c159 bl[159] br[159] wl[2] vdd gnd cell_6t
Xbit_r3_c159 bl[159] br[159] wl[3] vdd gnd cell_6t
Xbit_r4_c159 bl[159] br[159] wl[4] vdd gnd cell_6t
Xbit_r5_c159 bl[159] br[159] wl[5] vdd gnd cell_6t
Xbit_r6_c159 bl[159] br[159] wl[6] vdd gnd cell_6t
Xbit_r7_c159 bl[159] br[159] wl[7] vdd gnd cell_6t
Xbit_r8_c159 bl[159] br[159] wl[8] vdd gnd cell_6t
Xbit_r9_c159 bl[159] br[159] wl[9] vdd gnd cell_6t
Xbit_r10_c159 bl[159] br[159] wl[10] vdd gnd cell_6t
Xbit_r11_c159 bl[159] br[159] wl[11] vdd gnd cell_6t
Xbit_r12_c159 bl[159] br[159] wl[12] vdd gnd cell_6t
Xbit_r13_c159 bl[159] br[159] wl[13] vdd gnd cell_6t
Xbit_r14_c159 bl[159] br[159] wl[14] vdd gnd cell_6t
Xbit_r15_c159 bl[159] br[159] wl[15] vdd gnd cell_6t
Xbit_r16_c159 bl[159] br[159] wl[16] vdd gnd cell_6t
Xbit_r17_c159 bl[159] br[159] wl[17] vdd gnd cell_6t
Xbit_r18_c159 bl[159] br[159] wl[18] vdd gnd cell_6t
Xbit_r19_c159 bl[159] br[159] wl[19] vdd gnd cell_6t
Xbit_r20_c159 bl[159] br[159] wl[20] vdd gnd cell_6t
Xbit_r21_c159 bl[159] br[159] wl[21] vdd gnd cell_6t
Xbit_r22_c159 bl[159] br[159] wl[22] vdd gnd cell_6t
Xbit_r23_c159 bl[159] br[159] wl[23] vdd gnd cell_6t
Xbit_r24_c159 bl[159] br[159] wl[24] vdd gnd cell_6t
Xbit_r25_c159 bl[159] br[159] wl[25] vdd gnd cell_6t
Xbit_r26_c159 bl[159] br[159] wl[26] vdd gnd cell_6t
Xbit_r27_c159 bl[159] br[159] wl[27] vdd gnd cell_6t
Xbit_r28_c159 bl[159] br[159] wl[28] vdd gnd cell_6t
Xbit_r29_c159 bl[159] br[159] wl[29] vdd gnd cell_6t
Xbit_r30_c159 bl[159] br[159] wl[30] vdd gnd cell_6t
Xbit_r31_c159 bl[159] br[159] wl[31] vdd gnd cell_6t
Xbit_r32_c159 bl[159] br[159] wl[32] vdd gnd cell_6t
Xbit_r33_c159 bl[159] br[159] wl[33] vdd gnd cell_6t
Xbit_r34_c159 bl[159] br[159] wl[34] vdd gnd cell_6t
Xbit_r35_c159 bl[159] br[159] wl[35] vdd gnd cell_6t
Xbit_r36_c159 bl[159] br[159] wl[36] vdd gnd cell_6t
Xbit_r37_c159 bl[159] br[159] wl[37] vdd gnd cell_6t
Xbit_r38_c159 bl[159] br[159] wl[38] vdd gnd cell_6t
Xbit_r39_c159 bl[159] br[159] wl[39] vdd gnd cell_6t
Xbit_r40_c159 bl[159] br[159] wl[40] vdd gnd cell_6t
Xbit_r41_c159 bl[159] br[159] wl[41] vdd gnd cell_6t
Xbit_r42_c159 bl[159] br[159] wl[42] vdd gnd cell_6t
Xbit_r43_c159 bl[159] br[159] wl[43] vdd gnd cell_6t
Xbit_r44_c159 bl[159] br[159] wl[44] vdd gnd cell_6t
Xbit_r45_c159 bl[159] br[159] wl[45] vdd gnd cell_6t
Xbit_r46_c159 bl[159] br[159] wl[46] vdd gnd cell_6t
Xbit_r47_c159 bl[159] br[159] wl[47] vdd gnd cell_6t
Xbit_r48_c159 bl[159] br[159] wl[48] vdd gnd cell_6t
Xbit_r49_c159 bl[159] br[159] wl[49] vdd gnd cell_6t
Xbit_r50_c159 bl[159] br[159] wl[50] vdd gnd cell_6t
Xbit_r51_c159 bl[159] br[159] wl[51] vdd gnd cell_6t
Xbit_r52_c159 bl[159] br[159] wl[52] vdd gnd cell_6t
Xbit_r53_c159 bl[159] br[159] wl[53] vdd gnd cell_6t
Xbit_r54_c159 bl[159] br[159] wl[54] vdd gnd cell_6t
Xbit_r55_c159 bl[159] br[159] wl[55] vdd gnd cell_6t
Xbit_r56_c159 bl[159] br[159] wl[56] vdd gnd cell_6t
Xbit_r57_c159 bl[159] br[159] wl[57] vdd gnd cell_6t
Xbit_r58_c159 bl[159] br[159] wl[58] vdd gnd cell_6t
Xbit_r59_c159 bl[159] br[159] wl[59] vdd gnd cell_6t
Xbit_r60_c159 bl[159] br[159] wl[60] vdd gnd cell_6t
Xbit_r61_c159 bl[159] br[159] wl[61] vdd gnd cell_6t
Xbit_r62_c159 bl[159] br[159] wl[62] vdd gnd cell_6t
Xbit_r63_c159 bl[159] br[159] wl[63] vdd gnd cell_6t
Xbit_r64_c159 bl[159] br[159] wl[64] vdd gnd cell_6t
Xbit_r65_c159 bl[159] br[159] wl[65] vdd gnd cell_6t
Xbit_r66_c159 bl[159] br[159] wl[66] vdd gnd cell_6t
Xbit_r67_c159 bl[159] br[159] wl[67] vdd gnd cell_6t
Xbit_r68_c159 bl[159] br[159] wl[68] vdd gnd cell_6t
Xbit_r69_c159 bl[159] br[159] wl[69] vdd gnd cell_6t
Xbit_r70_c159 bl[159] br[159] wl[70] vdd gnd cell_6t
Xbit_r71_c159 bl[159] br[159] wl[71] vdd gnd cell_6t
Xbit_r72_c159 bl[159] br[159] wl[72] vdd gnd cell_6t
Xbit_r73_c159 bl[159] br[159] wl[73] vdd gnd cell_6t
Xbit_r74_c159 bl[159] br[159] wl[74] vdd gnd cell_6t
Xbit_r75_c159 bl[159] br[159] wl[75] vdd gnd cell_6t
Xbit_r76_c159 bl[159] br[159] wl[76] vdd gnd cell_6t
Xbit_r77_c159 bl[159] br[159] wl[77] vdd gnd cell_6t
Xbit_r78_c159 bl[159] br[159] wl[78] vdd gnd cell_6t
Xbit_r79_c159 bl[159] br[159] wl[79] vdd gnd cell_6t
Xbit_r80_c159 bl[159] br[159] wl[80] vdd gnd cell_6t
Xbit_r81_c159 bl[159] br[159] wl[81] vdd gnd cell_6t
Xbit_r82_c159 bl[159] br[159] wl[82] vdd gnd cell_6t
Xbit_r83_c159 bl[159] br[159] wl[83] vdd gnd cell_6t
Xbit_r84_c159 bl[159] br[159] wl[84] vdd gnd cell_6t
Xbit_r85_c159 bl[159] br[159] wl[85] vdd gnd cell_6t
Xbit_r86_c159 bl[159] br[159] wl[86] vdd gnd cell_6t
Xbit_r87_c159 bl[159] br[159] wl[87] vdd gnd cell_6t
Xbit_r88_c159 bl[159] br[159] wl[88] vdd gnd cell_6t
Xbit_r89_c159 bl[159] br[159] wl[89] vdd gnd cell_6t
Xbit_r90_c159 bl[159] br[159] wl[90] vdd gnd cell_6t
Xbit_r91_c159 bl[159] br[159] wl[91] vdd gnd cell_6t
Xbit_r92_c159 bl[159] br[159] wl[92] vdd gnd cell_6t
Xbit_r93_c159 bl[159] br[159] wl[93] vdd gnd cell_6t
Xbit_r94_c159 bl[159] br[159] wl[94] vdd gnd cell_6t
Xbit_r95_c159 bl[159] br[159] wl[95] vdd gnd cell_6t
Xbit_r96_c159 bl[159] br[159] wl[96] vdd gnd cell_6t
Xbit_r97_c159 bl[159] br[159] wl[97] vdd gnd cell_6t
Xbit_r98_c159 bl[159] br[159] wl[98] vdd gnd cell_6t
Xbit_r99_c159 bl[159] br[159] wl[99] vdd gnd cell_6t
Xbit_r100_c159 bl[159] br[159] wl[100] vdd gnd cell_6t
Xbit_r101_c159 bl[159] br[159] wl[101] vdd gnd cell_6t
Xbit_r102_c159 bl[159] br[159] wl[102] vdd gnd cell_6t
Xbit_r103_c159 bl[159] br[159] wl[103] vdd gnd cell_6t
Xbit_r104_c159 bl[159] br[159] wl[104] vdd gnd cell_6t
Xbit_r105_c159 bl[159] br[159] wl[105] vdd gnd cell_6t
Xbit_r106_c159 bl[159] br[159] wl[106] vdd gnd cell_6t
Xbit_r107_c159 bl[159] br[159] wl[107] vdd gnd cell_6t
Xbit_r108_c159 bl[159] br[159] wl[108] vdd gnd cell_6t
Xbit_r109_c159 bl[159] br[159] wl[109] vdd gnd cell_6t
Xbit_r110_c159 bl[159] br[159] wl[110] vdd gnd cell_6t
Xbit_r111_c159 bl[159] br[159] wl[111] vdd gnd cell_6t
Xbit_r112_c159 bl[159] br[159] wl[112] vdd gnd cell_6t
Xbit_r113_c159 bl[159] br[159] wl[113] vdd gnd cell_6t
Xbit_r114_c159 bl[159] br[159] wl[114] vdd gnd cell_6t
Xbit_r115_c159 bl[159] br[159] wl[115] vdd gnd cell_6t
Xbit_r116_c159 bl[159] br[159] wl[116] vdd gnd cell_6t
Xbit_r117_c159 bl[159] br[159] wl[117] vdd gnd cell_6t
Xbit_r118_c159 bl[159] br[159] wl[118] vdd gnd cell_6t
Xbit_r119_c159 bl[159] br[159] wl[119] vdd gnd cell_6t
Xbit_r120_c159 bl[159] br[159] wl[120] vdd gnd cell_6t
Xbit_r121_c159 bl[159] br[159] wl[121] vdd gnd cell_6t
Xbit_r122_c159 bl[159] br[159] wl[122] vdd gnd cell_6t
Xbit_r123_c159 bl[159] br[159] wl[123] vdd gnd cell_6t
Xbit_r124_c159 bl[159] br[159] wl[124] vdd gnd cell_6t
Xbit_r125_c159 bl[159] br[159] wl[125] vdd gnd cell_6t
Xbit_r126_c159 bl[159] br[159] wl[126] vdd gnd cell_6t
Xbit_r127_c159 bl[159] br[159] wl[127] vdd gnd cell_6t
Xbit_r0_c160 bl[160] br[160] wl[0] vdd gnd cell_6t
Xbit_r1_c160 bl[160] br[160] wl[1] vdd gnd cell_6t
Xbit_r2_c160 bl[160] br[160] wl[2] vdd gnd cell_6t
Xbit_r3_c160 bl[160] br[160] wl[3] vdd gnd cell_6t
Xbit_r4_c160 bl[160] br[160] wl[4] vdd gnd cell_6t
Xbit_r5_c160 bl[160] br[160] wl[5] vdd gnd cell_6t
Xbit_r6_c160 bl[160] br[160] wl[6] vdd gnd cell_6t
Xbit_r7_c160 bl[160] br[160] wl[7] vdd gnd cell_6t
Xbit_r8_c160 bl[160] br[160] wl[8] vdd gnd cell_6t
Xbit_r9_c160 bl[160] br[160] wl[9] vdd gnd cell_6t
Xbit_r10_c160 bl[160] br[160] wl[10] vdd gnd cell_6t
Xbit_r11_c160 bl[160] br[160] wl[11] vdd gnd cell_6t
Xbit_r12_c160 bl[160] br[160] wl[12] vdd gnd cell_6t
Xbit_r13_c160 bl[160] br[160] wl[13] vdd gnd cell_6t
Xbit_r14_c160 bl[160] br[160] wl[14] vdd gnd cell_6t
Xbit_r15_c160 bl[160] br[160] wl[15] vdd gnd cell_6t
Xbit_r16_c160 bl[160] br[160] wl[16] vdd gnd cell_6t
Xbit_r17_c160 bl[160] br[160] wl[17] vdd gnd cell_6t
Xbit_r18_c160 bl[160] br[160] wl[18] vdd gnd cell_6t
Xbit_r19_c160 bl[160] br[160] wl[19] vdd gnd cell_6t
Xbit_r20_c160 bl[160] br[160] wl[20] vdd gnd cell_6t
Xbit_r21_c160 bl[160] br[160] wl[21] vdd gnd cell_6t
Xbit_r22_c160 bl[160] br[160] wl[22] vdd gnd cell_6t
Xbit_r23_c160 bl[160] br[160] wl[23] vdd gnd cell_6t
Xbit_r24_c160 bl[160] br[160] wl[24] vdd gnd cell_6t
Xbit_r25_c160 bl[160] br[160] wl[25] vdd gnd cell_6t
Xbit_r26_c160 bl[160] br[160] wl[26] vdd gnd cell_6t
Xbit_r27_c160 bl[160] br[160] wl[27] vdd gnd cell_6t
Xbit_r28_c160 bl[160] br[160] wl[28] vdd gnd cell_6t
Xbit_r29_c160 bl[160] br[160] wl[29] vdd gnd cell_6t
Xbit_r30_c160 bl[160] br[160] wl[30] vdd gnd cell_6t
Xbit_r31_c160 bl[160] br[160] wl[31] vdd gnd cell_6t
Xbit_r32_c160 bl[160] br[160] wl[32] vdd gnd cell_6t
Xbit_r33_c160 bl[160] br[160] wl[33] vdd gnd cell_6t
Xbit_r34_c160 bl[160] br[160] wl[34] vdd gnd cell_6t
Xbit_r35_c160 bl[160] br[160] wl[35] vdd gnd cell_6t
Xbit_r36_c160 bl[160] br[160] wl[36] vdd gnd cell_6t
Xbit_r37_c160 bl[160] br[160] wl[37] vdd gnd cell_6t
Xbit_r38_c160 bl[160] br[160] wl[38] vdd gnd cell_6t
Xbit_r39_c160 bl[160] br[160] wl[39] vdd gnd cell_6t
Xbit_r40_c160 bl[160] br[160] wl[40] vdd gnd cell_6t
Xbit_r41_c160 bl[160] br[160] wl[41] vdd gnd cell_6t
Xbit_r42_c160 bl[160] br[160] wl[42] vdd gnd cell_6t
Xbit_r43_c160 bl[160] br[160] wl[43] vdd gnd cell_6t
Xbit_r44_c160 bl[160] br[160] wl[44] vdd gnd cell_6t
Xbit_r45_c160 bl[160] br[160] wl[45] vdd gnd cell_6t
Xbit_r46_c160 bl[160] br[160] wl[46] vdd gnd cell_6t
Xbit_r47_c160 bl[160] br[160] wl[47] vdd gnd cell_6t
Xbit_r48_c160 bl[160] br[160] wl[48] vdd gnd cell_6t
Xbit_r49_c160 bl[160] br[160] wl[49] vdd gnd cell_6t
Xbit_r50_c160 bl[160] br[160] wl[50] vdd gnd cell_6t
Xbit_r51_c160 bl[160] br[160] wl[51] vdd gnd cell_6t
Xbit_r52_c160 bl[160] br[160] wl[52] vdd gnd cell_6t
Xbit_r53_c160 bl[160] br[160] wl[53] vdd gnd cell_6t
Xbit_r54_c160 bl[160] br[160] wl[54] vdd gnd cell_6t
Xbit_r55_c160 bl[160] br[160] wl[55] vdd gnd cell_6t
Xbit_r56_c160 bl[160] br[160] wl[56] vdd gnd cell_6t
Xbit_r57_c160 bl[160] br[160] wl[57] vdd gnd cell_6t
Xbit_r58_c160 bl[160] br[160] wl[58] vdd gnd cell_6t
Xbit_r59_c160 bl[160] br[160] wl[59] vdd gnd cell_6t
Xbit_r60_c160 bl[160] br[160] wl[60] vdd gnd cell_6t
Xbit_r61_c160 bl[160] br[160] wl[61] vdd gnd cell_6t
Xbit_r62_c160 bl[160] br[160] wl[62] vdd gnd cell_6t
Xbit_r63_c160 bl[160] br[160] wl[63] vdd gnd cell_6t
Xbit_r64_c160 bl[160] br[160] wl[64] vdd gnd cell_6t
Xbit_r65_c160 bl[160] br[160] wl[65] vdd gnd cell_6t
Xbit_r66_c160 bl[160] br[160] wl[66] vdd gnd cell_6t
Xbit_r67_c160 bl[160] br[160] wl[67] vdd gnd cell_6t
Xbit_r68_c160 bl[160] br[160] wl[68] vdd gnd cell_6t
Xbit_r69_c160 bl[160] br[160] wl[69] vdd gnd cell_6t
Xbit_r70_c160 bl[160] br[160] wl[70] vdd gnd cell_6t
Xbit_r71_c160 bl[160] br[160] wl[71] vdd gnd cell_6t
Xbit_r72_c160 bl[160] br[160] wl[72] vdd gnd cell_6t
Xbit_r73_c160 bl[160] br[160] wl[73] vdd gnd cell_6t
Xbit_r74_c160 bl[160] br[160] wl[74] vdd gnd cell_6t
Xbit_r75_c160 bl[160] br[160] wl[75] vdd gnd cell_6t
Xbit_r76_c160 bl[160] br[160] wl[76] vdd gnd cell_6t
Xbit_r77_c160 bl[160] br[160] wl[77] vdd gnd cell_6t
Xbit_r78_c160 bl[160] br[160] wl[78] vdd gnd cell_6t
Xbit_r79_c160 bl[160] br[160] wl[79] vdd gnd cell_6t
Xbit_r80_c160 bl[160] br[160] wl[80] vdd gnd cell_6t
Xbit_r81_c160 bl[160] br[160] wl[81] vdd gnd cell_6t
Xbit_r82_c160 bl[160] br[160] wl[82] vdd gnd cell_6t
Xbit_r83_c160 bl[160] br[160] wl[83] vdd gnd cell_6t
Xbit_r84_c160 bl[160] br[160] wl[84] vdd gnd cell_6t
Xbit_r85_c160 bl[160] br[160] wl[85] vdd gnd cell_6t
Xbit_r86_c160 bl[160] br[160] wl[86] vdd gnd cell_6t
Xbit_r87_c160 bl[160] br[160] wl[87] vdd gnd cell_6t
Xbit_r88_c160 bl[160] br[160] wl[88] vdd gnd cell_6t
Xbit_r89_c160 bl[160] br[160] wl[89] vdd gnd cell_6t
Xbit_r90_c160 bl[160] br[160] wl[90] vdd gnd cell_6t
Xbit_r91_c160 bl[160] br[160] wl[91] vdd gnd cell_6t
Xbit_r92_c160 bl[160] br[160] wl[92] vdd gnd cell_6t
Xbit_r93_c160 bl[160] br[160] wl[93] vdd gnd cell_6t
Xbit_r94_c160 bl[160] br[160] wl[94] vdd gnd cell_6t
Xbit_r95_c160 bl[160] br[160] wl[95] vdd gnd cell_6t
Xbit_r96_c160 bl[160] br[160] wl[96] vdd gnd cell_6t
Xbit_r97_c160 bl[160] br[160] wl[97] vdd gnd cell_6t
Xbit_r98_c160 bl[160] br[160] wl[98] vdd gnd cell_6t
Xbit_r99_c160 bl[160] br[160] wl[99] vdd gnd cell_6t
Xbit_r100_c160 bl[160] br[160] wl[100] vdd gnd cell_6t
Xbit_r101_c160 bl[160] br[160] wl[101] vdd gnd cell_6t
Xbit_r102_c160 bl[160] br[160] wl[102] vdd gnd cell_6t
Xbit_r103_c160 bl[160] br[160] wl[103] vdd gnd cell_6t
Xbit_r104_c160 bl[160] br[160] wl[104] vdd gnd cell_6t
Xbit_r105_c160 bl[160] br[160] wl[105] vdd gnd cell_6t
Xbit_r106_c160 bl[160] br[160] wl[106] vdd gnd cell_6t
Xbit_r107_c160 bl[160] br[160] wl[107] vdd gnd cell_6t
Xbit_r108_c160 bl[160] br[160] wl[108] vdd gnd cell_6t
Xbit_r109_c160 bl[160] br[160] wl[109] vdd gnd cell_6t
Xbit_r110_c160 bl[160] br[160] wl[110] vdd gnd cell_6t
Xbit_r111_c160 bl[160] br[160] wl[111] vdd gnd cell_6t
Xbit_r112_c160 bl[160] br[160] wl[112] vdd gnd cell_6t
Xbit_r113_c160 bl[160] br[160] wl[113] vdd gnd cell_6t
Xbit_r114_c160 bl[160] br[160] wl[114] vdd gnd cell_6t
Xbit_r115_c160 bl[160] br[160] wl[115] vdd gnd cell_6t
Xbit_r116_c160 bl[160] br[160] wl[116] vdd gnd cell_6t
Xbit_r117_c160 bl[160] br[160] wl[117] vdd gnd cell_6t
Xbit_r118_c160 bl[160] br[160] wl[118] vdd gnd cell_6t
Xbit_r119_c160 bl[160] br[160] wl[119] vdd gnd cell_6t
Xbit_r120_c160 bl[160] br[160] wl[120] vdd gnd cell_6t
Xbit_r121_c160 bl[160] br[160] wl[121] vdd gnd cell_6t
Xbit_r122_c160 bl[160] br[160] wl[122] vdd gnd cell_6t
Xbit_r123_c160 bl[160] br[160] wl[123] vdd gnd cell_6t
Xbit_r124_c160 bl[160] br[160] wl[124] vdd gnd cell_6t
Xbit_r125_c160 bl[160] br[160] wl[125] vdd gnd cell_6t
Xbit_r126_c160 bl[160] br[160] wl[126] vdd gnd cell_6t
Xbit_r127_c160 bl[160] br[160] wl[127] vdd gnd cell_6t
Xbit_r0_c161 bl[161] br[161] wl[0] vdd gnd cell_6t
Xbit_r1_c161 bl[161] br[161] wl[1] vdd gnd cell_6t
Xbit_r2_c161 bl[161] br[161] wl[2] vdd gnd cell_6t
Xbit_r3_c161 bl[161] br[161] wl[3] vdd gnd cell_6t
Xbit_r4_c161 bl[161] br[161] wl[4] vdd gnd cell_6t
Xbit_r5_c161 bl[161] br[161] wl[5] vdd gnd cell_6t
Xbit_r6_c161 bl[161] br[161] wl[6] vdd gnd cell_6t
Xbit_r7_c161 bl[161] br[161] wl[7] vdd gnd cell_6t
Xbit_r8_c161 bl[161] br[161] wl[8] vdd gnd cell_6t
Xbit_r9_c161 bl[161] br[161] wl[9] vdd gnd cell_6t
Xbit_r10_c161 bl[161] br[161] wl[10] vdd gnd cell_6t
Xbit_r11_c161 bl[161] br[161] wl[11] vdd gnd cell_6t
Xbit_r12_c161 bl[161] br[161] wl[12] vdd gnd cell_6t
Xbit_r13_c161 bl[161] br[161] wl[13] vdd gnd cell_6t
Xbit_r14_c161 bl[161] br[161] wl[14] vdd gnd cell_6t
Xbit_r15_c161 bl[161] br[161] wl[15] vdd gnd cell_6t
Xbit_r16_c161 bl[161] br[161] wl[16] vdd gnd cell_6t
Xbit_r17_c161 bl[161] br[161] wl[17] vdd gnd cell_6t
Xbit_r18_c161 bl[161] br[161] wl[18] vdd gnd cell_6t
Xbit_r19_c161 bl[161] br[161] wl[19] vdd gnd cell_6t
Xbit_r20_c161 bl[161] br[161] wl[20] vdd gnd cell_6t
Xbit_r21_c161 bl[161] br[161] wl[21] vdd gnd cell_6t
Xbit_r22_c161 bl[161] br[161] wl[22] vdd gnd cell_6t
Xbit_r23_c161 bl[161] br[161] wl[23] vdd gnd cell_6t
Xbit_r24_c161 bl[161] br[161] wl[24] vdd gnd cell_6t
Xbit_r25_c161 bl[161] br[161] wl[25] vdd gnd cell_6t
Xbit_r26_c161 bl[161] br[161] wl[26] vdd gnd cell_6t
Xbit_r27_c161 bl[161] br[161] wl[27] vdd gnd cell_6t
Xbit_r28_c161 bl[161] br[161] wl[28] vdd gnd cell_6t
Xbit_r29_c161 bl[161] br[161] wl[29] vdd gnd cell_6t
Xbit_r30_c161 bl[161] br[161] wl[30] vdd gnd cell_6t
Xbit_r31_c161 bl[161] br[161] wl[31] vdd gnd cell_6t
Xbit_r32_c161 bl[161] br[161] wl[32] vdd gnd cell_6t
Xbit_r33_c161 bl[161] br[161] wl[33] vdd gnd cell_6t
Xbit_r34_c161 bl[161] br[161] wl[34] vdd gnd cell_6t
Xbit_r35_c161 bl[161] br[161] wl[35] vdd gnd cell_6t
Xbit_r36_c161 bl[161] br[161] wl[36] vdd gnd cell_6t
Xbit_r37_c161 bl[161] br[161] wl[37] vdd gnd cell_6t
Xbit_r38_c161 bl[161] br[161] wl[38] vdd gnd cell_6t
Xbit_r39_c161 bl[161] br[161] wl[39] vdd gnd cell_6t
Xbit_r40_c161 bl[161] br[161] wl[40] vdd gnd cell_6t
Xbit_r41_c161 bl[161] br[161] wl[41] vdd gnd cell_6t
Xbit_r42_c161 bl[161] br[161] wl[42] vdd gnd cell_6t
Xbit_r43_c161 bl[161] br[161] wl[43] vdd gnd cell_6t
Xbit_r44_c161 bl[161] br[161] wl[44] vdd gnd cell_6t
Xbit_r45_c161 bl[161] br[161] wl[45] vdd gnd cell_6t
Xbit_r46_c161 bl[161] br[161] wl[46] vdd gnd cell_6t
Xbit_r47_c161 bl[161] br[161] wl[47] vdd gnd cell_6t
Xbit_r48_c161 bl[161] br[161] wl[48] vdd gnd cell_6t
Xbit_r49_c161 bl[161] br[161] wl[49] vdd gnd cell_6t
Xbit_r50_c161 bl[161] br[161] wl[50] vdd gnd cell_6t
Xbit_r51_c161 bl[161] br[161] wl[51] vdd gnd cell_6t
Xbit_r52_c161 bl[161] br[161] wl[52] vdd gnd cell_6t
Xbit_r53_c161 bl[161] br[161] wl[53] vdd gnd cell_6t
Xbit_r54_c161 bl[161] br[161] wl[54] vdd gnd cell_6t
Xbit_r55_c161 bl[161] br[161] wl[55] vdd gnd cell_6t
Xbit_r56_c161 bl[161] br[161] wl[56] vdd gnd cell_6t
Xbit_r57_c161 bl[161] br[161] wl[57] vdd gnd cell_6t
Xbit_r58_c161 bl[161] br[161] wl[58] vdd gnd cell_6t
Xbit_r59_c161 bl[161] br[161] wl[59] vdd gnd cell_6t
Xbit_r60_c161 bl[161] br[161] wl[60] vdd gnd cell_6t
Xbit_r61_c161 bl[161] br[161] wl[61] vdd gnd cell_6t
Xbit_r62_c161 bl[161] br[161] wl[62] vdd gnd cell_6t
Xbit_r63_c161 bl[161] br[161] wl[63] vdd gnd cell_6t
Xbit_r64_c161 bl[161] br[161] wl[64] vdd gnd cell_6t
Xbit_r65_c161 bl[161] br[161] wl[65] vdd gnd cell_6t
Xbit_r66_c161 bl[161] br[161] wl[66] vdd gnd cell_6t
Xbit_r67_c161 bl[161] br[161] wl[67] vdd gnd cell_6t
Xbit_r68_c161 bl[161] br[161] wl[68] vdd gnd cell_6t
Xbit_r69_c161 bl[161] br[161] wl[69] vdd gnd cell_6t
Xbit_r70_c161 bl[161] br[161] wl[70] vdd gnd cell_6t
Xbit_r71_c161 bl[161] br[161] wl[71] vdd gnd cell_6t
Xbit_r72_c161 bl[161] br[161] wl[72] vdd gnd cell_6t
Xbit_r73_c161 bl[161] br[161] wl[73] vdd gnd cell_6t
Xbit_r74_c161 bl[161] br[161] wl[74] vdd gnd cell_6t
Xbit_r75_c161 bl[161] br[161] wl[75] vdd gnd cell_6t
Xbit_r76_c161 bl[161] br[161] wl[76] vdd gnd cell_6t
Xbit_r77_c161 bl[161] br[161] wl[77] vdd gnd cell_6t
Xbit_r78_c161 bl[161] br[161] wl[78] vdd gnd cell_6t
Xbit_r79_c161 bl[161] br[161] wl[79] vdd gnd cell_6t
Xbit_r80_c161 bl[161] br[161] wl[80] vdd gnd cell_6t
Xbit_r81_c161 bl[161] br[161] wl[81] vdd gnd cell_6t
Xbit_r82_c161 bl[161] br[161] wl[82] vdd gnd cell_6t
Xbit_r83_c161 bl[161] br[161] wl[83] vdd gnd cell_6t
Xbit_r84_c161 bl[161] br[161] wl[84] vdd gnd cell_6t
Xbit_r85_c161 bl[161] br[161] wl[85] vdd gnd cell_6t
Xbit_r86_c161 bl[161] br[161] wl[86] vdd gnd cell_6t
Xbit_r87_c161 bl[161] br[161] wl[87] vdd gnd cell_6t
Xbit_r88_c161 bl[161] br[161] wl[88] vdd gnd cell_6t
Xbit_r89_c161 bl[161] br[161] wl[89] vdd gnd cell_6t
Xbit_r90_c161 bl[161] br[161] wl[90] vdd gnd cell_6t
Xbit_r91_c161 bl[161] br[161] wl[91] vdd gnd cell_6t
Xbit_r92_c161 bl[161] br[161] wl[92] vdd gnd cell_6t
Xbit_r93_c161 bl[161] br[161] wl[93] vdd gnd cell_6t
Xbit_r94_c161 bl[161] br[161] wl[94] vdd gnd cell_6t
Xbit_r95_c161 bl[161] br[161] wl[95] vdd gnd cell_6t
Xbit_r96_c161 bl[161] br[161] wl[96] vdd gnd cell_6t
Xbit_r97_c161 bl[161] br[161] wl[97] vdd gnd cell_6t
Xbit_r98_c161 bl[161] br[161] wl[98] vdd gnd cell_6t
Xbit_r99_c161 bl[161] br[161] wl[99] vdd gnd cell_6t
Xbit_r100_c161 bl[161] br[161] wl[100] vdd gnd cell_6t
Xbit_r101_c161 bl[161] br[161] wl[101] vdd gnd cell_6t
Xbit_r102_c161 bl[161] br[161] wl[102] vdd gnd cell_6t
Xbit_r103_c161 bl[161] br[161] wl[103] vdd gnd cell_6t
Xbit_r104_c161 bl[161] br[161] wl[104] vdd gnd cell_6t
Xbit_r105_c161 bl[161] br[161] wl[105] vdd gnd cell_6t
Xbit_r106_c161 bl[161] br[161] wl[106] vdd gnd cell_6t
Xbit_r107_c161 bl[161] br[161] wl[107] vdd gnd cell_6t
Xbit_r108_c161 bl[161] br[161] wl[108] vdd gnd cell_6t
Xbit_r109_c161 bl[161] br[161] wl[109] vdd gnd cell_6t
Xbit_r110_c161 bl[161] br[161] wl[110] vdd gnd cell_6t
Xbit_r111_c161 bl[161] br[161] wl[111] vdd gnd cell_6t
Xbit_r112_c161 bl[161] br[161] wl[112] vdd gnd cell_6t
Xbit_r113_c161 bl[161] br[161] wl[113] vdd gnd cell_6t
Xbit_r114_c161 bl[161] br[161] wl[114] vdd gnd cell_6t
Xbit_r115_c161 bl[161] br[161] wl[115] vdd gnd cell_6t
Xbit_r116_c161 bl[161] br[161] wl[116] vdd gnd cell_6t
Xbit_r117_c161 bl[161] br[161] wl[117] vdd gnd cell_6t
Xbit_r118_c161 bl[161] br[161] wl[118] vdd gnd cell_6t
Xbit_r119_c161 bl[161] br[161] wl[119] vdd gnd cell_6t
Xbit_r120_c161 bl[161] br[161] wl[120] vdd gnd cell_6t
Xbit_r121_c161 bl[161] br[161] wl[121] vdd gnd cell_6t
Xbit_r122_c161 bl[161] br[161] wl[122] vdd gnd cell_6t
Xbit_r123_c161 bl[161] br[161] wl[123] vdd gnd cell_6t
Xbit_r124_c161 bl[161] br[161] wl[124] vdd gnd cell_6t
Xbit_r125_c161 bl[161] br[161] wl[125] vdd gnd cell_6t
Xbit_r126_c161 bl[161] br[161] wl[126] vdd gnd cell_6t
Xbit_r127_c161 bl[161] br[161] wl[127] vdd gnd cell_6t
Xbit_r0_c162 bl[162] br[162] wl[0] vdd gnd cell_6t
Xbit_r1_c162 bl[162] br[162] wl[1] vdd gnd cell_6t
Xbit_r2_c162 bl[162] br[162] wl[2] vdd gnd cell_6t
Xbit_r3_c162 bl[162] br[162] wl[3] vdd gnd cell_6t
Xbit_r4_c162 bl[162] br[162] wl[4] vdd gnd cell_6t
Xbit_r5_c162 bl[162] br[162] wl[5] vdd gnd cell_6t
Xbit_r6_c162 bl[162] br[162] wl[6] vdd gnd cell_6t
Xbit_r7_c162 bl[162] br[162] wl[7] vdd gnd cell_6t
Xbit_r8_c162 bl[162] br[162] wl[8] vdd gnd cell_6t
Xbit_r9_c162 bl[162] br[162] wl[9] vdd gnd cell_6t
Xbit_r10_c162 bl[162] br[162] wl[10] vdd gnd cell_6t
Xbit_r11_c162 bl[162] br[162] wl[11] vdd gnd cell_6t
Xbit_r12_c162 bl[162] br[162] wl[12] vdd gnd cell_6t
Xbit_r13_c162 bl[162] br[162] wl[13] vdd gnd cell_6t
Xbit_r14_c162 bl[162] br[162] wl[14] vdd gnd cell_6t
Xbit_r15_c162 bl[162] br[162] wl[15] vdd gnd cell_6t
Xbit_r16_c162 bl[162] br[162] wl[16] vdd gnd cell_6t
Xbit_r17_c162 bl[162] br[162] wl[17] vdd gnd cell_6t
Xbit_r18_c162 bl[162] br[162] wl[18] vdd gnd cell_6t
Xbit_r19_c162 bl[162] br[162] wl[19] vdd gnd cell_6t
Xbit_r20_c162 bl[162] br[162] wl[20] vdd gnd cell_6t
Xbit_r21_c162 bl[162] br[162] wl[21] vdd gnd cell_6t
Xbit_r22_c162 bl[162] br[162] wl[22] vdd gnd cell_6t
Xbit_r23_c162 bl[162] br[162] wl[23] vdd gnd cell_6t
Xbit_r24_c162 bl[162] br[162] wl[24] vdd gnd cell_6t
Xbit_r25_c162 bl[162] br[162] wl[25] vdd gnd cell_6t
Xbit_r26_c162 bl[162] br[162] wl[26] vdd gnd cell_6t
Xbit_r27_c162 bl[162] br[162] wl[27] vdd gnd cell_6t
Xbit_r28_c162 bl[162] br[162] wl[28] vdd gnd cell_6t
Xbit_r29_c162 bl[162] br[162] wl[29] vdd gnd cell_6t
Xbit_r30_c162 bl[162] br[162] wl[30] vdd gnd cell_6t
Xbit_r31_c162 bl[162] br[162] wl[31] vdd gnd cell_6t
Xbit_r32_c162 bl[162] br[162] wl[32] vdd gnd cell_6t
Xbit_r33_c162 bl[162] br[162] wl[33] vdd gnd cell_6t
Xbit_r34_c162 bl[162] br[162] wl[34] vdd gnd cell_6t
Xbit_r35_c162 bl[162] br[162] wl[35] vdd gnd cell_6t
Xbit_r36_c162 bl[162] br[162] wl[36] vdd gnd cell_6t
Xbit_r37_c162 bl[162] br[162] wl[37] vdd gnd cell_6t
Xbit_r38_c162 bl[162] br[162] wl[38] vdd gnd cell_6t
Xbit_r39_c162 bl[162] br[162] wl[39] vdd gnd cell_6t
Xbit_r40_c162 bl[162] br[162] wl[40] vdd gnd cell_6t
Xbit_r41_c162 bl[162] br[162] wl[41] vdd gnd cell_6t
Xbit_r42_c162 bl[162] br[162] wl[42] vdd gnd cell_6t
Xbit_r43_c162 bl[162] br[162] wl[43] vdd gnd cell_6t
Xbit_r44_c162 bl[162] br[162] wl[44] vdd gnd cell_6t
Xbit_r45_c162 bl[162] br[162] wl[45] vdd gnd cell_6t
Xbit_r46_c162 bl[162] br[162] wl[46] vdd gnd cell_6t
Xbit_r47_c162 bl[162] br[162] wl[47] vdd gnd cell_6t
Xbit_r48_c162 bl[162] br[162] wl[48] vdd gnd cell_6t
Xbit_r49_c162 bl[162] br[162] wl[49] vdd gnd cell_6t
Xbit_r50_c162 bl[162] br[162] wl[50] vdd gnd cell_6t
Xbit_r51_c162 bl[162] br[162] wl[51] vdd gnd cell_6t
Xbit_r52_c162 bl[162] br[162] wl[52] vdd gnd cell_6t
Xbit_r53_c162 bl[162] br[162] wl[53] vdd gnd cell_6t
Xbit_r54_c162 bl[162] br[162] wl[54] vdd gnd cell_6t
Xbit_r55_c162 bl[162] br[162] wl[55] vdd gnd cell_6t
Xbit_r56_c162 bl[162] br[162] wl[56] vdd gnd cell_6t
Xbit_r57_c162 bl[162] br[162] wl[57] vdd gnd cell_6t
Xbit_r58_c162 bl[162] br[162] wl[58] vdd gnd cell_6t
Xbit_r59_c162 bl[162] br[162] wl[59] vdd gnd cell_6t
Xbit_r60_c162 bl[162] br[162] wl[60] vdd gnd cell_6t
Xbit_r61_c162 bl[162] br[162] wl[61] vdd gnd cell_6t
Xbit_r62_c162 bl[162] br[162] wl[62] vdd gnd cell_6t
Xbit_r63_c162 bl[162] br[162] wl[63] vdd gnd cell_6t
Xbit_r64_c162 bl[162] br[162] wl[64] vdd gnd cell_6t
Xbit_r65_c162 bl[162] br[162] wl[65] vdd gnd cell_6t
Xbit_r66_c162 bl[162] br[162] wl[66] vdd gnd cell_6t
Xbit_r67_c162 bl[162] br[162] wl[67] vdd gnd cell_6t
Xbit_r68_c162 bl[162] br[162] wl[68] vdd gnd cell_6t
Xbit_r69_c162 bl[162] br[162] wl[69] vdd gnd cell_6t
Xbit_r70_c162 bl[162] br[162] wl[70] vdd gnd cell_6t
Xbit_r71_c162 bl[162] br[162] wl[71] vdd gnd cell_6t
Xbit_r72_c162 bl[162] br[162] wl[72] vdd gnd cell_6t
Xbit_r73_c162 bl[162] br[162] wl[73] vdd gnd cell_6t
Xbit_r74_c162 bl[162] br[162] wl[74] vdd gnd cell_6t
Xbit_r75_c162 bl[162] br[162] wl[75] vdd gnd cell_6t
Xbit_r76_c162 bl[162] br[162] wl[76] vdd gnd cell_6t
Xbit_r77_c162 bl[162] br[162] wl[77] vdd gnd cell_6t
Xbit_r78_c162 bl[162] br[162] wl[78] vdd gnd cell_6t
Xbit_r79_c162 bl[162] br[162] wl[79] vdd gnd cell_6t
Xbit_r80_c162 bl[162] br[162] wl[80] vdd gnd cell_6t
Xbit_r81_c162 bl[162] br[162] wl[81] vdd gnd cell_6t
Xbit_r82_c162 bl[162] br[162] wl[82] vdd gnd cell_6t
Xbit_r83_c162 bl[162] br[162] wl[83] vdd gnd cell_6t
Xbit_r84_c162 bl[162] br[162] wl[84] vdd gnd cell_6t
Xbit_r85_c162 bl[162] br[162] wl[85] vdd gnd cell_6t
Xbit_r86_c162 bl[162] br[162] wl[86] vdd gnd cell_6t
Xbit_r87_c162 bl[162] br[162] wl[87] vdd gnd cell_6t
Xbit_r88_c162 bl[162] br[162] wl[88] vdd gnd cell_6t
Xbit_r89_c162 bl[162] br[162] wl[89] vdd gnd cell_6t
Xbit_r90_c162 bl[162] br[162] wl[90] vdd gnd cell_6t
Xbit_r91_c162 bl[162] br[162] wl[91] vdd gnd cell_6t
Xbit_r92_c162 bl[162] br[162] wl[92] vdd gnd cell_6t
Xbit_r93_c162 bl[162] br[162] wl[93] vdd gnd cell_6t
Xbit_r94_c162 bl[162] br[162] wl[94] vdd gnd cell_6t
Xbit_r95_c162 bl[162] br[162] wl[95] vdd gnd cell_6t
Xbit_r96_c162 bl[162] br[162] wl[96] vdd gnd cell_6t
Xbit_r97_c162 bl[162] br[162] wl[97] vdd gnd cell_6t
Xbit_r98_c162 bl[162] br[162] wl[98] vdd gnd cell_6t
Xbit_r99_c162 bl[162] br[162] wl[99] vdd gnd cell_6t
Xbit_r100_c162 bl[162] br[162] wl[100] vdd gnd cell_6t
Xbit_r101_c162 bl[162] br[162] wl[101] vdd gnd cell_6t
Xbit_r102_c162 bl[162] br[162] wl[102] vdd gnd cell_6t
Xbit_r103_c162 bl[162] br[162] wl[103] vdd gnd cell_6t
Xbit_r104_c162 bl[162] br[162] wl[104] vdd gnd cell_6t
Xbit_r105_c162 bl[162] br[162] wl[105] vdd gnd cell_6t
Xbit_r106_c162 bl[162] br[162] wl[106] vdd gnd cell_6t
Xbit_r107_c162 bl[162] br[162] wl[107] vdd gnd cell_6t
Xbit_r108_c162 bl[162] br[162] wl[108] vdd gnd cell_6t
Xbit_r109_c162 bl[162] br[162] wl[109] vdd gnd cell_6t
Xbit_r110_c162 bl[162] br[162] wl[110] vdd gnd cell_6t
Xbit_r111_c162 bl[162] br[162] wl[111] vdd gnd cell_6t
Xbit_r112_c162 bl[162] br[162] wl[112] vdd gnd cell_6t
Xbit_r113_c162 bl[162] br[162] wl[113] vdd gnd cell_6t
Xbit_r114_c162 bl[162] br[162] wl[114] vdd gnd cell_6t
Xbit_r115_c162 bl[162] br[162] wl[115] vdd gnd cell_6t
Xbit_r116_c162 bl[162] br[162] wl[116] vdd gnd cell_6t
Xbit_r117_c162 bl[162] br[162] wl[117] vdd gnd cell_6t
Xbit_r118_c162 bl[162] br[162] wl[118] vdd gnd cell_6t
Xbit_r119_c162 bl[162] br[162] wl[119] vdd gnd cell_6t
Xbit_r120_c162 bl[162] br[162] wl[120] vdd gnd cell_6t
Xbit_r121_c162 bl[162] br[162] wl[121] vdd gnd cell_6t
Xbit_r122_c162 bl[162] br[162] wl[122] vdd gnd cell_6t
Xbit_r123_c162 bl[162] br[162] wl[123] vdd gnd cell_6t
Xbit_r124_c162 bl[162] br[162] wl[124] vdd gnd cell_6t
Xbit_r125_c162 bl[162] br[162] wl[125] vdd gnd cell_6t
Xbit_r126_c162 bl[162] br[162] wl[126] vdd gnd cell_6t
Xbit_r127_c162 bl[162] br[162] wl[127] vdd gnd cell_6t
Xbit_r0_c163 bl[163] br[163] wl[0] vdd gnd cell_6t
Xbit_r1_c163 bl[163] br[163] wl[1] vdd gnd cell_6t
Xbit_r2_c163 bl[163] br[163] wl[2] vdd gnd cell_6t
Xbit_r3_c163 bl[163] br[163] wl[3] vdd gnd cell_6t
Xbit_r4_c163 bl[163] br[163] wl[4] vdd gnd cell_6t
Xbit_r5_c163 bl[163] br[163] wl[5] vdd gnd cell_6t
Xbit_r6_c163 bl[163] br[163] wl[6] vdd gnd cell_6t
Xbit_r7_c163 bl[163] br[163] wl[7] vdd gnd cell_6t
Xbit_r8_c163 bl[163] br[163] wl[8] vdd gnd cell_6t
Xbit_r9_c163 bl[163] br[163] wl[9] vdd gnd cell_6t
Xbit_r10_c163 bl[163] br[163] wl[10] vdd gnd cell_6t
Xbit_r11_c163 bl[163] br[163] wl[11] vdd gnd cell_6t
Xbit_r12_c163 bl[163] br[163] wl[12] vdd gnd cell_6t
Xbit_r13_c163 bl[163] br[163] wl[13] vdd gnd cell_6t
Xbit_r14_c163 bl[163] br[163] wl[14] vdd gnd cell_6t
Xbit_r15_c163 bl[163] br[163] wl[15] vdd gnd cell_6t
Xbit_r16_c163 bl[163] br[163] wl[16] vdd gnd cell_6t
Xbit_r17_c163 bl[163] br[163] wl[17] vdd gnd cell_6t
Xbit_r18_c163 bl[163] br[163] wl[18] vdd gnd cell_6t
Xbit_r19_c163 bl[163] br[163] wl[19] vdd gnd cell_6t
Xbit_r20_c163 bl[163] br[163] wl[20] vdd gnd cell_6t
Xbit_r21_c163 bl[163] br[163] wl[21] vdd gnd cell_6t
Xbit_r22_c163 bl[163] br[163] wl[22] vdd gnd cell_6t
Xbit_r23_c163 bl[163] br[163] wl[23] vdd gnd cell_6t
Xbit_r24_c163 bl[163] br[163] wl[24] vdd gnd cell_6t
Xbit_r25_c163 bl[163] br[163] wl[25] vdd gnd cell_6t
Xbit_r26_c163 bl[163] br[163] wl[26] vdd gnd cell_6t
Xbit_r27_c163 bl[163] br[163] wl[27] vdd gnd cell_6t
Xbit_r28_c163 bl[163] br[163] wl[28] vdd gnd cell_6t
Xbit_r29_c163 bl[163] br[163] wl[29] vdd gnd cell_6t
Xbit_r30_c163 bl[163] br[163] wl[30] vdd gnd cell_6t
Xbit_r31_c163 bl[163] br[163] wl[31] vdd gnd cell_6t
Xbit_r32_c163 bl[163] br[163] wl[32] vdd gnd cell_6t
Xbit_r33_c163 bl[163] br[163] wl[33] vdd gnd cell_6t
Xbit_r34_c163 bl[163] br[163] wl[34] vdd gnd cell_6t
Xbit_r35_c163 bl[163] br[163] wl[35] vdd gnd cell_6t
Xbit_r36_c163 bl[163] br[163] wl[36] vdd gnd cell_6t
Xbit_r37_c163 bl[163] br[163] wl[37] vdd gnd cell_6t
Xbit_r38_c163 bl[163] br[163] wl[38] vdd gnd cell_6t
Xbit_r39_c163 bl[163] br[163] wl[39] vdd gnd cell_6t
Xbit_r40_c163 bl[163] br[163] wl[40] vdd gnd cell_6t
Xbit_r41_c163 bl[163] br[163] wl[41] vdd gnd cell_6t
Xbit_r42_c163 bl[163] br[163] wl[42] vdd gnd cell_6t
Xbit_r43_c163 bl[163] br[163] wl[43] vdd gnd cell_6t
Xbit_r44_c163 bl[163] br[163] wl[44] vdd gnd cell_6t
Xbit_r45_c163 bl[163] br[163] wl[45] vdd gnd cell_6t
Xbit_r46_c163 bl[163] br[163] wl[46] vdd gnd cell_6t
Xbit_r47_c163 bl[163] br[163] wl[47] vdd gnd cell_6t
Xbit_r48_c163 bl[163] br[163] wl[48] vdd gnd cell_6t
Xbit_r49_c163 bl[163] br[163] wl[49] vdd gnd cell_6t
Xbit_r50_c163 bl[163] br[163] wl[50] vdd gnd cell_6t
Xbit_r51_c163 bl[163] br[163] wl[51] vdd gnd cell_6t
Xbit_r52_c163 bl[163] br[163] wl[52] vdd gnd cell_6t
Xbit_r53_c163 bl[163] br[163] wl[53] vdd gnd cell_6t
Xbit_r54_c163 bl[163] br[163] wl[54] vdd gnd cell_6t
Xbit_r55_c163 bl[163] br[163] wl[55] vdd gnd cell_6t
Xbit_r56_c163 bl[163] br[163] wl[56] vdd gnd cell_6t
Xbit_r57_c163 bl[163] br[163] wl[57] vdd gnd cell_6t
Xbit_r58_c163 bl[163] br[163] wl[58] vdd gnd cell_6t
Xbit_r59_c163 bl[163] br[163] wl[59] vdd gnd cell_6t
Xbit_r60_c163 bl[163] br[163] wl[60] vdd gnd cell_6t
Xbit_r61_c163 bl[163] br[163] wl[61] vdd gnd cell_6t
Xbit_r62_c163 bl[163] br[163] wl[62] vdd gnd cell_6t
Xbit_r63_c163 bl[163] br[163] wl[63] vdd gnd cell_6t
Xbit_r64_c163 bl[163] br[163] wl[64] vdd gnd cell_6t
Xbit_r65_c163 bl[163] br[163] wl[65] vdd gnd cell_6t
Xbit_r66_c163 bl[163] br[163] wl[66] vdd gnd cell_6t
Xbit_r67_c163 bl[163] br[163] wl[67] vdd gnd cell_6t
Xbit_r68_c163 bl[163] br[163] wl[68] vdd gnd cell_6t
Xbit_r69_c163 bl[163] br[163] wl[69] vdd gnd cell_6t
Xbit_r70_c163 bl[163] br[163] wl[70] vdd gnd cell_6t
Xbit_r71_c163 bl[163] br[163] wl[71] vdd gnd cell_6t
Xbit_r72_c163 bl[163] br[163] wl[72] vdd gnd cell_6t
Xbit_r73_c163 bl[163] br[163] wl[73] vdd gnd cell_6t
Xbit_r74_c163 bl[163] br[163] wl[74] vdd gnd cell_6t
Xbit_r75_c163 bl[163] br[163] wl[75] vdd gnd cell_6t
Xbit_r76_c163 bl[163] br[163] wl[76] vdd gnd cell_6t
Xbit_r77_c163 bl[163] br[163] wl[77] vdd gnd cell_6t
Xbit_r78_c163 bl[163] br[163] wl[78] vdd gnd cell_6t
Xbit_r79_c163 bl[163] br[163] wl[79] vdd gnd cell_6t
Xbit_r80_c163 bl[163] br[163] wl[80] vdd gnd cell_6t
Xbit_r81_c163 bl[163] br[163] wl[81] vdd gnd cell_6t
Xbit_r82_c163 bl[163] br[163] wl[82] vdd gnd cell_6t
Xbit_r83_c163 bl[163] br[163] wl[83] vdd gnd cell_6t
Xbit_r84_c163 bl[163] br[163] wl[84] vdd gnd cell_6t
Xbit_r85_c163 bl[163] br[163] wl[85] vdd gnd cell_6t
Xbit_r86_c163 bl[163] br[163] wl[86] vdd gnd cell_6t
Xbit_r87_c163 bl[163] br[163] wl[87] vdd gnd cell_6t
Xbit_r88_c163 bl[163] br[163] wl[88] vdd gnd cell_6t
Xbit_r89_c163 bl[163] br[163] wl[89] vdd gnd cell_6t
Xbit_r90_c163 bl[163] br[163] wl[90] vdd gnd cell_6t
Xbit_r91_c163 bl[163] br[163] wl[91] vdd gnd cell_6t
Xbit_r92_c163 bl[163] br[163] wl[92] vdd gnd cell_6t
Xbit_r93_c163 bl[163] br[163] wl[93] vdd gnd cell_6t
Xbit_r94_c163 bl[163] br[163] wl[94] vdd gnd cell_6t
Xbit_r95_c163 bl[163] br[163] wl[95] vdd gnd cell_6t
Xbit_r96_c163 bl[163] br[163] wl[96] vdd gnd cell_6t
Xbit_r97_c163 bl[163] br[163] wl[97] vdd gnd cell_6t
Xbit_r98_c163 bl[163] br[163] wl[98] vdd gnd cell_6t
Xbit_r99_c163 bl[163] br[163] wl[99] vdd gnd cell_6t
Xbit_r100_c163 bl[163] br[163] wl[100] vdd gnd cell_6t
Xbit_r101_c163 bl[163] br[163] wl[101] vdd gnd cell_6t
Xbit_r102_c163 bl[163] br[163] wl[102] vdd gnd cell_6t
Xbit_r103_c163 bl[163] br[163] wl[103] vdd gnd cell_6t
Xbit_r104_c163 bl[163] br[163] wl[104] vdd gnd cell_6t
Xbit_r105_c163 bl[163] br[163] wl[105] vdd gnd cell_6t
Xbit_r106_c163 bl[163] br[163] wl[106] vdd gnd cell_6t
Xbit_r107_c163 bl[163] br[163] wl[107] vdd gnd cell_6t
Xbit_r108_c163 bl[163] br[163] wl[108] vdd gnd cell_6t
Xbit_r109_c163 bl[163] br[163] wl[109] vdd gnd cell_6t
Xbit_r110_c163 bl[163] br[163] wl[110] vdd gnd cell_6t
Xbit_r111_c163 bl[163] br[163] wl[111] vdd gnd cell_6t
Xbit_r112_c163 bl[163] br[163] wl[112] vdd gnd cell_6t
Xbit_r113_c163 bl[163] br[163] wl[113] vdd gnd cell_6t
Xbit_r114_c163 bl[163] br[163] wl[114] vdd gnd cell_6t
Xbit_r115_c163 bl[163] br[163] wl[115] vdd gnd cell_6t
Xbit_r116_c163 bl[163] br[163] wl[116] vdd gnd cell_6t
Xbit_r117_c163 bl[163] br[163] wl[117] vdd gnd cell_6t
Xbit_r118_c163 bl[163] br[163] wl[118] vdd gnd cell_6t
Xbit_r119_c163 bl[163] br[163] wl[119] vdd gnd cell_6t
Xbit_r120_c163 bl[163] br[163] wl[120] vdd gnd cell_6t
Xbit_r121_c163 bl[163] br[163] wl[121] vdd gnd cell_6t
Xbit_r122_c163 bl[163] br[163] wl[122] vdd gnd cell_6t
Xbit_r123_c163 bl[163] br[163] wl[123] vdd gnd cell_6t
Xbit_r124_c163 bl[163] br[163] wl[124] vdd gnd cell_6t
Xbit_r125_c163 bl[163] br[163] wl[125] vdd gnd cell_6t
Xbit_r126_c163 bl[163] br[163] wl[126] vdd gnd cell_6t
Xbit_r127_c163 bl[163] br[163] wl[127] vdd gnd cell_6t
Xbit_r0_c164 bl[164] br[164] wl[0] vdd gnd cell_6t
Xbit_r1_c164 bl[164] br[164] wl[1] vdd gnd cell_6t
Xbit_r2_c164 bl[164] br[164] wl[2] vdd gnd cell_6t
Xbit_r3_c164 bl[164] br[164] wl[3] vdd gnd cell_6t
Xbit_r4_c164 bl[164] br[164] wl[4] vdd gnd cell_6t
Xbit_r5_c164 bl[164] br[164] wl[5] vdd gnd cell_6t
Xbit_r6_c164 bl[164] br[164] wl[6] vdd gnd cell_6t
Xbit_r7_c164 bl[164] br[164] wl[7] vdd gnd cell_6t
Xbit_r8_c164 bl[164] br[164] wl[8] vdd gnd cell_6t
Xbit_r9_c164 bl[164] br[164] wl[9] vdd gnd cell_6t
Xbit_r10_c164 bl[164] br[164] wl[10] vdd gnd cell_6t
Xbit_r11_c164 bl[164] br[164] wl[11] vdd gnd cell_6t
Xbit_r12_c164 bl[164] br[164] wl[12] vdd gnd cell_6t
Xbit_r13_c164 bl[164] br[164] wl[13] vdd gnd cell_6t
Xbit_r14_c164 bl[164] br[164] wl[14] vdd gnd cell_6t
Xbit_r15_c164 bl[164] br[164] wl[15] vdd gnd cell_6t
Xbit_r16_c164 bl[164] br[164] wl[16] vdd gnd cell_6t
Xbit_r17_c164 bl[164] br[164] wl[17] vdd gnd cell_6t
Xbit_r18_c164 bl[164] br[164] wl[18] vdd gnd cell_6t
Xbit_r19_c164 bl[164] br[164] wl[19] vdd gnd cell_6t
Xbit_r20_c164 bl[164] br[164] wl[20] vdd gnd cell_6t
Xbit_r21_c164 bl[164] br[164] wl[21] vdd gnd cell_6t
Xbit_r22_c164 bl[164] br[164] wl[22] vdd gnd cell_6t
Xbit_r23_c164 bl[164] br[164] wl[23] vdd gnd cell_6t
Xbit_r24_c164 bl[164] br[164] wl[24] vdd gnd cell_6t
Xbit_r25_c164 bl[164] br[164] wl[25] vdd gnd cell_6t
Xbit_r26_c164 bl[164] br[164] wl[26] vdd gnd cell_6t
Xbit_r27_c164 bl[164] br[164] wl[27] vdd gnd cell_6t
Xbit_r28_c164 bl[164] br[164] wl[28] vdd gnd cell_6t
Xbit_r29_c164 bl[164] br[164] wl[29] vdd gnd cell_6t
Xbit_r30_c164 bl[164] br[164] wl[30] vdd gnd cell_6t
Xbit_r31_c164 bl[164] br[164] wl[31] vdd gnd cell_6t
Xbit_r32_c164 bl[164] br[164] wl[32] vdd gnd cell_6t
Xbit_r33_c164 bl[164] br[164] wl[33] vdd gnd cell_6t
Xbit_r34_c164 bl[164] br[164] wl[34] vdd gnd cell_6t
Xbit_r35_c164 bl[164] br[164] wl[35] vdd gnd cell_6t
Xbit_r36_c164 bl[164] br[164] wl[36] vdd gnd cell_6t
Xbit_r37_c164 bl[164] br[164] wl[37] vdd gnd cell_6t
Xbit_r38_c164 bl[164] br[164] wl[38] vdd gnd cell_6t
Xbit_r39_c164 bl[164] br[164] wl[39] vdd gnd cell_6t
Xbit_r40_c164 bl[164] br[164] wl[40] vdd gnd cell_6t
Xbit_r41_c164 bl[164] br[164] wl[41] vdd gnd cell_6t
Xbit_r42_c164 bl[164] br[164] wl[42] vdd gnd cell_6t
Xbit_r43_c164 bl[164] br[164] wl[43] vdd gnd cell_6t
Xbit_r44_c164 bl[164] br[164] wl[44] vdd gnd cell_6t
Xbit_r45_c164 bl[164] br[164] wl[45] vdd gnd cell_6t
Xbit_r46_c164 bl[164] br[164] wl[46] vdd gnd cell_6t
Xbit_r47_c164 bl[164] br[164] wl[47] vdd gnd cell_6t
Xbit_r48_c164 bl[164] br[164] wl[48] vdd gnd cell_6t
Xbit_r49_c164 bl[164] br[164] wl[49] vdd gnd cell_6t
Xbit_r50_c164 bl[164] br[164] wl[50] vdd gnd cell_6t
Xbit_r51_c164 bl[164] br[164] wl[51] vdd gnd cell_6t
Xbit_r52_c164 bl[164] br[164] wl[52] vdd gnd cell_6t
Xbit_r53_c164 bl[164] br[164] wl[53] vdd gnd cell_6t
Xbit_r54_c164 bl[164] br[164] wl[54] vdd gnd cell_6t
Xbit_r55_c164 bl[164] br[164] wl[55] vdd gnd cell_6t
Xbit_r56_c164 bl[164] br[164] wl[56] vdd gnd cell_6t
Xbit_r57_c164 bl[164] br[164] wl[57] vdd gnd cell_6t
Xbit_r58_c164 bl[164] br[164] wl[58] vdd gnd cell_6t
Xbit_r59_c164 bl[164] br[164] wl[59] vdd gnd cell_6t
Xbit_r60_c164 bl[164] br[164] wl[60] vdd gnd cell_6t
Xbit_r61_c164 bl[164] br[164] wl[61] vdd gnd cell_6t
Xbit_r62_c164 bl[164] br[164] wl[62] vdd gnd cell_6t
Xbit_r63_c164 bl[164] br[164] wl[63] vdd gnd cell_6t
Xbit_r64_c164 bl[164] br[164] wl[64] vdd gnd cell_6t
Xbit_r65_c164 bl[164] br[164] wl[65] vdd gnd cell_6t
Xbit_r66_c164 bl[164] br[164] wl[66] vdd gnd cell_6t
Xbit_r67_c164 bl[164] br[164] wl[67] vdd gnd cell_6t
Xbit_r68_c164 bl[164] br[164] wl[68] vdd gnd cell_6t
Xbit_r69_c164 bl[164] br[164] wl[69] vdd gnd cell_6t
Xbit_r70_c164 bl[164] br[164] wl[70] vdd gnd cell_6t
Xbit_r71_c164 bl[164] br[164] wl[71] vdd gnd cell_6t
Xbit_r72_c164 bl[164] br[164] wl[72] vdd gnd cell_6t
Xbit_r73_c164 bl[164] br[164] wl[73] vdd gnd cell_6t
Xbit_r74_c164 bl[164] br[164] wl[74] vdd gnd cell_6t
Xbit_r75_c164 bl[164] br[164] wl[75] vdd gnd cell_6t
Xbit_r76_c164 bl[164] br[164] wl[76] vdd gnd cell_6t
Xbit_r77_c164 bl[164] br[164] wl[77] vdd gnd cell_6t
Xbit_r78_c164 bl[164] br[164] wl[78] vdd gnd cell_6t
Xbit_r79_c164 bl[164] br[164] wl[79] vdd gnd cell_6t
Xbit_r80_c164 bl[164] br[164] wl[80] vdd gnd cell_6t
Xbit_r81_c164 bl[164] br[164] wl[81] vdd gnd cell_6t
Xbit_r82_c164 bl[164] br[164] wl[82] vdd gnd cell_6t
Xbit_r83_c164 bl[164] br[164] wl[83] vdd gnd cell_6t
Xbit_r84_c164 bl[164] br[164] wl[84] vdd gnd cell_6t
Xbit_r85_c164 bl[164] br[164] wl[85] vdd gnd cell_6t
Xbit_r86_c164 bl[164] br[164] wl[86] vdd gnd cell_6t
Xbit_r87_c164 bl[164] br[164] wl[87] vdd gnd cell_6t
Xbit_r88_c164 bl[164] br[164] wl[88] vdd gnd cell_6t
Xbit_r89_c164 bl[164] br[164] wl[89] vdd gnd cell_6t
Xbit_r90_c164 bl[164] br[164] wl[90] vdd gnd cell_6t
Xbit_r91_c164 bl[164] br[164] wl[91] vdd gnd cell_6t
Xbit_r92_c164 bl[164] br[164] wl[92] vdd gnd cell_6t
Xbit_r93_c164 bl[164] br[164] wl[93] vdd gnd cell_6t
Xbit_r94_c164 bl[164] br[164] wl[94] vdd gnd cell_6t
Xbit_r95_c164 bl[164] br[164] wl[95] vdd gnd cell_6t
Xbit_r96_c164 bl[164] br[164] wl[96] vdd gnd cell_6t
Xbit_r97_c164 bl[164] br[164] wl[97] vdd gnd cell_6t
Xbit_r98_c164 bl[164] br[164] wl[98] vdd gnd cell_6t
Xbit_r99_c164 bl[164] br[164] wl[99] vdd gnd cell_6t
Xbit_r100_c164 bl[164] br[164] wl[100] vdd gnd cell_6t
Xbit_r101_c164 bl[164] br[164] wl[101] vdd gnd cell_6t
Xbit_r102_c164 bl[164] br[164] wl[102] vdd gnd cell_6t
Xbit_r103_c164 bl[164] br[164] wl[103] vdd gnd cell_6t
Xbit_r104_c164 bl[164] br[164] wl[104] vdd gnd cell_6t
Xbit_r105_c164 bl[164] br[164] wl[105] vdd gnd cell_6t
Xbit_r106_c164 bl[164] br[164] wl[106] vdd gnd cell_6t
Xbit_r107_c164 bl[164] br[164] wl[107] vdd gnd cell_6t
Xbit_r108_c164 bl[164] br[164] wl[108] vdd gnd cell_6t
Xbit_r109_c164 bl[164] br[164] wl[109] vdd gnd cell_6t
Xbit_r110_c164 bl[164] br[164] wl[110] vdd gnd cell_6t
Xbit_r111_c164 bl[164] br[164] wl[111] vdd gnd cell_6t
Xbit_r112_c164 bl[164] br[164] wl[112] vdd gnd cell_6t
Xbit_r113_c164 bl[164] br[164] wl[113] vdd gnd cell_6t
Xbit_r114_c164 bl[164] br[164] wl[114] vdd gnd cell_6t
Xbit_r115_c164 bl[164] br[164] wl[115] vdd gnd cell_6t
Xbit_r116_c164 bl[164] br[164] wl[116] vdd gnd cell_6t
Xbit_r117_c164 bl[164] br[164] wl[117] vdd gnd cell_6t
Xbit_r118_c164 bl[164] br[164] wl[118] vdd gnd cell_6t
Xbit_r119_c164 bl[164] br[164] wl[119] vdd gnd cell_6t
Xbit_r120_c164 bl[164] br[164] wl[120] vdd gnd cell_6t
Xbit_r121_c164 bl[164] br[164] wl[121] vdd gnd cell_6t
Xbit_r122_c164 bl[164] br[164] wl[122] vdd gnd cell_6t
Xbit_r123_c164 bl[164] br[164] wl[123] vdd gnd cell_6t
Xbit_r124_c164 bl[164] br[164] wl[124] vdd gnd cell_6t
Xbit_r125_c164 bl[164] br[164] wl[125] vdd gnd cell_6t
Xbit_r126_c164 bl[164] br[164] wl[126] vdd gnd cell_6t
Xbit_r127_c164 bl[164] br[164] wl[127] vdd gnd cell_6t
Xbit_r0_c165 bl[165] br[165] wl[0] vdd gnd cell_6t
Xbit_r1_c165 bl[165] br[165] wl[1] vdd gnd cell_6t
Xbit_r2_c165 bl[165] br[165] wl[2] vdd gnd cell_6t
Xbit_r3_c165 bl[165] br[165] wl[3] vdd gnd cell_6t
Xbit_r4_c165 bl[165] br[165] wl[4] vdd gnd cell_6t
Xbit_r5_c165 bl[165] br[165] wl[5] vdd gnd cell_6t
Xbit_r6_c165 bl[165] br[165] wl[6] vdd gnd cell_6t
Xbit_r7_c165 bl[165] br[165] wl[7] vdd gnd cell_6t
Xbit_r8_c165 bl[165] br[165] wl[8] vdd gnd cell_6t
Xbit_r9_c165 bl[165] br[165] wl[9] vdd gnd cell_6t
Xbit_r10_c165 bl[165] br[165] wl[10] vdd gnd cell_6t
Xbit_r11_c165 bl[165] br[165] wl[11] vdd gnd cell_6t
Xbit_r12_c165 bl[165] br[165] wl[12] vdd gnd cell_6t
Xbit_r13_c165 bl[165] br[165] wl[13] vdd gnd cell_6t
Xbit_r14_c165 bl[165] br[165] wl[14] vdd gnd cell_6t
Xbit_r15_c165 bl[165] br[165] wl[15] vdd gnd cell_6t
Xbit_r16_c165 bl[165] br[165] wl[16] vdd gnd cell_6t
Xbit_r17_c165 bl[165] br[165] wl[17] vdd gnd cell_6t
Xbit_r18_c165 bl[165] br[165] wl[18] vdd gnd cell_6t
Xbit_r19_c165 bl[165] br[165] wl[19] vdd gnd cell_6t
Xbit_r20_c165 bl[165] br[165] wl[20] vdd gnd cell_6t
Xbit_r21_c165 bl[165] br[165] wl[21] vdd gnd cell_6t
Xbit_r22_c165 bl[165] br[165] wl[22] vdd gnd cell_6t
Xbit_r23_c165 bl[165] br[165] wl[23] vdd gnd cell_6t
Xbit_r24_c165 bl[165] br[165] wl[24] vdd gnd cell_6t
Xbit_r25_c165 bl[165] br[165] wl[25] vdd gnd cell_6t
Xbit_r26_c165 bl[165] br[165] wl[26] vdd gnd cell_6t
Xbit_r27_c165 bl[165] br[165] wl[27] vdd gnd cell_6t
Xbit_r28_c165 bl[165] br[165] wl[28] vdd gnd cell_6t
Xbit_r29_c165 bl[165] br[165] wl[29] vdd gnd cell_6t
Xbit_r30_c165 bl[165] br[165] wl[30] vdd gnd cell_6t
Xbit_r31_c165 bl[165] br[165] wl[31] vdd gnd cell_6t
Xbit_r32_c165 bl[165] br[165] wl[32] vdd gnd cell_6t
Xbit_r33_c165 bl[165] br[165] wl[33] vdd gnd cell_6t
Xbit_r34_c165 bl[165] br[165] wl[34] vdd gnd cell_6t
Xbit_r35_c165 bl[165] br[165] wl[35] vdd gnd cell_6t
Xbit_r36_c165 bl[165] br[165] wl[36] vdd gnd cell_6t
Xbit_r37_c165 bl[165] br[165] wl[37] vdd gnd cell_6t
Xbit_r38_c165 bl[165] br[165] wl[38] vdd gnd cell_6t
Xbit_r39_c165 bl[165] br[165] wl[39] vdd gnd cell_6t
Xbit_r40_c165 bl[165] br[165] wl[40] vdd gnd cell_6t
Xbit_r41_c165 bl[165] br[165] wl[41] vdd gnd cell_6t
Xbit_r42_c165 bl[165] br[165] wl[42] vdd gnd cell_6t
Xbit_r43_c165 bl[165] br[165] wl[43] vdd gnd cell_6t
Xbit_r44_c165 bl[165] br[165] wl[44] vdd gnd cell_6t
Xbit_r45_c165 bl[165] br[165] wl[45] vdd gnd cell_6t
Xbit_r46_c165 bl[165] br[165] wl[46] vdd gnd cell_6t
Xbit_r47_c165 bl[165] br[165] wl[47] vdd gnd cell_6t
Xbit_r48_c165 bl[165] br[165] wl[48] vdd gnd cell_6t
Xbit_r49_c165 bl[165] br[165] wl[49] vdd gnd cell_6t
Xbit_r50_c165 bl[165] br[165] wl[50] vdd gnd cell_6t
Xbit_r51_c165 bl[165] br[165] wl[51] vdd gnd cell_6t
Xbit_r52_c165 bl[165] br[165] wl[52] vdd gnd cell_6t
Xbit_r53_c165 bl[165] br[165] wl[53] vdd gnd cell_6t
Xbit_r54_c165 bl[165] br[165] wl[54] vdd gnd cell_6t
Xbit_r55_c165 bl[165] br[165] wl[55] vdd gnd cell_6t
Xbit_r56_c165 bl[165] br[165] wl[56] vdd gnd cell_6t
Xbit_r57_c165 bl[165] br[165] wl[57] vdd gnd cell_6t
Xbit_r58_c165 bl[165] br[165] wl[58] vdd gnd cell_6t
Xbit_r59_c165 bl[165] br[165] wl[59] vdd gnd cell_6t
Xbit_r60_c165 bl[165] br[165] wl[60] vdd gnd cell_6t
Xbit_r61_c165 bl[165] br[165] wl[61] vdd gnd cell_6t
Xbit_r62_c165 bl[165] br[165] wl[62] vdd gnd cell_6t
Xbit_r63_c165 bl[165] br[165] wl[63] vdd gnd cell_6t
Xbit_r64_c165 bl[165] br[165] wl[64] vdd gnd cell_6t
Xbit_r65_c165 bl[165] br[165] wl[65] vdd gnd cell_6t
Xbit_r66_c165 bl[165] br[165] wl[66] vdd gnd cell_6t
Xbit_r67_c165 bl[165] br[165] wl[67] vdd gnd cell_6t
Xbit_r68_c165 bl[165] br[165] wl[68] vdd gnd cell_6t
Xbit_r69_c165 bl[165] br[165] wl[69] vdd gnd cell_6t
Xbit_r70_c165 bl[165] br[165] wl[70] vdd gnd cell_6t
Xbit_r71_c165 bl[165] br[165] wl[71] vdd gnd cell_6t
Xbit_r72_c165 bl[165] br[165] wl[72] vdd gnd cell_6t
Xbit_r73_c165 bl[165] br[165] wl[73] vdd gnd cell_6t
Xbit_r74_c165 bl[165] br[165] wl[74] vdd gnd cell_6t
Xbit_r75_c165 bl[165] br[165] wl[75] vdd gnd cell_6t
Xbit_r76_c165 bl[165] br[165] wl[76] vdd gnd cell_6t
Xbit_r77_c165 bl[165] br[165] wl[77] vdd gnd cell_6t
Xbit_r78_c165 bl[165] br[165] wl[78] vdd gnd cell_6t
Xbit_r79_c165 bl[165] br[165] wl[79] vdd gnd cell_6t
Xbit_r80_c165 bl[165] br[165] wl[80] vdd gnd cell_6t
Xbit_r81_c165 bl[165] br[165] wl[81] vdd gnd cell_6t
Xbit_r82_c165 bl[165] br[165] wl[82] vdd gnd cell_6t
Xbit_r83_c165 bl[165] br[165] wl[83] vdd gnd cell_6t
Xbit_r84_c165 bl[165] br[165] wl[84] vdd gnd cell_6t
Xbit_r85_c165 bl[165] br[165] wl[85] vdd gnd cell_6t
Xbit_r86_c165 bl[165] br[165] wl[86] vdd gnd cell_6t
Xbit_r87_c165 bl[165] br[165] wl[87] vdd gnd cell_6t
Xbit_r88_c165 bl[165] br[165] wl[88] vdd gnd cell_6t
Xbit_r89_c165 bl[165] br[165] wl[89] vdd gnd cell_6t
Xbit_r90_c165 bl[165] br[165] wl[90] vdd gnd cell_6t
Xbit_r91_c165 bl[165] br[165] wl[91] vdd gnd cell_6t
Xbit_r92_c165 bl[165] br[165] wl[92] vdd gnd cell_6t
Xbit_r93_c165 bl[165] br[165] wl[93] vdd gnd cell_6t
Xbit_r94_c165 bl[165] br[165] wl[94] vdd gnd cell_6t
Xbit_r95_c165 bl[165] br[165] wl[95] vdd gnd cell_6t
Xbit_r96_c165 bl[165] br[165] wl[96] vdd gnd cell_6t
Xbit_r97_c165 bl[165] br[165] wl[97] vdd gnd cell_6t
Xbit_r98_c165 bl[165] br[165] wl[98] vdd gnd cell_6t
Xbit_r99_c165 bl[165] br[165] wl[99] vdd gnd cell_6t
Xbit_r100_c165 bl[165] br[165] wl[100] vdd gnd cell_6t
Xbit_r101_c165 bl[165] br[165] wl[101] vdd gnd cell_6t
Xbit_r102_c165 bl[165] br[165] wl[102] vdd gnd cell_6t
Xbit_r103_c165 bl[165] br[165] wl[103] vdd gnd cell_6t
Xbit_r104_c165 bl[165] br[165] wl[104] vdd gnd cell_6t
Xbit_r105_c165 bl[165] br[165] wl[105] vdd gnd cell_6t
Xbit_r106_c165 bl[165] br[165] wl[106] vdd gnd cell_6t
Xbit_r107_c165 bl[165] br[165] wl[107] vdd gnd cell_6t
Xbit_r108_c165 bl[165] br[165] wl[108] vdd gnd cell_6t
Xbit_r109_c165 bl[165] br[165] wl[109] vdd gnd cell_6t
Xbit_r110_c165 bl[165] br[165] wl[110] vdd gnd cell_6t
Xbit_r111_c165 bl[165] br[165] wl[111] vdd gnd cell_6t
Xbit_r112_c165 bl[165] br[165] wl[112] vdd gnd cell_6t
Xbit_r113_c165 bl[165] br[165] wl[113] vdd gnd cell_6t
Xbit_r114_c165 bl[165] br[165] wl[114] vdd gnd cell_6t
Xbit_r115_c165 bl[165] br[165] wl[115] vdd gnd cell_6t
Xbit_r116_c165 bl[165] br[165] wl[116] vdd gnd cell_6t
Xbit_r117_c165 bl[165] br[165] wl[117] vdd gnd cell_6t
Xbit_r118_c165 bl[165] br[165] wl[118] vdd gnd cell_6t
Xbit_r119_c165 bl[165] br[165] wl[119] vdd gnd cell_6t
Xbit_r120_c165 bl[165] br[165] wl[120] vdd gnd cell_6t
Xbit_r121_c165 bl[165] br[165] wl[121] vdd gnd cell_6t
Xbit_r122_c165 bl[165] br[165] wl[122] vdd gnd cell_6t
Xbit_r123_c165 bl[165] br[165] wl[123] vdd gnd cell_6t
Xbit_r124_c165 bl[165] br[165] wl[124] vdd gnd cell_6t
Xbit_r125_c165 bl[165] br[165] wl[125] vdd gnd cell_6t
Xbit_r126_c165 bl[165] br[165] wl[126] vdd gnd cell_6t
Xbit_r127_c165 bl[165] br[165] wl[127] vdd gnd cell_6t
Xbit_r0_c166 bl[166] br[166] wl[0] vdd gnd cell_6t
Xbit_r1_c166 bl[166] br[166] wl[1] vdd gnd cell_6t
Xbit_r2_c166 bl[166] br[166] wl[2] vdd gnd cell_6t
Xbit_r3_c166 bl[166] br[166] wl[3] vdd gnd cell_6t
Xbit_r4_c166 bl[166] br[166] wl[4] vdd gnd cell_6t
Xbit_r5_c166 bl[166] br[166] wl[5] vdd gnd cell_6t
Xbit_r6_c166 bl[166] br[166] wl[6] vdd gnd cell_6t
Xbit_r7_c166 bl[166] br[166] wl[7] vdd gnd cell_6t
Xbit_r8_c166 bl[166] br[166] wl[8] vdd gnd cell_6t
Xbit_r9_c166 bl[166] br[166] wl[9] vdd gnd cell_6t
Xbit_r10_c166 bl[166] br[166] wl[10] vdd gnd cell_6t
Xbit_r11_c166 bl[166] br[166] wl[11] vdd gnd cell_6t
Xbit_r12_c166 bl[166] br[166] wl[12] vdd gnd cell_6t
Xbit_r13_c166 bl[166] br[166] wl[13] vdd gnd cell_6t
Xbit_r14_c166 bl[166] br[166] wl[14] vdd gnd cell_6t
Xbit_r15_c166 bl[166] br[166] wl[15] vdd gnd cell_6t
Xbit_r16_c166 bl[166] br[166] wl[16] vdd gnd cell_6t
Xbit_r17_c166 bl[166] br[166] wl[17] vdd gnd cell_6t
Xbit_r18_c166 bl[166] br[166] wl[18] vdd gnd cell_6t
Xbit_r19_c166 bl[166] br[166] wl[19] vdd gnd cell_6t
Xbit_r20_c166 bl[166] br[166] wl[20] vdd gnd cell_6t
Xbit_r21_c166 bl[166] br[166] wl[21] vdd gnd cell_6t
Xbit_r22_c166 bl[166] br[166] wl[22] vdd gnd cell_6t
Xbit_r23_c166 bl[166] br[166] wl[23] vdd gnd cell_6t
Xbit_r24_c166 bl[166] br[166] wl[24] vdd gnd cell_6t
Xbit_r25_c166 bl[166] br[166] wl[25] vdd gnd cell_6t
Xbit_r26_c166 bl[166] br[166] wl[26] vdd gnd cell_6t
Xbit_r27_c166 bl[166] br[166] wl[27] vdd gnd cell_6t
Xbit_r28_c166 bl[166] br[166] wl[28] vdd gnd cell_6t
Xbit_r29_c166 bl[166] br[166] wl[29] vdd gnd cell_6t
Xbit_r30_c166 bl[166] br[166] wl[30] vdd gnd cell_6t
Xbit_r31_c166 bl[166] br[166] wl[31] vdd gnd cell_6t
Xbit_r32_c166 bl[166] br[166] wl[32] vdd gnd cell_6t
Xbit_r33_c166 bl[166] br[166] wl[33] vdd gnd cell_6t
Xbit_r34_c166 bl[166] br[166] wl[34] vdd gnd cell_6t
Xbit_r35_c166 bl[166] br[166] wl[35] vdd gnd cell_6t
Xbit_r36_c166 bl[166] br[166] wl[36] vdd gnd cell_6t
Xbit_r37_c166 bl[166] br[166] wl[37] vdd gnd cell_6t
Xbit_r38_c166 bl[166] br[166] wl[38] vdd gnd cell_6t
Xbit_r39_c166 bl[166] br[166] wl[39] vdd gnd cell_6t
Xbit_r40_c166 bl[166] br[166] wl[40] vdd gnd cell_6t
Xbit_r41_c166 bl[166] br[166] wl[41] vdd gnd cell_6t
Xbit_r42_c166 bl[166] br[166] wl[42] vdd gnd cell_6t
Xbit_r43_c166 bl[166] br[166] wl[43] vdd gnd cell_6t
Xbit_r44_c166 bl[166] br[166] wl[44] vdd gnd cell_6t
Xbit_r45_c166 bl[166] br[166] wl[45] vdd gnd cell_6t
Xbit_r46_c166 bl[166] br[166] wl[46] vdd gnd cell_6t
Xbit_r47_c166 bl[166] br[166] wl[47] vdd gnd cell_6t
Xbit_r48_c166 bl[166] br[166] wl[48] vdd gnd cell_6t
Xbit_r49_c166 bl[166] br[166] wl[49] vdd gnd cell_6t
Xbit_r50_c166 bl[166] br[166] wl[50] vdd gnd cell_6t
Xbit_r51_c166 bl[166] br[166] wl[51] vdd gnd cell_6t
Xbit_r52_c166 bl[166] br[166] wl[52] vdd gnd cell_6t
Xbit_r53_c166 bl[166] br[166] wl[53] vdd gnd cell_6t
Xbit_r54_c166 bl[166] br[166] wl[54] vdd gnd cell_6t
Xbit_r55_c166 bl[166] br[166] wl[55] vdd gnd cell_6t
Xbit_r56_c166 bl[166] br[166] wl[56] vdd gnd cell_6t
Xbit_r57_c166 bl[166] br[166] wl[57] vdd gnd cell_6t
Xbit_r58_c166 bl[166] br[166] wl[58] vdd gnd cell_6t
Xbit_r59_c166 bl[166] br[166] wl[59] vdd gnd cell_6t
Xbit_r60_c166 bl[166] br[166] wl[60] vdd gnd cell_6t
Xbit_r61_c166 bl[166] br[166] wl[61] vdd gnd cell_6t
Xbit_r62_c166 bl[166] br[166] wl[62] vdd gnd cell_6t
Xbit_r63_c166 bl[166] br[166] wl[63] vdd gnd cell_6t
Xbit_r64_c166 bl[166] br[166] wl[64] vdd gnd cell_6t
Xbit_r65_c166 bl[166] br[166] wl[65] vdd gnd cell_6t
Xbit_r66_c166 bl[166] br[166] wl[66] vdd gnd cell_6t
Xbit_r67_c166 bl[166] br[166] wl[67] vdd gnd cell_6t
Xbit_r68_c166 bl[166] br[166] wl[68] vdd gnd cell_6t
Xbit_r69_c166 bl[166] br[166] wl[69] vdd gnd cell_6t
Xbit_r70_c166 bl[166] br[166] wl[70] vdd gnd cell_6t
Xbit_r71_c166 bl[166] br[166] wl[71] vdd gnd cell_6t
Xbit_r72_c166 bl[166] br[166] wl[72] vdd gnd cell_6t
Xbit_r73_c166 bl[166] br[166] wl[73] vdd gnd cell_6t
Xbit_r74_c166 bl[166] br[166] wl[74] vdd gnd cell_6t
Xbit_r75_c166 bl[166] br[166] wl[75] vdd gnd cell_6t
Xbit_r76_c166 bl[166] br[166] wl[76] vdd gnd cell_6t
Xbit_r77_c166 bl[166] br[166] wl[77] vdd gnd cell_6t
Xbit_r78_c166 bl[166] br[166] wl[78] vdd gnd cell_6t
Xbit_r79_c166 bl[166] br[166] wl[79] vdd gnd cell_6t
Xbit_r80_c166 bl[166] br[166] wl[80] vdd gnd cell_6t
Xbit_r81_c166 bl[166] br[166] wl[81] vdd gnd cell_6t
Xbit_r82_c166 bl[166] br[166] wl[82] vdd gnd cell_6t
Xbit_r83_c166 bl[166] br[166] wl[83] vdd gnd cell_6t
Xbit_r84_c166 bl[166] br[166] wl[84] vdd gnd cell_6t
Xbit_r85_c166 bl[166] br[166] wl[85] vdd gnd cell_6t
Xbit_r86_c166 bl[166] br[166] wl[86] vdd gnd cell_6t
Xbit_r87_c166 bl[166] br[166] wl[87] vdd gnd cell_6t
Xbit_r88_c166 bl[166] br[166] wl[88] vdd gnd cell_6t
Xbit_r89_c166 bl[166] br[166] wl[89] vdd gnd cell_6t
Xbit_r90_c166 bl[166] br[166] wl[90] vdd gnd cell_6t
Xbit_r91_c166 bl[166] br[166] wl[91] vdd gnd cell_6t
Xbit_r92_c166 bl[166] br[166] wl[92] vdd gnd cell_6t
Xbit_r93_c166 bl[166] br[166] wl[93] vdd gnd cell_6t
Xbit_r94_c166 bl[166] br[166] wl[94] vdd gnd cell_6t
Xbit_r95_c166 bl[166] br[166] wl[95] vdd gnd cell_6t
Xbit_r96_c166 bl[166] br[166] wl[96] vdd gnd cell_6t
Xbit_r97_c166 bl[166] br[166] wl[97] vdd gnd cell_6t
Xbit_r98_c166 bl[166] br[166] wl[98] vdd gnd cell_6t
Xbit_r99_c166 bl[166] br[166] wl[99] vdd gnd cell_6t
Xbit_r100_c166 bl[166] br[166] wl[100] vdd gnd cell_6t
Xbit_r101_c166 bl[166] br[166] wl[101] vdd gnd cell_6t
Xbit_r102_c166 bl[166] br[166] wl[102] vdd gnd cell_6t
Xbit_r103_c166 bl[166] br[166] wl[103] vdd gnd cell_6t
Xbit_r104_c166 bl[166] br[166] wl[104] vdd gnd cell_6t
Xbit_r105_c166 bl[166] br[166] wl[105] vdd gnd cell_6t
Xbit_r106_c166 bl[166] br[166] wl[106] vdd gnd cell_6t
Xbit_r107_c166 bl[166] br[166] wl[107] vdd gnd cell_6t
Xbit_r108_c166 bl[166] br[166] wl[108] vdd gnd cell_6t
Xbit_r109_c166 bl[166] br[166] wl[109] vdd gnd cell_6t
Xbit_r110_c166 bl[166] br[166] wl[110] vdd gnd cell_6t
Xbit_r111_c166 bl[166] br[166] wl[111] vdd gnd cell_6t
Xbit_r112_c166 bl[166] br[166] wl[112] vdd gnd cell_6t
Xbit_r113_c166 bl[166] br[166] wl[113] vdd gnd cell_6t
Xbit_r114_c166 bl[166] br[166] wl[114] vdd gnd cell_6t
Xbit_r115_c166 bl[166] br[166] wl[115] vdd gnd cell_6t
Xbit_r116_c166 bl[166] br[166] wl[116] vdd gnd cell_6t
Xbit_r117_c166 bl[166] br[166] wl[117] vdd gnd cell_6t
Xbit_r118_c166 bl[166] br[166] wl[118] vdd gnd cell_6t
Xbit_r119_c166 bl[166] br[166] wl[119] vdd gnd cell_6t
Xbit_r120_c166 bl[166] br[166] wl[120] vdd gnd cell_6t
Xbit_r121_c166 bl[166] br[166] wl[121] vdd gnd cell_6t
Xbit_r122_c166 bl[166] br[166] wl[122] vdd gnd cell_6t
Xbit_r123_c166 bl[166] br[166] wl[123] vdd gnd cell_6t
Xbit_r124_c166 bl[166] br[166] wl[124] vdd gnd cell_6t
Xbit_r125_c166 bl[166] br[166] wl[125] vdd gnd cell_6t
Xbit_r126_c166 bl[166] br[166] wl[126] vdd gnd cell_6t
Xbit_r127_c166 bl[166] br[166] wl[127] vdd gnd cell_6t
Xbit_r0_c167 bl[167] br[167] wl[0] vdd gnd cell_6t
Xbit_r1_c167 bl[167] br[167] wl[1] vdd gnd cell_6t
Xbit_r2_c167 bl[167] br[167] wl[2] vdd gnd cell_6t
Xbit_r3_c167 bl[167] br[167] wl[3] vdd gnd cell_6t
Xbit_r4_c167 bl[167] br[167] wl[4] vdd gnd cell_6t
Xbit_r5_c167 bl[167] br[167] wl[5] vdd gnd cell_6t
Xbit_r6_c167 bl[167] br[167] wl[6] vdd gnd cell_6t
Xbit_r7_c167 bl[167] br[167] wl[7] vdd gnd cell_6t
Xbit_r8_c167 bl[167] br[167] wl[8] vdd gnd cell_6t
Xbit_r9_c167 bl[167] br[167] wl[9] vdd gnd cell_6t
Xbit_r10_c167 bl[167] br[167] wl[10] vdd gnd cell_6t
Xbit_r11_c167 bl[167] br[167] wl[11] vdd gnd cell_6t
Xbit_r12_c167 bl[167] br[167] wl[12] vdd gnd cell_6t
Xbit_r13_c167 bl[167] br[167] wl[13] vdd gnd cell_6t
Xbit_r14_c167 bl[167] br[167] wl[14] vdd gnd cell_6t
Xbit_r15_c167 bl[167] br[167] wl[15] vdd gnd cell_6t
Xbit_r16_c167 bl[167] br[167] wl[16] vdd gnd cell_6t
Xbit_r17_c167 bl[167] br[167] wl[17] vdd gnd cell_6t
Xbit_r18_c167 bl[167] br[167] wl[18] vdd gnd cell_6t
Xbit_r19_c167 bl[167] br[167] wl[19] vdd gnd cell_6t
Xbit_r20_c167 bl[167] br[167] wl[20] vdd gnd cell_6t
Xbit_r21_c167 bl[167] br[167] wl[21] vdd gnd cell_6t
Xbit_r22_c167 bl[167] br[167] wl[22] vdd gnd cell_6t
Xbit_r23_c167 bl[167] br[167] wl[23] vdd gnd cell_6t
Xbit_r24_c167 bl[167] br[167] wl[24] vdd gnd cell_6t
Xbit_r25_c167 bl[167] br[167] wl[25] vdd gnd cell_6t
Xbit_r26_c167 bl[167] br[167] wl[26] vdd gnd cell_6t
Xbit_r27_c167 bl[167] br[167] wl[27] vdd gnd cell_6t
Xbit_r28_c167 bl[167] br[167] wl[28] vdd gnd cell_6t
Xbit_r29_c167 bl[167] br[167] wl[29] vdd gnd cell_6t
Xbit_r30_c167 bl[167] br[167] wl[30] vdd gnd cell_6t
Xbit_r31_c167 bl[167] br[167] wl[31] vdd gnd cell_6t
Xbit_r32_c167 bl[167] br[167] wl[32] vdd gnd cell_6t
Xbit_r33_c167 bl[167] br[167] wl[33] vdd gnd cell_6t
Xbit_r34_c167 bl[167] br[167] wl[34] vdd gnd cell_6t
Xbit_r35_c167 bl[167] br[167] wl[35] vdd gnd cell_6t
Xbit_r36_c167 bl[167] br[167] wl[36] vdd gnd cell_6t
Xbit_r37_c167 bl[167] br[167] wl[37] vdd gnd cell_6t
Xbit_r38_c167 bl[167] br[167] wl[38] vdd gnd cell_6t
Xbit_r39_c167 bl[167] br[167] wl[39] vdd gnd cell_6t
Xbit_r40_c167 bl[167] br[167] wl[40] vdd gnd cell_6t
Xbit_r41_c167 bl[167] br[167] wl[41] vdd gnd cell_6t
Xbit_r42_c167 bl[167] br[167] wl[42] vdd gnd cell_6t
Xbit_r43_c167 bl[167] br[167] wl[43] vdd gnd cell_6t
Xbit_r44_c167 bl[167] br[167] wl[44] vdd gnd cell_6t
Xbit_r45_c167 bl[167] br[167] wl[45] vdd gnd cell_6t
Xbit_r46_c167 bl[167] br[167] wl[46] vdd gnd cell_6t
Xbit_r47_c167 bl[167] br[167] wl[47] vdd gnd cell_6t
Xbit_r48_c167 bl[167] br[167] wl[48] vdd gnd cell_6t
Xbit_r49_c167 bl[167] br[167] wl[49] vdd gnd cell_6t
Xbit_r50_c167 bl[167] br[167] wl[50] vdd gnd cell_6t
Xbit_r51_c167 bl[167] br[167] wl[51] vdd gnd cell_6t
Xbit_r52_c167 bl[167] br[167] wl[52] vdd gnd cell_6t
Xbit_r53_c167 bl[167] br[167] wl[53] vdd gnd cell_6t
Xbit_r54_c167 bl[167] br[167] wl[54] vdd gnd cell_6t
Xbit_r55_c167 bl[167] br[167] wl[55] vdd gnd cell_6t
Xbit_r56_c167 bl[167] br[167] wl[56] vdd gnd cell_6t
Xbit_r57_c167 bl[167] br[167] wl[57] vdd gnd cell_6t
Xbit_r58_c167 bl[167] br[167] wl[58] vdd gnd cell_6t
Xbit_r59_c167 bl[167] br[167] wl[59] vdd gnd cell_6t
Xbit_r60_c167 bl[167] br[167] wl[60] vdd gnd cell_6t
Xbit_r61_c167 bl[167] br[167] wl[61] vdd gnd cell_6t
Xbit_r62_c167 bl[167] br[167] wl[62] vdd gnd cell_6t
Xbit_r63_c167 bl[167] br[167] wl[63] vdd gnd cell_6t
Xbit_r64_c167 bl[167] br[167] wl[64] vdd gnd cell_6t
Xbit_r65_c167 bl[167] br[167] wl[65] vdd gnd cell_6t
Xbit_r66_c167 bl[167] br[167] wl[66] vdd gnd cell_6t
Xbit_r67_c167 bl[167] br[167] wl[67] vdd gnd cell_6t
Xbit_r68_c167 bl[167] br[167] wl[68] vdd gnd cell_6t
Xbit_r69_c167 bl[167] br[167] wl[69] vdd gnd cell_6t
Xbit_r70_c167 bl[167] br[167] wl[70] vdd gnd cell_6t
Xbit_r71_c167 bl[167] br[167] wl[71] vdd gnd cell_6t
Xbit_r72_c167 bl[167] br[167] wl[72] vdd gnd cell_6t
Xbit_r73_c167 bl[167] br[167] wl[73] vdd gnd cell_6t
Xbit_r74_c167 bl[167] br[167] wl[74] vdd gnd cell_6t
Xbit_r75_c167 bl[167] br[167] wl[75] vdd gnd cell_6t
Xbit_r76_c167 bl[167] br[167] wl[76] vdd gnd cell_6t
Xbit_r77_c167 bl[167] br[167] wl[77] vdd gnd cell_6t
Xbit_r78_c167 bl[167] br[167] wl[78] vdd gnd cell_6t
Xbit_r79_c167 bl[167] br[167] wl[79] vdd gnd cell_6t
Xbit_r80_c167 bl[167] br[167] wl[80] vdd gnd cell_6t
Xbit_r81_c167 bl[167] br[167] wl[81] vdd gnd cell_6t
Xbit_r82_c167 bl[167] br[167] wl[82] vdd gnd cell_6t
Xbit_r83_c167 bl[167] br[167] wl[83] vdd gnd cell_6t
Xbit_r84_c167 bl[167] br[167] wl[84] vdd gnd cell_6t
Xbit_r85_c167 bl[167] br[167] wl[85] vdd gnd cell_6t
Xbit_r86_c167 bl[167] br[167] wl[86] vdd gnd cell_6t
Xbit_r87_c167 bl[167] br[167] wl[87] vdd gnd cell_6t
Xbit_r88_c167 bl[167] br[167] wl[88] vdd gnd cell_6t
Xbit_r89_c167 bl[167] br[167] wl[89] vdd gnd cell_6t
Xbit_r90_c167 bl[167] br[167] wl[90] vdd gnd cell_6t
Xbit_r91_c167 bl[167] br[167] wl[91] vdd gnd cell_6t
Xbit_r92_c167 bl[167] br[167] wl[92] vdd gnd cell_6t
Xbit_r93_c167 bl[167] br[167] wl[93] vdd gnd cell_6t
Xbit_r94_c167 bl[167] br[167] wl[94] vdd gnd cell_6t
Xbit_r95_c167 bl[167] br[167] wl[95] vdd gnd cell_6t
Xbit_r96_c167 bl[167] br[167] wl[96] vdd gnd cell_6t
Xbit_r97_c167 bl[167] br[167] wl[97] vdd gnd cell_6t
Xbit_r98_c167 bl[167] br[167] wl[98] vdd gnd cell_6t
Xbit_r99_c167 bl[167] br[167] wl[99] vdd gnd cell_6t
Xbit_r100_c167 bl[167] br[167] wl[100] vdd gnd cell_6t
Xbit_r101_c167 bl[167] br[167] wl[101] vdd gnd cell_6t
Xbit_r102_c167 bl[167] br[167] wl[102] vdd gnd cell_6t
Xbit_r103_c167 bl[167] br[167] wl[103] vdd gnd cell_6t
Xbit_r104_c167 bl[167] br[167] wl[104] vdd gnd cell_6t
Xbit_r105_c167 bl[167] br[167] wl[105] vdd gnd cell_6t
Xbit_r106_c167 bl[167] br[167] wl[106] vdd gnd cell_6t
Xbit_r107_c167 bl[167] br[167] wl[107] vdd gnd cell_6t
Xbit_r108_c167 bl[167] br[167] wl[108] vdd gnd cell_6t
Xbit_r109_c167 bl[167] br[167] wl[109] vdd gnd cell_6t
Xbit_r110_c167 bl[167] br[167] wl[110] vdd gnd cell_6t
Xbit_r111_c167 bl[167] br[167] wl[111] vdd gnd cell_6t
Xbit_r112_c167 bl[167] br[167] wl[112] vdd gnd cell_6t
Xbit_r113_c167 bl[167] br[167] wl[113] vdd gnd cell_6t
Xbit_r114_c167 bl[167] br[167] wl[114] vdd gnd cell_6t
Xbit_r115_c167 bl[167] br[167] wl[115] vdd gnd cell_6t
Xbit_r116_c167 bl[167] br[167] wl[116] vdd gnd cell_6t
Xbit_r117_c167 bl[167] br[167] wl[117] vdd gnd cell_6t
Xbit_r118_c167 bl[167] br[167] wl[118] vdd gnd cell_6t
Xbit_r119_c167 bl[167] br[167] wl[119] vdd gnd cell_6t
Xbit_r120_c167 bl[167] br[167] wl[120] vdd gnd cell_6t
Xbit_r121_c167 bl[167] br[167] wl[121] vdd gnd cell_6t
Xbit_r122_c167 bl[167] br[167] wl[122] vdd gnd cell_6t
Xbit_r123_c167 bl[167] br[167] wl[123] vdd gnd cell_6t
Xbit_r124_c167 bl[167] br[167] wl[124] vdd gnd cell_6t
Xbit_r125_c167 bl[167] br[167] wl[125] vdd gnd cell_6t
Xbit_r126_c167 bl[167] br[167] wl[126] vdd gnd cell_6t
Xbit_r127_c167 bl[167] br[167] wl[127] vdd gnd cell_6t
Xbit_r0_c168 bl[168] br[168] wl[0] vdd gnd cell_6t
Xbit_r1_c168 bl[168] br[168] wl[1] vdd gnd cell_6t
Xbit_r2_c168 bl[168] br[168] wl[2] vdd gnd cell_6t
Xbit_r3_c168 bl[168] br[168] wl[3] vdd gnd cell_6t
Xbit_r4_c168 bl[168] br[168] wl[4] vdd gnd cell_6t
Xbit_r5_c168 bl[168] br[168] wl[5] vdd gnd cell_6t
Xbit_r6_c168 bl[168] br[168] wl[6] vdd gnd cell_6t
Xbit_r7_c168 bl[168] br[168] wl[7] vdd gnd cell_6t
Xbit_r8_c168 bl[168] br[168] wl[8] vdd gnd cell_6t
Xbit_r9_c168 bl[168] br[168] wl[9] vdd gnd cell_6t
Xbit_r10_c168 bl[168] br[168] wl[10] vdd gnd cell_6t
Xbit_r11_c168 bl[168] br[168] wl[11] vdd gnd cell_6t
Xbit_r12_c168 bl[168] br[168] wl[12] vdd gnd cell_6t
Xbit_r13_c168 bl[168] br[168] wl[13] vdd gnd cell_6t
Xbit_r14_c168 bl[168] br[168] wl[14] vdd gnd cell_6t
Xbit_r15_c168 bl[168] br[168] wl[15] vdd gnd cell_6t
Xbit_r16_c168 bl[168] br[168] wl[16] vdd gnd cell_6t
Xbit_r17_c168 bl[168] br[168] wl[17] vdd gnd cell_6t
Xbit_r18_c168 bl[168] br[168] wl[18] vdd gnd cell_6t
Xbit_r19_c168 bl[168] br[168] wl[19] vdd gnd cell_6t
Xbit_r20_c168 bl[168] br[168] wl[20] vdd gnd cell_6t
Xbit_r21_c168 bl[168] br[168] wl[21] vdd gnd cell_6t
Xbit_r22_c168 bl[168] br[168] wl[22] vdd gnd cell_6t
Xbit_r23_c168 bl[168] br[168] wl[23] vdd gnd cell_6t
Xbit_r24_c168 bl[168] br[168] wl[24] vdd gnd cell_6t
Xbit_r25_c168 bl[168] br[168] wl[25] vdd gnd cell_6t
Xbit_r26_c168 bl[168] br[168] wl[26] vdd gnd cell_6t
Xbit_r27_c168 bl[168] br[168] wl[27] vdd gnd cell_6t
Xbit_r28_c168 bl[168] br[168] wl[28] vdd gnd cell_6t
Xbit_r29_c168 bl[168] br[168] wl[29] vdd gnd cell_6t
Xbit_r30_c168 bl[168] br[168] wl[30] vdd gnd cell_6t
Xbit_r31_c168 bl[168] br[168] wl[31] vdd gnd cell_6t
Xbit_r32_c168 bl[168] br[168] wl[32] vdd gnd cell_6t
Xbit_r33_c168 bl[168] br[168] wl[33] vdd gnd cell_6t
Xbit_r34_c168 bl[168] br[168] wl[34] vdd gnd cell_6t
Xbit_r35_c168 bl[168] br[168] wl[35] vdd gnd cell_6t
Xbit_r36_c168 bl[168] br[168] wl[36] vdd gnd cell_6t
Xbit_r37_c168 bl[168] br[168] wl[37] vdd gnd cell_6t
Xbit_r38_c168 bl[168] br[168] wl[38] vdd gnd cell_6t
Xbit_r39_c168 bl[168] br[168] wl[39] vdd gnd cell_6t
Xbit_r40_c168 bl[168] br[168] wl[40] vdd gnd cell_6t
Xbit_r41_c168 bl[168] br[168] wl[41] vdd gnd cell_6t
Xbit_r42_c168 bl[168] br[168] wl[42] vdd gnd cell_6t
Xbit_r43_c168 bl[168] br[168] wl[43] vdd gnd cell_6t
Xbit_r44_c168 bl[168] br[168] wl[44] vdd gnd cell_6t
Xbit_r45_c168 bl[168] br[168] wl[45] vdd gnd cell_6t
Xbit_r46_c168 bl[168] br[168] wl[46] vdd gnd cell_6t
Xbit_r47_c168 bl[168] br[168] wl[47] vdd gnd cell_6t
Xbit_r48_c168 bl[168] br[168] wl[48] vdd gnd cell_6t
Xbit_r49_c168 bl[168] br[168] wl[49] vdd gnd cell_6t
Xbit_r50_c168 bl[168] br[168] wl[50] vdd gnd cell_6t
Xbit_r51_c168 bl[168] br[168] wl[51] vdd gnd cell_6t
Xbit_r52_c168 bl[168] br[168] wl[52] vdd gnd cell_6t
Xbit_r53_c168 bl[168] br[168] wl[53] vdd gnd cell_6t
Xbit_r54_c168 bl[168] br[168] wl[54] vdd gnd cell_6t
Xbit_r55_c168 bl[168] br[168] wl[55] vdd gnd cell_6t
Xbit_r56_c168 bl[168] br[168] wl[56] vdd gnd cell_6t
Xbit_r57_c168 bl[168] br[168] wl[57] vdd gnd cell_6t
Xbit_r58_c168 bl[168] br[168] wl[58] vdd gnd cell_6t
Xbit_r59_c168 bl[168] br[168] wl[59] vdd gnd cell_6t
Xbit_r60_c168 bl[168] br[168] wl[60] vdd gnd cell_6t
Xbit_r61_c168 bl[168] br[168] wl[61] vdd gnd cell_6t
Xbit_r62_c168 bl[168] br[168] wl[62] vdd gnd cell_6t
Xbit_r63_c168 bl[168] br[168] wl[63] vdd gnd cell_6t
Xbit_r64_c168 bl[168] br[168] wl[64] vdd gnd cell_6t
Xbit_r65_c168 bl[168] br[168] wl[65] vdd gnd cell_6t
Xbit_r66_c168 bl[168] br[168] wl[66] vdd gnd cell_6t
Xbit_r67_c168 bl[168] br[168] wl[67] vdd gnd cell_6t
Xbit_r68_c168 bl[168] br[168] wl[68] vdd gnd cell_6t
Xbit_r69_c168 bl[168] br[168] wl[69] vdd gnd cell_6t
Xbit_r70_c168 bl[168] br[168] wl[70] vdd gnd cell_6t
Xbit_r71_c168 bl[168] br[168] wl[71] vdd gnd cell_6t
Xbit_r72_c168 bl[168] br[168] wl[72] vdd gnd cell_6t
Xbit_r73_c168 bl[168] br[168] wl[73] vdd gnd cell_6t
Xbit_r74_c168 bl[168] br[168] wl[74] vdd gnd cell_6t
Xbit_r75_c168 bl[168] br[168] wl[75] vdd gnd cell_6t
Xbit_r76_c168 bl[168] br[168] wl[76] vdd gnd cell_6t
Xbit_r77_c168 bl[168] br[168] wl[77] vdd gnd cell_6t
Xbit_r78_c168 bl[168] br[168] wl[78] vdd gnd cell_6t
Xbit_r79_c168 bl[168] br[168] wl[79] vdd gnd cell_6t
Xbit_r80_c168 bl[168] br[168] wl[80] vdd gnd cell_6t
Xbit_r81_c168 bl[168] br[168] wl[81] vdd gnd cell_6t
Xbit_r82_c168 bl[168] br[168] wl[82] vdd gnd cell_6t
Xbit_r83_c168 bl[168] br[168] wl[83] vdd gnd cell_6t
Xbit_r84_c168 bl[168] br[168] wl[84] vdd gnd cell_6t
Xbit_r85_c168 bl[168] br[168] wl[85] vdd gnd cell_6t
Xbit_r86_c168 bl[168] br[168] wl[86] vdd gnd cell_6t
Xbit_r87_c168 bl[168] br[168] wl[87] vdd gnd cell_6t
Xbit_r88_c168 bl[168] br[168] wl[88] vdd gnd cell_6t
Xbit_r89_c168 bl[168] br[168] wl[89] vdd gnd cell_6t
Xbit_r90_c168 bl[168] br[168] wl[90] vdd gnd cell_6t
Xbit_r91_c168 bl[168] br[168] wl[91] vdd gnd cell_6t
Xbit_r92_c168 bl[168] br[168] wl[92] vdd gnd cell_6t
Xbit_r93_c168 bl[168] br[168] wl[93] vdd gnd cell_6t
Xbit_r94_c168 bl[168] br[168] wl[94] vdd gnd cell_6t
Xbit_r95_c168 bl[168] br[168] wl[95] vdd gnd cell_6t
Xbit_r96_c168 bl[168] br[168] wl[96] vdd gnd cell_6t
Xbit_r97_c168 bl[168] br[168] wl[97] vdd gnd cell_6t
Xbit_r98_c168 bl[168] br[168] wl[98] vdd gnd cell_6t
Xbit_r99_c168 bl[168] br[168] wl[99] vdd gnd cell_6t
Xbit_r100_c168 bl[168] br[168] wl[100] vdd gnd cell_6t
Xbit_r101_c168 bl[168] br[168] wl[101] vdd gnd cell_6t
Xbit_r102_c168 bl[168] br[168] wl[102] vdd gnd cell_6t
Xbit_r103_c168 bl[168] br[168] wl[103] vdd gnd cell_6t
Xbit_r104_c168 bl[168] br[168] wl[104] vdd gnd cell_6t
Xbit_r105_c168 bl[168] br[168] wl[105] vdd gnd cell_6t
Xbit_r106_c168 bl[168] br[168] wl[106] vdd gnd cell_6t
Xbit_r107_c168 bl[168] br[168] wl[107] vdd gnd cell_6t
Xbit_r108_c168 bl[168] br[168] wl[108] vdd gnd cell_6t
Xbit_r109_c168 bl[168] br[168] wl[109] vdd gnd cell_6t
Xbit_r110_c168 bl[168] br[168] wl[110] vdd gnd cell_6t
Xbit_r111_c168 bl[168] br[168] wl[111] vdd gnd cell_6t
Xbit_r112_c168 bl[168] br[168] wl[112] vdd gnd cell_6t
Xbit_r113_c168 bl[168] br[168] wl[113] vdd gnd cell_6t
Xbit_r114_c168 bl[168] br[168] wl[114] vdd gnd cell_6t
Xbit_r115_c168 bl[168] br[168] wl[115] vdd gnd cell_6t
Xbit_r116_c168 bl[168] br[168] wl[116] vdd gnd cell_6t
Xbit_r117_c168 bl[168] br[168] wl[117] vdd gnd cell_6t
Xbit_r118_c168 bl[168] br[168] wl[118] vdd gnd cell_6t
Xbit_r119_c168 bl[168] br[168] wl[119] vdd gnd cell_6t
Xbit_r120_c168 bl[168] br[168] wl[120] vdd gnd cell_6t
Xbit_r121_c168 bl[168] br[168] wl[121] vdd gnd cell_6t
Xbit_r122_c168 bl[168] br[168] wl[122] vdd gnd cell_6t
Xbit_r123_c168 bl[168] br[168] wl[123] vdd gnd cell_6t
Xbit_r124_c168 bl[168] br[168] wl[124] vdd gnd cell_6t
Xbit_r125_c168 bl[168] br[168] wl[125] vdd gnd cell_6t
Xbit_r126_c168 bl[168] br[168] wl[126] vdd gnd cell_6t
Xbit_r127_c168 bl[168] br[168] wl[127] vdd gnd cell_6t
Xbit_r0_c169 bl[169] br[169] wl[0] vdd gnd cell_6t
Xbit_r1_c169 bl[169] br[169] wl[1] vdd gnd cell_6t
Xbit_r2_c169 bl[169] br[169] wl[2] vdd gnd cell_6t
Xbit_r3_c169 bl[169] br[169] wl[3] vdd gnd cell_6t
Xbit_r4_c169 bl[169] br[169] wl[4] vdd gnd cell_6t
Xbit_r5_c169 bl[169] br[169] wl[5] vdd gnd cell_6t
Xbit_r6_c169 bl[169] br[169] wl[6] vdd gnd cell_6t
Xbit_r7_c169 bl[169] br[169] wl[7] vdd gnd cell_6t
Xbit_r8_c169 bl[169] br[169] wl[8] vdd gnd cell_6t
Xbit_r9_c169 bl[169] br[169] wl[9] vdd gnd cell_6t
Xbit_r10_c169 bl[169] br[169] wl[10] vdd gnd cell_6t
Xbit_r11_c169 bl[169] br[169] wl[11] vdd gnd cell_6t
Xbit_r12_c169 bl[169] br[169] wl[12] vdd gnd cell_6t
Xbit_r13_c169 bl[169] br[169] wl[13] vdd gnd cell_6t
Xbit_r14_c169 bl[169] br[169] wl[14] vdd gnd cell_6t
Xbit_r15_c169 bl[169] br[169] wl[15] vdd gnd cell_6t
Xbit_r16_c169 bl[169] br[169] wl[16] vdd gnd cell_6t
Xbit_r17_c169 bl[169] br[169] wl[17] vdd gnd cell_6t
Xbit_r18_c169 bl[169] br[169] wl[18] vdd gnd cell_6t
Xbit_r19_c169 bl[169] br[169] wl[19] vdd gnd cell_6t
Xbit_r20_c169 bl[169] br[169] wl[20] vdd gnd cell_6t
Xbit_r21_c169 bl[169] br[169] wl[21] vdd gnd cell_6t
Xbit_r22_c169 bl[169] br[169] wl[22] vdd gnd cell_6t
Xbit_r23_c169 bl[169] br[169] wl[23] vdd gnd cell_6t
Xbit_r24_c169 bl[169] br[169] wl[24] vdd gnd cell_6t
Xbit_r25_c169 bl[169] br[169] wl[25] vdd gnd cell_6t
Xbit_r26_c169 bl[169] br[169] wl[26] vdd gnd cell_6t
Xbit_r27_c169 bl[169] br[169] wl[27] vdd gnd cell_6t
Xbit_r28_c169 bl[169] br[169] wl[28] vdd gnd cell_6t
Xbit_r29_c169 bl[169] br[169] wl[29] vdd gnd cell_6t
Xbit_r30_c169 bl[169] br[169] wl[30] vdd gnd cell_6t
Xbit_r31_c169 bl[169] br[169] wl[31] vdd gnd cell_6t
Xbit_r32_c169 bl[169] br[169] wl[32] vdd gnd cell_6t
Xbit_r33_c169 bl[169] br[169] wl[33] vdd gnd cell_6t
Xbit_r34_c169 bl[169] br[169] wl[34] vdd gnd cell_6t
Xbit_r35_c169 bl[169] br[169] wl[35] vdd gnd cell_6t
Xbit_r36_c169 bl[169] br[169] wl[36] vdd gnd cell_6t
Xbit_r37_c169 bl[169] br[169] wl[37] vdd gnd cell_6t
Xbit_r38_c169 bl[169] br[169] wl[38] vdd gnd cell_6t
Xbit_r39_c169 bl[169] br[169] wl[39] vdd gnd cell_6t
Xbit_r40_c169 bl[169] br[169] wl[40] vdd gnd cell_6t
Xbit_r41_c169 bl[169] br[169] wl[41] vdd gnd cell_6t
Xbit_r42_c169 bl[169] br[169] wl[42] vdd gnd cell_6t
Xbit_r43_c169 bl[169] br[169] wl[43] vdd gnd cell_6t
Xbit_r44_c169 bl[169] br[169] wl[44] vdd gnd cell_6t
Xbit_r45_c169 bl[169] br[169] wl[45] vdd gnd cell_6t
Xbit_r46_c169 bl[169] br[169] wl[46] vdd gnd cell_6t
Xbit_r47_c169 bl[169] br[169] wl[47] vdd gnd cell_6t
Xbit_r48_c169 bl[169] br[169] wl[48] vdd gnd cell_6t
Xbit_r49_c169 bl[169] br[169] wl[49] vdd gnd cell_6t
Xbit_r50_c169 bl[169] br[169] wl[50] vdd gnd cell_6t
Xbit_r51_c169 bl[169] br[169] wl[51] vdd gnd cell_6t
Xbit_r52_c169 bl[169] br[169] wl[52] vdd gnd cell_6t
Xbit_r53_c169 bl[169] br[169] wl[53] vdd gnd cell_6t
Xbit_r54_c169 bl[169] br[169] wl[54] vdd gnd cell_6t
Xbit_r55_c169 bl[169] br[169] wl[55] vdd gnd cell_6t
Xbit_r56_c169 bl[169] br[169] wl[56] vdd gnd cell_6t
Xbit_r57_c169 bl[169] br[169] wl[57] vdd gnd cell_6t
Xbit_r58_c169 bl[169] br[169] wl[58] vdd gnd cell_6t
Xbit_r59_c169 bl[169] br[169] wl[59] vdd gnd cell_6t
Xbit_r60_c169 bl[169] br[169] wl[60] vdd gnd cell_6t
Xbit_r61_c169 bl[169] br[169] wl[61] vdd gnd cell_6t
Xbit_r62_c169 bl[169] br[169] wl[62] vdd gnd cell_6t
Xbit_r63_c169 bl[169] br[169] wl[63] vdd gnd cell_6t
Xbit_r64_c169 bl[169] br[169] wl[64] vdd gnd cell_6t
Xbit_r65_c169 bl[169] br[169] wl[65] vdd gnd cell_6t
Xbit_r66_c169 bl[169] br[169] wl[66] vdd gnd cell_6t
Xbit_r67_c169 bl[169] br[169] wl[67] vdd gnd cell_6t
Xbit_r68_c169 bl[169] br[169] wl[68] vdd gnd cell_6t
Xbit_r69_c169 bl[169] br[169] wl[69] vdd gnd cell_6t
Xbit_r70_c169 bl[169] br[169] wl[70] vdd gnd cell_6t
Xbit_r71_c169 bl[169] br[169] wl[71] vdd gnd cell_6t
Xbit_r72_c169 bl[169] br[169] wl[72] vdd gnd cell_6t
Xbit_r73_c169 bl[169] br[169] wl[73] vdd gnd cell_6t
Xbit_r74_c169 bl[169] br[169] wl[74] vdd gnd cell_6t
Xbit_r75_c169 bl[169] br[169] wl[75] vdd gnd cell_6t
Xbit_r76_c169 bl[169] br[169] wl[76] vdd gnd cell_6t
Xbit_r77_c169 bl[169] br[169] wl[77] vdd gnd cell_6t
Xbit_r78_c169 bl[169] br[169] wl[78] vdd gnd cell_6t
Xbit_r79_c169 bl[169] br[169] wl[79] vdd gnd cell_6t
Xbit_r80_c169 bl[169] br[169] wl[80] vdd gnd cell_6t
Xbit_r81_c169 bl[169] br[169] wl[81] vdd gnd cell_6t
Xbit_r82_c169 bl[169] br[169] wl[82] vdd gnd cell_6t
Xbit_r83_c169 bl[169] br[169] wl[83] vdd gnd cell_6t
Xbit_r84_c169 bl[169] br[169] wl[84] vdd gnd cell_6t
Xbit_r85_c169 bl[169] br[169] wl[85] vdd gnd cell_6t
Xbit_r86_c169 bl[169] br[169] wl[86] vdd gnd cell_6t
Xbit_r87_c169 bl[169] br[169] wl[87] vdd gnd cell_6t
Xbit_r88_c169 bl[169] br[169] wl[88] vdd gnd cell_6t
Xbit_r89_c169 bl[169] br[169] wl[89] vdd gnd cell_6t
Xbit_r90_c169 bl[169] br[169] wl[90] vdd gnd cell_6t
Xbit_r91_c169 bl[169] br[169] wl[91] vdd gnd cell_6t
Xbit_r92_c169 bl[169] br[169] wl[92] vdd gnd cell_6t
Xbit_r93_c169 bl[169] br[169] wl[93] vdd gnd cell_6t
Xbit_r94_c169 bl[169] br[169] wl[94] vdd gnd cell_6t
Xbit_r95_c169 bl[169] br[169] wl[95] vdd gnd cell_6t
Xbit_r96_c169 bl[169] br[169] wl[96] vdd gnd cell_6t
Xbit_r97_c169 bl[169] br[169] wl[97] vdd gnd cell_6t
Xbit_r98_c169 bl[169] br[169] wl[98] vdd gnd cell_6t
Xbit_r99_c169 bl[169] br[169] wl[99] vdd gnd cell_6t
Xbit_r100_c169 bl[169] br[169] wl[100] vdd gnd cell_6t
Xbit_r101_c169 bl[169] br[169] wl[101] vdd gnd cell_6t
Xbit_r102_c169 bl[169] br[169] wl[102] vdd gnd cell_6t
Xbit_r103_c169 bl[169] br[169] wl[103] vdd gnd cell_6t
Xbit_r104_c169 bl[169] br[169] wl[104] vdd gnd cell_6t
Xbit_r105_c169 bl[169] br[169] wl[105] vdd gnd cell_6t
Xbit_r106_c169 bl[169] br[169] wl[106] vdd gnd cell_6t
Xbit_r107_c169 bl[169] br[169] wl[107] vdd gnd cell_6t
Xbit_r108_c169 bl[169] br[169] wl[108] vdd gnd cell_6t
Xbit_r109_c169 bl[169] br[169] wl[109] vdd gnd cell_6t
Xbit_r110_c169 bl[169] br[169] wl[110] vdd gnd cell_6t
Xbit_r111_c169 bl[169] br[169] wl[111] vdd gnd cell_6t
Xbit_r112_c169 bl[169] br[169] wl[112] vdd gnd cell_6t
Xbit_r113_c169 bl[169] br[169] wl[113] vdd gnd cell_6t
Xbit_r114_c169 bl[169] br[169] wl[114] vdd gnd cell_6t
Xbit_r115_c169 bl[169] br[169] wl[115] vdd gnd cell_6t
Xbit_r116_c169 bl[169] br[169] wl[116] vdd gnd cell_6t
Xbit_r117_c169 bl[169] br[169] wl[117] vdd gnd cell_6t
Xbit_r118_c169 bl[169] br[169] wl[118] vdd gnd cell_6t
Xbit_r119_c169 bl[169] br[169] wl[119] vdd gnd cell_6t
Xbit_r120_c169 bl[169] br[169] wl[120] vdd gnd cell_6t
Xbit_r121_c169 bl[169] br[169] wl[121] vdd gnd cell_6t
Xbit_r122_c169 bl[169] br[169] wl[122] vdd gnd cell_6t
Xbit_r123_c169 bl[169] br[169] wl[123] vdd gnd cell_6t
Xbit_r124_c169 bl[169] br[169] wl[124] vdd gnd cell_6t
Xbit_r125_c169 bl[169] br[169] wl[125] vdd gnd cell_6t
Xbit_r126_c169 bl[169] br[169] wl[126] vdd gnd cell_6t
Xbit_r127_c169 bl[169] br[169] wl[127] vdd gnd cell_6t
Xbit_r0_c170 bl[170] br[170] wl[0] vdd gnd cell_6t
Xbit_r1_c170 bl[170] br[170] wl[1] vdd gnd cell_6t
Xbit_r2_c170 bl[170] br[170] wl[2] vdd gnd cell_6t
Xbit_r3_c170 bl[170] br[170] wl[3] vdd gnd cell_6t
Xbit_r4_c170 bl[170] br[170] wl[4] vdd gnd cell_6t
Xbit_r5_c170 bl[170] br[170] wl[5] vdd gnd cell_6t
Xbit_r6_c170 bl[170] br[170] wl[6] vdd gnd cell_6t
Xbit_r7_c170 bl[170] br[170] wl[7] vdd gnd cell_6t
Xbit_r8_c170 bl[170] br[170] wl[8] vdd gnd cell_6t
Xbit_r9_c170 bl[170] br[170] wl[9] vdd gnd cell_6t
Xbit_r10_c170 bl[170] br[170] wl[10] vdd gnd cell_6t
Xbit_r11_c170 bl[170] br[170] wl[11] vdd gnd cell_6t
Xbit_r12_c170 bl[170] br[170] wl[12] vdd gnd cell_6t
Xbit_r13_c170 bl[170] br[170] wl[13] vdd gnd cell_6t
Xbit_r14_c170 bl[170] br[170] wl[14] vdd gnd cell_6t
Xbit_r15_c170 bl[170] br[170] wl[15] vdd gnd cell_6t
Xbit_r16_c170 bl[170] br[170] wl[16] vdd gnd cell_6t
Xbit_r17_c170 bl[170] br[170] wl[17] vdd gnd cell_6t
Xbit_r18_c170 bl[170] br[170] wl[18] vdd gnd cell_6t
Xbit_r19_c170 bl[170] br[170] wl[19] vdd gnd cell_6t
Xbit_r20_c170 bl[170] br[170] wl[20] vdd gnd cell_6t
Xbit_r21_c170 bl[170] br[170] wl[21] vdd gnd cell_6t
Xbit_r22_c170 bl[170] br[170] wl[22] vdd gnd cell_6t
Xbit_r23_c170 bl[170] br[170] wl[23] vdd gnd cell_6t
Xbit_r24_c170 bl[170] br[170] wl[24] vdd gnd cell_6t
Xbit_r25_c170 bl[170] br[170] wl[25] vdd gnd cell_6t
Xbit_r26_c170 bl[170] br[170] wl[26] vdd gnd cell_6t
Xbit_r27_c170 bl[170] br[170] wl[27] vdd gnd cell_6t
Xbit_r28_c170 bl[170] br[170] wl[28] vdd gnd cell_6t
Xbit_r29_c170 bl[170] br[170] wl[29] vdd gnd cell_6t
Xbit_r30_c170 bl[170] br[170] wl[30] vdd gnd cell_6t
Xbit_r31_c170 bl[170] br[170] wl[31] vdd gnd cell_6t
Xbit_r32_c170 bl[170] br[170] wl[32] vdd gnd cell_6t
Xbit_r33_c170 bl[170] br[170] wl[33] vdd gnd cell_6t
Xbit_r34_c170 bl[170] br[170] wl[34] vdd gnd cell_6t
Xbit_r35_c170 bl[170] br[170] wl[35] vdd gnd cell_6t
Xbit_r36_c170 bl[170] br[170] wl[36] vdd gnd cell_6t
Xbit_r37_c170 bl[170] br[170] wl[37] vdd gnd cell_6t
Xbit_r38_c170 bl[170] br[170] wl[38] vdd gnd cell_6t
Xbit_r39_c170 bl[170] br[170] wl[39] vdd gnd cell_6t
Xbit_r40_c170 bl[170] br[170] wl[40] vdd gnd cell_6t
Xbit_r41_c170 bl[170] br[170] wl[41] vdd gnd cell_6t
Xbit_r42_c170 bl[170] br[170] wl[42] vdd gnd cell_6t
Xbit_r43_c170 bl[170] br[170] wl[43] vdd gnd cell_6t
Xbit_r44_c170 bl[170] br[170] wl[44] vdd gnd cell_6t
Xbit_r45_c170 bl[170] br[170] wl[45] vdd gnd cell_6t
Xbit_r46_c170 bl[170] br[170] wl[46] vdd gnd cell_6t
Xbit_r47_c170 bl[170] br[170] wl[47] vdd gnd cell_6t
Xbit_r48_c170 bl[170] br[170] wl[48] vdd gnd cell_6t
Xbit_r49_c170 bl[170] br[170] wl[49] vdd gnd cell_6t
Xbit_r50_c170 bl[170] br[170] wl[50] vdd gnd cell_6t
Xbit_r51_c170 bl[170] br[170] wl[51] vdd gnd cell_6t
Xbit_r52_c170 bl[170] br[170] wl[52] vdd gnd cell_6t
Xbit_r53_c170 bl[170] br[170] wl[53] vdd gnd cell_6t
Xbit_r54_c170 bl[170] br[170] wl[54] vdd gnd cell_6t
Xbit_r55_c170 bl[170] br[170] wl[55] vdd gnd cell_6t
Xbit_r56_c170 bl[170] br[170] wl[56] vdd gnd cell_6t
Xbit_r57_c170 bl[170] br[170] wl[57] vdd gnd cell_6t
Xbit_r58_c170 bl[170] br[170] wl[58] vdd gnd cell_6t
Xbit_r59_c170 bl[170] br[170] wl[59] vdd gnd cell_6t
Xbit_r60_c170 bl[170] br[170] wl[60] vdd gnd cell_6t
Xbit_r61_c170 bl[170] br[170] wl[61] vdd gnd cell_6t
Xbit_r62_c170 bl[170] br[170] wl[62] vdd gnd cell_6t
Xbit_r63_c170 bl[170] br[170] wl[63] vdd gnd cell_6t
Xbit_r64_c170 bl[170] br[170] wl[64] vdd gnd cell_6t
Xbit_r65_c170 bl[170] br[170] wl[65] vdd gnd cell_6t
Xbit_r66_c170 bl[170] br[170] wl[66] vdd gnd cell_6t
Xbit_r67_c170 bl[170] br[170] wl[67] vdd gnd cell_6t
Xbit_r68_c170 bl[170] br[170] wl[68] vdd gnd cell_6t
Xbit_r69_c170 bl[170] br[170] wl[69] vdd gnd cell_6t
Xbit_r70_c170 bl[170] br[170] wl[70] vdd gnd cell_6t
Xbit_r71_c170 bl[170] br[170] wl[71] vdd gnd cell_6t
Xbit_r72_c170 bl[170] br[170] wl[72] vdd gnd cell_6t
Xbit_r73_c170 bl[170] br[170] wl[73] vdd gnd cell_6t
Xbit_r74_c170 bl[170] br[170] wl[74] vdd gnd cell_6t
Xbit_r75_c170 bl[170] br[170] wl[75] vdd gnd cell_6t
Xbit_r76_c170 bl[170] br[170] wl[76] vdd gnd cell_6t
Xbit_r77_c170 bl[170] br[170] wl[77] vdd gnd cell_6t
Xbit_r78_c170 bl[170] br[170] wl[78] vdd gnd cell_6t
Xbit_r79_c170 bl[170] br[170] wl[79] vdd gnd cell_6t
Xbit_r80_c170 bl[170] br[170] wl[80] vdd gnd cell_6t
Xbit_r81_c170 bl[170] br[170] wl[81] vdd gnd cell_6t
Xbit_r82_c170 bl[170] br[170] wl[82] vdd gnd cell_6t
Xbit_r83_c170 bl[170] br[170] wl[83] vdd gnd cell_6t
Xbit_r84_c170 bl[170] br[170] wl[84] vdd gnd cell_6t
Xbit_r85_c170 bl[170] br[170] wl[85] vdd gnd cell_6t
Xbit_r86_c170 bl[170] br[170] wl[86] vdd gnd cell_6t
Xbit_r87_c170 bl[170] br[170] wl[87] vdd gnd cell_6t
Xbit_r88_c170 bl[170] br[170] wl[88] vdd gnd cell_6t
Xbit_r89_c170 bl[170] br[170] wl[89] vdd gnd cell_6t
Xbit_r90_c170 bl[170] br[170] wl[90] vdd gnd cell_6t
Xbit_r91_c170 bl[170] br[170] wl[91] vdd gnd cell_6t
Xbit_r92_c170 bl[170] br[170] wl[92] vdd gnd cell_6t
Xbit_r93_c170 bl[170] br[170] wl[93] vdd gnd cell_6t
Xbit_r94_c170 bl[170] br[170] wl[94] vdd gnd cell_6t
Xbit_r95_c170 bl[170] br[170] wl[95] vdd gnd cell_6t
Xbit_r96_c170 bl[170] br[170] wl[96] vdd gnd cell_6t
Xbit_r97_c170 bl[170] br[170] wl[97] vdd gnd cell_6t
Xbit_r98_c170 bl[170] br[170] wl[98] vdd gnd cell_6t
Xbit_r99_c170 bl[170] br[170] wl[99] vdd gnd cell_6t
Xbit_r100_c170 bl[170] br[170] wl[100] vdd gnd cell_6t
Xbit_r101_c170 bl[170] br[170] wl[101] vdd gnd cell_6t
Xbit_r102_c170 bl[170] br[170] wl[102] vdd gnd cell_6t
Xbit_r103_c170 bl[170] br[170] wl[103] vdd gnd cell_6t
Xbit_r104_c170 bl[170] br[170] wl[104] vdd gnd cell_6t
Xbit_r105_c170 bl[170] br[170] wl[105] vdd gnd cell_6t
Xbit_r106_c170 bl[170] br[170] wl[106] vdd gnd cell_6t
Xbit_r107_c170 bl[170] br[170] wl[107] vdd gnd cell_6t
Xbit_r108_c170 bl[170] br[170] wl[108] vdd gnd cell_6t
Xbit_r109_c170 bl[170] br[170] wl[109] vdd gnd cell_6t
Xbit_r110_c170 bl[170] br[170] wl[110] vdd gnd cell_6t
Xbit_r111_c170 bl[170] br[170] wl[111] vdd gnd cell_6t
Xbit_r112_c170 bl[170] br[170] wl[112] vdd gnd cell_6t
Xbit_r113_c170 bl[170] br[170] wl[113] vdd gnd cell_6t
Xbit_r114_c170 bl[170] br[170] wl[114] vdd gnd cell_6t
Xbit_r115_c170 bl[170] br[170] wl[115] vdd gnd cell_6t
Xbit_r116_c170 bl[170] br[170] wl[116] vdd gnd cell_6t
Xbit_r117_c170 bl[170] br[170] wl[117] vdd gnd cell_6t
Xbit_r118_c170 bl[170] br[170] wl[118] vdd gnd cell_6t
Xbit_r119_c170 bl[170] br[170] wl[119] vdd gnd cell_6t
Xbit_r120_c170 bl[170] br[170] wl[120] vdd gnd cell_6t
Xbit_r121_c170 bl[170] br[170] wl[121] vdd gnd cell_6t
Xbit_r122_c170 bl[170] br[170] wl[122] vdd gnd cell_6t
Xbit_r123_c170 bl[170] br[170] wl[123] vdd gnd cell_6t
Xbit_r124_c170 bl[170] br[170] wl[124] vdd gnd cell_6t
Xbit_r125_c170 bl[170] br[170] wl[125] vdd gnd cell_6t
Xbit_r126_c170 bl[170] br[170] wl[126] vdd gnd cell_6t
Xbit_r127_c170 bl[170] br[170] wl[127] vdd gnd cell_6t
Xbit_r0_c171 bl[171] br[171] wl[0] vdd gnd cell_6t
Xbit_r1_c171 bl[171] br[171] wl[1] vdd gnd cell_6t
Xbit_r2_c171 bl[171] br[171] wl[2] vdd gnd cell_6t
Xbit_r3_c171 bl[171] br[171] wl[3] vdd gnd cell_6t
Xbit_r4_c171 bl[171] br[171] wl[4] vdd gnd cell_6t
Xbit_r5_c171 bl[171] br[171] wl[5] vdd gnd cell_6t
Xbit_r6_c171 bl[171] br[171] wl[6] vdd gnd cell_6t
Xbit_r7_c171 bl[171] br[171] wl[7] vdd gnd cell_6t
Xbit_r8_c171 bl[171] br[171] wl[8] vdd gnd cell_6t
Xbit_r9_c171 bl[171] br[171] wl[9] vdd gnd cell_6t
Xbit_r10_c171 bl[171] br[171] wl[10] vdd gnd cell_6t
Xbit_r11_c171 bl[171] br[171] wl[11] vdd gnd cell_6t
Xbit_r12_c171 bl[171] br[171] wl[12] vdd gnd cell_6t
Xbit_r13_c171 bl[171] br[171] wl[13] vdd gnd cell_6t
Xbit_r14_c171 bl[171] br[171] wl[14] vdd gnd cell_6t
Xbit_r15_c171 bl[171] br[171] wl[15] vdd gnd cell_6t
Xbit_r16_c171 bl[171] br[171] wl[16] vdd gnd cell_6t
Xbit_r17_c171 bl[171] br[171] wl[17] vdd gnd cell_6t
Xbit_r18_c171 bl[171] br[171] wl[18] vdd gnd cell_6t
Xbit_r19_c171 bl[171] br[171] wl[19] vdd gnd cell_6t
Xbit_r20_c171 bl[171] br[171] wl[20] vdd gnd cell_6t
Xbit_r21_c171 bl[171] br[171] wl[21] vdd gnd cell_6t
Xbit_r22_c171 bl[171] br[171] wl[22] vdd gnd cell_6t
Xbit_r23_c171 bl[171] br[171] wl[23] vdd gnd cell_6t
Xbit_r24_c171 bl[171] br[171] wl[24] vdd gnd cell_6t
Xbit_r25_c171 bl[171] br[171] wl[25] vdd gnd cell_6t
Xbit_r26_c171 bl[171] br[171] wl[26] vdd gnd cell_6t
Xbit_r27_c171 bl[171] br[171] wl[27] vdd gnd cell_6t
Xbit_r28_c171 bl[171] br[171] wl[28] vdd gnd cell_6t
Xbit_r29_c171 bl[171] br[171] wl[29] vdd gnd cell_6t
Xbit_r30_c171 bl[171] br[171] wl[30] vdd gnd cell_6t
Xbit_r31_c171 bl[171] br[171] wl[31] vdd gnd cell_6t
Xbit_r32_c171 bl[171] br[171] wl[32] vdd gnd cell_6t
Xbit_r33_c171 bl[171] br[171] wl[33] vdd gnd cell_6t
Xbit_r34_c171 bl[171] br[171] wl[34] vdd gnd cell_6t
Xbit_r35_c171 bl[171] br[171] wl[35] vdd gnd cell_6t
Xbit_r36_c171 bl[171] br[171] wl[36] vdd gnd cell_6t
Xbit_r37_c171 bl[171] br[171] wl[37] vdd gnd cell_6t
Xbit_r38_c171 bl[171] br[171] wl[38] vdd gnd cell_6t
Xbit_r39_c171 bl[171] br[171] wl[39] vdd gnd cell_6t
Xbit_r40_c171 bl[171] br[171] wl[40] vdd gnd cell_6t
Xbit_r41_c171 bl[171] br[171] wl[41] vdd gnd cell_6t
Xbit_r42_c171 bl[171] br[171] wl[42] vdd gnd cell_6t
Xbit_r43_c171 bl[171] br[171] wl[43] vdd gnd cell_6t
Xbit_r44_c171 bl[171] br[171] wl[44] vdd gnd cell_6t
Xbit_r45_c171 bl[171] br[171] wl[45] vdd gnd cell_6t
Xbit_r46_c171 bl[171] br[171] wl[46] vdd gnd cell_6t
Xbit_r47_c171 bl[171] br[171] wl[47] vdd gnd cell_6t
Xbit_r48_c171 bl[171] br[171] wl[48] vdd gnd cell_6t
Xbit_r49_c171 bl[171] br[171] wl[49] vdd gnd cell_6t
Xbit_r50_c171 bl[171] br[171] wl[50] vdd gnd cell_6t
Xbit_r51_c171 bl[171] br[171] wl[51] vdd gnd cell_6t
Xbit_r52_c171 bl[171] br[171] wl[52] vdd gnd cell_6t
Xbit_r53_c171 bl[171] br[171] wl[53] vdd gnd cell_6t
Xbit_r54_c171 bl[171] br[171] wl[54] vdd gnd cell_6t
Xbit_r55_c171 bl[171] br[171] wl[55] vdd gnd cell_6t
Xbit_r56_c171 bl[171] br[171] wl[56] vdd gnd cell_6t
Xbit_r57_c171 bl[171] br[171] wl[57] vdd gnd cell_6t
Xbit_r58_c171 bl[171] br[171] wl[58] vdd gnd cell_6t
Xbit_r59_c171 bl[171] br[171] wl[59] vdd gnd cell_6t
Xbit_r60_c171 bl[171] br[171] wl[60] vdd gnd cell_6t
Xbit_r61_c171 bl[171] br[171] wl[61] vdd gnd cell_6t
Xbit_r62_c171 bl[171] br[171] wl[62] vdd gnd cell_6t
Xbit_r63_c171 bl[171] br[171] wl[63] vdd gnd cell_6t
Xbit_r64_c171 bl[171] br[171] wl[64] vdd gnd cell_6t
Xbit_r65_c171 bl[171] br[171] wl[65] vdd gnd cell_6t
Xbit_r66_c171 bl[171] br[171] wl[66] vdd gnd cell_6t
Xbit_r67_c171 bl[171] br[171] wl[67] vdd gnd cell_6t
Xbit_r68_c171 bl[171] br[171] wl[68] vdd gnd cell_6t
Xbit_r69_c171 bl[171] br[171] wl[69] vdd gnd cell_6t
Xbit_r70_c171 bl[171] br[171] wl[70] vdd gnd cell_6t
Xbit_r71_c171 bl[171] br[171] wl[71] vdd gnd cell_6t
Xbit_r72_c171 bl[171] br[171] wl[72] vdd gnd cell_6t
Xbit_r73_c171 bl[171] br[171] wl[73] vdd gnd cell_6t
Xbit_r74_c171 bl[171] br[171] wl[74] vdd gnd cell_6t
Xbit_r75_c171 bl[171] br[171] wl[75] vdd gnd cell_6t
Xbit_r76_c171 bl[171] br[171] wl[76] vdd gnd cell_6t
Xbit_r77_c171 bl[171] br[171] wl[77] vdd gnd cell_6t
Xbit_r78_c171 bl[171] br[171] wl[78] vdd gnd cell_6t
Xbit_r79_c171 bl[171] br[171] wl[79] vdd gnd cell_6t
Xbit_r80_c171 bl[171] br[171] wl[80] vdd gnd cell_6t
Xbit_r81_c171 bl[171] br[171] wl[81] vdd gnd cell_6t
Xbit_r82_c171 bl[171] br[171] wl[82] vdd gnd cell_6t
Xbit_r83_c171 bl[171] br[171] wl[83] vdd gnd cell_6t
Xbit_r84_c171 bl[171] br[171] wl[84] vdd gnd cell_6t
Xbit_r85_c171 bl[171] br[171] wl[85] vdd gnd cell_6t
Xbit_r86_c171 bl[171] br[171] wl[86] vdd gnd cell_6t
Xbit_r87_c171 bl[171] br[171] wl[87] vdd gnd cell_6t
Xbit_r88_c171 bl[171] br[171] wl[88] vdd gnd cell_6t
Xbit_r89_c171 bl[171] br[171] wl[89] vdd gnd cell_6t
Xbit_r90_c171 bl[171] br[171] wl[90] vdd gnd cell_6t
Xbit_r91_c171 bl[171] br[171] wl[91] vdd gnd cell_6t
Xbit_r92_c171 bl[171] br[171] wl[92] vdd gnd cell_6t
Xbit_r93_c171 bl[171] br[171] wl[93] vdd gnd cell_6t
Xbit_r94_c171 bl[171] br[171] wl[94] vdd gnd cell_6t
Xbit_r95_c171 bl[171] br[171] wl[95] vdd gnd cell_6t
Xbit_r96_c171 bl[171] br[171] wl[96] vdd gnd cell_6t
Xbit_r97_c171 bl[171] br[171] wl[97] vdd gnd cell_6t
Xbit_r98_c171 bl[171] br[171] wl[98] vdd gnd cell_6t
Xbit_r99_c171 bl[171] br[171] wl[99] vdd gnd cell_6t
Xbit_r100_c171 bl[171] br[171] wl[100] vdd gnd cell_6t
Xbit_r101_c171 bl[171] br[171] wl[101] vdd gnd cell_6t
Xbit_r102_c171 bl[171] br[171] wl[102] vdd gnd cell_6t
Xbit_r103_c171 bl[171] br[171] wl[103] vdd gnd cell_6t
Xbit_r104_c171 bl[171] br[171] wl[104] vdd gnd cell_6t
Xbit_r105_c171 bl[171] br[171] wl[105] vdd gnd cell_6t
Xbit_r106_c171 bl[171] br[171] wl[106] vdd gnd cell_6t
Xbit_r107_c171 bl[171] br[171] wl[107] vdd gnd cell_6t
Xbit_r108_c171 bl[171] br[171] wl[108] vdd gnd cell_6t
Xbit_r109_c171 bl[171] br[171] wl[109] vdd gnd cell_6t
Xbit_r110_c171 bl[171] br[171] wl[110] vdd gnd cell_6t
Xbit_r111_c171 bl[171] br[171] wl[111] vdd gnd cell_6t
Xbit_r112_c171 bl[171] br[171] wl[112] vdd gnd cell_6t
Xbit_r113_c171 bl[171] br[171] wl[113] vdd gnd cell_6t
Xbit_r114_c171 bl[171] br[171] wl[114] vdd gnd cell_6t
Xbit_r115_c171 bl[171] br[171] wl[115] vdd gnd cell_6t
Xbit_r116_c171 bl[171] br[171] wl[116] vdd gnd cell_6t
Xbit_r117_c171 bl[171] br[171] wl[117] vdd gnd cell_6t
Xbit_r118_c171 bl[171] br[171] wl[118] vdd gnd cell_6t
Xbit_r119_c171 bl[171] br[171] wl[119] vdd gnd cell_6t
Xbit_r120_c171 bl[171] br[171] wl[120] vdd gnd cell_6t
Xbit_r121_c171 bl[171] br[171] wl[121] vdd gnd cell_6t
Xbit_r122_c171 bl[171] br[171] wl[122] vdd gnd cell_6t
Xbit_r123_c171 bl[171] br[171] wl[123] vdd gnd cell_6t
Xbit_r124_c171 bl[171] br[171] wl[124] vdd gnd cell_6t
Xbit_r125_c171 bl[171] br[171] wl[125] vdd gnd cell_6t
Xbit_r126_c171 bl[171] br[171] wl[126] vdd gnd cell_6t
Xbit_r127_c171 bl[171] br[171] wl[127] vdd gnd cell_6t
Xbit_r0_c172 bl[172] br[172] wl[0] vdd gnd cell_6t
Xbit_r1_c172 bl[172] br[172] wl[1] vdd gnd cell_6t
Xbit_r2_c172 bl[172] br[172] wl[2] vdd gnd cell_6t
Xbit_r3_c172 bl[172] br[172] wl[3] vdd gnd cell_6t
Xbit_r4_c172 bl[172] br[172] wl[4] vdd gnd cell_6t
Xbit_r5_c172 bl[172] br[172] wl[5] vdd gnd cell_6t
Xbit_r6_c172 bl[172] br[172] wl[6] vdd gnd cell_6t
Xbit_r7_c172 bl[172] br[172] wl[7] vdd gnd cell_6t
Xbit_r8_c172 bl[172] br[172] wl[8] vdd gnd cell_6t
Xbit_r9_c172 bl[172] br[172] wl[9] vdd gnd cell_6t
Xbit_r10_c172 bl[172] br[172] wl[10] vdd gnd cell_6t
Xbit_r11_c172 bl[172] br[172] wl[11] vdd gnd cell_6t
Xbit_r12_c172 bl[172] br[172] wl[12] vdd gnd cell_6t
Xbit_r13_c172 bl[172] br[172] wl[13] vdd gnd cell_6t
Xbit_r14_c172 bl[172] br[172] wl[14] vdd gnd cell_6t
Xbit_r15_c172 bl[172] br[172] wl[15] vdd gnd cell_6t
Xbit_r16_c172 bl[172] br[172] wl[16] vdd gnd cell_6t
Xbit_r17_c172 bl[172] br[172] wl[17] vdd gnd cell_6t
Xbit_r18_c172 bl[172] br[172] wl[18] vdd gnd cell_6t
Xbit_r19_c172 bl[172] br[172] wl[19] vdd gnd cell_6t
Xbit_r20_c172 bl[172] br[172] wl[20] vdd gnd cell_6t
Xbit_r21_c172 bl[172] br[172] wl[21] vdd gnd cell_6t
Xbit_r22_c172 bl[172] br[172] wl[22] vdd gnd cell_6t
Xbit_r23_c172 bl[172] br[172] wl[23] vdd gnd cell_6t
Xbit_r24_c172 bl[172] br[172] wl[24] vdd gnd cell_6t
Xbit_r25_c172 bl[172] br[172] wl[25] vdd gnd cell_6t
Xbit_r26_c172 bl[172] br[172] wl[26] vdd gnd cell_6t
Xbit_r27_c172 bl[172] br[172] wl[27] vdd gnd cell_6t
Xbit_r28_c172 bl[172] br[172] wl[28] vdd gnd cell_6t
Xbit_r29_c172 bl[172] br[172] wl[29] vdd gnd cell_6t
Xbit_r30_c172 bl[172] br[172] wl[30] vdd gnd cell_6t
Xbit_r31_c172 bl[172] br[172] wl[31] vdd gnd cell_6t
Xbit_r32_c172 bl[172] br[172] wl[32] vdd gnd cell_6t
Xbit_r33_c172 bl[172] br[172] wl[33] vdd gnd cell_6t
Xbit_r34_c172 bl[172] br[172] wl[34] vdd gnd cell_6t
Xbit_r35_c172 bl[172] br[172] wl[35] vdd gnd cell_6t
Xbit_r36_c172 bl[172] br[172] wl[36] vdd gnd cell_6t
Xbit_r37_c172 bl[172] br[172] wl[37] vdd gnd cell_6t
Xbit_r38_c172 bl[172] br[172] wl[38] vdd gnd cell_6t
Xbit_r39_c172 bl[172] br[172] wl[39] vdd gnd cell_6t
Xbit_r40_c172 bl[172] br[172] wl[40] vdd gnd cell_6t
Xbit_r41_c172 bl[172] br[172] wl[41] vdd gnd cell_6t
Xbit_r42_c172 bl[172] br[172] wl[42] vdd gnd cell_6t
Xbit_r43_c172 bl[172] br[172] wl[43] vdd gnd cell_6t
Xbit_r44_c172 bl[172] br[172] wl[44] vdd gnd cell_6t
Xbit_r45_c172 bl[172] br[172] wl[45] vdd gnd cell_6t
Xbit_r46_c172 bl[172] br[172] wl[46] vdd gnd cell_6t
Xbit_r47_c172 bl[172] br[172] wl[47] vdd gnd cell_6t
Xbit_r48_c172 bl[172] br[172] wl[48] vdd gnd cell_6t
Xbit_r49_c172 bl[172] br[172] wl[49] vdd gnd cell_6t
Xbit_r50_c172 bl[172] br[172] wl[50] vdd gnd cell_6t
Xbit_r51_c172 bl[172] br[172] wl[51] vdd gnd cell_6t
Xbit_r52_c172 bl[172] br[172] wl[52] vdd gnd cell_6t
Xbit_r53_c172 bl[172] br[172] wl[53] vdd gnd cell_6t
Xbit_r54_c172 bl[172] br[172] wl[54] vdd gnd cell_6t
Xbit_r55_c172 bl[172] br[172] wl[55] vdd gnd cell_6t
Xbit_r56_c172 bl[172] br[172] wl[56] vdd gnd cell_6t
Xbit_r57_c172 bl[172] br[172] wl[57] vdd gnd cell_6t
Xbit_r58_c172 bl[172] br[172] wl[58] vdd gnd cell_6t
Xbit_r59_c172 bl[172] br[172] wl[59] vdd gnd cell_6t
Xbit_r60_c172 bl[172] br[172] wl[60] vdd gnd cell_6t
Xbit_r61_c172 bl[172] br[172] wl[61] vdd gnd cell_6t
Xbit_r62_c172 bl[172] br[172] wl[62] vdd gnd cell_6t
Xbit_r63_c172 bl[172] br[172] wl[63] vdd gnd cell_6t
Xbit_r64_c172 bl[172] br[172] wl[64] vdd gnd cell_6t
Xbit_r65_c172 bl[172] br[172] wl[65] vdd gnd cell_6t
Xbit_r66_c172 bl[172] br[172] wl[66] vdd gnd cell_6t
Xbit_r67_c172 bl[172] br[172] wl[67] vdd gnd cell_6t
Xbit_r68_c172 bl[172] br[172] wl[68] vdd gnd cell_6t
Xbit_r69_c172 bl[172] br[172] wl[69] vdd gnd cell_6t
Xbit_r70_c172 bl[172] br[172] wl[70] vdd gnd cell_6t
Xbit_r71_c172 bl[172] br[172] wl[71] vdd gnd cell_6t
Xbit_r72_c172 bl[172] br[172] wl[72] vdd gnd cell_6t
Xbit_r73_c172 bl[172] br[172] wl[73] vdd gnd cell_6t
Xbit_r74_c172 bl[172] br[172] wl[74] vdd gnd cell_6t
Xbit_r75_c172 bl[172] br[172] wl[75] vdd gnd cell_6t
Xbit_r76_c172 bl[172] br[172] wl[76] vdd gnd cell_6t
Xbit_r77_c172 bl[172] br[172] wl[77] vdd gnd cell_6t
Xbit_r78_c172 bl[172] br[172] wl[78] vdd gnd cell_6t
Xbit_r79_c172 bl[172] br[172] wl[79] vdd gnd cell_6t
Xbit_r80_c172 bl[172] br[172] wl[80] vdd gnd cell_6t
Xbit_r81_c172 bl[172] br[172] wl[81] vdd gnd cell_6t
Xbit_r82_c172 bl[172] br[172] wl[82] vdd gnd cell_6t
Xbit_r83_c172 bl[172] br[172] wl[83] vdd gnd cell_6t
Xbit_r84_c172 bl[172] br[172] wl[84] vdd gnd cell_6t
Xbit_r85_c172 bl[172] br[172] wl[85] vdd gnd cell_6t
Xbit_r86_c172 bl[172] br[172] wl[86] vdd gnd cell_6t
Xbit_r87_c172 bl[172] br[172] wl[87] vdd gnd cell_6t
Xbit_r88_c172 bl[172] br[172] wl[88] vdd gnd cell_6t
Xbit_r89_c172 bl[172] br[172] wl[89] vdd gnd cell_6t
Xbit_r90_c172 bl[172] br[172] wl[90] vdd gnd cell_6t
Xbit_r91_c172 bl[172] br[172] wl[91] vdd gnd cell_6t
Xbit_r92_c172 bl[172] br[172] wl[92] vdd gnd cell_6t
Xbit_r93_c172 bl[172] br[172] wl[93] vdd gnd cell_6t
Xbit_r94_c172 bl[172] br[172] wl[94] vdd gnd cell_6t
Xbit_r95_c172 bl[172] br[172] wl[95] vdd gnd cell_6t
Xbit_r96_c172 bl[172] br[172] wl[96] vdd gnd cell_6t
Xbit_r97_c172 bl[172] br[172] wl[97] vdd gnd cell_6t
Xbit_r98_c172 bl[172] br[172] wl[98] vdd gnd cell_6t
Xbit_r99_c172 bl[172] br[172] wl[99] vdd gnd cell_6t
Xbit_r100_c172 bl[172] br[172] wl[100] vdd gnd cell_6t
Xbit_r101_c172 bl[172] br[172] wl[101] vdd gnd cell_6t
Xbit_r102_c172 bl[172] br[172] wl[102] vdd gnd cell_6t
Xbit_r103_c172 bl[172] br[172] wl[103] vdd gnd cell_6t
Xbit_r104_c172 bl[172] br[172] wl[104] vdd gnd cell_6t
Xbit_r105_c172 bl[172] br[172] wl[105] vdd gnd cell_6t
Xbit_r106_c172 bl[172] br[172] wl[106] vdd gnd cell_6t
Xbit_r107_c172 bl[172] br[172] wl[107] vdd gnd cell_6t
Xbit_r108_c172 bl[172] br[172] wl[108] vdd gnd cell_6t
Xbit_r109_c172 bl[172] br[172] wl[109] vdd gnd cell_6t
Xbit_r110_c172 bl[172] br[172] wl[110] vdd gnd cell_6t
Xbit_r111_c172 bl[172] br[172] wl[111] vdd gnd cell_6t
Xbit_r112_c172 bl[172] br[172] wl[112] vdd gnd cell_6t
Xbit_r113_c172 bl[172] br[172] wl[113] vdd gnd cell_6t
Xbit_r114_c172 bl[172] br[172] wl[114] vdd gnd cell_6t
Xbit_r115_c172 bl[172] br[172] wl[115] vdd gnd cell_6t
Xbit_r116_c172 bl[172] br[172] wl[116] vdd gnd cell_6t
Xbit_r117_c172 bl[172] br[172] wl[117] vdd gnd cell_6t
Xbit_r118_c172 bl[172] br[172] wl[118] vdd gnd cell_6t
Xbit_r119_c172 bl[172] br[172] wl[119] vdd gnd cell_6t
Xbit_r120_c172 bl[172] br[172] wl[120] vdd gnd cell_6t
Xbit_r121_c172 bl[172] br[172] wl[121] vdd gnd cell_6t
Xbit_r122_c172 bl[172] br[172] wl[122] vdd gnd cell_6t
Xbit_r123_c172 bl[172] br[172] wl[123] vdd gnd cell_6t
Xbit_r124_c172 bl[172] br[172] wl[124] vdd gnd cell_6t
Xbit_r125_c172 bl[172] br[172] wl[125] vdd gnd cell_6t
Xbit_r126_c172 bl[172] br[172] wl[126] vdd gnd cell_6t
Xbit_r127_c172 bl[172] br[172] wl[127] vdd gnd cell_6t
Xbit_r0_c173 bl[173] br[173] wl[0] vdd gnd cell_6t
Xbit_r1_c173 bl[173] br[173] wl[1] vdd gnd cell_6t
Xbit_r2_c173 bl[173] br[173] wl[2] vdd gnd cell_6t
Xbit_r3_c173 bl[173] br[173] wl[3] vdd gnd cell_6t
Xbit_r4_c173 bl[173] br[173] wl[4] vdd gnd cell_6t
Xbit_r5_c173 bl[173] br[173] wl[5] vdd gnd cell_6t
Xbit_r6_c173 bl[173] br[173] wl[6] vdd gnd cell_6t
Xbit_r7_c173 bl[173] br[173] wl[7] vdd gnd cell_6t
Xbit_r8_c173 bl[173] br[173] wl[8] vdd gnd cell_6t
Xbit_r9_c173 bl[173] br[173] wl[9] vdd gnd cell_6t
Xbit_r10_c173 bl[173] br[173] wl[10] vdd gnd cell_6t
Xbit_r11_c173 bl[173] br[173] wl[11] vdd gnd cell_6t
Xbit_r12_c173 bl[173] br[173] wl[12] vdd gnd cell_6t
Xbit_r13_c173 bl[173] br[173] wl[13] vdd gnd cell_6t
Xbit_r14_c173 bl[173] br[173] wl[14] vdd gnd cell_6t
Xbit_r15_c173 bl[173] br[173] wl[15] vdd gnd cell_6t
Xbit_r16_c173 bl[173] br[173] wl[16] vdd gnd cell_6t
Xbit_r17_c173 bl[173] br[173] wl[17] vdd gnd cell_6t
Xbit_r18_c173 bl[173] br[173] wl[18] vdd gnd cell_6t
Xbit_r19_c173 bl[173] br[173] wl[19] vdd gnd cell_6t
Xbit_r20_c173 bl[173] br[173] wl[20] vdd gnd cell_6t
Xbit_r21_c173 bl[173] br[173] wl[21] vdd gnd cell_6t
Xbit_r22_c173 bl[173] br[173] wl[22] vdd gnd cell_6t
Xbit_r23_c173 bl[173] br[173] wl[23] vdd gnd cell_6t
Xbit_r24_c173 bl[173] br[173] wl[24] vdd gnd cell_6t
Xbit_r25_c173 bl[173] br[173] wl[25] vdd gnd cell_6t
Xbit_r26_c173 bl[173] br[173] wl[26] vdd gnd cell_6t
Xbit_r27_c173 bl[173] br[173] wl[27] vdd gnd cell_6t
Xbit_r28_c173 bl[173] br[173] wl[28] vdd gnd cell_6t
Xbit_r29_c173 bl[173] br[173] wl[29] vdd gnd cell_6t
Xbit_r30_c173 bl[173] br[173] wl[30] vdd gnd cell_6t
Xbit_r31_c173 bl[173] br[173] wl[31] vdd gnd cell_6t
Xbit_r32_c173 bl[173] br[173] wl[32] vdd gnd cell_6t
Xbit_r33_c173 bl[173] br[173] wl[33] vdd gnd cell_6t
Xbit_r34_c173 bl[173] br[173] wl[34] vdd gnd cell_6t
Xbit_r35_c173 bl[173] br[173] wl[35] vdd gnd cell_6t
Xbit_r36_c173 bl[173] br[173] wl[36] vdd gnd cell_6t
Xbit_r37_c173 bl[173] br[173] wl[37] vdd gnd cell_6t
Xbit_r38_c173 bl[173] br[173] wl[38] vdd gnd cell_6t
Xbit_r39_c173 bl[173] br[173] wl[39] vdd gnd cell_6t
Xbit_r40_c173 bl[173] br[173] wl[40] vdd gnd cell_6t
Xbit_r41_c173 bl[173] br[173] wl[41] vdd gnd cell_6t
Xbit_r42_c173 bl[173] br[173] wl[42] vdd gnd cell_6t
Xbit_r43_c173 bl[173] br[173] wl[43] vdd gnd cell_6t
Xbit_r44_c173 bl[173] br[173] wl[44] vdd gnd cell_6t
Xbit_r45_c173 bl[173] br[173] wl[45] vdd gnd cell_6t
Xbit_r46_c173 bl[173] br[173] wl[46] vdd gnd cell_6t
Xbit_r47_c173 bl[173] br[173] wl[47] vdd gnd cell_6t
Xbit_r48_c173 bl[173] br[173] wl[48] vdd gnd cell_6t
Xbit_r49_c173 bl[173] br[173] wl[49] vdd gnd cell_6t
Xbit_r50_c173 bl[173] br[173] wl[50] vdd gnd cell_6t
Xbit_r51_c173 bl[173] br[173] wl[51] vdd gnd cell_6t
Xbit_r52_c173 bl[173] br[173] wl[52] vdd gnd cell_6t
Xbit_r53_c173 bl[173] br[173] wl[53] vdd gnd cell_6t
Xbit_r54_c173 bl[173] br[173] wl[54] vdd gnd cell_6t
Xbit_r55_c173 bl[173] br[173] wl[55] vdd gnd cell_6t
Xbit_r56_c173 bl[173] br[173] wl[56] vdd gnd cell_6t
Xbit_r57_c173 bl[173] br[173] wl[57] vdd gnd cell_6t
Xbit_r58_c173 bl[173] br[173] wl[58] vdd gnd cell_6t
Xbit_r59_c173 bl[173] br[173] wl[59] vdd gnd cell_6t
Xbit_r60_c173 bl[173] br[173] wl[60] vdd gnd cell_6t
Xbit_r61_c173 bl[173] br[173] wl[61] vdd gnd cell_6t
Xbit_r62_c173 bl[173] br[173] wl[62] vdd gnd cell_6t
Xbit_r63_c173 bl[173] br[173] wl[63] vdd gnd cell_6t
Xbit_r64_c173 bl[173] br[173] wl[64] vdd gnd cell_6t
Xbit_r65_c173 bl[173] br[173] wl[65] vdd gnd cell_6t
Xbit_r66_c173 bl[173] br[173] wl[66] vdd gnd cell_6t
Xbit_r67_c173 bl[173] br[173] wl[67] vdd gnd cell_6t
Xbit_r68_c173 bl[173] br[173] wl[68] vdd gnd cell_6t
Xbit_r69_c173 bl[173] br[173] wl[69] vdd gnd cell_6t
Xbit_r70_c173 bl[173] br[173] wl[70] vdd gnd cell_6t
Xbit_r71_c173 bl[173] br[173] wl[71] vdd gnd cell_6t
Xbit_r72_c173 bl[173] br[173] wl[72] vdd gnd cell_6t
Xbit_r73_c173 bl[173] br[173] wl[73] vdd gnd cell_6t
Xbit_r74_c173 bl[173] br[173] wl[74] vdd gnd cell_6t
Xbit_r75_c173 bl[173] br[173] wl[75] vdd gnd cell_6t
Xbit_r76_c173 bl[173] br[173] wl[76] vdd gnd cell_6t
Xbit_r77_c173 bl[173] br[173] wl[77] vdd gnd cell_6t
Xbit_r78_c173 bl[173] br[173] wl[78] vdd gnd cell_6t
Xbit_r79_c173 bl[173] br[173] wl[79] vdd gnd cell_6t
Xbit_r80_c173 bl[173] br[173] wl[80] vdd gnd cell_6t
Xbit_r81_c173 bl[173] br[173] wl[81] vdd gnd cell_6t
Xbit_r82_c173 bl[173] br[173] wl[82] vdd gnd cell_6t
Xbit_r83_c173 bl[173] br[173] wl[83] vdd gnd cell_6t
Xbit_r84_c173 bl[173] br[173] wl[84] vdd gnd cell_6t
Xbit_r85_c173 bl[173] br[173] wl[85] vdd gnd cell_6t
Xbit_r86_c173 bl[173] br[173] wl[86] vdd gnd cell_6t
Xbit_r87_c173 bl[173] br[173] wl[87] vdd gnd cell_6t
Xbit_r88_c173 bl[173] br[173] wl[88] vdd gnd cell_6t
Xbit_r89_c173 bl[173] br[173] wl[89] vdd gnd cell_6t
Xbit_r90_c173 bl[173] br[173] wl[90] vdd gnd cell_6t
Xbit_r91_c173 bl[173] br[173] wl[91] vdd gnd cell_6t
Xbit_r92_c173 bl[173] br[173] wl[92] vdd gnd cell_6t
Xbit_r93_c173 bl[173] br[173] wl[93] vdd gnd cell_6t
Xbit_r94_c173 bl[173] br[173] wl[94] vdd gnd cell_6t
Xbit_r95_c173 bl[173] br[173] wl[95] vdd gnd cell_6t
Xbit_r96_c173 bl[173] br[173] wl[96] vdd gnd cell_6t
Xbit_r97_c173 bl[173] br[173] wl[97] vdd gnd cell_6t
Xbit_r98_c173 bl[173] br[173] wl[98] vdd gnd cell_6t
Xbit_r99_c173 bl[173] br[173] wl[99] vdd gnd cell_6t
Xbit_r100_c173 bl[173] br[173] wl[100] vdd gnd cell_6t
Xbit_r101_c173 bl[173] br[173] wl[101] vdd gnd cell_6t
Xbit_r102_c173 bl[173] br[173] wl[102] vdd gnd cell_6t
Xbit_r103_c173 bl[173] br[173] wl[103] vdd gnd cell_6t
Xbit_r104_c173 bl[173] br[173] wl[104] vdd gnd cell_6t
Xbit_r105_c173 bl[173] br[173] wl[105] vdd gnd cell_6t
Xbit_r106_c173 bl[173] br[173] wl[106] vdd gnd cell_6t
Xbit_r107_c173 bl[173] br[173] wl[107] vdd gnd cell_6t
Xbit_r108_c173 bl[173] br[173] wl[108] vdd gnd cell_6t
Xbit_r109_c173 bl[173] br[173] wl[109] vdd gnd cell_6t
Xbit_r110_c173 bl[173] br[173] wl[110] vdd gnd cell_6t
Xbit_r111_c173 bl[173] br[173] wl[111] vdd gnd cell_6t
Xbit_r112_c173 bl[173] br[173] wl[112] vdd gnd cell_6t
Xbit_r113_c173 bl[173] br[173] wl[113] vdd gnd cell_6t
Xbit_r114_c173 bl[173] br[173] wl[114] vdd gnd cell_6t
Xbit_r115_c173 bl[173] br[173] wl[115] vdd gnd cell_6t
Xbit_r116_c173 bl[173] br[173] wl[116] vdd gnd cell_6t
Xbit_r117_c173 bl[173] br[173] wl[117] vdd gnd cell_6t
Xbit_r118_c173 bl[173] br[173] wl[118] vdd gnd cell_6t
Xbit_r119_c173 bl[173] br[173] wl[119] vdd gnd cell_6t
Xbit_r120_c173 bl[173] br[173] wl[120] vdd gnd cell_6t
Xbit_r121_c173 bl[173] br[173] wl[121] vdd gnd cell_6t
Xbit_r122_c173 bl[173] br[173] wl[122] vdd gnd cell_6t
Xbit_r123_c173 bl[173] br[173] wl[123] vdd gnd cell_6t
Xbit_r124_c173 bl[173] br[173] wl[124] vdd gnd cell_6t
Xbit_r125_c173 bl[173] br[173] wl[125] vdd gnd cell_6t
Xbit_r126_c173 bl[173] br[173] wl[126] vdd gnd cell_6t
Xbit_r127_c173 bl[173] br[173] wl[127] vdd gnd cell_6t
Xbit_r0_c174 bl[174] br[174] wl[0] vdd gnd cell_6t
Xbit_r1_c174 bl[174] br[174] wl[1] vdd gnd cell_6t
Xbit_r2_c174 bl[174] br[174] wl[2] vdd gnd cell_6t
Xbit_r3_c174 bl[174] br[174] wl[3] vdd gnd cell_6t
Xbit_r4_c174 bl[174] br[174] wl[4] vdd gnd cell_6t
Xbit_r5_c174 bl[174] br[174] wl[5] vdd gnd cell_6t
Xbit_r6_c174 bl[174] br[174] wl[6] vdd gnd cell_6t
Xbit_r7_c174 bl[174] br[174] wl[7] vdd gnd cell_6t
Xbit_r8_c174 bl[174] br[174] wl[8] vdd gnd cell_6t
Xbit_r9_c174 bl[174] br[174] wl[9] vdd gnd cell_6t
Xbit_r10_c174 bl[174] br[174] wl[10] vdd gnd cell_6t
Xbit_r11_c174 bl[174] br[174] wl[11] vdd gnd cell_6t
Xbit_r12_c174 bl[174] br[174] wl[12] vdd gnd cell_6t
Xbit_r13_c174 bl[174] br[174] wl[13] vdd gnd cell_6t
Xbit_r14_c174 bl[174] br[174] wl[14] vdd gnd cell_6t
Xbit_r15_c174 bl[174] br[174] wl[15] vdd gnd cell_6t
Xbit_r16_c174 bl[174] br[174] wl[16] vdd gnd cell_6t
Xbit_r17_c174 bl[174] br[174] wl[17] vdd gnd cell_6t
Xbit_r18_c174 bl[174] br[174] wl[18] vdd gnd cell_6t
Xbit_r19_c174 bl[174] br[174] wl[19] vdd gnd cell_6t
Xbit_r20_c174 bl[174] br[174] wl[20] vdd gnd cell_6t
Xbit_r21_c174 bl[174] br[174] wl[21] vdd gnd cell_6t
Xbit_r22_c174 bl[174] br[174] wl[22] vdd gnd cell_6t
Xbit_r23_c174 bl[174] br[174] wl[23] vdd gnd cell_6t
Xbit_r24_c174 bl[174] br[174] wl[24] vdd gnd cell_6t
Xbit_r25_c174 bl[174] br[174] wl[25] vdd gnd cell_6t
Xbit_r26_c174 bl[174] br[174] wl[26] vdd gnd cell_6t
Xbit_r27_c174 bl[174] br[174] wl[27] vdd gnd cell_6t
Xbit_r28_c174 bl[174] br[174] wl[28] vdd gnd cell_6t
Xbit_r29_c174 bl[174] br[174] wl[29] vdd gnd cell_6t
Xbit_r30_c174 bl[174] br[174] wl[30] vdd gnd cell_6t
Xbit_r31_c174 bl[174] br[174] wl[31] vdd gnd cell_6t
Xbit_r32_c174 bl[174] br[174] wl[32] vdd gnd cell_6t
Xbit_r33_c174 bl[174] br[174] wl[33] vdd gnd cell_6t
Xbit_r34_c174 bl[174] br[174] wl[34] vdd gnd cell_6t
Xbit_r35_c174 bl[174] br[174] wl[35] vdd gnd cell_6t
Xbit_r36_c174 bl[174] br[174] wl[36] vdd gnd cell_6t
Xbit_r37_c174 bl[174] br[174] wl[37] vdd gnd cell_6t
Xbit_r38_c174 bl[174] br[174] wl[38] vdd gnd cell_6t
Xbit_r39_c174 bl[174] br[174] wl[39] vdd gnd cell_6t
Xbit_r40_c174 bl[174] br[174] wl[40] vdd gnd cell_6t
Xbit_r41_c174 bl[174] br[174] wl[41] vdd gnd cell_6t
Xbit_r42_c174 bl[174] br[174] wl[42] vdd gnd cell_6t
Xbit_r43_c174 bl[174] br[174] wl[43] vdd gnd cell_6t
Xbit_r44_c174 bl[174] br[174] wl[44] vdd gnd cell_6t
Xbit_r45_c174 bl[174] br[174] wl[45] vdd gnd cell_6t
Xbit_r46_c174 bl[174] br[174] wl[46] vdd gnd cell_6t
Xbit_r47_c174 bl[174] br[174] wl[47] vdd gnd cell_6t
Xbit_r48_c174 bl[174] br[174] wl[48] vdd gnd cell_6t
Xbit_r49_c174 bl[174] br[174] wl[49] vdd gnd cell_6t
Xbit_r50_c174 bl[174] br[174] wl[50] vdd gnd cell_6t
Xbit_r51_c174 bl[174] br[174] wl[51] vdd gnd cell_6t
Xbit_r52_c174 bl[174] br[174] wl[52] vdd gnd cell_6t
Xbit_r53_c174 bl[174] br[174] wl[53] vdd gnd cell_6t
Xbit_r54_c174 bl[174] br[174] wl[54] vdd gnd cell_6t
Xbit_r55_c174 bl[174] br[174] wl[55] vdd gnd cell_6t
Xbit_r56_c174 bl[174] br[174] wl[56] vdd gnd cell_6t
Xbit_r57_c174 bl[174] br[174] wl[57] vdd gnd cell_6t
Xbit_r58_c174 bl[174] br[174] wl[58] vdd gnd cell_6t
Xbit_r59_c174 bl[174] br[174] wl[59] vdd gnd cell_6t
Xbit_r60_c174 bl[174] br[174] wl[60] vdd gnd cell_6t
Xbit_r61_c174 bl[174] br[174] wl[61] vdd gnd cell_6t
Xbit_r62_c174 bl[174] br[174] wl[62] vdd gnd cell_6t
Xbit_r63_c174 bl[174] br[174] wl[63] vdd gnd cell_6t
Xbit_r64_c174 bl[174] br[174] wl[64] vdd gnd cell_6t
Xbit_r65_c174 bl[174] br[174] wl[65] vdd gnd cell_6t
Xbit_r66_c174 bl[174] br[174] wl[66] vdd gnd cell_6t
Xbit_r67_c174 bl[174] br[174] wl[67] vdd gnd cell_6t
Xbit_r68_c174 bl[174] br[174] wl[68] vdd gnd cell_6t
Xbit_r69_c174 bl[174] br[174] wl[69] vdd gnd cell_6t
Xbit_r70_c174 bl[174] br[174] wl[70] vdd gnd cell_6t
Xbit_r71_c174 bl[174] br[174] wl[71] vdd gnd cell_6t
Xbit_r72_c174 bl[174] br[174] wl[72] vdd gnd cell_6t
Xbit_r73_c174 bl[174] br[174] wl[73] vdd gnd cell_6t
Xbit_r74_c174 bl[174] br[174] wl[74] vdd gnd cell_6t
Xbit_r75_c174 bl[174] br[174] wl[75] vdd gnd cell_6t
Xbit_r76_c174 bl[174] br[174] wl[76] vdd gnd cell_6t
Xbit_r77_c174 bl[174] br[174] wl[77] vdd gnd cell_6t
Xbit_r78_c174 bl[174] br[174] wl[78] vdd gnd cell_6t
Xbit_r79_c174 bl[174] br[174] wl[79] vdd gnd cell_6t
Xbit_r80_c174 bl[174] br[174] wl[80] vdd gnd cell_6t
Xbit_r81_c174 bl[174] br[174] wl[81] vdd gnd cell_6t
Xbit_r82_c174 bl[174] br[174] wl[82] vdd gnd cell_6t
Xbit_r83_c174 bl[174] br[174] wl[83] vdd gnd cell_6t
Xbit_r84_c174 bl[174] br[174] wl[84] vdd gnd cell_6t
Xbit_r85_c174 bl[174] br[174] wl[85] vdd gnd cell_6t
Xbit_r86_c174 bl[174] br[174] wl[86] vdd gnd cell_6t
Xbit_r87_c174 bl[174] br[174] wl[87] vdd gnd cell_6t
Xbit_r88_c174 bl[174] br[174] wl[88] vdd gnd cell_6t
Xbit_r89_c174 bl[174] br[174] wl[89] vdd gnd cell_6t
Xbit_r90_c174 bl[174] br[174] wl[90] vdd gnd cell_6t
Xbit_r91_c174 bl[174] br[174] wl[91] vdd gnd cell_6t
Xbit_r92_c174 bl[174] br[174] wl[92] vdd gnd cell_6t
Xbit_r93_c174 bl[174] br[174] wl[93] vdd gnd cell_6t
Xbit_r94_c174 bl[174] br[174] wl[94] vdd gnd cell_6t
Xbit_r95_c174 bl[174] br[174] wl[95] vdd gnd cell_6t
Xbit_r96_c174 bl[174] br[174] wl[96] vdd gnd cell_6t
Xbit_r97_c174 bl[174] br[174] wl[97] vdd gnd cell_6t
Xbit_r98_c174 bl[174] br[174] wl[98] vdd gnd cell_6t
Xbit_r99_c174 bl[174] br[174] wl[99] vdd gnd cell_6t
Xbit_r100_c174 bl[174] br[174] wl[100] vdd gnd cell_6t
Xbit_r101_c174 bl[174] br[174] wl[101] vdd gnd cell_6t
Xbit_r102_c174 bl[174] br[174] wl[102] vdd gnd cell_6t
Xbit_r103_c174 bl[174] br[174] wl[103] vdd gnd cell_6t
Xbit_r104_c174 bl[174] br[174] wl[104] vdd gnd cell_6t
Xbit_r105_c174 bl[174] br[174] wl[105] vdd gnd cell_6t
Xbit_r106_c174 bl[174] br[174] wl[106] vdd gnd cell_6t
Xbit_r107_c174 bl[174] br[174] wl[107] vdd gnd cell_6t
Xbit_r108_c174 bl[174] br[174] wl[108] vdd gnd cell_6t
Xbit_r109_c174 bl[174] br[174] wl[109] vdd gnd cell_6t
Xbit_r110_c174 bl[174] br[174] wl[110] vdd gnd cell_6t
Xbit_r111_c174 bl[174] br[174] wl[111] vdd gnd cell_6t
Xbit_r112_c174 bl[174] br[174] wl[112] vdd gnd cell_6t
Xbit_r113_c174 bl[174] br[174] wl[113] vdd gnd cell_6t
Xbit_r114_c174 bl[174] br[174] wl[114] vdd gnd cell_6t
Xbit_r115_c174 bl[174] br[174] wl[115] vdd gnd cell_6t
Xbit_r116_c174 bl[174] br[174] wl[116] vdd gnd cell_6t
Xbit_r117_c174 bl[174] br[174] wl[117] vdd gnd cell_6t
Xbit_r118_c174 bl[174] br[174] wl[118] vdd gnd cell_6t
Xbit_r119_c174 bl[174] br[174] wl[119] vdd gnd cell_6t
Xbit_r120_c174 bl[174] br[174] wl[120] vdd gnd cell_6t
Xbit_r121_c174 bl[174] br[174] wl[121] vdd gnd cell_6t
Xbit_r122_c174 bl[174] br[174] wl[122] vdd gnd cell_6t
Xbit_r123_c174 bl[174] br[174] wl[123] vdd gnd cell_6t
Xbit_r124_c174 bl[174] br[174] wl[124] vdd gnd cell_6t
Xbit_r125_c174 bl[174] br[174] wl[125] vdd gnd cell_6t
Xbit_r126_c174 bl[174] br[174] wl[126] vdd gnd cell_6t
Xbit_r127_c174 bl[174] br[174] wl[127] vdd gnd cell_6t
Xbit_r0_c175 bl[175] br[175] wl[0] vdd gnd cell_6t
Xbit_r1_c175 bl[175] br[175] wl[1] vdd gnd cell_6t
Xbit_r2_c175 bl[175] br[175] wl[2] vdd gnd cell_6t
Xbit_r3_c175 bl[175] br[175] wl[3] vdd gnd cell_6t
Xbit_r4_c175 bl[175] br[175] wl[4] vdd gnd cell_6t
Xbit_r5_c175 bl[175] br[175] wl[5] vdd gnd cell_6t
Xbit_r6_c175 bl[175] br[175] wl[6] vdd gnd cell_6t
Xbit_r7_c175 bl[175] br[175] wl[7] vdd gnd cell_6t
Xbit_r8_c175 bl[175] br[175] wl[8] vdd gnd cell_6t
Xbit_r9_c175 bl[175] br[175] wl[9] vdd gnd cell_6t
Xbit_r10_c175 bl[175] br[175] wl[10] vdd gnd cell_6t
Xbit_r11_c175 bl[175] br[175] wl[11] vdd gnd cell_6t
Xbit_r12_c175 bl[175] br[175] wl[12] vdd gnd cell_6t
Xbit_r13_c175 bl[175] br[175] wl[13] vdd gnd cell_6t
Xbit_r14_c175 bl[175] br[175] wl[14] vdd gnd cell_6t
Xbit_r15_c175 bl[175] br[175] wl[15] vdd gnd cell_6t
Xbit_r16_c175 bl[175] br[175] wl[16] vdd gnd cell_6t
Xbit_r17_c175 bl[175] br[175] wl[17] vdd gnd cell_6t
Xbit_r18_c175 bl[175] br[175] wl[18] vdd gnd cell_6t
Xbit_r19_c175 bl[175] br[175] wl[19] vdd gnd cell_6t
Xbit_r20_c175 bl[175] br[175] wl[20] vdd gnd cell_6t
Xbit_r21_c175 bl[175] br[175] wl[21] vdd gnd cell_6t
Xbit_r22_c175 bl[175] br[175] wl[22] vdd gnd cell_6t
Xbit_r23_c175 bl[175] br[175] wl[23] vdd gnd cell_6t
Xbit_r24_c175 bl[175] br[175] wl[24] vdd gnd cell_6t
Xbit_r25_c175 bl[175] br[175] wl[25] vdd gnd cell_6t
Xbit_r26_c175 bl[175] br[175] wl[26] vdd gnd cell_6t
Xbit_r27_c175 bl[175] br[175] wl[27] vdd gnd cell_6t
Xbit_r28_c175 bl[175] br[175] wl[28] vdd gnd cell_6t
Xbit_r29_c175 bl[175] br[175] wl[29] vdd gnd cell_6t
Xbit_r30_c175 bl[175] br[175] wl[30] vdd gnd cell_6t
Xbit_r31_c175 bl[175] br[175] wl[31] vdd gnd cell_6t
Xbit_r32_c175 bl[175] br[175] wl[32] vdd gnd cell_6t
Xbit_r33_c175 bl[175] br[175] wl[33] vdd gnd cell_6t
Xbit_r34_c175 bl[175] br[175] wl[34] vdd gnd cell_6t
Xbit_r35_c175 bl[175] br[175] wl[35] vdd gnd cell_6t
Xbit_r36_c175 bl[175] br[175] wl[36] vdd gnd cell_6t
Xbit_r37_c175 bl[175] br[175] wl[37] vdd gnd cell_6t
Xbit_r38_c175 bl[175] br[175] wl[38] vdd gnd cell_6t
Xbit_r39_c175 bl[175] br[175] wl[39] vdd gnd cell_6t
Xbit_r40_c175 bl[175] br[175] wl[40] vdd gnd cell_6t
Xbit_r41_c175 bl[175] br[175] wl[41] vdd gnd cell_6t
Xbit_r42_c175 bl[175] br[175] wl[42] vdd gnd cell_6t
Xbit_r43_c175 bl[175] br[175] wl[43] vdd gnd cell_6t
Xbit_r44_c175 bl[175] br[175] wl[44] vdd gnd cell_6t
Xbit_r45_c175 bl[175] br[175] wl[45] vdd gnd cell_6t
Xbit_r46_c175 bl[175] br[175] wl[46] vdd gnd cell_6t
Xbit_r47_c175 bl[175] br[175] wl[47] vdd gnd cell_6t
Xbit_r48_c175 bl[175] br[175] wl[48] vdd gnd cell_6t
Xbit_r49_c175 bl[175] br[175] wl[49] vdd gnd cell_6t
Xbit_r50_c175 bl[175] br[175] wl[50] vdd gnd cell_6t
Xbit_r51_c175 bl[175] br[175] wl[51] vdd gnd cell_6t
Xbit_r52_c175 bl[175] br[175] wl[52] vdd gnd cell_6t
Xbit_r53_c175 bl[175] br[175] wl[53] vdd gnd cell_6t
Xbit_r54_c175 bl[175] br[175] wl[54] vdd gnd cell_6t
Xbit_r55_c175 bl[175] br[175] wl[55] vdd gnd cell_6t
Xbit_r56_c175 bl[175] br[175] wl[56] vdd gnd cell_6t
Xbit_r57_c175 bl[175] br[175] wl[57] vdd gnd cell_6t
Xbit_r58_c175 bl[175] br[175] wl[58] vdd gnd cell_6t
Xbit_r59_c175 bl[175] br[175] wl[59] vdd gnd cell_6t
Xbit_r60_c175 bl[175] br[175] wl[60] vdd gnd cell_6t
Xbit_r61_c175 bl[175] br[175] wl[61] vdd gnd cell_6t
Xbit_r62_c175 bl[175] br[175] wl[62] vdd gnd cell_6t
Xbit_r63_c175 bl[175] br[175] wl[63] vdd gnd cell_6t
Xbit_r64_c175 bl[175] br[175] wl[64] vdd gnd cell_6t
Xbit_r65_c175 bl[175] br[175] wl[65] vdd gnd cell_6t
Xbit_r66_c175 bl[175] br[175] wl[66] vdd gnd cell_6t
Xbit_r67_c175 bl[175] br[175] wl[67] vdd gnd cell_6t
Xbit_r68_c175 bl[175] br[175] wl[68] vdd gnd cell_6t
Xbit_r69_c175 bl[175] br[175] wl[69] vdd gnd cell_6t
Xbit_r70_c175 bl[175] br[175] wl[70] vdd gnd cell_6t
Xbit_r71_c175 bl[175] br[175] wl[71] vdd gnd cell_6t
Xbit_r72_c175 bl[175] br[175] wl[72] vdd gnd cell_6t
Xbit_r73_c175 bl[175] br[175] wl[73] vdd gnd cell_6t
Xbit_r74_c175 bl[175] br[175] wl[74] vdd gnd cell_6t
Xbit_r75_c175 bl[175] br[175] wl[75] vdd gnd cell_6t
Xbit_r76_c175 bl[175] br[175] wl[76] vdd gnd cell_6t
Xbit_r77_c175 bl[175] br[175] wl[77] vdd gnd cell_6t
Xbit_r78_c175 bl[175] br[175] wl[78] vdd gnd cell_6t
Xbit_r79_c175 bl[175] br[175] wl[79] vdd gnd cell_6t
Xbit_r80_c175 bl[175] br[175] wl[80] vdd gnd cell_6t
Xbit_r81_c175 bl[175] br[175] wl[81] vdd gnd cell_6t
Xbit_r82_c175 bl[175] br[175] wl[82] vdd gnd cell_6t
Xbit_r83_c175 bl[175] br[175] wl[83] vdd gnd cell_6t
Xbit_r84_c175 bl[175] br[175] wl[84] vdd gnd cell_6t
Xbit_r85_c175 bl[175] br[175] wl[85] vdd gnd cell_6t
Xbit_r86_c175 bl[175] br[175] wl[86] vdd gnd cell_6t
Xbit_r87_c175 bl[175] br[175] wl[87] vdd gnd cell_6t
Xbit_r88_c175 bl[175] br[175] wl[88] vdd gnd cell_6t
Xbit_r89_c175 bl[175] br[175] wl[89] vdd gnd cell_6t
Xbit_r90_c175 bl[175] br[175] wl[90] vdd gnd cell_6t
Xbit_r91_c175 bl[175] br[175] wl[91] vdd gnd cell_6t
Xbit_r92_c175 bl[175] br[175] wl[92] vdd gnd cell_6t
Xbit_r93_c175 bl[175] br[175] wl[93] vdd gnd cell_6t
Xbit_r94_c175 bl[175] br[175] wl[94] vdd gnd cell_6t
Xbit_r95_c175 bl[175] br[175] wl[95] vdd gnd cell_6t
Xbit_r96_c175 bl[175] br[175] wl[96] vdd gnd cell_6t
Xbit_r97_c175 bl[175] br[175] wl[97] vdd gnd cell_6t
Xbit_r98_c175 bl[175] br[175] wl[98] vdd gnd cell_6t
Xbit_r99_c175 bl[175] br[175] wl[99] vdd gnd cell_6t
Xbit_r100_c175 bl[175] br[175] wl[100] vdd gnd cell_6t
Xbit_r101_c175 bl[175] br[175] wl[101] vdd gnd cell_6t
Xbit_r102_c175 bl[175] br[175] wl[102] vdd gnd cell_6t
Xbit_r103_c175 bl[175] br[175] wl[103] vdd gnd cell_6t
Xbit_r104_c175 bl[175] br[175] wl[104] vdd gnd cell_6t
Xbit_r105_c175 bl[175] br[175] wl[105] vdd gnd cell_6t
Xbit_r106_c175 bl[175] br[175] wl[106] vdd gnd cell_6t
Xbit_r107_c175 bl[175] br[175] wl[107] vdd gnd cell_6t
Xbit_r108_c175 bl[175] br[175] wl[108] vdd gnd cell_6t
Xbit_r109_c175 bl[175] br[175] wl[109] vdd gnd cell_6t
Xbit_r110_c175 bl[175] br[175] wl[110] vdd gnd cell_6t
Xbit_r111_c175 bl[175] br[175] wl[111] vdd gnd cell_6t
Xbit_r112_c175 bl[175] br[175] wl[112] vdd gnd cell_6t
Xbit_r113_c175 bl[175] br[175] wl[113] vdd gnd cell_6t
Xbit_r114_c175 bl[175] br[175] wl[114] vdd gnd cell_6t
Xbit_r115_c175 bl[175] br[175] wl[115] vdd gnd cell_6t
Xbit_r116_c175 bl[175] br[175] wl[116] vdd gnd cell_6t
Xbit_r117_c175 bl[175] br[175] wl[117] vdd gnd cell_6t
Xbit_r118_c175 bl[175] br[175] wl[118] vdd gnd cell_6t
Xbit_r119_c175 bl[175] br[175] wl[119] vdd gnd cell_6t
Xbit_r120_c175 bl[175] br[175] wl[120] vdd gnd cell_6t
Xbit_r121_c175 bl[175] br[175] wl[121] vdd gnd cell_6t
Xbit_r122_c175 bl[175] br[175] wl[122] vdd gnd cell_6t
Xbit_r123_c175 bl[175] br[175] wl[123] vdd gnd cell_6t
Xbit_r124_c175 bl[175] br[175] wl[124] vdd gnd cell_6t
Xbit_r125_c175 bl[175] br[175] wl[125] vdd gnd cell_6t
Xbit_r126_c175 bl[175] br[175] wl[126] vdd gnd cell_6t
Xbit_r127_c175 bl[175] br[175] wl[127] vdd gnd cell_6t
Xbit_r0_c176 bl[176] br[176] wl[0] vdd gnd cell_6t
Xbit_r1_c176 bl[176] br[176] wl[1] vdd gnd cell_6t
Xbit_r2_c176 bl[176] br[176] wl[2] vdd gnd cell_6t
Xbit_r3_c176 bl[176] br[176] wl[3] vdd gnd cell_6t
Xbit_r4_c176 bl[176] br[176] wl[4] vdd gnd cell_6t
Xbit_r5_c176 bl[176] br[176] wl[5] vdd gnd cell_6t
Xbit_r6_c176 bl[176] br[176] wl[6] vdd gnd cell_6t
Xbit_r7_c176 bl[176] br[176] wl[7] vdd gnd cell_6t
Xbit_r8_c176 bl[176] br[176] wl[8] vdd gnd cell_6t
Xbit_r9_c176 bl[176] br[176] wl[9] vdd gnd cell_6t
Xbit_r10_c176 bl[176] br[176] wl[10] vdd gnd cell_6t
Xbit_r11_c176 bl[176] br[176] wl[11] vdd gnd cell_6t
Xbit_r12_c176 bl[176] br[176] wl[12] vdd gnd cell_6t
Xbit_r13_c176 bl[176] br[176] wl[13] vdd gnd cell_6t
Xbit_r14_c176 bl[176] br[176] wl[14] vdd gnd cell_6t
Xbit_r15_c176 bl[176] br[176] wl[15] vdd gnd cell_6t
Xbit_r16_c176 bl[176] br[176] wl[16] vdd gnd cell_6t
Xbit_r17_c176 bl[176] br[176] wl[17] vdd gnd cell_6t
Xbit_r18_c176 bl[176] br[176] wl[18] vdd gnd cell_6t
Xbit_r19_c176 bl[176] br[176] wl[19] vdd gnd cell_6t
Xbit_r20_c176 bl[176] br[176] wl[20] vdd gnd cell_6t
Xbit_r21_c176 bl[176] br[176] wl[21] vdd gnd cell_6t
Xbit_r22_c176 bl[176] br[176] wl[22] vdd gnd cell_6t
Xbit_r23_c176 bl[176] br[176] wl[23] vdd gnd cell_6t
Xbit_r24_c176 bl[176] br[176] wl[24] vdd gnd cell_6t
Xbit_r25_c176 bl[176] br[176] wl[25] vdd gnd cell_6t
Xbit_r26_c176 bl[176] br[176] wl[26] vdd gnd cell_6t
Xbit_r27_c176 bl[176] br[176] wl[27] vdd gnd cell_6t
Xbit_r28_c176 bl[176] br[176] wl[28] vdd gnd cell_6t
Xbit_r29_c176 bl[176] br[176] wl[29] vdd gnd cell_6t
Xbit_r30_c176 bl[176] br[176] wl[30] vdd gnd cell_6t
Xbit_r31_c176 bl[176] br[176] wl[31] vdd gnd cell_6t
Xbit_r32_c176 bl[176] br[176] wl[32] vdd gnd cell_6t
Xbit_r33_c176 bl[176] br[176] wl[33] vdd gnd cell_6t
Xbit_r34_c176 bl[176] br[176] wl[34] vdd gnd cell_6t
Xbit_r35_c176 bl[176] br[176] wl[35] vdd gnd cell_6t
Xbit_r36_c176 bl[176] br[176] wl[36] vdd gnd cell_6t
Xbit_r37_c176 bl[176] br[176] wl[37] vdd gnd cell_6t
Xbit_r38_c176 bl[176] br[176] wl[38] vdd gnd cell_6t
Xbit_r39_c176 bl[176] br[176] wl[39] vdd gnd cell_6t
Xbit_r40_c176 bl[176] br[176] wl[40] vdd gnd cell_6t
Xbit_r41_c176 bl[176] br[176] wl[41] vdd gnd cell_6t
Xbit_r42_c176 bl[176] br[176] wl[42] vdd gnd cell_6t
Xbit_r43_c176 bl[176] br[176] wl[43] vdd gnd cell_6t
Xbit_r44_c176 bl[176] br[176] wl[44] vdd gnd cell_6t
Xbit_r45_c176 bl[176] br[176] wl[45] vdd gnd cell_6t
Xbit_r46_c176 bl[176] br[176] wl[46] vdd gnd cell_6t
Xbit_r47_c176 bl[176] br[176] wl[47] vdd gnd cell_6t
Xbit_r48_c176 bl[176] br[176] wl[48] vdd gnd cell_6t
Xbit_r49_c176 bl[176] br[176] wl[49] vdd gnd cell_6t
Xbit_r50_c176 bl[176] br[176] wl[50] vdd gnd cell_6t
Xbit_r51_c176 bl[176] br[176] wl[51] vdd gnd cell_6t
Xbit_r52_c176 bl[176] br[176] wl[52] vdd gnd cell_6t
Xbit_r53_c176 bl[176] br[176] wl[53] vdd gnd cell_6t
Xbit_r54_c176 bl[176] br[176] wl[54] vdd gnd cell_6t
Xbit_r55_c176 bl[176] br[176] wl[55] vdd gnd cell_6t
Xbit_r56_c176 bl[176] br[176] wl[56] vdd gnd cell_6t
Xbit_r57_c176 bl[176] br[176] wl[57] vdd gnd cell_6t
Xbit_r58_c176 bl[176] br[176] wl[58] vdd gnd cell_6t
Xbit_r59_c176 bl[176] br[176] wl[59] vdd gnd cell_6t
Xbit_r60_c176 bl[176] br[176] wl[60] vdd gnd cell_6t
Xbit_r61_c176 bl[176] br[176] wl[61] vdd gnd cell_6t
Xbit_r62_c176 bl[176] br[176] wl[62] vdd gnd cell_6t
Xbit_r63_c176 bl[176] br[176] wl[63] vdd gnd cell_6t
Xbit_r64_c176 bl[176] br[176] wl[64] vdd gnd cell_6t
Xbit_r65_c176 bl[176] br[176] wl[65] vdd gnd cell_6t
Xbit_r66_c176 bl[176] br[176] wl[66] vdd gnd cell_6t
Xbit_r67_c176 bl[176] br[176] wl[67] vdd gnd cell_6t
Xbit_r68_c176 bl[176] br[176] wl[68] vdd gnd cell_6t
Xbit_r69_c176 bl[176] br[176] wl[69] vdd gnd cell_6t
Xbit_r70_c176 bl[176] br[176] wl[70] vdd gnd cell_6t
Xbit_r71_c176 bl[176] br[176] wl[71] vdd gnd cell_6t
Xbit_r72_c176 bl[176] br[176] wl[72] vdd gnd cell_6t
Xbit_r73_c176 bl[176] br[176] wl[73] vdd gnd cell_6t
Xbit_r74_c176 bl[176] br[176] wl[74] vdd gnd cell_6t
Xbit_r75_c176 bl[176] br[176] wl[75] vdd gnd cell_6t
Xbit_r76_c176 bl[176] br[176] wl[76] vdd gnd cell_6t
Xbit_r77_c176 bl[176] br[176] wl[77] vdd gnd cell_6t
Xbit_r78_c176 bl[176] br[176] wl[78] vdd gnd cell_6t
Xbit_r79_c176 bl[176] br[176] wl[79] vdd gnd cell_6t
Xbit_r80_c176 bl[176] br[176] wl[80] vdd gnd cell_6t
Xbit_r81_c176 bl[176] br[176] wl[81] vdd gnd cell_6t
Xbit_r82_c176 bl[176] br[176] wl[82] vdd gnd cell_6t
Xbit_r83_c176 bl[176] br[176] wl[83] vdd gnd cell_6t
Xbit_r84_c176 bl[176] br[176] wl[84] vdd gnd cell_6t
Xbit_r85_c176 bl[176] br[176] wl[85] vdd gnd cell_6t
Xbit_r86_c176 bl[176] br[176] wl[86] vdd gnd cell_6t
Xbit_r87_c176 bl[176] br[176] wl[87] vdd gnd cell_6t
Xbit_r88_c176 bl[176] br[176] wl[88] vdd gnd cell_6t
Xbit_r89_c176 bl[176] br[176] wl[89] vdd gnd cell_6t
Xbit_r90_c176 bl[176] br[176] wl[90] vdd gnd cell_6t
Xbit_r91_c176 bl[176] br[176] wl[91] vdd gnd cell_6t
Xbit_r92_c176 bl[176] br[176] wl[92] vdd gnd cell_6t
Xbit_r93_c176 bl[176] br[176] wl[93] vdd gnd cell_6t
Xbit_r94_c176 bl[176] br[176] wl[94] vdd gnd cell_6t
Xbit_r95_c176 bl[176] br[176] wl[95] vdd gnd cell_6t
Xbit_r96_c176 bl[176] br[176] wl[96] vdd gnd cell_6t
Xbit_r97_c176 bl[176] br[176] wl[97] vdd gnd cell_6t
Xbit_r98_c176 bl[176] br[176] wl[98] vdd gnd cell_6t
Xbit_r99_c176 bl[176] br[176] wl[99] vdd gnd cell_6t
Xbit_r100_c176 bl[176] br[176] wl[100] vdd gnd cell_6t
Xbit_r101_c176 bl[176] br[176] wl[101] vdd gnd cell_6t
Xbit_r102_c176 bl[176] br[176] wl[102] vdd gnd cell_6t
Xbit_r103_c176 bl[176] br[176] wl[103] vdd gnd cell_6t
Xbit_r104_c176 bl[176] br[176] wl[104] vdd gnd cell_6t
Xbit_r105_c176 bl[176] br[176] wl[105] vdd gnd cell_6t
Xbit_r106_c176 bl[176] br[176] wl[106] vdd gnd cell_6t
Xbit_r107_c176 bl[176] br[176] wl[107] vdd gnd cell_6t
Xbit_r108_c176 bl[176] br[176] wl[108] vdd gnd cell_6t
Xbit_r109_c176 bl[176] br[176] wl[109] vdd gnd cell_6t
Xbit_r110_c176 bl[176] br[176] wl[110] vdd gnd cell_6t
Xbit_r111_c176 bl[176] br[176] wl[111] vdd gnd cell_6t
Xbit_r112_c176 bl[176] br[176] wl[112] vdd gnd cell_6t
Xbit_r113_c176 bl[176] br[176] wl[113] vdd gnd cell_6t
Xbit_r114_c176 bl[176] br[176] wl[114] vdd gnd cell_6t
Xbit_r115_c176 bl[176] br[176] wl[115] vdd gnd cell_6t
Xbit_r116_c176 bl[176] br[176] wl[116] vdd gnd cell_6t
Xbit_r117_c176 bl[176] br[176] wl[117] vdd gnd cell_6t
Xbit_r118_c176 bl[176] br[176] wl[118] vdd gnd cell_6t
Xbit_r119_c176 bl[176] br[176] wl[119] vdd gnd cell_6t
Xbit_r120_c176 bl[176] br[176] wl[120] vdd gnd cell_6t
Xbit_r121_c176 bl[176] br[176] wl[121] vdd gnd cell_6t
Xbit_r122_c176 bl[176] br[176] wl[122] vdd gnd cell_6t
Xbit_r123_c176 bl[176] br[176] wl[123] vdd gnd cell_6t
Xbit_r124_c176 bl[176] br[176] wl[124] vdd gnd cell_6t
Xbit_r125_c176 bl[176] br[176] wl[125] vdd gnd cell_6t
Xbit_r126_c176 bl[176] br[176] wl[126] vdd gnd cell_6t
Xbit_r127_c176 bl[176] br[176] wl[127] vdd gnd cell_6t
Xbit_r0_c177 bl[177] br[177] wl[0] vdd gnd cell_6t
Xbit_r1_c177 bl[177] br[177] wl[1] vdd gnd cell_6t
Xbit_r2_c177 bl[177] br[177] wl[2] vdd gnd cell_6t
Xbit_r3_c177 bl[177] br[177] wl[3] vdd gnd cell_6t
Xbit_r4_c177 bl[177] br[177] wl[4] vdd gnd cell_6t
Xbit_r5_c177 bl[177] br[177] wl[5] vdd gnd cell_6t
Xbit_r6_c177 bl[177] br[177] wl[6] vdd gnd cell_6t
Xbit_r7_c177 bl[177] br[177] wl[7] vdd gnd cell_6t
Xbit_r8_c177 bl[177] br[177] wl[8] vdd gnd cell_6t
Xbit_r9_c177 bl[177] br[177] wl[9] vdd gnd cell_6t
Xbit_r10_c177 bl[177] br[177] wl[10] vdd gnd cell_6t
Xbit_r11_c177 bl[177] br[177] wl[11] vdd gnd cell_6t
Xbit_r12_c177 bl[177] br[177] wl[12] vdd gnd cell_6t
Xbit_r13_c177 bl[177] br[177] wl[13] vdd gnd cell_6t
Xbit_r14_c177 bl[177] br[177] wl[14] vdd gnd cell_6t
Xbit_r15_c177 bl[177] br[177] wl[15] vdd gnd cell_6t
Xbit_r16_c177 bl[177] br[177] wl[16] vdd gnd cell_6t
Xbit_r17_c177 bl[177] br[177] wl[17] vdd gnd cell_6t
Xbit_r18_c177 bl[177] br[177] wl[18] vdd gnd cell_6t
Xbit_r19_c177 bl[177] br[177] wl[19] vdd gnd cell_6t
Xbit_r20_c177 bl[177] br[177] wl[20] vdd gnd cell_6t
Xbit_r21_c177 bl[177] br[177] wl[21] vdd gnd cell_6t
Xbit_r22_c177 bl[177] br[177] wl[22] vdd gnd cell_6t
Xbit_r23_c177 bl[177] br[177] wl[23] vdd gnd cell_6t
Xbit_r24_c177 bl[177] br[177] wl[24] vdd gnd cell_6t
Xbit_r25_c177 bl[177] br[177] wl[25] vdd gnd cell_6t
Xbit_r26_c177 bl[177] br[177] wl[26] vdd gnd cell_6t
Xbit_r27_c177 bl[177] br[177] wl[27] vdd gnd cell_6t
Xbit_r28_c177 bl[177] br[177] wl[28] vdd gnd cell_6t
Xbit_r29_c177 bl[177] br[177] wl[29] vdd gnd cell_6t
Xbit_r30_c177 bl[177] br[177] wl[30] vdd gnd cell_6t
Xbit_r31_c177 bl[177] br[177] wl[31] vdd gnd cell_6t
Xbit_r32_c177 bl[177] br[177] wl[32] vdd gnd cell_6t
Xbit_r33_c177 bl[177] br[177] wl[33] vdd gnd cell_6t
Xbit_r34_c177 bl[177] br[177] wl[34] vdd gnd cell_6t
Xbit_r35_c177 bl[177] br[177] wl[35] vdd gnd cell_6t
Xbit_r36_c177 bl[177] br[177] wl[36] vdd gnd cell_6t
Xbit_r37_c177 bl[177] br[177] wl[37] vdd gnd cell_6t
Xbit_r38_c177 bl[177] br[177] wl[38] vdd gnd cell_6t
Xbit_r39_c177 bl[177] br[177] wl[39] vdd gnd cell_6t
Xbit_r40_c177 bl[177] br[177] wl[40] vdd gnd cell_6t
Xbit_r41_c177 bl[177] br[177] wl[41] vdd gnd cell_6t
Xbit_r42_c177 bl[177] br[177] wl[42] vdd gnd cell_6t
Xbit_r43_c177 bl[177] br[177] wl[43] vdd gnd cell_6t
Xbit_r44_c177 bl[177] br[177] wl[44] vdd gnd cell_6t
Xbit_r45_c177 bl[177] br[177] wl[45] vdd gnd cell_6t
Xbit_r46_c177 bl[177] br[177] wl[46] vdd gnd cell_6t
Xbit_r47_c177 bl[177] br[177] wl[47] vdd gnd cell_6t
Xbit_r48_c177 bl[177] br[177] wl[48] vdd gnd cell_6t
Xbit_r49_c177 bl[177] br[177] wl[49] vdd gnd cell_6t
Xbit_r50_c177 bl[177] br[177] wl[50] vdd gnd cell_6t
Xbit_r51_c177 bl[177] br[177] wl[51] vdd gnd cell_6t
Xbit_r52_c177 bl[177] br[177] wl[52] vdd gnd cell_6t
Xbit_r53_c177 bl[177] br[177] wl[53] vdd gnd cell_6t
Xbit_r54_c177 bl[177] br[177] wl[54] vdd gnd cell_6t
Xbit_r55_c177 bl[177] br[177] wl[55] vdd gnd cell_6t
Xbit_r56_c177 bl[177] br[177] wl[56] vdd gnd cell_6t
Xbit_r57_c177 bl[177] br[177] wl[57] vdd gnd cell_6t
Xbit_r58_c177 bl[177] br[177] wl[58] vdd gnd cell_6t
Xbit_r59_c177 bl[177] br[177] wl[59] vdd gnd cell_6t
Xbit_r60_c177 bl[177] br[177] wl[60] vdd gnd cell_6t
Xbit_r61_c177 bl[177] br[177] wl[61] vdd gnd cell_6t
Xbit_r62_c177 bl[177] br[177] wl[62] vdd gnd cell_6t
Xbit_r63_c177 bl[177] br[177] wl[63] vdd gnd cell_6t
Xbit_r64_c177 bl[177] br[177] wl[64] vdd gnd cell_6t
Xbit_r65_c177 bl[177] br[177] wl[65] vdd gnd cell_6t
Xbit_r66_c177 bl[177] br[177] wl[66] vdd gnd cell_6t
Xbit_r67_c177 bl[177] br[177] wl[67] vdd gnd cell_6t
Xbit_r68_c177 bl[177] br[177] wl[68] vdd gnd cell_6t
Xbit_r69_c177 bl[177] br[177] wl[69] vdd gnd cell_6t
Xbit_r70_c177 bl[177] br[177] wl[70] vdd gnd cell_6t
Xbit_r71_c177 bl[177] br[177] wl[71] vdd gnd cell_6t
Xbit_r72_c177 bl[177] br[177] wl[72] vdd gnd cell_6t
Xbit_r73_c177 bl[177] br[177] wl[73] vdd gnd cell_6t
Xbit_r74_c177 bl[177] br[177] wl[74] vdd gnd cell_6t
Xbit_r75_c177 bl[177] br[177] wl[75] vdd gnd cell_6t
Xbit_r76_c177 bl[177] br[177] wl[76] vdd gnd cell_6t
Xbit_r77_c177 bl[177] br[177] wl[77] vdd gnd cell_6t
Xbit_r78_c177 bl[177] br[177] wl[78] vdd gnd cell_6t
Xbit_r79_c177 bl[177] br[177] wl[79] vdd gnd cell_6t
Xbit_r80_c177 bl[177] br[177] wl[80] vdd gnd cell_6t
Xbit_r81_c177 bl[177] br[177] wl[81] vdd gnd cell_6t
Xbit_r82_c177 bl[177] br[177] wl[82] vdd gnd cell_6t
Xbit_r83_c177 bl[177] br[177] wl[83] vdd gnd cell_6t
Xbit_r84_c177 bl[177] br[177] wl[84] vdd gnd cell_6t
Xbit_r85_c177 bl[177] br[177] wl[85] vdd gnd cell_6t
Xbit_r86_c177 bl[177] br[177] wl[86] vdd gnd cell_6t
Xbit_r87_c177 bl[177] br[177] wl[87] vdd gnd cell_6t
Xbit_r88_c177 bl[177] br[177] wl[88] vdd gnd cell_6t
Xbit_r89_c177 bl[177] br[177] wl[89] vdd gnd cell_6t
Xbit_r90_c177 bl[177] br[177] wl[90] vdd gnd cell_6t
Xbit_r91_c177 bl[177] br[177] wl[91] vdd gnd cell_6t
Xbit_r92_c177 bl[177] br[177] wl[92] vdd gnd cell_6t
Xbit_r93_c177 bl[177] br[177] wl[93] vdd gnd cell_6t
Xbit_r94_c177 bl[177] br[177] wl[94] vdd gnd cell_6t
Xbit_r95_c177 bl[177] br[177] wl[95] vdd gnd cell_6t
Xbit_r96_c177 bl[177] br[177] wl[96] vdd gnd cell_6t
Xbit_r97_c177 bl[177] br[177] wl[97] vdd gnd cell_6t
Xbit_r98_c177 bl[177] br[177] wl[98] vdd gnd cell_6t
Xbit_r99_c177 bl[177] br[177] wl[99] vdd gnd cell_6t
Xbit_r100_c177 bl[177] br[177] wl[100] vdd gnd cell_6t
Xbit_r101_c177 bl[177] br[177] wl[101] vdd gnd cell_6t
Xbit_r102_c177 bl[177] br[177] wl[102] vdd gnd cell_6t
Xbit_r103_c177 bl[177] br[177] wl[103] vdd gnd cell_6t
Xbit_r104_c177 bl[177] br[177] wl[104] vdd gnd cell_6t
Xbit_r105_c177 bl[177] br[177] wl[105] vdd gnd cell_6t
Xbit_r106_c177 bl[177] br[177] wl[106] vdd gnd cell_6t
Xbit_r107_c177 bl[177] br[177] wl[107] vdd gnd cell_6t
Xbit_r108_c177 bl[177] br[177] wl[108] vdd gnd cell_6t
Xbit_r109_c177 bl[177] br[177] wl[109] vdd gnd cell_6t
Xbit_r110_c177 bl[177] br[177] wl[110] vdd gnd cell_6t
Xbit_r111_c177 bl[177] br[177] wl[111] vdd gnd cell_6t
Xbit_r112_c177 bl[177] br[177] wl[112] vdd gnd cell_6t
Xbit_r113_c177 bl[177] br[177] wl[113] vdd gnd cell_6t
Xbit_r114_c177 bl[177] br[177] wl[114] vdd gnd cell_6t
Xbit_r115_c177 bl[177] br[177] wl[115] vdd gnd cell_6t
Xbit_r116_c177 bl[177] br[177] wl[116] vdd gnd cell_6t
Xbit_r117_c177 bl[177] br[177] wl[117] vdd gnd cell_6t
Xbit_r118_c177 bl[177] br[177] wl[118] vdd gnd cell_6t
Xbit_r119_c177 bl[177] br[177] wl[119] vdd gnd cell_6t
Xbit_r120_c177 bl[177] br[177] wl[120] vdd gnd cell_6t
Xbit_r121_c177 bl[177] br[177] wl[121] vdd gnd cell_6t
Xbit_r122_c177 bl[177] br[177] wl[122] vdd gnd cell_6t
Xbit_r123_c177 bl[177] br[177] wl[123] vdd gnd cell_6t
Xbit_r124_c177 bl[177] br[177] wl[124] vdd gnd cell_6t
Xbit_r125_c177 bl[177] br[177] wl[125] vdd gnd cell_6t
Xbit_r126_c177 bl[177] br[177] wl[126] vdd gnd cell_6t
Xbit_r127_c177 bl[177] br[177] wl[127] vdd gnd cell_6t
Xbit_r0_c178 bl[178] br[178] wl[0] vdd gnd cell_6t
Xbit_r1_c178 bl[178] br[178] wl[1] vdd gnd cell_6t
Xbit_r2_c178 bl[178] br[178] wl[2] vdd gnd cell_6t
Xbit_r3_c178 bl[178] br[178] wl[3] vdd gnd cell_6t
Xbit_r4_c178 bl[178] br[178] wl[4] vdd gnd cell_6t
Xbit_r5_c178 bl[178] br[178] wl[5] vdd gnd cell_6t
Xbit_r6_c178 bl[178] br[178] wl[6] vdd gnd cell_6t
Xbit_r7_c178 bl[178] br[178] wl[7] vdd gnd cell_6t
Xbit_r8_c178 bl[178] br[178] wl[8] vdd gnd cell_6t
Xbit_r9_c178 bl[178] br[178] wl[9] vdd gnd cell_6t
Xbit_r10_c178 bl[178] br[178] wl[10] vdd gnd cell_6t
Xbit_r11_c178 bl[178] br[178] wl[11] vdd gnd cell_6t
Xbit_r12_c178 bl[178] br[178] wl[12] vdd gnd cell_6t
Xbit_r13_c178 bl[178] br[178] wl[13] vdd gnd cell_6t
Xbit_r14_c178 bl[178] br[178] wl[14] vdd gnd cell_6t
Xbit_r15_c178 bl[178] br[178] wl[15] vdd gnd cell_6t
Xbit_r16_c178 bl[178] br[178] wl[16] vdd gnd cell_6t
Xbit_r17_c178 bl[178] br[178] wl[17] vdd gnd cell_6t
Xbit_r18_c178 bl[178] br[178] wl[18] vdd gnd cell_6t
Xbit_r19_c178 bl[178] br[178] wl[19] vdd gnd cell_6t
Xbit_r20_c178 bl[178] br[178] wl[20] vdd gnd cell_6t
Xbit_r21_c178 bl[178] br[178] wl[21] vdd gnd cell_6t
Xbit_r22_c178 bl[178] br[178] wl[22] vdd gnd cell_6t
Xbit_r23_c178 bl[178] br[178] wl[23] vdd gnd cell_6t
Xbit_r24_c178 bl[178] br[178] wl[24] vdd gnd cell_6t
Xbit_r25_c178 bl[178] br[178] wl[25] vdd gnd cell_6t
Xbit_r26_c178 bl[178] br[178] wl[26] vdd gnd cell_6t
Xbit_r27_c178 bl[178] br[178] wl[27] vdd gnd cell_6t
Xbit_r28_c178 bl[178] br[178] wl[28] vdd gnd cell_6t
Xbit_r29_c178 bl[178] br[178] wl[29] vdd gnd cell_6t
Xbit_r30_c178 bl[178] br[178] wl[30] vdd gnd cell_6t
Xbit_r31_c178 bl[178] br[178] wl[31] vdd gnd cell_6t
Xbit_r32_c178 bl[178] br[178] wl[32] vdd gnd cell_6t
Xbit_r33_c178 bl[178] br[178] wl[33] vdd gnd cell_6t
Xbit_r34_c178 bl[178] br[178] wl[34] vdd gnd cell_6t
Xbit_r35_c178 bl[178] br[178] wl[35] vdd gnd cell_6t
Xbit_r36_c178 bl[178] br[178] wl[36] vdd gnd cell_6t
Xbit_r37_c178 bl[178] br[178] wl[37] vdd gnd cell_6t
Xbit_r38_c178 bl[178] br[178] wl[38] vdd gnd cell_6t
Xbit_r39_c178 bl[178] br[178] wl[39] vdd gnd cell_6t
Xbit_r40_c178 bl[178] br[178] wl[40] vdd gnd cell_6t
Xbit_r41_c178 bl[178] br[178] wl[41] vdd gnd cell_6t
Xbit_r42_c178 bl[178] br[178] wl[42] vdd gnd cell_6t
Xbit_r43_c178 bl[178] br[178] wl[43] vdd gnd cell_6t
Xbit_r44_c178 bl[178] br[178] wl[44] vdd gnd cell_6t
Xbit_r45_c178 bl[178] br[178] wl[45] vdd gnd cell_6t
Xbit_r46_c178 bl[178] br[178] wl[46] vdd gnd cell_6t
Xbit_r47_c178 bl[178] br[178] wl[47] vdd gnd cell_6t
Xbit_r48_c178 bl[178] br[178] wl[48] vdd gnd cell_6t
Xbit_r49_c178 bl[178] br[178] wl[49] vdd gnd cell_6t
Xbit_r50_c178 bl[178] br[178] wl[50] vdd gnd cell_6t
Xbit_r51_c178 bl[178] br[178] wl[51] vdd gnd cell_6t
Xbit_r52_c178 bl[178] br[178] wl[52] vdd gnd cell_6t
Xbit_r53_c178 bl[178] br[178] wl[53] vdd gnd cell_6t
Xbit_r54_c178 bl[178] br[178] wl[54] vdd gnd cell_6t
Xbit_r55_c178 bl[178] br[178] wl[55] vdd gnd cell_6t
Xbit_r56_c178 bl[178] br[178] wl[56] vdd gnd cell_6t
Xbit_r57_c178 bl[178] br[178] wl[57] vdd gnd cell_6t
Xbit_r58_c178 bl[178] br[178] wl[58] vdd gnd cell_6t
Xbit_r59_c178 bl[178] br[178] wl[59] vdd gnd cell_6t
Xbit_r60_c178 bl[178] br[178] wl[60] vdd gnd cell_6t
Xbit_r61_c178 bl[178] br[178] wl[61] vdd gnd cell_6t
Xbit_r62_c178 bl[178] br[178] wl[62] vdd gnd cell_6t
Xbit_r63_c178 bl[178] br[178] wl[63] vdd gnd cell_6t
Xbit_r64_c178 bl[178] br[178] wl[64] vdd gnd cell_6t
Xbit_r65_c178 bl[178] br[178] wl[65] vdd gnd cell_6t
Xbit_r66_c178 bl[178] br[178] wl[66] vdd gnd cell_6t
Xbit_r67_c178 bl[178] br[178] wl[67] vdd gnd cell_6t
Xbit_r68_c178 bl[178] br[178] wl[68] vdd gnd cell_6t
Xbit_r69_c178 bl[178] br[178] wl[69] vdd gnd cell_6t
Xbit_r70_c178 bl[178] br[178] wl[70] vdd gnd cell_6t
Xbit_r71_c178 bl[178] br[178] wl[71] vdd gnd cell_6t
Xbit_r72_c178 bl[178] br[178] wl[72] vdd gnd cell_6t
Xbit_r73_c178 bl[178] br[178] wl[73] vdd gnd cell_6t
Xbit_r74_c178 bl[178] br[178] wl[74] vdd gnd cell_6t
Xbit_r75_c178 bl[178] br[178] wl[75] vdd gnd cell_6t
Xbit_r76_c178 bl[178] br[178] wl[76] vdd gnd cell_6t
Xbit_r77_c178 bl[178] br[178] wl[77] vdd gnd cell_6t
Xbit_r78_c178 bl[178] br[178] wl[78] vdd gnd cell_6t
Xbit_r79_c178 bl[178] br[178] wl[79] vdd gnd cell_6t
Xbit_r80_c178 bl[178] br[178] wl[80] vdd gnd cell_6t
Xbit_r81_c178 bl[178] br[178] wl[81] vdd gnd cell_6t
Xbit_r82_c178 bl[178] br[178] wl[82] vdd gnd cell_6t
Xbit_r83_c178 bl[178] br[178] wl[83] vdd gnd cell_6t
Xbit_r84_c178 bl[178] br[178] wl[84] vdd gnd cell_6t
Xbit_r85_c178 bl[178] br[178] wl[85] vdd gnd cell_6t
Xbit_r86_c178 bl[178] br[178] wl[86] vdd gnd cell_6t
Xbit_r87_c178 bl[178] br[178] wl[87] vdd gnd cell_6t
Xbit_r88_c178 bl[178] br[178] wl[88] vdd gnd cell_6t
Xbit_r89_c178 bl[178] br[178] wl[89] vdd gnd cell_6t
Xbit_r90_c178 bl[178] br[178] wl[90] vdd gnd cell_6t
Xbit_r91_c178 bl[178] br[178] wl[91] vdd gnd cell_6t
Xbit_r92_c178 bl[178] br[178] wl[92] vdd gnd cell_6t
Xbit_r93_c178 bl[178] br[178] wl[93] vdd gnd cell_6t
Xbit_r94_c178 bl[178] br[178] wl[94] vdd gnd cell_6t
Xbit_r95_c178 bl[178] br[178] wl[95] vdd gnd cell_6t
Xbit_r96_c178 bl[178] br[178] wl[96] vdd gnd cell_6t
Xbit_r97_c178 bl[178] br[178] wl[97] vdd gnd cell_6t
Xbit_r98_c178 bl[178] br[178] wl[98] vdd gnd cell_6t
Xbit_r99_c178 bl[178] br[178] wl[99] vdd gnd cell_6t
Xbit_r100_c178 bl[178] br[178] wl[100] vdd gnd cell_6t
Xbit_r101_c178 bl[178] br[178] wl[101] vdd gnd cell_6t
Xbit_r102_c178 bl[178] br[178] wl[102] vdd gnd cell_6t
Xbit_r103_c178 bl[178] br[178] wl[103] vdd gnd cell_6t
Xbit_r104_c178 bl[178] br[178] wl[104] vdd gnd cell_6t
Xbit_r105_c178 bl[178] br[178] wl[105] vdd gnd cell_6t
Xbit_r106_c178 bl[178] br[178] wl[106] vdd gnd cell_6t
Xbit_r107_c178 bl[178] br[178] wl[107] vdd gnd cell_6t
Xbit_r108_c178 bl[178] br[178] wl[108] vdd gnd cell_6t
Xbit_r109_c178 bl[178] br[178] wl[109] vdd gnd cell_6t
Xbit_r110_c178 bl[178] br[178] wl[110] vdd gnd cell_6t
Xbit_r111_c178 bl[178] br[178] wl[111] vdd gnd cell_6t
Xbit_r112_c178 bl[178] br[178] wl[112] vdd gnd cell_6t
Xbit_r113_c178 bl[178] br[178] wl[113] vdd gnd cell_6t
Xbit_r114_c178 bl[178] br[178] wl[114] vdd gnd cell_6t
Xbit_r115_c178 bl[178] br[178] wl[115] vdd gnd cell_6t
Xbit_r116_c178 bl[178] br[178] wl[116] vdd gnd cell_6t
Xbit_r117_c178 bl[178] br[178] wl[117] vdd gnd cell_6t
Xbit_r118_c178 bl[178] br[178] wl[118] vdd gnd cell_6t
Xbit_r119_c178 bl[178] br[178] wl[119] vdd gnd cell_6t
Xbit_r120_c178 bl[178] br[178] wl[120] vdd gnd cell_6t
Xbit_r121_c178 bl[178] br[178] wl[121] vdd gnd cell_6t
Xbit_r122_c178 bl[178] br[178] wl[122] vdd gnd cell_6t
Xbit_r123_c178 bl[178] br[178] wl[123] vdd gnd cell_6t
Xbit_r124_c178 bl[178] br[178] wl[124] vdd gnd cell_6t
Xbit_r125_c178 bl[178] br[178] wl[125] vdd gnd cell_6t
Xbit_r126_c178 bl[178] br[178] wl[126] vdd gnd cell_6t
Xbit_r127_c178 bl[178] br[178] wl[127] vdd gnd cell_6t
Xbit_r0_c179 bl[179] br[179] wl[0] vdd gnd cell_6t
Xbit_r1_c179 bl[179] br[179] wl[1] vdd gnd cell_6t
Xbit_r2_c179 bl[179] br[179] wl[2] vdd gnd cell_6t
Xbit_r3_c179 bl[179] br[179] wl[3] vdd gnd cell_6t
Xbit_r4_c179 bl[179] br[179] wl[4] vdd gnd cell_6t
Xbit_r5_c179 bl[179] br[179] wl[5] vdd gnd cell_6t
Xbit_r6_c179 bl[179] br[179] wl[6] vdd gnd cell_6t
Xbit_r7_c179 bl[179] br[179] wl[7] vdd gnd cell_6t
Xbit_r8_c179 bl[179] br[179] wl[8] vdd gnd cell_6t
Xbit_r9_c179 bl[179] br[179] wl[9] vdd gnd cell_6t
Xbit_r10_c179 bl[179] br[179] wl[10] vdd gnd cell_6t
Xbit_r11_c179 bl[179] br[179] wl[11] vdd gnd cell_6t
Xbit_r12_c179 bl[179] br[179] wl[12] vdd gnd cell_6t
Xbit_r13_c179 bl[179] br[179] wl[13] vdd gnd cell_6t
Xbit_r14_c179 bl[179] br[179] wl[14] vdd gnd cell_6t
Xbit_r15_c179 bl[179] br[179] wl[15] vdd gnd cell_6t
Xbit_r16_c179 bl[179] br[179] wl[16] vdd gnd cell_6t
Xbit_r17_c179 bl[179] br[179] wl[17] vdd gnd cell_6t
Xbit_r18_c179 bl[179] br[179] wl[18] vdd gnd cell_6t
Xbit_r19_c179 bl[179] br[179] wl[19] vdd gnd cell_6t
Xbit_r20_c179 bl[179] br[179] wl[20] vdd gnd cell_6t
Xbit_r21_c179 bl[179] br[179] wl[21] vdd gnd cell_6t
Xbit_r22_c179 bl[179] br[179] wl[22] vdd gnd cell_6t
Xbit_r23_c179 bl[179] br[179] wl[23] vdd gnd cell_6t
Xbit_r24_c179 bl[179] br[179] wl[24] vdd gnd cell_6t
Xbit_r25_c179 bl[179] br[179] wl[25] vdd gnd cell_6t
Xbit_r26_c179 bl[179] br[179] wl[26] vdd gnd cell_6t
Xbit_r27_c179 bl[179] br[179] wl[27] vdd gnd cell_6t
Xbit_r28_c179 bl[179] br[179] wl[28] vdd gnd cell_6t
Xbit_r29_c179 bl[179] br[179] wl[29] vdd gnd cell_6t
Xbit_r30_c179 bl[179] br[179] wl[30] vdd gnd cell_6t
Xbit_r31_c179 bl[179] br[179] wl[31] vdd gnd cell_6t
Xbit_r32_c179 bl[179] br[179] wl[32] vdd gnd cell_6t
Xbit_r33_c179 bl[179] br[179] wl[33] vdd gnd cell_6t
Xbit_r34_c179 bl[179] br[179] wl[34] vdd gnd cell_6t
Xbit_r35_c179 bl[179] br[179] wl[35] vdd gnd cell_6t
Xbit_r36_c179 bl[179] br[179] wl[36] vdd gnd cell_6t
Xbit_r37_c179 bl[179] br[179] wl[37] vdd gnd cell_6t
Xbit_r38_c179 bl[179] br[179] wl[38] vdd gnd cell_6t
Xbit_r39_c179 bl[179] br[179] wl[39] vdd gnd cell_6t
Xbit_r40_c179 bl[179] br[179] wl[40] vdd gnd cell_6t
Xbit_r41_c179 bl[179] br[179] wl[41] vdd gnd cell_6t
Xbit_r42_c179 bl[179] br[179] wl[42] vdd gnd cell_6t
Xbit_r43_c179 bl[179] br[179] wl[43] vdd gnd cell_6t
Xbit_r44_c179 bl[179] br[179] wl[44] vdd gnd cell_6t
Xbit_r45_c179 bl[179] br[179] wl[45] vdd gnd cell_6t
Xbit_r46_c179 bl[179] br[179] wl[46] vdd gnd cell_6t
Xbit_r47_c179 bl[179] br[179] wl[47] vdd gnd cell_6t
Xbit_r48_c179 bl[179] br[179] wl[48] vdd gnd cell_6t
Xbit_r49_c179 bl[179] br[179] wl[49] vdd gnd cell_6t
Xbit_r50_c179 bl[179] br[179] wl[50] vdd gnd cell_6t
Xbit_r51_c179 bl[179] br[179] wl[51] vdd gnd cell_6t
Xbit_r52_c179 bl[179] br[179] wl[52] vdd gnd cell_6t
Xbit_r53_c179 bl[179] br[179] wl[53] vdd gnd cell_6t
Xbit_r54_c179 bl[179] br[179] wl[54] vdd gnd cell_6t
Xbit_r55_c179 bl[179] br[179] wl[55] vdd gnd cell_6t
Xbit_r56_c179 bl[179] br[179] wl[56] vdd gnd cell_6t
Xbit_r57_c179 bl[179] br[179] wl[57] vdd gnd cell_6t
Xbit_r58_c179 bl[179] br[179] wl[58] vdd gnd cell_6t
Xbit_r59_c179 bl[179] br[179] wl[59] vdd gnd cell_6t
Xbit_r60_c179 bl[179] br[179] wl[60] vdd gnd cell_6t
Xbit_r61_c179 bl[179] br[179] wl[61] vdd gnd cell_6t
Xbit_r62_c179 bl[179] br[179] wl[62] vdd gnd cell_6t
Xbit_r63_c179 bl[179] br[179] wl[63] vdd gnd cell_6t
Xbit_r64_c179 bl[179] br[179] wl[64] vdd gnd cell_6t
Xbit_r65_c179 bl[179] br[179] wl[65] vdd gnd cell_6t
Xbit_r66_c179 bl[179] br[179] wl[66] vdd gnd cell_6t
Xbit_r67_c179 bl[179] br[179] wl[67] vdd gnd cell_6t
Xbit_r68_c179 bl[179] br[179] wl[68] vdd gnd cell_6t
Xbit_r69_c179 bl[179] br[179] wl[69] vdd gnd cell_6t
Xbit_r70_c179 bl[179] br[179] wl[70] vdd gnd cell_6t
Xbit_r71_c179 bl[179] br[179] wl[71] vdd gnd cell_6t
Xbit_r72_c179 bl[179] br[179] wl[72] vdd gnd cell_6t
Xbit_r73_c179 bl[179] br[179] wl[73] vdd gnd cell_6t
Xbit_r74_c179 bl[179] br[179] wl[74] vdd gnd cell_6t
Xbit_r75_c179 bl[179] br[179] wl[75] vdd gnd cell_6t
Xbit_r76_c179 bl[179] br[179] wl[76] vdd gnd cell_6t
Xbit_r77_c179 bl[179] br[179] wl[77] vdd gnd cell_6t
Xbit_r78_c179 bl[179] br[179] wl[78] vdd gnd cell_6t
Xbit_r79_c179 bl[179] br[179] wl[79] vdd gnd cell_6t
Xbit_r80_c179 bl[179] br[179] wl[80] vdd gnd cell_6t
Xbit_r81_c179 bl[179] br[179] wl[81] vdd gnd cell_6t
Xbit_r82_c179 bl[179] br[179] wl[82] vdd gnd cell_6t
Xbit_r83_c179 bl[179] br[179] wl[83] vdd gnd cell_6t
Xbit_r84_c179 bl[179] br[179] wl[84] vdd gnd cell_6t
Xbit_r85_c179 bl[179] br[179] wl[85] vdd gnd cell_6t
Xbit_r86_c179 bl[179] br[179] wl[86] vdd gnd cell_6t
Xbit_r87_c179 bl[179] br[179] wl[87] vdd gnd cell_6t
Xbit_r88_c179 bl[179] br[179] wl[88] vdd gnd cell_6t
Xbit_r89_c179 bl[179] br[179] wl[89] vdd gnd cell_6t
Xbit_r90_c179 bl[179] br[179] wl[90] vdd gnd cell_6t
Xbit_r91_c179 bl[179] br[179] wl[91] vdd gnd cell_6t
Xbit_r92_c179 bl[179] br[179] wl[92] vdd gnd cell_6t
Xbit_r93_c179 bl[179] br[179] wl[93] vdd gnd cell_6t
Xbit_r94_c179 bl[179] br[179] wl[94] vdd gnd cell_6t
Xbit_r95_c179 bl[179] br[179] wl[95] vdd gnd cell_6t
Xbit_r96_c179 bl[179] br[179] wl[96] vdd gnd cell_6t
Xbit_r97_c179 bl[179] br[179] wl[97] vdd gnd cell_6t
Xbit_r98_c179 bl[179] br[179] wl[98] vdd gnd cell_6t
Xbit_r99_c179 bl[179] br[179] wl[99] vdd gnd cell_6t
Xbit_r100_c179 bl[179] br[179] wl[100] vdd gnd cell_6t
Xbit_r101_c179 bl[179] br[179] wl[101] vdd gnd cell_6t
Xbit_r102_c179 bl[179] br[179] wl[102] vdd gnd cell_6t
Xbit_r103_c179 bl[179] br[179] wl[103] vdd gnd cell_6t
Xbit_r104_c179 bl[179] br[179] wl[104] vdd gnd cell_6t
Xbit_r105_c179 bl[179] br[179] wl[105] vdd gnd cell_6t
Xbit_r106_c179 bl[179] br[179] wl[106] vdd gnd cell_6t
Xbit_r107_c179 bl[179] br[179] wl[107] vdd gnd cell_6t
Xbit_r108_c179 bl[179] br[179] wl[108] vdd gnd cell_6t
Xbit_r109_c179 bl[179] br[179] wl[109] vdd gnd cell_6t
Xbit_r110_c179 bl[179] br[179] wl[110] vdd gnd cell_6t
Xbit_r111_c179 bl[179] br[179] wl[111] vdd gnd cell_6t
Xbit_r112_c179 bl[179] br[179] wl[112] vdd gnd cell_6t
Xbit_r113_c179 bl[179] br[179] wl[113] vdd gnd cell_6t
Xbit_r114_c179 bl[179] br[179] wl[114] vdd gnd cell_6t
Xbit_r115_c179 bl[179] br[179] wl[115] vdd gnd cell_6t
Xbit_r116_c179 bl[179] br[179] wl[116] vdd gnd cell_6t
Xbit_r117_c179 bl[179] br[179] wl[117] vdd gnd cell_6t
Xbit_r118_c179 bl[179] br[179] wl[118] vdd gnd cell_6t
Xbit_r119_c179 bl[179] br[179] wl[119] vdd gnd cell_6t
Xbit_r120_c179 bl[179] br[179] wl[120] vdd gnd cell_6t
Xbit_r121_c179 bl[179] br[179] wl[121] vdd gnd cell_6t
Xbit_r122_c179 bl[179] br[179] wl[122] vdd gnd cell_6t
Xbit_r123_c179 bl[179] br[179] wl[123] vdd gnd cell_6t
Xbit_r124_c179 bl[179] br[179] wl[124] vdd gnd cell_6t
Xbit_r125_c179 bl[179] br[179] wl[125] vdd gnd cell_6t
Xbit_r126_c179 bl[179] br[179] wl[126] vdd gnd cell_6t
Xbit_r127_c179 bl[179] br[179] wl[127] vdd gnd cell_6t
Xbit_r0_c180 bl[180] br[180] wl[0] vdd gnd cell_6t
Xbit_r1_c180 bl[180] br[180] wl[1] vdd gnd cell_6t
Xbit_r2_c180 bl[180] br[180] wl[2] vdd gnd cell_6t
Xbit_r3_c180 bl[180] br[180] wl[3] vdd gnd cell_6t
Xbit_r4_c180 bl[180] br[180] wl[4] vdd gnd cell_6t
Xbit_r5_c180 bl[180] br[180] wl[5] vdd gnd cell_6t
Xbit_r6_c180 bl[180] br[180] wl[6] vdd gnd cell_6t
Xbit_r7_c180 bl[180] br[180] wl[7] vdd gnd cell_6t
Xbit_r8_c180 bl[180] br[180] wl[8] vdd gnd cell_6t
Xbit_r9_c180 bl[180] br[180] wl[9] vdd gnd cell_6t
Xbit_r10_c180 bl[180] br[180] wl[10] vdd gnd cell_6t
Xbit_r11_c180 bl[180] br[180] wl[11] vdd gnd cell_6t
Xbit_r12_c180 bl[180] br[180] wl[12] vdd gnd cell_6t
Xbit_r13_c180 bl[180] br[180] wl[13] vdd gnd cell_6t
Xbit_r14_c180 bl[180] br[180] wl[14] vdd gnd cell_6t
Xbit_r15_c180 bl[180] br[180] wl[15] vdd gnd cell_6t
Xbit_r16_c180 bl[180] br[180] wl[16] vdd gnd cell_6t
Xbit_r17_c180 bl[180] br[180] wl[17] vdd gnd cell_6t
Xbit_r18_c180 bl[180] br[180] wl[18] vdd gnd cell_6t
Xbit_r19_c180 bl[180] br[180] wl[19] vdd gnd cell_6t
Xbit_r20_c180 bl[180] br[180] wl[20] vdd gnd cell_6t
Xbit_r21_c180 bl[180] br[180] wl[21] vdd gnd cell_6t
Xbit_r22_c180 bl[180] br[180] wl[22] vdd gnd cell_6t
Xbit_r23_c180 bl[180] br[180] wl[23] vdd gnd cell_6t
Xbit_r24_c180 bl[180] br[180] wl[24] vdd gnd cell_6t
Xbit_r25_c180 bl[180] br[180] wl[25] vdd gnd cell_6t
Xbit_r26_c180 bl[180] br[180] wl[26] vdd gnd cell_6t
Xbit_r27_c180 bl[180] br[180] wl[27] vdd gnd cell_6t
Xbit_r28_c180 bl[180] br[180] wl[28] vdd gnd cell_6t
Xbit_r29_c180 bl[180] br[180] wl[29] vdd gnd cell_6t
Xbit_r30_c180 bl[180] br[180] wl[30] vdd gnd cell_6t
Xbit_r31_c180 bl[180] br[180] wl[31] vdd gnd cell_6t
Xbit_r32_c180 bl[180] br[180] wl[32] vdd gnd cell_6t
Xbit_r33_c180 bl[180] br[180] wl[33] vdd gnd cell_6t
Xbit_r34_c180 bl[180] br[180] wl[34] vdd gnd cell_6t
Xbit_r35_c180 bl[180] br[180] wl[35] vdd gnd cell_6t
Xbit_r36_c180 bl[180] br[180] wl[36] vdd gnd cell_6t
Xbit_r37_c180 bl[180] br[180] wl[37] vdd gnd cell_6t
Xbit_r38_c180 bl[180] br[180] wl[38] vdd gnd cell_6t
Xbit_r39_c180 bl[180] br[180] wl[39] vdd gnd cell_6t
Xbit_r40_c180 bl[180] br[180] wl[40] vdd gnd cell_6t
Xbit_r41_c180 bl[180] br[180] wl[41] vdd gnd cell_6t
Xbit_r42_c180 bl[180] br[180] wl[42] vdd gnd cell_6t
Xbit_r43_c180 bl[180] br[180] wl[43] vdd gnd cell_6t
Xbit_r44_c180 bl[180] br[180] wl[44] vdd gnd cell_6t
Xbit_r45_c180 bl[180] br[180] wl[45] vdd gnd cell_6t
Xbit_r46_c180 bl[180] br[180] wl[46] vdd gnd cell_6t
Xbit_r47_c180 bl[180] br[180] wl[47] vdd gnd cell_6t
Xbit_r48_c180 bl[180] br[180] wl[48] vdd gnd cell_6t
Xbit_r49_c180 bl[180] br[180] wl[49] vdd gnd cell_6t
Xbit_r50_c180 bl[180] br[180] wl[50] vdd gnd cell_6t
Xbit_r51_c180 bl[180] br[180] wl[51] vdd gnd cell_6t
Xbit_r52_c180 bl[180] br[180] wl[52] vdd gnd cell_6t
Xbit_r53_c180 bl[180] br[180] wl[53] vdd gnd cell_6t
Xbit_r54_c180 bl[180] br[180] wl[54] vdd gnd cell_6t
Xbit_r55_c180 bl[180] br[180] wl[55] vdd gnd cell_6t
Xbit_r56_c180 bl[180] br[180] wl[56] vdd gnd cell_6t
Xbit_r57_c180 bl[180] br[180] wl[57] vdd gnd cell_6t
Xbit_r58_c180 bl[180] br[180] wl[58] vdd gnd cell_6t
Xbit_r59_c180 bl[180] br[180] wl[59] vdd gnd cell_6t
Xbit_r60_c180 bl[180] br[180] wl[60] vdd gnd cell_6t
Xbit_r61_c180 bl[180] br[180] wl[61] vdd gnd cell_6t
Xbit_r62_c180 bl[180] br[180] wl[62] vdd gnd cell_6t
Xbit_r63_c180 bl[180] br[180] wl[63] vdd gnd cell_6t
Xbit_r64_c180 bl[180] br[180] wl[64] vdd gnd cell_6t
Xbit_r65_c180 bl[180] br[180] wl[65] vdd gnd cell_6t
Xbit_r66_c180 bl[180] br[180] wl[66] vdd gnd cell_6t
Xbit_r67_c180 bl[180] br[180] wl[67] vdd gnd cell_6t
Xbit_r68_c180 bl[180] br[180] wl[68] vdd gnd cell_6t
Xbit_r69_c180 bl[180] br[180] wl[69] vdd gnd cell_6t
Xbit_r70_c180 bl[180] br[180] wl[70] vdd gnd cell_6t
Xbit_r71_c180 bl[180] br[180] wl[71] vdd gnd cell_6t
Xbit_r72_c180 bl[180] br[180] wl[72] vdd gnd cell_6t
Xbit_r73_c180 bl[180] br[180] wl[73] vdd gnd cell_6t
Xbit_r74_c180 bl[180] br[180] wl[74] vdd gnd cell_6t
Xbit_r75_c180 bl[180] br[180] wl[75] vdd gnd cell_6t
Xbit_r76_c180 bl[180] br[180] wl[76] vdd gnd cell_6t
Xbit_r77_c180 bl[180] br[180] wl[77] vdd gnd cell_6t
Xbit_r78_c180 bl[180] br[180] wl[78] vdd gnd cell_6t
Xbit_r79_c180 bl[180] br[180] wl[79] vdd gnd cell_6t
Xbit_r80_c180 bl[180] br[180] wl[80] vdd gnd cell_6t
Xbit_r81_c180 bl[180] br[180] wl[81] vdd gnd cell_6t
Xbit_r82_c180 bl[180] br[180] wl[82] vdd gnd cell_6t
Xbit_r83_c180 bl[180] br[180] wl[83] vdd gnd cell_6t
Xbit_r84_c180 bl[180] br[180] wl[84] vdd gnd cell_6t
Xbit_r85_c180 bl[180] br[180] wl[85] vdd gnd cell_6t
Xbit_r86_c180 bl[180] br[180] wl[86] vdd gnd cell_6t
Xbit_r87_c180 bl[180] br[180] wl[87] vdd gnd cell_6t
Xbit_r88_c180 bl[180] br[180] wl[88] vdd gnd cell_6t
Xbit_r89_c180 bl[180] br[180] wl[89] vdd gnd cell_6t
Xbit_r90_c180 bl[180] br[180] wl[90] vdd gnd cell_6t
Xbit_r91_c180 bl[180] br[180] wl[91] vdd gnd cell_6t
Xbit_r92_c180 bl[180] br[180] wl[92] vdd gnd cell_6t
Xbit_r93_c180 bl[180] br[180] wl[93] vdd gnd cell_6t
Xbit_r94_c180 bl[180] br[180] wl[94] vdd gnd cell_6t
Xbit_r95_c180 bl[180] br[180] wl[95] vdd gnd cell_6t
Xbit_r96_c180 bl[180] br[180] wl[96] vdd gnd cell_6t
Xbit_r97_c180 bl[180] br[180] wl[97] vdd gnd cell_6t
Xbit_r98_c180 bl[180] br[180] wl[98] vdd gnd cell_6t
Xbit_r99_c180 bl[180] br[180] wl[99] vdd gnd cell_6t
Xbit_r100_c180 bl[180] br[180] wl[100] vdd gnd cell_6t
Xbit_r101_c180 bl[180] br[180] wl[101] vdd gnd cell_6t
Xbit_r102_c180 bl[180] br[180] wl[102] vdd gnd cell_6t
Xbit_r103_c180 bl[180] br[180] wl[103] vdd gnd cell_6t
Xbit_r104_c180 bl[180] br[180] wl[104] vdd gnd cell_6t
Xbit_r105_c180 bl[180] br[180] wl[105] vdd gnd cell_6t
Xbit_r106_c180 bl[180] br[180] wl[106] vdd gnd cell_6t
Xbit_r107_c180 bl[180] br[180] wl[107] vdd gnd cell_6t
Xbit_r108_c180 bl[180] br[180] wl[108] vdd gnd cell_6t
Xbit_r109_c180 bl[180] br[180] wl[109] vdd gnd cell_6t
Xbit_r110_c180 bl[180] br[180] wl[110] vdd gnd cell_6t
Xbit_r111_c180 bl[180] br[180] wl[111] vdd gnd cell_6t
Xbit_r112_c180 bl[180] br[180] wl[112] vdd gnd cell_6t
Xbit_r113_c180 bl[180] br[180] wl[113] vdd gnd cell_6t
Xbit_r114_c180 bl[180] br[180] wl[114] vdd gnd cell_6t
Xbit_r115_c180 bl[180] br[180] wl[115] vdd gnd cell_6t
Xbit_r116_c180 bl[180] br[180] wl[116] vdd gnd cell_6t
Xbit_r117_c180 bl[180] br[180] wl[117] vdd gnd cell_6t
Xbit_r118_c180 bl[180] br[180] wl[118] vdd gnd cell_6t
Xbit_r119_c180 bl[180] br[180] wl[119] vdd gnd cell_6t
Xbit_r120_c180 bl[180] br[180] wl[120] vdd gnd cell_6t
Xbit_r121_c180 bl[180] br[180] wl[121] vdd gnd cell_6t
Xbit_r122_c180 bl[180] br[180] wl[122] vdd gnd cell_6t
Xbit_r123_c180 bl[180] br[180] wl[123] vdd gnd cell_6t
Xbit_r124_c180 bl[180] br[180] wl[124] vdd gnd cell_6t
Xbit_r125_c180 bl[180] br[180] wl[125] vdd gnd cell_6t
Xbit_r126_c180 bl[180] br[180] wl[126] vdd gnd cell_6t
Xbit_r127_c180 bl[180] br[180] wl[127] vdd gnd cell_6t
Xbit_r0_c181 bl[181] br[181] wl[0] vdd gnd cell_6t
Xbit_r1_c181 bl[181] br[181] wl[1] vdd gnd cell_6t
Xbit_r2_c181 bl[181] br[181] wl[2] vdd gnd cell_6t
Xbit_r3_c181 bl[181] br[181] wl[3] vdd gnd cell_6t
Xbit_r4_c181 bl[181] br[181] wl[4] vdd gnd cell_6t
Xbit_r5_c181 bl[181] br[181] wl[5] vdd gnd cell_6t
Xbit_r6_c181 bl[181] br[181] wl[6] vdd gnd cell_6t
Xbit_r7_c181 bl[181] br[181] wl[7] vdd gnd cell_6t
Xbit_r8_c181 bl[181] br[181] wl[8] vdd gnd cell_6t
Xbit_r9_c181 bl[181] br[181] wl[9] vdd gnd cell_6t
Xbit_r10_c181 bl[181] br[181] wl[10] vdd gnd cell_6t
Xbit_r11_c181 bl[181] br[181] wl[11] vdd gnd cell_6t
Xbit_r12_c181 bl[181] br[181] wl[12] vdd gnd cell_6t
Xbit_r13_c181 bl[181] br[181] wl[13] vdd gnd cell_6t
Xbit_r14_c181 bl[181] br[181] wl[14] vdd gnd cell_6t
Xbit_r15_c181 bl[181] br[181] wl[15] vdd gnd cell_6t
Xbit_r16_c181 bl[181] br[181] wl[16] vdd gnd cell_6t
Xbit_r17_c181 bl[181] br[181] wl[17] vdd gnd cell_6t
Xbit_r18_c181 bl[181] br[181] wl[18] vdd gnd cell_6t
Xbit_r19_c181 bl[181] br[181] wl[19] vdd gnd cell_6t
Xbit_r20_c181 bl[181] br[181] wl[20] vdd gnd cell_6t
Xbit_r21_c181 bl[181] br[181] wl[21] vdd gnd cell_6t
Xbit_r22_c181 bl[181] br[181] wl[22] vdd gnd cell_6t
Xbit_r23_c181 bl[181] br[181] wl[23] vdd gnd cell_6t
Xbit_r24_c181 bl[181] br[181] wl[24] vdd gnd cell_6t
Xbit_r25_c181 bl[181] br[181] wl[25] vdd gnd cell_6t
Xbit_r26_c181 bl[181] br[181] wl[26] vdd gnd cell_6t
Xbit_r27_c181 bl[181] br[181] wl[27] vdd gnd cell_6t
Xbit_r28_c181 bl[181] br[181] wl[28] vdd gnd cell_6t
Xbit_r29_c181 bl[181] br[181] wl[29] vdd gnd cell_6t
Xbit_r30_c181 bl[181] br[181] wl[30] vdd gnd cell_6t
Xbit_r31_c181 bl[181] br[181] wl[31] vdd gnd cell_6t
Xbit_r32_c181 bl[181] br[181] wl[32] vdd gnd cell_6t
Xbit_r33_c181 bl[181] br[181] wl[33] vdd gnd cell_6t
Xbit_r34_c181 bl[181] br[181] wl[34] vdd gnd cell_6t
Xbit_r35_c181 bl[181] br[181] wl[35] vdd gnd cell_6t
Xbit_r36_c181 bl[181] br[181] wl[36] vdd gnd cell_6t
Xbit_r37_c181 bl[181] br[181] wl[37] vdd gnd cell_6t
Xbit_r38_c181 bl[181] br[181] wl[38] vdd gnd cell_6t
Xbit_r39_c181 bl[181] br[181] wl[39] vdd gnd cell_6t
Xbit_r40_c181 bl[181] br[181] wl[40] vdd gnd cell_6t
Xbit_r41_c181 bl[181] br[181] wl[41] vdd gnd cell_6t
Xbit_r42_c181 bl[181] br[181] wl[42] vdd gnd cell_6t
Xbit_r43_c181 bl[181] br[181] wl[43] vdd gnd cell_6t
Xbit_r44_c181 bl[181] br[181] wl[44] vdd gnd cell_6t
Xbit_r45_c181 bl[181] br[181] wl[45] vdd gnd cell_6t
Xbit_r46_c181 bl[181] br[181] wl[46] vdd gnd cell_6t
Xbit_r47_c181 bl[181] br[181] wl[47] vdd gnd cell_6t
Xbit_r48_c181 bl[181] br[181] wl[48] vdd gnd cell_6t
Xbit_r49_c181 bl[181] br[181] wl[49] vdd gnd cell_6t
Xbit_r50_c181 bl[181] br[181] wl[50] vdd gnd cell_6t
Xbit_r51_c181 bl[181] br[181] wl[51] vdd gnd cell_6t
Xbit_r52_c181 bl[181] br[181] wl[52] vdd gnd cell_6t
Xbit_r53_c181 bl[181] br[181] wl[53] vdd gnd cell_6t
Xbit_r54_c181 bl[181] br[181] wl[54] vdd gnd cell_6t
Xbit_r55_c181 bl[181] br[181] wl[55] vdd gnd cell_6t
Xbit_r56_c181 bl[181] br[181] wl[56] vdd gnd cell_6t
Xbit_r57_c181 bl[181] br[181] wl[57] vdd gnd cell_6t
Xbit_r58_c181 bl[181] br[181] wl[58] vdd gnd cell_6t
Xbit_r59_c181 bl[181] br[181] wl[59] vdd gnd cell_6t
Xbit_r60_c181 bl[181] br[181] wl[60] vdd gnd cell_6t
Xbit_r61_c181 bl[181] br[181] wl[61] vdd gnd cell_6t
Xbit_r62_c181 bl[181] br[181] wl[62] vdd gnd cell_6t
Xbit_r63_c181 bl[181] br[181] wl[63] vdd gnd cell_6t
Xbit_r64_c181 bl[181] br[181] wl[64] vdd gnd cell_6t
Xbit_r65_c181 bl[181] br[181] wl[65] vdd gnd cell_6t
Xbit_r66_c181 bl[181] br[181] wl[66] vdd gnd cell_6t
Xbit_r67_c181 bl[181] br[181] wl[67] vdd gnd cell_6t
Xbit_r68_c181 bl[181] br[181] wl[68] vdd gnd cell_6t
Xbit_r69_c181 bl[181] br[181] wl[69] vdd gnd cell_6t
Xbit_r70_c181 bl[181] br[181] wl[70] vdd gnd cell_6t
Xbit_r71_c181 bl[181] br[181] wl[71] vdd gnd cell_6t
Xbit_r72_c181 bl[181] br[181] wl[72] vdd gnd cell_6t
Xbit_r73_c181 bl[181] br[181] wl[73] vdd gnd cell_6t
Xbit_r74_c181 bl[181] br[181] wl[74] vdd gnd cell_6t
Xbit_r75_c181 bl[181] br[181] wl[75] vdd gnd cell_6t
Xbit_r76_c181 bl[181] br[181] wl[76] vdd gnd cell_6t
Xbit_r77_c181 bl[181] br[181] wl[77] vdd gnd cell_6t
Xbit_r78_c181 bl[181] br[181] wl[78] vdd gnd cell_6t
Xbit_r79_c181 bl[181] br[181] wl[79] vdd gnd cell_6t
Xbit_r80_c181 bl[181] br[181] wl[80] vdd gnd cell_6t
Xbit_r81_c181 bl[181] br[181] wl[81] vdd gnd cell_6t
Xbit_r82_c181 bl[181] br[181] wl[82] vdd gnd cell_6t
Xbit_r83_c181 bl[181] br[181] wl[83] vdd gnd cell_6t
Xbit_r84_c181 bl[181] br[181] wl[84] vdd gnd cell_6t
Xbit_r85_c181 bl[181] br[181] wl[85] vdd gnd cell_6t
Xbit_r86_c181 bl[181] br[181] wl[86] vdd gnd cell_6t
Xbit_r87_c181 bl[181] br[181] wl[87] vdd gnd cell_6t
Xbit_r88_c181 bl[181] br[181] wl[88] vdd gnd cell_6t
Xbit_r89_c181 bl[181] br[181] wl[89] vdd gnd cell_6t
Xbit_r90_c181 bl[181] br[181] wl[90] vdd gnd cell_6t
Xbit_r91_c181 bl[181] br[181] wl[91] vdd gnd cell_6t
Xbit_r92_c181 bl[181] br[181] wl[92] vdd gnd cell_6t
Xbit_r93_c181 bl[181] br[181] wl[93] vdd gnd cell_6t
Xbit_r94_c181 bl[181] br[181] wl[94] vdd gnd cell_6t
Xbit_r95_c181 bl[181] br[181] wl[95] vdd gnd cell_6t
Xbit_r96_c181 bl[181] br[181] wl[96] vdd gnd cell_6t
Xbit_r97_c181 bl[181] br[181] wl[97] vdd gnd cell_6t
Xbit_r98_c181 bl[181] br[181] wl[98] vdd gnd cell_6t
Xbit_r99_c181 bl[181] br[181] wl[99] vdd gnd cell_6t
Xbit_r100_c181 bl[181] br[181] wl[100] vdd gnd cell_6t
Xbit_r101_c181 bl[181] br[181] wl[101] vdd gnd cell_6t
Xbit_r102_c181 bl[181] br[181] wl[102] vdd gnd cell_6t
Xbit_r103_c181 bl[181] br[181] wl[103] vdd gnd cell_6t
Xbit_r104_c181 bl[181] br[181] wl[104] vdd gnd cell_6t
Xbit_r105_c181 bl[181] br[181] wl[105] vdd gnd cell_6t
Xbit_r106_c181 bl[181] br[181] wl[106] vdd gnd cell_6t
Xbit_r107_c181 bl[181] br[181] wl[107] vdd gnd cell_6t
Xbit_r108_c181 bl[181] br[181] wl[108] vdd gnd cell_6t
Xbit_r109_c181 bl[181] br[181] wl[109] vdd gnd cell_6t
Xbit_r110_c181 bl[181] br[181] wl[110] vdd gnd cell_6t
Xbit_r111_c181 bl[181] br[181] wl[111] vdd gnd cell_6t
Xbit_r112_c181 bl[181] br[181] wl[112] vdd gnd cell_6t
Xbit_r113_c181 bl[181] br[181] wl[113] vdd gnd cell_6t
Xbit_r114_c181 bl[181] br[181] wl[114] vdd gnd cell_6t
Xbit_r115_c181 bl[181] br[181] wl[115] vdd gnd cell_6t
Xbit_r116_c181 bl[181] br[181] wl[116] vdd gnd cell_6t
Xbit_r117_c181 bl[181] br[181] wl[117] vdd gnd cell_6t
Xbit_r118_c181 bl[181] br[181] wl[118] vdd gnd cell_6t
Xbit_r119_c181 bl[181] br[181] wl[119] vdd gnd cell_6t
Xbit_r120_c181 bl[181] br[181] wl[120] vdd gnd cell_6t
Xbit_r121_c181 bl[181] br[181] wl[121] vdd gnd cell_6t
Xbit_r122_c181 bl[181] br[181] wl[122] vdd gnd cell_6t
Xbit_r123_c181 bl[181] br[181] wl[123] vdd gnd cell_6t
Xbit_r124_c181 bl[181] br[181] wl[124] vdd gnd cell_6t
Xbit_r125_c181 bl[181] br[181] wl[125] vdd gnd cell_6t
Xbit_r126_c181 bl[181] br[181] wl[126] vdd gnd cell_6t
Xbit_r127_c181 bl[181] br[181] wl[127] vdd gnd cell_6t
Xbit_r0_c182 bl[182] br[182] wl[0] vdd gnd cell_6t
Xbit_r1_c182 bl[182] br[182] wl[1] vdd gnd cell_6t
Xbit_r2_c182 bl[182] br[182] wl[2] vdd gnd cell_6t
Xbit_r3_c182 bl[182] br[182] wl[3] vdd gnd cell_6t
Xbit_r4_c182 bl[182] br[182] wl[4] vdd gnd cell_6t
Xbit_r5_c182 bl[182] br[182] wl[5] vdd gnd cell_6t
Xbit_r6_c182 bl[182] br[182] wl[6] vdd gnd cell_6t
Xbit_r7_c182 bl[182] br[182] wl[7] vdd gnd cell_6t
Xbit_r8_c182 bl[182] br[182] wl[8] vdd gnd cell_6t
Xbit_r9_c182 bl[182] br[182] wl[9] vdd gnd cell_6t
Xbit_r10_c182 bl[182] br[182] wl[10] vdd gnd cell_6t
Xbit_r11_c182 bl[182] br[182] wl[11] vdd gnd cell_6t
Xbit_r12_c182 bl[182] br[182] wl[12] vdd gnd cell_6t
Xbit_r13_c182 bl[182] br[182] wl[13] vdd gnd cell_6t
Xbit_r14_c182 bl[182] br[182] wl[14] vdd gnd cell_6t
Xbit_r15_c182 bl[182] br[182] wl[15] vdd gnd cell_6t
Xbit_r16_c182 bl[182] br[182] wl[16] vdd gnd cell_6t
Xbit_r17_c182 bl[182] br[182] wl[17] vdd gnd cell_6t
Xbit_r18_c182 bl[182] br[182] wl[18] vdd gnd cell_6t
Xbit_r19_c182 bl[182] br[182] wl[19] vdd gnd cell_6t
Xbit_r20_c182 bl[182] br[182] wl[20] vdd gnd cell_6t
Xbit_r21_c182 bl[182] br[182] wl[21] vdd gnd cell_6t
Xbit_r22_c182 bl[182] br[182] wl[22] vdd gnd cell_6t
Xbit_r23_c182 bl[182] br[182] wl[23] vdd gnd cell_6t
Xbit_r24_c182 bl[182] br[182] wl[24] vdd gnd cell_6t
Xbit_r25_c182 bl[182] br[182] wl[25] vdd gnd cell_6t
Xbit_r26_c182 bl[182] br[182] wl[26] vdd gnd cell_6t
Xbit_r27_c182 bl[182] br[182] wl[27] vdd gnd cell_6t
Xbit_r28_c182 bl[182] br[182] wl[28] vdd gnd cell_6t
Xbit_r29_c182 bl[182] br[182] wl[29] vdd gnd cell_6t
Xbit_r30_c182 bl[182] br[182] wl[30] vdd gnd cell_6t
Xbit_r31_c182 bl[182] br[182] wl[31] vdd gnd cell_6t
Xbit_r32_c182 bl[182] br[182] wl[32] vdd gnd cell_6t
Xbit_r33_c182 bl[182] br[182] wl[33] vdd gnd cell_6t
Xbit_r34_c182 bl[182] br[182] wl[34] vdd gnd cell_6t
Xbit_r35_c182 bl[182] br[182] wl[35] vdd gnd cell_6t
Xbit_r36_c182 bl[182] br[182] wl[36] vdd gnd cell_6t
Xbit_r37_c182 bl[182] br[182] wl[37] vdd gnd cell_6t
Xbit_r38_c182 bl[182] br[182] wl[38] vdd gnd cell_6t
Xbit_r39_c182 bl[182] br[182] wl[39] vdd gnd cell_6t
Xbit_r40_c182 bl[182] br[182] wl[40] vdd gnd cell_6t
Xbit_r41_c182 bl[182] br[182] wl[41] vdd gnd cell_6t
Xbit_r42_c182 bl[182] br[182] wl[42] vdd gnd cell_6t
Xbit_r43_c182 bl[182] br[182] wl[43] vdd gnd cell_6t
Xbit_r44_c182 bl[182] br[182] wl[44] vdd gnd cell_6t
Xbit_r45_c182 bl[182] br[182] wl[45] vdd gnd cell_6t
Xbit_r46_c182 bl[182] br[182] wl[46] vdd gnd cell_6t
Xbit_r47_c182 bl[182] br[182] wl[47] vdd gnd cell_6t
Xbit_r48_c182 bl[182] br[182] wl[48] vdd gnd cell_6t
Xbit_r49_c182 bl[182] br[182] wl[49] vdd gnd cell_6t
Xbit_r50_c182 bl[182] br[182] wl[50] vdd gnd cell_6t
Xbit_r51_c182 bl[182] br[182] wl[51] vdd gnd cell_6t
Xbit_r52_c182 bl[182] br[182] wl[52] vdd gnd cell_6t
Xbit_r53_c182 bl[182] br[182] wl[53] vdd gnd cell_6t
Xbit_r54_c182 bl[182] br[182] wl[54] vdd gnd cell_6t
Xbit_r55_c182 bl[182] br[182] wl[55] vdd gnd cell_6t
Xbit_r56_c182 bl[182] br[182] wl[56] vdd gnd cell_6t
Xbit_r57_c182 bl[182] br[182] wl[57] vdd gnd cell_6t
Xbit_r58_c182 bl[182] br[182] wl[58] vdd gnd cell_6t
Xbit_r59_c182 bl[182] br[182] wl[59] vdd gnd cell_6t
Xbit_r60_c182 bl[182] br[182] wl[60] vdd gnd cell_6t
Xbit_r61_c182 bl[182] br[182] wl[61] vdd gnd cell_6t
Xbit_r62_c182 bl[182] br[182] wl[62] vdd gnd cell_6t
Xbit_r63_c182 bl[182] br[182] wl[63] vdd gnd cell_6t
Xbit_r64_c182 bl[182] br[182] wl[64] vdd gnd cell_6t
Xbit_r65_c182 bl[182] br[182] wl[65] vdd gnd cell_6t
Xbit_r66_c182 bl[182] br[182] wl[66] vdd gnd cell_6t
Xbit_r67_c182 bl[182] br[182] wl[67] vdd gnd cell_6t
Xbit_r68_c182 bl[182] br[182] wl[68] vdd gnd cell_6t
Xbit_r69_c182 bl[182] br[182] wl[69] vdd gnd cell_6t
Xbit_r70_c182 bl[182] br[182] wl[70] vdd gnd cell_6t
Xbit_r71_c182 bl[182] br[182] wl[71] vdd gnd cell_6t
Xbit_r72_c182 bl[182] br[182] wl[72] vdd gnd cell_6t
Xbit_r73_c182 bl[182] br[182] wl[73] vdd gnd cell_6t
Xbit_r74_c182 bl[182] br[182] wl[74] vdd gnd cell_6t
Xbit_r75_c182 bl[182] br[182] wl[75] vdd gnd cell_6t
Xbit_r76_c182 bl[182] br[182] wl[76] vdd gnd cell_6t
Xbit_r77_c182 bl[182] br[182] wl[77] vdd gnd cell_6t
Xbit_r78_c182 bl[182] br[182] wl[78] vdd gnd cell_6t
Xbit_r79_c182 bl[182] br[182] wl[79] vdd gnd cell_6t
Xbit_r80_c182 bl[182] br[182] wl[80] vdd gnd cell_6t
Xbit_r81_c182 bl[182] br[182] wl[81] vdd gnd cell_6t
Xbit_r82_c182 bl[182] br[182] wl[82] vdd gnd cell_6t
Xbit_r83_c182 bl[182] br[182] wl[83] vdd gnd cell_6t
Xbit_r84_c182 bl[182] br[182] wl[84] vdd gnd cell_6t
Xbit_r85_c182 bl[182] br[182] wl[85] vdd gnd cell_6t
Xbit_r86_c182 bl[182] br[182] wl[86] vdd gnd cell_6t
Xbit_r87_c182 bl[182] br[182] wl[87] vdd gnd cell_6t
Xbit_r88_c182 bl[182] br[182] wl[88] vdd gnd cell_6t
Xbit_r89_c182 bl[182] br[182] wl[89] vdd gnd cell_6t
Xbit_r90_c182 bl[182] br[182] wl[90] vdd gnd cell_6t
Xbit_r91_c182 bl[182] br[182] wl[91] vdd gnd cell_6t
Xbit_r92_c182 bl[182] br[182] wl[92] vdd gnd cell_6t
Xbit_r93_c182 bl[182] br[182] wl[93] vdd gnd cell_6t
Xbit_r94_c182 bl[182] br[182] wl[94] vdd gnd cell_6t
Xbit_r95_c182 bl[182] br[182] wl[95] vdd gnd cell_6t
Xbit_r96_c182 bl[182] br[182] wl[96] vdd gnd cell_6t
Xbit_r97_c182 bl[182] br[182] wl[97] vdd gnd cell_6t
Xbit_r98_c182 bl[182] br[182] wl[98] vdd gnd cell_6t
Xbit_r99_c182 bl[182] br[182] wl[99] vdd gnd cell_6t
Xbit_r100_c182 bl[182] br[182] wl[100] vdd gnd cell_6t
Xbit_r101_c182 bl[182] br[182] wl[101] vdd gnd cell_6t
Xbit_r102_c182 bl[182] br[182] wl[102] vdd gnd cell_6t
Xbit_r103_c182 bl[182] br[182] wl[103] vdd gnd cell_6t
Xbit_r104_c182 bl[182] br[182] wl[104] vdd gnd cell_6t
Xbit_r105_c182 bl[182] br[182] wl[105] vdd gnd cell_6t
Xbit_r106_c182 bl[182] br[182] wl[106] vdd gnd cell_6t
Xbit_r107_c182 bl[182] br[182] wl[107] vdd gnd cell_6t
Xbit_r108_c182 bl[182] br[182] wl[108] vdd gnd cell_6t
Xbit_r109_c182 bl[182] br[182] wl[109] vdd gnd cell_6t
Xbit_r110_c182 bl[182] br[182] wl[110] vdd gnd cell_6t
Xbit_r111_c182 bl[182] br[182] wl[111] vdd gnd cell_6t
Xbit_r112_c182 bl[182] br[182] wl[112] vdd gnd cell_6t
Xbit_r113_c182 bl[182] br[182] wl[113] vdd gnd cell_6t
Xbit_r114_c182 bl[182] br[182] wl[114] vdd gnd cell_6t
Xbit_r115_c182 bl[182] br[182] wl[115] vdd gnd cell_6t
Xbit_r116_c182 bl[182] br[182] wl[116] vdd gnd cell_6t
Xbit_r117_c182 bl[182] br[182] wl[117] vdd gnd cell_6t
Xbit_r118_c182 bl[182] br[182] wl[118] vdd gnd cell_6t
Xbit_r119_c182 bl[182] br[182] wl[119] vdd gnd cell_6t
Xbit_r120_c182 bl[182] br[182] wl[120] vdd gnd cell_6t
Xbit_r121_c182 bl[182] br[182] wl[121] vdd gnd cell_6t
Xbit_r122_c182 bl[182] br[182] wl[122] vdd gnd cell_6t
Xbit_r123_c182 bl[182] br[182] wl[123] vdd gnd cell_6t
Xbit_r124_c182 bl[182] br[182] wl[124] vdd gnd cell_6t
Xbit_r125_c182 bl[182] br[182] wl[125] vdd gnd cell_6t
Xbit_r126_c182 bl[182] br[182] wl[126] vdd gnd cell_6t
Xbit_r127_c182 bl[182] br[182] wl[127] vdd gnd cell_6t
Xbit_r0_c183 bl[183] br[183] wl[0] vdd gnd cell_6t
Xbit_r1_c183 bl[183] br[183] wl[1] vdd gnd cell_6t
Xbit_r2_c183 bl[183] br[183] wl[2] vdd gnd cell_6t
Xbit_r3_c183 bl[183] br[183] wl[3] vdd gnd cell_6t
Xbit_r4_c183 bl[183] br[183] wl[4] vdd gnd cell_6t
Xbit_r5_c183 bl[183] br[183] wl[5] vdd gnd cell_6t
Xbit_r6_c183 bl[183] br[183] wl[6] vdd gnd cell_6t
Xbit_r7_c183 bl[183] br[183] wl[7] vdd gnd cell_6t
Xbit_r8_c183 bl[183] br[183] wl[8] vdd gnd cell_6t
Xbit_r9_c183 bl[183] br[183] wl[9] vdd gnd cell_6t
Xbit_r10_c183 bl[183] br[183] wl[10] vdd gnd cell_6t
Xbit_r11_c183 bl[183] br[183] wl[11] vdd gnd cell_6t
Xbit_r12_c183 bl[183] br[183] wl[12] vdd gnd cell_6t
Xbit_r13_c183 bl[183] br[183] wl[13] vdd gnd cell_6t
Xbit_r14_c183 bl[183] br[183] wl[14] vdd gnd cell_6t
Xbit_r15_c183 bl[183] br[183] wl[15] vdd gnd cell_6t
Xbit_r16_c183 bl[183] br[183] wl[16] vdd gnd cell_6t
Xbit_r17_c183 bl[183] br[183] wl[17] vdd gnd cell_6t
Xbit_r18_c183 bl[183] br[183] wl[18] vdd gnd cell_6t
Xbit_r19_c183 bl[183] br[183] wl[19] vdd gnd cell_6t
Xbit_r20_c183 bl[183] br[183] wl[20] vdd gnd cell_6t
Xbit_r21_c183 bl[183] br[183] wl[21] vdd gnd cell_6t
Xbit_r22_c183 bl[183] br[183] wl[22] vdd gnd cell_6t
Xbit_r23_c183 bl[183] br[183] wl[23] vdd gnd cell_6t
Xbit_r24_c183 bl[183] br[183] wl[24] vdd gnd cell_6t
Xbit_r25_c183 bl[183] br[183] wl[25] vdd gnd cell_6t
Xbit_r26_c183 bl[183] br[183] wl[26] vdd gnd cell_6t
Xbit_r27_c183 bl[183] br[183] wl[27] vdd gnd cell_6t
Xbit_r28_c183 bl[183] br[183] wl[28] vdd gnd cell_6t
Xbit_r29_c183 bl[183] br[183] wl[29] vdd gnd cell_6t
Xbit_r30_c183 bl[183] br[183] wl[30] vdd gnd cell_6t
Xbit_r31_c183 bl[183] br[183] wl[31] vdd gnd cell_6t
Xbit_r32_c183 bl[183] br[183] wl[32] vdd gnd cell_6t
Xbit_r33_c183 bl[183] br[183] wl[33] vdd gnd cell_6t
Xbit_r34_c183 bl[183] br[183] wl[34] vdd gnd cell_6t
Xbit_r35_c183 bl[183] br[183] wl[35] vdd gnd cell_6t
Xbit_r36_c183 bl[183] br[183] wl[36] vdd gnd cell_6t
Xbit_r37_c183 bl[183] br[183] wl[37] vdd gnd cell_6t
Xbit_r38_c183 bl[183] br[183] wl[38] vdd gnd cell_6t
Xbit_r39_c183 bl[183] br[183] wl[39] vdd gnd cell_6t
Xbit_r40_c183 bl[183] br[183] wl[40] vdd gnd cell_6t
Xbit_r41_c183 bl[183] br[183] wl[41] vdd gnd cell_6t
Xbit_r42_c183 bl[183] br[183] wl[42] vdd gnd cell_6t
Xbit_r43_c183 bl[183] br[183] wl[43] vdd gnd cell_6t
Xbit_r44_c183 bl[183] br[183] wl[44] vdd gnd cell_6t
Xbit_r45_c183 bl[183] br[183] wl[45] vdd gnd cell_6t
Xbit_r46_c183 bl[183] br[183] wl[46] vdd gnd cell_6t
Xbit_r47_c183 bl[183] br[183] wl[47] vdd gnd cell_6t
Xbit_r48_c183 bl[183] br[183] wl[48] vdd gnd cell_6t
Xbit_r49_c183 bl[183] br[183] wl[49] vdd gnd cell_6t
Xbit_r50_c183 bl[183] br[183] wl[50] vdd gnd cell_6t
Xbit_r51_c183 bl[183] br[183] wl[51] vdd gnd cell_6t
Xbit_r52_c183 bl[183] br[183] wl[52] vdd gnd cell_6t
Xbit_r53_c183 bl[183] br[183] wl[53] vdd gnd cell_6t
Xbit_r54_c183 bl[183] br[183] wl[54] vdd gnd cell_6t
Xbit_r55_c183 bl[183] br[183] wl[55] vdd gnd cell_6t
Xbit_r56_c183 bl[183] br[183] wl[56] vdd gnd cell_6t
Xbit_r57_c183 bl[183] br[183] wl[57] vdd gnd cell_6t
Xbit_r58_c183 bl[183] br[183] wl[58] vdd gnd cell_6t
Xbit_r59_c183 bl[183] br[183] wl[59] vdd gnd cell_6t
Xbit_r60_c183 bl[183] br[183] wl[60] vdd gnd cell_6t
Xbit_r61_c183 bl[183] br[183] wl[61] vdd gnd cell_6t
Xbit_r62_c183 bl[183] br[183] wl[62] vdd gnd cell_6t
Xbit_r63_c183 bl[183] br[183] wl[63] vdd gnd cell_6t
Xbit_r64_c183 bl[183] br[183] wl[64] vdd gnd cell_6t
Xbit_r65_c183 bl[183] br[183] wl[65] vdd gnd cell_6t
Xbit_r66_c183 bl[183] br[183] wl[66] vdd gnd cell_6t
Xbit_r67_c183 bl[183] br[183] wl[67] vdd gnd cell_6t
Xbit_r68_c183 bl[183] br[183] wl[68] vdd gnd cell_6t
Xbit_r69_c183 bl[183] br[183] wl[69] vdd gnd cell_6t
Xbit_r70_c183 bl[183] br[183] wl[70] vdd gnd cell_6t
Xbit_r71_c183 bl[183] br[183] wl[71] vdd gnd cell_6t
Xbit_r72_c183 bl[183] br[183] wl[72] vdd gnd cell_6t
Xbit_r73_c183 bl[183] br[183] wl[73] vdd gnd cell_6t
Xbit_r74_c183 bl[183] br[183] wl[74] vdd gnd cell_6t
Xbit_r75_c183 bl[183] br[183] wl[75] vdd gnd cell_6t
Xbit_r76_c183 bl[183] br[183] wl[76] vdd gnd cell_6t
Xbit_r77_c183 bl[183] br[183] wl[77] vdd gnd cell_6t
Xbit_r78_c183 bl[183] br[183] wl[78] vdd gnd cell_6t
Xbit_r79_c183 bl[183] br[183] wl[79] vdd gnd cell_6t
Xbit_r80_c183 bl[183] br[183] wl[80] vdd gnd cell_6t
Xbit_r81_c183 bl[183] br[183] wl[81] vdd gnd cell_6t
Xbit_r82_c183 bl[183] br[183] wl[82] vdd gnd cell_6t
Xbit_r83_c183 bl[183] br[183] wl[83] vdd gnd cell_6t
Xbit_r84_c183 bl[183] br[183] wl[84] vdd gnd cell_6t
Xbit_r85_c183 bl[183] br[183] wl[85] vdd gnd cell_6t
Xbit_r86_c183 bl[183] br[183] wl[86] vdd gnd cell_6t
Xbit_r87_c183 bl[183] br[183] wl[87] vdd gnd cell_6t
Xbit_r88_c183 bl[183] br[183] wl[88] vdd gnd cell_6t
Xbit_r89_c183 bl[183] br[183] wl[89] vdd gnd cell_6t
Xbit_r90_c183 bl[183] br[183] wl[90] vdd gnd cell_6t
Xbit_r91_c183 bl[183] br[183] wl[91] vdd gnd cell_6t
Xbit_r92_c183 bl[183] br[183] wl[92] vdd gnd cell_6t
Xbit_r93_c183 bl[183] br[183] wl[93] vdd gnd cell_6t
Xbit_r94_c183 bl[183] br[183] wl[94] vdd gnd cell_6t
Xbit_r95_c183 bl[183] br[183] wl[95] vdd gnd cell_6t
Xbit_r96_c183 bl[183] br[183] wl[96] vdd gnd cell_6t
Xbit_r97_c183 bl[183] br[183] wl[97] vdd gnd cell_6t
Xbit_r98_c183 bl[183] br[183] wl[98] vdd gnd cell_6t
Xbit_r99_c183 bl[183] br[183] wl[99] vdd gnd cell_6t
Xbit_r100_c183 bl[183] br[183] wl[100] vdd gnd cell_6t
Xbit_r101_c183 bl[183] br[183] wl[101] vdd gnd cell_6t
Xbit_r102_c183 bl[183] br[183] wl[102] vdd gnd cell_6t
Xbit_r103_c183 bl[183] br[183] wl[103] vdd gnd cell_6t
Xbit_r104_c183 bl[183] br[183] wl[104] vdd gnd cell_6t
Xbit_r105_c183 bl[183] br[183] wl[105] vdd gnd cell_6t
Xbit_r106_c183 bl[183] br[183] wl[106] vdd gnd cell_6t
Xbit_r107_c183 bl[183] br[183] wl[107] vdd gnd cell_6t
Xbit_r108_c183 bl[183] br[183] wl[108] vdd gnd cell_6t
Xbit_r109_c183 bl[183] br[183] wl[109] vdd gnd cell_6t
Xbit_r110_c183 bl[183] br[183] wl[110] vdd gnd cell_6t
Xbit_r111_c183 bl[183] br[183] wl[111] vdd gnd cell_6t
Xbit_r112_c183 bl[183] br[183] wl[112] vdd gnd cell_6t
Xbit_r113_c183 bl[183] br[183] wl[113] vdd gnd cell_6t
Xbit_r114_c183 bl[183] br[183] wl[114] vdd gnd cell_6t
Xbit_r115_c183 bl[183] br[183] wl[115] vdd gnd cell_6t
Xbit_r116_c183 bl[183] br[183] wl[116] vdd gnd cell_6t
Xbit_r117_c183 bl[183] br[183] wl[117] vdd gnd cell_6t
Xbit_r118_c183 bl[183] br[183] wl[118] vdd gnd cell_6t
Xbit_r119_c183 bl[183] br[183] wl[119] vdd gnd cell_6t
Xbit_r120_c183 bl[183] br[183] wl[120] vdd gnd cell_6t
Xbit_r121_c183 bl[183] br[183] wl[121] vdd gnd cell_6t
Xbit_r122_c183 bl[183] br[183] wl[122] vdd gnd cell_6t
Xbit_r123_c183 bl[183] br[183] wl[123] vdd gnd cell_6t
Xbit_r124_c183 bl[183] br[183] wl[124] vdd gnd cell_6t
Xbit_r125_c183 bl[183] br[183] wl[125] vdd gnd cell_6t
Xbit_r126_c183 bl[183] br[183] wl[126] vdd gnd cell_6t
Xbit_r127_c183 bl[183] br[183] wl[127] vdd gnd cell_6t
Xbit_r0_c184 bl[184] br[184] wl[0] vdd gnd cell_6t
Xbit_r1_c184 bl[184] br[184] wl[1] vdd gnd cell_6t
Xbit_r2_c184 bl[184] br[184] wl[2] vdd gnd cell_6t
Xbit_r3_c184 bl[184] br[184] wl[3] vdd gnd cell_6t
Xbit_r4_c184 bl[184] br[184] wl[4] vdd gnd cell_6t
Xbit_r5_c184 bl[184] br[184] wl[5] vdd gnd cell_6t
Xbit_r6_c184 bl[184] br[184] wl[6] vdd gnd cell_6t
Xbit_r7_c184 bl[184] br[184] wl[7] vdd gnd cell_6t
Xbit_r8_c184 bl[184] br[184] wl[8] vdd gnd cell_6t
Xbit_r9_c184 bl[184] br[184] wl[9] vdd gnd cell_6t
Xbit_r10_c184 bl[184] br[184] wl[10] vdd gnd cell_6t
Xbit_r11_c184 bl[184] br[184] wl[11] vdd gnd cell_6t
Xbit_r12_c184 bl[184] br[184] wl[12] vdd gnd cell_6t
Xbit_r13_c184 bl[184] br[184] wl[13] vdd gnd cell_6t
Xbit_r14_c184 bl[184] br[184] wl[14] vdd gnd cell_6t
Xbit_r15_c184 bl[184] br[184] wl[15] vdd gnd cell_6t
Xbit_r16_c184 bl[184] br[184] wl[16] vdd gnd cell_6t
Xbit_r17_c184 bl[184] br[184] wl[17] vdd gnd cell_6t
Xbit_r18_c184 bl[184] br[184] wl[18] vdd gnd cell_6t
Xbit_r19_c184 bl[184] br[184] wl[19] vdd gnd cell_6t
Xbit_r20_c184 bl[184] br[184] wl[20] vdd gnd cell_6t
Xbit_r21_c184 bl[184] br[184] wl[21] vdd gnd cell_6t
Xbit_r22_c184 bl[184] br[184] wl[22] vdd gnd cell_6t
Xbit_r23_c184 bl[184] br[184] wl[23] vdd gnd cell_6t
Xbit_r24_c184 bl[184] br[184] wl[24] vdd gnd cell_6t
Xbit_r25_c184 bl[184] br[184] wl[25] vdd gnd cell_6t
Xbit_r26_c184 bl[184] br[184] wl[26] vdd gnd cell_6t
Xbit_r27_c184 bl[184] br[184] wl[27] vdd gnd cell_6t
Xbit_r28_c184 bl[184] br[184] wl[28] vdd gnd cell_6t
Xbit_r29_c184 bl[184] br[184] wl[29] vdd gnd cell_6t
Xbit_r30_c184 bl[184] br[184] wl[30] vdd gnd cell_6t
Xbit_r31_c184 bl[184] br[184] wl[31] vdd gnd cell_6t
Xbit_r32_c184 bl[184] br[184] wl[32] vdd gnd cell_6t
Xbit_r33_c184 bl[184] br[184] wl[33] vdd gnd cell_6t
Xbit_r34_c184 bl[184] br[184] wl[34] vdd gnd cell_6t
Xbit_r35_c184 bl[184] br[184] wl[35] vdd gnd cell_6t
Xbit_r36_c184 bl[184] br[184] wl[36] vdd gnd cell_6t
Xbit_r37_c184 bl[184] br[184] wl[37] vdd gnd cell_6t
Xbit_r38_c184 bl[184] br[184] wl[38] vdd gnd cell_6t
Xbit_r39_c184 bl[184] br[184] wl[39] vdd gnd cell_6t
Xbit_r40_c184 bl[184] br[184] wl[40] vdd gnd cell_6t
Xbit_r41_c184 bl[184] br[184] wl[41] vdd gnd cell_6t
Xbit_r42_c184 bl[184] br[184] wl[42] vdd gnd cell_6t
Xbit_r43_c184 bl[184] br[184] wl[43] vdd gnd cell_6t
Xbit_r44_c184 bl[184] br[184] wl[44] vdd gnd cell_6t
Xbit_r45_c184 bl[184] br[184] wl[45] vdd gnd cell_6t
Xbit_r46_c184 bl[184] br[184] wl[46] vdd gnd cell_6t
Xbit_r47_c184 bl[184] br[184] wl[47] vdd gnd cell_6t
Xbit_r48_c184 bl[184] br[184] wl[48] vdd gnd cell_6t
Xbit_r49_c184 bl[184] br[184] wl[49] vdd gnd cell_6t
Xbit_r50_c184 bl[184] br[184] wl[50] vdd gnd cell_6t
Xbit_r51_c184 bl[184] br[184] wl[51] vdd gnd cell_6t
Xbit_r52_c184 bl[184] br[184] wl[52] vdd gnd cell_6t
Xbit_r53_c184 bl[184] br[184] wl[53] vdd gnd cell_6t
Xbit_r54_c184 bl[184] br[184] wl[54] vdd gnd cell_6t
Xbit_r55_c184 bl[184] br[184] wl[55] vdd gnd cell_6t
Xbit_r56_c184 bl[184] br[184] wl[56] vdd gnd cell_6t
Xbit_r57_c184 bl[184] br[184] wl[57] vdd gnd cell_6t
Xbit_r58_c184 bl[184] br[184] wl[58] vdd gnd cell_6t
Xbit_r59_c184 bl[184] br[184] wl[59] vdd gnd cell_6t
Xbit_r60_c184 bl[184] br[184] wl[60] vdd gnd cell_6t
Xbit_r61_c184 bl[184] br[184] wl[61] vdd gnd cell_6t
Xbit_r62_c184 bl[184] br[184] wl[62] vdd gnd cell_6t
Xbit_r63_c184 bl[184] br[184] wl[63] vdd gnd cell_6t
Xbit_r64_c184 bl[184] br[184] wl[64] vdd gnd cell_6t
Xbit_r65_c184 bl[184] br[184] wl[65] vdd gnd cell_6t
Xbit_r66_c184 bl[184] br[184] wl[66] vdd gnd cell_6t
Xbit_r67_c184 bl[184] br[184] wl[67] vdd gnd cell_6t
Xbit_r68_c184 bl[184] br[184] wl[68] vdd gnd cell_6t
Xbit_r69_c184 bl[184] br[184] wl[69] vdd gnd cell_6t
Xbit_r70_c184 bl[184] br[184] wl[70] vdd gnd cell_6t
Xbit_r71_c184 bl[184] br[184] wl[71] vdd gnd cell_6t
Xbit_r72_c184 bl[184] br[184] wl[72] vdd gnd cell_6t
Xbit_r73_c184 bl[184] br[184] wl[73] vdd gnd cell_6t
Xbit_r74_c184 bl[184] br[184] wl[74] vdd gnd cell_6t
Xbit_r75_c184 bl[184] br[184] wl[75] vdd gnd cell_6t
Xbit_r76_c184 bl[184] br[184] wl[76] vdd gnd cell_6t
Xbit_r77_c184 bl[184] br[184] wl[77] vdd gnd cell_6t
Xbit_r78_c184 bl[184] br[184] wl[78] vdd gnd cell_6t
Xbit_r79_c184 bl[184] br[184] wl[79] vdd gnd cell_6t
Xbit_r80_c184 bl[184] br[184] wl[80] vdd gnd cell_6t
Xbit_r81_c184 bl[184] br[184] wl[81] vdd gnd cell_6t
Xbit_r82_c184 bl[184] br[184] wl[82] vdd gnd cell_6t
Xbit_r83_c184 bl[184] br[184] wl[83] vdd gnd cell_6t
Xbit_r84_c184 bl[184] br[184] wl[84] vdd gnd cell_6t
Xbit_r85_c184 bl[184] br[184] wl[85] vdd gnd cell_6t
Xbit_r86_c184 bl[184] br[184] wl[86] vdd gnd cell_6t
Xbit_r87_c184 bl[184] br[184] wl[87] vdd gnd cell_6t
Xbit_r88_c184 bl[184] br[184] wl[88] vdd gnd cell_6t
Xbit_r89_c184 bl[184] br[184] wl[89] vdd gnd cell_6t
Xbit_r90_c184 bl[184] br[184] wl[90] vdd gnd cell_6t
Xbit_r91_c184 bl[184] br[184] wl[91] vdd gnd cell_6t
Xbit_r92_c184 bl[184] br[184] wl[92] vdd gnd cell_6t
Xbit_r93_c184 bl[184] br[184] wl[93] vdd gnd cell_6t
Xbit_r94_c184 bl[184] br[184] wl[94] vdd gnd cell_6t
Xbit_r95_c184 bl[184] br[184] wl[95] vdd gnd cell_6t
Xbit_r96_c184 bl[184] br[184] wl[96] vdd gnd cell_6t
Xbit_r97_c184 bl[184] br[184] wl[97] vdd gnd cell_6t
Xbit_r98_c184 bl[184] br[184] wl[98] vdd gnd cell_6t
Xbit_r99_c184 bl[184] br[184] wl[99] vdd gnd cell_6t
Xbit_r100_c184 bl[184] br[184] wl[100] vdd gnd cell_6t
Xbit_r101_c184 bl[184] br[184] wl[101] vdd gnd cell_6t
Xbit_r102_c184 bl[184] br[184] wl[102] vdd gnd cell_6t
Xbit_r103_c184 bl[184] br[184] wl[103] vdd gnd cell_6t
Xbit_r104_c184 bl[184] br[184] wl[104] vdd gnd cell_6t
Xbit_r105_c184 bl[184] br[184] wl[105] vdd gnd cell_6t
Xbit_r106_c184 bl[184] br[184] wl[106] vdd gnd cell_6t
Xbit_r107_c184 bl[184] br[184] wl[107] vdd gnd cell_6t
Xbit_r108_c184 bl[184] br[184] wl[108] vdd gnd cell_6t
Xbit_r109_c184 bl[184] br[184] wl[109] vdd gnd cell_6t
Xbit_r110_c184 bl[184] br[184] wl[110] vdd gnd cell_6t
Xbit_r111_c184 bl[184] br[184] wl[111] vdd gnd cell_6t
Xbit_r112_c184 bl[184] br[184] wl[112] vdd gnd cell_6t
Xbit_r113_c184 bl[184] br[184] wl[113] vdd gnd cell_6t
Xbit_r114_c184 bl[184] br[184] wl[114] vdd gnd cell_6t
Xbit_r115_c184 bl[184] br[184] wl[115] vdd gnd cell_6t
Xbit_r116_c184 bl[184] br[184] wl[116] vdd gnd cell_6t
Xbit_r117_c184 bl[184] br[184] wl[117] vdd gnd cell_6t
Xbit_r118_c184 bl[184] br[184] wl[118] vdd gnd cell_6t
Xbit_r119_c184 bl[184] br[184] wl[119] vdd gnd cell_6t
Xbit_r120_c184 bl[184] br[184] wl[120] vdd gnd cell_6t
Xbit_r121_c184 bl[184] br[184] wl[121] vdd gnd cell_6t
Xbit_r122_c184 bl[184] br[184] wl[122] vdd gnd cell_6t
Xbit_r123_c184 bl[184] br[184] wl[123] vdd gnd cell_6t
Xbit_r124_c184 bl[184] br[184] wl[124] vdd gnd cell_6t
Xbit_r125_c184 bl[184] br[184] wl[125] vdd gnd cell_6t
Xbit_r126_c184 bl[184] br[184] wl[126] vdd gnd cell_6t
Xbit_r127_c184 bl[184] br[184] wl[127] vdd gnd cell_6t
Xbit_r0_c185 bl[185] br[185] wl[0] vdd gnd cell_6t
Xbit_r1_c185 bl[185] br[185] wl[1] vdd gnd cell_6t
Xbit_r2_c185 bl[185] br[185] wl[2] vdd gnd cell_6t
Xbit_r3_c185 bl[185] br[185] wl[3] vdd gnd cell_6t
Xbit_r4_c185 bl[185] br[185] wl[4] vdd gnd cell_6t
Xbit_r5_c185 bl[185] br[185] wl[5] vdd gnd cell_6t
Xbit_r6_c185 bl[185] br[185] wl[6] vdd gnd cell_6t
Xbit_r7_c185 bl[185] br[185] wl[7] vdd gnd cell_6t
Xbit_r8_c185 bl[185] br[185] wl[8] vdd gnd cell_6t
Xbit_r9_c185 bl[185] br[185] wl[9] vdd gnd cell_6t
Xbit_r10_c185 bl[185] br[185] wl[10] vdd gnd cell_6t
Xbit_r11_c185 bl[185] br[185] wl[11] vdd gnd cell_6t
Xbit_r12_c185 bl[185] br[185] wl[12] vdd gnd cell_6t
Xbit_r13_c185 bl[185] br[185] wl[13] vdd gnd cell_6t
Xbit_r14_c185 bl[185] br[185] wl[14] vdd gnd cell_6t
Xbit_r15_c185 bl[185] br[185] wl[15] vdd gnd cell_6t
Xbit_r16_c185 bl[185] br[185] wl[16] vdd gnd cell_6t
Xbit_r17_c185 bl[185] br[185] wl[17] vdd gnd cell_6t
Xbit_r18_c185 bl[185] br[185] wl[18] vdd gnd cell_6t
Xbit_r19_c185 bl[185] br[185] wl[19] vdd gnd cell_6t
Xbit_r20_c185 bl[185] br[185] wl[20] vdd gnd cell_6t
Xbit_r21_c185 bl[185] br[185] wl[21] vdd gnd cell_6t
Xbit_r22_c185 bl[185] br[185] wl[22] vdd gnd cell_6t
Xbit_r23_c185 bl[185] br[185] wl[23] vdd gnd cell_6t
Xbit_r24_c185 bl[185] br[185] wl[24] vdd gnd cell_6t
Xbit_r25_c185 bl[185] br[185] wl[25] vdd gnd cell_6t
Xbit_r26_c185 bl[185] br[185] wl[26] vdd gnd cell_6t
Xbit_r27_c185 bl[185] br[185] wl[27] vdd gnd cell_6t
Xbit_r28_c185 bl[185] br[185] wl[28] vdd gnd cell_6t
Xbit_r29_c185 bl[185] br[185] wl[29] vdd gnd cell_6t
Xbit_r30_c185 bl[185] br[185] wl[30] vdd gnd cell_6t
Xbit_r31_c185 bl[185] br[185] wl[31] vdd gnd cell_6t
Xbit_r32_c185 bl[185] br[185] wl[32] vdd gnd cell_6t
Xbit_r33_c185 bl[185] br[185] wl[33] vdd gnd cell_6t
Xbit_r34_c185 bl[185] br[185] wl[34] vdd gnd cell_6t
Xbit_r35_c185 bl[185] br[185] wl[35] vdd gnd cell_6t
Xbit_r36_c185 bl[185] br[185] wl[36] vdd gnd cell_6t
Xbit_r37_c185 bl[185] br[185] wl[37] vdd gnd cell_6t
Xbit_r38_c185 bl[185] br[185] wl[38] vdd gnd cell_6t
Xbit_r39_c185 bl[185] br[185] wl[39] vdd gnd cell_6t
Xbit_r40_c185 bl[185] br[185] wl[40] vdd gnd cell_6t
Xbit_r41_c185 bl[185] br[185] wl[41] vdd gnd cell_6t
Xbit_r42_c185 bl[185] br[185] wl[42] vdd gnd cell_6t
Xbit_r43_c185 bl[185] br[185] wl[43] vdd gnd cell_6t
Xbit_r44_c185 bl[185] br[185] wl[44] vdd gnd cell_6t
Xbit_r45_c185 bl[185] br[185] wl[45] vdd gnd cell_6t
Xbit_r46_c185 bl[185] br[185] wl[46] vdd gnd cell_6t
Xbit_r47_c185 bl[185] br[185] wl[47] vdd gnd cell_6t
Xbit_r48_c185 bl[185] br[185] wl[48] vdd gnd cell_6t
Xbit_r49_c185 bl[185] br[185] wl[49] vdd gnd cell_6t
Xbit_r50_c185 bl[185] br[185] wl[50] vdd gnd cell_6t
Xbit_r51_c185 bl[185] br[185] wl[51] vdd gnd cell_6t
Xbit_r52_c185 bl[185] br[185] wl[52] vdd gnd cell_6t
Xbit_r53_c185 bl[185] br[185] wl[53] vdd gnd cell_6t
Xbit_r54_c185 bl[185] br[185] wl[54] vdd gnd cell_6t
Xbit_r55_c185 bl[185] br[185] wl[55] vdd gnd cell_6t
Xbit_r56_c185 bl[185] br[185] wl[56] vdd gnd cell_6t
Xbit_r57_c185 bl[185] br[185] wl[57] vdd gnd cell_6t
Xbit_r58_c185 bl[185] br[185] wl[58] vdd gnd cell_6t
Xbit_r59_c185 bl[185] br[185] wl[59] vdd gnd cell_6t
Xbit_r60_c185 bl[185] br[185] wl[60] vdd gnd cell_6t
Xbit_r61_c185 bl[185] br[185] wl[61] vdd gnd cell_6t
Xbit_r62_c185 bl[185] br[185] wl[62] vdd gnd cell_6t
Xbit_r63_c185 bl[185] br[185] wl[63] vdd gnd cell_6t
Xbit_r64_c185 bl[185] br[185] wl[64] vdd gnd cell_6t
Xbit_r65_c185 bl[185] br[185] wl[65] vdd gnd cell_6t
Xbit_r66_c185 bl[185] br[185] wl[66] vdd gnd cell_6t
Xbit_r67_c185 bl[185] br[185] wl[67] vdd gnd cell_6t
Xbit_r68_c185 bl[185] br[185] wl[68] vdd gnd cell_6t
Xbit_r69_c185 bl[185] br[185] wl[69] vdd gnd cell_6t
Xbit_r70_c185 bl[185] br[185] wl[70] vdd gnd cell_6t
Xbit_r71_c185 bl[185] br[185] wl[71] vdd gnd cell_6t
Xbit_r72_c185 bl[185] br[185] wl[72] vdd gnd cell_6t
Xbit_r73_c185 bl[185] br[185] wl[73] vdd gnd cell_6t
Xbit_r74_c185 bl[185] br[185] wl[74] vdd gnd cell_6t
Xbit_r75_c185 bl[185] br[185] wl[75] vdd gnd cell_6t
Xbit_r76_c185 bl[185] br[185] wl[76] vdd gnd cell_6t
Xbit_r77_c185 bl[185] br[185] wl[77] vdd gnd cell_6t
Xbit_r78_c185 bl[185] br[185] wl[78] vdd gnd cell_6t
Xbit_r79_c185 bl[185] br[185] wl[79] vdd gnd cell_6t
Xbit_r80_c185 bl[185] br[185] wl[80] vdd gnd cell_6t
Xbit_r81_c185 bl[185] br[185] wl[81] vdd gnd cell_6t
Xbit_r82_c185 bl[185] br[185] wl[82] vdd gnd cell_6t
Xbit_r83_c185 bl[185] br[185] wl[83] vdd gnd cell_6t
Xbit_r84_c185 bl[185] br[185] wl[84] vdd gnd cell_6t
Xbit_r85_c185 bl[185] br[185] wl[85] vdd gnd cell_6t
Xbit_r86_c185 bl[185] br[185] wl[86] vdd gnd cell_6t
Xbit_r87_c185 bl[185] br[185] wl[87] vdd gnd cell_6t
Xbit_r88_c185 bl[185] br[185] wl[88] vdd gnd cell_6t
Xbit_r89_c185 bl[185] br[185] wl[89] vdd gnd cell_6t
Xbit_r90_c185 bl[185] br[185] wl[90] vdd gnd cell_6t
Xbit_r91_c185 bl[185] br[185] wl[91] vdd gnd cell_6t
Xbit_r92_c185 bl[185] br[185] wl[92] vdd gnd cell_6t
Xbit_r93_c185 bl[185] br[185] wl[93] vdd gnd cell_6t
Xbit_r94_c185 bl[185] br[185] wl[94] vdd gnd cell_6t
Xbit_r95_c185 bl[185] br[185] wl[95] vdd gnd cell_6t
Xbit_r96_c185 bl[185] br[185] wl[96] vdd gnd cell_6t
Xbit_r97_c185 bl[185] br[185] wl[97] vdd gnd cell_6t
Xbit_r98_c185 bl[185] br[185] wl[98] vdd gnd cell_6t
Xbit_r99_c185 bl[185] br[185] wl[99] vdd gnd cell_6t
Xbit_r100_c185 bl[185] br[185] wl[100] vdd gnd cell_6t
Xbit_r101_c185 bl[185] br[185] wl[101] vdd gnd cell_6t
Xbit_r102_c185 bl[185] br[185] wl[102] vdd gnd cell_6t
Xbit_r103_c185 bl[185] br[185] wl[103] vdd gnd cell_6t
Xbit_r104_c185 bl[185] br[185] wl[104] vdd gnd cell_6t
Xbit_r105_c185 bl[185] br[185] wl[105] vdd gnd cell_6t
Xbit_r106_c185 bl[185] br[185] wl[106] vdd gnd cell_6t
Xbit_r107_c185 bl[185] br[185] wl[107] vdd gnd cell_6t
Xbit_r108_c185 bl[185] br[185] wl[108] vdd gnd cell_6t
Xbit_r109_c185 bl[185] br[185] wl[109] vdd gnd cell_6t
Xbit_r110_c185 bl[185] br[185] wl[110] vdd gnd cell_6t
Xbit_r111_c185 bl[185] br[185] wl[111] vdd gnd cell_6t
Xbit_r112_c185 bl[185] br[185] wl[112] vdd gnd cell_6t
Xbit_r113_c185 bl[185] br[185] wl[113] vdd gnd cell_6t
Xbit_r114_c185 bl[185] br[185] wl[114] vdd gnd cell_6t
Xbit_r115_c185 bl[185] br[185] wl[115] vdd gnd cell_6t
Xbit_r116_c185 bl[185] br[185] wl[116] vdd gnd cell_6t
Xbit_r117_c185 bl[185] br[185] wl[117] vdd gnd cell_6t
Xbit_r118_c185 bl[185] br[185] wl[118] vdd gnd cell_6t
Xbit_r119_c185 bl[185] br[185] wl[119] vdd gnd cell_6t
Xbit_r120_c185 bl[185] br[185] wl[120] vdd gnd cell_6t
Xbit_r121_c185 bl[185] br[185] wl[121] vdd gnd cell_6t
Xbit_r122_c185 bl[185] br[185] wl[122] vdd gnd cell_6t
Xbit_r123_c185 bl[185] br[185] wl[123] vdd gnd cell_6t
Xbit_r124_c185 bl[185] br[185] wl[124] vdd gnd cell_6t
Xbit_r125_c185 bl[185] br[185] wl[125] vdd gnd cell_6t
Xbit_r126_c185 bl[185] br[185] wl[126] vdd gnd cell_6t
Xbit_r127_c185 bl[185] br[185] wl[127] vdd gnd cell_6t
Xbit_r0_c186 bl[186] br[186] wl[0] vdd gnd cell_6t
Xbit_r1_c186 bl[186] br[186] wl[1] vdd gnd cell_6t
Xbit_r2_c186 bl[186] br[186] wl[2] vdd gnd cell_6t
Xbit_r3_c186 bl[186] br[186] wl[3] vdd gnd cell_6t
Xbit_r4_c186 bl[186] br[186] wl[4] vdd gnd cell_6t
Xbit_r5_c186 bl[186] br[186] wl[5] vdd gnd cell_6t
Xbit_r6_c186 bl[186] br[186] wl[6] vdd gnd cell_6t
Xbit_r7_c186 bl[186] br[186] wl[7] vdd gnd cell_6t
Xbit_r8_c186 bl[186] br[186] wl[8] vdd gnd cell_6t
Xbit_r9_c186 bl[186] br[186] wl[9] vdd gnd cell_6t
Xbit_r10_c186 bl[186] br[186] wl[10] vdd gnd cell_6t
Xbit_r11_c186 bl[186] br[186] wl[11] vdd gnd cell_6t
Xbit_r12_c186 bl[186] br[186] wl[12] vdd gnd cell_6t
Xbit_r13_c186 bl[186] br[186] wl[13] vdd gnd cell_6t
Xbit_r14_c186 bl[186] br[186] wl[14] vdd gnd cell_6t
Xbit_r15_c186 bl[186] br[186] wl[15] vdd gnd cell_6t
Xbit_r16_c186 bl[186] br[186] wl[16] vdd gnd cell_6t
Xbit_r17_c186 bl[186] br[186] wl[17] vdd gnd cell_6t
Xbit_r18_c186 bl[186] br[186] wl[18] vdd gnd cell_6t
Xbit_r19_c186 bl[186] br[186] wl[19] vdd gnd cell_6t
Xbit_r20_c186 bl[186] br[186] wl[20] vdd gnd cell_6t
Xbit_r21_c186 bl[186] br[186] wl[21] vdd gnd cell_6t
Xbit_r22_c186 bl[186] br[186] wl[22] vdd gnd cell_6t
Xbit_r23_c186 bl[186] br[186] wl[23] vdd gnd cell_6t
Xbit_r24_c186 bl[186] br[186] wl[24] vdd gnd cell_6t
Xbit_r25_c186 bl[186] br[186] wl[25] vdd gnd cell_6t
Xbit_r26_c186 bl[186] br[186] wl[26] vdd gnd cell_6t
Xbit_r27_c186 bl[186] br[186] wl[27] vdd gnd cell_6t
Xbit_r28_c186 bl[186] br[186] wl[28] vdd gnd cell_6t
Xbit_r29_c186 bl[186] br[186] wl[29] vdd gnd cell_6t
Xbit_r30_c186 bl[186] br[186] wl[30] vdd gnd cell_6t
Xbit_r31_c186 bl[186] br[186] wl[31] vdd gnd cell_6t
Xbit_r32_c186 bl[186] br[186] wl[32] vdd gnd cell_6t
Xbit_r33_c186 bl[186] br[186] wl[33] vdd gnd cell_6t
Xbit_r34_c186 bl[186] br[186] wl[34] vdd gnd cell_6t
Xbit_r35_c186 bl[186] br[186] wl[35] vdd gnd cell_6t
Xbit_r36_c186 bl[186] br[186] wl[36] vdd gnd cell_6t
Xbit_r37_c186 bl[186] br[186] wl[37] vdd gnd cell_6t
Xbit_r38_c186 bl[186] br[186] wl[38] vdd gnd cell_6t
Xbit_r39_c186 bl[186] br[186] wl[39] vdd gnd cell_6t
Xbit_r40_c186 bl[186] br[186] wl[40] vdd gnd cell_6t
Xbit_r41_c186 bl[186] br[186] wl[41] vdd gnd cell_6t
Xbit_r42_c186 bl[186] br[186] wl[42] vdd gnd cell_6t
Xbit_r43_c186 bl[186] br[186] wl[43] vdd gnd cell_6t
Xbit_r44_c186 bl[186] br[186] wl[44] vdd gnd cell_6t
Xbit_r45_c186 bl[186] br[186] wl[45] vdd gnd cell_6t
Xbit_r46_c186 bl[186] br[186] wl[46] vdd gnd cell_6t
Xbit_r47_c186 bl[186] br[186] wl[47] vdd gnd cell_6t
Xbit_r48_c186 bl[186] br[186] wl[48] vdd gnd cell_6t
Xbit_r49_c186 bl[186] br[186] wl[49] vdd gnd cell_6t
Xbit_r50_c186 bl[186] br[186] wl[50] vdd gnd cell_6t
Xbit_r51_c186 bl[186] br[186] wl[51] vdd gnd cell_6t
Xbit_r52_c186 bl[186] br[186] wl[52] vdd gnd cell_6t
Xbit_r53_c186 bl[186] br[186] wl[53] vdd gnd cell_6t
Xbit_r54_c186 bl[186] br[186] wl[54] vdd gnd cell_6t
Xbit_r55_c186 bl[186] br[186] wl[55] vdd gnd cell_6t
Xbit_r56_c186 bl[186] br[186] wl[56] vdd gnd cell_6t
Xbit_r57_c186 bl[186] br[186] wl[57] vdd gnd cell_6t
Xbit_r58_c186 bl[186] br[186] wl[58] vdd gnd cell_6t
Xbit_r59_c186 bl[186] br[186] wl[59] vdd gnd cell_6t
Xbit_r60_c186 bl[186] br[186] wl[60] vdd gnd cell_6t
Xbit_r61_c186 bl[186] br[186] wl[61] vdd gnd cell_6t
Xbit_r62_c186 bl[186] br[186] wl[62] vdd gnd cell_6t
Xbit_r63_c186 bl[186] br[186] wl[63] vdd gnd cell_6t
Xbit_r64_c186 bl[186] br[186] wl[64] vdd gnd cell_6t
Xbit_r65_c186 bl[186] br[186] wl[65] vdd gnd cell_6t
Xbit_r66_c186 bl[186] br[186] wl[66] vdd gnd cell_6t
Xbit_r67_c186 bl[186] br[186] wl[67] vdd gnd cell_6t
Xbit_r68_c186 bl[186] br[186] wl[68] vdd gnd cell_6t
Xbit_r69_c186 bl[186] br[186] wl[69] vdd gnd cell_6t
Xbit_r70_c186 bl[186] br[186] wl[70] vdd gnd cell_6t
Xbit_r71_c186 bl[186] br[186] wl[71] vdd gnd cell_6t
Xbit_r72_c186 bl[186] br[186] wl[72] vdd gnd cell_6t
Xbit_r73_c186 bl[186] br[186] wl[73] vdd gnd cell_6t
Xbit_r74_c186 bl[186] br[186] wl[74] vdd gnd cell_6t
Xbit_r75_c186 bl[186] br[186] wl[75] vdd gnd cell_6t
Xbit_r76_c186 bl[186] br[186] wl[76] vdd gnd cell_6t
Xbit_r77_c186 bl[186] br[186] wl[77] vdd gnd cell_6t
Xbit_r78_c186 bl[186] br[186] wl[78] vdd gnd cell_6t
Xbit_r79_c186 bl[186] br[186] wl[79] vdd gnd cell_6t
Xbit_r80_c186 bl[186] br[186] wl[80] vdd gnd cell_6t
Xbit_r81_c186 bl[186] br[186] wl[81] vdd gnd cell_6t
Xbit_r82_c186 bl[186] br[186] wl[82] vdd gnd cell_6t
Xbit_r83_c186 bl[186] br[186] wl[83] vdd gnd cell_6t
Xbit_r84_c186 bl[186] br[186] wl[84] vdd gnd cell_6t
Xbit_r85_c186 bl[186] br[186] wl[85] vdd gnd cell_6t
Xbit_r86_c186 bl[186] br[186] wl[86] vdd gnd cell_6t
Xbit_r87_c186 bl[186] br[186] wl[87] vdd gnd cell_6t
Xbit_r88_c186 bl[186] br[186] wl[88] vdd gnd cell_6t
Xbit_r89_c186 bl[186] br[186] wl[89] vdd gnd cell_6t
Xbit_r90_c186 bl[186] br[186] wl[90] vdd gnd cell_6t
Xbit_r91_c186 bl[186] br[186] wl[91] vdd gnd cell_6t
Xbit_r92_c186 bl[186] br[186] wl[92] vdd gnd cell_6t
Xbit_r93_c186 bl[186] br[186] wl[93] vdd gnd cell_6t
Xbit_r94_c186 bl[186] br[186] wl[94] vdd gnd cell_6t
Xbit_r95_c186 bl[186] br[186] wl[95] vdd gnd cell_6t
Xbit_r96_c186 bl[186] br[186] wl[96] vdd gnd cell_6t
Xbit_r97_c186 bl[186] br[186] wl[97] vdd gnd cell_6t
Xbit_r98_c186 bl[186] br[186] wl[98] vdd gnd cell_6t
Xbit_r99_c186 bl[186] br[186] wl[99] vdd gnd cell_6t
Xbit_r100_c186 bl[186] br[186] wl[100] vdd gnd cell_6t
Xbit_r101_c186 bl[186] br[186] wl[101] vdd gnd cell_6t
Xbit_r102_c186 bl[186] br[186] wl[102] vdd gnd cell_6t
Xbit_r103_c186 bl[186] br[186] wl[103] vdd gnd cell_6t
Xbit_r104_c186 bl[186] br[186] wl[104] vdd gnd cell_6t
Xbit_r105_c186 bl[186] br[186] wl[105] vdd gnd cell_6t
Xbit_r106_c186 bl[186] br[186] wl[106] vdd gnd cell_6t
Xbit_r107_c186 bl[186] br[186] wl[107] vdd gnd cell_6t
Xbit_r108_c186 bl[186] br[186] wl[108] vdd gnd cell_6t
Xbit_r109_c186 bl[186] br[186] wl[109] vdd gnd cell_6t
Xbit_r110_c186 bl[186] br[186] wl[110] vdd gnd cell_6t
Xbit_r111_c186 bl[186] br[186] wl[111] vdd gnd cell_6t
Xbit_r112_c186 bl[186] br[186] wl[112] vdd gnd cell_6t
Xbit_r113_c186 bl[186] br[186] wl[113] vdd gnd cell_6t
Xbit_r114_c186 bl[186] br[186] wl[114] vdd gnd cell_6t
Xbit_r115_c186 bl[186] br[186] wl[115] vdd gnd cell_6t
Xbit_r116_c186 bl[186] br[186] wl[116] vdd gnd cell_6t
Xbit_r117_c186 bl[186] br[186] wl[117] vdd gnd cell_6t
Xbit_r118_c186 bl[186] br[186] wl[118] vdd gnd cell_6t
Xbit_r119_c186 bl[186] br[186] wl[119] vdd gnd cell_6t
Xbit_r120_c186 bl[186] br[186] wl[120] vdd gnd cell_6t
Xbit_r121_c186 bl[186] br[186] wl[121] vdd gnd cell_6t
Xbit_r122_c186 bl[186] br[186] wl[122] vdd gnd cell_6t
Xbit_r123_c186 bl[186] br[186] wl[123] vdd gnd cell_6t
Xbit_r124_c186 bl[186] br[186] wl[124] vdd gnd cell_6t
Xbit_r125_c186 bl[186] br[186] wl[125] vdd gnd cell_6t
Xbit_r126_c186 bl[186] br[186] wl[126] vdd gnd cell_6t
Xbit_r127_c186 bl[186] br[186] wl[127] vdd gnd cell_6t
Xbit_r0_c187 bl[187] br[187] wl[0] vdd gnd cell_6t
Xbit_r1_c187 bl[187] br[187] wl[1] vdd gnd cell_6t
Xbit_r2_c187 bl[187] br[187] wl[2] vdd gnd cell_6t
Xbit_r3_c187 bl[187] br[187] wl[3] vdd gnd cell_6t
Xbit_r4_c187 bl[187] br[187] wl[4] vdd gnd cell_6t
Xbit_r5_c187 bl[187] br[187] wl[5] vdd gnd cell_6t
Xbit_r6_c187 bl[187] br[187] wl[6] vdd gnd cell_6t
Xbit_r7_c187 bl[187] br[187] wl[7] vdd gnd cell_6t
Xbit_r8_c187 bl[187] br[187] wl[8] vdd gnd cell_6t
Xbit_r9_c187 bl[187] br[187] wl[9] vdd gnd cell_6t
Xbit_r10_c187 bl[187] br[187] wl[10] vdd gnd cell_6t
Xbit_r11_c187 bl[187] br[187] wl[11] vdd gnd cell_6t
Xbit_r12_c187 bl[187] br[187] wl[12] vdd gnd cell_6t
Xbit_r13_c187 bl[187] br[187] wl[13] vdd gnd cell_6t
Xbit_r14_c187 bl[187] br[187] wl[14] vdd gnd cell_6t
Xbit_r15_c187 bl[187] br[187] wl[15] vdd gnd cell_6t
Xbit_r16_c187 bl[187] br[187] wl[16] vdd gnd cell_6t
Xbit_r17_c187 bl[187] br[187] wl[17] vdd gnd cell_6t
Xbit_r18_c187 bl[187] br[187] wl[18] vdd gnd cell_6t
Xbit_r19_c187 bl[187] br[187] wl[19] vdd gnd cell_6t
Xbit_r20_c187 bl[187] br[187] wl[20] vdd gnd cell_6t
Xbit_r21_c187 bl[187] br[187] wl[21] vdd gnd cell_6t
Xbit_r22_c187 bl[187] br[187] wl[22] vdd gnd cell_6t
Xbit_r23_c187 bl[187] br[187] wl[23] vdd gnd cell_6t
Xbit_r24_c187 bl[187] br[187] wl[24] vdd gnd cell_6t
Xbit_r25_c187 bl[187] br[187] wl[25] vdd gnd cell_6t
Xbit_r26_c187 bl[187] br[187] wl[26] vdd gnd cell_6t
Xbit_r27_c187 bl[187] br[187] wl[27] vdd gnd cell_6t
Xbit_r28_c187 bl[187] br[187] wl[28] vdd gnd cell_6t
Xbit_r29_c187 bl[187] br[187] wl[29] vdd gnd cell_6t
Xbit_r30_c187 bl[187] br[187] wl[30] vdd gnd cell_6t
Xbit_r31_c187 bl[187] br[187] wl[31] vdd gnd cell_6t
Xbit_r32_c187 bl[187] br[187] wl[32] vdd gnd cell_6t
Xbit_r33_c187 bl[187] br[187] wl[33] vdd gnd cell_6t
Xbit_r34_c187 bl[187] br[187] wl[34] vdd gnd cell_6t
Xbit_r35_c187 bl[187] br[187] wl[35] vdd gnd cell_6t
Xbit_r36_c187 bl[187] br[187] wl[36] vdd gnd cell_6t
Xbit_r37_c187 bl[187] br[187] wl[37] vdd gnd cell_6t
Xbit_r38_c187 bl[187] br[187] wl[38] vdd gnd cell_6t
Xbit_r39_c187 bl[187] br[187] wl[39] vdd gnd cell_6t
Xbit_r40_c187 bl[187] br[187] wl[40] vdd gnd cell_6t
Xbit_r41_c187 bl[187] br[187] wl[41] vdd gnd cell_6t
Xbit_r42_c187 bl[187] br[187] wl[42] vdd gnd cell_6t
Xbit_r43_c187 bl[187] br[187] wl[43] vdd gnd cell_6t
Xbit_r44_c187 bl[187] br[187] wl[44] vdd gnd cell_6t
Xbit_r45_c187 bl[187] br[187] wl[45] vdd gnd cell_6t
Xbit_r46_c187 bl[187] br[187] wl[46] vdd gnd cell_6t
Xbit_r47_c187 bl[187] br[187] wl[47] vdd gnd cell_6t
Xbit_r48_c187 bl[187] br[187] wl[48] vdd gnd cell_6t
Xbit_r49_c187 bl[187] br[187] wl[49] vdd gnd cell_6t
Xbit_r50_c187 bl[187] br[187] wl[50] vdd gnd cell_6t
Xbit_r51_c187 bl[187] br[187] wl[51] vdd gnd cell_6t
Xbit_r52_c187 bl[187] br[187] wl[52] vdd gnd cell_6t
Xbit_r53_c187 bl[187] br[187] wl[53] vdd gnd cell_6t
Xbit_r54_c187 bl[187] br[187] wl[54] vdd gnd cell_6t
Xbit_r55_c187 bl[187] br[187] wl[55] vdd gnd cell_6t
Xbit_r56_c187 bl[187] br[187] wl[56] vdd gnd cell_6t
Xbit_r57_c187 bl[187] br[187] wl[57] vdd gnd cell_6t
Xbit_r58_c187 bl[187] br[187] wl[58] vdd gnd cell_6t
Xbit_r59_c187 bl[187] br[187] wl[59] vdd gnd cell_6t
Xbit_r60_c187 bl[187] br[187] wl[60] vdd gnd cell_6t
Xbit_r61_c187 bl[187] br[187] wl[61] vdd gnd cell_6t
Xbit_r62_c187 bl[187] br[187] wl[62] vdd gnd cell_6t
Xbit_r63_c187 bl[187] br[187] wl[63] vdd gnd cell_6t
Xbit_r64_c187 bl[187] br[187] wl[64] vdd gnd cell_6t
Xbit_r65_c187 bl[187] br[187] wl[65] vdd gnd cell_6t
Xbit_r66_c187 bl[187] br[187] wl[66] vdd gnd cell_6t
Xbit_r67_c187 bl[187] br[187] wl[67] vdd gnd cell_6t
Xbit_r68_c187 bl[187] br[187] wl[68] vdd gnd cell_6t
Xbit_r69_c187 bl[187] br[187] wl[69] vdd gnd cell_6t
Xbit_r70_c187 bl[187] br[187] wl[70] vdd gnd cell_6t
Xbit_r71_c187 bl[187] br[187] wl[71] vdd gnd cell_6t
Xbit_r72_c187 bl[187] br[187] wl[72] vdd gnd cell_6t
Xbit_r73_c187 bl[187] br[187] wl[73] vdd gnd cell_6t
Xbit_r74_c187 bl[187] br[187] wl[74] vdd gnd cell_6t
Xbit_r75_c187 bl[187] br[187] wl[75] vdd gnd cell_6t
Xbit_r76_c187 bl[187] br[187] wl[76] vdd gnd cell_6t
Xbit_r77_c187 bl[187] br[187] wl[77] vdd gnd cell_6t
Xbit_r78_c187 bl[187] br[187] wl[78] vdd gnd cell_6t
Xbit_r79_c187 bl[187] br[187] wl[79] vdd gnd cell_6t
Xbit_r80_c187 bl[187] br[187] wl[80] vdd gnd cell_6t
Xbit_r81_c187 bl[187] br[187] wl[81] vdd gnd cell_6t
Xbit_r82_c187 bl[187] br[187] wl[82] vdd gnd cell_6t
Xbit_r83_c187 bl[187] br[187] wl[83] vdd gnd cell_6t
Xbit_r84_c187 bl[187] br[187] wl[84] vdd gnd cell_6t
Xbit_r85_c187 bl[187] br[187] wl[85] vdd gnd cell_6t
Xbit_r86_c187 bl[187] br[187] wl[86] vdd gnd cell_6t
Xbit_r87_c187 bl[187] br[187] wl[87] vdd gnd cell_6t
Xbit_r88_c187 bl[187] br[187] wl[88] vdd gnd cell_6t
Xbit_r89_c187 bl[187] br[187] wl[89] vdd gnd cell_6t
Xbit_r90_c187 bl[187] br[187] wl[90] vdd gnd cell_6t
Xbit_r91_c187 bl[187] br[187] wl[91] vdd gnd cell_6t
Xbit_r92_c187 bl[187] br[187] wl[92] vdd gnd cell_6t
Xbit_r93_c187 bl[187] br[187] wl[93] vdd gnd cell_6t
Xbit_r94_c187 bl[187] br[187] wl[94] vdd gnd cell_6t
Xbit_r95_c187 bl[187] br[187] wl[95] vdd gnd cell_6t
Xbit_r96_c187 bl[187] br[187] wl[96] vdd gnd cell_6t
Xbit_r97_c187 bl[187] br[187] wl[97] vdd gnd cell_6t
Xbit_r98_c187 bl[187] br[187] wl[98] vdd gnd cell_6t
Xbit_r99_c187 bl[187] br[187] wl[99] vdd gnd cell_6t
Xbit_r100_c187 bl[187] br[187] wl[100] vdd gnd cell_6t
Xbit_r101_c187 bl[187] br[187] wl[101] vdd gnd cell_6t
Xbit_r102_c187 bl[187] br[187] wl[102] vdd gnd cell_6t
Xbit_r103_c187 bl[187] br[187] wl[103] vdd gnd cell_6t
Xbit_r104_c187 bl[187] br[187] wl[104] vdd gnd cell_6t
Xbit_r105_c187 bl[187] br[187] wl[105] vdd gnd cell_6t
Xbit_r106_c187 bl[187] br[187] wl[106] vdd gnd cell_6t
Xbit_r107_c187 bl[187] br[187] wl[107] vdd gnd cell_6t
Xbit_r108_c187 bl[187] br[187] wl[108] vdd gnd cell_6t
Xbit_r109_c187 bl[187] br[187] wl[109] vdd gnd cell_6t
Xbit_r110_c187 bl[187] br[187] wl[110] vdd gnd cell_6t
Xbit_r111_c187 bl[187] br[187] wl[111] vdd gnd cell_6t
Xbit_r112_c187 bl[187] br[187] wl[112] vdd gnd cell_6t
Xbit_r113_c187 bl[187] br[187] wl[113] vdd gnd cell_6t
Xbit_r114_c187 bl[187] br[187] wl[114] vdd gnd cell_6t
Xbit_r115_c187 bl[187] br[187] wl[115] vdd gnd cell_6t
Xbit_r116_c187 bl[187] br[187] wl[116] vdd gnd cell_6t
Xbit_r117_c187 bl[187] br[187] wl[117] vdd gnd cell_6t
Xbit_r118_c187 bl[187] br[187] wl[118] vdd gnd cell_6t
Xbit_r119_c187 bl[187] br[187] wl[119] vdd gnd cell_6t
Xbit_r120_c187 bl[187] br[187] wl[120] vdd gnd cell_6t
Xbit_r121_c187 bl[187] br[187] wl[121] vdd gnd cell_6t
Xbit_r122_c187 bl[187] br[187] wl[122] vdd gnd cell_6t
Xbit_r123_c187 bl[187] br[187] wl[123] vdd gnd cell_6t
Xbit_r124_c187 bl[187] br[187] wl[124] vdd gnd cell_6t
Xbit_r125_c187 bl[187] br[187] wl[125] vdd gnd cell_6t
Xbit_r126_c187 bl[187] br[187] wl[126] vdd gnd cell_6t
Xbit_r127_c187 bl[187] br[187] wl[127] vdd gnd cell_6t
Xbit_r0_c188 bl[188] br[188] wl[0] vdd gnd cell_6t
Xbit_r1_c188 bl[188] br[188] wl[1] vdd gnd cell_6t
Xbit_r2_c188 bl[188] br[188] wl[2] vdd gnd cell_6t
Xbit_r3_c188 bl[188] br[188] wl[3] vdd gnd cell_6t
Xbit_r4_c188 bl[188] br[188] wl[4] vdd gnd cell_6t
Xbit_r5_c188 bl[188] br[188] wl[5] vdd gnd cell_6t
Xbit_r6_c188 bl[188] br[188] wl[6] vdd gnd cell_6t
Xbit_r7_c188 bl[188] br[188] wl[7] vdd gnd cell_6t
Xbit_r8_c188 bl[188] br[188] wl[8] vdd gnd cell_6t
Xbit_r9_c188 bl[188] br[188] wl[9] vdd gnd cell_6t
Xbit_r10_c188 bl[188] br[188] wl[10] vdd gnd cell_6t
Xbit_r11_c188 bl[188] br[188] wl[11] vdd gnd cell_6t
Xbit_r12_c188 bl[188] br[188] wl[12] vdd gnd cell_6t
Xbit_r13_c188 bl[188] br[188] wl[13] vdd gnd cell_6t
Xbit_r14_c188 bl[188] br[188] wl[14] vdd gnd cell_6t
Xbit_r15_c188 bl[188] br[188] wl[15] vdd gnd cell_6t
Xbit_r16_c188 bl[188] br[188] wl[16] vdd gnd cell_6t
Xbit_r17_c188 bl[188] br[188] wl[17] vdd gnd cell_6t
Xbit_r18_c188 bl[188] br[188] wl[18] vdd gnd cell_6t
Xbit_r19_c188 bl[188] br[188] wl[19] vdd gnd cell_6t
Xbit_r20_c188 bl[188] br[188] wl[20] vdd gnd cell_6t
Xbit_r21_c188 bl[188] br[188] wl[21] vdd gnd cell_6t
Xbit_r22_c188 bl[188] br[188] wl[22] vdd gnd cell_6t
Xbit_r23_c188 bl[188] br[188] wl[23] vdd gnd cell_6t
Xbit_r24_c188 bl[188] br[188] wl[24] vdd gnd cell_6t
Xbit_r25_c188 bl[188] br[188] wl[25] vdd gnd cell_6t
Xbit_r26_c188 bl[188] br[188] wl[26] vdd gnd cell_6t
Xbit_r27_c188 bl[188] br[188] wl[27] vdd gnd cell_6t
Xbit_r28_c188 bl[188] br[188] wl[28] vdd gnd cell_6t
Xbit_r29_c188 bl[188] br[188] wl[29] vdd gnd cell_6t
Xbit_r30_c188 bl[188] br[188] wl[30] vdd gnd cell_6t
Xbit_r31_c188 bl[188] br[188] wl[31] vdd gnd cell_6t
Xbit_r32_c188 bl[188] br[188] wl[32] vdd gnd cell_6t
Xbit_r33_c188 bl[188] br[188] wl[33] vdd gnd cell_6t
Xbit_r34_c188 bl[188] br[188] wl[34] vdd gnd cell_6t
Xbit_r35_c188 bl[188] br[188] wl[35] vdd gnd cell_6t
Xbit_r36_c188 bl[188] br[188] wl[36] vdd gnd cell_6t
Xbit_r37_c188 bl[188] br[188] wl[37] vdd gnd cell_6t
Xbit_r38_c188 bl[188] br[188] wl[38] vdd gnd cell_6t
Xbit_r39_c188 bl[188] br[188] wl[39] vdd gnd cell_6t
Xbit_r40_c188 bl[188] br[188] wl[40] vdd gnd cell_6t
Xbit_r41_c188 bl[188] br[188] wl[41] vdd gnd cell_6t
Xbit_r42_c188 bl[188] br[188] wl[42] vdd gnd cell_6t
Xbit_r43_c188 bl[188] br[188] wl[43] vdd gnd cell_6t
Xbit_r44_c188 bl[188] br[188] wl[44] vdd gnd cell_6t
Xbit_r45_c188 bl[188] br[188] wl[45] vdd gnd cell_6t
Xbit_r46_c188 bl[188] br[188] wl[46] vdd gnd cell_6t
Xbit_r47_c188 bl[188] br[188] wl[47] vdd gnd cell_6t
Xbit_r48_c188 bl[188] br[188] wl[48] vdd gnd cell_6t
Xbit_r49_c188 bl[188] br[188] wl[49] vdd gnd cell_6t
Xbit_r50_c188 bl[188] br[188] wl[50] vdd gnd cell_6t
Xbit_r51_c188 bl[188] br[188] wl[51] vdd gnd cell_6t
Xbit_r52_c188 bl[188] br[188] wl[52] vdd gnd cell_6t
Xbit_r53_c188 bl[188] br[188] wl[53] vdd gnd cell_6t
Xbit_r54_c188 bl[188] br[188] wl[54] vdd gnd cell_6t
Xbit_r55_c188 bl[188] br[188] wl[55] vdd gnd cell_6t
Xbit_r56_c188 bl[188] br[188] wl[56] vdd gnd cell_6t
Xbit_r57_c188 bl[188] br[188] wl[57] vdd gnd cell_6t
Xbit_r58_c188 bl[188] br[188] wl[58] vdd gnd cell_6t
Xbit_r59_c188 bl[188] br[188] wl[59] vdd gnd cell_6t
Xbit_r60_c188 bl[188] br[188] wl[60] vdd gnd cell_6t
Xbit_r61_c188 bl[188] br[188] wl[61] vdd gnd cell_6t
Xbit_r62_c188 bl[188] br[188] wl[62] vdd gnd cell_6t
Xbit_r63_c188 bl[188] br[188] wl[63] vdd gnd cell_6t
Xbit_r64_c188 bl[188] br[188] wl[64] vdd gnd cell_6t
Xbit_r65_c188 bl[188] br[188] wl[65] vdd gnd cell_6t
Xbit_r66_c188 bl[188] br[188] wl[66] vdd gnd cell_6t
Xbit_r67_c188 bl[188] br[188] wl[67] vdd gnd cell_6t
Xbit_r68_c188 bl[188] br[188] wl[68] vdd gnd cell_6t
Xbit_r69_c188 bl[188] br[188] wl[69] vdd gnd cell_6t
Xbit_r70_c188 bl[188] br[188] wl[70] vdd gnd cell_6t
Xbit_r71_c188 bl[188] br[188] wl[71] vdd gnd cell_6t
Xbit_r72_c188 bl[188] br[188] wl[72] vdd gnd cell_6t
Xbit_r73_c188 bl[188] br[188] wl[73] vdd gnd cell_6t
Xbit_r74_c188 bl[188] br[188] wl[74] vdd gnd cell_6t
Xbit_r75_c188 bl[188] br[188] wl[75] vdd gnd cell_6t
Xbit_r76_c188 bl[188] br[188] wl[76] vdd gnd cell_6t
Xbit_r77_c188 bl[188] br[188] wl[77] vdd gnd cell_6t
Xbit_r78_c188 bl[188] br[188] wl[78] vdd gnd cell_6t
Xbit_r79_c188 bl[188] br[188] wl[79] vdd gnd cell_6t
Xbit_r80_c188 bl[188] br[188] wl[80] vdd gnd cell_6t
Xbit_r81_c188 bl[188] br[188] wl[81] vdd gnd cell_6t
Xbit_r82_c188 bl[188] br[188] wl[82] vdd gnd cell_6t
Xbit_r83_c188 bl[188] br[188] wl[83] vdd gnd cell_6t
Xbit_r84_c188 bl[188] br[188] wl[84] vdd gnd cell_6t
Xbit_r85_c188 bl[188] br[188] wl[85] vdd gnd cell_6t
Xbit_r86_c188 bl[188] br[188] wl[86] vdd gnd cell_6t
Xbit_r87_c188 bl[188] br[188] wl[87] vdd gnd cell_6t
Xbit_r88_c188 bl[188] br[188] wl[88] vdd gnd cell_6t
Xbit_r89_c188 bl[188] br[188] wl[89] vdd gnd cell_6t
Xbit_r90_c188 bl[188] br[188] wl[90] vdd gnd cell_6t
Xbit_r91_c188 bl[188] br[188] wl[91] vdd gnd cell_6t
Xbit_r92_c188 bl[188] br[188] wl[92] vdd gnd cell_6t
Xbit_r93_c188 bl[188] br[188] wl[93] vdd gnd cell_6t
Xbit_r94_c188 bl[188] br[188] wl[94] vdd gnd cell_6t
Xbit_r95_c188 bl[188] br[188] wl[95] vdd gnd cell_6t
Xbit_r96_c188 bl[188] br[188] wl[96] vdd gnd cell_6t
Xbit_r97_c188 bl[188] br[188] wl[97] vdd gnd cell_6t
Xbit_r98_c188 bl[188] br[188] wl[98] vdd gnd cell_6t
Xbit_r99_c188 bl[188] br[188] wl[99] vdd gnd cell_6t
Xbit_r100_c188 bl[188] br[188] wl[100] vdd gnd cell_6t
Xbit_r101_c188 bl[188] br[188] wl[101] vdd gnd cell_6t
Xbit_r102_c188 bl[188] br[188] wl[102] vdd gnd cell_6t
Xbit_r103_c188 bl[188] br[188] wl[103] vdd gnd cell_6t
Xbit_r104_c188 bl[188] br[188] wl[104] vdd gnd cell_6t
Xbit_r105_c188 bl[188] br[188] wl[105] vdd gnd cell_6t
Xbit_r106_c188 bl[188] br[188] wl[106] vdd gnd cell_6t
Xbit_r107_c188 bl[188] br[188] wl[107] vdd gnd cell_6t
Xbit_r108_c188 bl[188] br[188] wl[108] vdd gnd cell_6t
Xbit_r109_c188 bl[188] br[188] wl[109] vdd gnd cell_6t
Xbit_r110_c188 bl[188] br[188] wl[110] vdd gnd cell_6t
Xbit_r111_c188 bl[188] br[188] wl[111] vdd gnd cell_6t
Xbit_r112_c188 bl[188] br[188] wl[112] vdd gnd cell_6t
Xbit_r113_c188 bl[188] br[188] wl[113] vdd gnd cell_6t
Xbit_r114_c188 bl[188] br[188] wl[114] vdd gnd cell_6t
Xbit_r115_c188 bl[188] br[188] wl[115] vdd gnd cell_6t
Xbit_r116_c188 bl[188] br[188] wl[116] vdd gnd cell_6t
Xbit_r117_c188 bl[188] br[188] wl[117] vdd gnd cell_6t
Xbit_r118_c188 bl[188] br[188] wl[118] vdd gnd cell_6t
Xbit_r119_c188 bl[188] br[188] wl[119] vdd gnd cell_6t
Xbit_r120_c188 bl[188] br[188] wl[120] vdd gnd cell_6t
Xbit_r121_c188 bl[188] br[188] wl[121] vdd gnd cell_6t
Xbit_r122_c188 bl[188] br[188] wl[122] vdd gnd cell_6t
Xbit_r123_c188 bl[188] br[188] wl[123] vdd gnd cell_6t
Xbit_r124_c188 bl[188] br[188] wl[124] vdd gnd cell_6t
Xbit_r125_c188 bl[188] br[188] wl[125] vdd gnd cell_6t
Xbit_r126_c188 bl[188] br[188] wl[126] vdd gnd cell_6t
Xbit_r127_c188 bl[188] br[188] wl[127] vdd gnd cell_6t
Xbit_r0_c189 bl[189] br[189] wl[0] vdd gnd cell_6t
Xbit_r1_c189 bl[189] br[189] wl[1] vdd gnd cell_6t
Xbit_r2_c189 bl[189] br[189] wl[2] vdd gnd cell_6t
Xbit_r3_c189 bl[189] br[189] wl[3] vdd gnd cell_6t
Xbit_r4_c189 bl[189] br[189] wl[4] vdd gnd cell_6t
Xbit_r5_c189 bl[189] br[189] wl[5] vdd gnd cell_6t
Xbit_r6_c189 bl[189] br[189] wl[6] vdd gnd cell_6t
Xbit_r7_c189 bl[189] br[189] wl[7] vdd gnd cell_6t
Xbit_r8_c189 bl[189] br[189] wl[8] vdd gnd cell_6t
Xbit_r9_c189 bl[189] br[189] wl[9] vdd gnd cell_6t
Xbit_r10_c189 bl[189] br[189] wl[10] vdd gnd cell_6t
Xbit_r11_c189 bl[189] br[189] wl[11] vdd gnd cell_6t
Xbit_r12_c189 bl[189] br[189] wl[12] vdd gnd cell_6t
Xbit_r13_c189 bl[189] br[189] wl[13] vdd gnd cell_6t
Xbit_r14_c189 bl[189] br[189] wl[14] vdd gnd cell_6t
Xbit_r15_c189 bl[189] br[189] wl[15] vdd gnd cell_6t
Xbit_r16_c189 bl[189] br[189] wl[16] vdd gnd cell_6t
Xbit_r17_c189 bl[189] br[189] wl[17] vdd gnd cell_6t
Xbit_r18_c189 bl[189] br[189] wl[18] vdd gnd cell_6t
Xbit_r19_c189 bl[189] br[189] wl[19] vdd gnd cell_6t
Xbit_r20_c189 bl[189] br[189] wl[20] vdd gnd cell_6t
Xbit_r21_c189 bl[189] br[189] wl[21] vdd gnd cell_6t
Xbit_r22_c189 bl[189] br[189] wl[22] vdd gnd cell_6t
Xbit_r23_c189 bl[189] br[189] wl[23] vdd gnd cell_6t
Xbit_r24_c189 bl[189] br[189] wl[24] vdd gnd cell_6t
Xbit_r25_c189 bl[189] br[189] wl[25] vdd gnd cell_6t
Xbit_r26_c189 bl[189] br[189] wl[26] vdd gnd cell_6t
Xbit_r27_c189 bl[189] br[189] wl[27] vdd gnd cell_6t
Xbit_r28_c189 bl[189] br[189] wl[28] vdd gnd cell_6t
Xbit_r29_c189 bl[189] br[189] wl[29] vdd gnd cell_6t
Xbit_r30_c189 bl[189] br[189] wl[30] vdd gnd cell_6t
Xbit_r31_c189 bl[189] br[189] wl[31] vdd gnd cell_6t
Xbit_r32_c189 bl[189] br[189] wl[32] vdd gnd cell_6t
Xbit_r33_c189 bl[189] br[189] wl[33] vdd gnd cell_6t
Xbit_r34_c189 bl[189] br[189] wl[34] vdd gnd cell_6t
Xbit_r35_c189 bl[189] br[189] wl[35] vdd gnd cell_6t
Xbit_r36_c189 bl[189] br[189] wl[36] vdd gnd cell_6t
Xbit_r37_c189 bl[189] br[189] wl[37] vdd gnd cell_6t
Xbit_r38_c189 bl[189] br[189] wl[38] vdd gnd cell_6t
Xbit_r39_c189 bl[189] br[189] wl[39] vdd gnd cell_6t
Xbit_r40_c189 bl[189] br[189] wl[40] vdd gnd cell_6t
Xbit_r41_c189 bl[189] br[189] wl[41] vdd gnd cell_6t
Xbit_r42_c189 bl[189] br[189] wl[42] vdd gnd cell_6t
Xbit_r43_c189 bl[189] br[189] wl[43] vdd gnd cell_6t
Xbit_r44_c189 bl[189] br[189] wl[44] vdd gnd cell_6t
Xbit_r45_c189 bl[189] br[189] wl[45] vdd gnd cell_6t
Xbit_r46_c189 bl[189] br[189] wl[46] vdd gnd cell_6t
Xbit_r47_c189 bl[189] br[189] wl[47] vdd gnd cell_6t
Xbit_r48_c189 bl[189] br[189] wl[48] vdd gnd cell_6t
Xbit_r49_c189 bl[189] br[189] wl[49] vdd gnd cell_6t
Xbit_r50_c189 bl[189] br[189] wl[50] vdd gnd cell_6t
Xbit_r51_c189 bl[189] br[189] wl[51] vdd gnd cell_6t
Xbit_r52_c189 bl[189] br[189] wl[52] vdd gnd cell_6t
Xbit_r53_c189 bl[189] br[189] wl[53] vdd gnd cell_6t
Xbit_r54_c189 bl[189] br[189] wl[54] vdd gnd cell_6t
Xbit_r55_c189 bl[189] br[189] wl[55] vdd gnd cell_6t
Xbit_r56_c189 bl[189] br[189] wl[56] vdd gnd cell_6t
Xbit_r57_c189 bl[189] br[189] wl[57] vdd gnd cell_6t
Xbit_r58_c189 bl[189] br[189] wl[58] vdd gnd cell_6t
Xbit_r59_c189 bl[189] br[189] wl[59] vdd gnd cell_6t
Xbit_r60_c189 bl[189] br[189] wl[60] vdd gnd cell_6t
Xbit_r61_c189 bl[189] br[189] wl[61] vdd gnd cell_6t
Xbit_r62_c189 bl[189] br[189] wl[62] vdd gnd cell_6t
Xbit_r63_c189 bl[189] br[189] wl[63] vdd gnd cell_6t
Xbit_r64_c189 bl[189] br[189] wl[64] vdd gnd cell_6t
Xbit_r65_c189 bl[189] br[189] wl[65] vdd gnd cell_6t
Xbit_r66_c189 bl[189] br[189] wl[66] vdd gnd cell_6t
Xbit_r67_c189 bl[189] br[189] wl[67] vdd gnd cell_6t
Xbit_r68_c189 bl[189] br[189] wl[68] vdd gnd cell_6t
Xbit_r69_c189 bl[189] br[189] wl[69] vdd gnd cell_6t
Xbit_r70_c189 bl[189] br[189] wl[70] vdd gnd cell_6t
Xbit_r71_c189 bl[189] br[189] wl[71] vdd gnd cell_6t
Xbit_r72_c189 bl[189] br[189] wl[72] vdd gnd cell_6t
Xbit_r73_c189 bl[189] br[189] wl[73] vdd gnd cell_6t
Xbit_r74_c189 bl[189] br[189] wl[74] vdd gnd cell_6t
Xbit_r75_c189 bl[189] br[189] wl[75] vdd gnd cell_6t
Xbit_r76_c189 bl[189] br[189] wl[76] vdd gnd cell_6t
Xbit_r77_c189 bl[189] br[189] wl[77] vdd gnd cell_6t
Xbit_r78_c189 bl[189] br[189] wl[78] vdd gnd cell_6t
Xbit_r79_c189 bl[189] br[189] wl[79] vdd gnd cell_6t
Xbit_r80_c189 bl[189] br[189] wl[80] vdd gnd cell_6t
Xbit_r81_c189 bl[189] br[189] wl[81] vdd gnd cell_6t
Xbit_r82_c189 bl[189] br[189] wl[82] vdd gnd cell_6t
Xbit_r83_c189 bl[189] br[189] wl[83] vdd gnd cell_6t
Xbit_r84_c189 bl[189] br[189] wl[84] vdd gnd cell_6t
Xbit_r85_c189 bl[189] br[189] wl[85] vdd gnd cell_6t
Xbit_r86_c189 bl[189] br[189] wl[86] vdd gnd cell_6t
Xbit_r87_c189 bl[189] br[189] wl[87] vdd gnd cell_6t
Xbit_r88_c189 bl[189] br[189] wl[88] vdd gnd cell_6t
Xbit_r89_c189 bl[189] br[189] wl[89] vdd gnd cell_6t
Xbit_r90_c189 bl[189] br[189] wl[90] vdd gnd cell_6t
Xbit_r91_c189 bl[189] br[189] wl[91] vdd gnd cell_6t
Xbit_r92_c189 bl[189] br[189] wl[92] vdd gnd cell_6t
Xbit_r93_c189 bl[189] br[189] wl[93] vdd gnd cell_6t
Xbit_r94_c189 bl[189] br[189] wl[94] vdd gnd cell_6t
Xbit_r95_c189 bl[189] br[189] wl[95] vdd gnd cell_6t
Xbit_r96_c189 bl[189] br[189] wl[96] vdd gnd cell_6t
Xbit_r97_c189 bl[189] br[189] wl[97] vdd gnd cell_6t
Xbit_r98_c189 bl[189] br[189] wl[98] vdd gnd cell_6t
Xbit_r99_c189 bl[189] br[189] wl[99] vdd gnd cell_6t
Xbit_r100_c189 bl[189] br[189] wl[100] vdd gnd cell_6t
Xbit_r101_c189 bl[189] br[189] wl[101] vdd gnd cell_6t
Xbit_r102_c189 bl[189] br[189] wl[102] vdd gnd cell_6t
Xbit_r103_c189 bl[189] br[189] wl[103] vdd gnd cell_6t
Xbit_r104_c189 bl[189] br[189] wl[104] vdd gnd cell_6t
Xbit_r105_c189 bl[189] br[189] wl[105] vdd gnd cell_6t
Xbit_r106_c189 bl[189] br[189] wl[106] vdd gnd cell_6t
Xbit_r107_c189 bl[189] br[189] wl[107] vdd gnd cell_6t
Xbit_r108_c189 bl[189] br[189] wl[108] vdd gnd cell_6t
Xbit_r109_c189 bl[189] br[189] wl[109] vdd gnd cell_6t
Xbit_r110_c189 bl[189] br[189] wl[110] vdd gnd cell_6t
Xbit_r111_c189 bl[189] br[189] wl[111] vdd gnd cell_6t
Xbit_r112_c189 bl[189] br[189] wl[112] vdd gnd cell_6t
Xbit_r113_c189 bl[189] br[189] wl[113] vdd gnd cell_6t
Xbit_r114_c189 bl[189] br[189] wl[114] vdd gnd cell_6t
Xbit_r115_c189 bl[189] br[189] wl[115] vdd gnd cell_6t
Xbit_r116_c189 bl[189] br[189] wl[116] vdd gnd cell_6t
Xbit_r117_c189 bl[189] br[189] wl[117] vdd gnd cell_6t
Xbit_r118_c189 bl[189] br[189] wl[118] vdd gnd cell_6t
Xbit_r119_c189 bl[189] br[189] wl[119] vdd gnd cell_6t
Xbit_r120_c189 bl[189] br[189] wl[120] vdd gnd cell_6t
Xbit_r121_c189 bl[189] br[189] wl[121] vdd gnd cell_6t
Xbit_r122_c189 bl[189] br[189] wl[122] vdd gnd cell_6t
Xbit_r123_c189 bl[189] br[189] wl[123] vdd gnd cell_6t
Xbit_r124_c189 bl[189] br[189] wl[124] vdd gnd cell_6t
Xbit_r125_c189 bl[189] br[189] wl[125] vdd gnd cell_6t
Xbit_r126_c189 bl[189] br[189] wl[126] vdd gnd cell_6t
Xbit_r127_c189 bl[189] br[189] wl[127] vdd gnd cell_6t
Xbit_r0_c190 bl[190] br[190] wl[0] vdd gnd cell_6t
Xbit_r1_c190 bl[190] br[190] wl[1] vdd gnd cell_6t
Xbit_r2_c190 bl[190] br[190] wl[2] vdd gnd cell_6t
Xbit_r3_c190 bl[190] br[190] wl[3] vdd gnd cell_6t
Xbit_r4_c190 bl[190] br[190] wl[4] vdd gnd cell_6t
Xbit_r5_c190 bl[190] br[190] wl[5] vdd gnd cell_6t
Xbit_r6_c190 bl[190] br[190] wl[6] vdd gnd cell_6t
Xbit_r7_c190 bl[190] br[190] wl[7] vdd gnd cell_6t
Xbit_r8_c190 bl[190] br[190] wl[8] vdd gnd cell_6t
Xbit_r9_c190 bl[190] br[190] wl[9] vdd gnd cell_6t
Xbit_r10_c190 bl[190] br[190] wl[10] vdd gnd cell_6t
Xbit_r11_c190 bl[190] br[190] wl[11] vdd gnd cell_6t
Xbit_r12_c190 bl[190] br[190] wl[12] vdd gnd cell_6t
Xbit_r13_c190 bl[190] br[190] wl[13] vdd gnd cell_6t
Xbit_r14_c190 bl[190] br[190] wl[14] vdd gnd cell_6t
Xbit_r15_c190 bl[190] br[190] wl[15] vdd gnd cell_6t
Xbit_r16_c190 bl[190] br[190] wl[16] vdd gnd cell_6t
Xbit_r17_c190 bl[190] br[190] wl[17] vdd gnd cell_6t
Xbit_r18_c190 bl[190] br[190] wl[18] vdd gnd cell_6t
Xbit_r19_c190 bl[190] br[190] wl[19] vdd gnd cell_6t
Xbit_r20_c190 bl[190] br[190] wl[20] vdd gnd cell_6t
Xbit_r21_c190 bl[190] br[190] wl[21] vdd gnd cell_6t
Xbit_r22_c190 bl[190] br[190] wl[22] vdd gnd cell_6t
Xbit_r23_c190 bl[190] br[190] wl[23] vdd gnd cell_6t
Xbit_r24_c190 bl[190] br[190] wl[24] vdd gnd cell_6t
Xbit_r25_c190 bl[190] br[190] wl[25] vdd gnd cell_6t
Xbit_r26_c190 bl[190] br[190] wl[26] vdd gnd cell_6t
Xbit_r27_c190 bl[190] br[190] wl[27] vdd gnd cell_6t
Xbit_r28_c190 bl[190] br[190] wl[28] vdd gnd cell_6t
Xbit_r29_c190 bl[190] br[190] wl[29] vdd gnd cell_6t
Xbit_r30_c190 bl[190] br[190] wl[30] vdd gnd cell_6t
Xbit_r31_c190 bl[190] br[190] wl[31] vdd gnd cell_6t
Xbit_r32_c190 bl[190] br[190] wl[32] vdd gnd cell_6t
Xbit_r33_c190 bl[190] br[190] wl[33] vdd gnd cell_6t
Xbit_r34_c190 bl[190] br[190] wl[34] vdd gnd cell_6t
Xbit_r35_c190 bl[190] br[190] wl[35] vdd gnd cell_6t
Xbit_r36_c190 bl[190] br[190] wl[36] vdd gnd cell_6t
Xbit_r37_c190 bl[190] br[190] wl[37] vdd gnd cell_6t
Xbit_r38_c190 bl[190] br[190] wl[38] vdd gnd cell_6t
Xbit_r39_c190 bl[190] br[190] wl[39] vdd gnd cell_6t
Xbit_r40_c190 bl[190] br[190] wl[40] vdd gnd cell_6t
Xbit_r41_c190 bl[190] br[190] wl[41] vdd gnd cell_6t
Xbit_r42_c190 bl[190] br[190] wl[42] vdd gnd cell_6t
Xbit_r43_c190 bl[190] br[190] wl[43] vdd gnd cell_6t
Xbit_r44_c190 bl[190] br[190] wl[44] vdd gnd cell_6t
Xbit_r45_c190 bl[190] br[190] wl[45] vdd gnd cell_6t
Xbit_r46_c190 bl[190] br[190] wl[46] vdd gnd cell_6t
Xbit_r47_c190 bl[190] br[190] wl[47] vdd gnd cell_6t
Xbit_r48_c190 bl[190] br[190] wl[48] vdd gnd cell_6t
Xbit_r49_c190 bl[190] br[190] wl[49] vdd gnd cell_6t
Xbit_r50_c190 bl[190] br[190] wl[50] vdd gnd cell_6t
Xbit_r51_c190 bl[190] br[190] wl[51] vdd gnd cell_6t
Xbit_r52_c190 bl[190] br[190] wl[52] vdd gnd cell_6t
Xbit_r53_c190 bl[190] br[190] wl[53] vdd gnd cell_6t
Xbit_r54_c190 bl[190] br[190] wl[54] vdd gnd cell_6t
Xbit_r55_c190 bl[190] br[190] wl[55] vdd gnd cell_6t
Xbit_r56_c190 bl[190] br[190] wl[56] vdd gnd cell_6t
Xbit_r57_c190 bl[190] br[190] wl[57] vdd gnd cell_6t
Xbit_r58_c190 bl[190] br[190] wl[58] vdd gnd cell_6t
Xbit_r59_c190 bl[190] br[190] wl[59] vdd gnd cell_6t
Xbit_r60_c190 bl[190] br[190] wl[60] vdd gnd cell_6t
Xbit_r61_c190 bl[190] br[190] wl[61] vdd gnd cell_6t
Xbit_r62_c190 bl[190] br[190] wl[62] vdd gnd cell_6t
Xbit_r63_c190 bl[190] br[190] wl[63] vdd gnd cell_6t
Xbit_r64_c190 bl[190] br[190] wl[64] vdd gnd cell_6t
Xbit_r65_c190 bl[190] br[190] wl[65] vdd gnd cell_6t
Xbit_r66_c190 bl[190] br[190] wl[66] vdd gnd cell_6t
Xbit_r67_c190 bl[190] br[190] wl[67] vdd gnd cell_6t
Xbit_r68_c190 bl[190] br[190] wl[68] vdd gnd cell_6t
Xbit_r69_c190 bl[190] br[190] wl[69] vdd gnd cell_6t
Xbit_r70_c190 bl[190] br[190] wl[70] vdd gnd cell_6t
Xbit_r71_c190 bl[190] br[190] wl[71] vdd gnd cell_6t
Xbit_r72_c190 bl[190] br[190] wl[72] vdd gnd cell_6t
Xbit_r73_c190 bl[190] br[190] wl[73] vdd gnd cell_6t
Xbit_r74_c190 bl[190] br[190] wl[74] vdd gnd cell_6t
Xbit_r75_c190 bl[190] br[190] wl[75] vdd gnd cell_6t
Xbit_r76_c190 bl[190] br[190] wl[76] vdd gnd cell_6t
Xbit_r77_c190 bl[190] br[190] wl[77] vdd gnd cell_6t
Xbit_r78_c190 bl[190] br[190] wl[78] vdd gnd cell_6t
Xbit_r79_c190 bl[190] br[190] wl[79] vdd gnd cell_6t
Xbit_r80_c190 bl[190] br[190] wl[80] vdd gnd cell_6t
Xbit_r81_c190 bl[190] br[190] wl[81] vdd gnd cell_6t
Xbit_r82_c190 bl[190] br[190] wl[82] vdd gnd cell_6t
Xbit_r83_c190 bl[190] br[190] wl[83] vdd gnd cell_6t
Xbit_r84_c190 bl[190] br[190] wl[84] vdd gnd cell_6t
Xbit_r85_c190 bl[190] br[190] wl[85] vdd gnd cell_6t
Xbit_r86_c190 bl[190] br[190] wl[86] vdd gnd cell_6t
Xbit_r87_c190 bl[190] br[190] wl[87] vdd gnd cell_6t
Xbit_r88_c190 bl[190] br[190] wl[88] vdd gnd cell_6t
Xbit_r89_c190 bl[190] br[190] wl[89] vdd gnd cell_6t
Xbit_r90_c190 bl[190] br[190] wl[90] vdd gnd cell_6t
Xbit_r91_c190 bl[190] br[190] wl[91] vdd gnd cell_6t
Xbit_r92_c190 bl[190] br[190] wl[92] vdd gnd cell_6t
Xbit_r93_c190 bl[190] br[190] wl[93] vdd gnd cell_6t
Xbit_r94_c190 bl[190] br[190] wl[94] vdd gnd cell_6t
Xbit_r95_c190 bl[190] br[190] wl[95] vdd gnd cell_6t
Xbit_r96_c190 bl[190] br[190] wl[96] vdd gnd cell_6t
Xbit_r97_c190 bl[190] br[190] wl[97] vdd gnd cell_6t
Xbit_r98_c190 bl[190] br[190] wl[98] vdd gnd cell_6t
Xbit_r99_c190 bl[190] br[190] wl[99] vdd gnd cell_6t
Xbit_r100_c190 bl[190] br[190] wl[100] vdd gnd cell_6t
Xbit_r101_c190 bl[190] br[190] wl[101] vdd gnd cell_6t
Xbit_r102_c190 bl[190] br[190] wl[102] vdd gnd cell_6t
Xbit_r103_c190 bl[190] br[190] wl[103] vdd gnd cell_6t
Xbit_r104_c190 bl[190] br[190] wl[104] vdd gnd cell_6t
Xbit_r105_c190 bl[190] br[190] wl[105] vdd gnd cell_6t
Xbit_r106_c190 bl[190] br[190] wl[106] vdd gnd cell_6t
Xbit_r107_c190 bl[190] br[190] wl[107] vdd gnd cell_6t
Xbit_r108_c190 bl[190] br[190] wl[108] vdd gnd cell_6t
Xbit_r109_c190 bl[190] br[190] wl[109] vdd gnd cell_6t
Xbit_r110_c190 bl[190] br[190] wl[110] vdd gnd cell_6t
Xbit_r111_c190 bl[190] br[190] wl[111] vdd gnd cell_6t
Xbit_r112_c190 bl[190] br[190] wl[112] vdd gnd cell_6t
Xbit_r113_c190 bl[190] br[190] wl[113] vdd gnd cell_6t
Xbit_r114_c190 bl[190] br[190] wl[114] vdd gnd cell_6t
Xbit_r115_c190 bl[190] br[190] wl[115] vdd gnd cell_6t
Xbit_r116_c190 bl[190] br[190] wl[116] vdd gnd cell_6t
Xbit_r117_c190 bl[190] br[190] wl[117] vdd gnd cell_6t
Xbit_r118_c190 bl[190] br[190] wl[118] vdd gnd cell_6t
Xbit_r119_c190 bl[190] br[190] wl[119] vdd gnd cell_6t
Xbit_r120_c190 bl[190] br[190] wl[120] vdd gnd cell_6t
Xbit_r121_c190 bl[190] br[190] wl[121] vdd gnd cell_6t
Xbit_r122_c190 bl[190] br[190] wl[122] vdd gnd cell_6t
Xbit_r123_c190 bl[190] br[190] wl[123] vdd gnd cell_6t
Xbit_r124_c190 bl[190] br[190] wl[124] vdd gnd cell_6t
Xbit_r125_c190 bl[190] br[190] wl[125] vdd gnd cell_6t
Xbit_r126_c190 bl[190] br[190] wl[126] vdd gnd cell_6t
Xbit_r127_c190 bl[190] br[190] wl[127] vdd gnd cell_6t
Xbit_r0_c191 bl[191] br[191] wl[0] vdd gnd cell_6t
Xbit_r1_c191 bl[191] br[191] wl[1] vdd gnd cell_6t
Xbit_r2_c191 bl[191] br[191] wl[2] vdd gnd cell_6t
Xbit_r3_c191 bl[191] br[191] wl[3] vdd gnd cell_6t
Xbit_r4_c191 bl[191] br[191] wl[4] vdd gnd cell_6t
Xbit_r5_c191 bl[191] br[191] wl[5] vdd gnd cell_6t
Xbit_r6_c191 bl[191] br[191] wl[6] vdd gnd cell_6t
Xbit_r7_c191 bl[191] br[191] wl[7] vdd gnd cell_6t
Xbit_r8_c191 bl[191] br[191] wl[8] vdd gnd cell_6t
Xbit_r9_c191 bl[191] br[191] wl[9] vdd gnd cell_6t
Xbit_r10_c191 bl[191] br[191] wl[10] vdd gnd cell_6t
Xbit_r11_c191 bl[191] br[191] wl[11] vdd gnd cell_6t
Xbit_r12_c191 bl[191] br[191] wl[12] vdd gnd cell_6t
Xbit_r13_c191 bl[191] br[191] wl[13] vdd gnd cell_6t
Xbit_r14_c191 bl[191] br[191] wl[14] vdd gnd cell_6t
Xbit_r15_c191 bl[191] br[191] wl[15] vdd gnd cell_6t
Xbit_r16_c191 bl[191] br[191] wl[16] vdd gnd cell_6t
Xbit_r17_c191 bl[191] br[191] wl[17] vdd gnd cell_6t
Xbit_r18_c191 bl[191] br[191] wl[18] vdd gnd cell_6t
Xbit_r19_c191 bl[191] br[191] wl[19] vdd gnd cell_6t
Xbit_r20_c191 bl[191] br[191] wl[20] vdd gnd cell_6t
Xbit_r21_c191 bl[191] br[191] wl[21] vdd gnd cell_6t
Xbit_r22_c191 bl[191] br[191] wl[22] vdd gnd cell_6t
Xbit_r23_c191 bl[191] br[191] wl[23] vdd gnd cell_6t
Xbit_r24_c191 bl[191] br[191] wl[24] vdd gnd cell_6t
Xbit_r25_c191 bl[191] br[191] wl[25] vdd gnd cell_6t
Xbit_r26_c191 bl[191] br[191] wl[26] vdd gnd cell_6t
Xbit_r27_c191 bl[191] br[191] wl[27] vdd gnd cell_6t
Xbit_r28_c191 bl[191] br[191] wl[28] vdd gnd cell_6t
Xbit_r29_c191 bl[191] br[191] wl[29] vdd gnd cell_6t
Xbit_r30_c191 bl[191] br[191] wl[30] vdd gnd cell_6t
Xbit_r31_c191 bl[191] br[191] wl[31] vdd gnd cell_6t
Xbit_r32_c191 bl[191] br[191] wl[32] vdd gnd cell_6t
Xbit_r33_c191 bl[191] br[191] wl[33] vdd gnd cell_6t
Xbit_r34_c191 bl[191] br[191] wl[34] vdd gnd cell_6t
Xbit_r35_c191 bl[191] br[191] wl[35] vdd gnd cell_6t
Xbit_r36_c191 bl[191] br[191] wl[36] vdd gnd cell_6t
Xbit_r37_c191 bl[191] br[191] wl[37] vdd gnd cell_6t
Xbit_r38_c191 bl[191] br[191] wl[38] vdd gnd cell_6t
Xbit_r39_c191 bl[191] br[191] wl[39] vdd gnd cell_6t
Xbit_r40_c191 bl[191] br[191] wl[40] vdd gnd cell_6t
Xbit_r41_c191 bl[191] br[191] wl[41] vdd gnd cell_6t
Xbit_r42_c191 bl[191] br[191] wl[42] vdd gnd cell_6t
Xbit_r43_c191 bl[191] br[191] wl[43] vdd gnd cell_6t
Xbit_r44_c191 bl[191] br[191] wl[44] vdd gnd cell_6t
Xbit_r45_c191 bl[191] br[191] wl[45] vdd gnd cell_6t
Xbit_r46_c191 bl[191] br[191] wl[46] vdd gnd cell_6t
Xbit_r47_c191 bl[191] br[191] wl[47] vdd gnd cell_6t
Xbit_r48_c191 bl[191] br[191] wl[48] vdd gnd cell_6t
Xbit_r49_c191 bl[191] br[191] wl[49] vdd gnd cell_6t
Xbit_r50_c191 bl[191] br[191] wl[50] vdd gnd cell_6t
Xbit_r51_c191 bl[191] br[191] wl[51] vdd gnd cell_6t
Xbit_r52_c191 bl[191] br[191] wl[52] vdd gnd cell_6t
Xbit_r53_c191 bl[191] br[191] wl[53] vdd gnd cell_6t
Xbit_r54_c191 bl[191] br[191] wl[54] vdd gnd cell_6t
Xbit_r55_c191 bl[191] br[191] wl[55] vdd gnd cell_6t
Xbit_r56_c191 bl[191] br[191] wl[56] vdd gnd cell_6t
Xbit_r57_c191 bl[191] br[191] wl[57] vdd gnd cell_6t
Xbit_r58_c191 bl[191] br[191] wl[58] vdd gnd cell_6t
Xbit_r59_c191 bl[191] br[191] wl[59] vdd gnd cell_6t
Xbit_r60_c191 bl[191] br[191] wl[60] vdd gnd cell_6t
Xbit_r61_c191 bl[191] br[191] wl[61] vdd gnd cell_6t
Xbit_r62_c191 bl[191] br[191] wl[62] vdd gnd cell_6t
Xbit_r63_c191 bl[191] br[191] wl[63] vdd gnd cell_6t
Xbit_r64_c191 bl[191] br[191] wl[64] vdd gnd cell_6t
Xbit_r65_c191 bl[191] br[191] wl[65] vdd gnd cell_6t
Xbit_r66_c191 bl[191] br[191] wl[66] vdd gnd cell_6t
Xbit_r67_c191 bl[191] br[191] wl[67] vdd gnd cell_6t
Xbit_r68_c191 bl[191] br[191] wl[68] vdd gnd cell_6t
Xbit_r69_c191 bl[191] br[191] wl[69] vdd gnd cell_6t
Xbit_r70_c191 bl[191] br[191] wl[70] vdd gnd cell_6t
Xbit_r71_c191 bl[191] br[191] wl[71] vdd gnd cell_6t
Xbit_r72_c191 bl[191] br[191] wl[72] vdd gnd cell_6t
Xbit_r73_c191 bl[191] br[191] wl[73] vdd gnd cell_6t
Xbit_r74_c191 bl[191] br[191] wl[74] vdd gnd cell_6t
Xbit_r75_c191 bl[191] br[191] wl[75] vdd gnd cell_6t
Xbit_r76_c191 bl[191] br[191] wl[76] vdd gnd cell_6t
Xbit_r77_c191 bl[191] br[191] wl[77] vdd gnd cell_6t
Xbit_r78_c191 bl[191] br[191] wl[78] vdd gnd cell_6t
Xbit_r79_c191 bl[191] br[191] wl[79] vdd gnd cell_6t
Xbit_r80_c191 bl[191] br[191] wl[80] vdd gnd cell_6t
Xbit_r81_c191 bl[191] br[191] wl[81] vdd gnd cell_6t
Xbit_r82_c191 bl[191] br[191] wl[82] vdd gnd cell_6t
Xbit_r83_c191 bl[191] br[191] wl[83] vdd gnd cell_6t
Xbit_r84_c191 bl[191] br[191] wl[84] vdd gnd cell_6t
Xbit_r85_c191 bl[191] br[191] wl[85] vdd gnd cell_6t
Xbit_r86_c191 bl[191] br[191] wl[86] vdd gnd cell_6t
Xbit_r87_c191 bl[191] br[191] wl[87] vdd gnd cell_6t
Xbit_r88_c191 bl[191] br[191] wl[88] vdd gnd cell_6t
Xbit_r89_c191 bl[191] br[191] wl[89] vdd gnd cell_6t
Xbit_r90_c191 bl[191] br[191] wl[90] vdd gnd cell_6t
Xbit_r91_c191 bl[191] br[191] wl[91] vdd gnd cell_6t
Xbit_r92_c191 bl[191] br[191] wl[92] vdd gnd cell_6t
Xbit_r93_c191 bl[191] br[191] wl[93] vdd gnd cell_6t
Xbit_r94_c191 bl[191] br[191] wl[94] vdd gnd cell_6t
Xbit_r95_c191 bl[191] br[191] wl[95] vdd gnd cell_6t
Xbit_r96_c191 bl[191] br[191] wl[96] vdd gnd cell_6t
Xbit_r97_c191 bl[191] br[191] wl[97] vdd gnd cell_6t
Xbit_r98_c191 bl[191] br[191] wl[98] vdd gnd cell_6t
Xbit_r99_c191 bl[191] br[191] wl[99] vdd gnd cell_6t
Xbit_r100_c191 bl[191] br[191] wl[100] vdd gnd cell_6t
Xbit_r101_c191 bl[191] br[191] wl[101] vdd gnd cell_6t
Xbit_r102_c191 bl[191] br[191] wl[102] vdd gnd cell_6t
Xbit_r103_c191 bl[191] br[191] wl[103] vdd gnd cell_6t
Xbit_r104_c191 bl[191] br[191] wl[104] vdd gnd cell_6t
Xbit_r105_c191 bl[191] br[191] wl[105] vdd gnd cell_6t
Xbit_r106_c191 bl[191] br[191] wl[106] vdd gnd cell_6t
Xbit_r107_c191 bl[191] br[191] wl[107] vdd gnd cell_6t
Xbit_r108_c191 bl[191] br[191] wl[108] vdd gnd cell_6t
Xbit_r109_c191 bl[191] br[191] wl[109] vdd gnd cell_6t
Xbit_r110_c191 bl[191] br[191] wl[110] vdd gnd cell_6t
Xbit_r111_c191 bl[191] br[191] wl[111] vdd gnd cell_6t
Xbit_r112_c191 bl[191] br[191] wl[112] vdd gnd cell_6t
Xbit_r113_c191 bl[191] br[191] wl[113] vdd gnd cell_6t
Xbit_r114_c191 bl[191] br[191] wl[114] vdd gnd cell_6t
Xbit_r115_c191 bl[191] br[191] wl[115] vdd gnd cell_6t
Xbit_r116_c191 bl[191] br[191] wl[116] vdd gnd cell_6t
Xbit_r117_c191 bl[191] br[191] wl[117] vdd gnd cell_6t
Xbit_r118_c191 bl[191] br[191] wl[118] vdd gnd cell_6t
Xbit_r119_c191 bl[191] br[191] wl[119] vdd gnd cell_6t
Xbit_r120_c191 bl[191] br[191] wl[120] vdd gnd cell_6t
Xbit_r121_c191 bl[191] br[191] wl[121] vdd gnd cell_6t
Xbit_r122_c191 bl[191] br[191] wl[122] vdd gnd cell_6t
Xbit_r123_c191 bl[191] br[191] wl[123] vdd gnd cell_6t
Xbit_r124_c191 bl[191] br[191] wl[124] vdd gnd cell_6t
Xbit_r125_c191 bl[191] br[191] wl[125] vdd gnd cell_6t
Xbit_r126_c191 bl[191] br[191] wl[126] vdd gnd cell_6t
Xbit_r127_c191 bl[191] br[191] wl[127] vdd gnd cell_6t
Xbit_r0_c192 bl[192] br[192] wl[0] vdd gnd cell_6t
Xbit_r1_c192 bl[192] br[192] wl[1] vdd gnd cell_6t
Xbit_r2_c192 bl[192] br[192] wl[2] vdd gnd cell_6t
Xbit_r3_c192 bl[192] br[192] wl[3] vdd gnd cell_6t
Xbit_r4_c192 bl[192] br[192] wl[4] vdd gnd cell_6t
Xbit_r5_c192 bl[192] br[192] wl[5] vdd gnd cell_6t
Xbit_r6_c192 bl[192] br[192] wl[6] vdd gnd cell_6t
Xbit_r7_c192 bl[192] br[192] wl[7] vdd gnd cell_6t
Xbit_r8_c192 bl[192] br[192] wl[8] vdd gnd cell_6t
Xbit_r9_c192 bl[192] br[192] wl[9] vdd gnd cell_6t
Xbit_r10_c192 bl[192] br[192] wl[10] vdd gnd cell_6t
Xbit_r11_c192 bl[192] br[192] wl[11] vdd gnd cell_6t
Xbit_r12_c192 bl[192] br[192] wl[12] vdd gnd cell_6t
Xbit_r13_c192 bl[192] br[192] wl[13] vdd gnd cell_6t
Xbit_r14_c192 bl[192] br[192] wl[14] vdd gnd cell_6t
Xbit_r15_c192 bl[192] br[192] wl[15] vdd gnd cell_6t
Xbit_r16_c192 bl[192] br[192] wl[16] vdd gnd cell_6t
Xbit_r17_c192 bl[192] br[192] wl[17] vdd gnd cell_6t
Xbit_r18_c192 bl[192] br[192] wl[18] vdd gnd cell_6t
Xbit_r19_c192 bl[192] br[192] wl[19] vdd gnd cell_6t
Xbit_r20_c192 bl[192] br[192] wl[20] vdd gnd cell_6t
Xbit_r21_c192 bl[192] br[192] wl[21] vdd gnd cell_6t
Xbit_r22_c192 bl[192] br[192] wl[22] vdd gnd cell_6t
Xbit_r23_c192 bl[192] br[192] wl[23] vdd gnd cell_6t
Xbit_r24_c192 bl[192] br[192] wl[24] vdd gnd cell_6t
Xbit_r25_c192 bl[192] br[192] wl[25] vdd gnd cell_6t
Xbit_r26_c192 bl[192] br[192] wl[26] vdd gnd cell_6t
Xbit_r27_c192 bl[192] br[192] wl[27] vdd gnd cell_6t
Xbit_r28_c192 bl[192] br[192] wl[28] vdd gnd cell_6t
Xbit_r29_c192 bl[192] br[192] wl[29] vdd gnd cell_6t
Xbit_r30_c192 bl[192] br[192] wl[30] vdd gnd cell_6t
Xbit_r31_c192 bl[192] br[192] wl[31] vdd gnd cell_6t
Xbit_r32_c192 bl[192] br[192] wl[32] vdd gnd cell_6t
Xbit_r33_c192 bl[192] br[192] wl[33] vdd gnd cell_6t
Xbit_r34_c192 bl[192] br[192] wl[34] vdd gnd cell_6t
Xbit_r35_c192 bl[192] br[192] wl[35] vdd gnd cell_6t
Xbit_r36_c192 bl[192] br[192] wl[36] vdd gnd cell_6t
Xbit_r37_c192 bl[192] br[192] wl[37] vdd gnd cell_6t
Xbit_r38_c192 bl[192] br[192] wl[38] vdd gnd cell_6t
Xbit_r39_c192 bl[192] br[192] wl[39] vdd gnd cell_6t
Xbit_r40_c192 bl[192] br[192] wl[40] vdd gnd cell_6t
Xbit_r41_c192 bl[192] br[192] wl[41] vdd gnd cell_6t
Xbit_r42_c192 bl[192] br[192] wl[42] vdd gnd cell_6t
Xbit_r43_c192 bl[192] br[192] wl[43] vdd gnd cell_6t
Xbit_r44_c192 bl[192] br[192] wl[44] vdd gnd cell_6t
Xbit_r45_c192 bl[192] br[192] wl[45] vdd gnd cell_6t
Xbit_r46_c192 bl[192] br[192] wl[46] vdd gnd cell_6t
Xbit_r47_c192 bl[192] br[192] wl[47] vdd gnd cell_6t
Xbit_r48_c192 bl[192] br[192] wl[48] vdd gnd cell_6t
Xbit_r49_c192 bl[192] br[192] wl[49] vdd gnd cell_6t
Xbit_r50_c192 bl[192] br[192] wl[50] vdd gnd cell_6t
Xbit_r51_c192 bl[192] br[192] wl[51] vdd gnd cell_6t
Xbit_r52_c192 bl[192] br[192] wl[52] vdd gnd cell_6t
Xbit_r53_c192 bl[192] br[192] wl[53] vdd gnd cell_6t
Xbit_r54_c192 bl[192] br[192] wl[54] vdd gnd cell_6t
Xbit_r55_c192 bl[192] br[192] wl[55] vdd gnd cell_6t
Xbit_r56_c192 bl[192] br[192] wl[56] vdd gnd cell_6t
Xbit_r57_c192 bl[192] br[192] wl[57] vdd gnd cell_6t
Xbit_r58_c192 bl[192] br[192] wl[58] vdd gnd cell_6t
Xbit_r59_c192 bl[192] br[192] wl[59] vdd gnd cell_6t
Xbit_r60_c192 bl[192] br[192] wl[60] vdd gnd cell_6t
Xbit_r61_c192 bl[192] br[192] wl[61] vdd gnd cell_6t
Xbit_r62_c192 bl[192] br[192] wl[62] vdd gnd cell_6t
Xbit_r63_c192 bl[192] br[192] wl[63] vdd gnd cell_6t
Xbit_r64_c192 bl[192] br[192] wl[64] vdd gnd cell_6t
Xbit_r65_c192 bl[192] br[192] wl[65] vdd gnd cell_6t
Xbit_r66_c192 bl[192] br[192] wl[66] vdd gnd cell_6t
Xbit_r67_c192 bl[192] br[192] wl[67] vdd gnd cell_6t
Xbit_r68_c192 bl[192] br[192] wl[68] vdd gnd cell_6t
Xbit_r69_c192 bl[192] br[192] wl[69] vdd gnd cell_6t
Xbit_r70_c192 bl[192] br[192] wl[70] vdd gnd cell_6t
Xbit_r71_c192 bl[192] br[192] wl[71] vdd gnd cell_6t
Xbit_r72_c192 bl[192] br[192] wl[72] vdd gnd cell_6t
Xbit_r73_c192 bl[192] br[192] wl[73] vdd gnd cell_6t
Xbit_r74_c192 bl[192] br[192] wl[74] vdd gnd cell_6t
Xbit_r75_c192 bl[192] br[192] wl[75] vdd gnd cell_6t
Xbit_r76_c192 bl[192] br[192] wl[76] vdd gnd cell_6t
Xbit_r77_c192 bl[192] br[192] wl[77] vdd gnd cell_6t
Xbit_r78_c192 bl[192] br[192] wl[78] vdd gnd cell_6t
Xbit_r79_c192 bl[192] br[192] wl[79] vdd gnd cell_6t
Xbit_r80_c192 bl[192] br[192] wl[80] vdd gnd cell_6t
Xbit_r81_c192 bl[192] br[192] wl[81] vdd gnd cell_6t
Xbit_r82_c192 bl[192] br[192] wl[82] vdd gnd cell_6t
Xbit_r83_c192 bl[192] br[192] wl[83] vdd gnd cell_6t
Xbit_r84_c192 bl[192] br[192] wl[84] vdd gnd cell_6t
Xbit_r85_c192 bl[192] br[192] wl[85] vdd gnd cell_6t
Xbit_r86_c192 bl[192] br[192] wl[86] vdd gnd cell_6t
Xbit_r87_c192 bl[192] br[192] wl[87] vdd gnd cell_6t
Xbit_r88_c192 bl[192] br[192] wl[88] vdd gnd cell_6t
Xbit_r89_c192 bl[192] br[192] wl[89] vdd gnd cell_6t
Xbit_r90_c192 bl[192] br[192] wl[90] vdd gnd cell_6t
Xbit_r91_c192 bl[192] br[192] wl[91] vdd gnd cell_6t
Xbit_r92_c192 bl[192] br[192] wl[92] vdd gnd cell_6t
Xbit_r93_c192 bl[192] br[192] wl[93] vdd gnd cell_6t
Xbit_r94_c192 bl[192] br[192] wl[94] vdd gnd cell_6t
Xbit_r95_c192 bl[192] br[192] wl[95] vdd gnd cell_6t
Xbit_r96_c192 bl[192] br[192] wl[96] vdd gnd cell_6t
Xbit_r97_c192 bl[192] br[192] wl[97] vdd gnd cell_6t
Xbit_r98_c192 bl[192] br[192] wl[98] vdd gnd cell_6t
Xbit_r99_c192 bl[192] br[192] wl[99] vdd gnd cell_6t
Xbit_r100_c192 bl[192] br[192] wl[100] vdd gnd cell_6t
Xbit_r101_c192 bl[192] br[192] wl[101] vdd gnd cell_6t
Xbit_r102_c192 bl[192] br[192] wl[102] vdd gnd cell_6t
Xbit_r103_c192 bl[192] br[192] wl[103] vdd gnd cell_6t
Xbit_r104_c192 bl[192] br[192] wl[104] vdd gnd cell_6t
Xbit_r105_c192 bl[192] br[192] wl[105] vdd gnd cell_6t
Xbit_r106_c192 bl[192] br[192] wl[106] vdd gnd cell_6t
Xbit_r107_c192 bl[192] br[192] wl[107] vdd gnd cell_6t
Xbit_r108_c192 bl[192] br[192] wl[108] vdd gnd cell_6t
Xbit_r109_c192 bl[192] br[192] wl[109] vdd gnd cell_6t
Xbit_r110_c192 bl[192] br[192] wl[110] vdd gnd cell_6t
Xbit_r111_c192 bl[192] br[192] wl[111] vdd gnd cell_6t
Xbit_r112_c192 bl[192] br[192] wl[112] vdd gnd cell_6t
Xbit_r113_c192 bl[192] br[192] wl[113] vdd gnd cell_6t
Xbit_r114_c192 bl[192] br[192] wl[114] vdd gnd cell_6t
Xbit_r115_c192 bl[192] br[192] wl[115] vdd gnd cell_6t
Xbit_r116_c192 bl[192] br[192] wl[116] vdd gnd cell_6t
Xbit_r117_c192 bl[192] br[192] wl[117] vdd gnd cell_6t
Xbit_r118_c192 bl[192] br[192] wl[118] vdd gnd cell_6t
Xbit_r119_c192 bl[192] br[192] wl[119] vdd gnd cell_6t
Xbit_r120_c192 bl[192] br[192] wl[120] vdd gnd cell_6t
Xbit_r121_c192 bl[192] br[192] wl[121] vdd gnd cell_6t
Xbit_r122_c192 bl[192] br[192] wl[122] vdd gnd cell_6t
Xbit_r123_c192 bl[192] br[192] wl[123] vdd gnd cell_6t
Xbit_r124_c192 bl[192] br[192] wl[124] vdd gnd cell_6t
Xbit_r125_c192 bl[192] br[192] wl[125] vdd gnd cell_6t
Xbit_r126_c192 bl[192] br[192] wl[126] vdd gnd cell_6t
Xbit_r127_c192 bl[192] br[192] wl[127] vdd gnd cell_6t
Xbit_r0_c193 bl[193] br[193] wl[0] vdd gnd cell_6t
Xbit_r1_c193 bl[193] br[193] wl[1] vdd gnd cell_6t
Xbit_r2_c193 bl[193] br[193] wl[2] vdd gnd cell_6t
Xbit_r3_c193 bl[193] br[193] wl[3] vdd gnd cell_6t
Xbit_r4_c193 bl[193] br[193] wl[4] vdd gnd cell_6t
Xbit_r5_c193 bl[193] br[193] wl[5] vdd gnd cell_6t
Xbit_r6_c193 bl[193] br[193] wl[6] vdd gnd cell_6t
Xbit_r7_c193 bl[193] br[193] wl[7] vdd gnd cell_6t
Xbit_r8_c193 bl[193] br[193] wl[8] vdd gnd cell_6t
Xbit_r9_c193 bl[193] br[193] wl[9] vdd gnd cell_6t
Xbit_r10_c193 bl[193] br[193] wl[10] vdd gnd cell_6t
Xbit_r11_c193 bl[193] br[193] wl[11] vdd gnd cell_6t
Xbit_r12_c193 bl[193] br[193] wl[12] vdd gnd cell_6t
Xbit_r13_c193 bl[193] br[193] wl[13] vdd gnd cell_6t
Xbit_r14_c193 bl[193] br[193] wl[14] vdd gnd cell_6t
Xbit_r15_c193 bl[193] br[193] wl[15] vdd gnd cell_6t
Xbit_r16_c193 bl[193] br[193] wl[16] vdd gnd cell_6t
Xbit_r17_c193 bl[193] br[193] wl[17] vdd gnd cell_6t
Xbit_r18_c193 bl[193] br[193] wl[18] vdd gnd cell_6t
Xbit_r19_c193 bl[193] br[193] wl[19] vdd gnd cell_6t
Xbit_r20_c193 bl[193] br[193] wl[20] vdd gnd cell_6t
Xbit_r21_c193 bl[193] br[193] wl[21] vdd gnd cell_6t
Xbit_r22_c193 bl[193] br[193] wl[22] vdd gnd cell_6t
Xbit_r23_c193 bl[193] br[193] wl[23] vdd gnd cell_6t
Xbit_r24_c193 bl[193] br[193] wl[24] vdd gnd cell_6t
Xbit_r25_c193 bl[193] br[193] wl[25] vdd gnd cell_6t
Xbit_r26_c193 bl[193] br[193] wl[26] vdd gnd cell_6t
Xbit_r27_c193 bl[193] br[193] wl[27] vdd gnd cell_6t
Xbit_r28_c193 bl[193] br[193] wl[28] vdd gnd cell_6t
Xbit_r29_c193 bl[193] br[193] wl[29] vdd gnd cell_6t
Xbit_r30_c193 bl[193] br[193] wl[30] vdd gnd cell_6t
Xbit_r31_c193 bl[193] br[193] wl[31] vdd gnd cell_6t
Xbit_r32_c193 bl[193] br[193] wl[32] vdd gnd cell_6t
Xbit_r33_c193 bl[193] br[193] wl[33] vdd gnd cell_6t
Xbit_r34_c193 bl[193] br[193] wl[34] vdd gnd cell_6t
Xbit_r35_c193 bl[193] br[193] wl[35] vdd gnd cell_6t
Xbit_r36_c193 bl[193] br[193] wl[36] vdd gnd cell_6t
Xbit_r37_c193 bl[193] br[193] wl[37] vdd gnd cell_6t
Xbit_r38_c193 bl[193] br[193] wl[38] vdd gnd cell_6t
Xbit_r39_c193 bl[193] br[193] wl[39] vdd gnd cell_6t
Xbit_r40_c193 bl[193] br[193] wl[40] vdd gnd cell_6t
Xbit_r41_c193 bl[193] br[193] wl[41] vdd gnd cell_6t
Xbit_r42_c193 bl[193] br[193] wl[42] vdd gnd cell_6t
Xbit_r43_c193 bl[193] br[193] wl[43] vdd gnd cell_6t
Xbit_r44_c193 bl[193] br[193] wl[44] vdd gnd cell_6t
Xbit_r45_c193 bl[193] br[193] wl[45] vdd gnd cell_6t
Xbit_r46_c193 bl[193] br[193] wl[46] vdd gnd cell_6t
Xbit_r47_c193 bl[193] br[193] wl[47] vdd gnd cell_6t
Xbit_r48_c193 bl[193] br[193] wl[48] vdd gnd cell_6t
Xbit_r49_c193 bl[193] br[193] wl[49] vdd gnd cell_6t
Xbit_r50_c193 bl[193] br[193] wl[50] vdd gnd cell_6t
Xbit_r51_c193 bl[193] br[193] wl[51] vdd gnd cell_6t
Xbit_r52_c193 bl[193] br[193] wl[52] vdd gnd cell_6t
Xbit_r53_c193 bl[193] br[193] wl[53] vdd gnd cell_6t
Xbit_r54_c193 bl[193] br[193] wl[54] vdd gnd cell_6t
Xbit_r55_c193 bl[193] br[193] wl[55] vdd gnd cell_6t
Xbit_r56_c193 bl[193] br[193] wl[56] vdd gnd cell_6t
Xbit_r57_c193 bl[193] br[193] wl[57] vdd gnd cell_6t
Xbit_r58_c193 bl[193] br[193] wl[58] vdd gnd cell_6t
Xbit_r59_c193 bl[193] br[193] wl[59] vdd gnd cell_6t
Xbit_r60_c193 bl[193] br[193] wl[60] vdd gnd cell_6t
Xbit_r61_c193 bl[193] br[193] wl[61] vdd gnd cell_6t
Xbit_r62_c193 bl[193] br[193] wl[62] vdd gnd cell_6t
Xbit_r63_c193 bl[193] br[193] wl[63] vdd gnd cell_6t
Xbit_r64_c193 bl[193] br[193] wl[64] vdd gnd cell_6t
Xbit_r65_c193 bl[193] br[193] wl[65] vdd gnd cell_6t
Xbit_r66_c193 bl[193] br[193] wl[66] vdd gnd cell_6t
Xbit_r67_c193 bl[193] br[193] wl[67] vdd gnd cell_6t
Xbit_r68_c193 bl[193] br[193] wl[68] vdd gnd cell_6t
Xbit_r69_c193 bl[193] br[193] wl[69] vdd gnd cell_6t
Xbit_r70_c193 bl[193] br[193] wl[70] vdd gnd cell_6t
Xbit_r71_c193 bl[193] br[193] wl[71] vdd gnd cell_6t
Xbit_r72_c193 bl[193] br[193] wl[72] vdd gnd cell_6t
Xbit_r73_c193 bl[193] br[193] wl[73] vdd gnd cell_6t
Xbit_r74_c193 bl[193] br[193] wl[74] vdd gnd cell_6t
Xbit_r75_c193 bl[193] br[193] wl[75] vdd gnd cell_6t
Xbit_r76_c193 bl[193] br[193] wl[76] vdd gnd cell_6t
Xbit_r77_c193 bl[193] br[193] wl[77] vdd gnd cell_6t
Xbit_r78_c193 bl[193] br[193] wl[78] vdd gnd cell_6t
Xbit_r79_c193 bl[193] br[193] wl[79] vdd gnd cell_6t
Xbit_r80_c193 bl[193] br[193] wl[80] vdd gnd cell_6t
Xbit_r81_c193 bl[193] br[193] wl[81] vdd gnd cell_6t
Xbit_r82_c193 bl[193] br[193] wl[82] vdd gnd cell_6t
Xbit_r83_c193 bl[193] br[193] wl[83] vdd gnd cell_6t
Xbit_r84_c193 bl[193] br[193] wl[84] vdd gnd cell_6t
Xbit_r85_c193 bl[193] br[193] wl[85] vdd gnd cell_6t
Xbit_r86_c193 bl[193] br[193] wl[86] vdd gnd cell_6t
Xbit_r87_c193 bl[193] br[193] wl[87] vdd gnd cell_6t
Xbit_r88_c193 bl[193] br[193] wl[88] vdd gnd cell_6t
Xbit_r89_c193 bl[193] br[193] wl[89] vdd gnd cell_6t
Xbit_r90_c193 bl[193] br[193] wl[90] vdd gnd cell_6t
Xbit_r91_c193 bl[193] br[193] wl[91] vdd gnd cell_6t
Xbit_r92_c193 bl[193] br[193] wl[92] vdd gnd cell_6t
Xbit_r93_c193 bl[193] br[193] wl[93] vdd gnd cell_6t
Xbit_r94_c193 bl[193] br[193] wl[94] vdd gnd cell_6t
Xbit_r95_c193 bl[193] br[193] wl[95] vdd gnd cell_6t
Xbit_r96_c193 bl[193] br[193] wl[96] vdd gnd cell_6t
Xbit_r97_c193 bl[193] br[193] wl[97] vdd gnd cell_6t
Xbit_r98_c193 bl[193] br[193] wl[98] vdd gnd cell_6t
Xbit_r99_c193 bl[193] br[193] wl[99] vdd gnd cell_6t
Xbit_r100_c193 bl[193] br[193] wl[100] vdd gnd cell_6t
Xbit_r101_c193 bl[193] br[193] wl[101] vdd gnd cell_6t
Xbit_r102_c193 bl[193] br[193] wl[102] vdd gnd cell_6t
Xbit_r103_c193 bl[193] br[193] wl[103] vdd gnd cell_6t
Xbit_r104_c193 bl[193] br[193] wl[104] vdd gnd cell_6t
Xbit_r105_c193 bl[193] br[193] wl[105] vdd gnd cell_6t
Xbit_r106_c193 bl[193] br[193] wl[106] vdd gnd cell_6t
Xbit_r107_c193 bl[193] br[193] wl[107] vdd gnd cell_6t
Xbit_r108_c193 bl[193] br[193] wl[108] vdd gnd cell_6t
Xbit_r109_c193 bl[193] br[193] wl[109] vdd gnd cell_6t
Xbit_r110_c193 bl[193] br[193] wl[110] vdd gnd cell_6t
Xbit_r111_c193 bl[193] br[193] wl[111] vdd gnd cell_6t
Xbit_r112_c193 bl[193] br[193] wl[112] vdd gnd cell_6t
Xbit_r113_c193 bl[193] br[193] wl[113] vdd gnd cell_6t
Xbit_r114_c193 bl[193] br[193] wl[114] vdd gnd cell_6t
Xbit_r115_c193 bl[193] br[193] wl[115] vdd gnd cell_6t
Xbit_r116_c193 bl[193] br[193] wl[116] vdd gnd cell_6t
Xbit_r117_c193 bl[193] br[193] wl[117] vdd gnd cell_6t
Xbit_r118_c193 bl[193] br[193] wl[118] vdd gnd cell_6t
Xbit_r119_c193 bl[193] br[193] wl[119] vdd gnd cell_6t
Xbit_r120_c193 bl[193] br[193] wl[120] vdd gnd cell_6t
Xbit_r121_c193 bl[193] br[193] wl[121] vdd gnd cell_6t
Xbit_r122_c193 bl[193] br[193] wl[122] vdd gnd cell_6t
Xbit_r123_c193 bl[193] br[193] wl[123] vdd gnd cell_6t
Xbit_r124_c193 bl[193] br[193] wl[124] vdd gnd cell_6t
Xbit_r125_c193 bl[193] br[193] wl[125] vdd gnd cell_6t
Xbit_r126_c193 bl[193] br[193] wl[126] vdd gnd cell_6t
Xbit_r127_c193 bl[193] br[193] wl[127] vdd gnd cell_6t
Xbit_r0_c194 bl[194] br[194] wl[0] vdd gnd cell_6t
Xbit_r1_c194 bl[194] br[194] wl[1] vdd gnd cell_6t
Xbit_r2_c194 bl[194] br[194] wl[2] vdd gnd cell_6t
Xbit_r3_c194 bl[194] br[194] wl[3] vdd gnd cell_6t
Xbit_r4_c194 bl[194] br[194] wl[4] vdd gnd cell_6t
Xbit_r5_c194 bl[194] br[194] wl[5] vdd gnd cell_6t
Xbit_r6_c194 bl[194] br[194] wl[6] vdd gnd cell_6t
Xbit_r7_c194 bl[194] br[194] wl[7] vdd gnd cell_6t
Xbit_r8_c194 bl[194] br[194] wl[8] vdd gnd cell_6t
Xbit_r9_c194 bl[194] br[194] wl[9] vdd gnd cell_6t
Xbit_r10_c194 bl[194] br[194] wl[10] vdd gnd cell_6t
Xbit_r11_c194 bl[194] br[194] wl[11] vdd gnd cell_6t
Xbit_r12_c194 bl[194] br[194] wl[12] vdd gnd cell_6t
Xbit_r13_c194 bl[194] br[194] wl[13] vdd gnd cell_6t
Xbit_r14_c194 bl[194] br[194] wl[14] vdd gnd cell_6t
Xbit_r15_c194 bl[194] br[194] wl[15] vdd gnd cell_6t
Xbit_r16_c194 bl[194] br[194] wl[16] vdd gnd cell_6t
Xbit_r17_c194 bl[194] br[194] wl[17] vdd gnd cell_6t
Xbit_r18_c194 bl[194] br[194] wl[18] vdd gnd cell_6t
Xbit_r19_c194 bl[194] br[194] wl[19] vdd gnd cell_6t
Xbit_r20_c194 bl[194] br[194] wl[20] vdd gnd cell_6t
Xbit_r21_c194 bl[194] br[194] wl[21] vdd gnd cell_6t
Xbit_r22_c194 bl[194] br[194] wl[22] vdd gnd cell_6t
Xbit_r23_c194 bl[194] br[194] wl[23] vdd gnd cell_6t
Xbit_r24_c194 bl[194] br[194] wl[24] vdd gnd cell_6t
Xbit_r25_c194 bl[194] br[194] wl[25] vdd gnd cell_6t
Xbit_r26_c194 bl[194] br[194] wl[26] vdd gnd cell_6t
Xbit_r27_c194 bl[194] br[194] wl[27] vdd gnd cell_6t
Xbit_r28_c194 bl[194] br[194] wl[28] vdd gnd cell_6t
Xbit_r29_c194 bl[194] br[194] wl[29] vdd gnd cell_6t
Xbit_r30_c194 bl[194] br[194] wl[30] vdd gnd cell_6t
Xbit_r31_c194 bl[194] br[194] wl[31] vdd gnd cell_6t
Xbit_r32_c194 bl[194] br[194] wl[32] vdd gnd cell_6t
Xbit_r33_c194 bl[194] br[194] wl[33] vdd gnd cell_6t
Xbit_r34_c194 bl[194] br[194] wl[34] vdd gnd cell_6t
Xbit_r35_c194 bl[194] br[194] wl[35] vdd gnd cell_6t
Xbit_r36_c194 bl[194] br[194] wl[36] vdd gnd cell_6t
Xbit_r37_c194 bl[194] br[194] wl[37] vdd gnd cell_6t
Xbit_r38_c194 bl[194] br[194] wl[38] vdd gnd cell_6t
Xbit_r39_c194 bl[194] br[194] wl[39] vdd gnd cell_6t
Xbit_r40_c194 bl[194] br[194] wl[40] vdd gnd cell_6t
Xbit_r41_c194 bl[194] br[194] wl[41] vdd gnd cell_6t
Xbit_r42_c194 bl[194] br[194] wl[42] vdd gnd cell_6t
Xbit_r43_c194 bl[194] br[194] wl[43] vdd gnd cell_6t
Xbit_r44_c194 bl[194] br[194] wl[44] vdd gnd cell_6t
Xbit_r45_c194 bl[194] br[194] wl[45] vdd gnd cell_6t
Xbit_r46_c194 bl[194] br[194] wl[46] vdd gnd cell_6t
Xbit_r47_c194 bl[194] br[194] wl[47] vdd gnd cell_6t
Xbit_r48_c194 bl[194] br[194] wl[48] vdd gnd cell_6t
Xbit_r49_c194 bl[194] br[194] wl[49] vdd gnd cell_6t
Xbit_r50_c194 bl[194] br[194] wl[50] vdd gnd cell_6t
Xbit_r51_c194 bl[194] br[194] wl[51] vdd gnd cell_6t
Xbit_r52_c194 bl[194] br[194] wl[52] vdd gnd cell_6t
Xbit_r53_c194 bl[194] br[194] wl[53] vdd gnd cell_6t
Xbit_r54_c194 bl[194] br[194] wl[54] vdd gnd cell_6t
Xbit_r55_c194 bl[194] br[194] wl[55] vdd gnd cell_6t
Xbit_r56_c194 bl[194] br[194] wl[56] vdd gnd cell_6t
Xbit_r57_c194 bl[194] br[194] wl[57] vdd gnd cell_6t
Xbit_r58_c194 bl[194] br[194] wl[58] vdd gnd cell_6t
Xbit_r59_c194 bl[194] br[194] wl[59] vdd gnd cell_6t
Xbit_r60_c194 bl[194] br[194] wl[60] vdd gnd cell_6t
Xbit_r61_c194 bl[194] br[194] wl[61] vdd gnd cell_6t
Xbit_r62_c194 bl[194] br[194] wl[62] vdd gnd cell_6t
Xbit_r63_c194 bl[194] br[194] wl[63] vdd gnd cell_6t
Xbit_r64_c194 bl[194] br[194] wl[64] vdd gnd cell_6t
Xbit_r65_c194 bl[194] br[194] wl[65] vdd gnd cell_6t
Xbit_r66_c194 bl[194] br[194] wl[66] vdd gnd cell_6t
Xbit_r67_c194 bl[194] br[194] wl[67] vdd gnd cell_6t
Xbit_r68_c194 bl[194] br[194] wl[68] vdd gnd cell_6t
Xbit_r69_c194 bl[194] br[194] wl[69] vdd gnd cell_6t
Xbit_r70_c194 bl[194] br[194] wl[70] vdd gnd cell_6t
Xbit_r71_c194 bl[194] br[194] wl[71] vdd gnd cell_6t
Xbit_r72_c194 bl[194] br[194] wl[72] vdd gnd cell_6t
Xbit_r73_c194 bl[194] br[194] wl[73] vdd gnd cell_6t
Xbit_r74_c194 bl[194] br[194] wl[74] vdd gnd cell_6t
Xbit_r75_c194 bl[194] br[194] wl[75] vdd gnd cell_6t
Xbit_r76_c194 bl[194] br[194] wl[76] vdd gnd cell_6t
Xbit_r77_c194 bl[194] br[194] wl[77] vdd gnd cell_6t
Xbit_r78_c194 bl[194] br[194] wl[78] vdd gnd cell_6t
Xbit_r79_c194 bl[194] br[194] wl[79] vdd gnd cell_6t
Xbit_r80_c194 bl[194] br[194] wl[80] vdd gnd cell_6t
Xbit_r81_c194 bl[194] br[194] wl[81] vdd gnd cell_6t
Xbit_r82_c194 bl[194] br[194] wl[82] vdd gnd cell_6t
Xbit_r83_c194 bl[194] br[194] wl[83] vdd gnd cell_6t
Xbit_r84_c194 bl[194] br[194] wl[84] vdd gnd cell_6t
Xbit_r85_c194 bl[194] br[194] wl[85] vdd gnd cell_6t
Xbit_r86_c194 bl[194] br[194] wl[86] vdd gnd cell_6t
Xbit_r87_c194 bl[194] br[194] wl[87] vdd gnd cell_6t
Xbit_r88_c194 bl[194] br[194] wl[88] vdd gnd cell_6t
Xbit_r89_c194 bl[194] br[194] wl[89] vdd gnd cell_6t
Xbit_r90_c194 bl[194] br[194] wl[90] vdd gnd cell_6t
Xbit_r91_c194 bl[194] br[194] wl[91] vdd gnd cell_6t
Xbit_r92_c194 bl[194] br[194] wl[92] vdd gnd cell_6t
Xbit_r93_c194 bl[194] br[194] wl[93] vdd gnd cell_6t
Xbit_r94_c194 bl[194] br[194] wl[94] vdd gnd cell_6t
Xbit_r95_c194 bl[194] br[194] wl[95] vdd gnd cell_6t
Xbit_r96_c194 bl[194] br[194] wl[96] vdd gnd cell_6t
Xbit_r97_c194 bl[194] br[194] wl[97] vdd gnd cell_6t
Xbit_r98_c194 bl[194] br[194] wl[98] vdd gnd cell_6t
Xbit_r99_c194 bl[194] br[194] wl[99] vdd gnd cell_6t
Xbit_r100_c194 bl[194] br[194] wl[100] vdd gnd cell_6t
Xbit_r101_c194 bl[194] br[194] wl[101] vdd gnd cell_6t
Xbit_r102_c194 bl[194] br[194] wl[102] vdd gnd cell_6t
Xbit_r103_c194 bl[194] br[194] wl[103] vdd gnd cell_6t
Xbit_r104_c194 bl[194] br[194] wl[104] vdd gnd cell_6t
Xbit_r105_c194 bl[194] br[194] wl[105] vdd gnd cell_6t
Xbit_r106_c194 bl[194] br[194] wl[106] vdd gnd cell_6t
Xbit_r107_c194 bl[194] br[194] wl[107] vdd gnd cell_6t
Xbit_r108_c194 bl[194] br[194] wl[108] vdd gnd cell_6t
Xbit_r109_c194 bl[194] br[194] wl[109] vdd gnd cell_6t
Xbit_r110_c194 bl[194] br[194] wl[110] vdd gnd cell_6t
Xbit_r111_c194 bl[194] br[194] wl[111] vdd gnd cell_6t
Xbit_r112_c194 bl[194] br[194] wl[112] vdd gnd cell_6t
Xbit_r113_c194 bl[194] br[194] wl[113] vdd gnd cell_6t
Xbit_r114_c194 bl[194] br[194] wl[114] vdd gnd cell_6t
Xbit_r115_c194 bl[194] br[194] wl[115] vdd gnd cell_6t
Xbit_r116_c194 bl[194] br[194] wl[116] vdd gnd cell_6t
Xbit_r117_c194 bl[194] br[194] wl[117] vdd gnd cell_6t
Xbit_r118_c194 bl[194] br[194] wl[118] vdd gnd cell_6t
Xbit_r119_c194 bl[194] br[194] wl[119] vdd gnd cell_6t
Xbit_r120_c194 bl[194] br[194] wl[120] vdd gnd cell_6t
Xbit_r121_c194 bl[194] br[194] wl[121] vdd gnd cell_6t
Xbit_r122_c194 bl[194] br[194] wl[122] vdd gnd cell_6t
Xbit_r123_c194 bl[194] br[194] wl[123] vdd gnd cell_6t
Xbit_r124_c194 bl[194] br[194] wl[124] vdd gnd cell_6t
Xbit_r125_c194 bl[194] br[194] wl[125] vdd gnd cell_6t
Xbit_r126_c194 bl[194] br[194] wl[126] vdd gnd cell_6t
Xbit_r127_c194 bl[194] br[194] wl[127] vdd gnd cell_6t
Xbit_r0_c195 bl[195] br[195] wl[0] vdd gnd cell_6t
Xbit_r1_c195 bl[195] br[195] wl[1] vdd gnd cell_6t
Xbit_r2_c195 bl[195] br[195] wl[2] vdd gnd cell_6t
Xbit_r3_c195 bl[195] br[195] wl[3] vdd gnd cell_6t
Xbit_r4_c195 bl[195] br[195] wl[4] vdd gnd cell_6t
Xbit_r5_c195 bl[195] br[195] wl[5] vdd gnd cell_6t
Xbit_r6_c195 bl[195] br[195] wl[6] vdd gnd cell_6t
Xbit_r7_c195 bl[195] br[195] wl[7] vdd gnd cell_6t
Xbit_r8_c195 bl[195] br[195] wl[8] vdd gnd cell_6t
Xbit_r9_c195 bl[195] br[195] wl[9] vdd gnd cell_6t
Xbit_r10_c195 bl[195] br[195] wl[10] vdd gnd cell_6t
Xbit_r11_c195 bl[195] br[195] wl[11] vdd gnd cell_6t
Xbit_r12_c195 bl[195] br[195] wl[12] vdd gnd cell_6t
Xbit_r13_c195 bl[195] br[195] wl[13] vdd gnd cell_6t
Xbit_r14_c195 bl[195] br[195] wl[14] vdd gnd cell_6t
Xbit_r15_c195 bl[195] br[195] wl[15] vdd gnd cell_6t
Xbit_r16_c195 bl[195] br[195] wl[16] vdd gnd cell_6t
Xbit_r17_c195 bl[195] br[195] wl[17] vdd gnd cell_6t
Xbit_r18_c195 bl[195] br[195] wl[18] vdd gnd cell_6t
Xbit_r19_c195 bl[195] br[195] wl[19] vdd gnd cell_6t
Xbit_r20_c195 bl[195] br[195] wl[20] vdd gnd cell_6t
Xbit_r21_c195 bl[195] br[195] wl[21] vdd gnd cell_6t
Xbit_r22_c195 bl[195] br[195] wl[22] vdd gnd cell_6t
Xbit_r23_c195 bl[195] br[195] wl[23] vdd gnd cell_6t
Xbit_r24_c195 bl[195] br[195] wl[24] vdd gnd cell_6t
Xbit_r25_c195 bl[195] br[195] wl[25] vdd gnd cell_6t
Xbit_r26_c195 bl[195] br[195] wl[26] vdd gnd cell_6t
Xbit_r27_c195 bl[195] br[195] wl[27] vdd gnd cell_6t
Xbit_r28_c195 bl[195] br[195] wl[28] vdd gnd cell_6t
Xbit_r29_c195 bl[195] br[195] wl[29] vdd gnd cell_6t
Xbit_r30_c195 bl[195] br[195] wl[30] vdd gnd cell_6t
Xbit_r31_c195 bl[195] br[195] wl[31] vdd gnd cell_6t
Xbit_r32_c195 bl[195] br[195] wl[32] vdd gnd cell_6t
Xbit_r33_c195 bl[195] br[195] wl[33] vdd gnd cell_6t
Xbit_r34_c195 bl[195] br[195] wl[34] vdd gnd cell_6t
Xbit_r35_c195 bl[195] br[195] wl[35] vdd gnd cell_6t
Xbit_r36_c195 bl[195] br[195] wl[36] vdd gnd cell_6t
Xbit_r37_c195 bl[195] br[195] wl[37] vdd gnd cell_6t
Xbit_r38_c195 bl[195] br[195] wl[38] vdd gnd cell_6t
Xbit_r39_c195 bl[195] br[195] wl[39] vdd gnd cell_6t
Xbit_r40_c195 bl[195] br[195] wl[40] vdd gnd cell_6t
Xbit_r41_c195 bl[195] br[195] wl[41] vdd gnd cell_6t
Xbit_r42_c195 bl[195] br[195] wl[42] vdd gnd cell_6t
Xbit_r43_c195 bl[195] br[195] wl[43] vdd gnd cell_6t
Xbit_r44_c195 bl[195] br[195] wl[44] vdd gnd cell_6t
Xbit_r45_c195 bl[195] br[195] wl[45] vdd gnd cell_6t
Xbit_r46_c195 bl[195] br[195] wl[46] vdd gnd cell_6t
Xbit_r47_c195 bl[195] br[195] wl[47] vdd gnd cell_6t
Xbit_r48_c195 bl[195] br[195] wl[48] vdd gnd cell_6t
Xbit_r49_c195 bl[195] br[195] wl[49] vdd gnd cell_6t
Xbit_r50_c195 bl[195] br[195] wl[50] vdd gnd cell_6t
Xbit_r51_c195 bl[195] br[195] wl[51] vdd gnd cell_6t
Xbit_r52_c195 bl[195] br[195] wl[52] vdd gnd cell_6t
Xbit_r53_c195 bl[195] br[195] wl[53] vdd gnd cell_6t
Xbit_r54_c195 bl[195] br[195] wl[54] vdd gnd cell_6t
Xbit_r55_c195 bl[195] br[195] wl[55] vdd gnd cell_6t
Xbit_r56_c195 bl[195] br[195] wl[56] vdd gnd cell_6t
Xbit_r57_c195 bl[195] br[195] wl[57] vdd gnd cell_6t
Xbit_r58_c195 bl[195] br[195] wl[58] vdd gnd cell_6t
Xbit_r59_c195 bl[195] br[195] wl[59] vdd gnd cell_6t
Xbit_r60_c195 bl[195] br[195] wl[60] vdd gnd cell_6t
Xbit_r61_c195 bl[195] br[195] wl[61] vdd gnd cell_6t
Xbit_r62_c195 bl[195] br[195] wl[62] vdd gnd cell_6t
Xbit_r63_c195 bl[195] br[195] wl[63] vdd gnd cell_6t
Xbit_r64_c195 bl[195] br[195] wl[64] vdd gnd cell_6t
Xbit_r65_c195 bl[195] br[195] wl[65] vdd gnd cell_6t
Xbit_r66_c195 bl[195] br[195] wl[66] vdd gnd cell_6t
Xbit_r67_c195 bl[195] br[195] wl[67] vdd gnd cell_6t
Xbit_r68_c195 bl[195] br[195] wl[68] vdd gnd cell_6t
Xbit_r69_c195 bl[195] br[195] wl[69] vdd gnd cell_6t
Xbit_r70_c195 bl[195] br[195] wl[70] vdd gnd cell_6t
Xbit_r71_c195 bl[195] br[195] wl[71] vdd gnd cell_6t
Xbit_r72_c195 bl[195] br[195] wl[72] vdd gnd cell_6t
Xbit_r73_c195 bl[195] br[195] wl[73] vdd gnd cell_6t
Xbit_r74_c195 bl[195] br[195] wl[74] vdd gnd cell_6t
Xbit_r75_c195 bl[195] br[195] wl[75] vdd gnd cell_6t
Xbit_r76_c195 bl[195] br[195] wl[76] vdd gnd cell_6t
Xbit_r77_c195 bl[195] br[195] wl[77] vdd gnd cell_6t
Xbit_r78_c195 bl[195] br[195] wl[78] vdd gnd cell_6t
Xbit_r79_c195 bl[195] br[195] wl[79] vdd gnd cell_6t
Xbit_r80_c195 bl[195] br[195] wl[80] vdd gnd cell_6t
Xbit_r81_c195 bl[195] br[195] wl[81] vdd gnd cell_6t
Xbit_r82_c195 bl[195] br[195] wl[82] vdd gnd cell_6t
Xbit_r83_c195 bl[195] br[195] wl[83] vdd gnd cell_6t
Xbit_r84_c195 bl[195] br[195] wl[84] vdd gnd cell_6t
Xbit_r85_c195 bl[195] br[195] wl[85] vdd gnd cell_6t
Xbit_r86_c195 bl[195] br[195] wl[86] vdd gnd cell_6t
Xbit_r87_c195 bl[195] br[195] wl[87] vdd gnd cell_6t
Xbit_r88_c195 bl[195] br[195] wl[88] vdd gnd cell_6t
Xbit_r89_c195 bl[195] br[195] wl[89] vdd gnd cell_6t
Xbit_r90_c195 bl[195] br[195] wl[90] vdd gnd cell_6t
Xbit_r91_c195 bl[195] br[195] wl[91] vdd gnd cell_6t
Xbit_r92_c195 bl[195] br[195] wl[92] vdd gnd cell_6t
Xbit_r93_c195 bl[195] br[195] wl[93] vdd gnd cell_6t
Xbit_r94_c195 bl[195] br[195] wl[94] vdd gnd cell_6t
Xbit_r95_c195 bl[195] br[195] wl[95] vdd gnd cell_6t
Xbit_r96_c195 bl[195] br[195] wl[96] vdd gnd cell_6t
Xbit_r97_c195 bl[195] br[195] wl[97] vdd gnd cell_6t
Xbit_r98_c195 bl[195] br[195] wl[98] vdd gnd cell_6t
Xbit_r99_c195 bl[195] br[195] wl[99] vdd gnd cell_6t
Xbit_r100_c195 bl[195] br[195] wl[100] vdd gnd cell_6t
Xbit_r101_c195 bl[195] br[195] wl[101] vdd gnd cell_6t
Xbit_r102_c195 bl[195] br[195] wl[102] vdd gnd cell_6t
Xbit_r103_c195 bl[195] br[195] wl[103] vdd gnd cell_6t
Xbit_r104_c195 bl[195] br[195] wl[104] vdd gnd cell_6t
Xbit_r105_c195 bl[195] br[195] wl[105] vdd gnd cell_6t
Xbit_r106_c195 bl[195] br[195] wl[106] vdd gnd cell_6t
Xbit_r107_c195 bl[195] br[195] wl[107] vdd gnd cell_6t
Xbit_r108_c195 bl[195] br[195] wl[108] vdd gnd cell_6t
Xbit_r109_c195 bl[195] br[195] wl[109] vdd gnd cell_6t
Xbit_r110_c195 bl[195] br[195] wl[110] vdd gnd cell_6t
Xbit_r111_c195 bl[195] br[195] wl[111] vdd gnd cell_6t
Xbit_r112_c195 bl[195] br[195] wl[112] vdd gnd cell_6t
Xbit_r113_c195 bl[195] br[195] wl[113] vdd gnd cell_6t
Xbit_r114_c195 bl[195] br[195] wl[114] vdd gnd cell_6t
Xbit_r115_c195 bl[195] br[195] wl[115] vdd gnd cell_6t
Xbit_r116_c195 bl[195] br[195] wl[116] vdd gnd cell_6t
Xbit_r117_c195 bl[195] br[195] wl[117] vdd gnd cell_6t
Xbit_r118_c195 bl[195] br[195] wl[118] vdd gnd cell_6t
Xbit_r119_c195 bl[195] br[195] wl[119] vdd gnd cell_6t
Xbit_r120_c195 bl[195] br[195] wl[120] vdd gnd cell_6t
Xbit_r121_c195 bl[195] br[195] wl[121] vdd gnd cell_6t
Xbit_r122_c195 bl[195] br[195] wl[122] vdd gnd cell_6t
Xbit_r123_c195 bl[195] br[195] wl[123] vdd gnd cell_6t
Xbit_r124_c195 bl[195] br[195] wl[124] vdd gnd cell_6t
Xbit_r125_c195 bl[195] br[195] wl[125] vdd gnd cell_6t
Xbit_r126_c195 bl[195] br[195] wl[126] vdd gnd cell_6t
Xbit_r127_c195 bl[195] br[195] wl[127] vdd gnd cell_6t
Xbit_r0_c196 bl[196] br[196] wl[0] vdd gnd cell_6t
Xbit_r1_c196 bl[196] br[196] wl[1] vdd gnd cell_6t
Xbit_r2_c196 bl[196] br[196] wl[2] vdd gnd cell_6t
Xbit_r3_c196 bl[196] br[196] wl[3] vdd gnd cell_6t
Xbit_r4_c196 bl[196] br[196] wl[4] vdd gnd cell_6t
Xbit_r5_c196 bl[196] br[196] wl[5] vdd gnd cell_6t
Xbit_r6_c196 bl[196] br[196] wl[6] vdd gnd cell_6t
Xbit_r7_c196 bl[196] br[196] wl[7] vdd gnd cell_6t
Xbit_r8_c196 bl[196] br[196] wl[8] vdd gnd cell_6t
Xbit_r9_c196 bl[196] br[196] wl[9] vdd gnd cell_6t
Xbit_r10_c196 bl[196] br[196] wl[10] vdd gnd cell_6t
Xbit_r11_c196 bl[196] br[196] wl[11] vdd gnd cell_6t
Xbit_r12_c196 bl[196] br[196] wl[12] vdd gnd cell_6t
Xbit_r13_c196 bl[196] br[196] wl[13] vdd gnd cell_6t
Xbit_r14_c196 bl[196] br[196] wl[14] vdd gnd cell_6t
Xbit_r15_c196 bl[196] br[196] wl[15] vdd gnd cell_6t
Xbit_r16_c196 bl[196] br[196] wl[16] vdd gnd cell_6t
Xbit_r17_c196 bl[196] br[196] wl[17] vdd gnd cell_6t
Xbit_r18_c196 bl[196] br[196] wl[18] vdd gnd cell_6t
Xbit_r19_c196 bl[196] br[196] wl[19] vdd gnd cell_6t
Xbit_r20_c196 bl[196] br[196] wl[20] vdd gnd cell_6t
Xbit_r21_c196 bl[196] br[196] wl[21] vdd gnd cell_6t
Xbit_r22_c196 bl[196] br[196] wl[22] vdd gnd cell_6t
Xbit_r23_c196 bl[196] br[196] wl[23] vdd gnd cell_6t
Xbit_r24_c196 bl[196] br[196] wl[24] vdd gnd cell_6t
Xbit_r25_c196 bl[196] br[196] wl[25] vdd gnd cell_6t
Xbit_r26_c196 bl[196] br[196] wl[26] vdd gnd cell_6t
Xbit_r27_c196 bl[196] br[196] wl[27] vdd gnd cell_6t
Xbit_r28_c196 bl[196] br[196] wl[28] vdd gnd cell_6t
Xbit_r29_c196 bl[196] br[196] wl[29] vdd gnd cell_6t
Xbit_r30_c196 bl[196] br[196] wl[30] vdd gnd cell_6t
Xbit_r31_c196 bl[196] br[196] wl[31] vdd gnd cell_6t
Xbit_r32_c196 bl[196] br[196] wl[32] vdd gnd cell_6t
Xbit_r33_c196 bl[196] br[196] wl[33] vdd gnd cell_6t
Xbit_r34_c196 bl[196] br[196] wl[34] vdd gnd cell_6t
Xbit_r35_c196 bl[196] br[196] wl[35] vdd gnd cell_6t
Xbit_r36_c196 bl[196] br[196] wl[36] vdd gnd cell_6t
Xbit_r37_c196 bl[196] br[196] wl[37] vdd gnd cell_6t
Xbit_r38_c196 bl[196] br[196] wl[38] vdd gnd cell_6t
Xbit_r39_c196 bl[196] br[196] wl[39] vdd gnd cell_6t
Xbit_r40_c196 bl[196] br[196] wl[40] vdd gnd cell_6t
Xbit_r41_c196 bl[196] br[196] wl[41] vdd gnd cell_6t
Xbit_r42_c196 bl[196] br[196] wl[42] vdd gnd cell_6t
Xbit_r43_c196 bl[196] br[196] wl[43] vdd gnd cell_6t
Xbit_r44_c196 bl[196] br[196] wl[44] vdd gnd cell_6t
Xbit_r45_c196 bl[196] br[196] wl[45] vdd gnd cell_6t
Xbit_r46_c196 bl[196] br[196] wl[46] vdd gnd cell_6t
Xbit_r47_c196 bl[196] br[196] wl[47] vdd gnd cell_6t
Xbit_r48_c196 bl[196] br[196] wl[48] vdd gnd cell_6t
Xbit_r49_c196 bl[196] br[196] wl[49] vdd gnd cell_6t
Xbit_r50_c196 bl[196] br[196] wl[50] vdd gnd cell_6t
Xbit_r51_c196 bl[196] br[196] wl[51] vdd gnd cell_6t
Xbit_r52_c196 bl[196] br[196] wl[52] vdd gnd cell_6t
Xbit_r53_c196 bl[196] br[196] wl[53] vdd gnd cell_6t
Xbit_r54_c196 bl[196] br[196] wl[54] vdd gnd cell_6t
Xbit_r55_c196 bl[196] br[196] wl[55] vdd gnd cell_6t
Xbit_r56_c196 bl[196] br[196] wl[56] vdd gnd cell_6t
Xbit_r57_c196 bl[196] br[196] wl[57] vdd gnd cell_6t
Xbit_r58_c196 bl[196] br[196] wl[58] vdd gnd cell_6t
Xbit_r59_c196 bl[196] br[196] wl[59] vdd gnd cell_6t
Xbit_r60_c196 bl[196] br[196] wl[60] vdd gnd cell_6t
Xbit_r61_c196 bl[196] br[196] wl[61] vdd gnd cell_6t
Xbit_r62_c196 bl[196] br[196] wl[62] vdd gnd cell_6t
Xbit_r63_c196 bl[196] br[196] wl[63] vdd gnd cell_6t
Xbit_r64_c196 bl[196] br[196] wl[64] vdd gnd cell_6t
Xbit_r65_c196 bl[196] br[196] wl[65] vdd gnd cell_6t
Xbit_r66_c196 bl[196] br[196] wl[66] vdd gnd cell_6t
Xbit_r67_c196 bl[196] br[196] wl[67] vdd gnd cell_6t
Xbit_r68_c196 bl[196] br[196] wl[68] vdd gnd cell_6t
Xbit_r69_c196 bl[196] br[196] wl[69] vdd gnd cell_6t
Xbit_r70_c196 bl[196] br[196] wl[70] vdd gnd cell_6t
Xbit_r71_c196 bl[196] br[196] wl[71] vdd gnd cell_6t
Xbit_r72_c196 bl[196] br[196] wl[72] vdd gnd cell_6t
Xbit_r73_c196 bl[196] br[196] wl[73] vdd gnd cell_6t
Xbit_r74_c196 bl[196] br[196] wl[74] vdd gnd cell_6t
Xbit_r75_c196 bl[196] br[196] wl[75] vdd gnd cell_6t
Xbit_r76_c196 bl[196] br[196] wl[76] vdd gnd cell_6t
Xbit_r77_c196 bl[196] br[196] wl[77] vdd gnd cell_6t
Xbit_r78_c196 bl[196] br[196] wl[78] vdd gnd cell_6t
Xbit_r79_c196 bl[196] br[196] wl[79] vdd gnd cell_6t
Xbit_r80_c196 bl[196] br[196] wl[80] vdd gnd cell_6t
Xbit_r81_c196 bl[196] br[196] wl[81] vdd gnd cell_6t
Xbit_r82_c196 bl[196] br[196] wl[82] vdd gnd cell_6t
Xbit_r83_c196 bl[196] br[196] wl[83] vdd gnd cell_6t
Xbit_r84_c196 bl[196] br[196] wl[84] vdd gnd cell_6t
Xbit_r85_c196 bl[196] br[196] wl[85] vdd gnd cell_6t
Xbit_r86_c196 bl[196] br[196] wl[86] vdd gnd cell_6t
Xbit_r87_c196 bl[196] br[196] wl[87] vdd gnd cell_6t
Xbit_r88_c196 bl[196] br[196] wl[88] vdd gnd cell_6t
Xbit_r89_c196 bl[196] br[196] wl[89] vdd gnd cell_6t
Xbit_r90_c196 bl[196] br[196] wl[90] vdd gnd cell_6t
Xbit_r91_c196 bl[196] br[196] wl[91] vdd gnd cell_6t
Xbit_r92_c196 bl[196] br[196] wl[92] vdd gnd cell_6t
Xbit_r93_c196 bl[196] br[196] wl[93] vdd gnd cell_6t
Xbit_r94_c196 bl[196] br[196] wl[94] vdd gnd cell_6t
Xbit_r95_c196 bl[196] br[196] wl[95] vdd gnd cell_6t
Xbit_r96_c196 bl[196] br[196] wl[96] vdd gnd cell_6t
Xbit_r97_c196 bl[196] br[196] wl[97] vdd gnd cell_6t
Xbit_r98_c196 bl[196] br[196] wl[98] vdd gnd cell_6t
Xbit_r99_c196 bl[196] br[196] wl[99] vdd gnd cell_6t
Xbit_r100_c196 bl[196] br[196] wl[100] vdd gnd cell_6t
Xbit_r101_c196 bl[196] br[196] wl[101] vdd gnd cell_6t
Xbit_r102_c196 bl[196] br[196] wl[102] vdd gnd cell_6t
Xbit_r103_c196 bl[196] br[196] wl[103] vdd gnd cell_6t
Xbit_r104_c196 bl[196] br[196] wl[104] vdd gnd cell_6t
Xbit_r105_c196 bl[196] br[196] wl[105] vdd gnd cell_6t
Xbit_r106_c196 bl[196] br[196] wl[106] vdd gnd cell_6t
Xbit_r107_c196 bl[196] br[196] wl[107] vdd gnd cell_6t
Xbit_r108_c196 bl[196] br[196] wl[108] vdd gnd cell_6t
Xbit_r109_c196 bl[196] br[196] wl[109] vdd gnd cell_6t
Xbit_r110_c196 bl[196] br[196] wl[110] vdd gnd cell_6t
Xbit_r111_c196 bl[196] br[196] wl[111] vdd gnd cell_6t
Xbit_r112_c196 bl[196] br[196] wl[112] vdd gnd cell_6t
Xbit_r113_c196 bl[196] br[196] wl[113] vdd gnd cell_6t
Xbit_r114_c196 bl[196] br[196] wl[114] vdd gnd cell_6t
Xbit_r115_c196 bl[196] br[196] wl[115] vdd gnd cell_6t
Xbit_r116_c196 bl[196] br[196] wl[116] vdd gnd cell_6t
Xbit_r117_c196 bl[196] br[196] wl[117] vdd gnd cell_6t
Xbit_r118_c196 bl[196] br[196] wl[118] vdd gnd cell_6t
Xbit_r119_c196 bl[196] br[196] wl[119] vdd gnd cell_6t
Xbit_r120_c196 bl[196] br[196] wl[120] vdd gnd cell_6t
Xbit_r121_c196 bl[196] br[196] wl[121] vdd gnd cell_6t
Xbit_r122_c196 bl[196] br[196] wl[122] vdd gnd cell_6t
Xbit_r123_c196 bl[196] br[196] wl[123] vdd gnd cell_6t
Xbit_r124_c196 bl[196] br[196] wl[124] vdd gnd cell_6t
Xbit_r125_c196 bl[196] br[196] wl[125] vdd gnd cell_6t
Xbit_r126_c196 bl[196] br[196] wl[126] vdd gnd cell_6t
Xbit_r127_c196 bl[196] br[196] wl[127] vdd gnd cell_6t
Xbit_r0_c197 bl[197] br[197] wl[0] vdd gnd cell_6t
Xbit_r1_c197 bl[197] br[197] wl[1] vdd gnd cell_6t
Xbit_r2_c197 bl[197] br[197] wl[2] vdd gnd cell_6t
Xbit_r3_c197 bl[197] br[197] wl[3] vdd gnd cell_6t
Xbit_r4_c197 bl[197] br[197] wl[4] vdd gnd cell_6t
Xbit_r5_c197 bl[197] br[197] wl[5] vdd gnd cell_6t
Xbit_r6_c197 bl[197] br[197] wl[6] vdd gnd cell_6t
Xbit_r7_c197 bl[197] br[197] wl[7] vdd gnd cell_6t
Xbit_r8_c197 bl[197] br[197] wl[8] vdd gnd cell_6t
Xbit_r9_c197 bl[197] br[197] wl[9] vdd gnd cell_6t
Xbit_r10_c197 bl[197] br[197] wl[10] vdd gnd cell_6t
Xbit_r11_c197 bl[197] br[197] wl[11] vdd gnd cell_6t
Xbit_r12_c197 bl[197] br[197] wl[12] vdd gnd cell_6t
Xbit_r13_c197 bl[197] br[197] wl[13] vdd gnd cell_6t
Xbit_r14_c197 bl[197] br[197] wl[14] vdd gnd cell_6t
Xbit_r15_c197 bl[197] br[197] wl[15] vdd gnd cell_6t
Xbit_r16_c197 bl[197] br[197] wl[16] vdd gnd cell_6t
Xbit_r17_c197 bl[197] br[197] wl[17] vdd gnd cell_6t
Xbit_r18_c197 bl[197] br[197] wl[18] vdd gnd cell_6t
Xbit_r19_c197 bl[197] br[197] wl[19] vdd gnd cell_6t
Xbit_r20_c197 bl[197] br[197] wl[20] vdd gnd cell_6t
Xbit_r21_c197 bl[197] br[197] wl[21] vdd gnd cell_6t
Xbit_r22_c197 bl[197] br[197] wl[22] vdd gnd cell_6t
Xbit_r23_c197 bl[197] br[197] wl[23] vdd gnd cell_6t
Xbit_r24_c197 bl[197] br[197] wl[24] vdd gnd cell_6t
Xbit_r25_c197 bl[197] br[197] wl[25] vdd gnd cell_6t
Xbit_r26_c197 bl[197] br[197] wl[26] vdd gnd cell_6t
Xbit_r27_c197 bl[197] br[197] wl[27] vdd gnd cell_6t
Xbit_r28_c197 bl[197] br[197] wl[28] vdd gnd cell_6t
Xbit_r29_c197 bl[197] br[197] wl[29] vdd gnd cell_6t
Xbit_r30_c197 bl[197] br[197] wl[30] vdd gnd cell_6t
Xbit_r31_c197 bl[197] br[197] wl[31] vdd gnd cell_6t
Xbit_r32_c197 bl[197] br[197] wl[32] vdd gnd cell_6t
Xbit_r33_c197 bl[197] br[197] wl[33] vdd gnd cell_6t
Xbit_r34_c197 bl[197] br[197] wl[34] vdd gnd cell_6t
Xbit_r35_c197 bl[197] br[197] wl[35] vdd gnd cell_6t
Xbit_r36_c197 bl[197] br[197] wl[36] vdd gnd cell_6t
Xbit_r37_c197 bl[197] br[197] wl[37] vdd gnd cell_6t
Xbit_r38_c197 bl[197] br[197] wl[38] vdd gnd cell_6t
Xbit_r39_c197 bl[197] br[197] wl[39] vdd gnd cell_6t
Xbit_r40_c197 bl[197] br[197] wl[40] vdd gnd cell_6t
Xbit_r41_c197 bl[197] br[197] wl[41] vdd gnd cell_6t
Xbit_r42_c197 bl[197] br[197] wl[42] vdd gnd cell_6t
Xbit_r43_c197 bl[197] br[197] wl[43] vdd gnd cell_6t
Xbit_r44_c197 bl[197] br[197] wl[44] vdd gnd cell_6t
Xbit_r45_c197 bl[197] br[197] wl[45] vdd gnd cell_6t
Xbit_r46_c197 bl[197] br[197] wl[46] vdd gnd cell_6t
Xbit_r47_c197 bl[197] br[197] wl[47] vdd gnd cell_6t
Xbit_r48_c197 bl[197] br[197] wl[48] vdd gnd cell_6t
Xbit_r49_c197 bl[197] br[197] wl[49] vdd gnd cell_6t
Xbit_r50_c197 bl[197] br[197] wl[50] vdd gnd cell_6t
Xbit_r51_c197 bl[197] br[197] wl[51] vdd gnd cell_6t
Xbit_r52_c197 bl[197] br[197] wl[52] vdd gnd cell_6t
Xbit_r53_c197 bl[197] br[197] wl[53] vdd gnd cell_6t
Xbit_r54_c197 bl[197] br[197] wl[54] vdd gnd cell_6t
Xbit_r55_c197 bl[197] br[197] wl[55] vdd gnd cell_6t
Xbit_r56_c197 bl[197] br[197] wl[56] vdd gnd cell_6t
Xbit_r57_c197 bl[197] br[197] wl[57] vdd gnd cell_6t
Xbit_r58_c197 bl[197] br[197] wl[58] vdd gnd cell_6t
Xbit_r59_c197 bl[197] br[197] wl[59] vdd gnd cell_6t
Xbit_r60_c197 bl[197] br[197] wl[60] vdd gnd cell_6t
Xbit_r61_c197 bl[197] br[197] wl[61] vdd gnd cell_6t
Xbit_r62_c197 bl[197] br[197] wl[62] vdd gnd cell_6t
Xbit_r63_c197 bl[197] br[197] wl[63] vdd gnd cell_6t
Xbit_r64_c197 bl[197] br[197] wl[64] vdd gnd cell_6t
Xbit_r65_c197 bl[197] br[197] wl[65] vdd gnd cell_6t
Xbit_r66_c197 bl[197] br[197] wl[66] vdd gnd cell_6t
Xbit_r67_c197 bl[197] br[197] wl[67] vdd gnd cell_6t
Xbit_r68_c197 bl[197] br[197] wl[68] vdd gnd cell_6t
Xbit_r69_c197 bl[197] br[197] wl[69] vdd gnd cell_6t
Xbit_r70_c197 bl[197] br[197] wl[70] vdd gnd cell_6t
Xbit_r71_c197 bl[197] br[197] wl[71] vdd gnd cell_6t
Xbit_r72_c197 bl[197] br[197] wl[72] vdd gnd cell_6t
Xbit_r73_c197 bl[197] br[197] wl[73] vdd gnd cell_6t
Xbit_r74_c197 bl[197] br[197] wl[74] vdd gnd cell_6t
Xbit_r75_c197 bl[197] br[197] wl[75] vdd gnd cell_6t
Xbit_r76_c197 bl[197] br[197] wl[76] vdd gnd cell_6t
Xbit_r77_c197 bl[197] br[197] wl[77] vdd gnd cell_6t
Xbit_r78_c197 bl[197] br[197] wl[78] vdd gnd cell_6t
Xbit_r79_c197 bl[197] br[197] wl[79] vdd gnd cell_6t
Xbit_r80_c197 bl[197] br[197] wl[80] vdd gnd cell_6t
Xbit_r81_c197 bl[197] br[197] wl[81] vdd gnd cell_6t
Xbit_r82_c197 bl[197] br[197] wl[82] vdd gnd cell_6t
Xbit_r83_c197 bl[197] br[197] wl[83] vdd gnd cell_6t
Xbit_r84_c197 bl[197] br[197] wl[84] vdd gnd cell_6t
Xbit_r85_c197 bl[197] br[197] wl[85] vdd gnd cell_6t
Xbit_r86_c197 bl[197] br[197] wl[86] vdd gnd cell_6t
Xbit_r87_c197 bl[197] br[197] wl[87] vdd gnd cell_6t
Xbit_r88_c197 bl[197] br[197] wl[88] vdd gnd cell_6t
Xbit_r89_c197 bl[197] br[197] wl[89] vdd gnd cell_6t
Xbit_r90_c197 bl[197] br[197] wl[90] vdd gnd cell_6t
Xbit_r91_c197 bl[197] br[197] wl[91] vdd gnd cell_6t
Xbit_r92_c197 bl[197] br[197] wl[92] vdd gnd cell_6t
Xbit_r93_c197 bl[197] br[197] wl[93] vdd gnd cell_6t
Xbit_r94_c197 bl[197] br[197] wl[94] vdd gnd cell_6t
Xbit_r95_c197 bl[197] br[197] wl[95] vdd gnd cell_6t
Xbit_r96_c197 bl[197] br[197] wl[96] vdd gnd cell_6t
Xbit_r97_c197 bl[197] br[197] wl[97] vdd gnd cell_6t
Xbit_r98_c197 bl[197] br[197] wl[98] vdd gnd cell_6t
Xbit_r99_c197 bl[197] br[197] wl[99] vdd gnd cell_6t
Xbit_r100_c197 bl[197] br[197] wl[100] vdd gnd cell_6t
Xbit_r101_c197 bl[197] br[197] wl[101] vdd gnd cell_6t
Xbit_r102_c197 bl[197] br[197] wl[102] vdd gnd cell_6t
Xbit_r103_c197 bl[197] br[197] wl[103] vdd gnd cell_6t
Xbit_r104_c197 bl[197] br[197] wl[104] vdd gnd cell_6t
Xbit_r105_c197 bl[197] br[197] wl[105] vdd gnd cell_6t
Xbit_r106_c197 bl[197] br[197] wl[106] vdd gnd cell_6t
Xbit_r107_c197 bl[197] br[197] wl[107] vdd gnd cell_6t
Xbit_r108_c197 bl[197] br[197] wl[108] vdd gnd cell_6t
Xbit_r109_c197 bl[197] br[197] wl[109] vdd gnd cell_6t
Xbit_r110_c197 bl[197] br[197] wl[110] vdd gnd cell_6t
Xbit_r111_c197 bl[197] br[197] wl[111] vdd gnd cell_6t
Xbit_r112_c197 bl[197] br[197] wl[112] vdd gnd cell_6t
Xbit_r113_c197 bl[197] br[197] wl[113] vdd gnd cell_6t
Xbit_r114_c197 bl[197] br[197] wl[114] vdd gnd cell_6t
Xbit_r115_c197 bl[197] br[197] wl[115] vdd gnd cell_6t
Xbit_r116_c197 bl[197] br[197] wl[116] vdd gnd cell_6t
Xbit_r117_c197 bl[197] br[197] wl[117] vdd gnd cell_6t
Xbit_r118_c197 bl[197] br[197] wl[118] vdd gnd cell_6t
Xbit_r119_c197 bl[197] br[197] wl[119] vdd gnd cell_6t
Xbit_r120_c197 bl[197] br[197] wl[120] vdd gnd cell_6t
Xbit_r121_c197 bl[197] br[197] wl[121] vdd gnd cell_6t
Xbit_r122_c197 bl[197] br[197] wl[122] vdd gnd cell_6t
Xbit_r123_c197 bl[197] br[197] wl[123] vdd gnd cell_6t
Xbit_r124_c197 bl[197] br[197] wl[124] vdd gnd cell_6t
Xbit_r125_c197 bl[197] br[197] wl[125] vdd gnd cell_6t
Xbit_r126_c197 bl[197] br[197] wl[126] vdd gnd cell_6t
Xbit_r127_c197 bl[197] br[197] wl[127] vdd gnd cell_6t
Xbit_r0_c198 bl[198] br[198] wl[0] vdd gnd cell_6t
Xbit_r1_c198 bl[198] br[198] wl[1] vdd gnd cell_6t
Xbit_r2_c198 bl[198] br[198] wl[2] vdd gnd cell_6t
Xbit_r3_c198 bl[198] br[198] wl[3] vdd gnd cell_6t
Xbit_r4_c198 bl[198] br[198] wl[4] vdd gnd cell_6t
Xbit_r5_c198 bl[198] br[198] wl[5] vdd gnd cell_6t
Xbit_r6_c198 bl[198] br[198] wl[6] vdd gnd cell_6t
Xbit_r7_c198 bl[198] br[198] wl[7] vdd gnd cell_6t
Xbit_r8_c198 bl[198] br[198] wl[8] vdd gnd cell_6t
Xbit_r9_c198 bl[198] br[198] wl[9] vdd gnd cell_6t
Xbit_r10_c198 bl[198] br[198] wl[10] vdd gnd cell_6t
Xbit_r11_c198 bl[198] br[198] wl[11] vdd gnd cell_6t
Xbit_r12_c198 bl[198] br[198] wl[12] vdd gnd cell_6t
Xbit_r13_c198 bl[198] br[198] wl[13] vdd gnd cell_6t
Xbit_r14_c198 bl[198] br[198] wl[14] vdd gnd cell_6t
Xbit_r15_c198 bl[198] br[198] wl[15] vdd gnd cell_6t
Xbit_r16_c198 bl[198] br[198] wl[16] vdd gnd cell_6t
Xbit_r17_c198 bl[198] br[198] wl[17] vdd gnd cell_6t
Xbit_r18_c198 bl[198] br[198] wl[18] vdd gnd cell_6t
Xbit_r19_c198 bl[198] br[198] wl[19] vdd gnd cell_6t
Xbit_r20_c198 bl[198] br[198] wl[20] vdd gnd cell_6t
Xbit_r21_c198 bl[198] br[198] wl[21] vdd gnd cell_6t
Xbit_r22_c198 bl[198] br[198] wl[22] vdd gnd cell_6t
Xbit_r23_c198 bl[198] br[198] wl[23] vdd gnd cell_6t
Xbit_r24_c198 bl[198] br[198] wl[24] vdd gnd cell_6t
Xbit_r25_c198 bl[198] br[198] wl[25] vdd gnd cell_6t
Xbit_r26_c198 bl[198] br[198] wl[26] vdd gnd cell_6t
Xbit_r27_c198 bl[198] br[198] wl[27] vdd gnd cell_6t
Xbit_r28_c198 bl[198] br[198] wl[28] vdd gnd cell_6t
Xbit_r29_c198 bl[198] br[198] wl[29] vdd gnd cell_6t
Xbit_r30_c198 bl[198] br[198] wl[30] vdd gnd cell_6t
Xbit_r31_c198 bl[198] br[198] wl[31] vdd gnd cell_6t
Xbit_r32_c198 bl[198] br[198] wl[32] vdd gnd cell_6t
Xbit_r33_c198 bl[198] br[198] wl[33] vdd gnd cell_6t
Xbit_r34_c198 bl[198] br[198] wl[34] vdd gnd cell_6t
Xbit_r35_c198 bl[198] br[198] wl[35] vdd gnd cell_6t
Xbit_r36_c198 bl[198] br[198] wl[36] vdd gnd cell_6t
Xbit_r37_c198 bl[198] br[198] wl[37] vdd gnd cell_6t
Xbit_r38_c198 bl[198] br[198] wl[38] vdd gnd cell_6t
Xbit_r39_c198 bl[198] br[198] wl[39] vdd gnd cell_6t
Xbit_r40_c198 bl[198] br[198] wl[40] vdd gnd cell_6t
Xbit_r41_c198 bl[198] br[198] wl[41] vdd gnd cell_6t
Xbit_r42_c198 bl[198] br[198] wl[42] vdd gnd cell_6t
Xbit_r43_c198 bl[198] br[198] wl[43] vdd gnd cell_6t
Xbit_r44_c198 bl[198] br[198] wl[44] vdd gnd cell_6t
Xbit_r45_c198 bl[198] br[198] wl[45] vdd gnd cell_6t
Xbit_r46_c198 bl[198] br[198] wl[46] vdd gnd cell_6t
Xbit_r47_c198 bl[198] br[198] wl[47] vdd gnd cell_6t
Xbit_r48_c198 bl[198] br[198] wl[48] vdd gnd cell_6t
Xbit_r49_c198 bl[198] br[198] wl[49] vdd gnd cell_6t
Xbit_r50_c198 bl[198] br[198] wl[50] vdd gnd cell_6t
Xbit_r51_c198 bl[198] br[198] wl[51] vdd gnd cell_6t
Xbit_r52_c198 bl[198] br[198] wl[52] vdd gnd cell_6t
Xbit_r53_c198 bl[198] br[198] wl[53] vdd gnd cell_6t
Xbit_r54_c198 bl[198] br[198] wl[54] vdd gnd cell_6t
Xbit_r55_c198 bl[198] br[198] wl[55] vdd gnd cell_6t
Xbit_r56_c198 bl[198] br[198] wl[56] vdd gnd cell_6t
Xbit_r57_c198 bl[198] br[198] wl[57] vdd gnd cell_6t
Xbit_r58_c198 bl[198] br[198] wl[58] vdd gnd cell_6t
Xbit_r59_c198 bl[198] br[198] wl[59] vdd gnd cell_6t
Xbit_r60_c198 bl[198] br[198] wl[60] vdd gnd cell_6t
Xbit_r61_c198 bl[198] br[198] wl[61] vdd gnd cell_6t
Xbit_r62_c198 bl[198] br[198] wl[62] vdd gnd cell_6t
Xbit_r63_c198 bl[198] br[198] wl[63] vdd gnd cell_6t
Xbit_r64_c198 bl[198] br[198] wl[64] vdd gnd cell_6t
Xbit_r65_c198 bl[198] br[198] wl[65] vdd gnd cell_6t
Xbit_r66_c198 bl[198] br[198] wl[66] vdd gnd cell_6t
Xbit_r67_c198 bl[198] br[198] wl[67] vdd gnd cell_6t
Xbit_r68_c198 bl[198] br[198] wl[68] vdd gnd cell_6t
Xbit_r69_c198 bl[198] br[198] wl[69] vdd gnd cell_6t
Xbit_r70_c198 bl[198] br[198] wl[70] vdd gnd cell_6t
Xbit_r71_c198 bl[198] br[198] wl[71] vdd gnd cell_6t
Xbit_r72_c198 bl[198] br[198] wl[72] vdd gnd cell_6t
Xbit_r73_c198 bl[198] br[198] wl[73] vdd gnd cell_6t
Xbit_r74_c198 bl[198] br[198] wl[74] vdd gnd cell_6t
Xbit_r75_c198 bl[198] br[198] wl[75] vdd gnd cell_6t
Xbit_r76_c198 bl[198] br[198] wl[76] vdd gnd cell_6t
Xbit_r77_c198 bl[198] br[198] wl[77] vdd gnd cell_6t
Xbit_r78_c198 bl[198] br[198] wl[78] vdd gnd cell_6t
Xbit_r79_c198 bl[198] br[198] wl[79] vdd gnd cell_6t
Xbit_r80_c198 bl[198] br[198] wl[80] vdd gnd cell_6t
Xbit_r81_c198 bl[198] br[198] wl[81] vdd gnd cell_6t
Xbit_r82_c198 bl[198] br[198] wl[82] vdd gnd cell_6t
Xbit_r83_c198 bl[198] br[198] wl[83] vdd gnd cell_6t
Xbit_r84_c198 bl[198] br[198] wl[84] vdd gnd cell_6t
Xbit_r85_c198 bl[198] br[198] wl[85] vdd gnd cell_6t
Xbit_r86_c198 bl[198] br[198] wl[86] vdd gnd cell_6t
Xbit_r87_c198 bl[198] br[198] wl[87] vdd gnd cell_6t
Xbit_r88_c198 bl[198] br[198] wl[88] vdd gnd cell_6t
Xbit_r89_c198 bl[198] br[198] wl[89] vdd gnd cell_6t
Xbit_r90_c198 bl[198] br[198] wl[90] vdd gnd cell_6t
Xbit_r91_c198 bl[198] br[198] wl[91] vdd gnd cell_6t
Xbit_r92_c198 bl[198] br[198] wl[92] vdd gnd cell_6t
Xbit_r93_c198 bl[198] br[198] wl[93] vdd gnd cell_6t
Xbit_r94_c198 bl[198] br[198] wl[94] vdd gnd cell_6t
Xbit_r95_c198 bl[198] br[198] wl[95] vdd gnd cell_6t
Xbit_r96_c198 bl[198] br[198] wl[96] vdd gnd cell_6t
Xbit_r97_c198 bl[198] br[198] wl[97] vdd gnd cell_6t
Xbit_r98_c198 bl[198] br[198] wl[98] vdd gnd cell_6t
Xbit_r99_c198 bl[198] br[198] wl[99] vdd gnd cell_6t
Xbit_r100_c198 bl[198] br[198] wl[100] vdd gnd cell_6t
Xbit_r101_c198 bl[198] br[198] wl[101] vdd gnd cell_6t
Xbit_r102_c198 bl[198] br[198] wl[102] vdd gnd cell_6t
Xbit_r103_c198 bl[198] br[198] wl[103] vdd gnd cell_6t
Xbit_r104_c198 bl[198] br[198] wl[104] vdd gnd cell_6t
Xbit_r105_c198 bl[198] br[198] wl[105] vdd gnd cell_6t
Xbit_r106_c198 bl[198] br[198] wl[106] vdd gnd cell_6t
Xbit_r107_c198 bl[198] br[198] wl[107] vdd gnd cell_6t
Xbit_r108_c198 bl[198] br[198] wl[108] vdd gnd cell_6t
Xbit_r109_c198 bl[198] br[198] wl[109] vdd gnd cell_6t
Xbit_r110_c198 bl[198] br[198] wl[110] vdd gnd cell_6t
Xbit_r111_c198 bl[198] br[198] wl[111] vdd gnd cell_6t
Xbit_r112_c198 bl[198] br[198] wl[112] vdd gnd cell_6t
Xbit_r113_c198 bl[198] br[198] wl[113] vdd gnd cell_6t
Xbit_r114_c198 bl[198] br[198] wl[114] vdd gnd cell_6t
Xbit_r115_c198 bl[198] br[198] wl[115] vdd gnd cell_6t
Xbit_r116_c198 bl[198] br[198] wl[116] vdd gnd cell_6t
Xbit_r117_c198 bl[198] br[198] wl[117] vdd gnd cell_6t
Xbit_r118_c198 bl[198] br[198] wl[118] vdd gnd cell_6t
Xbit_r119_c198 bl[198] br[198] wl[119] vdd gnd cell_6t
Xbit_r120_c198 bl[198] br[198] wl[120] vdd gnd cell_6t
Xbit_r121_c198 bl[198] br[198] wl[121] vdd gnd cell_6t
Xbit_r122_c198 bl[198] br[198] wl[122] vdd gnd cell_6t
Xbit_r123_c198 bl[198] br[198] wl[123] vdd gnd cell_6t
Xbit_r124_c198 bl[198] br[198] wl[124] vdd gnd cell_6t
Xbit_r125_c198 bl[198] br[198] wl[125] vdd gnd cell_6t
Xbit_r126_c198 bl[198] br[198] wl[126] vdd gnd cell_6t
Xbit_r127_c198 bl[198] br[198] wl[127] vdd gnd cell_6t
Xbit_r0_c199 bl[199] br[199] wl[0] vdd gnd cell_6t
Xbit_r1_c199 bl[199] br[199] wl[1] vdd gnd cell_6t
Xbit_r2_c199 bl[199] br[199] wl[2] vdd gnd cell_6t
Xbit_r3_c199 bl[199] br[199] wl[3] vdd gnd cell_6t
Xbit_r4_c199 bl[199] br[199] wl[4] vdd gnd cell_6t
Xbit_r5_c199 bl[199] br[199] wl[5] vdd gnd cell_6t
Xbit_r6_c199 bl[199] br[199] wl[6] vdd gnd cell_6t
Xbit_r7_c199 bl[199] br[199] wl[7] vdd gnd cell_6t
Xbit_r8_c199 bl[199] br[199] wl[8] vdd gnd cell_6t
Xbit_r9_c199 bl[199] br[199] wl[9] vdd gnd cell_6t
Xbit_r10_c199 bl[199] br[199] wl[10] vdd gnd cell_6t
Xbit_r11_c199 bl[199] br[199] wl[11] vdd gnd cell_6t
Xbit_r12_c199 bl[199] br[199] wl[12] vdd gnd cell_6t
Xbit_r13_c199 bl[199] br[199] wl[13] vdd gnd cell_6t
Xbit_r14_c199 bl[199] br[199] wl[14] vdd gnd cell_6t
Xbit_r15_c199 bl[199] br[199] wl[15] vdd gnd cell_6t
Xbit_r16_c199 bl[199] br[199] wl[16] vdd gnd cell_6t
Xbit_r17_c199 bl[199] br[199] wl[17] vdd gnd cell_6t
Xbit_r18_c199 bl[199] br[199] wl[18] vdd gnd cell_6t
Xbit_r19_c199 bl[199] br[199] wl[19] vdd gnd cell_6t
Xbit_r20_c199 bl[199] br[199] wl[20] vdd gnd cell_6t
Xbit_r21_c199 bl[199] br[199] wl[21] vdd gnd cell_6t
Xbit_r22_c199 bl[199] br[199] wl[22] vdd gnd cell_6t
Xbit_r23_c199 bl[199] br[199] wl[23] vdd gnd cell_6t
Xbit_r24_c199 bl[199] br[199] wl[24] vdd gnd cell_6t
Xbit_r25_c199 bl[199] br[199] wl[25] vdd gnd cell_6t
Xbit_r26_c199 bl[199] br[199] wl[26] vdd gnd cell_6t
Xbit_r27_c199 bl[199] br[199] wl[27] vdd gnd cell_6t
Xbit_r28_c199 bl[199] br[199] wl[28] vdd gnd cell_6t
Xbit_r29_c199 bl[199] br[199] wl[29] vdd gnd cell_6t
Xbit_r30_c199 bl[199] br[199] wl[30] vdd gnd cell_6t
Xbit_r31_c199 bl[199] br[199] wl[31] vdd gnd cell_6t
Xbit_r32_c199 bl[199] br[199] wl[32] vdd gnd cell_6t
Xbit_r33_c199 bl[199] br[199] wl[33] vdd gnd cell_6t
Xbit_r34_c199 bl[199] br[199] wl[34] vdd gnd cell_6t
Xbit_r35_c199 bl[199] br[199] wl[35] vdd gnd cell_6t
Xbit_r36_c199 bl[199] br[199] wl[36] vdd gnd cell_6t
Xbit_r37_c199 bl[199] br[199] wl[37] vdd gnd cell_6t
Xbit_r38_c199 bl[199] br[199] wl[38] vdd gnd cell_6t
Xbit_r39_c199 bl[199] br[199] wl[39] vdd gnd cell_6t
Xbit_r40_c199 bl[199] br[199] wl[40] vdd gnd cell_6t
Xbit_r41_c199 bl[199] br[199] wl[41] vdd gnd cell_6t
Xbit_r42_c199 bl[199] br[199] wl[42] vdd gnd cell_6t
Xbit_r43_c199 bl[199] br[199] wl[43] vdd gnd cell_6t
Xbit_r44_c199 bl[199] br[199] wl[44] vdd gnd cell_6t
Xbit_r45_c199 bl[199] br[199] wl[45] vdd gnd cell_6t
Xbit_r46_c199 bl[199] br[199] wl[46] vdd gnd cell_6t
Xbit_r47_c199 bl[199] br[199] wl[47] vdd gnd cell_6t
Xbit_r48_c199 bl[199] br[199] wl[48] vdd gnd cell_6t
Xbit_r49_c199 bl[199] br[199] wl[49] vdd gnd cell_6t
Xbit_r50_c199 bl[199] br[199] wl[50] vdd gnd cell_6t
Xbit_r51_c199 bl[199] br[199] wl[51] vdd gnd cell_6t
Xbit_r52_c199 bl[199] br[199] wl[52] vdd gnd cell_6t
Xbit_r53_c199 bl[199] br[199] wl[53] vdd gnd cell_6t
Xbit_r54_c199 bl[199] br[199] wl[54] vdd gnd cell_6t
Xbit_r55_c199 bl[199] br[199] wl[55] vdd gnd cell_6t
Xbit_r56_c199 bl[199] br[199] wl[56] vdd gnd cell_6t
Xbit_r57_c199 bl[199] br[199] wl[57] vdd gnd cell_6t
Xbit_r58_c199 bl[199] br[199] wl[58] vdd gnd cell_6t
Xbit_r59_c199 bl[199] br[199] wl[59] vdd gnd cell_6t
Xbit_r60_c199 bl[199] br[199] wl[60] vdd gnd cell_6t
Xbit_r61_c199 bl[199] br[199] wl[61] vdd gnd cell_6t
Xbit_r62_c199 bl[199] br[199] wl[62] vdd gnd cell_6t
Xbit_r63_c199 bl[199] br[199] wl[63] vdd gnd cell_6t
Xbit_r64_c199 bl[199] br[199] wl[64] vdd gnd cell_6t
Xbit_r65_c199 bl[199] br[199] wl[65] vdd gnd cell_6t
Xbit_r66_c199 bl[199] br[199] wl[66] vdd gnd cell_6t
Xbit_r67_c199 bl[199] br[199] wl[67] vdd gnd cell_6t
Xbit_r68_c199 bl[199] br[199] wl[68] vdd gnd cell_6t
Xbit_r69_c199 bl[199] br[199] wl[69] vdd gnd cell_6t
Xbit_r70_c199 bl[199] br[199] wl[70] vdd gnd cell_6t
Xbit_r71_c199 bl[199] br[199] wl[71] vdd gnd cell_6t
Xbit_r72_c199 bl[199] br[199] wl[72] vdd gnd cell_6t
Xbit_r73_c199 bl[199] br[199] wl[73] vdd gnd cell_6t
Xbit_r74_c199 bl[199] br[199] wl[74] vdd gnd cell_6t
Xbit_r75_c199 bl[199] br[199] wl[75] vdd gnd cell_6t
Xbit_r76_c199 bl[199] br[199] wl[76] vdd gnd cell_6t
Xbit_r77_c199 bl[199] br[199] wl[77] vdd gnd cell_6t
Xbit_r78_c199 bl[199] br[199] wl[78] vdd gnd cell_6t
Xbit_r79_c199 bl[199] br[199] wl[79] vdd gnd cell_6t
Xbit_r80_c199 bl[199] br[199] wl[80] vdd gnd cell_6t
Xbit_r81_c199 bl[199] br[199] wl[81] vdd gnd cell_6t
Xbit_r82_c199 bl[199] br[199] wl[82] vdd gnd cell_6t
Xbit_r83_c199 bl[199] br[199] wl[83] vdd gnd cell_6t
Xbit_r84_c199 bl[199] br[199] wl[84] vdd gnd cell_6t
Xbit_r85_c199 bl[199] br[199] wl[85] vdd gnd cell_6t
Xbit_r86_c199 bl[199] br[199] wl[86] vdd gnd cell_6t
Xbit_r87_c199 bl[199] br[199] wl[87] vdd gnd cell_6t
Xbit_r88_c199 bl[199] br[199] wl[88] vdd gnd cell_6t
Xbit_r89_c199 bl[199] br[199] wl[89] vdd gnd cell_6t
Xbit_r90_c199 bl[199] br[199] wl[90] vdd gnd cell_6t
Xbit_r91_c199 bl[199] br[199] wl[91] vdd gnd cell_6t
Xbit_r92_c199 bl[199] br[199] wl[92] vdd gnd cell_6t
Xbit_r93_c199 bl[199] br[199] wl[93] vdd gnd cell_6t
Xbit_r94_c199 bl[199] br[199] wl[94] vdd gnd cell_6t
Xbit_r95_c199 bl[199] br[199] wl[95] vdd gnd cell_6t
Xbit_r96_c199 bl[199] br[199] wl[96] vdd gnd cell_6t
Xbit_r97_c199 bl[199] br[199] wl[97] vdd gnd cell_6t
Xbit_r98_c199 bl[199] br[199] wl[98] vdd gnd cell_6t
Xbit_r99_c199 bl[199] br[199] wl[99] vdd gnd cell_6t
Xbit_r100_c199 bl[199] br[199] wl[100] vdd gnd cell_6t
Xbit_r101_c199 bl[199] br[199] wl[101] vdd gnd cell_6t
Xbit_r102_c199 bl[199] br[199] wl[102] vdd gnd cell_6t
Xbit_r103_c199 bl[199] br[199] wl[103] vdd gnd cell_6t
Xbit_r104_c199 bl[199] br[199] wl[104] vdd gnd cell_6t
Xbit_r105_c199 bl[199] br[199] wl[105] vdd gnd cell_6t
Xbit_r106_c199 bl[199] br[199] wl[106] vdd gnd cell_6t
Xbit_r107_c199 bl[199] br[199] wl[107] vdd gnd cell_6t
Xbit_r108_c199 bl[199] br[199] wl[108] vdd gnd cell_6t
Xbit_r109_c199 bl[199] br[199] wl[109] vdd gnd cell_6t
Xbit_r110_c199 bl[199] br[199] wl[110] vdd gnd cell_6t
Xbit_r111_c199 bl[199] br[199] wl[111] vdd gnd cell_6t
Xbit_r112_c199 bl[199] br[199] wl[112] vdd gnd cell_6t
Xbit_r113_c199 bl[199] br[199] wl[113] vdd gnd cell_6t
Xbit_r114_c199 bl[199] br[199] wl[114] vdd gnd cell_6t
Xbit_r115_c199 bl[199] br[199] wl[115] vdd gnd cell_6t
Xbit_r116_c199 bl[199] br[199] wl[116] vdd gnd cell_6t
Xbit_r117_c199 bl[199] br[199] wl[117] vdd gnd cell_6t
Xbit_r118_c199 bl[199] br[199] wl[118] vdd gnd cell_6t
Xbit_r119_c199 bl[199] br[199] wl[119] vdd gnd cell_6t
Xbit_r120_c199 bl[199] br[199] wl[120] vdd gnd cell_6t
Xbit_r121_c199 bl[199] br[199] wl[121] vdd gnd cell_6t
Xbit_r122_c199 bl[199] br[199] wl[122] vdd gnd cell_6t
Xbit_r123_c199 bl[199] br[199] wl[123] vdd gnd cell_6t
Xbit_r124_c199 bl[199] br[199] wl[124] vdd gnd cell_6t
Xbit_r125_c199 bl[199] br[199] wl[125] vdd gnd cell_6t
Xbit_r126_c199 bl[199] br[199] wl[126] vdd gnd cell_6t
Xbit_r127_c199 bl[199] br[199] wl[127] vdd gnd cell_6t
Xbit_r0_c200 bl[200] br[200] wl[0] vdd gnd cell_6t
Xbit_r1_c200 bl[200] br[200] wl[1] vdd gnd cell_6t
Xbit_r2_c200 bl[200] br[200] wl[2] vdd gnd cell_6t
Xbit_r3_c200 bl[200] br[200] wl[3] vdd gnd cell_6t
Xbit_r4_c200 bl[200] br[200] wl[4] vdd gnd cell_6t
Xbit_r5_c200 bl[200] br[200] wl[5] vdd gnd cell_6t
Xbit_r6_c200 bl[200] br[200] wl[6] vdd gnd cell_6t
Xbit_r7_c200 bl[200] br[200] wl[7] vdd gnd cell_6t
Xbit_r8_c200 bl[200] br[200] wl[8] vdd gnd cell_6t
Xbit_r9_c200 bl[200] br[200] wl[9] vdd gnd cell_6t
Xbit_r10_c200 bl[200] br[200] wl[10] vdd gnd cell_6t
Xbit_r11_c200 bl[200] br[200] wl[11] vdd gnd cell_6t
Xbit_r12_c200 bl[200] br[200] wl[12] vdd gnd cell_6t
Xbit_r13_c200 bl[200] br[200] wl[13] vdd gnd cell_6t
Xbit_r14_c200 bl[200] br[200] wl[14] vdd gnd cell_6t
Xbit_r15_c200 bl[200] br[200] wl[15] vdd gnd cell_6t
Xbit_r16_c200 bl[200] br[200] wl[16] vdd gnd cell_6t
Xbit_r17_c200 bl[200] br[200] wl[17] vdd gnd cell_6t
Xbit_r18_c200 bl[200] br[200] wl[18] vdd gnd cell_6t
Xbit_r19_c200 bl[200] br[200] wl[19] vdd gnd cell_6t
Xbit_r20_c200 bl[200] br[200] wl[20] vdd gnd cell_6t
Xbit_r21_c200 bl[200] br[200] wl[21] vdd gnd cell_6t
Xbit_r22_c200 bl[200] br[200] wl[22] vdd gnd cell_6t
Xbit_r23_c200 bl[200] br[200] wl[23] vdd gnd cell_6t
Xbit_r24_c200 bl[200] br[200] wl[24] vdd gnd cell_6t
Xbit_r25_c200 bl[200] br[200] wl[25] vdd gnd cell_6t
Xbit_r26_c200 bl[200] br[200] wl[26] vdd gnd cell_6t
Xbit_r27_c200 bl[200] br[200] wl[27] vdd gnd cell_6t
Xbit_r28_c200 bl[200] br[200] wl[28] vdd gnd cell_6t
Xbit_r29_c200 bl[200] br[200] wl[29] vdd gnd cell_6t
Xbit_r30_c200 bl[200] br[200] wl[30] vdd gnd cell_6t
Xbit_r31_c200 bl[200] br[200] wl[31] vdd gnd cell_6t
Xbit_r32_c200 bl[200] br[200] wl[32] vdd gnd cell_6t
Xbit_r33_c200 bl[200] br[200] wl[33] vdd gnd cell_6t
Xbit_r34_c200 bl[200] br[200] wl[34] vdd gnd cell_6t
Xbit_r35_c200 bl[200] br[200] wl[35] vdd gnd cell_6t
Xbit_r36_c200 bl[200] br[200] wl[36] vdd gnd cell_6t
Xbit_r37_c200 bl[200] br[200] wl[37] vdd gnd cell_6t
Xbit_r38_c200 bl[200] br[200] wl[38] vdd gnd cell_6t
Xbit_r39_c200 bl[200] br[200] wl[39] vdd gnd cell_6t
Xbit_r40_c200 bl[200] br[200] wl[40] vdd gnd cell_6t
Xbit_r41_c200 bl[200] br[200] wl[41] vdd gnd cell_6t
Xbit_r42_c200 bl[200] br[200] wl[42] vdd gnd cell_6t
Xbit_r43_c200 bl[200] br[200] wl[43] vdd gnd cell_6t
Xbit_r44_c200 bl[200] br[200] wl[44] vdd gnd cell_6t
Xbit_r45_c200 bl[200] br[200] wl[45] vdd gnd cell_6t
Xbit_r46_c200 bl[200] br[200] wl[46] vdd gnd cell_6t
Xbit_r47_c200 bl[200] br[200] wl[47] vdd gnd cell_6t
Xbit_r48_c200 bl[200] br[200] wl[48] vdd gnd cell_6t
Xbit_r49_c200 bl[200] br[200] wl[49] vdd gnd cell_6t
Xbit_r50_c200 bl[200] br[200] wl[50] vdd gnd cell_6t
Xbit_r51_c200 bl[200] br[200] wl[51] vdd gnd cell_6t
Xbit_r52_c200 bl[200] br[200] wl[52] vdd gnd cell_6t
Xbit_r53_c200 bl[200] br[200] wl[53] vdd gnd cell_6t
Xbit_r54_c200 bl[200] br[200] wl[54] vdd gnd cell_6t
Xbit_r55_c200 bl[200] br[200] wl[55] vdd gnd cell_6t
Xbit_r56_c200 bl[200] br[200] wl[56] vdd gnd cell_6t
Xbit_r57_c200 bl[200] br[200] wl[57] vdd gnd cell_6t
Xbit_r58_c200 bl[200] br[200] wl[58] vdd gnd cell_6t
Xbit_r59_c200 bl[200] br[200] wl[59] vdd gnd cell_6t
Xbit_r60_c200 bl[200] br[200] wl[60] vdd gnd cell_6t
Xbit_r61_c200 bl[200] br[200] wl[61] vdd gnd cell_6t
Xbit_r62_c200 bl[200] br[200] wl[62] vdd gnd cell_6t
Xbit_r63_c200 bl[200] br[200] wl[63] vdd gnd cell_6t
Xbit_r64_c200 bl[200] br[200] wl[64] vdd gnd cell_6t
Xbit_r65_c200 bl[200] br[200] wl[65] vdd gnd cell_6t
Xbit_r66_c200 bl[200] br[200] wl[66] vdd gnd cell_6t
Xbit_r67_c200 bl[200] br[200] wl[67] vdd gnd cell_6t
Xbit_r68_c200 bl[200] br[200] wl[68] vdd gnd cell_6t
Xbit_r69_c200 bl[200] br[200] wl[69] vdd gnd cell_6t
Xbit_r70_c200 bl[200] br[200] wl[70] vdd gnd cell_6t
Xbit_r71_c200 bl[200] br[200] wl[71] vdd gnd cell_6t
Xbit_r72_c200 bl[200] br[200] wl[72] vdd gnd cell_6t
Xbit_r73_c200 bl[200] br[200] wl[73] vdd gnd cell_6t
Xbit_r74_c200 bl[200] br[200] wl[74] vdd gnd cell_6t
Xbit_r75_c200 bl[200] br[200] wl[75] vdd gnd cell_6t
Xbit_r76_c200 bl[200] br[200] wl[76] vdd gnd cell_6t
Xbit_r77_c200 bl[200] br[200] wl[77] vdd gnd cell_6t
Xbit_r78_c200 bl[200] br[200] wl[78] vdd gnd cell_6t
Xbit_r79_c200 bl[200] br[200] wl[79] vdd gnd cell_6t
Xbit_r80_c200 bl[200] br[200] wl[80] vdd gnd cell_6t
Xbit_r81_c200 bl[200] br[200] wl[81] vdd gnd cell_6t
Xbit_r82_c200 bl[200] br[200] wl[82] vdd gnd cell_6t
Xbit_r83_c200 bl[200] br[200] wl[83] vdd gnd cell_6t
Xbit_r84_c200 bl[200] br[200] wl[84] vdd gnd cell_6t
Xbit_r85_c200 bl[200] br[200] wl[85] vdd gnd cell_6t
Xbit_r86_c200 bl[200] br[200] wl[86] vdd gnd cell_6t
Xbit_r87_c200 bl[200] br[200] wl[87] vdd gnd cell_6t
Xbit_r88_c200 bl[200] br[200] wl[88] vdd gnd cell_6t
Xbit_r89_c200 bl[200] br[200] wl[89] vdd gnd cell_6t
Xbit_r90_c200 bl[200] br[200] wl[90] vdd gnd cell_6t
Xbit_r91_c200 bl[200] br[200] wl[91] vdd gnd cell_6t
Xbit_r92_c200 bl[200] br[200] wl[92] vdd gnd cell_6t
Xbit_r93_c200 bl[200] br[200] wl[93] vdd gnd cell_6t
Xbit_r94_c200 bl[200] br[200] wl[94] vdd gnd cell_6t
Xbit_r95_c200 bl[200] br[200] wl[95] vdd gnd cell_6t
Xbit_r96_c200 bl[200] br[200] wl[96] vdd gnd cell_6t
Xbit_r97_c200 bl[200] br[200] wl[97] vdd gnd cell_6t
Xbit_r98_c200 bl[200] br[200] wl[98] vdd gnd cell_6t
Xbit_r99_c200 bl[200] br[200] wl[99] vdd gnd cell_6t
Xbit_r100_c200 bl[200] br[200] wl[100] vdd gnd cell_6t
Xbit_r101_c200 bl[200] br[200] wl[101] vdd gnd cell_6t
Xbit_r102_c200 bl[200] br[200] wl[102] vdd gnd cell_6t
Xbit_r103_c200 bl[200] br[200] wl[103] vdd gnd cell_6t
Xbit_r104_c200 bl[200] br[200] wl[104] vdd gnd cell_6t
Xbit_r105_c200 bl[200] br[200] wl[105] vdd gnd cell_6t
Xbit_r106_c200 bl[200] br[200] wl[106] vdd gnd cell_6t
Xbit_r107_c200 bl[200] br[200] wl[107] vdd gnd cell_6t
Xbit_r108_c200 bl[200] br[200] wl[108] vdd gnd cell_6t
Xbit_r109_c200 bl[200] br[200] wl[109] vdd gnd cell_6t
Xbit_r110_c200 bl[200] br[200] wl[110] vdd gnd cell_6t
Xbit_r111_c200 bl[200] br[200] wl[111] vdd gnd cell_6t
Xbit_r112_c200 bl[200] br[200] wl[112] vdd gnd cell_6t
Xbit_r113_c200 bl[200] br[200] wl[113] vdd gnd cell_6t
Xbit_r114_c200 bl[200] br[200] wl[114] vdd gnd cell_6t
Xbit_r115_c200 bl[200] br[200] wl[115] vdd gnd cell_6t
Xbit_r116_c200 bl[200] br[200] wl[116] vdd gnd cell_6t
Xbit_r117_c200 bl[200] br[200] wl[117] vdd gnd cell_6t
Xbit_r118_c200 bl[200] br[200] wl[118] vdd gnd cell_6t
Xbit_r119_c200 bl[200] br[200] wl[119] vdd gnd cell_6t
Xbit_r120_c200 bl[200] br[200] wl[120] vdd gnd cell_6t
Xbit_r121_c200 bl[200] br[200] wl[121] vdd gnd cell_6t
Xbit_r122_c200 bl[200] br[200] wl[122] vdd gnd cell_6t
Xbit_r123_c200 bl[200] br[200] wl[123] vdd gnd cell_6t
Xbit_r124_c200 bl[200] br[200] wl[124] vdd gnd cell_6t
Xbit_r125_c200 bl[200] br[200] wl[125] vdd gnd cell_6t
Xbit_r126_c200 bl[200] br[200] wl[126] vdd gnd cell_6t
Xbit_r127_c200 bl[200] br[200] wl[127] vdd gnd cell_6t
Xbit_r0_c201 bl[201] br[201] wl[0] vdd gnd cell_6t
Xbit_r1_c201 bl[201] br[201] wl[1] vdd gnd cell_6t
Xbit_r2_c201 bl[201] br[201] wl[2] vdd gnd cell_6t
Xbit_r3_c201 bl[201] br[201] wl[3] vdd gnd cell_6t
Xbit_r4_c201 bl[201] br[201] wl[4] vdd gnd cell_6t
Xbit_r5_c201 bl[201] br[201] wl[5] vdd gnd cell_6t
Xbit_r6_c201 bl[201] br[201] wl[6] vdd gnd cell_6t
Xbit_r7_c201 bl[201] br[201] wl[7] vdd gnd cell_6t
Xbit_r8_c201 bl[201] br[201] wl[8] vdd gnd cell_6t
Xbit_r9_c201 bl[201] br[201] wl[9] vdd gnd cell_6t
Xbit_r10_c201 bl[201] br[201] wl[10] vdd gnd cell_6t
Xbit_r11_c201 bl[201] br[201] wl[11] vdd gnd cell_6t
Xbit_r12_c201 bl[201] br[201] wl[12] vdd gnd cell_6t
Xbit_r13_c201 bl[201] br[201] wl[13] vdd gnd cell_6t
Xbit_r14_c201 bl[201] br[201] wl[14] vdd gnd cell_6t
Xbit_r15_c201 bl[201] br[201] wl[15] vdd gnd cell_6t
Xbit_r16_c201 bl[201] br[201] wl[16] vdd gnd cell_6t
Xbit_r17_c201 bl[201] br[201] wl[17] vdd gnd cell_6t
Xbit_r18_c201 bl[201] br[201] wl[18] vdd gnd cell_6t
Xbit_r19_c201 bl[201] br[201] wl[19] vdd gnd cell_6t
Xbit_r20_c201 bl[201] br[201] wl[20] vdd gnd cell_6t
Xbit_r21_c201 bl[201] br[201] wl[21] vdd gnd cell_6t
Xbit_r22_c201 bl[201] br[201] wl[22] vdd gnd cell_6t
Xbit_r23_c201 bl[201] br[201] wl[23] vdd gnd cell_6t
Xbit_r24_c201 bl[201] br[201] wl[24] vdd gnd cell_6t
Xbit_r25_c201 bl[201] br[201] wl[25] vdd gnd cell_6t
Xbit_r26_c201 bl[201] br[201] wl[26] vdd gnd cell_6t
Xbit_r27_c201 bl[201] br[201] wl[27] vdd gnd cell_6t
Xbit_r28_c201 bl[201] br[201] wl[28] vdd gnd cell_6t
Xbit_r29_c201 bl[201] br[201] wl[29] vdd gnd cell_6t
Xbit_r30_c201 bl[201] br[201] wl[30] vdd gnd cell_6t
Xbit_r31_c201 bl[201] br[201] wl[31] vdd gnd cell_6t
Xbit_r32_c201 bl[201] br[201] wl[32] vdd gnd cell_6t
Xbit_r33_c201 bl[201] br[201] wl[33] vdd gnd cell_6t
Xbit_r34_c201 bl[201] br[201] wl[34] vdd gnd cell_6t
Xbit_r35_c201 bl[201] br[201] wl[35] vdd gnd cell_6t
Xbit_r36_c201 bl[201] br[201] wl[36] vdd gnd cell_6t
Xbit_r37_c201 bl[201] br[201] wl[37] vdd gnd cell_6t
Xbit_r38_c201 bl[201] br[201] wl[38] vdd gnd cell_6t
Xbit_r39_c201 bl[201] br[201] wl[39] vdd gnd cell_6t
Xbit_r40_c201 bl[201] br[201] wl[40] vdd gnd cell_6t
Xbit_r41_c201 bl[201] br[201] wl[41] vdd gnd cell_6t
Xbit_r42_c201 bl[201] br[201] wl[42] vdd gnd cell_6t
Xbit_r43_c201 bl[201] br[201] wl[43] vdd gnd cell_6t
Xbit_r44_c201 bl[201] br[201] wl[44] vdd gnd cell_6t
Xbit_r45_c201 bl[201] br[201] wl[45] vdd gnd cell_6t
Xbit_r46_c201 bl[201] br[201] wl[46] vdd gnd cell_6t
Xbit_r47_c201 bl[201] br[201] wl[47] vdd gnd cell_6t
Xbit_r48_c201 bl[201] br[201] wl[48] vdd gnd cell_6t
Xbit_r49_c201 bl[201] br[201] wl[49] vdd gnd cell_6t
Xbit_r50_c201 bl[201] br[201] wl[50] vdd gnd cell_6t
Xbit_r51_c201 bl[201] br[201] wl[51] vdd gnd cell_6t
Xbit_r52_c201 bl[201] br[201] wl[52] vdd gnd cell_6t
Xbit_r53_c201 bl[201] br[201] wl[53] vdd gnd cell_6t
Xbit_r54_c201 bl[201] br[201] wl[54] vdd gnd cell_6t
Xbit_r55_c201 bl[201] br[201] wl[55] vdd gnd cell_6t
Xbit_r56_c201 bl[201] br[201] wl[56] vdd gnd cell_6t
Xbit_r57_c201 bl[201] br[201] wl[57] vdd gnd cell_6t
Xbit_r58_c201 bl[201] br[201] wl[58] vdd gnd cell_6t
Xbit_r59_c201 bl[201] br[201] wl[59] vdd gnd cell_6t
Xbit_r60_c201 bl[201] br[201] wl[60] vdd gnd cell_6t
Xbit_r61_c201 bl[201] br[201] wl[61] vdd gnd cell_6t
Xbit_r62_c201 bl[201] br[201] wl[62] vdd gnd cell_6t
Xbit_r63_c201 bl[201] br[201] wl[63] vdd gnd cell_6t
Xbit_r64_c201 bl[201] br[201] wl[64] vdd gnd cell_6t
Xbit_r65_c201 bl[201] br[201] wl[65] vdd gnd cell_6t
Xbit_r66_c201 bl[201] br[201] wl[66] vdd gnd cell_6t
Xbit_r67_c201 bl[201] br[201] wl[67] vdd gnd cell_6t
Xbit_r68_c201 bl[201] br[201] wl[68] vdd gnd cell_6t
Xbit_r69_c201 bl[201] br[201] wl[69] vdd gnd cell_6t
Xbit_r70_c201 bl[201] br[201] wl[70] vdd gnd cell_6t
Xbit_r71_c201 bl[201] br[201] wl[71] vdd gnd cell_6t
Xbit_r72_c201 bl[201] br[201] wl[72] vdd gnd cell_6t
Xbit_r73_c201 bl[201] br[201] wl[73] vdd gnd cell_6t
Xbit_r74_c201 bl[201] br[201] wl[74] vdd gnd cell_6t
Xbit_r75_c201 bl[201] br[201] wl[75] vdd gnd cell_6t
Xbit_r76_c201 bl[201] br[201] wl[76] vdd gnd cell_6t
Xbit_r77_c201 bl[201] br[201] wl[77] vdd gnd cell_6t
Xbit_r78_c201 bl[201] br[201] wl[78] vdd gnd cell_6t
Xbit_r79_c201 bl[201] br[201] wl[79] vdd gnd cell_6t
Xbit_r80_c201 bl[201] br[201] wl[80] vdd gnd cell_6t
Xbit_r81_c201 bl[201] br[201] wl[81] vdd gnd cell_6t
Xbit_r82_c201 bl[201] br[201] wl[82] vdd gnd cell_6t
Xbit_r83_c201 bl[201] br[201] wl[83] vdd gnd cell_6t
Xbit_r84_c201 bl[201] br[201] wl[84] vdd gnd cell_6t
Xbit_r85_c201 bl[201] br[201] wl[85] vdd gnd cell_6t
Xbit_r86_c201 bl[201] br[201] wl[86] vdd gnd cell_6t
Xbit_r87_c201 bl[201] br[201] wl[87] vdd gnd cell_6t
Xbit_r88_c201 bl[201] br[201] wl[88] vdd gnd cell_6t
Xbit_r89_c201 bl[201] br[201] wl[89] vdd gnd cell_6t
Xbit_r90_c201 bl[201] br[201] wl[90] vdd gnd cell_6t
Xbit_r91_c201 bl[201] br[201] wl[91] vdd gnd cell_6t
Xbit_r92_c201 bl[201] br[201] wl[92] vdd gnd cell_6t
Xbit_r93_c201 bl[201] br[201] wl[93] vdd gnd cell_6t
Xbit_r94_c201 bl[201] br[201] wl[94] vdd gnd cell_6t
Xbit_r95_c201 bl[201] br[201] wl[95] vdd gnd cell_6t
Xbit_r96_c201 bl[201] br[201] wl[96] vdd gnd cell_6t
Xbit_r97_c201 bl[201] br[201] wl[97] vdd gnd cell_6t
Xbit_r98_c201 bl[201] br[201] wl[98] vdd gnd cell_6t
Xbit_r99_c201 bl[201] br[201] wl[99] vdd gnd cell_6t
Xbit_r100_c201 bl[201] br[201] wl[100] vdd gnd cell_6t
Xbit_r101_c201 bl[201] br[201] wl[101] vdd gnd cell_6t
Xbit_r102_c201 bl[201] br[201] wl[102] vdd gnd cell_6t
Xbit_r103_c201 bl[201] br[201] wl[103] vdd gnd cell_6t
Xbit_r104_c201 bl[201] br[201] wl[104] vdd gnd cell_6t
Xbit_r105_c201 bl[201] br[201] wl[105] vdd gnd cell_6t
Xbit_r106_c201 bl[201] br[201] wl[106] vdd gnd cell_6t
Xbit_r107_c201 bl[201] br[201] wl[107] vdd gnd cell_6t
Xbit_r108_c201 bl[201] br[201] wl[108] vdd gnd cell_6t
Xbit_r109_c201 bl[201] br[201] wl[109] vdd gnd cell_6t
Xbit_r110_c201 bl[201] br[201] wl[110] vdd gnd cell_6t
Xbit_r111_c201 bl[201] br[201] wl[111] vdd gnd cell_6t
Xbit_r112_c201 bl[201] br[201] wl[112] vdd gnd cell_6t
Xbit_r113_c201 bl[201] br[201] wl[113] vdd gnd cell_6t
Xbit_r114_c201 bl[201] br[201] wl[114] vdd gnd cell_6t
Xbit_r115_c201 bl[201] br[201] wl[115] vdd gnd cell_6t
Xbit_r116_c201 bl[201] br[201] wl[116] vdd gnd cell_6t
Xbit_r117_c201 bl[201] br[201] wl[117] vdd gnd cell_6t
Xbit_r118_c201 bl[201] br[201] wl[118] vdd gnd cell_6t
Xbit_r119_c201 bl[201] br[201] wl[119] vdd gnd cell_6t
Xbit_r120_c201 bl[201] br[201] wl[120] vdd gnd cell_6t
Xbit_r121_c201 bl[201] br[201] wl[121] vdd gnd cell_6t
Xbit_r122_c201 bl[201] br[201] wl[122] vdd gnd cell_6t
Xbit_r123_c201 bl[201] br[201] wl[123] vdd gnd cell_6t
Xbit_r124_c201 bl[201] br[201] wl[124] vdd gnd cell_6t
Xbit_r125_c201 bl[201] br[201] wl[125] vdd gnd cell_6t
Xbit_r126_c201 bl[201] br[201] wl[126] vdd gnd cell_6t
Xbit_r127_c201 bl[201] br[201] wl[127] vdd gnd cell_6t
Xbit_r0_c202 bl[202] br[202] wl[0] vdd gnd cell_6t
Xbit_r1_c202 bl[202] br[202] wl[1] vdd gnd cell_6t
Xbit_r2_c202 bl[202] br[202] wl[2] vdd gnd cell_6t
Xbit_r3_c202 bl[202] br[202] wl[3] vdd gnd cell_6t
Xbit_r4_c202 bl[202] br[202] wl[4] vdd gnd cell_6t
Xbit_r5_c202 bl[202] br[202] wl[5] vdd gnd cell_6t
Xbit_r6_c202 bl[202] br[202] wl[6] vdd gnd cell_6t
Xbit_r7_c202 bl[202] br[202] wl[7] vdd gnd cell_6t
Xbit_r8_c202 bl[202] br[202] wl[8] vdd gnd cell_6t
Xbit_r9_c202 bl[202] br[202] wl[9] vdd gnd cell_6t
Xbit_r10_c202 bl[202] br[202] wl[10] vdd gnd cell_6t
Xbit_r11_c202 bl[202] br[202] wl[11] vdd gnd cell_6t
Xbit_r12_c202 bl[202] br[202] wl[12] vdd gnd cell_6t
Xbit_r13_c202 bl[202] br[202] wl[13] vdd gnd cell_6t
Xbit_r14_c202 bl[202] br[202] wl[14] vdd gnd cell_6t
Xbit_r15_c202 bl[202] br[202] wl[15] vdd gnd cell_6t
Xbit_r16_c202 bl[202] br[202] wl[16] vdd gnd cell_6t
Xbit_r17_c202 bl[202] br[202] wl[17] vdd gnd cell_6t
Xbit_r18_c202 bl[202] br[202] wl[18] vdd gnd cell_6t
Xbit_r19_c202 bl[202] br[202] wl[19] vdd gnd cell_6t
Xbit_r20_c202 bl[202] br[202] wl[20] vdd gnd cell_6t
Xbit_r21_c202 bl[202] br[202] wl[21] vdd gnd cell_6t
Xbit_r22_c202 bl[202] br[202] wl[22] vdd gnd cell_6t
Xbit_r23_c202 bl[202] br[202] wl[23] vdd gnd cell_6t
Xbit_r24_c202 bl[202] br[202] wl[24] vdd gnd cell_6t
Xbit_r25_c202 bl[202] br[202] wl[25] vdd gnd cell_6t
Xbit_r26_c202 bl[202] br[202] wl[26] vdd gnd cell_6t
Xbit_r27_c202 bl[202] br[202] wl[27] vdd gnd cell_6t
Xbit_r28_c202 bl[202] br[202] wl[28] vdd gnd cell_6t
Xbit_r29_c202 bl[202] br[202] wl[29] vdd gnd cell_6t
Xbit_r30_c202 bl[202] br[202] wl[30] vdd gnd cell_6t
Xbit_r31_c202 bl[202] br[202] wl[31] vdd gnd cell_6t
Xbit_r32_c202 bl[202] br[202] wl[32] vdd gnd cell_6t
Xbit_r33_c202 bl[202] br[202] wl[33] vdd gnd cell_6t
Xbit_r34_c202 bl[202] br[202] wl[34] vdd gnd cell_6t
Xbit_r35_c202 bl[202] br[202] wl[35] vdd gnd cell_6t
Xbit_r36_c202 bl[202] br[202] wl[36] vdd gnd cell_6t
Xbit_r37_c202 bl[202] br[202] wl[37] vdd gnd cell_6t
Xbit_r38_c202 bl[202] br[202] wl[38] vdd gnd cell_6t
Xbit_r39_c202 bl[202] br[202] wl[39] vdd gnd cell_6t
Xbit_r40_c202 bl[202] br[202] wl[40] vdd gnd cell_6t
Xbit_r41_c202 bl[202] br[202] wl[41] vdd gnd cell_6t
Xbit_r42_c202 bl[202] br[202] wl[42] vdd gnd cell_6t
Xbit_r43_c202 bl[202] br[202] wl[43] vdd gnd cell_6t
Xbit_r44_c202 bl[202] br[202] wl[44] vdd gnd cell_6t
Xbit_r45_c202 bl[202] br[202] wl[45] vdd gnd cell_6t
Xbit_r46_c202 bl[202] br[202] wl[46] vdd gnd cell_6t
Xbit_r47_c202 bl[202] br[202] wl[47] vdd gnd cell_6t
Xbit_r48_c202 bl[202] br[202] wl[48] vdd gnd cell_6t
Xbit_r49_c202 bl[202] br[202] wl[49] vdd gnd cell_6t
Xbit_r50_c202 bl[202] br[202] wl[50] vdd gnd cell_6t
Xbit_r51_c202 bl[202] br[202] wl[51] vdd gnd cell_6t
Xbit_r52_c202 bl[202] br[202] wl[52] vdd gnd cell_6t
Xbit_r53_c202 bl[202] br[202] wl[53] vdd gnd cell_6t
Xbit_r54_c202 bl[202] br[202] wl[54] vdd gnd cell_6t
Xbit_r55_c202 bl[202] br[202] wl[55] vdd gnd cell_6t
Xbit_r56_c202 bl[202] br[202] wl[56] vdd gnd cell_6t
Xbit_r57_c202 bl[202] br[202] wl[57] vdd gnd cell_6t
Xbit_r58_c202 bl[202] br[202] wl[58] vdd gnd cell_6t
Xbit_r59_c202 bl[202] br[202] wl[59] vdd gnd cell_6t
Xbit_r60_c202 bl[202] br[202] wl[60] vdd gnd cell_6t
Xbit_r61_c202 bl[202] br[202] wl[61] vdd gnd cell_6t
Xbit_r62_c202 bl[202] br[202] wl[62] vdd gnd cell_6t
Xbit_r63_c202 bl[202] br[202] wl[63] vdd gnd cell_6t
Xbit_r64_c202 bl[202] br[202] wl[64] vdd gnd cell_6t
Xbit_r65_c202 bl[202] br[202] wl[65] vdd gnd cell_6t
Xbit_r66_c202 bl[202] br[202] wl[66] vdd gnd cell_6t
Xbit_r67_c202 bl[202] br[202] wl[67] vdd gnd cell_6t
Xbit_r68_c202 bl[202] br[202] wl[68] vdd gnd cell_6t
Xbit_r69_c202 bl[202] br[202] wl[69] vdd gnd cell_6t
Xbit_r70_c202 bl[202] br[202] wl[70] vdd gnd cell_6t
Xbit_r71_c202 bl[202] br[202] wl[71] vdd gnd cell_6t
Xbit_r72_c202 bl[202] br[202] wl[72] vdd gnd cell_6t
Xbit_r73_c202 bl[202] br[202] wl[73] vdd gnd cell_6t
Xbit_r74_c202 bl[202] br[202] wl[74] vdd gnd cell_6t
Xbit_r75_c202 bl[202] br[202] wl[75] vdd gnd cell_6t
Xbit_r76_c202 bl[202] br[202] wl[76] vdd gnd cell_6t
Xbit_r77_c202 bl[202] br[202] wl[77] vdd gnd cell_6t
Xbit_r78_c202 bl[202] br[202] wl[78] vdd gnd cell_6t
Xbit_r79_c202 bl[202] br[202] wl[79] vdd gnd cell_6t
Xbit_r80_c202 bl[202] br[202] wl[80] vdd gnd cell_6t
Xbit_r81_c202 bl[202] br[202] wl[81] vdd gnd cell_6t
Xbit_r82_c202 bl[202] br[202] wl[82] vdd gnd cell_6t
Xbit_r83_c202 bl[202] br[202] wl[83] vdd gnd cell_6t
Xbit_r84_c202 bl[202] br[202] wl[84] vdd gnd cell_6t
Xbit_r85_c202 bl[202] br[202] wl[85] vdd gnd cell_6t
Xbit_r86_c202 bl[202] br[202] wl[86] vdd gnd cell_6t
Xbit_r87_c202 bl[202] br[202] wl[87] vdd gnd cell_6t
Xbit_r88_c202 bl[202] br[202] wl[88] vdd gnd cell_6t
Xbit_r89_c202 bl[202] br[202] wl[89] vdd gnd cell_6t
Xbit_r90_c202 bl[202] br[202] wl[90] vdd gnd cell_6t
Xbit_r91_c202 bl[202] br[202] wl[91] vdd gnd cell_6t
Xbit_r92_c202 bl[202] br[202] wl[92] vdd gnd cell_6t
Xbit_r93_c202 bl[202] br[202] wl[93] vdd gnd cell_6t
Xbit_r94_c202 bl[202] br[202] wl[94] vdd gnd cell_6t
Xbit_r95_c202 bl[202] br[202] wl[95] vdd gnd cell_6t
Xbit_r96_c202 bl[202] br[202] wl[96] vdd gnd cell_6t
Xbit_r97_c202 bl[202] br[202] wl[97] vdd gnd cell_6t
Xbit_r98_c202 bl[202] br[202] wl[98] vdd gnd cell_6t
Xbit_r99_c202 bl[202] br[202] wl[99] vdd gnd cell_6t
Xbit_r100_c202 bl[202] br[202] wl[100] vdd gnd cell_6t
Xbit_r101_c202 bl[202] br[202] wl[101] vdd gnd cell_6t
Xbit_r102_c202 bl[202] br[202] wl[102] vdd gnd cell_6t
Xbit_r103_c202 bl[202] br[202] wl[103] vdd gnd cell_6t
Xbit_r104_c202 bl[202] br[202] wl[104] vdd gnd cell_6t
Xbit_r105_c202 bl[202] br[202] wl[105] vdd gnd cell_6t
Xbit_r106_c202 bl[202] br[202] wl[106] vdd gnd cell_6t
Xbit_r107_c202 bl[202] br[202] wl[107] vdd gnd cell_6t
Xbit_r108_c202 bl[202] br[202] wl[108] vdd gnd cell_6t
Xbit_r109_c202 bl[202] br[202] wl[109] vdd gnd cell_6t
Xbit_r110_c202 bl[202] br[202] wl[110] vdd gnd cell_6t
Xbit_r111_c202 bl[202] br[202] wl[111] vdd gnd cell_6t
Xbit_r112_c202 bl[202] br[202] wl[112] vdd gnd cell_6t
Xbit_r113_c202 bl[202] br[202] wl[113] vdd gnd cell_6t
Xbit_r114_c202 bl[202] br[202] wl[114] vdd gnd cell_6t
Xbit_r115_c202 bl[202] br[202] wl[115] vdd gnd cell_6t
Xbit_r116_c202 bl[202] br[202] wl[116] vdd gnd cell_6t
Xbit_r117_c202 bl[202] br[202] wl[117] vdd gnd cell_6t
Xbit_r118_c202 bl[202] br[202] wl[118] vdd gnd cell_6t
Xbit_r119_c202 bl[202] br[202] wl[119] vdd gnd cell_6t
Xbit_r120_c202 bl[202] br[202] wl[120] vdd gnd cell_6t
Xbit_r121_c202 bl[202] br[202] wl[121] vdd gnd cell_6t
Xbit_r122_c202 bl[202] br[202] wl[122] vdd gnd cell_6t
Xbit_r123_c202 bl[202] br[202] wl[123] vdd gnd cell_6t
Xbit_r124_c202 bl[202] br[202] wl[124] vdd gnd cell_6t
Xbit_r125_c202 bl[202] br[202] wl[125] vdd gnd cell_6t
Xbit_r126_c202 bl[202] br[202] wl[126] vdd gnd cell_6t
Xbit_r127_c202 bl[202] br[202] wl[127] vdd gnd cell_6t
Xbit_r0_c203 bl[203] br[203] wl[0] vdd gnd cell_6t
Xbit_r1_c203 bl[203] br[203] wl[1] vdd gnd cell_6t
Xbit_r2_c203 bl[203] br[203] wl[2] vdd gnd cell_6t
Xbit_r3_c203 bl[203] br[203] wl[3] vdd gnd cell_6t
Xbit_r4_c203 bl[203] br[203] wl[4] vdd gnd cell_6t
Xbit_r5_c203 bl[203] br[203] wl[5] vdd gnd cell_6t
Xbit_r6_c203 bl[203] br[203] wl[6] vdd gnd cell_6t
Xbit_r7_c203 bl[203] br[203] wl[7] vdd gnd cell_6t
Xbit_r8_c203 bl[203] br[203] wl[8] vdd gnd cell_6t
Xbit_r9_c203 bl[203] br[203] wl[9] vdd gnd cell_6t
Xbit_r10_c203 bl[203] br[203] wl[10] vdd gnd cell_6t
Xbit_r11_c203 bl[203] br[203] wl[11] vdd gnd cell_6t
Xbit_r12_c203 bl[203] br[203] wl[12] vdd gnd cell_6t
Xbit_r13_c203 bl[203] br[203] wl[13] vdd gnd cell_6t
Xbit_r14_c203 bl[203] br[203] wl[14] vdd gnd cell_6t
Xbit_r15_c203 bl[203] br[203] wl[15] vdd gnd cell_6t
Xbit_r16_c203 bl[203] br[203] wl[16] vdd gnd cell_6t
Xbit_r17_c203 bl[203] br[203] wl[17] vdd gnd cell_6t
Xbit_r18_c203 bl[203] br[203] wl[18] vdd gnd cell_6t
Xbit_r19_c203 bl[203] br[203] wl[19] vdd gnd cell_6t
Xbit_r20_c203 bl[203] br[203] wl[20] vdd gnd cell_6t
Xbit_r21_c203 bl[203] br[203] wl[21] vdd gnd cell_6t
Xbit_r22_c203 bl[203] br[203] wl[22] vdd gnd cell_6t
Xbit_r23_c203 bl[203] br[203] wl[23] vdd gnd cell_6t
Xbit_r24_c203 bl[203] br[203] wl[24] vdd gnd cell_6t
Xbit_r25_c203 bl[203] br[203] wl[25] vdd gnd cell_6t
Xbit_r26_c203 bl[203] br[203] wl[26] vdd gnd cell_6t
Xbit_r27_c203 bl[203] br[203] wl[27] vdd gnd cell_6t
Xbit_r28_c203 bl[203] br[203] wl[28] vdd gnd cell_6t
Xbit_r29_c203 bl[203] br[203] wl[29] vdd gnd cell_6t
Xbit_r30_c203 bl[203] br[203] wl[30] vdd gnd cell_6t
Xbit_r31_c203 bl[203] br[203] wl[31] vdd gnd cell_6t
Xbit_r32_c203 bl[203] br[203] wl[32] vdd gnd cell_6t
Xbit_r33_c203 bl[203] br[203] wl[33] vdd gnd cell_6t
Xbit_r34_c203 bl[203] br[203] wl[34] vdd gnd cell_6t
Xbit_r35_c203 bl[203] br[203] wl[35] vdd gnd cell_6t
Xbit_r36_c203 bl[203] br[203] wl[36] vdd gnd cell_6t
Xbit_r37_c203 bl[203] br[203] wl[37] vdd gnd cell_6t
Xbit_r38_c203 bl[203] br[203] wl[38] vdd gnd cell_6t
Xbit_r39_c203 bl[203] br[203] wl[39] vdd gnd cell_6t
Xbit_r40_c203 bl[203] br[203] wl[40] vdd gnd cell_6t
Xbit_r41_c203 bl[203] br[203] wl[41] vdd gnd cell_6t
Xbit_r42_c203 bl[203] br[203] wl[42] vdd gnd cell_6t
Xbit_r43_c203 bl[203] br[203] wl[43] vdd gnd cell_6t
Xbit_r44_c203 bl[203] br[203] wl[44] vdd gnd cell_6t
Xbit_r45_c203 bl[203] br[203] wl[45] vdd gnd cell_6t
Xbit_r46_c203 bl[203] br[203] wl[46] vdd gnd cell_6t
Xbit_r47_c203 bl[203] br[203] wl[47] vdd gnd cell_6t
Xbit_r48_c203 bl[203] br[203] wl[48] vdd gnd cell_6t
Xbit_r49_c203 bl[203] br[203] wl[49] vdd gnd cell_6t
Xbit_r50_c203 bl[203] br[203] wl[50] vdd gnd cell_6t
Xbit_r51_c203 bl[203] br[203] wl[51] vdd gnd cell_6t
Xbit_r52_c203 bl[203] br[203] wl[52] vdd gnd cell_6t
Xbit_r53_c203 bl[203] br[203] wl[53] vdd gnd cell_6t
Xbit_r54_c203 bl[203] br[203] wl[54] vdd gnd cell_6t
Xbit_r55_c203 bl[203] br[203] wl[55] vdd gnd cell_6t
Xbit_r56_c203 bl[203] br[203] wl[56] vdd gnd cell_6t
Xbit_r57_c203 bl[203] br[203] wl[57] vdd gnd cell_6t
Xbit_r58_c203 bl[203] br[203] wl[58] vdd gnd cell_6t
Xbit_r59_c203 bl[203] br[203] wl[59] vdd gnd cell_6t
Xbit_r60_c203 bl[203] br[203] wl[60] vdd gnd cell_6t
Xbit_r61_c203 bl[203] br[203] wl[61] vdd gnd cell_6t
Xbit_r62_c203 bl[203] br[203] wl[62] vdd gnd cell_6t
Xbit_r63_c203 bl[203] br[203] wl[63] vdd gnd cell_6t
Xbit_r64_c203 bl[203] br[203] wl[64] vdd gnd cell_6t
Xbit_r65_c203 bl[203] br[203] wl[65] vdd gnd cell_6t
Xbit_r66_c203 bl[203] br[203] wl[66] vdd gnd cell_6t
Xbit_r67_c203 bl[203] br[203] wl[67] vdd gnd cell_6t
Xbit_r68_c203 bl[203] br[203] wl[68] vdd gnd cell_6t
Xbit_r69_c203 bl[203] br[203] wl[69] vdd gnd cell_6t
Xbit_r70_c203 bl[203] br[203] wl[70] vdd gnd cell_6t
Xbit_r71_c203 bl[203] br[203] wl[71] vdd gnd cell_6t
Xbit_r72_c203 bl[203] br[203] wl[72] vdd gnd cell_6t
Xbit_r73_c203 bl[203] br[203] wl[73] vdd gnd cell_6t
Xbit_r74_c203 bl[203] br[203] wl[74] vdd gnd cell_6t
Xbit_r75_c203 bl[203] br[203] wl[75] vdd gnd cell_6t
Xbit_r76_c203 bl[203] br[203] wl[76] vdd gnd cell_6t
Xbit_r77_c203 bl[203] br[203] wl[77] vdd gnd cell_6t
Xbit_r78_c203 bl[203] br[203] wl[78] vdd gnd cell_6t
Xbit_r79_c203 bl[203] br[203] wl[79] vdd gnd cell_6t
Xbit_r80_c203 bl[203] br[203] wl[80] vdd gnd cell_6t
Xbit_r81_c203 bl[203] br[203] wl[81] vdd gnd cell_6t
Xbit_r82_c203 bl[203] br[203] wl[82] vdd gnd cell_6t
Xbit_r83_c203 bl[203] br[203] wl[83] vdd gnd cell_6t
Xbit_r84_c203 bl[203] br[203] wl[84] vdd gnd cell_6t
Xbit_r85_c203 bl[203] br[203] wl[85] vdd gnd cell_6t
Xbit_r86_c203 bl[203] br[203] wl[86] vdd gnd cell_6t
Xbit_r87_c203 bl[203] br[203] wl[87] vdd gnd cell_6t
Xbit_r88_c203 bl[203] br[203] wl[88] vdd gnd cell_6t
Xbit_r89_c203 bl[203] br[203] wl[89] vdd gnd cell_6t
Xbit_r90_c203 bl[203] br[203] wl[90] vdd gnd cell_6t
Xbit_r91_c203 bl[203] br[203] wl[91] vdd gnd cell_6t
Xbit_r92_c203 bl[203] br[203] wl[92] vdd gnd cell_6t
Xbit_r93_c203 bl[203] br[203] wl[93] vdd gnd cell_6t
Xbit_r94_c203 bl[203] br[203] wl[94] vdd gnd cell_6t
Xbit_r95_c203 bl[203] br[203] wl[95] vdd gnd cell_6t
Xbit_r96_c203 bl[203] br[203] wl[96] vdd gnd cell_6t
Xbit_r97_c203 bl[203] br[203] wl[97] vdd gnd cell_6t
Xbit_r98_c203 bl[203] br[203] wl[98] vdd gnd cell_6t
Xbit_r99_c203 bl[203] br[203] wl[99] vdd gnd cell_6t
Xbit_r100_c203 bl[203] br[203] wl[100] vdd gnd cell_6t
Xbit_r101_c203 bl[203] br[203] wl[101] vdd gnd cell_6t
Xbit_r102_c203 bl[203] br[203] wl[102] vdd gnd cell_6t
Xbit_r103_c203 bl[203] br[203] wl[103] vdd gnd cell_6t
Xbit_r104_c203 bl[203] br[203] wl[104] vdd gnd cell_6t
Xbit_r105_c203 bl[203] br[203] wl[105] vdd gnd cell_6t
Xbit_r106_c203 bl[203] br[203] wl[106] vdd gnd cell_6t
Xbit_r107_c203 bl[203] br[203] wl[107] vdd gnd cell_6t
Xbit_r108_c203 bl[203] br[203] wl[108] vdd gnd cell_6t
Xbit_r109_c203 bl[203] br[203] wl[109] vdd gnd cell_6t
Xbit_r110_c203 bl[203] br[203] wl[110] vdd gnd cell_6t
Xbit_r111_c203 bl[203] br[203] wl[111] vdd gnd cell_6t
Xbit_r112_c203 bl[203] br[203] wl[112] vdd gnd cell_6t
Xbit_r113_c203 bl[203] br[203] wl[113] vdd gnd cell_6t
Xbit_r114_c203 bl[203] br[203] wl[114] vdd gnd cell_6t
Xbit_r115_c203 bl[203] br[203] wl[115] vdd gnd cell_6t
Xbit_r116_c203 bl[203] br[203] wl[116] vdd gnd cell_6t
Xbit_r117_c203 bl[203] br[203] wl[117] vdd gnd cell_6t
Xbit_r118_c203 bl[203] br[203] wl[118] vdd gnd cell_6t
Xbit_r119_c203 bl[203] br[203] wl[119] vdd gnd cell_6t
Xbit_r120_c203 bl[203] br[203] wl[120] vdd gnd cell_6t
Xbit_r121_c203 bl[203] br[203] wl[121] vdd gnd cell_6t
Xbit_r122_c203 bl[203] br[203] wl[122] vdd gnd cell_6t
Xbit_r123_c203 bl[203] br[203] wl[123] vdd gnd cell_6t
Xbit_r124_c203 bl[203] br[203] wl[124] vdd gnd cell_6t
Xbit_r125_c203 bl[203] br[203] wl[125] vdd gnd cell_6t
Xbit_r126_c203 bl[203] br[203] wl[126] vdd gnd cell_6t
Xbit_r127_c203 bl[203] br[203] wl[127] vdd gnd cell_6t
Xbit_r0_c204 bl[204] br[204] wl[0] vdd gnd cell_6t
Xbit_r1_c204 bl[204] br[204] wl[1] vdd gnd cell_6t
Xbit_r2_c204 bl[204] br[204] wl[2] vdd gnd cell_6t
Xbit_r3_c204 bl[204] br[204] wl[3] vdd gnd cell_6t
Xbit_r4_c204 bl[204] br[204] wl[4] vdd gnd cell_6t
Xbit_r5_c204 bl[204] br[204] wl[5] vdd gnd cell_6t
Xbit_r6_c204 bl[204] br[204] wl[6] vdd gnd cell_6t
Xbit_r7_c204 bl[204] br[204] wl[7] vdd gnd cell_6t
Xbit_r8_c204 bl[204] br[204] wl[8] vdd gnd cell_6t
Xbit_r9_c204 bl[204] br[204] wl[9] vdd gnd cell_6t
Xbit_r10_c204 bl[204] br[204] wl[10] vdd gnd cell_6t
Xbit_r11_c204 bl[204] br[204] wl[11] vdd gnd cell_6t
Xbit_r12_c204 bl[204] br[204] wl[12] vdd gnd cell_6t
Xbit_r13_c204 bl[204] br[204] wl[13] vdd gnd cell_6t
Xbit_r14_c204 bl[204] br[204] wl[14] vdd gnd cell_6t
Xbit_r15_c204 bl[204] br[204] wl[15] vdd gnd cell_6t
Xbit_r16_c204 bl[204] br[204] wl[16] vdd gnd cell_6t
Xbit_r17_c204 bl[204] br[204] wl[17] vdd gnd cell_6t
Xbit_r18_c204 bl[204] br[204] wl[18] vdd gnd cell_6t
Xbit_r19_c204 bl[204] br[204] wl[19] vdd gnd cell_6t
Xbit_r20_c204 bl[204] br[204] wl[20] vdd gnd cell_6t
Xbit_r21_c204 bl[204] br[204] wl[21] vdd gnd cell_6t
Xbit_r22_c204 bl[204] br[204] wl[22] vdd gnd cell_6t
Xbit_r23_c204 bl[204] br[204] wl[23] vdd gnd cell_6t
Xbit_r24_c204 bl[204] br[204] wl[24] vdd gnd cell_6t
Xbit_r25_c204 bl[204] br[204] wl[25] vdd gnd cell_6t
Xbit_r26_c204 bl[204] br[204] wl[26] vdd gnd cell_6t
Xbit_r27_c204 bl[204] br[204] wl[27] vdd gnd cell_6t
Xbit_r28_c204 bl[204] br[204] wl[28] vdd gnd cell_6t
Xbit_r29_c204 bl[204] br[204] wl[29] vdd gnd cell_6t
Xbit_r30_c204 bl[204] br[204] wl[30] vdd gnd cell_6t
Xbit_r31_c204 bl[204] br[204] wl[31] vdd gnd cell_6t
Xbit_r32_c204 bl[204] br[204] wl[32] vdd gnd cell_6t
Xbit_r33_c204 bl[204] br[204] wl[33] vdd gnd cell_6t
Xbit_r34_c204 bl[204] br[204] wl[34] vdd gnd cell_6t
Xbit_r35_c204 bl[204] br[204] wl[35] vdd gnd cell_6t
Xbit_r36_c204 bl[204] br[204] wl[36] vdd gnd cell_6t
Xbit_r37_c204 bl[204] br[204] wl[37] vdd gnd cell_6t
Xbit_r38_c204 bl[204] br[204] wl[38] vdd gnd cell_6t
Xbit_r39_c204 bl[204] br[204] wl[39] vdd gnd cell_6t
Xbit_r40_c204 bl[204] br[204] wl[40] vdd gnd cell_6t
Xbit_r41_c204 bl[204] br[204] wl[41] vdd gnd cell_6t
Xbit_r42_c204 bl[204] br[204] wl[42] vdd gnd cell_6t
Xbit_r43_c204 bl[204] br[204] wl[43] vdd gnd cell_6t
Xbit_r44_c204 bl[204] br[204] wl[44] vdd gnd cell_6t
Xbit_r45_c204 bl[204] br[204] wl[45] vdd gnd cell_6t
Xbit_r46_c204 bl[204] br[204] wl[46] vdd gnd cell_6t
Xbit_r47_c204 bl[204] br[204] wl[47] vdd gnd cell_6t
Xbit_r48_c204 bl[204] br[204] wl[48] vdd gnd cell_6t
Xbit_r49_c204 bl[204] br[204] wl[49] vdd gnd cell_6t
Xbit_r50_c204 bl[204] br[204] wl[50] vdd gnd cell_6t
Xbit_r51_c204 bl[204] br[204] wl[51] vdd gnd cell_6t
Xbit_r52_c204 bl[204] br[204] wl[52] vdd gnd cell_6t
Xbit_r53_c204 bl[204] br[204] wl[53] vdd gnd cell_6t
Xbit_r54_c204 bl[204] br[204] wl[54] vdd gnd cell_6t
Xbit_r55_c204 bl[204] br[204] wl[55] vdd gnd cell_6t
Xbit_r56_c204 bl[204] br[204] wl[56] vdd gnd cell_6t
Xbit_r57_c204 bl[204] br[204] wl[57] vdd gnd cell_6t
Xbit_r58_c204 bl[204] br[204] wl[58] vdd gnd cell_6t
Xbit_r59_c204 bl[204] br[204] wl[59] vdd gnd cell_6t
Xbit_r60_c204 bl[204] br[204] wl[60] vdd gnd cell_6t
Xbit_r61_c204 bl[204] br[204] wl[61] vdd gnd cell_6t
Xbit_r62_c204 bl[204] br[204] wl[62] vdd gnd cell_6t
Xbit_r63_c204 bl[204] br[204] wl[63] vdd gnd cell_6t
Xbit_r64_c204 bl[204] br[204] wl[64] vdd gnd cell_6t
Xbit_r65_c204 bl[204] br[204] wl[65] vdd gnd cell_6t
Xbit_r66_c204 bl[204] br[204] wl[66] vdd gnd cell_6t
Xbit_r67_c204 bl[204] br[204] wl[67] vdd gnd cell_6t
Xbit_r68_c204 bl[204] br[204] wl[68] vdd gnd cell_6t
Xbit_r69_c204 bl[204] br[204] wl[69] vdd gnd cell_6t
Xbit_r70_c204 bl[204] br[204] wl[70] vdd gnd cell_6t
Xbit_r71_c204 bl[204] br[204] wl[71] vdd gnd cell_6t
Xbit_r72_c204 bl[204] br[204] wl[72] vdd gnd cell_6t
Xbit_r73_c204 bl[204] br[204] wl[73] vdd gnd cell_6t
Xbit_r74_c204 bl[204] br[204] wl[74] vdd gnd cell_6t
Xbit_r75_c204 bl[204] br[204] wl[75] vdd gnd cell_6t
Xbit_r76_c204 bl[204] br[204] wl[76] vdd gnd cell_6t
Xbit_r77_c204 bl[204] br[204] wl[77] vdd gnd cell_6t
Xbit_r78_c204 bl[204] br[204] wl[78] vdd gnd cell_6t
Xbit_r79_c204 bl[204] br[204] wl[79] vdd gnd cell_6t
Xbit_r80_c204 bl[204] br[204] wl[80] vdd gnd cell_6t
Xbit_r81_c204 bl[204] br[204] wl[81] vdd gnd cell_6t
Xbit_r82_c204 bl[204] br[204] wl[82] vdd gnd cell_6t
Xbit_r83_c204 bl[204] br[204] wl[83] vdd gnd cell_6t
Xbit_r84_c204 bl[204] br[204] wl[84] vdd gnd cell_6t
Xbit_r85_c204 bl[204] br[204] wl[85] vdd gnd cell_6t
Xbit_r86_c204 bl[204] br[204] wl[86] vdd gnd cell_6t
Xbit_r87_c204 bl[204] br[204] wl[87] vdd gnd cell_6t
Xbit_r88_c204 bl[204] br[204] wl[88] vdd gnd cell_6t
Xbit_r89_c204 bl[204] br[204] wl[89] vdd gnd cell_6t
Xbit_r90_c204 bl[204] br[204] wl[90] vdd gnd cell_6t
Xbit_r91_c204 bl[204] br[204] wl[91] vdd gnd cell_6t
Xbit_r92_c204 bl[204] br[204] wl[92] vdd gnd cell_6t
Xbit_r93_c204 bl[204] br[204] wl[93] vdd gnd cell_6t
Xbit_r94_c204 bl[204] br[204] wl[94] vdd gnd cell_6t
Xbit_r95_c204 bl[204] br[204] wl[95] vdd gnd cell_6t
Xbit_r96_c204 bl[204] br[204] wl[96] vdd gnd cell_6t
Xbit_r97_c204 bl[204] br[204] wl[97] vdd gnd cell_6t
Xbit_r98_c204 bl[204] br[204] wl[98] vdd gnd cell_6t
Xbit_r99_c204 bl[204] br[204] wl[99] vdd gnd cell_6t
Xbit_r100_c204 bl[204] br[204] wl[100] vdd gnd cell_6t
Xbit_r101_c204 bl[204] br[204] wl[101] vdd gnd cell_6t
Xbit_r102_c204 bl[204] br[204] wl[102] vdd gnd cell_6t
Xbit_r103_c204 bl[204] br[204] wl[103] vdd gnd cell_6t
Xbit_r104_c204 bl[204] br[204] wl[104] vdd gnd cell_6t
Xbit_r105_c204 bl[204] br[204] wl[105] vdd gnd cell_6t
Xbit_r106_c204 bl[204] br[204] wl[106] vdd gnd cell_6t
Xbit_r107_c204 bl[204] br[204] wl[107] vdd gnd cell_6t
Xbit_r108_c204 bl[204] br[204] wl[108] vdd gnd cell_6t
Xbit_r109_c204 bl[204] br[204] wl[109] vdd gnd cell_6t
Xbit_r110_c204 bl[204] br[204] wl[110] vdd gnd cell_6t
Xbit_r111_c204 bl[204] br[204] wl[111] vdd gnd cell_6t
Xbit_r112_c204 bl[204] br[204] wl[112] vdd gnd cell_6t
Xbit_r113_c204 bl[204] br[204] wl[113] vdd gnd cell_6t
Xbit_r114_c204 bl[204] br[204] wl[114] vdd gnd cell_6t
Xbit_r115_c204 bl[204] br[204] wl[115] vdd gnd cell_6t
Xbit_r116_c204 bl[204] br[204] wl[116] vdd gnd cell_6t
Xbit_r117_c204 bl[204] br[204] wl[117] vdd gnd cell_6t
Xbit_r118_c204 bl[204] br[204] wl[118] vdd gnd cell_6t
Xbit_r119_c204 bl[204] br[204] wl[119] vdd gnd cell_6t
Xbit_r120_c204 bl[204] br[204] wl[120] vdd gnd cell_6t
Xbit_r121_c204 bl[204] br[204] wl[121] vdd gnd cell_6t
Xbit_r122_c204 bl[204] br[204] wl[122] vdd gnd cell_6t
Xbit_r123_c204 bl[204] br[204] wl[123] vdd gnd cell_6t
Xbit_r124_c204 bl[204] br[204] wl[124] vdd gnd cell_6t
Xbit_r125_c204 bl[204] br[204] wl[125] vdd gnd cell_6t
Xbit_r126_c204 bl[204] br[204] wl[126] vdd gnd cell_6t
Xbit_r127_c204 bl[204] br[204] wl[127] vdd gnd cell_6t
Xbit_r0_c205 bl[205] br[205] wl[0] vdd gnd cell_6t
Xbit_r1_c205 bl[205] br[205] wl[1] vdd gnd cell_6t
Xbit_r2_c205 bl[205] br[205] wl[2] vdd gnd cell_6t
Xbit_r3_c205 bl[205] br[205] wl[3] vdd gnd cell_6t
Xbit_r4_c205 bl[205] br[205] wl[4] vdd gnd cell_6t
Xbit_r5_c205 bl[205] br[205] wl[5] vdd gnd cell_6t
Xbit_r6_c205 bl[205] br[205] wl[6] vdd gnd cell_6t
Xbit_r7_c205 bl[205] br[205] wl[7] vdd gnd cell_6t
Xbit_r8_c205 bl[205] br[205] wl[8] vdd gnd cell_6t
Xbit_r9_c205 bl[205] br[205] wl[9] vdd gnd cell_6t
Xbit_r10_c205 bl[205] br[205] wl[10] vdd gnd cell_6t
Xbit_r11_c205 bl[205] br[205] wl[11] vdd gnd cell_6t
Xbit_r12_c205 bl[205] br[205] wl[12] vdd gnd cell_6t
Xbit_r13_c205 bl[205] br[205] wl[13] vdd gnd cell_6t
Xbit_r14_c205 bl[205] br[205] wl[14] vdd gnd cell_6t
Xbit_r15_c205 bl[205] br[205] wl[15] vdd gnd cell_6t
Xbit_r16_c205 bl[205] br[205] wl[16] vdd gnd cell_6t
Xbit_r17_c205 bl[205] br[205] wl[17] vdd gnd cell_6t
Xbit_r18_c205 bl[205] br[205] wl[18] vdd gnd cell_6t
Xbit_r19_c205 bl[205] br[205] wl[19] vdd gnd cell_6t
Xbit_r20_c205 bl[205] br[205] wl[20] vdd gnd cell_6t
Xbit_r21_c205 bl[205] br[205] wl[21] vdd gnd cell_6t
Xbit_r22_c205 bl[205] br[205] wl[22] vdd gnd cell_6t
Xbit_r23_c205 bl[205] br[205] wl[23] vdd gnd cell_6t
Xbit_r24_c205 bl[205] br[205] wl[24] vdd gnd cell_6t
Xbit_r25_c205 bl[205] br[205] wl[25] vdd gnd cell_6t
Xbit_r26_c205 bl[205] br[205] wl[26] vdd gnd cell_6t
Xbit_r27_c205 bl[205] br[205] wl[27] vdd gnd cell_6t
Xbit_r28_c205 bl[205] br[205] wl[28] vdd gnd cell_6t
Xbit_r29_c205 bl[205] br[205] wl[29] vdd gnd cell_6t
Xbit_r30_c205 bl[205] br[205] wl[30] vdd gnd cell_6t
Xbit_r31_c205 bl[205] br[205] wl[31] vdd gnd cell_6t
Xbit_r32_c205 bl[205] br[205] wl[32] vdd gnd cell_6t
Xbit_r33_c205 bl[205] br[205] wl[33] vdd gnd cell_6t
Xbit_r34_c205 bl[205] br[205] wl[34] vdd gnd cell_6t
Xbit_r35_c205 bl[205] br[205] wl[35] vdd gnd cell_6t
Xbit_r36_c205 bl[205] br[205] wl[36] vdd gnd cell_6t
Xbit_r37_c205 bl[205] br[205] wl[37] vdd gnd cell_6t
Xbit_r38_c205 bl[205] br[205] wl[38] vdd gnd cell_6t
Xbit_r39_c205 bl[205] br[205] wl[39] vdd gnd cell_6t
Xbit_r40_c205 bl[205] br[205] wl[40] vdd gnd cell_6t
Xbit_r41_c205 bl[205] br[205] wl[41] vdd gnd cell_6t
Xbit_r42_c205 bl[205] br[205] wl[42] vdd gnd cell_6t
Xbit_r43_c205 bl[205] br[205] wl[43] vdd gnd cell_6t
Xbit_r44_c205 bl[205] br[205] wl[44] vdd gnd cell_6t
Xbit_r45_c205 bl[205] br[205] wl[45] vdd gnd cell_6t
Xbit_r46_c205 bl[205] br[205] wl[46] vdd gnd cell_6t
Xbit_r47_c205 bl[205] br[205] wl[47] vdd gnd cell_6t
Xbit_r48_c205 bl[205] br[205] wl[48] vdd gnd cell_6t
Xbit_r49_c205 bl[205] br[205] wl[49] vdd gnd cell_6t
Xbit_r50_c205 bl[205] br[205] wl[50] vdd gnd cell_6t
Xbit_r51_c205 bl[205] br[205] wl[51] vdd gnd cell_6t
Xbit_r52_c205 bl[205] br[205] wl[52] vdd gnd cell_6t
Xbit_r53_c205 bl[205] br[205] wl[53] vdd gnd cell_6t
Xbit_r54_c205 bl[205] br[205] wl[54] vdd gnd cell_6t
Xbit_r55_c205 bl[205] br[205] wl[55] vdd gnd cell_6t
Xbit_r56_c205 bl[205] br[205] wl[56] vdd gnd cell_6t
Xbit_r57_c205 bl[205] br[205] wl[57] vdd gnd cell_6t
Xbit_r58_c205 bl[205] br[205] wl[58] vdd gnd cell_6t
Xbit_r59_c205 bl[205] br[205] wl[59] vdd gnd cell_6t
Xbit_r60_c205 bl[205] br[205] wl[60] vdd gnd cell_6t
Xbit_r61_c205 bl[205] br[205] wl[61] vdd gnd cell_6t
Xbit_r62_c205 bl[205] br[205] wl[62] vdd gnd cell_6t
Xbit_r63_c205 bl[205] br[205] wl[63] vdd gnd cell_6t
Xbit_r64_c205 bl[205] br[205] wl[64] vdd gnd cell_6t
Xbit_r65_c205 bl[205] br[205] wl[65] vdd gnd cell_6t
Xbit_r66_c205 bl[205] br[205] wl[66] vdd gnd cell_6t
Xbit_r67_c205 bl[205] br[205] wl[67] vdd gnd cell_6t
Xbit_r68_c205 bl[205] br[205] wl[68] vdd gnd cell_6t
Xbit_r69_c205 bl[205] br[205] wl[69] vdd gnd cell_6t
Xbit_r70_c205 bl[205] br[205] wl[70] vdd gnd cell_6t
Xbit_r71_c205 bl[205] br[205] wl[71] vdd gnd cell_6t
Xbit_r72_c205 bl[205] br[205] wl[72] vdd gnd cell_6t
Xbit_r73_c205 bl[205] br[205] wl[73] vdd gnd cell_6t
Xbit_r74_c205 bl[205] br[205] wl[74] vdd gnd cell_6t
Xbit_r75_c205 bl[205] br[205] wl[75] vdd gnd cell_6t
Xbit_r76_c205 bl[205] br[205] wl[76] vdd gnd cell_6t
Xbit_r77_c205 bl[205] br[205] wl[77] vdd gnd cell_6t
Xbit_r78_c205 bl[205] br[205] wl[78] vdd gnd cell_6t
Xbit_r79_c205 bl[205] br[205] wl[79] vdd gnd cell_6t
Xbit_r80_c205 bl[205] br[205] wl[80] vdd gnd cell_6t
Xbit_r81_c205 bl[205] br[205] wl[81] vdd gnd cell_6t
Xbit_r82_c205 bl[205] br[205] wl[82] vdd gnd cell_6t
Xbit_r83_c205 bl[205] br[205] wl[83] vdd gnd cell_6t
Xbit_r84_c205 bl[205] br[205] wl[84] vdd gnd cell_6t
Xbit_r85_c205 bl[205] br[205] wl[85] vdd gnd cell_6t
Xbit_r86_c205 bl[205] br[205] wl[86] vdd gnd cell_6t
Xbit_r87_c205 bl[205] br[205] wl[87] vdd gnd cell_6t
Xbit_r88_c205 bl[205] br[205] wl[88] vdd gnd cell_6t
Xbit_r89_c205 bl[205] br[205] wl[89] vdd gnd cell_6t
Xbit_r90_c205 bl[205] br[205] wl[90] vdd gnd cell_6t
Xbit_r91_c205 bl[205] br[205] wl[91] vdd gnd cell_6t
Xbit_r92_c205 bl[205] br[205] wl[92] vdd gnd cell_6t
Xbit_r93_c205 bl[205] br[205] wl[93] vdd gnd cell_6t
Xbit_r94_c205 bl[205] br[205] wl[94] vdd gnd cell_6t
Xbit_r95_c205 bl[205] br[205] wl[95] vdd gnd cell_6t
Xbit_r96_c205 bl[205] br[205] wl[96] vdd gnd cell_6t
Xbit_r97_c205 bl[205] br[205] wl[97] vdd gnd cell_6t
Xbit_r98_c205 bl[205] br[205] wl[98] vdd gnd cell_6t
Xbit_r99_c205 bl[205] br[205] wl[99] vdd gnd cell_6t
Xbit_r100_c205 bl[205] br[205] wl[100] vdd gnd cell_6t
Xbit_r101_c205 bl[205] br[205] wl[101] vdd gnd cell_6t
Xbit_r102_c205 bl[205] br[205] wl[102] vdd gnd cell_6t
Xbit_r103_c205 bl[205] br[205] wl[103] vdd gnd cell_6t
Xbit_r104_c205 bl[205] br[205] wl[104] vdd gnd cell_6t
Xbit_r105_c205 bl[205] br[205] wl[105] vdd gnd cell_6t
Xbit_r106_c205 bl[205] br[205] wl[106] vdd gnd cell_6t
Xbit_r107_c205 bl[205] br[205] wl[107] vdd gnd cell_6t
Xbit_r108_c205 bl[205] br[205] wl[108] vdd gnd cell_6t
Xbit_r109_c205 bl[205] br[205] wl[109] vdd gnd cell_6t
Xbit_r110_c205 bl[205] br[205] wl[110] vdd gnd cell_6t
Xbit_r111_c205 bl[205] br[205] wl[111] vdd gnd cell_6t
Xbit_r112_c205 bl[205] br[205] wl[112] vdd gnd cell_6t
Xbit_r113_c205 bl[205] br[205] wl[113] vdd gnd cell_6t
Xbit_r114_c205 bl[205] br[205] wl[114] vdd gnd cell_6t
Xbit_r115_c205 bl[205] br[205] wl[115] vdd gnd cell_6t
Xbit_r116_c205 bl[205] br[205] wl[116] vdd gnd cell_6t
Xbit_r117_c205 bl[205] br[205] wl[117] vdd gnd cell_6t
Xbit_r118_c205 bl[205] br[205] wl[118] vdd gnd cell_6t
Xbit_r119_c205 bl[205] br[205] wl[119] vdd gnd cell_6t
Xbit_r120_c205 bl[205] br[205] wl[120] vdd gnd cell_6t
Xbit_r121_c205 bl[205] br[205] wl[121] vdd gnd cell_6t
Xbit_r122_c205 bl[205] br[205] wl[122] vdd gnd cell_6t
Xbit_r123_c205 bl[205] br[205] wl[123] vdd gnd cell_6t
Xbit_r124_c205 bl[205] br[205] wl[124] vdd gnd cell_6t
Xbit_r125_c205 bl[205] br[205] wl[125] vdd gnd cell_6t
Xbit_r126_c205 bl[205] br[205] wl[126] vdd gnd cell_6t
Xbit_r127_c205 bl[205] br[205] wl[127] vdd gnd cell_6t
Xbit_r0_c206 bl[206] br[206] wl[0] vdd gnd cell_6t
Xbit_r1_c206 bl[206] br[206] wl[1] vdd gnd cell_6t
Xbit_r2_c206 bl[206] br[206] wl[2] vdd gnd cell_6t
Xbit_r3_c206 bl[206] br[206] wl[3] vdd gnd cell_6t
Xbit_r4_c206 bl[206] br[206] wl[4] vdd gnd cell_6t
Xbit_r5_c206 bl[206] br[206] wl[5] vdd gnd cell_6t
Xbit_r6_c206 bl[206] br[206] wl[6] vdd gnd cell_6t
Xbit_r7_c206 bl[206] br[206] wl[7] vdd gnd cell_6t
Xbit_r8_c206 bl[206] br[206] wl[8] vdd gnd cell_6t
Xbit_r9_c206 bl[206] br[206] wl[9] vdd gnd cell_6t
Xbit_r10_c206 bl[206] br[206] wl[10] vdd gnd cell_6t
Xbit_r11_c206 bl[206] br[206] wl[11] vdd gnd cell_6t
Xbit_r12_c206 bl[206] br[206] wl[12] vdd gnd cell_6t
Xbit_r13_c206 bl[206] br[206] wl[13] vdd gnd cell_6t
Xbit_r14_c206 bl[206] br[206] wl[14] vdd gnd cell_6t
Xbit_r15_c206 bl[206] br[206] wl[15] vdd gnd cell_6t
Xbit_r16_c206 bl[206] br[206] wl[16] vdd gnd cell_6t
Xbit_r17_c206 bl[206] br[206] wl[17] vdd gnd cell_6t
Xbit_r18_c206 bl[206] br[206] wl[18] vdd gnd cell_6t
Xbit_r19_c206 bl[206] br[206] wl[19] vdd gnd cell_6t
Xbit_r20_c206 bl[206] br[206] wl[20] vdd gnd cell_6t
Xbit_r21_c206 bl[206] br[206] wl[21] vdd gnd cell_6t
Xbit_r22_c206 bl[206] br[206] wl[22] vdd gnd cell_6t
Xbit_r23_c206 bl[206] br[206] wl[23] vdd gnd cell_6t
Xbit_r24_c206 bl[206] br[206] wl[24] vdd gnd cell_6t
Xbit_r25_c206 bl[206] br[206] wl[25] vdd gnd cell_6t
Xbit_r26_c206 bl[206] br[206] wl[26] vdd gnd cell_6t
Xbit_r27_c206 bl[206] br[206] wl[27] vdd gnd cell_6t
Xbit_r28_c206 bl[206] br[206] wl[28] vdd gnd cell_6t
Xbit_r29_c206 bl[206] br[206] wl[29] vdd gnd cell_6t
Xbit_r30_c206 bl[206] br[206] wl[30] vdd gnd cell_6t
Xbit_r31_c206 bl[206] br[206] wl[31] vdd gnd cell_6t
Xbit_r32_c206 bl[206] br[206] wl[32] vdd gnd cell_6t
Xbit_r33_c206 bl[206] br[206] wl[33] vdd gnd cell_6t
Xbit_r34_c206 bl[206] br[206] wl[34] vdd gnd cell_6t
Xbit_r35_c206 bl[206] br[206] wl[35] vdd gnd cell_6t
Xbit_r36_c206 bl[206] br[206] wl[36] vdd gnd cell_6t
Xbit_r37_c206 bl[206] br[206] wl[37] vdd gnd cell_6t
Xbit_r38_c206 bl[206] br[206] wl[38] vdd gnd cell_6t
Xbit_r39_c206 bl[206] br[206] wl[39] vdd gnd cell_6t
Xbit_r40_c206 bl[206] br[206] wl[40] vdd gnd cell_6t
Xbit_r41_c206 bl[206] br[206] wl[41] vdd gnd cell_6t
Xbit_r42_c206 bl[206] br[206] wl[42] vdd gnd cell_6t
Xbit_r43_c206 bl[206] br[206] wl[43] vdd gnd cell_6t
Xbit_r44_c206 bl[206] br[206] wl[44] vdd gnd cell_6t
Xbit_r45_c206 bl[206] br[206] wl[45] vdd gnd cell_6t
Xbit_r46_c206 bl[206] br[206] wl[46] vdd gnd cell_6t
Xbit_r47_c206 bl[206] br[206] wl[47] vdd gnd cell_6t
Xbit_r48_c206 bl[206] br[206] wl[48] vdd gnd cell_6t
Xbit_r49_c206 bl[206] br[206] wl[49] vdd gnd cell_6t
Xbit_r50_c206 bl[206] br[206] wl[50] vdd gnd cell_6t
Xbit_r51_c206 bl[206] br[206] wl[51] vdd gnd cell_6t
Xbit_r52_c206 bl[206] br[206] wl[52] vdd gnd cell_6t
Xbit_r53_c206 bl[206] br[206] wl[53] vdd gnd cell_6t
Xbit_r54_c206 bl[206] br[206] wl[54] vdd gnd cell_6t
Xbit_r55_c206 bl[206] br[206] wl[55] vdd gnd cell_6t
Xbit_r56_c206 bl[206] br[206] wl[56] vdd gnd cell_6t
Xbit_r57_c206 bl[206] br[206] wl[57] vdd gnd cell_6t
Xbit_r58_c206 bl[206] br[206] wl[58] vdd gnd cell_6t
Xbit_r59_c206 bl[206] br[206] wl[59] vdd gnd cell_6t
Xbit_r60_c206 bl[206] br[206] wl[60] vdd gnd cell_6t
Xbit_r61_c206 bl[206] br[206] wl[61] vdd gnd cell_6t
Xbit_r62_c206 bl[206] br[206] wl[62] vdd gnd cell_6t
Xbit_r63_c206 bl[206] br[206] wl[63] vdd gnd cell_6t
Xbit_r64_c206 bl[206] br[206] wl[64] vdd gnd cell_6t
Xbit_r65_c206 bl[206] br[206] wl[65] vdd gnd cell_6t
Xbit_r66_c206 bl[206] br[206] wl[66] vdd gnd cell_6t
Xbit_r67_c206 bl[206] br[206] wl[67] vdd gnd cell_6t
Xbit_r68_c206 bl[206] br[206] wl[68] vdd gnd cell_6t
Xbit_r69_c206 bl[206] br[206] wl[69] vdd gnd cell_6t
Xbit_r70_c206 bl[206] br[206] wl[70] vdd gnd cell_6t
Xbit_r71_c206 bl[206] br[206] wl[71] vdd gnd cell_6t
Xbit_r72_c206 bl[206] br[206] wl[72] vdd gnd cell_6t
Xbit_r73_c206 bl[206] br[206] wl[73] vdd gnd cell_6t
Xbit_r74_c206 bl[206] br[206] wl[74] vdd gnd cell_6t
Xbit_r75_c206 bl[206] br[206] wl[75] vdd gnd cell_6t
Xbit_r76_c206 bl[206] br[206] wl[76] vdd gnd cell_6t
Xbit_r77_c206 bl[206] br[206] wl[77] vdd gnd cell_6t
Xbit_r78_c206 bl[206] br[206] wl[78] vdd gnd cell_6t
Xbit_r79_c206 bl[206] br[206] wl[79] vdd gnd cell_6t
Xbit_r80_c206 bl[206] br[206] wl[80] vdd gnd cell_6t
Xbit_r81_c206 bl[206] br[206] wl[81] vdd gnd cell_6t
Xbit_r82_c206 bl[206] br[206] wl[82] vdd gnd cell_6t
Xbit_r83_c206 bl[206] br[206] wl[83] vdd gnd cell_6t
Xbit_r84_c206 bl[206] br[206] wl[84] vdd gnd cell_6t
Xbit_r85_c206 bl[206] br[206] wl[85] vdd gnd cell_6t
Xbit_r86_c206 bl[206] br[206] wl[86] vdd gnd cell_6t
Xbit_r87_c206 bl[206] br[206] wl[87] vdd gnd cell_6t
Xbit_r88_c206 bl[206] br[206] wl[88] vdd gnd cell_6t
Xbit_r89_c206 bl[206] br[206] wl[89] vdd gnd cell_6t
Xbit_r90_c206 bl[206] br[206] wl[90] vdd gnd cell_6t
Xbit_r91_c206 bl[206] br[206] wl[91] vdd gnd cell_6t
Xbit_r92_c206 bl[206] br[206] wl[92] vdd gnd cell_6t
Xbit_r93_c206 bl[206] br[206] wl[93] vdd gnd cell_6t
Xbit_r94_c206 bl[206] br[206] wl[94] vdd gnd cell_6t
Xbit_r95_c206 bl[206] br[206] wl[95] vdd gnd cell_6t
Xbit_r96_c206 bl[206] br[206] wl[96] vdd gnd cell_6t
Xbit_r97_c206 bl[206] br[206] wl[97] vdd gnd cell_6t
Xbit_r98_c206 bl[206] br[206] wl[98] vdd gnd cell_6t
Xbit_r99_c206 bl[206] br[206] wl[99] vdd gnd cell_6t
Xbit_r100_c206 bl[206] br[206] wl[100] vdd gnd cell_6t
Xbit_r101_c206 bl[206] br[206] wl[101] vdd gnd cell_6t
Xbit_r102_c206 bl[206] br[206] wl[102] vdd gnd cell_6t
Xbit_r103_c206 bl[206] br[206] wl[103] vdd gnd cell_6t
Xbit_r104_c206 bl[206] br[206] wl[104] vdd gnd cell_6t
Xbit_r105_c206 bl[206] br[206] wl[105] vdd gnd cell_6t
Xbit_r106_c206 bl[206] br[206] wl[106] vdd gnd cell_6t
Xbit_r107_c206 bl[206] br[206] wl[107] vdd gnd cell_6t
Xbit_r108_c206 bl[206] br[206] wl[108] vdd gnd cell_6t
Xbit_r109_c206 bl[206] br[206] wl[109] vdd gnd cell_6t
Xbit_r110_c206 bl[206] br[206] wl[110] vdd gnd cell_6t
Xbit_r111_c206 bl[206] br[206] wl[111] vdd gnd cell_6t
Xbit_r112_c206 bl[206] br[206] wl[112] vdd gnd cell_6t
Xbit_r113_c206 bl[206] br[206] wl[113] vdd gnd cell_6t
Xbit_r114_c206 bl[206] br[206] wl[114] vdd gnd cell_6t
Xbit_r115_c206 bl[206] br[206] wl[115] vdd gnd cell_6t
Xbit_r116_c206 bl[206] br[206] wl[116] vdd gnd cell_6t
Xbit_r117_c206 bl[206] br[206] wl[117] vdd gnd cell_6t
Xbit_r118_c206 bl[206] br[206] wl[118] vdd gnd cell_6t
Xbit_r119_c206 bl[206] br[206] wl[119] vdd gnd cell_6t
Xbit_r120_c206 bl[206] br[206] wl[120] vdd gnd cell_6t
Xbit_r121_c206 bl[206] br[206] wl[121] vdd gnd cell_6t
Xbit_r122_c206 bl[206] br[206] wl[122] vdd gnd cell_6t
Xbit_r123_c206 bl[206] br[206] wl[123] vdd gnd cell_6t
Xbit_r124_c206 bl[206] br[206] wl[124] vdd gnd cell_6t
Xbit_r125_c206 bl[206] br[206] wl[125] vdd gnd cell_6t
Xbit_r126_c206 bl[206] br[206] wl[126] vdd gnd cell_6t
Xbit_r127_c206 bl[206] br[206] wl[127] vdd gnd cell_6t
Xbit_r0_c207 bl[207] br[207] wl[0] vdd gnd cell_6t
Xbit_r1_c207 bl[207] br[207] wl[1] vdd gnd cell_6t
Xbit_r2_c207 bl[207] br[207] wl[2] vdd gnd cell_6t
Xbit_r3_c207 bl[207] br[207] wl[3] vdd gnd cell_6t
Xbit_r4_c207 bl[207] br[207] wl[4] vdd gnd cell_6t
Xbit_r5_c207 bl[207] br[207] wl[5] vdd gnd cell_6t
Xbit_r6_c207 bl[207] br[207] wl[6] vdd gnd cell_6t
Xbit_r7_c207 bl[207] br[207] wl[7] vdd gnd cell_6t
Xbit_r8_c207 bl[207] br[207] wl[8] vdd gnd cell_6t
Xbit_r9_c207 bl[207] br[207] wl[9] vdd gnd cell_6t
Xbit_r10_c207 bl[207] br[207] wl[10] vdd gnd cell_6t
Xbit_r11_c207 bl[207] br[207] wl[11] vdd gnd cell_6t
Xbit_r12_c207 bl[207] br[207] wl[12] vdd gnd cell_6t
Xbit_r13_c207 bl[207] br[207] wl[13] vdd gnd cell_6t
Xbit_r14_c207 bl[207] br[207] wl[14] vdd gnd cell_6t
Xbit_r15_c207 bl[207] br[207] wl[15] vdd gnd cell_6t
Xbit_r16_c207 bl[207] br[207] wl[16] vdd gnd cell_6t
Xbit_r17_c207 bl[207] br[207] wl[17] vdd gnd cell_6t
Xbit_r18_c207 bl[207] br[207] wl[18] vdd gnd cell_6t
Xbit_r19_c207 bl[207] br[207] wl[19] vdd gnd cell_6t
Xbit_r20_c207 bl[207] br[207] wl[20] vdd gnd cell_6t
Xbit_r21_c207 bl[207] br[207] wl[21] vdd gnd cell_6t
Xbit_r22_c207 bl[207] br[207] wl[22] vdd gnd cell_6t
Xbit_r23_c207 bl[207] br[207] wl[23] vdd gnd cell_6t
Xbit_r24_c207 bl[207] br[207] wl[24] vdd gnd cell_6t
Xbit_r25_c207 bl[207] br[207] wl[25] vdd gnd cell_6t
Xbit_r26_c207 bl[207] br[207] wl[26] vdd gnd cell_6t
Xbit_r27_c207 bl[207] br[207] wl[27] vdd gnd cell_6t
Xbit_r28_c207 bl[207] br[207] wl[28] vdd gnd cell_6t
Xbit_r29_c207 bl[207] br[207] wl[29] vdd gnd cell_6t
Xbit_r30_c207 bl[207] br[207] wl[30] vdd gnd cell_6t
Xbit_r31_c207 bl[207] br[207] wl[31] vdd gnd cell_6t
Xbit_r32_c207 bl[207] br[207] wl[32] vdd gnd cell_6t
Xbit_r33_c207 bl[207] br[207] wl[33] vdd gnd cell_6t
Xbit_r34_c207 bl[207] br[207] wl[34] vdd gnd cell_6t
Xbit_r35_c207 bl[207] br[207] wl[35] vdd gnd cell_6t
Xbit_r36_c207 bl[207] br[207] wl[36] vdd gnd cell_6t
Xbit_r37_c207 bl[207] br[207] wl[37] vdd gnd cell_6t
Xbit_r38_c207 bl[207] br[207] wl[38] vdd gnd cell_6t
Xbit_r39_c207 bl[207] br[207] wl[39] vdd gnd cell_6t
Xbit_r40_c207 bl[207] br[207] wl[40] vdd gnd cell_6t
Xbit_r41_c207 bl[207] br[207] wl[41] vdd gnd cell_6t
Xbit_r42_c207 bl[207] br[207] wl[42] vdd gnd cell_6t
Xbit_r43_c207 bl[207] br[207] wl[43] vdd gnd cell_6t
Xbit_r44_c207 bl[207] br[207] wl[44] vdd gnd cell_6t
Xbit_r45_c207 bl[207] br[207] wl[45] vdd gnd cell_6t
Xbit_r46_c207 bl[207] br[207] wl[46] vdd gnd cell_6t
Xbit_r47_c207 bl[207] br[207] wl[47] vdd gnd cell_6t
Xbit_r48_c207 bl[207] br[207] wl[48] vdd gnd cell_6t
Xbit_r49_c207 bl[207] br[207] wl[49] vdd gnd cell_6t
Xbit_r50_c207 bl[207] br[207] wl[50] vdd gnd cell_6t
Xbit_r51_c207 bl[207] br[207] wl[51] vdd gnd cell_6t
Xbit_r52_c207 bl[207] br[207] wl[52] vdd gnd cell_6t
Xbit_r53_c207 bl[207] br[207] wl[53] vdd gnd cell_6t
Xbit_r54_c207 bl[207] br[207] wl[54] vdd gnd cell_6t
Xbit_r55_c207 bl[207] br[207] wl[55] vdd gnd cell_6t
Xbit_r56_c207 bl[207] br[207] wl[56] vdd gnd cell_6t
Xbit_r57_c207 bl[207] br[207] wl[57] vdd gnd cell_6t
Xbit_r58_c207 bl[207] br[207] wl[58] vdd gnd cell_6t
Xbit_r59_c207 bl[207] br[207] wl[59] vdd gnd cell_6t
Xbit_r60_c207 bl[207] br[207] wl[60] vdd gnd cell_6t
Xbit_r61_c207 bl[207] br[207] wl[61] vdd gnd cell_6t
Xbit_r62_c207 bl[207] br[207] wl[62] vdd gnd cell_6t
Xbit_r63_c207 bl[207] br[207] wl[63] vdd gnd cell_6t
Xbit_r64_c207 bl[207] br[207] wl[64] vdd gnd cell_6t
Xbit_r65_c207 bl[207] br[207] wl[65] vdd gnd cell_6t
Xbit_r66_c207 bl[207] br[207] wl[66] vdd gnd cell_6t
Xbit_r67_c207 bl[207] br[207] wl[67] vdd gnd cell_6t
Xbit_r68_c207 bl[207] br[207] wl[68] vdd gnd cell_6t
Xbit_r69_c207 bl[207] br[207] wl[69] vdd gnd cell_6t
Xbit_r70_c207 bl[207] br[207] wl[70] vdd gnd cell_6t
Xbit_r71_c207 bl[207] br[207] wl[71] vdd gnd cell_6t
Xbit_r72_c207 bl[207] br[207] wl[72] vdd gnd cell_6t
Xbit_r73_c207 bl[207] br[207] wl[73] vdd gnd cell_6t
Xbit_r74_c207 bl[207] br[207] wl[74] vdd gnd cell_6t
Xbit_r75_c207 bl[207] br[207] wl[75] vdd gnd cell_6t
Xbit_r76_c207 bl[207] br[207] wl[76] vdd gnd cell_6t
Xbit_r77_c207 bl[207] br[207] wl[77] vdd gnd cell_6t
Xbit_r78_c207 bl[207] br[207] wl[78] vdd gnd cell_6t
Xbit_r79_c207 bl[207] br[207] wl[79] vdd gnd cell_6t
Xbit_r80_c207 bl[207] br[207] wl[80] vdd gnd cell_6t
Xbit_r81_c207 bl[207] br[207] wl[81] vdd gnd cell_6t
Xbit_r82_c207 bl[207] br[207] wl[82] vdd gnd cell_6t
Xbit_r83_c207 bl[207] br[207] wl[83] vdd gnd cell_6t
Xbit_r84_c207 bl[207] br[207] wl[84] vdd gnd cell_6t
Xbit_r85_c207 bl[207] br[207] wl[85] vdd gnd cell_6t
Xbit_r86_c207 bl[207] br[207] wl[86] vdd gnd cell_6t
Xbit_r87_c207 bl[207] br[207] wl[87] vdd gnd cell_6t
Xbit_r88_c207 bl[207] br[207] wl[88] vdd gnd cell_6t
Xbit_r89_c207 bl[207] br[207] wl[89] vdd gnd cell_6t
Xbit_r90_c207 bl[207] br[207] wl[90] vdd gnd cell_6t
Xbit_r91_c207 bl[207] br[207] wl[91] vdd gnd cell_6t
Xbit_r92_c207 bl[207] br[207] wl[92] vdd gnd cell_6t
Xbit_r93_c207 bl[207] br[207] wl[93] vdd gnd cell_6t
Xbit_r94_c207 bl[207] br[207] wl[94] vdd gnd cell_6t
Xbit_r95_c207 bl[207] br[207] wl[95] vdd gnd cell_6t
Xbit_r96_c207 bl[207] br[207] wl[96] vdd gnd cell_6t
Xbit_r97_c207 bl[207] br[207] wl[97] vdd gnd cell_6t
Xbit_r98_c207 bl[207] br[207] wl[98] vdd gnd cell_6t
Xbit_r99_c207 bl[207] br[207] wl[99] vdd gnd cell_6t
Xbit_r100_c207 bl[207] br[207] wl[100] vdd gnd cell_6t
Xbit_r101_c207 bl[207] br[207] wl[101] vdd gnd cell_6t
Xbit_r102_c207 bl[207] br[207] wl[102] vdd gnd cell_6t
Xbit_r103_c207 bl[207] br[207] wl[103] vdd gnd cell_6t
Xbit_r104_c207 bl[207] br[207] wl[104] vdd gnd cell_6t
Xbit_r105_c207 bl[207] br[207] wl[105] vdd gnd cell_6t
Xbit_r106_c207 bl[207] br[207] wl[106] vdd gnd cell_6t
Xbit_r107_c207 bl[207] br[207] wl[107] vdd gnd cell_6t
Xbit_r108_c207 bl[207] br[207] wl[108] vdd gnd cell_6t
Xbit_r109_c207 bl[207] br[207] wl[109] vdd gnd cell_6t
Xbit_r110_c207 bl[207] br[207] wl[110] vdd gnd cell_6t
Xbit_r111_c207 bl[207] br[207] wl[111] vdd gnd cell_6t
Xbit_r112_c207 bl[207] br[207] wl[112] vdd gnd cell_6t
Xbit_r113_c207 bl[207] br[207] wl[113] vdd gnd cell_6t
Xbit_r114_c207 bl[207] br[207] wl[114] vdd gnd cell_6t
Xbit_r115_c207 bl[207] br[207] wl[115] vdd gnd cell_6t
Xbit_r116_c207 bl[207] br[207] wl[116] vdd gnd cell_6t
Xbit_r117_c207 bl[207] br[207] wl[117] vdd gnd cell_6t
Xbit_r118_c207 bl[207] br[207] wl[118] vdd gnd cell_6t
Xbit_r119_c207 bl[207] br[207] wl[119] vdd gnd cell_6t
Xbit_r120_c207 bl[207] br[207] wl[120] vdd gnd cell_6t
Xbit_r121_c207 bl[207] br[207] wl[121] vdd gnd cell_6t
Xbit_r122_c207 bl[207] br[207] wl[122] vdd gnd cell_6t
Xbit_r123_c207 bl[207] br[207] wl[123] vdd gnd cell_6t
Xbit_r124_c207 bl[207] br[207] wl[124] vdd gnd cell_6t
Xbit_r125_c207 bl[207] br[207] wl[125] vdd gnd cell_6t
Xbit_r126_c207 bl[207] br[207] wl[126] vdd gnd cell_6t
Xbit_r127_c207 bl[207] br[207] wl[127] vdd gnd cell_6t
Xbit_r0_c208 bl[208] br[208] wl[0] vdd gnd cell_6t
Xbit_r1_c208 bl[208] br[208] wl[1] vdd gnd cell_6t
Xbit_r2_c208 bl[208] br[208] wl[2] vdd gnd cell_6t
Xbit_r3_c208 bl[208] br[208] wl[3] vdd gnd cell_6t
Xbit_r4_c208 bl[208] br[208] wl[4] vdd gnd cell_6t
Xbit_r5_c208 bl[208] br[208] wl[5] vdd gnd cell_6t
Xbit_r6_c208 bl[208] br[208] wl[6] vdd gnd cell_6t
Xbit_r7_c208 bl[208] br[208] wl[7] vdd gnd cell_6t
Xbit_r8_c208 bl[208] br[208] wl[8] vdd gnd cell_6t
Xbit_r9_c208 bl[208] br[208] wl[9] vdd gnd cell_6t
Xbit_r10_c208 bl[208] br[208] wl[10] vdd gnd cell_6t
Xbit_r11_c208 bl[208] br[208] wl[11] vdd gnd cell_6t
Xbit_r12_c208 bl[208] br[208] wl[12] vdd gnd cell_6t
Xbit_r13_c208 bl[208] br[208] wl[13] vdd gnd cell_6t
Xbit_r14_c208 bl[208] br[208] wl[14] vdd gnd cell_6t
Xbit_r15_c208 bl[208] br[208] wl[15] vdd gnd cell_6t
Xbit_r16_c208 bl[208] br[208] wl[16] vdd gnd cell_6t
Xbit_r17_c208 bl[208] br[208] wl[17] vdd gnd cell_6t
Xbit_r18_c208 bl[208] br[208] wl[18] vdd gnd cell_6t
Xbit_r19_c208 bl[208] br[208] wl[19] vdd gnd cell_6t
Xbit_r20_c208 bl[208] br[208] wl[20] vdd gnd cell_6t
Xbit_r21_c208 bl[208] br[208] wl[21] vdd gnd cell_6t
Xbit_r22_c208 bl[208] br[208] wl[22] vdd gnd cell_6t
Xbit_r23_c208 bl[208] br[208] wl[23] vdd gnd cell_6t
Xbit_r24_c208 bl[208] br[208] wl[24] vdd gnd cell_6t
Xbit_r25_c208 bl[208] br[208] wl[25] vdd gnd cell_6t
Xbit_r26_c208 bl[208] br[208] wl[26] vdd gnd cell_6t
Xbit_r27_c208 bl[208] br[208] wl[27] vdd gnd cell_6t
Xbit_r28_c208 bl[208] br[208] wl[28] vdd gnd cell_6t
Xbit_r29_c208 bl[208] br[208] wl[29] vdd gnd cell_6t
Xbit_r30_c208 bl[208] br[208] wl[30] vdd gnd cell_6t
Xbit_r31_c208 bl[208] br[208] wl[31] vdd gnd cell_6t
Xbit_r32_c208 bl[208] br[208] wl[32] vdd gnd cell_6t
Xbit_r33_c208 bl[208] br[208] wl[33] vdd gnd cell_6t
Xbit_r34_c208 bl[208] br[208] wl[34] vdd gnd cell_6t
Xbit_r35_c208 bl[208] br[208] wl[35] vdd gnd cell_6t
Xbit_r36_c208 bl[208] br[208] wl[36] vdd gnd cell_6t
Xbit_r37_c208 bl[208] br[208] wl[37] vdd gnd cell_6t
Xbit_r38_c208 bl[208] br[208] wl[38] vdd gnd cell_6t
Xbit_r39_c208 bl[208] br[208] wl[39] vdd gnd cell_6t
Xbit_r40_c208 bl[208] br[208] wl[40] vdd gnd cell_6t
Xbit_r41_c208 bl[208] br[208] wl[41] vdd gnd cell_6t
Xbit_r42_c208 bl[208] br[208] wl[42] vdd gnd cell_6t
Xbit_r43_c208 bl[208] br[208] wl[43] vdd gnd cell_6t
Xbit_r44_c208 bl[208] br[208] wl[44] vdd gnd cell_6t
Xbit_r45_c208 bl[208] br[208] wl[45] vdd gnd cell_6t
Xbit_r46_c208 bl[208] br[208] wl[46] vdd gnd cell_6t
Xbit_r47_c208 bl[208] br[208] wl[47] vdd gnd cell_6t
Xbit_r48_c208 bl[208] br[208] wl[48] vdd gnd cell_6t
Xbit_r49_c208 bl[208] br[208] wl[49] vdd gnd cell_6t
Xbit_r50_c208 bl[208] br[208] wl[50] vdd gnd cell_6t
Xbit_r51_c208 bl[208] br[208] wl[51] vdd gnd cell_6t
Xbit_r52_c208 bl[208] br[208] wl[52] vdd gnd cell_6t
Xbit_r53_c208 bl[208] br[208] wl[53] vdd gnd cell_6t
Xbit_r54_c208 bl[208] br[208] wl[54] vdd gnd cell_6t
Xbit_r55_c208 bl[208] br[208] wl[55] vdd gnd cell_6t
Xbit_r56_c208 bl[208] br[208] wl[56] vdd gnd cell_6t
Xbit_r57_c208 bl[208] br[208] wl[57] vdd gnd cell_6t
Xbit_r58_c208 bl[208] br[208] wl[58] vdd gnd cell_6t
Xbit_r59_c208 bl[208] br[208] wl[59] vdd gnd cell_6t
Xbit_r60_c208 bl[208] br[208] wl[60] vdd gnd cell_6t
Xbit_r61_c208 bl[208] br[208] wl[61] vdd gnd cell_6t
Xbit_r62_c208 bl[208] br[208] wl[62] vdd gnd cell_6t
Xbit_r63_c208 bl[208] br[208] wl[63] vdd gnd cell_6t
Xbit_r64_c208 bl[208] br[208] wl[64] vdd gnd cell_6t
Xbit_r65_c208 bl[208] br[208] wl[65] vdd gnd cell_6t
Xbit_r66_c208 bl[208] br[208] wl[66] vdd gnd cell_6t
Xbit_r67_c208 bl[208] br[208] wl[67] vdd gnd cell_6t
Xbit_r68_c208 bl[208] br[208] wl[68] vdd gnd cell_6t
Xbit_r69_c208 bl[208] br[208] wl[69] vdd gnd cell_6t
Xbit_r70_c208 bl[208] br[208] wl[70] vdd gnd cell_6t
Xbit_r71_c208 bl[208] br[208] wl[71] vdd gnd cell_6t
Xbit_r72_c208 bl[208] br[208] wl[72] vdd gnd cell_6t
Xbit_r73_c208 bl[208] br[208] wl[73] vdd gnd cell_6t
Xbit_r74_c208 bl[208] br[208] wl[74] vdd gnd cell_6t
Xbit_r75_c208 bl[208] br[208] wl[75] vdd gnd cell_6t
Xbit_r76_c208 bl[208] br[208] wl[76] vdd gnd cell_6t
Xbit_r77_c208 bl[208] br[208] wl[77] vdd gnd cell_6t
Xbit_r78_c208 bl[208] br[208] wl[78] vdd gnd cell_6t
Xbit_r79_c208 bl[208] br[208] wl[79] vdd gnd cell_6t
Xbit_r80_c208 bl[208] br[208] wl[80] vdd gnd cell_6t
Xbit_r81_c208 bl[208] br[208] wl[81] vdd gnd cell_6t
Xbit_r82_c208 bl[208] br[208] wl[82] vdd gnd cell_6t
Xbit_r83_c208 bl[208] br[208] wl[83] vdd gnd cell_6t
Xbit_r84_c208 bl[208] br[208] wl[84] vdd gnd cell_6t
Xbit_r85_c208 bl[208] br[208] wl[85] vdd gnd cell_6t
Xbit_r86_c208 bl[208] br[208] wl[86] vdd gnd cell_6t
Xbit_r87_c208 bl[208] br[208] wl[87] vdd gnd cell_6t
Xbit_r88_c208 bl[208] br[208] wl[88] vdd gnd cell_6t
Xbit_r89_c208 bl[208] br[208] wl[89] vdd gnd cell_6t
Xbit_r90_c208 bl[208] br[208] wl[90] vdd gnd cell_6t
Xbit_r91_c208 bl[208] br[208] wl[91] vdd gnd cell_6t
Xbit_r92_c208 bl[208] br[208] wl[92] vdd gnd cell_6t
Xbit_r93_c208 bl[208] br[208] wl[93] vdd gnd cell_6t
Xbit_r94_c208 bl[208] br[208] wl[94] vdd gnd cell_6t
Xbit_r95_c208 bl[208] br[208] wl[95] vdd gnd cell_6t
Xbit_r96_c208 bl[208] br[208] wl[96] vdd gnd cell_6t
Xbit_r97_c208 bl[208] br[208] wl[97] vdd gnd cell_6t
Xbit_r98_c208 bl[208] br[208] wl[98] vdd gnd cell_6t
Xbit_r99_c208 bl[208] br[208] wl[99] vdd gnd cell_6t
Xbit_r100_c208 bl[208] br[208] wl[100] vdd gnd cell_6t
Xbit_r101_c208 bl[208] br[208] wl[101] vdd gnd cell_6t
Xbit_r102_c208 bl[208] br[208] wl[102] vdd gnd cell_6t
Xbit_r103_c208 bl[208] br[208] wl[103] vdd gnd cell_6t
Xbit_r104_c208 bl[208] br[208] wl[104] vdd gnd cell_6t
Xbit_r105_c208 bl[208] br[208] wl[105] vdd gnd cell_6t
Xbit_r106_c208 bl[208] br[208] wl[106] vdd gnd cell_6t
Xbit_r107_c208 bl[208] br[208] wl[107] vdd gnd cell_6t
Xbit_r108_c208 bl[208] br[208] wl[108] vdd gnd cell_6t
Xbit_r109_c208 bl[208] br[208] wl[109] vdd gnd cell_6t
Xbit_r110_c208 bl[208] br[208] wl[110] vdd gnd cell_6t
Xbit_r111_c208 bl[208] br[208] wl[111] vdd gnd cell_6t
Xbit_r112_c208 bl[208] br[208] wl[112] vdd gnd cell_6t
Xbit_r113_c208 bl[208] br[208] wl[113] vdd gnd cell_6t
Xbit_r114_c208 bl[208] br[208] wl[114] vdd gnd cell_6t
Xbit_r115_c208 bl[208] br[208] wl[115] vdd gnd cell_6t
Xbit_r116_c208 bl[208] br[208] wl[116] vdd gnd cell_6t
Xbit_r117_c208 bl[208] br[208] wl[117] vdd gnd cell_6t
Xbit_r118_c208 bl[208] br[208] wl[118] vdd gnd cell_6t
Xbit_r119_c208 bl[208] br[208] wl[119] vdd gnd cell_6t
Xbit_r120_c208 bl[208] br[208] wl[120] vdd gnd cell_6t
Xbit_r121_c208 bl[208] br[208] wl[121] vdd gnd cell_6t
Xbit_r122_c208 bl[208] br[208] wl[122] vdd gnd cell_6t
Xbit_r123_c208 bl[208] br[208] wl[123] vdd gnd cell_6t
Xbit_r124_c208 bl[208] br[208] wl[124] vdd gnd cell_6t
Xbit_r125_c208 bl[208] br[208] wl[125] vdd gnd cell_6t
Xbit_r126_c208 bl[208] br[208] wl[126] vdd gnd cell_6t
Xbit_r127_c208 bl[208] br[208] wl[127] vdd gnd cell_6t
Xbit_r0_c209 bl[209] br[209] wl[0] vdd gnd cell_6t
Xbit_r1_c209 bl[209] br[209] wl[1] vdd gnd cell_6t
Xbit_r2_c209 bl[209] br[209] wl[2] vdd gnd cell_6t
Xbit_r3_c209 bl[209] br[209] wl[3] vdd gnd cell_6t
Xbit_r4_c209 bl[209] br[209] wl[4] vdd gnd cell_6t
Xbit_r5_c209 bl[209] br[209] wl[5] vdd gnd cell_6t
Xbit_r6_c209 bl[209] br[209] wl[6] vdd gnd cell_6t
Xbit_r7_c209 bl[209] br[209] wl[7] vdd gnd cell_6t
Xbit_r8_c209 bl[209] br[209] wl[8] vdd gnd cell_6t
Xbit_r9_c209 bl[209] br[209] wl[9] vdd gnd cell_6t
Xbit_r10_c209 bl[209] br[209] wl[10] vdd gnd cell_6t
Xbit_r11_c209 bl[209] br[209] wl[11] vdd gnd cell_6t
Xbit_r12_c209 bl[209] br[209] wl[12] vdd gnd cell_6t
Xbit_r13_c209 bl[209] br[209] wl[13] vdd gnd cell_6t
Xbit_r14_c209 bl[209] br[209] wl[14] vdd gnd cell_6t
Xbit_r15_c209 bl[209] br[209] wl[15] vdd gnd cell_6t
Xbit_r16_c209 bl[209] br[209] wl[16] vdd gnd cell_6t
Xbit_r17_c209 bl[209] br[209] wl[17] vdd gnd cell_6t
Xbit_r18_c209 bl[209] br[209] wl[18] vdd gnd cell_6t
Xbit_r19_c209 bl[209] br[209] wl[19] vdd gnd cell_6t
Xbit_r20_c209 bl[209] br[209] wl[20] vdd gnd cell_6t
Xbit_r21_c209 bl[209] br[209] wl[21] vdd gnd cell_6t
Xbit_r22_c209 bl[209] br[209] wl[22] vdd gnd cell_6t
Xbit_r23_c209 bl[209] br[209] wl[23] vdd gnd cell_6t
Xbit_r24_c209 bl[209] br[209] wl[24] vdd gnd cell_6t
Xbit_r25_c209 bl[209] br[209] wl[25] vdd gnd cell_6t
Xbit_r26_c209 bl[209] br[209] wl[26] vdd gnd cell_6t
Xbit_r27_c209 bl[209] br[209] wl[27] vdd gnd cell_6t
Xbit_r28_c209 bl[209] br[209] wl[28] vdd gnd cell_6t
Xbit_r29_c209 bl[209] br[209] wl[29] vdd gnd cell_6t
Xbit_r30_c209 bl[209] br[209] wl[30] vdd gnd cell_6t
Xbit_r31_c209 bl[209] br[209] wl[31] vdd gnd cell_6t
Xbit_r32_c209 bl[209] br[209] wl[32] vdd gnd cell_6t
Xbit_r33_c209 bl[209] br[209] wl[33] vdd gnd cell_6t
Xbit_r34_c209 bl[209] br[209] wl[34] vdd gnd cell_6t
Xbit_r35_c209 bl[209] br[209] wl[35] vdd gnd cell_6t
Xbit_r36_c209 bl[209] br[209] wl[36] vdd gnd cell_6t
Xbit_r37_c209 bl[209] br[209] wl[37] vdd gnd cell_6t
Xbit_r38_c209 bl[209] br[209] wl[38] vdd gnd cell_6t
Xbit_r39_c209 bl[209] br[209] wl[39] vdd gnd cell_6t
Xbit_r40_c209 bl[209] br[209] wl[40] vdd gnd cell_6t
Xbit_r41_c209 bl[209] br[209] wl[41] vdd gnd cell_6t
Xbit_r42_c209 bl[209] br[209] wl[42] vdd gnd cell_6t
Xbit_r43_c209 bl[209] br[209] wl[43] vdd gnd cell_6t
Xbit_r44_c209 bl[209] br[209] wl[44] vdd gnd cell_6t
Xbit_r45_c209 bl[209] br[209] wl[45] vdd gnd cell_6t
Xbit_r46_c209 bl[209] br[209] wl[46] vdd gnd cell_6t
Xbit_r47_c209 bl[209] br[209] wl[47] vdd gnd cell_6t
Xbit_r48_c209 bl[209] br[209] wl[48] vdd gnd cell_6t
Xbit_r49_c209 bl[209] br[209] wl[49] vdd gnd cell_6t
Xbit_r50_c209 bl[209] br[209] wl[50] vdd gnd cell_6t
Xbit_r51_c209 bl[209] br[209] wl[51] vdd gnd cell_6t
Xbit_r52_c209 bl[209] br[209] wl[52] vdd gnd cell_6t
Xbit_r53_c209 bl[209] br[209] wl[53] vdd gnd cell_6t
Xbit_r54_c209 bl[209] br[209] wl[54] vdd gnd cell_6t
Xbit_r55_c209 bl[209] br[209] wl[55] vdd gnd cell_6t
Xbit_r56_c209 bl[209] br[209] wl[56] vdd gnd cell_6t
Xbit_r57_c209 bl[209] br[209] wl[57] vdd gnd cell_6t
Xbit_r58_c209 bl[209] br[209] wl[58] vdd gnd cell_6t
Xbit_r59_c209 bl[209] br[209] wl[59] vdd gnd cell_6t
Xbit_r60_c209 bl[209] br[209] wl[60] vdd gnd cell_6t
Xbit_r61_c209 bl[209] br[209] wl[61] vdd gnd cell_6t
Xbit_r62_c209 bl[209] br[209] wl[62] vdd gnd cell_6t
Xbit_r63_c209 bl[209] br[209] wl[63] vdd gnd cell_6t
Xbit_r64_c209 bl[209] br[209] wl[64] vdd gnd cell_6t
Xbit_r65_c209 bl[209] br[209] wl[65] vdd gnd cell_6t
Xbit_r66_c209 bl[209] br[209] wl[66] vdd gnd cell_6t
Xbit_r67_c209 bl[209] br[209] wl[67] vdd gnd cell_6t
Xbit_r68_c209 bl[209] br[209] wl[68] vdd gnd cell_6t
Xbit_r69_c209 bl[209] br[209] wl[69] vdd gnd cell_6t
Xbit_r70_c209 bl[209] br[209] wl[70] vdd gnd cell_6t
Xbit_r71_c209 bl[209] br[209] wl[71] vdd gnd cell_6t
Xbit_r72_c209 bl[209] br[209] wl[72] vdd gnd cell_6t
Xbit_r73_c209 bl[209] br[209] wl[73] vdd gnd cell_6t
Xbit_r74_c209 bl[209] br[209] wl[74] vdd gnd cell_6t
Xbit_r75_c209 bl[209] br[209] wl[75] vdd gnd cell_6t
Xbit_r76_c209 bl[209] br[209] wl[76] vdd gnd cell_6t
Xbit_r77_c209 bl[209] br[209] wl[77] vdd gnd cell_6t
Xbit_r78_c209 bl[209] br[209] wl[78] vdd gnd cell_6t
Xbit_r79_c209 bl[209] br[209] wl[79] vdd gnd cell_6t
Xbit_r80_c209 bl[209] br[209] wl[80] vdd gnd cell_6t
Xbit_r81_c209 bl[209] br[209] wl[81] vdd gnd cell_6t
Xbit_r82_c209 bl[209] br[209] wl[82] vdd gnd cell_6t
Xbit_r83_c209 bl[209] br[209] wl[83] vdd gnd cell_6t
Xbit_r84_c209 bl[209] br[209] wl[84] vdd gnd cell_6t
Xbit_r85_c209 bl[209] br[209] wl[85] vdd gnd cell_6t
Xbit_r86_c209 bl[209] br[209] wl[86] vdd gnd cell_6t
Xbit_r87_c209 bl[209] br[209] wl[87] vdd gnd cell_6t
Xbit_r88_c209 bl[209] br[209] wl[88] vdd gnd cell_6t
Xbit_r89_c209 bl[209] br[209] wl[89] vdd gnd cell_6t
Xbit_r90_c209 bl[209] br[209] wl[90] vdd gnd cell_6t
Xbit_r91_c209 bl[209] br[209] wl[91] vdd gnd cell_6t
Xbit_r92_c209 bl[209] br[209] wl[92] vdd gnd cell_6t
Xbit_r93_c209 bl[209] br[209] wl[93] vdd gnd cell_6t
Xbit_r94_c209 bl[209] br[209] wl[94] vdd gnd cell_6t
Xbit_r95_c209 bl[209] br[209] wl[95] vdd gnd cell_6t
Xbit_r96_c209 bl[209] br[209] wl[96] vdd gnd cell_6t
Xbit_r97_c209 bl[209] br[209] wl[97] vdd gnd cell_6t
Xbit_r98_c209 bl[209] br[209] wl[98] vdd gnd cell_6t
Xbit_r99_c209 bl[209] br[209] wl[99] vdd gnd cell_6t
Xbit_r100_c209 bl[209] br[209] wl[100] vdd gnd cell_6t
Xbit_r101_c209 bl[209] br[209] wl[101] vdd gnd cell_6t
Xbit_r102_c209 bl[209] br[209] wl[102] vdd gnd cell_6t
Xbit_r103_c209 bl[209] br[209] wl[103] vdd gnd cell_6t
Xbit_r104_c209 bl[209] br[209] wl[104] vdd gnd cell_6t
Xbit_r105_c209 bl[209] br[209] wl[105] vdd gnd cell_6t
Xbit_r106_c209 bl[209] br[209] wl[106] vdd gnd cell_6t
Xbit_r107_c209 bl[209] br[209] wl[107] vdd gnd cell_6t
Xbit_r108_c209 bl[209] br[209] wl[108] vdd gnd cell_6t
Xbit_r109_c209 bl[209] br[209] wl[109] vdd gnd cell_6t
Xbit_r110_c209 bl[209] br[209] wl[110] vdd gnd cell_6t
Xbit_r111_c209 bl[209] br[209] wl[111] vdd gnd cell_6t
Xbit_r112_c209 bl[209] br[209] wl[112] vdd gnd cell_6t
Xbit_r113_c209 bl[209] br[209] wl[113] vdd gnd cell_6t
Xbit_r114_c209 bl[209] br[209] wl[114] vdd gnd cell_6t
Xbit_r115_c209 bl[209] br[209] wl[115] vdd gnd cell_6t
Xbit_r116_c209 bl[209] br[209] wl[116] vdd gnd cell_6t
Xbit_r117_c209 bl[209] br[209] wl[117] vdd gnd cell_6t
Xbit_r118_c209 bl[209] br[209] wl[118] vdd gnd cell_6t
Xbit_r119_c209 bl[209] br[209] wl[119] vdd gnd cell_6t
Xbit_r120_c209 bl[209] br[209] wl[120] vdd gnd cell_6t
Xbit_r121_c209 bl[209] br[209] wl[121] vdd gnd cell_6t
Xbit_r122_c209 bl[209] br[209] wl[122] vdd gnd cell_6t
Xbit_r123_c209 bl[209] br[209] wl[123] vdd gnd cell_6t
Xbit_r124_c209 bl[209] br[209] wl[124] vdd gnd cell_6t
Xbit_r125_c209 bl[209] br[209] wl[125] vdd gnd cell_6t
Xbit_r126_c209 bl[209] br[209] wl[126] vdd gnd cell_6t
Xbit_r127_c209 bl[209] br[209] wl[127] vdd gnd cell_6t
Xbit_r0_c210 bl[210] br[210] wl[0] vdd gnd cell_6t
Xbit_r1_c210 bl[210] br[210] wl[1] vdd gnd cell_6t
Xbit_r2_c210 bl[210] br[210] wl[2] vdd gnd cell_6t
Xbit_r3_c210 bl[210] br[210] wl[3] vdd gnd cell_6t
Xbit_r4_c210 bl[210] br[210] wl[4] vdd gnd cell_6t
Xbit_r5_c210 bl[210] br[210] wl[5] vdd gnd cell_6t
Xbit_r6_c210 bl[210] br[210] wl[6] vdd gnd cell_6t
Xbit_r7_c210 bl[210] br[210] wl[7] vdd gnd cell_6t
Xbit_r8_c210 bl[210] br[210] wl[8] vdd gnd cell_6t
Xbit_r9_c210 bl[210] br[210] wl[9] vdd gnd cell_6t
Xbit_r10_c210 bl[210] br[210] wl[10] vdd gnd cell_6t
Xbit_r11_c210 bl[210] br[210] wl[11] vdd gnd cell_6t
Xbit_r12_c210 bl[210] br[210] wl[12] vdd gnd cell_6t
Xbit_r13_c210 bl[210] br[210] wl[13] vdd gnd cell_6t
Xbit_r14_c210 bl[210] br[210] wl[14] vdd gnd cell_6t
Xbit_r15_c210 bl[210] br[210] wl[15] vdd gnd cell_6t
Xbit_r16_c210 bl[210] br[210] wl[16] vdd gnd cell_6t
Xbit_r17_c210 bl[210] br[210] wl[17] vdd gnd cell_6t
Xbit_r18_c210 bl[210] br[210] wl[18] vdd gnd cell_6t
Xbit_r19_c210 bl[210] br[210] wl[19] vdd gnd cell_6t
Xbit_r20_c210 bl[210] br[210] wl[20] vdd gnd cell_6t
Xbit_r21_c210 bl[210] br[210] wl[21] vdd gnd cell_6t
Xbit_r22_c210 bl[210] br[210] wl[22] vdd gnd cell_6t
Xbit_r23_c210 bl[210] br[210] wl[23] vdd gnd cell_6t
Xbit_r24_c210 bl[210] br[210] wl[24] vdd gnd cell_6t
Xbit_r25_c210 bl[210] br[210] wl[25] vdd gnd cell_6t
Xbit_r26_c210 bl[210] br[210] wl[26] vdd gnd cell_6t
Xbit_r27_c210 bl[210] br[210] wl[27] vdd gnd cell_6t
Xbit_r28_c210 bl[210] br[210] wl[28] vdd gnd cell_6t
Xbit_r29_c210 bl[210] br[210] wl[29] vdd gnd cell_6t
Xbit_r30_c210 bl[210] br[210] wl[30] vdd gnd cell_6t
Xbit_r31_c210 bl[210] br[210] wl[31] vdd gnd cell_6t
Xbit_r32_c210 bl[210] br[210] wl[32] vdd gnd cell_6t
Xbit_r33_c210 bl[210] br[210] wl[33] vdd gnd cell_6t
Xbit_r34_c210 bl[210] br[210] wl[34] vdd gnd cell_6t
Xbit_r35_c210 bl[210] br[210] wl[35] vdd gnd cell_6t
Xbit_r36_c210 bl[210] br[210] wl[36] vdd gnd cell_6t
Xbit_r37_c210 bl[210] br[210] wl[37] vdd gnd cell_6t
Xbit_r38_c210 bl[210] br[210] wl[38] vdd gnd cell_6t
Xbit_r39_c210 bl[210] br[210] wl[39] vdd gnd cell_6t
Xbit_r40_c210 bl[210] br[210] wl[40] vdd gnd cell_6t
Xbit_r41_c210 bl[210] br[210] wl[41] vdd gnd cell_6t
Xbit_r42_c210 bl[210] br[210] wl[42] vdd gnd cell_6t
Xbit_r43_c210 bl[210] br[210] wl[43] vdd gnd cell_6t
Xbit_r44_c210 bl[210] br[210] wl[44] vdd gnd cell_6t
Xbit_r45_c210 bl[210] br[210] wl[45] vdd gnd cell_6t
Xbit_r46_c210 bl[210] br[210] wl[46] vdd gnd cell_6t
Xbit_r47_c210 bl[210] br[210] wl[47] vdd gnd cell_6t
Xbit_r48_c210 bl[210] br[210] wl[48] vdd gnd cell_6t
Xbit_r49_c210 bl[210] br[210] wl[49] vdd gnd cell_6t
Xbit_r50_c210 bl[210] br[210] wl[50] vdd gnd cell_6t
Xbit_r51_c210 bl[210] br[210] wl[51] vdd gnd cell_6t
Xbit_r52_c210 bl[210] br[210] wl[52] vdd gnd cell_6t
Xbit_r53_c210 bl[210] br[210] wl[53] vdd gnd cell_6t
Xbit_r54_c210 bl[210] br[210] wl[54] vdd gnd cell_6t
Xbit_r55_c210 bl[210] br[210] wl[55] vdd gnd cell_6t
Xbit_r56_c210 bl[210] br[210] wl[56] vdd gnd cell_6t
Xbit_r57_c210 bl[210] br[210] wl[57] vdd gnd cell_6t
Xbit_r58_c210 bl[210] br[210] wl[58] vdd gnd cell_6t
Xbit_r59_c210 bl[210] br[210] wl[59] vdd gnd cell_6t
Xbit_r60_c210 bl[210] br[210] wl[60] vdd gnd cell_6t
Xbit_r61_c210 bl[210] br[210] wl[61] vdd gnd cell_6t
Xbit_r62_c210 bl[210] br[210] wl[62] vdd gnd cell_6t
Xbit_r63_c210 bl[210] br[210] wl[63] vdd gnd cell_6t
Xbit_r64_c210 bl[210] br[210] wl[64] vdd gnd cell_6t
Xbit_r65_c210 bl[210] br[210] wl[65] vdd gnd cell_6t
Xbit_r66_c210 bl[210] br[210] wl[66] vdd gnd cell_6t
Xbit_r67_c210 bl[210] br[210] wl[67] vdd gnd cell_6t
Xbit_r68_c210 bl[210] br[210] wl[68] vdd gnd cell_6t
Xbit_r69_c210 bl[210] br[210] wl[69] vdd gnd cell_6t
Xbit_r70_c210 bl[210] br[210] wl[70] vdd gnd cell_6t
Xbit_r71_c210 bl[210] br[210] wl[71] vdd gnd cell_6t
Xbit_r72_c210 bl[210] br[210] wl[72] vdd gnd cell_6t
Xbit_r73_c210 bl[210] br[210] wl[73] vdd gnd cell_6t
Xbit_r74_c210 bl[210] br[210] wl[74] vdd gnd cell_6t
Xbit_r75_c210 bl[210] br[210] wl[75] vdd gnd cell_6t
Xbit_r76_c210 bl[210] br[210] wl[76] vdd gnd cell_6t
Xbit_r77_c210 bl[210] br[210] wl[77] vdd gnd cell_6t
Xbit_r78_c210 bl[210] br[210] wl[78] vdd gnd cell_6t
Xbit_r79_c210 bl[210] br[210] wl[79] vdd gnd cell_6t
Xbit_r80_c210 bl[210] br[210] wl[80] vdd gnd cell_6t
Xbit_r81_c210 bl[210] br[210] wl[81] vdd gnd cell_6t
Xbit_r82_c210 bl[210] br[210] wl[82] vdd gnd cell_6t
Xbit_r83_c210 bl[210] br[210] wl[83] vdd gnd cell_6t
Xbit_r84_c210 bl[210] br[210] wl[84] vdd gnd cell_6t
Xbit_r85_c210 bl[210] br[210] wl[85] vdd gnd cell_6t
Xbit_r86_c210 bl[210] br[210] wl[86] vdd gnd cell_6t
Xbit_r87_c210 bl[210] br[210] wl[87] vdd gnd cell_6t
Xbit_r88_c210 bl[210] br[210] wl[88] vdd gnd cell_6t
Xbit_r89_c210 bl[210] br[210] wl[89] vdd gnd cell_6t
Xbit_r90_c210 bl[210] br[210] wl[90] vdd gnd cell_6t
Xbit_r91_c210 bl[210] br[210] wl[91] vdd gnd cell_6t
Xbit_r92_c210 bl[210] br[210] wl[92] vdd gnd cell_6t
Xbit_r93_c210 bl[210] br[210] wl[93] vdd gnd cell_6t
Xbit_r94_c210 bl[210] br[210] wl[94] vdd gnd cell_6t
Xbit_r95_c210 bl[210] br[210] wl[95] vdd gnd cell_6t
Xbit_r96_c210 bl[210] br[210] wl[96] vdd gnd cell_6t
Xbit_r97_c210 bl[210] br[210] wl[97] vdd gnd cell_6t
Xbit_r98_c210 bl[210] br[210] wl[98] vdd gnd cell_6t
Xbit_r99_c210 bl[210] br[210] wl[99] vdd gnd cell_6t
Xbit_r100_c210 bl[210] br[210] wl[100] vdd gnd cell_6t
Xbit_r101_c210 bl[210] br[210] wl[101] vdd gnd cell_6t
Xbit_r102_c210 bl[210] br[210] wl[102] vdd gnd cell_6t
Xbit_r103_c210 bl[210] br[210] wl[103] vdd gnd cell_6t
Xbit_r104_c210 bl[210] br[210] wl[104] vdd gnd cell_6t
Xbit_r105_c210 bl[210] br[210] wl[105] vdd gnd cell_6t
Xbit_r106_c210 bl[210] br[210] wl[106] vdd gnd cell_6t
Xbit_r107_c210 bl[210] br[210] wl[107] vdd gnd cell_6t
Xbit_r108_c210 bl[210] br[210] wl[108] vdd gnd cell_6t
Xbit_r109_c210 bl[210] br[210] wl[109] vdd gnd cell_6t
Xbit_r110_c210 bl[210] br[210] wl[110] vdd gnd cell_6t
Xbit_r111_c210 bl[210] br[210] wl[111] vdd gnd cell_6t
Xbit_r112_c210 bl[210] br[210] wl[112] vdd gnd cell_6t
Xbit_r113_c210 bl[210] br[210] wl[113] vdd gnd cell_6t
Xbit_r114_c210 bl[210] br[210] wl[114] vdd gnd cell_6t
Xbit_r115_c210 bl[210] br[210] wl[115] vdd gnd cell_6t
Xbit_r116_c210 bl[210] br[210] wl[116] vdd gnd cell_6t
Xbit_r117_c210 bl[210] br[210] wl[117] vdd gnd cell_6t
Xbit_r118_c210 bl[210] br[210] wl[118] vdd gnd cell_6t
Xbit_r119_c210 bl[210] br[210] wl[119] vdd gnd cell_6t
Xbit_r120_c210 bl[210] br[210] wl[120] vdd gnd cell_6t
Xbit_r121_c210 bl[210] br[210] wl[121] vdd gnd cell_6t
Xbit_r122_c210 bl[210] br[210] wl[122] vdd gnd cell_6t
Xbit_r123_c210 bl[210] br[210] wl[123] vdd gnd cell_6t
Xbit_r124_c210 bl[210] br[210] wl[124] vdd gnd cell_6t
Xbit_r125_c210 bl[210] br[210] wl[125] vdd gnd cell_6t
Xbit_r126_c210 bl[210] br[210] wl[126] vdd gnd cell_6t
Xbit_r127_c210 bl[210] br[210] wl[127] vdd gnd cell_6t
Xbit_r0_c211 bl[211] br[211] wl[0] vdd gnd cell_6t
Xbit_r1_c211 bl[211] br[211] wl[1] vdd gnd cell_6t
Xbit_r2_c211 bl[211] br[211] wl[2] vdd gnd cell_6t
Xbit_r3_c211 bl[211] br[211] wl[3] vdd gnd cell_6t
Xbit_r4_c211 bl[211] br[211] wl[4] vdd gnd cell_6t
Xbit_r5_c211 bl[211] br[211] wl[5] vdd gnd cell_6t
Xbit_r6_c211 bl[211] br[211] wl[6] vdd gnd cell_6t
Xbit_r7_c211 bl[211] br[211] wl[7] vdd gnd cell_6t
Xbit_r8_c211 bl[211] br[211] wl[8] vdd gnd cell_6t
Xbit_r9_c211 bl[211] br[211] wl[9] vdd gnd cell_6t
Xbit_r10_c211 bl[211] br[211] wl[10] vdd gnd cell_6t
Xbit_r11_c211 bl[211] br[211] wl[11] vdd gnd cell_6t
Xbit_r12_c211 bl[211] br[211] wl[12] vdd gnd cell_6t
Xbit_r13_c211 bl[211] br[211] wl[13] vdd gnd cell_6t
Xbit_r14_c211 bl[211] br[211] wl[14] vdd gnd cell_6t
Xbit_r15_c211 bl[211] br[211] wl[15] vdd gnd cell_6t
Xbit_r16_c211 bl[211] br[211] wl[16] vdd gnd cell_6t
Xbit_r17_c211 bl[211] br[211] wl[17] vdd gnd cell_6t
Xbit_r18_c211 bl[211] br[211] wl[18] vdd gnd cell_6t
Xbit_r19_c211 bl[211] br[211] wl[19] vdd gnd cell_6t
Xbit_r20_c211 bl[211] br[211] wl[20] vdd gnd cell_6t
Xbit_r21_c211 bl[211] br[211] wl[21] vdd gnd cell_6t
Xbit_r22_c211 bl[211] br[211] wl[22] vdd gnd cell_6t
Xbit_r23_c211 bl[211] br[211] wl[23] vdd gnd cell_6t
Xbit_r24_c211 bl[211] br[211] wl[24] vdd gnd cell_6t
Xbit_r25_c211 bl[211] br[211] wl[25] vdd gnd cell_6t
Xbit_r26_c211 bl[211] br[211] wl[26] vdd gnd cell_6t
Xbit_r27_c211 bl[211] br[211] wl[27] vdd gnd cell_6t
Xbit_r28_c211 bl[211] br[211] wl[28] vdd gnd cell_6t
Xbit_r29_c211 bl[211] br[211] wl[29] vdd gnd cell_6t
Xbit_r30_c211 bl[211] br[211] wl[30] vdd gnd cell_6t
Xbit_r31_c211 bl[211] br[211] wl[31] vdd gnd cell_6t
Xbit_r32_c211 bl[211] br[211] wl[32] vdd gnd cell_6t
Xbit_r33_c211 bl[211] br[211] wl[33] vdd gnd cell_6t
Xbit_r34_c211 bl[211] br[211] wl[34] vdd gnd cell_6t
Xbit_r35_c211 bl[211] br[211] wl[35] vdd gnd cell_6t
Xbit_r36_c211 bl[211] br[211] wl[36] vdd gnd cell_6t
Xbit_r37_c211 bl[211] br[211] wl[37] vdd gnd cell_6t
Xbit_r38_c211 bl[211] br[211] wl[38] vdd gnd cell_6t
Xbit_r39_c211 bl[211] br[211] wl[39] vdd gnd cell_6t
Xbit_r40_c211 bl[211] br[211] wl[40] vdd gnd cell_6t
Xbit_r41_c211 bl[211] br[211] wl[41] vdd gnd cell_6t
Xbit_r42_c211 bl[211] br[211] wl[42] vdd gnd cell_6t
Xbit_r43_c211 bl[211] br[211] wl[43] vdd gnd cell_6t
Xbit_r44_c211 bl[211] br[211] wl[44] vdd gnd cell_6t
Xbit_r45_c211 bl[211] br[211] wl[45] vdd gnd cell_6t
Xbit_r46_c211 bl[211] br[211] wl[46] vdd gnd cell_6t
Xbit_r47_c211 bl[211] br[211] wl[47] vdd gnd cell_6t
Xbit_r48_c211 bl[211] br[211] wl[48] vdd gnd cell_6t
Xbit_r49_c211 bl[211] br[211] wl[49] vdd gnd cell_6t
Xbit_r50_c211 bl[211] br[211] wl[50] vdd gnd cell_6t
Xbit_r51_c211 bl[211] br[211] wl[51] vdd gnd cell_6t
Xbit_r52_c211 bl[211] br[211] wl[52] vdd gnd cell_6t
Xbit_r53_c211 bl[211] br[211] wl[53] vdd gnd cell_6t
Xbit_r54_c211 bl[211] br[211] wl[54] vdd gnd cell_6t
Xbit_r55_c211 bl[211] br[211] wl[55] vdd gnd cell_6t
Xbit_r56_c211 bl[211] br[211] wl[56] vdd gnd cell_6t
Xbit_r57_c211 bl[211] br[211] wl[57] vdd gnd cell_6t
Xbit_r58_c211 bl[211] br[211] wl[58] vdd gnd cell_6t
Xbit_r59_c211 bl[211] br[211] wl[59] vdd gnd cell_6t
Xbit_r60_c211 bl[211] br[211] wl[60] vdd gnd cell_6t
Xbit_r61_c211 bl[211] br[211] wl[61] vdd gnd cell_6t
Xbit_r62_c211 bl[211] br[211] wl[62] vdd gnd cell_6t
Xbit_r63_c211 bl[211] br[211] wl[63] vdd gnd cell_6t
Xbit_r64_c211 bl[211] br[211] wl[64] vdd gnd cell_6t
Xbit_r65_c211 bl[211] br[211] wl[65] vdd gnd cell_6t
Xbit_r66_c211 bl[211] br[211] wl[66] vdd gnd cell_6t
Xbit_r67_c211 bl[211] br[211] wl[67] vdd gnd cell_6t
Xbit_r68_c211 bl[211] br[211] wl[68] vdd gnd cell_6t
Xbit_r69_c211 bl[211] br[211] wl[69] vdd gnd cell_6t
Xbit_r70_c211 bl[211] br[211] wl[70] vdd gnd cell_6t
Xbit_r71_c211 bl[211] br[211] wl[71] vdd gnd cell_6t
Xbit_r72_c211 bl[211] br[211] wl[72] vdd gnd cell_6t
Xbit_r73_c211 bl[211] br[211] wl[73] vdd gnd cell_6t
Xbit_r74_c211 bl[211] br[211] wl[74] vdd gnd cell_6t
Xbit_r75_c211 bl[211] br[211] wl[75] vdd gnd cell_6t
Xbit_r76_c211 bl[211] br[211] wl[76] vdd gnd cell_6t
Xbit_r77_c211 bl[211] br[211] wl[77] vdd gnd cell_6t
Xbit_r78_c211 bl[211] br[211] wl[78] vdd gnd cell_6t
Xbit_r79_c211 bl[211] br[211] wl[79] vdd gnd cell_6t
Xbit_r80_c211 bl[211] br[211] wl[80] vdd gnd cell_6t
Xbit_r81_c211 bl[211] br[211] wl[81] vdd gnd cell_6t
Xbit_r82_c211 bl[211] br[211] wl[82] vdd gnd cell_6t
Xbit_r83_c211 bl[211] br[211] wl[83] vdd gnd cell_6t
Xbit_r84_c211 bl[211] br[211] wl[84] vdd gnd cell_6t
Xbit_r85_c211 bl[211] br[211] wl[85] vdd gnd cell_6t
Xbit_r86_c211 bl[211] br[211] wl[86] vdd gnd cell_6t
Xbit_r87_c211 bl[211] br[211] wl[87] vdd gnd cell_6t
Xbit_r88_c211 bl[211] br[211] wl[88] vdd gnd cell_6t
Xbit_r89_c211 bl[211] br[211] wl[89] vdd gnd cell_6t
Xbit_r90_c211 bl[211] br[211] wl[90] vdd gnd cell_6t
Xbit_r91_c211 bl[211] br[211] wl[91] vdd gnd cell_6t
Xbit_r92_c211 bl[211] br[211] wl[92] vdd gnd cell_6t
Xbit_r93_c211 bl[211] br[211] wl[93] vdd gnd cell_6t
Xbit_r94_c211 bl[211] br[211] wl[94] vdd gnd cell_6t
Xbit_r95_c211 bl[211] br[211] wl[95] vdd gnd cell_6t
Xbit_r96_c211 bl[211] br[211] wl[96] vdd gnd cell_6t
Xbit_r97_c211 bl[211] br[211] wl[97] vdd gnd cell_6t
Xbit_r98_c211 bl[211] br[211] wl[98] vdd gnd cell_6t
Xbit_r99_c211 bl[211] br[211] wl[99] vdd gnd cell_6t
Xbit_r100_c211 bl[211] br[211] wl[100] vdd gnd cell_6t
Xbit_r101_c211 bl[211] br[211] wl[101] vdd gnd cell_6t
Xbit_r102_c211 bl[211] br[211] wl[102] vdd gnd cell_6t
Xbit_r103_c211 bl[211] br[211] wl[103] vdd gnd cell_6t
Xbit_r104_c211 bl[211] br[211] wl[104] vdd gnd cell_6t
Xbit_r105_c211 bl[211] br[211] wl[105] vdd gnd cell_6t
Xbit_r106_c211 bl[211] br[211] wl[106] vdd gnd cell_6t
Xbit_r107_c211 bl[211] br[211] wl[107] vdd gnd cell_6t
Xbit_r108_c211 bl[211] br[211] wl[108] vdd gnd cell_6t
Xbit_r109_c211 bl[211] br[211] wl[109] vdd gnd cell_6t
Xbit_r110_c211 bl[211] br[211] wl[110] vdd gnd cell_6t
Xbit_r111_c211 bl[211] br[211] wl[111] vdd gnd cell_6t
Xbit_r112_c211 bl[211] br[211] wl[112] vdd gnd cell_6t
Xbit_r113_c211 bl[211] br[211] wl[113] vdd gnd cell_6t
Xbit_r114_c211 bl[211] br[211] wl[114] vdd gnd cell_6t
Xbit_r115_c211 bl[211] br[211] wl[115] vdd gnd cell_6t
Xbit_r116_c211 bl[211] br[211] wl[116] vdd gnd cell_6t
Xbit_r117_c211 bl[211] br[211] wl[117] vdd gnd cell_6t
Xbit_r118_c211 bl[211] br[211] wl[118] vdd gnd cell_6t
Xbit_r119_c211 bl[211] br[211] wl[119] vdd gnd cell_6t
Xbit_r120_c211 bl[211] br[211] wl[120] vdd gnd cell_6t
Xbit_r121_c211 bl[211] br[211] wl[121] vdd gnd cell_6t
Xbit_r122_c211 bl[211] br[211] wl[122] vdd gnd cell_6t
Xbit_r123_c211 bl[211] br[211] wl[123] vdd gnd cell_6t
Xbit_r124_c211 bl[211] br[211] wl[124] vdd gnd cell_6t
Xbit_r125_c211 bl[211] br[211] wl[125] vdd gnd cell_6t
Xbit_r126_c211 bl[211] br[211] wl[126] vdd gnd cell_6t
Xbit_r127_c211 bl[211] br[211] wl[127] vdd gnd cell_6t
Xbit_r0_c212 bl[212] br[212] wl[0] vdd gnd cell_6t
Xbit_r1_c212 bl[212] br[212] wl[1] vdd gnd cell_6t
Xbit_r2_c212 bl[212] br[212] wl[2] vdd gnd cell_6t
Xbit_r3_c212 bl[212] br[212] wl[3] vdd gnd cell_6t
Xbit_r4_c212 bl[212] br[212] wl[4] vdd gnd cell_6t
Xbit_r5_c212 bl[212] br[212] wl[5] vdd gnd cell_6t
Xbit_r6_c212 bl[212] br[212] wl[6] vdd gnd cell_6t
Xbit_r7_c212 bl[212] br[212] wl[7] vdd gnd cell_6t
Xbit_r8_c212 bl[212] br[212] wl[8] vdd gnd cell_6t
Xbit_r9_c212 bl[212] br[212] wl[9] vdd gnd cell_6t
Xbit_r10_c212 bl[212] br[212] wl[10] vdd gnd cell_6t
Xbit_r11_c212 bl[212] br[212] wl[11] vdd gnd cell_6t
Xbit_r12_c212 bl[212] br[212] wl[12] vdd gnd cell_6t
Xbit_r13_c212 bl[212] br[212] wl[13] vdd gnd cell_6t
Xbit_r14_c212 bl[212] br[212] wl[14] vdd gnd cell_6t
Xbit_r15_c212 bl[212] br[212] wl[15] vdd gnd cell_6t
Xbit_r16_c212 bl[212] br[212] wl[16] vdd gnd cell_6t
Xbit_r17_c212 bl[212] br[212] wl[17] vdd gnd cell_6t
Xbit_r18_c212 bl[212] br[212] wl[18] vdd gnd cell_6t
Xbit_r19_c212 bl[212] br[212] wl[19] vdd gnd cell_6t
Xbit_r20_c212 bl[212] br[212] wl[20] vdd gnd cell_6t
Xbit_r21_c212 bl[212] br[212] wl[21] vdd gnd cell_6t
Xbit_r22_c212 bl[212] br[212] wl[22] vdd gnd cell_6t
Xbit_r23_c212 bl[212] br[212] wl[23] vdd gnd cell_6t
Xbit_r24_c212 bl[212] br[212] wl[24] vdd gnd cell_6t
Xbit_r25_c212 bl[212] br[212] wl[25] vdd gnd cell_6t
Xbit_r26_c212 bl[212] br[212] wl[26] vdd gnd cell_6t
Xbit_r27_c212 bl[212] br[212] wl[27] vdd gnd cell_6t
Xbit_r28_c212 bl[212] br[212] wl[28] vdd gnd cell_6t
Xbit_r29_c212 bl[212] br[212] wl[29] vdd gnd cell_6t
Xbit_r30_c212 bl[212] br[212] wl[30] vdd gnd cell_6t
Xbit_r31_c212 bl[212] br[212] wl[31] vdd gnd cell_6t
Xbit_r32_c212 bl[212] br[212] wl[32] vdd gnd cell_6t
Xbit_r33_c212 bl[212] br[212] wl[33] vdd gnd cell_6t
Xbit_r34_c212 bl[212] br[212] wl[34] vdd gnd cell_6t
Xbit_r35_c212 bl[212] br[212] wl[35] vdd gnd cell_6t
Xbit_r36_c212 bl[212] br[212] wl[36] vdd gnd cell_6t
Xbit_r37_c212 bl[212] br[212] wl[37] vdd gnd cell_6t
Xbit_r38_c212 bl[212] br[212] wl[38] vdd gnd cell_6t
Xbit_r39_c212 bl[212] br[212] wl[39] vdd gnd cell_6t
Xbit_r40_c212 bl[212] br[212] wl[40] vdd gnd cell_6t
Xbit_r41_c212 bl[212] br[212] wl[41] vdd gnd cell_6t
Xbit_r42_c212 bl[212] br[212] wl[42] vdd gnd cell_6t
Xbit_r43_c212 bl[212] br[212] wl[43] vdd gnd cell_6t
Xbit_r44_c212 bl[212] br[212] wl[44] vdd gnd cell_6t
Xbit_r45_c212 bl[212] br[212] wl[45] vdd gnd cell_6t
Xbit_r46_c212 bl[212] br[212] wl[46] vdd gnd cell_6t
Xbit_r47_c212 bl[212] br[212] wl[47] vdd gnd cell_6t
Xbit_r48_c212 bl[212] br[212] wl[48] vdd gnd cell_6t
Xbit_r49_c212 bl[212] br[212] wl[49] vdd gnd cell_6t
Xbit_r50_c212 bl[212] br[212] wl[50] vdd gnd cell_6t
Xbit_r51_c212 bl[212] br[212] wl[51] vdd gnd cell_6t
Xbit_r52_c212 bl[212] br[212] wl[52] vdd gnd cell_6t
Xbit_r53_c212 bl[212] br[212] wl[53] vdd gnd cell_6t
Xbit_r54_c212 bl[212] br[212] wl[54] vdd gnd cell_6t
Xbit_r55_c212 bl[212] br[212] wl[55] vdd gnd cell_6t
Xbit_r56_c212 bl[212] br[212] wl[56] vdd gnd cell_6t
Xbit_r57_c212 bl[212] br[212] wl[57] vdd gnd cell_6t
Xbit_r58_c212 bl[212] br[212] wl[58] vdd gnd cell_6t
Xbit_r59_c212 bl[212] br[212] wl[59] vdd gnd cell_6t
Xbit_r60_c212 bl[212] br[212] wl[60] vdd gnd cell_6t
Xbit_r61_c212 bl[212] br[212] wl[61] vdd gnd cell_6t
Xbit_r62_c212 bl[212] br[212] wl[62] vdd gnd cell_6t
Xbit_r63_c212 bl[212] br[212] wl[63] vdd gnd cell_6t
Xbit_r64_c212 bl[212] br[212] wl[64] vdd gnd cell_6t
Xbit_r65_c212 bl[212] br[212] wl[65] vdd gnd cell_6t
Xbit_r66_c212 bl[212] br[212] wl[66] vdd gnd cell_6t
Xbit_r67_c212 bl[212] br[212] wl[67] vdd gnd cell_6t
Xbit_r68_c212 bl[212] br[212] wl[68] vdd gnd cell_6t
Xbit_r69_c212 bl[212] br[212] wl[69] vdd gnd cell_6t
Xbit_r70_c212 bl[212] br[212] wl[70] vdd gnd cell_6t
Xbit_r71_c212 bl[212] br[212] wl[71] vdd gnd cell_6t
Xbit_r72_c212 bl[212] br[212] wl[72] vdd gnd cell_6t
Xbit_r73_c212 bl[212] br[212] wl[73] vdd gnd cell_6t
Xbit_r74_c212 bl[212] br[212] wl[74] vdd gnd cell_6t
Xbit_r75_c212 bl[212] br[212] wl[75] vdd gnd cell_6t
Xbit_r76_c212 bl[212] br[212] wl[76] vdd gnd cell_6t
Xbit_r77_c212 bl[212] br[212] wl[77] vdd gnd cell_6t
Xbit_r78_c212 bl[212] br[212] wl[78] vdd gnd cell_6t
Xbit_r79_c212 bl[212] br[212] wl[79] vdd gnd cell_6t
Xbit_r80_c212 bl[212] br[212] wl[80] vdd gnd cell_6t
Xbit_r81_c212 bl[212] br[212] wl[81] vdd gnd cell_6t
Xbit_r82_c212 bl[212] br[212] wl[82] vdd gnd cell_6t
Xbit_r83_c212 bl[212] br[212] wl[83] vdd gnd cell_6t
Xbit_r84_c212 bl[212] br[212] wl[84] vdd gnd cell_6t
Xbit_r85_c212 bl[212] br[212] wl[85] vdd gnd cell_6t
Xbit_r86_c212 bl[212] br[212] wl[86] vdd gnd cell_6t
Xbit_r87_c212 bl[212] br[212] wl[87] vdd gnd cell_6t
Xbit_r88_c212 bl[212] br[212] wl[88] vdd gnd cell_6t
Xbit_r89_c212 bl[212] br[212] wl[89] vdd gnd cell_6t
Xbit_r90_c212 bl[212] br[212] wl[90] vdd gnd cell_6t
Xbit_r91_c212 bl[212] br[212] wl[91] vdd gnd cell_6t
Xbit_r92_c212 bl[212] br[212] wl[92] vdd gnd cell_6t
Xbit_r93_c212 bl[212] br[212] wl[93] vdd gnd cell_6t
Xbit_r94_c212 bl[212] br[212] wl[94] vdd gnd cell_6t
Xbit_r95_c212 bl[212] br[212] wl[95] vdd gnd cell_6t
Xbit_r96_c212 bl[212] br[212] wl[96] vdd gnd cell_6t
Xbit_r97_c212 bl[212] br[212] wl[97] vdd gnd cell_6t
Xbit_r98_c212 bl[212] br[212] wl[98] vdd gnd cell_6t
Xbit_r99_c212 bl[212] br[212] wl[99] vdd gnd cell_6t
Xbit_r100_c212 bl[212] br[212] wl[100] vdd gnd cell_6t
Xbit_r101_c212 bl[212] br[212] wl[101] vdd gnd cell_6t
Xbit_r102_c212 bl[212] br[212] wl[102] vdd gnd cell_6t
Xbit_r103_c212 bl[212] br[212] wl[103] vdd gnd cell_6t
Xbit_r104_c212 bl[212] br[212] wl[104] vdd gnd cell_6t
Xbit_r105_c212 bl[212] br[212] wl[105] vdd gnd cell_6t
Xbit_r106_c212 bl[212] br[212] wl[106] vdd gnd cell_6t
Xbit_r107_c212 bl[212] br[212] wl[107] vdd gnd cell_6t
Xbit_r108_c212 bl[212] br[212] wl[108] vdd gnd cell_6t
Xbit_r109_c212 bl[212] br[212] wl[109] vdd gnd cell_6t
Xbit_r110_c212 bl[212] br[212] wl[110] vdd gnd cell_6t
Xbit_r111_c212 bl[212] br[212] wl[111] vdd gnd cell_6t
Xbit_r112_c212 bl[212] br[212] wl[112] vdd gnd cell_6t
Xbit_r113_c212 bl[212] br[212] wl[113] vdd gnd cell_6t
Xbit_r114_c212 bl[212] br[212] wl[114] vdd gnd cell_6t
Xbit_r115_c212 bl[212] br[212] wl[115] vdd gnd cell_6t
Xbit_r116_c212 bl[212] br[212] wl[116] vdd gnd cell_6t
Xbit_r117_c212 bl[212] br[212] wl[117] vdd gnd cell_6t
Xbit_r118_c212 bl[212] br[212] wl[118] vdd gnd cell_6t
Xbit_r119_c212 bl[212] br[212] wl[119] vdd gnd cell_6t
Xbit_r120_c212 bl[212] br[212] wl[120] vdd gnd cell_6t
Xbit_r121_c212 bl[212] br[212] wl[121] vdd gnd cell_6t
Xbit_r122_c212 bl[212] br[212] wl[122] vdd gnd cell_6t
Xbit_r123_c212 bl[212] br[212] wl[123] vdd gnd cell_6t
Xbit_r124_c212 bl[212] br[212] wl[124] vdd gnd cell_6t
Xbit_r125_c212 bl[212] br[212] wl[125] vdd gnd cell_6t
Xbit_r126_c212 bl[212] br[212] wl[126] vdd gnd cell_6t
Xbit_r127_c212 bl[212] br[212] wl[127] vdd gnd cell_6t
Xbit_r0_c213 bl[213] br[213] wl[0] vdd gnd cell_6t
Xbit_r1_c213 bl[213] br[213] wl[1] vdd gnd cell_6t
Xbit_r2_c213 bl[213] br[213] wl[2] vdd gnd cell_6t
Xbit_r3_c213 bl[213] br[213] wl[3] vdd gnd cell_6t
Xbit_r4_c213 bl[213] br[213] wl[4] vdd gnd cell_6t
Xbit_r5_c213 bl[213] br[213] wl[5] vdd gnd cell_6t
Xbit_r6_c213 bl[213] br[213] wl[6] vdd gnd cell_6t
Xbit_r7_c213 bl[213] br[213] wl[7] vdd gnd cell_6t
Xbit_r8_c213 bl[213] br[213] wl[8] vdd gnd cell_6t
Xbit_r9_c213 bl[213] br[213] wl[9] vdd gnd cell_6t
Xbit_r10_c213 bl[213] br[213] wl[10] vdd gnd cell_6t
Xbit_r11_c213 bl[213] br[213] wl[11] vdd gnd cell_6t
Xbit_r12_c213 bl[213] br[213] wl[12] vdd gnd cell_6t
Xbit_r13_c213 bl[213] br[213] wl[13] vdd gnd cell_6t
Xbit_r14_c213 bl[213] br[213] wl[14] vdd gnd cell_6t
Xbit_r15_c213 bl[213] br[213] wl[15] vdd gnd cell_6t
Xbit_r16_c213 bl[213] br[213] wl[16] vdd gnd cell_6t
Xbit_r17_c213 bl[213] br[213] wl[17] vdd gnd cell_6t
Xbit_r18_c213 bl[213] br[213] wl[18] vdd gnd cell_6t
Xbit_r19_c213 bl[213] br[213] wl[19] vdd gnd cell_6t
Xbit_r20_c213 bl[213] br[213] wl[20] vdd gnd cell_6t
Xbit_r21_c213 bl[213] br[213] wl[21] vdd gnd cell_6t
Xbit_r22_c213 bl[213] br[213] wl[22] vdd gnd cell_6t
Xbit_r23_c213 bl[213] br[213] wl[23] vdd gnd cell_6t
Xbit_r24_c213 bl[213] br[213] wl[24] vdd gnd cell_6t
Xbit_r25_c213 bl[213] br[213] wl[25] vdd gnd cell_6t
Xbit_r26_c213 bl[213] br[213] wl[26] vdd gnd cell_6t
Xbit_r27_c213 bl[213] br[213] wl[27] vdd gnd cell_6t
Xbit_r28_c213 bl[213] br[213] wl[28] vdd gnd cell_6t
Xbit_r29_c213 bl[213] br[213] wl[29] vdd gnd cell_6t
Xbit_r30_c213 bl[213] br[213] wl[30] vdd gnd cell_6t
Xbit_r31_c213 bl[213] br[213] wl[31] vdd gnd cell_6t
Xbit_r32_c213 bl[213] br[213] wl[32] vdd gnd cell_6t
Xbit_r33_c213 bl[213] br[213] wl[33] vdd gnd cell_6t
Xbit_r34_c213 bl[213] br[213] wl[34] vdd gnd cell_6t
Xbit_r35_c213 bl[213] br[213] wl[35] vdd gnd cell_6t
Xbit_r36_c213 bl[213] br[213] wl[36] vdd gnd cell_6t
Xbit_r37_c213 bl[213] br[213] wl[37] vdd gnd cell_6t
Xbit_r38_c213 bl[213] br[213] wl[38] vdd gnd cell_6t
Xbit_r39_c213 bl[213] br[213] wl[39] vdd gnd cell_6t
Xbit_r40_c213 bl[213] br[213] wl[40] vdd gnd cell_6t
Xbit_r41_c213 bl[213] br[213] wl[41] vdd gnd cell_6t
Xbit_r42_c213 bl[213] br[213] wl[42] vdd gnd cell_6t
Xbit_r43_c213 bl[213] br[213] wl[43] vdd gnd cell_6t
Xbit_r44_c213 bl[213] br[213] wl[44] vdd gnd cell_6t
Xbit_r45_c213 bl[213] br[213] wl[45] vdd gnd cell_6t
Xbit_r46_c213 bl[213] br[213] wl[46] vdd gnd cell_6t
Xbit_r47_c213 bl[213] br[213] wl[47] vdd gnd cell_6t
Xbit_r48_c213 bl[213] br[213] wl[48] vdd gnd cell_6t
Xbit_r49_c213 bl[213] br[213] wl[49] vdd gnd cell_6t
Xbit_r50_c213 bl[213] br[213] wl[50] vdd gnd cell_6t
Xbit_r51_c213 bl[213] br[213] wl[51] vdd gnd cell_6t
Xbit_r52_c213 bl[213] br[213] wl[52] vdd gnd cell_6t
Xbit_r53_c213 bl[213] br[213] wl[53] vdd gnd cell_6t
Xbit_r54_c213 bl[213] br[213] wl[54] vdd gnd cell_6t
Xbit_r55_c213 bl[213] br[213] wl[55] vdd gnd cell_6t
Xbit_r56_c213 bl[213] br[213] wl[56] vdd gnd cell_6t
Xbit_r57_c213 bl[213] br[213] wl[57] vdd gnd cell_6t
Xbit_r58_c213 bl[213] br[213] wl[58] vdd gnd cell_6t
Xbit_r59_c213 bl[213] br[213] wl[59] vdd gnd cell_6t
Xbit_r60_c213 bl[213] br[213] wl[60] vdd gnd cell_6t
Xbit_r61_c213 bl[213] br[213] wl[61] vdd gnd cell_6t
Xbit_r62_c213 bl[213] br[213] wl[62] vdd gnd cell_6t
Xbit_r63_c213 bl[213] br[213] wl[63] vdd gnd cell_6t
Xbit_r64_c213 bl[213] br[213] wl[64] vdd gnd cell_6t
Xbit_r65_c213 bl[213] br[213] wl[65] vdd gnd cell_6t
Xbit_r66_c213 bl[213] br[213] wl[66] vdd gnd cell_6t
Xbit_r67_c213 bl[213] br[213] wl[67] vdd gnd cell_6t
Xbit_r68_c213 bl[213] br[213] wl[68] vdd gnd cell_6t
Xbit_r69_c213 bl[213] br[213] wl[69] vdd gnd cell_6t
Xbit_r70_c213 bl[213] br[213] wl[70] vdd gnd cell_6t
Xbit_r71_c213 bl[213] br[213] wl[71] vdd gnd cell_6t
Xbit_r72_c213 bl[213] br[213] wl[72] vdd gnd cell_6t
Xbit_r73_c213 bl[213] br[213] wl[73] vdd gnd cell_6t
Xbit_r74_c213 bl[213] br[213] wl[74] vdd gnd cell_6t
Xbit_r75_c213 bl[213] br[213] wl[75] vdd gnd cell_6t
Xbit_r76_c213 bl[213] br[213] wl[76] vdd gnd cell_6t
Xbit_r77_c213 bl[213] br[213] wl[77] vdd gnd cell_6t
Xbit_r78_c213 bl[213] br[213] wl[78] vdd gnd cell_6t
Xbit_r79_c213 bl[213] br[213] wl[79] vdd gnd cell_6t
Xbit_r80_c213 bl[213] br[213] wl[80] vdd gnd cell_6t
Xbit_r81_c213 bl[213] br[213] wl[81] vdd gnd cell_6t
Xbit_r82_c213 bl[213] br[213] wl[82] vdd gnd cell_6t
Xbit_r83_c213 bl[213] br[213] wl[83] vdd gnd cell_6t
Xbit_r84_c213 bl[213] br[213] wl[84] vdd gnd cell_6t
Xbit_r85_c213 bl[213] br[213] wl[85] vdd gnd cell_6t
Xbit_r86_c213 bl[213] br[213] wl[86] vdd gnd cell_6t
Xbit_r87_c213 bl[213] br[213] wl[87] vdd gnd cell_6t
Xbit_r88_c213 bl[213] br[213] wl[88] vdd gnd cell_6t
Xbit_r89_c213 bl[213] br[213] wl[89] vdd gnd cell_6t
Xbit_r90_c213 bl[213] br[213] wl[90] vdd gnd cell_6t
Xbit_r91_c213 bl[213] br[213] wl[91] vdd gnd cell_6t
Xbit_r92_c213 bl[213] br[213] wl[92] vdd gnd cell_6t
Xbit_r93_c213 bl[213] br[213] wl[93] vdd gnd cell_6t
Xbit_r94_c213 bl[213] br[213] wl[94] vdd gnd cell_6t
Xbit_r95_c213 bl[213] br[213] wl[95] vdd gnd cell_6t
Xbit_r96_c213 bl[213] br[213] wl[96] vdd gnd cell_6t
Xbit_r97_c213 bl[213] br[213] wl[97] vdd gnd cell_6t
Xbit_r98_c213 bl[213] br[213] wl[98] vdd gnd cell_6t
Xbit_r99_c213 bl[213] br[213] wl[99] vdd gnd cell_6t
Xbit_r100_c213 bl[213] br[213] wl[100] vdd gnd cell_6t
Xbit_r101_c213 bl[213] br[213] wl[101] vdd gnd cell_6t
Xbit_r102_c213 bl[213] br[213] wl[102] vdd gnd cell_6t
Xbit_r103_c213 bl[213] br[213] wl[103] vdd gnd cell_6t
Xbit_r104_c213 bl[213] br[213] wl[104] vdd gnd cell_6t
Xbit_r105_c213 bl[213] br[213] wl[105] vdd gnd cell_6t
Xbit_r106_c213 bl[213] br[213] wl[106] vdd gnd cell_6t
Xbit_r107_c213 bl[213] br[213] wl[107] vdd gnd cell_6t
Xbit_r108_c213 bl[213] br[213] wl[108] vdd gnd cell_6t
Xbit_r109_c213 bl[213] br[213] wl[109] vdd gnd cell_6t
Xbit_r110_c213 bl[213] br[213] wl[110] vdd gnd cell_6t
Xbit_r111_c213 bl[213] br[213] wl[111] vdd gnd cell_6t
Xbit_r112_c213 bl[213] br[213] wl[112] vdd gnd cell_6t
Xbit_r113_c213 bl[213] br[213] wl[113] vdd gnd cell_6t
Xbit_r114_c213 bl[213] br[213] wl[114] vdd gnd cell_6t
Xbit_r115_c213 bl[213] br[213] wl[115] vdd gnd cell_6t
Xbit_r116_c213 bl[213] br[213] wl[116] vdd gnd cell_6t
Xbit_r117_c213 bl[213] br[213] wl[117] vdd gnd cell_6t
Xbit_r118_c213 bl[213] br[213] wl[118] vdd gnd cell_6t
Xbit_r119_c213 bl[213] br[213] wl[119] vdd gnd cell_6t
Xbit_r120_c213 bl[213] br[213] wl[120] vdd gnd cell_6t
Xbit_r121_c213 bl[213] br[213] wl[121] vdd gnd cell_6t
Xbit_r122_c213 bl[213] br[213] wl[122] vdd gnd cell_6t
Xbit_r123_c213 bl[213] br[213] wl[123] vdd gnd cell_6t
Xbit_r124_c213 bl[213] br[213] wl[124] vdd gnd cell_6t
Xbit_r125_c213 bl[213] br[213] wl[125] vdd gnd cell_6t
Xbit_r126_c213 bl[213] br[213] wl[126] vdd gnd cell_6t
Xbit_r127_c213 bl[213] br[213] wl[127] vdd gnd cell_6t
Xbit_r0_c214 bl[214] br[214] wl[0] vdd gnd cell_6t
Xbit_r1_c214 bl[214] br[214] wl[1] vdd gnd cell_6t
Xbit_r2_c214 bl[214] br[214] wl[2] vdd gnd cell_6t
Xbit_r3_c214 bl[214] br[214] wl[3] vdd gnd cell_6t
Xbit_r4_c214 bl[214] br[214] wl[4] vdd gnd cell_6t
Xbit_r5_c214 bl[214] br[214] wl[5] vdd gnd cell_6t
Xbit_r6_c214 bl[214] br[214] wl[6] vdd gnd cell_6t
Xbit_r7_c214 bl[214] br[214] wl[7] vdd gnd cell_6t
Xbit_r8_c214 bl[214] br[214] wl[8] vdd gnd cell_6t
Xbit_r9_c214 bl[214] br[214] wl[9] vdd gnd cell_6t
Xbit_r10_c214 bl[214] br[214] wl[10] vdd gnd cell_6t
Xbit_r11_c214 bl[214] br[214] wl[11] vdd gnd cell_6t
Xbit_r12_c214 bl[214] br[214] wl[12] vdd gnd cell_6t
Xbit_r13_c214 bl[214] br[214] wl[13] vdd gnd cell_6t
Xbit_r14_c214 bl[214] br[214] wl[14] vdd gnd cell_6t
Xbit_r15_c214 bl[214] br[214] wl[15] vdd gnd cell_6t
Xbit_r16_c214 bl[214] br[214] wl[16] vdd gnd cell_6t
Xbit_r17_c214 bl[214] br[214] wl[17] vdd gnd cell_6t
Xbit_r18_c214 bl[214] br[214] wl[18] vdd gnd cell_6t
Xbit_r19_c214 bl[214] br[214] wl[19] vdd gnd cell_6t
Xbit_r20_c214 bl[214] br[214] wl[20] vdd gnd cell_6t
Xbit_r21_c214 bl[214] br[214] wl[21] vdd gnd cell_6t
Xbit_r22_c214 bl[214] br[214] wl[22] vdd gnd cell_6t
Xbit_r23_c214 bl[214] br[214] wl[23] vdd gnd cell_6t
Xbit_r24_c214 bl[214] br[214] wl[24] vdd gnd cell_6t
Xbit_r25_c214 bl[214] br[214] wl[25] vdd gnd cell_6t
Xbit_r26_c214 bl[214] br[214] wl[26] vdd gnd cell_6t
Xbit_r27_c214 bl[214] br[214] wl[27] vdd gnd cell_6t
Xbit_r28_c214 bl[214] br[214] wl[28] vdd gnd cell_6t
Xbit_r29_c214 bl[214] br[214] wl[29] vdd gnd cell_6t
Xbit_r30_c214 bl[214] br[214] wl[30] vdd gnd cell_6t
Xbit_r31_c214 bl[214] br[214] wl[31] vdd gnd cell_6t
Xbit_r32_c214 bl[214] br[214] wl[32] vdd gnd cell_6t
Xbit_r33_c214 bl[214] br[214] wl[33] vdd gnd cell_6t
Xbit_r34_c214 bl[214] br[214] wl[34] vdd gnd cell_6t
Xbit_r35_c214 bl[214] br[214] wl[35] vdd gnd cell_6t
Xbit_r36_c214 bl[214] br[214] wl[36] vdd gnd cell_6t
Xbit_r37_c214 bl[214] br[214] wl[37] vdd gnd cell_6t
Xbit_r38_c214 bl[214] br[214] wl[38] vdd gnd cell_6t
Xbit_r39_c214 bl[214] br[214] wl[39] vdd gnd cell_6t
Xbit_r40_c214 bl[214] br[214] wl[40] vdd gnd cell_6t
Xbit_r41_c214 bl[214] br[214] wl[41] vdd gnd cell_6t
Xbit_r42_c214 bl[214] br[214] wl[42] vdd gnd cell_6t
Xbit_r43_c214 bl[214] br[214] wl[43] vdd gnd cell_6t
Xbit_r44_c214 bl[214] br[214] wl[44] vdd gnd cell_6t
Xbit_r45_c214 bl[214] br[214] wl[45] vdd gnd cell_6t
Xbit_r46_c214 bl[214] br[214] wl[46] vdd gnd cell_6t
Xbit_r47_c214 bl[214] br[214] wl[47] vdd gnd cell_6t
Xbit_r48_c214 bl[214] br[214] wl[48] vdd gnd cell_6t
Xbit_r49_c214 bl[214] br[214] wl[49] vdd gnd cell_6t
Xbit_r50_c214 bl[214] br[214] wl[50] vdd gnd cell_6t
Xbit_r51_c214 bl[214] br[214] wl[51] vdd gnd cell_6t
Xbit_r52_c214 bl[214] br[214] wl[52] vdd gnd cell_6t
Xbit_r53_c214 bl[214] br[214] wl[53] vdd gnd cell_6t
Xbit_r54_c214 bl[214] br[214] wl[54] vdd gnd cell_6t
Xbit_r55_c214 bl[214] br[214] wl[55] vdd gnd cell_6t
Xbit_r56_c214 bl[214] br[214] wl[56] vdd gnd cell_6t
Xbit_r57_c214 bl[214] br[214] wl[57] vdd gnd cell_6t
Xbit_r58_c214 bl[214] br[214] wl[58] vdd gnd cell_6t
Xbit_r59_c214 bl[214] br[214] wl[59] vdd gnd cell_6t
Xbit_r60_c214 bl[214] br[214] wl[60] vdd gnd cell_6t
Xbit_r61_c214 bl[214] br[214] wl[61] vdd gnd cell_6t
Xbit_r62_c214 bl[214] br[214] wl[62] vdd gnd cell_6t
Xbit_r63_c214 bl[214] br[214] wl[63] vdd gnd cell_6t
Xbit_r64_c214 bl[214] br[214] wl[64] vdd gnd cell_6t
Xbit_r65_c214 bl[214] br[214] wl[65] vdd gnd cell_6t
Xbit_r66_c214 bl[214] br[214] wl[66] vdd gnd cell_6t
Xbit_r67_c214 bl[214] br[214] wl[67] vdd gnd cell_6t
Xbit_r68_c214 bl[214] br[214] wl[68] vdd gnd cell_6t
Xbit_r69_c214 bl[214] br[214] wl[69] vdd gnd cell_6t
Xbit_r70_c214 bl[214] br[214] wl[70] vdd gnd cell_6t
Xbit_r71_c214 bl[214] br[214] wl[71] vdd gnd cell_6t
Xbit_r72_c214 bl[214] br[214] wl[72] vdd gnd cell_6t
Xbit_r73_c214 bl[214] br[214] wl[73] vdd gnd cell_6t
Xbit_r74_c214 bl[214] br[214] wl[74] vdd gnd cell_6t
Xbit_r75_c214 bl[214] br[214] wl[75] vdd gnd cell_6t
Xbit_r76_c214 bl[214] br[214] wl[76] vdd gnd cell_6t
Xbit_r77_c214 bl[214] br[214] wl[77] vdd gnd cell_6t
Xbit_r78_c214 bl[214] br[214] wl[78] vdd gnd cell_6t
Xbit_r79_c214 bl[214] br[214] wl[79] vdd gnd cell_6t
Xbit_r80_c214 bl[214] br[214] wl[80] vdd gnd cell_6t
Xbit_r81_c214 bl[214] br[214] wl[81] vdd gnd cell_6t
Xbit_r82_c214 bl[214] br[214] wl[82] vdd gnd cell_6t
Xbit_r83_c214 bl[214] br[214] wl[83] vdd gnd cell_6t
Xbit_r84_c214 bl[214] br[214] wl[84] vdd gnd cell_6t
Xbit_r85_c214 bl[214] br[214] wl[85] vdd gnd cell_6t
Xbit_r86_c214 bl[214] br[214] wl[86] vdd gnd cell_6t
Xbit_r87_c214 bl[214] br[214] wl[87] vdd gnd cell_6t
Xbit_r88_c214 bl[214] br[214] wl[88] vdd gnd cell_6t
Xbit_r89_c214 bl[214] br[214] wl[89] vdd gnd cell_6t
Xbit_r90_c214 bl[214] br[214] wl[90] vdd gnd cell_6t
Xbit_r91_c214 bl[214] br[214] wl[91] vdd gnd cell_6t
Xbit_r92_c214 bl[214] br[214] wl[92] vdd gnd cell_6t
Xbit_r93_c214 bl[214] br[214] wl[93] vdd gnd cell_6t
Xbit_r94_c214 bl[214] br[214] wl[94] vdd gnd cell_6t
Xbit_r95_c214 bl[214] br[214] wl[95] vdd gnd cell_6t
Xbit_r96_c214 bl[214] br[214] wl[96] vdd gnd cell_6t
Xbit_r97_c214 bl[214] br[214] wl[97] vdd gnd cell_6t
Xbit_r98_c214 bl[214] br[214] wl[98] vdd gnd cell_6t
Xbit_r99_c214 bl[214] br[214] wl[99] vdd gnd cell_6t
Xbit_r100_c214 bl[214] br[214] wl[100] vdd gnd cell_6t
Xbit_r101_c214 bl[214] br[214] wl[101] vdd gnd cell_6t
Xbit_r102_c214 bl[214] br[214] wl[102] vdd gnd cell_6t
Xbit_r103_c214 bl[214] br[214] wl[103] vdd gnd cell_6t
Xbit_r104_c214 bl[214] br[214] wl[104] vdd gnd cell_6t
Xbit_r105_c214 bl[214] br[214] wl[105] vdd gnd cell_6t
Xbit_r106_c214 bl[214] br[214] wl[106] vdd gnd cell_6t
Xbit_r107_c214 bl[214] br[214] wl[107] vdd gnd cell_6t
Xbit_r108_c214 bl[214] br[214] wl[108] vdd gnd cell_6t
Xbit_r109_c214 bl[214] br[214] wl[109] vdd gnd cell_6t
Xbit_r110_c214 bl[214] br[214] wl[110] vdd gnd cell_6t
Xbit_r111_c214 bl[214] br[214] wl[111] vdd gnd cell_6t
Xbit_r112_c214 bl[214] br[214] wl[112] vdd gnd cell_6t
Xbit_r113_c214 bl[214] br[214] wl[113] vdd gnd cell_6t
Xbit_r114_c214 bl[214] br[214] wl[114] vdd gnd cell_6t
Xbit_r115_c214 bl[214] br[214] wl[115] vdd gnd cell_6t
Xbit_r116_c214 bl[214] br[214] wl[116] vdd gnd cell_6t
Xbit_r117_c214 bl[214] br[214] wl[117] vdd gnd cell_6t
Xbit_r118_c214 bl[214] br[214] wl[118] vdd gnd cell_6t
Xbit_r119_c214 bl[214] br[214] wl[119] vdd gnd cell_6t
Xbit_r120_c214 bl[214] br[214] wl[120] vdd gnd cell_6t
Xbit_r121_c214 bl[214] br[214] wl[121] vdd gnd cell_6t
Xbit_r122_c214 bl[214] br[214] wl[122] vdd gnd cell_6t
Xbit_r123_c214 bl[214] br[214] wl[123] vdd gnd cell_6t
Xbit_r124_c214 bl[214] br[214] wl[124] vdd gnd cell_6t
Xbit_r125_c214 bl[214] br[214] wl[125] vdd gnd cell_6t
Xbit_r126_c214 bl[214] br[214] wl[126] vdd gnd cell_6t
Xbit_r127_c214 bl[214] br[214] wl[127] vdd gnd cell_6t
Xbit_r0_c215 bl[215] br[215] wl[0] vdd gnd cell_6t
Xbit_r1_c215 bl[215] br[215] wl[1] vdd gnd cell_6t
Xbit_r2_c215 bl[215] br[215] wl[2] vdd gnd cell_6t
Xbit_r3_c215 bl[215] br[215] wl[3] vdd gnd cell_6t
Xbit_r4_c215 bl[215] br[215] wl[4] vdd gnd cell_6t
Xbit_r5_c215 bl[215] br[215] wl[5] vdd gnd cell_6t
Xbit_r6_c215 bl[215] br[215] wl[6] vdd gnd cell_6t
Xbit_r7_c215 bl[215] br[215] wl[7] vdd gnd cell_6t
Xbit_r8_c215 bl[215] br[215] wl[8] vdd gnd cell_6t
Xbit_r9_c215 bl[215] br[215] wl[9] vdd gnd cell_6t
Xbit_r10_c215 bl[215] br[215] wl[10] vdd gnd cell_6t
Xbit_r11_c215 bl[215] br[215] wl[11] vdd gnd cell_6t
Xbit_r12_c215 bl[215] br[215] wl[12] vdd gnd cell_6t
Xbit_r13_c215 bl[215] br[215] wl[13] vdd gnd cell_6t
Xbit_r14_c215 bl[215] br[215] wl[14] vdd gnd cell_6t
Xbit_r15_c215 bl[215] br[215] wl[15] vdd gnd cell_6t
Xbit_r16_c215 bl[215] br[215] wl[16] vdd gnd cell_6t
Xbit_r17_c215 bl[215] br[215] wl[17] vdd gnd cell_6t
Xbit_r18_c215 bl[215] br[215] wl[18] vdd gnd cell_6t
Xbit_r19_c215 bl[215] br[215] wl[19] vdd gnd cell_6t
Xbit_r20_c215 bl[215] br[215] wl[20] vdd gnd cell_6t
Xbit_r21_c215 bl[215] br[215] wl[21] vdd gnd cell_6t
Xbit_r22_c215 bl[215] br[215] wl[22] vdd gnd cell_6t
Xbit_r23_c215 bl[215] br[215] wl[23] vdd gnd cell_6t
Xbit_r24_c215 bl[215] br[215] wl[24] vdd gnd cell_6t
Xbit_r25_c215 bl[215] br[215] wl[25] vdd gnd cell_6t
Xbit_r26_c215 bl[215] br[215] wl[26] vdd gnd cell_6t
Xbit_r27_c215 bl[215] br[215] wl[27] vdd gnd cell_6t
Xbit_r28_c215 bl[215] br[215] wl[28] vdd gnd cell_6t
Xbit_r29_c215 bl[215] br[215] wl[29] vdd gnd cell_6t
Xbit_r30_c215 bl[215] br[215] wl[30] vdd gnd cell_6t
Xbit_r31_c215 bl[215] br[215] wl[31] vdd gnd cell_6t
Xbit_r32_c215 bl[215] br[215] wl[32] vdd gnd cell_6t
Xbit_r33_c215 bl[215] br[215] wl[33] vdd gnd cell_6t
Xbit_r34_c215 bl[215] br[215] wl[34] vdd gnd cell_6t
Xbit_r35_c215 bl[215] br[215] wl[35] vdd gnd cell_6t
Xbit_r36_c215 bl[215] br[215] wl[36] vdd gnd cell_6t
Xbit_r37_c215 bl[215] br[215] wl[37] vdd gnd cell_6t
Xbit_r38_c215 bl[215] br[215] wl[38] vdd gnd cell_6t
Xbit_r39_c215 bl[215] br[215] wl[39] vdd gnd cell_6t
Xbit_r40_c215 bl[215] br[215] wl[40] vdd gnd cell_6t
Xbit_r41_c215 bl[215] br[215] wl[41] vdd gnd cell_6t
Xbit_r42_c215 bl[215] br[215] wl[42] vdd gnd cell_6t
Xbit_r43_c215 bl[215] br[215] wl[43] vdd gnd cell_6t
Xbit_r44_c215 bl[215] br[215] wl[44] vdd gnd cell_6t
Xbit_r45_c215 bl[215] br[215] wl[45] vdd gnd cell_6t
Xbit_r46_c215 bl[215] br[215] wl[46] vdd gnd cell_6t
Xbit_r47_c215 bl[215] br[215] wl[47] vdd gnd cell_6t
Xbit_r48_c215 bl[215] br[215] wl[48] vdd gnd cell_6t
Xbit_r49_c215 bl[215] br[215] wl[49] vdd gnd cell_6t
Xbit_r50_c215 bl[215] br[215] wl[50] vdd gnd cell_6t
Xbit_r51_c215 bl[215] br[215] wl[51] vdd gnd cell_6t
Xbit_r52_c215 bl[215] br[215] wl[52] vdd gnd cell_6t
Xbit_r53_c215 bl[215] br[215] wl[53] vdd gnd cell_6t
Xbit_r54_c215 bl[215] br[215] wl[54] vdd gnd cell_6t
Xbit_r55_c215 bl[215] br[215] wl[55] vdd gnd cell_6t
Xbit_r56_c215 bl[215] br[215] wl[56] vdd gnd cell_6t
Xbit_r57_c215 bl[215] br[215] wl[57] vdd gnd cell_6t
Xbit_r58_c215 bl[215] br[215] wl[58] vdd gnd cell_6t
Xbit_r59_c215 bl[215] br[215] wl[59] vdd gnd cell_6t
Xbit_r60_c215 bl[215] br[215] wl[60] vdd gnd cell_6t
Xbit_r61_c215 bl[215] br[215] wl[61] vdd gnd cell_6t
Xbit_r62_c215 bl[215] br[215] wl[62] vdd gnd cell_6t
Xbit_r63_c215 bl[215] br[215] wl[63] vdd gnd cell_6t
Xbit_r64_c215 bl[215] br[215] wl[64] vdd gnd cell_6t
Xbit_r65_c215 bl[215] br[215] wl[65] vdd gnd cell_6t
Xbit_r66_c215 bl[215] br[215] wl[66] vdd gnd cell_6t
Xbit_r67_c215 bl[215] br[215] wl[67] vdd gnd cell_6t
Xbit_r68_c215 bl[215] br[215] wl[68] vdd gnd cell_6t
Xbit_r69_c215 bl[215] br[215] wl[69] vdd gnd cell_6t
Xbit_r70_c215 bl[215] br[215] wl[70] vdd gnd cell_6t
Xbit_r71_c215 bl[215] br[215] wl[71] vdd gnd cell_6t
Xbit_r72_c215 bl[215] br[215] wl[72] vdd gnd cell_6t
Xbit_r73_c215 bl[215] br[215] wl[73] vdd gnd cell_6t
Xbit_r74_c215 bl[215] br[215] wl[74] vdd gnd cell_6t
Xbit_r75_c215 bl[215] br[215] wl[75] vdd gnd cell_6t
Xbit_r76_c215 bl[215] br[215] wl[76] vdd gnd cell_6t
Xbit_r77_c215 bl[215] br[215] wl[77] vdd gnd cell_6t
Xbit_r78_c215 bl[215] br[215] wl[78] vdd gnd cell_6t
Xbit_r79_c215 bl[215] br[215] wl[79] vdd gnd cell_6t
Xbit_r80_c215 bl[215] br[215] wl[80] vdd gnd cell_6t
Xbit_r81_c215 bl[215] br[215] wl[81] vdd gnd cell_6t
Xbit_r82_c215 bl[215] br[215] wl[82] vdd gnd cell_6t
Xbit_r83_c215 bl[215] br[215] wl[83] vdd gnd cell_6t
Xbit_r84_c215 bl[215] br[215] wl[84] vdd gnd cell_6t
Xbit_r85_c215 bl[215] br[215] wl[85] vdd gnd cell_6t
Xbit_r86_c215 bl[215] br[215] wl[86] vdd gnd cell_6t
Xbit_r87_c215 bl[215] br[215] wl[87] vdd gnd cell_6t
Xbit_r88_c215 bl[215] br[215] wl[88] vdd gnd cell_6t
Xbit_r89_c215 bl[215] br[215] wl[89] vdd gnd cell_6t
Xbit_r90_c215 bl[215] br[215] wl[90] vdd gnd cell_6t
Xbit_r91_c215 bl[215] br[215] wl[91] vdd gnd cell_6t
Xbit_r92_c215 bl[215] br[215] wl[92] vdd gnd cell_6t
Xbit_r93_c215 bl[215] br[215] wl[93] vdd gnd cell_6t
Xbit_r94_c215 bl[215] br[215] wl[94] vdd gnd cell_6t
Xbit_r95_c215 bl[215] br[215] wl[95] vdd gnd cell_6t
Xbit_r96_c215 bl[215] br[215] wl[96] vdd gnd cell_6t
Xbit_r97_c215 bl[215] br[215] wl[97] vdd gnd cell_6t
Xbit_r98_c215 bl[215] br[215] wl[98] vdd gnd cell_6t
Xbit_r99_c215 bl[215] br[215] wl[99] vdd gnd cell_6t
Xbit_r100_c215 bl[215] br[215] wl[100] vdd gnd cell_6t
Xbit_r101_c215 bl[215] br[215] wl[101] vdd gnd cell_6t
Xbit_r102_c215 bl[215] br[215] wl[102] vdd gnd cell_6t
Xbit_r103_c215 bl[215] br[215] wl[103] vdd gnd cell_6t
Xbit_r104_c215 bl[215] br[215] wl[104] vdd gnd cell_6t
Xbit_r105_c215 bl[215] br[215] wl[105] vdd gnd cell_6t
Xbit_r106_c215 bl[215] br[215] wl[106] vdd gnd cell_6t
Xbit_r107_c215 bl[215] br[215] wl[107] vdd gnd cell_6t
Xbit_r108_c215 bl[215] br[215] wl[108] vdd gnd cell_6t
Xbit_r109_c215 bl[215] br[215] wl[109] vdd gnd cell_6t
Xbit_r110_c215 bl[215] br[215] wl[110] vdd gnd cell_6t
Xbit_r111_c215 bl[215] br[215] wl[111] vdd gnd cell_6t
Xbit_r112_c215 bl[215] br[215] wl[112] vdd gnd cell_6t
Xbit_r113_c215 bl[215] br[215] wl[113] vdd gnd cell_6t
Xbit_r114_c215 bl[215] br[215] wl[114] vdd gnd cell_6t
Xbit_r115_c215 bl[215] br[215] wl[115] vdd gnd cell_6t
Xbit_r116_c215 bl[215] br[215] wl[116] vdd gnd cell_6t
Xbit_r117_c215 bl[215] br[215] wl[117] vdd gnd cell_6t
Xbit_r118_c215 bl[215] br[215] wl[118] vdd gnd cell_6t
Xbit_r119_c215 bl[215] br[215] wl[119] vdd gnd cell_6t
Xbit_r120_c215 bl[215] br[215] wl[120] vdd gnd cell_6t
Xbit_r121_c215 bl[215] br[215] wl[121] vdd gnd cell_6t
Xbit_r122_c215 bl[215] br[215] wl[122] vdd gnd cell_6t
Xbit_r123_c215 bl[215] br[215] wl[123] vdd gnd cell_6t
Xbit_r124_c215 bl[215] br[215] wl[124] vdd gnd cell_6t
Xbit_r125_c215 bl[215] br[215] wl[125] vdd gnd cell_6t
Xbit_r126_c215 bl[215] br[215] wl[126] vdd gnd cell_6t
Xbit_r127_c215 bl[215] br[215] wl[127] vdd gnd cell_6t
Xbit_r0_c216 bl[216] br[216] wl[0] vdd gnd cell_6t
Xbit_r1_c216 bl[216] br[216] wl[1] vdd gnd cell_6t
Xbit_r2_c216 bl[216] br[216] wl[2] vdd gnd cell_6t
Xbit_r3_c216 bl[216] br[216] wl[3] vdd gnd cell_6t
Xbit_r4_c216 bl[216] br[216] wl[4] vdd gnd cell_6t
Xbit_r5_c216 bl[216] br[216] wl[5] vdd gnd cell_6t
Xbit_r6_c216 bl[216] br[216] wl[6] vdd gnd cell_6t
Xbit_r7_c216 bl[216] br[216] wl[7] vdd gnd cell_6t
Xbit_r8_c216 bl[216] br[216] wl[8] vdd gnd cell_6t
Xbit_r9_c216 bl[216] br[216] wl[9] vdd gnd cell_6t
Xbit_r10_c216 bl[216] br[216] wl[10] vdd gnd cell_6t
Xbit_r11_c216 bl[216] br[216] wl[11] vdd gnd cell_6t
Xbit_r12_c216 bl[216] br[216] wl[12] vdd gnd cell_6t
Xbit_r13_c216 bl[216] br[216] wl[13] vdd gnd cell_6t
Xbit_r14_c216 bl[216] br[216] wl[14] vdd gnd cell_6t
Xbit_r15_c216 bl[216] br[216] wl[15] vdd gnd cell_6t
Xbit_r16_c216 bl[216] br[216] wl[16] vdd gnd cell_6t
Xbit_r17_c216 bl[216] br[216] wl[17] vdd gnd cell_6t
Xbit_r18_c216 bl[216] br[216] wl[18] vdd gnd cell_6t
Xbit_r19_c216 bl[216] br[216] wl[19] vdd gnd cell_6t
Xbit_r20_c216 bl[216] br[216] wl[20] vdd gnd cell_6t
Xbit_r21_c216 bl[216] br[216] wl[21] vdd gnd cell_6t
Xbit_r22_c216 bl[216] br[216] wl[22] vdd gnd cell_6t
Xbit_r23_c216 bl[216] br[216] wl[23] vdd gnd cell_6t
Xbit_r24_c216 bl[216] br[216] wl[24] vdd gnd cell_6t
Xbit_r25_c216 bl[216] br[216] wl[25] vdd gnd cell_6t
Xbit_r26_c216 bl[216] br[216] wl[26] vdd gnd cell_6t
Xbit_r27_c216 bl[216] br[216] wl[27] vdd gnd cell_6t
Xbit_r28_c216 bl[216] br[216] wl[28] vdd gnd cell_6t
Xbit_r29_c216 bl[216] br[216] wl[29] vdd gnd cell_6t
Xbit_r30_c216 bl[216] br[216] wl[30] vdd gnd cell_6t
Xbit_r31_c216 bl[216] br[216] wl[31] vdd gnd cell_6t
Xbit_r32_c216 bl[216] br[216] wl[32] vdd gnd cell_6t
Xbit_r33_c216 bl[216] br[216] wl[33] vdd gnd cell_6t
Xbit_r34_c216 bl[216] br[216] wl[34] vdd gnd cell_6t
Xbit_r35_c216 bl[216] br[216] wl[35] vdd gnd cell_6t
Xbit_r36_c216 bl[216] br[216] wl[36] vdd gnd cell_6t
Xbit_r37_c216 bl[216] br[216] wl[37] vdd gnd cell_6t
Xbit_r38_c216 bl[216] br[216] wl[38] vdd gnd cell_6t
Xbit_r39_c216 bl[216] br[216] wl[39] vdd gnd cell_6t
Xbit_r40_c216 bl[216] br[216] wl[40] vdd gnd cell_6t
Xbit_r41_c216 bl[216] br[216] wl[41] vdd gnd cell_6t
Xbit_r42_c216 bl[216] br[216] wl[42] vdd gnd cell_6t
Xbit_r43_c216 bl[216] br[216] wl[43] vdd gnd cell_6t
Xbit_r44_c216 bl[216] br[216] wl[44] vdd gnd cell_6t
Xbit_r45_c216 bl[216] br[216] wl[45] vdd gnd cell_6t
Xbit_r46_c216 bl[216] br[216] wl[46] vdd gnd cell_6t
Xbit_r47_c216 bl[216] br[216] wl[47] vdd gnd cell_6t
Xbit_r48_c216 bl[216] br[216] wl[48] vdd gnd cell_6t
Xbit_r49_c216 bl[216] br[216] wl[49] vdd gnd cell_6t
Xbit_r50_c216 bl[216] br[216] wl[50] vdd gnd cell_6t
Xbit_r51_c216 bl[216] br[216] wl[51] vdd gnd cell_6t
Xbit_r52_c216 bl[216] br[216] wl[52] vdd gnd cell_6t
Xbit_r53_c216 bl[216] br[216] wl[53] vdd gnd cell_6t
Xbit_r54_c216 bl[216] br[216] wl[54] vdd gnd cell_6t
Xbit_r55_c216 bl[216] br[216] wl[55] vdd gnd cell_6t
Xbit_r56_c216 bl[216] br[216] wl[56] vdd gnd cell_6t
Xbit_r57_c216 bl[216] br[216] wl[57] vdd gnd cell_6t
Xbit_r58_c216 bl[216] br[216] wl[58] vdd gnd cell_6t
Xbit_r59_c216 bl[216] br[216] wl[59] vdd gnd cell_6t
Xbit_r60_c216 bl[216] br[216] wl[60] vdd gnd cell_6t
Xbit_r61_c216 bl[216] br[216] wl[61] vdd gnd cell_6t
Xbit_r62_c216 bl[216] br[216] wl[62] vdd gnd cell_6t
Xbit_r63_c216 bl[216] br[216] wl[63] vdd gnd cell_6t
Xbit_r64_c216 bl[216] br[216] wl[64] vdd gnd cell_6t
Xbit_r65_c216 bl[216] br[216] wl[65] vdd gnd cell_6t
Xbit_r66_c216 bl[216] br[216] wl[66] vdd gnd cell_6t
Xbit_r67_c216 bl[216] br[216] wl[67] vdd gnd cell_6t
Xbit_r68_c216 bl[216] br[216] wl[68] vdd gnd cell_6t
Xbit_r69_c216 bl[216] br[216] wl[69] vdd gnd cell_6t
Xbit_r70_c216 bl[216] br[216] wl[70] vdd gnd cell_6t
Xbit_r71_c216 bl[216] br[216] wl[71] vdd gnd cell_6t
Xbit_r72_c216 bl[216] br[216] wl[72] vdd gnd cell_6t
Xbit_r73_c216 bl[216] br[216] wl[73] vdd gnd cell_6t
Xbit_r74_c216 bl[216] br[216] wl[74] vdd gnd cell_6t
Xbit_r75_c216 bl[216] br[216] wl[75] vdd gnd cell_6t
Xbit_r76_c216 bl[216] br[216] wl[76] vdd gnd cell_6t
Xbit_r77_c216 bl[216] br[216] wl[77] vdd gnd cell_6t
Xbit_r78_c216 bl[216] br[216] wl[78] vdd gnd cell_6t
Xbit_r79_c216 bl[216] br[216] wl[79] vdd gnd cell_6t
Xbit_r80_c216 bl[216] br[216] wl[80] vdd gnd cell_6t
Xbit_r81_c216 bl[216] br[216] wl[81] vdd gnd cell_6t
Xbit_r82_c216 bl[216] br[216] wl[82] vdd gnd cell_6t
Xbit_r83_c216 bl[216] br[216] wl[83] vdd gnd cell_6t
Xbit_r84_c216 bl[216] br[216] wl[84] vdd gnd cell_6t
Xbit_r85_c216 bl[216] br[216] wl[85] vdd gnd cell_6t
Xbit_r86_c216 bl[216] br[216] wl[86] vdd gnd cell_6t
Xbit_r87_c216 bl[216] br[216] wl[87] vdd gnd cell_6t
Xbit_r88_c216 bl[216] br[216] wl[88] vdd gnd cell_6t
Xbit_r89_c216 bl[216] br[216] wl[89] vdd gnd cell_6t
Xbit_r90_c216 bl[216] br[216] wl[90] vdd gnd cell_6t
Xbit_r91_c216 bl[216] br[216] wl[91] vdd gnd cell_6t
Xbit_r92_c216 bl[216] br[216] wl[92] vdd gnd cell_6t
Xbit_r93_c216 bl[216] br[216] wl[93] vdd gnd cell_6t
Xbit_r94_c216 bl[216] br[216] wl[94] vdd gnd cell_6t
Xbit_r95_c216 bl[216] br[216] wl[95] vdd gnd cell_6t
Xbit_r96_c216 bl[216] br[216] wl[96] vdd gnd cell_6t
Xbit_r97_c216 bl[216] br[216] wl[97] vdd gnd cell_6t
Xbit_r98_c216 bl[216] br[216] wl[98] vdd gnd cell_6t
Xbit_r99_c216 bl[216] br[216] wl[99] vdd gnd cell_6t
Xbit_r100_c216 bl[216] br[216] wl[100] vdd gnd cell_6t
Xbit_r101_c216 bl[216] br[216] wl[101] vdd gnd cell_6t
Xbit_r102_c216 bl[216] br[216] wl[102] vdd gnd cell_6t
Xbit_r103_c216 bl[216] br[216] wl[103] vdd gnd cell_6t
Xbit_r104_c216 bl[216] br[216] wl[104] vdd gnd cell_6t
Xbit_r105_c216 bl[216] br[216] wl[105] vdd gnd cell_6t
Xbit_r106_c216 bl[216] br[216] wl[106] vdd gnd cell_6t
Xbit_r107_c216 bl[216] br[216] wl[107] vdd gnd cell_6t
Xbit_r108_c216 bl[216] br[216] wl[108] vdd gnd cell_6t
Xbit_r109_c216 bl[216] br[216] wl[109] vdd gnd cell_6t
Xbit_r110_c216 bl[216] br[216] wl[110] vdd gnd cell_6t
Xbit_r111_c216 bl[216] br[216] wl[111] vdd gnd cell_6t
Xbit_r112_c216 bl[216] br[216] wl[112] vdd gnd cell_6t
Xbit_r113_c216 bl[216] br[216] wl[113] vdd gnd cell_6t
Xbit_r114_c216 bl[216] br[216] wl[114] vdd gnd cell_6t
Xbit_r115_c216 bl[216] br[216] wl[115] vdd gnd cell_6t
Xbit_r116_c216 bl[216] br[216] wl[116] vdd gnd cell_6t
Xbit_r117_c216 bl[216] br[216] wl[117] vdd gnd cell_6t
Xbit_r118_c216 bl[216] br[216] wl[118] vdd gnd cell_6t
Xbit_r119_c216 bl[216] br[216] wl[119] vdd gnd cell_6t
Xbit_r120_c216 bl[216] br[216] wl[120] vdd gnd cell_6t
Xbit_r121_c216 bl[216] br[216] wl[121] vdd gnd cell_6t
Xbit_r122_c216 bl[216] br[216] wl[122] vdd gnd cell_6t
Xbit_r123_c216 bl[216] br[216] wl[123] vdd gnd cell_6t
Xbit_r124_c216 bl[216] br[216] wl[124] vdd gnd cell_6t
Xbit_r125_c216 bl[216] br[216] wl[125] vdd gnd cell_6t
Xbit_r126_c216 bl[216] br[216] wl[126] vdd gnd cell_6t
Xbit_r127_c216 bl[216] br[216] wl[127] vdd gnd cell_6t
Xbit_r0_c217 bl[217] br[217] wl[0] vdd gnd cell_6t
Xbit_r1_c217 bl[217] br[217] wl[1] vdd gnd cell_6t
Xbit_r2_c217 bl[217] br[217] wl[2] vdd gnd cell_6t
Xbit_r3_c217 bl[217] br[217] wl[3] vdd gnd cell_6t
Xbit_r4_c217 bl[217] br[217] wl[4] vdd gnd cell_6t
Xbit_r5_c217 bl[217] br[217] wl[5] vdd gnd cell_6t
Xbit_r6_c217 bl[217] br[217] wl[6] vdd gnd cell_6t
Xbit_r7_c217 bl[217] br[217] wl[7] vdd gnd cell_6t
Xbit_r8_c217 bl[217] br[217] wl[8] vdd gnd cell_6t
Xbit_r9_c217 bl[217] br[217] wl[9] vdd gnd cell_6t
Xbit_r10_c217 bl[217] br[217] wl[10] vdd gnd cell_6t
Xbit_r11_c217 bl[217] br[217] wl[11] vdd gnd cell_6t
Xbit_r12_c217 bl[217] br[217] wl[12] vdd gnd cell_6t
Xbit_r13_c217 bl[217] br[217] wl[13] vdd gnd cell_6t
Xbit_r14_c217 bl[217] br[217] wl[14] vdd gnd cell_6t
Xbit_r15_c217 bl[217] br[217] wl[15] vdd gnd cell_6t
Xbit_r16_c217 bl[217] br[217] wl[16] vdd gnd cell_6t
Xbit_r17_c217 bl[217] br[217] wl[17] vdd gnd cell_6t
Xbit_r18_c217 bl[217] br[217] wl[18] vdd gnd cell_6t
Xbit_r19_c217 bl[217] br[217] wl[19] vdd gnd cell_6t
Xbit_r20_c217 bl[217] br[217] wl[20] vdd gnd cell_6t
Xbit_r21_c217 bl[217] br[217] wl[21] vdd gnd cell_6t
Xbit_r22_c217 bl[217] br[217] wl[22] vdd gnd cell_6t
Xbit_r23_c217 bl[217] br[217] wl[23] vdd gnd cell_6t
Xbit_r24_c217 bl[217] br[217] wl[24] vdd gnd cell_6t
Xbit_r25_c217 bl[217] br[217] wl[25] vdd gnd cell_6t
Xbit_r26_c217 bl[217] br[217] wl[26] vdd gnd cell_6t
Xbit_r27_c217 bl[217] br[217] wl[27] vdd gnd cell_6t
Xbit_r28_c217 bl[217] br[217] wl[28] vdd gnd cell_6t
Xbit_r29_c217 bl[217] br[217] wl[29] vdd gnd cell_6t
Xbit_r30_c217 bl[217] br[217] wl[30] vdd gnd cell_6t
Xbit_r31_c217 bl[217] br[217] wl[31] vdd gnd cell_6t
Xbit_r32_c217 bl[217] br[217] wl[32] vdd gnd cell_6t
Xbit_r33_c217 bl[217] br[217] wl[33] vdd gnd cell_6t
Xbit_r34_c217 bl[217] br[217] wl[34] vdd gnd cell_6t
Xbit_r35_c217 bl[217] br[217] wl[35] vdd gnd cell_6t
Xbit_r36_c217 bl[217] br[217] wl[36] vdd gnd cell_6t
Xbit_r37_c217 bl[217] br[217] wl[37] vdd gnd cell_6t
Xbit_r38_c217 bl[217] br[217] wl[38] vdd gnd cell_6t
Xbit_r39_c217 bl[217] br[217] wl[39] vdd gnd cell_6t
Xbit_r40_c217 bl[217] br[217] wl[40] vdd gnd cell_6t
Xbit_r41_c217 bl[217] br[217] wl[41] vdd gnd cell_6t
Xbit_r42_c217 bl[217] br[217] wl[42] vdd gnd cell_6t
Xbit_r43_c217 bl[217] br[217] wl[43] vdd gnd cell_6t
Xbit_r44_c217 bl[217] br[217] wl[44] vdd gnd cell_6t
Xbit_r45_c217 bl[217] br[217] wl[45] vdd gnd cell_6t
Xbit_r46_c217 bl[217] br[217] wl[46] vdd gnd cell_6t
Xbit_r47_c217 bl[217] br[217] wl[47] vdd gnd cell_6t
Xbit_r48_c217 bl[217] br[217] wl[48] vdd gnd cell_6t
Xbit_r49_c217 bl[217] br[217] wl[49] vdd gnd cell_6t
Xbit_r50_c217 bl[217] br[217] wl[50] vdd gnd cell_6t
Xbit_r51_c217 bl[217] br[217] wl[51] vdd gnd cell_6t
Xbit_r52_c217 bl[217] br[217] wl[52] vdd gnd cell_6t
Xbit_r53_c217 bl[217] br[217] wl[53] vdd gnd cell_6t
Xbit_r54_c217 bl[217] br[217] wl[54] vdd gnd cell_6t
Xbit_r55_c217 bl[217] br[217] wl[55] vdd gnd cell_6t
Xbit_r56_c217 bl[217] br[217] wl[56] vdd gnd cell_6t
Xbit_r57_c217 bl[217] br[217] wl[57] vdd gnd cell_6t
Xbit_r58_c217 bl[217] br[217] wl[58] vdd gnd cell_6t
Xbit_r59_c217 bl[217] br[217] wl[59] vdd gnd cell_6t
Xbit_r60_c217 bl[217] br[217] wl[60] vdd gnd cell_6t
Xbit_r61_c217 bl[217] br[217] wl[61] vdd gnd cell_6t
Xbit_r62_c217 bl[217] br[217] wl[62] vdd gnd cell_6t
Xbit_r63_c217 bl[217] br[217] wl[63] vdd gnd cell_6t
Xbit_r64_c217 bl[217] br[217] wl[64] vdd gnd cell_6t
Xbit_r65_c217 bl[217] br[217] wl[65] vdd gnd cell_6t
Xbit_r66_c217 bl[217] br[217] wl[66] vdd gnd cell_6t
Xbit_r67_c217 bl[217] br[217] wl[67] vdd gnd cell_6t
Xbit_r68_c217 bl[217] br[217] wl[68] vdd gnd cell_6t
Xbit_r69_c217 bl[217] br[217] wl[69] vdd gnd cell_6t
Xbit_r70_c217 bl[217] br[217] wl[70] vdd gnd cell_6t
Xbit_r71_c217 bl[217] br[217] wl[71] vdd gnd cell_6t
Xbit_r72_c217 bl[217] br[217] wl[72] vdd gnd cell_6t
Xbit_r73_c217 bl[217] br[217] wl[73] vdd gnd cell_6t
Xbit_r74_c217 bl[217] br[217] wl[74] vdd gnd cell_6t
Xbit_r75_c217 bl[217] br[217] wl[75] vdd gnd cell_6t
Xbit_r76_c217 bl[217] br[217] wl[76] vdd gnd cell_6t
Xbit_r77_c217 bl[217] br[217] wl[77] vdd gnd cell_6t
Xbit_r78_c217 bl[217] br[217] wl[78] vdd gnd cell_6t
Xbit_r79_c217 bl[217] br[217] wl[79] vdd gnd cell_6t
Xbit_r80_c217 bl[217] br[217] wl[80] vdd gnd cell_6t
Xbit_r81_c217 bl[217] br[217] wl[81] vdd gnd cell_6t
Xbit_r82_c217 bl[217] br[217] wl[82] vdd gnd cell_6t
Xbit_r83_c217 bl[217] br[217] wl[83] vdd gnd cell_6t
Xbit_r84_c217 bl[217] br[217] wl[84] vdd gnd cell_6t
Xbit_r85_c217 bl[217] br[217] wl[85] vdd gnd cell_6t
Xbit_r86_c217 bl[217] br[217] wl[86] vdd gnd cell_6t
Xbit_r87_c217 bl[217] br[217] wl[87] vdd gnd cell_6t
Xbit_r88_c217 bl[217] br[217] wl[88] vdd gnd cell_6t
Xbit_r89_c217 bl[217] br[217] wl[89] vdd gnd cell_6t
Xbit_r90_c217 bl[217] br[217] wl[90] vdd gnd cell_6t
Xbit_r91_c217 bl[217] br[217] wl[91] vdd gnd cell_6t
Xbit_r92_c217 bl[217] br[217] wl[92] vdd gnd cell_6t
Xbit_r93_c217 bl[217] br[217] wl[93] vdd gnd cell_6t
Xbit_r94_c217 bl[217] br[217] wl[94] vdd gnd cell_6t
Xbit_r95_c217 bl[217] br[217] wl[95] vdd gnd cell_6t
Xbit_r96_c217 bl[217] br[217] wl[96] vdd gnd cell_6t
Xbit_r97_c217 bl[217] br[217] wl[97] vdd gnd cell_6t
Xbit_r98_c217 bl[217] br[217] wl[98] vdd gnd cell_6t
Xbit_r99_c217 bl[217] br[217] wl[99] vdd gnd cell_6t
Xbit_r100_c217 bl[217] br[217] wl[100] vdd gnd cell_6t
Xbit_r101_c217 bl[217] br[217] wl[101] vdd gnd cell_6t
Xbit_r102_c217 bl[217] br[217] wl[102] vdd gnd cell_6t
Xbit_r103_c217 bl[217] br[217] wl[103] vdd gnd cell_6t
Xbit_r104_c217 bl[217] br[217] wl[104] vdd gnd cell_6t
Xbit_r105_c217 bl[217] br[217] wl[105] vdd gnd cell_6t
Xbit_r106_c217 bl[217] br[217] wl[106] vdd gnd cell_6t
Xbit_r107_c217 bl[217] br[217] wl[107] vdd gnd cell_6t
Xbit_r108_c217 bl[217] br[217] wl[108] vdd gnd cell_6t
Xbit_r109_c217 bl[217] br[217] wl[109] vdd gnd cell_6t
Xbit_r110_c217 bl[217] br[217] wl[110] vdd gnd cell_6t
Xbit_r111_c217 bl[217] br[217] wl[111] vdd gnd cell_6t
Xbit_r112_c217 bl[217] br[217] wl[112] vdd gnd cell_6t
Xbit_r113_c217 bl[217] br[217] wl[113] vdd gnd cell_6t
Xbit_r114_c217 bl[217] br[217] wl[114] vdd gnd cell_6t
Xbit_r115_c217 bl[217] br[217] wl[115] vdd gnd cell_6t
Xbit_r116_c217 bl[217] br[217] wl[116] vdd gnd cell_6t
Xbit_r117_c217 bl[217] br[217] wl[117] vdd gnd cell_6t
Xbit_r118_c217 bl[217] br[217] wl[118] vdd gnd cell_6t
Xbit_r119_c217 bl[217] br[217] wl[119] vdd gnd cell_6t
Xbit_r120_c217 bl[217] br[217] wl[120] vdd gnd cell_6t
Xbit_r121_c217 bl[217] br[217] wl[121] vdd gnd cell_6t
Xbit_r122_c217 bl[217] br[217] wl[122] vdd gnd cell_6t
Xbit_r123_c217 bl[217] br[217] wl[123] vdd gnd cell_6t
Xbit_r124_c217 bl[217] br[217] wl[124] vdd gnd cell_6t
Xbit_r125_c217 bl[217] br[217] wl[125] vdd gnd cell_6t
Xbit_r126_c217 bl[217] br[217] wl[126] vdd gnd cell_6t
Xbit_r127_c217 bl[217] br[217] wl[127] vdd gnd cell_6t
Xbit_r0_c218 bl[218] br[218] wl[0] vdd gnd cell_6t
Xbit_r1_c218 bl[218] br[218] wl[1] vdd gnd cell_6t
Xbit_r2_c218 bl[218] br[218] wl[2] vdd gnd cell_6t
Xbit_r3_c218 bl[218] br[218] wl[3] vdd gnd cell_6t
Xbit_r4_c218 bl[218] br[218] wl[4] vdd gnd cell_6t
Xbit_r5_c218 bl[218] br[218] wl[5] vdd gnd cell_6t
Xbit_r6_c218 bl[218] br[218] wl[6] vdd gnd cell_6t
Xbit_r7_c218 bl[218] br[218] wl[7] vdd gnd cell_6t
Xbit_r8_c218 bl[218] br[218] wl[8] vdd gnd cell_6t
Xbit_r9_c218 bl[218] br[218] wl[9] vdd gnd cell_6t
Xbit_r10_c218 bl[218] br[218] wl[10] vdd gnd cell_6t
Xbit_r11_c218 bl[218] br[218] wl[11] vdd gnd cell_6t
Xbit_r12_c218 bl[218] br[218] wl[12] vdd gnd cell_6t
Xbit_r13_c218 bl[218] br[218] wl[13] vdd gnd cell_6t
Xbit_r14_c218 bl[218] br[218] wl[14] vdd gnd cell_6t
Xbit_r15_c218 bl[218] br[218] wl[15] vdd gnd cell_6t
Xbit_r16_c218 bl[218] br[218] wl[16] vdd gnd cell_6t
Xbit_r17_c218 bl[218] br[218] wl[17] vdd gnd cell_6t
Xbit_r18_c218 bl[218] br[218] wl[18] vdd gnd cell_6t
Xbit_r19_c218 bl[218] br[218] wl[19] vdd gnd cell_6t
Xbit_r20_c218 bl[218] br[218] wl[20] vdd gnd cell_6t
Xbit_r21_c218 bl[218] br[218] wl[21] vdd gnd cell_6t
Xbit_r22_c218 bl[218] br[218] wl[22] vdd gnd cell_6t
Xbit_r23_c218 bl[218] br[218] wl[23] vdd gnd cell_6t
Xbit_r24_c218 bl[218] br[218] wl[24] vdd gnd cell_6t
Xbit_r25_c218 bl[218] br[218] wl[25] vdd gnd cell_6t
Xbit_r26_c218 bl[218] br[218] wl[26] vdd gnd cell_6t
Xbit_r27_c218 bl[218] br[218] wl[27] vdd gnd cell_6t
Xbit_r28_c218 bl[218] br[218] wl[28] vdd gnd cell_6t
Xbit_r29_c218 bl[218] br[218] wl[29] vdd gnd cell_6t
Xbit_r30_c218 bl[218] br[218] wl[30] vdd gnd cell_6t
Xbit_r31_c218 bl[218] br[218] wl[31] vdd gnd cell_6t
Xbit_r32_c218 bl[218] br[218] wl[32] vdd gnd cell_6t
Xbit_r33_c218 bl[218] br[218] wl[33] vdd gnd cell_6t
Xbit_r34_c218 bl[218] br[218] wl[34] vdd gnd cell_6t
Xbit_r35_c218 bl[218] br[218] wl[35] vdd gnd cell_6t
Xbit_r36_c218 bl[218] br[218] wl[36] vdd gnd cell_6t
Xbit_r37_c218 bl[218] br[218] wl[37] vdd gnd cell_6t
Xbit_r38_c218 bl[218] br[218] wl[38] vdd gnd cell_6t
Xbit_r39_c218 bl[218] br[218] wl[39] vdd gnd cell_6t
Xbit_r40_c218 bl[218] br[218] wl[40] vdd gnd cell_6t
Xbit_r41_c218 bl[218] br[218] wl[41] vdd gnd cell_6t
Xbit_r42_c218 bl[218] br[218] wl[42] vdd gnd cell_6t
Xbit_r43_c218 bl[218] br[218] wl[43] vdd gnd cell_6t
Xbit_r44_c218 bl[218] br[218] wl[44] vdd gnd cell_6t
Xbit_r45_c218 bl[218] br[218] wl[45] vdd gnd cell_6t
Xbit_r46_c218 bl[218] br[218] wl[46] vdd gnd cell_6t
Xbit_r47_c218 bl[218] br[218] wl[47] vdd gnd cell_6t
Xbit_r48_c218 bl[218] br[218] wl[48] vdd gnd cell_6t
Xbit_r49_c218 bl[218] br[218] wl[49] vdd gnd cell_6t
Xbit_r50_c218 bl[218] br[218] wl[50] vdd gnd cell_6t
Xbit_r51_c218 bl[218] br[218] wl[51] vdd gnd cell_6t
Xbit_r52_c218 bl[218] br[218] wl[52] vdd gnd cell_6t
Xbit_r53_c218 bl[218] br[218] wl[53] vdd gnd cell_6t
Xbit_r54_c218 bl[218] br[218] wl[54] vdd gnd cell_6t
Xbit_r55_c218 bl[218] br[218] wl[55] vdd gnd cell_6t
Xbit_r56_c218 bl[218] br[218] wl[56] vdd gnd cell_6t
Xbit_r57_c218 bl[218] br[218] wl[57] vdd gnd cell_6t
Xbit_r58_c218 bl[218] br[218] wl[58] vdd gnd cell_6t
Xbit_r59_c218 bl[218] br[218] wl[59] vdd gnd cell_6t
Xbit_r60_c218 bl[218] br[218] wl[60] vdd gnd cell_6t
Xbit_r61_c218 bl[218] br[218] wl[61] vdd gnd cell_6t
Xbit_r62_c218 bl[218] br[218] wl[62] vdd gnd cell_6t
Xbit_r63_c218 bl[218] br[218] wl[63] vdd gnd cell_6t
Xbit_r64_c218 bl[218] br[218] wl[64] vdd gnd cell_6t
Xbit_r65_c218 bl[218] br[218] wl[65] vdd gnd cell_6t
Xbit_r66_c218 bl[218] br[218] wl[66] vdd gnd cell_6t
Xbit_r67_c218 bl[218] br[218] wl[67] vdd gnd cell_6t
Xbit_r68_c218 bl[218] br[218] wl[68] vdd gnd cell_6t
Xbit_r69_c218 bl[218] br[218] wl[69] vdd gnd cell_6t
Xbit_r70_c218 bl[218] br[218] wl[70] vdd gnd cell_6t
Xbit_r71_c218 bl[218] br[218] wl[71] vdd gnd cell_6t
Xbit_r72_c218 bl[218] br[218] wl[72] vdd gnd cell_6t
Xbit_r73_c218 bl[218] br[218] wl[73] vdd gnd cell_6t
Xbit_r74_c218 bl[218] br[218] wl[74] vdd gnd cell_6t
Xbit_r75_c218 bl[218] br[218] wl[75] vdd gnd cell_6t
Xbit_r76_c218 bl[218] br[218] wl[76] vdd gnd cell_6t
Xbit_r77_c218 bl[218] br[218] wl[77] vdd gnd cell_6t
Xbit_r78_c218 bl[218] br[218] wl[78] vdd gnd cell_6t
Xbit_r79_c218 bl[218] br[218] wl[79] vdd gnd cell_6t
Xbit_r80_c218 bl[218] br[218] wl[80] vdd gnd cell_6t
Xbit_r81_c218 bl[218] br[218] wl[81] vdd gnd cell_6t
Xbit_r82_c218 bl[218] br[218] wl[82] vdd gnd cell_6t
Xbit_r83_c218 bl[218] br[218] wl[83] vdd gnd cell_6t
Xbit_r84_c218 bl[218] br[218] wl[84] vdd gnd cell_6t
Xbit_r85_c218 bl[218] br[218] wl[85] vdd gnd cell_6t
Xbit_r86_c218 bl[218] br[218] wl[86] vdd gnd cell_6t
Xbit_r87_c218 bl[218] br[218] wl[87] vdd gnd cell_6t
Xbit_r88_c218 bl[218] br[218] wl[88] vdd gnd cell_6t
Xbit_r89_c218 bl[218] br[218] wl[89] vdd gnd cell_6t
Xbit_r90_c218 bl[218] br[218] wl[90] vdd gnd cell_6t
Xbit_r91_c218 bl[218] br[218] wl[91] vdd gnd cell_6t
Xbit_r92_c218 bl[218] br[218] wl[92] vdd gnd cell_6t
Xbit_r93_c218 bl[218] br[218] wl[93] vdd gnd cell_6t
Xbit_r94_c218 bl[218] br[218] wl[94] vdd gnd cell_6t
Xbit_r95_c218 bl[218] br[218] wl[95] vdd gnd cell_6t
Xbit_r96_c218 bl[218] br[218] wl[96] vdd gnd cell_6t
Xbit_r97_c218 bl[218] br[218] wl[97] vdd gnd cell_6t
Xbit_r98_c218 bl[218] br[218] wl[98] vdd gnd cell_6t
Xbit_r99_c218 bl[218] br[218] wl[99] vdd gnd cell_6t
Xbit_r100_c218 bl[218] br[218] wl[100] vdd gnd cell_6t
Xbit_r101_c218 bl[218] br[218] wl[101] vdd gnd cell_6t
Xbit_r102_c218 bl[218] br[218] wl[102] vdd gnd cell_6t
Xbit_r103_c218 bl[218] br[218] wl[103] vdd gnd cell_6t
Xbit_r104_c218 bl[218] br[218] wl[104] vdd gnd cell_6t
Xbit_r105_c218 bl[218] br[218] wl[105] vdd gnd cell_6t
Xbit_r106_c218 bl[218] br[218] wl[106] vdd gnd cell_6t
Xbit_r107_c218 bl[218] br[218] wl[107] vdd gnd cell_6t
Xbit_r108_c218 bl[218] br[218] wl[108] vdd gnd cell_6t
Xbit_r109_c218 bl[218] br[218] wl[109] vdd gnd cell_6t
Xbit_r110_c218 bl[218] br[218] wl[110] vdd gnd cell_6t
Xbit_r111_c218 bl[218] br[218] wl[111] vdd gnd cell_6t
Xbit_r112_c218 bl[218] br[218] wl[112] vdd gnd cell_6t
Xbit_r113_c218 bl[218] br[218] wl[113] vdd gnd cell_6t
Xbit_r114_c218 bl[218] br[218] wl[114] vdd gnd cell_6t
Xbit_r115_c218 bl[218] br[218] wl[115] vdd gnd cell_6t
Xbit_r116_c218 bl[218] br[218] wl[116] vdd gnd cell_6t
Xbit_r117_c218 bl[218] br[218] wl[117] vdd gnd cell_6t
Xbit_r118_c218 bl[218] br[218] wl[118] vdd gnd cell_6t
Xbit_r119_c218 bl[218] br[218] wl[119] vdd gnd cell_6t
Xbit_r120_c218 bl[218] br[218] wl[120] vdd gnd cell_6t
Xbit_r121_c218 bl[218] br[218] wl[121] vdd gnd cell_6t
Xbit_r122_c218 bl[218] br[218] wl[122] vdd gnd cell_6t
Xbit_r123_c218 bl[218] br[218] wl[123] vdd gnd cell_6t
Xbit_r124_c218 bl[218] br[218] wl[124] vdd gnd cell_6t
Xbit_r125_c218 bl[218] br[218] wl[125] vdd gnd cell_6t
Xbit_r126_c218 bl[218] br[218] wl[126] vdd gnd cell_6t
Xbit_r127_c218 bl[218] br[218] wl[127] vdd gnd cell_6t
Xbit_r0_c219 bl[219] br[219] wl[0] vdd gnd cell_6t
Xbit_r1_c219 bl[219] br[219] wl[1] vdd gnd cell_6t
Xbit_r2_c219 bl[219] br[219] wl[2] vdd gnd cell_6t
Xbit_r3_c219 bl[219] br[219] wl[3] vdd gnd cell_6t
Xbit_r4_c219 bl[219] br[219] wl[4] vdd gnd cell_6t
Xbit_r5_c219 bl[219] br[219] wl[5] vdd gnd cell_6t
Xbit_r6_c219 bl[219] br[219] wl[6] vdd gnd cell_6t
Xbit_r7_c219 bl[219] br[219] wl[7] vdd gnd cell_6t
Xbit_r8_c219 bl[219] br[219] wl[8] vdd gnd cell_6t
Xbit_r9_c219 bl[219] br[219] wl[9] vdd gnd cell_6t
Xbit_r10_c219 bl[219] br[219] wl[10] vdd gnd cell_6t
Xbit_r11_c219 bl[219] br[219] wl[11] vdd gnd cell_6t
Xbit_r12_c219 bl[219] br[219] wl[12] vdd gnd cell_6t
Xbit_r13_c219 bl[219] br[219] wl[13] vdd gnd cell_6t
Xbit_r14_c219 bl[219] br[219] wl[14] vdd gnd cell_6t
Xbit_r15_c219 bl[219] br[219] wl[15] vdd gnd cell_6t
Xbit_r16_c219 bl[219] br[219] wl[16] vdd gnd cell_6t
Xbit_r17_c219 bl[219] br[219] wl[17] vdd gnd cell_6t
Xbit_r18_c219 bl[219] br[219] wl[18] vdd gnd cell_6t
Xbit_r19_c219 bl[219] br[219] wl[19] vdd gnd cell_6t
Xbit_r20_c219 bl[219] br[219] wl[20] vdd gnd cell_6t
Xbit_r21_c219 bl[219] br[219] wl[21] vdd gnd cell_6t
Xbit_r22_c219 bl[219] br[219] wl[22] vdd gnd cell_6t
Xbit_r23_c219 bl[219] br[219] wl[23] vdd gnd cell_6t
Xbit_r24_c219 bl[219] br[219] wl[24] vdd gnd cell_6t
Xbit_r25_c219 bl[219] br[219] wl[25] vdd gnd cell_6t
Xbit_r26_c219 bl[219] br[219] wl[26] vdd gnd cell_6t
Xbit_r27_c219 bl[219] br[219] wl[27] vdd gnd cell_6t
Xbit_r28_c219 bl[219] br[219] wl[28] vdd gnd cell_6t
Xbit_r29_c219 bl[219] br[219] wl[29] vdd gnd cell_6t
Xbit_r30_c219 bl[219] br[219] wl[30] vdd gnd cell_6t
Xbit_r31_c219 bl[219] br[219] wl[31] vdd gnd cell_6t
Xbit_r32_c219 bl[219] br[219] wl[32] vdd gnd cell_6t
Xbit_r33_c219 bl[219] br[219] wl[33] vdd gnd cell_6t
Xbit_r34_c219 bl[219] br[219] wl[34] vdd gnd cell_6t
Xbit_r35_c219 bl[219] br[219] wl[35] vdd gnd cell_6t
Xbit_r36_c219 bl[219] br[219] wl[36] vdd gnd cell_6t
Xbit_r37_c219 bl[219] br[219] wl[37] vdd gnd cell_6t
Xbit_r38_c219 bl[219] br[219] wl[38] vdd gnd cell_6t
Xbit_r39_c219 bl[219] br[219] wl[39] vdd gnd cell_6t
Xbit_r40_c219 bl[219] br[219] wl[40] vdd gnd cell_6t
Xbit_r41_c219 bl[219] br[219] wl[41] vdd gnd cell_6t
Xbit_r42_c219 bl[219] br[219] wl[42] vdd gnd cell_6t
Xbit_r43_c219 bl[219] br[219] wl[43] vdd gnd cell_6t
Xbit_r44_c219 bl[219] br[219] wl[44] vdd gnd cell_6t
Xbit_r45_c219 bl[219] br[219] wl[45] vdd gnd cell_6t
Xbit_r46_c219 bl[219] br[219] wl[46] vdd gnd cell_6t
Xbit_r47_c219 bl[219] br[219] wl[47] vdd gnd cell_6t
Xbit_r48_c219 bl[219] br[219] wl[48] vdd gnd cell_6t
Xbit_r49_c219 bl[219] br[219] wl[49] vdd gnd cell_6t
Xbit_r50_c219 bl[219] br[219] wl[50] vdd gnd cell_6t
Xbit_r51_c219 bl[219] br[219] wl[51] vdd gnd cell_6t
Xbit_r52_c219 bl[219] br[219] wl[52] vdd gnd cell_6t
Xbit_r53_c219 bl[219] br[219] wl[53] vdd gnd cell_6t
Xbit_r54_c219 bl[219] br[219] wl[54] vdd gnd cell_6t
Xbit_r55_c219 bl[219] br[219] wl[55] vdd gnd cell_6t
Xbit_r56_c219 bl[219] br[219] wl[56] vdd gnd cell_6t
Xbit_r57_c219 bl[219] br[219] wl[57] vdd gnd cell_6t
Xbit_r58_c219 bl[219] br[219] wl[58] vdd gnd cell_6t
Xbit_r59_c219 bl[219] br[219] wl[59] vdd gnd cell_6t
Xbit_r60_c219 bl[219] br[219] wl[60] vdd gnd cell_6t
Xbit_r61_c219 bl[219] br[219] wl[61] vdd gnd cell_6t
Xbit_r62_c219 bl[219] br[219] wl[62] vdd gnd cell_6t
Xbit_r63_c219 bl[219] br[219] wl[63] vdd gnd cell_6t
Xbit_r64_c219 bl[219] br[219] wl[64] vdd gnd cell_6t
Xbit_r65_c219 bl[219] br[219] wl[65] vdd gnd cell_6t
Xbit_r66_c219 bl[219] br[219] wl[66] vdd gnd cell_6t
Xbit_r67_c219 bl[219] br[219] wl[67] vdd gnd cell_6t
Xbit_r68_c219 bl[219] br[219] wl[68] vdd gnd cell_6t
Xbit_r69_c219 bl[219] br[219] wl[69] vdd gnd cell_6t
Xbit_r70_c219 bl[219] br[219] wl[70] vdd gnd cell_6t
Xbit_r71_c219 bl[219] br[219] wl[71] vdd gnd cell_6t
Xbit_r72_c219 bl[219] br[219] wl[72] vdd gnd cell_6t
Xbit_r73_c219 bl[219] br[219] wl[73] vdd gnd cell_6t
Xbit_r74_c219 bl[219] br[219] wl[74] vdd gnd cell_6t
Xbit_r75_c219 bl[219] br[219] wl[75] vdd gnd cell_6t
Xbit_r76_c219 bl[219] br[219] wl[76] vdd gnd cell_6t
Xbit_r77_c219 bl[219] br[219] wl[77] vdd gnd cell_6t
Xbit_r78_c219 bl[219] br[219] wl[78] vdd gnd cell_6t
Xbit_r79_c219 bl[219] br[219] wl[79] vdd gnd cell_6t
Xbit_r80_c219 bl[219] br[219] wl[80] vdd gnd cell_6t
Xbit_r81_c219 bl[219] br[219] wl[81] vdd gnd cell_6t
Xbit_r82_c219 bl[219] br[219] wl[82] vdd gnd cell_6t
Xbit_r83_c219 bl[219] br[219] wl[83] vdd gnd cell_6t
Xbit_r84_c219 bl[219] br[219] wl[84] vdd gnd cell_6t
Xbit_r85_c219 bl[219] br[219] wl[85] vdd gnd cell_6t
Xbit_r86_c219 bl[219] br[219] wl[86] vdd gnd cell_6t
Xbit_r87_c219 bl[219] br[219] wl[87] vdd gnd cell_6t
Xbit_r88_c219 bl[219] br[219] wl[88] vdd gnd cell_6t
Xbit_r89_c219 bl[219] br[219] wl[89] vdd gnd cell_6t
Xbit_r90_c219 bl[219] br[219] wl[90] vdd gnd cell_6t
Xbit_r91_c219 bl[219] br[219] wl[91] vdd gnd cell_6t
Xbit_r92_c219 bl[219] br[219] wl[92] vdd gnd cell_6t
Xbit_r93_c219 bl[219] br[219] wl[93] vdd gnd cell_6t
Xbit_r94_c219 bl[219] br[219] wl[94] vdd gnd cell_6t
Xbit_r95_c219 bl[219] br[219] wl[95] vdd gnd cell_6t
Xbit_r96_c219 bl[219] br[219] wl[96] vdd gnd cell_6t
Xbit_r97_c219 bl[219] br[219] wl[97] vdd gnd cell_6t
Xbit_r98_c219 bl[219] br[219] wl[98] vdd gnd cell_6t
Xbit_r99_c219 bl[219] br[219] wl[99] vdd gnd cell_6t
Xbit_r100_c219 bl[219] br[219] wl[100] vdd gnd cell_6t
Xbit_r101_c219 bl[219] br[219] wl[101] vdd gnd cell_6t
Xbit_r102_c219 bl[219] br[219] wl[102] vdd gnd cell_6t
Xbit_r103_c219 bl[219] br[219] wl[103] vdd gnd cell_6t
Xbit_r104_c219 bl[219] br[219] wl[104] vdd gnd cell_6t
Xbit_r105_c219 bl[219] br[219] wl[105] vdd gnd cell_6t
Xbit_r106_c219 bl[219] br[219] wl[106] vdd gnd cell_6t
Xbit_r107_c219 bl[219] br[219] wl[107] vdd gnd cell_6t
Xbit_r108_c219 bl[219] br[219] wl[108] vdd gnd cell_6t
Xbit_r109_c219 bl[219] br[219] wl[109] vdd gnd cell_6t
Xbit_r110_c219 bl[219] br[219] wl[110] vdd gnd cell_6t
Xbit_r111_c219 bl[219] br[219] wl[111] vdd gnd cell_6t
Xbit_r112_c219 bl[219] br[219] wl[112] vdd gnd cell_6t
Xbit_r113_c219 bl[219] br[219] wl[113] vdd gnd cell_6t
Xbit_r114_c219 bl[219] br[219] wl[114] vdd gnd cell_6t
Xbit_r115_c219 bl[219] br[219] wl[115] vdd gnd cell_6t
Xbit_r116_c219 bl[219] br[219] wl[116] vdd gnd cell_6t
Xbit_r117_c219 bl[219] br[219] wl[117] vdd gnd cell_6t
Xbit_r118_c219 bl[219] br[219] wl[118] vdd gnd cell_6t
Xbit_r119_c219 bl[219] br[219] wl[119] vdd gnd cell_6t
Xbit_r120_c219 bl[219] br[219] wl[120] vdd gnd cell_6t
Xbit_r121_c219 bl[219] br[219] wl[121] vdd gnd cell_6t
Xbit_r122_c219 bl[219] br[219] wl[122] vdd gnd cell_6t
Xbit_r123_c219 bl[219] br[219] wl[123] vdd gnd cell_6t
Xbit_r124_c219 bl[219] br[219] wl[124] vdd gnd cell_6t
Xbit_r125_c219 bl[219] br[219] wl[125] vdd gnd cell_6t
Xbit_r126_c219 bl[219] br[219] wl[126] vdd gnd cell_6t
Xbit_r127_c219 bl[219] br[219] wl[127] vdd gnd cell_6t
Xbit_r0_c220 bl[220] br[220] wl[0] vdd gnd cell_6t
Xbit_r1_c220 bl[220] br[220] wl[1] vdd gnd cell_6t
Xbit_r2_c220 bl[220] br[220] wl[2] vdd gnd cell_6t
Xbit_r3_c220 bl[220] br[220] wl[3] vdd gnd cell_6t
Xbit_r4_c220 bl[220] br[220] wl[4] vdd gnd cell_6t
Xbit_r5_c220 bl[220] br[220] wl[5] vdd gnd cell_6t
Xbit_r6_c220 bl[220] br[220] wl[6] vdd gnd cell_6t
Xbit_r7_c220 bl[220] br[220] wl[7] vdd gnd cell_6t
Xbit_r8_c220 bl[220] br[220] wl[8] vdd gnd cell_6t
Xbit_r9_c220 bl[220] br[220] wl[9] vdd gnd cell_6t
Xbit_r10_c220 bl[220] br[220] wl[10] vdd gnd cell_6t
Xbit_r11_c220 bl[220] br[220] wl[11] vdd gnd cell_6t
Xbit_r12_c220 bl[220] br[220] wl[12] vdd gnd cell_6t
Xbit_r13_c220 bl[220] br[220] wl[13] vdd gnd cell_6t
Xbit_r14_c220 bl[220] br[220] wl[14] vdd gnd cell_6t
Xbit_r15_c220 bl[220] br[220] wl[15] vdd gnd cell_6t
Xbit_r16_c220 bl[220] br[220] wl[16] vdd gnd cell_6t
Xbit_r17_c220 bl[220] br[220] wl[17] vdd gnd cell_6t
Xbit_r18_c220 bl[220] br[220] wl[18] vdd gnd cell_6t
Xbit_r19_c220 bl[220] br[220] wl[19] vdd gnd cell_6t
Xbit_r20_c220 bl[220] br[220] wl[20] vdd gnd cell_6t
Xbit_r21_c220 bl[220] br[220] wl[21] vdd gnd cell_6t
Xbit_r22_c220 bl[220] br[220] wl[22] vdd gnd cell_6t
Xbit_r23_c220 bl[220] br[220] wl[23] vdd gnd cell_6t
Xbit_r24_c220 bl[220] br[220] wl[24] vdd gnd cell_6t
Xbit_r25_c220 bl[220] br[220] wl[25] vdd gnd cell_6t
Xbit_r26_c220 bl[220] br[220] wl[26] vdd gnd cell_6t
Xbit_r27_c220 bl[220] br[220] wl[27] vdd gnd cell_6t
Xbit_r28_c220 bl[220] br[220] wl[28] vdd gnd cell_6t
Xbit_r29_c220 bl[220] br[220] wl[29] vdd gnd cell_6t
Xbit_r30_c220 bl[220] br[220] wl[30] vdd gnd cell_6t
Xbit_r31_c220 bl[220] br[220] wl[31] vdd gnd cell_6t
Xbit_r32_c220 bl[220] br[220] wl[32] vdd gnd cell_6t
Xbit_r33_c220 bl[220] br[220] wl[33] vdd gnd cell_6t
Xbit_r34_c220 bl[220] br[220] wl[34] vdd gnd cell_6t
Xbit_r35_c220 bl[220] br[220] wl[35] vdd gnd cell_6t
Xbit_r36_c220 bl[220] br[220] wl[36] vdd gnd cell_6t
Xbit_r37_c220 bl[220] br[220] wl[37] vdd gnd cell_6t
Xbit_r38_c220 bl[220] br[220] wl[38] vdd gnd cell_6t
Xbit_r39_c220 bl[220] br[220] wl[39] vdd gnd cell_6t
Xbit_r40_c220 bl[220] br[220] wl[40] vdd gnd cell_6t
Xbit_r41_c220 bl[220] br[220] wl[41] vdd gnd cell_6t
Xbit_r42_c220 bl[220] br[220] wl[42] vdd gnd cell_6t
Xbit_r43_c220 bl[220] br[220] wl[43] vdd gnd cell_6t
Xbit_r44_c220 bl[220] br[220] wl[44] vdd gnd cell_6t
Xbit_r45_c220 bl[220] br[220] wl[45] vdd gnd cell_6t
Xbit_r46_c220 bl[220] br[220] wl[46] vdd gnd cell_6t
Xbit_r47_c220 bl[220] br[220] wl[47] vdd gnd cell_6t
Xbit_r48_c220 bl[220] br[220] wl[48] vdd gnd cell_6t
Xbit_r49_c220 bl[220] br[220] wl[49] vdd gnd cell_6t
Xbit_r50_c220 bl[220] br[220] wl[50] vdd gnd cell_6t
Xbit_r51_c220 bl[220] br[220] wl[51] vdd gnd cell_6t
Xbit_r52_c220 bl[220] br[220] wl[52] vdd gnd cell_6t
Xbit_r53_c220 bl[220] br[220] wl[53] vdd gnd cell_6t
Xbit_r54_c220 bl[220] br[220] wl[54] vdd gnd cell_6t
Xbit_r55_c220 bl[220] br[220] wl[55] vdd gnd cell_6t
Xbit_r56_c220 bl[220] br[220] wl[56] vdd gnd cell_6t
Xbit_r57_c220 bl[220] br[220] wl[57] vdd gnd cell_6t
Xbit_r58_c220 bl[220] br[220] wl[58] vdd gnd cell_6t
Xbit_r59_c220 bl[220] br[220] wl[59] vdd gnd cell_6t
Xbit_r60_c220 bl[220] br[220] wl[60] vdd gnd cell_6t
Xbit_r61_c220 bl[220] br[220] wl[61] vdd gnd cell_6t
Xbit_r62_c220 bl[220] br[220] wl[62] vdd gnd cell_6t
Xbit_r63_c220 bl[220] br[220] wl[63] vdd gnd cell_6t
Xbit_r64_c220 bl[220] br[220] wl[64] vdd gnd cell_6t
Xbit_r65_c220 bl[220] br[220] wl[65] vdd gnd cell_6t
Xbit_r66_c220 bl[220] br[220] wl[66] vdd gnd cell_6t
Xbit_r67_c220 bl[220] br[220] wl[67] vdd gnd cell_6t
Xbit_r68_c220 bl[220] br[220] wl[68] vdd gnd cell_6t
Xbit_r69_c220 bl[220] br[220] wl[69] vdd gnd cell_6t
Xbit_r70_c220 bl[220] br[220] wl[70] vdd gnd cell_6t
Xbit_r71_c220 bl[220] br[220] wl[71] vdd gnd cell_6t
Xbit_r72_c220 bl[220] br[220] wl[72] vdd gnd cell_6t
Xbit_r73_c220 bl[220] br[220] wl[73] vdd gnd cell_6t
Xbit_r74_c220 bl[220] br[220] wl[74] vdd gnd cell_6t
Xbit_r75_c220 bl[220] br[220] wl[75] vdd gnd cell_6t
Xbit_r76_c220 bl[220] br[220] wl[76] vdd gnd cell_6t
Xbit_r77_c220 bl[220] br[220] wl[77] vdd gnd cell_6t
Xbit_r78_c220 bl[220] br[220] wl[78] vdd gnd cell_6t
Xbit_r79_c220 bl[220] br[220] wl[79] vdd gnd cell_6t
Xbit_r80_c220 bl[220] br[220] wl[80] vdd gnd cell_6t
Xbit_r81_c220 bl[220] br[220] wl[81] vdd gnd cell_6t
Xbit_r82_c220 bl[220] br[220] wl[82] vdd gnd cell_6t
Xbit_r83_c220 bl[220] br[220] wl[83] vdd gnd cell_6t
Xbit_r84_c220 bl[220] br[220] wl[84] vdd gnd cell_6t
Xbit_r85_c220 bl[220] br[220] wl[85] vdd gnd cell_6t
Xbit_r86_c220 bl[220] br[220] wl[86] vdd gnd cell_6t
Xbit_r87_c220 bl[220] br[220] wl[87] vdd gnd cell_6t
Xbit_r88_c220 bl[220] br[220] wl[88] vdd gnd cell_6t
Xbit_r89_c220 bl[220] br[220] wl[89] vdd gnd cell_6t
Xbit_r90_c220 bl[220] br[220] wl[90] vdd gnd cell_6t
Xbit_r91_c220 bl[220] br[220] wl[91] vdd gnd cell_6t
Xbit_r92_c220 bl[220] br[220] wl[92] vdd gnd cell_6t
Xbit_r93_c220 bl[220] br[220] wl[93] vdd gnd cell_6t
Xbit_r94_c220 bl[220] br[220] wl[94] vdd gnd cell_6t
Xbit_r95_c220 bl[220] br[220] wl[95] vdd gnd cell_6t
Xbit_r96_c220 bl[220] br[220] wl[96] vdd gnd cell_6t
Xbit_r97_c220 bl[220] br[220] wl[97] vdd gnd cell_6t
Xbit_r98_c220 bl[220] br[220] wl[98] vdd gnd cell_6t
Xbit_r99_c220 bl[220] br[220] wl[99] vdd gnd cell_6t
Xbit_r100_c220 bl[220] br[220] wl[100] vdd gnd cell_6t
Xbit_r101_c220 bl[220] br[220] wl[101] vdd gnd cell_6t
Xbit_r102_c220 bl[220] br[220] wl[102] vdd gnd cell_6t
Xbit_r103_c220 bl[220] br[220] wl[103] vdd gnd cell_6t
Xbit_r104_c220 bl[220] br[220] wl[104] vdd gnd cell_6t
Xbit_r105_c220 bl[220] br[220] wl[105] vdd gnd cell_6t
Xbit_r106_c220 bl[220] br[220] wl[106] vdd gnd cell_6t
Xbit_r107_c220 bl[220] br[220] wl[107] vdd gnd cell_6t
Xbit_r108_c220 bl[220] br[220] wl[108] vdd gnd cell_6t
Xbit_r109_c220 bl[220] br[220] wl[109] vdd gnd cell_6t
Xbit_r110_c220 bl[220] br[220] wl[110] vdd gnd cell_6t
Xbit_r111_c220 bl[220] br[220] wl[111] vdd gnd cell_6t
Xbit_r112_c220 bl[220] br[220] wl[112] vdd gnd cell_6t
Xbit_r113_c220 bl[220] br[220] wl[113] vdd gnd cell_6t
Xbit_r114_c220 bl[220] br[220] wl[114] vdd gnd cell_6t
Xbit_r115_c220 bl[220] br[220] wl[115] vdd gnd cell_6t
Xbit_r116_c220 bl[220] br[220] wl[116] vdd gnd cell_6t
Xbit_r117_c220 bl[220] br[220] wl[117] vdd gnd cell_6t
Xbit_r118_c220 bl[220] br[220] wl[118] vdd gnd cell_6t
Xbit_r119_c220 bl[220] br[220] wl[119] vdd gnd cell_6t
Xbit_r120_c220 bl[220] br[220] wl[120] vdd gnd cell_6t
Xbit_r121_c220 bl[220] br[220] wl[121] vdd gnd cell_6t
Xbit_r122_c220 bl[220] br[220] wl[122] vdd gnd cell_6t
Xbit_r123_c220 bl[220] br[220] wl[123] vdd gnd cell_6t
Xbit_r124_c220 bl[220] br[220] wl[124] vdd gnd cell_6t
Xbit_r125_c220 bl[220] br[220] wl[125] vdd gnd cell_6t
Xbit_r126_c220 bl[220] br[220] wl[126] vdd gnd cell_6t
Xbit_r127_c220 bl[220] br[220] wl[127] vdd gnd cell_6t
Xbit_r0_c221 bl[221] br[221] wl[0] vdd gnd cell_6t
Xbit_r1_c221 bl[221] br[221] wl[1] vdd gnd cell_6t
Xbit_r2_c221 bl[221] br[221] wl[2] vdd gnd cell_6t
Xbit_r3_c221 bl[221] br[221] wl[3] vdd gnd cell_6t
Xbit_r4_c221 bl[221] br[221] wl[4] vdd gnd cell_6t
Xbit_r5_c221 bl[221] br[221] wl[5] vdd gnd cell_6t
Xbit_r6_c221 bl[221] br[221] wl[6] vdd gnd cell_6t
Xbit_r7_c221 bl[221] br[221] wl[7] vdd gnd cell_6t
Xbit_r8_c221 bl[221] br[221] wl[8] vdd gnd cell_6t
Xbit_r9_c221 bl[221] br[221] wl[9] vdd gnd cell_6t
Xbit_r10_c221 bl[221] br[221] wl[10] vdd gnd cell_6t
Xbit_r11_c221 bl[221] br[221] wl[11] vdd gnd cell_6t
Xbit_r12_c221 bl[221] br[221] wl[12] vdd gnd cell_6t
Xbit_r13_c221 bl[221] br[221] wl[13] vdd gnd cell_6t
Xbit_r14_c221 bl[221] br[221] wl[14] vdd gnd cell_6t
Xbit_r15_c221 bl[221] br[221] wl[15] vdd gnd cell_6t
Xbit_r16_c221 bl[221] br[221] wl[16] vdd gnd cell_6t
Xbit_r17_c221 bl[221] br[221] wl[17] vdd gnd cell_6t
Xbit_r18_c221 bl[221] br[221] wl[18] vdd gnd cell_6t
Xbit_r19_c221 bl[221] br[221] wl[19] vdd gnd cell_6t
Xbit_r20_c221 bl[221] br[221] wl[20] vdd gnd cell_6t
Xbit_r21_c221 bl[221] br[221] wl[21] vdd gnd cell_6t
Xbit_r22_c221 bl[221] br[221] wl[22] vdd gnd cell_6t
Xbit_r23_c221 bl[221] br[221] wl[23] vdd gnd cell_6t
Xbit_r24_c221 bl[221] br[221] wl[24] vdd gnd cell_6t
Xbit_r25_c221 bl[221] br[221] wl[25] vdd gnd cell_6t
Xbit_r26_c221 bl[221] br[221] wl[26] vdd gnd cell_6t
Xbit_r27_c221 bl[221] br[221] wl[27] vdd gnd cell_6t
Xbit_r28_c221 bl[221] br[221] wl[28] vdd gnd cell_6t
Xbit_r29_c221 bl[221] br[221] wl[29] vdd gnd cell_6t
Xbit_r30_c221 bl[221] br[221] wl[30] vdd gnd cell_6t
Xbit_r31_c221 bl[221] br[221] wl[31] vdd gnd cell_6t
Xbit_r32_c221 bl[221] br[221] wl[32] vdd gnd cell_6t
Xbit_r33_c221 bl[221] br[221] wl[33] vdd gnd cell_6t
Xbit_r34_c221 bl[221] br[221] wl[34] vdd gnd cell_6t
Xbit_r35_c221 bl[221] br[221] wl[35] vdd gnd cell_6t
Xbit_r36_c221 bl[221] br[221] wl[36] vdd gnd cell_6t
Xbit_r37_c221 bl[221] br[221] wl[37] vdd gnd cell_6t
Xbit_r38_c221 bl[221] br[221] wl[38] vdd gnd cell_6t
Xbit_r39_c221 bl[221] br[221] wl[39] vdd gnd cell_6t
Xbit_r40_c221 bl[221] br[221] wl[40] vdd gnd cell_6t
Xbit_r41_c221 bl[221] br[221] wl[41] vdd gnd cell_6t
Xbit_r42_c221 bl[221] br[221] wl[42] vdd gnd cell_6t
Xbit_r43_c221 bl[221] br[221] wl[43] vdd gnd cell_6t
Xbit_r44_c221 bl[221] br[221] wl[44] vdd gnd cell_6t
Xbit_r45_c221 bl[221] br[221] wl[45] vdd gnd cell_6t
Xbit_r46_c221 bl[221] br[221] wl[46] vdd gnd cell_6t
Xbit_r47_c221 bl[221] br[221] wl[47] vdd gnd cell_6t
Xbit_r48_c221 bl[221] br[221] wl[48] vdd gnd cell_6t
Xbit_r49_c221 bl[221] br[221] wl[49] vdd gnd cell_6t
Xbit_r50_c221 bl[221] br[221] wl[50] vdd gnd cell_6t
Xbit_r51_c221 bl[221] br[221] wl[51] vdd gnd cell_6t
Xbit_r52_c221 bl[221] br[221] wl[52] vdd gnd cell_6t
Xbit_r53_c221 bl[221] br[221] wl[53] vdd gnd cell_6t
Xbit_r54_c221 bl[221] br[221] wl[54] vdd gnd cell_6t
Xbit_r55_c221 bl[221] br[221] wl[55] vdd gnd cell_6t
Xbit_r56_c221 bl[221] br[221] wl[56] vdd gnd cell_6t
Xbit_r57_c221 bl[221] br[221] wl[57] vdd gnd cell_6t
Xbit_r58_c221 bl[221] br[221] wl[58] vdd gnd cell_6t
Xbit_r59_c221 bl[221] br[221] wl[59] vdd gnd cell_6t
Xbit_r60_c221 bl[221] br[221] wl[60] vdd gnd cell_6t
Xbit_r61_c221 bl[221] br[221] wl[61] vdd gnd cell_6t
Xbit_r62_c221 bl[221] br[221] wl[62] vdd gnd cell_6t
Xbit_r63_c221 bl[221] br[221] wl[63] vdd gnd cell_6t
Xbit_r64_c221 bl[221] br[221] wl[64] vdd gnd cell_6t
Xbit_r65_c221 bl[221] br[221] wl[65] vdd gnd cell_6t
Xbit_r66_c221 bl[221] br[221] wl[66] vdd gnd cell_6t
Xbit_r67_c221 bl[221] br[221] wl[67] vdd gnd cell_6t
Xbit_r68_c221 bl[221] br[221] wl[68] vdd gnd cell_6t
Xbit_r69_c221 bl[221] br[221] wl[69] vdd gnd cell_6t
Xbit_r70_c221 bl[221] br[221] wl[70] vdd gnd cell_6t
Xbit_r71_c221 bl[221] br[221] wl[71] vdd gnd cell_6t
Xbit_r72_c221 bl[221] br[221] wl[72] vdd gnd cell_6t
Xbit_r73_c221 bl[221] br[221] wl[73] vdd gnd cell_6t
Xbit_r74_c221 bl[221] br[221] wl[74] vdd gnd cell_6t
Xbit_r75_c221 bl[221] br[221] wl[75] vdd gnd cell_6t
Xbit_r76_c221 bl[221] br[221] wl[76] vdd gnd cell_6t
Xbit_r77_c221 bl[221] br[221] wl[77] vdd gnd cell_6t
Xbit_r78_c221 bl[221] br[221] wl[78] vdd gnd cell_6t
Xbit_r79_c221 bl[221] br[221] wl[79] vdd gnd cell_6t
Xbit_r80_c221 bl[221] br[221] wl[80] vdd gnd cell_6t
Xbit_r81_c221 bl[221] br[221] wl[81] vdd gnd cell_6t
Xbit_r82_c221 bl[221] br[221] wl[82] vdd gnd cell_6t
Xbit_r83_c221 bl[221] br[221] wl[83] vdd gnd cell_6t
Xbit_r84_c221 bl[221] br[221] wl[84] vdd gnd cell_6t
Xbit_r85_c221 bl[221] br[221] wl[85] vdd gnd cell_6t
Xbit_r86_c221 bl[221] br[221] wl[86] vdd gnd cell_6t
Xbit_r87_c221 bl[221] br[221] wl[87] vdd gnd cell_6t
Xbit_r88_c221 bl[221] br[221] wl[88] vdd gnd cell_6t
Xbit_r89_c221 bl[221] br[221] wl[89] vdd gnd cell_6t
Xbit_r90_c221 bl[221] br[221] wl[90] vdd gnd cell_6t
Xbit_r91_c221 bl[221] br[221] wl[91] vdd gnd cell_6t
Xbit_r92_c221 bl[221] br[221] wl[92] vdd gnd cell_6t
Xbit_r93_c221 bl[221] br[221] wl[93] vdd gnd cell_6t
Xbit_r94_c221 bl[221] br[221] wl[94] vdd gnd cell_6t
Xbit_r95_c221 bl[221] br[221] wl[95] vdd gnd cell_6t
Xbit_r96_c221 bl[221] br[221] wl[96] vdd gnd cell_6t
Xbit_r97_c221 bl[221] br[221] wl[97] vdd gnd cell_6t
Xbit_r98_c221 bl[221] br[221] wl[98] vdd gnd cell_6t
Xbit_r99_c221 bl[221] br[221] wl[99] vdd gnd cell_6t
Xbit_r100_c221 bl[221] br[221] wl[100] vdd gnd cell_6t
Xbit_r101_c221 bl[221] br[221] wl[101] vdd gnd cell_6t
Xbit_r102_c221 bl[221] br[221] wl[102] vdd gnd cell_6t
Xbit_r103_c221 bl[221] br[221] wl[103] vdd gnd cell_6t
Xbit_r104_c221 bl[221] br[221] wl[104] vdd gnd cell_6t
Xbit_r105_c221 bl[221] br[221] wl[105] vdd gnd cell_6t
Xbit_r106_c221 bl[221] br[221] wl[106] vdd gnd cell_6t
Xbit_r107_c221 bl[221] br[221] wl[107] vdd gnd cell_6t
Xbit_r108_c221 bl[221] br[221] wl[108] vdd gnd cell_6t
Xbit_r109_c221 bl[221] br[221] wl[109] vdd gnd cell_6t
Xbit_r110_c221 bl[221] br[221] wl[110] vdd gnd cell_6t
Xbit_r111_c221 bl[221] br[221] wl[111] vdd gnd cell_6t
Xbit_r112_c221 bl[221] br[221] wl[112] vdd gnd cell_6t
Xbit_r113_c221 bl[221] br[221] wl[113] vdd gnd cell_6t
Xbit_r114_c221 bl[221] br[221] wl[114] vdd gnd cell_6t
Xbit_r115_c221 bl[221] br[221] wl[115] vdd gnd cell_6t
Xbit_r116_c221 bl[221] br[221] wl[116] vdd gnd cell_6t
Xbit_r117_c221 bl[221] br[221] wl[117] vdd gnd cell_6t
Xbit_r118_c221 bl[221] br[221] wl[118] vdd gnd cell_6t
Xbit_r119_c221 bl[221] br[221] wl[119] vdd gnd cell_6t
Xbit_r120_c221 bl[221] br[221] wl[120] vdd gnd cell_6t
Xbit_r121_c221 bl[221] br[221] wl[121] vdd gnd cell_6t
Xbit_r122_c221 bl[221] br[221] wl[122] vdd gnd cell_6t
Xbit_r123_c221 bl[221] br[221] wl[123] vdd gnd cell_6t
Xbit_r124_c221 bl[221] br[221] wl[124] vdd gnd cell_6t
Xbit_r125_c221 bl[221] br[221] wl[125] vdd gnd cell_6t
Xbit_r126_c221 bl[221] br[221] wl[126] vdd gnd cell_6t
Xbit_r127_c221 bl[221] br[221] wl[127] vdd gnd cell_6t
Xbit_r0_c222 bl[222] br[222] wl[0] vdd gnd cell_6t
Xbit_r1_c222 bl[222] br[222] wl[1] vdd gnd cell_6t
Xbit_r2_c222 bl[222] br[222] wl[2] vdd gnd cell_6t
Xbit_r3_c222 bl[222] br[222] wl[3] vdd gnd cell_6t
Xbit_r4_c222 bl[222] br[222] wl[4] vdd gnd cell_6t
Xbit_r5_c222 bl[222] br[222] wl[5] vdd gnd cell_6t
Xbit_r6_c222 bl[222] br[222] wl[6] vdd gnd cell_6t
Xbit_r7_c222 bl[222] br[222] wl[7] vdd gnd cell_6t
Xbit_r8_c222 bl[222] br[222] wl[8] vdd gnd cell_6t
Xbit_r9_c222 bl[222] br[222] wl[9] vdd gnd cell_6t
Xbit_r10_c222 bl[222] br[222] wl[10] vdd gnd cell_6t
Xbit_r11_c222 bl[222] br[222] wl[11] vdd gnd cell_6t
Xbit_r12_c222 bl[222] br[222] wl[12] vdd gnd cell_6t
Xbit_r13_c222 bl[222] br[222] wl[13] vdd gnd cell_6t
Xbit_r14_c222 bl[222] br[222] wl[14] vdd gnd cell_6t
Xbit_r15_c222 bl[222] br[222] wl[15] vdd gnd cell_6t
Xbit_r16_c222 bl[222] br[222] wl[16] vdd gnd cell_6t
Xbit_r17_c222 bl[222] br[222] wl[17] vdd gnd cell_6t
Xbit_r18_c222 bl[222] br[222] wl[18] vdd gnd cell_6t
Xbit_r19_c222 bl[222] br[222] wl[19] vdd gnd cell_6t
Xbit_r20_c222 bl[222] br[222] wl[20] vdd gnd cell_6t
Xbit_r21_c222 bl[222] br[222] wl[21] vdd gnd cell_6t
Xbit_r22_c222 bl[222] br[222] wl[22] vdd gnd cell_6t
Xbit_r23_c222 bl[222] br[222] wl[23] vdd gnd cell_6t
Xbit_r24_c222 bl[222] br[222] wl[24] vdd gnd cell_6t
Xbit_r25_c222 bl[222] br[222] wl[25] vdd gnd cell_6t
Xbit_r26_c222 bl[222] br[222] wl[26] vdd gnd cell_6t
Xbit_r27_c222 bl[222] br[222] wl[27] vdd gnd cell_6t
Xbit_r28_c222 bl[222] br[222] wl[28] vdd gnd cell_6t
Xbit_r29_c222 bl[222] br[222] wl[29] vdd gnd cell_6t
Xbit_r30_c222 bl[222] br[222] wl[30] vdd gnd cell_6t
Xbit_r31_c222 bl[222] br[222] wl[31] vdd gnd cell_6t
Xbit_r32_c222 bl[222] br[222] wl[32] vdd gnd cell_6t
Xbit_r33_c222 bl[222] br[222] wl[33] vdd gnd cell_6t
Xbit_r34_c222 bl[222] br[222] wl[34] vdd gnd cell_6t
Xbit_r35_c222 bl[222] br[222] wl[35] vdd gnd cell_6t
Xbit_r36_c222 bl[222] br[222] wl[36] vdd gnd cell_6t
Xbit_r37_c222 bl[222] br[222] wl[37] vdd gnd cell_6t
Xbit_r38_c222 bl[222] br[222] wl[38] vdd gnd cell_6t
Xbit_r39_c222 bl[222] br[222] wl[39] vdd gnd cell_6t
Xbit_r40_c222 bl[222] br[222] wl[40] vdd gnd cell_6t
Xbit_r41_c222 bl[222] br[222] wl[41] vdd gnd cell_6t
Xbit_r42_c222 bl[222] br[222] wl[42] vdd gnd cell_6t
Xbit_r43_c222 bl[222] br[222] wl[43] vdd gnd cell_6t
Xbit_r44_c222 bl[222] br[222] wl[44] vdd gnd cell_6t
Xbit_r45_c222 bl[222] br[222] wl[45] vdd gnd cell_6t
Xbit_r46_c222 bl[222] br[222] wl[46] vdd gnd cell_6t
Xbit_r47_c222 bl[222] br[222] wl[47] vdd gnd cell_6t
Xbit_r48_c222 bl[222] br[222] wl[48] vdd gnd cell_6t
Xbit_r49_c222 bl[222] br[222] wl[49] vdd gnd cell_6t
Xbit_r50_c222 bl[222] br[222] wl[50] vdd gnd cell_6t
Xbit_r51_c222 bl[222] br[222] wl[51] vdd gnd cell_6t
Xbit_r52_c222 bl[222] br[222] wl[52] vdd gnd cell_6t
Xbit_r53_c222 bl[222] br[222] wl[53] vdd gnd cell_6t
Xbit_r54_c222 bl[222] br[222] wl[54] vdd gnd cell_6t
Xbit_r55_c222 bl[222] br[222] wl[55] vdd gnd cell_6t
Xbit_r56_c222 bl[222] br[222] wl[56] vdd gnd cell_6t
Xbit_r57_c222 bl[222] br[222] wl[57] vdd gnd cell_6t
Xbit_r58_c222 bl[222] br[222] wl[58] vdd gnd cell_6t
Xbit_r59_c222 bl[222] br[222] wl[59] vdd gnd cell_6t
Xbit_r60_c222 bl[222] br[222] wl[60] vdd gnd cell_6t
Xbit_r61_c222 bl[222] br[222] wl[61] vdd gnd cell_6t
Xbit_r62_c222 bl[222] br[222] wl[62] vdd gnd cell_6t
Xbit_r63_c222 bl[222] br[222] wl[63] vdd gnd cell_6t
Xbit_r64_c222 bl[222] br[222] wl[64] vdd gnd cell_6t
Xbit_r65_c222 bl[222] br[222] wl[65] vdd gnd cell_6t
Xbit_r66_c222 bl[222] br[222] wl[66] vdd gnd cell_6t
Xbit_r67_c222 bl[222] br[222] wl[67] vdd gnd cell_6t
Xbit_r68_c222 bl[222] br[222] wl[68] vdd gnd cell_6t
Xbit_r69_c222 bl[222] br[222] wl[69] vdd gnd cell_6t
Xbit_r70_c222 bl[222] br[222] wl[70] vdd gnd cell_6t
Xbit_r71_c222 bl[222] br[222] wl[71] vdd gnd cell_6t
Xbit_r72_c222 bl[222] br[222] wl[72] vdd gnd cell_6t
Xbit_r73_c222 bl[222] br[222] wl[73] vdd gnd cell_6t
Xbit_r74_c222 bl[222] br[222] wl[74] vdd gnd cell_6t
Xbit_r75_c222 bl[222] br[222] wl[75] vdd gnd cell_6t
Xbit_r76_c222 bl[222] br[222] wl[76] vdd gnd cell_6t
Xbit_r77_c222 bl[222] br[222] wl[77] vdd gnd cell_6t
Xbit_r78_c222 bl[222] br[222] wl[78] vdd gnd cell_6t
Xbit_r79_c222 bl[222] br[222] wl[79] vdd gnd cell_6t
Xbit_r80_c222 bl[222] br[222] wl[80] vdd gnd cell_6t
Xbit_r81_c222 bl[222] br[222] wl[81] vdd gnd cell_6t
Xbit_r82_c222 bl[222] br[222] wl[82] vdd gnd cell_6t
Xbit_r83_c222 bl[222] br[222] wl[83] vdd gnd cell_6t
Xbit_r84_c222 bl[222] br[222] wl[84] vdd gnd cell_6t
Xbit_r85_c222 bl[222] br[222] wl[85] vdd gnd cell_6t
Xbit_r86_c222 bl[222] br[222] wl[86] vdd gnd cell_6t
Xbit_r87_c222 bl[222] br[222] wl[87] vdd gnd cell_6t
Xbit_r88_c222 bl[222] br[222] wl[88] vdd gnd cell_6t
Xbit_r89_c222 bl[222] br[222] wl[89] vdd gnd cell_6t
Xbit_r90_c222 bl[222] br[222] wl[90] vdd gnd cell_6t
Xbit_r91_c222 bl[222] br[222] wl[91] vdd gnd cell_6t
Xbit_r92_c222 bl[222] br[222] wl[92] vdd gnd cell_6t
Xbit_r93_c222 bl[222] br[222] wl[93] vdd gnd cell_6t
Xbit_r94_c222 bl[222] br[222] wl[94] vdd gnd cell_6t
Xbit_r95_c222 bl[222] br[222] wl[95] vdd gnd cell_6t
Xbit_r96_c222 bl[222] br[222] wl[96] vdd gnd cell_6t
Xbit_r97_c222 bl[222] br[222] wl[97] vdd gnd cell_6t
Xbit_r98_c222 bl[222] br[222] wl[98] vdd gnd cell_6t
Xbit_r99_c222 bl[222] br[222] wl[99] vdd gnd cell_6t
Xbit_r100_c222 bl[222] br[222] wl[100] vdd gnd cell_6t
Xbit_r101_c222 bl[222] br[222] wl[101] vdd gnd cell_6t
Xbit_r102_c222 bl[222] br[222] wl[102] vdd gnd cell_6t
Xbit_r103_c222 bl[222] br[222] wl[103] vdd gnd cell_6t
Xbit_r104_c222 bl[222] br[222] wl[104] vdd gnd cell_6t
Xbit_r105_c222 bl[222] br[222] wl[105] vdd gnd cell_6t
Xbit_r106_c222 bl[222] br[222] wl[106] vdd gnd cell_6t
Xbit_r107_c222 bl[222] br[222] wl[107] vdd gnd cell_6t
Xbit_r108_c222 bl[222] br[222] wl[108] vdd gnd cell_6t
Xbit_r109_c222 bl[222] br[222] wl[109] vdd gnd cell_6t
Xbit_r110_c222 bl[222] br[222] wl[110] vdd gnd cell_6t
Xbit_r111_c222 bl[222] br[222] wl[111] vdd gnd cell_6t
Xbit_r112_c222 bl[222] br[222] wl[112] vdd gnd cell_6t
Xbit_r113_c222 bl[222] br[222] wl[113] vdd gnd cell_6t
Xbit_r114_c222 bl[222] br[222] wl[114] vdd gnd cell_6t
Xbit_r115_c222 bl[222] br[222] wl[115] vdd gnd cell_6t
Xbit_r116_c222 bl[222] br[222] wl[116] vdd gnd cell_6t
Xbit_r117_c222 bl[222] br[222] wl[117] vdd gnd cell_6t
Xbit_r118_c222 bl[222] br[222] wl[118] vdd gnd cell_6t
Xbit_r119_c222 bl[222] br[222] wl[119] vdd gnd cell_6t
Xbit_r120_c222 bl[222] br[222] wl[120] vdd gnd cell_6t
Xbit_r121_c222 bl[222] br[222] wl[121] vdd gnd cell_6t
Xbit_r122_c222 bl[222] br[222] wl[122] vdd gnd cell_6t
Xbit_r123_c222 bl[222] br[222] wl[123] vdd gnd cell_6t
Xbit_r124_c222 bl[222] br[222] wl[124] vdd gnd cell_6t
Xbit_r125_c222 bl[222] br[222] wl[125] vdd gnd cell_6t
Xbit_r126_c222 bl[222] br[222] wl[126] vdd gnd cell_6t
Xbit_r127_c222 bl[222] br[222] wl[127] vdd gnd cell_6t
Xbit_r0_c223 bl[223] br[223] wl[0] vdd gnd cell_6t
Xbit_r1_c223 bl[223] br[223] wl[1] vdd gnd cell_6t
Xbit_r2_c223 bl[223] br[223] wl[2] vdd gnd cell_6t
Xbit_r3_c223 bl[223] br[223] wl[3] vdd gnd cell_6t
Xbit_r4_c223 bl[223] br[223] wl[4] vdd gnd cell_6t
Xbit_r5_c223 bl[223] br[223] wl[5] vdd gnd cell_6t
Xbit_r6_c223 bl[223] br[223] wl[6] vdd gnd cell_6t
Xbit_r7_c223 bl[223] br[223] wl[7] vdd gnd cell_6t
Xbit_r8_c223 bl[223] br[223] wl[8] vdd gnd cell_6t
Xbit_r9_c223 bl[223] br[223] wl[9] vdd gnd cell_6t
Xbit_r10_c223 bl[223] br[223] wl[10] vdd gnd cell_6t
Xbit_r11_c223 bl[223] br[223] wl[11] vdd gnd cell_6t
Xbit_r12_c223 bl[223] br[223] wl[12] vdd gnd cell_6t
Xbit_r13_c223 bl[223] br[223] wl[13] vdd gnd cell_6t
Xbit_r14_c223 bl[223] br[223] wl[14] vdd gnd cell_6t
Xbit_r15_c223 bl[223] br[223] wl[15] vdd gnd cell_6t
Xbit_r16_c223 bl[223] br[223] wl[16] vdd gnd cell_6t
Xbit_r17_c223 bl[223] br[223] wl[17] vdd gnd cell_6t
Xbit_r18_c223 bl[223] br[223] wl[18] vdd gnd cell_6t
Xbit_r19_c223 bl[223] br[223] wl[19] vdd gnd cell_6t
Xbit_r20_c223 bl[223] br[223] wl[20] vdd gnd cell_6t
Xbit_r21_c223 bl[223] br[223] wl[21] vdd gnd cell_6t
Xbit_r22_c223 bl[223] br[223] wl[22] vdd gnd cell_6t
Xbit_r23_c223 bl[223] br[223] wl[23] vdd gnd cell_6t
Xbit_r24_c223 bl[223] br[223] wl[24] vdd gnd cell_6t
Xbit_r25_c223 bl[223] br[223] wl[25] vdd gnd cell_6t
Xbit_r26_c223 bl[223] br[223] wl[26] vdd gnd cell_6t
Xbit_r27_c223 bl[223] br[223] wl[27] vdd gnd cell_6t
Xbit_r28_c223 bl[223] br[223] wl[28] vdd gnd cell_6t
Xbit_r29_c223 bl[223] br[223] wl[29] vdd gnd cell_6t
Xbit_r30_c223 bl[223] br[223] wl[30] vdd gnd cell_6t
Xbit_r31_c223 bl[223] br[223] wl[31] vdd gnd cell_6t
Xbit_r32_c223 bl[223] br[223] wl[32] vdd gnd cell_6t
Xbit_r33_c223 bl[223] br[223] wl[33] vdd gnd cell_6t
Xbit_r34_c223 bl[223] br[223] wl[34] vdd gnd cell_6t
Xbit_r35_c223 bl[223] br[223] wl[35] vdd gnd cell_6t
Xbit_r36_c223 bl[223] br[223] wl[36] vdd gnd cell_6t
Xbit_r37_c223 bl[223] br[223] wl[37] vdd gnd cell_6t
Xbit_r38_c223 bl[223] br[223] wl[38] vdd gnd cell_6t
Xbit_r39_c223 bl[223] br[223] wl[39] vdd gnd cell_6t
Xbit_r40_c223 bl[223] br[223] wl[40] vdd gnd cell_6t
Xbit_r41_c223 bl[223] br[223] wl[41] vdd gnd cell_6t
Xbit_r42_c223 bl[223] br[223] wl[42] vdd gnd cell_6t
Xbit_r43_c223 bl[223] br[223] wl[43] vdd gnd cell_6t
Xbit_r44_c223 bl[223] br[223] wl[44] vdd gnd cell_6t
Xbit_r45_c223 bl[223] br[223] wl[45] vdd gnd cell_6t
Xbit_r46_c223 bl[223] br[223] wl[46] vdd gnd cell_6t
Xbit_r47_c223 bl[223] br[223] wl[47] vdd gnd cell_6t
Xbit_r48_c223 bl[223] br[223] wl[48] vdd gnd cell_6t
Xbit_r49_c223 bl[223] br[223] wl[49] vdd gnd cell_6t
Xbit_r50_c223 bl[223] br[223] wl[50] vdd gnd cell_6t
Xbit_r51_c223 bl[223] br[223] wl[51] vdd gnd cell_6t
Xbit_r52_c223 bl[223] br[223] wl[52] vdd gnd cell_6t
Xbit_r53_c223 bl[223] br[223] wl[53] vdd gnd cell_6t
Xbit_r54_c223 bl[223] br[223] wl[54] vdd gnd cell_6t
Xbit_r55_c223 bl[223] br[223] wl[55] vdd gnd cell_6t
Xbit_r56_c223 bl[223] br[223] wl[56] vdd gnd cell_6t
Xbit_r57_c223 bl[223] br[223] wl[57] vdd gnd cell_6t
Xbit_r58_c223 bl[223] br[223] wl[58] vdd gnd cell_6t
Xbit_r59_c223 bl[223] br[223] wl[59] vdd gnd cell_6t
Xbit_r60_c223 bl[223] br[223] wl[60] vdd gnd cell_6t
Xbit_r61_c223 bl[223] br[223] wl[61] vdd gnd cell_6t
Xbit_r62_c223 bl[223] br[223] wl[62] vdd gnd cell_6t
Xbit_r63_c223 bl[223] br[223] wl[63] vdd gnd cell_6t
Xbit_r64_c223 bl[223] br[223] wl[64] vdd gnd cell_6t
Xbit_r65_c223 bl[223] br[223] wl[65] vdd gnd cell_6t
Xbit_r66_c223 bl[223] br[223] wl[66] vdd gnd cell_6t
Xbit_r67_c223 bl[223] br[223] wl[67] vdd gnd cell_6t
Xbit_r68_c223 bl[223] br[223] wl[68] vdd gnd cell_6t
Xbit_r69_c223 bl[223] br[223] wl[69] vdd gnd cell_6t
Xbit_r70_c223 bl[223] br[223] wl[70] vdd gnd cell_6t
Xbit_r71_c223 bl[223] br[223] wl[71] vdd gnd cell_6t
Xbit_r72_c223 bl[223] br[223] wl[72] vdd gnd cell_6t
Xbit_r73_c223 bl[223] br[223] wl[73] vdd gnd cell_6t
Xbit_r74_c223 bl[223] br[223] wl[74] vdd gnd cell_6t
Xbit_r75_c223 bl[223] br[223] wl[75] vdd gnd cell_6t
Xbit_r76_c223 bl[223] br[223] wl[76] vdd gnd cell_6t
Xbit_r77_c223 bl[223] br[223] wl[77] vdd gnd cell_6t
Xbit_r78_c223 bl[223] br[223] wl[78] vdd gnd cell_6t
Xbit_r79_c223 bl[223] br[223] wl[79] vdd gnd cell_6t
Xbit_r80_c223 bl[223] br[223] wl[80] vdd gnd cell_6t
Xbit_r81_c223 bl[223] br[223] wl[81] vdd gnd cell_6t
Xbit_r82_c223 bl[223] br[223] wl[82] vdd gnd cell_6t
Xbit_r83_c223 bl[223] br[223] wl[83] vdd gnd cell_6t
Xbit_r84_c223 bl[223] br[223] wl[84] vdd gnd cell_6t
Xbit_r85_c223 bl[223] br[223] wl[85] vdd gnd cell_6t
Xbit_r86_c223 bl[223] br[223] wl[86] vdd gnd cell_6t
Xbit_r87_c223 bl[223] br[223] wl[87] vdd gnd cell_6t
Xbit_r88_c223 bl[223] br[223] wl[88] vdd gnd cell_6t
Xbit_r89_c223 bl[223] br[223] wl[89] vdd gnd cell_6t
Xbit_r90_c223 bl[223] br[223] wl[90] vdd gnd cell_6t
Xbit_r91_c223 bl[223] br[223] wl[91] vdd gnd cell_6t
Xbit_r92_c223 bl[223] br[223] wl[92] vdd gnd cell_6t
Xbit_r93_c223 bl[223] br[223] wl[93] vdd gnd cell_6t
Xbit_r94_c223 bl[223] br[223] wl[94] vdd gnd cell_6t
Xbit_r95_c223 bl[223] br[223] wl[95] vdd gnd cell_6t
Xbit_r96_c223 bl[223] br[223] wl[96] vdd gnd cell_6t
Xbit_r97_c223 bl[223] br[223] wl[97] vdd gnd cell_6t
Xbit_r98_c223 bl[223] br[223] wl[98] vdd gnd cell_6t
Xbit_r99_c223 bl[223] br[223] wl[99] vdd gnd cell_6t
Xbit_r100_c223 bl[223] br[223] wl[100] vdd gnd cell_6t
Xbit_r101_c223 bl[223] br[223] wl[101] vdd gnd cell_6t
Xbit_r102_c223 bl[223] br[223] wl[102] vdd gnd cell_6t
Xbit_r103_c223 bl[223] br[223] wl[103] vdd gnd cell_6t
Xbit_r104_c223 bl[223] br[223] wl[104] vdd gnd cell_6t
Xbit_r105_c223 bl[223] br[223] wl[105] vdd gnd cell_6t
Xbit_r106_c223 bl[223] br[223] wl[106] vdd gnd cell_6t
Xbit_r107_c223 bl[223] br[223] wl[107] vdd gnd cell_6t
Xbit_r108_c223 bl[223] br[223] wl[108] vdd gnd cell_6t
Xbit_r109_c223 bl[223] br[223] wl[109] vdd gnd cell_6t
Xbit_r110_c223 bl[223] br[223] wl[110] vdd gnd cell_6t
Xbit_r111_c223 bl[223] br[223] wl[111] vdd gnd cell_6t
Xbit_r112_c223 bl[223] br[223] wl[112] vdd gnd cell_6t
Xbit_r113_c223 bl[223] br[223] wl[113] vdd gnd cell_6t
Xbit_r114_c223 bl[223] br[223] wl[114] vdd gnd cell_6t
Xbit_r115_c223 bl[223] br[223] wl[115] vdd gnd cell_6t
Xbit_r116_c223 bl[223] br[223] wl[116] vdd gnd cell_6t
Xbit_r117_c223 bl[223] br[223] wl[117] vdd gnd cell_6t
Xbit_r118_c223 bl[223] br[223] wl[118] vdd gnd cell_6t
Xbit_r119_c223 bl[223] br[223] wl[119] vdd gnd cell_6t
Xbit_r120_c223 bl[223] br[223] wl[120] vdd gnd cell_6t
Xbit_r121_c223 bl[223] br[223] wl[121] vdd gnd cell_6t
Xbit_r122_c223 bl[223] br[223] wl[122] vdd gnd cell_6t
Xbit_r123_c223 bl[223] br[223] wl[123] vdd gnd cell_6t
Xbit_r124_c223 bl[223] br[223] wl[124] vdd gnd cell_6t
Xbit_r125_c223 bl[223] br[223] wl[125] vdd gnd cell_6t
Xbit_r126_c223 bl[223] br[223] wl[126] vdd gnd cell_6t
Xbit_r127_c223 bl[223] br[223] wl[127] vdd gnd cell_6t
Xbit_r0_c224 bl[224] br[224] wl[0] vdd gnd cell_6t
Xbit_r1_c224 bl[224] br[224] wl[1] vdd gnd cell_6t
Xbit_r2_c224 bl[224] br[224] wl[2] vdd gnd cell_6t
Xbit_r3_c224 bl[224] br[224] wl[3] vdd gnd cell_6t
Xbit_r4_c224 bl[224] br[224] wl[4] vdd gnd cell_6t
Xbit_r5_c224 bl[224] br[224] wl[5] vdd gnd cell_6t
Xbit_r6_c224 bl[224] br[224] wl[6] vdd gnd cell_6t
Xbit_r7_c224 bl[224] br[224] wl[7] vdd gnd cell_6t
Xbit_r8_c224 bl[224] br[224] wl[8] vdd gnd cell_6t
Xbit_r9_c224 bl[224] br[224] wl[9] vdd gnd cell_6t
Xbit_r10_c224 bl[224] br[224] wl[10] vdd gnd cell_6t
Xbit_r11_c224 bl[224] br[224] wl[11] vdd gnd cell_6t
Xbit_r12_c224 bl[224] br[224] wl[12] vdd gnd cell_6t
Xbit_r13_c224 bl[224] br[224] wl[13] vdd gnd cell_6t
Xbit_r14_c224 bl[224] br[224] wl[14] vdd gnd cell_6t
Xbit_r15_c224 bl[224] br[224] wl[15] vdd gnd cell_6t
Xbit_r16_c224 bl[224] br[224] wl[16] vdd gnd cell_6t
Xbit_r17_c224 bl[224] br[224] wl[17] vdd gnd cell_6t
Xbit_r18_c224 bl[224] br[224] wl[18] vdd gnd cell_6t
Xbit_r19_c224 bl[224] br[224] wl[19] vdd gnd cell_6t
Xbit_r20_c224 bl[224] br[224] wl[20] vdd gnd cell_6t
Xbit_r21_c224 bl[224] br[224] wl[21] vdd gnd cell_6t
Xbit_r22_c224 bl[224] br[224] wl[22] vdd gnd cell_6t
Xbit_r23_c224 bl[224] br[224] wl[23] vdd gnd cell_6t
Xbit_r24_c224 bl[224] br[224] wl[24] vdd gnd cell_6t
Xbit_r25_c224 bl[224] br[224] wl[25] vdd gnd cell_6t
Xbit_r26_c224 bl[224] br[224] wl[26] vdd gnd cell_6t
Xbit_r27_c224 bl[224] br[224] wl[27] vdd gnd cell_6t
Xbit_r28_c224 bl[224] br[224] wl[28] vdd gnd cell_6t
Xbit_r29_c224 bl[224] br[224] wl[29] vdd gnd cell_6t
Xbit_r30_c224 bl[224] br[224] wl[30] vdd gnd cell_6t
Xbit_r31_c224 bl[224] br[224] wl[31] vdd gnd cell_6t
Xbit_r32_c224 bl[224] br[224] wl[32] vdd gnd cell_6t
Xbit_r33_c224 bl[224] br[224] wl[33] vdd gnd cell_6t
Xbit_r34_c224 bl[224] br[224] wl[34] vdd gnd cell_6t
Xbit_r35_c224 bl[224] br[224] wl[35] vdd gnd cell_6t
Xbit_r36_c224 bl[224] br[224] wl[36] vdd gnd cell_6t
Xbit_r37_c224 bl[224] br[224] wl[37] vdd gnd cell_6t
Xbit_r38_c224 bl[224] br[224] wl[38] vdd gnd cell_6t
Xbit_r39_c224 bl[224] br[224] wl[39] vdd gnd cell_6t
Xbit_r40_c224 bl[224] br[224] wl[40] vdd gnd cell_6t
Xbit_r41_c224 bl[224] br[224] wl[41] vdd gnd cell_6t
Xbit_r42_c224 bl[224] br[224] wl[42] vdd gnd cell_6t
Xbit_r43_c224 bl[224] br[224] wl[43] vdd gnd cell_6t
Xbit_r44_c224 bl[224] br[224] wl[44] vdd gnd cell_6t
Xbit_r45_c224 bl[224] br[224] wl[45] vdd gnd cell_6t
Xbit_r46_c224 bl[224] br[224] wl[46] vdd gnd cell_6t
Xbit_r47_c224 bl[224] br[224] wl[47] vdd gnd cell_6t
Xbit_r48_c224 bl[224] br[224] wl[48] vdd gnd cell_6t
Xbit_r49_c224 bl[224] br[224] wl[49] vdd gnd cell_6t
Xbit_r50_c224 bl[224] br[224] wl[50] vdd gnd cell_6t
Xbit_r51_c224 bl[224] br[224] wl[51] vdd gnd cell_6t
Xbit_r52_c224 bl[224] br[224] wl[52] vdd gnd cell_6t
Xbit_r53_c224 bl[224] br[224] wl[53] vdd gnd cell_6t
Xbit_r54_c224 bl[224] br[224] wl[54] vdd gnd cell_6t
Xbit_r55_c224 bl[224] br[224] wl[55] vdd gnd cell_6t
Xbit_r56_c224 bl[224] br[224] wl[56] vdd gnd cell_6t
Xbit_r57_c224 bl[224] br[224] wl[57] vdd gnd cell_6t
Xbit_r58_c224 bl[224] br[224] wl[58] vdd gnd cell_6t
Xbit_r59_c224 bl[224] br[224] wl[59] vdd gnd cell_6t
Xbit_r60_c224 bl[224] br[224] wl[60] vdd gnd cell_6t
Xbit_r61_c224 bl[224] br[224] wl[61] vdd gnd cell_6t
Xbit_r62_c224 bl[224] br[224] wl[62] vdd gnd cell_6t
Xbit_r63_c224 bl[224] br[224] wl[63] vdd gnd cell_6t
Xbit_r64_c224 bl[224] br[224] wl[64] vdd gnd cell_6t
Xbit_r65_c224 bl[224] br[224] wl[65] vdd gnd cell_6t
Xbit_r66_c224 bl[224] br[224] wl[66] vdd gnd cell_6t
Xbit_r67_c224 bl[224] br[224] wl[67] vdd gnd cell_6t
Xbit_r68_c224 bl[224] br[224] wl[68] vdd gnd cell_6t
Xbit_r69_c224 bl[224] br[224] wl[69] vdd gnd cell_6t
Xbit_r70_c224 bl[224] br[224] wl[70] vdd gnd cell_6t
Xbit_r71_c224 bl[224] br[224] wl[71] vdd gnd cell_6t
Xbit_r72_c224 bl[224] br[224] wl[72] vdd gnd cell_6t
Xbit_r73_c224 bl[224] br[224] wl[73] vdd gnd cell_6t
Xbit_r74_c224 bl[224] br[224] wl[74] vdd gnd cell_6t
Xbit_r75_c224 bl[224] br[224] wl[75] vdd gnd cell_6t
Xbit_r76_c224 bl[224] br[224] wl[76] vdd gnd cell_6t
Xbit_r77_c224 bl[224] br[224] wl[77] vdd gnd cell_6t
Xbit_r78_c224 bl[224] br[224] wl[78] vdd gnd cell_6t
Xbit_r79_c224 bl[224] br[224] wl[79] vdd gnd cell_6t
Xbit_r80_c224 bl[224] br[224] wl[80] vdd gnd cell_6t
Xbit_r81_c224 bl[224] br[224] wl[81] vdd gnd cell_6t
Xbit_r82_c224 bl[224] br[224] wl[82] vdd gnd cell_6t
Xbit_r83_c224 bl[224] br[224] wl[83] vdd gnd cell_6t
Xbit_r84_c224 bl[224] br[224] wl[84] vdd gnd cell_6t
Xbit_r85_c224 bl[224] br[224] wl[85] vdd gnd cell_6t
Xbit_r86_c224 bl[224] br[224] wl[86] vdd gnd cell_6t
Xbit_r87_c224 bl[224] br[224] wl[87] vdd gnd cell_6t
Xbit_r88_c224 bl[224] br[224] wl[88] vdd gnd cell_6t
Xbit_r89_c224 bl[224] br[224] wl[89] vdd gnd cell_6t
Xbit_r90_c224 bl[224] br[224] wl[90] vdd gnd cell_6t
Xbit_r91_c224 bl[224] br[224] wl[91] vdd gnd cell_6t
Xbit_r92_c224 bl[224] br[224] wl[92] vdd gnd cell_6t
Xbit_r93_c224 bl[224] br[224] wl[93] vdd gnd cell_6t
Xbit_r94_c224 bl[224] br[224] wl[94] vdd gnd cell_6t
Xbit_r95_c224 bl[224] br[224] wl[95] vdd gnd cell_6t
Xbit_r96_c224 bl[224] br[224] wl[96] vdd gnd cell_6t
Xbit_r97_c224 bl[224] br[224] wl[97] vdd gnd cell_6t
Xbit_r98_c224 bl[224] br[224] wl[98] vdd gnd cell_6t
Xbit_r99_c224 bl[224] br[224] wl[99] vdd gnd cell_6t
Xbit_r100_c224 bl[224] br[224] wl[100] vdd gnd cell_6t
Xbit_r101_c224 bl[224] br[224] wl[101] vdd gnd cell_6t
Xbit_r102_c224 bl[224] br[224] wl[102] vdd gnd cell_6t
Xbit_r103_c224 bl[224] br[224] wl[103] vdd gnd cell_6t
Xbit_r104_c224 bl[224] br[224] wl[104] vdd gnd cell_6t
Xbit_r105_c224 bl[224] br[224] wl[105] vdd gnd cell_6t
Xbit_r106_c224 bl[224] br[224] wl[106] vdd gnd cell_6t
Xbit_r107_c224 bl[224] br[224] wl[107] vdd gnd cell_6t
Xbit_r108_c224 bl[224] br[224] wl[108] vdd gnd cell_6t
Xbit_r109_c224 bl[224] br[224] wl[109] vdd gnd cell_6t
Xbit_r110_c224 bl[224] br[224] wl[110] vdd gnd cell_6t
Xbit_r111_c224 bl[224] br[224] wl[111] vdd gnd cell_6t
Xbit_r112_c224 bl[224] br[224] wl[112] vdd gnd cell_6t
Xbit_r113_c224 bl[224] br[224] wl[113] vdd gnd cell_6t
Xbit_r114_c224 bl[224] br[224] wl[114] vdd gnd cell_6t
Xbit_r115_c224 bl[224] br[224] wl[115] vdd gnd cell_6t
Xbit_r116_c224 bl[224] br[224] wl[116] vdd gnd cell_6t
Xbit_r117_c224 bl[224] br[224] wl[117] vdd gnd cell_6t
Xbit_r118_c224 bl[224] br[224] wl[118] vdd gnd cell_6t
Xbit_r119_c224 bl[224] br[224] wl[119] vdd gnd cell_6t
Xbit_r120_c224 bl[224] br[224] wl[120] vdd gnd cell_6t
Xbit_r121_c224 bl[224] br[224] wl[121] vdd gnd cell_6t
Xbit_r122_c224 bl[224] br[224] wl[122] vdd gnd cell_6t
Xbit_r123_c224 bl[224] br[224] wl[123] vdd gnd cell_6t
Xbit_r124_c224 bl[224] br[224] wl[124] vdd gnd cell_6t
Xbit_r125_c224 bl[224] br[224] wl[125] vdd gnd cell_6t
Xbit_r126_c224 bl[224] br[224] wl[126] vdd gnd cell_6t
Xbit_r127_c224 bl[224] br[224] wl[127] vdd gnd cell_6t
Xbit_r0_c225 bl[225] br[225] wl[0] vdd gnd cell_6t
Xbit_r1_c225 bl[225] br[225] wl[1] vdd gnd cell_6t
Xbit_r2_c225 bl[225] br[225] wl[2] vdd gnd cell_6t
Xbit_r3_c225 bl[225] br[225] wl[3] vdd gnd cell_6t
Xbit_r4_c225 bl[225] br[225] wl[4] vdd gnd cell_6t
Xbit_r5_c225 bl[225] br[225] wl[5] vdd gnd cell_6t
Xbit_r6_c225 bl[225] br[225] wl[6] vdd gnd cell_6t
Xbit_r7_c225 bl[225] br[225] wl[7] vdd gnd cell_6t
Xbit_r8_c225 bl[225] br[225] wl[8] vdd gnd cell_6t
Xbit_r9_c225 bl[225] br[225] wl[9] vdd gnd cell_6t
Xbit_r10_c225 bl[225] br[225] wl[10] vdd gnd cell_6t
Xbit_r11_c225 bl[225] br[225] wl[11] vdd gnd cell_6t
Xbit_r12_c225 bl[225] br[225] wl[12] vdd gnd cell_6t
Xbit_r13_c225 bl[225] br[225] wl[13] vdd gnd cell_6t
Xbit_r14_c225 bl[225] br[225] wl[14] vdd gnd cell_6t
Xbit_r15_c225 bl[225] br[225] wl[15] vdd gnd cell_6t
Xbit_r16_c225 bl[225] br[225] wl[16] vdd gnd cell_6t
Xbit_r17_c225 bl[225] br[225] wl[17] vdd gnd cell_6t
Xbit_r18_c225 bl[225] br[225] wl[18] vdd gnd cell_6t
Xbit_r19_c225 bl[225] br[225] wl[19] vdd gnd cell_6t
Xbit_r20_c225 bl[225] br[225] wl[20] vdd gnd cell_6t
Xbit_r21_c225 bl[225] br[225] wl[21] vdd gnd cell_6t
Xbit_r22_c225 bl[225] br[225] wl[22] vdd gnd cell_6t
Xbit_r23_c225 bl[225] br[225] wl[23] vdd gnd cell_6t
Xbit_r24_c225 bl[225] br[225] wl[24] vdd gnd cell_6t
Xbit_r25_c225 bl[225] br[225] wl[25] vdd gnd cell_6t
Xbit_r26_c225 bl[225] br[225] wl[26] vdd gnd cell_6t
Xbit_r27_c225 bl[225] br[225] wl[27] vdd gnd cell_6t
Xbit_r28_c225 bl[225] br[225] wl[28] vdd gnd cell_6t
Xbit_r29_c225 bl[225] br[225] wl[29] vdd gnd cell_6t
Xbit_r30_c225 bl[225] br[225] wl[30] vdd gnd cell_6t
Xbit_r31_c225 bl[225] br[225] wl[31] vdd gnd cell_6t
Xbit_r32_c225 bl[225] br[225] wl[32] vdd gnd cell_6t
Xbit_r33_c225 bl[225] br[225] wl[33] vdd gnd cell_6t
Xbit_r34_c225 bl[225] br[225] wl[34] vdd gnd cell_6t
Xbit_r35_c225 bl[225] br[225] wl[35] vdd gnd cell_6t
Xbit_r36_c225 bl[225] br[225] wl[36] vdd gnd cell_6t
Xbit_r37_c225 bl[225] br[225] wl[37] vdd gnd cell_6t
Xbit_r38_c225 bl[225] br[225] wl[38] vdd gnd cell_6t
Xbit_r39_c225 bl[225] br[225] wl[39] vdd gnd cell_6t
Xbit_r40_c225 bl[225] br[225] wl[40] vdd gnd cell_6t
Xbit_r41_c225 bl[225] br[225] wl[41] vdd gnd cell_6t
Xbit_r42_c225 bl[225] br[225] wl[42] vdd gnd cell_6t
Xbit_r43_c225 bl[225] br[225] wl[43] vdd gnd cell_6t
Xbit_r44_c225 bl[225] br[225] wl[44] vdd gnd cell_6t
Xbit_r45_c225 bl[225] br[225] wl[45] vdd gnd cell_6t
Xbit_r46_c225 bl[225] br[225] wl[46] vdd gnd cell_6t
Xbit_r47_c225 bl[225] br[225] wl[47] vdd gnd cell_6t
Xbit_r48_c225 bl[225] br[225] wl[48] vdd gnd cell_6t
Xbit_r49_c225 bl[225] br[225] wl[49] vdd gnd cell_6t
Xbit_r50_c225 bl[225] br[225] wl[50] vdd gnd cell_6t
Xbit_r51_c225 bl[225] br[225] wl[51] vdd gnd cell_6t
Xbit_r52_c225 bl[225] br[225] wl[52] vdd gnd cell_6t
Xbit_r53_c225 bl[225] br[225] wl[53] vdd gnd cell_6t
Xbit_r54_c225 bl[225] br[225] wl[54] vdd gnd cell_6t
Xbit_r55_c225 bl[225] br[225] wl[55] vdd gnd cell_6t
Xbit_r56_c225 bl[225] br[225] wl[56] vdd gnd cell_6t
Xbit_r57_c225 bl[225] br[225] wl[57] vdd gnd cell_6t
Xbit_r58_c225 bl[225] br[225] wl[58] vdd gnd cell_6t
Xbit_r59_c225 bl[225] br[225] wl[59] vdd gnd cell_6t
Xbit_r60_c225 bl[225] br[225] wl[60] vdd gnd cell_6t
Xbit_r61_c225 bl[225] br[225] wl[61] vdd gnd cell_6t
Xbit_r62_c225 bl[225] br[225] wl[62] vdd gnd cell_6t
Xbit_r63_c225 bl[225] br[225] wl[63] vdd gnd cell_6t
Xbit_r64_c225 bl[225] br[225] wl[64] vdd gnd cell_6t
Xbit_r65_c225 bl[225] br[225] wl[65] vdd gnd cell_6t
Xbit_r66_c225 bl[225] br[225] wl[66] vdd gnd cell_6t
Xbit_r67_c225 bl[225] br[225] wl[67] vdd gnd cell_6t
Xbit_r68_c225 bl[225] br[225] wl[68] vdd gnd cell_6t
Xbit_r69_c225 bl[225] br[225] wl[69] vdd gnd cell_6t
Xbit_r70_c225 bl[225] br[225] wl[70] vdd gnd cell_6t
Xbit_r71_c225 bl[225] br[225] wl[71] vdd gnd cell_6t
Xbit_r72_c225 bl[225] br[225] wl[72] vdd gnd cell_6t
Xbit_r73_c225 bl[225] br[225] wl[73] vdd gnd cell_6t
Xbit_r74_c225 bl[225] br[225] wl[74] vdd gnd cell_6t
Xbit_r75_c225 bl[225] br[225] wl[75] vdd gnd cell_6t
Xbit_r76_c225 bl[225] br[225] wl[76] vdd gnd cell_6t
Xbit_r77_c225 bl[225] br[225] wl[77] vdd gnd cell_6t
Xbit_r78_c225 bl[225] br[225] wl[78] vdd gnd cell_6t
Xbit_r79_c225 bl[225] br[225] wl[79] vdd gnd cell_6t
Xbit_r80_c225 bl[225] br[225] wl[80] vdd gnd cell_6t
Xbit_r81_c225 bl[225] br[225] wl[81] vdd gnd cell_6t
Xbit_r82_c225 bl[225] br[225] wl[82] vdd gnd cell_6t
Xbit_r83_c225 bl[225] br[225] wl[83] vdd gnd cell_6t
Xbit_r84_c225 bl[225] br[225] wl[84] vdd gnd cell_6t
Xbit_r85_c225 bl[225] br[225] wl[85] vdd gnd cell_6t
Xbit_r86_c225 bl[225] br[225] wl[86] vdd gnd cell_6t
Xbit_r87_c225 bl[225] br[225] wl[87] vdd gnd cell_6t
Xbit_r88_c225 bl[225] br[225] wl[88] vdd gnd cell_6t
Xbit_r89_c225 bl[225] br[225] wl[89] vdd gnd cell_6t
Xbit_r90_c225 bl[225] br[225] wl[90] vdd gnd cell_6t
Xbit_r91_c225 bl[225] br[225] wl[91] vdd gnd cell_6t
Xbit_r92_c225 bl[225] br[225] wl[92] vdd gnd cell_6t
Xbit_r93_c225 bl[225] br[225] wl[93] vdd gnd cell_6t
Xbit_r94_c225 bl[225] br[225] wl[94] vdd gnd cell_6t
Xbit_r95_c225 bl[225] br[225] wl[95] vdd gnd cell_6t
Xbit_r96_c225 bl[225] br[225] wl[96] vdd gnd cell_6t
Xbit_r97_c225 bl[225] br[225] wl[97] vdd gnd cell_6t
Xbit_r98_c225 bl[225] br[225] wl[98] vdd gnd cell_6t
Xbit_r99_c225 bl[225] br[225] wl[99] vdd gnd cell_6t
Xbit_r100_c225 bl[225] br[225] wl[100] vdd gnd cell_6t
Xbit_r101_c225 bl[225] br[225] wl[101] vdd gnd cell_6t
Xbit_r102_c225 bl[225] br[225] wl[102] vdd gnd cell_6t
Xbit_r103_c225 bl[225] br[225] wl[103] vdd gnd cell_6t
Xbit_r104_c225 bl[225] br[225] wl[104] vdd gnd cell_6t
Xbit_r105_c225 bl[225] br[225] wl[105] vdd gnd cell_6t
Xbit_r106_c225 bl[225] br[225] wl[106] vdd gnd cell_6t
Xbit_r107_c225 bl[225] br[225] wl[107] vdd gnd cell_6t
Xbit_r108_c225 bl[225] br[225] wl[108] vdd gnd cell_6t
Xbit_r109_c225 bl[225] br[225] wl[109] vdd gnd cell_6t
Xbit_r110_c225 bl[225] br[225] wl[110] vdd gnd cell_6t
Xbit_r111_c225 bl[225] br[225] wl[111] vdd gnd cell_6t
Xbit_r112_c225 bl[225] br[225] wl[112] vdd gnd cell_6t
Xbit_r113_c225 bl[225] br[225] wl[113] vdd gnd cell_6t
Xbit_r114_c225 bl[225] br[225] wl[114] vdd gnd cell_6t
Xbit_r115_c225 bl[225] br[225] wl[115] vdd gnd cell_6t
Xbit_r116_c225 bl[225] br[225] wl[116] vdd gnd cell_6t
Xbit_r117_c225 bl[225] br[225] wl[117] vdd gnd cell_6t
Xbit_r118_c225 bl[225] br[225] wl[118] vdd gnd cell_6t
Xbit_r119_c225 bl[225] br[225] wl[119] vdd gnd cell_6t
Xbit_r120_c225 bl[225] br[225] wl[120] vdd gnd cell_6t
Xbit_r121_c225 bl[225] br[225] wl[121] vdd gnd cell_6t
Xbit_r122_c225 bl[225] br[225] wl[122] vdd gnd cell_6t
Xbit_r123_c225 bl[225] br[225] wl[123] vdd gnd cell_6t
Xbit_r124_c225 bl[225] br[225] wl[124] vdd gnd cell_6t
Xbit_r125_c225 bl[225] br[225] wl[125] vdd gnd cell_6t
Xbit_r126_c225 bl[225] br[225] wl[126] vdd gnd cell_6t
Xbit_r127_c225 bl[225] br[225] wl[127] vdd gnd cell_6t
Xbit_r0_c226 bl[226] br[226] wl[0] vdd gnd cell_6t
Xbit_r1_c226 bl[226] br[226] wl[1] vdd gnd cell_6t
Xbit_r2_c226 bl[226] br[226] wl[2] vdd gnd cell_6t
Xbit_r3_c226 bl[226] br[226] wl[3] vdd gnd cell_6t
Xbit_r4_c226 bl[226] br[226] wl[4] vdd gnd cell_6t
Xbit_r5_c226 bl[226] br[226] wl[5] vdd gnd cell_6t
Xbit_r6_c226 bl[226] br[226] wl[6] vdd gnd cell_6t
Xbit_r7_c226 bl[226] br[226] wl[7] vdd gnd cell_6t
Xbit_r8_c226 bl[226] br[226] wl[8] vdd gnd cell_6t
Xbit_r9_c226 bl[226] br[226] wl[9] vdd gnd cell_6t
Xbit_r10_c226 bl[226] br[226] wl[10] vdd gnd cell_6t
Xbit_r11_c226 bl[226] br[226] wl[11] vdd gnd cell_6t
Xbit_r12_c226 bl[226] br[226] wl[12] vdd gnd cell_6t
Xbit_r13_c226 bl[226] br[226] wl[13] vdd gnd cell_6t
Xbit_r14_c226 bl[226] br[226] wl[14] vdd gnd cell_6t
Xbit_r15_c226 bl[226] br[226] wl[15] vdd gnd cell_6t
Xbit_r16_c226 bl[226] br[226] wl[16] vdd gnd cell_6t
Xbit_r17_c226 bl[226] br[226] wl[17] vdd gnd cell_6t
Xbit_r18_c226 bl[226] br[226] wl[18] vdd gnd cell_6t
Xbit_r19_c226 bl[226] br[226] wl[19] vdd gnd cell_6t
Xbit_r20_c226 bl[226] br[226] wl[20] vdd gnd cell_6t
Xbit_r21_c226 bl[226] br[226] wl[21] vdd gnd cell_6t
Xbit_r22_c226 bl[226] br[226] wl[22] vdd gnd cell_6t
Xbit_r23_c226 bl[226] br[226] wl[23] vdd gnd cell_6t
Xbit_r24_c226 bl[226] br[226] wl[24] vdd gnd cell_6t
Xbit_r25_c226 bl[226] br[226] wl[25] vdd gnd cell_6t
Xbit_r26_c226 bl[226] br[226] wl[26] vdd gnd cell_6t
Xbit_r27_c226 bl[226] br[226] wl[27] vdd gnd cell_6t
Xbit_r28_c226 bl[226] br[226] wl[28] vdd gnd cell_6t
Xbit_r29_c226 bl[226] br[226] wl[29] vdd gnd cell_6t
Xbit_r30_c226 bl[226] br[226] wl[30] vdd gnd cell_6t
Xbit_r31_c226 bl[226] br[226] wl[31] vdd gnd cell_6t
Xbit_r32_c226 bl[226] br[226] wl[32] vdd gnd cell_6t
Xbit_r33_c226 bl[226] br[226] wl[33] vdd gnd cell_6t
Xbit_r34_c226 bl[226] br[226] wl[34] vdd gnd cell_6t
Xbit_r35_c226 bl[226] br[226] wl[35] vdd gnd cell_6t
Xbit_r36_c226 bl[226] br[226] wl[36] vdd gnd cell_6t
Xbit_r37_c226 bl[226] br[226] wl[37] vdd gnd cell_6t
Xbit_r38_c226 bl[226] br[226] wl[38] vdd gnd cell_6t
Xbit_r39_c226 bl[226] br[226] wl[39] vdd gnd cell_6t
Xbit_r40_c226 bl[226] br[226] wl[40] vdd gnd cell_6t
Xbit_r41_c226 bl[226] br[226] wl[41] vdd gnd cell_6t
Xbit_r42_c226 bl[226] br[226] wl[42] vdd gnd cell_6t
Xbit_r43_c226 bl[226] br[226] wl[43] vdd gnd cell_6t
Xbit_r44_c226 bl[226] br[226] wl[44] vdd gnd cell_6t
Xbit_r45_c226 bl[226] br[226] wl[45] vdd gnd cell_6t
Xbit_r46_c226 bl[226] br[226] wl[46] vdd gnd cell_6t
Xbit_r47_c226 bl[226] br[226] wl[47] vdd gnd cell_6t
Xbit_r48_c226 bl[226] br[226] wl[48] vdd gnd cell_6t
Xbit_r49_c226 bl[226] br[226] wl[49] vdd gnd cell_6t
Xbit_r50_c226 bl[226] br[226] wl[50] vdd gnd cell_6t
Xbit_r51_c226 bl[226] br[226] wl[51] vdd gnd cell_6t
Xbit_r52_c226 bl[226] br[226] wl[52] vdd gnd cell_6t
Xbit_r53_c226 bl[226] br[226] wl[53] vdd gnd cell_6t
Xbit_r54_c226 bl[226] br[226] wl[54] vdd gnd cell_6t
Xbit_r55_c226 bl[226] br[226] wl[55] vdd gnd cell_6t
Xbit_r56_c226 bl[226] br[226] wl[56] vdd gnd cell_6t
Xbit_r57_c226 bl[226] br[226] wl[57] vdd gnd cell_6t
Xbit_r58_c226 bl[226] br[226] wl[58] vdd gnd cell_6t
Xbit_r59_c226 bl[226] br[226] wl[59] vdd gnd cell_6t
Xbit_r60_c226 bl[226] br[226] wl[60] vdd gnd cell_6t
Xbit_r61_c226 bl[226] br[226] wl[61] vdd gnd cell_6t
Xbit_r62_c226 bl[226] br[226] wl[62] vdd gnd cell_6t
Xbit_r63_c226 bl[226] br[226] wl[63] vdd gnd cell_6t
Xbit_r64_c226 bl[226] br[226] wl[64] vdd gnd cell_6t
Xbit_r65_c226 bl[226] br[226] wl[65] vdd gnd cell_6t
Xbit_r66_c226 bl[226] br[226] wl[66] vdd gnd cell_6t
Xbit_r67_c226 bl[226] br[226] wl[67] vdd gnd cell_6t
Xbit_r68_c226 bl[226] br[226] wl[68] vdd gnd cell_6t
Xbit_r69_c226 bl[226] br[226] wl[69] vdd gnd cell_6t
Xbit_r70_c226 bl[226] br[226] wl[70] vdd gnd cell_6t
Xbit_r71_c226 bl[226] br[226] wl[71] vdd gnd cell_6t
Xbit_r72_c226 bl[226] br[226] wl[72] vdd gnd cell_6t
Xbit_r73_c226 bl[226] br[226] wl[73] vdd gnd cell_6t
Xbit_r74_c226 bl[226] br[226] wl[74] vdd gnd cell_6t
Xbit_r75_c226 bl[226] br[226] wl[75] vdd gnd cell_6t
Xbit_r76_c226 bl[226] br[226] wl[76] vdd gnd cell_6t
Xbit_r77_c226 bl[226] br[226] wl[77] vdd gnd cell_6t
Xbit_r78_c226 bl[226] br[226] wl[78] vdd gnd cell_6t
Xbit_r79_c226 bl[226] br[226] wl[79] vdd gnd cell_6t
Xbit_r80_c226 bl[226] br[226] wl[80] vdd gnd cell_6t
Xbit_r81_c226 bl[226] br[226] wl[81] vdd gnd cell_6t
Xbit_r82_c226 bl[226] br[226] wl[82] vdd gnd cell_6t
Xbit_r83_c226 bl[226] br[226] wl[83] vdd gnd cell_6t
Xbit_r84_c226 bl[226] br[226] wl[84] vdd gnd cell_6t
Xbit_r85_c226 bl[226] br[226] wl[85] vdd gnd cell_6t
Xbit_r86_c226 bl[226] br[226] wl[86] vdd gnd cell_6t
Xbit_r87_c226 bl[226] br[226] wl[87] vdd gnd cell_6t
Xbit_r88_c226 bl[226] br[226] wl[88] vdd gnd cell_6t
Xbit_r89_c226 bl[226] br[226] wl[89] vdd gnd cell_6t
Xbit_r90_c226 bl[226] br[226] wl[90] vdd gnd cell_6t
Xbit_r91_c226 bl[226] br[226] wl[91] vdd gnd cell_6t
Xbit_r92_c226 bl[226] br[226] wl[92] vdd gnd cell_6t
Xbit_r93_c226 bl[226] br[226] wl[93] vdd gnd cell_6t
Xbit_r94_c226 bl[226] br[226] wl[94] vdd gnd cell_6t
Xbit_r95_c226 bl[226] br[226] wl[95] vdd gnd cell_6t
Xbit_r96_c226 bl[226] br[226] wl[96] vdd gnd cell_6t
Xbit_r97_c226 bl[226] br[226] wl[97] vdd gnd cell_6t
Xbit_r98_c226 bl[226] br[226] wl[98] vdd gnd cell_6t
Xbit_r99_c226 bl[226] br[226] wl[99] vdd gnd cell_6t
Xbit_r100_c226 bl[226] br[226] wl[100] vdd gnd cell_6t
Xbit_r101_c226 bl[226] br[226] wl[101] vdd gnd cell_6t
Xbit_r102_c226 bl[226] br[226] wl[102] vdd gnd cell_6t
Xbit_r103_c226 bl[226] br[226] wl[103] vdd gnd cell_6t
Xbit_r104_c226 bl[226] br[226] wl[104] vdd gnd cell_6t
Xbit_r105_c226 bl[226] br[226] wl[105] vdd gnd cell_6t
Xbit_r106_c226 bl[226] br[226] wl[106] vdd gnd cell_6t
Xbit_r107_c226 bl[226] br[226] wl[107] vdd gnd cell_6t
Xbit_r108_c226 bl[226] br[226] wl[108] vdd gnd cell_6t
Xbit_r109_c226 bl[226] br[226] wl[109] vdd gnd cell_6t
Xbit_r110_c226 bl[226] br[226] wl[110] vdd gnd cell_6t
Xbit_r111_c226 bl[226] br[226] wl[111] vdd gnd cell_6t
Xbit_r112_c226 bl[226] br[226] wl[112] vdd gnd cell_6t
Xbit_r113_c226 bl[226] br[226] wl[113] vdd gnd cell_6t
Xbit_r114_c226 bl[226] br[226] wl[114] vdd gnd cell_6t
Xbit_r115_c226 bl[226] br[226] wl[115] vdd gnd cell_6t
Xbit_r116_c226 bl[226] br[226] wl[116] vdd gnd cell_6t
Xbit_r117_c226 bl[226] br[226] wl[117] vdd gnd cell_6t
Xbit_r118_c226 bl[226] br[226] wl[118] vdd gnd cell_6t
Xbit_r119_c226 bl[226] br[226] wl[119] vdd gnd cell_6t
Xbit_r120_c226 bl[226] br[226] wl[120] vdd gnd cell_6t
Xbit_r121_c226 bl[226] br[226] wl[121] vdd gnd cell_6t
Xbit_r122_c226 bl[226] br[226] wl[122] vdd gnd cell_6t
Xbit_r123_c226 bl[226] br[226] wl[123] vdd gnd cell_6t
Xbit_r124_c226 bl[226] br[226] wl[124] vdd gnd cell_6t
Xbit_r125_c226 bl[226] br[226] wl[125] vdd gnd cell_6t
Xbit_r126_c226 bl[226] br[226] wl[126] vdd gnd cell_6t
Xbit_r127_c226 bl[226] br[226] wl[127] vdd gnd cell_6t
Xbit_r0_c227 bl[227] br[227] wl[0] vdd gnd cell_6t
Xbit_r1_c227 bl[227] br[227] wl[1] vdd gnd cell_6t
Xbit_r2_c227 bl[227] br[227] wl[2] vdd gnd cell_6t
Xbit_r3_c227 bl[227] br[227] wl[3] vdd gnd cell_6t
Xbit_r4_c227 bl[227] br[227] wl[4] vdd gnd cell_6t
Xbit_r5_c227 bl[227] br[227] wl[5] vdd gnd cell_6t
Xbit_r6_c227 bl[227] br[227] wl[6] vdd gnd cell_6t
Xbit_r7_c227 bl[227] br[227] wl[7] vdd gnd cell_6t
Xbit_r8_c227 bl[227] br[227] wl[8] vdd gnd cell_6t
Xbit_r9_c227 bl[227] br[227] wl[9] vdd gnd cell_6t
Xbit_r10_c227 bl[227] br[227] wl[10] vdd gnd cell_6t
Xbit_r11_c227 bl[227] br[227] wl[11] vdd gnd cell_6t
Xbit_r12_c227 bl[227] br[227] wl[12] vdd gnd cell_6t
Xbit_r13_c227 bl[227] br[227] wl[13] vdd gnd cell_6t
Xbit_r14_c227 bl[227] br[227] wl[14] vdd gnd cell_6t
Xbit_r15_c227 bl[227] br[227] wl[15] vdd gnd cell_6t
Xbit_r16_c227 bl[227] br[227] wl[16] vdd gnd cell_6t
Xbit_r17_c227 bl[227] br[227] wl[17] vdd gnd cell_6t
Xbit_r18_c227 bl[227] br[227] wl[18] vdd gnd cell_6t
Xbit_r19_c227 bl[227] br[227] wl[19] vdd gnd cell_6t
Xbit_r20_c227 bl[227] br[227] wl[20] vdd gnd cell_6t
Xbit_r21_c227 bl[227] br[227] wl[21] vdd gnd cell_6t
Xbit_r22_c227 bl[227] br[227] wl[22] vdd gnd cell_6t
Xbit_r23_c227 bl[227] br[227] wl[23] vdd gnd cell_6t
Xbit_r24_c227 bl[227] br[227] wl[24] vdd gnd cell_6t
Xbit_r25_c227 bl[227] br[227] wl[25] vdd gnd cell_6t
Xbit_r26_c227 bl[227] br[227] wl[26] vdd gnd cell_6t
Xbit_r27_c227 bl[227] br[227] wl[27] vdd gnd cell_6t
Xbit_r28_c227 bl[227] br[227] wl[28] vdd gnd cell_6t
Xbit_r29_c227 bl[227] br[227] wl[29] vdd gnd cell_6t
Xbit_r30_c227 bl[227] br[227] wl[30] vdd gnd cell_6t
Xbit_r31_c227 bl[227] br[227] wl[31] vdd gnd cell_6t
Xbit_r32_c227 bl[227] br[227] wl[32] vdd gnd cell_6t
Xbit_r33_c227 bl[227] br[227] wl[33] vdd gnd cell_6t
Xbit_r34_c227 bl[227] br[227] wl[34] vdd gnd cell_6t
Xbit_r35_c227 bl[227] br[227] wl[35] vdd gnd cell_6t
Xbit_r36_c227 bl[227] br[227] wl[36] vdd gnd cell_6t
Xbit_r37_c227 bl[227] br[227] wl[37] vdd gnd cell_6t
Xbit_r38_c227 bl[227] br[227] wl[38] vdd gnd cell_6t
Xbit_r39_c227 bl[227] br[227] wl[39] vdd gnd cell_6t
Xbit_r40_c227 bl[227] br[227] wl[40] vdd gnd cell_6t
Xbit_r41_c227 bl[227] br[227] wl[41] vdd gnd cell_6t
Xbit_r42_c227 bl[227] br[227] wl[42] vdd gnd cell_6t
Xbit_r43_c227 bl[227] br[227] wl[43] vdd gnd cell_6t
Xbit_r44_c227 bl[227] br[227] wl[44] vdd gnd cell_6t
Xbit_r45_c227 bl[227] br[227] wl[45] vdd gnd cell_6t
Xbit_r46_c227 bl[227] br[227] wl[46] vdd gnd cell_6t
Xbit_r47_c227 bl[227] br[227] wl[47] vdd gnd cell_6t
Xbit_r48_c227 bl[227] br[227] wl[48] vdd gnd cell_6t
Xbit_r49_c227 bl[227] br[227] wl[49] vdd gnd cell_6t
Xbit_r50_c227 bl[227] br[227] wl[50] vdd gnd cell_6t
Xbit_r51_c227 bl[227] br[227] wl[51] vdd gnd cell_6t
Xbit_r52_c227 bl[227] br[227] wl[52] vdd gnd cell_6t
Xbit_r53_c227 bl[227] br[227] wl[53] vdd gnd cell_6t
Xbit_r54_c227 bl[227] br[227] wl[54] vdd gnd cell_6t
Xbit_r55_c227 bl[227] br[227] wl[55] vdd gnd cell_6t
Xbit_r56_c227 bl[227] br[227] wl[56] vdd gnd cell_6t
Xbit_r57_c227 bl[227] br[227] wl[57] vdd gnd cell_6t
Xbit_r58_c227 bl[227] br[227] wl[58] vdd gnd cell_6t
Xbit_r59_c227 bl[227] br[227] wl[59] vdd gnd cell_6t
Xbit_r60_c227 bl[227] br[227] wl[60] vdd gnd cell_6t
Xbit_r61_c227 bl[227] br[227] wl[61] vdd gnd cell_6t
Xbit_r62_c227 bl[227] br[227] wl[62] vdd gnd cell_6t
Xbit_r63_c227 bl[227] br[227] wl[63] vdd gnd cell_6t
Xbit_r64_c227 bl[227] br[227] wl[64] vdd gnd cell_6t
Xbit_r65_c227 bl[227] br[227] wl[65] vdd gnd cell_6t
Xbit_r66_c227 bl[227] br[227] wl[66] vdd gnd cell_6t
Xbit_r67_c227 bl[227] br[227] wl[67] vdd gnd cell_6t
Xbit_r68_c227 bl[227] br[227] wl[68] vdd gnd cell_6t
Xbit_r69_c227 bl[227] br[227] wl[69] vdd gnd cell_6t
Xbit_r70_c227 bl[227] br[227] wl[70] vdd gnd cell_6t
Xbit_r71_c227 bl[227] br[227] wl[71] vdd gnd cell_6t
Xbit_r72_c227 bl[227] br[227] wl[72] vdd gnd cell_6t
Xbit_r73_c227 bl[227] br[227] wl[73] vdd gnd cell_6t
Xbit_r74_c227 bl[227] br[227] wl[74] vdd gnd cell_6t
Xbit_r75_c227 bl[227] br[227] wl[75] vdd gnd cell_6t
Xbit_r76_c227 bl[227] br[227] wl[76] vdd gnd cell_6t
Xbit_r77_c227 bl[227] br[227] wl[77] vdd gnd cell_6t
Xbit_r78_c227 bl[227] br[227] wl[78] vdd gnd cell_6t
Xbit_r79_c227 bl[227] br[227] wl[79] vdd gnd cell_6t
Xbit_r80_c227 bl[227] br[227] wl[80] vdd gnd cell_6t
Xbit_r81_c227 bl[227] br[227] wl[81] vdd gnd cell_6t
Xbit_r82_c227 bl[227] br[227] wl[82] vdd gnd cell_6t
Xbit_r83_c227 bl[227] br[227] wl[83] vdd gnd cell_6t
Xbit_r84_c227 bl[227] br[227] wl[84] vdd gnd cell_6t
Xbit_r85_c227 bl[227] br[227] wl[85] vdd gnd cell_6t
Xbit_r86_c227 bl[227] br[227] wl[86] vdd gnd cell_6t
Xbit_r87_c227 bl[227] br[227] wl[87] vdd gnd cell_6t
Xbit_r88_c227 bl[227] br[227] wl[88] vdd gnd cell_6t
Xbit_r89_c227 bl[227] br[227] wl[89] vdd gnd cell_6t
Xbit_r90_c227 bl[227] br[227] wl[90] vdd gnd cell_6t
Xbit_r91_c227 bl[227] br[227] wl[91] vdd gnd cell_6t
Xbit_r92_c227 bl[227] br[227] wl[92] vdd gnd cell_6t
Xbit_r93_c227 bl[227] br[227] wl[93] vdd gnd cell_6t
Xbit_r94_c227 bl[227] br[227] wl[94] vdd gnd cell_6t
Xbit_r95_c227 bl[227] br[227] wl[95] vdd gnd cell_6t
Xbit_r96_c227 bl[227] br[227] wl[96] vdd gnd cell_6t
Xbit_r97_c227 bl[227] br[227] wl[97] vdd gnd cell_6t
Xbit_r98_c227 bl[227] br[227] wl[98] vdd gnd cell_6t
Xbit_r99_c227 bl[227] br[227] wl[99] vdd gnd cell_6t
Xbit_r100_c227 bl[227] br[227] wl[100] vdd gnd cell_6t
Xbit_r101_c227 bl[227] br[227] wl[101] vdd gnd cell_6t
Xbit_r102_c227 bl[227] br[227] wl[102] vdd gnd cell_6t
Xbit_r103_c227 bl[227] br[227] wl[103] vdd gnd cell_6t
Xbit_r104_c227 bl[227] br[227] wl[104] vdd gnd cell_6t
Xbit_r105_c227 bl[227] br[227] wl[105] vdd gnd cell_6t
Xbit_r106_c227 bl[227] br[227] wl[106] vdd gnd cell_6t
Xbit_r107_c227 bl[227] br[227] wl[107] vdd gnd cell_6t
Xbit_r108_c227 bl[227] br[227] wl[108] vdd gnd cell_6t
Xbit_r109_c227 bl[227] br[227] wl[109] vdd gnd cell_6t
Xbit_r110_c227 bl[227] br[227] wl[110] vdd gnd cell_6t
Xbit_r111_c227 bl[227] br[227] wl[111] vdd gnd cell_6t
Xbit_r112_c227 bl[227] br[227] wl[112] vdd gnd cell_6t
Xbit_r113_c227 bl[227] br[227] wl[113] vdd gnd cell_6t
Xbit_r114_c227 bl[227] br[227] wl[114] vdd gnd cell_6t
Xbit_r115_c227 bl[227] br[227] wl[115] vdd gnd cell_6t
Xbit_r116_c227 bl[227] br[227] wl[116] vdd gnd cell_6t
Xbit_r117_c227 bl[227] br[227] wl[117] vdd gnd cell_6t
Xbit_r118_c227 bl[227] br[227] wl[118] vdd gnd cell_6t
Xbit_r119_c227 bl[227] br[227] wl[119] vdd gnd cell_6t
Xbit_r120_c227 bl[227] br[227] wl[120] vdd gnd cell_6t
Xbit_r121_c227 bl[227] br[227] wl[121] vdd gnd cell_6t
Xbit_r122_c227 bl[227] br[227] wl[122] vdd gnd cell_6t
Xbit_r123_c227 bl[227] br[227] wl[123] vdd gnd cell_6t
Xbit_r124_c227 bl[227] br[227] wl[124] vdd gnd cell_6t
Xbit_r125_c227 bl[227] br[227] wl[125] vdd gnd cell_6t
Xbit_r126_c227 bl[227] br[227] wl[126] vdd gnd cell_6t
Xbit_r127_c227 bl[227] br[227] wl[127] vdd gnd cell_6t
Xbit_r0_c228 bl[228] br[228] wl[0] vdd gnd cell_6t
Xbit_r1_c228 bl[228] br[228] wl[1] vdd gnd cell_6t
Xbit_r2_c228 bl[228] br[228] wl[2] vdd gnd cell_6t
Xbit_r3_c228 bl[228] br[228] wl[3] vdd gnd cell_6t
Xbit_r4_c228 bl[228] br[228] wl[4] vdd gnd cell_6t
Xbit_r5_c228 bl[228] br[228] wl[5] vdd gnd cell_6t
Xbit_r6_c228 bl[228] br[228] wl[6] vdd gnd cell_6t
Xbit_r7_c228 bl[228] br[228] wl[7] vdd gnd cell_6t
Xbit_r8_c228 bl[228] br[228] wl[8] vdd gnd cell_6t
Xbit_r9_c228 bl[228] br[228] wl[9] vdd gnd cell_6t
Xbit_r10_c228 bl[228] br[228] wl[10] vdd gnd cell_6t
Xbit_r11_c228 bl[228] br[228] wl[11] vdd gnd cell_6t
Xbit_r12_c228 bl[228] br[228] wl[12] vdd gnd cell_6t
Xbit_r13_c228 bl[228] br[228] wl[13] vdd gnd cell_6t
Xbit_r14_c228 bl[228] br[228] wl[14] vdd gnd cell_6t
Xbit_r15_c228 bl[228] br[228] wl[15] vdd gnd cell_6t
Xbit_r16_c228 bl[228] br[228] wl[16] vdd gnd cell_6t
Xbit_r17_c228 bl[228] br[228] wl[17] vdd gnd cell_6t
Xbit_r18_c228 bl[228] br[228] wl[18] vdd gnd cell_6t
Xbit_r19_c228 bl[228] br[228] wl[19] vdd gnd cell_6t
Xbit_r20_c228 bl[228] br[228] wl[20] vdd gnd cell_6t
Xbit_r21_c228 bl[228] br[228] wl[21] vdd gnd cell_6t
Xbit_r22_c228 bl[228] br[228] wl[22] vdd gnd cell_6t
Xbit_r23_c228 bl[228] br[228] wl[23] vdd gnd cell_6t
Xbit_r24_c228 bl[228] br[228] wl[24] vdd gnd cell_6t
Xbit_r25_c228 bl[228] br[228] wl[25] vdd gnd cell_6t
Xbit_r26_c228 bl[228] br[228] wl[26] vdd gnd cell_6t
Xbit_r27_c228 bl[228] br[228] wl[27] vdd gnd cell_6t
Xbit_r28_c228 bl[228] br[228] wl[28] vdd gnd cell_6t
Xbit_r29_c228 bl[228] br[228] wl[29] vdd gnd cell_6t
Xbit_r30_c228 bl[228] br[228] wl[30] vdd gnd cell_6t
Xbit_r31_c228 bl[228] br[228] wl[31] vdd gnd cell_6t
Xbit_r32_c228 bl[228] br[228] wl[32] vdd gnd cell_6t
Xbit_r33_c228 bl[228] br[228] wl[33] vdd gnd cell_6t
Xbit_r34_c228 bl[228] br[228] wl[34] vdd gnd cell_6t
Xbit_r35_c228 bl[228] br[228] wl[35] vdd gnd cell_6t
Xbit_r36_c228 bl[228] br[228] wl[36] vdd gnd cell_6t
Xbit_r37_c228 bl[228] br[228] wl[37] vdd gnd cell_6t
Xbit_r38_c228 bl[228] br[228] wl[38] vdd gnd cell_6t
Xbit_r39_c228 bl[228] br[228] wl[39] vdd gnd cell_6t
Xbit_r40_c228 bl[228] br[228] wl[40] vdd gnd cell_6t
Xbit_r41_c228 bl[228] br[228] wl[41] vdd gnd cell_6t
Xbit_r42_c228 bl[228] br[228] wl[42] vdd gnd cell_6t
Xbit_r43_c228 bl[228] br[228] wl[43] vdd gnd cell_6t
Xbit_r44_c228 bl[228] br[228] wl[44] vdd gnd cell_6t
Xbit_r45_c228 bl[228] br[228] wl[45] vdd gnd cell_6t
Xbit_r46_c228 bl[228] br[228] wl[46] vdd gnd cell_6t
Xbit_r47_c228 bl[228] br[228] wl[47] vdd gnd cell_6t
Xbit_r48_c228 bl[228] br[228] wl[48] vdd gnd cell_6t
Xbit_r49_c228 bl[228] br[228] wl[49] vdd gnd cell_6t
Xbit_r50_c228 bl[228] br[228] wl[50] vdd gnd cell_6t
Xbit_r51_c228 bl[228] br[228] wl[51] vdd gnd cell_6t
Xbit_r52_c228 bl[228] br[228] wl[52] vdd gnd cell_6t
Xbit_r53_c228 bl[228] br[228] wl[53] vdd gnd cell_6t
Xbit_r54_c228 bl[228] br[228] wl[54] vdd gnd cell_6t
Xbit_r55_c228 bl[228] br[228] wl[55] vdd gnd cell_6t
Xbit_r56_c228 bl[228] br[228] wl[56] vdd gnd cell_6t
Xbit_r57_c228 bl[228] br[228] wl[57] vdd gnd cell_6t
Xbit_r58_c228 bl[228] br[228] wl[58] vdd gnd cell_6t
Xbit_r59_c228 bl[228] br[228] wl[59] vdd gnd cell_6t
Xbit_r60_c228 bl[228] br[228] wl[60] vdd gnd cell_6t
Xbit_r61_c228 bl[228] br[228] wl[61] vdd gnd cell_6t
Xbit_r62_c228 bl[228] br[228] wl[62] vdd gnd cell_6t
Xbit_r63_c228 bl[228] br[228] wl[63] vdd gnd cell_6t
Xbit_r64_c228 bl[228] br[228] wl[64] vdd gnd cell_6t
Xbit_r65_c228 bl[228] br[228] wl[65] vdd gnd cell_6t
Xbit_r66_c228 bl[228] br[228] wl[66] vdd gnd cell_6t
Xbit_r67_c228 bl[228] br[228] wl[67] vdd gnd cell_6t
Xbit_r68_c228 bl[228] br[228] wl[68] vdd gnd cell_6t
Xbit_r69_c228 bl[228] br[228] wl[69] vdd gnd cell_6t
Xbit_r70_c228 bl[228] br[228] wl[70] vdd gnd cell_6t
Xbit_r71_c228 bl[228] br[228] wl[71] vdd gnd cell_6t
Xbit_r72_c228 bl[228] br[228] wl[72] vdd gnd cell_6t
Xbit_r73_c228 bl[228] br[228] wl[73] vdd gnd cell_6t
Xbit_r74_c228 bl[228] br[228] wl[74] vdd gnd cell_6t
Xbit_r75_c228 bl[228] br[228] wl[75] vdd gnd cell_6t
Xbit_r76_c228 bl[228] br[228] wl[76] vdd gnd cell_6t
Xbit_r77_c228 bl[228] br[228] wl[77] vdd gnd cell_6t
Xbit_r78_c228 bl[228] br[228] wl[78] vdd gnd cell_6t
Xbit_r79_c228 bl[228] br[228] wl[79] vdd gnd cell_6t
Xbit_r80_c228 bl[228] br[228] wl[80] vdd gnd cell_6t
Xbit_r81_c228 bl[228] br[228] wl[81] vdd gnd cell_6t
Xbit_r82_c228 bl[228] br[228] wl[82] vdd gnd cell_6t
Xbit_r83_c228 bl[228] br[228] wl[83] vdd gnd cell_6t
Xbit_r84_c228 bl[228] br[228] wl[84] vdd gnd cell_6t
Xbit_r85_c228 bl[228] br[228] wl[85] vdd gnd cell_6t
Xbit_r86_c228 bl[228] br[228] wl[86] vdd gnd cell_6t
Xbit_r87_c228 bl[228] br[228] wl[87] vdd gnd cell_6t
Xbit_r88_c228 bl[228] br[228] wl[88] vdd gnd cell_6t
Xbit_r89_c228 bl[228] br[228] wl[89] vdd gnd cell_6t
Xbit_r90_c228 bl[228] br[228] wl[90] vdd gnd cell_6t
Xbit_r91_c228 bl[228] br[228] wl[91] vdd gnd cell_6t
Xbit_r92_c228 bl[228] br[228] wl[92] vdd gnd cell_6t
Xbit_r93_c228 bl[228] br[228] wl[93] vdd gnd cell_6t
Xbit_r94_c228 bl[228] br[228] wl[94] vdd gnd cell_6t
Xbit_r95_c228 bl[228] br[228] wl[95] vdd gnd cell_6t
Xbit_r96_c228 bl[228] br[228] wl[96] vdd gnd cell_6t
Xbit_r97_c228 bl[228] br[228] wl[97] vdd gnd cell_6t
Xbit_r98_c228 bl[228] br[228] wl[98] vdd gnd cell_6t
Xbit_r99_c228 bl[228] br[228] wl[99] vdd gnd cell_6t
Xbit_r100_c228 bl[228] br[228] wl[100] vdd gnd cell_6t
Xbit_r101_c228 bl[228] br[228] wl[101] vdd gnd cell_6t
Xbit_r102_c228 bl[228] br[228] wl[102] vdd gnd cell_6t
Xbit_r103_c228 bl[228] br[228] wl[103] vdd gnd cell_6t
Xbit_r104_c228 bl[228] br[228] wl[104] vdd gnd cell_6t
Xbit_r105_c228 bl[228] br[228] wl[105] vdd gnd cell_6t
Xbit_r106_c228 bl[228] br[228] wl[106] vdd gnd cell_6t
Xbit_r107_c228 bl[228] br[228] wl[107] vdd gnd cell_6t
Xbit_r108_c228 bl[228] br[228] wl[108] vdd gnd cell_6t
Xbit_r109_c228 bl[228] br[228] wl[109] vdd gnd cell_6t
Xbit_r110_c228 bl[228] br[228] wl[110] vdd gnd cell_6t
Xbit_r111_c228 bl[228] br[228] wl[111] vdd gnd cell_6t
Xbit_r112_c228 bl[228] br[228] wl[112] vdd gnd cell_6t
Xbit_r113_c228 bl[228] br[228] wl[113] vdd gnd cell_6t
Xbit_r114_c228 bl[228] br[228] wl[114] vdd gnd cell_6t
Xbit_r115_c228 bl[228] br[228] wl[115] vdd gnd cell_6t
Xbit_r116_c228 bl[228] br[228] wl[116] vdd gnd cell_6t
Xbit_r117_c228 bl[228] br[228] wl[117] vdd gnd cell_6t
Xbit_r118_c228 bl[228] br[228] wl[118] vdd gnd cell_6t
Xbit_r119_c228 bl[228] br[228] wl[119] vdd gnd cell_6t
Xbit_r120_c228 bl[228] br[228] wl[120] vdd gnd cell_6t
Xbit_r121_c228 bl[228] br[228] wl[121] vdd gnd cell_6t
Xbit_r122_c228 bl[228] br[228] wl[122] vdd gnd cell_6t
Xbit_r123_c228 bl[228] br[228] wl[123] vdd gnd cell_6t
Xbit_r124_c228 bl[228] br[228] wl[124] vdd gnd cell_6t
Xbit_r125_c228 bl[228] br[228] wl[125] vdd gnd cell_6t
Xbit_r126_c228 bl[228] br[228] wl[126] vdd gnd cell_6t
Xbit_r127_c228 bl[228] br[228] wl[127] vdd gnd cell_6t
Xbit_r0_c229 bl[229] br[229] wl[0] vdd gnd cell_6t
Xbit_r1_c229 bl[229] br[229] wl[1] vdd gnd cell_6t
Xbit_r2_c229 bl[229] br[229] wl[2] vdd gnd cell_6t
Xbit_r3_c229 bl[229] br[229] wl[3] vdd gnd cell_6t
Xbit_r4_c229 bl[229] br[229] wl[4] vdd gnd cell_6t
Xbit_r5_c229 bl[229] br[229] wl[5] vdd gnd cell_6t
Xbit_r6_c229 bl[229] br[229] wl[6] vdd gnd cell_6t
Xbit_r7_c229 bl[229] br[229] wl[7] vdd gnd cell_6t
Xbit_r8_c229 bl[229] br[229] wl[8] vdd gnd cell_6t
Xbit_r9_c229 bl[229] br[229] wl[9] vdd gnd cell_6t
Xbit_r10_c229 bl[229] br[229] wl[10] vdd gnd cell_6t
Xbit_r11_c229 bl[229] br[229] wl[11] vdd gnd cell_6t
Xbit_r12_c229 bl[229] br[229] wl[12] vdd gnd cell_6t
Xbit_r13_c229 bl[229] br[229] wl[13] vdd gnd cell_6t
Xbit_r14_c229 bl[229] br[229] wl[14] vdd gnd cell_6t
Xbit_r15_c229 bl[229] br[229] wl[15] vdd gnd cell_6t
Xbit_r16_c229 bl[229] br[229] wl[16] vdd gnd cell_6t
Xbit_r17_c229 bl[229] br[229] wl[17] vdd gnd cell_6t
Xbit_r18_c229 bl[229] br[229] wl[18] vdd gnd cell_6t
Xbit_r19_c229 bl[229] br[229] wl[19] vdd gnd cell_6t
Xbit_r20_c229 bl[229] br[229] wl[20] vdd gnd cell_6t
Xbit_r21_c229 bl[229] br[229] wl[21] vdd gnd cell_6t
Xbit_r22_c229 bl[229] br[229] wl[22] vdd gnd cell_6t
Xbit_r23_c229 bl[229] br[229] wl[23] vdd gnd cell_6t
Xbit_r24_c229 bl[229] br[229] wl[24] vdd gnd cell_6t
Xbit_r25_c229 bl[229] br[229] wl[25] vdd gnd cell_6t
Xbit_r26_c229 bl[229] br[229] wl[26] vdd gnd cell_6t
Xbit_r27_c229 bl[229] br[229] wl[27] vdd gnd cell_6t
Xbit_r28_c229 bl[229] br[229] wl[28] vdd gnd cell_6t
Xbit_r29_c229 bl[229] br[229] wl[29] vdd gnd cell_6t
Xbit_r30_c229 bl[229] br[229] wl[30] vdd gnd cell_6t
Xbit_r31_c229 bl[229] br[229] wl[31] vdd gnd cell_6t
Xbit_r32_c229 bl[229] br[229] wl[32] vdd gnd cell_6t
Xbit_r33_c229 bl[229] br[229] wl[33] vdd gnd cell_6t
Xbit_r34_c229 bl[229] br[229] wl[34] vdd gnd cell_6t
Xbit_r35_c229 bl[229] br[229] wl[35] vdd gnd cell_6t
Xbit_r36_c229 bl[229] br[229] wl[36] vdd gnd cell_6t
Xbit_r37_c229 bl[229] br[229] wl[37] vdd gnd cell_6t
Xbit_r38_c229 bl[229] br[229] wl[38] vdd gnd cell_6t
Xbit_r39_c229 bl[229] br[229] wl[39] vdd gnd cell_6t
Xbit_r40_c229 bl[229] br[229] wl[40] vdd gnd cell_6t
Xbit_r41_c229 bl[229] br[229] wl[41] vdd gnd cell_6t
Xbit_r42_c229 bl[229] br[229] wl[42] vdd gnd cell_6t
Xbit_r43_c229 bl[229] br[229] wl[43] vdd gnd cell_6t
Xbit_r44_c229 bl[229] br[229] wl[44] vdd gnd cell_6t
Xbit_r45_c229 bl[229] br[229] wl[45] vdd gnd cell_6t
Xbit_r46_c229 bl[229] br[229] wl[46] vdd gnd cell_6t
Xbit_r47_c229 bl[229] br[229] wl[47] vdd gnd cell_6t
Xbit_r48_c229 bl[229] br[229] wl[48] vdd gnd cell_6t
Xbit_r49_c229 bl[229] br[229] wl[49] vdd gnd cell_6t
Xbit_r50_c229 bl[229] br[229] wl[50] vdd gnd cell_6t
Xbit_r51_c229 bl[229] br[229] wl[51] vdd gnd cell_6t
Xbit_r52_c229 bl[229] br[229] wl[52] vdd gnd cell_6t
Xbit_r53_c229 bl[229] br[229] wl[53] vdd gnd cell_6t
Xbit_r54_c229 bl[229] br[229] wl[54] vdd gnd cell_6t
Xbit_r55_c229 bl[229] br[229] wl[55] vdd gnd cell_6t
Xbit_r56_c229 bl[229] br[229] wl[56] vdd gnd cell_6t
Xbit_r57_c229 bl[229] br[229] wl[57] vdd gnd cell_6t
Xbit_r58_c229 bl[229] br[229] wl[58] vdd gnd cell_6t
Xbit_r59_c229 bl[229] br[229] wl[59] vdd gnd cell_6t
Xbit_r60_c229 bl[229] br[229] wl[60] vdd gnd cell_6t
Xbit_r61_c229 bl[229] br[229] wl[61] vdd gnd cell_6t
Xbit_r62_c229 bl[229] br[229] wl[62] vdd gnd cell_6t
Xbit_r63_c229 bl[229] br[229] wl[63] vdd gnd cell_6t
Xbit_r64_c229 bl[229] br[229] wl[64] vdd gnd cell_6t
Xbit_r65_c229 bl[229] br[229] wl[65] vdd gnd cell_6t
Xbit_r66_c229 bl[229] br[229] wl[66] vdd gnd cell_6t
Xbit_r67_c229 bl[229] br[229] wl[67] vdd gnd cell_6t
Xbit_r68_c229 bl[229] br[229] wl[68] vdd gnd cell_6t
Xbit_r69_c229 bl[229] br[229] wl[69] vdd gnd cell_6t
Xbit_r70_c229 bl[229] br[229] wl[70] vdd gnd cell_6t
Xbit_r71_c229 bl[229] br[229] wl[71] vdd gnd cell_6t
Xbit_r72_c229 bl[229] br[229] wl[72] vdd gnd cell_6t
Xbit_r73_c229 bl[229] br[229] wl[73] vdd gnd cell_6t
Xbit_r74_c229 bl[229] br[229] wl[74] vdd gnd cell_6t
Xbit_r75_c229 bl[229] br[229] wl[75] vdd gnd cell_6t
Xbit_r76_c229 bl[229] br[229] wl[76] vdd gnd cell_6t
Xbit_r77_c229 bl[229] br[229] wl[77] vdd gnd cell_6t
Xbit_r78_c229 bl[229] br[229] wl[78] vdd gnd cell_6t
Xbit_r79_c229 bl[229] br[229] wl[79] vdd gnd cell_6t
Xbit_r80_c229 bl[229] br[229] wl[80] vdd gnd cell_6t
Xbit_r81_c229 bl[229] br[229] wl[81] vdd gnd cell_6t
Xbit_r82_c229 bl[229] br[229] wl[82] vdd gnd cell_6t
Xbit_r83_c229 bl[229] br[229] wl[83] vdd gnd cell_6t
Xbit_r84_c229 bl[229] br[229] wl[84] vdd gnd cell_6t
Xbit_r85_c229 bl[229] br[229] wl[85] vdd gnd cell_6t
Xbit_r86_c229 bl[229] br[229] wl[86] vdd gnd cell_6t
Xbit_r87_c229 bl[229] br[229] wl[87] vdd gnd cell_6t
Xbit_r88_c229 bl[229] br[229] wl[88] vdd gnd cell_6t
Xbit_r89_c229 bl[229] br[229] wl[89] vdd gnd cell_6t
Xbit_r90_c229 bl[229] br[229] wl[90] vdd gnd cell_6t
Xbit_r91_c229 bl[229] br[229] wl[91] vdd gnd cell_6t
Xbit_r92_c229 bl[229] br[229] wl[92] vdd gnd cell_6t
Xbit_r93_c229 bl[229] br[229] wl[93] vdd gnd cell_6t
Xbit_r94_c229 bl[229] br[229] wl[94] vdd gnd cell_6t
Xbit_r95_c229 bl[229] br[229] wl[95] vdd gnd cell_6t
Xbit_r96_c229 bl[229] br[229] wl[96] vdd gnd cell_6t
Xbit_r97_c229 bl[229] br[229] wl[97] vdd gnd cell_6t
Xbit_r98_c229 bl[229] br[229] wl[98] vdd gnd cell_6t
Xbit_r99_c229 bl[229] br[229] wl[99] vdd gnd cell_6t
Xbit_r100_c229 bl[229] br[229] wl[100] vdd gnd cell_6t
Xbit_r101_c229 bl[229] br[229] wl[101] vdd gnd cell_6t
Xbit_r102_c229 bl[229] br[229] wl[102] vdd gnd cell_6t
Xbit_r103_c229 bl[229] br[229] wl[103] vdd gnd cell_6t
Xbit_r104_c229 bl[229] br[229] wl[104] vdd gnd cell_6t
Xbit_r105_c229 bl[229] br[229] wl[105] vdd gnd cell_6t
Xbit_r106_c229 bl[229] br[229] wl[106] vdd gnd cell_6t
Xbit_r107_c229 bl[229] br[229] wl[107] vdd gnd cell_6t
Xbit_r108_c229 bl[229] br[229] wl[108] vdd gnd cell_6t
Xbit_r109_c229 bl[229] br[229] wl[109] vdd gnd cell_6t
Xbit_r110_c229 bl[229] br[229] wl[110] vdd gnd cell_6t
Xbit_r111_c229 bl[229] br[229] wl[111] vdd gnd cell_6t
Xbit_r112_c229 bl[229] br[229] wl[112] vdd gnd cell_6t
Xbit_r113_c229 bl[229] br[229] wl[113] vdd gnd cell_6t
Xbit_r114_c229 bl[229] br[229] wl[114] vdd gnd cell_6t
Xbit_r115_c229 bl[229] br[229] wl[115] vdd gnd cell_6t
Xbit_r116_c229 bl[229] br[229] wl[116] vdd gnd cell_6t
Xbit_r117_c229 bl[229] br[229] wl[117] vdd gnd cell_6t
Xbit_r118_c229 bl[229] br[229] wl[118] vdd gnd cell_6t
Xbit_r119_c229 bl[229] br[229] wl[119] vdd gnd cell_6t
Xbit_r120_c229 bl[229] br[229] wl[120] vdd gnd cell_6t
Xbit_r121_c229 bl[229] br[229] wl[121] vdd gnd cell_6t
Xbit_r122_c229 bl[229] br[229] wl[122] vdd gnd cell_6t
Xbit_r123_c229 bl[229] br[229] wl[123] vdd gnd cell_6t
Xbit_r124_c229 bl[229] br[229] wl[124] vdd gnd cell_6t
Xbit_r125_c229 bl[229] br[229] wl[125] vdd gnd cell_6t
Xbit_r126_c229 bl[229] br[229] wl[126] vdd gnd cell_6t
Xbit_r127_c229 bl[229] br[229] wl[127] vdd gnd cell_6t
Xbit_r0_c230 bl[230] br[230] wl[0] vdd gnd cell_6t
Xbit_r1_c230 bl[230] br[230] wl[1] vdd gnd cell_6t
Xbit_r2_c230 bl[230] br[230] wl[2] vdd gnd cell_6t
Xbit_r3_c230 bl[230] br[230] wl[3] vdd gnd cell_6t
Xbit_r4_c230 bl[230] br[230] wl[4] vdd gnd cell_6t
Xbit_r5_c230 bl[230] br[230] wl[5] vdd gnd cell_6t
Xbit_r6_c230 bl[230] br[230] wl[6] vdd gnd cell_6t
Xbit_r7_c230 bl[230] br[230] wl[7] vdd gnd cell_6t
Xbit_r8_c230 bl[230] br[230] wl[8] vdd gnd cell_6t
Xbit_r9_c230 bl[230] br[230] wl[9] vdd gnd cell_6t
Xbit_r10_c230 bl[230] br[230] wl[10] vdd gnd cell_6t
Xbit_r11_c230 bl[230] br[230] wl[11] vdd gnd cell_6t
Xbit_r12_c230 bl[230] br[230] wl[12] vdd gnd cell_6t
Xbit_r13_c230 bl[230] br[230] wl[13] vdd gnd cell_6t
Xbit_r14_c230 bl[230] br[230] wl[14] vdd gnd cell_6t
Xbit_r15_c230 bl[230] br[230] wl[15] vdd gnd cell_6t
Xbit_r16_c230 bl[230] br[230] wl[16] vdd gnd cell_6t
Xbit_r17_c230 bl[230] br[230] wl[17] vdd gnd cell_6t
Xbit_r18_c230 bl[230] br[230] wl[18] vdd gnd cell_6t
Xbit_r19_c230 bl[230] br[230] wl[19] vdd gnd cell_6t
Xbit_r20_c230 bl[230] br[230] wl[20] vdd gnd cell_6t
Xbit_r21_c230 bl[230] br[230] wl[21] vdd gnd cell_6t
Xbit_r22_c230 bl[230] br[230] wl[22] vdd gnd cell_6t
Xbit_r23_c230 bl[230] br[230] wl[23] vdd gnd cell_6t
Xbit_r24_c230 bl[230] br[230] wl[24] vdd gnd cell_6t
Xbit_r25_c230 bl[230] br[230] wl[25] vdd gnd cell_6t
Xbit_r26_c230 bl[230] br[230] wl[26] vdd gnd cell_6t
Xbit_r27_c230 bl[230] br[230] wl[27] vdd gnd cell_6t
Xbit_r28_c230 bl[230] br[230] wl[28] vdd gnd cell_6t
Xbit_r29_c230 bl[230] br[230] wl[29] vdd gnd cell_6t
Xbit_r30_c230 bl[230] br[230] wl[30] vdd gnd cell_6t
Xbit_r31_c230 bl[230] br[230] wl[31] vdd gnd cell_6t
Xbit_r32_c230 bl[230] br[230] wl[32] vdd gnd cell_6t
Xbit_r33_c230 bl[230] br[230] wl[33] vdd gnd cell_6t
Xbit_r34_c230 bl[230] br[230] wl[34] vdd gnd cell_6t
Xbit_r35_c230 bl[230] br[230] wl[35] vdd gnd cell_6t
Xbit_r36_c230 bl[230] br[230] wl[36] vdd gnd cell_6t
Xbit_r37_c230 bl[230] br[230] wl[37] vdd gnd cell_6t
Xbit_r38_c230 bl[230] br[230] wl[38] vdd gnd cell_6t
Xbit_r39_c230 bl[230] br[230] wl[39] vdd gnd cell_6t
Xbit_r40_c230 bl[230] br[230] wl[40] vdd gnd cell_6t
Xbit_r41_c230 bl[230] br[230] wl[41] vdd gnd cell_6t
Xbit_r42_c230 bl[230] br[230] wl[42] vdd gnd cell_6t
Xbit_r43_c230 bl[230] br[230] wl[43] vdd gnd cell_6t
Xbit_r44_c230 bl[230] br[230] wl[44] vdd gnd cell_6t
Xbit_r45_c230 bl[230] br[230] wl[45] vdd gnd cell_6t
Xbit_r46_c230 bl[230] br[230] wl[46] vdd gnd cell_6t
Xbit_r47_c230 bl[230] br[230] wl[47] vdd gnd cell_6t
Xbit_r48_c230 bl[230] br[230] wl[48] vdd gnd cell_6t
Xbit_r49_c230 bl[230] br[230] wl[49] vdd gnd cell_6t
Xbit_r50_c230 bl[230] br[230] wl[50] vdd gnd cell_6t
Xbit_r51_c230 bl[230] br[230] wl[51] vdd gnd cell_6t
Xbit_r52_c230 bl[230] br[230] wl[52] vdd gnd cell_6t
Xbit_r53_c230 bl[230] br[230] wl[53] vdd gnd cell_6t
Xbit_r54_c230 bl[230] br[230] wl[54] vdd gnd cell_6t
Xbit_r55_c230 bl[230] br[230] wl[55] vdd gnd cell_6t
Xbit_r56_c230 bl[230] br[230] wl[56] vdd gnd cell_6t
Xbit_r57_c230 bl[230] br[230] wl[57] vdd gnd cell_6t
Xbit_r58_c230 bl[230] br[230] wl[58] vdd gnd cell_6t
Xbit_r59_c230 bl[230] br[230] wl[59] vdd gnd cell_6t
Xbit_r60_c230 bl[230] br[230] wl[60] vdd gnd cell_6t
Xbit_r61_c230 bl[230] br[230] wl[61] vdd gnd cell_6t
Xbit_r62_c230 bl[230] br[230] wl[62] vdd gnd cell_6t
Xbit_r63_c230 bl[230] br[230] wl[63] vdd gnd cell_6t
Xbit_r64_c230 bl[230] br[230] wl[64] vdd gnd cell_6t
Xbit_r65_c230 bl[230] br[230] wl[65] vdd gnd cell_6t
Xbit_r66_c230 bl[230] br[230] wl[66] vdd gnd cell_6t
Xbit_r67_c230 bl[230] br[230] wl[67] vdd gnd cell_6t
Xbit_r68_c230 bl[230] br[230] wl[68] vdd gnd cell_6t
Xbit_r69_c230 bl[230] br[230] wl[69] vdd gnd cell_6t
Xbit_r70_c230 bl[230] br[230] wl[70] vdd gnd cell_6t
Xbit_r71_c230 bl[230] br[230] wl[71] vdd gnd cell_6t
Xbit_r72_c230 bl[230] br[230] wl[72] vdd gnd cell_6t
Xbit_r73_c230 bl[230] br[230] wl[73] vdd gnd cell_6t
Xbit_r74_c230 bl[230] br[230] wl[74] vdd gnd cell_6t
Xbit_r75_c230 bl[230] br[230] wl[75] vdd gnd cell_6t
Xbit_r76_c230 bl[230] br[230] wl[76] vdd gnd cell_6t
Xbit_r77_c230 bl[230] br[230] wl[77] vdd gnd cell_6t
Xbit_r78_c230 bl[230] br[230] wl[78] vdd gnd cell_6t
Xbit_r79_c230 bl[230] br[230] wl[79] vdd gnd cell_6t
Xbit_r80_c230 bl[230] br[230] wl[80] vdd gnd cell_6t
Xbit_r81_c230 bl[230] br[230] wl[81] vdd gnd cell_6t
Xbit_r82_c230 bl[230] br[230] wl[82] vdd gnd cell_6t
Xbit_r83_c230 bl[230] br[230] wl[83] vdd gnd cell_6t
Xbit_r84_c230 bl[230] br[230] wl[84] vdd gnd cell_6t
Xbit_r85_c230 bl[230] br[230] wl[85] vdd gnd cell_6t
Xbit_r86_c230 bl[230] br[230] wl[86] vdd gnd cell_6t
Xbit_r87_c230 bl[230] br[230] wl[87] vdd gnd cell_6t
Xbit_r88_c230 bl[230] br[230] wl[88] vdd gnd cell_6t
Xbit_r89_c230 bl[230] br[230] wl[89] vdd gnd cell_6t
Xbit_r90_c230 bl[230] br[230] wl[90] vdd gnd cell_6t
Xbit_r91_c230 bl[230] br[230] wl[91] vdd gnd cell_6t
Xbit_r92_c230 bl[230] br[230] wl[92] vdd gnd cell_6t
Xbit_r93_c230 bl[230] br[230] wl[93] vdd gnd cell_6t
Xbit_r94_c230 bl[230] br[230] wl[94] vdd gnd cell_6t
Xbit_r95_c230 bl[230] br[230] wl[95] vdd gnd cell_6t
Xbit_r96_c230 bl[230] br[230] wl[96] vdd gnd cell_6t
Xbit_r97_c230 bl[230] br[230] wl[97] vdd gnd cell_6t
Xbit_r98_c230 bl[230] br[230] wl[98] vdd gnd cell_6t
Xbit_r99_c230 bl[230] br[230] wl[99] vdd gnd cell_6t
Xbit_r100_c230 bl[230] br[230] wl[100] vdd gnd cell_6t
Xbit_r101_c230 bl[230] br[230] wl[101] vdd gnd cell_6t
Xbit_r102_c230 bl[230] br[230] wl[102] vdd gnd cell_6t
Xbit_r103_c230 bl[230] br[230] wl[103] vdd gnd cell_6t
Xbit_r104_c230 bl[230] br[230] wl[104] vdd gnd cell_6t
Xbit_r105_c230 bl[230] br[230] wl[105] vdd gnd cell_6t
Xbit_r106_c230 bl[230] br[230] wl[106] vdd gnd cell_6t
Xbit_r107_c230 bl[230] br[230] wl[107] vdd gnd cell_6t
Xbit_r108_c230 bl[230] br[230] wl[108] vdd gnd cell_6t
Xbit_r109_c230 bl[230] br[230] wl[109] vdd gnd cell_6t
Xbit_r110_c230 bl[230] br[230] wl[110] vdd gnd cell_6t
Xbit_r111_c230 bl[230] br[230] wl[111] vdd gnd cell_6t
Xbit_r112_c230 bl[230] br[230] wl[112] vdd gnd cell_6t
Xbit_r113_c230 bl[230] br[230] wl[113] vdd gnd cell_6t
Xbit_r114_c230 bl[230] br[230] wl[114] vdd gnd cell_6t
Xbit_r115_c230 bl[230] br[230] wl[115] vdd gnd cell_6t
Xbit_r116_c230 bl[230] br[230] wl[116] vdd gnd cell_6t
Xbit_r117_c230 bl[230] br[230] wl[117] vdd gnd cell_6t
Xbit_r118_c230 bl[230] br[230] wl[118] vdd gnd cell_6t
Xbit_r119_c230 bl[230] br[230] wl[119] vdd gnd cell_6t
Xbit_r120_c230 bl[230] br[230] wl[120] vdd gnd cell_6t
Xbit_r121_c230 bl[230] br[230] wl[121] vdd gnd cell_6t
Xbit_r122_c230 bl[230] br[230] wl[122] vdd gnd cell_6t
Xbit_r123_c230 bl[230] br[230] wl[123] vdd gnd cell_6t
Xbit_r124_c230 bl[230] br[230] wl[124] vdd gnd cell_6t
Xbit_r125_c230 bl[230] br[230] wl[125] vdd gnd cell_6t
Xbit_r126_c230 bl[230] br[230] wl[126] vdd gnd cell_6t
Xbit_r127_c230 bl[230] br[230] wl[127] vdd gnd cell_6t
Xbit_r0_c231 bl[231] br[231] wl[0] vdd gnd cell_6t
Xbit_r1_c231 bl[231] br[231] wl[1] vdd gnd cell_6t
Xbit_r2_c231 bl[231] br[231] wl[2] vdd gnd cell_6t
Xbit_r3_c231 bl[231] br[231] wl[3] vdd gnd cell_6t
Xbit_r4_c231 bl[231] br[231] wl[4] vdd gnd cell_6t
Xbit_r5_c231 bl[231] br[231] wl[5] vdd gnd cell_6t
Xbit_r6_c231 bl[231] br[231] wl[6] vdd gnd cell_6t
Xbit_r7_c231 bl[231] br[231] wl[7] vdd gnd cell_6t
Xbit_r8_c231 bl[231] br[231] wl[8] vdd gnd cell_6t
Xbit_r9_c231 bl[231] br[231] wl[9] vdd gnd cell_6t
Xbit_r10_c231 bl[231] br[231] wl[10] vdd gnd cell_6t
Xbit_r11_c231 bl[231] br[231] wl[11] vdd gnd cell_6t
Xbit_r12_c231 bl[231] br[231] wl[12] vdd gnd cell_6t
Xbit_r13_c231 bl[231] br[231] wl[13] vdd gnd cell_6t
Xbit_r14_c231 bl[231] br[231] wl[14] vdd gnd cell_6t
Xbit_r15_c231 bl[231] br[231] wl[15] vdd gnd cell_6t
Xbit_r16_c231 bl[231] br[231] wl[16] vdd gnd cell_6t
Xbit_r17_c231 bl[231] br[231] wl[17] vdd gnd cell_6t
Xbit_r18_c231 bl[231] br[231] wl[18] vdd gnd cell_6t
Xbit_r19_c231 bl[231] br[231] wl[19] vdd gnd cell_6t
Xbit_r20_c231 bl[231] br[231] wl[20] vdd gnd cell_6t
Xbit_r21_c231 bl[231] br[231] wl[21] vdd gnd cell_6t
Xbit_r22_c231 bl[231] br[231] wl[22] vdd gnd cell_6t
Xbit_r23_c231 bl[231] br[231] wl[23] vdd gnd cell_6t
Xbit_r24_c231 bl[231] br[231] wl[24] vdd gnd cell_6t
Xbit_r25_c231 bl[231] br[231] wl[25] vdd gnd cell_6t
Xbit_r26_c231 bl[231] br[231] wl[26] vdd gnd cell_6t
Xbit_r27_c231 bl[231] br[231] wl[27] vdd gnd cell_6t
Xbit_r28_c231 bl[231] br[231] wl[28] vdd gnd cell_6t
Xbit_r29_c231 bl[231] br[231] wl[29] vdd gnd cell_6t
Xbit_r30_c231 bl[231] br[231] wl[30] vdd gnd cell_6t
Xbit_r31_c231 bl[231] br[231] wl[31] vdd gnd cell_6t
Xbit_r32_c231 bl[231] br[231] wl[32] vdd gnd cell_6t
Xbit_r33_c231 bl[231] br[231] wl[33] vdd gnd cell_6t
Xbit_r34_c231 bl[231] br[231] wl[34] vdd gnd cell_6t
Xbit_r35_c231 bl[231] br[231] wl[35] vdd gnd cell_6t
Xbit_r36_c231 bl[231] br[231] wl[36] vdd gnd cell_6t
Xbit_r37_c231 bl[231] br[231] wl[37] vdd gnd cell_6t
Xbit_r38_c231 bl[231] br[231] wl[38] vdd gnd cell_6t
Xbit_r39_c231 bl[231] br[231] wl[39] vdd gnd cell_6t
Xbit_r40_c231 bl[231] br[231] wl[40] vdd gnd cell_6t
Xbit_r41_c231 bl[231] br[231] wl[41] vdd gnd cell_6t
Xbit_r42_c231 bl[231] br[231] wl[42] vdd gnd cell_6t
Xbit_r43_c231 bl[231] br[231] wl[43] vdd gnd cell_6t
Xbit_r44_c231 bl[231] br[231] wl[44] vdd gnd cell_6t
Xbit_r45_c231 bl[231] br[231] wl[45] vdd gnd cell_6t
Xbit_r46_c231 bl[231] br[231] wl[46] vdd gnd cell_6t
Xbit_r47_c231 bl[231] br[231] wl[47] vdd gnd cell_6t
Xbit_r48_c231 bl[231] br[231] wl[48] vdd gnd cell_6t
Xbit_r49_c231 bl[231] br[231] wl[49] vdd gnd cell_6t
Xbit_r50_c231 bl[231] br[231] wl[50] vdd gnd cell_6t
Xbit_r51_c231 bl[231] br[231] wl[51] vdd gnd cell_6t
Xbit_r52_c231 bl[231] br[231] wl[52] vdd gnd cell_6t
Xbit_r53_c231 bl[231] br[231] wl[53] vdd gnd cell_6t
Xbit_r54_c231 bl[231] br[231] wl[54] vdd gnd cell_6t
Xbit_r55_c231 bl[231] br[231] wl[55] vdd gnd cell_6t
Xbit_r56_c231 bl[231] br[231] wl[56] vdd gnd cell_6t
Xbit_r57_c231 bl[231] br[231] wl[57] vdd gnd cell_6t
Xbit_r58_c231 bl[231] br[231] wl[58] vdd gnd cell_6t
Xbit_r59_c231 bl[231] br[231] wl[59] vdd gnd cell_6t
Xbit_r60_c231 bl[231] br[231] wl[60] vdd gnd cell_6t
Xbit_r61_c231 bl[231] br[231] wl[61] vdd gnd cell_6t
Xbit_r62_c231 bl[231] br[231] wl[62] vdd gnd cell_6t
Xbit_r63_c231 bl[231] br[231] wl[63] vdd gnd cell_6t
Xbit_r64_c231 bl[231] br[231] wl[64] vdd gnd cell_6t
Xbit_r65_c231 bl[231] br[231] wl[65] vdd gnd cell_6t
Xbit_r66_c231 bl[231] br[231] wl[66] vdd gnd cell_6t
Xbit_r67_c231 bl[231] br[231] wl[67] vdd gnd cell_6t
Xbit_r68_c231 bl[231] br[231] wl[68] vdd gnd cell_6t
Xbit_r69_c231 bl[231] br[231] wl[69] vdd gnd cell_6t
Xbit_r70_c231 bl[231] br[231] wl[70] vdd gnd cell_6t
Xbit_r71_c231 bl[231] br[231] wl[71] vdd gnd cell_6t
Xbit_r72_c231 bl[231] br[231] wl[72] vdd gnd cell_6t
Xbit_r73_c231 bl[231] br[231] wl[73] vdd gnd cell_6t
Xbit_r74_c231 bl[231] br[231] wl[74] vdd gnd cell_6t
Xbit_r75_c231 bl[231] br[231] wl[75] vdd gnd cell_6t
Xbit_r76_c231 bl[231] br[231] wl[76] vdd gnd cell_6t
Xbit_r77_c231 bl[231] br[231] wl[77] vdd gnd cell_6t
Xbit_r78_c231 bl[231] br[231] wl[78] vdd gnd cell_6t
Xbit_r79_c231 bl[231] br[231] wl[79] vdd gnd cell_6t
Xbit_r80_c231 bl[231] br[231] wl[80] vdd gnd cell_6t
Xbit_r81_c231 bl[231] br[231] wl[81] vdd gnd cell_6t
Xbit_r82_c231 bl[231] br[231] wl[82] vdd gnd cell_6t
Xbit_r83_c231 bl[231] br[231] wl[83] vdd gnd cell_6t
Xbit_r84_c231 bl[231] br[231] wl[84] vdd gnd cell_6t
Xbit_r85_c231 bl[231] br[231] wl[85] vdd gnd cell_6t
Xbit_r86_c231 bl[231] br[231] wl[86] vdd gnd cell_6t
Xbit_r87_c231 bl[231] br[231] wl[87] vdd gnd cell_6t
Xbit_r88_c231 bl[231] br[231] wl[88] vdd gnd cell_6t
Xbit_r89_c231 bl[231] br[231] wl[89] vdd gnd cell_6t
Xbit_r90_c231 bl[231] br[231] wl[90] vdd gnd cell_6t
Xbit_r91_c231 bl[231] br[231] wl[91] vdd gnd cell_6t
Xbit_r92_c231 bl[231] br[231] wl[92] vdd gnd cell_6t
Xbit_r93_c231 bl[231] br[231] wl[93] vdd gnd cell_6t
Xbit_r94_c231 bl[231] br[231] wl[94] vdd gnd cell_6t
Xbit_r95_c231 bl[231] br[231] wl[95] vdd gnd cell_6t
Xbit_r96_c231 bl[231] br[231] wl[96] vdd gnd cell_6t
Xbit_r97_c231 bl[231] br[231] wl[97] vdd gnd cell_6t
Xbit_r98_c231 bl[231] br[231] wl[98] vdd gnd cell_6t
Xbit_r99_c231 bl[231] br[231] wl[99] vdd gnd cell_6t
Xbit_r100_c231 bl[231] br[231] wl[100] vdd gnd cell_6t
Xbit_r101_c231 bl[231] br[231] wl[101] vdd gnd cell_6t
Xbit_r102_c231 bl[231] br[231] wl[102] vdd gnd cell_6t
Xbit_r103_c231 bl[231] br[231] wl[103] vdd gnd cell_6t
Xbit_r104_c231 bl[231] br[231] wl[104] vdd gnd cell_6t
Xbit_r105_c231 bl[231] br[231] wl[105] vdd gnd cell_6t
Xbit_r106_c231 bl[231] br[231] wl[106] vdd gnd cell_6t
Xbit_r107_c231 bl[231] br[231] wl[107] vdd gnd cell_6t
Xbit_r108_c231 bl[231] br[231] wl[108] vdd gnd cell_6t
Xbit_r109_c231 bl[231] br[231] wl[109] vdd gnd cell_6t
Xbit_r110_c231 bl[231] br[231] wl[110] vdd gnd cell_6t
Xbit_r111_c231 bl[231] br[231] wl[111] vdd gnd cell_6t
Xbit_r112_c231 bl[231] br[231] wl[112] vdd gnd cell_6t
Xbit_r113_c231 bl[231] br[231] wl[113] vdd gnd cell_6t
Xbit_r114_c231 bl[231] br[231] wl[114] vdd gnd cell_6t
Xbit_r115_c231 bl[231] br[231] wl[115] vdd gnd cell_6t
Xbit_r116_c231 bl[231] br[231] wl[116] vdd gnd cell_6t
Xbit_r117_c231 bl[231] br[231] wl[117] vdd gnd cell_6t
Xbit_r118_c231 bl[231] br[231] wl[118] vdd gnd cell_6t
Xbit_r119_c231 bl[231] br[231] wl[119] vdd gnd cell_6t
Xbit_r120_c231 bl[231] br[231] wl[120] vdd gnd cell_6t
Xbit_r121_c231 bl[231] br[231] wl[121] vdd gnd cell_6t
Xbit_r122_c231 bl[231] br[231] wl[122] vdd gnd cell_6t
Xbit_r123_c231 bl[231] br[231] wl[123] vdd gnd cell_6t
Xbit_r124_c231 bl[231] br[231] wl[124] vdd gnd cell_6t
Xbit_r125_c231 bl[231] br[231] wl[125] vdd gnd cell_6t
Xbit_r126_c231 bl[231] br[231] wl[126] vdd gnd cell_6t
Xbit_r127_c231 bl[231] br[231] wl[127] vdd gnd cell_6t
Xbit_r0_c232 bl[232] br[232] wl[0] vdd gnd cell_6t
Xbit_r1_c232 bl[232] br[232] wl[1] vdd gnd cell_6t
Xbit_r2_c232 bl[232] br[232] wl[2] vdd gnd cell_6t
Xbit_r3_c232 bl[232] br[232] wl[3] vdd gnd cell_6t
Xbit_r4_c232 bl[232] br[232] wl[4] vdd gnd cell_6t
Xbit_r5_c232 bl[232] br[232] wl[5] vdd gnd cell_6t
Xbit_r6_c232 bl[232] br[232] wl[6] vdd gnd cell_6t
Xbit_r7_c232 bl[232] br[232] wl[7] vdd gnd cell_6t
Xbit_r8_c232 bl[232] br[232] wl[8] vdd gnd cell_6t
Xbit_r9_c232 bl[232] br[232] wl[9] vdd gnd cell_6t
Xbit_r10_c232 bl[232] br[232] wl[10] vdd gnd cell_6t
Xbit_r11_c232 bl[232] br[232] wl[11] vdd gnd cell_6t
Xbit_r12_c232 bl[232] br[232] wl[12] vdd gnd cell_6t
Xbit_r13_c232 bl[232] br[232] wl[13] vdd gnd cell_6t
Xbit_r14_c232 bl[232] br[232] wl[14] vdd gnd cell_6t
Xbit_r15_c232 bl[232] br[232] wl[15] vdd gnd cell_6t
Xbit_r16_c232 bl[232] br[232] wl[16] vdd gnd cell_6t
Xbit_r17_c232 bl[232] br[232] wl[17] vdd gnd cell_6t
Xbit_r18_c232 bl[232] br[232] wl[18] vdd gnd cell_6t
Xbit_r19_c232 bl[232] br[232] wl[19] vdd gnd cell_6t
Xbit_r20_c232 bl[232] br[232] wl[20] vdd gnd cell_6t
Xbit_r21_c232 bl[232] br[232] wl[21] vdd gnd cell_6t
Xbit_r22_c232 bl[232] br[232] wl[22] vdd gnd cell_6t
Xbit_r23_c232 bl[232] br[232] wl[23] vdd gnd cell_6t
Xbit_r24_c232 bl[232] br[232] wl[24] vdd gnd cell_6t
Xbit_r25_c232 bl[232] br[232] wl[25] vdd gnd cell_6t
Xbit_r26_c232 bl[232] br[232] wl[26] vdd gnd cell_6t
Xbit_r27_c232 bl[232] br[232] wl[27] vdd gnd cell_6t
Xbit_r28_c232 bl[232] br[232] wl[28] vdd gnd cell_6t
Xbit_r29_c232 bl[232] br[232] wl[29] vdd gnd cell_6t
Xbit_r30_c232 bl[232] br[232] wl[30] vdd gnd cell_6t
Xbit_r31_c232 bl[232] br[232] wl[31] vdd gnd cell_6t
Xbit_r32_c232 bl[232] br[232] wl[32] vdd gnd cell_6t
Xbit_r33_c232 bl[232] br[232] wl[33] vdd gnd cell_6t
Xbit_r34_c232 bl[232] br[232] wl[34] vdd gnd cell_6t
Xbit_r35_c232 bl[232] br[232] wl[35] vdd gnd cell_6t
Xbit_r36_c232 bl[232] br[232] wl[36] vdd gnd cell_6t
Xbit_r37_c232 bl[232] br[232] wl[37] vdd gnd cell_6t
Xbit_r38_c232 bl[232] br[232] wl[38] vdd gnd cell_6t
Xbit_r39_c232 bl[232] br[232] wl[39] vdd gnd cell_6t
Xbit_r40_c232 bl[232] br[232] wl[40] vdd gnd cell_6t
Xbit_r41_c232 bl[232] br[232] wl[41] vdd gnd cell_6t
Xbit_r42_c232 bl[232] br[232] wl[42] vdd gnd cell_6t
Xbit_r43_c232 bl[232] br[232] wl[43] vdd gnd cell_6t
Xbit_r44_c232 bl[232] br[232] wl[44] vdd gnd cell_6t
Xbit_r45_c232 bl[232] br[232] wl[45] vdd gnd cell_6t
Xbit_r46_c232 bl[232] br[232] wl[46] vdd gnd cell_6t
Xbit_r47_c232 bl[232] br[232] wl[47] vdd gnd cell_6t
Xbit_r48_c232 bl[232] br[232] wl[48] vdd gnd cell_6t
Xbit_r49_c232 bl[232] br[232] wl[49] vdd gnd cell_6t
Xbit_r50_c232 bl[232] br[232] wl[50] vdd gnd cell_6t
Xbit_r51_c232 bl[232] br[232] wl[51] vdd gnd cell_6t
Xbit_r52_c232 bl[232] br[232] wl[52] vdd gnd cell_6t
Xbit_r53_c232 bl[232] br[232] wl[53] vdd gnd cell_6t
Xbit_r54_c232 bl[232] br[232] wl[54] vdd gnd cell_6t
Xbit_r55_c232 bl[232] br[232] wl[55] vdd gnd cell_6t
Xbit_r56_c232 bl[232] br[232] wl[56] vdd gnd cell_6t
Xbit_r57_c232 bl[232] br[232] wl[57] vdd gnd cell_6t
Xbit_r58_c232 bl[232] br[232] wl[58] vdd gnd cell_6t
Xbit_r59_c232 bl[232] br[232] wl[59] vdd gnd cell_6t
Xbit_r60_c232 bl[232] br[232] wl[60] vdd gnd cell_6t
Xbit_r61_c232 bl[232] br[232] wl[61] vdd gnd cell_6t
Xbit_r62_c232 bl[232] br[232] wl[62] vdd gnd cell_6t
Xbit_r63_c232 bl[232] br[232] wl[63] vdd gnd cell_6t
Xbit_r64_c232 bl[232] br[232] wl[64] vdd gnd cell_6t
Xbit_r65_c232 bl[232] br[232] wl[65] vdd gnd cell_6t
Xbit_r66_c232 bl[232] br[232] wl[66] vdd gnd cell_6t
Xbit_r67_c232 bl[232] br[232] wl[67] vdd gnd cell_6t
Xbit_r68_c232 bl[232] br[232] wl[68] vdd gnd cell_6t
Xbit_r69_c232 bl[232] br[232] wl[69] vdd gnd cell_6t
Xbit_r70_c232 bl[232] br[232] wl[70] vdd gnd cell_6t
Xbit_r71_c232 bl[232] br[232] wl[71] vdd gnd cell_6t
Xbit_r72_c232 bl[232] br[232] wl[72] vdd gnd cell_6t
Xbit_r73_c232 bl[232] br[232] wl[73] vdd gnd cell_6t
Xbit_r74_c232 bl[232] br[232] wl[74] vdd gnd cell_6t
Xbit_r75_c232 bl[232] br[232] wl[75] vdd gnd cell_6t
Xbit_r76_c232 bl[232] br[232] wl[76] vdd gnd cell_6t
Xbit_r77_c232 bl[232] br[232] wl[77] vdd gnd cell_6t
Xbit_r78_c232 bl[232] br[232] wl[78] vdd gnd cell_6t
Xbit_r79_c232 bl[232] br[232] wl[79] vdd gnd cell_6t
Xbit_r80_c232 bl[232] br[232] wl[80] vdd gnd cell_6t
Xbit_r81_c232 bl[232] br[232] wl[81] vdd gnd cell_6t
Xbit_r82_c232 bl[232] br[232] wl[82] vdd gnd cell_6t
Xbit_r83_c232 bl[232] br[232] wl[83] vdd gnd cell_6t
Xbit_r84_c232 bl[232] br[232] wl[84] vdd gnd cell_6t
Xbit_r85_c232 bl[232] br[232] wl[85] vdd gnd cell_6t
Xbit_r86_c232 bl[232] br[232] wl[86] vdd gnd cell_6t
Xbit_r87_c232 bl[232] br[232] wl[87] vdd gnd cell_6t
Xbit_r88_c232 bl[232] br[232] wl[88] vdd gnd cell_6t
Xbit_r89_c232 bl[232] br[232] wl[89] vdd gnd cell_6t
Xbit_r90_c232 bl[232] br[232] wl[90] vdd gnd cell_6t
Xbit_r91_c232 bl[232] br[232] wl[91] vdd gnd cell_6t
Xbit_r92_c232 bl[232] br[232] wl[92] vdd gnd cell_6t
Xbit_r93_c232 bl[232] br[232] wl[93] vdd gnd cell_6t
Xbit_r94_c232 bl[232] br[232] wl[94] vdd gnd cell_6t
Xbit_r95_c232 bl[232] br[232] wl[95] vdd gnd cell_6t
Xbit_r96_c232 bl[232] br[232] wl[96] vdd gnd cell_6t
Xbit_r97_c232 bl[232] br[232] wl[97] vdd gnd cell_6t
Xbit_r98_c232 bl[232] br[232] wl[98] vdd gnd cell_6t
Xbit_r99_c232 bl[232] br[232] wl[99] vdd gnd cell_6t
Xbit_r100_c232 bl[232] br[232] wl[100] vdd gnd cell_6t
Xbit_r101_c232 bl[232] br[232] wl[101] vdd gnd cell_6t
Xbit_r102_c232 bl[232] br[232] wl[102] vdd gnd cell_6t
Xbit_r103_c232 bl[232] br[232] wl[103] vdd gnd cell_6t
Xbit_r104_c232 bl[232] br[232] wl[104] vdd gnd cell_6t
Xbit_r105_c232 bl[232] br[232] wl[105] vdd gnd cell_6t
Xbit_r106_c232 bl[232] br[232] wl[106] vdd gnd cell_6t
Xbit_r107_c232 bl[232] br[232] wl[107] vdd gnd cell_6t
Xbit_r108_c232 bl[232] br[232] wl[108] vdd gnd cell_6t
Xbit_r109_c232 bl[232] br[232] wl[109] vdd gnd cell_6t
Xbit_r110_c232 bl[232] br[232] wl[110] vdd gnd cell_6t
Xbit_r111_c232 bl[232] br[232] wl[111] vdd gnd cell_6t
Xbit_r112_c232 bl[232] br[232] wl[112] vdd gnd cell_6t
Xbit_r113_c232 bl[232] br[232] wl[113] vdd gnd cell_6t
Xbit_r114_c232 bl[232] br[232] wl[114] vdd gnd cell_6t
Xbit_r115_c232 bl[232] br[232] wl[115] vdd gnd cell_6t
Xbit_r116_c232 bl[232] br[232] wl[116] vdd gnd cell_6t
Xbit_r117_c232 bl[232] br[232] wl[117] vdd gnd cell_6t
Xbit_r118_c232 bl[232] br[232] wl[118] vdd gnd cell_6t
Xbit_r119_c232 bl[232] br[232] wl[119] vdd gnd cell_6t
Xbit_r120_c232 bl[232] br[232] wl[120] vdd gnd cell_6t
Xbit_r121_c232 bl[232] br[232] wl[121] vdd gnd cell_6t
Xbit_r122_c232 bl[232] br[232] wl[122] vdd gnd cell_6t
Xbit_r123_c232 bl[232] br[232] wl[123] vdd gnd cell_6t
Xbit_r124_c232 bl[232] br[232] wl[124] vdd gnd cell_6t
Xbit_r125_c232 bl[232] br[232] wl[125] vdd gnd cell_6t
Xbit_r126_c232 bl[232] br[232] wl[126] vdd gnd cell_6t
Xbit_r127_c232 bl[232] br[232] wl[127] vdd gnd cell_6t
Xbit_r0_c233 bl[233] br[233] wl[0] vdd gnd cell_6t
Xbit_r1_c233 bl[233] br[233] wl[1] vdd gnd cell_6t
Xbit_r2_c233 bl[233] br[233] wl[2] vdd gnd cell_6t
Xbit_r3_c233 bl[233] br[233] wl[3] vdd gnd cell_6t
Xbit_r4_c233 bl[233] br[233] wl[4] vdd gnd cell_6t
Xbit_r5_c233 bl[233] br[233] wl[5] vdd gnd cell_6t
Xbit_r6_c233 bl[233] br[233] wl[6] vdd gnd cell_6t
Xbit_r7_c233 bl[233] br[233] wl[7] vdd gnd cell_6t
Xbit_r8_c233 bl[233] br[233] wl[8] vdd gnd cell_6t
Xbit_r9_c233 bl[233] br[233] wl[9] vdd gnd cell_6t
Xbit_r10_c233 bl[233] br[233] wl[10] vdd gnd cell_6t
Xbit_r11_c233 bl[233] br[233] wl[11] vdd gnd cell_6t
Xbit_r12_c233 bl[233] br[233] wl[12] vdd gnd cell_6t
Xbit_r13_c233 bl[233] br[233] wl[13] vdd gnd cell_6t
Xbit_r14_c233 bl[233] br[233] wl[14] vdd gnd cell_6t
Xbit_r15_c233 bl[233] br[233] wl[15] vdd gnd cell_6t
Xbit_r16_c233 bl[233] br[233] wl[16] vdd gnd cell_6t
Xbit_r17_c233 bl[233] br[233] wl[17] vdd gnd cell_6t
Xbit_r18_c233 bl[233] br[233] wl[18] vdd gnd cell_6t
Xbit_r19_c233 bl[233] br[233] wl[19] vdd gnd cell_6t
Xbit_r20_c233 bl[233] br[233] wl[20] vdd gnd cell_6t
Xbit_r21_c233 bl[233] br[233] wl[21] vdd gnd cell_6t
Xbit_r22_c233 bl[233] br[233] wl[22] vdd gnd cell_6t
Xbit_r23_c233 bl[233] br[233] wl[23] vdd gnd cell_6t
Xbit_r24_c233 bl[233] br[233] wl[24] vdd gnd cell_6t
Xbit_r25_c233 bl[233] br[233] wl[25] vdd gnd cell_6t
Xbit_r26_c233 bl[233] br[233] wl[26] vdd gnd cell_6t
Xbit_r27_c233 bl[233] br[233] wl[27] vdd gnd cell_6t
Xbit_r28_c233 bl[233] br[233] wl[28] vdd gnd cell_6t
Xbit_r29_c233 bl[233] br[233] wl[29] vdd gnd cell_6t
Xbit_r30_c233 bl[233] br[233] wl[30] vdd gnd cell_6t
Xbit_r31_c233 bl[233] br[233] wl[31] vdd gnd cell_6t
Xbit_r32_c233 bl[233] br[233] wl[32] vdd gnd cell_6t
Xbit_r33_c233 bl[233] br[233] wl[33] vdd gnd cell_6t
Xbit_r34_c233 bl[233] br[233] wl[34] vdd gnd cell_6t
Xbit_r35_c233 bl[233] br[233] wl[35] vdd gnd cell_6t
Xbit_r36_c233 bl[233] br[233] wl[36] vdd gnd cell_6t
Xbit_r37_c233 bl[233] br[233] wl[37] vdd gnd cell_6t
Xbit_r38_c233 bl[233] br[233] wl[38] vdd gnd cell_6t
Xbit_r39_c233 bl[233] br[233] wl[39] vdd gnd cell_6t
Xbit_r40_c233 bl[233] br[233] wl[40] vdd gnd cell_6t
Xbit_r41_c233 bl[233] br[233] wl[41] vdd gnd cell_6t
Xbit_r42_c233 bl[233] br[233] wl[42] vdd gnd cell_6t
Xbit_r43_c233 bl[233] br[233] wl[43] vdd gnd cell_6t
Xbit_r44_c233 bl[233] br[233] wl[44] vdd gnd cell_6t
Xbit_r45_c233 bl[233] br[233] wl[45] vdd gnd cell_6t
Xbit_r46_c233 bl[233] br[233] wl[46] vdd gnd cell_6t
Xbit_r47_c233 bl[233] br[233] wl[47] vdd gnd cell_6t
Xbit_r48_c233 bl[233] br[233] wl[48] vdd gnd cell_6t
Xbit_r49_c233 bl[233] br[233] wl[49] vdd gnd cell_6t
Xbit_r50_c233 bl[233] br[233] wl[50] vdd gnd cell_6t
Xbit_r51_c233 bl[233] br[233] wl[51] vdd gnd cell_6t
Xbit_r52_c233 bl[233] br[233] wl[52] vdd gnd cell_6t
Xbit_r53_c233 bl[233] br[233] wl[53] vdd gnd cell_6t
Xbit_r54_c233 bl[233] br[233] wl[54] vdd gnd cell_6t
Xbit_r55_c233 bl[233] br[233] wl[55] vdd gnd cell_6t
Xbit_r56_c233 bl[233] br[233] wl[56] vdd gnd cell_6t
Xbit_r57_c233 bl[233] br[233] wl[57] vdd gnd cell_6t
Xbit_r58_c233 bl[233] br[233] wl[58] vdd gnd cell_6t
Xbit_r59_c233 bl[233] br[233] wl[59] vdd gnd cell_6t
Xbit_r60_c233 bl[233] br[233] wl[60] vdd gnd cell_6t
Xbit_r61_c233 bl[233] br[233] wl[61] vdd gnd cell_6t
Xbit_r62_c233 bl[233] br[233] wl[62] vdd gnd cell_6t
Xbit_r63_c233 bl[233] br[233] wl[63] vdd gnd cell_6t
Xbit_r64_c233 bl[233] br[233] wl[64] vdd gnd cell_6t
Xbit_r65_c233 bl[233] br[233] wl[65] vdd gnd cell_6t
Xbit_r66_c233 bl[233] br[233] wl[66] vdd gnd cell_6t
Xbit_r67_c233 bl[233] br[233] wl[67] vdd gnd cell_6t
Xbit_r68_c233 bl[233] br[233] wl[68] vdd gnd cell_6t
Xbit_r69_c233 bl[233] br[233] wl[69] vdd gnd cell_6t
Xbit_r70_c233 bl[233] br[233] wl[70] vdd gnd cell_6t
Xbit_r71_c233 bl[233] br[233] wl[71] vdd gnd cell_6t
Xbit_r72_c233 bl[233] br[233] wl[72] vdd gnd cell_6t
Xbit_r73_c233 bl[233] br[233] wl[73] vdd gnd cell_6t
Xbit_r74_c233 bl[233] br[233] wl[74] vdd gnd cell_6t
Xbit_r75_c233 bl[233] br[233] wl[75] vdd gnd cell_6t
Xbit_r76_c233 bl[233] br[233] wl[76] vdd gnd cell_6t
Xbit_r77_c233 bl[233] br[233] wl[77] vdd gnd cell_6t
Xbit_r78_c233 bl[233] br[233] wl[78] vdd gnd cell_6t
Xbit_r79_c233 bl[233] br[233] wl[79] vdd gnd cell_6t
Xbit_r80_c233 bl[233] br[233] wl[80] vdd gnd cell_6t
Xbit_r81_c233 bl[233] br[233] wl[81] vdd gnd cell_6t
Xbit_r82_c233 bl[233] br[233] wl[82] vdd gnd cell_6t
Xbit_r83_c233 bl[233] br[233] wl[83] vdd gnd cell_6t
Xbit_r84_c233 bl[233] br[233] wl[84] vdd gnd cell_6t
Xbit_r85_c233 bl[233] br[233] wl[85] vdd gnd cell_6t
Xbit_r86_c233 bl[233] br[233] wl[86] vdd gnd cell_6t
Xbit_r87_c233 bl[233] br[233] wl[87] vdd gnd cell_6t
Xbit_r88_c233 bl[233] br[233] wl[88] vdd gnd cell_6t
Xbit_r89_c233 bl[233] br[233] wl[89] vdd gnd cell_6t
Xbit_r90_c233 bl[233] br[233] wl[90] vdd gnd cell_6t
Xbit_r91_c233 bl[233] br[233] wl[91] vdd gnd cell_6t
Xbit_r92_c233 bl[233] br[233] wl[92] vdd gnd cell_6t
Xbit_r93_c233 bl[233] br[233] wl[93] vdd gnd cell_6t
Xbit_r94_c233 bl[233] br[233] wl[94] vdd gnd cell_6t
Xbit_r95_c233 bl[233] br[233] wl[95] vdd gnd cell_6t
Xbit_r96_c233 bl[233] br[233] wl[96] vdd gnd cell_6t
Xbit_r97_c233 bl[233] br[233] wl[97] vdd gnd cell_6t
Xbit_r98_c233 bl[233] br[233] wl[98] vdd gnd cell_6t
Xbit_r99_c233 bl[233] br[233] wl[99] vdd gnd cell_6t
Xbit_r100_c233 bl[233] br[233] wl[100] vdd gnd cell_6t
Xbit_r101_c233 bl[233] br[233] wl[101] vdd gnd cell_6t
Xbit_r102_c233 bl[233] br[233] wl[102] vdd gnd cell_6t
Xbit_r103_c233 bl[233] br[233] wl[103] vdd gnd cell_6t
Xbit_r104_c233 bl[233] br[233] wl[104] vdd gnd cell_6t
Xbit_r105_c233 bl[233] br[233] wl[105] vdd gnd cell_6t
Xbit_r106_c233 bl[233] br[233] wl[106] vdd gnd cell_6t
Xbit_r107_c233 bl[233] br[233] wl[107] vdd gnd cell_6t
Xbit_r108_c233 bl[233] br[233] wl[108] vdd gnd cell_6t
Xbit_r109_c233 bl[233] br[233] wl[109] vdd gnd cell_6t
Xbit_r110_c233 bl[233] br[233] wl[110] vdd gnd cell_6t
Xbit_r111_c233 bl[233] br[233] wl[111] vdd gnd cell_6t
Xbit_r112_c233 bl[233] br[233] wl[112] vdd gnd cell_6t
Xbit_r113_c233 bl[233] br[233] wl[113] vdd gnd cell_6t
Xbit_r114_c233 bl[233] br[233] wl[114] vdd gnd cell_6t
Xbit_r115_c233 bl[233] br[233] wl[115] vdd gnd cell_6t
Xbit_r116_c233 bl[233] br[233] wl[116] vdd gnd cell_6t
Xbit_r117_c233 bl[233] br[233] wl[117] vdd gnd cell_6t
Xbit_r118_c233 bl[233] br[233] wl[118] vdd gnd cell_6t
Xbit_r119_c233 bl[233] br[233] wl[119] vdd gnd cell_6t
Xbit_r120_c233 bl[233] br[233] wl[120] vdd gnd cell_6t
Xbit_r121_c233 bl[233] br[233] wl[121] vdd gnd cell_6t
Xbit_r122_c233 bl[233] br[233] wl[122] vdd gnd cell_6t
Xbit_r123_c233 bl[233] br[233] wl[123] vdd gnd cell_6t
Xbit_r124_c233 bl[233] br[233] wl[124] vdd gnd cell_6t
Xbit_r125_c233 bl[233] br[233] wl[125] vdd gnd cell_6t
Xbit_r126_c233 bl[233] br[233] wl[126] vdd gnd cell_6t
Xbit_r127_c233 bl[233] br[233] wl[127] vdd gnd cell_6t
Xbit_r0_c234 bl[234] br[234] wl[0] vdd gnd cell_6t
Xbit_r1_c234 bl[234] br[234] wl[1] vdd gnd cell_6t
Xbit_r2_c234 bl[234] br[234] wl[2] vdd gnd cell_6t
Xbit_r3_c234 bl[234] br[234] wl[3] vdd gnd cell_6t
Xbit_r4_c234 bl[234] br[234] wl[4] vdd gnd cell_6t
Xbit_r5_c234 bl[234] br[234] wl[5] vdd gnd cell_6t
Xbit_r6_c234 bl[234] br[234] wl[6] vdd gnd cell_6t
Xbit_r7_c234 bl[234] br[234] wl[7] vdd gnd cell_6t
Xbit_r8_c234 bl[234] br[234] wl[8] vdd gnd cell_6t
Xbit_r9_c234 bl[234] br[234] wl[9] vdd gnd cell_6t
Xbit_r10_c234 bl[234] br[234] wl[10] vdd gnd cell_6t
Xbit_r11_c234 bl[234] br[234] wl[11] vdd gnd cell_6t
Xbit_r12_c234 bl[234] br[234] wl[12] vdd gnd cell_6t
Xbit_r13_c234 bl[234] br[234] wl[13] vdd gnd cell_6t
Xbit_r14_c234 bl[234] br[234] wl[14] vdd gnd cell_6t
Xbit_r15_c234 bl[234] br[234] wl[15] vdd gnd cell_6t
Xbit_r16_c234 bl[234] br[234] wl[16] vdd gnd cell_6t
Xbit_r17_c234 bl[234] br[234] wl[17] vdd gnd cell_6t
Xbit_r18_c234 bl[234] br[234] wl[18] vdd gnd cell_6t
Xbit_r19_c234 bl[234] br[234] wl[19] vdd gnd cell_6t
Xbit_r20_c234 bl[234] br[234] wl[20] vdd gnd cell_6t
Xbit_r21_c234 bl[234] br[234] wl[21] vdd gnd cell_6t
Xbit_r22_c234 bl[234] br[234] wl[22] vdd gnd cell_6t
Xbit_r23_c234 bl[234] br[234] wl[23] vdd gnd cell_6t
Xbit_r24_c234 bl[234] br[234] wl[24] vdd gnd cell_6t
Xbit_r25_c234 bl[234] br[234] wl[25] vdd gnd cell_6t
Xbit_r26_c234 bl[234] br[234] wl[26] vdd gnd cell_6t
Xbit_r27_c234 bl[234] br[234] wl[27] vdd gnd cell_6t
Xbit_r28_c234 bl[234] br[234] wl[28] vdd gnd cell_6t
Xbit_r29_c234 bl[234] br[234] wl[29] vdd gnd cell_6t
Xbit_r30_c234 bl[234] br[234] wl[30] vdd gnd cell_6t
Xbit_r31_c234 bl[234] br[234] wl[31] vdd gnd cell_6t
Xbit_r32_c234 bl[234] br[234] wl[32] vdd gnd cell_6t
Xbit_r33_c234 bl[234] br[234] wl[33] vdd gnd cell_6t
Xbit_r34_c234 bl[234] br[234] wl[34] vdd gnd cell_6t
Xbit_r35_c234 bl[234] br[234] wl[35] vdd gnd cell_6t
Xbit_r36_c234 bl[234] br[234] wl[36] vdd gnd cell_6t
Xbit_r37_c234 bl[234] br[234] wl[37] vdd gnd cell_6t
Xbit_r38_c234 bl[234] br[234] wl[38] vdd gnd cell_6t
Xbit_r39_c234 bl[234] br[234] wl[39] vdd gnd cell_6t
Xbit_r40_c234 bl[234] br[234] wl[40] vdd gnd cell_6t
Xbit_r41_c234 bl[234] br[234] wl[41] vdd gnd cell_6t
Xbit_r42_c234 bl[234] br[234] wl[42] vdd gnd cell_6t
Xbit_r43_c234 bl[234] br[234] wl[43] vdd gnd cell_6t
Xbit_r44_c234 bl[234] br[234] wl[44] vdd gnd cell_6t
Xbit_r45_c234 bl[234] br[234] wl[45] vdd gnd cell_6t
Xbit_r46_c234 bl[234] br[234] wl[46] vdd gnd cell_6t
Xbit_r47_c234 bl[234] br[234] wl[47] vdd gnd cell_6t
Xbit_r48_c234 bl[234] br[234] wl[48] vdd gnd cell_6t
Xbit_r49_c234 bl[234] br[234] wl[49] vdd gnd cell_6t
Xbit_r50_c234 bl[234] br[234] wl[50] vdd gnd cell_6t
Xbit_r51_c234 bl[234] br[234] wl[51] vdd gnd cell_6t
Xbit_r52_c234 bl[234] br[234] wl[52] vdd gnd cell_6t
Xbit_r53_c234 bl[234] br[234] wl[53] vdd gnd cell_6t
Xbit_r54_c234 bl[234] br[234] wl[54] vdd gnd cell_6t
Xbit_r55_c234 bl[234] br[234] wl[55] vdd gnd cell_6t
Xbit_r56_c234 bl[234] br[234] wl[56] vdd gnd cell_6t
Xbit_r57_c234 bl[234] br[234] wl[57] vdd gnd cell_6t
Xbit_r58_c234 bl[234] br[234] wl[58] vdd gnd cell_6t
Xbit_r59_c234 bl[234] br[234] wl[59] vdd gnd cell_6t
Xbit_r60_c234 bl[234] br[234] wl[60] vdd gnd cell_6t
Xbit_r61_c234 bl[234] br[234] wl[61] vdd gnd cell_6t
Xbit_r62_c234 bl[234] br[234] wl[62] vdd gnd cell_6t
Xbit_r63_c234 bl[234] br[234] wl[63] vdd gnd cell_6t
Xbit_r64_c234 bl[234] br[234] wl[64] vdd gnd cell_6t
Xbit_r65_c234 bl[234] br[234] wl[65] vdd gnd cell_6t
Xbit_r66_c234 bl[234] br[234] wl[66] vdd gnd cell_6t
Xbit_r67_c234 bl[234] br[234] wl[67] vdd gnd cell_6t
Xbit_r68_c234 bl[234] br[234] wl[68] vdd gnd cell_6t
Xbit_r69_c234 bl[234] br[234] wl[69] vdd gnd cell_6t
Xbit_r70_c234 bl[234] br[234] wl[70] vdd gnd cell_6t
Xbit_r71_c234 bl[234] br[234] wl[71] vdd gnd cell_6t
Xbit_r72_c234 bl[234] br[234] wl[72] vdd gnd cell_6t
Xbit_r73_c234 bl[234] br[234] wl[73] vdd gnd cell_6t
Xbit_r74_c234 bl[234] br[234] wl[74] vdd gnd cell_6t
Xbit_r75_c234 bl[234] br[234] wl[75] vdd gnd cell_6t
Xbit_r76_c234 bl[234] br[234] wl[76] vdd gnd cell_6t
Xbit_r77_c234 bl[234] br[234] wl[77] vdd gnd cell_6t
Xbit_r78_c234 bl[234] br[234] wl[78] vdd gnd cell_6t
Xbit_r79_c234 bl[234] br[234] wl[79] vdd gnd cell_6t
Xbit_r80_c234 bl[234] br[234] wl[80] vdd gnd cell_6t
Xbit_r81_c234 bl[234] br[234] wl[81] vdd gnd cell_6t
Xbit_r82_c234 bl[234] br[234] wl[82] vdd gnd cell_6t
Xbit_r83_c234 bl[234] br[234] wl[83] vdd gnd cell_6t
Xbit_r84_c234 bl[234] br[234] wl[84] vdd gnd cell_6t
Xbit_r85_c234 bl[234] br[234] wl[85] vdd gnd cell_6t
Xbit_r86_c234 bl[234] br[234] wl[86] vdd gnd cell_6t
Xbit_r87_c234 bl[234] br[234] wl[87] vdd gnd cell_6t
Xbit_r88_c234 bl[234] br[234] wl[88] vdd gnd cell_6t
Xbit_r89_c234 bl[234] br[234] wl[89] vdd gnd cell_6t
Xbit_r90_c234 bl[234] br[234] wl[90] vdd gnd cell_6t
Xbit_r91_c234 bl[234] br[234] wl[91] vdd gnd cell_6t
Xbit_r92_c234 bl[234] br[234] wl[92] vdd gnd cell_6t
Xbit_r93_c234 bl[234] br[234] wl[93] vdd gnd cell_6t
Xbit_r94_c234 bl[234] br[234] wl[94] vdd gnd cell_6t
Xbit_r95_c234 bl[234] br[234] wl[95] vdd gnd cell_6t
Xbit_r96_c234 bl[234] br[234] wl[96] vdd gnd cell_6t
Xbit_r97_c234 bl[234] br[234] wl[97] vdd gnd cell_6t
Xbit_r98_c234 bl[234] br[234] wl[98] vdd gnd cell_6t
Xbit_r99_c234 bl[234] br[234] wl[99] vdd gnd cell_6t
Xbit_r100_c234 bl[234] br[234] wl[100] vdd gnd cell_6t
Xbit_r101_c234 bl[234] br[234] wl[101] vdd gnd cell_6t
Xbit_r102_c234 bl[234] br[234] wl[102] vdd gnd cell_6t
Xbit_r103_c234 bl[234] br[234] wl[103] vdd gnd cell_6t
Xbit_r104_c234 bl[234] br[234] wl[104] vdd gnd cell_6t
Xbit_r105_c234 bl[234] br[234] wl[105] vdd gnd cell_6t
Xbit_r106_c234 bl[234] br[234] wl[106] vdd gnd cell_6t
Xbit_r107_c234 bl[234] br[234] wl[107] vdd gnd cell_6t
Xbit_r108_c234 bl[234] br[234] wl[108] vdd gnd cell_6t
Xbit_r109_c234 bl[234] br[234] wl[109] vdd gnd cell_6t
Xbit_r110_c234 bl[234] br[234] wl[110] vdd gnd cell_6t
Xbit_r111_c234 bl[234] br[234] wl[111] vdd gnd cell_6t
Xbit_r112_c234 bl[234] br[234] wl[112] vdd gnd cell_6t
Xbit_r113_c234 bl[234] br[234] wl[113] vdd gnd cell_6t
Xbit_r114_c234 bl[234] br[234] wl[114] vdd gnd cell_6t
Xbit_r115_c234 bl[234] br[234] wl[115] vdd gnd cell_6t
Xbit_r116_c234 bl[234] br[234] wl[116] vdd gnd cell_6t
Xbit_r117_c234 bl[234] br[234] wl[117] vdd gnd cell_6t
Xbit_r118_c234 bl[234] br[234] wl[118] vdd gnd cell_6t
Xbit_r119_c234 bl[234] br[234] wl[119] vdd gnd cell_6t
Xbit_r120_c234 bl[234] br[234] wl[120] vdd gnd cell_6t
Xbit_r121_c234 bl[234] br[234] wl[121] vdd gnd cell_6t
Xbit_r122_c234 bl[234] br[234] wl[122] vdd gnd cell_6t
Xbit_r123_c234 bl[234] br[234] wl[123] vdd gnd cell_6t
Xbit_r124_c234 bl[234] br[234] wl[124] vdd gnd cell_6t
Xbit_r125_c234 bl[234] br[234] wl[125] vdd gnd cell_6t
Xbit_r126_c234 bl[234] br[234] wl[126] vdd gnd cell_6t
Xbit_r127_c234 bl[234] br[234] wl[127] vdd gnd cell_6t
Xbit_r0_c235 bl[235] br[235] wl[0] vdd gnd cell_6t
Xbit_r1_c235 bl[235] br[235] wl[1] vdd gnd cell_6t
Xbit_r2_c235 bl[235] br[235] wl[2] vdd gnd cell_6t
Xbit_r3_c235 bl[235] br[235] wl[3] vdd gnd cell_6t
Xbit_r4_c235 bl[235] br[235] wl[4] vdd gnd cell_6t
Xbit_r5_c235 bl[235] br[235] wl[5] vdd gnd cell_6t
Xbit_r6_c235 bl[235] br[235] wl[6] vdd gnd cell_6t
Xbit_r7_c235 bl[235] br[235] wl[7] vdd gnd cell_6t
Xbit_r8_c235 bl[235] br[235] wl[8] vdd gnd cell_6t
Xbit_r9_c235 bl[235] br[235] wl[9] vdd gnd cell_6t
Xbit_r10_c235 bl[235] br[235] wl[10] vdd gnd cell_6t
Xbit_r11_c235 bl[235] br[235] wl[11] vdd gnd cell_6t
Xbit_r12_c235 bl[235] br[235] wl[12] vdd gnd cell_6t
Xbit_r13_c235 bl[235] br[235] wl[13] vdd gnd cell_6t
Xbit_r14_c235 bl[235] br[235] wl[14] vdd gnd cell_6t
Xbit_r15_c235 bl[235] br[235] wl[15] vdd gnd cell_6t
Xbit_r16_c235 bl[235] br[235] wl[16] vdd gnd cell_6t
Xbit_r17_c235 bl[235] br[235] wl[17] vdd gnd cell_6t
Xbit_r18_c235 bl[235] br[235] wl[18] vdd gnd cell_6t
Xbit_r19_c235 bl[235] br[235] wl[19] vdd gnd cell_6t
Xbit_r20_c235 bl[235] br[235] wl[20] vdd gnd cell_6t
Xbit_r21_c235 bl[235] br[235] wl[21] vdd gnd cell_6t
Xbit_r22_c235 bl[235] br[235] wl[22] vdd gnd cell_6t
Xbit_r23_c235 bl[235] br[235] wl[23] vdd gnd cell_6t
Xbit_r24_c235 bl[235] br[235] wl[24] vdd gnd cell_6t
Xbit_r25_c235 bl[235] br[235] wl[25] vdd gnd cell_6t
Xbit_r26_c235 bl[235] br[235] wl[26] vdd gnd cell_6t
Xbit_r27_c235 bl[235] br[235] wl[27] vdd gnd cell_6t
Xbit_r28_c235 bl[235] br[235] wl[28] vdd gnd cell_6t
Xbit_r29_c235 bl[235] br[235] wl[29] vdd gnd cell_6t
Xbit_r30_c235 bl[235] br[235] wl[30] vdd gnd cell_6t
Xbit_r31_c235 bl[235] br[235] wl[31] vdd gnd cell_6t
Xbit_r32_c235 bl[235] br[235] wl[32] vdd gnd cell_6t
Xbit_r33_c235 bl[235] br[235] wl[33] vdd gnd cell_6t
Xbit_r34_c235 bl[235] br[235] wl[34] vdd gnd cell_6t
Xbit_r35_c235 bl[235] br[235] wl[35] vdd gnd cell_6t
Xbit_r36_c235 bl[235] br[235] wl[36] vdd gnd cell_6t
Xbit_r37_c235 bl[235] br[235] wl[37] vdd gnd cell_6t
Xbit_r38_c235 bl[235] br[235] wl[38] vdd gnd cell_6t
Xbit_r39_c235 bl[235] br[235] wl[39] vdd gnd cell_6t
Xbit_r40_c235 bl[235] br[235] wl[40] vdd gnd cell_6t
Xbit_r41_c235 bl[235] br[235] wl[41] vdd gnd cell_6t
Xbit_r42_c235 bl[235] br[235] wl[42] vdd gnd cell_6t
Xbit_r43_c235 bl[235] br[235] wl[43] vdd gnd cell_6t
Xbit_r44_c235 bl[235] br[235] wl[44] vdd gnd cell_6t
Xbit_r45_c235 bl[235] br[235] wl[45] vdd gnd cell_6t
Xbit_r46_c235 bl[235] br[235] wl[46] vdd gnd cell_6t
Xbit_r47_c235 bl[235] br[235] wl[47] vdd gnd cell_6t
Xbit_r48_c235 bl[235] br[235] wl[48] vdd gnd cell_6t
Xbit_r49_c235 bl[235] br[235] wl[49] vdd gnd cell_6t
Xbit_r50_c235 bl[235] br[235] wl[50] vdd gnd cell_6t
Xbit_r51_c235 bl[235] br[235] wl[51] vdd gnd cell_6t
Xbit_r52_c235 bl[235] br[235] wl[52] vdd gnd cell_6t
Xbit_r53_c235 bl[235] br[235] wl[53] vdd gnd cell_6t
Xbit_r54_c235 bl[235] br[235] wl[54] vdd gnd cell_6t
Xbit_r55_c235 bl[235] br[235] wl[55] vdd gnd cell_6t
Xbit_r56_c235 bl[235] br[235] wl[56] vdd gnd cell_6t
Xbit_r57_c235 bl[235] br[235] wl[57] vdd gnd cell_6t
Xbit_r58_c235 bl[235] br[235] wl[58] vdd gnd cell_6t
Xbit_r59_c235 bl[235] br[235] wl[59] vdd gnd cell_6t
Xbit_r60_c235 bl[235] br[235] wl[60] vdd gnd cell_6t
Xbit_r61_c235 bl[235] br[235] wl[61] vdd gnd cell_6t
Xbit_r62_c235 bl[235] br[235] wl[62] vdd gnd cell_6t
Xbit_r63_c235 bl[235] br[235] wl[63] vdd gnd cell_6t
Xbit_r64_c235 bl[235] br[235] wl[64] vdd gnd cell_6t
Xbit_r65_c235 bl[235] br[235] wl[65] vdd gnd cell_6t
Xbit_r66_c235 bl[235] br[235] wl[66] vdd gnd cell_6t
Xbit_r67_c235 bl[235] br[235] wl[67] vdd gnd cell_6t
Xbit_r68_c235 bl[235] br[235] wl[68] vdd gnd cell_6t
Xbit_r69_c235 bl[235] br[235] wl[69] vdd gnd cell_6t
Xbit_r70_c235 bl[235] br[235] wl[70] vdd gnd cell_6t
Xbit_r71_c235 bl[235] br[235] wl[71] vdd gnd cell_6t
Xbit_r72_c235 bl[235] br[235] wl[72] vdd gnd cell_6t
Xbit_r73_c235 bl[235] br[235] wl[73] vdd gnd cell_6t
Xbit_r74_c235 bl[235] br[235] wl[74] vdd gnd cell_6t
Xbit_r75_c235 bl[235] br[235] wl[75] vdd gnd cell_6t
Xbit_r76_c235 bl[235] br[235] wl[76] vdd gnd cell_6t
Xbit_r77_c235 bl[235] br[235] wl[77] vdd gnd cell_6t
Xbit_r78_c235 bl[235] br[235] wl[78] vdd gnd cell_6t
Xbit_r79_c235 bl[235] br[235] wl[79] vdd gnd cell_6t
Xbit_r80_c235 bl[235] br[235] wl[80] vdd gnd cell_6t
Xbit_r81_c235 bl[235] br[235] wl[81] vdd gnd cell_6t
Xbit_r82_c235 bl[235] br[235] wl[82] vdd gnd cell_6t
Xbit_r83_c235 bl[235] br[235] wl[83] vdd gnd cell_6t
Xbit_r84_c235 bl[235] br[235] wl[84] vdd gnd cell_6t
Xbit_r85_c235 bl[235] br[235] wl[85] vdd gnd cell_6t
Xbit_r86_c235 bl[235] br[235] wl[86] vdd gnd cell_6t
Xbit_r87_c235 bl[235] br[235] wl[87] vdd gnd cell_6t
Xbit_r88_c235 bl[235] br[235] wl[88] vdd gnd cell_6t
Xbit_r89_c235 bl[235] br[235] wl[89] vdd gnd cell_6t
Xbit_r90_c235 bl[235] br[235] wl[90] vdd gnd cell_6t
Xbit_r91_c235 bl[235] br[235] wl[91] vdd gnd cell_6t
Xbit_r92_c235 bl[235] br[235] wl[92] vdd gnd cell_6t
Xbit_r93_c235 bl[235] br[235] wl[93] vdd gnd cell_6t
Xbit_r94_c235 bl[235] br[235] wl[94] vdd gnd cell_6t
Xbit_r95_c235 bl[235] br[235] wl[95] vdd gnd cell_6t
Xbit_r96_c235 bl[235] br[235] wl[96] vdd gnd cell_6t
Xbit_r97_c235 bl[235] br[235] wl[97] vdd gnd cell_6t
Xbit_r98_c235 bl[235] br[235] wl[98] vdd gnd cell_6t
Xbit_r99_c235 bl[235] br[235] wl[99] vdd gnd cell_6t
Xbit_r100_c235 bl[235] br[235] wl[100] vdd gnd cell_6t
Xbit_r101_c235 bl[235] br[235] wl[101] vdd gnd cell_6t
Xbit_r102_c235 bl[235] br[235] wl[102] vdd gnd cell_6t
Xbit_r103_c235 bl[235] br[235] wl[103] vdd gnd cell_6t
Xbit_r104_c235 bl[235] br[235] wl[104] vdd gnd cell_6t
Xbit_r105_c235 bl[235] br[235] wl[105] vdd gnd cell_6t
Xbit_r106_c235 bl[235] br[235] wl[106] vdd gnd cell_6t
Xbit_r107_c235 bl[235] br[235] wl[107] vdd gnd cell_6t
Xbit_r108_c235 bl[235] br[235] wl[108] vdd gnd cell_6t
Xbit_r109_c235 bl[235] br[235] wl[109] vdd gnd cell_6t
Xbit_r110_c235 bl[235] br[235] wl[110] vdd gnd cell_6t
Xbit_r111_c235 bl[235] br[235] wl[111] vdd gnd cell_6t
Xbit_r112_c235 bl[235] br[235] wl[112] vdd gnd cell_6t
Xbit_r113_c235 bl[235] br[235] wl[113] vdd gnd cell_6t
Xbit_r114_c235 bl[235] br[235] wl[114] vdd gnd cell_6t
Xbit_r115_c235 bl[235] br[235] wl[115] vdd gnd cell_6t
Xbit_r116_c235 bl[235] br[235] wl[116] vdd gnd cell_6t
Xbit_r117_c235 bl[235] br[235] wl[117] vdd gnd cell_6t
Xbit_r118_c235 bl[235] br[235] wl[118] vdd gnd cell_6t
Xbit_r119_c235 bl[235] br[235] wl[119] vdd gnd cell_6t
Xbit_r120_c235 bl[235] br[235] wl[120] vdd gnd cell_6t
Xbit_r121_c235 bl[235] br[235] wl[121] vdd gnd cell_6t
Xbit_r122_c235 bl[235] br[235] wl[122] vdd gnd cell_6t
Xbit_r123_c235 bl[235] br[235] wl[123] vdd gnd cell_6t
Xbit_r124_c235 bl[235] br[235] wl[124] vdd gnd cell_6t
Xbit_r125_c235 bl[235] br[235] wl[125] vdd gnd cell_6t
Xbit_r126_c235 bl[235] br[235] wl[126] vdd gnd cell_6t
Xbit_r127_c235 bl[235] br[235] wl[127] vdd gnd cell_6t
Xbit_r0_c236 bl[236] br[236] wl[0] vdd gnd cell_6t
Xbit_r1_c236 bl[236] br[236] wl[1] vdd gnd cell_6t
Xbit_r2_c236 bl[236] br[236] wl[2] vdd gnd cell_6t
Xbit_r3_c236 bl[236] br[236] wl[3] vdd gnd cell_6t
Xbit_r4_c236 bl[236] br[236] wl[4] vdd gnd cell_6t
Xbit_r5_c236 bl[236] br[236] wl[5] vdd gnd cell_6t
Xbit_r6_c236 bl[236] br[236] wl[6] vdd gnd cell_6t
Xbit_r7_c236 bl[236] br[236] wl[7] vdd gnd cell_6t
Xbit_r8_c236 bl[236] br[236] wl[8] vdd gnd cell_6t
Xbit_r9_c236 bl[236] br[236] wl[9] vdd gnd cell_6t
Xbit_r10_c236 bl[236] br[236] wl[10] vdd gnd cell_6t
Xbit_r11_c236 bl[236] br[236] wl[11] vdd gnd cell_6t
Xbit_r12_c236 bl[236] br[236] wl[12] vdd gnd cell_6t
Xbit_r13_c236 bl[236] br[236] wl[13] vdd gnd cell_6t
Xbit_r14_c236 bl[236] br[236] wl[14] vdd gnd cell_6t
Xbit_r15_c236 bl[236] br[236] wl[15] vdd gnd cell_6t
Xbit_r16_c236 bl[236] br[236] wl[16] vdd gnd cell_6t
Xbit_r17_c236 bl[236] br[236] wl[17] vdd gnd cell_6t
Xbit_r18_c236 bl[236] br[236] wl[18] vdd gnd cell_6t
Xbit_r19_c236 bl[236] br[236] wl[19] vdd gnd cell_6t
Xbit_r20_c236 bl[236] br[236] wl[20] vdd gnd cell_6t
Xbit_r21_c236 bl[236] br[236] wl[21] vdd gnd cell_6t
Xbit_r22_c236 bl[236] br[236] wl[22] vdd gnd cell_6t
Xbit_r23_c236 bl[236] br[236] wl[23] vdd gnd cell_6t
Xbit_r24_c236 bl[236] br[236] wl[24] vdd gnd cell_6t
Xbit_r25_c236 bl[236] br[236] wl[25] vdd gnd cell_6t
Xbit_r26_c236 bl[236] br[236] wl[26] vdd gnd cell_6t
Xbit_r27_c236 bl[236] br[236] wl[27] vdd gnd cell_6t
Xbit_r28_c236 bl[236] br[236] wl[28] vdd gnd cell_6t
Xbit_r29_c236 bl[236] br[236] wl[29] vdd gnd cell_6t
Xbit_r30_c236 bl[236] br[236] wl[30] vdd gnd cell_6t
Xbit_r31_c236 bl[236] br[236] wl[31] vdd gnd cell_6t
Xbit_r32_c236 bl[236] br[236] wl[32] vdd gnd cell_6t
Xbit_r33_c236 bl[236] br[236] wl[33] vdd gnd cell_6t
Xbit_r34_c236 bl[236] br[236] wl[34] vdd gnd cell_6t
Xbit_r35_c236 bl[236] br[236] wl[35] vdd gnd cell_6t
Xbit_r36_c236 bl[236] br[236] wl[36] vdd gnd cell_6t
Xbit_r37_c236 bl[236] br[236] wl[37] vdd gnd cell_6t
Xbit_r38_c236 bl[236] br[236] wl[38] vdd gnd cell_6t
Xbit_r39_c236 bl[236] br[236] wl[39] vdd gnd cell_6t
Xbit_r40_c236 bl[236] br[236] wl[40] vdd gnd cell_6t
Xbit_r41_c236 bl[236] br[236] wl[41] vdd gnd cell_6t
Xbit_r42_c236 bl[236] br[236] wl[42] vdd gnd cell_6t
Xbit_r43_c236 bl[236] br[236] wl[43] vdd gnd cell_6t
Xbit_r44_c236 bl[236] br[236] wl[44] vdd gnd cell_6t
Xbit_r45_c236 bl[236] br[236] wl[45] vdd gnd cell_6t
Xbit_r46_c236 bl[236] br[236] wl[46] vdd gnd cell_6t
Xbit_r47_c236 bl[236] br[236] wl[47] vdd gnd cell_6t
Xbit_r48_c236 bl[236] br[236] wl[48] vdd gnd cell_6t
Xbit_r49_c236 bl[236] br[236] wl[49] vdd gnd cell_6t
Xbit_r50_c236 bl[236] br[236] wl[50] vdd gnd cell_6t
Xbit_r51_c236 bl[236] br[236] wl[51] vdd gnd cell_6t
Xbit_r52_c236 bl[236] br[236] wl[52] vdd gnd cell_6t
Xbit_r53_c236 bl[236] br[236] wl[53] vdd gnd cell_6t
Xbit_r54_c236 bl[236] br[236] wl[54] vdd gnd cell_6t
Xbit_r55_c236 bl[236] br[236] wl[55] vdd gnd cell_6t
Xbit_r56_c236 bl[236] br[236] wl[56] vdd gnd cell_6t
Xbit_r57_c236 bl[236] br[236] wl[57] vdd gnd cell_6t
Xbit_r58_c236 bl[236] br[236] wl[58] vdd gnd cell_6t
Xbit_r59_c236 bl[236] br[236] wl[59] vdd gnd cell_6t
Xbit_r60_c236 bl[236] br[236] wl[60] vdd gnd cell_6t
Xbit_r61_c236 bl[236] br[236] wl[61] vdd gnd cell_6t
Xbit_r62_c236 bl[236] br[236] wl[62] vdd gnd cell_6t
Xbit_r63_c236 bl[236] br[236] wl[63] vdd gnd cell_6t
Xbit_r64_c236 bl[236] br[236] wl[64] vdd gnd cell_6t
Xbit_r65_c236 bl[236] br[236] wl[65] vdd gnd cell_6t
Xbit_r66_c236 bl[236] br[236] wl[66] vdd gnd cell_6t
Xbit_r67_c236 bl[236] br[236] wl[67] vdd gnd cell_6t
Xbit_r68_c236 bl[236] br[236] wl[68] vdd gnd cell_6t
Xbit_r69_c236 bl[236] br[236] wl[69] vdd gnd cell_6t
Xbit_r70_c236 bl[236] br[236] wl[70] vdd gnd cell_6t
Xbit_r71_c236 bl[236] br[236] wl[71] vdd gnd cell_6t
Xbit_r72_c236 bl[236] br[236] wl[72] vdd gnd cell_6t
Xbit_r73_c236 bl[236] br[236] wl[73] vdd gnd cell_6t
Xbit_r74_c236 bl[236] br[236] wl[74] vdd gnd cell_6t
Xbit_r75_c236 bl[236] br[236] wl[75] vdd gnd cell_6t
Xbit_r76_c236 bl[236] br[236] wl[76] vdd gnd cell_6t
Xbit_r77_c236 bl[236] br[236] wl[77] vdd gnd cell_6t
Xbit_r78_c236 bl[236] br[236] wl[78] vdd gnd cell_6t
Xbit_r79_c236 bl[236] br[236] wl[79] vdd gnd cell_6t
Xbit_r80_c236 bl[236] br[236] wl[80] vdd gnd cell_6t
Xbit_r81_c236 bl[236] br[236] wl[81] vdd gnd cell_6t
Xbit_r82_c236 bl[236] br[236] wl[82] vdd gnd cell_6t
Xbit_r83_c236 bl[236] br[236] wl[83] vdd gnd cell_6t
Xbit_r84_c236 bl[236] br[236] wl[84] vdd gnd cell_6t
Xbit_r85_c236 bl[236] br[236] wl[85] vdd gnd cell_6t
Xbit_r86_c236 bl[236] br[236] wl[86] vdd gnd cell_6t
Xbit_r87_c236 bl[236] br[236] wl[87] vdd gnd cell_6t
Xbit_r88_c236 bl[236] br[236] wl[88] vdd gnd cell_6t
Xbit_r89_c236 bl[236] br[236] wl[89] vdd gnd cell_6t
Xbit_r90_c236 bl[236] br[236] wl[90] vdd gnd cell_6t
Xbit_r91_c236 bl[236] br[236] wl[91] vdd gnd cell_6t
Xbit_r92_c236 bl[236] br[236] wl[92] vdd gnd cell_6t
Xbit_r93_c236 bl[236] br[236] wl[93] vdd gnd cell_6t
Xbit_r94_c236 bl[236] br[236] wl[94] vdd gnd cell_6t
Xbit_r95_c236 bl[236] br[236] wl[95] vdd gnd cell_6t
Xbit_r96_c236 bl[236] br[236] wl[96] vdd gnd cell_6t
Xbit_r97_c236 bl[236] br[236] wl[97] vdd gnd cell_6t
Xbit_r98_c236 bl[236] br[236] wl[98] vdd gnd cell_6t
Xbit_r99_c236 bl[236] br[236] wl[99] vdd gnd cell_6t
Xbit_r100_c236 bl[236] br[236] wl[100] vdd gnd cell_6t
Xbit_r101_c236 bl[236] br[236] wl[101] vdd gnd cell_6t
Xbit_r102_c236 bl[236] br[236] wl[102] vdd gnd cell_6t
Xbit_r103_c236 bl[236] br[236] wl[103] vdd gnd cell_6t
Xbit_r104_c236 bl[236] br[236] wl[104] vdd gnd cell_6t
Xbit_r105_c236 bl[236] br[236] wl[105] vdd gnd cell_6t
Xbit_r106_c236 bl[236] br[236] wl[106] vdd gnd cell_6t
Xbit_r107_c236 bl[236] br[236] wl[107] vdd gnd cell_6t
Xbit_r108_c236 bl[236] br[236] wl[108] vdd gnd cell_6t
Xbit_r109_c236 bl[236] br[236] wl[109] vdd gnd cell_6t
Xbit_r110_c236 bl[236] br[236] wl[110] vdd gnd cell_6t
Xbit_r111_c236 bl[236] br[236] wl[111] vdd gnd cell_6t
Xbit_r112_c236 bl[236] br[236] wl[112] vdd gnd cell_6t
Xbit_r113_c236 bl[236] br[236] wl[113] vdd gnd cell_6t
Xbit_r114_c236 bl[236] br[236] wl[114] vdd gnd cell_6t
Xbit_r115_c236 bl[236] br[236] wl[115] vdd gnd cell_6t
Xbit_r116_c236 bl[236] br[236] wl[116] vdd gnd cell_6t
Xbit_r117_c236 bl[236] br[236] wl[117] vdd gnd cell_6t
Xbit_r118_c236 bl[236] br[236] wl[118] vdd gnd cell_6t
Xbit_r119_c236 bl[236] br[236] wl[119] vdd gnd cell_6t
Xbit_r120_c236 bl[236] br[236] wl[120] vdd gnd cell_6t
Xbit_r121_c236 bl[236] br[236] wl[121] vdd gnd cell_6t
Xbit_r122_c236 bl[236] br[236] wl[122] vdd gnd cell_6t
Xbit_r123_c236 bl[236] br[236] wl[123] vdd gnd cell_6t
Xbit_r124_c236 bl[236] br[236] wl[124] vdd gnd cell_6t
Xbit_r125_c236 bl[236] br[236] wl[125] vdd gnd cell_6t
Xbit_r126_c236 bl[236] br[236] wl[126] vdd gnd cell_6t
Xbit_r127_c236 bl[236] br[236] wl[127] vdd gnd cell_6t
Xbit_r0_c237 bl[237] br[237] wl[0] vdd gnd cell_6t
Xbit_r1_c237 bl[237] br[237] wl[1] vdd gnd cell_6t
Xbit_r2_c237 bl[237] br[237] wl[2] vdd gnd cell_6t
Xbit_r3_c237 bl[237] br[237] wl[3] vdd gnd cell_6t
Xbit_r4_c237 bl[237] br[237] wl[4] vdd gnd cell_6t
Xbit_r5_c237 bl[237] br[237] wl[5] vdd gnd cell_6t
Xbit_r6_c237 bl[237] br[237] wl[6] vdd gnd cell_6t
Xbit_r7_c237 bl[237] br[237] wl[7] vdd gnd cell_6t
Xbit_r8_c237 bl[237] br[237] wl[8] vdd gnd cell_6t
Xbit_r9_c237 bl[237] br[237] wl[9] vdd gnd cell_6t
Xbit_r10_c237 bl[237] br[237] wl[10] vdd gnd cell_6t
Xbit_r11_c237 bl[237] br[237] wl[11] vdd gnd cell_6t
Xbit_r12_c237 bl[237] br[237] wl[12] vdd gnd cell_6t
Xbit_r13_c237 bl[237] br[237] wl[13] vdd gnd cell_6t
Xbit_r14_c237 bl[237] br[237] wl[14] vdd gnd cell_6t
Xbit_r15_c237 bl[237] br[237] wl[15] vdd gnd cell_6t
Xbit_r16_c237 bl[237] br[237] wl[16] vdd gnd cell_6t
Xbit_r17_c237 bl[237] br[237] wl[17] vdd gnd cell_6t
Xbit_r18_c237 bl[237] br[237] wl[18] vdd gnd cell_6t
Xbit_r19_c237 bl[237] br[237] wl[19] vdd gnd cell_6t
Xbit_r20_c237 bl[237] br[237] wl[20] vdd gnd cell_6t
Xbit_r21_c237 bl[237] br[237] wl[21] vdd gnd cell_6t
Xbit_r22_c237 bl[237] br[237] wl[22] vdd gnd cell_6t
Xbit_r23_c237 bl[237] br[237] wl[23] vdd gnd cell_6t
Xbit_r24_c237 bl[237] br[237] wl[24] vdd gnd cell_6t
Xbit_r25_c237 bl[237] br[237] wl[25] vdd gnd cell_6t
Xbit_r26_c237 bl[237] br[237] wl[26] vdd gnd cell_6t
Xbit_r27_c237 bl[237] br[237] wl[27] vdd gnd cell_6t
Xbit_r28_c237 bl[237] br[237] wl[28] vdd gnd cell_6t
Xbit_r29_c237 bl[237] br[237] wl[29] vdd gnd cell_6t
Xbit_r30_c237 bl[237] br[237] wl[30] vdd gnd cell_6t
Xbit_r31_c237 bl[237] br[237] wl[31] vdd gnd cell_6t
Xbit_r32_c237 bl[237] br[237] wl[32] vdd gnd cell_6t
Xbit_r33_c237 bl[237] br[237] wl[33] vdd gnd cell_6t
Xbit_r34_c237 bl[237] br[237] wl[34] vdd gnd cell_6t
Xbit_r35_c237 bl[237] br[237] wl[35] vdd gnd cell_6t
Xbit_r36_c237 bl[237] br[237] wl[36] vdd gnd cell_6t
Xbit_r37_c237 bl[237] br[237] wl[37] vdd gnd cell_6t
Xbit_r38_c237 bl[237] br[237] wl[38] vdd gnd cell_6t
Xbit_r39_c237 bl[237] br[237] wl[39] vdd gnd cell_6t
Xbit_r40_c237 bl[237] br[237] wl[40] vdd gnd cell_6t
Xbit_r41_c237 bl[237] br[237] wl[41] vdd gnd cell_6t
Xbit_r42_c237 bl[237] br[237] wl[42] vdd gnd cell_6t
Xbit_r43_c237 bl[237] br[237] wl[43] vdd gnd cell_6t
Xbit_r44_c237 bl[237] br[237] wl[44] vdd gnd cell_6t
Xbit_r45_c237 bl[237] br[237] wl[45] vdd gnd cell_6t
Xbit_r46_c237 bl[237] br[237] wl[46] vdd gnd cell_6t
Xbit_r47_c237 bl[237] br[237] wl[47] vdd gnd cell_6t
Xbit_r48_c237 bl[237] br[237] wl[48] vdd gnd cell_6t
Xbit_r49_c237 bl[237] br[237] wl[49] vdd gnd cell_6t
Xbit_r50_c237 bl[237] br[237] wl[50] vdd gnd cell_6t
Xbit_r51_c237 bl[237] br[237] wl[51] vdd gnd cell_6t
Xbit_r52_c237 bl[237] br[237] wl[52] vdd gnd cell_6t
Xbit_r53_c237 bl[237] br[237] wl[53] vdd gnd cell_6t
Xbit_r54_c237 bl[237] br[237] wl[54] vdd gnd cell_6t
Xbit_r55_c237 bl[237] br[237] wl[55] vdd gnd cell_6t
Xbit_r56_c237 bl[237] br[237] wl[56] vdd gnd cell_6t
Xbit_r57_c237 bl[237] br[237] wl[57] vdd gnd cell_6t
Xbit_r58_c237 bl[237] br[237] wl[58] vdd gnd cell_6t
Xbit_r59_c237 bl[237] br[237] wl[59] vdd gnd cell_6t
Xbit_r60_c237 bl[237] br[237] wl[60] vdd gnd cell_6t
Xbit_r61_c237 bl[237] br[237] wl[61] vdd gnd cell_6t
Xbit_r62_c237 bl[237] br[237] wl[62] vdd gnd cell_6t
Xbit_r63_c237 bl[237] br[237] wl[63] vdd gnd cell_6t
Xbit_r64_c237 bl[237] br[237] wl[64] vdd gnd cell_6t
Xbit_r65_c237 bl[237] br[237] wl[65] vdd gnd cell_6t
Xbit_r66_c237 bl[237] br[237] wl[66] vdd gnd cell_6t
Xbit_r67_c237 bl[237] br[237] wl[67] vdd gnd cell_6t
Xbit_r68_c237 bl[237] br[237] wl[68] vdd gnd cell_6t
Xbit_r69_c237 bl[237] br[237] wl[69] vdd gnd cell_6t
Xbit_r70_c237 bl[237] br[237] wl[70] vdd gnd cell_6t
Xbit_r71_c237 bl[237] br[237] wl[71] vdd gnd cell_6t
Xbit_r72_c237 bl[237] br[237] wl[72] vdd gnd cell_6t
Xbit_r73_c237 bl[237] br[237] wl[73] vdd gnd cell_6t
Xbit_r74_c237 bl[237] br[237] wl[74] vdd gnd cell_6t
Xbit_r75_c237 bl[237] br[237] wl[75] vdd gnd cell_6t
Xbit_r76_c237 bl[237] br[237] wl[76] vdd gnd cell_6t
Xbit_r77_c237 bl[237] br[237] wl[77] vdd gnd cell_6t
Xbit_r78_c237 bl[237] br[237] wl[78] vdd gnd cell_6t
Xbit_r79_c237 bl[237] br[237] wl[79] vdd gnd cell_6t
Xbit_r80_c237 bl[237] br[237] wl[80] vdd gnd cell_6t
Xbit_r81_c237 bl[237] br[237] wl[81] vdd gnd cell_6t
Xbit_r82_c237 bl[237] br[237] wl[82] vdd gnd cell_6t
Xbit_r83_c237 bl[237] br[237] wl[83] vdd gnd cell_6t
Xbit_r84_c237 bl[237] br[237] wl[84] vdd gnd cell_6t
Xbit_r85_c237 bl[237] br[237] wl[85] vdd gnd cell_6t
Xbit_r86_c237 bl[237] br[237] wl[86] vdd gnd cell_6t
Xbit_r87_c237 bl[237] br[237] wl[87] vdd gnd cell_6t
Xbit_r88_c237 bl[237] br[237] wl[88] vdd gnd cell_6t
Xbit_r89_c237 bl[237] br[237] wl[89] vdd gnd cell_6t
Xbit_r90_c237 bl[237] br[237] wl[90] vdd gnd cell_6t
Xbit_r91_c237 bl[237] br[237] wl[91] vdd gnd cell_6t
Xbit_r92_c237 bl[237] br[237] wl[92] vdd gnd cell_6t
Xbit_r93_c237 bl[237] br[237] wl[93] vdd gnd cell_6t
Xbit_r94_c237 bl[237] br[237] wl[94] vdd gnd cell_6t
Xbit_r95_c237 bl[237] br[237] wl[95] vdd gnd cell_6t
Xbit_r96_c237 bl[237] br[237] wl[96] vdd gnd cell_6t
Xbit_r97_c237 bl[237] br[237] wl[97] vdd gnd cell_6t
Xbit_r98_c237 bl[237] br[237] wl[98] vdd gnd cell_6t
Xbit_r99_c237 bl[237] br[237] wl[99] vdd gnd cell_6t
Xbit_r100_c237 bl[237] br[237] wl[100] vdd gnd cell_6t
Xbit_r101_c237 bl[237] br[237] wl[101] vdd gnd cell_6t
Xbit_r102_c237 bl[237] br[237] wl[102] vdd gnd cell_6t
Xbit_r103_c237 bl[237] br[237] wl[103] vdd gnd cell_6t
Xbit_r104_c237 bl[237] br[237] wl[104] vdd gnd cell_6t
Xbit_r105_c237 bl[237] br[237] wl[105] vdd gnd cell_6t
Xbit_r106_c237 bl[237] br[237] wl[106] vdd gnd cell_6t
Xbit_r107_c237 bl[237] br[237] wl[107] vdd gnd cell_6t
Xbit_r108_c237 bl[237] br[237] wl[108] vdd gnd cell_6t
Xbit_r109_c237 bl[237] br[237] wl[109] vdd gnd cell_6t
Xbit_r110_c237 bl[237] br[237] wl[110] vdd gnd cell_6t
Xbit_r111_c237 bl[237] br[237] wl[111] vdd gnd cell_6t
Xbit_r112_c237 bl[237] br[237] wl[112] vdd gnd cell_6t
Xbit_r113_c237 bl[237] br[237] wl[113] vdd gnd cell_6t
Xbit_r114_c237 bl[237] br[237] wl[114] vdd gnd cell_6t
Xbit_r115_c237 bl[237] br[237] wl[115] vdd gnd cell_6t
Xbit_r116_c237 bl[237] br[237] wl[116] vdd gnd cell_6t
Xbit_r117_c237 bl[237] br[237] wl[117] vdd gnd cell_6t
Xbit_r118_c237 bl[237] br[237] wl[118] vdd gnd cell_6t
Xbit_r119_c237 bl[237] br[237] wl[119] vdd gnd cell_6t
Xbit_r120_c237 bl[237] br[237] wl[120] vdd gnd cell_6t
Xbit_r121_c237 bl[237] br[237] wl[121] vdd gnd cell_6t
Xbit_r122_c237 bl[237] br[237] wl[122] vdd gnd cell_6t
Xbit_r123_c237 bl[237] br[237] wl[123] vdd gnd cell_6t
Xbit_r124_c237 bl[237] br[237] wl[124] vdd gnd cell_6t
Xbit_r125_c237 bl[237] br[237] wl[125] vdd gnd cell_6t
Xbit_r126_c237 bl[237] br[237] wl[126] vdd gnd cell_6t
Xbit_r127_c237 bl[237] br[237] wl[127] vdd gnd cell_6t
Xbit_r0_c238 bl[238] br[238] wl[0] vdd gnd cell_6t
Xbit_r1_c238 bl[238] br[238] wl[1] vdd gnd cell_6t
Xbit_r2_c238 bl[238] br[238] wl[2] vdd gnd cell_6t
Xbit_r3_c238 bl[238] br[238] wl[3] vdd gnd cell_6t
Xbit_r4_c238 bl[238] br[238] wl[4] vdd gnd cell_6t
Xbit_r5_c238 bl[238] br[238] wl[5] vdd gnd cell_6t
Xbit_r6_c238 bl[238] br[238] wl[6] vdd gnd cell_6t
Xbit_r7_c238 bl[238] br[238] wl[7] vdd gnd cell_6t
Xbit_r8_c238 bl[238] br[238] wl[8] vdd gnd cell_6t
Xbit_r9_c238 bl[238] br[238] wl[9] vdd gnd cell_6t
Xbit_r10_c238 bl[238] br[238] wl[10] vdd gnd cell_6t
Xbit_r11_c238 bl[238] br[238] wl[11] vdd gnd cell_6t
Xbit_r12_c238 bl[238] br[238] wl[12] vdd gnd cell_6t
Xbit_r13_c238 bl[238] br[238] wl[13] vdd gnd cell_6t
Xbit_r14_c238 bl[238] br[238] wl[14] vdd gnd cell_6t
Xbit_r15_c238 bl[238] br[238] wl[15] vdd gnd cell_6t
Xbit_r16_c238 bl[238] br[238] wl[16] vdd gnd cell_6t
Xbit_r17_c238 bl[238] br[238] wl[17] vdd gnd cell_6t
Xbit_r18_c238 bl[238] br[238] wl[18] vdd gnd cell_6t
Xbit_r19_c238 bl[238] br[238] wl[19] vdd gnd cell_6t
Xbit_r20_c238 bl[238] br[238] wl[20] vdd gnd cell_6t
Xbit_r21_c238 bl[238] br[238] wl[21] vdd gnd cell_6t
Xbit_r22_c238 bl[238] br[238] wl[22] vdd gnd cell_6t
Xbit_r23_c238 bl[238] br[238] wl[23] vdd gnd cell_6t
Xbit_r24_c238 bl[238] br[238] wl[24] vdd gnd cell_6t
Xbit_r25_c238 bl[238] br[238] wl[25] vdd gnd cell_6t
Xbit_r26_c238 bl[238] br[238] wl[26] vdd gnd cell_6t
Xbit_r27_c238 bl[238] br[238] wl[27] vdd gnd cell_6t
Xbit_r28_c238 bl[238] br[238] wl[28] vdd gnd cell_6t
Xbit_r29_c238 bl[238] br[238] wl[29] vdd gnd cell_6t
Xbit_r30_c238 bl[238] br[238] wl[30] vdd gnd cell_6t
Xbit_r31_c238 bl[238] br[238] wl[31] vdd gnd cell_6t
Xbit_r32_c238 bl[238] br[238] wl[32] vdd gnd cell_6t
Xbit_r33_c238 bl[238] br[238] wl[33] vdd gnd cell_6t
Xbit_r34_c238 bl[238] br[238] wl[34] vdd gnd cell_6t
Xbit_r35_c238 bl[238] br[238] wl[35] vdd gnd cell_6t
Xbit_r36_c238 bl[238] br[238] wl[36] vdd gnd cell_6t
Xbit_r37_c238 bl[238] br[238] wl[37] vdd gnd cell_6t
Xbit_r38_c238 bl[238] br[238] wl[38] vdd gnd cell_6t
Xbit_r39_c238 bl[238] br[238] wl[39] vdd gnd cell_6t
Xbit_r40_c238 bl[238] br[238] wl[40] vdd gnd cell_6t
Xbit_r41_c238 bl[238] br[238] wl[41] vdd gnd cell_6t
Xbit_r42_c238 bl[238] br[238] wl[42] vdd gnd cell_6t
Xbit_r43_c238 bl[238] br[238] wl[43] vdd gnd cell_6t
Xbit_r44_c238 bl[238] br[238] wl[44] vdd gnd cell_6t
Xbit_r45_c238 bl[238] br[238] wl[45] vdd gnd cell_6t
Xbit_r46_c238 bl[238] br[238] wl[46] vdd gnd cell_6t
Xbit_r47_c238 bl[238] br[238] wl[47] vdd gnd cell_6t
Xbit_r48_c238 bl[238] br[238] wl[48] vdd gnd cell_6t
Xbit_r49_c238 bl[238] br[238] wl[49] vdd gnd cell_6t
Xbit_r50_c238 bl[238] br[238] wl[50] vdd gnd cell_6t
Xbit_r51_c238 bl[238] br[238] wl[51] vdd gnd cell_6t
Xbit_r52_c238 bl[238] br[238] wl[52] vdd gnd cell_6t
Xbit_r53_c238 bl[238] br[238] wl[53] vdd gnd cell_6t
Xbit_r54_c238 bl[238] br[238] wl[54] vdd gnd cell_6t
Xbit_r55_c238 bl[238] br[238] wl[55] vdd gnd cell_6t
Xbit_r56_c238 bl[238] br[238] wl[56] vdd gnd cell_6t
Xbit_r57_c238 bl[238] br[238] wl[57] vdd gnd cell_6t
Xbit_r58_c238 bl[238] br[238] wl[58] vdd gnd cell_6t
Xbit_r59_c238 bl[238] br[238] wl[59] vdd gnd cell_6t
Xbit_r60_c238 bl[238] br[238] wl[60] vdd gnd cell_6t
Xbit_r61_c238 bl[238] br[238] wl[61] vdd gnd cell_6t
Xbit_r62_c238 bl[238] br[238] wl[62] vdd gnd cell_6t
Xbit_r63_c238 bl[238] br[238] wl[63] vdd gnd cell_6t
Xbit_r64_c238 bl[238] br[238] wl[64] vdd gnd cell_6t
Xbit_r65_c238 bl[238] br[238] wl[65] vdd gnd cell_6t
Xbit_r66_c238 bl[238] br[238] wl[66] vdd gnd cell_6t
Xbit_r67_c238 bl[238] br[238] wl[67] vdd gnd cell_6t
Xbit_r68_c238 bl[238] br[238] wl[68] vdd gnd cell_6t
Xbit_r69_c238 bl[238] br[238] wl[69] vdd gnd cell_6t
Xbit_r70_c238 bl[238] br[238] wl[70] vdd gnd cell_6t
Xbit_r71_c238 bl[238] br[238] wl[71] vdd gnd cell_6t
Xbit_r72_c238 bl[238] br[238] wl[72] vdd gnd cell_6t
Xbit_r73_c238 bl[238] br[238] wl[73] vdd gnd cell_6t
Xbit_r74_c238 bl[238] br[238] wl[74] vdd gnd cell_6t
Xbit_r75_c238 bl[238] br[238] wl[75] vdd gnd cell_6t
Xbit_r76_c238 bl[238] br[238] wl[76] vdd gnd cell_6t
Xbit_r77_c238 bl[238] br[238] wl[77] vdd gnd cell_6t
Xbit_r78_c238 bl[238] br[238] wl[78] vdd gnd cell_6t
Xbit_r79_c238 bl[238] br[238] wl[79] vdd gnd cell_6t
Xbit_r80_c238 bl[238] br[238] wl[80] vdd gnd cell_6t
Xbit_r81_c238 bl[238] br[238] wl[81] vdd gnd cell_6t
Xbit_r82_c238 bl[238] br[238] wl[82] vdd gnd cell_6t
Xbit_r83_c238 bl[238] br[238] wl[83] vdd gnd cell_6t
Xbit_r84_c238 bl[238] br[238] wl[84] vdd gnd cell_6t
Xbit_r85_c238 bl[238] br[238] wl[85] vdd gnd cell_6t
Xbit_r86_c238 bl[238] br[238] wl[86] vdd gnd cell_6t
Xbit_r87_c238 bl[238] br[238] wl[87] vdd gnd cell_6t
Xbit_r88_c238 bl[238] br[238] wl[88] vdd gnd cell_6t
Xbit_r89_c238 bl[238] br[238] wl[89] vdd gnd cell_6t
Xbit_r90_c238 bl[238] br[238] wl[90] vdd gnd cell_6t
Xbit_r91_c238 bl[238] br[238] wl[91] vdd gnd cell_6t
Xbit_r92_c238 bl[238] br[238] wl[92] vdd gnd cell_6t
Xbit_r93_c238 bl[238] br[238] wl[93] vdd gnd cell_6t
Xbit_r94_c238 bl[238] br[238] wl[94] vdd gnd cell_6t
Xbit_r95_c238 bl[238] br[238] wl[95] vdd gnd cell_6t
Xbit_r96_c238 bl[238] br[238] wl[96] vdd gnd cell_6t
Xbit_r97_c238 bl[238] br[238] wl[97] vdd gnd cell_6t
Xbit_r98_c238 bl[238] br[238] wl[98] vdd gnd cell_6t
Xbit_r99_c238 bl[238] br[238] wl[99] vdd gnd cell_6t
Xbit_r100_c238 bl[238] br[238] wl[100] vdd gnd cell_6t
Xbit_r101_c238 bl[238] br[238] wl[101] vdd gnd cell_6t
Xbit_r102_c238 bl[238] br[238] wl[102] vdd gnd cell_6t
Xbit_r103_c238 bl[238] br[238] wl[103] vdd gnd cell_6t
Xbit_r104_c238 bl[238] br[238] wl[104] vdd gnd cell_6t
Xbit_r105_c238 bl[238] br[238] wl[105] vdd gnd cell_6t
Xbit_r106_c238 bl[238] br[238] wl[106] vdd gnd cell_6t
Xbit_r107_c238 bl[238] br[238] wl[107] vdd gnd cell_6t
Xbit_r108_c238 bl[238] br[238] wl[108] vdd gnd cell_6t
Xbit_r109_c238 bl[238] br[238] wl[109] vdd gnd cell_6t
Xbit_r110_c238 bl[238] br[238] wl[110] vdd gnd cell_6t
Xbit_r111_c238 bl[238] br[238] wl[111] vdd gnd cell_6t
Xbit_r112_c238 bl[238] br[238] wl[112] vdd gnd cell_6t
Xbit_r113_c238 bl[238] br[238] wl[113] vdd gnd cell_6t
Xbit_r114_c238 bl[238] br[238] wl[114] vdd gnd cell_6t
Xbit_r115_c238 bl[238] br[238] wl[115] vdd gnd cell_6t
Xbit_r116_c238 bl[238] br[238] wl[116] vdd gnd cell_6t
Xbit_r117_c238 bl[238] br[238] wl[117] vdd gnd cell_6t
Xbit_r118_c238 bl[238] br[238] wl[118] vdd gnd cell_6t
Xbit_r119_c238 bl[238] br[238] wl[119] vdd gnd cell_6t
Xbit_r120_c238 bl[238] br[238] wl[120] vdd gnd cell_6t
Xbit_r121_c238 bl[238] br[238] wl[121] vdd gnd cell_6t
Xbit_r122_c238 bl[238] br[238] wl[122] vdd gnd cell_6t
Xbit_r123_c238 bl[238] br[238] wl[123] vdd gnd cell_6t
Xbit_r124_c238 bl[238] br[238] wl[124] vdd gnd cell_6t
Xbit_r125_c238 bl[238] br[238] wl[125] vdd gnd cell_6t
Xbit_r126_c238 bl[238] br[238] wl[126] vdd gnd cell_6t
Xbit_r127_c238 bl[238] br[238] wl[127] vdd gnd cell_6t
Xbit_r0_c239 bl[239] br[239] wl[0] vdd gnd cell_6t
Xbit_r1_c239 bl[239] br[239] wl[1] vdd gnd cell_6t
Xbit_r2_c239 bl[239] br[239] wl[2] vdd gnd cell_6t
Xbit_r3_c239 bl[239] br[239] wl[3] vdd gnd cell_6t
Xbit_r4_c239 bl[239] br[239] wl[4] vdd gnd cell_6t
Xbit_r5_c239 bl[239] br[239] wl[5] vdd gnd cell_6t
Xbit_r6_c239 bl[239] br[239] wl[6] vdd gnd cell_6t
Xbit_r7_c239 bl[239] br[239] wl[7] vdd gnd cell_6t
Xbit_r8_c239 bl[239] br[239] wl[8] vdd gnd cell_6t
Xbit_r9_c239 bl[239] br[239] wl[9] vdd gnd cell_6t
Xbit_r10_c239 bl[239] br[239] wl[10] vdd gnd cell_6t
Xbit_r11_c239 bl[239] br[239] wl[11] vdd gnd cell_6t
Xbit_r12_c239 bl[239] br[239] wl[12] vdd gnd cell_6t
Xbit_r13_c239 bl[239] br[239] wl[13] vdd gnd cell_6t
Xbit_r14_c239 bl[239] br[239] wl[14] vdd gnd cell_6t
Xbit_r15_c239 bl[239] br[239] wl[15] vdd gnd cell_6t
Xbit_r16_c239 bl[239] br[239] wl[16] vdd gnd cell_6t
Xbit_r17_c239 bl[239] br[239] wl[17] vdd gnd cell_6t
Xbit_r18_c239 bl[239] br[239] wl[18] vdd gnd cell_6t
Xbit_r19_c239 bl[239] br[239] wl[19] vdd gnd cell_6t
Xbit_r20_c239 bl[239] br[239] wl[20] vdd gnd cell_6t
Xbit_r21_c239 bl[239] br[239] wl[21] vdd gnd cell_6t
Xbit_r22_c239 bl[239] br[239] wl[22] vdd gnd cell_6t
Xbit_r23_c239 bl[239] br[239] wl[23] vdd gnd cell_6t
Xbit_r24_c239 bl[239] br[239] wl[24] vdd gnd cell_6t
Xbit_r25_c239 bl[239] br[239] wl[25] vdd gnd cell_6t
Xbit_r26_c239 bl[239] br[239] wl[26] vdd gnd cell_6t
Xbit_r27_c239 bl[239] br[239] wl[27] vdd gnd cell_6t
Xbit_r28_c239 bl[239] br[239] wl[28] vdd gnd cell_6t
Xbit_r29_c239 bl[239] br[239] wl[29] vdd gnd cell_6t
Xbit_r30_c239 bl[239] br[239] wl[30] vdd gnd cell_6t
Xbit_r31_c239 bl[239] br[239] wl[31] vdd gnd cell_6t
Xbit_r32_c239 bl[239] br[239] wl[32] vdd gnd cell_6t
Xbit_r33_c239 bl[239] br[239] wl[33] vdd gnd cell_6t
Xbit_r34_c239 bl[239] br[239] wl[34] vdd gnd cell_6t
Xbit_r35_c239 bl[239] br[239] wl[35] vdd gnd cell_6t
Xbit_r36_c239 bl[239] br[239] wl[36] vdd gnd cell_6t
Xbit_r37_c239 bl[239] br[239] wl[37] vdd gnd cell_6t
Xbit_r38_c239 bl[239] br[239] wl[38] vdd gnd cell_6t
Xbit_r39_c239 bl[239] br[239] wl[39] vdd gnd cell_6t
Xbit_r40_c239 bl[239] br[239] wl[40] vdd gnd cell_6t
Xbit_r41_c239 bl[239] br[239] wl[41] vdd gnd cell_6t
Xbit_r42_c239 bl[239] br[239] wl[42] vdd gnd cell_6t
Xbit_r43_c239 bl[239] br[239] wl[43] vdd gnd cell_6t
Xbit_r44_c239 bl[239] br[239] wl[44] vdd gnd cell_6t
Xbit_r45_c239 bl[239] br[239] wl[45] vdd gnd cell_6t
Xbit_r46_c239 bl[239] br[239] wl[46] vdd gnd cell_6t
Xbit_r47_c239 bl[239] br[239] wl[47] vdd gnd cell_6t
Xbit_r48_c239 bl[239] br[239] wl[48] vdd gnd cell_6t
Xbit_r49_c239 bl[239] br[239] wl[49] vdd gnd cell_6t
Xbit_r50_c239 bl[239] br[239] wl[50] vdd gnd cell_6t
Xbit_r51_c239 bl[239] br[239] wl[51] vdd gnd cell_6t
Xbit_r52_c239 bl[239] br[239] wl[52] vdd gnd cell_6t
Xbit_r53_c239 bl[239] br[239] wl[53] vdd gnd cell_6t
Xbit_r54_c239 bl[239] br[239] wl[54] vdd gnd cell_6t
Xbit_r55_c239 bl[239] br[239] wl[55] vdd gnd cell_6t
Xbit_r56_c239 bl[239] br[239] wl[56] vdd gnd cell_6t
Xbit_r57_c239 bl[239] br[239] wl[57] vdd gnd cell_6t
Xbit_r58_c239 bl[239] br[239] wl[58] vdd gnd cell_6t
Xbit_r59_c239 bl[239] br[239] wl[59] vdd gnd cell_6t
Xbit_r60_c239 bl[239] br[239] wl[60] vdd gnd cell_6t
Xbit_r61_c239 bl[239] br[239] wl[61] vdd gnd cell_6t
Xbit_r62_c239 bl[239] br[239] wl[62] vdd gnd cell_6t
Xbit_r63_c239 bl[239] br[239] wl[63] vdd gnd cell_6t
Xbit_r64_c239 bl[239] br[239] wl[64] vdd gnd cell_6t
Xbit_r65_c239 bl[239] br[239] wl[65] vdd gnd cell_6t
Xbit_r66_c239 bl[239] br[239] wl[66] vdd gnd cell_6t
Xbit_r67_c239 bl[239] br[239] wl[67] vdd gnd cell_6t
Xbit_r68_c239 bl[239] br[239] wl[68] vdd gnd cell_6t
Xbit_r69_c239 bl[239] br[239] wl[69] vdd gnd cell_6t
Xbit_r70_c239 bl[239] br[239] wl[70] vdd gnd cell_6t
Xbit_r71_c239 bl[239] br[239] wl[71] vdd gnd cell_6t
Xbit_r72_c239 bl[239] br[239] wl[72] vdd gnd cell_6t
Xbit_r73_c239 bl[239] br[239] wl[73] vdd gnd cell_6t
Xbit_r74_c239 bl[239] br[239] wl[74] vdd gnd cell_6t
Xbit_r75_c239 bl[239] br[239] wl[75] vdd gnd cell_6t
Xbit_r76_c239 bl[239] br[239] wl[76] vdd gnd cell_6t
Xbit_r77_c239 bl[239] br[239] wl[77] vdd gnd cell_6t
Xbit_r78_c239 bl[239] br[239] wl[78] vdd gnd cell_6t
Xbit_r79_c239 bl[239] br[239] wl[79] vdd gnd cell_6t
Xbit_r80_c239 bl[239] br[239] wl[80] vdd gnd cell_6t
Xbit_r81_c239 bl[239] br[239] wl[81] vdd gnd cell_6t
Xbit_r82_c239 bl[239] br[239] wl[82] vdd gnd cell_6t
Xbit_r83_c239 bl[239] br[239] wl[83] vdd gnd cell_6t
Xbit_r84_c239 bl[239] br[239] wl[84] vdd gnd cell_6t
Xbit_r85_c239 bl[239] br[239] wl[85] vdd gnd cell_6t
Xbit_r86_c239 bl[239] br[239] wl[86] vdd gnd cell_6t
Xbit_r87_c239 bl[239] br[239] wl[87] vdd gnd cell_6t
Xbit_r88_c239 bl[239] br[239] wl[88] vdd gnd cell_6t
Xbit_r89_c239 bl[239] br[239] wl[89] vdd gnd cell_6t
Xbit_r90_c239 bl[239] br[239] wl[90] vdd gnd cell_6t
Xbit_r91_c239 bl[239] br[239] wl[91] vdd gnd cell_6t
Xbit_r92_c239 bl[239] br[239] wl[92] vdd gnd cell_6t
Xbit_r93_c239 bl[239] br[239] wl[93] vdd gnd cell_6t
Xbit_r94_c239 bl[239] br[239] wl[94] vdd gnd cell_6t
Xbit_r95_c239 bl[239] br[239] wl[95] vdd gnd cell_6t
Xbit_r96_c239 bl[239] br[239] wl[96] vdd gnd cell_6t
Xbit_r97_c239 bl[239] br[239] wl[97] vdd gnd cell_6t
Xbit_r98_c239 bl[239] br[239] wl[98] vdd gnd cell_6t
Xbit_r99_c239 bl[239] br[239] wl[99] vdd gnd cell_6t
Xbit_r100_c239 bl[239] br[239] wl[100] vdd gnd cell_6t
Xbit_r101_c239 bl[239] br[239] wl[101] vdd gnd cell_6t
Xbit_r102_c239 bl[239] br[239] wl[102] vdd gnd cell_6t
Xbit_r103_c239 bl[239] br[239] wl[103] vdd gnd cell_6t
Xbit_r104_c239 bl[239] br[239] wl[104] vdd gnd cell_6t
Xbit_r105_c239 bl[239] br[239] wl[105] vdd gnd cell_6t
Xbit_r106_c239 bl[239] br[239] wl[106] vdd gnd cell_6t
Xbit_r107_c239 bl[239] br[239] wl[107] vdd gnd cell_6t
Xbit_r108_c239 bl[239] br[239] wl[108] vdd gnd cell_6t
Xbit_r109_c239 bl[239] br[239] wl[109] vdd gnd cell_6t
Xbit_r110_c239 bl[239] br[239] wl[110] vdd gnd cell_6t
Xbit_r111_c239 bl[239] br[239] wl[111] vdd gnd cell_6t
Xbit_r112_c239 bl[239] br[239] wl[112] vdd gnd cell_6t
Xbit_r113_c239 bl[239] br[239] wl[113] vdd gnd cell_6t
Xbit_r114_c239 bl[239] br[239] wl[114] vdd gnd cell_6t
Xbit_r115_c239 bl[239] br[239] wl[115] vdd gnd cell_6t
Xbit_r116_c239 bl[239] br[239] wl[116] vdd gnd cell_6t
Xbit_r117_c239 bl[239] br[239] wl[117] vdd gnd cell_6t
Xbit_r118_c239 bl[239] br[239] wl[118] vdd gnd cell_6t
Xbit_r119_c239 bl[239] br[239] wl[119] vdd gnd cell_6t
Xbit_r120_c239 bl[239] br[239] wl[120] vdd gnd cell_6t
Xbit_r121_c239 bl[239] br[239] wl[121] vdd gnd cell_6t
Xbit_r122_c239 bl[239] br[239] wl[122] vdd gnd cell_6t
Xbit_r123_c239 bl[239] br[239] wl[123] vdd gnd cell_6t
Xbit_r124_c239 bl[239] br[239] wl[124] vdd gnd cell_6t
Xbit_r125_c239 bl[239] br[239] wl[125] vdd gnd cell_6t
Xbit_r126_c239 bl[239] br[239] wl[126] vdd gnd cell_6t
Xbit_r127_c239 bl[239] br[239] wl[127] vdd gnd cell_6t
Xbit_r0_c240 bl[240] br[240] wl[0] vdd gnd cell_6t
Xbit_r1_c240 bl[240] br[240] wl[1] vdd gnd cell_6t
Xbit_r2_c240 bl[240] br[240] wl[2] vdd gnd cell_6t
Xbit_r3_c240 bl[240] br[240] wl[3] vdd gnd cell_6t
Xbit_r4_c240 bl[240] br[240] wl[4] vdd gnd cell_6t
Xbit_r5_c240 bl[240] br[240] wl[5] vdd gnd cell_6t
Xbit_r6_c240 bl[240] br[240] wl[6] vdd gnd cell_6t
Xbit_r7_c240 bl[240] br[240] wl[7] vdd gnd cell_6t
Xbit_r8_c240 bl[240] br[240] wl[8] vdd gnd cell_6t
Xbit_r9_c240 bl[240] br[240] wl[9] vdd gnd cell_6t
Xbit_r10_c240 bl[240] br[240] wl[10] vdd gnd cell_6t
Xbit_r11_c240 bl[240] br[240] wl[11] vdd gnd cell_6t
Xbit_r12_c240 bl[240] br[240] wl[12] vdd gnd cell_6t
Xbit_r13_c240 bl[240] br[240] wl[13] vdd gnd cell_6t
Xbit_r14_c240 bl[240] br[240] wl[14] vdd gnd cell_6t
Xbit_r15_c240 bl[240] br[240] wl[15] vdd gnd cell_6t
Xbit_r16_c240 bl[240] br[240] wl[16] vdd gnd cell_6t
Xbit_r17_c240 bl[240] br[240] wl[17] vdd gnd cell_6t
Xbit_r18_c240 bl[240] br[240] wl[18] vdd gnd cell_6t
Xbit_r19_c240 bl[240] br[240] wl[19] vdd gnd cell_6t
Xbit_r20_c240 bl[240] br[240] wl[20] vdd gnd cell_6t
Xbit_r21_c240 bl[240] br[240] wl[21] vdd gnd cell_6t
Xbit_r22_c240 bl[240] br[240] wl[22] vdd gnd cell_6t
Xbit_r23_c240 bl[240] br[240] wl[23] vdd gnd cell_6t
Xbit_r24_c240 bl[240] br[240] wl[24] vdd gnd cell_6t
Xbit_r25_c240 bl[240] br[240] wl[25] vdd gnd cell_6t
Xbit_r26_c240 bl[240] br[240] wl[26] vdd gnd cell_6t
Xbit_r27_c240 bl[240] br[240] wl[27] vdd gnd cell_6t
Xbit_r28_c240 bl[240] br[240] wl[28] vdd gnd cell_6t
Xbit_r29_c240 bl[240] br[240] wl[29] vdd gnd cell_6t
Xbit_r30_c240 bl[240] br[240] wl[30] vdd gnd cell_6t
Xbit_r31_c240 bl[240] br[240] wl[31] vdd gnd cell_6t
Xbit_r32_c240 bl[240] br[240] wl[32] vdd gnd cell_6t
Xbit_r33_c240 bl[240] br[240] wl[33] vdd gnd cell_6t
Xbit_r34_c240 bl[240] br[240] wl[34] vdd gnd cell_6t
Xbit_r35_c240 bl[240] br[240] wl[35] vdd gnd cell_6t
Xbit_r36_c240 bl[240] br[240] wl[36] vdd gnd cell_6t
Xbit_r37_c240 bl[240] br[240] wl[37] vdd gnd cell_6t
Xbit_r38_c240 bl[240] br[240] wl[38] vdd gnd cell_6t
Xbit_r39_c240 bl[240] br[240] wl[39] vdd gnd cell_6t
Xbit_r40_c240 bl[240] br[240] wl[40] vdd gnd cell_6t
Xbit_r41_c240 bl[240] br[240] wl[41] vdd gnd cell_6t
Xbit_r42_c240 bl[240] br[240] wl[42] vdd gnd cell_6t
Xbit_r43_c240 bl[240] br[240] wl[43] vdd gnd cell_6t
Xbit_r44_c240 bl[240] br[240] wl[44] vdd gnd cell_6t
Xbit_r45_c240 bl[240] br[240] wl[45] vdd gnd cell_6t
Xbit_r46_c240 bl[240] br[240] wl[46] vdd gnd cell_6t
Xbit_r47_c240 bl[240] br[240] wl[47] vdd gnd cell_6t
Xbit_r48_c240 bl[240] br[240] wl[48] vdd gnd cell_6t
Xbit_r49_c240 bl[240] br[240] wl[49] vdd gnd cell_6t
Xbit_r50_c240 bl[240] br[240] wl[50] vdd gnd cell_6t
Xbit_r51_c240 bl[240] br[240] wl[51] vdd gnd cell_6t
Xbit_r52_c240 bl[240] br[240] wl[52] vdd gnd cell_6t
Xbit_r53_c240 bl[240] br[240] wl[53] vdd gnd cell_6t
Xbit_r54_c240 bl[240] br[240] wl[54] vdd gnd cell_6t
Xbit_r55_c240 bl[240] br[240] wl[55] vdd gnd cell_6t
Xbit_r56_c240 bl[240] br[240] wl[56] vdd gnd cell_6t
Xbit_r57_c240 bl[240] br[240] wl[57] vdd gnd cell_6t
Xbit_r58_c240 bl[240] br[240] wl[58] vdd gnd cell_6t
Xbit_r59_c240 bl[240] br[240] wl[59] vdd gnd cell_6t
Xbit_r60_c240 bl[240] br[240] wl[60] vdd gnd cell_6t
Xbit_r61_c240 bl[240] br[240] wl[61] vdd gnd cell_6t
Xbit_r62_c240 bl[240] br[240] wl[62] vdd gnd cell_6t
Xbit_r63_c240 bl[240] br[240] wl[63] vdd gnd cell_6t
Xbit_r64_c240 bl[240] br[240] wl[64] vdd gnd cell_6t
Xbit_r65_c240 bl[240] br[240] wl[65] vdd gnd cell_6t
Xbit_r66_c240 bl[240] br[240] wl[66] vdd gnd cell_6t
Xbit_r67_c240 bl[240] br[240] wl[67] vdd gnd cell_6t
Xbit_r68_c240 bl[240] br[240] wl[68] vdd gnd cell_6t
Xbit_r69_c240 bl[240] br[240] wl[69] vdd gnd cell_6t
Xbit_r70_c240 bl[240] br[240] wl[70] vdd gnd cell_6t
Xbit_r71_c240 bl[240] br[240] wl[71] vdd gnd cell_6t
Xbit_r72_c240 bl[240] br[240] wl[72] vdd gnd cell_6t
Xbit_r73_c240 bl[240] br[240] wl[73] vdd gnd cell_6t
Xbit_r74_c240 bl[240] br[240] wl[74] vdd gnd cell_6t
Xbit_r75_c240 bl[240] br[240] wl[75] vdd gnd cell_6t
Xbit_r76_c240 bl[240] br[240] wl[76] vdd gnd cell_6t
Xbit_r77_c240 bl[240] br[240] wl[77] vdd gnd cell_6t
Xbit_r78_c240 bl[240] br[240] wl[78] vdd gnd cell_6t
Xbit_r79_c240 bl[240] br[240] wl[79] vdd gnd cell_6t
Xbit_r80_c240 bl[240] br[240] wl[80] vdd gnd cell_6t
Xbit_r81_c240 bl[240] br[240] wl[81] vdd gnd cell_6t
Xbit_r82_c240 bl[240] br[240] wl[82] vdd gnd cell_6t
Xbit_r83_c240 bl[240] br[240] wl[83] vdd gnd cell_6t
Xbit_r84_c240 bl[240] br[240] wl[84] vdd gnd cell_6t
Xbit_r85_c240 bl[240] br[240] wl[85] vdd gnd cell_6t
Xbit_r86_c240 bl[240] br[240] wl[86] vdd gnd cell_6t
Xbit_r87_c240 bl[240] br[240] wl[87] vdd gnd cell_6t
Xbit_r88_c240 bl[240] br[240] wl[88] vdd gnd cell_6t
Xbit_r89_c240 bl[240] br[240] wl[89] vdd gnd cell_6t
Xbit_r90_c240 bl[240] br[240] wl[90] vdd gnd cell_6t
Xbit_r91_c240 bl[240] br[240] wl[91] vdd gnd cell_6t
Xbit_r92_c240 bl[240] br[240] wl[92] vdd gnd cell_6t
Xbit_r93_c240 bl[240] br[240] wl[93] vdd gnd cell_6t
Xbit_r94_c240 bl[240] br[240] wl[94] vdd gnd cell_6t
Xbit_r95_c240 bl[240] br[240] wl[95] vdd gnd cell_6t
Xbit_r96_c240 bl[240] br[240] wl[96] vdd gnd cell_6t
Xbit_r97_c240 bl[240] br[240] wl[97] vdd gnd cell_6t
Xbit_r98_c240 bl[240] br[240] wl[98] vdd gnd cell_6t
Xbit_r99_c240 bl[240] br[240] wl[99] vdd gnd cell_6t
Xbit_r100_c240 bl[240] br[240] wl[100] vdd gnd cell_6t
Xbit_r101_c240 bl[240] br[240] wl[101] vdd gnd cell_6t
Xbit_r102_c240 bl[240] br[240] wl[102] vdd gnd cell_6t
Xbit_r103_c240 bl[240] br[240] wl[103] vdd gnd cell_6t
Xbit_r104_c240 bl[240] br[240] wl[104] vdd gnd cell_6t
Xbit_r105_c240 bl[240] br[240] wl[105] vdd gnd cell_6t
Xbit_r106_c240 bl[240] br[240] wl[106] vdd gnd cell_6t
Xbit_r107_c240 bl[240] br[240] wl[107] vdd gnd cell_6t
Xbit_r108_c240 bl[240] br[240] wl[108] vdd gnd cell_6t
Xbit_r109_c240 bl[240] br[240] wl[109] vdd gnd cell_6t
Xbit_r110_c240 bl[240] br[240] wl[110] vdd gnd cell_6t
Xbit_r111_c240 bl[240] br[240] wl[111] vdd gnd cell_6t
Xbit_r112_c240 bl[240] br[240] wl[112] vdd gnd cell_6t
Xbit_r113_c240 bl[240] br[240] wl[113] vdd gnd cell_6t
Xbit_r114_c240 bl[240] br[240] wl[114] vdd gnd cell_6t
Xbit_r115_c240 bl[240] br[240] wl[115] vdd gnd cell_6t
Xbit_r116_c240 bl[240] br[240] wl[116] vdd gnd cell_6t
Xbit_r117_c240 bl[240] br[240] wl[117] vdd gnd cell_6t
Xbit_r118_c240 bl[240] br[240] wl[118] vdd gnd cell_6t
Xbit_r119_c240 bl[240] br[240] wl[119] vdd gnd cell_6t
Xbit_r120_c240 bl[240] br[240] wl[120] vdd gnd cell_6t
Xbit_r121_c240 bl[240] br[240] wl[121] vdd gnd cell_6t
Xbit_r122_c240 bl[240] br[240] wl[122] vdd gnd cell_6t
Xbit_r123_c240 bl[240] br[240] wl[123] vdd gnd cell_6t
Xbit_r124_c240 bl[240] br[240] wl[124] vdd gnd cell_6t
Xbit_r125_c240 bl[240] br[240] wl[125] vdd gnd cell_6t
Xbit_r126_c240 bl[240] br[240] wl[126] vdd gnd cell_6t
Xbit_r127_c240 bl[240] br[240] wl[127] vdd gnd cell_6t
Xbit_r0_c241 bl[241] br[241] wl[0] vdd gnd cell_6t
Xbit_r1_c241 bl[241] br[241] wl[1] vdd gnd cell_6t
Xbit_r2_c241 bl[241] br[241] wl[2] vdd gnd cell_6t
Xbit_r3_c241 bl[241] br[241] wl[3] vdd gnd cell_6t
Xbit_r4_c241 bl[241] br[241] wl[4] vdd gnd cell_6t
Xbit_r5_c241 bl[241] br[241] wl[5] vdd gnd cell_6t
Xbit_r6_c241 bl[241] br[241] wl[6] vdd gnd cell_6t
Xbit_r7_c241 bl[241] br[241] wl[7] vdd gnd cell_6t
Xbit_r8_c241 bl[241] br[241] wl[8] vdd gnd cell_6t
Xbit_r9_c241 bl[241] br[241] wl[9] vdd gnd cell_6t
Xbit_r10_c241 bl[241] br[241] wl[10] vdd gnd cell_6t
Xbit_r11_c241 bl[241] br[241] wl[11] vdd gnd cell_6t
Xbit_r12_c241 bl[241] br[241] wl[12] vdd gnd cell_6t
Xbit_r13_c241 bl[241] br[241] wl[13] vdd gnd cell_6t
Xbit_r14_c241 bl[241] br[241] wl[14] vdd gnd cell_6t
Xbit_r15_c241 bl[241] br[241] wl[15] vdd gnd cell_6t
Xbit_r16_c241 bl[241] br[241] wl[16] vdd gnd cell_6t
Xbit_r17_c241 bl[241] br[241] wl[17] vdd gnd cell_6t
Xbit_r18_c241 bl[241] br[241] wl[18] vdd gnd cell_6t
Xbit_r19_c241 bl[241] br[241] wl[19] vdd gnd cell_6t
Xbit_r20_c241 bl[241] br[241] wl[20] vdd gnd cell_6t
Xbit_r21_c241 bl[241] br[241] wl[21] vdd gnd cell_6t
Xbit_r22_c241 bl[241] br[241] wl[22] vdd gnd cell_6t
Xbit_r23_c241 bl[241] br[241] wl[23] vdd gnd cell_6t
Xbit_r24_c241 bl[241] br[241] wl[24] vdd gnd cell_6t
Xbit_r25_c241 bl[241] br[241] wl[25] vdd gnd cell_6t
Xbit_r26_c241 bl[241] br[241] wl[26] vdd gnd cell_6t
Xbit_r27_c241 bl[241] br[241] wl[27] vdd gnd cell_6t
Xbit_r28_c241 bl[241] br[241] wl[28] vdd gnd cell_6t
Xbit_r29_c241 bl[241] br[241] wl[29] vdd gnd cell_6t
Xbit_r30_c241 bl[241] br[241] wl[30] vdd gnd cell_6t
Xbit_r31_c241 bl[241] br[241] wl[31] vdd gnd cell_6t
Xbit_r32_c241 bl[241] br[241] wl[32] vdd gnd cell_6t
Xbit_r33_c241 bl[241] br[241] wl[33] vdd gnd cell_6t
Xbit_r34_c241 bl[241] br[241] wl[34] vdd gnd cell_6t
Xbit_r35_c241 bl[241] br[241] wl[35] vdd gnd cell_6t
Xbit_r36_c241 bl[241] br[241] wl[36] vdd gnd cell_6t
Xbit_r37_c241 bl[241] br[241] wl[37] vdd gnd cell_6t
Xbit_r38_c241 bl[241] br[241] wl[38] vdd gnd cell_6t
Xbit_r39_c241 bl[241] br[241] wl[39] vdd gnd cell_6t
Xbit_r40_c241 bl[241] br[241] wl[40] vdd gnd cell_6t
Xbit_r41_c241 bl[241] br[241] wl[41] vdd gnd cell_6t
Xbit_r42_c241 bl[241] br[241] wl[42] vdd gnd cell_6t
Xbit_r43_c241 bl[241] br[241] wl[43] vdd gnd cell_6t
Xbit_r44_c241 bl[241] br[241] wl[44] vdd gnd cell_6t
Xbit_r45_c241 bl[241] br[241] wl[45] vdd gnd cell_6t
Xbit_r46_c241 bl[241] br[241] wl[46] vdd gnd cell_6t
Xbit_r47_c241 bl[241] br[241] wl[47] vdd gnd cell_6t
Xbit_r48_c241 bl[241] br[241] wl[48] vdd gnd cell_6t
Xbit_r49_c241 bl[241] br[241] wl[49] vdd gnd cell_6t
Xbit_r50_c241 bl[241] br[241] wl[50] vdd gnd cell_6t
Xbit_r51_c241 bl[241] br[241] wl[51] vdd gnd cell_6t
Xbit_r52_c241 bl[241] br[241] wl[52] vdd gnd cell_6t
Xbit_r53_c241 bl[241] br[241] wl[53] vdd gnd cell_6t
Xbit_r54_c241 bl[241] br[241] wl[54] vdd gnd cell_6t
Xbit_r55_c241 bl[241] br[241] wl[55] vdd gnd cell_6t
Xbit_r56_c241 bl[241] br[241] wl[56] vdd gnd cell_6t
Xbit_r57_c241 bl[241] br[241] wl[57] vdd gnd cell_6t
Xbit_r58_c241 bl[241] br[241] wl[58] vdd gnd cell_6t
Xbit_r59_c241 bl[241] br[241] wl[59] vdd gnd cell_6t
Xbit_r60_c241 bl[241] br[241] wl[60] vdd gnd cell_6t
Xbit_r61_c241 bl[241] br[241] wl[61] vdd gnd cell_6t
Xbit_r62_c241 bl[241] br[241] wl[62] vdd gnd cell_6t
Xbit_r63_c241 bl[241] br[241] wl[63] vdd gnd cell_6t
Xbit_r64_c241 bl[241] br[241] wl[64] vdd gnd cell_6t
Xbit_r65_c241 bl[241] br[241] wl[65] vdd gnd cell_6t
Xbit_r66_c241 bl[241] br[241] wl[66] vdd gnd cell_6t
Xbit_r67_c241 bl[241] br[241] wl[67] vdd gnd cell_6t
Xbit_r68_c241 bl[241] br[241] wl[68] vdd gnd cell_6t
Xbit_r69_c241 bl[241] br[241] wl[69] vdd gnd cell_6t
Xbit_r70_c241 bl[241] br[241] wl[70] vdd gnd cell_6t
Xbit_r71_c241 bl[241] br[241] wl[71] vdd gnd cell_6t
Xbit_r72_c241 bl[241] br[241] wl[72] vdd gnd cell_6t
Xbit_r73_c241 bl[241] br[241] wl[73] vdd gnd cell_6t
Xbit_r74_c241 bl[241] br[241] wl[74] vdd gnd cell_6t
Xbit_r75_c241 bl[241] br[241] wl[75] vdd gnd cell_6t
Xbit_r76_c241 bl[241] br[241] wl[76] vdd gnd cell_6t
Xbit_r77_c241 bl[241] br[241] wl[77] vdd gnd cell_6t
Xbit_r78_c241 bl[241] br[241] wl[78] vdd gnd cell_6t
Xbit_r79_c241 bl[241] br[241] wl[79] vdd gnd cell_6t
Xbit_r80_c241 bl[241] br[241] wl[80] vdd gnd cell_6t
Xbit_r81_c241 bl[241] br[241] wl[81] vdd gnd cell_6t
Xbit_r82_c241 bl[241] br[241] wl[82] vdd gnd cell_6t
Xbit_r83_c241 bl[241] br[241] wl[83] vdd gnd cell_6t
Xbit_r84_c241 bl[241] br[241] wl[84] vdd gnd cell_6t
Xbit_r85_c241 bl[241] br[241] wl[85] vdd gnd cell_6t
Xbit_r86_c241 bl[241] br[241] wl[86] vdd gnd cell_6t
Xbit_r87_c241 bl[241] br[241] wl[87] vdd gnd cell_6t
Xbit_r88_c241 bl[241] br[241] wl[88] vdd gnd cell_6t
Xbit_r89_c241 bl[241] br[241] wl[89] vdd gnd cell_6t
Xbit_r90_c241 bl[241] br[241] wl[90] vdd gnd cell_6t
Xbit_r91_c241 bl[241] br[241] wl[91] vdd gnd cell_6t
Xbit_r92_c241 bl[241] br[241] wl[92] vdd gnd cell_6t
Xbit_r93_c241 bl[241] br[241] wl[93] vdd gnd cell_6t
Xbit_r94_c241 bl[241] br[241] wl[94] vdd gnd cell_6t
Xbit_r95_c241 bl[241] br[241] wl[95] vdd gnd cell_6t
Xbit_r96_c241 bl[241] br[241] wl[96] vdd gnd cell_6t
Xbit_r97_c241 bl[241] br[241] wl[97] vdd gnd cell_6t
Xbit_r98_c241 bl[241] br[241] wl[98] vdd gnd cell_6t
Xbit_r99_c241 bl[241] br[241] wl[99] vdd gnd cell_6t
Xbit_r100_c241 bl[241] br[241] wl[100] vdd gnd cell_6t
Xbit_r101_c241 bl[241] br[241] wl[101] vdd gnd cell_6t
Xbit_r102_c241 bl[241] br[241] wl[102] vdd gnd cell_6t
Xbit_r103_c241 bl[241] br[241] wl[103] vdd gnd cell_6t
Xbit_r104_c241 bl[241] br[241] wl[104] vdd gnd cell_6t
Xbit_r105_c241 bl[241] br[241] wl[105] vdd gnd cell_6t
Xbit_r106_c241 bl[241] br[241] wl[106] vdd gnd cell_6t
Xbit_r107_c241 bl[241] br[241] wl[107] vdd gnd cell_6t
Xbit_r108_c241 bl[241] br[241] wl[108] vdd gnd cell_6t
Xbit_r109_c241 bl[241] br[241] wl[109] vdd gnd cell_6t
Xbit_r110_c241 bl[241] br[241] wl[110] vdd gnd cell_6t
Xbit_r111_c241 bl[241] br[241] wl[111] vdd gnd cell_6t
Xbit_r112_c241 bl[241] br[241] wl[112] vdd gnd cell_6t
Xbit_r113_c241 bl[241] br[241] wl[113] vdd gnd cell_6t
Xbit_r114_c241 bl[241] br[241] wl[114] vdd gnd cell_6t
Xbit_r115_c241 bl[241] br[241] wl[115] vdd gnd cell_6t
Xbit_r116_c241 bl[241] br[241] wl[116] vdd gnd cell_6t
Xbit_r117_c241 bl[241] br[241] wl[117] vdd gnd cell_6t
Xbit_r118_c241 bl[241] br[241] wl[118] vdd gnd cell_6t
Xbit_r119_c241 bl[241] br[241] wl[119] vdd gnd cell_6t
Xbit_r120_c241 bl[241] br[241] wl[120] vdd gnd cell_6t
Xbit_r121_c241 bl[241] br[241] wl[121] vdd gnd cell_6t
Xbit_r122_c241 bl[241] br[241] wl[122] vdd gnd cell_6t
Xbit_r123_c241 bl[241] br[241] wl[123] vdd gnd cell_6t
Xbit_r124_c241 bl[241] br[241] wl[124] vdd gnd cell_6t
Xbit_r125_c241 bl[241] br[241] wl[125] vdd gnd cell_6t
Xbit_r126_c241 bl[241] br[241] wl[126] vdd gnd cell_6t
Xbit_r127_c241 bl[241] br[241] wl[127] vdd gnd cell_6t
Xbit_r0_c242 bl[242] br[242] wl[0] vdd gnd cell_6t
Xbit_r1_c242 bl[242] br[242] wl[1] vdd gnd cell_6t
Xbit_r2_c242 bl[242] br[242] wl[2] vdd gnd cell_6t
Xbit_r3_c242 bl[242] br[242] wl[3] vdd gnd cell_6t
Xbit_r4_c242 bl[242] br[242] wl[4] vdd gnd cell_6t
Xbit_r5_c242 bl[242] br[242] wl[5] vdd gnd cell_6t
Xbit_r6_c242 bl[242] br[242] wl[6] vdd gnd cell_6t
Xbit_r7_c242 bl[242] br[242] wl[7] vdd gnd cell_6t
Xbit_r8_c242 bl[242] br[242] wl[8] vdd gnd cell_6t
Xbit_r9_c242 bl[242] br[242] wl[9] vdd gnd cell_6t
Xbit_r10_c242 bl[242] br[242] wl[10] vdd gnd cell_6t
Xbit_r11_c242 bl[242] br[242] wl[11] vdd gnd cell_6t
Xbit_r12_c242 bl[242] br[242] wl[12] vdd gnd cell_6t
Xbit_r13_c242 bl[242] br[242] wl[13] vdd gnd cell_6t
Xbit_r14_c242 bl[242] br[242] wl[14] vdd gnd cell_6t
Xbit_r15_c242 bl[242] br[242] wl[15] vdd gnd cell_6t
Xbit_r16_c242 bl[242] br[242] wl[16] vdd gnd cell_6t
Xbit_r17_c242 bl[242] br[242] wl[17] vdd gnd cell_6t
Xbit_r18_c242 bl[242] br[242] wl[18] vdd gnd cell_6t
Xbit_r19_c242 bl[242] br[242] wl[19] vdd gnd cell_6t
Xbit_r20_c242 bl[242] br[242] wl[20] vdd gnd cell_6t
Xbit_r21_c242 bl[242] br[242] wl[21] vdd gnd cell_6t
Xbit_r22_c242 bl[242] br[242] wl[22] vdd gnd cell_6t
Xbit_r23_c242 bl[242] br[242] wl[23] vdd gnd cell_6t
Xbit_r24_c242 bl[242] br[242] wl[24] vdd gnd cell_6t
Xbit_r25_c242 bl[242] br[242] wl[25] vdd gnd cell_6t
Xbit_r26_c242 bl[242] br[242] wl[26] vdd gnd cell_6t
Xbit_r27_c242 bl[242] br[242] wl[27] vdd gnd cell_6t
Xbit_r28_c242 bl[242] br[242] wl[28] vdd gnd cell_6t
Xbit_r29_c242 bl[242] br[242] wl[29] vdd gnd cell_6t
Xbit_r30_c242 bl[242] br[242] wl[30] vdd gnd cell_6t
Xbit_r31_c242 bl[242] br[242] wl[31] vdd gnd cell_6t
Xbit_r32_c242 bl[242] br[242] wl[32] vdd gnd cell_6t
Xbit_r33_c242 bl[242] br[242] wl[33] vdd gnd cell_6t
Xbit_r34_c242 bl[242] br[242] wl[34] vdd gnd cell_6t
Xbit_r35_c242 bl[242] br[242] wl[35] vdd gnd cell_6t
Xbit_r36_c242 bl[242] br[242] wl[36] vdd gnd cell_6t
Xbit_r37_c242 bl[242] br[242] wl[37] vdd gnd cell_6t
Xbit_r38_c242 bl[242] br[242] wl[38] vdd gnd cell_6t
Xbit_r39_c242 bl[242] br[242] wl[39] vdd gnd cell_6t
Xbit_r40_c242 bl[242] br[242] wl[40] vdd gnd cell_6t
Xbit_r41_c242 bl[242] br[242] wl[41] vdd gnd cell_6t
Xbit_r42_c242 bl[242] br[242] wl[42] vdd gnd cell_6t
Xbit_r43_c242 bl[242] br[242] wl[43] vdd gnd cell_6t
Xbit_r44_c242 bl[242] br[242] wl[44] vdd gnd cell_6t
Xbit_r45_c242 bl[242] br[242] wl[45] vdd gnd cell_6t
Xbit_r46_c242 bl[242] br[242] wl[46] vdd gnd cell_6t
Xbit_r47_c242 bl[242] br[242] wl[47] vdd gnd cell_6t
Xbit_r48_c242 bl[242] br[242] wl[48] vdd gnd cell_6t
Xbit_r49_c242 bl[242] br[242] wl[49] vdd gnd cell_6t
Xbit_r50_c242 bl[242] br[242] wl[50] vdd gnd cell_6t
Xbit_r51_c242 bl[242] br[242] wl[51] vdd gnd cell_6t
Xbit_r52_c242 bl[242] br[242] wl[52] vdd gnd cell_6t
Xbit_r53_c242 bl[242] br[242] wl[53] vdd gnd cell_6t
Xbit_r54_c242 bl[242] br[242] wl[54] vdd gnd cell_6t
Xbit_r55_c242 bl[242] br[242] wl[55] vdd gnd cell_6t
Xbit_r56_c242 bl[242] br[242] wl[56] vdd gnd cell_6t
Xbit_r57_c242 bl[242] br[242] wl[57] vdd gnd cell_6t
Xbit_r58_c242 bl[242] br[242] wl[58] vdd gnd cell_6t
Xbit_r59_c242 bl[242] br[242] wl[59] vdd gnd cell_6t
Xbit_r60_c242 bl[242] br[242] wl[60] vdd gnd cell_6t
Xbit_r61_c242 bl[242] br[242] wl[61] vdd gnd cell_6t
Xbit_r62_c242 bl[242] br[242] wl[62] vdd gnd cell_6t
Xbit_r63_c242 bl[242] br[242] wl[63] vdd gnd cell_6t
Xbit_r64_c242 bl[242] br[242] wl[64] vdd gnd cell_6t
Xbit_r65_c242 bl[242] br[242] wl[65] vdd gnd cell_6t
Xbit_r66_c242 bl[242] br[242] wl[66] vdd gnd cell_6t
Xbit_r67_c242 bl[242] br[242] wl[67] vdd gnd cell_6t
Xbit_r68_c242 bl[242] br[242] wl[68] vdd gnd cell_6t
Xbit_r69_c242 bl[242] br[242] wl[69] vdd gnd cell_6t
Xbit_r70_c242 bl[242] br[242] wl[70] vdd gnd cell_6t
Xbit_r71_c242 bl[242] br[242] wl[71] vdd gnd cell_6t
Xbit_r72_c242 bl[242] br[242] wl[72] vdd gnd cell_6t
Xbit_r73_c242 bl[242] br[242] wl[73] vdd gnd cell_6t
Xbit_r74_c242 bl[242] br[242] wl[74] vdd gnd cell_6t
Xbit_r75_c242 bl[242] br[242] wl[75] vdd gnd cell_6t
Xbit_r76_c242 bl[242] br[242] wl[76] vdd gnd cell_6t
Xbit_r77_c242 bl[242] br[242] wl[77] vdd gnd cell_6t
Xbit_r78_c242 bl[242] br[242] wl[78] vdd gnd cell_6t
Xbit_r79_c242 bl[242] br[242] wl[79] vdd gnd cell_6t
Xbit_r80_c242 bl[242] br[242] wl[80] vdd gnd cell_6t
Xbit_r81_c242 bl[242] br[242] wl[81] vdd gnd cell_6t
Xbit_r82_c242 bl[242] br[242] wl[82] vdd gnd cell_6t
Xbit_r83_c242 bl[242] br[242] wl[83] vdd gnd cell_6t
Xbit_r84_c242 bl[242] br[242] wl[84] vdd gnd cell_6t
Xbit_r85_c242 bl[242] br[242] wl[85] vdd gnd cell_6t
Xbit_r86_c242 bl[242] br[242] wl[86] vdd gnd cell_6t
Xbit_r87_c242 bl[242] br[242] wl[87] vdd gnd cell_6t
Xbit_r88_c242 bl[242] br[242] wl[88] vdd gnd cell_6t
Xbit_r89_c242 bl[242] br[242] wl[89] vdd gnd cell_6t
Xbit_r90_c242 bl[242] br[242] wl[90] vdd gnd cell_6t
Xbit_r91_c242 bl[242] br[242] wl[91] vdd gnd cell_6t
Xbit_r92_c242 bl[242] br[242] wl[92] vdd gnd cell_6t
Xbit_r93_c242 bl[242] br[242] wl[93] vdd gnd cell_6t
Xbit_r94_c242 bl[242] br[242] wl[94] vdd gnd cell_6t
Xbit_r95_c242 bl[242] br[242] wl[95] vdd gnd cell_6t
Xbit_r96_c242 bl[242] br[242] wl[96] vdd gnd cell_6t
Xbit_r97_c242 bl[242] br[242] wl[97] vdd gnd cell_6t
Xbit_r98_c242 bl[242] br[242] wl[98] vdd gnd cell_6t
Xbit_r99_c242 bl[242] br[242] wl[99] vdd gnd cell_6t
Xbit_r100_c242 bl[242] br[242] wl[100] vdd gnd cell_6t
Xbit_r101_c242 bl[242] br[242] wl[101] vdd gnd cell_6t
Xbit_r102_c242 bl[242] br[242] wl[102] vdd gnd cell_6t
Xbit_r103_c242 bl[242] br[242] wl[103] vdd gnd cell_6t
Xbit_r104_c242 bl[242] br[242] wl[104] vdd gnd cell_6t
Xbit_r105_c242 bl[242] br[242] wl[105] vdd gnd cell_6t
Xbit_r106_c242 bl[242] br[242] wl[106] vdd gnd cell_6t
Xbit_r107_c242 bl[242] br[242] wl[107] vdd gnd cell_6t
Xbit_r108_c242 bl[242] br[242] wl[108] vdd gnd cell_6t
Xbit_r109_c242 bl[242] br[242] wl[109] vdd gnd cell_6t
Xbit_r110_c242 bl[242] br[242] wl[110] vdd gnd cell_6t
Xbit_r111_c242 bl[242] br[242] wl[111] vdd gnd cell_6t
Xbit_r112_c242 bl[242] br[242] wl[112] vdd gnd cell_6t
Xbit_r113_c242 bl[242] br[242] wl[113] vdd gnd cell_6t
Xbit_r114_c242 bl[242] br[242] wl[114] vdd gnd cell_6t
Xbit_r115_c242 bl[242] br[242] wl[115] vdd gnd cell_6t
Xbit_r116_c242 bl[242] br[242] wl[116] vdd gnd cell_6t
Xbit_r117_c242 bl[242] br[242] wl[117] vdd gnd cell_6t
Xbit_r118_c242 bl[242] br[242] wl[118] vdd gnd cell_6t
Xbit_r119_c242 bl[242] br[242] wl[119] vdd gnd cell_6t
Xbit_r120_c242 bl[242] br[242] wl[120] vdd gnd cell_6t
Xbit_r121_c242 bl[242] br[242] wl[121] vdd gnd cell_6t
Xbit_r122_c242 bl[242] br[242] wl[122] vdd gnd cell_6t
Xbit_r123_c242 bl[242] br[242] wl[123] vdd gnd cell_6t
Xbit_r124_c242 bl[242] br[242] wl[124] vdd gnd cell_6t
Xbit_r125_c242 bl[242] br[242] wl[125] vdd gnd cell_6t
Xbit_r126_c242 bl[242] br[242] wl[126] vdd gnd cell_6t
Xbit_r127_c242 bl[242] br[242] wl[127] vdd gnd cell_6t
Xbit_r0_c243 bl[243] br[243] wl[0] vdd gnd cell_6t
Xbit_r1_c243 bl[243] br[243] wl[1] vdd gnd cell_6t
Xbit_r2_c243 bl[243] br[243] wl[2] vdd gnd cell_6t
Xbit_r3_c243 bl[243] br[243] wl[3] vdd gnd cell_6t
Xbit_r4_c243 bl[243] br[243] wl[4] vdd gnd cell_6t
Xbit_r5_c243 bl[243] br[243] wl[5] vdd gnd cell_6t
Xbit_r6_c243 bl[243] br[243] wl[6] vdd gnd cell_6t
Xbit_r7_c243 bl[243] br[243] wl[7] vdd gnd cell_6t
Xbit_r8_c243 bl[243] br[243] wl[8] vdd gnd cell_6t
Xbit_r9_c243 bl[243] br[243] wl[9] vdd gnd cell_6t
Xbit_r10_c243 bl[243] br[243] wl[10] vdd gnd cell_6t
Xbit_r11_c243 bl[243] br[243] wl[11] vdd gnd cell_6t
Xbit_r12_c243 bl[243] br[243] wl[12] vdd gnd cell_6t
Xbit_r13_c243 bl[243] br[243] wl[13] vdd gnd cell_6t
Xbit_r14_c243 bl[243] br[243] wl[14] vdd gnd cell_6t
Xbit_r15_c243 bl[243] br[243] wl[15] vdd gnd cell_6t
Xbit_r16_c243 bl[243] br[243] wl[16] vdd gnd cell_6t
Xbit_r17_c243 bl[243] br[243] wl[17] vdd gnd cell_6t
Xbit_r18_c243 bl[243] br[243] wl[18] vdd gnd cell_6t
Xbit_r19_c243 bl[243] br[243] wl[19] vdd gnd cell_6t
Xbit_r20_c243 bl[243] br[243] wl[20] vdd gnd cell_6t
Xbit_r21_c243 bl[243] br[243] wl[21] vdd gnd cell_6t
Xbit_r22_c243 bl[243] br[243] wl[22] vdd gnd cell_6t
Xbit_r23_c243 bl[243] br[243] wl[23] vdd gnd cell_6t
Xbit_r24_c243 bl[243] br[243] wl[24] vdd gnd cell_6t
Xbit_r25_c243 bl[243] br[243] wl[25] vdd gnd cell_6t
Xbit_r26_c243 bl[243] br[243] wl[26] vdd gnd cell_6t
Xbit_r27_c243 bl[243] br[243] wl[27] vdd gnd cell_6t
Xbit_r28_c243 bl[243] br[243] wl[28] vdd gnd cell_6t
Xbit_r29_c243 bl[243] br[243] wl[29] vdd gnd cell_6t
Xbit_r30_c243 bl[243] br[243] wl[30] vdd gnd cell_6t
Xbit_r31_c243 bl[243] br[243] wl[31] vdd gnd cell_6t
Xbit_r32_c243 bl[243] br[243] wl[32] vdd gnd cell_6t
Xbit_r33_c243 bl[243] br[243] wl[33] vdd gnd cell_6t
Xbit_r34_c243 bl[243] br[243] wl[34] vdd gnd cell_6t
Xbit_r35_c243 bl[243] br[243] wl[35] vdd gnd cell_6t
Xbit_r36_c243 bl[243] br[243] wl[36] vdd gnd cell_6t
Xbit_r37_c243 bl[243] br[243] wl[37] vdd gnd cell_6t
Xbit_r38_c243 bl[243] br[243] wl[38] vdd gnd cell_6t
Xbit_r39_c243 bl[243] br[243] wl[39] vdd gnd cell_6t
Xbit_r40_c243 bl[243] br[243] wl[40] vdd gnd cell_6t
Xbit_r41_c243 bl[243] br[243] wl[41] vdd gnd cell_6t
Xbit_r42_c243 bl[243] br[243] wl[42] vdd gnd cell_6t
Xbit_r43_c243 bl[243] br[243] wl[43] vdd gnd cell_6t
Xbit_r44_c243 bl[243] br[243] wl[44] vdd gnd cell_6t
Xbit_r45_c243 bl[243] br[243] wl[45] vdd gnd cell_6t
Xbit_r46_c243 bl[243] br[243] wl[46] vdd gnd cell_6t
Xbit_r47_c243 bl[243] br[243] wl[47] vdd gnd cell_6t
Xbit_r48_c243 bl[243] br[243] wl[48] vdd gnd cell_6t
Xbit_r49_c243 bl[243] br[243] wl[49] vdd gnd cell_6t
Xbit_r50_c243 bl[243] br[243] wl[50] vdd gnd cell_6t
Xbit_r51_c243 bl[243] br[243] wl[51] vdd gnd cell_6t
Xbit_r52_c243 bl[243] br[243] wl[52] vdd gnd cell_6t
Xbit_r53_c243 bl[243] br[243] wl[53] vdd gnd cell_6t
Xbit_r54_c243 bl[243] br[243] wl[54] vdd gnd cell_6t
Xbit_r55_c243 bl[243] br[243] wl[55] vdd gnd cell_6t
Xbit_r56_c243 bl[243] br[243] wl[56] vdd gnd cell_6t
Xbit_r57_c243 bl[243] br[243] wl[57] vdd gnd cell_6t
Xbit_r58_c243 bl[243] br[243] wl[58] vdd gnd cell_6t
Xbit_r59_c243 bl[243] br[243] wl[59] vdd gnd cell_6t
Xbit_r60_c243 bl[243] br[243] wl[60] vdd gnd cell_6t
Xbit_r61_c243 bl[243] br[243] wl[61] vdd gnd cell_6t
Xbit_r62_c243 bl[243] br[243] wl[62] vdd gnd cell_6t
Xbit_r63_c243 bl[243] br[243] wl[63] vdd gnd cell_6t
Xbit_r64_c243 bl[243] br[243] wl[64] vdd gnd cell_6t
Xbit_r65_c243 bl[243] br[243] wl[65] vdd gnd cell_6t
Xbit_r66_c243 bl[243] br[243] wl[66] vdd gnd cell_6t
Xbit_r67_c243 bl[243] br[243] wl[67] vdd gnd cell_6t
Xbit_r68_c243 bl[243] br[243] wl[68] vdd gnd cell_6t
Xbit_r69_c243 bl[243] br[243] wl[69] vdd gnd cell_6t
Xbit_r70_c243 bl[243] br[243] wl[70] vdd gnd cell_6t
Xbit_r71_c243 bl[243] br[243] wl[71] vdd gnd cell_6t
Xbit_r72_c243 bl[243] br[243] wl[72] vdd gnd cell_6t
Xbit_r73_c243 bl[243] br[243] wl[73] vdd gnd cell_6t
Xbit_r74_c243 bl[243] br[243] wl[74] vdd gnd cell_6t
Xbit_r75_c243 bl[243] br[243] wl[75] vdd gnd cell_6t
Xbit_r76_c243 bl[243] br[243] wl[76] vdd gnd cell_6t
Xbit_r77_c243 bl[243] br[243] wl[77] vdd gnd cell_6t
Xbit_r78_c243 bl[243] br[243] wl[78] vdd gnd cell_6t
Xbit_r79_c243 bl[243] br[243] wl[79] vdd gnd cell_6t
Xbit_r80_c243 bl[243] br[243] wl[80] vdd gnd cell_6t
Xbit_r81_c243 bl[243] br[243] wl[81] vdd gnd cell_6t
Xbit_r82_c243 bl[243] br[243] wl[82] vdd gnd cell_6t
Xbit_r83_c243 bl[243] br[243] wl[83] vdd gnd cell_6t
Xbit_r84_c243 bl[243] br[243] wl[84] vdd gnd cell_6t
Xbit_r85_c243 bl[243] br[243] wl[85] vdd gnd cell_6t
Xbit_r86_c243 bl[243] br[243] wl[86] vdd gnd cell_6t
Xbit_r87_c243 bl[243] br[243] wl[87] vdd gnd cell_6t
Xbit_r88_c243 bl[243] br[243] wl[88] vdd gnd cell_6t
Xbit_r89_c243 bl[243] br[243] wl[89] vdd gnd cell_6t
Xbit_r90_c243 bl[243] br[243] wl[90] vdd gnd cell_6t
Xbit_r91_c243 bl[243] br[243] wl[91] vdd gnd cell_6t
Xbit_r92_c243 bl[243] br[243] wl[92] vdd gnd cell_6t
Xbit_r93_c243 bl[243] br[243] wl[93] vdd gnd cell_6t
Xbit_r94_c243 bl[243] br[243] wl[94] vdd gnd cell_6t
Xbit_r95_c243 bl[243] br[243] wl[95] vdd gnd cell_6t
Xbit_r96_c243 bl[243] br[243] wl[96] vdd gnd cell_6t
Xbit_r97_c243 bl[243] br[243] wl[97] vdd gnd cell_6t
Xbit_r98_c243 bl[243] br[243] wl[98] vdd gnd cell_6t
Xbit_r99_c243 bl[243] br[243] wl[99] vdd gnd cell_6t
Xbit_r100_c243 bl[243] br[243] wl[100] vdd gnd cell_6t
Xbit_r101_c243 bl[243] br[243] wl[101] vdd gnd cell_6t
Xbit_r102_c243 bl[243] br[243] wl[102] vdd gnd cell_6t
Xbit_r103_c243 bl[243] br[243] wl[103] vdd gnd cell_6t
Xbit_r104_c243 bl[243] br[243] wl[104] vdd gnd cell_6t
Xbit_r105_c243 bl[243] br[243] wl[105] vdd gnd cell_6t
Xbit_r106_c243 bl[243] br[243] wl[106] vdd gnd cell_6t
Xbit_r107_c243 bl[243] br[243] wl[107] vdd gnd cell_6t
Xbit_r108_c243 bl[243] br[243] wl[108] vdd gnd cell_6t
Xbit_r109_c243 bl[243] br[243] wl[109] vdd gnd cell_6t
Xbit_r110_c243 bl[243] br[243] wl[110] vdd gnd cell_6t
Xbit_r111_c243 bl[243] br[243] wl[111] vdd gnd cell_6t
Xbit_r112_c243 bl[243] br[243] wl[112] vdd gnd cell_6t
Xbit_r113_c243 bl[243] br[243] wl[113] vdd gnd cell_6t
Xbit_r114_c243 bl[243] br[243] wl[114] vdd gnd cell_6t
Xbit_r115_c243 bl[243] br[243] wl[115] vdd gnd cell_6t
Xbit_r116_c243 bl[243] br[243] wl[116] vdd gnd cell_6t
Xbit_r117_c243 bl[243] br[243] wl[117] vdd gnd cell_6t
Xbit_r118_c243 bl[243] br[243] wl[118] vdd gnd cell_6t
Xbit_r119_c243 bl[243] br[243] wl[119] vdd gnd cell_6t
Xbit_r120_c243 bl[243] br[243] wl[120] vdd gnd cell_6t
Xbit_r121_c243 bl[243] br[243] wl[121] vdd gnd cell_6t
Xbit_r122_c243 bl[243] br[243] wl[122] vdd gnd cell_6t
Xbit_r123_c243 bl[243] br[243] wl[123] vdd gnd cell_6t
Xbit_r124_c243 bl[243] br[243] wl[124] vdd gnd cell_6t
Xbit_r125_c243 bl[243] br[243] wl[125] vdd gnd cell_6t
Xbit_r126_c243 bl[243] br[243] wl[126] vdd gnd cell_6t
Xbit_r127_c243 bl[243] br[243] wl[127] vdd gnd cell_6t
Xbit_r0_c244 bl[244] br[244] wl[0] vdd gnd cell_6t
Xbit_r1_c244 bl[244] br[244] wl[1] vdd gnd cell_6t
Xbit_r2_c244 bl[244] br[244] wl[2] vdd gnd cell_6t
Xbit_r3_c244 bl[244] br[244] wl[3] vdd gnd cell_6t
Xbit_r4_c244 bl[244] br[244] wl[4] vdd gnd cell_6t
Xbit_r5_c244 bl[244] br[244] wl[5] vdd gnd cell_6t
Xbit_r6_c244 bl[244] br[244] wl[6] vdd gnd cell_6t
Xbit_r7_c244 bl[244] br[244] wl[7] vdd gnd cell_6t
Xbit_r8_c244 bl[244] br[244] wl[8] vdd gnd cell_6t
Xbit_r9_c244 bl[244] br[244] wl[9] vdd gnd cell_6t
Xbit_r10_c244 bl[244] br[244] wl[10] vdd gnd cell_6t
Xbit_r11_c244 bl[244] br[244] wl[11] vdd gnd cell_6t
Xbit_r12_c244 bl[244] br[244] wl[12] vdd gnd cell_6t
Xbit_r13_c244 bl[244] br[244] wl[13] vdd gnd cell_6t
Xbit_r14_c244 bl[244] br[244] wl[14] vdd gnd cell_6t
Xbit_r15_c244 bl[244] br[244] wl[15] vdd gnd cell_6t
Xbit_r16_c244 bl[244] br[244] wl[16] vdd gnd cell_6t
Xbit_r17_c244 bl[244] br[244] wl[17] vdd gnd cell_6t
Xbit_r18_c244 bl[244] br[244] wl[18] vdd gnd cell_6t
Xbit_r19_c244 bl[244] br[244] wl[19] vdd gnd cell_6t
Xbit_r20_c244 bl[244] br[244] wl[20] vdd gnd cell_6t
Xbit_r21_c244 bl[244] br[244] wl[21] vdd gnd cell_6t
Xbit_r22_c244 bl[244] br[244] wl[22] vdd gnd cell_6t
Xbit_r23_c244 bl[244] br[244] wl[23] vdd gnd cell_6t
Xbit_r24_c244 bl[244] br[244] wl[24] vdd gnd cell_6t
Xbit_r25_c244 bl[244] br[244] wl[25] vdd gnd cell_6t
Xbit_r26_c244 bl[244] br[244] wl[26] vdd gnd cell_6t
Xbit_r27_c244 bl[244] br[244] wl[27] vdd gnd cell_6t
Xbit_r28_c244 bl[244] br[244] wl[28] vdd gnd cell_6t
Xbit_r29_c244 bl[244] br[244] wl[29] vdd gnd cell_6t
Xbit_r30_c244 bl[244] br[244] wl[30] vdd gnd cell_6t
Xbit_r31_c244 bl[244] br[244] wl[31] vdd gnd cell_6t
Xbit_r32_c244 bl[244] br[244] wl[32] vdd gnd cell_6t
Xbit_r33_c244 bl[244] br[244] wl[33] vdd gnd cell_6t
Xbit_r34_c244 bl[244] br[244] wl[34] vdd gnd cell_6t
Xbit_r35_c244 bl[244] br[244] wl[35] vdd gnd cell_6t
Xbit_r36_c244 bl[244] br[244] wl[36] vdd gnd cell_6t
Xbit_r37_c244 bl[244] br[244] wl[37] vdd gnd cell_6t
Xbit_r38_c244 bl[244] br[244] wl[38] vdd gnd cell_6t
Xbit_r39_c244 bl[244] br[244] wl[39] vdd gnd cell_6t
Xbit_r40_c244 bl[244] br[244] wl[40] vdd gnd cell_6t
Xbit_r41_c244 bl[244] br[244] wl[41] vdd gnd cell_6t
Xbit_r42_c244 bl[244] br[244] wl[42] vdd gnd cell_6t
Xbit_r43_c244 bl[244] br[244] wl[43] vdd gnd cell_6t
Xbit_r44_c244 bl[244] br[244] wl[44] vdd gnd cell_6t
Xbit_r45_c244 bl[244] br[244] wl[45] vdd gnd cell_6t
Xbit_r46_c244 bl[244] br[244] wl[46] vdd gnd cell_6t
Xbit_r47_c244 bl[244] br[244] wl[47] vdd gnd cell_6t
Xbit_r48_c244 bl[244] br[244] wl[48] vdd gnd cell_6t
Xbit_r49_c244 bl[244] br[244] wl[49] vdd gnd cell_6t
Xbit_r50_c244 bl[244] br[244] wl[50] vdd gnd cell_6t
Xbit_r51_c244 bl[244] br[244] wl[51] vdd gnd cell_6t
Xbit_r52_c244 bl[244] br[244] wl[52] vdd gnd cell_6t
Xbit_r53_c244 bl[244] br[244] wl[53] vdd gnd cell_6t
Xbit_r54_c244 bl[244] br[244] wl[54] vdd gnd cell_6t
Xbit_r55_c244 bl[244] br[244] wl[55] vdd gnd cell_6t
Xbit_r56_c244 bl[244] br[244] wl[56] vdd gnd cell_6t
Xbit_r57_c244 bl[244] br[244] wl[57] vdd gnd cell_6t
Xbit_r58_c244 bl[244] br[244] wl[58] vdd gnd cell_6t
Xbit_r59_c244 bl[244] br[244] wl[59] vdd gnd cell_6t
Xbit_r60_c244 bl[244] br[244] wl[60] vdd gnd cell_6t
Xbit_r61_c244 bl[244] br[244] wl[61] vdd gnd cell_6t
Xbit_r62_c244 bl[244] br[244] wl[62] vdd gnd cell_6t
Xbit_r63_c244 bl[244] br[244] wl[63] vdd gnd cell_6t
Xbit_r64_c244 bl[244] br[244] wl[64] vdd gnd cell_6t
Xbit_r65_c244 bl[244] br[244] wl[65] vdd gnd cell_6t
Xbit_r66_c244 bl[244] br[244] wl[66] vdd gnd cell_6t
Xbit_r67_c244 bl[244] br[244] wl[67] vdd gnd cell_6t
Xbit_r68_c244 bl[244] br[244] wl[68] vdd gnd cell_6t
Xbit_r69_c244 bl[244] br[244] wl[69] vdd gnd cell_6t
Xbit_r70_c244 bl[244] br[244] wl[70] vdd gnd cell_6t
Xbit_r71_c244 bl[244] br[244] wl[71] vdd gnd cell_6t
Xbit_r72_c244 bl[244] br[244] wl[72] vdd gnd cell_6t
Xbit_r73_c244 bl[244] br[244] wl[73] vdd gnd cell_6t
Xbit_r74_c244 bl[244] br[244] wl[74] vdd gnd cell_6t
Xbit_r75_c244 bl[244] br[244] wl[75] vdd gnd cell_6t
Xbit_r76_c244 bl[244] br[244] wl[76] vdd gnd cell_6t
Xbit_r77_c244 bl[244] br[244] wl[77] vdd gnd cell_6t
Xbit_r78_c244 bl[244] br[244] wl[78] vdd gnd cell_6t
Xbit_r79_c244 bl[244] br[244] wl[79] vdd gnd cell_6t
Xbit_r80_c244 bl[244] br[244] wl[80] vdd gnd cell_6t
Xbit_r81_c244 bl[244] br[244] wl[81] vdd gnd cell_6t
Xbit_r82_c244 bl[244] br[244] wl[82] vdd gnd cell_6t
Xbit_r83_c244 bl[244] br[244] wl[83] vdd gnd cell_6t
Xbit_r84_c244 bl[244] br[244] wl[84] vdd gnd cell_6t
Xbit_r85_c244 bl[244] br[244] wl[85] vdd gnd cell_6t
Xbit_r86_c244 bl[244] br[244] wl[86] vdd gnd cell_6t
Xbit_r87_c244 bl[244] br[244] wl[87] vdd gnd cell_6t
Xbit_r88_c244 bl[244] br[244] wl[88] vdd gnd cell_6t
Xbit_r89_c244 bl[244] br[244] wl[89] vdd gnd cell_6t
Xbit_r90_c244 bl[244] br[244] wl[90] vdd gnd cell_6t
Xbit_r91_c244 bl[244] br[244] wl[91] vdd gnd cell_6t
Xbit_r92_c244 bl[244] br[244] wl[92] vdd gnd cell_6t
Xbit_r93_c244 bl[244] br[244] wl[93] vdd gnd cell_6t
Xbit_r94_c244 bl[244] br[244] wl[94] vdd gnd cell_6t
Xbit_r95_c244 bl[244] br[244] wl[95] vdd gnd cell_6t
Xbit_r96_c244 bl[244] br[244] wl[96] vdd gnd cell_6t
Xbit_r97_c244 bl[244] br[244] wl[97] vdd gnd cell_6t
Xbit_r98_c244 bl[244] br[244] wl[98] vdd gnd cell_6t
Xbit_r99_c244 bl[244] br[244] wl[99] vdd gnd cell_6t
Xbit_r100_c244 bl[244] br[244] wl[100] vdd gnd cell_6t
Xbit_r101_c244 bl[244] br[244] wl[101] vdd gnd cell_6t
Xbit_r102_c244 bl[244] br[244] wl[102] vdd gnd cell_6t
Xbit_r103_c244 bl[244] br[244] wl[103] vdd gnd cell_6t
Xbit_r104_c244 bl[244] br[244] wl[104] vdd gnd cell_6t
Xbit_r105_c244 bl[244] br[244] wl[105] vdd gnd cell_6t
Xbit_r106_c244 bl[244] br[244] wl[106] vdd gnd cell_6t
Xbit_r107_c244 bl[244] br[244] wl[107] vdd gnd cell_6t
Xbit_r108_c244 bl[244] br[244] wl[108] vdd gnd cell_6t
Xbit_r109_c244 bl[244] br[244] wl[109] vdd gnd cell_6t
Xbit_r110_c244 bl[244] br[244] wl[110] vdd gnd cell_6t
Xbit_r111_c244 bl[244] br[244] wl[111] vdd gnd cell_6t
Xbit_r112_c244 bl[244] br[244] wl[112] vdd gnd cell_6t
Xbit_r113_c244 bl[244] br[244] wl[113] vdd gnd cell_6t
Xbit_r114_c244 bl[244] br[244] wl[114] vdd gnd cell_6t
Xbit_r115_c244 bl[244] br[244] wl[115] vdd gnd cell_6t
Xbit_r116_c244 bl[244] br[244] wl[116] vdd gnd cell_6t
Xbit_r117_c244 bl[244] br[244] wl[117] vdd gnd cell_6t
Xbit_r118_c244 bl[244] br[244] wl[118] vdd gnd cell_6t
Xbit_r119_c244 bl[244] br[244] wl[119] vdd gnd cell_6t
Xbit_r120_c244 bl[244] br[244] wl[120] vdd gnd cell_6t
Xbit_r121_c244 bl[244] br[244] wl[121] vdd gnd cell_6t
Xbit_r122_c244 bl[244] br[244] wl[122] vdd gnd cell_6t
Xbit_r123_c244 bl[244] br[244] wl[123] vdd gnd cell_6t
Xbit_r124_c244 bl[244] br[244] wl[124] vdd gnd cell_6t
Xbit_r125_c244 bl[244] br[244] wl[125] vdd gnd cell_6t
Xbit_r126_c244 bl[244] br[244] wl[126] vdd gnd cell_6t
Xbit_r127_c244 bl[244] br[244] wl[127] vdd gnd cell_6t
Xbit_r0_c245 bl[245] br[245] wl[0] vdd gnd cell_6t
Xbit_r1_c245 bl[245] br[245] wl[1] vdd gnd cell_6t
Xbit_r2_c245 bl[245] br[245] wl[2] vdd gnd cell_6t
Xbit_r3_c245 bl[245] br[245] wl[3] vdd gnd cell_6t
Xbit_r4_c245 bl[245] br[245] wl[4] vdd gnd cell_6t
Xbit_r5_c245 bl[245] br[245] wl[5] vdd gnd cell_6t
Xbit_r6_c245 bl[245] br[245] wl[6] vdd gnd cell_6t
Xbit_r7_c245 bl[245] br[245] wl[7] vdd gnd cell_6t
Xbit_r8_c245 bl[245] br[245] wl[8] vdd gnd cell_6t
Xbit_r9_c245 bl[245] br[245] wl[9] vdd gnd cell_6t
Xbit_r10_c245 bl[245] br[245] wl[10] vdd gnd cell_6t
Xbit_r11_c245 bl[245] br[245] wl[11] vdd gnd cell_6t
Xbit_r12_c245 bl[245] br[245] wl[12] vdd gnd cell_6t
Xbit_r13_c245 bl[245] br[245] wl[13] vdd gnd cell_6t
Xbit_r14_c245 bl[245] br[245] wl[14] vdd gnd cell_6t
Xbit_r15_c245 bl[245] br[245] wl[15] vdd gnd cell_6t
Xbit_r16_c245 bl[245] br[245] wl[16] vdd gnd cell_6t
Xbit_r17_c245 bl[245] br[245] wl[17] vdd gnd cell_6t
Xbit_r18_c245 bl[245] br[245] wl[18] vdd gnd cell_6t
Xbit_r19_c245 bl[245] br[245] wl[19] vdd gnd cell_6t
Xbit_r20_c245 bl[245] br[245] wl[20] vdd gnd cell_6t
Xbit_r21_c245 bl[245] br[245] wl[21] vdd gnd cell_6t
Xbit_r22_c245 bl[245] br[245] wl[22] vdd gnd cell_6t
Xbit_r23_c245 bl[245] br[245] wl[23] vdd gnd cell_6t
Xbit_r24_c245 bl[245] br[245] wl[24] vdd gnd cell_6t
Xbit_r25_c245 bl[245] br[245] wl[25] vdd gnd cell_6t
Xbit_r26_c245 bl[245] br[245] wl[26] vdd gnd cell_6t
Xbit_r27_c245 bl[245] br[245] wl[27] vdd gnd cell_6t
Xbit_r28_c245 bl[245] br[245] wl[28] vdd gnd cell_6t
Xbit_r29_c245 bl[245] br[245] wl[29] vdd gnd cell_6t
Xbit_r30_c245 bl[245] br[245] wl[30] vdd gnd cell_6t
Xbit_r31_c245 bl[245] br[245] wl[31] vdd gnd cell_6t
Xbit_r32_c245 bl[245] br[245] wl[32] vdd gnd cell_6t
Xbit_r33_c245 bl[245] br[245] wl[33] vdd gnd cell_6t
Xbit_r34_c245 bl[245] br[245] wl[34] vdd gnd cell_6t
Xbit_r35_c245 bl[245] br[245] wl[35] vdd gnd cell_6t
Xbit_r36_c245 bl[245] br[245] wl[36] vdd gnd cell_6t
Xbit_r37_c245 bl[245] br[245] wl[37] vdd gnd cell_6t
Xbit_r38_c245 bl[245] br[245] wl[38] vdd gnd cell_6t
Xbit_r39_c245 bl[245] br[245] wl[39] vdd gnd cell_6t
Xbit_r40_c245 bl[245] br[245] wl[40] vdd gnd cell_6t
Xbit_r41_c245 bl[245] br[245] wl[41] vdd gnd cell_6t
Xbit_r42_c245 bl[245] br[245] wl[42] vdd gnd cell_6t
Xbit_r43_c245 bl[245] br[245] wl[43] vdd gnd cell_6t
Xbit_r44_c245 bl[245] br[245] wl[44] vdd gnd cell_6t
Xbit_r45_c245 bl[245] br[245] wl[45] vdd gnd cell_6t
Xbit_r46_c245 bl[245] br[245] wl[46] vdd gnd cell_6t
Xbit_r47_c245 bl[245] br[245] wl[47] vdd gnd cell_6t
Xbit_r48_c245 bl[245] br[245] wl[48] vdd gnd cell_6t
Xbit_r49_c245 bl[245] br[245] wl[49] vdd gnd cell_6t
Xbit_r50_c245 bl[245] br[245] wl[50] vdd gnd cell_6t
Xbit_r51_c245 bl[245] br[245] wl[51] vdd gnd cell_6t
Xbit_r52_c245 bl[245] br[245] wl[52] vdd gnd cell_6t
Xbit_r53_c245 bl[245] br[245] wl[53] vdd gnd cell_6t
Xbit_r54_c245 bl[245] br[245] wl[54] vdd gnd cell_6t
Xbit_r55_c245 bl[245] br[245] wl[55] vdd gnd cell_6t
Xbit_r56_c245 bl[245] br[245] wl[56] vdd gnd cell_6t
Xbit_r57_c245 bl[245] br[245] wl[57] vdd gnd cell_6t
Xbit_r58_c245 bl[245] br[245] wl[58] vdd gnd cell_6t
Xbit_r59_c245 bl[245] br[245] wl[59] vdd gnd cell_6t
Xbit_r60_c245 bl[245] br[245] wl[60] vdd gnd cell_6t
Xbit_r61_c245 bl[245] br[245] wl[61] vdd gnd cell_6t
Xbit_r62_c245 bl[245] br[245] wl[62] vdd gnd cell_6t
Xbit_r63_c245 bl[245] br[245] wl[63] vdd gnd cell_6t
Xbit_r64_c245 bl[245] br[245] wl[64] vdd gnd cell_6t
Xbit_r65_c245 bl[245] br[245] wl[65] vdd gnd cell_6t
Xbit_r66_c245 bl[245] br[245] wl[66] vdd gnd cell_6t
Xbit_r67_c245 bl[245] br[245] wl[67] vdd gnd cell_6t
Xbit_r68_c245 bl[245] br[245] wl[68] vdd gnd cell_6t
Xbit_r69_c245 bl[245] br[245] wl[69] vdd gnd cell_6t
Xbit_r70_c245 bl[245] br[245] wl[70] vdd gnd cell_6t
Xbit_r71_c245 bl[245] br[245] wl[71] vdd gnd cell_6t
Xbit_r72_c245 bl[245] br[245] wl[72] vdd gnd cell_6t
Xbit_r73_c245 bl[245] br[245] wl[73] vdd gnd cell_6t
Xbit_r74_c245 bl[245] br[245] wl[74] vdd gnd cell_6t
Xbit_r75_c245 bl[245] br[245] wl[75] vdd gnd cell_6t
Xbit_r76_c245 bl[245] br[245] wl[76] vdd gnd cell_6t
Xbit_r77_c245 bl[245] br[245] wl[77] vdd gnd cell_6t
Xbit_r78_c245 bl[245] br[245] wl[78] vdd gnd cell_6t
Xbit_r79_c245 bl[245] br[245] wl[79] vdd gnd cell_6t
Xbit_r80_c245 bl[245] br[245] wl[80] vdd gnd cell_6t
Xbit_r81_c245 bl[245] br[245] wl[81] vdd gnd cell_6t
Xbit_r82_c245 bl[245] br[245] wl[82] vdd gnd cell_6t
Xbit_r83_c245 bl[245] br[245] wl[83] vdd gnd cell_6t
Xbit_r84_c245 bl[245] br[245] wl[84] vdd gnd cell_6t
Xbit_r85_c245 bl[245] br[245] wl[85] vdd gnd cell_6t
Xbit_r86_c245 bl[245] br[245] wl[86] vdd gnd cell_6t
Xbit_r87_c245 bl[245] br[245] wl[87] vdd gnd cell_6t
Xbit_r88_c245 bl[245] br[245] wl[88] vdd gnd cell_6t
Xbit_r89_c245 bl[245] br[245] wl[89] vdd gnd cell_6t
Xbit_r90_c245 bl[245] br[245] wl[90] vdd gnd cell_6t
Xbit_r91_c245 bl[245] br[245] wl[91] vdd gnd cell_6t
Xbit_r92_c245 bl[245] br[245] wl[92] vdd gnd cell_6t
Xbit_r93_c245 bl[245] br[245] wl[93] vdd gnd cell_6t
Xbit_r94_c245 bl[245] br[245] wl[94] vdd gnd cell_6t
Xbit_r95_c245 bl[245] br[245] wl[95] vdd gnd cell_6t
Xbit_r96_c245 bl[245] br[245] wl[96] vdd gnd cell_6t
Xbit_r97_c245 bl[245] br[245] wl[97] vdd gnd cell_6t
Xbit_r98_c245 bl[245] br[245] wl[98] vdd gnd cell_6t
Xbit_r99_c245 bl[245] br[245] wl[99] vdd gnd cell_6t
Xbit_r100_c245 bl[245] br[245] wl[100] vdd gnd cell_6t
Xbit_r101_c245 bl[245] br[245] wl[101] vdd gnd cell_6t
Xbit_r102_c245 bl[245] br[245] wl[102] vdd gnd cell_6t
Xbit_r103_c245 bl[245] br[245] wl[103] vdd gnd cell_6t
Xbit_r104_c245 bl[245] br[245] wl[104] vdd gnd cell_6t
Xbit_r105_c245 bl[245] br[245] wl[105] vdd gnd cell_6t
Xbit_r106_c245 bl[245] br[245] wl[106] vdd gnd cell_6t
Xbit_r107_c245 bl[245] br[245] wl[107] vdd gnd cell_6t
Xbit_r108_c245 bl[245] br[245] wl[108] vdd gnd cell_6t
Xbit_r109_c245 bl[245] br[245] wl[109] vdd gnd cell_6t
Xbit_r110_c245 bl[245] br[245] wl[110] vdd gnd cell_6t
Xbit_r111_c245 bl[245] br[245] wl[111] vdd gnd cell_6t
Xbit_r112_c245 bl[245] br[245] wl[112] vdd gnd cell_6t
Xbit_r113_c245 bl[245] br[245] wl[113] vdd gnd cell_6t
Xbit_r114_c245 bl[245] br[245] wl[114] vdd gnd cell_6t
Xbit_r115_c245 bl[245] br[245] wl[115] vdd gnd cell_6t
Xbit_r116_c245 bl[245] br[245] wl[116] vdd gnd cell_6t
Xbit_r117_c245 bl[245] br[245] wl[117] vdd gnd cell_6t
Xbit_r118_c245 bl[245] br[245] wl[118] vdd gnd cell_6t
Xbit_r119_c245 bl[245] br[245] wl[119] vdd gnd cell_6t
Xbit_r120_c245 bl[245] br[245] wl[120] vdd gnd cell_6t
Xbit_r121_c245 bl[245] br[245] wl[121] vdd gnd cell_6t
Xbit_r122_c245 bl[245] br[245] wl[122] vdd gnd cell_6t
Xbit_r123_c245 bl[245] br[245] wl[123] vdd gnd cell_6t
Xbit_r124_c245 bl[245] br[245] wl[124] vdd gnd cell_6t
Xbit_r125_c245 bl[245] br[245] wl[125] vdd gnd cell_6t
Xbit_r126_c245 bl[245] br[245] wl[126] vdd gnd cell_6t
Xbit_r127_c245 bl[245] br[245] wl[127] vdd gnd cell_6t
Xbit_r0_c246 bl[246] br[246] wl[0] vdd gnd cell_6t
Xbit_r1_c246 bl[246] br[246] wl[1] vdd gnd cell_6t
Xbit_r2_c246 bl[246] br[246] wl[2] vdd gnd cell_6t
Xbit_r3_c246 bl[246] br[246] wl[3] vdd gnd cell_6t
Xbit_r4_c246 bl[246] br[246] wl[4] vdd gnd cell_6t
Xbit_r5_c246 bl[246] br[246] wl[5] vdd gnd cell_6t
Xbit_r6_c246 bl[246] br[246] wl[6] vdd gnd cell_6t
Xbit_r7_c246 bl[246] br[246] wl[7] vdd gnd cell_6t
Xbit_r8_c246 bl[246] br[246] wl[8] vdd gnd cell_6t
Xbit_r9_c246 bl[246] br[246] wl[9] vdd gnd cell_6t
Xbit_r10_c246 bl[246] br[246] wl[10] vdd gnd cell_6t
Xbit_r11_c246 bl[246] br[246] wl[11] vdd gnd cell_6t
Xbit_r12_c246 bl[246] br[246] wl[12] vdd gnd cell_6t
Xbit_r13_c246 bl[246] br[246] wl[13] vdd gnd cell_6t
Xbit_r14_c246 bl[246] br[246] wl[14] vdd gnd cell_6t
Xbit_r15_c246 bl[246] br[246] wl[15] vdd gnd cell_6t
Xbit_r16_c246 bl[246] br[246] wl[16] vdd gnd cell_6t
Xbit_r17_c246 bl[246] br[246] wl[17] vdd gnd cell_6t
Xbit_r18_c246 bl[246] br[246] wl[18] vdd gnd cell_6t
Xbit_r19_c246 bl[246] br[246] wl[19] vdd gnd cell_6t
Xbit_r20_c246 bl[246] br[246] wl[20] vdd gnd cell_6t
Xbit_r21_c246 bl[246] br[246] wl[21] vdd gnd cell_6t
Xbit_r22_c246 bl[246] br[246] wl[22] vdd gnd cell_6t
Xbit_r23_c246 bl[246] br[246] wl[23] vdd gnd cell_6t
Xbit_r24_c246 bl[246] br[246] wl[24] vdd gnd cell_6t
Xbit_r25_c246 bl[246] br[246] wl[25] vdd gnd cell_6t
Xbit_r26_c246 bl[246] br[246] wl[26] vdd gnd cell_6t
Xbit_r27_c246 bl[246] br[246] wl[27] vdd gnd cell_6t
Xbit_r28_c246 bl[246] br[246] wl[28] vdd gnd cell_6t
Xbit_r29_c246 bl[246] br[246] wl[29] vdd gnd cell_6t
Xbit_r30_c246 bl[246] br[246] wl[30] vdd gnd cell_6t
Xbit_r31_c246 bl[246] br[246] wl[31] vdd gnd cell_6t
Xbit_r32_c246 bl[246] br[246] wl[32] vdd gnd cell_6t
Xbit_r33_c246 bl[246] br[246] wl[33] vdd gnd cell_6t
Xbit_r34_c246 bl[246] br[246] wl[34] vdd gnd cell_6t
Xbit_r35_c246 bl[246] br[246] wl[35] vdd gnd cell_6t
Xbit_r36_c246 bl[246] br[246] wl[36] vdd gnd cell_6t
Xbit_r37_c246 bl[246] br[246] wl[37] vdd gnd cell_6t
Xbit_r38_c246 bl[246] br[246] wl[38] vdd gnd cell_6t
Xbit_r39_c246 bl[246] br[246] wl[39] vdd gnd cell_6t
Xbit_r40_c246 bl[246] br[246] wl[40] vdd gnd cell_6t
Xbit_r41_c246 bl[246] br[246] wl[41] vdd gnd cell_6t
Xbit_r42_c246 bl[246] br[246] wl[42] vdd gnd cell_6t
Xbit_r43_c246 bl[246] br[246] wl[43] vdd gnd cell_6t
Xbit_r44_c246 bl[246] br[246] wl[44] vdd gnd cell_6t
Xbit_r45_c246 bl[246] br[246] wl[45] vdd gnd cell_6t
Xbit_r46_c246 bl[246] br[246] wl[46] vdd gnd cell_6t
Xbit_r47_c246 bl[246] br[246] wl[47] vdd gnd cell_6t
Xbit_r48_c246 bl[246] br[246] wl[48] vdd gnd cell_6t
Xbit_r49_c246 bl[246] br[246] wl[49] vdd gnd cell_6t
Xbit_r50_c246 bl[246] br[246] wl[50] vdd gnd cell_6t
Xbit_r51_c246 bl[246] br[246] wl[51] vdd gnd cell_6t
Xbit_r52_c246 bl[246] br[246] wl[52] vdd gnd cell_6t
Xbit_r53_c246 bl[246] br[246] wl[53] vdd gnd cell_6t
Xbit_r54_c246 bl[246] br[246] wl[54] vdd gnd cell_6t
Xbit_r55_c246 bl[246] br[246] wl[55] vdd gnd cell_6t
Xbit_r56_c246 bl[246] br[246] wl[56] vdd gnd cell_6t
Xbit_r57_c246 bl[246] br[246] wl[57] vdd gnd cell_6t
Xbit_r58_c246 bl[246] br[246] wl[58] vdd gnd cell_6t
Xbit_r59_c246 bl[246] br[246] wl[59] vdd gnd cell_6t
Xbit_r60_c246 bl[246] br[246] wl[60] vdd gnd cell_6t
Xbit_r61_c246 bl[246] br[246] wl[61] vdd gnd cell_6t
Xbit_r62_c246 bl[246] br[246] wl[62] vdd gnd cell_6t
Xbit_r63_c246 bl[246] br[246] wl[63] vdd gnd cell_6t
Xbit_r64_c246 bl[246] br[246] wl[64] vdd gnd cell_6t
Xbit_r65_c246 bl[246] br[246] wl[65] vdd gnd cell_6t
Xbit_r66_c246 bl[246] br[246] wl[66] vdd gnd cell_6t
Xbit_r67_c246 bl[246] br[246] wl[67] vdd gnd cell_6t
Xbit_r68_c246 bl[246] br[246] wl[68] vdd gnd cell_6t
Xbit_r69_c246 bl[246] br[246] wl[69] vdd gnd cell_6t
Xbit_r70_c246 bl[246] br[246] wl[70] vdd gnd cell_6t
Xbit_r71_c246 bl[246] br[246] wl[71] vdd gnd cell_6t
Xbit_r72_c246 bl[246] br[246] wl[72] vdd gnd cell_6t
Xbit_r73_c246 bl[246] br[246] wl[73] vdd gnd cell_6t
Xbit_r74_c246 bl[246] br[246] wl[74] vdd gnd cell_6t
Xbit_r75_c246 bl[246] br[246] wl[75] vdd gnd cell_6t
Xbit_r76_c246 bl[246] br[246] wl[76] vdd gnd cell_6t
Xbit_r77_c246 bl[246] br[246] wl[77] vdd gnd cell_6t
Xbit_r78_c246 bl[246] br[246] wl[78] vdd gnd cell_6t
Xbit_r79_c246 bl[246] br[246] wl[79] vdd gnd cell_6t
Xbit_r80_c246 bl[246] br[246] wl[80] vdd gnd cell_6t
Xbit_r81_c246 bl[246] br[246] wl[81] vdd gnd cell_6t
Xbit_r82_c246 bl[246] br[246] wl[82] vdd gnd cell_6t
Xbit_r83_c246 bl[246] br[246] wl[83] vdd gnd cell_6t
Xbit_r84_c246 bl[246] br[246] wl[84] vdd gnd cell_6t
Xbit_r85_c246 bl[246] br[246] wl[85] vdd gnd cell_6t
Xbit_r86_c246 bl[246] br[246] wl[86] vdd gnd cell_6t
Xbit_r87_c246 bl[246] br[246] wl[87] vdd gnd cell_6t
Xbit_r88_c246 bl[246] br[246] wl[88] vdd gnd cell_6t
Xbit_r89_c246 bl[246] br[246] wl[89] vdd gnd cell_6t
Xbit_r90_c246 bl[246] br[246] wl[90] vdd gnd cell_6t
Xbit_r91_c246 bl[246] br[246] wl[91] vdd gnd cell_6t
Xbit_r92_c246 bl[246] br[246] wl[92] vdd gnd cell_6t
Xbit_r93_c246 bl[246] br[246] wl[93] vdd gnd cell_6t
Xbit_r94_c246 bl[246] br[246] wl[94] vdd gnd cell_6t
Xbit_r95_c246 bl[246] br[246] wl[95] vdd gnd cell_6t
Xbit_r96_c246 bl[246] br[246] wl[96] vdd gnd cell_6t
Xbit_r97_c246 bl[246] br[246] wl[97] vdd gnd cell_6t
Xbit_r98_c246 bl[246] br[246] wl[98] vdd gnd cell_6t
Xbit_r99_c246 bl[246] br[246] wl[99] vdd gnd cell_6t
Xbit_r100_c246 bl[246] br[246] wl[100] vdd gnd cell_6t
Xbit_r101_c246 bl[246] br[246] wl[101] vdd gnd cell_6t
Xbit_r102_c246 bl[246] br[246] wl[102] vdd gnd cell_6t
Xbit_r103_c246 bl[246] br[246] wl[103] vdd gnd cell_6t
Xbit_r104_c246 bl[246] br[246] wl[104] vdd gnd cell_6t
Xbit_r105_c246 bl[246] br[246] wl[105] vdd gnd cell_6t
Xbit_r106_c246 bl[246] br[246] wl[106] vdd gnd cell_6t
Xbit_r107_c246 bl[246] br[246] wl[107] vdd gnd cell_6t
Xbit_r108_c246 bl[246] br[246] wl[108] vdd gnd cell_6t
Xbit_r109_c246 bl[246] br[246] wl[109] vdd gnd cell_6t
Xbit_r110_c246 bl[246] br[246] wl[110] vdd gnd cell_6t
Xbit_r111_c246 bl[246] br[246] wl[111] vdd gnd cell_6t
Xbit_r112_c246 bl[246] br[246] wl[112] vdd gnd cell_6t
Xbit_r113_c246 bl[246] br[246] wl[113] vdd gnd cell_6t
Xbit_r114_c246 bl[246] br[246] wl[114] vdd gnd cell_6t
Xbit_r115_c246 bl[246] br[246] wl[115] vdd gnd cell_6t
Xbit_r116_c246 bl[246] br[246] wl[116] vdd gnd cell_6t
Xbit_r117_c246 bl[246] br[246] wl[117] vdd gnd cell_6t
Xbit_r118_c246 bl[246] br[246] wl[118] vdd gnd cell_6t
Xbit_r119_c246 bl[246] br[246] wl[119] vdd gnd cell_6t
Xbit_r120_c246 bl[246] br[246] wl[120] vdd gnd cell_6t
Xbit_r121_c246 bl[246] br[246] wl[121] vdd gnd cell_6t
Xbit_r122_c246 bl[246] br[246] wl[122] vdd gnd cell_6t
Xbit_r123_c246 bl[246] br[246] wl[123] vdd gnd cell_6t
Xbit_r124_c246 bl[246] br[246] wl[124] vdd gnd cell_6t
Xbit_r125_c246 bl[246] br[246] wl[125] vdd gnd cell_6t
Xbit_r126_c246 bl[246] br[246] wl[126] vdd gnd cell_6t
Xbit_r127_c246 bl[246] br[246] wl[127] vdd gnd cell_6t
Xbit_r0_c247 bl[247] br[247] wl[0] vdd gnd cell_6t
Xbit_r1_c247 bl[247] br[247] wl[1] vdd gnd cell_6t
Xbit_r2_c247 bl[247] br[247] wl[2] vdd gnd cell_6t
Xbit_r3_c247 bl[247] br[247] wl[3] vdd gnd cell_6t
Xbit_r4_c247 bl[247] br[247] wl[4] vdd gnd cell_6t
Xbit_r5_c247 bl[247] br[247] wl[5] vdd gnd cell_6t
Xbit_r6_c247 bl[247] br[247] wl[6] vdd gnd cell_6t
Xbit_r7_c247 bl[247] br[247] wl[7] vdd gnd cell_6t
Xbit_r8_c247 bl[247] br[247] wl[8] vdd gnd cell_6t
Xbit_r9_c247 bl[247] br[247] wl[9] vdd gnd cell_6t
Xbit_r10_c247 bl[247] br[247] wl[10] vdd gnd cell_6t
Xbit_r11_c247 bl[247] br[247] wl[11] vdd gnd cell_6t
Xbit_r12_c247 bl[247] br[247] wl[12] vdd gnd cell_6t
Xbit_r13_c247 bl[247] br[247] wl[13] vdd gnd cell_6t
Xbit_r14_c247 bl[247] br[247] wl[14] vdd gnd cell_6t
Xbit_r15_c247 bl[247] br[247] wl[15] vdd gnd cell_6t
Xbit_r16_c247 bl[247] br[247] wl[16] vdd gnd cell_6t
Xbit_r17_c247 bl[247] br[247] wl[17] vdd gnd cell_6t
Xbit_r18_c247 bl[247] br[247] wl[18] vdd gnd cell_6t
Xbit_r19_c247 bl[247] br[247] wl[19] vdd gnd cell_6t
Xbit_r20_c247 bl[247] br[247] wl[20] vdd gnd cell_6t
Xbit_r21_c247 bl[247] br[247] wl[21] vdd gnd cell_6t
Xbit_r22_c247 bl[247] br[247] wl[22] vdd gnd cell_6t
Xbit_r23_c247 bl[247] br[247] wl[23] vdd gnd cell_6t
Xbit_r24_c247 bl[247] br[247] wl[24] vdd gnd cell_6t
Xbit_r25_c247 bl[247] br[247] wl[25] vdd gnd cell_6t
Xbit_r26_c247 bl[247] br[247] wl[26] vdd gnd cell_6t
Xbit_r27_c247 bl[247] br[247] wl[27] vdd gnd cell_6t
Xbit_r28_c247 bl[247] br[247] wl[28] vdd gnd cell_6t
Xbit_r29_c247 bl[247] br[247] wl[29] vdd gnd cell_6t
Xbit_r30_c247 bl[247] br[247] wl[30] vdd gnd cell_6t
Xbit_r31_c247 bl[247] br[247] wl[31] vdd gnd cell_6t
Xbit_r32_c247 bl[247] br[247] wl[32] vdd gnd cell_6t
Xbit_r33_c247 bl[247] br[247] wl[33] vdd gnd cell_6t
Xbit_r34_c247 bl[247] br[247] wl[34] vdd gnd cell_6t
Xbit_r35_c247 bl[247] br[247] wl[35] vdd gnd cell_6t
Xbit_r36_c247 bl[247] br[247] wl[36] vdd gnd cell_6t
Xbit_r37_c247 bl[247] br[247] wl[37] vdd gnd cell_6t
Xbit_r38_c247 bl[247] br[247] wl[38] vdd gnd cell_6t
Xbit_r39_c247 bl[247] br[247] wl[39] vdd gnd cell_6t
Xbit_r40_c247 bl[247] br[247] wl[40] vdd gnd cell_6t
Xbit_r41_c247 bl[247] br[247] wl[41] vdd gnd cell_6t
Xbit_r42_c247 bl[247] br[247] wl[42] vdd gnd cell_6t
Xbit_r43_c247 bl[247] br[247] wl[43] vdd gnd cell_6t
Xbit_r44_c247 bl[247] br[247] wl[44] vdd gnd cell_6t
Xbit_r45_c247 bl[247] br[247] wl[45] vdd gnd cell_6t
Xbit_r46_c247 bl[247] br[247] wl[46] vdd gnd cell_6t
Xbit_r47_c247 bl[247] br[247] wl[47] vdd gnd cell_6t
Xbit_r48_c247 bl[247] br[247] wl[48] vdd gnd cell_6t
Xbit_r49_c247 bl[247] br[247] wl[49] vdd gnd cell_6t
Xbit_r50_c247 bl[247] br[247] wl[50] vdd gnd cell_6t
Xbit_r51_c247 bl[247] br[247] wl[51] vdd gnd cell_6t
Xbit_r52_c247 bl[247] br[247] wl[52] vdd gnd cell_6t
Xbit_r53_c247 bl[247] br[247] wl[53] vdd gnd cell_6t
Xbit_r54_c247 bl[247] br[247] wl[54] vdd gnd cell_6t
Xbit_r55_c247 bl[247] br[247] wl[55] vdd gnd cell_6t
Xbit_r56_c247 bl[247] br[247] wl[56] vdd gnd cell_6t
Xbit_r57_c247 bl[247] br[247] wl[57] vdd gnd cell_6t
Xbit_r58_c247 bl[247] br[247] wl[58] vdd gnd cell_6t
Xbit_r59_c247 bl[247] br[247] wl[59] vdd gnd cell_6t
Xbit_r60_c247 bl[247] br[247] wl[60] vdd gnd cell_6t
Xbit_r61_c247 bl[247] br[247] wl[61] vdd gnd cell_6t
Xbit_r62_c247 bl[247] br[247] wl[62] vdd gnd cell_6t
Xbit_r63_c247 bl[247] br[247] wl[63] vdd gnd cell_6t
Xbit_r64_c247 bl[247] br[247] wl[64] vdd gnd cell_6t
Xbit_r65_c247 bl[247] br[247] wl[65] vdd gnd cell_6t
Xbit_r66_c247 bl[247] br[247] wl[66] vdd gnd cell_6t
Xbit_r67_c247 bl[247] br[247] wl[67] vdd gnd cell_6t
Xbit_r68_c247 bl[247] br[247] wl[68] vdd gnd cell_6t
Xbit_r69_c247 bl[247] br[247] wl[69] vdd gnd cell_6t
Xbit_r70_c247 bl[247] br[247] wl[70] vdd gnd cell_6t
Xbit_r71_c247 bl[247] br[247] wl[71] vdd gnd cell_6t
Xbit_r72_c247 bl[247] br[247] wl[72] vdd gnd cell_6t
Xbit_r73_c247 bl[247] br[247] wl[73] vdd gnd cell_6t
Xbit_r74_c247 bl[247] br[247] wl[74] vdd gnd cell_6t
Xbit_r75_c247 bl[247] br[247] wl[75] vdd gnd cell_6t
Xbit_r76_c247 bl[247] br[247] wl[76] vdd gnd cell_6t
Xbit_r77_c247 bl[247] br[247] wl[77] vdd gnd cell_6t
Xbit_r78_c247 bl[247] br[247] wl[78] vdd gnd cell_6t
Xbit_r79_c247 bl[247] br[247] wl[79] vdd gnd cell_6t
Xbit_r80_c247 bl[247] br[247] wl[80] vdd gnd cell_6t
Xbit_r81_c247 bl[247] br[247] wl[81] vdd gnd cell_6t
Xbit_r82_c247 bl[247] br[247] wl[82] vdd gnd cell_6t
Xbit_r83_c247 bl[247] br[247] wl[83] vdd gnd cell_6t
Xbit_r84_c247 bl[247] br[247] wl[84] vdd gnd cell_6t
Xbit_r85_c247 bl[247] br[247] wl[85] vdd gnd cell_6t
Xbit_r86_c247 bl[247] br[247] wl[86] vdd gnd cell_6t
Xbit_r87_c247 bl[247] br[247] wl[87] vdd gnd cell_6t
Xbit_r88_c247 bl[247] br[247] wl[88] vdd gnd cell_6t
Xbit_r89_c247 bl[247] br[247] wl[89] vdd gnd cell_6t
Xbit_r90_c247 bl[247] br[247] wl[90] vdd gnd cell_6t
Xbit_r91_c247 bl[247] br[247] wl[91] vdd gnd cell_6t
Xbit_r92_c247 bl[247] br[247] wl[92] vdd gnd cell_6t
Xbit_r93_c247 bl[247] br[247] wl[93] vdd gnd cell_6t
Xbit_r94_c247 bl[247] br[247] wl[94] vdd gnd cell_6t
Xbit_r95_c247 bl[247] br[247] wl[95] vdd gnd cell_6t
Xbit_r96_c247 bl[247] br[247] wl[96] vdd gnd cell_6t
Xbit_r97_c247 bl[247] br[247] wl[97] vdd gnd cell_6t
Xbit_r98_c247 bl[247] br[247] wl[98] vdd gnd cell_6t
Xbit_r99_c247 bl[247] br[247] wl[99] vdd gnd cell_6t
Xbit_r100_c247 bl[247] br[247] wl[100] vdd gnd cell_6t
Xbit_r101_c247 bl[247] br[247] wl[101] vdd gnd cell_6t
Xbit_r102_c247 bl[247] br[247] wl[102] vdd gnd cell_6t
Xbit_r103_c247 bl[247] br[247] wl[103] vdd gnd cell_6t
Xbit_r104_c247 bl[247] br[247] wl[104] vdd gnd cell_6t
Xbit_r105_c247 bl[247] br[247] wl[105] vdd gnd cell_6t
Xbit_r106_c247 bl[247] br[247] wl[106] vdd gnd cell_6t
Xbit_r107_c247 bl[247] br[247] wl[107] vdd gnd cell_6t
Xbit_r108_c247 bl[247] br[247] wl[108] vdd gnd cell_6t
Xbit_r109_c247 bl[247] br[247] wl[109] vdd gnd cell_6t
Xbit_r110_c247 bl[247] br[247] wl[110] vdd gnd cell_6t
Xbit_r111_c247 bl[247] br[247] wl[111] vdd gnd cell_6t
Xbit_r112_c247 bl[247] br[247] wl[112] vdd gnd cell_6t
Xbit_r113_c247 bl[247] br[247] wl[113] vdd gnd cell_6t
Xbit_r114_c247 bl[247] br[247] wl[114] vdd gnd cell_6t
Xbit_r115_c247 bl[247] br[247] wl[115] vdd gnd cell_6t
Xbit_r116_c247 bl[247] br[247] wl[116] vdd gnd cell_6t
Xbit_r117_c247 bl[247] br[247] wl[117] vdd gnd cell_6t
Xbit_r118_c247 bl[247] br[247] wl[118] vdd gnd cell_6t
Xbit_r119_c247 bl[247] br[247] wl[119] vdd gnd cell_6t
Xbit_r120_c247 bl[247] br[247] wl[120] vdd gnd cell_6t
Xbit_r121_c247 bl[247] br[247] wl[121] vdd gnd cell_6t
Xbit_r122_c247 bl[247] br[247] wl[122] vdd gnd cell_6t
Xbit_r123_c247 bl[247] br[247] wl[123] vdd gnd cell_6t
Xbit_r124_c247 bl[247] br[247] wl[124] vdd gnd cell_6t
Xbit_r125_c247 bl[247] br[247] wl[125] vdd gnd cell_6t
Xbit_r126_c247 bl[247] br[247] wl[126] vdd gnd cell_6t
Xbit_r127_c247 bl[247] br[247] wl[127] vdd gnd cell_6t
Xbit_r0_c248 bl[248] br[248] wl[0] vdd gnd cell_6t
Xbit_r1_c248 bl[248] br[248] wl[1] vdd gnd cell_6t
Xbit_r2_c248 bl[248] br[248] wl[2] vdd gnd cell_6t
Xbit_r3_c248 bl[248] br[248] wl[3] vdd gnd cell_6t
Xbit_r4_c248 bl[248] br[248] wl[4] vdd gnd cell_6t
Xbit_r5_c248 bl[248] br[248] wl[5] vdd gnd cell_6t
Xbit_r6_c248 bl[248] br[248] wl[6] vdd gnd cell_6t
Xbit_r7_c248 bl[248] br[248] wl[7] vdd gnd cell_6t
Xbit_r8_c248 bl[248] br[248] wl[8] vdd gnd cell_6t
Xbit_r9_c248 bl[248] br[248] wl[9] vdd gnd cell_6t
Xbit_r10_c248 bl[248] br[248] wl[10] vdd gnd cell_6t
Xbit_r11_c248 bl[248] br[248] wl[11] vdd gnd cell_6t
Xbit_r12_c248 bl[248] br[248] wl[12] vdd gnd cell_6t
Xbit_r13_c248 bl[248] br[248] wl[13] vdd gnd cell_6t
Xbit_r14_c248 bl[248] br[248] wl[14] vdd gnd cell_6t
Xbit_r15_c248 bl[248] br[248] wl[15] vdd gnd cell_6t
Xbit_r16_c248 bl[248] br[248] wl[16] vdd gnd cell_6t
Xbit_r17_c248 bl[248] br[248] wl[17] vdd gnd cell_6t
Xbit_r18_c248 bl[248] br[248] wl[18] vdd gnd cell_6t
Xbit_r19_c248 bl[248] br[248] wl[19] vdd gnd cell_6t
Xbit_r20_c248 bl[248] br[248] wl[20] vdd gnd cell_6t
Xbit_r21_c248 bl[248] br[248] wl[21] vdd gnd cell_6t
Xbit_r22_c248 bl[248] br[248] wl[22] vdd gnd cell_6t
Xbit_r23_c248 bl[248] br[248] wl[23] vdd gnd cell_6t
Xbit_r24_c248 bl[248] br[248] wl[24] vdd gnd cell_6t
Xbit_r25_c248 bl[248] br[248] wl[25] vdd gnd cell_6t
Xbit_r26_c248 bl[248] br[248] wl[26] vdd gnd cell_6t
Xbit_r27_c248 bl[248] br[248] wl[27] vdd gnd cell_6t
Xbit_r28_c248 bl[248] br[248] wl[28] vdd gnd cell_6t
Xbit_r29_c248 bl[248] br[248] wl[29] vdd gnd cell_6t
Xbit_r30_c248 bl[248] br[248] wl[30] vdd gnd cell_6t
Xbit_r31_c248 bl[248] br[248] wl[31] vdd gnd cell_6t
Xbit_r32_c248 bl[248] br[248] wl[32] vdd gnd cell_6t
Xbit_r33_c248 bl[248] br[248] wl[33] vdd gnd cell_6t
Xbit_r34_c248 bl[248] br[248] wl[34] vdd gnd cell_6t
Xbit_r35_c248 bl[248] br[248] wl[35] vdd gnd cell_6t
Xbit_r36_c248 bl[248] br[248] wl[36] vdd gnd cell_6t
Xbit_r37_c248 bl[248] br[248] wl[37] vdd gnd cell_6t
Xbit_r38_c248 bl[248] br[248] wl[38] vdd gnd cell_6t
Xbit_r39_c248 bl[248] br[248] wl[39] vdd gnd cell_6t
Xbit_r40_c248 bl[248] br[248] wl[40] vdd gnd cell_6t
Xbit_r41_c248 bl[248] br[248] wl[41] vdd gnd cell_6t
Xbit_r42_c248 bl[248] br[248] wl[42] vdd gnd cell_6t
Xbit_r43_c248 bl[248] br[248] wl[43] vdd gnd cell_6t
Xbit_r44_c248 bl[248] br[248] wl[44] vdd gnd cell_6t
Xbit_r45_c248 bl[248] br[248] wl[45] vdd gnd cell_6t
Xbit_r46_c248 bl[248] br[248] wl[46] vdd gnd cell_6t
Xbit_r47_c248 bl[248] br[248] wl[47] vdd gnd cell_6t
Xbit_r48_c248 bl[248] br[248] wl[48] vdd gnd cell_6t
Xbit_r49_c248 bl[248] br[248] wl[49] vdd gnd cell_6t
Xbit_r50_c248 bl[248] br[248] wl[50] vdd gnd cell_6t
Xbit_r51_c248 bl[248] br[248] wl[51] vdd gnd cell_6t
Xbit_r52_c248 bl[248] br[248] wl[52] vdd gnd cell_6t
Xbit_r53_c248 bl[248] br[248] wl[53] vdd gnd cell_6t
Xbit_r54_c248 bl[248] br[248] wl[54] vdd gnd cell_6t
Xbit_r55_c248 bl[248] br[248] wl[55] vdd gnd cell_6t
Xbit_r56_c248 bl[248] br[248] wl[56] vdd gnd cell_6t
Xbit_r57_c248 bl[248] br[248] wl[57] vdd gnd cell_6t
Xbit_r58_c248 bl[248] br[248] wl[58] vdd gnd cell_6t
Xbit_r59_c248 bl[248] br[248] wl[59] vdd gnd cell_6t
Xbit_r60_c248 bl[248] br[248] wl[60] vdd gnd cell_6t
Xbit_r61_c248 bl[248] br[248] wl[61] vdd gnd cell_6t
Xbit_r62_c248 bl[248] br[248] wl[62] vdd gnd cell_6t
Xbit_r63_c248 bl[248] br[248] wl[63] vdd gnd cell_6t
Xbit_r64_c248 bl[248] br[248] wl[64] vdd gnd cell_6t
Xbit_r65_c248 bl[248] br[248] wl[65] vdd gnd cell_6t
Xbit_r66_c248 bl[248] br[248] wl[66] vdd gnd cell_6t
Xbit_r67_c248 bl[248] br[248] wl[67] vdd gnd cell_6t
Xbit_r68_c248 bl[248] br[248] wl[68] vdd gnd cell_6t
Xbit_r69_c248 bl[248] br[248] wl[69] vdd gnd cell_6t
Xbit_r70_c248 bl[248] br[248] wl[70] vdd gnd cell_6t
Xbit_r71_c248 bl[248] br[248] wl[71] vdd gnd cell_6t
Xbit_r72_c248 bl[248] br[248] wl[72] vdd gnd cell_6t
Xbit_r73_c248 bl[248] br[248] wl[73] vdd gnd cell_6t
Xbit_r74_c248 bl[248] br[248] wl[74] vdd gnd cell_6t
Xbit_r75_c248 bl[248] br[248] wl[75] vdd gnd cell_6t
Xbit_r76_c248 bl[248] br[248] wl[76] vdd gnd cell_6t
Xbit_r77_c248 bl[248] br[248] wl[77] vdd gnd cell_6t
Xbit_r78_c248 bl[248] br[248] wl[78] vdd gnd cell_6t
Xbit_r79_c248 bl[248] br[248] wl[79] vdd gnd cell_6t
Xbit_r80_c248 bl[248] br[248] wl[80] vdd gnd cell_6t
Xbit_r81_c248 bl[248] br[248] wl[81] vdd gnd cell_6t
Xbit_r82_c248 bl[248] br[248] wl[82] vdd gnd cell_6t
Xbit_r83_c248 bl[248] br[248] wl[83] vdd gnd cell_6t
Xbit_r84_c248 bl[248] br[248] wl[84] vdd gnd cell_6t
Xbit_r85_c248 bl[248] br[248] wl[85] vdd gnd cell_6t
Xbit_r86_c248 bl[248] br[248] wl[86] vdd gnd cell_6t
Xbit_r87_c248 bl[248] br[248] wl[87] vdd gnd cell_6t
Xbit_r88_c248 bl[248] br[248] wl[88] vdd gnd cell_6t
Xbit_r89_c248 bl[248] br[248] wl[89] vdd gnd cell_6t
Xbit_r90_c248 bl[248] br[248] wl[90] vdd gnd cell_6t
Xbit_r91_c248 bl[248] br[248] wl[91] vdd gnd cell_6t
Xbit_r92_c248 bl[248] br[248] wl[92] vdd gnd cell_6t
Xbit_r93_c248 bl[248] br[248] wl[93] vdd gnd cell_6t
Xbit_r94_c248 bl[248] br[248] wl[94] vdd gnd cell_6t
Xbit_r95_c248 bl[248] br[248] wl[95] vdd gnd cell_6t
Xbit_r96_c248 bl[248] br[248] wl[96] vdd gnd cell_6t
Xbit_r97_c248 bl[248] br[248] wl[97] vdd gnd cell_6t
Xbit_r98_c248 bl[248] br[248] wl[98] vdd gnd cell_6t
Xbit_r99_c248 bl[248] br[248] wl[99] vdd gnd cell_6t
Xbit_r100_c248 bl[248] br[248] wl[100] vdd gnd cell_6t
Xbit_r101_c248 bl[248] br[248] wl[101] vdd gnd cell_6t
Xbit_r102_c248 bl[248] br[248] wl[102] vdd gnd cell_6t
Xbit_r103_c248 bl[248] br[248] wl[103] vdd gnd cell_6t
Xbit_r104_c248 bl[248] br[248] wl[104] vdd gnd cell_6t
Xbit_r105_c248 bl[248] br[248] wl[105] vdd gnd cell_6t
Xbit_r106_c248 bl[248] br[248] wl[106] vdd gnd cell_6t
Xbit_r107_c248 bl[248] br[248] wl[107] vdd gnd cell_6t
Xbit_r108_c248 bl[248] br[248] wl[108] vdd gnd cell_6t
Xbit_r109_c248 bl[248] br[248] wl[109] vdd gnd cell_6t
Xbit_r110_c248 bl[248] br[248] wl[110] vdd gnd cell_6t
Xbit_r111_c248 bl[248] br[248] wl[111] vdd gnd cell_6t
Xbit_r112_c248 bl[248] br[248] wl[112] vdd gnd cell_6t
Xbit_r113_c248 bl[248] br[248] wl[113] vdd gnd cell_6t
Xbit_r114_c248 bl[248] br[248] wl[114] vdd gnd cell_6t
Xbit_r115_c248 bl[248] br[248] wl[115] vdd gnd cell_6t
Xbit_r116_c248 bl[248] br[248] wl[116] vdd gnd cell_6t
Xbit_r117_c248 bl[248] br[248] wl[117] vdd gnd cell_6t
Xbit_r118_c248 bl[248] br[248] wl[118] vdd gnd cell_6t
Xbit_r119_c248 bl[248] br[248] wl[119] vdd gnd cell_6t
Xbit_r120_c248 bl[248] br[248] wl[120] vdd gnd cell_6t
Xbit_r121_c248 bl[248] br[248] wl[121] vdd gnd cell_6t
Xbit_r122_c248 bl[248] br[248] wl[122] vdd gnd cell_6t
Xbit_r123_c248 bl[248] br[248] wl[123] vdd gnd cell_6t
Xbit_r124_c248 bl[248] br[248] wl[124] vdd gnd cell_6t
Xbit_r125_c248 bl[248] br[248] wl[125] vdd gnd cell_6t
Xbit_r126_c248 bl[248] br[248] wl[126] vdd gnd cell_6t
Xbit_r127_c248 bl[248] br[248] wl[127] vdd gnd cell_6t
Xbit_r0_c249 bl[249] br[249] wl[0] vdd gnd cell_6t
Xbit_r1_c249 bl[249] br[249] wl[1] vdd gnd cell_6t
Xbit_r2_c249 bl[249] br[249] wl[2] vdd gnd cell_6t
Xbit_r3_c249 bl[249] br[249] wl[3] vdd gnd cell_6t
Xbit_r4_c249 bl[249] br[249] wl[4] vdd gnd cell_6t
Xbit_r5_c249 bl[249] br[249] wl[5] vdd gnd cell_6t
Xbit_r6_c249 bl[249] br[249] wl[6] vdd gnd cell_6t
Xbit_r7_c249 bl[249] br[249] wl[7] vdd gnd cell_6t
Xbit_r8_c249 bl[249] br[249] wl[8] vdd gnd cell_6t
Xbit_r9_c249 bl[249] br[249] wl[9] vdd gnd cell_6t
Xbit_r10_c249 bl[249] br[249] wl[10] vdd gnd cell_6t
Xbit_r11_c249 bl[249] br[249] wl[11] vdd gnd cell_6t
Xbit_r12_c249 bl[249] br[249] wl[12] vdd gnd cell_6t
Xbit_r13_c249 bl[249] br[249] wl[13] vdd gnd cell_6t
Xbit_r14_c249 bl[249] br[249] wl[14] vdd gnd cell_6t
Xbit_r15_c249 bl[249] br[249] wl[15] vdd gnd cell_6t
Xbit_r16_c249 bl[249] br[249] wl[16] vdd gnd cell_6t
Xbit_r17_c249 bl[249] br[249] wl[17] vdd gnd cell_6t
Xbit_r18_c249 bl[249] br[249] wl[18] vdd gnd cell_6t
Xbit_r19_c249 bl[249] br[249] wl[19] vdd gnd cell_6t
Xbit_r20_c249 bl[249] br[249] wl[20] vdd gnd cell_6t
Xbit_r21_c249 bl[249] br[249] wl[21] vdd gnd cell_6t
Xbit_r22_c249 bl[249] br[249] wl[22] vdd gnd cell_6t
Xbit_r23_c249 bl[249] br[249] wl[23] vdd gnd cell_6t
Xbit_r24_c249 bl[249] br[249] wl[24] vdd gnd cell_6t
Xbit_r25_c249 bl[249] br[249] wl[25] vdd gnd cell_6t
Xbit_r26_c249 bl[249] br[249] wl[26] vdd gnd cell_6t
Xbit_r27_c249 bl[249] br[249] wl[27] vdd gnd cell_6t
Xbit_r28_c249 bl[249] br[249] wl[28] vdd gnd cell_6t
Xbit_r29_c249 bl[249] br[249] wl[29] vdd gnd cell_6t
Xbit_r30_c249 bl[249] br[249] wl[30] vdd gnd cell_6t
Xbit_r31_c249 bl[249] br[249] wl[31] vdd gnd cell_6t
Xbit_r32_c249 bl[249] br[249] wl[32] vdd gnd cell_6t
Xbit_r33_c249 bl[249] br[249] wl[33] vdd gnd cell_6t
Xbit_r34_c249 bl[249] br[249] wl[34] vdd gnd cell_6t
Xbit_r35_c249 bl[249] br[249] wl[35] vdd gnd cell_6t
Xbit_r36_c249 bl[249] br[249] wl[36] vdd gnd cell_6t
Xbit_r37_c249 bl[249] br[249] wl[37] vdd gnd cell_6t
Xbit_r38_c249 bl[249] br[249] wl[38] vdd gnd cell_6t
Xbit_r39_c249 bl[249] br[249] wl[39] vdd gnd cell_6t
Xbit_r40_c249 bl[249] br[249] wl[40] vdd gnd cell_6t
Xbit_r41_c249 bl[249] br[249] wl[41] vdd gnd cell_6t
Xbit_r42_c249 bl[249] br[249] wl[42] vdd gnd cell_6t
Xbit_r43_c249 bl[249] br[249] wl[43] vdd gnd cell_6t
Xbit_r44_c249 bl[249] br[249] wl[44] vdd gnd cell_6t
Xbit_r45_c249 bl[249] br[249] wl[45] vdd gnd cell_6t
Xbit_r46_c249 bl[249] br[249] wl[46] vdd gnd cell_6t
Xbit_r47_c249 bl[249] br[249] wl[47] vdd gnd cell_6t
Xbit_r48_c249 bl[249] br[249] wl[48] vdd gnd cell_6t
Xbit_r49_c249 bl[249] br[249] wl[49] vdd gnd cell_6t
Xbit_r50_c249 bl[249] br[249] wl[50] vdd gnd cell_6t
Xbit_r51_c249 bl[249] br[249] wl[51] vdd gnd cell_6t
Xbit_r52_c249 bl[249] br[249] wl[52] vdd gnd cell_6t
Xbit_r53_c249 bl[249] br[249] wl[53] vdd gnd cell_6t
Xbit_r54_c249 bl[249] br[249] wl[54] vdd gnd cell_6t
Xbit_r55_c249 bl[249] br[249] wl[55] vdd gnd cell_6t
Xbit_r56_c249 bl[249] br[249] wl[56] vdd gnd cell_6t
Xbit_r57_c249 bl[249] br[249] wl[57] vdd gnd cell_6t
Xbit_r58_c249 bl[249] br[249] wl[58] vdd gnd cell_6t
Xbit_r59_c249 bl[249] br[249] wl[59] vdd gnd cell_6t
Xbit_r60_c249 bl[249] br[249] wl[60] vdd gnd cell_6t
Xbit_r61_c249 bl[249] br[249] wl[61] vdd gnd cell_6t
Xbit_r62_c249 bl[249] br[249] wl[62] vdd gnd cell_6t
Xbit_r63_c249 bl[249] br[249] wl[63] vdd gnd cell_6t
Xbit_r64_c249 bl[249] br[249] wl[64] vdd gnd cell_6t
Xbit_r65_c249 bl[249] br[249] wl[65] vdd gnd cell_6t
Xbit_r66_c249 bl[249] br[249] wl[66] vdd gnd cell_6t
Xbit_r67_c249 bl[249] br[249] wl[67] vdd gnd cell_6t
Xbit_r68_c249 bl[249] br[249] wl[68] vdd gnd cell_6t
Xbit_r69_c249 bl[249] br[249] wl[69] vdd gnd cell_6t
Xbit_r70_c249 bl[249] br[249] wl[70] vdd gnd cell_6t
Xbit_r71_c249 bl[249] br[249] wl[71] vdd gnd cell_6t
Xbit_r72_c249 bl[249] br[249] wl[72] vdd gnd cell_6t
Xbit_r73_c249 bl[249] br[249] wl[73] vdd gnd cell_6t
Xbit_r74_c249 bl[249] br[249] wl[74] vdd gnd cell_6t
Xbit_r75_c249 bl[249] br[249] wl[75] vdd gnd cell_6t
Xbit_r76_c249 bl[249] br[249] wl[76] vdd gnd cell_6t
Xbit_r77_c249 bl[249] br[249] wl[77] vdd gnd cell_6t
Xbit_r78_c249 bl[249] br[249] wl[78] vdd gnd cell_6t
Xbit_r79_c249 bl[249] br[249] wl[79] vdd gnd cell_6t
Xbit_r80_c249 bl[249] br[249] wl[80] vdd gnd cell_6t
Xbit_r81_c249 bl[249] br[249] wl[81] vdd gnd cell_6t
Xbit_r82_c249 bl[249] br[249] wl[82] vdd gnd cell_6t
Xbit_r83_c249 bl[249] br[249] wl[83] vdd gnd cell_6t
Xbit_r84_c249 bl[249] br[249] wl[84] vdd gnd cell_6t
Xbit_r85_c249 bl[249] br[249] wl[85] vdd gnd cell_6t
Xbit_r86_c249 bl[249] br[249] wl[86] vdd gnd cell_6t
Xbit_r87_c249 bl[249] br[249] wl[87] vdd gnd cell_6t
Xbit_r88_c249 bl[249] br[249] wl[88] vdd gnd cell_6t
Xbit_r89_c249 bl[249] br[249] wl[89] vdd gnd cell_6t
Xbit_r90_c249 bl[249] br[249] wl[90] vdd gnd cell_6t
Xbit_r91_c249 bl[249] br[249] wl[91] vdd gnd cell_6t
Xbit_r92_c249 bl[249] br[249] wl[92] vdd gnd cell_6t
Xbit_r93_c249 bl[249] br[249] wl[93] vdd gnd cell_6t
Xbit_r94_c249 bl[249] br[249] wl[94] vdd gnd cell_6t
Xbit_r95_c249 bl[249] br[249] wl[95] vdd gnd cell_6t
Xbit_r96_c249 bl[249] br[249] wl[96] vdd gnd cell_6t
Xbit_r97_c249 bl[249] br[249] wl[97] vdd gnd cell_6t
Xbit_r98_c249 bl[249] br[249] wl[98] vdd gnd cell_6t
Xbit_r99_c249 bl[249] br[249] wl[99] vdd gnd cell_6t
Xbit_r100_c249 bl[249] br[249] wl[100] vdd gnd cell_6t
Xbit_r101_c249 bl[249] br[249] wl[101] vdd gnd cell_6t
Xbit_r102_c249 bl[249] br[249] wl[102] vdd gnd cell_6t
Xbit_r103_c249 bl[249] br[249] wl[103] vdd gnd cell_6t
Xbit_r104_c249 bl[249] br[249] wl[104] vdd gnd cell_6t
Xbit_r105_c249 bl[249] br[249] wl[105] vdd gnd cell_6t
Xbit_r106_c249 bl[249] br[249] wl[106] vdd gnd cell_6t
Xbit_r107_c249 bl[249] br[249] wl[107] vdd gnd cell_6t
Xbit_r108_c249 bl[249] br[249] wl[108] vdd gnd cell_6t
Xbit_r109_c249 bl[249] br[249] wl[109] vdd gnd cell_6t
Xbit_r110_c249 bl[249] br[249] wl[110] vdd gnd cell_6t
Xbit_r111_c249 bl[249] br[249] wl[111] vdd gnd cell_6t
Xbit_r112_c249 bl[249] br[249] wl[112] vdd gnd cell_6t
Xbit_r113_c249 bl[249] br[249] wl[113] vdd gnd cell_6t
Xbit_r114_c249 bl[249] br[249] wl[114] vdd gnd cell_6t
Xbit_r115_c249 bl[249] br[249] wl[115] vdd gnd cell_6t
Xbit_r116_c249 bl[249] br[249] wl[116] vdd gnd cell_6t
Xbit_r117_c249 bl[249] br[249] wl[117] vdd gnd cell_6t
Xbit_r118_c249 bl[249] br[249] wl[118] vdd gnd cell_6t
Xbit_r119_c249 bl[249] br[249] wl[119] vdd gnd cell_6t
Xbit_r120_c249 bl[249] br[249] wl[120] vdd gnd cell_6t
Xbit_r121_c249 bl[249] br[249] wl[121] vdd gnd cell_6t
Xbit_r122_c249 bl[249] br[249] wl[122] vdd gnd cell_6t
Xbit_r123_c249 bl[249] br[249] wl[123] vdd gnd cell_6t
Xbit_r124_c249 bl[249] br[249] wl[124] vdd gnd cell_6t
Xbit_r125_c249 bl[249] br[249] wl[125] vdd gnd cell_6t
Xbit_r126_c249 bl[249] br[249] wl[126] vdd gnd cell_6t
Xbit_r127_c249 bl[249] br[249] wl[127] vdd gnd cell_6t
Xbit_r0_c250 bl[250] br[250] wl[0] vdd gnd cell_6t
Xbit_r1_c250 bl[250] br[250] wl[1] vdd gnd cell_6t
Xbit_r2_c250 bl[250] br[250] wl[2] vdd gnd cell_6t
Xbit_r3_c250 bl[250] br[250] wl[3] vdd gnd cell_6t
Xbit_r4_c250 bl[250] br[250] wl[4] vdd gnd cell_6t
Xbit_r5_c250 bl[250] br[250] wl[5] vdd gnd cell_6t
Xbit_r6_c250 bl[250] br[250] wl[6] vdd gnd cell_6t
Xbit_r7_c250 bl[250] br[250] wl[7] vdd gnd cell_6t
Xbit_r8_c250 bl[250] br[250] wl[8] vdd gnd cell_6t
Xbit_r9_c250 bl[250] br[250] wl[9] vdd gnd cell_6t
Xbit_r10_c250 bl[250] br[250] wl[10] vdd gnd cell_6t
Xbit_r11_c250 bl[250] br[250] wl[11] vdd gnd cell_6t
Xbit_r12_c250 bl[250] br[250] wl[12] vdd gnd cell_6t
Xbit_r13_c250 bl[250] br[250] wl[13] vdd gnd cell_6t
Xbit_r14_c250 bl[250] br[250] wl[14] vdd gnd cell_6t
Xbit_r15_c250 bl[250] br[250] wl[15] vdd gnd cell_6t
Xbit_r16_c250 bl[250] br[250] wl[16] vdd gnd cell_6t
Xbit_r17_c250 bl[250] br[250] wl[17] vdd gnd cell_6t
Xbit_r18_c250 bl[250] br[250] wl[18] vdd gnd cell_6t
Xbit_r19_c250 bl[250] br[250] wl[19] vdd gnd cell_6t
Xbit_r20_c250 bl[250] br[250] wl[20] vdd gnd cell_6t
Xbit_r21_c250 bl[250] br[250] wl[21] vdd gnd cell_6t
Xbit_r22_c250 bl[250] br[250] wl[22] vdd gnd cell_6t
Xbit_r23_c250 bl[250] br[250] wl[23] vdd gnd cell_6t
Xbit_r24_c250 bl[250] br[250] wl[24] vdd gnd cell_6t
Xbit_r25_c250 bl[250] br[250] wl[25] vdd gnd cell_6t
Xbit_r26_c250 bl[250] br[250] wl[26] vdd gnd cell_6t
Xbit_r27_c250 bl[250] br[250] wl[27] vdd gnd cell_6t
Xbit_r28_c250 bl[250] br[250] wl[28] vdd gnd cell_6t
Xbit_r29_c250 bl[250] br[250] wl[29] vdd gnd cell_6t
Xbit_r30_c250 bl[250] br[250] wl[30] vdd gnd cell_6t
Xbit_r31_c250 bl[250] br[250] wl[31] vdd gnd cell_6t
Xbit_r32_c250 bl[250] br[250] wl[32] vdd gnd cell_6t
Xbit_r33_c250 bl[250] br[250] wl[33] vdd gnd cell_6t
Xbit_r34_c250 bl[250] br[250] wl[34] vdd gnd cell_6t
Xbit_r35_c250 bl[250] br[250] wl[35] vdd gnd cell_6t
Xbit_r36_c250 bl[250] br[250] wl[36] vdd gnd cell_6t
Xbit_r37_c250 bl[250] br[250] wl[37] vdd gnd cell_6t
Xbit_r38_c250 bl[250] br[250] wl[38] vdd gnd cell_6t
Xbit_r39_c250 bl[250] br[250] wl[39] vdd gnd cell_6t
Xbit_r40_c250 bl[250] br[250] wl[40] vdd gnd cell_6t
Xbit_r41_c250 bl[250] br[250] wl[41] vdd gnd cell_6t
Xbit_r42_c250 bl[250] br[250] wl[42] vdd gnd cell_6t
Xbit_r43_c250 bl[250] br[250] wl[43] vdd gnd cell_6t
Xbit_r44_c250 bl[250] br[250] wl[44] vdd gnd cell_6t
Xbit_r45_c250 bl[250] br[250] wl[45] vdd gnd cell_6t
Xbit_r46_c250 bl[250] br[250] wl[46] vdd gnd cell_6t
Xbit_r47_c250 bl[250] br[250] wl[47] vdd gnd cell_6t
Xbit_r48_c250 bl[250] br[250] wl[48] vdd gnd cell_6t
Xbit_r49_c250 bl[250] br[250] wl[49] vdd gnd cell_6t
Xbit_r50_c250 bl[250] br[250] wl[50] vdd gnd cell_6t
Xbit_r51_c250 bl[250] br[250] wl[51] vdd gnd cell_6t
Xbit_r52_c250 bl[250] br[250] wl[52] vdd gnd cell_6t
Xbit_r53_c250 bl[250] br[250] wl[53] vdd gnd cell_6t
Xbit_r54_c250 bl[250] br[250] wl[54] vdd gnd cell_6t
Xbit_r55_c250 bl[250] br[250] wl[55] vdd gnd cell_6t
Xbit_r56_c250 bl[250] br[250] wl[56] vdd gnd cell_6t
Xbit_r57_c250 bl[250] br[250] wl[57] vdd gnd cell_6t
Xbit_r58_c250 bl[250] br[250] wl[58] vdd gnd cell_6t
Xbit_r59_c250 bl[250] br[250] wl[59] vdd gnd cell_6t
Xbit_r60_c250 bl[250] br[250] wl[60] vdd gnd cell_6t
Xbit_r61_c250 bl[250] br[250] wl[61] vdd gnd cell_6t
Xbit_r62_c250 bl[250] br[250] wl[62] vdd gnd cell_6t
Xbit_r63_c250 bl[250] br[250] wl[63] vdd gnd cell_6t
Xbit_r64_c250 bl[250] br[250] wl[64] vdd gnd cell_6t
Xbit_r65_c250 bl[250] br[250] wl[65] vdd gnd cell_6t
Xbit_r66_c250 bl[250] br[250] wl[66] vdd gnd cell_6t
Xbit_r67_c250 bl[250] br[250] wl[67] vdd gnd cell_6t
Xbit_r68_c250 bl[250] br[250] wl[68] vdd gnd cell_6t
Xbit_r69_c250 bl[250] br[250] wl[69] vdd gnd cell_6t
Xbit_r70_c250 bl[250] br[250] wl[70] vdd gnd cell_6t
Xbit_r71_c250 bl[250] br[250] wl[71] vdd gnd cell_6t
Xbit_r72_c250 bl[250] br[250] wl[72] vdd gnd cell_6t
Xbit_r73_c250 bl[250] br[250] wl[73] vdd gnd cell_6t
Xbit_r74_c250 bl[250] br[250] wl[74] vdd gnd cell_6t
Xbit_r75_c250 bl[250] br[250] wl[75] vdd gnd cell_6t
Xbit_r76_c250 bl[250] br[250] wl[76] vdd gnd cell_6t
Xbit_r77_c250 bl[250] br[250] wl[77] vdd gnd cell_6t
Xbit_r78_c250 bl[250] br[250] wl[78] vdd gnd cell_6t
Xbit_r79_c250 bl[250] br[250] wl[79] vdd gnd cell_6t
Xbit_r80_c250 bl[250] br[250] wl[80] vdd gnd cell_6t
Xbit_r81_c250 bl[250] br[250] wl[81] vdd gnd cell_6t
Xbit_r82_c250 bl[250] br[250] wl[82] vdd gnd cell_6t
Xbit_r83_c250 bl[250] br[250] wl[83] vdd gnd cell_6t
Xbit_r84_c250 bl[250] br[250] wl[84] vdd gnd cell_6t
Xbit_r85_c250 bl[250] br[250] wl[85] vdd gnd cell_6t
Xbit_r86_c250 bl[250] br[250] wl[86] vdd gnd cell_6t
Xbit_r87_c250 bl[250] br[250] wl[87] vdd gnd cell_6t
Xbit_r88_c250 bl[250] br[250] wl[88] vdd gnd cell_6t
Xbit_r89_c250 bl[250] br[250] wl[89] vdd gnd cell_6t
Xbit_r90_c250 bl[250] br[250] wl[90] vdd gnd cell_6t
Xbit_r91_c250 bl[250] br[250] wl[91] vdd gnd cell_6t
Xbit_r92_c250 bl[250] br[250] wl[92] vdd gnd cell_6t
Xbit_r93_c250 bl[250] br[250] wl[93] vdd gnd cell_6t
Xbit_r94_c250 bl[250] br[250] wl[94] vdd gnd cell_6t
Xbit_r95_c250 bl[250] br[250] wl[95] vdd gnd cell_6t
Xbit_r96_c250 bl[250] br[250] wl[96] vdd gnd cell_6t
Xbit_r97_c250 bl[250] br[250] wl[97] vdd gnd cell_6t
Xbit_r98_c250 bl[250] br[250] wl[98] vdd gnd cell_6t
Xbit_r99_c250 bl[250] br[250] wl[99] vdd gnd cell_6t
Xbit_r100_c250 bl[250] br[250] wl[100] vdd gnd cell_6t
Xbit_r101_c250 bl[250] br[250] wl[101] vdd gnd cell_6t
Xbit_r102_c250 bl[250] br[250] wl[102] vdd gnd cell_6t
Xbit_r103_c250 bl[250] br[250] wl[103] vdd gnd cell_6t
Xbit_r104_c250 bl[250] br[250] wl[104] vdd gnd cell_6t
Xbit_r105_c250 bl[250] br[250] wl[105] vdd gnd cell_6t
Xbit_r106_c250 bl[250] br[250] wl[106] vdd gnd cell_6t
Xbit_r107_c250 bl[250] br[250] wl[107] vdd gnd cell_6t
Xbit_r108_c250 bl[250] br[250] wl[108] vdd gnd cell_6t
Xbit_r109_c250 bl[250] br[250] wl[109] vdd gnd cell_6t
Xbit_r110_c250 bl[250] br[250] wl[110] vdd gnd cell_6t
Xbit_r111_c250 bl[250] br[250] wl[111] vdd gnd cell_6t
Xbit_r112_c250 bl[250] br[250] wl[112] vdd gnd cell_6t
Xbit_r113_c250 bl[250] br[250] wl[113] vdd gnd cell_6t
Xbit_r114_c250 bl[250] br[250] wl[114] vdd gnd cell_6t
Xbit_r115_c250 bl[250] br[250] wl[115] vdd gnd cell_6t
Xbit_r116_c250 bl[250] br[250] wl[116] vdd gnd cell_6t
Xbit_r117_c250 bl[250] br[250] wl[117] vdd gnd cell_6t
Xbit_r118_c250 bl[250] br[250] wl[118] vdd gnd cell_6t
Xbit_r119_c250 bl[250] br[250] wl[119] vdd gnd cell_6t
Xbit_r120_c250 bl[250] br[250] wl[120] vdd gnd cell_6t
Xbit_r121_c250 bl[250] br[250] wl[121] vdd gnd cell_6t
Xbit_r122_c250 bl[250] br[250] wl[122] vdd gnd cell_6t
Xbit_r123_c250 bl[250] br[250] wl[123] vdd gnd cell_6t
Xbit_r124_c250 bl[250] br[250] wl[124] vdd gnd cell_6t
Xbit_r125_c250 bl[250] br[250] wl[125] vdd gnd cell_6t
Xbit_r126_c250 bl[250] br[250] wl[126] vdd gnd cell_6t
Xbit_r127_c250 bl[250] br[250] wl[127] vdd gnd cell_6t
Xbit_r0_c251 bl[251] br[251] wl[0] vdd gnd cell_6t
Xbit_r1_c251 bl[251] br[251] wl[1] vdd gnd cell_6t
Xbit_r2_c251 bl[251] br[251] wl[2] vdd gnd cell_6t
Xbit_r3_c251 bl[251] br[251] wl[3] vdd gnd cell_6t
Xbit_r4_c251 bl[251] br[251] wl[4] vdd gnd cell_6t
Xbit_r5_c251 bl[251] br[251] wl[5] vdd gnd cell_6t
Xbit_r6_c251 bl[251] br[251] wl[6] vdd gnd cell_6t
Xbit_r7_c251 bl[251] br[251] wl[7] vdd gnd cell_6t
Xbit_r8_c251 bl[251] br[251] wl[8] vdd gnd cell_6t
Xbit_r9_c251 bl[251] br[251] wl[9] vdd gnd cell_6t
Xbit_r10_c251 bl[251] br[251] wl[10] vdd gnd cell_6t
Xbit_r11_c251 bl[251] br[251] wl[11] vdd gnd cell_6t
Xbit_r12_c251 bl[251] br[251] wl[12] vdd gnd cell_6t
Xbit_r13_c251 bl[251] br[251] wl[13] vdd gnd cell_6t
Xbit_r14_c251 bl[251] br[251] wl[14] vdd gnd cell_6t
Xbit_r15_c251 bl[251] br[251] wl[15] vdd gnd cell_6t
Xbit_r16_c251 bl[251] br[251] wl[16] vdd gnd cell_6t
Xbit_r17_c251 bl[251] br[251] wl[17] vdd gnd cell_6t
Xbit_r18_c251 bl[251] br[251] wl[18] vdd gnd cell_6t
Xbit_r19_c251 bl[251] br[251] wl[19] vdd gnd cell_6t
Xbit_r20_c251 bl[251] br[251] wl[20] vdd gnd cell_6t
Xbit_r21_c251 bl[251] br[251] wl[21] vdd gnd cell_6t
Xbit_r22_c251 bl[251] br[251] wl[22] vdd gnd cell_6t
Xbit_r23_c251 bl[251] br[251] wl[23] vdd gnd cell_6t
Xbit_r24_c251 bl[251] br[251] wl[24] vdd gnd cell_6t
Xbit_r25_c251 bl[251] br[251] wl[25] vdd gnd cell_6t
Xbit_r26_c251 bl[251] br[251] wl[26] vdd gnd cell_6t
Xbit_r27_c251 bl[251] br[251] wl[27] vdd gnd cell_6t
Xbit_r28_c251 bl[251] br[251] wl[28] vdd gnd cell_6t
Xbit_r29_c251 bl[251] br[251] wl[29] vdd gnd cell_6t
Xbit_r30_c251 bl[251] br[251] wl[30] vdd gnd cell_6t
Xbit_r31_c251 bl[251] br[251] wl[31] vdd gnd cell_6t
Xbit_r32_c251 bl[251] br[251] wl[32] vdd gnd cell_6t
Xbit_r33_c251 bl[251] br[251] wl[33] vdd gnd cell_6t
Xbit_r34_c251 bl[251] br[251] wl[34] vdd gnd cell_6t
Xbit_r35_c251 bl[251] br[251] wl[35] vdd gnd cell_6t
Xbit_r36_c251 bl[251] br[251] wl[36] vdd gnd cell_6t
Xbit_r37_c251 bl[251] br[251] wl[37] vdd gnd cell_6t
Xbit_r38_c251 bl[251] br[251] wl[38] vdd gnd cell_6t
Xbit_r39_c251 bl[251] br[251] wl[39] vdd gnd cell_6t
Xbit_r40_c251 bl[251] br[251] wl[40] vdd gnd cell_6t
Xbit_r41_c251 bl[251] br[251] wl[41] vdd gnd cell_6t
Xbit_r42_c251 bl[251] br[251] wl[42] vdd gnd cell_6t
Xbit_r43_c251 bl[251] br[251] wl[43] vdd gnd cell_6t
Xbit_r44_c251 bl[251] br[251] wl[44] vdd gnd cell_6t
Xbit_r45_c251 bl[251] br[251] wl[45] vdd gnd cell_6t
Xbit_r46_c251 bl[251] br[251] wl[46] vdd gnd cell_6t
Xbit_r47_c251 bl[251] br[251] wl[47] vdd gnd cell_6t
Xbit_r48_c251 bl[251] br[251] wl[48] vdd gnd cell_6t
Xbit_r49_c251 bl[251] br[251] wl[49] vdd gnd cell_6t
Xbit_r50_c251 bl[251] br[251] wl[50] vdd gnd cell_6t
Xbit_r51_c251 bl[251] br[251] wl[51] vdd gnd cell_6t
Xbit_r52_c251 bl[251] br[251] wl[52] vdd gnd cell_6t
Xbit_r53_c251 bl[251] br[251] wl[53] vdd gnd cell_6t
Xbit_r54_c251 bl[251] br[251] wl[54] vdd gnd cell_6t
Xbit_r55_c251 bl[251] br[251] wl[55] vdd gnd cell_6t
Xbit_r56_c251 bl[251] br[251] wl[56] vdd gnd cell_6t
Xbit_r57_c251 bl[251] br[251] wl[57] vdd gnd cell_6t
Xbit_r58_c251 bl[251] br[251] wl[58] vdd gnd cell_6t
Xbit_r59_c251 bl[251] br[251] wl[59] vdd gnd cell_6t
Xbit_r60_c251 bl[251] br[251] wl[60] vdd gnd cell_6t
Xbit_r61_c251 bl[251] br[251] wl[61] vdd gnd cell_6t
Xbit_r62_c251 bl[251] br[251] wl[62] vdd gnd cell_6t
Xbit_r63_c251 bl[251] br[251] wl[63] vdd gnd cell_6t
Xbit_r64_c251 bl[251] br[251] wl[64] vdd gnd cell_6t
Xbit_r65_c251 bl[251] br[251] wl[65] vdd gnd cell_6t
Xbit_r66_c251 bl[251] br[251] wl[66] vdd gnd cell_6t
Xbit_r67_c251 bl[251] br[251] wl[67] vdd gnd cell_6t
Xbit_r68_c251 bl[251] br[251] wl[68] vdd gnd cell_6t
Xbit_r69_c251 bl[251] br[251] wl[69] vdd gnd cell_6t
Xbit_r70_c251 bl[251] br[251] wl[70] vdd gnd cell_6t
Xbit_r71_c251 bl[251] br[251] wl[71] vdd gnd cell_6t
Xbit_r72_c251 bl[251] br[251] wl[72] vdd gnd cell_6t
Xbit_r73_c251 bl[251] br[251] wl[73] vdd gnd cell_6t
Xbit_r74_c251 bl[251] br[251] wl[74] vdd gnd cell_6t
Xbit_r75_c251 bl[251] br[251] wl[75] vdd gnd cell_6t
Xbit_r76_c251 bl[251] br[251] wl[76] vdd gnd cell_6t
Xbit_r77_c251 bl[251] br[251] wl[77] vdd gnd cell_6t
Xbit_r78_c251 bl[251] br[251] wl[78] vdd gnd cell_6t
Xbit_r79_c251 bl[251] br[251] wl[79] vdd gnd cell_6t
Xbit_r80_c251 bl[251] br[251] wl[80] vdd gnd cell_6t
Xbit_r81_c251 bl[251] br[251] wl[81] vdd gnd cell_6t
Xbit_r82_c251 bl[251] br[251] wl[82] vdd gnd cell_6t
Xbit_r83_c251 bl[251] br[251] wl[83] vdd gnd cell_6t
Xbit_r84_c251 bl[251] br[251] wl[84] vdd gnd cell_6t
Xbit_r85_c251 bl[251] br[251] wl[85] vdd gnd cell_6t
Xbit_r86_c251 bl[251] br[251] wl[86] vdd gnd cell_6t
Xbit_r87_c251 bl[251] br[251] wl[87] vdd gnd cell_6t
Xbit_r88_c251 bl[251] br[251] wl[88] vdd gnd cell_6t
Xbit_r89_c251 bl[251] br[251] wl[89] vdd gnd cell_6t
Xbit_r90_c251 bl[251] br[251] wl[90] vdd gnd cell_6t
Xbit_r91_c251 bl[251] br[251] wl[91] vdd gnd cell_6t
Xbit_r92_c251 bl[251] br[251] wl[92] vdd gnd cell_6t
Xbit_r93_c251 bl[251] br[251] wl[93] vdd gnd cell_6t
Xbit_r94_c251 bl[251] br[251] wl[94] vdd gnd cell_6t
Xbit_r95_c251 bl[251] br[251] wl[95] vdd gnd cell_6t
Xbit_r96_c251 bl[251] br[251] wl[96] vdd gnd cell_6t
Xbit_r97_c251 bl[251] br[251] wl[97] vdd gnd cell_6t
Xbit_r98_c251 bl[251] br[251] wl[98] vdd gnd cell_6t
Xbit_r99_c251 bl[251] br[251] wl[99] vdd gnd cell_6t
Xbit_r100_c251 bl[251] br[251] wl[100] vdd gnd cell_6t
Xbit_r101_c251 bl[251] br[251] wl[101] vdd gnd cell_6t
Xbit_r102_c251 bl[251] br[251] wl[102] vdd gnd cell_6t
Xbit_r103_c251 bl[251] br[251] wl[103] vdd gnd cell_6t
Xbit_r104_c251 bl[251] br[251] wl[104] vdd gnd cell_6t
Xbit_r105_c251 bl[251] br[251] wl[105] vdd gnd cell_6t
Xbit_r106_c251 bl[251] br[251] wl[106] vdd gnd cell_6t
Xbit_r107_c251 bl[251] br[251] wl[107] vdd gnd cell_6t
Xbit_r108_c251 bl[251] br[251] wl[108] vdd gnd cell_6t
Xbit_r109_c251 bl[251] br[251] wl[109] vdd gnd cell_6t
Xbit_r110_c251 bl[251] br[251] wl[110] vdd gnd cell_6t
Xbit_r111_c251 bl[251] br[251] wl[111] vdd gnd cell_6t
Xbit_r112_c251 bl[251] br[251] wl[112] vdd gnd cell_6t
Xbit_r113_c251 bl[251] br[251] wl[113] vdd gnd cell_6t
Xbit_r114_c251 bl[251] br[251] wl[114] vdd gnd cell_6t
Xbit_r115_c251 bl[251] br[251] wl[115] vdd gnd cell_6t
Xbit_r116_c251 bl[251] br[251] wl[116] vdd gnd cell_6t
Xbit_r117_c251 bl[251] br[251] wl[117] vdd gnd cell_6t
Xbit_r118_c251 bl[251] br[251] wl[118] vdd gnd cell_6t
Xbit_r119_c251 bl[251] br[251] wl[119] vdd gnd cell_6t
Xbit_r120_c251 bl[251] br[251] wl[120] vdd gnd cell_6t
Xbit_r121_c251 bl[251] br[251] wl[121] vdd gnd cell_6t
Xbit_r122_c251 bl[251] br[251] wl[122] vdd gnd cell_6t
Xbit_r123_c251 bl[251] br[251] wl[123] vdd gnd cell_6t
Xbit_r124_c251 bl[251] br[251] wl[124] vdd gnd cell_6t
Xbit_r125_c251 bl[251] br[251] wl[125] vdd gnd cell_6t
Xbit_r126_c251 bl[251] br[251] wl[126] vdd gnd cell_6t
Xbit_r127_c251 bl[251] br[251] wl[127] vdd gnd cell_6t
Xbit_r0_c252 bl[252] br[252] wl[0] vdd gnd cell_6t
Xbit_r1_c252 bl[252] br[252] wl[1] vdd gnd cell_6t
Xbit_r2_c252 bl[252] br[252] wl[2] vdd gnd cell_6t
Xbit_r3_c252 bl[252] br[252] wl[3] vdd gnd cell_6t
Xbit_r4_c252 bl[252] br[252] wl[4] vdd gnd cell_6t
Xbit_r5_c252 bl[252] br[252] wl[5] vdd gnd cell_6t
Xbit_r6_c252 bl[252] br[252] wl[6] vdd gnd cell_6t
Xbit_r7_c252 bl[252] br[252] wl[7] vdd gnd cell_6t
Xbit_r8_c252 bl[252] br[252] wl[8] vdd gnd cell_6t
Xbit_r9_c252 bl[252] br[252] wl[9] vdd gnd cell_6t
Xbit_r10_c252 bl[252] br[252] wl[10] vdd gnd cell_6t
Xbit_r11_c252 bl[252] br[252] wl[11] vdd gnd cell_6t
Xbit_r12_c252 bl[252] br[252] wl[12] vdd gnd cell_6t
Xbit_r13_c252 bl[252] br[252] wl[13] vdd gnd cell_6t
Xbit_r14_c252 bl[252] br[252] wl[14] vdd gnd cell_6t
Xbit_r15_c252 bl[252] br[252] wl[15] vdd gnd cell_6t
Xbit_r16_c252 bl[252] br[252] wl[16] vdd gnd cell_6t
Xbit_r17_c252 bl[252] br[252] wl[17] vdd gnd cell_6t
Xbit_r18_c252 bl[252] br[252] wl[18] vdd gnd cell_6t
Xbit_r19_c252 bl[252] br[252] wl[19] vdd gnd cell_6t
Xbit_r20_c252 bl[252] br[252] wl[20] vdd gnd cell_6t
Xbit_r21_c252 bl[252] br[252] wl[21] vdd gnd cell_6t
Xbit_r22_c252 bl[252] br[252] wl[22] vdd gnd cell_6t
Xbit_r23_c252 bl[252] br[252] wl[23] vdd gnd cell_6t
Xbit_r24_c252 bl[252] br[252] wl[24] vdd gnd cell_6t
Xbit_r25_c252 bl[252] br[252] wl[25] vdd gnd cell_6t
Xbit_r26_c252 bl[252] br[252] wl[26] vdd gnd cell_6t
Xbit_r27_c252 bl[252] br[252] wl[27] vdd gnd cell_6t
Xbit_r28_c252 bl[252] br[252] wl[28] vdd gnd cell_6t
Xbit_r29_c252 bl[252] br[252] wl[29] vdd gnd cell_6t
Xbit_r30_c252 bl[252] br[252] wl[30] vdd gnd cell_6t
Xbit_r31_c252 bl[252] br[252] wl[31] vdd gnd cell_6t
Xbit_r32_c252 bl[252] br[252] wl[32] vdd gnd cell_6t
Xbit_r33_c252 bl[252] br[252] wl[33] vdd gnd cell_6t
Xbit_r34_c252 bl[252] br[252] wl[34] vdd gnd cell_6t
Xbit_r35_c252 bl[252] br[252] wl[35] vdd gnd cell_6t
Xbit_r36_c252 bl[252] br[252] wl[36] vdd gnd cell_6t
Xbit_r37_c252 bl[252] br[252] wl[37] vdd gnd cell_6t
Xbit_r38_c252 bl[252] br[252] wl[38] vdd gnd cell_6t
Xbit_r39_c252 bl[252] br[252] wl[39] vdd gnd cell_6t
Xbit_r40_c252 bl[252] br[252] wl[40] vdd gnd cell_6t
Xbit_r41_c252 bl[252] br[252] wl[41] vdd gnd cell_6t
Xbit_r42_c252 bl[252] br[252] wl[42] vdd gnd cell_6t
Xbit_r43_c252 bl[252] br[252] wl[43] vdd gnd cell_6t
Xbit_r44_c252 bl[252] br[252] wl[44] vdd gnd cell_6t
Xbit_r45_c252 bl[252] br[252] wl[45] vdd gnd cell_6t
Xbit_r46_c252 bl[252] br[252] wl[46] vdd gnd cell_6t
Xbit_r47_c252 bl[252] br[252] wl[47] vdd gnd cell_6t
Xbit_r48_c252 bl[252] br[252] wl[48] vdd gnd cell_6t
Xbit_r49_c252 bl[252] br[252] wl[49] vdd gnd cell_6t
Xbit_r50_c252 bl[252] br[252] wl[50] vdd gnd cell_6t
Xbit_r51_c252 bl[252] br[252] wl[51] vdd gnd cell_6t
Xbit_r52_c252 bl[252] br[252] wl[52] vdd gnd cell_6t
Xbit_r53_c252 bl[252] br[252] wl[53] vdd gnd cell_6t
Xbit_r54_c252 bl[252] br[252] wl[54] vdd gnd cell_6t
Xbit_r55_c252 bl[252] br[252] wl[55] vdd gnd cell_6t
Xbit_r56_c252 bl[252] br[252] wl[56] vdd gnd cell_6t
Xbit_r57_c252 bl[252] br[252] wl[57] vdd gnd cell_6t
Xbit_r58_c252 bl[252] br[252] wl[58] vdd gnd cell_6t
Xbit_r59_c252 bl[252] br[252] wl[59] vdd gnd cell_6t
Xbit_r60_c252 bl[252] br[252] wl[60] vdd gnd cell_6t
Xbit_r61_c252 bl[252] br[252] wl[61] vdd gnd cell_6t
Xbit_r62_c252 bl[252] br[252] wl[62] vdd gnd cell_6t
Xbit_r63_c252 bl[252] br[252] wl[63] vdd gnd cell_6t
Xbit_r64_c252 bl[252] br[252] wl[64] vdd gnd cell_6t
Xbit_r65_c252 bl[252] br[252] wl[65] vdd gnd cell_6t
Xbit_r66_c252 bl[252] br[252] wl[66] vdd gnd cell_6t
Xbit_r67_c252 bl[252] br[252] wl[67] vdd gnd cell_6t
Xbit_r68_c252 bl[252] br[252] wl[68] vdd gnd cell_6t
Xbit_r69_c252 bl[252] br[252] wl[69] vdd gnd cell_6t
Xbit_r70_c252 bl[252] br[252] wl[70] vdd gnd cell_6t
Xbit_r71_c252 bl[252] br[252] wl[71] vdd gnd cell_6t
Xbit_r72_c252 bl[252] br[252] wl[72] vdd gnd cell_6t
Xbit_r73_c252 bl[252] br[252] wl[73] vdd gnd cell_6t
Xbit_r74_c252 bl[252] br[252] wl[74] vdd gnd cell_6t
Xbit_r75_c252 bl[252] br[252] wl[75] vdd gnd cell_6t
Xbit_r76_c252 bl[252] br[252] wl[76] vdd gnd cell_6t
Xbit_r77_c252 bl[252] br[252] wl[77] vdd gnd cell_6t
Xbit_r78_c252 bl[252] br[252] wl[78] vdd gnd cell_6t
Xbit_r79_c252 bl[252] br[252] wl[79] vdd gnd cell_6t
Xbit_r80_c252 bl[252] br[252] wl[80] vdd gnd cell_6t
Xbit_r81_c252 bl[252] br[252] wl[81] vdd gnd cell_6t
Xbit_r82_c252 bl[252] br[252] wl[82] vdd gnd cell_6t
Xbit_r83_c252 bl[252] br[252] wl[83] vdd gnd cell_6t
Xbit_r84_c252 bl[252] br[252] wl[84] vdd gnd cell_6t
Xbit_r85_c252 bl[252] br[252] wl[85] vdd gnd cell_6t
Xbit_r86_c252 bl[252] br[252] wl[86] vdd gnd cell_6t
Xbit_r87_c252 bl[252] br[252] wl[87] vdd gnd cell_6t
Xbit_r88_c252 bl[252] br[252] wl[88] vdd gnd cell_6t
Xbit_r89_c252 bl[252] br[252] wl[89] vdd gnd cell_6t
Xbit_r90_c252 bl[252] br[252] wl[90] vdd gnd cell_6t
Xbit_r91_c252 bl[252] br[252] wl[91] vdd gnd cell_6t
Xbit_r92_c252 bl[252] br[252] wl[92] vdd gnd cell_6t
Xbit_r93_c252 bl[252] br[252] wl[93] vdd gnd cell_6t
Xbit_r94_c252 bl[252] br[252] wl[94] vdd gnd cell_6t
Xbit_r95_c252 bl[252] br[252] wl[95] vdd gnd cell_6t
Xbit_r96_c252 bl[252] br[252] wl[96] vdd gnd cell_6t
Xbit_r97_c252 bl[252] br[252] wl[97] vdd gnd cell_6t
Xbit_r98_c252 bl[252] br[252] wl[98] vdd gnd cell_6t
Xbit_r99_c252 bl[252] br[252] wl[99] vdd gnd cell_6t
Xbit_r100_c252 bl[252] br[252] wl[100] vdd gnd cell_6t
Xbit_r101_c252 bl[252] br[252] wl[101] vdd gnd cell_6t
Xbit_r102_c252 bl[252] br[252] wl[102] vdd gnd cell_6t
Xbit_r103_c252 bl[252] br[252] wl[103] vdd gnd cell_6t
Xbit_r104_c252 bl[252] br[252] wl[104] vdd gnd cell_6t
Xbit_r105_c252 bl[252] br[252] wl[105] vdd gnd cell_6t
Xbit_r106_c252 bl[252] br[252] wl[106] vdd gnd cell_6t
Xbit_r107_c252 bl[252] br[252] wl[107] vdd gnd cell_6t
Xbit_r108_c252 bl[252] br[252] wl[108] vdd gnd cell_6t
Xbit_r109_c252 bl[252] br[252] wl[109] vdd gnd cell_6t
Xbit_r110_c252 bl[252] br[252] wl[110] vdd gnd cell_6t
Xbit_r111_c252 bl[252] br[252] wl[111] vdd gnd cell_6t
Xbit_r112_c252 bl[252] br[252] wl[112] vdd gnd cell_6t
Xbit_r113_c252 bl[252] br[252] wl[113] vdd gnd cell_6t
Xbit_r114_c252 bl[252] br[252] wl[114] vdd gnd cell_6t
Xbit_r115_c252 bl[252] br[252] wl[115] vdd gnd cell_6t
Xbit_r116_c252 bl[252] br[252] wl[116] vdd gnd cell_6t
Xbit_r117_c252 bl[252] br[252] wl[117] vdd gnd cell_6t
Xbit_r118_c252 bl[252] br[252] wl[118] vdd gnd cell_6t
Xbit_r119_c252 bl[252] br[252] wl[119] vdd gnd cell_6t
Xbit_r120_c252 bl[252] br[252] wl[120] vdd gnd cell_6t
Xbit_r121_c252 bl[252] br[252] wl[121] vdd gnd cell_6t
Xbit_r122_c252 bl[252] br[252] wl[122] vdd gnd cell_6t
Xbit_r123_c252 bl[252] br[252] wl[123] vdd gnd cell_6t
Xbit_r124_c252 bl[252] br[252] wl[124] vdd gnd cell_6t
Xbit_r125_c252 bl[252] br[252] wl[125] vdd gnd cell_6t
Xbit_r126_c252 bl[252] br[252] wl[126] vdd gnd cell_6t
Xbit_r127_c252 bl[252] br[252] wl[127] vdd gnd cell_6t
Xbit_r0_c253 bl[253] br[253] wl[0] vdd gnd cell_6t
Xbit_r1_c253 bl[253] br[253] wl[1] vdd gnd cell_6t
Xbit_r2_c253 bl[253] br[253] wl[2] vdd gnd cell_6t
Xbit_r3_c253 bl[253] br[253] wl[3] vdd gnd cell_6t
Xbit_r4_c253 bl[253] br[253] wl[4] vdd gnd cell_6t
Xbit_r5_c253 bl[253] br[253] wl[5] vdd gnd cell_6t
Xbit_r6_c253 bl[253] br[253] wl[6] vdd gnd cell_6t
Xbit_r7_c253 bl[253] br[253] wl[7] vdd gnd cell_6t
Xbit_r8_c253 bl[253] br[253] wl[8] vdd gnd cell_6t
Xbit_r9_c253 bl[253] br[253] wl[9] vdd gnd cell_6t
Xbit_r10_c253 bl[253] br[253] wl[10] vdd gnd cell_6t
Xbit_r11_c253 bl[253] br[253] wl[11] vdd gnd cell_6t
Xbit_r12_c253 bl[253] br[253] wl[12] vdd gnd cell_6t
Xbit_r13_c253 bl[253] br[253] wl[13] vdd gnd cell_6t
Xbit_r14_c253 bl[253] br[253] wl[14] vdd gnd cell_6t
Xbit_r15_c253 bl[253] br[253] wl[15] vdd gnd cell_6t
Xbit_r16_c253 bl[253] br[253] wl[16] vdd gnd cell_6t
Xbit_r17_c253 bl[253] br[253] wl[17] vdd gnd cell_6t
Xbit_r18_c253 bl[253] br[253] wl[18] vdd gnd cell_6t
Xbit_r19_c253 bl[253] br[253] wl[19] vdd gnd cell_6t
Xbit_r20_c253 bl[253] br[253] wl[20] vdd gnd cell_6t
Xbit_r21_c253 bl[253] br[253] wl[21] vdd gnd cell_6t
Xbit_r22_c253 bl[253] br[253] wl[22] vdd gnd cell_6t
Xbit_r23_c253 bl[253] br[253] wl[23] vdd gnd cell_6t
Xbit_r24_c253 bl[253] br[253] wl[24] vdd gnd cell_6t
Xbit_r25_c253 bl[253] br[253] wl[25] vdd gnd cell_6t
Xbit_r26_c253 bl[253] br[253] wl[26] vdd gnd cell_6t
Xbit_r27_c253 bl[253] br[253] wl[27] vdd gnd cell_6t
Xbit_r28_c253 bl[253] br[253] wl[28] vdd gnd cell_6t
Xbit_r29_c253 bl[253] br[253] wl[29] vdd gnd cell_6t
Xbit_r30_c253 bl[253] br[253] wl[30] vdd gnd cell_6t
Xbit_r31_c253 bl[253] br[253] wl[31] vdd gnd cell_6t
Xbit_r32_c253 bl[253] br[253] wl[32] vdd gnd cell_6t
Xbit_r33_c253 bl[253] br[253] wl[33] vdd gnd cell_6t
Xbit_r34_c253 bl[253] br[253] wl[34] vdd gnd cell_6t
Xbit_r35_c253 bl[253] br[253] wl[35] vdd gnd cell_6t
Xbit_r36_c253 bl[253] br[253] wl[36] vdd gnd cell_6t
Xbit_r37_c253 bl[253] br[253] wl[37] vdd gnd cell_6t
Xbit_r38_c253 bl[253] br[253] wl[38] vdd gnd cell_6t
Xbit_r39_c253 bl[253] br[253] wl[39] vdd gnd cell_6t
Xbit_r40_c253 bl[253] br[253] wl[40] vdd gnd cell_6t
Xbit_r41_c253 bl[253] br[253] wl[41] vdd gnd cell_6t
Xbit_r42_c253 bl[253] br[253] wl[42] vdd gnd cell_6t
Xbit_r43_c253 bl[253] br[253] wl[43] vdd gnd cell_6t
Xbit_r44_c253 bl[253] br[253] wl[44] vdd gnd cell_6t
Xbit_r45_c253 bl[253] br[253] wl[45] vdd gnd cell_6t
Xbit_r46_c253 bl[253] br[253] wl[46] vdd gnd cell_6t
Xbit_r47_c253 bl[253] br[253] wl[47] vdd gnd cell_6t
Xbit_r48_c253 bl[253] br[253] wl[48] vdd gnd cell_6t
Xbit_r49_c253 bl[253] br[253] wl[49] vdd gnd cell_6t
Xbit_r50_c253 bl[253] br[253] wl[50] vdd gnd cell_6t
Xbit_r51_c253 bl[253] br[253] wl[51] vdd gnd cell_6t
Xbit_r52_c253 bl[253] br[253] wl[52] vdd gnd cell_6t
Xbit_r53_c253 bl[253] br[253] wl[53] vdd gnd cell_6t
Xbit_r54_c253 bl[253] br[253] wl[54] vdd gnd cell_6t
Xbit_r55_c253 bl[253] br[253] wl[55] vdd gnd cell_6t
Xbit_r56_c253 bl[253] br[253] wl[56] vdd gnd cell_6t
Xbit_r57_c253 bl[253] br[253] wl[57] vdd gnd cell_6t
Xbit_r58_c253 bl[253] br[253] wl[58] vdd gnd cell_6t
Xbit_r59_c253 bl[253] br[253] wl[59] vdd gnd cell_6t
Xbit_r60_c253 bl[253] br[253] wl[60] vdd gnd cell_6t
Xbit_r61_c253 bl[253] br[253] wl[61] vdd gnd cell_6t
Xbit_r62_c253 bl[253] br[253] wl[62] vdd gnd cell_6t
Xbit_r63_c253 bl[253] br[253] wl[63] vdd gnd cell_6t
Xbit_r64_c253 bl[253] br[253] wl[64] vdd gnd cell_6t
Xbit_r65_c253 bl[253] br[253] wl[65] vdd gnd cell_6t
Xbit_r66_c253 bl[253] br[253] wl[66] vdd gnd cell_6t
Xbit_r67_c253 bl[253] br[253] wl[67] vdd gnd cell_6t
Xbit_r68_c253 bl[253] br[253] wl[68] vdd gnd cell_6t
Xbit_r69_c253 bl[253] br[253] wl[69] vdd gnd cell_6t
Xbit_r70_c253 bl[253] br[253] wl[70] vdd gnd cell_6t
Xbit_r71_c253 bl[253] br[253] wl[71] vdd gnd cell_6t
Xbit_r72_c253 bl[253] br[253] wl[72] vdd gnd cell_6t
Xbit_r73_c253 bl[253] br[253] wl[73] vdd gnd cell_6t
Xbit_r74_c253 bl[253] br[253] wl[74] vdd gnd cell_6t
Xbit_r75_c253 bl[253] br[253] wl[75] vdd gnd cell_6t
Xbit_r76_c253 bl[253] br[253] wl[76] vdd gnd cell_6t
Xbit_r77_c253 bl[253] br[253] wl[77] vdd gnd cell_6t
Xbit_r78_c253 bl[253] br[253] wl[78] vdd gnd cell_6t
Xbit_r79_c253 bl[253] br[253] wl[79] vdd gnd cell_6t
Xbit_r80_c253 bl[253] br[253] wl[80] vdd gnd cell_6t
Xbit_r81_c253 bl[253] br[253] wl[81] vdd gnd cell_6t
Xbit_r82_c253 bl[253] br[253] wl[82] vdd gnd cell_6t
Xbit_r83_c253 bl[253] br[253] wl[83] vdd gnd cell_6t
Xbit_r84_c253 bl[253] br[253] wl[84] vdd gnd cell_6t
Xbit_r85_c253 bl[253] br[253] wl[85] vdd gnd cell_6t
Xbit_r86_c253 bl[253] br[253] wl[86] vdd gnd cell_6t
Xbit_r87_c253 bl[253] br[253] wl[87] vdd gnd cell_6t
Xbit_r88_c253 bl[253] br[253] wl[88] vdd gnd cell_6t
Xbit_r89_c253 bl[253] br[253] wl[89] vdd gnd cell_6t
Xbit_r90_c253 bl[253] br[253] wl[90] vdd gnd cell_6t
Xbit_r91_c253 bl[253] br[253] wl[91] vdd gnd cell_6t
Xbit_r92_c253 bl[253] br[253] wl[92] vdd gnd cell_6t
Xbit_r93_c253 bl[253] br[253] wl[93] vdd gnd cell_6t
Xbit_r94_c253 bl[253] br[253] wl[94] vdd gnd cell_6t
Xbit_r95_c253 bl[253] br[253] wl[95] vdd gnd cell_6t
Xbit_r96_c253 bl[253] br[253] wl[96] vdd gnd cell_6t
Xbit_r97_c253 bl[253] br[253] wl[97] vdd gnd cell_6t
Xbit_r98_c253 bl[253] br[253] wl[98] vdd gnd cell_6t
Xbit_r99_c253 bl[253] br[253] wl[99] vdd gnd cell_6t
Xbit_r100_c253 bl[253] br[253] wl[100] vdd gnd cell_6t
Xbit_r101_c253 bl[253] br[253] wl[101] vdd gnd cell_6t
Xbit_r102_c253 bl[253] br[253] wl[102] vdd gnd cell_6t
Xbit_r103_c253 bl[253] br[253] wl[103] vdd gnd cell_6t
Xbit_r104_c253 bl[253] br[253] wl[104] vdd gnd cell_6t
Xbit_r105_c253 bl[253] br[253] wl[105] vdd gnd cell_6t
Xbit_r106_c253 bl[253] br[253] wl[106] vdd gnd cell_6t
Xbit_r107_c253 bl[253] br[253] wl[107] vdd gnd cell_6t
Xbit_r108_c253 bl[253] br[253] wl[108] vdd gnd cell_6t
Xbit_r109_c253 bl[253] br[253] wl[109] vdd gnd cell_6t
Xbit_r110_c253 bl[253] br[253] wl[110] vdd gnd cell_6t
Xbit_r111_c253 bl[253] br[253] wl[111] vdd gnd cell_6t
Xbit_r112_c253 bl[253] br[253] wl[112] vdd gnd cell_6t
Xbit_r113_c253 bl[253] br[253] wl[113] vdd gnd cell_6t
Xbit_r114_c253 bl[253] br[253] wl[114] vdd gnd cell_6t
Xbit_r115_c253 bl[253] br[253] wl[115] vdd gnd cell_6t
Xbit_r116_c253 bl[253] br[253] wl[116] vdd gnd cell_6t
Xbit_r117_c253 bl[253] br[253] wl[117] vdd gnd cell_6t
Xbit_r118_c253 bl[253] br[253] wl[118] vdd gnd cell_6t
Xbit_r119_c253 bl[253] br[253] wl[119] vdd gnd cell_6t
Xbit_r120_c253 bl[253] br[253] wl[120] vdd gnd cell_6t
Xbit_r121_c253 bl[253] br[253] wl[121] vdd gnd cell_6t
Xbit_r122_c253 bl[253] br[253] wl[122] vdd gnd cell_6t
Xbit_r123_c253 bl[253] br[253] wl[123] vdd gnd cell_6t
Xbit_r124_c253 bl[253] br[253] wl[124] vdd gnd cell_6t
Xbit_r125_c253 bl[253] br[253] wl[125] vdd gnd cell_6t
Xbit_r126_c253 bl[253] br[253] wl[126] vdd gnd cell_6t
Xbit_r127_c253 bl[253] br[253] wl[127] vdd gnd cell_6t
Xbit_r0_c254 bl[254] br[254] wl[0] vdd gnd cell_6t
Xbit_r1_c254 bl[254] br[254] wl[1] vdd gnd cell_6t
Xbit_r2_c254 bl[254] br[254] wl[2] vdd gnd cell_6t
Xbit_r3_c254 bl[254] br[254] wl[3] vdd gnd cell_6t
Xbit_r4_c254 bl[254] br[254] wl[4] vdd gnd cell_6t
Xbit_r5_c254 bl[254] br[254] wl[5] vdd gnd cell_6t
Xbit_r6_c254 bl[254] br[254] wl[6] vdd gnd cell_6t
Xbit_r7_c254 bl[254] br[254] wl[7] vdd gnd cell_6t
Xbit_r8_c254 bl[254] br[254] wl[8] vdd gnd cell_6t
Xbit_r9_c254 bl[254] br[254] wl[9] vdd gnd cell_6t
Xbit_r10_c254 bl[254] br[254] wl[10] vdd gnd cell_6t
Xbit_r11_c254 bl[254] br[254] wl[11] vdd gnd cell_6t
Xbit_r12_c254 bl[254] br[254] wl[12] vdd gnd cell_6t
Xbit_r13_c254 bl[254] br[254] wl[13] vdd gnd cell_6t
Xbit_r14_c254 bl[254] br[254] wl[14] vdd gnd cell_6t
Xbit_r15_c254 bl[254] br[254] wl[15] vdd gnd cell_6t
Xbit_r16_c254 bl[254] br[254] wl[16] vdd gnd cell_6t
Xbit_r17_c254 bl[254] br[254] wl[17] vdd gnd cell_6t
Xbit_r18_c254 bl[254] br[254] wl[18] vdd gnd cell_6t
Xbit_r19_c254 bl[254] br[254] wl[19] vdd gnd cell_6t
Xbit_r20_c254 bl[254] br[254] wl[20] vdd gnd cell_6t
Xbit_r21_c254 bl[254] br[254] wl[21] vdd gnd cell_6t
Xbit_r22_c254 bl[254] br[254] wl[22] vdd gnd cell_6t
Xbit_r23_c254 bl[254] br[254] wl[23] vdd gnd cell_6t
Xbit_r24_c254 bl[254] br[254] wl[24] vdd gnd cell_6t
Xbit_r25_c254 bl[254] br[254] wl[25] vdd gnd cell_6t
Xbit_r26_c254 bl[254] br[254] wl[26] vdd gnd cell_6t
Xbit_r27_c254 bl[254] br[254] wl[27] vdd gnd cell_6t
Xbit_r28_c254 bl[254] br[254] wl[28] vdd gnd cell_6t
Xbit_r29_c254 bl[254] br[254] wl[29] vdd gnd cell_6t
Xbit_r30_c254 bl[254] br[254] wl[30] vdd gnd cell_6t
Xbit_r31_c254 bl[254] br[254] wl[31] vdd gnd cell_6t
Xbit_r32_c254 bl[254] br[254] wl[32] vdd gnd cell_6t
Xbit_r33_c254 bl[254] br[254] wl[33] vdd gnd cell_6t
Xbit_r34_c254 bl[254] br[254] wl[34] vdd gnd cell_6t
Xbit_r35_c254 bl[254] br[254] wl[35] vdd gnd cell_6t
Xbit_r36_c254 bl[254] br[254] wl[36] vdd gnd cell_6t
Xbit_r37_c254 bl[254] br[254] wl[37] vdd gnd cell_6t
Xbit_r38_c254 bl[254] br[254] wl[38] vdd gnd cell_6t
Xbit_r39_c254 bl[254] br[254] wl[39] vdd gnd cell_6t
Xbit_r40_c254 bl[254] br[254] wl[40] vdd gnd cell_6t
Xbit_r41_c254 bl[254] br[254] wl[41] vdd gnd cell_6t
Xbit_r42_c254 bl[254] br[254] wl[42] vdd gnd cell_6t
Xbit_r43_c254 bl[254] br[254] wl[43] vdd gnd cell_6t
Xbit_r44_c254 bl[254] br[254] wl[44] vdd gnd cell_6t
Xbit_r45_c254 bl[254] br[254] wl[45] vdd gnd cell_6t
Xbit_r46_c254 bl[254] br[254] wl[46] vdd gnd cell_6t
Xbit_r47_c254 bl[254] br[254] wl[47] vdd gnd cell_6t
Xbit_r48_c254 bl[254] br[254] wl[48] vdd gnd cell_6t
Xbit_r49_c254 bl[254] br[254] wl[49] vdd gnd cell_6t
Xbit_r50_c254 bl[254] br[254] wl[50] vdd gnd cell_6t
Xbit_r51_c254 bl[254] br[254] wl[51] vdd gnd cell_6t
Xbit_r52_c254 bl[254] br[254] wl[52] vdd gnd cell_6t
Xbit_r53_c254 bl[254] br[254] wl[53] vdd gnd cell_6t
Xbit_r54_c254 bl[254] br[254] wl[54] vdd gnd cell_6t
Xbit_r55_c254 bl[254] br[254] wl[55] vdd gnd cell_6t
Xbit_r56_c254 bl[254] br[254] wl[56] vdd gnd cell_6t
Xbit_r57_c254 bl[254] br[254] wl[57] vdd gnd cell_6t
Xbit_r58_c254 bl[254] br[254] wl[58] vdd gnd cell_6t
Xbit_r59_c254 bl[254] br[254] wl[59] vdd gnd cell_6t
Xbit_r60_c254 bl[254] br[254] wl[60] vdd gnd cell_6t
Xbit_r61_c254 bl[254] br[254] wl[61] vdd gnd cell_6t
Xbit_r62_c254 bl[254] br[254] wl[62] vdd gnd cell_6t
Xbit_r63_c254 bl[254] br[254] wl[63] vdd gnd cell_6t
Xbit_r64_c254 bl[254] br[254] wl[64] vdd gnd cell_6t
Xbit_r65_c254 bl[254] br[254] wl[65] vdd gnd cell_6t
Xbit_r66_c254 bl[254] br[254] wl[66] vdd gnd cell_6t
Xbit_r67_c254 bl[254] br[254] wl[67] vdd gnd cell_6t
Xbit_r68_c254 bl[254] br[254] wl[68] vdd gnd cell_6t
Xbit_r69_c254 bl[254] br[254] wl[69] vdd gnd cell_6t
Xbit_r70_c254 bl[254] br[254] wl[70] vdd gnd cell_6t
Xbit_r71_c254 bl[254] br[254] wl[71] vdd gnd cell_6t
Xbit_r72_c254 bl[254] br[254] wl[72] vdd gnd cell_6t
Xbit_r73_c254 bl[254] br[254] wl[73] vdd gnd cell_6t
Xbit_r74_c254 bl[254] br[254] wl[74] vdd gnd cell_6t
Xbit_r75_c254 bl[254] br[254] wl[75] vdd gnd cell_6t
Xbit_r76_c254 bl[254] br[254] wl[76] vdd gnd cell_6t
Xbit_r77_c254 bl[254] br[254] wl[77] vdd gnd cell_6t
Xbit_r78_c254 bl[254] br[254] wl[78] vdd gnd cell_6t
Xbit_r79_c254 bl[254] br[254] wl[79] vdd gnd cell_6t
Xbit_r80_c254 bl[254] br[254] wl[80] vdd gnd cell_6t
Xbit_r81_c254 bl[254] br[254] wl[81] vdd gnd cell_6t
Xbit_r82_c254 bl[254] br[254] wl[82] vdd gnd cell_6t
Xbit_r83_c254 bl[254] br[254] wl[83] vdd gnd cell_6t
Xbit_r84_c254 bl[254] br[254] wl[84] vdd gnd cell_6t
Xbit_r85_c254 bl[254] br[254] wl[85] vdd gnd cell_6t
Xbit_r86_c254 bl[254] br[254] wl[86] vdd gnd cell_6t
Xbit_r87_c254 bl[254] br[254] wl[87] vdd gnd cell_6t
Xbit_r88_c254 bl[254] br[254] wl[88] vdd gnd cell_6t
Xbit_r89_c254 bl[254] br[254] wl[89] vdd gnd cell_6t
Xbit_r90_c254 bl[254] br[254] wl[90] vdd gnd cell_6t
Xbit_r91_c254 bl[254] br[254] wl[91] vdd gnd cell_6t
Xbit_r92_c254 bl[254] br[254] wl[92] vdd gnd cell_6t
Xbit_r93_c254 bl[254] br[254] wl[93] vdd gnd cell_6t
Xbit_r94_c254 bl[254] br[254] wl[94] vdd gnd cell_6t
Xbit_r95_c254 bl[254] br[254] wl[95] vdd gnd cell_6t
Xbit_r96_c254 bl[254] br[254] wl[96] vdd gnd cell_6t
Xbit_r97_c254 bl[254] br[254] wl[97] vdd gnd cell_6t
Xbit_r98_c254 bl[254] br[254] wl[98] vdd gnd cell_6t
Xbit_r99_c254 bl[254] br[254] wl[99] vdd gnd cell_6t
Xbit_r100_c254 bl[254] br[254] wl[100] vdd gnd cell_6t
Xbit_r101_c254 bl[254] br[254] wl[101] vdd gnd cell_6t
Xbit_r102_c254 bl[254] br[254] wl[102] vdd gnd cell_6t
Xbit_r103_c254 bl[254] br[254] wl[103] vdd gnd cell_6t
Xbit_r104_c254 bl[254] br[254] wl[104] vdd gnd cell_6t
Xbit_r105_c254 bl[254] br[254] wl[105] vdd gnd cell_6t
Xbit_r106_c254 bl[254] br[254] wl[106] vdd gnd cell_6t
Xbit_r107_c254 bl[254] br[254] wl[107] vdd gnd cell_6t
Xbit_r108_c254 bl[254] br[254] wl[108] vdd gnd cell_6t
Xbit_r109_c254 bl[254] br[254] wl[109] vdd gnd cell_6t
Xbit_r110_c254 bl[254] br[254] wl[110] vdd gnd cell_6t
Xbit_r111_c254 bl[254] br[254] wl[111] vdd gnd cell_6t
Xbit_r112_c254 bl[254] br[254] wl[112] vdd gnd cell_6t
Xbit_r113_c254 bl[254] br[254] wl[113] vdd gnd cell_6t
Xbit_r114_c254 bl[254] br[254] wl[114] vdd gnd cell_6t
Xbit_r115_c254 bl[254] br[254] wl[115] vdd gnd cell_6t
Xbit_r116_c254 bl[254] br[254] wl[116] vdd gnd cell_6t
Xbit_r117_c254 bl[254] br[254] wl[117] vdd gnd cell_6t
Xbit_r118_c254 bl[254] br[254] wl[118] vdd gnd cell_6t
Xbit_r119_c254 bl[254] br[254] wl[119] vdd gnd cell_6t
Xbit_r120_c254 bl[254] br[254] wl[120] vdd gnd cell_6t
Xbit_r121_c254 bl[254] br[254] wl[121] vdd gnd cell_6t
Xbit_r122_c254 bl[254] br[254] wl[122] vdd gnd cell_6t
Xbit_r123_c254 bl[254] br[254] wl[123] vdd gnd cell_6t
Xbit_r124_c254 bl[254] br[254] wl[124] vdd gnd cell_6t
Xbit_r125_c254 bl[254] br[254] wl[125] vdd gnd cell_6t
Xbit_r126_c254 bl[254] br[254] wl[126] vdd gnd cell_6t
Xbit_r127_c254 bl[254] br[254] wl[127] vdd gnd cell_6t
Xbit_r0_c255 bl[255] br[255] wl[0] vdd gnd cell_6t
Xbit_r1_c255 bl[255] br[255] wl[1] vdd gnd cell_6t
Xbit_r2_c255 bl[255] br[255] wl[2] vdd gnd cell_6t
Xbit_r3_c255 bl[255] br[255] wl[3] vdd gnd cell_6t
Xbit_r4_c255 bl[255] br[255] wl[4] vdd gnd cell_6t
Xbit_r5_c255 bl[255] br[255] wl[5] vdd gnd cell_6t
Xbit_r6_c255 bl[255] br[255] wl[6] vdd gnd cell_6t
Xbit_r7_c255 bl[255] br[255] wl[7] vdd gnd cell_6t
Xbit_r8_c255 bl[255] br[255] wl[8] vdd gnd cell_6t
Xbit_r9_c255 bl[255] br[255] wl[9] vdd gnd cell_6t
Xbit_r10_c255 bl[255] br[255] wl[10] vdd gnd cell_6t
Xbit_r11_c255 bl[255] br[255] wl[11] vdd gnd cell_6t
Xbit_r12_c255 bl[255] br[255] wl[12] vdd gnd cell_6t
Xbit_r13_c255 bl[255] br[255] wl[13] vdd gnd cell_6t
Xbit_r14_c255 bl[255] br[255] wl[14] vdd gnd cell_6t
Xbit_r15_c255 bl[255] br[255] wl[15] vdd gnd cell_6t
Xbit_r16_c255 bl[255] br[255] wl[16] vdd gnd cell_6t
Xbit_r17_c255 bl[255] br[255] wl[17] vdd gnd cell_6t
Xbit_r18_c255 bl[255] br[255] wl[18] vdd gnd cell_6t
Xbit_r19_c255 bl[255] br[255] wl[19] vdd gnd cell_6t
Xbit_r20_c255 bl[255] br[255] wl[20] vdd gnd cell_6t
Xbit_r21_c255 bl[255] br[255] wl[21] vdd gnd cell_6t
Xbit_r22_c255 bl[255] br[255] wl[22] vdd gnd cell_6t
Xbit_r23_c255 bl[255] br[255] wl[23] vdd gnd cell_6t
Xbit_r24_c255 bl[255] br[255] wl[24] vdd gnd cell_6t
Xbit_r25_c255 bl[255] br[255] wl[25] vdd gnd cell_6t
Xbit_r26_c255 bl[255] br[255] wl[26] vdd gnd cell_6t
Xbit_r27_c255 bl[255] br[255] wl[27] vdd gnd cell_6t
Xbit_r28_c255 bl[255] br[255] wl[28] vdd gnd cell_6t
Xbit_r29_c255 bl[255] br[255] wl[29] vdd gnd cell_6t
Xbit_r30_c255 bl[255] br[255] wl[30] vdd gnd cell_6t
Xbit_r31_c255 bl[255] br[255] wl[31] vdd gnd cell_6t
Xbit_r32_c255 bl[255] br[255] wl[32] vdd gnd cell_6t
Xbit_r33_c255 bl[255] br[255] wl[33] vdd gnd cell_6t
Xbit_r34_c255 bl[255] br[255] wl[34] vdd gnd cell_6t
Xbit_r35_c255 bl[255] br[255] wl[35] vdd gnd cell_6t
Xbit_r36_c255 bl[255] br[255] wl[36] vdd gnd cell_6t
Xbit_r37_c255 bl[255] br[255] wl[37] vdd gnd cell_6t
Xbit_r38_c255 bl[255] br[255] wl[38] vdd gnd cell_6t
Xbit_r39_c255 bl[255] br[255] wl[39] vdd gnd cell_6t
Xbit_r40_c255 bl[255] br[255] wl[40] vdd gnd cell_6t
Xbit_r41_c255 bl[255] br[255] wl[41] vdd gnd cell_6t
Xbit_r42_c255 bl[255] br[255] wl[42] vdd gnd cell_6t
Xbit_r43_c255 bl[255] br[255] wl[43] vdd gnd cell_6t
Xbit_r44_c255 bl[255] br[255] wl[44] vdd gnd cell_6t
Xbit_r45_c255 bl[255] br[255] wl[45] vdd gnd cell_6t
Xbit_r46_c255 bl[255] br[255] wl[46] vdd gnd cell_6t
Xbit_r47_c255 bl[255] br[255] wl[47] vdd gnd cell_6t
Xbit_r48_c255 bl[255] br[255] wl[48] vdd gnd cell_6t
Xbit_r49_c255 bl[255] br[255] wl[49] vdd gnd cell_6t
Xbit_r50_c255 bl[255] br[255] wl[50] vdd gnd cell_6t
Xbit_r51_c255 bl[255] br[255] wl[51] vdd gnd cell_6t
Xbit_r52_c255 bl[255] br[255] wl[52] vdd gnd cell_6t
Xbit_r53_c255 bl[255] br[255] wl[53] vdd gnd cell_6t
Xbit_r54_c255 bl[255] br[255] wl[54] vdd gnd cell_6t
Xbit_r55_c255 bl[255] br[255] wl[55] vdd gnd cell_6t
Xbit_r56_c255 bl[255] br[255] wl[56] vdd gnd cell_6t
Xbit_r57_c255 bl[255] br[255] wl[57] vdd gnd cell_6t
Xbit_r58_c255 bl[255] br[255] wl[58] vdd gnd cell_6t
Xbit_r59_c255 bl[255] br[255] wl[59] vdd gnd cell_6t
Xbit_r60_c255 bl[255] br[255] wl[60] vdd gnd cell_6t
Xbit_r61_c255 bl[255] br[255] wl[61] vdd gnd cell_6t
Xbit_r62_c255 bl[255] br[255] wl[62] vdd gnd cell_6t
Xbit_r63_c255 bl[255] br[255] wl[63] vdd gnd cell_6t
Xbit_r64_c255 bl[255] br[255] wl[64] vdd gnd cell_6t
Xbit_r65_c255 bl[255] br[255] wl[65] vdd gnd cell_6t
Xbit_r66_c255 bl[255] br[255] wl[66] vdd gnd cell_6t
Xbit_r67_c255 bl[255] br[255] wl[67] vdd gnd cell_6t
Xbit_r68_c255 bl[255] br[255] wl[68] vdd gnd cell_6t
Xbit_r69_c255 bl[255] br[255] wl[69] vdd gnd cell_6t
Xbit_r70_c255 bl[255] br[255] wl[70] vdd gnd cell_6t
Xbit_r71_c255 bl[255] br[255] wl[71] vdd gnd cell_6t
Xbit_r72_c255 bl[255] br[255] wl[72] vdd gnd cell_6t
Xbit_r73_c255 bl[255] br[255] wl[73] vdd gnd cell_6t
Xbit_r74_c255 bl[255] br[255] wl[74] vdd gnd cell_6t
Xbit_r75_c255 bl[255] br[255] wl[75] vdd gnd cell_6t
Xbit_r76_c255 bl[255] br[255] wl[76] vdd gnd cell_6t
Xbit_r77_c255 bl[255] br[255] wl[77] vdd gnd cell_6t
Xbit_r78_c255 bl[255] br[255] wl[78] vdd gnd cell_6t
Xbit_r79_c255 bl[255] br[255] wl[79] vdd gnd cell_6t
Xbit_r80_c255 bl[255] br[255] wl[80] vdd gnd cell_6t
Xbit_r81_c255 bl[255] br[255] wl[81] vdd gnd cell_6t
Xbit_r82_c255 bl[255] br[255] wl[82] vdd gnd cell_6t
Xbit_r83_c255 bl[255] br[255] wl[83] vdd gnd cell_6t
Xbit_r84_c255 bl[255] br[255] wl[84] vdd gnd cell_6t
Xbit_r85_c255 bl[255] br[255] wl[85] vdd gnd cell_6t
Xbit_r86_c255 bl[255] br[255] wl[86] vdd gnd cell_6t
Xbit_r87_c255 bl[255] br[255] wl[87] vdd gnd cell_6t
Xbit_r88_c255 bl[255] br[255] wl[88] vdd gnd cell_6t
Xbit_r89_c255 bl[255] br[255] wl[89] vdd gnd cell_6t
Xbit_r90_c255 bl[255] br[255] wl[90] vdd gnd cell_6t
Xbit_r91_c255 bl[255] br[255] wl[91] vdd gnd cell_6t
Xbit_r92_c255 bl[255] br[255] wl[92] vdd gnd cell_6t
Xbit_r93_c255 bl[255] br[255] wl[93] vdd gnd cell_6t
Xbit_r94_c255 bl[255] br[255] wl[94] vdd gnd cell_6t
Xbit_r95_c255 bl[255] br[255] wl[95] vdd gnd cell_6t
Xbit_r96_c255 bl[255] br[255] wl[96] vdd gnd cell_6t
Xbit_r97_c255 bl[255] br[255] wl[97] vdd gnd cell_6t
Xbit_r98_c255 bl[255] br[255] wl[98] vdd gnd cell_6t
Xbit_r99_c255 bl[255] br[255] wl[99] vdd gnd cell_6t
Xbit_r100_c255 bl[255] br[255] wl[100] vdd gnd cell_6t
Xbit_r101_c255 bl[255] br[255] wl[101] vdd gnd cell_6t
Xbit_r102_c255 bl[255] br[255] wl[102] vdd gnd cell_6t
Xbit_r103_c255 bl[255] br[255] wl[103] vdd gnd cell_6t
Xbit_r104_c255 bl[255] br[255] wl[104] vdd gnd cell_6t
Xbit_r105_c255 bl[255] br[255] wl[105] vdd gnd cell_6t
Xbit_r106_c255 bl[255] br[255] wl[106] vdd gnd cell_6t
Xbit_r107_c255 bl[255] br[255] wl[107] vdd gnd cell_6t
Xbit_r108_c255 bl[255] br[255] wl[108] vdd gnd cell_6t
Xbit_r109_c255 bl[255] br[255] wl[109] vdd gnd cell_6t
Xbit_r110_c255 bl[255] br[255] wl[110] vdd gnd cell_6t
Xbit_r111_c255 bl[255] br[255] wl[111] vdd gnd cell_6t
Xbit_r112_c255 bl[255] br[255] wl[112] vdd gnd cell_6t
Xbit_r113_c255 bl[255] br[255] wl[113] vdd gnd cell_6t
Xbit_r114_c255 bl[255] br[255] wl[114] vdd gnd cell_6t
Xbit_r115_c255 bl[255] br[255] wl[115] vdd gnd cell_6t
Xbit_r116_c255 bl[255] br[255] wl[116] vdd gnd cell_6t
Xbit_r117_c255 bl[255] br[255] wl[117] vdd gnd cell_6t
Xbit_r118_c255 bl[255] br[255] wl[118] vdd gnd cell_6t
Xbit_r119_c255 bl[255] br[255] wl[119] vdd gnd cell_6t
Xbit_r120_c255 bl[255] br[255] wl[120] vdd gnd cell_6t
Xbit_r121_c255 bl[255] br[255] wl[121] vdd gnd cell_6t
Xbit_r122_c255 bl[255] br[255] wl[122] vdd gnd cell_6t
Xbit_r123_c255 bl[255] br[255] wl[123] vdd gnd cell_6t
Xbit_r124_c255 bl[255] br[255] wl[124] vdd gnd cell_6t
Xbit_r125_c255 bl[255] br[255] wl[125] vdd gnd cell_6t
Xbit_r126_c255 bl[255] br[255] wl[126] vdd gnd cell_6t
Xbit_r127_c255 bl[255] br[255] wl[127] vdd gnd cell_6t
.ENDS bitcell_array

* ptx M{0} {1} p m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p

.SUBCKT precharge bl br en vdd
Mlower_pmos bl en BR vdd p m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mupper_pmos1 bl en vdd vdd p m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mupper_pmos2 br en vdd vdd p m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
.ENDS precharge

.SUBCKT precharge_array bl[0] br[0] bl[1] br[1] bl[2] br[2] bl[3] br[3] bl[4] br[4] bl[5] br[5] bl[6] br[6] bl[7] br[7] bl[8] br[8] bl[9] br[9] bl[10] br[10] bl[11] br[11] bl[12] br[12] bl[13] br[13] bl[14] br[14] bl[15] br[15] bl[16] br[16] bl[17] br[17] bl[18] br[18] bl[19] br[19] bl[20] br[20] bl[21] br[21] bl[22] br[22] bl[23] br[23] bl[24] br[24] bl[25] br[25] bl[26] br[26] bl[27] br[27] bl[28] br[28] bl[29] br[29] bl[30] br[30] bl[31] br[31] bl[32] br[32] bl[33] br[33] bl[34] br[34] bl[35] br[35] bl[36] br[36] bl[37] br[37] bl[38] br[38] bl[39] br[39] bl[40] br[40] bl[41] br[41] bl[42] br[42] bl[43] br[43] bl[44] br[44] bl[45] br[45] bl[46] br[46] bl[47] br[47] bl[48] br[48] bl[49] br[49] bl[50] br[50] bl[51] br[51] bl[52] br[52] bl[53] br[53] bl[54] br[54] bl[55] br[55] bl[56] br[56] bl[57] br[57] bl[58] br[58] bl[59] br[59] bl[60] br[60] bl[61] br[61] bl[62] br[62] bl[63] br[63] bl[64] br[64] bl[65] br[65] bl[66] br[66] bl[67] br[67] bl[68] br[68] bl[69] br[69] bl[70] br[70] bl[71] br[71] bl[72] br[72] bl[73] br[73] bl[74] br[74] bl[75] br[75] bl[76] br[76] bl[77] br[77] bl[78] br[78] bl[79] br[79] bl[80] br[80] bl[81] br[81] bl[82] br[82] bl[83] br[83] bl[84] br[84] bl[85] br[85] bl[86] br[86] bl[87] br[87] bl[88] br[88] bl[89] br[89] bl[90] br[90] bl[91] br[91] bl[92] br[92] bl[93] br[93] bl[94] br[94] bl[95] br[95] bl[96] br[96] bl[97] br[97] bl[98] br[98] bl[99] br[99] bl[100] br[100] bl[101] br[101] bl[102] br[102] bl[103] br[103] bl[104] br[104] bl[105] br[105] bl[106] br[106] bl[107] br[107] bl[108] br[108] bl[109] br[109] bl[110] br[110] bl[111] br[111] bl[112] br[112] bl[113] br[113] bl[114] br[114] bl[115] br[115] bl[116] br[116] bl[117] br[117] bl[118] br[118] bl[119] br[119] bl[120] br[120] bl[121] br[121] bl[122] br[122] bl[123] br[123] bl[124] br[124] bl[125] br[125] bl[126] br[126] bl[127] br[127] bl[128] br[128] bl[129] br[129] bl[130] br[130] bl[131] br[131] bl[132] br[132] bl[133] br[133] bl[134] br[134] bl[135] br[135] bl[136] br[136] bl[137] br[137] bl[138] br[138] bl[139] br[139] bl[140] br[140] bl[141] br[141] bl[142] br[142] bl[143] br[143] bl[144] br[144] bl[145] br[145] bl[146] br[146] bl[147] br[147] bl[148] br[148] bl[149] br[149] bl[150] br[150] bl[151] br[151] bl[152] br[152] bl[153] br[153] bl[154] br[154] bl[155] br[155] bl[156] br[156] bl[157] br[157] bl[158] br[158] bl[159] br[159] bl[160] br[160] bl[161] br[161] bl[162] br[162] bl[163] br[163] bl[164] br[164] bl[165] br[165] bl[166] br[166] bl[167] br[167] bl[168] br[168] bl[169] br[169] bl[170] br[170] bl[171] br[171] bl[172] br[172] bl[173] br[173] bl[174] br[174] bl[175] br[175] bl[176] br[176] bl[177] br[177] bl[178] br[178] bl[179] br[179] bl[180] br[180] bl[181] br[181] bl[182] br[182] bl[183] br[183] bl[184] br[184] bl[185] br[185] bl[186] br[186] bl[187] br[187] bl[188] br[188] bl[189] br[189] bl[190] br[190] bl[191] br[191] bl[192] br[192] bl[193] br[193] bl[194] br[194] bl[195] br[195] bl[196] br[196] bl[197] br[197] bl[198] br[198] bl[199] br[199] bl[200] br[200] bl[201] br[201] bl[202] br[202] bl[203] br[203] bl[204] br[204] bl[205] br[205] bl[206] br[206] bl[207] br[207] bl[208] br[208] bl[209] br[209] bl[210] br[210] bl[211] br[211] bl[212] br[212] bl[213] br[213] bl[214] br[214] bl[215] br[215] bl[216] br[216] bl[217] br[217] bl[218] br[218] bl[219] br[219] bl[220] br[220] bl[221] br[221] bl[222] br[222] bl[223] br[223] bl[224] br[224] bl[225] br[225] bl[226] br[226] bl[227] br[227] bl[228] br[228] bl[229] br[229] bl[230] br[230] bl[231] br[231] bl[232] br[232] bl[233] br[233] bl[234] br[234] bl[235] br[235] bl[236] br[236] bl[237] br[237] bl[238] br[238] bl[239] br[239] bl[240] br[240] bl[241] br[241] bl[242] br[242] bl[243] br[243] bl[244] br[244] bl[245] br[245] bl[246] br[246] bl[247] br[247] bl[248] br[248] bl[249] br[249] bl[250] br[250] bl[251] br[251] bl[252] br[252] bl[253] br[253] bl[254] br[254] bl[255] br[255] en vdd
Xpre_column_0 bl[0] br[0] en vdd precharge
Xpre_column_1 bl[1] br[1] en vdd precharge
Xpre_column_2 bl[2] br[2] en vdd precharge
Xpre_column_3 bl[3] br[3] en vdd precharge
Xpre_column_4 bl[4] br[4] en vdd precharge
Xpre_column_5 bl[5] br[5] en vdd precharge
Xpre_column_6 bl[6] br[6] en vdd precharge
Xpre_column_7 bl[7] br[7] en vdd precharge
Xpre_column_8 bl[8] br[8] en vdd precharge
Xpre_column_9 bl[9] br[9] en vdd precharge
Xpre_column_10 bl[10] br[10] en vdd precharge
Xpre_column_11 bl[11] br[11] en vdd precharge
Xpre_column_12 bl[12] br[12] en vdd precharge
Xpre_column_13 bl[13] br[13] en vdd precharge
Xpre_column_14 bl[14] br[14] en vdd precharge
Xpre_column_15 bl[15] br[15] en vdd precharge
Xpre_column_16 bl[16] br[16] en vdd precharge
Xpre_column_17 bl[17] br[17] en vdd precharge
Xpre_column_18 bl[18] br[18] en vdd precharge
Xpre_column_19 bl[19] br[19] en vdd precharge
Xpre_column_20 bl[20] br[20] en vdd precharge
Xpre_column_21 bl[21] br[21] en vdd precharge
Xpre_column_22 bl[22] br[22] en vdd precharge
Xpre_column_23 bl[23] br[23] en vdd precharge
Xpre_column_24 bl[24] br[24] en vdd precharge
Xpre_column_25 bl[25] br[25] en vdd precharge
Xpre_column_26 bl[26] br[26] en vdd precharge
Xpre_column_27 bl[27] br[27] en vdd precharge
Xpre_column_28 bl[28] br[28] en vdd precharge
Xpre_column_29 bl[29] br[29] en vdd precharge
Xpre_column_30 bl[30] br[30] en vdd precharge
Xpre_column_31 bl[31] br[31] en vdd precharge
Xpre_column_32 bl[32] br[32] en vdd precharge
Xpre_column_33 bl[33] br[33] en vdd precharge
Xpre_column_34 bl[34] br[34] en vdd precharge
Xpre_column_35 bl[35] br[35] en vdd precharge
Xpre_column_36 bl[36] br[36] en vdd precharge
Xpre_column_37 bl[37] br[37] en vdd precharge
Xpre_column_38 bl[38] br[38] en vdd precharge
Xpre_column_39 bl[39] br[39] en vdd precharge
Xpre_column_40 bl[40] br[40] en vdd precharge
Xpre_column_41 bl[41] br[41] en vdd precharge
Xpre_column_42 bl[42] br[42] en vdd precharge
Xpre_column_43 bl[43] br[43] en vdd precharge
Xpre_column_44 bl[44] br[44] en vdd precharge
Xpre_column_45 bl[45] br[45] en vdd precharge
Xpre_column_46 bl[46] br[46] en vdd precharge
Xpre_column_47 bl[47] br[47] en vdd precharge
Xpre_column_48 bl[48] br[48] en vdd precharge
Xpre_column_49 bl[49] br[49] en vdd precharge
Xpre_column_50 bl[50] br[50] en vdd precharge
Xpre_column_51 bl[51] br[51] en vdd precharge
Xpre_column_52 bl[52] br[52] en vdd precharge
Xpre_column_53 bl[53] br[53] en vdd precharge
Xpre_column_54 bl[54] br[54] en vdd precharge
Xpre_column_55 bl[55] br[55] en vdd precharge
Xpre_column_56 bl[56] br[56] en vdd precharge
Xpre_column_57 bl[57] br[57] en vdd precharge
Xpre_column_58 bl[58] br[58] en vdd precharge
Xpre_column_59 bl[59] br[59] en vdd precharge
Xpre_column_60 bl[60] br[60] en vdd precharge
Xpre_column_61 bl[61] br[61] en vdd precharge
Xpre_column_62 bl[62] br[62] en vdd precharge
Xpre_column_63 bl[63] br[63] en vdd precharge
Xpre_column_64 bl[64] br[64] en vdd precharge
Xpre_column_65 bl[65] br[65] en vdd precharge
Xpre_column_66 bl[66] br[66] en vdd precharge
Xpre_column_67 bl[67] br[67] en vdd precharge
Xpre_column_68 bl[68] br[68] en vdd precharge
Xpre_column_69 bl[69] br[69] en vdd precharge
Xpre_column_70 bl[70] br[70] en vdd precharge
Xpre_column_71 bl[71] br[71] en vdd precharge
Xpre_column_72 bl[72] br[72] en vdd precharge
Xpre_column_73 bl[73] br[73] en vdd precharge
Xpre_column_74 bl[74] br[74] en vdd precharge
Xpre_column_75 bl[75] br[75] en vdd precharge
Xpre_column_76 bl[76] br[76] en vdd precharge
Xpre_column_77 bl[77] br[77] en vdd precharge
Xpre_column_78 bl[78] br[78] en vdd precharge
Xpre_column_79 bl[79] br[79] en vdd precharge
Xpre_column_80 bl[80] br[80] en vdd precharge
Xpre_column_81 bl[81] br[81] en vdd precharge
Xpre_column_82 bl[82] br[82] en vdd precharge
Xpre_column_83 bl[83] br[83] en vdd precharge
Xpre_column_84 bl[84] br[84] en vdd precharge
Xpre_column_85 bl[85] br[85] en vdd precharge
Xpre_column_86 bl[86] br[86] en vdd precharge
Xpre_column_87 bl[87] br[87] en vdd precharge
Xpre_column_88 bl[88] br[88] en vdd precharge
Xpre_column_89 bl[89] br[89] en vdd precharge
Xpre_column_90 bl[90] br[90] en vdd precharge
Xpre_column_91 bl[91] br[91] en vdd precharge
Xpre_column_92 bl[92] br[92] en vdd precharge
Xpre_column_93 bl[93] br[93] en vdd precharge
Xpre_column_94 bl[94] br[94] en vdd precharge
Xpre_column_95 bl[95] br[95] en vdd precharge
Xpre_column_96 bl[96] br[96] en vdd precharge
Xpre_column_97 bl[97] br[97] en vdd precharge
Xpre_column_98 bl[98] br[98] en vdd precharge
Xpre_column_99 bl[99] br[99] en vdd precharge
Xpre_column_100 bl[100] br[100] en vdd precharge
Xpre_column_101 bl[101] br[101] en vdd precharge
Xpre_column_102 bl[102] br[102] en vdd precharge
Xpre_column_103 bl[103] br[103] en vdd precharge
Xpre_column_104 bl[104] br[104] en vdd precharge
Xpre_column_105 bl[105] br[105] en vdd precharge
Xpre_column_106 bl[106] br[106] en vdd precharge
Xpre_column_107 bl[107] br[107] en vdd precharge
Xpre_column_108 bl[108] br[108] en vdd precharge
Xpre_column_109 bl[109] br[109] en vdd precharge
Xpre_column_110 bl[110] br[110] en vdd precharge
Xpre_column_111 bl[111] br[111] en vdd precharge
Xpre_column_112 bl[112] br[112] en vdd precharge
Xpre_column_113 bl[113] br[113] en vdd precharge
Xpre_column_114 bl[114] br[114] en vdd precharge
Xpre_column_115 bl[115] br[115] en vdd precharge
Xpre_column_116 bl[116] br[116] en vdd precharge
Xpre_column_117 bl[117] br[117] en vdd precharge
Xpre_column_118 bl[118] br[118] en vdd precharge
Xpre_column_119 bl[119] br[119] en vdd precharge
Xpre_column_120 bl[120] br[120] en vdd precharge
Xpre_column_121 bl[121] br[121] en vdd precharge
Xpre_column_122 bl[122] br[122] en vdd precharge
Xpre_column_123 bl[123] br[123] en vdd precharge
Xpre_column_124 bl[124] br[124] en vdd precharge
Xpre_column_125 bl[125] br[125] en vdd precharge
Xpre_column_126 bl[126] br[126] en vdd precharge
Xpre_column_127 bl[127] br[127] en vdd precharge
Xpre_column_128 bl[128] br[128] en vdd precharge
Xpre_column_129 bl[129] br[129] en vdd precharge
Xpre_column_130 bl[130] br[130] en vdd precharge
Xpre_column_131 bl[131] br[131] en vdd precharge
Xpre_column_132 bl[132] br[132] en vdd precharge
Xpre_column_133 bl[133] br[133] en vdd precharge
Xpre_column_134 bl[134] br[134] en vdd precharge
Xpre_column_135 bl[135] br[135] en vdd precharge
Xpre_column_136 bl[136] br[136] en vdd precharge
Xpre_column_137 bl[137] br[137] en vdd precharge
Xpre_column_138 bl[138] br[138] en vdd precharge
Xpre_column_139 bl[139] br[139] en vdd precharge
Xpre_column_140 bl[140] br[140] en vdd precharge
Xpre_column_141 bl[141] br[141] en vdd precharge
Xpre_column_142 bl[142] br[142] en vdd precharge
Xpre_column_143 bl[143] br[143] en vdd precharge
Xpre_column_144 bl[144] br[144] en vdd precharge
Xpre_column_145 bl[145] br[145] en vdd precharge
Xpre_column_146 bl[146] br[146] en vdd precharge
Xpre_column_147 bl[147] br[147] en vdd precharge
Xpre_column_148 bl[148] br[148] en vdd precharge
Xpre_column_149 bl[149] br[149] en vdd precharge
Xpre_column_150 bl[150] br[150] en vdd precharge
Xpre_column_151 bl[151] br[151] en vdd precharge
Xpre_column_152 bl[152] br[152] en vdd precharge
Xpre_column_153 bl[153] br[153] en vdd precharge
Xpre_column_154 bl[154] br[154] en vdd precharge
Xpre_column_155 bl[155] br[155] en vdd precharge
Xpre_column_156 bl[156] br[156] en vdd precharge
Xpre_column_157 bl[157] br[157] en vdd precharge
Xpre_column_158 bl[158] br[158] en vdd precharge
Xpre_column_159 bl[159] br[159] en vdd precharge
Xpre_column_160 bl[160] br[160] en vdd precharge
Xpre_column_161 bl[161] br[161] en vdd precharge
Xpre_column_162 bl[162] br[162] en vdd precharge
Xpre_column_163 bl[163] br[163] en vdd precharge
Xpre_column_164 bl[164] br[164] en vdd precharge
Xpre_column_165 bl[165] br[165] en vdd precharge
Xpre_column_166 bl[166] br[166] en vdd precharge
Xpre_column_167 bl[167] br[167] en vdd precharge
Xpre_column_168 bl[168] br[168] en vdd precharge
Xpre_column_169 bl[169] br[169] en vdd precharge
Xpre_column_170 bl[170] br[170] en vdd precharge
Xpre_column_171 bl[171] br[171] en vdd precharge
Xpre_column_172 bl[172] br[172] en vdd precharge
Xpre_column_173 bl[173] br[173] en vdd precharge
Xpre_column_174 bl[174] br[174] en vdd precharge
Xpre_column_175 bl[175] br[175] en vdd precharge
Xpre_column_176 bl[176] br[176] en vdd precharge
Xpre_column_177 bl[177] br[177] en vdd precharge
Xpre_column_178 bl[178] br[178] en vdd precharge
Xpre_column_179 bl[179] br[179] en vdd precharge
Xpre_column_180 bl[180] br[180] en vdd precharge
Xpre_column_181 bl[181] br[181] en vdd precharge
Xpre_column_182 bl[182] br[182] en vdd precharge
Xpre_column_183 bl[183] br[183] en vdd precharge
Xpre_column_184 bl[184] br[184] en vdd precharge
Xpre_column_185 bl[185] br[185] en vdd precharge
Xpre_column_186 bl[186] br[186] en vdd precharge
Xpre_column_187 bl[187] br[187] en vdd precharge
Xpre_column_188 bl[188] br[188] en vdd precharge
Xpre_column_189 bl[189] br[189] en vdd precharge
Xpre_column_190 bl[190] br[190] en vdd precharge
Xpre_column_191 bl[191] br[191] en vdd precharge
Xpre_column_192 bl[192] br[192] en vdd precharge
Xpre_column_193 bl[193] br[193] en vdd precharge
Xpre_column_194 bl[194] br[194] en vdd precharge
Xpre_column_195 bl[195] br[195] en vdd precharge
Xpre_column_196 bl[196] br[196] en vdd precharge
Xpre_column_197 bl[197] br[197] en vdd precharge
Xpre_column_198 bl[198] br[198] en vdd precharge
Xpre_column_199 bl[199] br[199] en vdd precharge
Xpre_column_200 bl[200] br[200] en vdd precharge
Xpre_column_201 bl[201] br[201] en vdd precharge
Xpre_column_202 bl[202] br[202] en vdd precharge
Xpre_column_203 bl[203] br[203] en vdd precharge
Xpre_column_204 bl[204] br[204] en vdd precharge
Xpre_column_205 bl[205] br[205] en vdd precharge
Xpre_column_206 bl[206] br[206] en vdd precharge
Xpre_column_207 bl[207] br[207] en vdd precharge
Xpre_column_208 bl[208] br[208] en vdd precharge
Xpre_column_209 bl[209] br[209] en vdd precharge
Xpre_column_210 bl[210] br[210] en vdd precharge
Xpre_column_211 bl[211] br[211] en vdd precharge
Xpre_column_212 bl[212] br[212] en vdd precharge
Xpre_column_213 bl[213] br[213] en vdd precharge
Xpre_column_214 bl[214] br[214] en vdd precharge
Xpre_column_215 bl[215] br[215] en vdd precharge
Xpre_column_216 bl[216] br[216] en vdd precharge
Xpre_column_217 bl[217] br[217] en vdd precharge
Xpre_column_218 bl[218] br[218] en vdd precharge
Xpre_column_219 bl[219] br[219] en vdd precharge
Xpre_column_220 bl[220] br[220] en vdd precharge
Xpre_column_221 bl[221] br[221] en vdd precharge
Xpre_column_222 bl[222] br[222] en vdd precharge
Xpre_column_223 bl[223] br[223] en vdd precharge
Xpre_column_224 bl[224] br[224] en vdd precharge
Xpre_column_225 bl[225] br[225] en vdd precharge
Xpre_column_226 bl[226] br[226] en vdd precharge
Xpre_column_227 bl[227] br[227] en vdd precharge
Xpre_column_228 bl[228] br[228] en vdd precharge
Xpre_column_229 bl[229] br[229] en vdd precharge
Xpre_column_230 bl[230] br[230] en vdd precharge
Xpre_column_231 bl[231] br[231] en vdd precharge
Xpre_column_232 bl[232] br[232] en vdd precharge
Xpre_column_233 bl[233] br[233] en vdd precharge
Xpre_column_234 bl[234] br[234] en vdd precharge
Xpre_column_235 bl[235] br[235] en vdd precharge
Xpre_column_236 bl[236] br[236] en vdd precharge
Xpre_column_237 bl[237] br[237] en vdd precharge
Xpre_column_238 bl[238] br[238] en vdd precharge
Xpre_column_239 bl[239] br[239] en vdd precharge
Xpre_column_240 bl[240] br[240] en vdd precharge
Xpre_column_241 bl[241] br[241] en vdd precharge
Xpre_column_242 bl[242] br[242] en vdd precharge
Xpre_column_243 bl[243] br[243] en vdd precharge
Xpre_column_244 bl[244] br[244] en vdd precharge
Xpre_column_245 bl[245] br[245] en vdd precharge
Xpre_column_246 bl[246] br[246] en vdd precharge
Xpre_column_247 bl[247] br[247] en vdd precharge
Xpre_column_248 bl[248] br[248] en vdd precharge
Xpre_column_249 bl[249] br[249] en vdd precharge
Xpre_column_250 bl[250] br[250] en vdd precharge
Xpre_column_251 bl[251] br[251] en vdd precharge
Xpre_column_252 bl[252] br[252] en vdd precharge
Xpre_column_253 bl[253] br[253] en vdd precharge
Xpre_column_254 bl[254] br[254] en vdd precharge
Xpre_column_255 bl[255] br[255] en vdd precharge
.ENDS precharge_array

* ptx M{0} {1} n m=1 w=9.6u l=0.6u pd=20.4u ps=20.4u as=14.4p ad=14.4p

.SUBCKT single_level_column_mux_8 bl br bl_out br_out sel gnd
Mmux_tx1 bl sel bl_out gnd n m=1 w=9.6u l=0.6u pd=20.4u ps=20.4u as=14.4p ad=14.4p
Mmux_tx2 br sel br_out gnd n m=1 w=9.6u l=0.6u pd=20.4u ps=20.4u as=14.4p ad=14.4p
.ENDS single_level_column_mux_8

.SUBCKT columnmux_array bl[0] br[0] bl[1] br[1] bl[2] br[2] bl[3] br[3] bl[4] br[4] bl[5] br[5] bl[6] br[6] bl[7] br[7] bl[8] br[8] bl[9] br[9] bl[10] br[10] bl[11] br[11] bl[12] br[12] bl[13] br[13] bl[14] br[14] bl[15] br[15] bl[16] br[16] bl[17] br[17] bl[18] br[18] bl[19] br[19] bl[20] br[20] bl[21] br[21] bl[22] br[22] bl[23] br[23] bl[24] br[24] bl[25] br[25] bl[26] br[26] bl[27] br[27] bl[28] br[28] bl[29] br[29] bl[30] br[30] bl[31] br[31] bl[32] br[32] bl[33] br[33] bl[34] br[34] bl[35] br[35] bl[36] br[36] bl[37] br[37] bl[38] br[38] bl[39] br[39] bl[40] br[40] bl[41] br[41] bl[42] br[42] bl[43] br[43] bl[44] br[44] bl[45] br[45] bl[46] br[46] bl[47] br[47] bl[48] br[48] bl[49] br[49] bl[50] br[50] bl[51] br[51] bl[52] br[52] bl[53] br[53] bl[54] br[54] bl[55] br[55] bl[56] br[56] bl[57] br[57] bl[58] br[58] bl[59] br[59] bl[60] br[60] bl[61] br[61] bl[62] br[62] bl[63] br[63] bl[64] br[64] bl[65] br[65] bl[66] br[66] bl[67] br[67] bl[68] br[68] bl[69] br[69] bl[70] br[70] bl[71] br[71] bl[72] br[72] bl[73] br[73] bl[74] br[74] bl[75] br[75] bl[76] br[76] bl[77] br[77] bl[78] br[78] bl[79] br[79] bl[80] br[80] bl[81] br[81] bl[82] br[82] bl[83] br[83] bl[84] br[84] bl[85] br[85] bl[86] br[86] bl[87] br[87] bl[88] br[88] bl[89] br[89] bl[90] br[90] bl[91] br[91] bl[92] br[92] bl[93] br[93] bl[94] br[94] bl[95] br[95] bl[96] br[96] bl[97] br[97] bl[98] br[98] bl[99] br[99] bl[100] br[100] bl[101] br[101] bl[102] br[102] bl[103] br[103] bl[104] br[104] bl[105] br[105] bl[106] br[106] bl[107] br[107] bl[108] br[108] bl[109] br[109] bl[110] br[110] bl[111] br[111] bl[112] br[112] bl[113] br[113] bl[114] br[114] bl[115] br[115] bl[116] br[116] bl[117] br[117] bl[118] br[118] bl[119] br[119] bl[120] br[120] bl[121] br[121] bl[122] br[122] bl[123] br[123] bl[124] br[124] bl[125] br[125] bl[126] br[126] bl[127] br[127] bl[128] br[128] bl[129] br[129] bl[130] br[130] bl[131] br[131] bl[132] br[132] bl[133] br[133] bl[134] br[134] bl[135] br[135] bl[136] br[136] bl[137] br[137] bl[138] br[138] bl[139] br[139] bl[140] br[140] bl[141] br[141] bl[142] br[142] bl[143] br[143] bl[144] br[144] bl[145] br[145] bl[146] br[146] bl[147] br[147] bl[148] br[148] bl[149] br[149] bl[150] br[150] bl[151] br[151] bl[152] br[152] bl[153] br[153] bl[154] br[154] bl[155] br[155] bl[156] br[156] bl[157] br[157] bl[158] br[158] bl[159] br[159] bl[160] br[160] bl[161] br[161] bl[162] br[162] bl[163] br[163] bl[164] br[164] bl[165] br[165] bl[166] br[166] bl[167] br[167] bl[168] br[168] bl[169] br[169] bl[170] br[170] bl[171] br[171] bl[172] br[172] bl[173] br[173] bl[174] br[174] bl[175] br[175] bl[176] br[176] bl[177] br[177] bl[178] br[178] bl[179] br[179] bl[180] br[180] bl[181] br[181] bl[182] br[182] bl[183] br[183] bl[184] br[184] bl[185] br[185] bl[186] br[186] bl[187] br[187] bl[188] br[188] bl[189] br[189] bl[190] br[190] bl[191] br[191] bl[192] br[192] bl[193] br[193] bl[194] br[194] bl[195] br[195] bl[196] br[196] bl[197] br[197] bl[198] br[198] bl[199] br[199] bl[200] br[200] bl[201] br[201] bl[202] br[202] bl[203] br[203] bl[204] br[204] bl[205] br[205] bl[206] br[206] bl[207] br[207] bl[208] br[208] bl[209] br[209] bl[210] br[210] bl[211] br[211] bl[212] br[212] bl[213] br[213] bl[214] br[214] bl[215] br[215] bl[216] br[216] bl[217] br[217] bl[218] br[218] bl[219] br[219] bl[220] br[220] bl[221] br[221] bl[222] br[222] bl[223] br[223] bl[224] br[224] bl[225] br[225] bl[226] br[226] bl[227] br[227] bl[228] br[228] bl[229] br[229] bl[230] br[230] bl[231] br[231] bl[232] br[232] bl[233] br[233] bl[234] br[234] bl[235] br[235] bl[236] br[236] bl[237] br[237] bl[238] br[238] bl[239] br[239] bl[240] br[240] bl[241] br[241] bl[242] br[242] bl[243] br[243] bl[244] br[244] bl[245] br[245] bl[246] br[246] bl[247] br[247] bl[248] br[248] bl[249] br[249] bl[250] br[250] bl[251] br[251] bl[252] br[252] bl[253] br[253] bl[254] br[254] bl[255] br[255] sel[0] sel[1] bl_out[0] br_out[0] bl_out[1] br_out[1] bl_out[2] br_out[2] bl_out[3] br_out[3] bl_out[4] br_out[4] bl_out[5] br_out[5] bl_out[6] br_out[6] bl_out[7] br_out[7] bl_out[8] br_out[8] bl_out[9] br_out[9] bl_out[10] br_out[10] bl_out[11] br_out[11] bl_out[12] br_out[12] bl_out[13] br_out[13] bl_out[14] br_out[14] bl_out[15] br_out[15] bl_out[16] br_out[16] bl_out[17] br_out[17] bl_out[18] br_out[18] bl_out[19] br_out[19] bl_out[20] br_out[20] bl_out[21] br_out[21] bl_out[22] br_out[22] bl_out[23] br_out[23] bl_out[24] br_out[24] bl_out[25] br_out[25] bl_out[26] br_out[26] bl_out[27] br_out[27] bl_out[28] br_out[28] bl_out[29] br_out[29] bl_out[30] br_out[30] bl_out[31] br_out[31] bl_out[32] br_out[32] bl_out[33] br_out[33] bl_out[34] br_out[34] bl_out[35] br_out[35] bl_out[36] br_out[36] bl_out[37] br_out[37] bl_out[38] br_out[38] bl_out[39] br_out[39] bl_out[40] br_out[40] bl_out[41] br_out[41] bl_out[42] br_out[42] bl_out[43] br_out[43] bl_out[44] br_out[44] bl_out[45] br_out[45] bl_out[46] br_out[46] bl_out[47] br_out[47] bl_out[48] br_out[48] bl_out[49] br_out[49] bl_out[50] br_out[50] bl_out[51] br_out[51] bl_out[52] br_out[52] bl_out[53] br_out[53] bl_out[54] br_out[54] bl_out[55] br_out[55] bl_out[56] br_out[56] bl_out[57] br_out[57] bl_out[58] br_out[58] bl_out[59] br_out[59] bl_out[60] br_out[60] bl_out[61] br_out[61] bl_out[62] br_out[62] bl_out[63] br_out[63] bl_out[64] br_out[64] bl_out[65] br_out[65] bl_out[66] br_out[66] bl_out[67] br_out[67] bl_out[68] br_out[68] bl_out[69] br_out[69] bl_out[70] br_out[70] bl_out[71] br_out[71] bl_out[72] br_out[72] bl_out[73] br_out[73] bl_out[74] br_out[74] bl_out[75] br_out[75] bl_out[76] br_out[76] bl_out[77] br_out[77] bl_out[78] br_out[78] bl_out[79] br_out[79] bl_out[80] br_out[80] bl_out[81] br_out[81] bl_out[82] br_out[82] bl_out[83] br_out[83] bl_out[84] br_out[84] bl_out[85] br_out[85] bl_out[86] br_out[86] bl_out[87] br_out[87] bl_out[88] br_out[88] bl_out[89] br_out[89] bl_out[90] br_out[90] bl_out[91] br_out[91] bl_out[92] br_out[92] bl_out[93] br_out[93] bl_out[94] br_out[94] bl_out[95] br_out[95] bl_out[96] br_out[96] bl_out[97] br_out[97] bl_out[98] br_out[98] bl_out[99] br_out[99] bl_out[100] br_out[100] bl_out[101] br_out[101] bl_out[102] br_out[102] bl_out[103] br_out[103] bl_out[104] br_out[104] bl_out[105] br_out[105] bl_out[106] br_out[106] bl_out[107] br_out[107] bl_out[108] br_out[108] bl_out[109] br_out[109] bl_out[110] br_out[110] bl_out[111] br_out[111] bl_out[112] br_out[112] bl_out[113] br_out[113] bl_out[114] br_out[114] bl_out[115] br_out[115] bl_out[116] br_out[116] bl_out[117] br_out[117] bl_out[118] br_out[118] bl_out[119] br_out[119] bl_out[120] br_out[120] bl_out[121] br_out[121] bl_out[122] br_out[122] bl_out[123] br_out[123] bl_out[124] br_out[124] bl_out[125] br_out[125] bl_out[126] br_out[126] bl_out[127] br_out[127] gnd
XXMUX0 bl[0] br[0] bl_out[0] br_out[0] sel[0] gnd single_level_column_mux_8
XXMUX1 bl[1] br[1] bl_out[0] br_out[0] sel[1] gnd single_level_column_mux_8
XXMUX2 bl[2] br[2] bl_out[1] br_out[1] sel[0] gnd single_level_column_mux_8
XXMUX3 bl[3] br[3] bl_out[1] br_out[1] sel[1] gnd single_level_column_mux_8
XXMUX4 bl[4] br[4] bl_out[2] br_out[2] sel[0] gnd single_level_column_mux_8
XXMUX5 bl[5] br[5] bl_out[2] br_out[2] sel[1] gnd single_level_column_mux_8
XXMUX6 bl[6] br[6] bl_out[3] br_out[3] sel[0] gnd single_level_column_mux_8
XXMUX7 bl[7] br[7] bl_out[3] br_out[3] sel[1] gnd single_level_column_mux_8
XXMUX8 bl[8] br[8] bl_out[4] br_out[4] sel[0] gnd single_level_column_mux_8
XXMUX9 bl[9] br[9] bl_out[4] br_out[4] sel[1] gnd single_level_column_mux_8
XXMUX10 bl[10] br[10] bl_out[5] br_out[5] sel[0] gnd single_level_column_mux_8
XXMUX11 bl[11] br[11] bl_out[5] br_out[5] sel[1] gnd single_level_column_mux_8
XXMUX12 bl[12] br[12] bl_out[6] br_out[6] sel[0] gnd single_level_column_mux_8
XXMUX13 bl[13] br[13] bl_out[6] br_out[6] sel[1] gnd single_level_column_mux_8
XXMUX14 bl[14] br[14] bl_out[7] br_out[7] sel[0] gnd single_level_column_mux_8
XXMUX15 bl[15] br[15] bl_out[7] br_out[7] sel[1] gnd single_level_column_mux_8
XXMUX16 bl[16] br[16] bl_out[8] br_out[8] sel[0] gnd single_level_column_mux_8
XXMUX17 bl[17] br[17] bl_out[8] br_out[8] sel[1] gnd single_level_column_mux_8
XXMUX18 bl[18] br[18] bl_out[9] br_out[9] sel[0] gnd single_level_column_mux_8
XXMUX19 bl[19] br[19] bl_out[9] br_out[9] sel[1] gnd single_level_column_mux_8
XXMUX20 bl[20] br[20] bl_out[10] br_out[10] sel[0] gnd single_level_column_mux_8
XXMUX21 bl[21] br[21] bl_out[10] br_out[10] sel[1] gnd single_level_column_mux_8
XXMUX22 bl[22] br[22] bl_out[11] br_out[11] sel[0] gnd single_level_column_mux_8
XXMUX23 bl[23] br[23] bl_out[11] br_out[11] sel[1] gnd single_level_column_mux_8
XXMUX24 bl[24] br[24] bl_out[12] br_out[12] sel[0] gnd single_level_column_mux_8
XXMUX25 bl[25] br[25] bl_out[12] br_out[12] sel[1] gnd single_level_column_mux_8
XXMUX26 bl[26] br[26] bl_out[13] br_out[13] sel[0] gnd single_level_column_mux_8
XXMUX27 bl[27] br[27] bl_out[13] br_out[13] sel[1] gnd single_level_column_mux_8
XXMUX28 bl[28] br[28] bl_out[14] br_out[14] sel[0] gnd single_level_column_mux_8
XXMUX29 bl[29] br[29] bl_out[14] br_out[14] sel[1] gnd single_level_column_mux_8
XXMUX30 bl[30] br[30] bl_out[15] br_out[15] sel[0] gnd single_level_column_mux_8
XXMUX31 bl[31] br[31] bl_out[15] br_out[15] sel[1] gnd single_level_column_mux_8
XXMUX32 bl[32] br[32] bl_out[16] br_out[16] sel[0] gnd single_level_column_mux_8
XXMUX33 bl[33] br[33] bl_out[16] br_out[16] sel[1] gnd single_level_column_mux_8
XXMUX34 bl[34] br[34] bl_out[17] br_out[17] sel[0] gnd single_level_column_mux_8
XXMUX35 bl[35] br[35] bl_out[17] br_out[17] sel[1] gnd single_level_column_mux_8
XXMUX36 bl[36] br[36] bl_out[18] br_out[18] sel[0] gnd single_level_column_mux_8
XXMUX37 bl[37] br[37] bl_out[18] br_out[18] sel[1] gnd single_level_column_mux_8
XXMUX38 bl[38] br[38] bl_out[19] br_out[19] sel[0] gnd single_level_column_mux_8
XXMUX39 bl[39] br[39] bl_out[19] br_out[19] sel[1] gnd single_level_column_mux_8
XXMUX40 bl[40] br[40] bl_out[20] br_out[20] sel[0] gnd single_level_column_mux_8
XXMUX41 bl[41] br[41] bl_out[20] br_out[20] sel[1] gnd single_level_column_mux_8
XXMUX42 bl[42] br[42] bl_out[21] br_out[21] sel[0] gnd single_level_column_mux_8
XXMUX43 bl[43] br[43] bl_out[21] br_out[21] sel[1] gnd single_level_column_mux_8
XXMUX44 bl[44] br[44] bl_out[22] br_out[22] sel[0] gnd single_level_column_mux_8
XXMUX45 bl[45] br[45] bl_out[22] br_out[22] sel[1] gnd single_level_column_mux_8
XXMUX46 bl[46] br[46] bl_out[23] br_out[23] sel[0] gnd single_level_column_mux_8
XXMUX47 bl[47] br[47] bl_out[23] br_out[23] sel[1] gnd single_level_column_mux_8
XXMUX48 bl[48] br[48] bl_out[24] br_out[24] sel[0] gnd single_level_column_mux_8
XXMUX49 bl[49] br[49] bl_out[24] br_out[24] sel[1] gnd single_level_column_mux_8
XXMUX50 bl[50] br[50] bl_out[25] br_out[25] sel[0] gnd single_level_column_mux_8
XXMUX51 bl[51] br[51] bl_out[25] br_out[25] sel[1] gnd single_level_column_mux_8
XXMUX52 bl[52] br[52] bl_out[26] br_out[26] sel[0] gnd single_level_column_mux_8
XXMUX53 bl[53] br[53] bl_out[26] br_out[26] sel[1] gnd single_level_column_mux_8
XXMUX54 bl[54] br[54] bl_out[27] br_out[27] sel[0] gnd single_level_column_mux_8
XXMUX55 bl[55] br[55] bl_out[27] br_out[27] sel[1] gnd single_level_column_mux_8
XXMUX56 bl[56] br[56] bl_out[28] br_out[28] sel[0] gnd single_level_column_mux_8
XXMUX57 bl[57] br[57] bl_out[28] br_out[28] sel[1] gnd single_level_column_mux_8
XXMUX58 bl[58] br[58] bl_out[29] br_out[29] sel[0] gnd single_level_column_mux_8
XXMUX59 bl[59] br[59] bl_out[29] br_out[29] sel[1] gnd single_level_column_mux_8
XXMUX60 bl[60] br[60] bl_out[30] br_out[30] sel[0] gnd single_level_column_mux_8
XXMUX61 bl[61] br[61] bl_out[30] br_out[30] sel[1] gnd single_level_column_mux_8
XXMUX62 bl[62] br[62] bl_out[31] br_out[31] sel[0] gnd single_level_column_mux_8
XXMUX63 bl[63] br[63] bl_out[31] br_out[31] sel[1] gnd single_level_column_mux_8
XXMUX64 bl[64] br[64] bl_out[32] br_out[32] sel[0] gnd single_level_column_mux_8
XXMUX65 bl[65] br[65] bl_out[32] br_out[32] sel[1] gnd single_level_column_mux_8
XXMUX66 bl[66] br[66] bl_out[33] br_out[33] sel[0] gnd single_level_column_mux_8
XXMUX67 bl[67] br[67] bl_out[33] br_out[33] sel[1] gnd single_level_column_mux_8
XXMUX68 bl[68] br[68] bl_out[34] br_out[34] sel[0] gnd single_level_column_mux_8
XXMUX69 bl[69] br[69] bl_out[34] br_out[34] sel[1] gnd single_level_column_mux_8
XXMUX70 bl[70] br[70] bl_out[35] br_out[35] sel[0] gnd single_level_column_mux_8
XXMUX71 bl[71] br[71] bl_out[35] br_out[35] sel[1] gnd single_level_column_mux_8
XXMUX72 bl[72] br[72] bl_out[36] br_out[36] sel[0] gnd single_level_column_mux_8
XXMUX73 bl[73] br[73] bl_out[36] br_out[36] sel[1] gnd single_level_column_mux_8
XXMUX74 bl[74] br[74] bl_out[37] br_out[37] sel[0] gnd single_level_column_mux_8
XXMUX75 bl[75] br[75] bl_out[37] br_out[37] sel[1] gnd single_level_column_mux_8
XXMUX76 bl[76] br[76] bl_out[38] br_out[38] sel[0] gnd single_level_column_mux_8
XXMUX77 bl[77] br[77] bl_out[38] br_out[38] sel[1] gnd single_level_column_mux_8
XXMUX78 bl[78] br[78] bl_out[39] br_out[39] sel[0] gnd single_level_column_mux_8
XXMUX79 bl[79] br[79] bl_out[39] br_out[39] sel[1] gnd single_level_column_mux_8
XXMUX80 bl[80] br[80] bl_out[40] br_out[40] sel[0] gnd single_level_column_mux_8
XXMUX81 bl[81] br[81] bl_out[40] br_out[40] sel[1] gnd single_level_column_mux_8
XXMUX82 bl[82] br[82] bl_out[41] br_out[41] sel[0] gnd single_level_column_mux_8
XXMUX83 bl[83] br[83] bl_out[41] br_out[41] sel[1] gnd single_level_column_mux_8
XXMUX84 bl[84] br[84] bl_out[42] br_out[42] sel[0] gnd single_level_column_mux_8
XXMUX85 bl[85] br[85] bl_out[42] br_out[42] sel[1] gnd single_level_column_mux_8
XXMUX86 bl[86] br[86] bl_out[43] br_out[43] sel[0] gnd single_level_column_mux_8
XXMUX87 bl[87] br[87] bl_out[43] br_out[43] sel[1] gnd single_level_column_mux_8
XXMUX88 bl[88] br[88] bl_out[44] br_out[44] sel[0] gnd single_level_column_mux_8
XXMUX89 bl[89] br[89] bl_out[44] br_out[44] sel[1] gnd single_level_column_mux_8
XXMUX90 bl[90] br[90] bl_out[45] br_out[45] sel[0] gnd single_level_column_mux_8
XXMUX91 bl[91] br[91] bl_out[45] br_out[45] sel[1] gnd single_level_column_mux_8
XXMUX92 bl[92] br[92] bl_out[46] br_out[46] sel[0] gnd single_level_column_mux_8
XXMUX93 bl[93] br[93] bl_out[46] br_out[46] sel[1] gnd single_level_column_mux_8
XXMUX94 bl[94] br[94] bl_out[47] br_out[47] sel[0] gnd single_level_column_mux_8
XXMUX95 bl[95] br[95] bl_out[47] br_out[47] sel[1] gnd single_level_column_mux_8
XXMUX96 bl[96] br[96] bl_out[48] br_out[48] sel[0] gnd single_level_column_mux_8
XXMUX97 bl[97] br[97] bl_out[48] br_out[48] sel[1] gnd single_level_column_mux_8
XXMUX98 bl[98] br[98] bl_out[49] br_out[49] sel[0] gnd single_level_column_mux_8
XXMUX99 bl[99] br[99] bl_out[49] br_out[49] sel[1] gnd single_level_column_mux_8
XXMUX100 bl[100] br[100] bl_out[50] br_out[50] sel[0] gnd single_level_column_mux_8
XXMUX101 bl[101] br[101] bl_out[50] br_out[50] sel[1] gnd single_level_column_mux_8
XXMUX102 bl[102] br[102] bl_out[51] br_out[51] sel[0] gnd single_level_column_mux_8
XXMUX103 bl[103] br[103] bl_out[51] br_out[51] sel[1] gnd single_level_column_mux_8
XXMUX104 bl[104] br[104] bl_out[52] br_out[52] sel[0] gnd single_level_column_mux_8
XXMUX105 bl[105] br[105] bl_out[52] br_out[52] sel[1] gnd single_level_column_mux_8
XXMUX106 bl[106] br[106] bl_out[53] br_out[53] sel[0] gnd single_level_column_mux_8
XXMUX107 bl[107] br[107] bl_out[53] br_out[53] sel[1] gnd single_level_column_mux_8
XXMUX108 bl[108] br[108] bl_out[54] br_out[54] sel[0] gnd single_level_column_mux_8
XXMUX109 bl[109] br[109] bl_out[54] br_out[54] sel[1] gnd single_level_column_mux_8
XXMUX110 bl[110] br[110] bl_out[55] br_out[55] sel[0] gnd single_level_column_mux_8
XXMUX111 bl[111] br[111] bl_out[55] br_out[55] sel[1] gnd single_level_column_mux_8
XXMUX112 bl[112] br[112] bl_out[56] br_out[56] sel[0] gnd single_level_column_mux_8
XXMUX113 bl[113] br[113] bl_out[56] br_out[56] sel[1] gnd single_level_column_mux_8
XXMUX114 bl[114] br[114] bl_out[57] br_out[57] sel[0] gnd single_level_column_mux_8
XXMUX115 bl[115] br[115] bl_out[57] br_out[57] sel[1] gnd single_level_column_mux_8
XXMUX116 bl[116] br[116] bl_out[58] br_out[58] sel[0] gnd single_level_column_mux_8
XXMUX117 bl[117] br[117] bl_out[58] br_out[58] sel[1] gnd single_level_column_mux_8
XXMUX118 bl[118] br[118] bl_out[59] br_out[59] sel[0] gnd single_level_column_mux_8
XXMUX119 bl[119] br[119] bl_out[59] br_out[59] sel[1] gnd single_level_column_mux_8
XXMUX120 bl[120] br[120] bl_out[60] br_out[60] sel[0] gnd single_level_column_mux_8
XXMUX121 bl[121] br[121] bl_out[60] br_out[60] sel[1] gnd single_level_column_mux_8
XXMUX122 bl[122] br[122] bl_out[61] br_out[61] sel[0] gnd single_level_column_mux_8
XXMUX123 bl[123] br[123] bl_out[61] br_out[61] sel[1] gnd single_level_column_mux_8
XXMUX124 bl[124] br[124] bl_out[62] br_out[62] sel[0] gnd single_level_column_mux_8
XXMUX125 bl[125] br[125] bl_out[62] br_out[62] sel[1] gnd single_level_column_mux_8
XXMUX126 bl[126] br[126] bl_out[63] br_out[63] sel[0] gnd single_level_column_mux_8
XXMUX127 bl[127] br[127] bl_out[63] br_out[63] sel[1] gnd single_level_column_mux_8
XXMUX128 bl[128] br[128] bl_out[64] br_out[64] sel[0] gnd single_level_column_mux_8
XXMUX129 bl[129] br[129] bl_out[64] br_out[64] sel[1] gnd single_level_column_mux_8
XXMUX130 bl[130] br[130] bl_out[65] br_out[65] sel[0] gnd single_level_column_mux_8
XXMUX131 bl[131] br[131] bl_out[65] br_out[65] sel[1] gnd single_level_column_mux_8
XXMUX132 bl[132] br[132] bl_out[66] br_out[66] sel[0] gnd single_level_column_mux_8
XXMUX133 bl[133] br[133] bl_out[66] br_out[66] sel[1] gnd single_level_column_mux_8
XXMUX134 bl[134] br[134] bl_out[67] br_out[67] sel[0] gnd single_level_column_mux_8
XXMUX135 bl[135] br[135] bl_out[67] br_out[67] sel[1] gnd single_level_column_mux_8
XXMUX136 bl[136] br[136] bl_out[68] br_out[68] sel[0] gnd single_level_column_mux_8
XXMUX137 bl[137] br[137] bl_out[68] br_out[68] sel[1] gnd single_level_column_mux_8
XXMUX138 bl[138] br[138] bl_out[69] br_out[69] sel[0] gnd single_level_column_mux_8
XXMUX139 bl[139] br[139] bl_out[69] br_out[69] sel[1] gnd single_level_column_mux_8
XXMUX140 bl[140] br[140] bl_out[70] br_out[70] sel[0] gnd single_level_column_mux_8
XXMUX141 bl[141] br[141] bl_out[70] br_out[70] sel[1] gnd single_level_column_mux_8
XXMUX142 bl[142] br[142] bl_out[71] br_out[71] sel[0] gnd single_level_column_mux_8
XXMUX143 bl[143] br[143] bl_out[71] br_out[71] sel[1] gnd single_level_column_mux_8
XXMUX144 bl[144] br[144] bl_out[72] br_out[72] sel[0] gnd single_level_column_mux_8
XXMUX145 bl[145] br[145] bl_out[72] br_out[72] sel[1] gnd single_level_column_mux_8
XXMUX146 bl[146] br[146] bl_out[73] br_out[73] sel[0] gnd single_level_column_mux_8
XXMUX147 bl[147] br[147] bl_out[73] br_out[73] sel[1] gnd single_level_column_mux_8
XXMUX148 bl[148] br[148] bl_out[74] br_out[74] sel[0] gnd single_level_column_mux_8
XXMUX149 bl[149] br[149] bl_out[74] br_out[74] sel[1] gnd single_level_column_mux_8
XXMUX150 bl[150] br[150] bl_out[75] br_out[75] sel[0] gnd single_level_column_mux_8
XXMUX151 bl[151] br[151] bl_out[75] br_out[75] sel[1] gnd single_level_column_mux_8
XXMUX152 bl[152] br[152] bl_out[76] br_out[76] sel[0] gnd single_level_column_mux_8
XXMUX153 bl[153] br[153] bl_out[76] br_out[76] sel[1] gnd single_level_column_mux_8
XXMUX154 bl[154] br[154] bl_out[77] br_out[77] sel[0] gnd single_level_column_mux_8
XXMUX155 bl[155] br[155] bl_out[77] br_out[77] sel[1] gnd single_level_column_mux_8
XXMUX156 bl[156] br[156] bl_out[78] br_out[78] sel[0] gnd single_level_column_mux_8
XXMUX157 bl[157] br[157] bl_out[78] br_out[78] sel[1] gnd single_level_column_mux_8
XXMUX158 bl[158] br[158] bl_out[79] br_out[79] sel[0] gnd single_level_column_mux_8
XXMUX159 bl[159] br[159] bl_out[79] br_out[79] sel[1] gnd single_level_column_mux_8
XXMUX160 bl[160] br[160] bl_out[80] br_out[80] sel[0] gnd single_level_column_mux_8
XXMUX161 bl[161] br[161] bl_out[80] br_out[80] sel[1] gnd single_level_column_mux_8
XXMUX162 bl[162] br[162] bl_out[81] br_out[81] sel[0] gnd single_level_column_mux_8
XXMUX163 bl[163] br[163] bl_out[81] br_out[81] sel[1] gnd single_level_column_mux_8
XXMUX164 bl[164] br[164] bl_out[82] br_out[82] sel[0] gnd single_level_column_mux_8
XXMUX165 bl[165] br[165] bl_out[82] br_out[82] sel[1] gnd single_level_column_mux_8
XXMUX166 bl[166] br[166] bl_out[83] br_out[83] sel[0] gnd single_level_column_mux_8
XXMUX167 bl[167] br[167] bl_out[83] br_out[83] sel[1] gnd single_level_column_mux_8
XXMUX168 bl[168] br[168] bl_out[84] br_out[84] sel[0] gnd single_level_column_mux_8
XXMUX169 bl[169] br[169] bl_out[84] br_out[84] sel[1] gnd single_level_column_mux_8
XXMUX170 bl[170] br[170] bl_out[85] br_out[85] sel[0] gnd single_level_column_mux_8
XXMUX171 bl[171] br[171] bl_out[85] br_out[85] sel[1] gnd single_level_column_mux_8
XXMUX172 bl[172] br[172] bl_out[86] br_out[86] sel[0] gnd single_level_column_mux_8
XXMUX173 bl[173] br[173] bl_out[86] br_out[86] sel[1] gnd single_level_column_mux_8
XXMUX174 bl[174] br[174] bl_out[87] br_out[87] sel[0] gnd single_level_column_mux_8
XXMUX175 bl[175] br[175] bl_out[87] br_out[87] sel[1] gnd single_level_column_mux_8
XXMUX176 bl[176] br[176] bl_out[88] br_out[88] sel[0] gnd single_level_column_mux_8
XXMUX177 bl[177] br[177] bl_out[88] br_out[88] sel[1] gnd single_level_column_mux_8
XXMUX178 bl[178] br[178] bl_out[89] br_out[89] sel[0] gnd single_level_column_mux_8
XXMUX179 bl[179] br[179] bl_out[89] br_out[89] sel[1] gnd single_level_column_mux_8
XXMUX180 bl[180] br[180] bl_out[90] br_out[90] sel[0] gnd single_level_column_mux_8
XXMUX181 bl[181] br[181] bl_out[90] br_out[90] sel[1] gnd single_level_column_mux_8
XXMUX182 bl[182] br[182] bl_out[91] br_out[91] sel[0] gnd single_level_column_mux_8
XXMUX183 bl[183] br[183] bl_out[91] br_out[91] sel[1] gnd single_level_column_mux_8
XXMUX184 bl[184] br[184] bl_out[92] br_out[92] sel[0] gnd single_level_column_mux_8
XXMUX185 bl[185] br[185] bl_out[92] br_out[92] sel[1] gnd single_level_column_mux_8
XXMUX186 bl[186] br[186] bl_out[93] br_out[93] sel[0] gnd single_level_column_mux_8
XXMUX187 bl[187] br[187] bl_out[93] br_out[93] sel[1] gnd single_level_column_mux_8
XXMUX188 bl[188] br[188] bl_out[94] br_out[94] sel[0] gnd single_level_column_mux_8
XXMUX189 bl[189] br[189] bl_out[94] br_out[94] sel[1] gnd single_level_column_mux_8
XXMUX190 bl[190] br[190] bl_out[95] br_out[95] sel[0] gnd single_level_column_mux_8
XXMUX191 bl[191] br[191] bl_out[95] br_out[95] sel[1] gnd single_level_column_mux_8
XXMUX192 bl[192] br[192] bl_out[96] br_out[96] sel[0] gnd single_level_column_mux_8
XXMUX193 bl[193] br[193] bl_out[96] br_out[96] sel[1] gnd single_level_column_mux_8
XXMUX194 bl[194] br[194] bl_out[97] br_out[97] sel[0] gnd single_level_column_mux_8
XXMUX195 bl[195] br[195] bl_out[97] br_out[97] sel[1] gnd single_level_column_mux_8
XXMUX196 bl[196] br[196] bl_out[98] br_out[98] sel[0] gnd single_level_column_mux_8
XXMUX197 bl[197] br[197] bl_out[98] br_out[98] sel[1] gnd single_level_column_mux_8
XXMUX198 bl[198] br[198] bl_out[99] br_out[99] sel[0] gnd single_level_column_mux_8
XXMUX199 bl[199] br[199] bl_out[99] br_out[99] sel[1] gnd single_level_column_mux_8
XXMUX200 bl[200] br[200] bl_out[100] br_out[100] sel[0] gnd single_level_column_mux_8
XXMUX201 bl[201] br[201] bl_out[100] br_out[100] sel[1] gnd single_level_column_mux_8
XXMUX202 bl[202] br[202] bl_out[101] br_out[101] sel[0] gnd single_level_column_mux_8
XXMUX203 bl[203] br[203] bl_out[101] br_out[101] sel[1] gnd single_level_column_mux_8
XXMUX204 bl[204] br[204] bl_out[102] br_out[102] sel[0] gnd single_level_column_mux_8
XXMUX205 bl[205] br[205] bl_out[102] br_out[102] sel[1] gnd single_level_column_mux_8
XXMUX206 bl[206] br[206] bl_out[103] br_out[103] sel[0] gnd single_level_column_mux_8
XXMUX207 bl[207] br[207] bl_out[103] br_out[103] sel[1] gnd single_level_column_mux_8
XXMUX208 bl[208] br[208] bl_out[104] br_out[104] sel[0] gnd single_level_column_mux_8
XXMUX209 bl[209] br[209] bl_out[104] br_out[104] sel[1] gnd single_level_column_mux_8
XXMUX210 bl[210] br[210] bl_out[105] br_out[105] sel[0] gnd single_level_column_mux_8
XXMUX211 bl[211] br[211] bl_out[105] br_out[105] sel[1] gnd single_level_column_mux_8
XXMUX212 bl[212] br[212] bl_out[106] br_out[106] sel[0] gnd single_level_column_mux_8
XXMUX213 bl[213] br[213] bl_out[106] br_out[106] sel[1] gnd single_level_column_mux_8
XXMUX214 bl[214] br[214] bl_out[107] br_out[107] sel[0] gnd single_level_column_mux_8
XXMUX215 bl[215] br[215] bl_out[107] br_out[107] sel[1] gnd single_level_column_mux_8
XXMUX216 bl[216] br[216] bl_out[108] br_out[108] sel[0] gnd single_level_column_mux_8
XXMUX217 bl[217] br[217] bl_out[108] br_out[108] sel[1] gnd single_level_column_mux_8
XXMUX218 bl[218] br[218] bl_out[109] br_out[109] sel[0] gnd single_level_column_mux_8
XXMUX219 bl[219] br[219] bl_out[109] br_out[109] sel[1] gnd single_level_column_mux_8
XXMUX220 bl[220] br[220] bl_out[110] br_out[110] sel[0] gnd single_level_column_mux_8
XXMUX221 bl[221] br[221] bl_out[110] br_out[110] sel[1] gnd single_level_column_mux_8
XXMUX222 bl[222] br[222] bl_out[111] br_out[111] sel[0] gnd single_level_column_mux_8
XXMUX223 bl[223] br[223] bl_out[111] br_out[111] sel[1] gnd single_level_column_mux_8
XXMUX224 bl[224] br[224] bl_out[112] br_out[112] sel[0] gnd single_level_column_mux_8
XXMUX225 bl[225] br[225] bl_out[112] br_out[112] sel[1] gnd single_level_column_mux_8
XXMUX226 bl[226] br[226] bl_out[113] br_out[113] sel[0] gnd single_level_column_mux_8
XXMUX227 bl[227] br[227] bl_out[113] br_out[113] sel[1] gnd single_level_column_mux_8
XXMUX228 bl[228] br[228] bl_out[114] br_out[114] sel[0] gnd single_level_column_mux_8
XXMUX229 bl[229] br[229] bl_out[114] br_out[114] sel[1] gnd single_level_column_mux_8
XXMUX230 bl[230] br[230] bl_out[115] br_out[115] sel[0] gnd single_level_column_mux_8
XXMUX231 bl[231] br[231] bl_out[115] br_out[115] sel[1] gnd single_level_column_mux_8
XXMUX232 bl[232] br[232] bl_out[116] br_out[116] sel[0] gnd single_level_column_mux_8
XXMUX233 bl[233] br[233] bl_out[116] br_out[116] sel[1] gnd single_level_column_mux_8
XXMUX234 bl[234] br[234] bl_out[117] br_out[117] sel[0] gnd single_level_column_mux_8
XXMUX235 bl[235] br[235] bl_out[117] br_out[117] sel[1] gnd single_level_column_mux_8
XXMUX236 bl[236] br[236] bl_out[118] br_out[118] sel[0] gnd single_level_column_mux_8
XXMUX237 bl[237] br[237] bl_out[118] br_out[118] sel[1] gnd single_level_column_mux_8
XXMUX238 bl[238] br[238] bl_out[119] br_out[119] sel[0] gnd single_level_column_mux_8
XXMUX239 bl[239] br[239] bl_out[119] br_out[119] sel[1] gnd single_level_column_mux_8
XXMUX240 bl[240] br[240] bl_out[120] br_out[120] sel[0] gnd single_level_column_mux_8
XXMUX241 bl[241] br[241] bl_out[120] br_out[120] sel[1] gnd single_level_column_mux_8
XXMUX242 bl[242] br[242] bl_out[121] br_out[121] sel[0] gnd single_level_column_mux_8
XXMUX243 bl[243] br[243] bl_out[121] br_out[121] sel[1] gnd single_level_column_mux_8
XXMUX244 bl[244] br[244] bl_out[122] br_out[122] sel[0] gnd single_level_column_mux_8
XXMUX245 bl[245] br[245] bl_out[122] br_out[122] sel[1] gnd single_level_column_mux_8
XXMUX246 bl[246] br[246] bl_out[123] br_out[123] sel[0] gnd single_level_column_mux_8
XXMUX247 bl[247] br[247] bl_out[123] br_out[123] sel[1] gnd single_level_column_mux_8
XXMUX248 bl[248] br[248] bl_out[124] br_out[124] sel[0] gnd single_level_column_mux_8
XXMUX249 bl[249] br[249] bl_out[124] br_out[124] sel[1] gnd single_level_column_mux_8
XXMUX250 bl[250] br[250] bl_out[125] br_out[125] sel[0] gnd single_level_column_mux_8
XXMUX251 bl[251] br[251] bl_out[125] br_out[125] sel[1] gnd single_level_column_mux_8
XXMUX252 bl[252] br[252] bl_out[126] br_out[126] sel[0] gnd single_level_column_mux_8
XXMUX253 bl[253] br[253] bl_out[126] br_out[126] sel[1] gnd single_level_column_mux_8
XXMUX254 bl[254] br[254] bl_out[127] br_out[127] sel[0] gnd single_level_column_mux_8
XXMUX255 bl[255] br[255] bl_out[127] br_out[127] sel[1] gnd single_level_column_mux_8
.ENDS columnmux_array
*********************** "sense_amp" ******************************

.SUBCKT sense_amp bl br dout en vdd gnd
M_1 dout net_1 vdd vdd p W='5.4*1u' L=0.6u
M_2 dout net_1 net_2 gnd n W='2.7*1u' L=0.6u
M_3 net_1 dout vdd vdd p W='5.4*1u' L=0.6u
M_4 net_1 dout net_2 gnd n W='2.7*1u' L=0.6u
M_5 bl en dout vdd p W='7.2*1u' L=0.6u
M_6 br en net_1 vdd p W='7.2*1u' L=0.6u
M_7 net_2 en gnd gnd n W='2.7*1u' L=0.6u
.ENDS	 sense_amp


.SUBCKT sense_amp_array data[0] bl[0] br[0] data[1] bl[2] br[2] data[2] bl[4] br[4] data[3] bl[6] br[6] data[4] bl[8] br[8] data[5] bl[10] br[10] data[6] bl[12] br[12] data[7] bl[14] br[14] data[8] bl[16] br[16] data[9] bl[18] br[18] data[10] bl[20] br[20] data[11] bl[22] br[22] data[12] bl[24] br[24] data[13] bl[26] br[26] data[14] bl[28] br[28] data[15] bl[30] br[30] data[16] bl[32] br[32] data[17] bl[34] br[34] data[18] bl[36] br[36] data[19] bl[38] br[38] data[20] bl[40] br[40] data[21] bl[42] br[42] data[22] bl[44] br[44] data[23] bl[46] br[46] data[24] bl[48] br[48] data[25] bl[50] br[50] data[26] bl[52] br[52] data[27] bl[54] br[54] data[28] bl[56] br[56] data[29] bl[58] br[58] data[30] bl[60] br[60] data[31] bl[62] br[62] data[32] bl[64] br[64] data[33] bl[66] br[66] data[34] bl[68] br[68] data[35] bl[70] br[70] data[36] bl[72] br[72] data[37] bl[74] br[74] data[38] bl[76] br[76] data[39] bl[78] br[78] data[40] bl[80] br[80] data[41] bl[82] br[82] data[42] bl[84] br[84] data[43] bl[86] br[86] data[44] bl[88] br[88] data[45] bl[90] br[90] data[46] bl[92] br[92] data[47] bl[94] br[94] data[48] bl[96] br[96] data[49] bl[98] br[98] data[50] bl[100] br[100] data[51] bl[102] br[102] data[52] bl[104] br[104] data[53] bl[106] br[106] data[54] bl[108] br[108] data[55] bl[110] br[110] data[56] bl[112] br[112] data[57] bl[114] br[114] data[58] bl[116] br[116] data[59] bl[118] br[118] data[60] bl[120] br[120] data[61] bl[122] br[122] data[62] bl[124] br[124] data[63] bl[126] br[126] data[64] bl[128] br[128] data[65] bl[130] br[130] data[66] bl[132] br[132] data[67] bl[134] br[134] data[68] bl[136] br[136] data[69] bl[138] br[138] data[70] bl[140] br[140] data[71] bl[142] br[142] data[72] bl[144] br[144] data[73] bl[146] br[146] data[74] bl[148] br[148] data[75] bl[150] br[150] data[76] bl[152] br[152] data[77] bl[154] br[154] data[78] bl[156] br[156] data[79] bl[158] br[158] data[80] bl[160] br[160] data[81] bl[162] br[162] data[82] bl[164] br[164] data[83] bl[166] br[166] data[84] bl[168] br[168] data[85] bl[170] br[170] data[86] bl[172] br[172] data[87] bl[174] br[174] data[88] bl[176] br[176] data[89] bl[178] br[178] data[90] bl[180] br[180] data[91] bl[182] br[182] data[92] bl[184] br[184] data[93] bl[186] br[186] data[94] bl[188] br[188] data[95] bl[190] br[190] data[96] bl[192] br[192] data[97] bl[194] br[194] data[98] bl[196] br[196] data[99] bl[198] br[198] data[100] bl[200] br[200] data[101] bl[202] br[202] data[102] bl[204] br[204] data[103] bl[206] br[206] data[104] bl[208] br[208] data[105] bl[210] br[210] data[106] bl[212] br[212] data[107] bl[214] br[214] data[108] bl[216] br[216] data[109] bl[218] br[218] data[110] bl[220] br[220] data[111] bl[222] br[222] data[112] bl[224] br[224] data[113] bl[226] br[226] data[114] bl[228] br[228] data[115] bl[230] br[230] data[116] bl[232] br[232] data[117] bl[234] br[234] data[118] bl[236] br[236] data[119] bl[238] br[238] data[120] bl[240] br[240] data[121] bl[242] br[242] data[122] bl[244] br[244] data[123] bl[246] br[246] data[124] bl[248] br[248] data[125] bl[250] br[250] data[126] bl[252] br[252] data[127] bl[254] br[254] en vdd gnd
Xsa_d0 bl[0] br[0] data[0] en vdd gnd sense_amp
Xsa_d2 bl[2] br[2] data[1] en vdd gnd sense_amp
Xsa_d4 bl[4] br[4] data[2] en vdd gnd sense_amp
Xsa_d6 bl[6] br[6] data[3] en vdd gnd sense_amp
Xsa_d8 bl[8] br[8] data[4] en vdd gnd sense_amp
Xsa_d10 bl[10] br[10] data[5] en vdd gnd sense_amp
Xsa_d12 bl[12] br[12] data[6] en vdd gnd sense_amp
Xsa_d14 bl[14] br[14] data[7] en vdd gnd sense_amp
Xsa_d16 bl[16] br[16] data[8] en vdd gnd sense_amp
Xsa_d18 bl[18] br[18] data[9] en vdd gnd sense_amp
Xsa_d20 bl[20] br[20] data[10] en vdd gnd sense_amp
Xsa_d22 bl[22] br[22] data[11] en vdd gnd sense_amp
Xsa_d24 bl[24] br[24] data[12] en vdd gnd sense_amp
Xsa_d26 bl[26] br[26] data[13] en vdd gnd sense_amp
Xsa_d28 bl[28] br[28] data[14] en vdd gnd sense_amp
Xsa_d30 bl[30] br[30] data[15] en vdd gnd sense_amp
Xsa_d32 bl[32] br[32] data[16] en vdd gnd sense_amp
Xsa_d34 bl[34] br[34] data[17] en vdd gnd sense_amp
Xsa_d36 bl[36] br[36] data[18] en vdd gnd sense_amp
Xsa_d38 bl[38] br[38] data[19] en vdd gnd sense_amp
Xsa_d40 bl[40] br[40] data[20] en vdd gnd sense_amp
Xsa_d42 bl[42] br[42] data[21] en vdd gnd sense_amp
Xsa_d44 bl[44] br[44] data[22] en vdd gnd sense_amp
Xsa_d46 bl[46] br[46] data[23] en vdd gnd sense_amp
Xsa_d48 bl[48] br[48] data[24] en vdd gnd sense_amp
Xsa_d50 bl[50] br[50] data[25] en vdd gnd sense_amp
Xsa_d52 bl[52] br[52] data[26] en vdd gnd sense_amp
Xsa_d54 bl[54] br[54] data[27] en vdd gnd sense_amp
Xsa_d56 bl[56] br[56] data[28] en vdd gnd sense_amp
Xsa_d58 bl[58] br[58] data[29] en vdd gnd sense_amp
Xsa_d60 bl[60] br[60] data[30] en vdd gnd sense_amp
Xsa_d62 bl[62] br[62] data[31] en vdd gnd sense_amp
Xsa_d64 bl[64] br[64] data[32] en vdd gnd sense_amp
Xsa_d66 bl[66] br[66] data[33] en vdd gnd sense_amp
Xsa_d68 bl[68] br[68] data[34] en vdd gnd sense_amp
Xsa_d70 bl[70] br[70] data[35] en vdd gnd sense_amp
Xsa_d72 bl[72] br[72] data[36] en vdd gnd sense_amp
Xsa_d74 bl[74] br[74] data[37] en vdd gnd sense_amp
Xsa_d76 bl[76] br[76] data[38] en vdd gnd sense_amp
Xsa_d78 bl[78] br[78] data[39] en vdd gnd sense_amp
Xsa_d80 bl[80] br[80] data[40] en vdd gnd sense_amp
Xsa_d82 bl[82] br[82] data[41] en vdd gnd sense_amp
Xsa_d84 bl[84] br[84] data[42] en vdd gnd sense_amp
Xsa_d86 bl[86] br[86] data[43] en vdd gnd sense_amp
Xsa_d88 bl[88] br[88] data[44] en vdd gnd sense_amp
Xsa_d90 bl[90] br[90] data[45] en vdd gnd sense_amp
Xsa_d92 bl[92] br[92] data[46] en vdd gnd sense_amp
Xsa_d94 bl[94] br[94] data[47] en vdd gnd sense_amp
Xsa_d96 bl[96] br[96] data[48] en vdd gnd sense_amp
Xsa_d98 bl[98] br[98] data[49] en vdd gnd sense_amp
Xsa_d100 bl[100] br[100] data[50] en vdd gnd sense_amp
Xsa_d102 bl[102] br[102] data[51] en vdd gnd sense_amp
Xsa_d104 bl[104] br[104] data[52] en vdd gnd sense_amp
Xsa_d106 bl[106] br[106] data[53] en vdd gnd sense_amp
Xsa_d108 bl[108] br[108] data[54] en vdd gnd sense_amp
Xsa_d110 bl[110] br[110] data[55] en vdd gnd sense_amp
Xsa_d112 bl[112] br[112] data[56] en vdd gnd sense_amp
Xsa_d114 bl[114] br[114] data[57] en vdd gnd sense_amp
Xsa_d116 bl[116] br[116] data[58] en vdd gnd sense_amp
Xsa_d118 bl[118] br[118] data[59] en vdd gnd sense_amp
Xsa_d120 bl[120] br[120] data[60] en vdd gnd sense_amp
Xsa_d122 bl[122] br[122] data[61] en vdd gnd sense_amp
Xsa_d124 bl[124] br[124] data[62] en vdd gnd sense_amp
Xsa_d126 bl[126] br[126] data[63] en vdd gnd sense_amp
Xsa_d128 bl[128] br[128] data[64] en vdd gnd sense_amp
Xsa_d130 bl[130] br[130] data[65] en vdd gnd sense_amp
Xsa_d132 bl[132] br[132] data[66] en vdd gnd sense_amp
Xsa_d134 bl[134] br[134] data[67] en vdd gnd sense_amp
Xsa_d136 bl[136] br[136] data[68] en vdd gnd sense_amp
Xsa_d138 bl[138] br[138] data[69] en vdd gnd sense_amp
Xsa_d140 bl[140] br[140] data[70] en vdd gnd sense_amp
Xsa_d142 bl[142] br[142] data[71] en vdd gnd sense_amp
Xsa_d144 bl[144] br[144] data[72] en vdd gnd sense_amp
Xsa_d146 bl[146] br[146] data[73] en vdd gnd sense_amp
Xsa_d148 bl[148] br[148] data[74] en vdd gnd sense_amp
Xsa_d150 bl[150] br[150] data[75] en vdd gnd sense_amp
Xsa_d152 bl[152] br[152] data[76] en vdd gnd sense_amp
Xsa_d154 bl[154] br[154] data[77] en vdd gnd sense_amp
Xsa_d156 bl[156] br[156] data[78] en vdd gnd sense_amp
Xsa_d158 bl[158] br[158] data[79] en vdd gnd sense_amp
Xsa_d160 bl[160] br[160] data[80] en vdd gnd sense_amp
Xsa_d162 bl[162] br[162] data[81] en vdd gnd sense_amp
Xsa_d164 bl[164] br[164] data[82] en vdd gnd sense_amp
Xsa_d166 bl[166] br[166] data[83] en vdd gnd sense_amp
Xsa_d168 bl[168] br[168] data[84] en vdd gnd sense_amp
Xsa_d170 bl[170] br[170] data[85] en vdd gnd sense_amp
Xsa_d172 bl[172] br[172] data[86] en vdd gnd sense_amp
Xsa_d174 bl[174] br[174] data[87] en vdd gnd sense_amp
Xsa_d176 bl[176] br[176] data[88] en vdd gnd sense_amp
Xsa_d178 bl[178] br[178] data[89] en vdd gnd sense_amp
Xsa_d180 bl[180] br[180] data[90] en vdd gnd sense_amp
Xsa_d182 bl[182] br[182] data[91] en vdd gnd sense_amp
Xsa_d184 bl[184] br[184] data[92] en vdd gnd sense_amp
Xsa_d186 bl[186] br[186] data[93] en vdd gnd sense_amp
Xsa_d188 bl[188] br[188] data[94] en vdd gnd sense_amp
Xsa_d190 bl[190] br[190] data[95] en vdd gnd sense_amp
Xsa_d192 bl[192] br[192] data[96] en vdd gnd sense_amp
Xsa_d194 bl[194] br[194] data[97] en vdd gnd sense_amp
Xsa_d196 bl[196] br[196] data[98] en vdd gnd sense_amp
Xsa_d198 bl[198] br[198] data[99] en vdd gnd sense_amp
Xsa_d200 bl[200] br[200] data[100] en vdd gnd sense_amp
Xsa_d202 bl[202] br[202] data[101] en vdd gnd sense_amp
Xsa_d204 bl[204] br[204] data[102] en vdd gnd sense_amp
Xsa_d206 bl[206] br[206] data[103] en vdd gnd sense_amp
Xsa_d208 bl[208] br[208] data[104] en vdd gnd sense_amp
Xsa_d210 bl[210] br[210] data[105] en vdd gnd sense_amp
Xsa_d212 bl[212] br[212] data[106] en vdd gnd sense_amp
Xsa_d214 bl[214] br[214] data[107] en vdd gnd sense_amp
Xsa_d216 bl[216] br[216] data[108] en vdd gnd sense_amp
Xsa_d218 bl[218] br[218] data[109] en vdd gnd sense_amp
Xsa_d220 bl[220] br[220] data[110] en vdd gnd sense_amp
Xsa_d222 bl[222] br[222] data[111] en vdd gnd sense_amp
Xsa_d224 bl[224] br[224] data[112] en vdd gnd sense_amp
Xsa_d226 bl[226] br[226] data[113] en vdd gnd sense_amp
Xsa_d228 bl[228] br[228] data[114] en vdd gnd sense_amp
Xsa_d230 bl[230] br[230] data[115] en vdd gnd sense_amp
Xsa_d232 bl[232] br[232] data[116] en vdd gnd sense_amp
Xsa_d234 bl[234] br[234] data[117] en vdd gnd sense_amp
Xsa_d236 bl[236] br[236] data[118] en vdd gnd sense_amp
Xsa_d238 bl[238] br[238] data[119] en vdd gnd sense_amp
Xsa_d240 bl[240] br[240] data[120] en vdd gnd sense_amp
Xsa_d242 bl[242] br[242] data[121] en vdd gnd sense_amp
Xsa_d244 bl[244] br[244] data[122] en vdd gnd sense_amp
Xsa_d246 bl[246] br[246] data[123] en vdd gnd sense_amp
Xsa_d248 bl[248] br[248] data[124] en vdd gnd sense_amp
Xsa_d250 bl[250] br[250] data[125] en vdd gnd sense_amp
Xsa_d252 bl[252] br[252] data[126] en vdd gnd sense_amp
Xsa_d254 bl[254] br[254] data[127] en vdd gnd sense_amp
.ENDS sense_amp_array
*********************** Write_Driver ******************************
.SUBCKT write_driver din bl br en vdd gnd

**** Inverter to conver Data_in to data_in_bar ******
M_1 net_3 din gnd gnd n W='1.2*1u' L=0.6u
M_2 net_3 din vdd vdd p W='2.1*1u' L=0.6u

**** 2input nand gate follwed by inverter to drive BL ******
M_3 net_2 en net_7 gnd n W='2.1*1u' L=0.6u
M_4 net_7 din gnd gnd n W='2.1*1u' L=0.6u
M_5 net_2 en vdd vdd p W='2.1*1u' L=0.6u
M_6 net_2 din vdd vdd p W='2.1*1u' L=0.6u


M_7 net_1 net_2 vdd vdd p W='2.1*1u' L=0.6u
M_8 net_1 net_2 gnd gnd n W='1.2*1u' L=0.6u

**** 2input nand gate follwed by inverter to drive BR******

M_9 net_4 en vdd vdd p W='2.1*1u' L=0.6u
M_10 net_4 en net_8 gnd n W='2.1*1u' L=0.6u
M_11 net_8 net_3 gnd gnd n W='2.1*1u' L=0.6u
M_12 net_4 net_3 vdd vdd p W='2.1*1u' L=0.6u

M_13 net_6 net_4 vdd vdd p W='2.1*1u' L=0.6u
M_14 net_6 net_4 gnd gnd n W='1.2*1u' L=0.6u

************************************************

M_15 bl net_6 net_5 gnd n W='3.6*1u' L=0.6u
M_16 br net_1 net_5 gnd n W='3.6*1u' L=0.6u
M_17 net_5 en gnd gnd n W='3.6*1u' L=0.6u



.ENDS	$ write_driver


.SUBCKT write_driver_array data[0] data[1] data[2] data[3] data[4] data[5] data[6] data[7] data[8] data[9] data[10] data[11] data[12] data[13] data[14] data[15] data[16] data[17] data[18] data[19] data[20] data[21] data[22] data[23] data[24] data[25] data[26] data[27] data[28] data[29] data[30] data[31] data[32] data[33] data[34] data[35] data[36] data[37] data[38] data[39] data[40] data[41] data[42] data[43] data[44] data[45] data[46] data[47] data[48] data[49] data[50] data[51] data[52] data[53] data[54] data[55] data[56] data[57] data[58] data[59] data[60] data[61] data[62] data[63] data[64] data[65] data[66] data[67] data[68] data[69] data[70] data[71] data[72] data[73] data[74] data[75] data[76] data[77] data[78] data[79] data[80] data[81] data[82] data[83] data[84] data[85] data[86] data[87] data[88] data[89] data[90] data[91] data[92] data[93] data[94] data[95] data[96] data[97] data[98] data[99] data[100] data[101] data[102] data[103] data[104] data[105] data[106] data[107] data[108] data[109] data[110] data[111] data[112] data[113] data[114] data[115] data[116] data[117] data[118] data[119] data[120] data[121] data[122] data[123] data[124] data[125] data[126] data[127] bl[0] br[0] bl[1] br[1] bl[2] br[2] bl[3] br[3] bl[4] br[4] bl[5] br[5] bl[6] br[6] bl[7] br[7] bl[8] br[8] bl[9] br[9] bl[10] br[10] bl[11] br[11] bl[12] br[12] bl[13] br[13] bl[14] br[14] bl[15] br[15] bl[16] br[16] bl[17] br[17] bl[18] br[18] bl[19] br[19] bl[20] br[20] bl[21] br[21] bl[22] br[22] bl[23] br[23] bl[24] br[24] bl[25] br[25] bl[26] br[26] bl[27] br[27] bl[28] br[28] bl[29] br[29] bl[30] br[30] bl[31] br[31] bl[32] br[32] bl[33] br[33] bl[34] br[34] bl[35] br[35] bl[36] br[36] bl[37] br[37] bl[38] br[38] bl[39] br[39] bl[40] br[40] bl[41] br[41] bl[42] br[42] bl[43] br[43] bl[44] br[44] bl[45] br[45] bl[46] br[46] bl[47] br[47] bl[48] br[48] bl[49] br[49] bl[50] br[50] bl[51] br[51] bl[52] br[52] bl[53] br[53] bl[54] br[54] bl[55] br[55] bl[56] br[56] bl[57] br[57] bl[58] br[58] bl[59] br[59] bl[60] br[60] bl[61] br[61] bl[62] br[62] bl[63] br[63] bl[64] br[64] bl[65] br[65] bl[66] br[66] bl[67] br[67] bl[68] br[68] bl[69] br[69] bl[70] br[70] bl[71] br[71] bl[72] br[72] bl[73] br[73] bl[74] br[74] bl[75] br[75] bl[76] br[76] bl[77] br[77] bl[78] br[78] bl[79] br[79] bl[80] br[80] bl[81] br[81] bl[82] br[82] bl[83] br[83] bl[84] br[84] bl[85] br[85] bl[86] br[86] bl[87] br[87] bl[88] br[88] bl[89] br[89] bl[90] br[90] bl[91] br[91] bl[92] br[92] bl[93] br[93] bl[94] br[94] bl[95] br[95] bl[96] br[96] bl[97] br[97] bl[98] br[98] bl[99] br[99] bl[100] br[100] bl[101] br[101] bl[102] br[102] bl[103] br[103] bl[104] br[104] bl[105] br[105] bl[106] br[106] bl[107] br[107] bl[108] br[108] bl[109] br[109] bl[110] br[110] bl[111] br[111] bl[112] br[112] bl[113] br[113] bl[114] br[114] bl[115] br[115] bl[116] br[116] bl[117] br[117] bl[118] br[118] bl[119] br[119] bl[120] br[120] bl[121] br[121] bl[122] br[122] bl[123] br[123] bl[124] br[124] bl[125] br[125] bl[126] br[126] bl[127] br[127] en vdd gnd
XXwrite_driver0 data[0] bl[0] br[0] en vdd gnd write_driver
XXwrite_driver2 data[1] bl[1] br[1] en vdd gnd write_driver
XXwrite_driver4 data[2] bl[2] br[2] en vdd gnd write_driver
XXwrite_driver6 data[3] bl[3] br[3] en vdd gnd write_driver
XXwrite_driver8 data[4] bl[4] br[4] en vdd gnd write_driver
XXwrite_driver10 data[5] bl[5] br[5] en vdd gnd write_driver
XXwrite_driver12 data[6] bl[6] br[6] en vdd gnd write_driver
XXwrite_driver14 data[7] bl[7] br[7] en vdd gnd write_driver
XXwrite_driver16 data[8] bl[8] br[8] en vdd gnd write_driver
XXwrite_driver18 data[9] bl[9] br[9] en vdd gnd write_driver
XXwrite_driver20 data[10] bl[10] br[10] en vdd gnd write_driver
XXwrite_driver22 data[11] bl[11] br[11] en vdd gnd write_driver
XXwrite_driver24 data[12] bl[12] br[12] en vdd gnd write_driver
XXwrite_driver26 data[13] bl[13] br[13] en vdd gnd write_driver
XXwrite_driver28 data[14] bl[14] br[14] en vdd gnd write_driver
XXwrite_driver30 data[15] bl[15] br[15] en vdd gnd write_driver
XXwrite_driver32 data[16] bl[16] br[16] en vdd gnd write_driver
XXwrite_driver34 data[17] bl[17] br[17] en vdd gnd write_driver
XXwrite_driver36 data[18] bl[18] br[18] en vdd gnd write_driver
XXwrite_driver38 data[19] bl[19] br[19] en vdd gnd write_driver
XXwrite_driver40 data[20] bl[20] br[20] en vdd gnd write_driver
XXwrite_driver42 data[21] bl[21] br[21] en vdd gnd write_driver
XXwrite_driver44 data[22] bl[22] br[22] en vdd gnd write_driver
XXwrite_driver46 data[23] bl[23] br[23] en vdd gnd write_driver
XXwrite_driver48 data[24] bl[24] br[24] en vdd gnd write_driver
XXwrite_driver50 data[25] bl[25] br[25] en vdd gnd write_driver
XXwrite_driver52 data[26] bl[26] br[26] en vdd gnd write_driver
XXwrite_driver54 data[27] bl[27] br[27] en vdd gnd write_driver
XXwrite_driver56 data[28] bl[28] br[28] en vdd gnd write_driver
XXwrite_driver58 data[29] bl[29] br[29] en vdd gnd write_driver
XXwrite_driver60 data[30] bl[30] br[30] en vdd gnd write_driver
XXwrite_driver62 data[31] bl[31] br[31] en vdd gnd write_driver
XXwrite_driver64 data[32] bl[32] br[32] en vdd gnd write_driver
XXwrite_driver66 data[33] bl[33] br[33] en vdd gnd write_driver
XXwrite_driver68 data[34] bl[34] br[34] en vdd gnd write_driver
XXwrite_driver70 data[35] bl[35] br[35] en vdd gnd write_driver
XXwrite_driver72 data[36] bl[36] br[36] en vdd gnd write_driver
XXwrite_driver74 data[37] bl[37] br[37] en vdd gnd write_driver
XXwrite_driver76 data[38] bl[38] br[38] en vdd gnd write_driver
XXwrite_driver78 data[39] bl[39] br[39] en vdd gnd write_driver
XXwrite_driver80 data[40] bl[40] br[40] en vdd gnd write_driver
XXwrite_driver82 data[41] bl[41] br[41] en vdd gnd write_driver
XXwrite_driver84 data[42] bl[42] br[42] en vdd gnd write_driver
XXwrite_driver86 data[43] bl[43] br[43] en vdd gnd write_driver
XXwrite_driver88 data[44] bl[44] br[44] en vdd gnd write_driver
XXwrite_driver90 data[45] bl[45] br[45] en vdd gnd write_driver
XXwrite_driver92 data[46] bl[46] br[46] en vdd gnd write_driver
XXwrite_driver94 data[47] bl[47] br[47] en vdd gnd write_driver
XXwrite_driver96 data[48] bl[48] br[48] en vdd gnd write_driver
XXwrite_driver98 data[49] bl[49] br[49] en vdd gnd write_driver
XXwrite_driver100 data[50] bl[50] br[50] en vdd gnd write_driver
XXwrite_driver102 data[51] bl[51] br[51] en vdd gnd write_driver
XXwrite_driver104 data[52] bl[52] br[52] en vdd gnd write_driver
XXwrite_driver106 data[53] bl[53] br[53] en vdd gnd write_driver
XXwrite_driver108 data[54] bl[54] br[54] en vdd gnd write_driver
XXwrite_driver110 data[55] bl[55] br[55] en vdd gnd write_driver
XXwrite_driver112 data[56] bl[56] br[56] en vdd gnd write_driver
XXwrite_driver114 data[57] bl[57] br[57] en vdd gnd write_driver
XXwrite_driver116 data[58] bl[58] br[58] en vdd gnd write_driver
XXwrite_driver118 data[59] bl[59] br[59] en vdd gnd write_driver
XXwrite_driver120 data[60] bl[60] br[60] en vdd gnd write_driver
XXwrite_driver122 data[61] bl[61] br[61] en vdd gnd write_driver
XXwrite_driver124 data[62] bl[62] br[62] en vdd gnd write_driver
XXwrite_driver126 data[63] bl[63] br[63] en vdd gnd write_driver
XXwrite_driver128 data[64] bl[64] br[64] en vdd gnd write_driver
XXwrite_driver130 data[65] bl[65] br[65] en vdd gnd write_driver
XXwrite_driver132 data[66] bl[66] br[66] en vdd gnd write_driver
XXwrite_driver134 data[67] bl[67] br[67] en vdd gnd write_driver
XXwrite_driver136 data[68] bl[68] br[68] en vdd gnd write_driver
XXwrite_driver138 data[69] bl[69] br[69] en vdd gnd write_driver
XXwrite_driver140 data[70] bl[70] br[70] en vdd gnd write_driver
XXwrite_driver142 data[71] bl[71] br[71] en vdd gnd write_driver
XXwrite_driver144 data[72] bl[72] br[72] en vdd gnd write_driver
XXwrite_driver146 data[73] bl[73] br[73] en vdd gnd write_driver
XXwrite_driver148 data[74] bl[74] br[74] en vdd gnd write_driver
XXwrite_driver150 data[75] bl[75] br[75] en vdd gnd write_driver
XXwrite_driver152 data[76] bl[76] br[76] en vdd gnd write_driver
XXwrite_driver154 data[77] bl[77] br[77] en vdd gnd write_driver
XXwrite_driver156 data[78] bl[78] br[78] en vdd gnd write_driver
XXwrite_driver158 data[79] bl[79] br[79] en vdd gnd write_driver
XXwrite_driver160 data[80] bl[80] br[80] en vdd gnd write_driver
XXwrite_driver162 data[81] bl[81] br[81] en vdd gnd write_driver
XXwrite_driver164 data[82] bl[82] br[82] en vdd gnd write_driver
XXwrite_driver166 data[83] bl[83] br[83] en vdd gnd write_driver
XXwrite_driver168 data[84] bl[84] br[84] en vdd gnd write_driver
XXwrite_driver170 data[85] bl[85] br[85] en vdd gnd write_driver
XXwrite_driver172 data[86] bl[86] br[86] en vdd gnd write_driver
XXwrite_driver174 data[87] bl[87] br[87] en vdd gnd write_driver
XXwrite_driver176 data[88] bl[88] br[88] en vdd gnd write_driver
XXwrite_driver178 data[89] bl[89] br[89] en vdd gnd write_driver
XXwrite_driver180 data[90] bl[90] br[90] en vdd gnd write_driver
XXwrite_driver182 data[91] bl[91] br[91] en vdd gnd write_driver
XXwrite_driver184 data[92] bl[92] br[92] en vdd gnd write_driver
XXwrite_driver186 data[93] bl[93] br[93] en vdd gnd write_driver
XXwrite_driver188 data[94] bl[94] br[94] en vdd gnd write_driver
XXwrite_driver190 data[95] bl[95] br[95] en vdd gnd write_driver
XXwrite_driver192 data[96] bl[96] br[96] en vdd gnd write_driver
XXwrite_driver194 data[97] bl[97] br[97] en vdd gnd write_driver
XXwrite_driver196 data[98] bl[98] br[98] en vdd gnd write_driver
XXwrite_driver198 data[99] bl[99] br[99] en vdd gnd write_driver
XXwrite_driver200 data[100] bl[100] br[100] en vdd gnd write_driver
XXwrite_driver202 data[101] bl[101] br[101] en vdd gnd write_driver
XXwrite_driver204 data[102] bl[102] br[102] en vdd gnd write_driver
XXwrite_driver206 data[103] bl[103] br[103] en vdd gnd write_driver
XXwrite_driver208 data[104] bl[104] br[104] en vdd gnd write_driver
XXwrite_driver210 data[105] bl[105] br[105] en vdd gnd write_driver
XXwrite_driver212 data[106] bl[106] br[106] en vdd gnd write_driver
XXwrite_driver214 data[107] bl[107] br[107] en vdd gnd write_driver
XXwrite_driver216 data[108] bl[108] br[108] en vdd gnd write_driver
XXwrite_driver218 data[109] bl[109] br[109] en vdd gnd write_driver
XXwrite_driver220 data[110] bl[110] br[110] en vdd gnd write_driver
XXwrite_driver222 data[111] bl[111] br[111] en vdd gnd write_driver
XXwrite_driver224 data[112] bl[112] br[112] en vdd gnd write_driver
XXwrite_driver226 data[113] bl[113] br[113] en vdd gnd write_driver
XXwrite_driver228 data[114] bl[114] br[114] en vdd gnd write_driver
XXwrite_driver230 data[115] bl[115] br[115] en vdd gnd write_driver
XXwrite_driver232 data[116] bl[116] br[116] en vdd gnd write_driver
XXwrite_driver234 data[117] bl[117] br[117] en vdd gnd write_driver
XXwrite_driver236 data[118] bl[118] br[118] en vdd gnd write_driver
XXwrite_driver238 data[119] bl[119] br[119] en vdd gnd write_driver
XXwrite_driver240 data[120] bl[120] br[120] en vdd gnd write_driver
XXwrite_driver242 data[121] bl[121] br[121] en vdd gnd write_driver
XXwrite_driver244 data[122] bl[122] br[122] en vdd gnd write_driver
XXwrite_driver246 data[123] bl[123] br[123] en vdd gnd write_driver
XXwrite_driver248 data[124] bl[124] br[124] en vdd gnd write_driver
XXwrite_driver250 data[125] bl[125] br[125] en vdd gnd write_driver
XXwrite_driver252 data[126] bl[126] br[126] en vdd gnd write_driver
XXwrite_driver254 data[127] bl[127] br[127] en vdd gnd write_driver
.ENDS write_driver_array

.SUBCKT pinv_8 A Z vdd gnd
Mpinv_pmos Z A vdd vdd p m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpinv_nmos Z A gnd gnd n m=1 w=1.2u l=0.6u pd=3.6u ps=3.6u as=1.8p ad=1.8p
.ENDS pinv_8

.SUBCKT pnand2_2 A B Z vdd gnd
Mpnand2_pmos1 vdd A Z vdd p m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpnand2_pmos2 Z B vdd vdd p m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpnand2_nmos1 Z B net1 gnd n m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpnand2_nmos2 net1 A gnd gnd n m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
.ENDS pnand2_2

.SUBCKT pnand3_2 A B C Z vdd gnd
Mpnand3_pmos1 vdd A Z vdd p m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpnand3_pmos2 Z B vdd vdd p m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpnand3_pmos3 Z C vdd vdd p m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpnand3_nmos1 Z C net1 gnd n m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpnand3_nmos2 net1 B net2 gnd n m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpnand3_nmos3 net2 A gnd gnd n m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
.ENDS pnand3_2

.SUBCKT pinv_9 A Z vdd gnd
Mpinv_pmos Z A vdd vdd p m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpinv_nmos Z A gnd gnd n m=1 w=1.2u l=0.6u pd=3.6u ps=3.6u as=1.8p ad=1.8p
.ENDS pinv_9

.SUBCKT pnand2_3 A B Z vdd gnd
Mpnand2_pmos1 vdd A Z vdd p m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpnand2_pmos2 Z B vdd vdd p m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpnand2_nmos1 Z B net1 gnd n m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpnand2_nmos2 net1 A gnd gnd n m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
.ENDS pnand2_3

.SUBCKT pre2x4 in[0] in[1] out[0] out[1] out[2] out[3] vdd gnd
XXpre_inv[0] in[0] inbar[0] vdd gnd pinv_9
XXpre_inv[1] in[1] inbar[1] vdd gnd pinv_9
XXpre_nand_inv[0] Z[0] out[0] vdd gnd pinv_9
XXpre_nand_inv[1] Z[1] out[1] vdd gnd pinv_9
XXpre_nand_inv[2] Z[2] out[2] vdd gnd pinv_9
XXpre_nand_inv[3] Z[3] out[3] vdd gnd pinv_9
XXpre2x4_nand[0] inbar[0] inbar[1] Z[0] vdd gnd pnand2_3
XXpre2x4_nand[1] in[0] inbar[1] Z[1] vdd gnd pnand2_3
XXpre2x4_nand[2] inbar[0] in[1] Z[2] vdd gnd pnand2_3
XXpre2x4_nand[3] in[0] in[1] Z[3] vdd gnd pnand2_3
.ENDS pre2x4

.SUBCKT pinv_10 A Z vdd gnd
Mpinv_pmos Z A vdd vdd p m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpinv_nmos Z A gnd gnd n m=1 w=1.2u l=0.6u pd=3.6u ps=3.6u as=1.8p ad=1.8p
.ENDS pinv_10

.SUBCKT pnand3_3 A B C Z vdd gnd
Mpnand3_pmos1 vdd A Z vdd p m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpnand3_pmos2 Z B vdd vdd p m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpnand3_pmos3 Z C vdd vdd p m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpnand3_nmos1 Z C net1 gnd n m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpnand3_nmos2 net1 B net2 gnd n m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpnand3_nmos3 net2 A gnd gnd n m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
.ENDS pnand3_3

.SUBCKT pre3x8 in[0] in[1] in[2] out[0] out[1] out[2] out[3] out[4] out[5] out[6] out[7] vdd gnd
XXpre_inv[0] in[0] inbar[0] vdd gnd pinv_10
XXpre_inv[1] in[1] inbar[1] vdd gnd pinv_10
XXpre_inv[2] in[2] inbar[2] vdd gnd pinv_10
XXpre_nand_inv[0] Z[0] out[0] vdd gnd pinv_10
XXpre_nand_inv[1] Z[1] out[1] vdd gnd pinv_10
XXpre_nand_inv[2] Z[2] out[2] vdd gnd pinv_10
XXpre_nand_inv[3] Z[3] out[3] vdd gnd pinv_10
XXpre_nand_inv[4] Z[4] out[4] vdd gnd pinv_10
XXpre_nand_inv[5] Z[5] out[5] vdd gnd pinv_10
XXpre_nand_inv[6] Z[6] out[6] vdd gnd pinv_10
XXpre_nand_inv[7] Z[7] out[7] vdd gnd pinv_10
XXpre3x8_nand[0] inbar[0] inbar[1] inbar[2] Z[0] vdd gnd pnand3_3
XXpre3x8_nand[1] in[0] inbar[1] inbar[2] Z[1] vdd gnd pnand3_3
XXpre3x8_nand[2] inbar[0] in[1] inbar[2] Z[2] vdd gnd pnand3_3
XXpre3x8_nand[3] in[0] in[1] inbar[2] Z[3] vdd gnd pnand3_3
XXpre3x8_nand[4] inbar[0] inbar[1] in[2] Z[4] vdd gnd pnand3_3
XXpre3x8_nand[5] in[0] inbar[1] in[2] Z[5] vdd gnd pnand3_3
XXpre3x8_nand[6] inbar[0] in[1] in[2] Z[6] vdd gnd pnand3_3
XXpre3x8_nand[7] in[0] in[1] in[2] Z[7] vdd gnd pnand3_3
.ENDS pre3x8

.SUBCKT hierarchical_decoder_128rows A[0] A[1] A[2] A[3] A[4] A[5] A[6] decode[0] decode[1] decode[2] decode[3] decode[4] decode[5] decode[6] decode[7] decode[8] decode[9] decode[10] decode[11] decode[12] decode[13] decode[14] decode[15] decode[16] decode[17] decode[18] decode[19] decode[20] decode[21] decode[22] decode[23] decode[24] decode[25] decode[26] decode[27] decode[28] decode[29] decode[30] decode[31] decode[32] decode[33] decode[34] decode[35] decode[36] decode[37] decode[38] decode[39] decode[40] decode[41] decode[42] decode[43] decode[44] decode[45] decode[46] decode[47] decode[48] decode[49] decode[50] decode[51] decode[52] decode[53] decode[54] decode[55] decode[56] decode[57] decode[58] decode[59] decode[60] decode[61] decode[62] decode[63] decode[64] decode[65] decode[66] decode[67] decode[68] decode[69] decode[70] decode[71] decode[72] decode[73] decode[74] decode[75] decode[76] decode[77] decode[78] decode[79] decode[80] decode[81] decode[82] decode[83] decode[84] decode[85] decode[86] decode[87] decode[88] decode[89] decode[90] decode[91] decode[92] decode[93] decode[94] decode[95] decode[96] decode[97] decode[98] decode[99] decode[100] decode[101] decode[102] decode[103] decode[104] decode[105] decode[106] decode[107] decode[108] decode[109] decode[110] decode[111] decode[112] decode[113] decode[114] decode[115] decode[116] decode[117] decode[118] decode[119] decode[120] decode[121] decode[122] decode[123] decode[124] decode[125] decode[126] decode[127] vdd gnd
Xpre[0] A[0] A[1] out[0] out[1] out[2] out[3] vdd gnd pre2x4
Xpre[1] A[2] A[3] out[4] out[5] out[6] out[7] vdd gnd pre2x4
Xpre3x8[0] A[4] A[5] A[6] out[8] out[9] out[10] out[11] out[12] out[13] out[14] out[15] vdd gnd pre3x8
XDEC_NAND[0] out[0] out[4] out[8] Z[0] vdd gnd pnand3_2
XDEC_NAND[1] out[0] out[4] out[9] Z[1] vdd gnd pnand3_2
XDEC_NAND[2] out[0] out[4] out[10] Z[2] vdd gnd pnand3_2
XDEC_NAND[3] out[0] out[4] out[11] Z[3] vdd gnd pnand3_2
XDEC_NAND[4] out[0] out[4] out[12] Z[4] vdd gnd pnand3_2
XDEC_NAND[5] out[0] out[4] out[13] Z[5] vdd gnd pnand3_2
XDEC_NAND[6] out[0] out[4] out[14] Z[6] vdd gnd pnand3_2
XDEC_NAND[7] out[0] out[4] out[15] Z[7] vdd gnd pnand3_2
XDEC_NAND[8] out[0] out[5] out[8] Z[8] vdd gnd pnand3_2
XDEC_NAND[9] out[0] out[5] out[9] Z[9] vdd gnd pnand3_2
XDEC_NAND[10] out[0] out[5] out[10] Z[10] vdd gnd pnand3_2
XDEC_NAND[11] out[0] out[5] out[11] Z[11] vdd gnd pnand3_2
XDEC_NAND[12] out[0] out[5] out[12] Z[12] vdd gnd pnand3_2
XDEC_NAND[13] out[0] out[5] out[13] Z[13] vdd gnd pnand3_2
XDEC_NAND[14] out[0] out[5] out[14] Z[14] vdd gnd pnand3_2
XDEC_NAND[15] out[0] out[5] out[15] Z[15] vdd gnd pnand3_2
XDEC_NAND[16] out[0] out[6] out[8] Z[16] vdd gnd pnand3_2
XDEC_NAND[17] out[0] out[6] out[9] Z[17] vdd gnd pnand3_2
XDEC_NAND[18] out[0] out[6] out[10] Z[18] vdd gnd pnand3_2
XDEC_NAND[19] out[0] out[6] out[11] Z[19] vdd gnd pnand3_2
XDEC_NAND[20] out[0] out[6] out[12] Z[20] vdd gnd pnand3_2
XDEC_NAND[21] out[0] out[6] out[13] Z[21] vdd gnd pnand3_2
XDEC_NAND[22] out[0] out[6] out[14] Z[22] vdd gnd pnand3_2
XDEC_NAND[23] out[0] out[6] out[15] Z[23] vdd gnd pnand3_2
XDEC_NAND[24] out[0] out[7] out[8] Z[24] vdd gnd pnand3_2
XDEC_NAND[25] out[0] out[7] out[9] Z[25] vdd gnd pnand3_2
XDEC_NAND[26] out[0] out[7] out[10] Z[26] vdd gnd pnand3_2
XDEC_NAND[27] out[0] out[7] out[11] Z[27] vdd gnd pnand3_2
XDEC_NAND[28] out[0] out[7] out[12] Z[28] vdd gnd pnand3_2
XDEC_NAND[29] out[0] out[7] out[13] Z[29] vdd gnd pnand3_2
XDEC_NAND[30] out[0] out[7] out[14] Z[30] vdd gnd pnand3_2
XDEC_NAND[31] out[0] out[7] out[15] Z[31] vdd gnd pnand3_2
XDEC_NAND[32] out[1] out[4] out[8] Z[32] vdd gnd pnand3_2
XDEC_NAND[33] out[1] out[4] out[9] Z[33] vdd gnd pnand3_2
XDEC_NAND[34] out[1] out[4] out[10] Z[34] vdd gnd pnand3_2
XDEC_NAND[35] out[1] out[4] out[11] Z[35] vdd gnd pnand3_2
XDEC_NAND[36] out[1] out[4] out[12] Z[36] vdd gnd pnand3_2
XDEC_NAND[37] out[1] out[4] out[13] Z[37] vdd gnd pnand3_2
XDEC_NAND[38] out[1] out[4] out[14] Z[38] vdd gnd pnand3_2
XDEC_NAND[39] out[1] out[4] out[15] Z[39] vdd gnd pnand3_2
XDEC_NAND[40] out[1] out[5] out[8] Z[40] vdd gnd pnand3_2
XDEC_NAND[41] out[1] out[5] out[9] Z[41] vdd gnd pnand3_2
XDEC_NAND[42] out[1] out[5] out[10] Z[42] vdd gnd pnand3_2
XDEC_NAND[43] out[1] out[5] out[11] Z[43] vdd gnd pnand3_2
XDEC_NAND[44] out[1] out[5] out[12] Z[44] vdd gnd pnand3_2
XDEC_NAND[45] out[1] out[5] out[13] Z[45] vdd gnd pnand3_2
XDEC_NAND[46] out[1] out[5] out[14] Z[46] vdd gnd pnand3_2
XDEC_NAND[47] out[1] out[5] out[15] Z[47] vdd gnd pnand3_2
XDEC_NAND[48] out[1] out[6] out[8] Z[48] vdd gnd pnand3_2
XDEC_NAND[49] out[1] out[6] out[9] Z[49] vdd gnd pnand3_2
XDEC_NAND[50] out[1] out[6] out[10] Z[50] vdd gnd pnand3_2
XDEC_NAND[51] out[1] out[6] out[11] Z[51] vdd gnd pnand3_2
XDEC_NAND[52] out[1] out[6] out[12] Z[52] vdd gnd pnand3_2
XDEC_NAND[53] out[1] out[6] out[13] Z[53] vdd gnd pnand3_2
XDEC_NAND[54] out[1] out[6] out[14] Z[54] vdd gnd pnand3_2
XDEC_NAND[55] out[1] out[6] out[15] Z[55] vdd gnd pnand3_2
XDEC_NAND[56] out[1] out[7] out[8] Z[56] vdd gnd pnand3_2
XDEC_NAND[57] out[1] out[7] out[9] Z[57] vdd gnd pnand3_2
XDEC_NAND[58] out[1] out[7] out[10] Z[58] vdd gnd pnand3_2
XDEC_NAND[59] out[1] out[7] out[11] Z[59] vdd gnd pnand3_2
XDEC_NAND[60] out[1] out[7] out[12] Z[60] vdd gnd pnand3_2
XDEC_NAND[61] out[1] out[7] out[13] Z[61] vdd gnd pnand3_2
XDEC_NAND[62] out[1] out[7] out[14] Z[62] vdd gnd pnand3_2
XDEC_NAND[63] out[1] out[7] out[15] Z[63] vdd gnd pnand3_2
XDEC_NAND[64] out[2] out[4] out[8] Z[64] vdd gnd pnand3_2
XDEC_NAND[65] out[2] out[4] out[9] Z[65] vdd gnd pnand3_2
XDEC_NAND[66] out[2] out[4] out[10] Z[66] vdd gnd pnand3_2
XDEC_NAND[67] out[2] out[4] out[11] Z[67] vdd gnd pnand3_2
XDEC_NAND[68] out[2] out[4] out[12] Z[68] vdd gnd pnand3_2
XDEC_NAND[69] out[2] out[4] out[13] Z[69] vdd gnd pnand3_2
XDEC_NAND[70] out[2] out[4] out[14] Z[70] vdd gnd pnand3_2
XDEC_NAND[71] out[2] out[4] out[15] Z[71] vdd gnd pnand3_2
XDEC_NAND[72] out[2] out[5] out[8] Z[72] vdd gnd pnand3_2
XDEC_NAND[73] out[2] out[5] out[9] Z[73] vdd gnd pnand3_2
XDEC_NAND[74] out[2] out[5] out[10] Z[74] vdd gnd pnand3_2
XDEC_NAND[75] out[2] out[5] out[11] Z[75] vdd gnd pnand3_2
XDEC_NAND[76] out[2] out[5] out[12] Z[76] vdd gnd pnand3_2
XDEC_NAND[77] out[2] out[5] out[13] Z[77] vdd gnd pnand3_2
XDEC_NAND[78] out[2] out[5] out[14] Z[78] vdd gnd pnand3_2
XDEC_NAND[79] out[2] out[5] out[15] Z[79] vdd gnd pnand3_2
XDEC_NAND[80] out[2] out[6] out[8] Z[80] vdd gnd pnand3_2
XDEC_NAND[81] out[2] out[6] out[9] Z[81] vdd gnd pnand3_2
XDEC_NAND[82] out[2] out[6] out[10] Z[82] vdd gnd pnand3_2
XDEC_NAND[83] out[2] out[6] out[11] Z[83] vdd gnd pnand3_2
XDEC_NAND[84] out[2] out[6] out[12] Z[84] vdd gnd pnand3_2
XDEC_NAND[85] out[2] out[6] out[13] Z[85] vdd gnd pnand3_2
XDEC_NAND[86] out[2] out[6] out[14] Z[86] vdd gnd pnand3_2
XDEC_NAND[87] out[2] out[6] out[15] Z[87] vdd gnd pnand3_2
XDEC_NAND[88] out[2] out[7] out[8] Z[88] vdd gnd pnand3_2
XDEC_NAND[89] out[2] out[7] out[9] Z[89] vdd gnd pnand3_2
XDEC_NAND[90] out[2] out[7] out[10] Z[90] vdd gnd pnand3_2
XDEC_NAND[91] out[2] out[7] out[11] Z[91] vdd gnd pnand3_2
XDEC_NAND[92] out[2] out[7] out[12] Z[92] vdd gnd pnand3_2
XDEC_NAND[93] out[2] out[7] out[13] Z[93] vdd gnd pnand3_2
XDEC_NAND[94] out[2] out[7] out[14] Z[94] vdd gnd pnand3_2
XDEC_NAND[95] out[2] out[7] out[15] Z[95] vdd gnd pnand3_2
XDEC_NAND[96] out[3] out[4] out[8] Z[96] vdd gnd pnand3_2
XDEC_NAND[97] out[3] out[4] out[9] Z[97] vdd gnd pnand3_2
XDEC_NAND[98] out[3] out[4] out[10] Z[98] vdd gnd pnand3_2
XDEC_NAND[99] out[3] out[4] out[11] Z[99] vdd gnd pnand3_2
XDEC_NAND[100] out[3] out[4] out[12] Z[100] vdd gnd pnand3_2
XDEC_NAND[101] out[3] out[4] out[13] Z[101] vdd gnd pnand3_2
XDEC_NAND[102] out[3] out[4] out[14] Z[102] vdd gnd pnand3_2
XDEC_NAND[103] out[3] out[4] out[15] Z[103] vdd gnd pnand3_2
XDEC_NAND[104] out[3] out[5] out[8] Z[104] vdd gnd pnand3_2
XDEC_NAND[105] out[3] out[5] out[9] Z[105] vdd gnd pnand3_2
XDEC_NAND[106] out[3] out[5] out[10] Z[106] vdd gnd pnand3_2
XDEC_NAND[107] out[3] out[5] out[11] Z[107] vdd gnd pnand3_2
XDEC_NAND[108] out[3] out[5] out[12] Z[108] vdd gnd pnand3_2
XDEC_NAND[109] out[3] out[5] out[13] Z[109] vdd gnd pnand3_2
XDEC_NAND[110] out[3] out[5] out[14] Z[110] vdd gnd pnand3_2
XDEC_NAND[111] out[3] out[5] out[15] Z[111] vdd gnd pnand3_2
XDEC_NAND[112] out[3] out[6] out[8] Z[112] vdd gnd pnand3_2
XDEC_NAND[113] out[3] out[6] out[9] Z[113] vdd gnd pnand3_2
XDEC_NAND[114] out[3] out[6] out[10] Z[114] vdd gnd pnand3_2
XDEC_NAND[115] out[3] out[6] out[11] Z[115] vdd gnd pnand3_2
XDEC_NAND[116] out[3] out[6] out[12] Z[116] vdd gnd pnand3_2
XDEC_NAND[117] out[3] out[6] out[13] Z[117] vdd gnd pnand3_2
XDEC_NAND[118] out[3] out[6] out[14] Z[118] vdd gnd pnand3_2
XDEC_NAND[119] out[3] out[6] out[15] Z[119] vdd gnd pnand3_2
XDEC_NAND[120] out[3] out[7] out[8] Z[120] vdd gnd pnand3_2
XDEC_NAND[121] out[3] out[7] out[9] Z[121] vdd gnd pnand3_2
XDEC_NAND[122] out[3] out[7] out[10] Z[122] vdd gnd pnand3_2
XDEC_NAND[123] out[3] out[7] out[11] Z[123] vdd gnd pnand3_2
XDEC_NAND[124] out[3] out[7] out[12] Z[124] vdd gnd pnand3_2
XDEC_NAND[125] out[3] out[7] out[13] Z[125] vdd gnd pnand3_2
XDEC_NAND[126] out[3] out[7] out[14] Z[126] vdd gnd pnand3_2
XDEC_NAND[127] out[3] out[7] out[15] Z[127] vdd gnd pnand3_2
XDEC_INV_[0] Z[0] decode[0] vdd gnd pinv_8
XDEC_INV_[1] Z[1] decode[1] vdd gnd pinv_8
XDEC_INV_[2] Z[2] decode[2] vdd gnd pinv_8
XDEC_INV_[3] Z[3] decode[3] vdd gnd pinv_8
XDEC_INV_[4] Z[4] decode[4] vdd gnd pinv_8
XDEC_INV_[5] Z[5] decode[5] vdd gnd pinv_8
XDEC_INV_[6] Z[6] decode[6] vdd gnd pinv_8
XDEC_INV_[7] Z[7] decode[7] vdd gnd pinv_8
XDEC_INV_[8] Z[8] decode[8] vdd gnd pinv_8
XDEC_INV_[9] Z[9] decode[9] vdd gnd pinv_8
XDEC_INV_[10] Z[10] decode[10] vdd gnd pinv_8
XDEC_INV_[11] Z[11] decode[11] vdd gnd pinv_8
XDEC_INV_[12] Z[12] decode[12] vdd gnd pinv_8
XDEC_INV_[13] Z[13] decode[13] vdd gnd pinv_8
XDEC_INV_[14] Z[14] decode[14] vdd gnd pinv_8
XDEC_INV_[15] Z[15] decode[15] vdd gnd pinv_8
XDEC_INV_[16] Z[16] decode[16] vdd gnd pinv_8
XDEC_INV_[17] Z[17] decode[17] vdd gnd pinv_8
XDEC_INV_[18] Z[18] decode[18] vdd gnd pinv_8
XDEC_INV_[19] Z[19] decode[19] vdd gnd pinv_8
XDEC_INV_[20] Z[20] decode[20] vdd gnd pinv_8
XDEC_INV_[21] Z[21] decode[21] vdd gnd pinv_8
XDEC_INV_[22] Z[22] decode[22] vdd gnd pinv_8
XDEC_INV_[23] Z[23] decode[23] vdd gnd pinv_8
XDEC_INV_[24] Z[24] decode[24] vdd gnd pinv_8
XDEC_INV_[25] Z[25] decode[25] vdd gnd pinv_8
XDEC_INV_[26] Z[26] decode[26] vdd gnd pinv_8
XDEC_INV_[27] Z[27] decode[27] vdd gnd pinv_8
XDEC_INV_[28] Z[28] decode[28] vdd gnd pinv_8
XDEC_INV_[29] Z[29] decode[29] vdd gnd pinv_8
XDEC_INV_[30] Z[30] decode[30] vdd gnd pinv_8
XDEC_INV_[31] Z[31] decode[31] vdd gnd pinv_8
XDEC_INV_[32] Z[32] decode[32] vdd gnd pinv_8
XDEC_INV_[33] Z[33] decode[33] vdd gnd pinv_8
XDEC_INV_[34] Z[34] decode[34] vdd gnd pinv_8
XDEC_INV_[35] Z[35] decode[35] vdd gnd pinv_8
XDEC_INV_[36] Z[36] decode[36] vdd gnd pinv_8
XDEC_INV_[37] Z[37] decode[37] vdd gnd pinv_8
XDEC_INV_[38] Z[38] decode[38] vdd gnd pinv_8
XDEC_INV_[39] Z[39] decode[39] vdd gnd pinv_8
XDEC_INV_[40] Z[40] decode[40] vdd gnd pinv_8
XDEC_INV_[41] Z[41] decode[41] vdd gnd pinv_8
XDEC_INV_[42] Z[42] decode[42] vdd gnd pinv_8
XDEC_INV_[43] Z[43] decode[43] vdd gnd pinv_8
XDEC_INV_[44] Z[44] decode[44] vdd gnd pinv_8
XDEC_INV_[45] Z[45] decode[45] vdd gnd pinv_8
XDEC_INV_[46] Z[46] decode[46] vdd gnd pinv_8
XDEC_INV_[47] Z[47] decode[47] vdd gnd pinv_8
XDEC_INV_[48] Z[48] decode[48] vdd gnd pinv_8
XDEC_INV_[49] Z[49] decode[49] vdd gnd pinv_8
XDEC_INV_[50] Z[50] decode[50] vdd gnd pinv_8
XDEC_INV_[51] Z[51] decode[51] vdd gnd pinv_8
XDEC_INV_[52] Z[52] decode[52] vdd gnd pinv_8
XDEC_INV_[53] Z[53] decode[53] vdd gnd pinv_8
XDEC_INV_[54] Z[54] decode[54] vdd gnd pinv_8
XDEC_INV_[55] Z[55] decode[55] vdd gnd pinv_8
XDEC_INV_[56] Z[56] decode[56] vdd gnd pinv_8
XDEC_INV_[57] Z[57] decode[57] vdd gnd pinv_8
XDEC_INV_[58] Z[58] decode[58] vdd gnd pinv_8
XDEC_INV_[59] Z[59] decode[59] vdd gnd pinv_8
XDEC_INV_[60] Z[60] decode[60] vdd gnd pinv_8
XDEC_INV_[61] Z[61] decode[61] vdd gnd pinv_8
XDEC_INV_[62] Z[62] decode[62] vdd gnd pinv_8
XDEC_INV_[63] Z[63] decode[63] vdd gnd pinv_8
XDEC_INV_[64] Z[64] decode[64] vdd gnd pinv_8
XDEC_INV_[65] Z[65] decode[65] vdd gnd pinv_8
XDEC_INV_[66] Z[66] decode[66] vdd gnd pinv_8
XDEC_INV_[67] Z[67] decode[67] vdd gnd pinv_8
XDEC_INV_[68] Z[68] decode[68] vdd gnd pinv_8
XDEC_INV_[69] Z[69] decode[69] vdd gnd pinv_8
XDEC_INV_[70] Z[70] decode[70] vdd gnd pinv_8
XDEC_INV_[71] Z[71] decode[71] vdd gnd pinv_8
XDEC_INV_[72] Z[72] decode[72] vdd gnd pinv_8
XDEC_INV_[73] Z[73] decode[73] vdd gnd pinv_8
XDEC_INV_[74] Z[74] decode[74] vdd gnd pinv_8
XDEC_INV_[75] Z[75] decode[75] vdd gnd pinv_8
XDEC_INV_[76] Z[76] decode[76] vdd gnd pinv_8
XDEC_INV_[77] Z[77] decode[77] vdd gnd pinv_8
XDEC_INV_[78] Z[78] decode[78] vdd gnd pinv_8
XDEC_INV_[79] Z[79] decode[79] vdd gnd pinv_8
XDEC_INV_[80] Z[80] decode[80] vdd gnd pinv_8
XDEC_INV_[81] Z[81] decode[81] vdd gnd pinv_8
XDEC_INV_[82] Z[82] decode[82] vdd gnd pinv_8
XDEC_INV_[83] Z[83] decode[83] vdd gnd pinv_8
XDEC_INV_[84] Z[84] decode[84] vdd gnd pinv_8
XDEC_INV_[85] Z[85] decode[85] vdd gnd pinv_8
XDEC_INV_[86] Z[86] decode[86] vdd gnd pinv_8
XDEC_INV_[87] Z[87] decode[87] vdd gnd pinv_8
XDEC_INV_[88] Z[88] decode[88] vdd gnd pinv_8
XDEC_INV_[89] Z[89] decode[89] vdd gnd pinv_8
XDEC_INV_[90] Z[90] decode[90] vdd gnd pinv_8
XDEC_INV_[91] Z[91] decode[91] vdd gnd pinv_8
XDEC_INV_[92] Z[92] decode[92] vdd gnd pinv_8
XDEC_INV_[93] Z[93] decode[93] vdd gnd pinv_8
XDEC_INV_[94] Z[94] decode[94] vdd gnd pinv_8
XDEC_INV_[95] Z[95] decode[95] vdd gnd pinv_8
XDEC_INV_[96] Z[96] decode[96] vdd gnd pinv_8
XDEC_INV_[97] Z[97] decode[97] vdd gnd pinv_8
XDEC_INV_[98] Z[98] decode[98] vdd gnd pinv_8
XDEC_INV_[99] Z[99] decode[99] vdd gnd pinv_8
XDEC_INV_[100] Z[100] decode[100] vdd gnd pinv_8
XDEC_INV_[101] Z[101] decode[101] vdd gnd pinv_8
XDEC_INV_[102] Z[102] decode[102] vdd gnd pinv_8
XDEC_INV_[103] Z[103] decode[103] vdd gnd pinv_8
XDEC_INV_[104] Z[104] decode[104] vdd gnd pinv_8
XDEC_INV_[105] Z[105] decode[105] vdd gnd pinv_8
XDEC_INV_[106] Z[106] decode[106] vdd gnd pinv_8
XDEC_INV_[107] Z[107] decode[107] vdd gnd pinv_8
XDEC_INV_[108] Z[108] decode[108] vdd gnd pinv_8
XDEC_INV_[109] Z[109] decode[109] vdd gnd pinv_8
XDEC_INV_[110] Z[110] decode[110] vdd gnd pinv_8
XDEC_INV_[111] Z[111] decode[111] vdd gnd pinv_8
XDEC_INV_[112] Z[112] decode[112] vdd gnd pinv_8
XDEC_INV_[113] Z[113] decode[113] vdd gnd pinv_8
XDEC_INV_[114] Z[114] decode[114] vdd gnd pinv_8
XDEC_INV_[115] Z[115] decode[115] vdd gnd pinv_8
XDEC_INV_[116] Z[116] decode[116] vdd gnd pinv_8
XDEC_INV_[117] Z[117] decode[117] vdd gnd pinv_8
XDEC_INV_[118] Z[118] decode[118] vdd gnd pinv_8
XDEC_INV_[119] Z[119] decode[119] vdd gnd pinv_8
XDEC_INV_[120] Z[120] decode[120] vdd gnd pinv_8
XDEC_INV_[121] Z[121] decode[121] vdd gnd pinv_8
XDEC_INV_[122] Z[122] decode[122] vdd gnd pinv_8
XDEC_INV_[123] Z[123] decode[123] vdd gnd pinv_8
XDEC_INV_[124] Z[124] decode[124] vdd gnd pinv_8
XDEC_INV_[125] Z[125] decode[125] vdd gnd pinv_8
XDEC_INV_[126] Z[126] decode[126] vdd gnd pinv_8
XDEC_INV_[127] Z[127] decode[127] vdd gnd pinv_8
.ENDS hierarchical_decoder_128rows

.SUBCKT msf_address din[0] din[1] din[2] din[3] din[4] din[5] din[6] din[7] dout[0] dout_bar[0] dout[1] dout_bar[1] dout[2] dout_bar[2] dout[3] dout_bar[3] dout[4] dout_bar[4] dout[5] dout_bar[5] dout[6] dout_bar[6] dout[7] dout_bar[7] clk vdd gnd
XXdff0 din[0] dout[0] dout_bar[0] clk vdd gnd ms_flop
XXdff1 din[1] dout[1] dout_bar[1] clk vdd gnd ms_flop
XXdff2 din[2] dout[2] dout_bar[2] clk vdd gnd ms_flop
XXdff3 din[3] dout[3] dout_bar[3] clk vdd gnd ms_flop
XXdff4 din[4] dout[4] dout_bar[4] clk vdd gnd ms_flop
XXdff5 din[5] dout[5] dout_bar[5] clk vdd gnd ms_flop
XXdff6 din[6] dout[6] dout_bar[6] clk vdd gnd ms_flop
XXdff7 din[7] dout[7] dout_bar[7] clk vdd gnd ms_flop
.ENDS msf_address

.SUBCKT msf_data_in din[0] din[1] din[2] din[3] din[4] din[5] din[6] din[7] din[8] din[9] din[10] din[11] din[12] din[13] din[14] din[15] din[16] din[17] din[18] din[19] din[20] din[21] din[22] din[23] din[24] din[25] din[26] din[27] din[28] din[29] din[30] din[31] din[32] din[33] din[34] din[35] din[36] din[37] din[38] din[39] din[40] din[41] din[42] din[43] din[44] din[45] din[46] din[47] din[48] din[49] din[50] din[51] din[52] din[53] din[54] din[55] din[56] din[57] din[58] din[59] din[60] din[61] din[62] din[63] din[64] din[65] din[66] din[67] din[68] din[69] din[70] din[71] din[72] din[73] din[74] din[75] din[76] din[77] din[78] din[79] din[80] din[81] din[82] din[83] din[84] din[85] din[86] din[87] din[88] din[89] din[90] din[91] din[92] din[93] din[94] din[95] din[96] din[97] din[98] din[99] din[100] din[101] din[102] din[103] din[104] din[105] din[106] din[107] din[108] din[109] din[110] din[111] din[112] din[113] din[114] din[115] din[116] din[117] din[118] din[119] din[120] din[121] din[122] din[123] din[124] din[125] din[126] din[127] dout[0] dout_bar[0] dout[1] dout_bar[1] dout[2] dout_bar[2] dout[3] dout_bar[3] dout[4] dout_bar[4] dout[5] dout_bar[5] dout[6] dout_bar[6] dout[7] dout_bar[7] dout[8] dout_bar[8] dout[9] dout_bar[9] dout[10] dout_bar[10] dout[11] dout_bar[11] dout[12] dout_bar[12] dout[13] dout_bar[13] dout[14] dout_bar[14] dout[15] dout_bar[15] dout[16] dout_bar[16] dout[17] dout_bar[17] dout[18] dout_bar[18] dout[19] dout_bar[19] dout[20] dout_bar[20] dout[21] dout_bar[21] dout[22] dout_bar[22] dout[23] dout_bar[23] dout[24] dout_bar[24] dout[25] dout_bar[25] dout[26] dout_bar[26] dout[27] dout_bar[27] dout[28] dout_bar[28] dout[29] dout_bar[29] dout[30] dout_bar[30] dout[31] dout_bar[31] dout[32] dout_bar[32] dout[33] dout_bar[33] dout[34] dout_bar[34] dout[35] dout_bar[35] dout[36] dout_bar[36] dout[37] dout_bar[37] dout[38] dout_bar[38] dout[39] dout_bar[39] dout[40] dout_bar[40] dout[41] dout_bar[41] dout[42] dout_bar[42] dout[43] dout_bar[43] dout[44] dout_bar[44] dout[45] dout_bar[45] dout[46] dout_bar[46] dout[47] dout_bar[47] dout[48] dout_bar[48] dout[49] dout_bar[49] dout[50] dout_bar[50] dout[51] dout_bar[51] dout[52] dout_bar[52] dout[53] dout_bar[53] dout[54] dout_bar[54] dout[55] dout_bar[55] dout[56] dout_bar[56] dout[57] dout_bar[57] dout[58] dout_bar[58] dout[59] dout_bar[59] dout[60] dout_bar[60] dout[61] dout_bar[61] dout[62] dout_bar[62] dout[63] dout_bar[63] dout[64] dout_bar[64] dout[65] dout_bar[65] dout[66] dout_bar[66] dout[67] dout_bar[67] dout[68] dout_bar[68] dout[69] dout_bar[69] dout[70] dout_bar[70] dout[71] dout_bar[71] dout[72] dout_bar[72] dout[73] dout_bar[73] dout[74] dout_bar[74] dout[75] dout_bar[75] dout[76] dout_bar[76] dout[77] dout_bar[77] dout[78] dout_bar[78] dout[79] dout_bar[79] dout[80] dout_bar[80] dout[81] dout_bar[81] dout[82] dout_bar[82] dout[83] dout_bar[83] dout[84] dout_bar[84] dout[85] dout_bar[85] dout[86] dout_bar[86] dout[87] dout_bar[87] dout[88] dout_bar[88] dout[89] dout_bar[89] dout[90] dout_bar[90] dout[91] dout_bar[91] dout[92] dout_bar[92] dout[93] dout_bar[93] dout[94] dout_bar[94] dout[95] dout_bar[95] dout[96] dout_bar[96] dout[97] dout_bar[97] dout[98] dout_bar[98] dout[99] dout_bar[99] dout[100] dout_bar[100] dout[101] dout_bar[101] dout[102] dout_bar[102] dout[103] dout_bar[103] dout[104] dout_bar[104] dout[105] dout_bar[105] dout[106] dout_bar[106] dout[107] dout_bar[107] dout[108] dout_bar[108] dout[109] dout_bar[109] dout[110] dout_bar[110] dout[111] dout_bar[111] dout[112] dout_bar[112] dout[113] dout_bar[113] dout[114] dout_bar[114] dout[115] dout_bar[115] dout[116] dout_bar[116] dout[117] dout_bar[117] dout[118] dout_bar[118] dout[119] dout_bar[119] dout[120] dout_bar[120] dout[121] dout_bar[121] dout[122] dout_bar[122] dout[123] dout_bar[123] dout[124] dout_bar[124] dout[125] dout_bar[125] dout[126] dout_bar[126] dout[127] dout_bar[127] clk vdd gnd
XXdff0 din[0] dout[0] dout_bar[0] clk vdd gnd ms_flop
XXdff2 din[1] dout[1] dout_bar[1] clk vdd gnd ms_flop
XXdff4 din[2] dout[2] dout_bar[2] clk vdd gnd ms_flop
XXdff6 din[3] dout[3] dout_bar[3] clk vdd gnd ms_flop
XXdff8 din[4] dout[4] dout_bar[4] clk vdd gnd ms_flop
XXdff10 din[5] dout[5] dout_bar[5] clk vdd gnd ms_flop
XXdff12 din[6] dout[6] dout_bar[6] clk vdd gnd ms_flop
XXdff14 din[7] dout[7] dout_bar[7] clk vdd gnd ms_flop
XXdff16 din[8] dout[8] dout_bar[8] clk vdd gnd ms_flop
XXdff18 din[9] dout[9] dout_bar[9] clk vdd gnd ms_flop
XXdff20 din[10] dout[10] dout_bar[10] clk vdd gnd ms_flop
XXdff22 din[11] dout[11] dout_bar[11] clk vdd gnd ms_flop
XXdff24 din[12] dout[12] dout_bar[12] clk vdd gnd ms_flop
XXdff26 din[13] dout[13] dout_bar[13] clk vdd gnd ms_flop
XXdff28 din[14] dout[14] dout_bar[14] clk vdd gnd ms_flop
XXdff30 din[15] dout[15] dout_bar[15] clk vdd gnd ms_flop
XXdff32 din[16] dout[16] dout_bar[16] clk vdd gnd ms_flop
XXdff34 din[17] dout[17] dout_bar[17] clk vdd gnd ms_flop
XXdff36 din[18] dout[18] dout_bar[18] clk vdd gnd ms_flop
XXdff38 din[19] dout[19] dout_bar[19] clk vdd gnd ms_flop
XXdff40 din[20] dout[20] dout_bar[20] clk vdd gnd ms_flop
XXdff42 din[21] dout[21] dout_bar[21] clk vdd gnd ms_flop
XXdff44 din[22] dout[22] dout_bar[22] clk vdd gnd ms_flop
XXdff46 din[23] dout[23] dout_bar[23] clk vdd gnd ms_flop
XXdff48 din[24] dout[24] dout_bar[24] clk vdd gnd ms_flop
XXdff50 din[25] dout[25] dout_bar[25] clk vdd gnd ms_flop
XXdff52 din[26] dout[26] dout_bar[26] clk vdd gnd ms_flop
XXdff54 din[27] dout[27] dout_bar[27] clk vdd gnd ms_flop
XXdff56 din[28] dout[28] dout_bar[28] clk vdd gnd ms_flop
XXdff58 din[29] dout[29] dout_bar[29] clk vdd gnd ms_flop
XXdff60 din[30] dout[30] dout_bar[30] clk vdd gnd ms_flop
XXdff62 din[31] dout[31] dout_bar[31] clk vdd gnd ms_flop
XXdff64 din[32] dout[32] dout_bar[32] clk vdd gnd ms_flop
XXdff66 din[33] dout[33] dout_bar[33] clk vdd gnd ms_flop
XXdff68 din[34] dout[34] dout_bar[34] clk vdd gnd ms_flop
XXdff70 din[35] dout[35] dout_bar[35] clk vdd gnd ms_flop
XXdff72 din[36] dout[36] dout_bar[36] clk vdd gnd ms_flop
XXdff74 din[37] dout[37] dout_bar[37] clk vdd gnd ms_flop
XXdff76 din[38] dout[38] dout_bar[38] clk vdd gnd ms_flop
XXdff78 din[39] dout[39] dout_bar[39] clk vdd gnd ms_flop
XXdff80 din[40] dout[40] dout_bar[40] clk vdd gnd ms_flop
XXdff82 din[41] dout[41] dout_bar[41] clk vdd gnd ms_flop
XXdff84 din[42] dout[42] dout_bar[42] clk vdd gnd ms_flop
XXdff86 din[43] dout[43] dout_bar[43] clk vdd gnd ms_flop
XXdff88 din[44] dout[44] dout_bar[44] clk vdd gnd ms_flop
XXdff90 din[45] dout[45] dout_bar[45] clk vdd gnd ms_flop
XXdff92 din[46] dout[46] dout_bar[46] clk vdd gnd ms_flop
XXdff94 din[47] dout[47] dout_bar[47] clk vdd gnd ms_flop
XXdff96 din[48] dout[48] dout_bar[48] clk vdd gnd ms_flop
XXdff98 din[49] dout[49] dout_bar[49] clk vdd gnd ms_flop
XXdff100 din[50] dout[50] dout_bar[50] clk vdd gnd ms_flop
XXdff102 din[51] dout[51] dout_bar[51] clk vdd gnd ms_flop
XXdff104 din[52] dout[52] dout_bar[52] clk vdd gnd ms_flop
XXdff106 din[53] dout[53] dout_bar[53] clk vdd gnd ms_flop
XXdff108 din[54] dout[54] dout_bar[54] clk vdd gnd ms_flop
XXdff110 din[55] dout[55] dout_bar[55] clk vdd gnd ms_flop
XXdff112 din[56] dout[56] dout_bar[56] clk vdd gnd ms_flop
XXdff114 din[57] dout[57] dout_bar[57] clk vdd gnd ms_flop
XXdff116 din[58] dout[58] dout_bar[58] clk vdd gnd ms_flop
XXdff118 din[59] dout[59] dout_bar[59] clk vdd gnd ms_flop
XXdff120 din[60] dout[60] dout_bar[60] clk vdd gnd ms_flop
XXdff122 din[61] dout[61] dout_bar[61] clk vdd gnd ms_flop
XXdff124 din[62] dout[62] dout_bar[62] clk vdd gnd ms_flop
XXdff126 din[63] dout[63] dout_bar[63] clk vdd gnd ms_flop
XXdff128 din[64] dout[64] dout_bar[64] clk vdd gnd ms_flop
XXdff130 din[65] dout[65] dout_bar[65] clk vdd gnd ms_flop
XXdff132 din[66] dout[66] dout_bar[66] clk vdd gnd ms_flop
XXdff134 din[67] dout[67] dout_bar[67] clk vdd gnd ms_flop
XXdff136 din[68] dout[68] dout_bar[68] clk vdd gnd ms_flop
XXdff138 din[69] dout[69] dout_bar[69] clk vdd gnd ms_flop
XXdff140 din[70] dout[70] dout_bar[70] clk vdd gnd ms_flop
XXdff142 din[71] dout[71] dout_bar[71] clk vdd gnd ms_flop
XXdff144 din[72] dout[72] dout_bar[72] clk vdd gnd ms_flop
XXdff146 din[73] dout[73] dout_bar[73] clk vdd gnd ms_flop
XXdff148 din[74] dout[74] dout_bar[74] clk vdd gnd ms_flop
XXdff150 din[75] dout[75] dout_bar[75] clk vdd gnd ms_flop
XXdff152 din[76] dout[76] dout_bar[76] clk vdd gnd ms_flop
XXdff154 din[77] dout[77] dout_bar[77] clk vdd gnd ms_flop
XXdff156 din[78] dout[78] dout_bar[78] clk vdd gnd ms_flop
XXdff158 din[79] dout[79] dout_bar[79] clk vdd gnd ms_flop
XXdff160 din[80] dout[80] dout_bar[80] clk vdd gnd ms_flop
XXdff162 din[81] dout[81] dout_bar[81] clk vdd gnd ms_flop
XXdff164 din[82] dout[82] dout_bar[82] clk vdd gnd ms_flop
XXdff166 din[83] dout[83] dout_bar[83] clk vdd gnd ms_flop
XXdff168 din[84] dout[84] dout_bar[84] clk vdd gnd ms_flop
XXdff170 din[85] dout[85] dout_bar[85] clk vdd gnd ms_flop
XXdff172 din[86] dout[86] dout_bar[86] clk vdd gnd ms_flop
XXdff174 din[87] dout[87] dout_bar[87] clk vdd gnd ms_flop
XXdff176 din[88] dout[88] dout_bar[88] clk vdd gnd ms_flop
XXdff178 din[89] dout[89] dout_bar[89] clk vdd gnd ms_flop
XXdff180 din[90] dout[90] dout_bar[90] clk vdd gnd ms_flop
XXdff182 din[91] dout[91] dout_bar[91] clk vdd gnd ms_flop
XXdff184 din[92] dout[92] dout_bar[92] clk vdd gnd ms_flop
XXdff186 din[93] dout[93] dout_bar[93] clk vdd gnd ms_flop
XXdff188 din[94] dout[94] dout_bar[94] clk vdd gnd ms_flop
XXdff190 din[95] dout[95] dout_bar[95] clk vdd gnd ms_flop
XXdff192 din[96] dout[96] dout_bar[96] clk vdd gnd ms_flop
XXdff194 din[97] dout[97] dout_bar[97] clk vdd gnd ms_flop
XXdff196 din[98] dout[98] dout_bar[98] clk vdd gnd ms_flop
XXdff198 din[99] dout[99] dout_bar[99] clk vdd gnd ms_flop
XXdff200 din[100] dout[100] dout_bar[100] clk vdd gnd ms_flop
XXdff202 din[101] dout[101] dout_bar[101] clk vdd gnd ms_flop
XXdff204 din[102] dout[102] dout_bar[102] clk vdd gnd ms_flop
XXdff206 din[103] dout[103] dout_bar[103] clk vdd gnd ms_flop
XXdff208 din[104] dout[104] dout_bar[104] clk vdd gnd ms_flop
XXdff210 din[105] dout[105] dout_bar[105] clk vdd gnd ms_flop
XXdff212 din[106] dout[106] dout_bar[106] clk vdd gnd ms_flop
XXdff214 din[107] dout[107] dout_bar[107] clk vdd gnd ms_flop
XXdff216 din[108] dout[108] dout_bar[108] clk vdd gnd ms_flop
XXdff218 din[109] dout[109] dout_bar[109] clk vdd gnd ms_flop
XXdff220 din[110] dout[110] dout_bar[110] clk vdd gnd ms_flop
XXdff222 din[111] dout[111] dout_bar[111] clk vdd gnd ms_flop
XXdff224 din[112] dout[112] dout_bar[112] clk vdd gnd ms_flop
XXdff226 din[113] dout[113] dout_bar[113] clk vdd gnd ms_flop
XXdff228 din[114] dout[114] dout_bar[114] clk vdd gnd ms_flop
XXdff230 din[115] dout[115] dout_bar[115] clk vdd gnd ms_flop
XXdff232 din[116] dout[116] dout_bar[116] clk vdd gnd ms_flop
XXdff234 din[117] dout[117] dout_bar[117] clk vdd gnd ms_flop
XXdff236 din[118] dout[118] dout_bar[118] clk vdd gnd ms_flop
XXdff238 din[119] dout[119] dout_bar[119] clk vdd gnd ms_flop
XXdff240 din[120] dout[120] dout_bar[120] clk vdd gnd ms_flop
XXdff242 din[121] dout[121] dout_bar[121] clk vdd gnd ms_flop
XXdff244 din[122] dout[122] dout_bar[122] clk vdd gnd ms_flop
XXdff246 din[123] dout[123] dout_bar[123] clk vdd gnd ms_flop
XXdff248 din[124] dout[124] dout_bar[124] clk vdd gnd ms_flop
XXdff250 din[125] dout[125] dout_bar[125] clk vdd gnd ms_flop
XXdff252 din[126] dout[126] dout_bar[126] clk vdd gnd ms_flop
XXdff254 din[127] dout[127] dout_bar[127] clk vdd gnd ms_flop
.ENDS msf_data_in
*********************** tri_gate ******************************

.SUBCKT tri_gate in out en en_bar vdd gnd

M_1 net_2 in_inv gnd gnd n W='1.2*1u' L=0.6u
M_2 net_3 in_inv vdd vdd p W='2.4*1u' L=0.6u
M_3 out en_bar net_3 vdd p W='2.4*1u' L=0.6u
M_4 out en net_2 gnd n W='1.2*1u' L=0.6u
M_5 in_inv in vdd vdd p W='2.4*1u' L=0.6u
M_6 in_inv in gnd gnd n W='1.2*1u' L=0.6u


.ENDS	

.SUBCKT tri_gate_array in[0] in[1] in[2] in[3] in[4] in[5] in[6] in[7] in[8] in[9] in[10] in[11] in[12] in[13] in[14] in[15] in[16] in[17] in[18] in[19] in[20] in[21] in[22] in[23] in[24] in[25] in[26] in[27] in[28] in[29] in[30] in[31] in[32] in[33] in[34] in[35] in[36] in[37] in[38] in[39] in[40] in[41] in[42] in[43] in[44] in[45] in[46] in[47] in[48] in[49] in[50] in[51] in[52] in[53] in[54] in[55] in[56] in[57] in[58] in[59] in[60] in[61] in[62] in[63] in[64] in[65] in[66] in[67] in[68] in[69] in[70] in[71] in[72] in[73] in[74] in[75] in[76] in[77] in[78] in[79] in[80] in[81] in[82] in[83] in[84] in[85] in[86] in[87] in[88] in[89] in[90] in[91] in[92] in[93] in[94] in[95] in[96] in[97] in[98] in[99] in[100] in[101] in[102] in[103] in[104] in[105] in[106] in[107] in[108] in[109] in[110] in[111] in[112] in[113] in[114] in[115] in[116] in[117] in[118] in[119] in[120] in[121] in[122] in[123] in[124] in[125] in[126] in[127] out[0] out[1] out[2] out[3] out[4] out[5] out[6] out[7] out[8] out[9] out[10] out[11] out[12] out[13] out[14] out[15] out[16] out[17] out[18] out[19] out[20] out[21] out[22] out[23] out[24] out[25] out[26] out[27] out[28] out[29] out[30] out[31] out[32] out[33] out[34] out[35] out[36] out[37] out[38] out[39] out[40] out[41] out[42] out[43] out[44] out[45] out[46] out[47] out[48] out[49] out[50] out[51] out[52] out[53] out[54] out[55] out[56] out[57] out[58] out[59] out[60] out[61] out[62] out[63] out[64] out[65] out[66] out[67] out[68] out[69] out[70] out[71] out[72] out[73] out[74] out[75] out[76] out[77] out[78] out[79] out[80] out[81] out[82] out[83] out[84] out[85] out[86] out[87] out[88] out[89] out[90] out[91] out[92] out[93] out[94] out[95] out[96] out[97] out[98] out[99] out[100] out[101] out[102] out[103] out[104] out[105] out[106] out[107] out[108] out[109] out[110] out[111] out[112] out[113] out[114] out[115] out[116] out[117] out[118] out[119] out[120] out[121] out[122] out[123] out[124] out[125] out[126] out[127] en en_bar vdd gnd
XXtri_gate0 in[0] out[0] en en_bar vdd gnd tri_gate
XXtri_gate2 in[1] out[1] en en_bar vdd gnd tri_gate
XXtri_gate4 in[2] out[2] en en_bar vdd gnd tri_gate
XXtri_gate6 in[3] out[3] en en_bar vdd gnd tri_gate
XXtri_gate8 in[4] out[4] en en_bar vdd gnd tri_gate
XXtri_gate10 in[5] out[5] en en_bar vdd gnd tri_gate
XXtri_gate12 in[6] out[6] en en_bar vdd gnd tri_gate
XXtri_gate14 in[7] out[7] en en_bar vdd gnd tri_gate
XXtri_gate16 in[8] out[8] en en_bar vdd gnd tri_gate
XXtri_gate18 in[9] out[9] en en_bar vdd gnd tri_gate
XXtri_gate20 in[10] out[10] en en_bar vdd gnd tri_gate
XXtri_gate22 in[11] out[11] en en_bar vdd gnd tri_gate
XXtri_gate24 in[12] out[12] en en_bar vdd gnd tri_gate
XXtri_gate26 in[13] out[13] en en_bar vdd gnd tri_gate
XXtri_gate28 in[14] out[14] en en_bar vdd gnd tri_gate
XXtri_gate30 in[15] out[15] en en_bar vdd gnd tri_gate
XXtri_gate32 in[16] out[16] en en_bar vdd gnd tri_gate
XXtri_gate34 in[17] out[17] en en_bar vdd gnd tri_gate
XXtri_gate36 in[18] out[18] en en_bar vdd gnd tri_gate
XXtri_gate38 in[19] out[19] en en_bar vdd gnd tri_gate
XXtri_gate40 in[20] out[20] en en_bar vdd gnd tri_gate
XXtri_gate42 in[21] out[21] en en_bar vdd gnd tri_gate
XXtri_gate44 in[22] out[22] en en_bar vdd gnd tri_gate
XXtri_gate46 in[23] out[23] en en_bar vdd gnd tri_gate
XXtri_gate48 in[24] out[24] en en_bar vdd gnd tri_gate
XXtri_gate50 in[25] out[25] en en_bar vdd gnd tri_gate
XXtri_gate52 in[26] out[26] en en_bar vdd gnd tri_gate
XXtri_gate54 in[27] out[27] en en_bar vdd gnd tri_gate
XXtri_gate56 in[28] out[28] en en_bar vdd gnd tri_gate
XXtri_gate58 in[29] out[29] en en_bar vdd gnd tri_gate
XXtri_gate60 in[30] out[30] en en_bar vdd gnd tri_gate
XXtri_gate62 in[31] out[31] en en_bar vdd gnd tri_gate
XXtri_gate64 in[32] out[32] en en_bar vdd gnd tri_gate
XXtri_gate66 in[33] out[33] en en_bar vdd gnd tri_gate
XXtri_gate68 in[34] out[34] en en_bar vdd gnd tri_gate
XXtri_gate70 in[35] out[35] en en_bar vdd gnd tri_gate
XXtri_gate72 in[36] out[36] en en_bar vdd gnd tri_gate
XXtri_gate74 in[37] out[37] en en_bar vdd gnd tri_gate
XXtri_gate76 in[38] out[38] en en_bar vdd gnd tri_gate
XXtri_gate78 in[39] out[39] en en_bar vdd gnd tri_gate
XXtri_gate80 in[40] out[40] en en_bar vdd gnd tri_gate
XXtri_gate82 in[41] out[41] en en_bar vdd gnd tri_gate
XXtri_gate84 in[42] out[42] en en_bar vdd gnd tri_gate
XXtri_gate86 in[43] out[43] en en_bar vdd gnd tri_gate
XXtri_gate88 in[44] out[44] en en_bar vdd gnd tri_gate
XXtri_gate90 in[45] out[45] en en_bar vdd gnd tri_gate
XXtri_gate92 in[46] out[46] en en_bar vdd gnd tri_gate
XXtri_gate94 in[47] out[47] en en_bar vdd gnd tri_gate
XXtri_gate96 in[48] out[48] en en_bar vdd gnd tri_gate
XXtri_gate98 in[49] out[49] en en_bar vdd gnd tri_gate
XXtri_gate100 in[50] out[50] en en_bar vdd gnd tri_gate
XXtri_gate102 in[51] out[51] en en_bar vdd gnd tri_gate
XXtri_gate104 in[52] out[52] en en_bar vdd gnd tri_gate
XXtri_gate106 in[53] out[53] en en_bar vdd gnd tri_gate
XXtri_gate108 in[54] out[54] en en_bar vdd gnd tri_gate
XXtri_gate110 in[55] out[55] en en_bar vdd gnd tri_gate
XXtri_gate112 in[56] out[56] en en_bar vdd gnd tri_gate
XXtri_gate114 in[57] out[57] en en_bar vdd gnd tri_gate
XXtri_gate116 in[58] out[58] en en_bar vdd gnd tri_gate
XXtri_gate118 in[59] out[59] en en_bar vdd gnd tri_gate
XXtri_gate120 in[60] out[60] en en_bar vdd gnd tri_gate
XXtri_gate122 in[61] out[61] en en_bar vdd gnd tri_gate
XXtri_gate124 in[62] out[62] en en_bar vdd gnd tri_gate
XXtri_gate126 in[63] out[63] en en_bar vdd gnd tri_gate
XXtri_gate128 in[64] out[64] en en_bar vdd gnd tri_gate
XXtri_gate130 in[65] out[65] en en_bar vdd gnd tri_gate
XXtri_gate132 in[66] out[66] en en_bar vdd gnd tri_gate
XXtri_gate134 in[67] out[67] en en_bar vdd gnd tri_gate
XXtri_gate136 in[68] out[68] en en_bar vdd gnd tri_gate
XXtri_gate138 in[69] out[69] en en_bar vdd gnd tri_gate
XXtri_gate140 in[70] out[70] en en_bar vdd gnd tri_gate
XXtri_gate142 in[71] out[71] en en_bar vdd gnd tri_gate
XXtri_gate144 in[72] out[72] en en_bar vdd gnd tri_gate
XXtri_gate146 in[73] out[73] en en_bar vdd gnd tri_gate
XXtri_gate148 in[74] out[74] en en_bar vdd gnd tri_gate
XXtri_gate150 in[75] out[75] en en_bar vdd gnd tri_gate
XXtri_gate152 in[76] out[76] en en_bar vdd gnd tri_gate
XXtri_gate154 in[77] out[77] en en_bar vdd gnd tri_gate
XXtri_gate156 in[78] out[78] en en_bar vdd gnd tri_gate
XXtri_gate158 in[79] out[79] en en_bar vdd gnd tri_gate
XXtri_gate160 in[80] out[80] en en_bar vdd gnd tri_gate
XXtri_gate162 in[81] out[81] en en_bar vdd gnd tri_gate
XXtri_gate164 in[82] out[82] en en_bar vdd gnd tri_gate
XXtri_gate166 in[83] out[83] en en_bar vdd gnd tri_gate
XXtri_gate168 in[84] out[84] en en_bar vdd gnd tri_gate
XXtri_gate170 in[85] out[85] en en_bar vdd gnd tri_gate
XXtri_gate172 in[86] out[86] en en_bar vdd gnd tri_gate
XXtri_gate174 in[87] out[87] en en_bar vdd gnd tri_gate
XXtri_gate176 in[88] out[88] en en_bar vdd gnd tri_gate
XXtri_gate178 in[89] out[89] en en_bar vdd gnd tri_gate
XXtri_gate180 in[90] out[90] en en_bar vdd gnd tri_gate
XXtri_gate182 in[91] out[91] en en_bar vdd gnd tri_gate
XXtri_gate184 in[92] out[92] en en_bar vdd gnd tri_gate
XXtri_gate186 in[93] out[93] en en_bar vdd gnd tri_gate
XXtri_gate188 in[94] out[94] en en_bar vdd gnd tri_gate
XXtri_gate190 in[95] out[95] en en_bar vdd gnd tri_gate
XXtri_gate192 in[96] out[96] en en_bar vdd gnd tri_gate
XXtri_gate194 in[97] out[97] en en_bar vdd gnd tri_gate
XXtri_gate196 in[98] out[98] en en_bar vdd gnd tri_gate
XXtri_gate198 in[99] out[99] en en_bar vdd gnd tri_gate
XXtri_gate200 in[100] out[100] en en_bar vdd gnd tri_gate
XXtri_gate202 in[101] out[101] en en_bar vdd gnd tri_gate
XXtri_gate204 in[102] out[102] en en_bar vdd gnd tri_gate
XXtri_gate206 in[103] out[103] en en_bar vdd gnd tri_gate
XXtri_gate208 in[104] out[104] en en_bar vdd gnd tri_gate
XXtri_gate210 in[105] out[105] en en_bar vdd gnd tri_gate
XXtri_gate212 in[106] out[106] en en_bar vdd gnd tri_gate
XXtri_gate214 in[107] out[107] en en_bar vdd gnd tri_gate
XXtri_gate216 in[108] out[108] en en_bar vdd gnd tri_gate
XXtri_gate218 in[109] out[109] en en_bar vdd gnd tri_gate
XXtri_gate220 in[110] out[110] en en_bar vdd gnd tri_gate
XXtri_gate222 in[111] out[111] en en_bar vdd gnd tri_gate
XXtri_gate224 in[112] out[112] en en_bar vdd gnd tri_gate
XXtri_gate226 in[113] out[113] en en_bar vdd gnd tri_gate
XXtri_gate228 in[114] out[114] en en_bar vdd gnd tri_gate
XXtri_gate230 in[115] out[115] en en_bar vdd gnd tri_gate
XXtri_gate232 in[116] out[116] en en_bar vdd gnd tri_gate
XXtri_gate234 in[117] out[117] en en_bar vdd gnd tri_gate
XXtri_gate236 in[118] out[118] en en_bar vdd gnd tri_gate
XXtri_gate238 in[119] out[119] en en_bar vdd gnd tri_gate
XXtri_gate240 in[120] out[120] en en_bar vdd gnd tri_gate
XXtri_gate242 in[121] out[121] en en_bar vdd gnd tri_gate
XXtri_gate244 in[122] out[122] en en_bar vdd gnd tri_gate
XXtri_gate246 in[123] out[123] en en_bar vdd gnd tri_gate
XXtri_gate248 in[124] out[124] en en_bar vdd gnd tri_gate
XXtri_gate250 in[125] out[125] en en_bar vdd gnd tri_gate
XXtri_gate252 in[126] out[126] en en_bar vdd gnd tri_gate
XXtri_gate254 in[127] out[127] en en_bar vdd gnd tri_gate
.ENDS tri_gate_array

.SUBCKT pinv_11 A Z vdd gnd
Mpinv_pmos Z A vdd vdd p m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpinv_nmos Z A gnd gnd n m=1 w=1.2u l=0.6u pd=3.6u ps=3.6u as=1.8p ad=1.8p
.ENDS pinv_11

.SUBCKT pinv_12 A Z vdd gnd
Mpinv_pmos Z A vdd vdd p m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpinv_nmos Z A gnd gnd n m=1 w=1.2u l=0.6u pd=3.6u ps=3.6u as=1.8p ad=1.8p
.ENDS pinv_12

.SUBCKT pnand2_4 A B Z vdd gnd
Mpnand2_pmos1 vdd A Z vdd p m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpnand2_pmos2 Z B vdd vdd p m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpnand2_nmos1 Z B net1 gnd n m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpnand2_nmos2 net1 A gnd gnd n m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
.ENDS pnand2_4

.SUBCKT wordline_driver in[0] in[1] in[2] in[3] in[4] in[5] in[6] in[7] in[8] in[9] in[10] in[11] in[12] in[13] in[14] in[15] in[16] in[17] in[18] in[19] in[20] in[21] in[22] in[23] in[24] in[25] in[26] in[27] in[28] in[29] in[30] in[31] in[32] in[33] in[34] in[35] in[36] in[37] in[38] in[39] in[40] in[41] in[42] in[43] in[44] in[45] in[46] in[47] in[48] in[49] in[50] in[51] in[52] in[53] in[54] in[55] in[56] in[57] in[58] in[59] in[60] in[61] in[62] in[63] in[64] in[65] in[66] in[67] in[68] in[69] in[70] in[71] in[72] in[73] in[74] in[75] in[76] in[77] in[78] in[79] in[80] in[81] in[82] in[83] in[84] in[85] in[86] in[87] in[88] in[89] in[90] in[91] in[92] in[93] in[94] in[95] in[96] in[97] in[98] in[99] in[100] in[101] in[102] in[103] in[104] in[105] in[106] in[107] in[108] in[109] in[110] in[111] in[112] in[113] in[114] in[115] in[116] in[117] in[118] in[119] in[120] in[121] in[122] in[123] in[124] in[125] in[126] in[127] wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55] wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63] wl[64] wl[65] wl[66] wl[67] wl[68] wl[69] wl[70] wl[71] wl[72] wl[73] wl[74] wl[75] wl[76] wl[77] wl[78] wl[79] wl[80] wl[81] wl[82] wl[83] wl[84] wl[85] wl[86] wl[87] wl[88] wl[89] wl[90] wl[91] wl[92] wl[93] wl[94] wl[95] wl[96] wl[97] wl[98] wl[99] wl[100] wl[101] wl[102] wl[103] wl[104] wl[105] wl[106] wl[107] wl[108] wl[109] wl[110] wl[111] wl[112] wl[113] wl[114] wl[115] wl[116] wl[117] wl[118] wl[119] wl[120] wl[121] wl[122] wl[123] wl[124] wl[125] wl[126] wl[127] en vdd gnd
Xwl_driver_inv_en0 en en_bar[0] vdd gnd pinv_12
Xwl_driver_nand0 en_bar[0] in[0] net[0] vdd gnd pnand2_4
Xwl_driver_inv0 net[0] wl[0] vdd gnd pinv_11
Xwl_driver_inv_en1 en en_bar[1] vdd gnd pinv_12
Xwl_driver_nand1 en_bar[1] in[1] net[1] vdd gnd pnand2_4
Xwl_driver_inv1 net[1] wl[1] vdd gnd pinv_11
Xwl_driver_inv_en2 en en_bar[2] vdd gnd pinv_12
Xwl_driver_nand2 en_bar[2] in[2] net[2] vdd gnd pnand2_4
Xwl_driver_inv2 net[2] wl[2] vdd gnd pinv_11
Xwl_driver_inv_en3 en en_bar[3] vdd gnd pinv_12
Xwl_driver_nand3 en_bar[3] in[3] net[3] vdd gnd pnand2_4
Xwl_driver_inv3 net[3] wl[3] vdd gnd pinv_11
Xwl_driver_inv_en4 en en_bar[4] vdd gnd pinv_12
Xwl_driver_nand4 en_bar[4] in[4] net[4] vdd gnd pnand2_4
Xwl_driver_inv4 net[4] wl[4] vdd gnd pinv_11
Xwl_driver_inv_en5 en en_bar[5] vdd gnd pinv_12
Xwl_driver_nand5 en_bar[5] in[5] net[5] vdd gnd pnand2_4
Xwl_driver_inv5 net[5] wl[5] vdd gnd pinv_11
Xwl_driver_inv_en6 en en_bar[6] vdd gnd pinv_12
Xwl_driver_nand6 en_bar[6] in[6] net[6] vdd gnd pnand2_4
Xwl_driver_inv6 net[6] wl[6] vdd gnd pinv_11
Xwl_driver_inv_en7 en en_bar[7] vdd gnd pinv_12
Xwl_driver_nand7 en_bar[7] in[7] net[7] vdd gnd pnand2_4
Xwl_driver_inv7 net[7] wl[7] vdd gnd pinv_11
Xwl_driver_inv_en8 en en_bar[8] vdd gnd pinv_12
Xwl_driver_nand8 en_bar[8] in[8] net[8] vdd gnd pnand2_4
Xwl_driver_inv8 net[8] wl[8] vdd gnd pinv_11
Xwl_driver_inv_en9 en en_bar[9] vdd gnd pinv_12
Xwl_driver_nand9 en_bar[9] in[9] net[9] vdd gnd pnand2_4
Xwl_driver_inv9 net[9] wl[9] vdd gnd pinv_11
Xwl_driver_inv_en10 en en_bar[10] vdd gnd pinv_12
Xwl_driver_nand10 en_bar[10] in[10] net[10] vdd gnd pnand2_4
Xwl_driver_inv10 net[10] wl[10] vdd gnd pinv_11
Xwl_driver_inv_en11 en en_bar[11] vdd gnd pinv_12
Xwl_driver_nand11 en_bar[11] in[11] net[11] vdd gnd pnand2_4
Xwl_driver_inv11 net[11] wl[11] vdd gnd pinv_11
Xwl_driver_inv_en12 en en_bar[12] vdd gnd pinv_12
Xwl_driver_nand12 en_bar[12] in[12] net[12] vdd gnd pnand2_4
Xwl_driver_inv12 net[12] wl[12] vdd gnd pinv_11
Xwl_driver_inv_en13 en en_bar[13] vdd gnd pinv_12
Xwl_driver_nand13 en_bar[13] in[13] net[13] vdd gnd pnand2_4
Xwl_driver_inv13 net[13] wl[13] vdd gnd pinv_11
Xwl_driver_inv_en14 en en_bar[14] vdd gnd pinv_12
Xwl_driver_nand14 en_bar[14] in[14] net[14] vdd gnd pnand2_4
Xwl_driver_inv14 net[14] wl[14] vdd gnd pinv_11
Xwl_driver_inv_en15 en en_bar[15] vdd gnd pinv_12
Xwl_driver_nand15 en_bar[15] in[15] net[15] vdd gnd pnand2_4
Xwl_driver_inv15 net[15] wl[15] vdd gnd pinv_11
Xwl_driver_inv_en16 en en_bar[16] vdd gnd pinv_12
Xwl_driver_nand16 en_bar[16] in[16] net[16] vdd gnd pnand2_4
Xwl_driver_inv16 net[16] wl[16] vdd gnd pinv_11
Xwl_driver_inv_en17 en en_bar[17] vdd gnd pinv_12
Xwl_driver_nand17 en_bar[17] in[17] net[17] vdd gnd pnand2_4
Xwl_driver_inv17 net[17] wl[17] vdd gnd pinv_11
Xwl_driver_inv_en18 en en_bar[18] vdd gnd pinv_12
Xwl_driver_nand18 en_bar[18] in[18] net[18] vdd gnd pnand2_4
Xwl_driver_inv18 net[18] wl[18] vdd gnd pinv_11
Xwl_driver_inv_en19 en en_bar[19] vdd gnd pinv_12
Xwl_driver_nand19 en_bar[19] in[19] net[19] vdd gnd pnand2_4
Xwl_driver_inv19 net[19] wl[19] vdd gnd pinv_11
Xwl_driver_inv_en20 en en_bar[20] vdd gnd pinv_12
Xwl_driver_nand20 en_bar[20] in[20] net[20] vdd gnd pnand2_4
Xwl_driver_inv20 net[20] wl[20] vdd gnd pinv_11
Xwl_driver_inv_en21 en en_bar[21] vdd gnd pinv_12
Xwl_driver_nand21 en_bar[21] in[21] net[21] vdd gnd pnand2_4
Xwl_driver_inv21 net[21] wl[21] vdd gnd pinv_11
Xwl_driver_inv_en22 en en_bar[22] vdd gnd pinv_12
Xwl_driver_nand22 en_bar[22] in[22] net[22] vdd gnd pnand2_4
Xwl_driver_inv22 net[22] wl[22] vdd gnd pinv_11
Xwl_driver_inv_en23 en en_bar[23] vdd gnd pinv_12
Xwl_driver_nand23 en_bar[23] in[23] net[23] vdd gnd pnand2_4
Xwl_driver_inv23 net[23] wl[23] vdd gnd pinv_11
Xwl_driver_inv_en24 en en_bar[24] vdd gnd pinv_12
Xwl_driver_nand24 en_bar[24] in[24] net[24] vdd gnd pnand2_4
Xwl_driver_inv24 net[24] wl[24] vdd gnd pinv_11
Xwl_driver_inv_en25 en en_bar[25] vdd gnd pinv_12
Xwl_driver_nand25 en_bar[25] in[25] net[25] vdd gnd pnand2_4
Xwl_driver_inv25 net[25] wl[25] vdd gnd pinv_11
Xwl_driver_inv_en26 en en_bar[26] vdd gnd pinv_12
Xwl_driver_nand26 en_bar[26] in[26] net[26] vdd gnd pnand2_4
Xwl_driver_inv26 net[26] wl[26] vdd gnd pinv_11
Xwl_driver_inv_en27 en en_bar[27] vdd gnd pinv_12
Xwl_driver_nand27 en_bar[27] in[27] net[27] vdd gnd pnand2_4
Xwl_driver_inv27 net[27] wl[27] vdd gnd pinv_11
Xwl_driver_inv_en28 en en_bar[28] vdd gnd pinv_12
Xwl_driver_nand28 en_bar[28] in[28] net[28] vdd gnd pnand2_4
Xwl_driver_inv28 net[28] wl[28] vdd gnd pinv_11
Xwl_driver_inv_en29 en en_bar[29] vdd gnd pinv_12
Xwl_driver_nand29 en_bar[29] in[29] net[29] vdd gnd pnand2_4
Xwl_driver_inv29 net[29] wl[29] vdd gnd pinv_11
Xwl_driver_inv_en30 en en_bar[30] vdd gnd pinv_12
Xwl_driver_nand30 en_bar[30] in[30] net[30] vdd gnd pnand2_4
Xwl_driver_inv30 net[30] wl[30] vdd gnd pinv_11
Xwl_driver_inv_en31 en en_bar[31] vdd gnd pinv_12
Xwl_driver_nand31 en_bar[31] in[31] net[31] vdd gnd pnand2_4
Xwl_driver_inv31 net[31] wl[31] vdd gnd pinv_11
Xwl_driver_inv_en32 en en_bar[32] vdd gnd pinv_12
Xwl_driver_nand32 en_bar[32] in[32] net[32] vdd gnd pnand2_4
Xwl_driver_inv32 net[32] wl[32] vdd gnd pinv_11
Xwl_driver_inv_en33 en en_bar[33] vdd gnd pinv_12
Xwl_driver_nand33 en_bar[33] in[33] net[33] vdd gnd pnand2_4
Xwl_driver_inv33 net[33] wl[33] vdd gnd pinv_11
Xwl_driver_inv_en34 en en_bar[34] vdd gnd pinv_12
Xwl_driver_nand34 en_bar[34] in[34] net[34] vdd gnd pnand2_4
Xwl_driver_inv34 net[34] wl[34] vdd gnd pinv_11
Xwl_driver_inv_en35 en en_bar[35] vdd gnd pinv_12
Xwl_driver_nand35 en_bar[35] in[35] net[35] vdd gnd pnand2_4
Xwl_driver_inv35 net[35] wl[35] vdd gnd pinv_11
Xwl_driver_inv_en36 en en_bar[36] vdd gnd pinv_12
Xwl_driver_nand36 en_bar[36] in[36] net[36] vdd gnd pnand2_4
Xwl_driver_inv36 net[36] wl[36] vdd gnd pinv_11
Xwl_driver_inv_en37 en en_bar[37] vdd gnd pinv_12
Xwl_driver_nand37 en_bar[37] in[37] net[37] vdd gnd pnand2_4
Xwl_driver_inv37 net[37] wl[37] vdd gnd pinv_11
Xwl_driver_inv_en38 en en_bar[38] vdd gnd pinv_12
Xwl_driver_nand38 en_bar[38] in[38] net[38] vdd gnd pnand2_4
Xwl_driver_inv38 net[38] wl[38] vdd gnd pinv_11
Xwl_driver_inv_en39 en en_bar[39] vdd gnd pinv_12
Xwl_driver_nand39 en_bar[39] in[39] net[39] vdd gnd pnand2_4
Xwl_driver_inv39 net[39] wl[39] vdd gnd pinv_11
Xwl_driver_inv_en40 en en_bar[40] vdd gnd pinv_12
Xwl_driver_nand40 en_bar[40] in[40] net[40] vdd gnd pnand2_4
Xwl_driver_inv40 net[40] wl[40] vdd gnd pinv_11
Xwl_driver_inv_en41 en en_bar[41] vdd gnd pinv_12
Xwl_driver_nand41 en_bar[41] in[41] net[41] vdd gnd pnand2_4
Xwl_driver_inv41 net[41] wl[41] vdd gnd pinv_11
Xwl_driver_inv_en42 en en_bar[42] vdd gnd pinv_12
Xwl_driver_nand42 en_bar[42] in[42] net[42] vdd gnd pnand2_4
Xwl_driver_inv42 net[42] wl[42] vdd gnd pinv_11
Xwl_driver_inv_en43 en en_bar[43] vdd gnd pinv_12
Xwl_driver_nand43 en_bar[43] in[43] net[43] vdd gnd pnand2_4
Xwl_driver_inv43 net[43] wl[43] vdd gnd pinv_11
Xwl_driver_inv_en44 en en_bar[44] vdd gnd pinv_12
Xwl_driver_nand44 en_bar[44] in[44] net[44] vdd gnd pnand2_4
Xwl_driver_inv44 net[44] wl[44] vdd gnd pinv_11
Xwl_driver_inv_en45 en en_bar[45] vdd gnd pinv_12
Xwl_driver_nand45 en_bar[45] in[45] net[45] vdd gnd pnand2_4
Xwl_driver_inv45 net[45] wl[45] vdd gnd pinv_11
Xwl_driver_inv_en46 en en_bar[46] vdd gnd pinv_12
Xwl_driver_nand46 en_bar[46] in[46] net[46] vdd gnd pnand2_4
Xwl_driver_inv46 net[46] wl[46] vdd gnd pinv_11
Xwl_driver_inv_en47 en en_bar[47] vdd gnd pinv_12
Xwl_driver_nand47 en_bar[47] in[47] net[47] vdd gnd pnand2_4
Xwl_driver_inv47 net[47] wl[47] vdd gnd pinv_11
Xwl_driver_inv_en48 en en_bar[48] vdd gnd pinv_12
Xwl_driver_nand48 en_bar[48] in[48] net[48] vdd gnd pnand2_4
Xwl_driver_inv48 net[48] wl[48] vdd gnd pinv_11
Xwl_driver_inv_en49 en en_bar[49] vdd gnd pinv_12
Xwl_driver_nand49 en_bar[49] in[49] net[49] vdd gnd pnand2_4
Xwl_driver_inv49 net[49] wl[49] vdd gnd pinv_11
Xwl_driver_inv_en50 en en_bar[50] vdd gnd pinv_12
Xwl_driver_nand50 en_bar[50] in[50] net[50] vdd gnd pnand2_4
Xwl_driver_inv50 net[50] wl[50] vdd gnd pinv_11
Xwl_driver_inv_en51 en en_bar[51] vdd gnd pinv_12
Xwl_driver_nand51 en_bar[51] in[51] net[51] vdd gnd pnand2_4
Xwl_driver_inv51 net[51] wl[51] vdd gnd pinv_11
Xwl_driver_inv_en52 en en_bar[52] vdd gnd pinv_12
Xwl_driver_nand52 en_bar[52] in[52] net[52] vdd gnd pnand2_4
Xwl_driver_inv52 net[52] wl[52] vdd gnd pinv_11
Xwl_driver_inv_en53 en en_bar[53] vdd gnd pinv_12
Xwl_driver_nand53 en_bar[53] in[53] net[53] vdd gnd pnand2_4
Xwl_driver_inv53 net[53] wl[53] vdd gnd pinv_11
Xwl_driver_inv_en54 en en_bar[54] vdd gnd pinv_12
Xwl_driver_nand54 en_bar[54] in[54] net[54] vdd gnd pnand2_4
Xwl_driver_inv54 net[54] wl[54] vdd gnd pinv_11
Xwl_driver_inv_en55 en en_bar[55] vdd gnd pinv_12
Xwl_driver_nand55 en_bar[55] in[55] net[55] vdd gnd pnand2_4
Xwl_driver_inv55 net[55] wl[55] vdd gnd pinv_11
Xwl_driver_inv_en56 en en_bar[56] vdd gnd pinv_12
Xwl_driver_nand56 en_bar[56] in[56] net[56] vdd gnd pnand2_4
Xwl_driver_inv56 net[56] wl[56] vdd gnd pinv_11
Xwl_driver_inv_en57 en en_bar[57] vdd gnd pinv_12
Xwl_driver_nand57 en_bar[57] in[57] net[57] vdd gnd pnand2_4
Xwl_driver_inv57 net[57] wl[57] vdd gnd pinv_11
Xwl_driver_inv_en58 en en_bar[58] vdd gnd pinv_12
Xwl_driver_nand58 en_bar[58] in[58] net[58] vdd gnd pnand2_4
Xwl_driver_inv58 net[58] wl[58] vdd gnd pinv_11
Xwl_driver_inv_en59 en en_bar[59] vdd gnd pinv_12
Xwl_driver_nand59 en_bar[59] in[59] net[59] vdd gnd pnand2_4
Xwl_driver_inv59 net[59] wl[59] vdd gnd pinv_11
Xwl_driver_inv_en60 en en_bar[60] vdd gnd pinv_12
Xwl_driver_nand60 en_bar[60] in[60] net[60] vdd gnd pnand2_4
Xwl_driver_inv60 net[60] wl[60] vdd gnd pinv_11
Xwl_driver_inv_en61 en en_bar[61] vdd gnd pinv_12
Xwl_driver_nand61 en_bar[61] in[61] net[61] vdd gnd pnand2_4
Xwl_driver_inv61 net[61] wl[61] vdd gnd pinv_11
Xwl_driver_inv_en62 en en_bar[62] vdd gnd pinv_12
Xwl_driver_nand62 en_bar[62] in[62] net[62] vdd gnd pnand2_4
Xwl_driver_inv62 net[62] wl[62] vdd gnd pinv_11
Xwl_driver_inv_en63 en en_bar[63] vdd gnd pinv_12
Xwl_driver_nand63 en_bar[63] in[63] net[63] vdd gnd pnand2_4
Xwl_driver_inv63 net[63] wl[63] vdd gnd pinv_11
Xwl_driver_inv_en64 en en_bar[64] vdd gnd pinv_12
Xwl_driver_nand64 en_bar[64] in[64] net[64] vdd gnd pnand2_4
Xwl_driver_inv64 net[64] wl[64] vdd gnd pinv_11
Xwl_driver_inv_en65 en en_bar[65] vdd gnd pinv_12
Xwl_driver_nand65 en_bar[65] in[65] net[65] vdd gnd pnand2_4
Xwl_driver_inv65 net[65] wl[65] vdd gnd pinv_11
Xwl_driver_inv_en66 en en_bar[66] vdd gnd pinv_12
Xwl_driver_nand66 en_bar[66] in[66] net[66] vdd gnd pnand2_4
Xwl_driver_inv66 net[66] wl[66] vdd gnd pinv_11
Xwl_driver_inv_en67 en en_bar[67] vdd gnd pinv_12
Xwl_driver_nand67 en_bar[67] in[67] net[67] vdd gnd pnand2_4
Xwl_driver_inv67 net[67] wl[67] vdd gnd pinv_11
Xwl_driver_inv_en68 en en_bar[68] vdd gnd pinv_12
Xwl_driver_nand68 en_bar[68] in[68] net[68] vdd gnd pnand2_4
Xwl_driver_inv68 net[68] wl[68] vdd gnd pinv_11
Xwl_driver_inv_en69 en en_bar[69] vdd gnd pinv_12
Xwl_driver_nand69 en_bar[69] in[69] net[69] vdd gnd pnand2_4
Xwl_driver_inv69 net[69] wl[69] vdd gnd pinv_11
Xwl_driver_inv_en70 en en_bar[70] vdd gnd pinv_12
Xwl_driver_nand70 en_bar[70] in[70] net[70] vdd gnd pnand2_4
Xwl_driver_inv70 net[70] wl[70] vdd gnd pinv_11
Xwl_driver_inv_en71 en en_bar[71] vdd gnd pinv_12
Xwl_driver_nand71 en_bar[71] in[71] net[71] vdd gnd pnand2_4
Xwl_driver_inv71 net[71] wl[71] vdd gnd pinv_11
Xwl_driver_inv_en72 en en_bar[72] vdd gnd pinv_12
Xwl_driver_nand72 en_bar[72] in[72] net[72] vdd gnd pnand2_4
Xwl_driver_inv72 net[72] wl[72] vdd gnd pinv_11
Xwl_driver_inv_en73 en en_bar[73] vdd gnd pinv_12
Xwl_driver_nand73 en_bar[73] in[73] net[73] vdd gnd pnand2_4
Xwl_driver_inv73 net[73] wl[73] vdd gnd pinv_11
Xwl_driver_inv_en74 en en_bar[74] vdd gnd pinv_12
Xwl_driver_nand74 en_bar[74] in[74] net[74] vdd gnd pnand2_4
Xwl_driver_inv74 net[74] wl[74] vdd gnd pinv_11
Xwl_driver_inv_en75 en en_bar[75] vdd gnd pinv_12
Xwl_driver_nand75 en_bar[75] in[75] net[75] vdd gnd pnand2_4
Xwl_driver_inv75 net[75] wl[75] vdd gnd pinv_11
Xwl_driver_inv_en76 en en_bar[76] vdd gnd pinv_12
Xwl_driver_nand76 en_bar[76] in[76] net[76] vdd gnd pnand2_4
Xwl_driver_inv76 net[76] wl[76] vdd gnd pinv_11
Xwl_driver_inv_en77 en en_bar[77] vdd gnd pinv_12
Xwl_driver_nand77 en_bar[77] in[77] net[77] vdd gnd pnand2_4
Xwl_driver_inv77 net[77] wl[77] vdd gnd pinv_11
Xwl_driver_inv_en78 en en_bar[78] vdd gnd pinv_12
Xwl_driver_nand78 en_bar[78] in[78] net[78] vdd gnd pnand2_4
Xwl_driver_inv78 net[78] wl[78] vdd gnd pinv_11
Xwl_driver_inv_en79 en en_bar[79] vdd gnd pinv_12
Xwl_driver_nand79 en_bar[79] in[79] net[79] vdd gnd pnand2_4
Xwl_driver_inv79 net[79] wl[79] vdd gnd pinv_11
Xwl_driver_inv_en80 en en_bar[80] vdd gnd pinv_12
Xwl_driver_nand80 en_bar[80] in[80] net[80] vdd gnd pnand2_4
Xwl_driver_inv80 net[80] wl[80] vdd gnd pinv_11
Xwl_driver_inv_en81 en en_bar[81] vdd gnd pinv_12
Xwl_driver_nand81 en_bar[81] in[81] net[81] vdd gnd pnand2_4
Xwl_driver_inv81 net[81] wl[81] vdd gnd pinv_11
Xwl_driver_inv_en82 en en_bar[82] vdd gnd pinv_12
Xwl_driver_nand82 en_bar[82] in[82] net[82] vdd gnd pnand2_4
Xwl_driver_inv82 net[82] wl[82] vdd gnd pinv_11
Xwl_driver_inv_en83 en en_bar[83] vdd gnd pinv_12
Xwl_driver_nand83 en_bar[83] in[83] net[83] vdd gnd pnand2_4
Xwl_driver_inv83 net[83] wl[83] vdd gnd pinv_11
Xwl_driver_inv_en84 en en_bar[84] vdd gnd pinv_12
Xwl_driver_nand84 en_bar[84] in[84] net[84] vdd gnd pnand2_4
Xwl_driver_inv84 net[84] wl[84] vdd gnd pinv_11
Xwl_driver_inv_en85 en en_bar[85] vdd gnd pinv_12
Xwl_driver_nand85 en_bar[85] in[85] net[85] vdd gnd pnand2_4
Xwl_driver_inv85 net[85] wl[85] vdd gnd pinv_11
Xwl_driver_inv_en86 en en_bar[86] vdd gnd pinv_12
Xwl_driver_nand86 en_bar[86] in[86] net[86] vdd gnd pnand2_4
Xwl_driver_inv86 net[86] wl[86] vdd gnd pinv_11
Xwl_driver_inv_en87 en en_bar[87] vdd gnd pinv_12
Xwl_driver_nand87 en_bar[87] in[87] net[87] vdd gnd pnand2_4
Xwl_driver_inv87 net[87] wl[87] vdd gnd pinv_11
Xwl_driver_inv_en88 en en_bar[88] vdd gnd pinv_12
Xwl_driver_nand88 en_bar[88] in[88] net[88] vdd gnd pnand2_4
Xwl_driver_inv88 net[88] wl[88] vdd gnd pinv_11
Xwl_driver_inv_en89 en en_bar[89] vdd gnd pinv_12
Xwl_driver_nand89 en_bar[89] in[89] net[89] vdd gnd pnand2_4
Xwl_driver_inv89 net[89] wl[89] vdd gnd pinv_11
Xwl_driver_inv_en90 en en_bar[90] vdd gnd pinv_12
Xwl_driver_nand90 en_bar[90] in[90] net[90] vdd gnd pnand2_4
Xwl_driver_inv90 net[90] wl[90] vdd gnd pinv_11
Xwl_driver_inv_en91 en en_bar[91] vdd gnd pinv_12
Xwl_driver_nand91 en_bar[91] in[91] net[91] vdd gnd pnand2_4
Xwl_driver_inv91 net[91] wl[91] vdd gnd pinv_11
Xwl_driver_inv_en92 en en_bar[92] vdd gnd pinv_12
Xwl_driver_nand92 en_bar[92] in[92] net[92] vdd gnd pnand2_4
Xwl_driver_inv92 net[92] wl[92] vdd gnd pinv_11
Xwl_driver_inv_en93 en en_bar[93] vdd gnd pinv_12
Xwl_driver_nand93 en_bar[93] in[93] net[93] vdd gnd pnand2_4
Xwl_driver_inv93 net[93] wl[93] vdd gnd pinv_11
Xwl_driver_inv_en94 en en_bar[94] vdd gnd pinv_12
Xwl_driver_nand94 en_bar[94] in[94] net[94] vdd gnd pnand2_4
Xwl_driver_inv94 net[94] wl[94] vdd gnd pinv_11
Xwl_driver_inv_en95 en en_bar[95] vdd gnd pinv_12
Xwl_driver_nand95 en_bar[95] in[95] net[95] vdd gnd pnand2_4
Xwl_driver_inv95 net[95] wl[95] vdd gnd pinv_11
Xwl_driver_inv_en96 en en_bar[96] vdd gnd pinv_12
Xwl_driver_nand96 en_bar[96] in[96] net[96] vdd gnd pnand2_4
Xwl_driver_inv96 net[96] wl[96] vdd gnd pinv_11
Xwl_driver_inv_en97 en en_bar[97] vdd gnd pinv_12
Xwl_driver_nand97 en_bar[97] in[97] net[97] vdd gnd pnand2_4
Xwl_driver_inv97 net[97] wl[97] vdd gnd pinv_11
Xwl_driver_inv_en98 en en_bar[98] vdd gnd pinv_12
Xwl_driver_nand98 en_bar[98] in[98] net[98] vdd gnd pnand2_4
Xwl_driver_inv98 net[98] wl[98] vdd gnd pinv_11
Xwl_driver_inv_en99 en en_bar[99] vdd gnd pinv_12
Xwl_driver_nand99 en_bar[99] in[99] net[99] vdd gnd pnand2_4
Xwl_driver_inv99 net[99] wl[99] vdd gnd pinv_11
Xwl_driver_inv_en100 en en_bar[100] vdd gnd pinv_12
Xwl_driver_nand100 en_bar[100] in[100] net[100] vdd gnd pnand2_4
Xwl_driver_inv100 net[100] wl[100] vdd gnd pinv_11
Xwl_driver_inv_en101 en en_bar[101] vdd gnd pinv_12
Xwl_driver_nand101 en_bar[101] in[101] net[101] vdd gnd pnand2_4
Xwl_driver_inv101 net[101] wl[101] vdd gnd pinv_11
Xwl_driver_inv_en102 en en_bar[102] vdd gnd pinv_12
Xwl_driver_nand102 en_bar[102] in[102] net[102] vdd gnd pnand2_4
Xwl_driver_inv102 net[102] wl[102] vdd gnd pinv_11
Xwl_driver_inv_en103 en en_bar[103] vdd gnd pinv_12
Xwl_driver_nand103 en_bar[103] in[103] net[103] vdd gnd pnand2_4
Xwl_driver_inv103 net[103] wl[103] vdd gnd pinv_11
Xwl_driver_inv_en104 en en_bar[104] vdd gnd pinv_12
Xwl_driver_nand104 en_bar[104] in[104] net[104] vdd gnd pnand2_4
Xwl_driver_inv104 net[104] wl[104] vdd gnd pinv_11
Xwl_driver_inv_en105 en en_bar[105] vdd gnd pinv_12
Xwl_driver_nand105 en_bar[105] in[105] net[105] vdd gnd pnand2_4
Xwl_driver_inv105 net[105] wl[105] vdd gnd pinv_11
Xwl_driver_inv_en106 en en_bar[106] vdd gnd pinv_12
Xwl_driver_nand106 en_bar[106] in[106] net[106] vdd gnd pnand2_4
Xwl_driver_inv106 net[106] wl[106] vdd gnd pinv_11
Xwl_driver_inv_en107 en en_bar[107] vdd gnd pinv_12
Xwl_driver_nand107 en_bar[107] in[107] net[107] vdd gnd pnand2_4
Xwl_driver_inv107 net[107] wl[107] vdd gnd pinv_11
Xwl_driver_inv_en108 en en_bar[108] vdd gnd pinv_12
Xwl_driver_nand108 en_bar[108] in[108] net[108] vdd gnd pnand2_4
Xwl_driver_inv108 net[108] wl[108] vdd gnd pinv_11
Xwl_driver_inv_en109 en en_bar[109] vdd gnd pinv_12
Xwl_driver_nand109 en_bar[109] in[109] net[109] vdd gnd pnand2_4
Xwl_driver_inv109 net[109] wl[109] vdd gnd pinv_11
Xwl_driver_inv_en110 en en_bar[110] vdd gnd pinv_12
Xwl_driver_nand110 en_bar[110] in[110] net[110] vdd gnd pnand2_4
Xwl_driver_inv110 net[110] wl[110] vdd gnd pinv_11
Xwl_driver_inv_en111 en en_bar[111] vdd gnd pinv_12
Xwl_driver_nand111 en_bar[111] in[111] net[111] vdd gnd pnand2_4
Xwl_driver_inv111 net[111] wl[111] vdd gnd pinv_11
Xwl_driver_inv_en112 en en_bar[112] vdd gnd pinv_12
Xwl_driver_nand112 en_bar[112] in[112] net[112] vdd gnd pnand2_4
Xwl_driver_inv112 net[112] wl[112] vdd gnd pinv_11
Xwl_driver_inv_en113 en en_bar[113] vdd gnd pinv_12
Xwl_driver_nand113 en_bar[113] in[113] net[113] vdd gnd pnand2_4
Xwl_driver_inv113 net[113] wl[113] vdd gnd pinv_11
Xwl_driver_inv_en114 en en_bar[114] vdd gnd pinv_12
Xwl_driver_nand114 en_bar[114] in[114] net[114] vdd gnd pnand2_4
Xwl_driver_inv114 net[114] wl[114] vdd gnd pinv_11
Xwl_driver_inv_en115 en en_bar[115] vdd gnd pinv_12
Xwl_driver_nand115 en_bar[115] in[115] net[115] vdd gnd pnand2_4
Xwl_driver_inv115 net[115] wl[115] vdd gnd pinv_11
Xwl_driver_inv_en116 en en_bar[116] vdd gnd pinv_12
Xwl_driver_nand116 en_bar[116] in[116] net[116] vdd gnd pnand2_4
Xwl_driver_inv116 net[116] wl[116] vdd gnd pinv_11
Xwl_driver_inv_en117 en en_bar[117] vdd gnd pinv_12
Xwl_driver_nand117 en_bar[117] in[117] net[117] vdd gnd pnand2_4
Xwl_driver_inv117 net[117] wl[117] vdd gnd pinv_11
Xwl_driver_inv_en118 en en_bar[118] vdd gnd pinv_12
Xwl_driver_nand118 en_bar[118] in[118] net[118] vdd gnd pnand2_4
Xwl_driver_inv118 net[118] wl[118] vdd gnd pinv_11
Xwl_driver_inv_en119 en en_bar[119] vdd gnd pinv_12
Xwl_driver_nand119 en_bar[119] in[119] net[119] vdd gnd pnand2_4
Xwl_driver_inv119 net[119] wl[119] vdd gnd pinv_11
Xwl_driver_inv_en120 en en_bar[120] vdd gnd pinv_12
Xwl_driver_nand120 en_bar[120] in[120] net[120] vdd gnd pnand2_4
Xwl_driver_inv120 net[120] wl[120] vdd gnd pinv_11
Xwl_driver_inv_en121 en en_bar[121] vdd gnd pinv_12
Xwl_driver_nand121 en_bar[121] in[121] net[121] vdd gnd pnand2_4
Xwl_driver_inv121 net[121] wl[121] vdd gnd pinv_11
Xwl_driver_inv_en122 en en_bar[122] vdd gnd pinv_12
Xwl_driver_nand122 en_bar[122] in[122] net[122] vdd gnd pnand2_4
Xwl_driver_inv122 net[122] wl[122] vdd gnd pinv_11
Xwl_driver_inv_en123 en en_bar[123] vdd gnd pinv_12
Xwl_driver_nand123 en_bar[123] in[123] net[123] vdd gnd pnand2_4
Xwl_driver_inv123 net[123] wl[123] vdd gnd pinv_11
Xwl_driver_inv_en124 en en_bar[124] vdd gnd pinv_12
Xwl_driver_nand124 en_bar[124] in[124] net[124] vdd gnd pnand2_4
Xwl_driver_inv124 net[124] wl[124] vdd gnd pinv_11
Xwl_driver_inv_en125 en en_bar[125] vdd gnd pinv_12
Xwl_driver_nand125 en_bar[125] in[125] net[125] vdd gnd pnand2_4
Xwl_driver_inv125 net[125] wl[125] vdd gnd pinv_11
Xwl_driver_inv_en126 en en_bar[126] vdd gnd pinv_12
Xwl_driver_nand126 en_bar[126] in[126] net[126] vdd gnd pnand2_4
Xwl_driver_inv126 net[126] wl[126] vdd gnd pinv_11
Xwl_driver_inv_en127 en en_bar[127] vdd gnd pinv_12
Xwl_driver_nand127 en_bar[127] in[127] net[127] vdd gnd pnand2_4
Xwl_driver_inv127 net[127] wl[127] vdd gnd pinv_11
.ENDS wordline_driver

.SUBCKT pinv_13 A Z vdd gnd
Mpinv_pmos Z A vdd vdd p m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpinv_nmos Z A gnd gnd n m=1 w=1.2u l=0.6u pd=3.6u ps=3.6u as=1.8p ad=1.8p
.ENDS pinv_13

.SUBCKT pinv_14 A Z vdd gnd
Mpinv_pmos Z A vdd vdd p m=3 w=3.15u l=0.6u pd=7.5u ps=7.5u as=4.725p ad=4.725p
Mpinv_nmos Z A gnd gnd n m=3 w=1.65u l=0.6u pd=4.5u ps=4.5u as=2.475p ad=2.475p
.ENDS pinv_14

.SUBCKT pnor2_2 A B Z vdd gnd
Mpnor2_pmos1 vdd A net1 vdd p m=1 w=3.6u l=0.6u pd=8.4u ps=8.4u as=5.4p ad=5.4p
Mpnor2_pmos2 net1 B Z vdd p m=1 w=3.6u l=0.6u pd=8.4u ps=8.4u as=5.4p ad=5.4p
Mpnor2_nmos1 Z A gnd gnd n m=1 w=1.2u l=0.6u pd=3.6u ps=3.6u as=1.8p ad=1.8p
Mpnor2_nmos2 Z B gnd gnd n m=1 w=1.2u l=0.6u pd=3.6u ps=3.6u as=1.8p ad=1.8p
.ENDS pnor2_2

.SUBCKT pnand2_5 A B Z vdd gnd
Mpnand2_pmos1 vdd A Z vdd p m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpnand2_pmos2 Z B vdd vdd p m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpnand2_nmos1 Z B net1 gnd n m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpnand2_nmos2 net1 A gnd gnd n m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
.ENDS pnand2_5

.SUBCKT bank DATA[0] DATA[1] DATA[2] DATA[3] DATA[4] DATA[5] DATA[6] DATA[7] DATA[8] DATA[9] DATA[10] DATA[11] DATA[12] DATA[13] DATA[14] DATA[15] DATA[16] DATA[17] DATA[18] DATA[19] DATA[20] DATA[21] DATA[22] DATA[23] DATA[24] DATA[25] DATA[26] DATA[27] DATA[28] DATA[29] DATA[30] DATA[31] DATA[32] DATA[33] DATA[34] DATA[35] DATA[36] DATA[37] DATA[38] DATA[39] DATA[40] DATA[41] DATA[42] DATA[43] DATA[44] DATA[45] DATA[46] DATA[47] DATA[48] DATA[49] DATA[50] DATA[51] DATA[52] DATA[53] DATA[54] DATA[55] DATA[56] DATA[57] DATA[58] DATA[59] DATA[60] DATA[61] DATA[62] DATA[63] DATA[64] DATA[65] DATA[66] DATA[67] DATA[68] DATA[69] DATA[70] DATA[71] DATA[72] DATA[73] DATA[74] DATA[75] DATA[76] DATA[77] DATA[78] DATA[79] DATA[80] DATA[81] DATA[82] DATA[83] DATA[84] DATA[85] DATA[86] DATA[87] DATA[88] DATA[89] DATA[90] DATA[91] DATA[92] DATA[93] DATA[94] DATA[95] DATA[96] DATA[97] DATA[98] DATA[99] DATA[100] DATA[101] DATA[102] DATA[103] DATA[104] DATA[105] DATA[106] DATA[107] DATA[108] DATA[109] DATA[110] DATA[111] DATA[112] DATA[113] DATA[114] DATA[115] DATA[116] DATA[117] DATA[118] DATA[119] DATA[120] DATA[121] DATA[122] DATA[123] DATA[124] DATA[125] DATA[126] DATA[127] ADDR[0] ADDR[1] ADDR[2] ADDR[3] ADDR[4] ADDR[5] ADDR[6] ADDR[7] bank_sel s_en w_en tri_en_bar tri_en clk_bar clk_buf vdd gnd
Xbitcell_array bl[0] br[0] bl[1] br[1] bl[2] br[2] bl[3] br[3] bl[4] br[4] bl[5] br[5] bl[6] br[6] bl[7] br[7] bl[8] br[8] bl[9] br[9] bl[10] br[10] bl[11] br[11] bl[12] br[12] bl[13] br[13] bl[14] br[14] bl[15] br[15] bl[16] br[16] bl[17] br[17] bl[18] br[18] bl[19] br[19] bl[20] br[20] bl[21] br[21] bl[22] br[22] bl[23] br[23] bl[24] br[24] bl[25] br[25] bl[26] br[26] bl[27] br[27] bl[28] br[28] bl[29] br[29] bl[30] br[30] bl[31] br[31] bl[32] br[32] bl[33] br[33] bl[34] br[34] bl[35] br[35] bl[36] br[36] bl[37] br[37] bl[38] br[38] bl[39] br[39] bl[40] br[40] bl[41] br[41] bl[42] br[42] bl[43] br[43] bl[44] br[44] bl[45] br[45] bl[46] br[46] bl[47] br[47] bl[48] br[48] bl[49] br[49] bl[50] br[50] bl[51] br[51] bl[52] br[52] bl[53] br[53] bl[54] br[54] bl[55] br[55] bl[56] br[56] bl[57] br[57] bl[58] br[58] bl[59] br[59] bl[60] br[60] bl[61] br[61] bl[62] br[62] bl[63] br[63] bl[64] br[64] bl[65] br[65] bl[66] br[66] bl[67] br[67] bl[68] br[68] bl[69] br[69] bl[70] br[70] bl[71] br[71] bl[72] br[72] bl[73] br[73] bl[74] br[74] bl[75] br[75] bl[76] br[76] bl[77] br[77] bl[78] br[78] bl[79] br[79] bl[80] br[80] bl[81] br[81] bl[82] br[82] bl[83] br[83] bl[84] br[84] bl[85] br[85] bl[86] br[86] bl[87] br[87] bl[88] br[88] bl[89] br[89] bl[90] br[90] bl[91] br[91] bl[92] br[92] bl[93] br[93] bl[94] br[94] bl[95] br[95] bl[96] br[96] bl[97] br[97] bl[98] br[98] bl[99] br[99] bl[100] br[100] bl[101] br[101] bl[102] br[102] bl[103] br[103] bl[104] br[104] bl[105] br[105] bl[106] br[106] bl[107] br[107] bl[108] br[108] bl[109] br[109] bl[110] br[110] bl[111] br[111] bl[112] br[112] bl[113] br[113] bl[114] br[114] bl[115] br[115] bl[116] br[116] bl[117] br[117] bl[118] br[118] bl[119] br[119] bl[120] br[120] bl[121] br[121] bl[122] br[122] bl[123] br[123] bl[124] br[124] bl[125] br[125] bl[126] br[126] bl[127] br[127] bl[128] br[128] bl[129] br[129] bl[130] br[130] bl[131] br[131] bl[132] br[132] bl[133] br[133] bl[134] br[134] bl[135] br[135] bl[136] br[136] bl[137] br[137] bl[138] br[138] bl[139] br[139] bl[140] br[140] bl[141] br[141] bl[142] br[142] bl[143] br[143] bl[144] br[144] bl[145] br[145] bl[146] br[146] bl[147] br[147] bl[148] br[148] bl[149] br[149] bl[150] br[150] bl[151] br[151] bl[152] br[152] bl[153] br[153] bl[154] br[154] bl[155] br[155] bl[156] br[156] bl[157] br[157] bl[158] br[158] bl[159] br[159] bl[160] br[160] bl[161] br[161] bl[162] br[162] bl[163] br[163] bl[164] br[164] bl[165] br[165] bl[166] br[166] bl[167] br[167] bl[168] br[168] bl[169] br[169] bl[170] br[170] bl[171] br[171] bl[172] br[172] bl[173] br[173] bl[174] br[174] bl[175] br[175] bl[176] br[176] bl[177] br[177] bl[178] br[178] bl[179] br[179] bl[180] br[180] bl[181] br[181] bl[182] br[182] bl[183] br[183] bl[184] br[184] bl[185] br[185] bl[186] br[186] bl[187] br[187] bl[188] br[188] bl[189] br[189] bl[190] br[190] bl[191] br[191] bl[192] br[192] bl[193] br[193] bl[194] br[194] bl[195] br[195] bl[196] br[196] bl[197] br[197] bl[198] br[198] bl[199] br[199] bl[200] br[200] bl[201] br[201] bl[202] br[202] bl[203] br[203] bl[204] br[204] bl[205] br[205] bl[206] br[206] bl[207] br[207] bl[208] br[208] bl[209] br[209] bl[210] br[210] bl[211] br[211] bl[212] br[212] bl[213] br[213] bl[214] br[214] bl[215] br[215] bl[216] br[216] bl[217] br[217] bl[218] br[218] bl[219] br[219] bl[220] br[220] bl[221] br[221] bl[222] br[222] bl[223] br[223] bl[224] br[224] bl[225] br[225] bl[226] br[226] bl[227] br[227] bl[228] br[228] bl[229] br[229] bl[230] br[230] bl[231] br[231] bl[232] br[232] bl[233] br[233] bl[234] br[234] bl[235] br[235] bl[236] br[236] bl[237] br[237] bl[238] br[238] bl[239] br[239] bl[240] br[240] bl[241] br[241] bl[242] br[242] bl[243] br[243] bl[244] br[244] bl[245] br[245] bl[246] br[246] bl[247] br[247] bl[248] br[248] bl[249] br[249] bl[250] br[250] bl[251] br[251] bl[252] br[252] bl[253] br[253] bl[254] br[254] bl[255] br[255] wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55] wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63] wl[64] wl[65] wl[66] wl[67] wl[68] wl[69] wl[70] wl[71] wl[72] wl[73] wl[74] wl[75] wl[76] wl[77] wl[78] wl[79] wl[80] wl[81] wl[82] wl[83] wl[84] wl[85] wl[86] wl[87] wl[88] wl[89] wl[90] wl[91] wl[92] wl[93] wl[94] wl[95] wl[96] wl[97] wl[98] wl[99] wl[100] wl[101] wl[102] wl[103] wl[104] wl[105] wl[106] wl[107] wl[108] wl[109] wl[110] wl[111] wl[112] wl[113] wl[114] wl[115] wl[116] wl[117] wl[118] wl[119] wl[120] wl[121] wl[122] wl[123] wl[124] wl[125] wl[126] wl[127] vdd gnd bitcell_array
Xprecharge_array bl[0] br[0] bl[1] br[1] bl[2] br[2] bl[3] br[3] bl[4] br[4] bl[5] br[5] bl[6] br[6] bl[7] br[7] bl[8] br[8] bl[9] br[9] bl[10] br[10] bl[11] br[11] bl[12] br[12] bl[13] br[13] bl[14] br[14] bl[15] br[15] bl[16] br[16] bl[17] br[17] bl[18] br[18] bl[19] br[19] bl[20] br[20] bl[21] br[21] bl[22] br[22] bl[23] br[23] bl[24] br[24] bl[25] br[25] bl[26] br[26] bl[27] br[27] bl[28] br[28] bl[29] br[29] bl[30] br[30] bl[31] br[31] bl[32] br[32] bl[33] br[33] bl[34] br[34] bl[35] br[35] bl[36] br[36] bl[37] br[37] bl[38] br[38] bl[39] br[39] bl[40] br[40] bl[41] br[41] bl[42] br[42] bl[43] br[43] bl[44] br[44] bl[45] br[45] bl[46] br[46] bl[47] br[47] bl[48] br[48] bl[49] br[49] bl[50] br[50] bl[51] br[51] bl[52] br[52] bl[53] br[53] bl[54] br[54] bl[55] br[55] bl[56] br[56] bl[57] br[57] bl[58] br[58] bl[59] br[59] bl[60] br[60] bl[61] br[61] bl[62] br[62] bl[63] br[63] bl[64] br[64] bl[65] br[65] bl[66] br[66] bl[67] br[67] bl[68] br[68] bl[69] br[69] bl[70] br[70] bl[71] br[71] bl[72] br[72] bl[73] br[73] bl[74] br[74] bl[75] br[75] bl[76] br[76] bl[77] br[77] bl[78] br[78] bl[79] br[79] bl[80] br[80] bl[81] br[81] bl[82] br[82] bl[83] br[83] bl[84] br[84] bl[85] br[85] bl[86] br[86] bl[87] br[87] bl[88] br[88] bl[89] br[89] bl[90] br[90] bl[91] br[91] bl[92] br[92] bl[93] br[93] bl[94] br[94] bl[95] br[95] bl[96] br[96] bl[97] br[97] bl[98] br[98] bl[99] br[99] bl[100] br[100] bl[101] br[101] bl[102] br[102] bl[103] br[103] bl[104] br[104] bl[105] br[105] bl[106] br[106] bl[107] br[107] bl[108] br[108] bl[109] br[109] bl[110] br[110] bl[111] br[111] bl[112] br[112] bl[113] br[113] bl[114] br[114] bl[115] br[115] bl[116] br[116] bl[117] br[117] bl[118] br[118] bl[119] br[119] bl[120] br[120] bl[121] br[121] bl[122] br[122] bl[123] br[123] bl[124] br[124] bl[125] br[125] bl[126] br[126] bl[127] br[127] bl[128] br[128] bl[129] br[129] bl[130] br[130] bl[131] br[131] bl[132] br[132] bl[133] br[133] bl[134] br[134] bl[135] br[135] bl[136] br[136] bl[137] br[137] bl[138] br[138] bl[139] br[139] bl[140] br[140] bl[141] br[141] bl[142] br[142] bl[143] br[143] bl[144] br[144] bl[145] br[145] bl[146] br[146] bl[147] br[147] bl[148] br[148] bl[149] br[149] bl[150] br[150] bl[151] br[151] bl[152] br[152] bl[153] br[153] bl[154] br[154] bl[155] br[155] bl[156] br[156] bl[157] br[157] bl[158] br[158] bl[159] br[159] bl[160] br[160] bl[161] br[161] bl[162] br[162] bl[163] br[163] bl[164] br[164] bl[165] br[165] bl[166] br[166] bl[167] br[167] bl[168] br[168] bl[169] br[169] bl[170] br[170] bl[171] br[171] bl[172] br[172] bl[173] br[173] bl[174] br[174] bl[175] br[175] bl[176] br[176] bl[177] br[177] bl[178] br[178] bl[179] br[179] bl[180] br[180] bl[181] br[181] bl[182] br[182] bl[183] br[183] bl[184] br[184] bl[185] br[185] bl[186] br[186] bl[187] br[187] bl[188] br[188] bl[189] br[189] bl[190] br[190] bl[191] br[191] bl[192] br[192] bl[193] br[193] bl[194] br[194] bl[195] br[195] bl[196] br[196] bl[197] br[197] bl[198] br[198] bl[199] br[199] bl[200] br[200] bl[201] br[201] bl[202] br[202] bl[203] br[203] bl[204] br[204] bl[205] br[205] bl[206] br[206] bl[207] br[207] bl[208] br[208] bl[209] br[209] bl[210] br[210] bl[211] br[211] bl[212] br[212] bl[213] br[213] bl[214] br[214] bl[215] br[215] bl[216] br[216] bl[217] br[217] bl[218] br[218] bl[219] br[219] bl[220] br[220] bl[221] br[221] bl[222] br[222] bl[223] br[223] bl[224] br[224] bl[225] br[225] bl[226] br[226] bl[227] br[227] bl[228] br[228] bl[229] br[229] bl[230] br[230] bl[231] br[231] bl[232] br[232] bl[233] br[233] bl[234] br[234] bl[235] br[235] bl[236] br[236] bl[237] br[237] bl[238] br[238] bl[239] br[239] bl[240] br[240] bl[241] br[241] bl[242] br[242] bl[243] br[243] bl[244] br[244] bl[245] br[245] bl[246] br[246] bl[247] br[247] bl[248] br[248] bl[249] br[249] bl[250] br[250] bl[251] br[251] bl[252] br[252] bl[253] br[253] bl[254] br[254] bl[255] br[255] gated_clk_bar vdd precharge_array
Xcolumn_mux_array bl[0] br[0] bl[1] br[1] bl[2] br[2] bl[3] br[3] bl[4] br[4] bl[5] br[5] bl[6] br[6] bl[7] br[7] bl[8] br[8] bl[9] br[9] bl[10] br[10] bl[11] br[11] bl[12] br[12] bl[13] br[13] bl[14] br[14] bl[15] br[15] bl[16] br[16] bl[17] br[17] bl[18] br[18] bl[19] br[19] bl[20] br[20] bl[21] br[21] bl[22] br[22] bl[23] br[23] bl[24] br[24] bl[25] br[25] bl[26] br[26] bl[27] br[27] bl[28] br[28] bl[29] br[29] bl[30] br[30] bl[31] br[31] bl[32] br[32] bl[33] br[33] bl[34] br[34] bl[35] br[35] bl[36] br[36] bl[37] br[37] bl[38] br[38] bl[39] br[39] bl[40] br[40] bl[41] br[41] bl[42] br[42] bl[43] br[43] bl[44] br[44] bl[45] br[45] bl[46] br[46] bl[47] br[47] bl[48] br[48] bl[49] br[49] bl[50] br[50] bl[51] br[51] bl[52] br[52] bl[53] br[53] bl[54] br[54] bl[55] br[55] bl[56] br[56] bl[57] br[57] bl[58] br[58] bl[59] br[59] bl[60] br[60] bl[61] br[61] bl[62] br[62] bl[63] br[63] bl[64] br[64] bl[65] br[65] bl[66] br[66] bl[67] br[67] bl[68] br[68] bl[69] br[69] bl[70] br[70] bl[71] br[71] bl[72] br[72] bl[73] br[73] bl[74] br[74] bl[75] br[75] bl[76] br[76] bl[77] br[77] bl[78] br[78] bl[79] br[79] bl[80] br[80] bl[81] br[81] bl[82] br[82] bl[83] br[83] bl[84] br[84] bl[85] br[85] bl[86] br[86] bl[87] br[87] bl[88] br[88] bl[89] br[89] bl[90] br[90] bl[91] br[91] bl[92] br[92] bl[93] br[93] bl[94] br[94] bl[95] br[95] bl[96] br[96] bl[97] br[97] bl[98] br[98] bl[99] br[99] bl[100] br[100] bl[101] br[101] bl[102] br[102] bl[103] br[103] bl[104] br[104] bl[105] br[105] bl[106] br[106] bl[107] br[107] bl[108] br[108] bl[109] br[109] bl[110] br[110] bl[111] br[111] bl[112] br[112] bl[113] br[113] bl[114] br[114] bl[115] br[115] bl[116] br[116] bl[117] br[117] bl[118] br[118] bl[119] br[119] bl[120] br[120] bl[121] br[121] bl[122] br[122] bl[123] br[123] bl[124] br[124] bl[125] br[125] bl[126] br[126] bl[127] br[127] bl[128] br[128] bl[129] br[129] bl[130] br[130] bl[131] br[131] bl[132] br[132] bl[133] br[133] bl[134] br[134] bl[135] br[135] bl[136] br[136] bl[137] br[137] bl[138] br[138] bl[139] br[139] bl[140] br[140] bl[141] br[141] bl[142] br[142] bl[143] br[143] bl[144] br[144] bl[145] br[145] bl[146] br[146] bl[147] br[147] bl[148] br[148] bl[149] br[149] bl[150] br[150] bl[151] br[151] bl[152] br[152] bl[153] br[153] bl[154] br[154] bl[155] br[155] bl[156] br[156] bl[157] br[157] bl[158] br[158] bl[159] br[159] bl[160] br[160] bl[161] br[161] bl[162] br[162] bl[163] br[163] bl[164] br[164] bl[165] br[165] bl[166] br[166] bl[167] br[167] bl[168] br[168] bl[169] br[169] bl[170] br[170] bl[171] br[171] bl[172] br[172] bl[173] br[173] bl[174] br[174] bl[175] br[175] bl[176] br[176] bl[177] br[177] bl[178] br[178] bl[179] br[179] bl[180] br[180] bl[181] br[181] bl[182] br[182] bl[183] br[183] bl[184] br[184] bl[185] br[185] bl[186] br[186] bl[187] br[187] bl[188] br[188] bl[189] br[189] bl[190] br[190] bl[191] br[191] bl[192] br[192] bl[193] br[193] bl[194] br[194] bl[195] br[195] bl[196] br[196] bl[197] br[197] bl[198] br[198] bl[199] br[199] bl[200] br[200] bl[201] br[201] bl[202] br[202] bl[203] br[203] bl[204] br[204] bl[205] br[205] bl[206] br[206] bl[207] br[207] bl[208] br[208] bl[209] br[209] bl[210] br[210] bl[211] br[211] bl[212] br[212] bl[213] br[213] bl[214] br[214] bl[215] br[215] bl[216] br[216] bl[217] br[217] bl[218] br[218] bl[219] br[219] bl[220] br[220] bl[221] br[221] bl[222] br[222] bl[223] br[223] bl[224] br[224] bl[225] br[225] bl[226] br[226] bl[227] br[227] bl[228] br[228] bl[229] br[229] bl[230] br[230] bl[231] br[231] bl[232] br[232] bl[233] br[233] bl[234] br[234] bl[235] br[235] bl[236] br[236] bl[237] br[237] bl[238] br[238] bl[239] br[239] bl[240] br[240] bl[241] br[241] bl[242] br[242] bl[243] br[243] bl[244] br[244] bl[245] br[245] bl[246] br[246] bl[247] br[247] bl[248] br[248] bl[249] br[249] bl[250] br[250] bl[251] br[251] bl[252] br[252] bl[253] br[253] bl[254] br[254] bl[255] br[255] sel[0] sel[1] bl_out[0] br_out[0] bl_out[1] br_out[1] bl_out[2] br_out[2] bl_out[3] br_out[3] bl_out[4] br_out[4] bl_out[5] br_out[5] bl_out[6] br_out[6] bl_out[7] br_out[7] bl_out[8] br_out[8] bl_out[9] br_out[9] bl_out[10] br_out[10] bl_out[11] br_out[11] bl_out[12] br_out[12] bl_out[13] br_out[13] bl_out[14] br_out[14] bl_out[15] br_out[15] bl_out[16] br_out[16] bl_out[17] br_out[17] bl_out[18] br_out[18] bl_out[19] br_out[19] bl_out[20] br_out[20] bl_out[21] br_out[21] bl_out[22] br_out[22] bl_out[23] br_out[23] bl_out[24] br_out[24] bl_out[25] br_out[25] bl_out[26] br_out[26] bl_out[27] br_out[27] bl_out[28] br_out[28] bl_out[29] br_out[29] bl_out[30] br_out[30] bl_out[31] br_out[31] bl_out[32] br_out[32] bl_out[33] br_out[33] bl_out[34] br_out[34] bl_out[35] br_out[35] bl_out[36] br_out[36] bl_out[37] br_out[37] bl_out[38] br_out[38] bl_out[39] br_out[39] bl_out[40] br_out[40] bl_out[41] br_out[41] bl_out[42] br_out[42] bl_out[43] br_out[43] bl_out[44] br_out[44] bl_out[45] br_out[45] bl_out[46] br_out[46] bl_out[47] br_out[47] bl_out[48] br_out[48] bl_out[49] br_out[49] bl_out[50] br_out[50] bl_out[51] br_out[51] bl_out[52] br_out[52] bl_out[53] br_out[53] bl_out[54] br_out[54] bl_out[55] br_out[55] bl_out[56] br_out[56] bl_out[57] br_out[57] bl_out[58] br_out[58] bl_out[59] br_out[59] bl_out[60] br_out[60] bl_out[61] br_out[61] bl_out[62] br_out[62] bl_out[63] br_out[63] bl_out[64] br_out[64] bl_out[65] br_out[65] bl_out[66] br_out[66] bl_out[67] br_out[67] bl_out[68] br_out[68] bl_out[69] br_out[69] bl_out[70] br_out[70] bl_out[71] br_out[71] bl_out[72] br_out[72] bl_out[73] br_out[73] bl_out[74] br_out[74] bl_out[75] br_out[75] bl_out[76] br_out[76] bl_out[77] br_out[77] bl_out[78] br_out[78] bl_out[79] br_out[79] bl_out[80] br_out[80] bl_out[81] br_out[81] bl_out[82] br_out[82] bl_out[83] br_out[83] bl_out[84] br_out[84] bl_out[85] br_out[85] bl_out[86] br_out[86] bl_out[87] br_out[87] bl_out[88] br_out[88] bl_out[89] br_out[89] bl_out[90] br_out[90] bl_out[91] br_out[91] bl_out[92] br_out[92] bl_out[93] br_out[93] bl_out[94] br_out[94] bl_out[95] br_out[95] bl_out[96] br_out[96] bl_out[97] br_out[97] bl_out[98] br_out[98] bl_out[99] br_out[99] bl_out[100] br_out[100] bl_out[101] br_out[101] bl_out[102] br_out[102] bl_out[103] br_out[103] bl_out[104] br_out[104] bl_out[105] br_out[105] bl_out[106] br_out[106] bl_out[107] br_out[107] bl_out[108] br_out[108] bl_out[109] br_out[109] bl_out[110] br_out[110] bl_out[111] br_out[111] bl_out[112] br_out[112] bl_out[113] br_out[113] bl_out[114] br_out[114] bl_out[115] br_out[115] bl_out[116] br_out[116] bl_out[117] br_out[117] bl_out[118] br_out[118] bl_out[119] br_out[119] bl_out[120] br_out[120] bl_out[121] br_out[121] bl_out[122] br_out[122] bl_out[123] br_out[123] bl_out[124] br_out[124] bl_out[125] br_out[125] bl_out[126] br_out[126] bl_out[127] br_out[127] gnd columnmux_array
Xsense_amp_array data_out[0] bl_out[0] br_out[0] data_out[1] bl_out[1] br_out[1] data_out[2] bl_out[2] br_out[2] data_out[3] bl_out[3] br_out[3] data_out[4] bl_out[4] br_out[4] data_out[5] bl_out[5] br_out[5] data_out[6] bl_out[6] br_out[6] data_out[7] bl_out[7] br_out[7] data_out[8] bl_out[8] br_out[8] data_out[9] bl_out[9] br_out[9] data_out[10] bl_out[10] br_out[10] data_out[11] bl_out[11] br_out[11] data_out[12] bl_out[12] br_out[12] data_out[13] bl_out[13] br_out[13] data_out[14] bl_out[14] br_out[14] data_out[15] bl_out[15] br_out[15] data_out[16] bl_out[16] br_out[16] data_out[17] bl_out[17] br_out[17] data_out[18] bl_out[18] br_out[18] data_out[19] bl_out[19] br_out[19] data_out[20] bl_out[20] br_out[20] data_out[21] bl_out[21] br_out[21] data_out[22] bl_out[22] br_out[22] data_out[23] bl_out[23] br_out[23] data_out[24] bl_out[24] br_out[24] data_out[25] bl_out[25] br_out[25] data_out[26] bl_out[26] br_out[26] data_out[27] bl_out[27] br_out[27] data_out[28] bl_out[28] br_out[28] data_out[29] bl_out[29] br_out[29] data_out[30] bl_out[30] br_out[30] data_out[31] bl_out[31] br_out[31] data_out[32] bl_out[32] br_out[32] data_out[33] bl_out[33] br_out[33] data_out[34] bl_out[34] br_out[34] data_out[35] bl_out[35] br_out[35] data_out[36] bl_out[36] br_out[36] data_out[37] bl_out[37] br_out[37] data_out[38] bl_out[38] br_out[38] data_out[39] bl_out[39] br_out[39] data_out[40] bl_out[40] br_out[40] data_out[41] bl_out[41] br_out[41] data_out[42] bl_out[42] br_out[42] data_out[43] bl_out[43] br_out[43] data_out[44] bl_out[44] br_out[44] data_out[45] bl_out[45] br_out[45] data_out[46] bl_out[46] br_out[46] data_out[47] bl_out[47] br_out[47] data_out[48] bl_out[48] br_out[48] data_out[49] bl_out[49] br_out[49] data_out[50] bl_out[50] br_out[50] data_out[51] bl_out[51] br_out[51] data_out[52] bl_out[52] br_out[52] data_out[53] bl_out[53] br_out[53] data_out[54] bl_out[54] br_out[54] data_out[55] bl_out[55] br_out[55] data_out[56] bl_out[56] br_out[56] data_out[57] bl_out[57] br_out[57] data_out[58] bl_out[58] br_out[58] data_out[59] bl_out[59] br_out[59] data_out[60] bl_out[60] br_out[60] data_out[61] bl_out[61] br_out[61] data_out[62] bl_out[62] br_out[62] data_out[63] bl_out[63] br_out[63] data_out[64] bl_out[64] br_out[64] data_out[65] bl_out[65] br_out[65] data_out[66] bl_out[66] br_out[66] data_out[67] bl_out[67] br_out[67] data_out[68] bl_out[68] br_out[68] data_out[69] bl_out[69] br_out[69] data_out[70] bl_out[70] br_out[70] data_out[71] bl_out[71] br_out[71] data_out[72] bl_out[72] br_out[72] data_out[73] bl_out[73] br_out[73] data_out[74] bl_out[74] br_out[74] data_out[75] bl_out[75] br_out[75] data_out[76] bl_out[76] br_out[76] data_out[77] bl_out[77] br_out[77] data_out[78] bl_out[78] br_out[78] data_out[79] bl_out[79] br_out[79] data_out[80] bl_out[80] br_out[80] data_out[81] bl_out[81] br_out[81] data_out[82] bl_out[82] br_out[82] data_out[83] bl_out[83] br_out[83] data_out[84] bl_out[84] br_out[84] data_out[85] bl_out[85] br_out[85] data_out[86] bl_out[86] br_out[86] data_out[87] bl_out[87] br_out[87] data_out[88] bl_out[88] br_out[88] data_out[89] bl_out[89] br_out[89] data_out[90] bl_out[90] br_out[90] data_out[91] bl_out[91] br_out[91] data_out[92] bl_out[92] br_out[92] data_out[93] bl_out[93] br_out[93] data_out[94] bl_out[94] br_out[94] data_out[95] bl_out[95] br_out[95] data_out[96] bl_out[96] br_out[96] data_out[97] bl_out[97] br_out[97] data_out[98] bl_out[98] br_out[98] data_out[99] bl_out[99] br_out[99] data_out[100] bl_out[100] br_out[100] data_out[101] bl_out[101] br_out[101] data_out[102] bl_out[102] br_out[102] data_out[103] bl_out[103] br_out[103] data_out[104] bl_out[104] br_out[104] data_out[105] bl_out[105] br_out[105] data_out[106] bl_out[106] br_out[106] data_out[107] bl_out[107] br_out[107] data_out[108] bl_out[108] br_out[108] data_out[109] bl_out[109] br_out[109] data_out[110] bl_out[110] br_out[110] data_out[111] bl_out[111] br_out[111] data_out[112] bl_out[112] br_out[112] data_out[113] bl_out[113] br_out[113] data_out[114] bl_out[114] br_out[114] data_out[115] bl_out[115] br_out[115] data_out[116] bl_out[116] br_out[116] data_out[117] bl_out[117] br_out[117] data_out[118] bl_out[118] br_out[118] data_out[119] bl_out[119] br_out[119] data_out[120] bl_out[120] br_out[120] data_out[121] bl_out[121] br_out[121] data_out[122] bl_out[122] br_out[122] data_out[123] bl_out[123] br_out[123] data_out[124] bl_out[124] br_out[124] data_out[125] bl_out[125] br_out[125] data_out[126] bl_out[126] br_out[126] data_out[127] bl_out[127] br_out[127] gated_s_en vdd gnd sense_amp_array
Xwrite_driver_array data_in[0] data_in[1] data_in[2] data_in[3] data_in[4] data_in[5] data_in[6] data_in[7] data_in[8] data_in[9] data_in[10] data_in[11] data_in[12] data_in[13] data_in[14] data_in[15] data_in[16] data_in[17] data_in[18] data_in[19] data_in[20] data_in[21] data_in[22] data_in[23] data_in[24] data_in[25] data_in[26] data_in[27] data_in[28] data_in[29] data_in[30] data_in[31] data_in[32] data_in[33] data_in[34] data_in[35] data_in[36] data_in[37] data_in[38] data_in[39] data_in[40] data_in[41] data_in[42] data_in[43] data_in[44] data_in[45] data_in[46] data_in[47] data_in[48] data_in[49] data_in[50] data_in[51] data_in[52] data_in[53] data_in[54] data_in[55] data_in[56] data_in[57] data_in[58] data_in[59] data_in[60] data_in[61] data_in[62] data_in[63] data_in[64] data_in[65] data_in[66] data_in[67] data_in[68] data_in[69] data_in[70] data_in[71] data_in[72] data_in[73] data_in[74] data_in[75] data_in[76] data_in[77] data_in[78] data_in[79] data_in[80] data_in[81] data_in[82] data_in[83] data_in[84] data_in[85] data_in[86] data_in[87] data_in[88] data_in[89] data_in[90] data_in[91] data_in[92] data_in[93] data_in[94] data_in[95] data_in[96] data_in[97] data_in[98] data_in[99] data_in[100] data_in[101] data_in[102] data_in[103] data_in[104] data_in[105] data_in[106] data_in[107] data_in[108] data_in[109] data_in[110] data_in[111] data_in[112] data_in[113] data_in[114] data_in[115] data_in[116] data_in[117] data_in[118] data_in[119] data_in[120] data_in[121] data_in[122] data_in[123] data_in[124] data_in[125] data_in[126] data_in[127] bl_out[0] br_out[0] bl_out[1] br_out[1] bl_out[2] br_out[2] bl_out[3] br_out[3] bl_out[4] br_out[4] bl_out[5] br_out[5] bl_out[6] br_out[6] bl_out[7] br_out[7] bl_out[8] br_out[8] bl_out[9] br_out[9] bl_out[10] br_out[10] bl_out[11] br_out[11] bl_out[12] br_out[12] bl_out[13] br_out[13] bl_out[14] br_out[14] bl_out[15] br_out[15] bl_out[16] br_out[16] bl_out[17] br_out[17] bl_out[18] br_out[18] bl_out[19] br_out[19] bl_out[20] br_out[20] bl_out[21] br_out[21] bl_out[22] br_out[22] bl_out[23] br_out[23] bl_out[24] br_out[24] bl_out[25] br_out[25] bl_out[26] br_out[26] bl_out[27] br_out[27] bl_out[28] br_out[28] bl_out[29] br_out[29] bl_out[30] br_out[30] bl_out[31] br_out[31] bl_out[32] br_out[32] bl_out[33] br_out[33] bl_out[34] br_out[34] bl_out[35] br_out[35] bl_out[36] br_out[36] bl_out[37] br_out[37] bl_out[38] br_out[38] bl_out[39] br_out[39] bl_out[40] br_out[40] bl_out[41] br_out[41] bl_out[42] br_out[42] bl_out[43] br_out[43] bl_out[44] br_out[44] bl_out[45] br_out[45] bl_out[46] br_out[46] bl_out[47] br_out[47] bl_out[48] br_out[48] bl_out[49] br_out[49] bl_out[50] br_out[50] bl_out[51] br_out[51] bl_out[52] br_out[52] bl_out[53] br_out[53] bl_out[54] br_out[54] bl_out[55] br_out[55] bl_out[56] br_out[56] bl_out[57] br_out[57] bl_out[58] br_out[58] bl_out[59] br_out[59] bl_out[60] br_out[60] bl_out[61] br_out[61] bl_out[62] br_out[62] bl_out[63] br_out[63] bl_out[64] br_out[64] bl_out[65] br_out[65] bl_out[66] br_out[66] bl_out[67] br_out[67] bl_out[68] br_out[68] bl_out[69] br_out[69] bl_out[70] br_out[70] bl_out[71] br_out[71] bl_out[72] br_out[72] bl_out[73] br_out[73] bl_out[74] br_out[74] bl_out[75] br_out[75] bl_out[76] br_out[76] bl_out[77] br_out[77] bl_out[78] br_out[78] bl_out[79] br_out[79] bl_out[80] br_out[80] bl_out[81] br_out[81] bl_out[82] br_out[82] bl_out[83] br_out[83] bl_out[84] br_out[84] bl_out[85] br_out[85] bl_out[86] br_out[86] bl_out[87] br_out[87] bl_out[88] br_out[88] bl_out[89] br_out[89] bl_out[90] br_out[90] bl_out[91] br_out[91] bl_out[92] br_out[92] bl_out[93] br_out[93] bl_out[94] br_out[94] bl_out[95] br_out[95] bl_out[96] br_out[96] bl_out[97] br_out[97] bl_out[98] br_out[98] bl_out[99] br_out[99] bl_out[100] br_out[100] bl_out[101] br_out[101] bl_out[102] br_out[102] bl_out[103] br_out[103] bl_out[104] br_out[104] bl_out[105] br_out[105] bl_out[106] br_out[106] bl_out[107] br_out[107] bl_out[108] br_out[108] bl_out[109] br_out[109] bl_out[110] br_out[110] bl_out[111] br_out[111] bl_out[112] br_out[112] bl_out[113] br_out[113] bl_out[114] br_out[114] bl_out[115] br_out[115] bl_out[116] br_out[116] bl_out[117] br_out[117] bl_out[118] br_out[118] bl_out[119] br_out[119] bl_out[120] br_out[120] bl_out[121] br_out[121] bl_out[122] br_out[122] bl_out[123] br_out[123] bl_out[124] br_out[124] bl_out[125] br_out[125] bl_out[126] br_out[126] bl_out[127] br_out[127] gated_w_en vdd gnd write_driver_array
Xdata_in_flop_array DATA[0] DATA[1] DATA[2] DATA[3] DATA[4] DATA[5] DATA[6] DATA[7] DATA[8] DATA[9] DATA[10] DATA[11] DATA[12] DATA[13] DATA[14] DATA[15] DATA[16] DATA[17] DATA[18] DATA[19] DATA[20] DATA[21] DATA[22] DATA[23] DATA[24] DATA[25] DATA[26] DATA[27] DATA[28] DATA[29] DATA[30] DATA[31] DATA[32] DATA[33] DATA[34] DATA[35] DATA[36] DATA[37] DATA[38] DATA[39] DATA[40] DATA[41] DATA[42] DATA[43] DATA[44] DATA[45] DATA[46] DATA[47] DATA[48] DATA[49] DATA[50] DATA[51] DATA[52] DATA[53] DATA[54] DATA[55] DATA[56] DATA[57] DATA[58] DATA[59] DATA[60] DATA[61] DATA[62] DATA[63] DATA[64] DATA[65] DATA[66] DATA[67] DATA[68] DATA[69] DATA[70] DATA[71] DATA[72] DATA[73] DATA[74] DATA[75] DATA[76] DATA[77] DATA[78] DATA[79] DATA[80] DATA[81] DATA[82] DATA[83] DATA[84] DATA[85] DATA[86] DATA[87] DATA[88] DATA[89] DATA[90] DATA[91] DATA[92] DATA[93] DATA[94] DATA[95] DATA[96] DATA[97] DATA[98] DATA[99] DATA[100] DATA[101] DATA[102] DATA[103] DATA[104] DATA[105] DATA[106] DATA[107] DATA[108] DATA[109] DATA[110] DATA[111] DATA[112] DATA[113] DATA[114] DATA[115] DATA[116] DATA[117] DATA[118] DATA[119] DATA[120] DATA[121] DATA[122] DATA[123] DATA[124] DATA[125] DATA[126] DATA[127] data_in[0] data_in_bar[0] data_in[1] data_in_bar[1] data_in[2] data_in_bar[2] data_in[3] data_in_bar[3] data_in[4] data_in_bar[4] data_in[5] data_in_bar[5] data_in[6] data_in_bar[6] data_in[7] data_in_bar[7] data_in[8] data_in_bar[8] data_in[9] data_in_bar[9] data_in[10] data_in_bar[10] data_in[11] data_in_bar[11] data_in[12] data_in_bar[12] data_in[13] data_in_bar[13] data_in[14] data_in_bar[14] data_in[15] data_in_bar[15] data_in[16] data_in_bar[16] data_in[17] data_in_bar[17] data_in[18] data_in_bar[18] data_in[19] data_in_bar[19] data_in[20] data_in_bar[20] data_in[21] data_in_bar[21] data_in[22] data_in_bar[22] data_in[23] data_in_bar[23] data_in[24] data_in_bar[24] data_in[25] data_in_bar[25] data_in[26] data_in_bar[26] data_in[27] data_in_bar[27] data_in[28] data_in_bar[28] data_in[29] data_in_bar[29] data_in[30] data_in_bar[30] data_in[31] data_in_bar[31] data_in[32] data_in_bar[32] data_in[33] data_in_bar[33] data_in[34] data_in_bar[34] data_in[35] data_in_bar[35] data_in[36] data_in_bar[36] data_in[37] data_in_bar[37] data_in[38] data_in_bar[38] data_in[39] data_in_bar[39] data_in[40] data_in_bar[40] data_in[41] data_in_bar[41] data_in[42] data_in_bar[42] data_in[43] data_in_bar[43] data_in[44] data_in_bar[44] data_in[45] data_in_bar[45] data_in[46] data_in_bar[46] data_in[47] data_in_bar[47] data_in[48] data_in_bar[48] data_in[49] data_in_bar[49] data_in[50] data_in_bar[50] data_in[51] data_in_bar[51] data_in[52] data_in_bar[52] data_in[53] data_in_bar[53] data_in[54] data_in_bar[54] data_in[55] data_in_bar[55] data_in[56] data_in_bar[56] data_in[57] data_in_bar[57] data_in[58] data_in_bar[58] data_in[59] data_in_bar[59] data_in[60] data_in_bar[60] data_in[61] data_in_bar[61] data_in[62] data_in_bar[62] data_in[63] data_in_bar[63] data_in[64] data_in_bar[64] data_in[65] data_in_bar[65] data_in[66] data_in_bar[66] data_in[67] data_in_bar[67] data_in[68] data_in_bar[68] data_in[69] data_in_bar[69] data_in[70] data_in_bar[70] data_in[71] data_in_bar[71] data_in[72] data_in_bar[72] data_in[73] data_in_bar[73] data_in[74] data_in_bar[74] data_in[75] data_in_bar[75] data_in[76] data_in_bar[76] data_in[77] data_in_bar[77] data_in[78] data_in_bar[78] data_in[79] data_in_bar[79] data_in[80] data_in_bar[80] data_in[81] data_in_bar[81] data_in[82] data_in_bar[82] data_in[83] data_in_bar[83] data_in[84] data_in_bar[84] data_in[85] data_in_bar[85] data_in[86] data_in_bar[86] data_in[87] data_in_bar[87] data_in[88] data_in_bar[88] data_in[89] data_in_bar[89] data_in[90] data_in_bar[90] data_in[91] data_in_bar[91] data_in[92] data_in_bar[92] data_in[93] data_in_bar[93] data_in[94] data_in_bar[94] data_in[95] data_in_bar[95] data_in[96] data_in_bar[96] data_in[97] data_in_bar[97] data_in[98] data_in_bar[98] data_in[99] data_in_bar[99] data_in[100] data_in_bar[100] data_in[101] data_in_bar[101] data_in[102] data_in_bar[102] data_in[103] data_in_bar[103] data_in[104] data_in_bar[104] data_in[105] data_in_bar[105] data_in[106] data_in_bar[106] data_in[107] data_in_bar[107] data_in[108] data_in_bar[108] data_in[109] data_in_bar[109] data_in[110] data_in_bar[110] data_in[111] data_in_bar[111] data_in[112] data_in_bar[112] data_in[113] data_in_bar[113] data_in[114] data_in_bar[114] data_in[115] data_in_bar[115] data_in[116] data_in_bar[116] data_in[117] data_in_bar[117] data_in[118] data_in_bar[118] data_in[119] data_in_bar[119] data_in[120] data_in_bar[120] data_in[121] data_in_bar[121] data_in[122] data_in_bar[122] data_in[123] data_in_bar[123] data_in[124] data_in_bar[124] data_in[125] data_in_bar[125] data_in[126] data_in_bar[126] data_in[127] data_in_bar[127] gated_clk_bar vdd gnd msf_data_in
Xtri_gate_array data_out[0] data_out[1] data_out[2] data_out[3] data_out[4] data_out[5] data_out[6] data_out[7] data_out[8] data_out[9] data_out[10] data_out[11] data_out[12] data_out[13] data_out[14] data_out[15] data_out[16] data_out[17] data_out[18] data_out[19] data_out[20] data_out[21] data_out[22] data_out[23] data_out[24] data_out[25] data_out[26] data_out[27] data_out[28] data_out[29] data_out[30] data_out[31] data_out[32] data_out[33] data_out[34] data_out[35] data_out[36] data_out[37] data_out[38] data_out[39] data_out[40] data_out[41] data_out[42] data_out[43] data_out[44] data_out[45] data_out[46] data_out[47] data_out[48] data_out[49] data_out[50] data_out[51] data_out[52] data_out[53] data_out[54] data_out[55] data_out[56] data_out[57] data_out[58] data_out[59] data_out[60] data_out[61] data_out[62] data_out[63] data_out[64] data_out[65] data_out[66] data_out[67] data_out[68] data_out[69] data_out[70] data_out[71] data_out[72] data_out[73] data_out[74] data_out[75] data_out[76] data_out[77] data_out[78] data_out[79] data_out[80] data_out[81] data_out[82] data_out[83] data_out[84] data_out[85] data_out[86] data_out[87] data_out[88] data_out[89] data_out[90] data_out[91] data_out[92] data_out[93] data_out[94] data_out[95] data_out[96] data_out[97] data_out[98] data_out[99] data_out[100] data_out[101] data_out[102] data_out[103] data_out[104] data_out[105] data_out[106] data_out[107] data_out[108] data_out[109] data_out[110] data_out[111] data_out[112] data_out[113] data_out[114] data_out[115] data_out[116] data_out[117] data_out[118] data_out[119] data_out[120] data_out[121] data_out[122] data_out[123] data_out[124] data_out[125] data_out[126] data_out[127] DATA[0] DATA[1] DATA[2] DATA[3] DATA[4] DATA[5] DATA[6] DATA[7] DATA[8] DATA[9] DATA[10] DATA[11] DATA[12] DATA[13] DATA[14] DATA[15] DATA[16] DATA[17] DATA[18] DATA[19] DATA[20] DATA[21] DATA[22] DATA[23] DATA[24] DATA[25] DATA[26] DATA[27] DATA[28] DATA[29] DATA[30] DATA[31] DATA[32] DATA[33] DATA[34] DATA[35] DATA[36] DATA[37] DATA[38] DATA[39] DATA[40] DATA[41] DATA[42] DATA[43] DATA[44] DATA[45] DATA[46] DATA[47] DATA[48] DATA[49] DATA[50] DATA[51] DATA[52] DATA[53] DATA[54] DATA[55] DATA[56] DATA[57] DATA[58] DATA[59] DATA[60] DATA[61] DATA[62] DATA[63] DATA[64] DATA[65] DATA[66] DATA[67] DATA[68] DATA[69] DATA[70] DATA[71] DATA[72] DATA[73] DATA[74] DATA[75] DATA[76] DATA[77] DATA[78] DATA[79] DATA[80] DATA[81] DATA[82] DATA[83] DATA[84] DATA[85] DATA[86] DATA[87] DATA[88] DATA[89] DATA[90] DATA[91] DATA[92] DATA[93] DATA[94] DATA[95] DATA[96] DATA[97] DATA[98] DATA[99] DATA[100] DATA[101] DATA[102] DATA[103] DATA[104] DATA[105] DATA[106] DATA[107] DATA[108] DATA[109] DATA[110] DATA[111] DATA[112] DATA[113] DATA[114] DATA[115] DATA[116] DATA[117] DATA[118] DATA[119] DATA[120] DATA[121] DATA[122] DATA[123] DATA[124] DATA[125] DATA[126] DATA[127] gated_tri_en gated_tri_en_bar vdd gnd tri_gate_array
Xrow_decoder A[0] A[1] A[2] A[3] A[4] A[5] A[6] dec_out[0] dec_out[1] dec_out[2] dec_out[3] dec_out[4] dec_out[5] dec_out[6] dec_out[7] dec_out[8] dec_out[9] dec_out[10] dec_out[11] dec_out[12] dec_out[13] dec_out[14] dec_out[15] dec_out[16] dec_out[17] dec_out[18] dec_out[19] dec_out[20] dec_out[21] dec_out[22] dec_out[23] dec_out[24] dec_out[25] dec_out[26] dec_out[27] dec_out[28] dec_out[29] dec_out[30] dec_out[31] dec_out[32] dec_out[33] dec_out[34] dec_out[35] dec_out[36] dec_out[37] dec_out[38] dec_out[39] dec_out[40] dec_out[41] dec_out[42] dec_out[43] dec_out[44] dec_out[45] dec_out[46] dec_out[47] dec_out[48] dec_out[49] dec_out[50] dec_out[51] dec_out[52] dec_out[53] dec_out[54] dec_out[55] dec_out[56] dec_out[57] dec_out[58] dec_out[59] dec_out[60] dec_out[61] dec_out[62] dec_out[63] dec_out[64] dec_out[65] dec_out[66] dec_out[67] dec_out[68] dec_out[69] dec_out[70] dec_out[71] dec_out[72] dec_out[73] dec_out[74] dec_out[75] dec_out[76] dec_out[77] dec_out[78] dec_out[79] dec_out[80] dec_out[81] dec_out[82] dec_out[83] dec_out[84] dec_out[85] dec_out[86] dec_out[87] dec_out[88] dec_out[89] dec_out[90] dec_out[91] dec_out[92] dec_out[93] dec_out[94] dec_out[95] dec_out[96] dec_out[97] dec_out[98] dec_out[99] dec_out[100] dec_out[101] dec_out[102] dec_out[103] dec_out[104] dec_out[105] dec_out[106] dec_out[107] dec_out[108] dec_out[109] dec_out[110] dec_out[111] dec_out[112] dec_out[113] dec_out[114] dec_out[115] dec_out[116] dec_out[117] dec_out[118] dec_out[119] dec_out[120] dec_out[121] dec_out[122] dec_out[123] dec_out[124] dec_out[125] dec_out[126] dec_out[127] vdd gnd hierarchical_decoder_128rows
Xwordline_driver dec_out[0] dec_out[1] dec_out[2] dec_out[3] dec_out[4] dec_out[5] dec_out[6] dec_out[7] dec_out[8] dec_out[9] dec_out[10] dec_out[11] dec_out[12] dec_out[13] dec_out[14] dec_out[15] dec_out[16] dec_out[17] dec_out[18] dec_out[19] dec_out[20] dec_out[21] dec_out[22] dec_out[23] dec_out[24] dec_out[25] dec_out[26] dec_out[27] dec_out[28] dec_out[29] dec_out[30] dec_out[31] dec_out[32] dec_out[33] dec_out[34] dec_out[35] dec_out[36] dec_out[37] dec_out[38] dec_out[39] dec_out[40] dec_out[41] dec_out[42] dec_out[43] dec_out[44] dec_out[45] dec_out[46] dec_out[47] dec_out[48] dec_out[49] dec_out[50] dec_out[51] dec_out[52] dec_out[53] dec_out[54] dec_out[55] dec_out[56] dec_out[57] dec_out[58] dec_out[59] dec_out[60] dec_out[61] dec_out[62] dec_out[63] dec_out[64] dec_out[65] dec_out[66] dec_out[67] dec_out[68] dec_out[69] dec_out[70] dec_out[71] dec_out[72] dec_out[73] dec_out[74] dec_out[75] dec_out[76] dec_out[77] dec_out[78] dec_out[79] dec_out[80] dec_out[81] dec_out[82] dec_out[83] dec_out[84] dec_out[85] dec_out[86] dec_out[87] dec_out[88] dec_out[89] dec_out[90] dec_out[91] dec_out[92] dec_out[93] dec_out[94] dec_out[95] dec_out[96] dec_out[97] dec_out[98] dec_out[99] dec_out[100] dec_out[101] dec_out[102] dec_out[103] dec_out[104] dec_out[105] dec_out[106] dec_out[107] dec_out[108] dec_out[109] dec_out[110] dec_out[111] dec_out[112] dec_out[113] dec_out[114] dec_out[115] dec_out[116] dec_out[117] dec_out[118] dec_out[119] dec_out[120] dec_out[121] dec_out[122] dec_out[123] dec_out[124] dec_out[125] dec_out[126] dec_out[127] wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55] wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63] wl[64] wl[65] wl[66] wl[67] wl[68] wl[69] wl[70] wl[71] wl[72] wl[73] wl[74] wl[75] wl[76] wl[77] wl[78] wl[79] wl[80] wl[81] wl[82] wl[83] wl[84] wl[85] wl[86] wl[87] wl[88] wl[89] wl[90] wl[91] wl[92] wl[93] wl[94] wl[95] wl[96] wl[97] wl[98] wl[99] wl[100] wl[101] wl[102] wl[103] wl[104] wl[105] wl[106] wl[107] wl[108] wl[109] wl[110] wl[111] wl[112] wl[113] wl[114] wl[115] wl[116] wl[117] wl[118] wl[119] wl[120] wl[121] wl[122] wl[123] wl[124] wl[125] wl[126] wl[127] gated_clk_buf vdd gnd wordline_driver
Xaddress_flop_array ADDR[0] ADDR[1] ADDR[2] ADDR[3] ADDR[4] ADDR[5] ADDR[6] ADDR[7] A[0] A_bar[0] A[1] A_bar[1] A[2] A_bar[2] A[3] A_bar[3] A[4] A_bar[4] A[5] A_bar[5] A[6] A_bar[6] sel[1] sel[0] gated_clk_buf vdd gnd msf_address
Xbank_sel_inv bank_sel bank_sel_bar vdd gnd pinv_13
Xnor_clk_buf clk_buf bank_sel_bar gated_clk_buf_temp_bar vdd gnd pnor2_2
Xinv_clk_buf gated_clk_buf_temp_bar gated_clk_buf vdd gnd pinv_14
Xnor_tri_en_bar tri_en_bar bank_sel_bar gated_tri_en_bar_temp_bar vdd gnd pnor2_2
Xinv_tri_en_bar gated_tri_en_bar_temp_bar gated_tri_en_bar vdd gnd pinv_14
Xnand_tri_en tri_en bank_sel gated_tri_en_temp_bar vdd gnd pnand2_5
Xinv_tri_en gated_tri_en_temp_bar gated_tri_en vdd gnd pinv_14
Xnand_clk_bar clk_bar bank_sel gated_clk_bar_temp_bar vdd gnd pnand2_5
Xinv_clk_bar gated_clk_bar_temp_bar gated_clk_bar vdd gnd pinv_14
Xnand_w_en w_en bank_sel gated_w_en_temp_bar vdd gnd pnand2_5
Xinv_w_en gated_w_en_temp_bar gated_w_en vdd gnd pinv_14
Xnand_s_en s_en bank_sel gated_s_en_temp_bar vdd gnd pnand2_5
Xinv_s_en gated_s_en_temp_bar gated_s_en vdd gnd pinv_14
.ENDS bank

.SUBCKT msb_address din[0] din[1] dout[0] dout_bar[0] dout[1] dout_bar[1] clk vdd gnd
XXdff0 din[0] dout[0] dout_bar[0] clk vdd gnd ms_flop
XXdff1 din[1] dout[1] dout_bar[1] clk vdd gnd ms_flop
.ENDS msb_address

.SUBCKT sram_1rw_128b_1024w_4bank_scn3me_subm DATA[0] DATA[1] DATA[2] DATA[3] DATA[4] DATA[5] DATA[6] DATA[7] DATA[8] DATA[9] DATA[10] DATA[11] DATA[12] DATA[13] DATA[14] DATA[15] DATA[16] DATA[17] DATA[18] DATA[19] DATA[20] DATA[21] DATA[22] DATA[23] DATA[24] DATA[25] DATA[26] DATA[27] DATA[28] DATA[29] DATA[30] DATA[31] DATA[32] DATA[33] DATA[34] DATA[35] DATA[36] DATA[37] DATA[38] DATA[39] DATA[40] DATA[41] DATA[42] DATA[43] DATA[44] DATA[45] DATA[46] DATA[47] DATA[48] DATA[49] DATA[50] DATA[51] DATA[52] DATA[53] DATA[54] DATA[55] DATA[56] DATA[57] DATA[58] DATA[59] DATA[60] DATA[61] DATA[62] DATA[63] DATA[64] DATA[65] DATA[66] DATA[67] DATA[68] DATA[69] DATA[70] DATA[71] DATA[72] DATA[73] DATA[74] DATA[75] DATA[76] DATA[77] DATA[78] DATA[79] DATA[80] DATA[81] DATA[82] DATA[83] DATA[84] DATA[85] DATA[86] DATA[87] DATA[88] DATA[89] DATA[90] DATA[91] DATA[92] DATA[93] DATA[94] DATA[95] DATA[96] DATA[97] DATA[98] DATA[99] DATA[100] DATA[101] DATA[102] DATA[103] DATA[104] DATA[105] DATA[106] DATA[107] DATA[108] DATA[109] DATA[110] DATA[111] DATA[112] DATA[113] DATA[114] DATA[115] DATA[116] DATA[117] DATA[118] DATA[119] DATA[120] DATA[121] DATA[122] DATA[123] DATA[124] DATA[125] DATA[126] DATA[127] ADDR[0] ADDR[1] ADDR[2] ADDR[3] ADDR[4] ADDR[5] ADDR[6] ADDR[7] ADDR[8] ADDR[9] CSb WEb OEb clk vdd gnd
Xbank0 DATA[0] DATA[1] DATA[2] DATA[3] DATA[4] DATA[5] DATA[6] DATA[7] DATA[8] DATA[9] DATA[10] DATA[11] DATA[12] DATA[13] DATA[14] DATA[15] DATA[16] DATA[17] DATA[18] DATA[19] DATA[20] DATA[21] DATA[22] DATA[23] DATA[24] DATA[25] DATA[26] DATA[27] DATA[28] DATA[29] DATA[30] DATA[31] DATA[32] DATA[33] DATA[34] DATA[35] DATA[36] DATA[37] DATA[38] DATA[39] DATA[40] DATA[41] DATA[42] DATA[43] DATA[44] DATA[45] DATA[46] DATA[47] DATA[48] DATA[49] DATA[50] DATA[51] DATA[52] DATA[53] DATA[54] DATA[55] DATA[56] DATA[57] DATA[58] DATA[59] DATA[60] DATA[61] DATA[62] DATA[63] DATA[64] DATA[65] DATA[66] DATA[67] DATA[68] DATA[69] DATA[70] DATA[71] DATA[72] DATA[73] DATA[74] DATA[75] DATA[76] DATA[77] DATA[78] DATA[79] DATA[80] DATA[81] DATA[82] DATA[83] DATA[84] DATA[85] DATA[86] DATA[87] DATA[88] DATA[89] DATA[90] DATA[91] DATA[92] DATA[93] DATA[94] DATA[95] DATA[96] DATA[97] DATA[98] DATA[99] DATA[100] DATA[101] DATA[102] DATA[103] DATA[104] DATA[105] DATA[106] DATA[107] DATA[108] DATA[109] DATA[110] DATA[111] DATA[112] DATA[113] DATA[114] DATA[115] DATA[116] DATA[117] DATA[118] DATA[119] DATA[120] DATA[121] DATA[122] DATA[123] DATA[124] DATA[125] DATA[126] DATA[127] ADDR[0] ADDR[1] ADDR[2] ADDR[3] ADDR[4] ADDR[5] ADDR[6] ADDR[7] bank_sel[0] s_en w_en tri_en_bar tri_en clk_bar clk_buf vdd gnd bank
Xbank1 DATA[0] DATA[1] DATA[2] DATA[3] DATA[4] DATA[5] DATA[6] DATA[7] DATA[8] DATA[9] DATA[10] DATA[11] DATA[12] DATA[13] DATA[14] DATA[15] DATA[16] DATA[17] DATA[18] DATA[19] DATA[20] DATA[21] DATA[22] DATA[23] DATA[24] DATA[25] DATA[26] DATA[27] DATA[28] DATA[29] DATA[30] DATA[31] DATA[32] DATA[33] DATA[34] DATA[35] DATA[36] DATA[37] DATA[38] DATA[39] DATA[40] DATA[41] DATA[42] DATA[43] DATA[44] DATA[45] DATA[46] DATA[47] DATA[48] DATA[49] DATA[50] DATA[51] DATA[52] DATA[53] DATA[54] DATA[55] DATA[56] DATA[57] DATA[58] DATA[59] DATA[60] DATA[61] DATA[62] DATA[63] DATA[64] DATA[65] DATA[66] DATA[67] DATA[68] DATA[69] DATA[70] DATA[71] DATA[72] DATA[73] DATA[74] DATA[75] DATA[76] DATA[77] DATA[78] DATA[79] DATA[80] DATA[81] DATA[82] DATA[83] DATA[84] DATA[85] DATA[86] DATA[87] DATA[88] DATA[89] DATA[90] DATA[91] DATA[92] DATA[93] DATA[94] DATA[95] DATA[96] DATA[97] DATA[98] DATA[99] DATA[100] DATA[101] DATA[102] DATA[103] DATA[104] DATA[105] DATA[106] DATA[107] DATA[108] DATA[109] DATA[110] DATA[111] DATA[112] DATA[113] DATA[114] DATA[115] DATA[116] DATA[117] DATA[118] DATA[119] DATA[120] DATA[121] DATA[122] DATA[123] DATA[124] DATA[125] DATA[126] DATA[127] ADDR[0] ADDR[1] ADDR[2] ADDR[3] ADDR[4] ADDR[5] ADDR[6] ADDR[7] bank_sel[1] s_en w_en tri_en_bar tri_en clk_bar clk_buf vdd gnd bank
Xbank2 DATA[0] DATA[1] DATA[2] DATA[3] DATA[4] DATA[5] DATA[6] DATA[7] DATA[8] DATA[9] DATA[10] DATA[11] DATA[12] DATA[13] DATA[14] DATA[15] DATA[16] DATA[17] DATA[18] DATA[19] DATA[20] DATA[21] DATA[22] DATA[23] DATA[24] DATA[25] DATA[26] DATA[27] DATA[28] DATA[29] DATA[30] DATA[31] DATA[32] DATA[33] DATA[34] DATA[35] DATA[36] DATA[37] DATA[38] DATA[39] DATA[40] DATA[41] DATA[42] DATA[43] DATA[44] DATA[45] DATA[46] DATA[47] DATA[48] DATA[49] DATA[50] DATA[51] DATA[52] DATA[53] DATA[54] DATA[55] DATA[56] DATA[57] DATA[58] DATA[59] DATA[60] DATA[61] DATA[62] DATA[63] DATA[64] DATA[65] DATA[66] DATA[67] DATA[68] DATA[69] DATA[70] DATA[71] DATA[72] DATA[73] DATA[74] DATA[75] DATA[76] DATA[77] DATA[78] DATA[79] DATA[80] DATA[81] DATA[82] DATA[83] DATA[84] DATA[85] DATA[86] DATA[87] DATA[88] DATA[89] DATA[90] DATA[91] DATA[92] DATA[93] DATA[94] DATA[95] DATA[96] DATA[97] DATA[98] DATA[99] DATA[100] DATA[101] DATA[102] DATA[103] DATA[104] DATA[105] DATA[106] DATA[107] DATA[108] DATA[109] DATA[110] DATA[111] DATA[112] DATA[113] DATA[114] DATA[115] DATA[116] DATA[117] DATA[118] DATA[119] DATA[120] DATA[121] DATA[122] DATA[123] DATA[124] DATA[125] DATA[126] DATA[127] ADDR[0] ADDR[1] ADDR[2] ADDR[3] ADDR[4] ADDR[5] ADDR[6] ADDR[7] bank_sel[2] s_en w_en tri_en_bar tri_en clk_bar clk_buf vdd gnd bank
Xbank3 DATA[0] DATA[1] DATA[2] DATA[3] DATA[4] DATA[5] DATA[6] DATA[7] DATA[8] DATA[9] DATA[10] DATA[11] DATA[12] DATA[13] DATA[14] DATA[15] DATA[16] DATA[17] DATA[18] DATA[19] DATA[20] DATA[21] DATA[22] DATA[23] DATA[24] DATA[25] DATA[26] DATA[27] DATA[28] DATA[29] DATA[30] DATA[31] DATA[32] DATA[33] DATA[34] DATA[35] DATA[36] DATA[37] DATA[38] DATA[39] DATA[40] DATA[41] DATA[42] DATA[43] DATA[44] DATA[45] DATA[46] DATA[47] DATA[48] DATA[49] DATA[50] DATA[51] DATA[52] DATA[53] DATA[54] DATA[55] DATA[56] DATA[57] DATA[58] DATA[59] DATA[60] DATA[61] DATA[62] DATA[63] DATA[64] DATA[65] DATA[66] DATA[67] DATA[68] DATA[69] DATA[70] DATA[71] DATA[72] DATA[73] DATA[74] DATA[75] DATA[76] DATA[77] DATA[78] DATA[79] DATA[80] DATA[81] DATA[82] DATA[83] DATA[84] DATA[85] DATA[86] DATA[87] DATA[88] DATA[89] DATA[90] DATA[91] DATA[92] DATA[93] DATA[94] DATA[95] DATA[96] DATA[97] DATA[98] DATA[99] DATA[100] DATA[101] DATA[102] DATA[103] DATA[104] DATA[105] DATA[106] DATA[107] DATA[108] DATA[109] DATA[110] DATA[111] DATA[112] DATA[113] DATA[114] DATA[115] DATA[116] DATA[117] DATA[118] DATA[119] DATA[120] DATA[121] DATA[122] DATA[123] DATA[124] DATA[125] DATA[126] DATA[127] ADDR[0] ADDR[1] ADDR[2] ADDR[3] ADDR[4] ADDR[5] ADDR[6] ADDR[7] bank_sel[3] s_en w_en tri_en_bar tri_en clk_bar clk_buf vdd gnd bank
Xcontrol CSb WEb OEb clk s_en w_en tri_en tri_en_bar clk_bar clk_buf vdd gnd control_logic
Xmsb_address ADDR[8] ADDR[9] msb[0] msb_bar[0] msb[1] msb_bar[1] clk_buf vdd gnd msb_address
Xmsb_decoder msb[0] msb[1] bank_sel[0] bank_sel[1] bank_sel[2] bank_sel[3] vdd gnd pre2x4
.ENDS sram_1rw_128b_1024w_4bank_scn3me_subm
