magic
tech sky130A
magscale 1 2
timestamp 1595931502
<< checkpaint >>
rect -1260 7033 3132 7037
rect -1260 -1022 3168 7033
<< metal1 >>
rect 879 5717 939 5773
rect 1433 5717 1493 5773
rect 624 5655 1872 5683
rect 751 3700 779 3766
rect 751 3672 851 3700
rect 728 3260 774 3514
rect 823 2384 851 3672
rect 953 3620 981 3766
rect 896 3592 981 3620
rect 1391 3620 1419 3766
rect 1593 3700 1621 3766
rect 1521 3672 1621 3700
rect 1391 3592 1476 3620
rect 896 2372 924 3592
rect 1448 2372 1476 3592
rect 1521 2384 1549 3672
rect 1598 3260 1644 3514
rect 823 1192 851 1258
rect 690 1164 851 1192
rect 66 252 94 1006
rect 530 252 558 1006
rect 690 252 718 1164
rect 896 1112 924 1258
rect 1448 1112 1476 1258
rect 1521 1192 1549 1258
rect 1521 1164 1806 1192
rect 896 1084 1182 1112
rect 1154 252 1182 1084
rect 1314 1084 1476 1112
rect 1314 252 1342 1084
rect 1778 252 1806 1164
<< metal3 >>
rect 851 5537 949 5635
rect 1423 5537 1521 5635
rect 837 5121 935 5219
rect 1437 5121 1535 5219
rect 952 4919 1050 5017
rect 1322 4919 1420 5017
rect 831 4587 929 4685
rect 1443 4587 1541 4685
rect 842 4150 940 4248
rect 1432 4150 1530 4248
rect 956 3357 1054 3455
rect 1318 3357 1416 3455
rect 956 3035 1054 3133
rect 1318 3035 1416 3133
rect 944 2197 1042 2295
rect 1330 2197 1428 2295
rect 1026 1423 1124 1521
rect 1248 1423 1346 1521
rect 624 1290 1872 1350
rect 0 951 1872 1011
rect 382 313 480 411
rect 768 313 866 411
rect 1630 313 1728 411
use sense_amp_array  sense_amp_array_0
timestamp 1595931502
transform 1 0 624 0 -1 3514
box -160 0 1284 2256
use write_driver_array  write_driver_array_0
timestamp 1595931502
transform 1 0 624 0 -1 5777
box -152 4 1276 2011
use precharge_array  precharge_array_0
timestamp 1595931502
transform 1 0 0 0 -1 1006
box 0 -12 1872 768
<< labels >>
rlabel metal3 s 1297 1472 1297 1472 4 gnd
rlabel metal3 s 891 4199 891 4199 4 gnd
rlabel metal3 s 1371 4968 1371 4968 4 gnd
rlabel metal3 s 1486 5170 1486 5170 4 gnd
rlabel metal3 s 886 5170 886 5170 4 gnd
rlabel metal3 s 1481 4199 1481 4199 4 gnd
rlabel metal3 s 1367 3406 1367 3406 4 gnd
rlabel metal3 s 1075 1472 1075 1472 4 gnd
rlabel metal3 s 1005 3406 1005 3406 4 gnd
rlabel metal3 s 1001 4968 1001 4968 4 gnd
rlabel metal1 s 751 3387 751 3387 4 dout_0
rlabel metal1 s 909 5745 909 5745 4 din_0
rlabel metal1 s 80 629 80 629 4 rbl_br
rlabel metal1 s 544 629 544 629 4 rbl_bl
rlabel metal3 s 993 2246 993 2246 4 vdd
rlabel metal3 s 1679 362 1679 362 4 vdd
rlabel metal3 s 1492 4636 1492 4636 4 vdd
rlabel metal3 s 1005 3084 1005 3084 4 vdd
rlabel metal3 s 1367 3084 1367 3084 4 vdd
rlabel metal3 s 431 362 431 362 4 vdd
rlabel metal3 s 900 5586 900 5586 4 vdd
rlabel metal3 s 880 4636 880 4636 4 vdd
rlabel metal3 s 817 362 817 362 4 vdd
rlabel metal3 s 1379 2246 1379 2246 4 vdd
rlabel metal3 s 1472 5586 1472 5586 4 vdd
rlabel metal1 s 1248 5669 1248 5669 4 w_en
rlabel metal3 s 1248 1320 1248 1320 4 s_en
rlabel metal1 s 1168 629 1168 629 4 br_0
rlabel metal1 s 1792 629 1792 629 4 bl_1
rlabel metal3 s 936 981 936 981 4 p_en_bar
rlabel metal1 s 1463 5745 1463 5745 4 din_1
rlabel metal1 s 1328 629 1328 629 4 br_1
rlabel metal1 s 1621 3387 1621 3387 4 dout_1
rlabel metal1 s 704 629 704 629 4 bl_0
<< properties >>
string FIXED_BBOX 0 0 1872 5777
<< end >>
