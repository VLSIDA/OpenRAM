magic
tech sky130A
magscale 1 2
timestamp 1595931502
<< checkpaint >>
rect -1309 -1311 3560 4139
<< locali >>
rect 0 2812 2264 2848
rect 0 1396 2264 1432
rect 0 -20 2264 16
<< metal1 >>
rect -32 2804 32 2856
rect -32 1388 32 1440
rect -32 -28 32 24
<< metal2 >>
rect -28 2806 28 2854
rect 137 2238 203 2290
rect -28 1390 28 1438
rect 137 538 203 590
rect -28 -26 28 22
rect 369 0 397 2828
rect 2074 2311 2102 2339
rect 1568 1929 1596 1957
rect 1568 871 1596 899
rect 2074 489 2102 517
<< metal3 >>
rect -49 2781 49 2879
rect -49 1365 49 1463
rect -49 -51 49 47
use contact_9  contact_9_3
timestamp 1595931502
transform 1 0 -33 0 1 1377
box 0 0 66 74
use contact_9  contact_9_2
timestamp 1595931502
transform 1 0 -33 0 1 -39
box 0 0 66 74
use contact_9  contact_9_1
timestamp 1595931502
transform 1 0 -33 0 1 1377
box 0 0 66 74
use contact_9  contact_9_0
timestamp 1595931502
transform 1 0 -33 0 1 2793
box 0 0 66 74
use contact_8  contact_8_3
timestamp 1595931502
transform 1 0 -32 0 1 1382
box 0 0 64 64
use contact_8  contact_8_2
timestamp 1595931502
transform 1 0 -32 0 1 -34
box 0 0 64 64
use contact_8  contact_8_1
timestamp 1595931502
transform 1 0 -32 0 1 1382
box 0 0 64 64
use contact_8  contact_8_0
timestamp 1595931502
transform 1 0 -32 0 1 2798
box 0 0 64 64
use contact_7  contact_7_3
timestamp 1595931502
transform 1 0 -29 0 1 1381
box 0 0 58 66
use contact_7  contact_7_2
timestamp 1595931502
transform 1 0 -29 0 1 -35
box 0 0 58 66
use contact_7  contact_7_1
timestamp 1595931502
transform 1 0 -29 0 1 1381
box 0 0 58 66
use contact_7  contact_7_0
timestamp 1595931502
transform 1 0 -29 0 1 2797
box 0 0 58 66
use dff_buf_0  dff_buf_0_0
timestamp 1595931502
transform 1 0 0 0 -1 2828
box -8 -20 2300 1471
use dff_buf_0  dff_buf_0_1
timestamp 1595931502
transform 1 0 0 0 1 0
box -8 -20 2300 1471
<< labels >>
rlabel metal3 s 0 2830 0 2830 4 gnd
rlabel metal3 s 0 -2 0 -2 4 gnd
rlabel metal2 s 2088 503 2088 503 4 dout_0
rlabel metal2 s 2088 2325 2088 2325 4 dout_1
rlabel metal2 s 170 564 170 564 4 din_0
rlabel metal2 s 170 2264 170 2264 4 din_1
rlabel metal2 s 383 1414 383 1414 4 clk
rlabel metal2 s 1582 1943 1582 1943 4 dout_bar_1
rlabel metal3 s 0 1414 0 1414 4 vdd
rlabel metal2 s 1582 885 1582 885 4 dout_bar_0
<< properties >>
string FIXED_BBOX 0 0 2264 2828
<< end >>
