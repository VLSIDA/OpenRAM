VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  dataBASE MICRONS 1000 ;
END UNITS
SITE  MacroSite
   CLASS Core ;
   SIZE 12145.0 by 43967.5 ;
END  MacroSite
MACRO sram_2_16_1_freepdk45
   CLASS BLOCK ;
   SIZE 12145.0 BY 43967.5 ;
   SYMMETRY X Y R90 ;
   SITE MacroSite ;
   PIN data[0]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  10260.0 67.5 10330.0 207.5 ;
      END
   END data[0]
   PIN data[1]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  10965.0 67.5 11035.0 207.5 ;
      END
   END data[1]
   PIN addr[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  67.5 8370.0 837.5 8440.0 ;
      END
   END addr[0]
   PIN addr[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  67.5 7665.0 837.5 7735.0 ;
      END
   END addr[1]
   PIN addr[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  67.5 6960.0 837.5 7030.0 ;
      END
   END addr[2]
   PIN addr[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  67.5 6255.0 837.5 6325.0 ;
      END
   END addr[3]
   PIN CSb
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  -2987.5 23757.5 -2917.5 23897.5 ;
      END
   END CSb
   PIN WEb
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  -2282.5 23757.5 -2212.5 23897.5 ;
      END
   END WEb
   PIN OEb
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  -3692.5 23757.5 -3622.5 23897.5 ;
      END
   END OEb
   PIN clk
      DIRECTION INPUT ;
      PORT
         LAYER metal1 ;
         RECT  -835.0 23757.5 -700.0 23947.5 ;
      END
   END clk
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal2 ;
         RECT  452.5 67.5 732.5 44035.0 ;
         LAYER metal2 ;
         RECT  11932.5 67.5 12212.5 44035.0 ;
         LAYER metal1 ;
         RECT  67.5 452.5 12212.5 732.5 ;
         LAYER metal1 ;
         RECT  67.5 43755.0 12212.5 44035.0 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal2 ;
         RECT  67.5 67.5 347.5 44035.0 ;
         LAYER metal2 ;
         RECT  11547.5 67.5 11827.5 44035.0 ;
         LAYER metal1 ;
         RECT  67.5 67.5 12212.5 347.5 ;
         LAYER metal1 ;
         RECT  67.5 43370.0 12212.5 43650.0 ;
      END
   END gnd
   OBS
   LAYER  metal1 ;
      RECT  4657.5 20522.5 4722.5 20587.5 ;
      RECT  4657.5 20250.0 4722.5 20315.0 ;
      RECT  4587.5 20522.5 4690.0 20587.5 ;
      RECT  4657.5 20282.5 4722.5 20555.0 ;
      RECT  4690.0 20250.0 4792.5 20315.0 ;
      RECT  8435.0 20522.5 8500.0 20587.5 ;
      RECT  8435.0 20035.0 8500.0 20100.0 ;
      RECT  7082.5 20522.5 8467.5 20587.5 ;
      RECT  8435.0 20067.5 8500.0 20555.0 ;
      RECT  8467.5 20035.0 9852.5 20100.0 ;
      RECT  4657.5 21957.5 4722.5 22022.5 ;
      RECT  4657.5 22230.0 4722.5 22295.0 ;
      RECT  4587.5 21957.5 4690.0 22022.5 ;
      RECT  4657.5 21990.0 4722.5 22262.5 ;
      RECT  4690.0 22230.0 4792.5 22295.0 ;
      RECT  8435.0 21957.5 8500.0 22022.5 ;
      RECT  8435.0 22445.0 8500.0 22510.0 ;
      RECT  7082.5 21957.5 8467.5 22022.5 ;
      RECT  8435.0 21990.0 8500.0 22477.5 ;
      RECT  8467.5 22445.0 9852.5 22510.0 ;
      RECT  4657.5 23212.5 4722.5 23277.5 ;
      RECT  4657.5 22940.0 4722.5 23005.0 ;
      RECT  4587.5 23212.5 4690.0 23277.5 ;
      RECT  4657.5 22972.5 4722.5 23245.0 ;
      RECT  4690.0 22940.0 4792.5 23005.0 ;
      RECT  8435.0 23212.5 8500.0 23277.5 ;
      RECT  8435.0 22725.0 8500.0 22790.0 ;
      RECT  7082.5 23212.5 8467.5 23277.5 ;
      RECT  8435.0 22757.5 8500.0 23245.0 ;
      RECT  8467.5 22725.0 9852.5 22790.0 ;
      RECT  4657.5 24647.5 4722.5 24712.5 ;
      RECT  4657.5 24920.0 4722.5 24985.0 ;
      RECT  4587.5 24647.5 4690.0 24712.5 ;
      RECT  4657.5 24680.0 4722.5 24952.5 ;
      RECT  4690.0 24920.0 4792.5 24985.0 ;
      RECT  8435.0 24647.5 8500.0 24712.5 ;
      RECT  8435.0 25135.0 8500.0 25200.0 ;
      RECT  7082.5 24647.5 8467.5 24712.5 ;
      RECT  8435.0 24680.0 8500.0 25167.5 ;
      RECT  8467.5 25135.0 9852.5 25200.0 ;
      RECT  4657.5 25902.5 4722.5 25967.5 ;
      RECT  4657.5 25630.0 4722.5 25695.0 ;
      RECT  4587.5 25902.5 4690.0 25967.5 ;
      RECT  4657.5 25662.5 4722.5 25935.0 ;
      RECT  4690.0 25630.0 4792.5 25695.0 ;
      RECT  8435.0 25902.5 8500.0 25967.5 ;
      RECT  8435.0 25415.0 8500.0 25480.0 ;
      RECT  7082.5 25902.5 8467.5 25967.5 ;
      RECT  8435.0 25447.5 8500.0 25935.0 ;
      RECT  8467.5 25415.0 9852.5 25480.0 ;
      RECT  4657.5 27337.5 4722.5 27402.5 ;
      RECT  4657.5 27610.0 4722.5 27675.0 ;
      RECT  4587.5 27337.5 4690.0 27402.5 ;
      RECT  4657.5 27370.0 4722.5 27642.5 ;
      RECT  4690.0 27610.0 4792.5 27675.0 ;
      RECT  8435.0 27337.5 8500.0 27402.5 ;
      RECT  8435.0 27825.0 8500.0 27890.0 ;
      RECT  7082.5 27337.5 8467.5 27402.5 ;
      RECT  8435.0 27370.0 8500.0 27857.5 ;
      RECT  8467.5 27825.0 9852.5 27890.0 ;
      RECT  4657.5 28592.5 4722.5 28657.5 ;
      RECT  4657.5 28320.0 4722.5 28385.0 ;
      RECT  4587.5 28592.5 4690.0 28657.5 ;
      RECT  4657.5 28352.5 4722.5 28625.0 ;
      RECT  4690.0 28320.0 4792.5 28385.0 ;
      RECT  8435.0 28592.5 8500.0 28657.5 ;
      RECT  8435.0 28105.0 8500.0 28170.0 ;
      RECT  7082.5 28592.5 8467.5 28657.5 ;
      RECT  8435.0 28137.5 8500.0 28625.0 ;
      RECT  8467.5 28105.0 9852.5 28170.0 ;
      RECT  4657.5 30027.5 4722.5 30092.5 ;
      RECT  4657.5 30300.0 4722.5 30365.0 ;
      RECT  4587.5 30027.5 4690.0 30092.5 ;
      RECT  4657.5 30060.0 4722.5 30332.5 ;
      RECT  4690.0 30300.0 4792.5 30365.0 ;
      RECT  8435.0 30027.5 8500.0 30092.5 ;
      RECT  8435.0 30515.0 8500.0 30580.0 ;
      RECT  7082.5 30027.5 8467.5 30092.5 ;
      RECT  8435.0 30060.0 8500.0 30547.5 ;
      RECT  8467.5 30515.0 9852.5 30580.0 ;
      RECT  4657.5 31282.5 4722.5 31347.5 ;
      RECT  4657.5 31010.0 4722.5 31075.0 ;
      RECT  4587.5 31282.5 4690.0 31347.5 ;
      RECT  4657.5 31042.5 4722.5 31315.0 ;
      RECT  4690.0 31010.0 4792.5 31075.0 ;
      RECT  8435.0 31282.5 8500.0 31347.5 ;
      RECT  8435.0 30795.0 8500.0 30860.0 ;
      RECT  7082.5 31282.5 8467.5 31347.5 ;
      RECT  8435.0 30827.5 8500.0 31315.0 ;
      RECT  8467.5 30795.0 9852.5 30860.0 ;
      RECT  4657.5 32717.5 4722.5 32782.5 ;
      RECT  4657.5 32990.0 4722.5 33055.0 ;
      RECT  4587.5 32717.5 4690.0 32782.5 ;
      RECT  4657.5 32750.0 4722.5 33022.5 ;
      RECT  4690.0 32990.0 4792.5 33055.0 ;
      RECT  8435.0 32717.5 8500.0 32782.5 ;
      RECT  8435.0 33205.0 8500.0 33270.0 ;
      RECT  7082.5 32717.5 8467.5 32782.5 ;
      RECT  8435.0 32750.0 8500.0 33237.5 ;
      RECT  8467.5 33205.0 9852.5 33270.0 ;
      RECT  4657.5 33972.5 4722.5 34037.5 ;
      RECT  4657.5 33700.0 4722.5 33765.0 ;
      RECT  4587.5 33972.5 4690.0 34037.5 ;
      RECT  4657.5 33732.5 4722.5 34005.0 ;
      RECT  4690.0 33700.0 4792.5 33765.0 ;
      RECT  8435.0 33972.5 8500.0 34037.5 ;
      RECT  8435.0 33485.0 8500.0 33550.0 ;
      RECT  7082.5 33972.5 8467.5 34037.5 ;
      RECT  8435.0 33517.5 8500.0 34005.0 ;
      RECT  8467.5 33485.0 9852.5 33550.0 ;
      RECT  4657.5 35407.5 4722.5 35472.5 ;
      RECT  4657.5 35680.0 4722.5 35745.0 ;
      RECT  4587.5 35407.5 4690.0 35472.5 ;
      RECT  4657.5 35440.0 4722.5 35712.5 ;
      RECT  4690.0 35680.0 4792.5 35745.0 ;
      RECT  8435.0 35407.5 8500.0 35472.5 ;
      RECT  8435.0 35895.0 8500.0 35960.0 ;
      RECT  7082.5 35407.5 8467.5 35472.5 ;
      RECT  8435.0 35440.0 8500.0 35927.5 ;
      RECT  8467.5 35895.0 9852.5 35960.0 ;
      RECT  4657.5 36662.5 4722.5 36727.5 ;
      RECT  4657.5 36390.0 4722.5 36455.0 ;
      RECT  4587.5 36662.5 4690.0 36727.5 ;
      RECT  4657.5 36422.5 4722.5 36695.0 ;
      RECT  4690.0 36390.0 4792.5 36455.0 ;
      RECT  8435.0 36662.5 8500.0 36727.5 ;
      RECT  8435.0 36175.0 8500.0 36240.0 ;
      RECT  7082.5 36662.5 8467.5 36727.5 ;
      RECT  8435.0 36207.5 8500.0 36695.0 ;
      RECT  8467.5 36175.0 9852.5 36240.0 ;
      RECT  4657.5 38097.5 4722.5 38162.5 ;
      RECT  4657.5 38370.0 4722.5 38435.0 ;
      RECT  4587.5 38097.5 4690.0 38162.5 ;
      RECT  4657.5 38130.0 4722.5 38402.5 ;
      RECT  4690.0 38370.0 4792.5 38435.0 ;
      RECT  8435.0 38097.5 8500.0 38162.5 ;
      RECT  8435.0 38585.0 8500.0 38650.0 ;
      RECT  7082.5 38097.5 8467.5 38162.5 ;
      RECT  8435.0 38130.0 8500.0 38617.5 ;
      RECT  8467.5 38585.0 9852.5 38650.0 ;
      RECT  4657.5 39352.5 4722.5 39417.5 ;
      RECT  4657.5 39080.0 4722.5 39145.0 ;
      RECT  4587.5 39352.5 4690.0 39417.5 ;
      RECT  4657.5 39112.5 4722.5 39385.0 ;
      RECT  4690.0 39080.0 4792.5 39145.0 ;
      RECT  8435.0 39352.5 8500.0 39417.5 ;
      RECT  8435.0 38865.0 8500.0 38930.0 ;
      RECT  7082.5 39352.5 8467.5 39417.5 ;
      RECT  8435.0 38897.5 8500.0 39385.0 ;
      RECT  8467.5 38865.0 9852.5 38930.0 ;
      RECT  4657.5 40787.5 4722.5 40852.5 ;
      RECT  4657.5 41060.0 4722.5 41125.0 ;
      RECT  4587.5 40787.5 4690.0 40852.5 ;
      RECT  4657.5 40820.0 4722.5 41092.5 ;
      RECT  4690.0 41060.0 4792.5 41125.0 ;
      RECT  8435.0 40787.5 8500.0 40852.5 ;
      RECT  8435.0 41275.0 8500.0 41340.0 ;
      RECT  7082.5 40787.5 8467.5 40852.5 ;
      RECT  8435.0 40820.0 8500.0 41307.5 ;
      RECT  8467.5 41275.0 9852.5 41340.0 ;
      RECT  7277.5 9340.0 7620.0 9405.0 ;
      RECT  7002.5 10685.0 7825.0 10750.0 ;
      RECT  7277.5 14720.0 8030.0 14785.0 ;
      RECT  7002.5 16065.0 8235.0 16130.0 ;
      RECT  207.5 9135.0 7277.5 9200.0 ;
      RECT  207.5 11825.0 7277.5 11890.0 ;
      RECT  207.5 14515.0 7277.5 14580.0 ;
      RECT  207.5 17205.0 7277.5 17270.0 ;
      RECT  592.5 10480.0 7277.5 10545.0 ;
      RECT  592.5 13170.0 7277.5 13235.0 ;
      RECT  592.5 15860.0 7277.5 15925.0 ;
      RECT  592.5 18550.0 7277.5 18615.0 ;
      RECT  7277.5 8372.5 7620.0 8437.5 ;
      RECT  7277.5 7667.5 7825.0 7732.5 ;
      RECT  7277.5 6962.5 8030.0 7027.5 ;
      RECT  7277.5 6257.5 8235.0 6322.5 ;
      RECT  207.5 8725.0 837.5 8790.0 ;
      RECT  207.5 8020.0 837.5 8085.0 ;
      RECT  207.5 7315.0 837.5 7380.0 ;
      RECT  207.5 6610.0 837.5 6675.0 ;
      RECT  207.5 5905.0 837.5 5970.0 ;
      RECT  4047.5 5700.0 4112.5 5765.0 ;
      RECT  4047.5 5732.5 4112.5 5937.5 ;
      RECT  592.5 5700.0 4080.0 5765.0 ;
      RECT  7007.5 5700.0 7072.5 5765.0 ;
      RECT  7007.5 5732.5 7072.5 5937.5 ;
      RECT  592.5 5700.0 7040.0 5765.0 ;
      RECT  2057.5 5700.0 2122.5 5765.0 ;
      RECT  2057.5 5732.5 2122.5 5937.5 ;
      RECT  592.5 5700.0 2090.0 5765.0 ;
      RECT  5017.5 5700.0 5082.5 5765.0 ;
      RECT  5017.5 5732.5 5082.5 5937.5 ;
      RECT  592.5 5700.0 5050.0 5765.0 ;
      RECT  9055.0 4632.5 9942.5 4697.5 ;
      RECT  8645.0 2447.5 9942.5 2512.5 ;
      RECT  8850.0 3995.0 9942.5 4060.0 ;
      RECT  9055.0 42425.0 9942.5 42490.0 ;
      RECT  9260.0 11135.0 9942.5 11200.0 ;
      RECT  9465.0 15160.0 9942.5 15225.0 ;
      RECT  1042.5 8930.0 1107.5 8995.0 ;
      RECT  1042.5 8757.5 1107.5 8962.5 ;
      RECT  1075.0 8930.0 8440.0 8995.0 ;
      RECT  5022.5 41620.0 8505.0 41685.0 ;
      RECT  9942.5 43110.0 12072.5 43175.0 ;
      RECT  9942.5 19732.5 12072.5 19797.5 ;
      RECT  9942.5 11265.0 12072.5 11330.0 ;
      RECT  9942.5 7637.5 12072.5 7702.5 ;
      RECT  9942.5 10597.5 12072.5 10662.5 ;
      RECT  9942.5 5647.5 12072.5 5712.5 ;
      RECT  9942.5 8607.5 12072.5 8672.5 ;
      RECT  9942.5 2577.5 12072.5 2642.5 ;
      RECT  592.5 21240.0 12072.5 21305.0 ;
      RECT  592.5 23930.0 12072.5 23995.0 ;
      RECT  592.5 26620.0 12072.5 26685.0 ;
      RECT  592.5 29310.0 12072.5 29375.0 ;
      RECT  592.5 32000.0 12072.5 32065.0 ;
      RECT  592.5 34690.0 12072.5 34755.0 ;
      RECT  592.5 37380.0 12072.5 37445.0 ;
      RECT  592.5 40070.0 12072.5 40135.0 ;
      RECT  9942.5 3865.0 11827.5 3930.0 ;
      RECT  9942.5 15290.0 11827.5 15355.0 ;
      RECT  9942.5 4792.5 11827.5 4857.5 ;
      RECT  9942.5 12067.5 11827.5 12132.5 ;
      RECT  207.5 19895.0 5247.5 19960.0 ;
      RECT  207.5 22585.0 5247.5 22650.0 ;
      RECT  207.5 25275.0 5247.5 25340.0 ;
      RECT  207.5 27965.0 5247.5 28030.0 ;
      RECT  207.5 30655.0 5247.5 30720.0 ;
      RECT  207.5 33345.0 5247.5 33410.0 ;
      RECT  207.5 36035.0 5247.5 36100.0 ;
      RECT  207.5 38725.0 5247.5 38790.0 ;
      RECT  207.5 41415.0 5247.5 41480.0 ;
      RECT  9942.5 19927.5 10647.5 21272.5 ;
      RECT  9942.5 22617.5 10647.5 21272.5 ;
      RECT  9942.5 22617.5 10647.5 23962.5 ;
      RECT  9942.5 25307.5 10647.5 23962.5 ;
      RECT  9942.5 25307.5 10647.5 26652.5 ;
      RECT  9942.5 27997.5 10647.5 26652.5 ;
      RECT  9942.5 27997.5 10647.5 29342.5 ;
      RECT  9942.5 30687.5 10647.5 29342.5 ;
      RECT  9942.5 30687.5 10647.5 32032.5 ;
      RECT  9942.5 33377.5 10647.5 32032.5 ;
      RECT  9942.5 33377.5 10647.5 34722.5 ;
      RECT  9942.5 36067.5 10647.5 34722.5 ;
      RECT  9942.5 36067.5 10647.5 37412.5 ;
      RECT  9942.5 38757.5 10647.5 37412.5 ;
      RECT  9942.5 38757.5 10647.5 40102.5 ;
      RECT  9942.5 41447.5 10647.5 40102.5 ;
      RECT  10647.5 19927.5 11352.5 21272.5 ;
      RECT  10647.5 22617.5 11352.5 21272.5 ;
      RECT  10647.5 22617.5 11352.5 23962.5 ;
      RECT  10647.5 25307.5 11352.5 23962.5 ;
      RECT  10647.5 25307.5 11352.5 26652.5 ;
      RECT  10647.5 27997.5 11352.5 26652.5 ;
      RECT  10647.5 27997.5 11352.5 29342.5 ;
      RECT  10647.5 30687.5 11352.5 29342.5 ;
      RECT  10647.5 30687.5 11352.5 32032.5 ;
      RECT  10647.5 33377.5 11352.5 32032.5 ;
      RECT  10647.5 33377.5 11352.5 34722.5 ;
      RECT  10647.5 36067.5 11352.5 34722.5 ;
      RECT  10647.5 36067.5 11352.5 37412.5 ;
      RECT  10647.5 38757.5 11352.5 37412.5 ;
      RECT  10647.5 38757.5 11352.5 40102.5 ;
      RECT  10647.5 41447.5 11352.5 40102.5 ;
      RECT  9852.5 20035.0 11442.5 20100.0 ;
      RECT  9852.5 22445.0 11442.5 22510.0 ;
      RECT  9852.5 22725.0 11442.5 22790.0 ;
      RECT  9852.5 25135.0 11442.5 25200.0 ;
      RECT  9852.5 25415.0 11442.5 25480.0 ;
      RECT  9852.5 27825.0 11442.5 27890.0 ;
      RECT  9852.5 28105.0 11442.5 28170.0 ;
      RECT  9852.5 30515.0 11442.5 30580.0 ;
      RECT  9852.5 30795.0 11442.5 30860.0 ;
      RECT  9852.5 33205.0 11442.5 33270.0 ;
      RECT  9852.5 33485.0 11442.5 33550.0 ;
      RECT  9852.5 35895.0 11442.5 35960.0 ;
      RECT  9852.5 36175.0 11442.5 36240.0 ;
      RECT  9852.5 38585.0 11442.5 38650.0 ;
      RECT  9852.5 38865.0 11442.5 38930.0 ;
      RECT  9852.5 41275.0 11442.5 41340.0 ;
      RECT  9852.5 21240.0 11442.5 21305.0 ;
      RECT  9852.5 23930.0 11442.5 23995.0 ;
      RECT  9852.5 26620.0 11442.5 26685.0 ;
      RECT  9852.5 29310.0 11442.5 29375.0 ;
      RECT  9852.5 32000.0 11442.5 32065.0 ;
      RECT  9852.5 34690.0 11442.5 34755.0 ;
      RECT  9852.5 37380.0 11442.5 37445.0 ;
      RECT  9852.5 40070.0 11442.5 40135.0 ;
      RECT  9852.5 19895.0 11442.5 19960.0 ;
      RECT  9852.5 22585.0 11442.5 22650.0 ;
      RECT  9852.5 25275.0 11442.5 25340.0 ;
      RECT  9852.5 27965.0 11442.5 28030.0 ;
      RECT  9852.5 30655.0 11442.5 30720.0 ;
      RECT  9852.5 33345.0 11442.5 33410.0 ;
      RECT  9852.5 36035.0 11442.5 36100.0 ;
      RECT  9852.5 38725.0 11442.5 38790.0 ;
      RECT  9852.5 41415.0 11442.5 41480.0 ;
      RECT  10295.0 42660.0 10360.0 43175.0 ;
      RECT  10105.0 42130.0 10170.0 42265.0 ;
      RECT  10295.0 42130.0 10360.0 42265.0 ;
      RECT  10295.0 42130.0 10360.0 42265.0 ;
      RECT  10105.0 42130.0 10170.0 42265.0 ;
      RECT  10105.0 42660.0 10170.0 42795.0 ;
      RECT  10295.0 42660.0 10360.0 42795.0 ;
      RECT  10295.0 42660.0 10360.0 42795.0 ;
      RECT  10105.0 42660.0 10170.0 42795.0 ;
      RECT  10295.0 42660.0 10360.0 42795.0 ;
      RECT  10485.0 42660.0 10550.0 42795.0 ;
      RECT  10485.0 42660.0 10550.0 42795.0 ;
      RECT  10295.0 42660.0 10360.0 42795.0 ;
      RECT  10275.0 42425.0 10140.0 42490.0 ;
      RECT  10295.0 42972.5 10360.0 43107.5 ;
      RECT  10105.0 42130.0 10170.0 42265.0 ;
      RECT  10295.0 42130.0 10360.0 42265.0 ;
      RECT  10105.0 42660.0 10170.0 42795.0 ;
      RECT  10485.0 42660.0 10550.0 42795.0 ;
      RECT  9942.5 42425.0 10647.5 42490.0 ;
      RECT  9942.5 43110.0 10647.5 43175.0 ;
      RECT  11000.0 42660.0 11065.0 43175.0 ;
      RECT  10810.0 42130.0 10875.0 42265.0 ;
      RECT  11000.0 42130.0 11065.0 42265.0 ;
      RECT  11000.0 42130.0 11065.0 42265.0 ;
      RECT  10810.0 42130.0 10875.0 42265.0 ;
      RECT  10810.0 42660.0 10875.0 42795.0 ;
      RECT  11000.0 42660.0 11065.0 42795.0 ;
      RECT  11000.0 42660.0 11065.0 42795.0 ;
      RECT  10810.0 42660.0 10875.0 42795.0 ;
      RECT  11000.0 42660.0 11065.0 42795.0 ;
      RECT  11190.0 42660.0 11255.0 42795.0 ;
      RECT  11190.0 42660.0 11255.0 42795.0 ;
      RECT  11000.0 42660.0 11065.0 42795.0 ;
      RECT  10980.0 42425.0 10845.0 42490.0 ;
      RECT  11000.0 42972.5 11065.0 43107.5 ;
      RECT  10810.0 42130.0 10875.0 42265.0 ;
      RECT  11000.0 42130.0 11065.0 42265.0 ;
      RECT  10810.0 42660.0 10875.0 42795.0 ;
      RECT  11190.0 42660.0 11255.0 42795.0 ;
      RECT  10647.5 42425.0 11352.5 42490.0 ;
      RECT  10647.5 43110.0 11352.5 43175.0 ;
      RECT  9942.5 42425.0 11352.5 42490.0 ;
      RECT  9942.5 43110.0 11352.5 43175.0 ;
      RECT  9942.5 15042.5 10647.5 19927.5 ;
      RECT  10647.5 15042.5 11352.5 19927.5 ;
      RECT  9942.5 15160.0 11352.5 15225.0 ;
      RECT  9942.5 19732.5 11352.5 19797.5 ;
      RECT  9942.5 15290.0 11352.5 15355.0 ;
      RECT  9942.5 10867.5 10647.5 15042.5 ;
      RECT  10647.5 10867.5 11352.5 15042.5 ;
      RECT  9942.5 11135.0 11352.5 11200.0 ;
      RECT  9942.5 11265.0 11352.5 11330.0 ;
      RECT  9942.5 12067.5 11352.5 12132.5 ;
      RECT  9942.5 4427.5 10647.5 10867.5 ;
      RECT  11352.5 4427.5 10647.5 10867.5 ;
      RECT  9942.5 4632.5 11352.5 4697.5 ;
      RECT  9942.5 7637.5 11352.5 7702.5 ;
      RECT  9942.5 10597.5 11352.5 10662.5 ;
      RECT  9942.5 5647.5 11352.5 5712.5 ;
      RECT  9942.5 8607.5 11352.5 8672.5 ;
      RECT  9942.5 4792.5 11352.5 4857.5 ;
      RECT  9942.5 4427.5 10647.5 1452.5 ;
      RECT  10647.5 4427.5 11352.5 1452.5 ;
      RECT  9942.5 4060.0 11352.5 3995.0 ;
      RECT  9942.5 2512.5 11352.5 2447.5 ;
      RECT  9942.5 2642.5 11352.5 2577.5 ;
      RECT  9942.5 3930.0 11352.5 3865.0 ;
      RECT  4077.5 20535.0 4142.5 20600.0 ;
      RECT  4077.5 20522.5 4142.5 20587.5 ;
      RECT  3860.0 20535.0 4110.0 20600.0 ;
      RECT  4077.5 20555.0 4142.5 20567.5 ;
      RECT  4110.0 20522.5 4357.5 20587.5 ;
      RECT  4077.5 21945.0 4142.5 22010.0 ;
      RECT  4077.5 21957.5 4142.5 22022.5 ;
      RECT  3860.0 21945.0 4110.0 22010.0 ;
      RECT  4077.5 21977.5 4142.5 21990.0 ;
      RECT  4110.0 21957.5 4357.5 22022.5 ;
      RECT  4077.5 23225.0 4142.5 23290.0 ;
      RECT  4077.5 23212.5 4142.5 23277.5 ;
      RECT  3860.0 23225.0 4110.0 23290.0 ;
      RECT  4077.5 23245.0 4142.5 23257.5 ;
      RECT  4110.0 23212.5 4357.5 23277.5 ;
      RECT  4077.5 24635.0 4142.5 24700.0 ;
      RECT  4077.5 24647.5 4142.5 24712.5 ;
      RECT  3860.0 24635.0 4110.0 24700.0 ;
      RECT  4077.5 24667.5 4142.5 24680.0 ;
      RECT  4110.0 24647.5 4357.5 24712.5 ;
      RECT  4077.5 25915.0 4142.5 25980.0 ;
      RECT  4077.5 25902.5 4142.5 25967.5 ;
      RECT  3860.0 25915.0 4110.0 25980.0 ;
      RECT  4077.5 25935.0 4142.5 25947.5 ;
      RECT  4110.0 25902.5 4357.5 25967.5 ;
      RECT  4077.5 27325.0 4142.5 27390.0 ;
      RECT  4077.5 27337.5 4142.5 27402.5 ;
      RECT  3860.0 27325.0 4110.0 27390.0 ;
      RECT  4077.5 27357.5 4142.5 27370.0 ;
      RECT  4110.0 27337.5 4357.5 27402.5 ;
      RECT  4077.5 28605.0 4142.5 28670.0 ;
      RECT  4077.5 28592.5 4142.5 28657.5 ;
      RECT  3860.0 28605.0 4110.0 28670.0 ;
      RECT  4077.5 28625.0 4142.5 28637.5 ;
      RECT  4110.0 28592.5 4357.5 28657.5 ;
      RECT  4077.5 30015.0 4142.5 30080.0 ;
      RECT  4077.5 30027.5 4142.5 30092.5 ;
      RECT  3860.0 30015.0 4110.0 30080.0 ;
      RECT  4077.5 30047.5 4142.5 30060.0 ;
      RECT  4110.0 30027.5 4357.5 30092.5 ;
      RECT  4077.5 31295.0 4142.5 31360.0 ;
      RECT  4077.5 31282.5 4142.5 31347.5 ;
      RECT  3860.0 31295.0 4110.0 31360.0 ;
      RECT  4077.5 31315.0 4142.5 31327.5 ;
      RECT  4110.0 31282.5 4357.5 31347.5 ;
      RECT  4077.5 32705.0 4142.5 32770.0 ;
      RECT  4077.5 32717.5 4142.5 32782.5 ;
      RECT  3860.0 32705.0 4110.0 32770.0 ;
      RECT  4077.5 32737.5 4142.5 32750.0 ;
      RECT  4110.0 32717.5 4357.5 32782.5 ;
      RECT  4077.5 33985.0 4142.5 34050.0 ;
      RECT  4077.5 33972.5 4142.5 34037.5 ;
      RECT  3860.0 33985.0 4110.0 34050.0 ;
      RECT  4077.5 34005.0 4142.5 34017.5 ;
      RECT  4110.0 33972.5 4357.5 34037.5 ;
      RECT  4077.5 35395.0 4142.5 35460.0 ;
      RECT  4077.5 35407.5 4142.5 35472.5 ;
      RECT  3860.0 35395.0 4110.0 35460.0 ;
      RECT  4077.5 35427.5 4142.5 35440.0 ;
      RECT  4110.0 35407.5 4357.5 35472.5 ;
      RECT  4077.5 36675.0 4142.5 36740.0 ;
      RECT  4077.5 36662.5 4142.5 36727.5 ;
      RECT  3860.0 36675.0 4110.0 36740.0 ;
      RECT  4077.5 36695.0 4142.5 36707.5 ;
      RECT  4110.0 36662.5 4357.5 36727.5 ;
      RECT  4077.5 38085.0 4142.5 38150.0 ;
      RECT  4077.5 38097.5 4142.5 38162.5 ;
      RECT  3860.0 38085.0 4110.0 38150.0 ;
      RECT  4077.5 38117.5 4142.5 38130.0 ;
      RECT  4110.0 38097.5 4357.5 38162.5 ;
      RECT  4077.5 39365.0 4142.5 39430.0 ;
      RECT  4077.5 39352.5 4142.5 39417.5 ;
      RECT  3860.0 39365.0 4110.0 39430.0 ;
      RECT  4077.5 39385.0 4142.5 39397.5 ;
      RECT  4110.0 39352.5 4357.5 39417.5 ;
      RECT  4077.5 40775.0 4142.5 40840.0 ;
      RECT  4077.5 40787.5 4142.5 40852.5 ;
      RECT  3860.0 40775.0 4110.0 40840.0 ;
      RECT  4077.5 40807.5 4142.5 40820.0 ;
      RECT  4110.0 40787.5 4357.5 40852.5 ;
      RECT  1947.5 9762.5 3312.5 9827.5 ;
      RECT  2122.5 11197.5 3312.5 11262.5 ;
      RECT  2297.5 12452.5 3312.5 12517.5 ;
      RECT  2472.5 13887.5 3312.5 13952.5 ;
      RECT  2647.5 15142.5 3312.5 15207.5 ;
      RECT  2822.5 16577.5 3312.5 16642.5 ;
      RECT  2997.5 17832.5 3312.5 17897.5 ;
      RECT  3172.5 19267.5 3312.5 19332.5 ;
      RECT  1947.5 20535.0 3372.5 20600.0 ;
      RECT  2647.5 20320.0 3630.0 20385.0 ;
      RECT  1947.5 21945.0 3372.5 22010.0 ;
      RECT  2822.5 22160.0 3630.0 22225.0 ;
      RECT  1947.5 23225.0 3372.5 23290.0 ;
      RECT  2997.5 23010.0 3630.0 23075.0 ;
      RECT  1947.5 24635.0 3372.5 24700.0 ;
      RECT  3172.5 24850.0 3630.0 24915.0 ;
      RECT  2122.5 25915.0 3372.5 25980.0 ;
      RECT  2647.5 25700.0 3630.0 25765.0 ;
      RECT  2122.5 27325.0 3372.5 27390.0 ;
      RECT  2822.5 27540.0 3630.0 27605.0 ;
      RECT  2122.5 28605.0 3372.5 28670.0 ;
      RECT  2997.5 28390.0 3630.0 28455.0 ;
      RECT  2122.5 30015.0 3372.5 30080.0 ;
      RECT  3172.5 30230.0 3630.0 30295.0 ;
      RECT  2297.5 31295.0 3372.5 31360.0 ;
      RECT  2647.5 31080.0 3630.0 31145.0 ;
      RECT  2297.5 32705.0 3372.5 32770.0 ;
      RECT  2822.5 32920.0 3630.0 32985.0 ;
      RECT  2297.5 33985.0 3372.5 34050.0 ;
      RECT  2997.5 33770.0 3630.0 33835.0 ;
      RECT  2297.5 35395.0 3372.5 35460.0 ;
      RECT  3172.5 35610.0 3630.0 35675.0 ;
      RECT  2472.5 36675.0 3372.5 36740.0 ;
      RECT  2647.5 36460.0 3630.0 36525.0 ;
      RECT  2472.5 38085.0 3372.5 38150.0 ;
      RECT  2822.5 38300.0 3630.0 38365.0 ;
      RECT  2472.5 39365.0 3372.5 39430.0 ;
      RECT  2997.5 39150.0 3630.0 39215.0 ;
      RECT  2472.5 40775.0 3372.5 40840.0 ;
      RECT  3172.5 40990.0 3630.0 41055.0 ;
      RECT  6135.0 9762.5 6070.0 9827.5 ;
      RECT  6135.0 10285.0 6070.0 10350.0 ;
      RECT  6372.5 9762.5 6102.5 9827.5 ;
      RECT  6135.0 9795.0 6070.0 10317.5 ;
      RECT  6102.5 10285.0 5857.5 10350.0 ;
      RECT  7242.5 9762.5 6602.5 9827.5 ;
      RECT  6135.0 11197.5 6070.0 11262.5 ;
      RECT  6135.0 11630.0 6070.0 11695.0 ;
      RECT  6372.5 11197.5 6102.5 11262.5 ;
      RECT  6135.0 11230.0 6070.0 11662.5 ;
      RECT  6102.5 11630.0 5582.5 11695.0 ;
      RECT  6967.5 11197.5 6602.5 11262.5 ;
      RECT  7242.5 11960.0 5307.5 12025.0 ;
      RECT  6967.5 13305.0 5032.5 13370.0 ;
      RECT  5857.5 9775.0 4732.5 9840.0 ;
      RECT  5582.5 9560.0 4475.0 9625.0 ;
      RECT  5307.5 11185.0 4732.5 11250.0 ;
      RECT  5582.5 11400.0 4475.0 11465.0 ;
      RECT  5857.5 12465.0 4732.5 12530.0 ;
      RECT  5032.5 12250.0 4475.0 12315.0 ;
      RECT  5307.5 13875.0 4732.5 13940.0 ;
      RECT  5032.5 14090.0 4475.0 14155.0 ;
      RECT  4027.5 9775.0 3962.5 9840.0 ;
      RECT  4027.5 9762.5 3962.5 9827.5 ;
      RECT  4245.0 9775.0 3995.0 9840.0 ;
      RECT  4027.5 9795.0 3962.5 9807.5 ;
      RECT  3995.0 9762.5 3747.5 9827.5 ;
      RECT  4027.5 11185.0 3962.5 11250.0 ;
      RECT  4027.5 11197.5 3962.5 11262.5 ;
      RECT  4245.0 11185.0 3995.0 11250.0 ;
      RECT  4027.5 11217.5 3962.5 11230.0 ;
      RECT  3995.0 11197.5 3747.5 11262.5 ;
      RECT  4027.5 12465.0 3962.5 12530.0 ;
      RECT  4027.5 12452.5 3962.5 12517.5 ;
      RECT  4245.0 12465.0 3995.0 12530.0 ;
      RECT  4027.5 12485.0 3962.5 12497.5 ;
      RECT  3995.0 12452.5 3747.5 12517.5 ;
      RECT  4027.5 13875.0 3962.5 13940.0 ;
      RECT  4027.5 13887.5 3962.5 13952.5 ;
      RECT  4245.0 13875.0 3995.0 13940.0 ;
      RECT  4027.5 13907.5 3962.5 13920.0 ;
      RECT  3995.0 13887.5 3747.5 13952.5 ;
      RECT  6300.0 10327.5 6235.0 10512.5 ;
      RECT  6300.0 9167.5 6235.0 9352.5 ;
      RECT  6660.0 9285.0 6595.0 9135.0 ;
      RECT  6660.0 10170.0 6595.0 10545.0 ;
      RECT  6470.0 9285.0 6405.0 10170.0 ;
      RECT  6660.0 10170.0 6595.0 10305.0 ;
      RECT  6470.0 10170.0 6405.0 10305.0 ;
      RECT  6470.0 10170.0 6405.0 10305.0 ;
      RECT  6660.0 10170.0 6595.0 10305.0 ;
      RECT  6660.0 9285.0 6595.0 9420.0 ;
      RECT  6470.0 9285.0 6405.0 9420.0 ;
      RECT  6470.0 9285.0 6405.0 9420.0 ;
      RECT  6660.0 9285.0 6595.0 9420.0 ;
      RECT  6300.0 10260.0 6235.0 10395.0 ;
      RECT  6300.0 9285.0 6235.0 9420.0 ;
      RECT  6602.5 9727.5 6537.5 9862.5 ;
      RECT  6602.5 9727.5 6537.5 9862.5 ;
      RECT  6437.5 9762.5 6372.5 9827.5 ;
      RECT  6727.5 10480.0 6167.5 10545.0 ;
      RECT  6727.5 9135.0 6167.5 9200.0 ;
      RECT  6300.0 10697.5 6235.0 10512.5 ;
      RECT  6300.0 11857.5 6235.0 11672.5 ;
      RECT  6660.0 11740.0 6595.0 11890.0 ;
      RECT  6660.0 10855.0 6595.0 10480.0 ;
      RECT  6470.0 11740.0 6405.0 10855.0 ;
      RECT  6660.0 10855.0 6595.0 10720.0 ;
      RECT  6470.0 10855.0 6405.0 10720.0 ;
      RECT  6470.0 10855.0 6405.0 10720.0 ;
      RECT  6660.0 10855.0 6595.0 10720.0 ;
      RECT  6660.0 11740.0 6595.0 11605.0 ;
      RECT  6470.0 11740.0 6405.0 11605.0 ;
      RECT  6470.0 11740.0 6405.0 11605.0 ;
      RECT  6660.0 11740.0 6595.0 11605.0 ;
      RECT  6300.0 10765.0 6235.0 10630.0 ;
      RECT  6300.0 11740.0 6235.0 11605.0 ;
      RECT  6602.5 11297.5 6537.5 11162.5 ;
      RECT  6602.5 11297.5 6537.5 11162.5 ;
      RECT  6437.5 11262.5 6372.5 11197.5 ;
      RECT  6727.5 10545.0 6167.5 10480.0 ;
      RECT  6727.5 11890.0 6167.5 11825.0 ;
      RECT  3445.0 10327.5 3380.0 10512.5 ;
      RECT  3445.0 9167.5 3380.0 9352.5 ;
      RECT  3805.0 9285.0 3740.0 9135.0 ;
      RECT  3805.0 10170.0 3740.0 10545.0 ;
      RECT  3615.0 9285.0 3550.0 10170.0 ;
      RECT  3805.0 10170.0 3740.0 10305.0 ;
      RECT  3615.0 10170.0 3550.0 10305.0 ;
      RECT  3615.0 10170.0 3550.0 10305.0 ;
      RECT  3805.0 10170.0 3740.0 10305.0 ;
      RECT  3805.0 9285.0 3740.0 9420.0 ;
      RECT  3615.0 9285.0 3550.0 9420.0 ;
      RECT  3615.0 9285.0 3550.0 9420.0 ;
      RECT  3805.0 9285.0 3740.0 9420.0 ;
      RECT  3445.0 10260.0 3380.0 10395.0 ;
      RECT  3445.0 9285.0 3380.0 9420.0 ;
      RECT  3747.5 9727.5 3682.5 9862.5 ;
      RECT  3747.5 9727.5 3682.5 9862.5 ;
      RECT  3582.5 9762.5 3517.5 9827.5 ;
      RECT  3872.5 10480.0 3312.5 10545.0 ;
      RECT  3872.5 9135.0 3312.5 9200.0 ;
      RECT  3445.0 10697.5 3380.0 10512.5 ;
      RECT  3445.0 11857.5 3380.0 11672.5 ;
      RECT  3805.0 11740.0 3740.0 11890.0 ;
      RECT  3805.0 10855.0 3740.0 10480.0 ;
      RECT  3615.0 11740.0 3550.0 10855.0 ;
      RECT  3805.0 10855.0 3740.0 10720.0 ;
      RECT  3615.0 10855.0 3550.0 10720.0 ;
      RECT  3615.0 10855.0 3550.0 10720.0 ;
      RECT  3805.0 10855.0 3740.0 10720.0 ;
      RECT  3805.0 11740.0 3740.0 11605.0 ;
      RECT  3615.0 11740.0 3550.0 11605.0 ;
      RECT  3615.0 11740.0 3550.0 11605.0 ;
      RECT  3805.0 11740.0 3740.0 11605.0 ;
      RECT  3445.0 10765.0 3380.0 10630.0 ;
      RECT  3445.0 11740.0 3380.0 11605.0 ;
      RECT  3747.5 11297.5 3682.5 11162.5 ;
      RECT  3747.5 11297.5 3682.5 11162.5 ;
      RECT  3582.5 11262.5 3517.5 11197.5 ;
      RECT  3872.5 10545.0 3312.5 10480.0 ;
      RECT  3872.5 11890.0 3312.5 11825.0 ;
      RECT  3445.0 13017.5 3380.0 13202.5 ;
      RECT  3445.0 11857.5 3380.0 12042.5 ;
      RECT  3805.0 11975.0 3740.0 11825.0 ;
      RECT  3805.0 12860.0 3740.0 13235.0 ;
      RECT  3615.0 11975.0 3550.0 12860.0 ;
      RECT  3805.0 12860.0 3740.0 12995.0 ;
      RECT  3615.0 12860.0 3550.0 12995.0 ;
      RECT  3615.0 12860.0 3550.0 12995.0 ;
      RECT  3805.0 12860.0 3740.0 12995.0 ;
      RECT  3805.0 11975.0 3740.0 12110.0 ;
      RECT  3615.0 11975.0 3550.0 12110.0 ;
      RECT  3615.0 11975.0 3550.0 12110.0 ;
      RECT  3805.0 11975.0 3740.0 12110.0 ;
      RECT  3445.0 12950.0 3380.0 13085.0 ;
      RECT  3445.0 11975.0 3380.0 12110.0 ;
      RECT  3747.5 12417.5 3682.5 12552.5 ;
      RECT  3747.5 12417.5 3682.5 12552.5 ;
      RECT  3582.5 12452.5 3517.5 12517.5 ;
      RECT  3872.5 13170.0 3312.5 13235.0 ;
      RECT  3872.5 11825.0 3312.5 11890.0 ;
      RECT  3445.0 13387.5 3380.0 13202.5 ;
      RECT  3445.0 14547.5 3380.0 14362.5 ;
      RECT  3805.0 14430.0 3740.0 14580.0 ;
      RECT  3805.0 13545.0 3740.0 13170.0 ;
      RECT  3615.0 14430.0 3550.0 13545.0 ;
      RECT  3805.0 13545.0 3740.0 13410.0 ;
      RECT  3615.0 13545.0 3550.0 13410.0 ;
      RECT  3615.0 13545.0 3550.0 13410.0 ;
      RECT  3805.0 13545.0 3740.0 13410.0 ;
      RECT  3805.0 14430.0 3740.0 14295.0 ;
      RECT  3615.0 14430.0 3550.0 14295.0 ;
      RECT  3615.0 14430.0 3550.0 14295.0 ;
      RECT  3805.0 14430.0 3740.0 14295.0 ;
      RECT  3445.0 13455.0 3380.0 13320.0 ;
      RECT  3445.0 14430.0 3380.0 14295.0 ;
      RECT  3747.5 13987.5 3682.5 13852.5 ;
      RECT  3747.5 13987.5 3682.5 13852.5 ;
      RECT  3582.5 13952.5 3517.5 13887.5 ;
      RECT  3872.5 13235.0 3312.5 13170.0 ;
      RECT  3872.5 14580.0 3312.5 14515.0 ;
      RECT  4725.0 9330.0 4660.0 9135.0 ;
      RECT  4725.0 10170.0 4660.0 10545.0 ;
      RECT  4345.0 10170.0 4280.0 10545.0 ;
      RECT  4175.0 10327.5 4110.0 10512.5 ;
      RECT  4175.0 9167.5 4110.0 9352.5 ;
      RECT  4725.0 10170.0 4660.0 10305.0 ;
      RECT  4535.0 10170.0 4470.0 10305.0 ;
      RECT  4535.0 10170.0 4470.0 10305.0 ;
      RECT  4725.0 10170.0 4660.0 10305.0 ;
      RECT  4535.0 10170.0 4470.0 10305.0 ;
      RECT  4345.0 10170.0 4280.0 10305.0 ;
      RECT  4345.0 10170.0 4280.0 10305.0 ;
      RECT  4535.0 10170.0 4470.0 10305.0 ;
      RECT  4725.0 9330.0 4660.0 9465.0 ;
      RECT  4535.0 9330.0 4470.0 9465.0 ;
      RECT  4535.0 9330.0 4470.0 9465.0 ;
      RECT  4725.0 9330.0 4660.0 9465.0 ;
      RECT  4535.0 9330.0 4470.0 9465.0 ;
      RECT  4345.0 9330.0 4280.0 9465.0 ;
      RECT  4345.0 9330.0 4280.0 9465.0 ;
      RECT  4535.0 9330.0 4470.0 9465.0 ;
      RECT  4175.0 10260.0 4110.0 10395.0 ;
      RECT  4175.0 9285.0 4110.0 9420.0 ;
      RECT  4340.0 9560.0 4475.0 9625.0 ;
      RECT  4597.5 9775.0 4732.5 9840.0 ;
      RECT  4535.0 10170.0 4470.0 10305.0 ;
      RECT  4345.0 9330.0 4280.0 9465.0 ;
      RECT  4245.0 9775.0 4380.0 9840.0 ;
      RECT  4732.5 9775.0 4597.5 9840.0 ;
      RECT  4475.0 9560.0 4340.0 9625.0 ;
      RECT  4380.0 9775.0 4245.0 9840.0 ;
      RECT  4792.5 10480.0 3872.5 10545.0 ;
      RECT  4792.5 9135.0 3872.5 9200.0 ;
      RECT  4725.0 11695.0 4660.0 11890.0 ;
      RECT  4725.0 10855.0 4660.0 10480.0 ;
      RECT  4345.0 10855.0 4280.0 10480.0 ;
      RECT  4175.0 10697.5 4110.0 10512.5 ;
      RECT  4175.0 11857.5 4110.0 11672.5 ;
      RECT  4725.0 10855.0 4660.0 10720.0 ;
      RECT  4535.0 10855.0 4470.0 10720.0 ;
      RECT  4535.0 10855.0 4470.0 10720.0 ;
      RECT  4725.0 10855.0 4660.0 10720.0 ;
      RECT  4535.0 10855.0 4470.0 10720.0 ;
      RECT  4345.0 10855.0 4280.0 10720.0 ;
      RECT  4345.0 10855.0 4280.0 10720.0 ;
      RECT  4535.0 10855.0 4470.0 10720.0 ;
      RECT  4725.0 11695.0 4660.0 11560.0 ;
      RECT  4535.0 11695.0 4470.0 11560.0 ;
      RECT  4535.0 11695.0 4470.0 11560.0 ;
      RECT  4725.0 11695.0 4660.0 11560.0 ;
      RECT  4535.0 11695.0 4470.0 11560.0 ;
      RECT  4345.0 11695.0 4280.0 11560.0 ;
      RECT  4345.0 11695.0 4280.0 11560.0 ;
      RECT  4535.0 11695.0 4470.0 11560.0 ;
      RECT  4175.0 10765.0 4110.0 10630.0 ;
      RECT  4175.0 11740.0 4110.0 11605.0 ;
      RECT  4340.0 11465.0 4475.0 11400.0 ;
      RECT  4597.5 11250.0 4732.5 11185.0 ;
      RECT  4535.0 10855.0 4470.0 10720.0 ;
      RECT  4345.0 11695.0 4280.0 11560.0 ;
      RECT  4245.0 11250.0 4380.0 11185.0 ;
      RECT  4732.5 11250.0 4597.5 11185.0 ;
      RECT  4475.0 11465.0 4340.0 11400.0 ;
      RECT  4380.0 11250.0 4245.0 11185.0 ;
      RECT  4792.5 10545.0 3872.5 10480.0 ;
      RECT  4792.5 11890.0 3872.5 11825.0 ;
      RECT  4725.0 12020.0 4660.0 11825.0 ;
      RECT  4725.0 12860.0 4660.0 13235.0 ;
      RECT  4345.0 12860.0 4280.0 13235.0 ;
      RECT  4175.0 13017.5 4110.0 13202.5 ;
      RECT  4175.0 11857.5 4110.0 12042.5 ;
      RECT  4725.0 12860.0 4660.0 12995.0 ;
      RECT  4535.0 12860.0 4470.0 12995.0 ;
      RECT  4535.0 12860.0 4470.0 12995.0 ;
      RECT  4725.0 12860.0 4660.0 12995.0 ;
      RECT  4535.0 12860.0 4470.0 12995.0 ;
      RECT  4345.0 12860.0 4280.0 12995.0 ;
      RECT  4345.0 12860.0 4280.0 12995.0 ;
      RECT  4535.0 12860.0 4470.0 12995.0 ;
      RECT  4725.0 12020.0 4660.0 12155.0 ;
      RECT  4535.0 12020.0 4470.0 12155.0 ;
      RECT  4535.0 12020.0 4470.0 12155.0 ;
      RECT  4725.0 12020.0 4660.0 12155.0 ;
      RECT  4535.0 12020.0 4470.0 12155.0 ;
      RECT  4345.0 12020.0 4280.0 12155.0 ;
      RECT  4345.0 12020.0 4280.0 12155.0 ;
      RECT  4535.0 12020.0 4470.0 12155.0 ;
      RECT  4175.0 12950.0 4110.0 13085.0 ;
      RECT  4175.0 11975.0 4110.0 12110.0 ;
      RECT  4340.0 12250.0 4475.0 12315.0 ;
      RECT  4597.5 12465.0 4732.5 12530.0 ;
      RECT  4535.0 12860.0 4470.0 12995.0 ;
      RECT  4345.0 12020.0 4280.0 12155.0 ;
      RECT  4245.0 12465.0 4380.0 12530.0 ;
      RECT  4732.5 12465.0 4597.5 12530.0 ;
      RECT  4475.0 12250.0 4340.0 12315.0 ;
      RECT  4380.0 12465.0 4245.0 12530.0 ;
      RECT  4792.5 13170.0 3872.5 13235.0 ;
      RECT  4792.5 11825.0 3872.5 11890.0 ;
      RECT  4725.0 14385.0 4660.0 14580.0 ;
      RECT  4725.0 13545.0 4660.0 13170.0 ;
      RECT  4345.0 13545.0 4280.0 13170.0 ;
      RECT  4175.0 13387.5 4110.0 13202.5 ;
      RECT  4175.0 14547.5 4110.0 14362.5 ;
      RECT  4725.0 13545.0 4660.0 13410.0 ;
      RECT  4535.0 13545.0 4470.0 13410.0 ;
      RECT  4535.0 13545.0 4470.0 13410.0 ;
      RECT  4725.0 13545.0 4660.0 13410.0 ;
      RECT  4535.0 13545.0 4470.0 13410.0 ;
      RECT  4345.0 13545.0 4280.0 13410.0 ;
      RECT  4345.0 13545.0 4280.0 13410.0 ;
      RECT  4535.0 13545.0 4470.0 13410.0 ;
      RECT  4725.0 14385.0 4660.0 14250.0 ;
      RECT  4535.0 14385.0 4470.0 14250.0 ;
      RECT  4535.0 14385.0 4470.0 14250.0 ;
      RECT  4725.0 14385.0 4660.0 14250.0 ;
      RECT  4535.0 14385.0 4470.0 14250.0 ;
      RECT  4345.0 14385.0 4280.0 14250.0 ;
      RECT  4345.0 14385.0 4280.0 14250.0 ;
      RECT  4535.0 14385.0 4470.0 14250.0 ;
      RECT  4175.0 13455.0 4110.0 13320.0 ;
      RECT  4175.0 14430.0 4110.0 14295.0 ;
      RECT  4340.0 14155.0 4475.0 14090.0 ;
      RECT  4597.5 13940.0 4732.5 13875.0 ;
      RECT  4535.0 13545.0 4470.0 13410.0 ;
      RECT  4345.0 14385.0 4280.0 14250.0 ;
      RECT  4245.0 13940.0 4380.0 13875.0 ;
      RECT  4732.5 13940.0 4597.5 13875.0 ;
      RECT  4475.0 14155.0 4340.0 14090.0 ;
      RECT  4380.0 13940.0 4245.0 13875.0 ;
      RECT  4792.5 13235.0 3872.5 13170.0 ;
      RECT  4792.5 14580.0 3872.5 14515.0 ;
      RECT  5790.0 10285.0 5925.0 10350.0 ;
      RECT  7175.0 9762.5 7310.0 9827.5 ;
      RECT  5515.0 11630.0 5650.0 11695.0 ;
      RECT  6900.0 11197.5 7035.0 11262.5 ;
      RECT  7175.0 11960.0 7310.0 12025.0 ;
      RECT  5240.0 11960.0 5375.0 12025.0 ;
      RECT  6900.0 13305.0 7035.0 13370.0 ;
      RECT  4965.0 13305.0 5100.0 13370.0 ;
      RECT  5790.0 9775.0 5925.0 9840.0 ;
      RECT  5515.0 9560.0 5650.0 9625.0 ;
      RECT  5240.0 11185.0 5375.0 11250.0 ;
      RECT  5515.0 11400.0 5650.0 11465.0 ;
      RECT  5790.0 12465.0 5925.0 12530.0 ;
      RECT  4965.0 12250.0 5100.0 12315.0 ;
      RECT  5240.0 13875.0 5375.0 13940.0 ;
      RECT  4965.0 14090.0 5100.0 14155.0 ;
      RECT  3517.5 9762.5 3312.5 9827.5 ;
      RECT  3517.5 11197.5 3312.5 11262.5 ;
      RECT  3517.5 12452.5 3312.5 12517.5 ;
      RECT  3517.5 13887.5 3312.5 13952.5 ;
      RECT  7277.5 10480.0 3312.5 10545.0 ;
      RECT  7277.5 13170.0 3312.5 13235.0 ;
      RECT  7277.5 9135.0 3312.5 9200.0 ;
      RECT  7277.5 11825.0 3312.5 11890.0 ;
      RECT  7277.5 14515.0 3312.5 14580.0 ;
      RECT  6135.0 15142.5 6070.0 15207.5 ;
      RECT  6135.0 15665.0 6070.0 15730.0 ;
      RECT  6372.5 15142.5 6102.5 15207.5 ;
      RECT  6135.0 15175.0 6070.0 15697.5 ;
      RECT  6102.5 15665.0 5857.5 15730.0 ;
      RECT  7242.5 15142.5 6602.5 15207.5 ;
      RECT  6135.0 16577.5 6070.0 16642.5 ;
      RECT  6135.0 17010.0 6070.0 17075.0 ;
      RECT  6372.5 16577.5 6102.5 16642.5 ;
      RECT  6135.0 16610.0 6070.0 17042.5 ;
      RECT  6102.5 17010.0 5582.5 17075.0 ;
      RECT  6967.5 16577.5 6602.5 16642.5 ;
      RECT  7242.5 17340.0 5307.5 17405.0 ;
      RECT  6967.5 18685.0 5032.5 18750.0 ;
      RECT  5857.5 15155.0 4732.5 15220.0 ;
      RECT  5582.5 14940.0 4475.0 15005.0 ;
      RECT  5307.5 16565.0 4732.5 16630.0 ;
      RECT  5582.5 16780.0 4475.0 16845.0 ;
      RECT  5857.5 17845.0 4732.5 17910.0 ;
      RECT  5032.5 17630.0 4475.0 17695.0 ;
      RECT  5307.5 19255.0 4732.5 19320.0 ;
      RECT  5032.5 19470.0 4475.0 19535.0 ;
      RECT  4027.5 15155.0 3962.5 15220.0 ;
      RECT  4027.5 15142.5 3962.5 15207.5 ;
      RECT  4245.0 15155.0 3995.0 15220.0 ;
      RECT  4027.5 15175.0 3962.5 15187.5 ;
      RECT  3995.0 15142.5 3747.5 15207.5 ;
      RECT  4027.5 16565.0 3962.5 16630.0 ;
      RECT  4027.5 16577.5 3962.5 16642.5 ;
      RECT  4245.0 16565.0 3995.0 16630.0 ;
      RECT  4027.5 16597.5 3962.5 16610.0 ;
      RECT  3995.0 16577.5 3747.5 16642.5 ;
      RECT  4027.5 17845.0 3962.5 17910.0 ;
      RECT  4027.5 17832.5 3962.5 17897.5 ;
      RECT  4245.0 17845.0 3995.0 17910.0 ;
      RECT  4027.5 17865.0 3962.5 17877.5 ;
      RECT  3995.0 17832.5 3747.5 17897.5 ;
      RECT  4027.5 19255.0 3962.5 19320.0 ;
      RECT  4027.5 19267.5 3962.5 19332.5 ;
      RECT  4245.0 19255.0 3995.0 19320.0 ;
      RECT  4027.5 19287.5 3962.5 19300.0 ;
      RECT  3995.0 19267.5 3747.5 19332.5 ;
      RECT  6300.0 15707.5 6235.0 15892.5 ;
      RECT  6300.0 14547.5 6235.0 14732.5 ;
      RECT  6660.0 14665.0 6595.0 14515.0 ;
      RECT  6660.0 15550.0 6595.0 15925.0 ;
      RECT  6470.0 14665.0 6405.0 15550.0 ;
      RECT  6660.0 15550.0 6595.0 15685.0 ;
      RECT  6470.0 15550.0 6405.0 15685.0 ;
      RECT  6470.0 15550.0 6405.0 15685.0 ;
      RECT  6660.0 15550.0 6595.0 15685.0 ;
      RECT  6660.0 14665.0 6595.0 14800.0 ;
      RECT  6470.0 14665.0 6405.0 14800.0 ;
      RECT  6470.0 14665.0 6405.0 14800.0 ;
      RECT  6660.0 14665.0 6595.0 14800.0 ;
      RECT  6300.0 15640.0 6235.0 15775.0 ;
      RECT  6300.0 14665.0 6235.0 14800.0 ;
      RECT  6602.5 15107.5 6537.5 15242.5 ;
      RECT  6602.5 15107.5 6537.5 15242.5 ;
      RECT  6437.5 15142.5 6372.5 15207.5 ;
      RECT  6727.5 15860.0 6167.5 15925.0 ;
      RECT  6727.5 14515.0 6167.5 14580.0 ;
      RECT  6300.0 16077.5 6235.0 15892.5 ;
      RECT  6300.0 17237.5 6235.0 17052.5 ;
      RECT  6660.0 17120.0 6595.0 17270.0 ;
      RECT  6660.0 16235.0 6595.0 15860.0 ;
      RECT  6470.0 17120.0 6405.0 16235.0 ;
      RECT  6660.0 16235.0 6595.0 16100.0 ;
      RECT  6470.0 16235.0 6405.0 16100.0 ;
      RECT  6470.0 16235.0 6405.0 16100.0 ;
      RECT  6660.0 16235.0 6595.0 16100.0 ;
      RECT  6660.0 17120.0 6595.0 16985.0 ;
      RECT  6470.0 17120.0 6405.0 16985.0 ;
      RECT  6470.0 17120.0 6405.0 16985.0 ;
      RECT  6660.0 17120.0 6595.0 16985.0 ;
      RECT  6300.0 16145.0 6235.0 16010.0 ;
      RECT  6300.0 17120.0 6235.0 16985.0 ;
      RECT  6602.5 16677.5 6537.5 16542.5 ;
      RECT  6602.5 16677.5 6537.5 16542.5 ;
      RECT  6437.5 16642.5 6372.5 16577.5 ;
      RECT  6727.5 15925.0 6167.5 15860.0 ;
      RECT  6727.5 17270.0 6167.5 17205.0 ;
      RECT  3445.0 15707.5 3380.0 15892.5 ;
      RECT  3445.0 14547.5 3380.0 14732.5 ;
      RECT  3805.0 14665.0 3740.0 14515.0 ;
      RECT  3805.0 15550.0 3740.0 15925.0 ;
      RECT  3615.0 14665.0 3550.0 15550.0 ;
      RECT  3805.0 15550.0 3740.0 15685.0 ;
      RECT  3615.0 15550.0 3550.0 15685.0 ;
      RECT  3615.0 15550.0 3550.0 15685.0 ;
      RECT  3805.0 15550.0 3740.0 15685.0 ;
      RECT  3805.0 14665.0 3740.0 14800.0 ;
      RECT  3615.0 14665.0 3550.0 14800.0 ;
      RECT  3615.0 14665.0 3550.0 14800.0 ;
      RECT  3805.0 14665.0 3740.0 14800.0 ;
      RECT  3445.0 15640.0 3380.0 15775.0 ;
      RECT  3445.0 14665.0 3380.0 14800.0 ;
      RECT  3747.5 15107.5 3682.5 15242.5 ;
      RECT  3747.5 15107.5 3682.5 15242.5 ;
      RECT  3582.5 15142.5 3517.5 15207.5 ;
      RECT  3872.5 15860.0 3312.5 15925.0 ;
      RECT  3872.5 14515.0 3312.5 14580.0 ;
      RECT  3445.0 16077.5 3380.0 15892.5 ;
      RECT  3445.0 17237.5 3380.0 17052.5 ;
      RECT  3805.0 17120.0 3740.0 17270.0 ;
      RECT  3805.0 16235.0 3740.0 15860.0 ;
      RECT  3615.0 17120.0 3550.0 16235.0 ;
      RECT  3805.0 16235.0 3740.0 16100.0 ;
      RECT  3615.0 16235.0 3550.0 16100.0 ;
      RECT  3615.0 16235.0 3550.0 16100.0 ;
      RECT  3805.0 16235.0 3740.0 16100.0 ;
      RECT  3805.0 17120.0 3740.0 16985.0 ;
      RECT  3615.0 17120.0 3550.0 16985.0 ;
      RECT  3615.0 17120.0 3550.0 16985.0 ;
      RECT  3805.0 17120.0 3740.0 16985.0 ;
      RECT  3445.0 16145.0 3380.0 16010.0 ;
      RECT  3445.0 17120.0 3380.0 16985.0 ;
      RECT  3747.5 16677.5 3682.5 16542.5 ;
      RECT  3747.5 16677.5 3682.5 16542.5 ;
      RECT  3582.5 16642.5 3517.5 16577.5 ;
      RECT  3872.5 15925.0 3312.5 15860.0 ;
      RECT  3872.5 17270.0 3312.5 17205.0 ;
      RECT  3445.0 18397.5 3380.0 18582.5 ;
      RECT  3445.0 17237.5 3380.0 17422.5 ;
      RECT  3805.0 17355.0 3740.0 17205.0 ;
      RECT  3805.0 18240.0 3740.0 18615.0 ;
      RECT  3615.0 17355.0 3550.0 18240.0 ;
      RECT  3805.0 18240.0 3740.0 18375.0 ;
      RECT  3615.0 18240.0 3550.0 18375.0 ;
      RECT  3615.0 18240.0 3550.0 18375.0 ;
      RECT  3805.0 18240.0 3740.0 18375.0 ;
      RECT  3805.0 17355.0 3740.0 17490.0 ;
      RECT  3615.0 17355.0 3550.0 17490.0 ;
      RECT  3615.0 17355.0 3550.0 17490.0 ;
      RECT  3805.0 17355.0 3740.0 17490.0 ;
      RECT  3445.0 18330.0 3380.0 18465.0 ;
      RECT  3445.0 17355.0 3380.0 17490.0 ;
      RECT  3747.5 17797.5 3682.5 17932.5 ;
      RECT  3747.5 17797.5 3682.5 17932.5 ;
      RECT  3582.5 17832.5 3517.5 17897.5 ;
      RECT  3872.5 18550.0 3312.5 18615.0 ;
      RECT  3872.5 17205.0 3312.5 17270.0 ;
      RECT  3445.0 18767.5 3380.0 18582.5 ;
      RECT  3445.0 19927.5 3380.0 19742.5 ;
      RECT  3805.0 19810.0 3740.0 19960.0 ;
      RECT  3805.0 18925.0 3740.0 18550.0 ;
      RECT  3615.0 19810.0 3550.0 18925.0 ;
      RECT  3805.0 18925.0 3740.0 18790.0 ;
      RECT  3615.0 18925.0 3550.0 18790.0 ;
      RECT  3615.0 18925.0 3550.0 18790.0 ;
      RECT  3805.0 18925.0 3740.0 18790.0 ;
      RECT  3805.0 19810.0 3740.0 19675.0 ;
      RECT  3615.0 19810.0 3550.0 19675.0 ;
      RECT  3615.0 19810.0 3550.0 19675.0 ;
      RECT  3805.0 19810.0 3740.0 19675.0 ;
      RECT  3445.0 18835.0 3380.0 18700.0 ;
      RECT  3445.0 19810.0 3380.0 19675.0 ;
      RECT  3747.5 19367.5 3682.5 19232.5 ;
      RECT  3747.5 19367.5 3682.5 19232.5 ;
      RECT  3582.5 19332.5 3517.5 19267.5 ;
      RECT  3872.5 18615.0 3312.5 18550.0 ;
      RECT  3872.5 19960.0 3312.5 19895.0 ;
      RECT  4725.0 14710.0 4660.0 14515.0 ;
      RECT  4725.0 15550.0 4660.0 15925.0 ;
      RECT  4345.0 15550.0 4280.0 15925.0 ;
      RECT  4175.0 15707.5 4110.0 15892.5 ;
      RECT  4175.0 14547.5 4110.0 14732.5 ;
      RECT  4725.0 15550.0 4660.0 15685.0 ;
      RECT  4535.0 15550.0 4470.0 15685.0 ;
      RECT  4535.0 15550.0 4470.0 15685.0 ;
      RECT  4725.0 15550.0 4660.0 15685.0 ;
      RECT  4535.0 15550.0 4470.0 15685.0 ;
      RECT  4345.0 15550.0 4280.0 15685.0 ;
      RECT  4345.0 15550.0 4280.0 15685.0 ;
      RECT  4535.0 15550.0 4470.0 15685.0 ;
      RECT  4725.0 14710.0 4660.0 14845.0 ;
      RECT  4535.0 14710.0 4470.0 14845.0 ;
      RECT  4535.0 14710.0 4470.0 14845.0 ;
      RECT  4725.0 14710.0 4660.0 14845.0 ;
      RECT  4535.0 14710.0 4470.0 14845.0 ;
      RECT  4345.0 14710.0 4280.0 14845.0 ;
      RECT  4345.0 14710.0 4280.0 14845.0 ;
      RECT  4535.0 14710.0 4470.0 14845.0 ;
      RECT  4175.0 15640.0 4110.0 15775.0 ;
      RECT  4175.0 14665.0 4110.0 14800.0 ;
      RECT  4340.0 14940.0 4475.0 15005.0 ;
      RECT  4597.5 15155.0 4732.5 15220.0 ;
      RECT  4535.0 15550.0 4470.0 15685.0 ;
      RECT  4345.0 14710.0 4280.0 14845.0 ;
      RECT  4245.0 15155.0 4380.0 15220.0 ;
      RECT  4732.5 15155.0 4597.5 15220.0 ;
      RECT  4475.0 14940.0 4340.0 15005.0 ;
      RECT  4380.0 15155.0 4245.0 15220.0 ;
      RECT  4792.5 15860.0 3872.5 15925.0 ;
      RECT  4792.5 14515.0 3872.5 14580.0 ;
      RECT  4725.0 17075.0 4660.0 17270.0 ;
      RECT  4725.0 16235.0 4660.0 15860.0 ;
      RECT  4345.0 16235.0 4280.0 15860.0 ;
      RECT  4175.0 16077.5 4110.0 15892.5 ;
      RECT  4175.0 17237.5 4110.0 17052.5 ;
      RECT  4725.0 16235.0 4660.0 16100.0 ;
      RECT  4535.0 16235.0 4470.0 16100.0 ;
      RECT  4535.0 16235.0 4470.0 16100.0 ;
      RECT  4725.0 16235.0 4660.0 16100.0 ;
      RECT  4535.0 16235.0 4470.0 16100.0 ;
      RECT  4345.0 16235.0 4280.0 16100.0 ;
      RECT  4345.0 16235.0 4280.0 16100.0 ;
      RECT  4535.0 16235.0 4470.0 16100.0 ;
      RECT  4725.0 17075.0 4660.0 16940.0 ;
      RECT  4535.0 17075.0 4470.0 16940.0 ;
      RECT  4535.0 17075.0 4470.0 16940.0 ;
      RECT  4725.0 17075.0 4660.0 16940.0 ;
      RECT  4535.0 17075.0 4470.0 16940.0 ;
      RECT  4345.0 17075.0 4280.0 16940.0 ;
      RECT  4345.0 17075.0 4280.0 16940.0 ;
      RECT  4535.0 17075.0 4470.0 16940.0 ;
      RECT  4175.0 16145.0 4110.0 16010.0 ;
      RECT  4175.0 17120.0 4110.0 16985.0 ;
      RECT  4340.0 16845.0 4475.0 16780.0 ;
      RECT  4597.5 16630.0 4732.5 16565.0 ;
      RECT  4535.0 16235.0 4470.0 16100.0 ;
      RECT  4345.0 17075.0 4280.0 16940.0 ;
      RECT  4245.0 16630.0 4380.0 16565.0 ;
      RECT  4732.5 16630.0 4597.5 16565.0 ;
      RECT  4475.0 16845.0 4340.0 16780.0 ;
      RECT  4380.0 16630.0 4245.0 16565.0 ;
      RECT  4792.5 15925.0 3872.5 15860.0 ;
      RECT  4792.5 17270.0 3872.5 17205.0 ;
      RECT  4725.0 17400.0 4660.0 17205.0 ;
      RECT  4725.0 18240.0 4660.0 18615.0 ;
      RECT  4345.0 18240.0 4280.0 18615.0 ;
      RECT  4175.0 18397.5 4110.0 18582.5 ;
      RECT  4175.0 17237.5 4110.0 17422.5 ;
      RECT  4725.0 18240.0 4660.0 18375.0 ;
      RECT  4535.0 18240.0 4470.0 18375.0 ;
      RECT  4535.0 18240.0 4470.0 18375.0 ;
      RECT  4725.0 18240.0 4660.0 18375.0 ;
      RECT  4535.0 18240.0 4470.0 18375.0 ;
      RECT  4345.0 18240.0 4280.0 18375.0 ;
      RECT  4345.0 18240.0 4280.0 18375.0 ;
      RECT  4535.0 18240.0 4470.0 18375.0 ;
      RECT  4725.0 17400.0 4660.0 17535.0 ;
      RECT  4535.0 17400.0 4470.0 17535.0 ;
      RECT  4535.0 17400.0 4470.0 17535.0 ;
      RECT  4725.0 17400.0 4660.0 17535.0 ;
      RECT  4535.0 17400.0 4470.0 17535.0 ;
      RECT  4345.0 17400.0 4280.0 17535.0 ;
      RECT  4345.0 17400.0 4280.0 17535.0 ;
      RECT  4535.0 17400.0 4470.0 17535.0 ;
      RECT  4175.0 18330.0 4110.0 18465.0 ;
      RECT  4175.0 17355.0 4110.0 17490.0 ;
      RECT  4340.0 17630.0 4475.0 17695.0 ;
      RECT  4597.5 17845.0 4732.5 17910.0 ;
      RECT  4535.0 18240.0 4470.0 18375.0 ;
      RECT  4345.0 17400.0 4280.0 17535.0 ;
      RECT  4245.0 17845.0 4380.0 17910.0 ;
      RECT  4732.5 17845.0 4597.5 17910.0 ;
      RECT  4475.0 17630.0 4340.0 17695.0 ;
      RECT  4380.0 17845.0 4245.0 17910.0 ;
      RECT  4792.5 18550.0 3872.5 18615.0 ;
      RECT  4792.5 17205.0 3872.5 17270.0 ;
      RECT  4725.0 19765.0 4660.0 19960.0 ;
      RECT  4725.0 18925.0 4660.0 18550.0 ;
      RECT  4345.0 18925.0 4280.0 18550.0 ;
      RECT  4175.0 18767.5 4110.0 18582.5 ;
      RECT  4175.0 19927.5 4110.0 19742.5 ;
      RECT  4725.0 18925.0 4660.0 18790.0 ;
      RECT  4535.0 18925.0 4470.0 18790.0 ;
      RECT  4535.0 18925.0 4470.0 18790.0 ;
      RECT  4725.0 18925.0 4660.0 18790.0 ;
      RECT  4535.0 18925.0 4470.0 18790.0 ;
      RECT  4345.0 18925.0 4280.0 18790.0 ;
      RECT  4345.0 18925.0 4280.0 18790.0 ;
      RECT  4535.0 18925.0 4470.0 18790.0 ;
      RECT  4725.0 19765.0 4660.0 19630.0 ;
      RECT  4535.0 19765.0 4470.0 19630.0 ;
      RECT  4535.0 19765.0 4470.0 19630.0 ;
      RECT  4725.0 19765.0 4660.0 19630.0 ;
      RECT  4535.0 19765.0 4470.0 19630.0 ;
      RECT  4345.0 19765.0 4280.0 19630.0 ;
      RECT  4345.0 19765.0 4280.0 19630.0 ;
      RECT  4535.0 19765.0 4470.0 19630.0 ;
      RECT  4175.0 18835.0 4110.0 18700.0 ;
      RECT  4175.0 19810.0 4110.0 19675.0 ;
      RECT  4340.0 19535.0 4475.0 19470.0 ;
      RECT  4597.5 19320.0 4732.5 19255.0 ;
      RECT  4535.0 18925.0 4470.0 18790.0 ;
      RECT  4345.0 19765.0 4280.0 19630.0 ;
      RECT  4245.0 19320.0 4380.0 19255.0 ;
      RECT  4732.5 19320.0 4597.5 19255.0 ;
      RECT  4475.0 19535.0 4340.0 19470.0 ;
      RECT  4380.0 19320.0 4245.0 19255.0 ;
      RECT  4792.5 18615.0 3872.5 18550.0 ;
      RECT  4792.5 19960.0 3872.5 19895.0 ;
      RECT  5790.0 15665.0 5925.0 15730.0 ;
      RECT  7175.0 15142.5 7310.0 15207.5 ;
      RECT  5515.0 17010.0 5650.0 17075.0 ;
      RECT  6900.0 16577.5 7035.0 16642.5 ;
      RECT  7175.0 17340.0 7310.0 17405.0 ;
      RECT  5240.0 17340.0 5375.0 17405.0 ;
      RECT  6900.0 18685.0 7035.0 18750.0 ;
      RECT  4965.0 18685.0 5100.0 18750.0 ;
      RECT  5790.0 15155.0 5925.0 15220.0 ;
      RECT  5515.0 14940.0 5650.0 15005.0 ;
      RECT  5240.0 16565.0 5375.0 16630.0 ;
      RECT  5515.0 16780.0 5650.0 16845.0 ;
      RECT  5790.0 17845.0 5925.0 17910.0 ;
      RECT  4965.0 17630.0 5100.0 17695.0 ;
      RECT  5240.0 19255.0 5375.0 19320.0 ;
      RECT  4965.0 19470.0 5100.0 19535.0 ;
      RECT  3517.5 15142.5 3312.5 15207.5 ;
      RECT  3517.5 16577.5 3312.5 16642.5 ;
      RECT  3517.5 17832.5 3312.5 17897.5 ;
      RECT  3517.5 19267.5 3312.5 19332.5 ;
      RECT  7277.5 15860.0 3312.5 15925.0 ;
      RECT  7277.5 18550.0 3312.5 18615.0 ;
      RECT  7277.5 14515.0 3312.5 14580.0 ;
      RECT  7277.5 17205.0 3312.5 17270.0 ;
      RECT  7277.5 19895.0 3312.5 19960.0 ;
      RECT  3380.0 20090.0 3445.0 19895.0 ;
      RECT  3380.0 20930.0 3445.0 21305.0 ;
      RECT  3760.0 20930.0 3825.0 21305.0 ;
      RECT  3930.0 21087.5 3995.0 21272.5 ;
      RECT  3930.0 19927.5 3995.0 20112.5 ;
      RECT  3380.0 20930.0 3445.0 21065.0 ;
      RECT  3570.0 20930.0 3635.0 21065.0 ;
      RECT  3570.0 20930.0 3635.0 21065.0 ;
      RECT  3380.0 20930.0 3445.0 21065.0 ;
      RECT  3570.0 20930.0 3635.0 21065.0 ;
      RECT  3760.0 20930.0 3825.0 21065.0 ;
      RECT  3760.0 20930.0 3825.0 21065.0 ;
      RECT  3570.0 20930.0 3635.0 21065.0 ;
      RECT  3380.0 20090.0 3445.0 20225.0 ;
      RECT  3570.0 20090.0 3635.0 20225.0 ;
      RECT  3570.0 20090.0 3635.0 20225.0 ;
      RECT  3380.0 20090.0 3445.0 20225.0 ;
      RECT  3570.0 20090.0 3635.0 20225.0 ;
      RECT  3760.0 20090.0 3825.0 20225.0 ;
      RECT  3760.0 20090.0 3825.0 20225.0 ;
      RECT  3570.0 20090.0 3635.0 20225.0 ;
      RECT  3930.0 21020.0 3995.0 21155.0 ;
      RECT  3930.0 20045.0 3995.0 20180.0 ;
      RECT  3765.0 20320.0 3630.0 20385.0 ;
      RECT  3507.5 20535.0 3372.5 20600.0 ;
      RECT  3570.0 20930.0 3635.0 21065.0 ;
      RECT  3760.0 20090.0 3825.0 20225.0 ;
      RECT  3860.0 20535.0 3725.0 20600.0 ;
      RECT  3372.5 20535.0 3507.5 20600.0 ;
      RECT  3630.0 20320.0 3765.0 20385.0 ;
      RECT  3725.0 20535.0 3860.0 20600.0 ;
      RECT  3312.5 21240.0 4232.5 21305.0 ;
      RECT  3312.5 19895.0 4232.5 19960.0 ;
      RECT  3380.0 22455.0 3445.0 22650.0 ;
      RECT  3380.0 21615.0 3445.0 21240.0 ;
      RECT  3760.0 21615.0 3825.0 21240.0 ;
      RECT  3930.0 21457.5 3995.0 21272.5 ;
      RECT  3930.0 22617.5 3995.0 22432.5 ;
      RECT  3380.0 21615.0 3445.0 21480.0 ;
      RECT  3570.0 21615.0 3635.0 21480.0 ;
      RECT  3570.0 21615.0 3635.0 21480.0 ;
      RECT  3380.0 21615.0 3445.0 21480.0 ;
      RECT  3570.0 21615.0 3635.0 21480.0 ;
      RECT  3760.0 21615.0 3825.0 21480.0 ;
      RECT  3760.0 21615.0 3825.0 21480.0 ;
      RECT  3570.0 21615.0 3635.0 21480.0 ;
      RECT  3380.0 22455.0 3445.0 22320.0 ;
      RECT  3570.0 22455.0 3635.0 22320.0 ;
      RECT  3570.0 22455.0 3635.0 22320.0 ;
      RECT  3380.0 22455.0 3445.0 22320.0 ;
      RECT  3570.0 22455.0 3635.0 22320.0 ;
      RECT  3760.0 22455.0 3825.0 22320.0 ;
      RECT  3760.0 22455.0 3825.0 22320.0 ;
      RECT  3570.0 22455.0 3635.0 22320.0 ;
      RECT  3930.0 21525.0 3995.0 21390.0 ;
      RECT  3930.0 22500.0 3995.0 22365.0 ;
      RECT  3765.0 22225.0 3630.0 22160.0 ;
      RECT  3507.5 22010.0 3372.5 21945.0 ;
      RECT  3570.0 21615.0 3635.0 21480.0 ;
      RECT  3760.0 22455.0 3825.0 22320.0 ;
      RECT  3860.0 22010.0 3725.0 21945.0 ;
      RECT  3372.5 22010.0 3507.5 21945.0 ;
      RECT  3630.0 22225.0 3765.0 22160.0 ;
      RECT  3725.0 22010.0 3860.0 21945.0 ;
      RECT  3312.5 21305.0 4232.5 21240.0 ;
      RECT  3312.5 22650.0 4232.5 22585.0 ;
      RECT  3380.0 22780.0 3445.0 22585.0 ;
      RECT  3380.0 23620.0 3445.0 23995.0 ;
      RECT  3760.0 23620.0 3825.0 23995.0 ;
      RECT  3930.0 23777.5 3995.0 23962.5 ;
      RECT  3930.0 22617.5 3995.0 22802.5 ;
      RECT  3380.0 23620.0 3445.0 23755.0 ;
      RECT  3570.0 23620.0 3635.0 23755.0 ;
      RECT  3570.0 23620.0 3635.0 23755.0 ;
      RECT  3380.0 23620.0 3445.0 23755.0 ;
      RECT  3570.0 23620.0 3635.0 23755.0 ;
      RECT  3760.0 23620.0 3825.0 23755.0 ;
      RECT  3760.0 23620.0 3825.0 23755.0 ;
      RECT  3570.0 23620.0 3635.0 23755.0 ;
      RECT  3380.0 22780.0 3445.0 22915.0 ;
      RECT  3570.0 22780.0 3635.0 22915.0 ;
      RECT  3570.0 22780.0 3635.0 22915.0 ;
      RECT  3380.0 22780.0 3445.0 22915.0 ;
      RECT  3570.0 22780.0 3635.0 22915.0 ;
      RECT  3760.0 22780.0 3825.0 22915.0 ;
      RECT  3760.0 22780.0 3825.0 22915.0 ;
      RECT  3570.0 22780.0 3635.0 22915.0 ;
      RECT  3930.0 23710.0 3995.0 23845.0 ;
      RECT  3930.0 22735.0 3995.0 22870.0 ;
      RECT  3765.0 23010.0 3630.0 23075.0 ;
      RECT  3507.5 23225.0 3372.5 23290.0 ;
      RECT  3570.0 23620.0 3635.0 23755.0 ;
      RECT  3760.0 22780.0 3825.0 22915.0 ;
      RECT  3860.0 23225.0 3725.0 23290.0 ;
      RECT  3372.5 23225.0 3507.5 23290.0 ;
      RECT  3630.0 23010.0 3765.0 23075.0 ;
      RECT  3725.0 23225.0 3860.0 23290.0 ;
      RECT  3312.5 23930.0 4232.5 23995.0 ;
      RECT  3312.5 22585.0 4232.5 22650.0 ;
      RECT  3380.0 25145.0 3445.0 25340.0 ;
      RECT  3380.0 24305.0 3445.0 23930.0 ;
      RECT  3760.0 24305.0 3825.0 23930.0 ;
      RECT  3930.0 24147.5 3995.0 23962.5 ;
      RECT  3930.0 25307.5 3995.0 25122.5 ;
      RECT  3380.0 24305.0 3445.0 24170.0 ;
      RECT  3570.0 24305.0 3635.0 24170.0 ;
      RECT  3570.0 24305.0 3635.0 24170.0 ;
      RECT  3380.0 24305.0 3445.0 24170.0 ;
      RECT  3570.0 24305.0 3635.0 24170.0 ;
      RECT  3760.0 24305.0 3825.0 24170.0 ;
      RECT  3760.0 24305.0 3825.0 24170.0 ;
      RECT  3570.0 24305.0 3635.0 24170.0 ;
      RECT  3380.0 25145.0 3445.0 25010.0 ;
      RECT  3570.0 25145.0 3635.0 25010.0 ;
      RECT  3570.0 25145.0 3635.0 25010.0 ;
      RECT  3380.0 25145.0 3445.0 25010.0 ;
      RECT  3570.0 25145.0 3635.0 25010.0 ;
      RECT  3760.0 25145.0 3825.0 25010.0 ;
      RECT  3760.0 25145.0 3825.0 25010.0 ;
      RECT  3570.0 25145.0 3635.0 25010.0 ;
      RECT  3930.0 24215.0 3995.0 24080.0 ;
      RECT  3930.0 25190.0 3995.0 25055.0 ;
      RECT  3765.0 24915.0 3630.0 24850.0 ;
      RECT  3507.5 24700.0 3372.5 24635.0 ;
      RECT  3570.0 24305.0 3635.0 24170.0 ;
      RECT  3760.0 25145.0 3825.0 25010.0 ;
      RECT  3860.0 24700.0 3725.0 24635.0 ;
      RECT  3372.5 24700.0 3507.5 24635.0 ;
      RECT  3630.0 24915.0 3765.0 24850.0 ;
      RECT  3725.0 24700.0 3860.0 24635.0 ;
      RECT  3312.5 23995.0 4232.5 23930.0 ;
      RECT  3312.5 25340.0 4232.5 25275.0 ;
      RECT  3380.0 25470.0 3445.0 25275.0 ;
      RECT  3380.0 26310.0 3445.0 26685.0 ;
      RECT  3760.0 26310.0 3825.0 26685.0 ;
      RECT  3930.0 26467.5 3995.0 26652.5 ;
      RECT  3930.0 25307.5 3995.0 25492.5 ;
      RECT  3380.0 26310.0 3445.0 26445.0 ;
      RECT  3570.0 26310.0 3635.0 26445.0 ;
      RECT  3570.0 26310.0 3635.0 26445.0 ;
      RECT  3380.0 26310.0 3445.0 26445.0 ;
      RECT  3570.0 26310.0 3635.0 26445.0 ;
      RECT  3760.0 26310.0 3825.0 26445.0 ;
      RECT  3760.0 26310.0 3825.0 26445.0 ;
      RECT  3570.0 26310.0 3635.0 26445.0 ;
      RECT  3380.0 25470.0 3445.0 25605.0 ;
      RECT  3570.0 25470.0 3635.0 25605.0 ;
      RECT  3570.0 25470.0 3635.0 25605.0 ;
      RECT  3380.0 25470.0 3445.0 25605.0 ;
      RECT  3570.0 25470.0 3635.0 25605.0 ;
      RECT  3760.0 25470.0 3825.0 25605.0 ;
      RECT  3760.0 25470.0 3825.0 25605.0 ;
      RECT  3570.0 25470.0 3635.0 25605.0 ;
      RECT  3930.0 26400.0 3995.0 26535.0 ;
      RECT  3930.0 25425.0 3995.0 25560.0 ;
      RECT  3765.0 25700.0 3630.0 25765.0 ;
      RECT  3507.5 25915.0 3372.5 25980.0 ;
      RECT  3570.0 26310.0 3635.0 26445.0 ;
      RECT  3760.0 25470.0 3825.0 25605.0 ;
      RECT  3860.0 25915.0 3725.0 25980.0 ;
      RECT  3372.5 25915.0 3507.5 25980.0 ;
      RECT  3630.0 25700.0 3765.0 25765.0 ;
      RECT  3725.0 25915.0 3860.0 25980.0 ;
      RECT  3312.5 26620.0 4232.5 26685.0 ;
      RECT  3312.5 25275.0 4232.5 25340.0 ;
      RECT  3380.0 27835.0 3445.0 28030.0 ;
      RECT  3380.0 26995.0 3445.0 26620.0 ;
      RECT  3760.0 26995.0 3825.0 26620.0 ;
      RECT  3930.0 26837.5 3995.0 26652.5 ;
      RECT  3930.0 27997.5 3995.0 27812.5 ;
      RECT  3380.0 26995.0 3445.0 26860.0 ;
      RECT  3570.0 26995.0 3635.0 26860.0 ;
      RECT  3570.0 26995.0 3635.0 26860.0 ;
      RECT  3380.0 26995.0 3445.0 26860.0 ;
      RECT  3570.0 26995.0 3635.0 26860.0 ;
      RECT  3760.0 26995.0 3825.0 26860.0 ;
      RECT  3760.0 26995.0 3825.0 26860.0 ;
      RECT  3570.0 26995.0 3635.0 26860.0 ;
      RECT  3380.0 27835.0 3445.0 27700.0 ;
      RECT  3570.0 27835.0 3635.0 27700.0 ;
      RECT  3570.0 27835.0 3635.0 27700.0 ;
      RECT  3380.0 27835.0 3445.0 27700.0 ;
      RECT  3570.0 27835.0 3635.0 27700.0 ;
      RECT  3760.0 27835.0 3825.0 27700.0 ;
      RECT  3760.0 27835.0 3825.0 27700.0 ;
      RECT  3570.0 27835.0 3635.0 27700.0 ;
      RECT  3930.0 26905.0 3995.0 26770.0 ;
      RECT  3930.0 27880.0 3995.0 27745.0 ;
      RECT  3765.0 27605.0 3630.0 27540.0 ;
      RECT  3507.5 27390.0 3372.5 27325.0 ;
      RECT  3570.0 26995.0 3635.0 26860.0 ;
      RECT  3760.0 27835.0 3825.0 27700.0 ;
      RECT  3860.0 27390.0 3725.0 27325.0 ;
      RECT  3372.5 27390.0 3507.5 27325.0 ;
      RECT  3630.0 27605.0 3765.0 27540.0 ;
      RECT  3725.0 27390.0 3860.0 27325.0 ;
      RECT  3312.5 26685.0 4232.5 26620.0 ;
      RECT  3312.5 28030.0 4232.5 27965.0 ;
      RECT  3380.0 28160.0 3445.0 27965.0 ;
      RECT  3380.0 29000.0 3445.0 29375.0 ;
      RECT  3760.0 29000.0 3825.0 29375.0 ;
      RECT  3930.0 29157.5 3995.0 29342.5 ;
      RECT  3930.0 27997.5 3995.0 28182.5 ;
      RECT  3380.0 29000.0 3445.0 29135.0 ;
      RECT  3570.0 29000.0 3635.0 29135.0 ;
      RECT  3570.0 29000.0 3635.0 29135.0 ;
      RECT  3380.0 29000.0 3445.0 29135.0 ;
      RECT  3570.0 29000.0 3635.0 29135.0 ;
      RECT  3760.0 29000.0 3825.0 29135.0 ;
      RECT  3760.0 29000.0 3825.0 29135.0 ;
      RECT  3570.0 29000.0 3635.0 29135.0 ;
      RECT  3380.0 28160.0 3445.0 28295.0 ;
      RECT  3570.0 28160.0 3635.0 28295.0 ;
      RECT  3570.0 28160.0 3635.0 28295.0 ;
      RECT  3380.0 28160.0 3445.0 28295.0 ;
      RECT  3570.0 28160.0 3635.0 28295.0 ;
      RECT  3760.0 28160.0 3825.0 28295.0 ;
      RECT  3760.0 28160.0 3825.0 28295.0 ;
      RECT  3570.0 28160.0 3635.0 28295.0 ;
      RECT  3930.0 29090.0 3995.0 29225.0 ;
      RECT  3930.0 28115.0 3995.0 28250.0 ;
      RECT  3765.0 28390.0 3630.0 28455.0 ;
      RECT  3507.5 28605.0 3372.5 28670.0 ;
      RECT  3570.0 29000.0 3635.0 29135.0 ;
      RECT  3760.0 28160.0 3825.0 28295.0 ;
      RECT  3860.0 28605.0 3725.0 28670.0 ;
      RECT  3372.5 28605.0 3507.5 28670.0 ;
      RECT  3630.0 28390.0 3765.0 28455.0 ;
      RECT  3725.0 28605.0 3860.0 28670.0 ;
      RECT  3312.5 29310.0 4232.5 29375.0 ;
      RECT  3312.5 27965.0 4232.5 28030.0 ;
      RECT  3380.0 30525.0 3445.0 30720.0 ;
      RECT  3380.0 29685.0 3445.0 29310.0 ;
      RECT  3760.0 29685.0 3825.0 29310.0 ;
      RECT  3930.0 29527.5 3995.0 29342.5 ;
      RECT  3930.0 30687.5 3995.0 30502.5 ;
      RECT  3380.0 29685.0 3445.0 29550.0 ;
      RECT  3570.0 29685.0 3635.0 29550.0 ;
      RECT  3570.0 29685.0 3635.0 29550.0 ;
      RECT  3380.0 29685.0 3445.0 29550.0 ;
      RECT  3570.0 29685.0 3635.0 29550.0 ;
      RECT  3760.0 29685.0 3825.0 29550.0 ;
      RECT  3760.0 29685.0 3825.0 29550.0 ;
      RECT  3570.0 29685.0 3635.0 29550.0 ;
      RECT  3380.0 30525.0 3445.0 30390.0 ;
      RECT  3570.0 30525.0 3635.0 30390.0 ;
      RECT  3570.0 30525.0 3635.0 30390.0 ;
      RECT  3380.0 30525.0 3445.0 30390.0 ;
      RECT  3570.0 30525.0 3635.0 30390.0 ;
      RECT  3760.0 30525.0 3825.0 30390.0 ;
      RECT  3760.0 30525.0 3825.0 30390.0 ;
      RECT  3570.0 30525.0 3635.0 30390.0 ;
      RECT  3930.0 29595.0 3995.0 29460.0 ;
      RECT  3930.0 30570.0 3995.0 30435.0 ;
      RECT  3765.0 30295.0 3630.0 30230.0 ;
      RECT  3507.5 30080.0 3372.5 30015.0 ;
      RECT  3570.0 29685.0 3635.0 29550.0 ;
      RECT  3760.0 30525.0 3825.0 30390.0 ;
      RECT  3860.0 30080.0 3725.0 30015.0 ;
      RECT  3372.5 30080.0 3507.5 30015.0 ;
      RECT  3630.0 30295.0 3765.0 30230.0 ;
      RECT  3725.0 30080.0 3860.0 30015.0 ;
      RECT  3312.5 29375.0 4232.5 29310.0 ;
      RECT  3312.5 30720.0 4232.5 30655.0 ;
      RECT  3380.0 30850.0 3445.0 30655.0 ;
      RECT  3380.0 31690.0 3445.0 32065.0 ;
      RECT  3760.0 31690.0 3825.0 32065.0 ;
      RECT  3930.0 31847.5 3995.0 32032.5 ;
      RECT  3930.0 30687.5 3995.0 30872.5 ;
      RECT  3380.0 31690.0 3445.0 31825.0 ;
      RECT  3570.0 31690.0 3635.0 31825.0 ;
      RECT  3570.0 31690.0 3635.0 31825.0 ;
      RECT  3380.0 31690.0 3445.0 31825.0 ;
      RECT  3570.0 31690.0 3635.0 31825.0 ;
      RECT  3760.0 31690.0 3825.0 31825.0 ;
      RECT  3760.0 31690.0 3825.0 31825.0 ;
      RECT  3570.0 31690.0 3635.0 31825.0 ;
      RECT  3380.0 30850.0 3445.0 30985.0 ;
      RECT  3570.0 30850.0 3635.0 30985.0 ;
      RECT  3570.0 30850.0 3635.0 30985.0 ;
      RECT  3380.0 30850.0 3445.0 30985.0 ;
      RECT  3570.0 30850.0 3635.0 30985.0 ;
      RECT  3760.0 30850.0 3825.0 30985.0 ;
      RECT  3760.0 30850.0 3825.0 30985.0 ;
      RECT  3570.0 30850.0 3635.0 30985.0 ;
      RECT  3930.0 31780.0 3995.0 31915.0 ;
      RECT  3930.0 30805.0 3995.0 30940.0 ;
      RECT  3765.0 31080.0 3630.0 31145.0 ;
      RECT  3507.5 31295.0 3372.5 31360.0 ;
      RECT  3570.0 31690.0 3635.0 31825.0 ;
      RECT  3760.0 30850.0 3825.0 30985.0 ;
      RECT  3860.0 31295.0 3725.0 31360.0 ;
      RECT  3372.5 31295.0 3507.5 31360.0 ;
      RECT  3630.0 31080.0 3765.0 31145.0 ;
      RECT  3725.0 31295.0 3860.0 31360.0 ;
      RECT  3312.5 32000.0 4232.5 32065.0 ;
      RECT  3312.5 30655.0 4232.5 30720.0 ;
      RECT  3380.0 33215.0 3445.0 33410.0 ;
      RECT  3380.0 32375.0 3445.0 32000.0 ;
      RECT  3760.0 32375.0 3825.0 32000.0 ;
      RECT  3930.0 32217.5 3995.0 32032.5 ;
      RECT  3930.0 33377.5 3995.0 33192.5 ;
      RECT  3380.0 32375.0 3445.0 32240.0 ;
      RECT  3570.0 32375.0 3635.0 32240.0 ;
      RECT  3570.0 32375.0 3635.0 32240.0 ;
      RECT  3380.0 32375.0 3445.0 32240.0 ;
      RECT  3570.0 32375.0 3635.0 32240.0 ;
      RECT  3760.0 32375.0 3825.0 32240.0 ;
      RECT  3760.0 32375.0 3825.0 32240.0 ;
      RECT  3570.0 32375.0 3635.0 32240.0 ;
      RECT  3380.0 33215.0 3445.0 33080.0 ;
      RECT  3570.0 33215.0 3635.0 33080.0 ;
      RECT  3570.0 33215.0 3635.0 33080.0 ;
      RECT  3380.0 33215.0 3445.0 33080.0 ;
      RECT  3570.0 33215.0 3635.0 33080.0 ;
      RECT  3760.0 33215.0 3825.0 33080.0 ;
      RECT  3760.0 33215.0 3825.0 33080.0 ;
      RECT  3570.0 33215.0 3635.0 33080.0 ;
      RECT  3930.0 32285.0 3995.0 32150.0 ;
      RECT  3930.0 33260.0 3995.0 33125.0 ;
      RECT  3765.0 32985.0 3630.0 32920.0 ;
      RECT  3507.5 32770.0 3372.5 32705.0 ;
      RECT  3570.0 32375.0 3635.0 32240.0 ;
      RECT  3760.0 33215.0 3825.0 33080.0 ;
      RECT  3860.0 32770.0 3725.0 32705.0 ;
      RECT  3372.5 32770.0 3507.5 32705.0 ;
      RECT  3630.0 32985.0 3765.0 32920.0 ;
      RECT  3725.0 32770.0 3860.0 32705.0 ;
      RECT  3312.5 32065.0 4232.5 32000.0 ;
      RECT  3312.5 33410.0 4232.5 33345.0 ;
      RECT  3380.0 33540.0 3445.0 33345.0 ;
      RECT  3380.0 34380.0 3445.0 34755.0 ;
      RECT  3760.0 34380.0 3825.0 34755.0 ;
      RECT  3930.0 34537.5 3995.0 34722.5 ;
      RECT  3930.0 33377.5 3995.0 33562.5 ;
      RECT  3380.0 34380.0 3445.0 34515.0 ;
      RECT  3570.0 34380.0 3635.0 34515.0 ;
      RECT  3570.0 34380.0 3635.0 34515.0 ;
      RECT  3380.0 34380.0 3445.0 34515.0 ;
      RECT  3570.0 34380.0 3635.0 34515.0 ;
      RECT  3760.0 34380.0 3825.0 34515.0 ;
      RECT  3760.0 34380.0 3825.0 34515.0 ;
      RECT  3570.0 34380.0 3635.0 34515.0 ;
      RECT  3380.0 33540.0 3445.0 33675.0 ;
      RECT  3570.0 33540.0 3635.0 33675.0 ;
      RECT  3570.0 33540.0 3635.0 33675.0 ;
      RECT  3380.0 33540.0 3445.0 33675.0 ;
      RECT  3570.0 33540.0 3635.0 33675.0 ;
      RECT  3760.0 33540.0 3825.0 33675.0 ;
      RECT  3760.0 33540.0 3825.0 33675.0 ;
      RECT  3570.0 33540.0 3635.0 33675.0 ;
      RECT  3930.0 34470.0 3995.0 34605.0 ;
      RECT  3930.0 33495.0 3995.0 33630.0 ;
      RECT  3765.0 33770.0 3630.0 33835.0 ;
      RECT  3507.5 33985.0 3372.5 34050.0 ;
      RECT  3570.0 34380.0 3635.0 34515.0 ;
      RECT  3760.0 33540.0 3825.0 33675.0 ;
      RECT  3860.0 33985.0 3725.0 34050.0 ;
      RECT  3372.5 33985.0 3507.5 34050.0 ;
      RECT  3630.0 33770.0 3765.0 33835.0 ;
      RECT  3725.0 33985.0 3860.0 34050.0 ;
      RECT  3312.5 34690.0 4232.5 34755.0 ;
      RECT  3312.5 33345.0 4232.5 33410.0 ;
      RECT  3380.0 35905.0 3445.0 36100.0 ;
      RECT  3380.0 35065.0 3445.0 34690.0 ;
      RECT  3760.0 35065.0 3825.0 34690.0 ;
      RECT  3930.0 34907.5 3995.0 34722.5 ;
      RECT  3930.0 36067.5 3995.0 35882.5 ;
      RECT  3380.0 35065.0 3445.0 34930.0 ;
      RECT  3570.0 35065.0 3635.0 34930.0 ;
      RECT  3570.0 35065.0 3635.0 34930.0 ;
      RECT  3380.0 35065.0 3445.0 34930.0 ;
      RECT  3570.0 35065.0 3635.0 34930.0 ;
      RECT  3760.0 35065.0 3825.0 34930.0 ;
      RECT  3760.0 35065.0 3825.0 34930.0 ;
      RECT  3570.0 35065.0 3635.0 34930.0 ;
      RECT  3380.0 35905.0 3445.0 35770.0 ;
      RECT  3570.0 35905.0 3635.0 35770.0 ;
      RECT  3570.0 35905.0 3635.0 35770.0 ;
      RECT  3380.0 35905.0 3445.0 35770.0 ;
      RECT  3570.0 35905.0 3635.0 35770.0 ;
      RECT  3760.0 35905.0 3825.0 35770.0 ;
      RECT  3760.0 35905.0 3825.0 35770.0 ;
      RECT  3570.0 35905.0 3635.0 35770.0 ;
      RECT  3930.0 34975.0 3995.0 34840.0 ;
      RECT  3930.0 35950.0 3995.0 35815.0 ;
      RECT  3765.0 35675.0 3630.0 35610.0 ;
      RECT  3507.5 35460.0 3372.5 35395.0 ;
      RECT  3570.0 35065.0 3635.0 34930.0 ;
      RECT  3760.0 35905.0 3825.0 35770.0 ;
      RECT  3860.0 35460.0 3725.0 35395.0 ;
      RECT  3372.5 35460.0 3507.5 35395.0 ;
      RECT  3630.0 35675.0 3765.0 35610.0 ;
      RECT  3725.0 35460.0 3860.0 35395.0 ;
      RECT  3312.5 34755.0 4232.5 34690.0 ;
      RECT  3312.5 36100.0 4232.5 36035.0 ;
      RECT  3380.0 36230.0 3445.0 36035.0 ;
      RECT  3380.0 37070.0 3445.0 37445.0 ;
      RECT  3760.0 37070.0 3825.0 37445.0 ;
      RECT  3930.0 37227.5 3995.0 37412.5 ;
      RECT  3930.0 36067.5 3995.0 36252.5 ;
      RECT  3380.0 37070.0 3445.0 37205.0 ;
      RECT  3570.0 37070.0 3635.0 37205.0 ;
      RECT  3570.0 37070.0 3635.0 37205.0 ;
      RECT  3380.0 37070.0 3445.0 37205.0 ;
      RECT  3570.0 37070.0 3635.0 37205.0 ;
      RECT  3760.0 37070.0 3825.0 37205.0 ;
      RECT  3760.0 37070.0 3825.0 37205.0 ;
      RECT  3570.0 37070.0 3635.0 37205.0 ;
      RECT  3380.0 36230.0 3445.0 36365.0 ;
      RECT  3570.0 36230.0 3635.0 36365.0 ;
      RECT  3570.0 36230.0 3635.0 36365.0 ;
      RECT  3380.0 36230.0 3445.0 36365.0 ;
      RECT  3570.0 36230.0 3635.0 36365.0 ;
      RECT  3760.0 36230.0 3825.0 36365.0 ;
      RECT  3760.0 36230.0 3825.0 36365.0 ;
      RECT  3570.0 36230.0 3635.0 36365.0 ;
      RECT  3930.0 37160.0 3995.0 37295.0 ;
      RECT  3930.0 36185.0 3995.0 36320.0 ;
      RECT  3765.0 36460.0 3630.0 36525.0 ;
      RECT  3507.5 36675.0 3372.5 36740.0 ;
      RECT  3570.0 37070.0 3635.0 37205.0 ;
      RECT  3760.0 36230.0 3825.0 36365.0 ;
      RECT  3860.0 36675.0 3725.0 36740.0 ;
      RECT  3372.5 36675.0 3507.5 36740.0 ;
      RECT  3630.0 36460.0 3765.0 36525.0 ;
      RECT  3725.0 36675.0 3860.0 36740.0 ;
      RECT  3312.5 37380.0 4232.5 37445.0 ;
      RECT  3312.5 36035.0 4232.5 36100.0 ;
      RECT  3380.0 38595.0 3445.0 38790.0 ;
      RECT  3380.0 37755.0 3445.0 37380.0 ;
      RECT  3760.0 37755.0 3825.0 37380.0 ;
      RECT  3930.0 37597.5 3995.0 37412.5 ;
      RECT  3930.0 38757.5 3995.0 38572.5 ;
      RECT  3380.0 37755.0 3445.0 37620.0 ;
      RECT  3570.0 37755.0 3635.0 37620.0 ;
      RECT  3570.0 37755.0 3635.0 37620.0 ;
      RECT  3380.0 37755.0 3445.0 37620.0 ;
      RECT  3570.0 37755.0 3635.0 37620.0 ;
      RECT  3760.0 37755.0 3825.0 37620.0 ;
      RECT  3760.0 37755.0 3825.0 37620.0 ;
      RECT  3570.0 37755.0 3635.0 37620.0 ;
      RECT  3380.0 38595.0 3445.0 38460.0 ;
      RECT  3570.0 38595.0 3635.0 38460.0 ;
      RECT  3570.0 38595.0 3635.0 38460.0 ;
      RECT  3380.0 38595.0 3445.0 38460.0 ;
      RECT  3570.0 38595.0 3635.0 38460.0 ;
      RECT  3760.0 38595.0 3825.0 38460.0 ;
      RECT  3760.0 38595.0 3825.0 38460.0 ;
      RECT  3570.0 38595.0 3635.0 38460.0 ;
      RECT  3930.0 37665.0 3995.0 37530.0 ;
      RECT  3930.0 38640.0 3995.0 38505.0 ;
      RECT  3765.0 38365.0 3630.0 38300.0 ;
      RECT  3507.5 38150.0 3372.5 38085.0 ;
      RECT  3570.0 37755.0 3635.0 37620.0 ;
      RECT  3760.0 38595.0 3825.0 38460.0 ;
      RECT  3860.0 38150.0 3725.0 38085.0 ;
      RECT  3372.5 38150.0 3507.5 38085.0 ;
      RECT  3630.0 38365.0 3765.0 38300.0 ;
      RECT  3725.0 38150.0 3860.0 38085.0 ;
      RECT  3312.5 37445.0 4232.5 37380.0 ;
      RECT  3312.5 38790.0 4232.5 38725.0 ;
      RECT  3380.0 38920.0 3445.0 38725.0 ;
      RECT  3380.0 39760.0 3445.0 40135.0 ;
      RECT  3760.0 39760.0 3825.0 40135.0 ;
      RECT  3930.0 39917.5 3995.0 40102.5 ;
      RECT  3930.0 38757.5 3995.0 38942.5 ;
      RECT  3380.0 39760.0 3445.0 39895.0 ;
      RECT  3570.0 39760.0 3635.0 39895.0 ;
      RECT  3570.0 39760.0 3635.0 39895.0 ;
      RECT  3380.0 39760.0 3445.0 39895.0 ;
      RECT  3570.0 39760.0 3635.0 39895.0 ;
      RECT  3760.0 39760.0 3825.0 39895.0 ;
      RECT  3760.0 39760.0 3825.0 39895.0 ;
      RECT  3570.0 39760.0 3635.0 39895.0 ;
      RECT  3380.0 38920.0 3445.0 39055.0 ;
      RECT  3570.0 38920.0 3635.0 39055.0 ;
      RECT  3570.0 38920.0 3635.0 39055.0 ;
      RECT  3380.0 38920.0 3445.0 39055.0 ;
      RECT  3570.0 38920.0 3635.0 39055.0 ;
      RECT  3760.0 38920.0 3825.0 39055.0 ;
      RECT  3760.0 38920.0 3825.0 39055.0 ;
      RECT  3570.0 38920.0 3635.0 39055.0 ;
      RECT  3930.0 39850.0 3995.0 39985.0 ;
      RECT  3930.0 38875.0 3995.0 39010.0 ;
      RECT  3765.0 39150.0 3630.0 39215.0 ;
      RECT  3507.5 39365.0 3372.5 39430.0 ;
      RECT  3570.0 39760.0 3635.0 39895.0 ;
      RECT  3760.0 38920.0 3825.0 39055.0 ;
      RECT  3860.0 39365.0 3725.0 39430.0 ;
      RECT  3372.5 39365.0 3507.5 39430.0 ;
      RECT  3630.0 39150.0 3765.0 39215.0 ;
      RECT  3725.0 39365.0 3860.0 39430.0 ;
      RECT  3312.5 40070.0 4232.5 40135.0 ;
      RECT  3312.5 38725.0 4232.5 38790.0 ;
      RECT  3380.0 41285.0 3445.0 41480.0 ;
      RECT  3380.0 40445.0 3445.0 40070.0 ;
      RECT  3760.0 40445.0 3825.0 40070.0 ;
      RECT  3930.0 40287.5 3995.0 40102.5 ;
      RECT  3930.0 41447.5 3995.0 41262.5 ;
      RECT  3380.0 40445.0 3445.0 40310.0 ;
      RECT  3570.0 40445.0 3635.0 40310.0 ;
      RECT  3570.0 40445.0 3635.0 40310.0 ;
      RECT  3380.0 40445.0 3445.0 40310.0 ;
      RECT  3570.0 40445.0 3635.0 40310.0 ;
      RECT  3760.0 40445.0 3825.0 40310.0 ;
      RECT  3760.0 40445.0 3825.0 40310.0 ;
      RECT  3570.0 40445.0 3635.0 40310.0 ;
      RECT  3380.0 41285.0 3445.0 41150.0 ;
      RECT  3570.0 41285.0 3635.0 41150.0 ;
      RECT  3570.0 41285.0 3635.0 41150.0 ;
      RECT  3380.0 41285.0 3445.0 41150.0 ;
      RECT  3570.0 41285.0 3635.0 41150.0 ;
      RECT  3760.0 41285.0 3825.0 41150.0 ;
      RECT  3760.0 41285.0 3825.0 41150.0 ;
      RECT  3570.0 41285.0 3635.0 41150.0 ;
      RECT  3930.0 40355.0 3995.0 40220.0 ;
      RECT  3930.0 41330.0 3995.0 41195.0 ;
      RECT  3765.0 41055.0 3630.0 40990.0 ;
      RECT  3507.5 40840.0 3372.5 40775.0 ;
      RECT  3570.0 40445.0 3635.0 40310.0 ;
      RECT  3760.0 41285.0 3825.0 41150.0 ;
      RECT  3860.0 40840.0 3725.0 40775.0 ;
      RECT  3372.5 40840.0 3507.5 40775.0 ;
      RECT  3630.0 41055.0 3765.0 40990.0 ;
      RECT  3725.0 40840.0 3860.0 40775.0 ;
      RECT  3312.5 40135.0 4232.5 40070.0 ;
      RECT  3312.5 41480.0 4232.5 41415.0 ;
      RECT  4660.0 21087.5 4725.0 21272.5 ;
      RECT  4660.0 19927.5 4725.0 20112.5 ;
      RECT  4300.0 20045.0 4365.0 19895.0 ;
      RECT  4300.0 20930.0 4365.0 21305.0 ;
      RECT  4490.0 20045.0 4555.0 20930.0 ;
      RECT  4300.0 20930.0 4365.0 21065.0 ;
      RECT  4490.0 20930.0 4555.0 21065.0 ;
      RECT  4490.0 20930.0 4555.0 21065.0 ;
      RECT  4300.0 20930.0 4365.0 21065.0 ;
      RECT  4300.0 20045.0 4365.0 20180.0 ;
      RECT  4490.0 20045.0 4555.0 20180.0 ;
      RECT  4490.0 20045.0 4555.0 20180.0 ;
      RECT  4300.0 20045.0 4365.0 20180.0 ;
      RECT  4660.0 21020.0 4725.0 21155.0 ;
      RECT  4660.0 20045.0 4725.0 20180.0 ;
      RECT  4357.5 20487.5 4422.5 20622.5 ;
      RECT  4357.5 20487.5 4422.5 20622.5 ;
      RECT  4522.5 20522.5 4587.5 20587.5 ;
      RECT  4232.5 21240.0 4792.5 21305.0 ;
      RECT  4232.5 19895.0 4792.5 19960.0 ;
      RECT  4660.0 21457.5 4725.0 21272.5 ;
      RECT  4660.0 22617.5 4725.0 22432.5 ;
      RECT  4300.0 22500.0 4365.0 22650.0 ;
      RECT  4300.0 21615.0 4365.0 21240.0 ;
      RECT  4490.0 22500.0 4555.0 21615.0 ;
      RECT  4300.0 21615.0 4365.0 21480.0 ;
      RECT  4490.0 21615.0 4555.0 21480.0 ;
      RECT  4490.0 21615.0 4555.0 21480.0 ;
      RECT  4300.0 21615.0 4365.0 21480.0 ;
      RECT  4300.0 22500.0 4365.0 22365.0 ;
      RECT  4490.0 22500.0 4555.0 22365.0 ;
      RECT  4490.0 22500.0 4555.0 22365.0 ;
      RECT  4300.0 22500.0 4365.0 22365.0 ;
      RECT  4660.0 21525.0 4725.0 21390.0 ;
      RECT  4660.0 22500.0 4725.0 22365.0 ;
      RECT  4357.5 22057.5 4422.5 21922.5 ;
      RECT  4357.5 22057.5 4422.5 21922.5 ;
      RECT  4522.5 22022.5 4587.5 21957.5 ;
      RECT  4232.5 21305.0 4792.5 21240.0 ;
      RECT  4232.5 22650.0 4792.5 22585.0 ;
      RECT  4660.0 23777.5 4725.0 23962.5 ;
      RECT  4660.0 22617.5 4725.0 22802.5 ;
      RECT  4300.0 22735.0 4365.0 22585.0 ;
      RECT  4300.0 23620.0 4365.0 23995.0 ;
      RECT  4490.0 22735.0 4555.0 23620.0 ;
      RECT  4300.0 23620.0 4365.0 23755.0 ;
      RECT  4490.0 23620.0 4555.0 23755.0 ;
      RECT  4490.0 23620.0 4555.0 23755.0 ;
      RECT  4300.0 23620.0 4365.0 23755.0 ;
      RECT  4300.0 22735.0 4365.0 22870.0 ;
      RECT  4490.0 22735.0 4555.0 22870.0 ;
      RECT  4490.0 22735.0 4555.0 22870.0 ;
      RECT  4300.0 22735.0 4365.0 22870.0 ;
      RECT  4660.0 23710.0 4725.0 23845.0 ;
      RECT  4660.0 22735.0 4725.0 22870.0 ;
      RECT  4357.5 23177.5 4422.5 23312.5 ;
      RECT  4357.5 23177.5 4422.5 23312.5 ;
      RECT  4522.5 23212.5 4587.5 23277.5 ;
      RECT  4232.5 23930.0 4792.5 23995.0 ;
      RECT  4232.5 22585.0 4792.5 22650.0 ;
      RECT  4660.0 24147.5 4725.0 23962.5 ;
      RECT  4660.0 25307.5 4725.0 25122.5 ;
      RECT  4300.0 25190.0 4365.0 25340.0 ;
      RECT  4300.0 24305.0 4365.0 23930.0 ;
      RECT  4490.0 25190.0 4555.0 24305.0 ;
      RECT  4300.0 24305.0 4365.0 24170.0 ;
      RECT  4490.0 24305.0 4555.0 24170.0 ;
      RECT  4490.0 24305.0 4555.0 24170.0 ;
      RECT  4300.0 24305.0 4365.0 24170.0 ;
      RECT  4300.0 25190.0 4365.0 25055.0 ;
      RECT  4490.0 25190.0 4555.0 25055.0 ;
      RECT  4490.0 25190.0 4555.0 25055.0 ;
      RECT  4300.0 25190.0 4365.0 25055.0 ;
      RECT  4660.0 24215.0 4725.0 24080.0 ;
      RECT  4660.0 25190.0 4725.0 25055.0 ;
      RECT  4357.5 24747.5 4422.5 24612.5 ;
      RECT  4357.5 24747.5 4422.5 24612.5 ;
      RECT  4522.5 24712.5 4587.5 24647.5 ;
      RECT  4232.5 23995.0 4792.5 23930.0 ;
      RECT  4232.5 25340.0 4792.5 25275.0 ;
      RECT  4660.0 26467.5 4725.0 26652.5 ;
      RECT  4660.0 25307.5 4725.0 25492.5 ;
      RECT  4300.0 25425.0 4365.0 25275.0 ;
      RECT  4300.0 26310.0 4365.0 26685.0 ;
      RECT  4490.0 25425.0 4555.0 26310.0 ;
      RECT  4300.0 26310.0 4365.0 26445.0 ;
      RECT  4490.0 26310.0 4555.0 26445.0 ;
      RECT  4490.0 26310.0 4555.0 26445.0 ;
      RECT  4300.0 26310.0 4365.0 26445.0 ;
      RECT  4300.0 25425.0 4365.0 25560.0 ;
      RECT  4490.0 25425.0 4555.0 25560.0 ;
      RECT  4490.0 25425.0 4555.0 25560.0 ;
      RECT  4300.0 25425.0 4365.0 25560.0 ;
      RECT  4660.0 26400.0 4725.0 26535.0 ;
      RECT  4660.0 25425.0 4725.0 25560.0 ;
      RECT  4357.5 25867.5 4422.5 26002.5 ;
      RECT  4357.5 25867.5 4422.5 26002.5 ;
      RECT  4522.5 25902.5 4587.5 25967.5 ;
      RECT  4232.5 26620.0 4792.5 26685.0 ;
      RECT  4232.5 25275.0 4792.5 25340.0 ;
      RECT  4660.0 26837.5 4725.0 26652.5 ;
      RECT  4660.0 27997.5 4725.0 27812.5 ;
      RECT  4300.0 27880.0 4365.0 28030.0 ;
      RECT  4300.0 26995.0 4365.0 26620.0 ;
      RECT  4490.0 27880.0 4555.0 26995.0 ;
      RECT  4300.0 26995.0 4365.0 26860.0 ;
      RECT  4490.0 26995.0 4555.0 26860.0 ;
      RECT  4490.0 26995.0 4555.0 26860.0 ;
      RECT  4300.0 26995.0 4365.0 26860.0 ;
      RECT  4300.0 27880.0 4365.0 27745.0 ;
      RECT  4490.0 27880.0 4555.0 27745.0 ;
      RECT  4490.0 27880.0 4555.0 27745.0 ;
      RECT  4300.0 27880.0 4365.0 27745.0 ;
      RECT  4660.0 26905.0 4725.0 26770.0 ;
      RECT  4660.0 27880.0 4725.0 27745.0 ;
      RECT  4357.5 27437.5 4422.5 27302.5 ;
      RECT  4357.5 27437.5 4422.5 27302.5 ;
      RECT  4522.5 27402.5 4587.5 27337.5 ;
      RECT  4232.5 26685.0 4792.5 26620.0 ;
      RECT  4232.5 28030.0 4792.5 27965.0 ;
      RECT  4660.0 29157.5 4725.0 29342.5 ;
      RECT  4660.0 27997.5 4725.0 28182.5 ;
      RECT  4300.0 28115.0 4365.0 27965.0 ;
      RECT  4300.0 29000.0 4365.0 29375.0 ;
      RECT  4490.0 28115.0 4555.0 29000.0 ;
      RECT  4300.0 29000.0 4365.0 29135.0 ;
      RECT  4490.0 29000.0 4555.0 29135.0 ;
      RECT  4490.0 29000.0 4555.0 29135.0 ;
      RECT  4300.0 29000.0 4365.0 29135.0 ;
      RECT  4300.0 28115.0 4365.0 28250.0 ;
      RECT  4490.0 28115.0 4555.0 28250.0 ;
      RECT  4490.0 28115.0 4555.0 28250.0 ;
      RECT  4300.0 28115.0 4365.0 28250.0 ;
      RECT  4660.0 29090.0 4725.0 29225.0 ;
      RECT  4660.0 28115.0 4725.0 28250.0 ;
      RECT  4357.5 28557.5 4422.5 28692.5 ;
      RECT  4357.5 28557.5 4422.5 28692.5 ;
      RECT  4522.5 28592.5 4587.5 28657.5 ;
      RECT  4232.5 29310.0 4792.5 29375.0 ;
      RECT  4232.5 27965.0 4792.5 28030.0 ;
      RECT  4660.0 29527.5 4725.0 29342.5 ;
      RECT  4660.0 30687.5 4725.0 30502.5 ;
      RECT  4300.0 30570.0 4365.0 30720.0 ;
      RECT  4300.0 29685.0 4365.0 29310.0 ;
      RECT  4490.0 30570.0 4555.0 29685.0 ;
      RECT  4300.0 29685.0 4365.0 29550.0 ;
      RECT  4490.0 29685.0 4555.0 29550.0 ;
      RECT  4490.0 29685.0 4555.0 29550.0 ;
      RECT  4300.0 29685.0 4365.0 29550.0 ;
      RECT  4300.0 30570.0 4365.0 30435.0 ;
      RECT  4490.0 30570.0 4555.0 30435.0 ;
      RECT  4490.0 30570.0 4555.0 30435.0 ;
      RECT  4300.0 30570.0 4365.0 30435.0 ;
      RECT  4660.0 29595.0 4725.0 29460.0 ;
      RECT  4660.0 30570.0 4725.0 30435.0 ;
      RECT  4357.5 30127.5 4422.5 29992.5 ;
      RECT  4357.5 30127.5 4422.5 29992.5 ;
      RECT  4522.5 30092.5 4587.5 30027.5 ;
      RECT  4232.5 29375.0 4792.5 29310.0 ;
      RECT  4232.5 30720.0 4792.5 30655.0 ;
      RECT  4660.0 31847.5 4725.0 32032.5 ;
      RECT  4660.0 30687.5 4725.0 30872.5 ;
      RECT  4300.0 30805.0 4365.0 30655.0 ;
      RECT  4300.0 31690.0 4365.0 32065.0 ;
      RECT  4490.0 30805.0 4555.0 31690.0 ;
      RECT  4300.0 31690.0 4365.0 31825.0 ;
      RECT  4490.0 31690.0 4555.0 31825.0 ;
      RECT  4490.0 31690.0 4555.0 31825.0 ;
      RECT  4300.0 31690.0 4365.0 31825.0 ;
      RECT  4300.0 30805.0 4365.0 30940.0 ;
      RECT  4490.0 30805.0 4555.0 30940.0 ;
      RECT  4490.0 30805.0 4555.0 30940.0 ;
      RECT  4300.0 30805.0 4365.0 30940.0 ;
      RECT  4660.0 31780.0 4725.0 31915.0 ;
      RECT  4660.0 30805.0 4725.0 30940.0 ;
      RECT  4357.5 31247.5 4422.5 31382.5 ;
      RECT  4357.5 31247.5 4422.5 31382.5 ;
      RECT  4522.5 31282.5 4587.5 31347.5 ;
      RECT  4232.5 32000.0 4792.5 32065.0 ;
      RECT  4232.5 30655.0 4792.5 30720.0 ;
      RECT  4660.0 32217.5 4725.0 32032.5 ;
      RECT  4660.0 33377.5 4725.0 33192.5 ;
      RECT  4300.0 33260.0 4365.0 33410.0 ;
      RECT  4300.0 32375.0 4365.0 32000.0 ;
      RECT  4490.0 33260.0 4555.0 32375.0 ;
      RECT  4300.0 32375.0 4365.0 32240.0 ;
      RECT  4490.0 32375.0 4555.0 32240.0 ;
      RECT  4490.0 32375.0 4555.0 32240.0 ;
      RECT  4300.0 32375.0 4365.0 32240.0 ;
      RECT  4300.0 33260.0 4365.0 33125.0 ;
      RECT  4490.0 33260.0 4555.0 33125.0 ;
      RECT  4490.0 33260.0 4555.0 33125.0 ;
      RECT  4300.0 33260.0 4365.0 33125.0 ;
      RECT  4660.0 32285.0 4725.0 32150.0 ;
      RECT  4660.0 33260.0 4725.0 33125.0 ;
      RECT  4357.5 32817.5 4422.5 32682.5 ;
      RECT  4357.5 32817.5 4422.5 32682.5 ;
      RECT  4522.5 32782.5 4587.5 32717.5 ;
      RECT  4232.5 32065.0 4792.5 32000.0 ;
      RECT  4232.5 33410.0 4792.5 33345.0 ;
      RECT  4660.0 34537.5 4725.0 34722.5 ;
      RECT  4660.0 33377.5 4725.0 33562.5 ;
      RECT  4300.0 33495.0 4365.0 33345.0 ;
      RECT  4300.0 34380.0 4365.0 34755.0 ;
      RECT  4490.0 33495.0 4555.0 34380.0 ;
      RECT  4300.0 34380.0 4365.0 34515.0 ;
      RECT  4490.0 34380.0 4555.0 34515.0 ;
      RECT  4490.0 34380.0 4555.0 34515.0 ;
      RECT  4300.0 34380.0 4365.0 34515.0 ;
      RECT  4300.0 33495.0 4365.0 33630.0 ;
      RECT  4490.0 33495.0 4555.0 33630.0 ;
      RECT  4490.0 33495.0 4555.0 33630.0 ;
      RECT  4300.0 33495.0 4365.0 33630.0 ;
      RECT  4660.0 34470.0 4725.0 34605.0 ;
      RECT  4660.0 33495.0 4725.0 33630.0 ;
      RECT  4357.5 33937.5 4422.5 34072.5 ;
      RECT  4357.5 33937.5 4422.5 34072.5 ;
      RECT  4522.5 33972.5 4587.5 34037.5 ;
      RECT  4232.5 34690.0 4792.5 34755.0 ;
      RECT  4232.5 33345.0 4792.5 33410.0 ;
      RECT  4660.0 34907.5 4725.0 34722.5 ;
      RECT  4660.0 36067.5 4725.0 35882.5 ;
      RECT  4300.0 35950.0 4365.0 36100.0 ;
      RECT  4300.0 35065.0 4365.0 34690.0 ;
      RECT  4490.0 35950.0 4555.0 35065.0 ;
      RECT  4300.0 35065.0 4365.0 34930.0 ;
      RECT  4490.0 35065.0 4555.0 34930.0 ;
      RECT  4490.0 35065.0 4555.0 34930.0 ;
      RECT  4300.0 35065.0 4365.0 34930.0 ;
      RECT  4300.0 35950.0 4365.0 35815.0 ;
      RECT  4490.0 35950.0 4555.0 35815.0 ;
      RECT  4490.0 35950.0 4555.0 35815.0 ;
      RECT  4300.0 35950.0 4365.0 35815.0 ;
      RECT  4660.0 34975.0 4725.0 34840.0 ;
      RECT  4660.0 35950.0 4725.0 35815.0 ;
      RECT  4357.5 35507.5 4422.5 35372.5 ;
      RECT  4357.5 35507.5 4422.5 35372.5 ;
      RECT  4522.5 35472.5 4587.5 35407.5 ;
      RECT  4232.5 34755.0 4792.5 34690.0 ;
      RECT  4232.5 36100.0 4792.5 36035.0 ;
      RECT  4660.0 37227.5 4725.0 37412.5 ;
      RECT  4660.0 36067.5 4725.0 36252.5 ;
      RECT  4300.0 36185.0 4365.0 36035.0 ;
      RECT  4300.0 37070.0 4365.0 37445.0 ;
      RECT  4490.0 36185.0 4555.0 37070.0 ;
      RECT  4300.0 37070.0 4365.0 37205.0 ;
      RECT  4490.0 37070.0 4555.0 37205.0 ;
      RECT  4490.0 37070.0 4555.0 37205.0 ;
      RECT  4300.0 37070.0 4365.0 37205.0 ;
      RECT  4300.0 36185.0 4365.0 36320.0 ;
      RECT  4490.0 36185.0 4555.0 36320.0 ;
      RECT  4490.0 36185.0 4555.0 36320.0 ;
      RECT  4300.0 36185.0 4365.0 36320.0 ;
      RECT  4660.0 37160.0 4725.0 37295.0 ;
      RECT  4660.0 36185.0 4725.0 36320.0 ;
      RECT  4357.5 36627.5 4422.5 36762.5 ;
      RECT  4357.5 36627.5 4422.5 36762.5 ;
      RECT  4522.5 36662.5 4587.5 36727.5 ;
      RECT  4232.5 37380.0 4792.5 37445.0 ;
      RECT  4232.5 36035.0 4792.5 36100.0 ;
      RECT  4660.0 37597.5 4725.0 37412.5 ;
      RECT  4660.0 38757.5 4725.0 38572.5 ;
      RECT  4300.0 38640.0 4365.0 38790.0 ;
      RECT  4300.0 37755.0 4365.0 37380.0 ;
      RECT  4490.0 38640.0 4555.0 37755.0 ;
      RECT  4300.0 37755.0 4365.0 37620.0 ;
      RECT  4490.0 37755.0 4555.0 37620.0 ;
      RECT  4490.0 37755.0 4555.0 37620.0 ;
      RECT  4300.0 37755.0 4365.0 37620.0 ;
      RECT  4300.0 38640.0 4365.0 38505.0 ;
      RECT  4490.0 38640.0 4555.0 38505.0 ;
      RECT  4490.0 38640.0 4555.0 38505.0 ;
      RECT  4300.0 38640.0 4365.0 38505.0 ;
      RECT  4660.0 37665.0 4725.0 37530.0 ;
      RECT  4660.0 38640.0 4725.0 38505.0 ;
      RECT  4357.5 38197.5 4422.5 38062.5 ;
      RECT  4357.5 38197.5 4422.5 38062.5 ;
      RECT  4522.5 38162.5 4587.5 38097.5 ;
      RECT  4232.5 37445.0 4792.5 37380.0 ;
      RECT  4232.5 38790.0 4792.5 38725.0 ;
      RECT  4660.0 39917.5 4725.0 40102.5 ;
      RECT  4660.0 38757.5 4725.0 38942.5 ;
      RECT  4300.0 38875.0 4365.0 38725.0 ;
      RECT  4300.0 39760.0 4365.0 40135.0 ;
      RECT  4490.0 38875.0 4555.0 39760.0 ;
      RECT  4300.0 39760.0 4365.0 39895.0 ;
      RECT  4490.0 39760.0 4555.0 39895.0 ;
      RECT  4490.0 39760.0 4555.0 39895.0 ;
      RECT  4300.0 39760.0 4365.0 39895.0 ;
      RECT  4300.0 38875.0 4365.0 39010.0 ;
      RECT  4490.0 38875.0 4555.0 39010.0 ;
      RECT  4490.0 38875.0 4555.0 39010.0 ;
      RECT  4300.0 38875.0 4365.0 39010.0 ;
      RECT  4660.0 39850.0 4725.0 39985.0 ;
      RECT  4660.0 38875.0 4725.0 39010.0 ;
      RECT  4357.5 39317.5 4422.5 39452.5 ;
      RECT  4357.5 39317.5 4422.5 39452.5 ;
      RECT  4522.5 39352.5 4587.5 39417.5 ;
      RECT  4232.5 40070.0 4792.5 40135.0 ;
      RECT  4232.5 38725.0 4792.5 38790.0 ;
      RECT  4660.0 40287.5 4725.0 40102.5 ;
      RECT  4660.0 41447.5 4725.0 41262.5 ;
      RECT  4300.0 41330.0 4365.0 41480.0 ;
      RECT  4300.0 40445.0 4365.0 40070.0 ;
      RECT  4490.0 41330.0 4555.0 40445.0 ;
      RECT  4300.0 40445.0 4365.0 40310.0 ;
      RECT  4490.0 40445.0 4555.0 40310.0 ;
      RECT  4490.0 40445.0 4555.0 40310.0 ;
      RECT  4300.0 40445.0 4365.0 40310.0 ;
      RECT  4300.0 41330.0 4365.0 41195.0 ;
      RECT  4490.0 41330.0 4555.0 41195.0 ;
      RECT  4490.0 41330.0 4555.0 41195.0 ;
      RECT  4300.0 41330.0 4365.0 41195.0 ;
      RECT  4660.0 40355.0 4725.0 40220.0 ;
      RECT  4660.0 41330.0 4725.0 41195.0 ;
      RECT  4357.5 40887.5 4422.5 40752.5 ;
      RECT  4357.5 40887.5 4422.5 40752.5 ;
      RECT  4522.5 40852.5 4587.5 40787.5 ;
      RECT  4232.5 40135.0 4792.5 40070.0 ;
      RECT  4232.5 41480.0 4792.5 41415.0 ;
      RECT  2015.0 9762.5 1880.0 9827.5 ;
      RECT  2190.0 11197.5 2055.0 11262.5 ;
      RECT  2365.0 12452.5 2230.0 12517.5 ;
      RECT  2540.0 13887.5 2405.0 13952.5 ;
      RECT  2715.0 15142.5 2580.0 15207.5 ;
      RECT  2890.0 16577.5 2755.0 16642.5 ;
      RECT  3065.0 17832.5 2930.0 17897.5 ;
      RECT  3240.0 19267.5 3105.0 19332.5 ;
      RECT  2015.0 20535.0 1880.0 20600.0 ;
      RECT  2715.0 20320.0 2580.0 20385.0 ;
      RECT  2015.0 21945.0 1880.0 22010.0 ;
      RECT  2890.0 22160.0 2755.0 22225.0 ;
      RECT  2015.0 23225.0 1880.0 23290.0 ;
      RECT  3065.0 23010.0 2930.0 23075.0 ;
      RECT  2015.0 24635.0 1880.0 24700.0 ;
      RECT  3240.0 24850.0 3105.0 24915.0 ;
      RECT  2190.0 25915.0 2055.0 25980.0 ;
      RECT  2715.0 25700.0 2580.0 25765.0 ;
      RECT  2190.0 27325.0 2055.0 27390.0 ;
      RECT  2890.0 27540.0 2755.0 27605.0 ;
      RECT  2190.0 28605.0 2055.0 28670.0 ;
      RECT  3065.0 28390.0 2930.0 28455.0 ;
      RECT  2190.0 30015.0 2055.0 30080.0 ;
      RECT  3240.0 30230.0 3105.0 30295.0 ;
      RECT  2365.0 31295.0 2230.0 31360.0 ;
      RECT  2715.0 31080.0 2580.0 31145.0 ;
      RECT  2365.0 32705.0 2230.0 32770.0 ;
      RECT  2890.0 32920.0 2755.0 32985.0 ;
      RECT  2365.0 33985.0 2230.0 34050.0 ;
      RECT  3065.0 33770.0 2930.0 33835.0 ;
      RECT  2365.0 35395.0 2230.0 35460.0 ;
      RECT  3240.0 35610.0 3105.0 35675.0 ;
      RECT  2540.0 36675.0 2405.0 36740.0 ;
      RECT  2715.0 36460.0 2580.0 36525.0 ;
      RECT  2540.0 38085.0 2405.0 38150.0 ;
      RECT  2890.0 38300.0 2755.0 38365.0 ;
      RECT  2540.0 39365.0 2405.0 39430.0 ;
      RECT  3065.0 39150.0 2930.0 39215.0 ;
      RECT  2540.0 40775.0 2405.0 40840.0 ;
      RECT  3240.0 40990.0 3105.0 41055.0 ;
      RECT  4522.5 20522.5 4587.5 20587.5 ;
      RECT  4522.5 21957.5 4587.5 22022.5 ;
      RECT  4522.5 23212.5 4587.5 23277.5 ;
      RECT  4522.5 24647.5 4587.5 24712.5 ;
      RECT  4522.5 25902.5 4587.5 25967.5 ;
      RECT  4522.5 27337.5 4587.5 27402.5 ;
      RECT  4522.5 28592.5 4587.5 28657.5 ;
      RECT  4522.5 30027.5 4587.5 30092.5 ;
      RECT  4522.5 31282.5 4587.5 31347.5 ;
      RECT  4522.5 32717.5 4587.5 32782.5 ;
      RECT  4522.5 33972.5 4587.5 34037.5 ;
      RECT  4522.5 35407.5 4587.5 35472.5 ;
      RECT  4522.5 36662.5 4587.5 36727.5 ;
      RECT  4522.5 38097.5 4587.5 38162.5 ;
      RECT  4522.5 39352.5 4587.5 39417.5 ;
      RECT  4522.5 40787.5 4587.5 40852.5 ;
      RECT  1912.5 10480.0 7277.5 10545.0 ;
      RECT  1912.5 13170.0 7277.5 13235.0 ;
      RECT  1912.5 15860.0 7277.5 15925.0 ;
      RECT  1912.5 18550.0 7277.5 18615.0 ;
      RECT  1912.5 21240.0 7277.5 21305.0 ;
      RECT  1912.5 23930.0 7277.5 23995.0 ;
      RECT  1912.5 26620.0 7277.5 26685.0 ;
      RECT  1912.5 29310.0 7277.5 29375.0 ;
      RECT  1912.5 32000.0 7277.5 32065.0 ;
      RECT  1912.5 34690.0 7277.5 34755.0 ;
      RECT  1912.5 37380.0 7277.5 37445.0 ;
      RECT  1912.5 40070.0 7277.5 40135.0 ;
      RECT  1912.5 9135.0 7277.5 9200.0 ;
      RECT  1912.5 11825.0 7277.5 11890.0 ;
      RECT  1912.5 14515.0 7277.5 14580.0 ;
      RECT  1912.5 17205.0 7277.5 17270.0 ;
      RECT  1912.5 19895.0 7277.5 19960.0 ;
      RECT  1912.5 22585.0 7277.5 22650.0 ;
      RECT  1912.5 25275.0 7277.5 25340.0 ;
      RECT  1912.5 27965.0 7277.5 28030.0 ;
      RECT  1912.5 30655.0 7277.5 30720.0 ;
      RECT  1912.5 33345.0 7277.5 33410.0 ;
      RECT  1912.5 36035.0 7277.5 36100.0 ;
      RECT  1912.5 38725.0 7277.5 38790.0 ;
      RECT  1912.5 41415.0 7277.5 41480.0 ;
      RECT  5022.5 20522.5 5372.5 20587.5 ;
      RECT  5537.5 20535.0 5602.5 20600.0 ;
      RECT  5537.5 20522.5 5602.5 20587.5 ;
      RECT  5537.5 20567.5 5602.5 20587.5 ;
      RECT  5570.0 20535.0 5867.5 20600.0 ;
      RECT  5867.5 20535.0 6002.5 20600.0 ;
      RECT  6572.5 20535.0 6637.5 20600.0 ;
      RECT  6572.5 20522.5 6637.5 20587.5 ;
      RECT  6355.0 20535.0 6605.0 20600.0 ;
      RECT  6572.5 20555.0 6637.5 20567.5 ;
      RECT  6605.0 20522.5 6852.5 20587.5 ;
      RECT  5022.5 21957.5 5372.5 22022.5 ;
      RECT  5537.5 21945.0 5602.5 22010.0 ;
      RECT  5537.5 21957.5 5602.5 22022.5 ;
      RECT  5537.5 21977.5 5602.5 22022.5 ;
      RECT  5570.0 21945.0 5867.5 22010.0 ;
      RECT  5867.5 21945.0 6002.5 22010.0 ;
      RECT  6572.5 21945.0 6637.5 22010.0 ;
      RECT  6572.5 21957.5 6637.5 22022.5 ;
      RECT  6355.0 21945.0 6605.0 22010.0 ;
      RECT  6572.5 21977.5 6637.5 21990.0 ;
      RECT  6605.0 21957.5 6852.5 22022.5 ;
      RECT  5022.5 23212.5 5372.5 23277.5 ;
      RECT  5537.5 23225.0 5602.5 23290.0 ;
      RECT  5537.5 23212.5 5602.5 23277.5 ;
      RECT  5537.5 23257.5 5602.5 23277.5 ;
      RECT  5570.0 23225.0 5867.5 23290.0 ;
      RECT  5867.5 23225.0 6002.5 23290.0 ;
      RECT  6572.5 23225.0 6637.5 23290.0 ;
      RECT  6572.5 23212.5 6637.5 23277.5 ;
      RECT  6355.0 23225.0 6605.0 23290.0 ;
      RECT  6572.5 23245.0 6637.5 23257.5 ;
      RECT  6605.0 23212.5 6852.5 23277.5 ;
      RECT  5022.5 24647.5 5372.5 24712.5 ;
      RECT  5537.5 24635.0 5602.5 24700.0 ;
      RECT  5537.5 24647.5 5602.5 24712.5 ;
      RECT  5537.5 24667.5 5602.5 24712.5 ;
      RECT  5570.0 24635.0 5867.5 24700.0 ;
      RECT  5867.5 24635.0 6002.5 24700.0 ;
      RECT  6572.5 24635.0 6637.5 24700.0 ;
      RECT  6572.5 24647.5 6637.5 24712.5 ;
      RECT  6355.0 24635.0 6605.0 24700.0 ;
      RECT  6572.5 24667.5 6637.5 24680.0 ;
      RECT  6605.0 24647.5 6852.5 24712.5 ;
      RECT  5022.5 25902.5 5372.5 25967.5 ;
      RECT  5537.5 25915.0 5602.5 25980.0 ;
      RECT  5537.5 25902.5 5602.5 25967.5 ;
      RECT  5537.5 25947.5 5602.5 25967.5 ;
      RECT  5570.0 25915.0 5867.5 25980.0 ;
      RECT  5867.5 25915.0 6002.5 25980.0 ;
      RECT  6572.5 25915.0 6637.5 25980.0 ;
      RECT  6572.5 25902.5 6637.5 25967.5 ;
      RECT  6355.0 25915.0 6605.0 25980.0 ;
      RECT  6572.5 25935.0 6637.5 25947.5 ;
      RECT  6605.0 25902.5 6852.5 25967.5 ;
      RECT  5022.5 27337.5 5372.5 27402.5 ;
      RECT  5537.5 27325.0 5602.5 27390.0 ;
      RECT  5537.5 27337.5 5602.5 27402.5 ;
      RECT  5537.5 27357.5 5602.5 27402.5 ;
      RECT  5570.0 27325.0 5867.5 27390.0 ;
      RECT  5867.5 27325.0 6002.5 27390.0 ;
      RECT  6572.5 27325.0 6637.5 27390.0 ;
      RECT  6572.5 27337.5 6637.5 27402.5 ;
      RECT  6355.0 27325.0 6605.0 27390.0 ;
      RECT  6572.5 27357.5 6637.5 27370.0 ;
      RECT  6605.0 27337.5 6852.5 27402.5 ;
      RECT  5022.5 28592.5 5372.5 28657.5 ;
      RECT  5537.5 28605.0 5602.5 28670.0 ;
      RECT  5537.5 28592.5 5602.5 28657.5 ;
      RECT  5537.5 28637.5 5602.5 28657.5 ;
      RECT  5570.0 28605.0 5867.5 28670.0 ;
      RECT  5867.5 28605.0 6002.5 28670.0 ;
      RECT  6572.5 28605.0 6637.5 28670.0 ;
      RECT  6572.5 28592.5 6637.5 28657.5 ;
      RECT  6355.0 28605.0 6605.0 28670.0 ;
      RECT  6572.5 28625.0 6637.5 28637.5 ;
      RECT  6605.0 28592.5 6852.5 28657.5 ;
      RECT  5022.5 30027.5 5372.5 30092.5 ;
      RECT  5537.5 30015.0 5602.5 30080.0 ;
      RECT  5537.5 30027.5 5602.5 30092.5 ;
      RECT  5537.5 30047.5 5602.5 30092.5 ;
      RECT  5570.0 30015.0 5867.5 30080.0 ;
      RECT  5867.5 30015.0 6002.5 30080.0 ;
      RECT  6572.5 30015.0 6637.5 30080.0 ;
      RECT  6572.5 30027.5 6637.5 30092.5 ;
      RECT  6355.0 30015.0 6605.0 30080.0 ;
      RECT  6572.5 30047.5 6637.5 30060.0 ;
      RECT  6605.0 30027.5 6852.5 30092.5 ;
      RECT  5022.5 31282.5 5372.5 31347.5 ;
      RECT  5537.5 31295.0 5602.5 31360.0 ;
      RECT  5537.5 31282.5 5602.5 31347.5 ;
      RECT  5537.5 31327.5 5602.5 31347.5 ;
      RECT  5570.0 31295.0 5867.5 31360.0 ;
      RECT  5867.5 31295.0 6002.5 31360.0 ;
      RECT  6572.5 31295.0 6637.5 31360.0 ;
      RECT  6572.5 31282.5 6637.5 31347.5 ;
      RECT  6355.0 31295.0 6605.0 31360.0 ;
      RECT  6572.5 31315.0 6637.5 31327.5 ;
      RECT  6605.0 31282.5 6852.5 31347.5 ;
      RECT  5022.5 32717.5 5372.5 32782.5 ;
      RECT  5537.5 32705.0 5602.5 32770.0 ;
      RECT  5537.5 32717.5 5602.5 32782.5 ;
      RECT  5537.5 32737.5 5602.5 32782.5 ;
      RECT  5570.0 32705.0 5867.5 32770.0 ;
      RECT  5867.5 32705.0 6002.5 32770.0 ;
      RECT  6572.5 32705.0 6637.5 32770.0 ;
      RECT  6572.5 32717.5 6637.5 32782.5 ;
      RECT  6355.0 32705.0 6605.0 32770.0 ;
      RECT  6572.5 32737.5 6637.5 32750.0 ;
      RECT  6605.0 32717.5 6852.5 32782.5 ;
      RECT  5022.5 33972.5 5372.5 34037.5 ;
      RECT  5537.5 33985.0 5602.5 34050.0 ;
      RECT  5537.5 33972.5 5602.5 34037.5 ;
      RECT  5537.5 34017.5 5602.5 34037.5 ;
      RECT  5570.0 33985.0 5867.5 34050.0 ;
      RECT  5867.5 33985.0 6002.5 34050.0 ;
      RECT  6572.5 33985.0 6637.5 34050.0 ;
      RECT  6572.5 33972.5 6637.5 34037.5 ;
      RECT  6355.0 33985.0 6605.0 34050.0 ;
      RECT  6572.5 34005.0 6637.5 34017.5 ;
      RECT  6605.0 33972.5 6852.5 34037.5 ;
      RECT  5022.5 35407.5 5372.5 35472.5 ;
      RECT  5537.5 35395.0 5602.5 35460.0 ;
      RECT  5537.5 35407.5 5602.5 35472.5 ;
      RECT  5537.5 35427.5 5602.5 35472.5 ;
      RECT  5570.0 35395.0 5867.5 35460.0 ;
      RECT  5867.5 35395.0 6002.5 35460.0 ;
      RECT  6572.5 35395.0 6637.5 35460.0 ;
      RECT  6572.5 35407.5 6637.5 35472.5 ;
      RECT  6355.0 35395.0 6605.0 35460.0 ;
      RECT  6572.5 35427.5 6637.5 35440.0 ;
      RECT  6605.0 35407.5 6852.5 35472.5 ;
      RECT  5022.5 36662.5 5372.5 36727.5 ;
      RECT  5537.5 36675.0 5602.5 36740.0 ;
      RECT  5537.5 36662.5 5602.5 36727.5 ;
      RECT  5537.5 36707.5 5602.5 36727.5 ;
      RECT  5570.0 36675.0 5867.5 36740.0 ;
      RECT  5867.5 36675.0 6002.5 36740.0 ;
      RECT  6572.5 36675.0 6637.5 36740.0 ;
      RECT  6572.5 36662.5 6637.5 36727.5 ;
      RECT  6355.0 36675.0 6605.0 36740.0 ;
      RECT  6572.5 36695.0 6637.5 36707.5 ;
      RECT  6605.0 36662.5 6852.5 36727.5 ;
      RECT  5022.5 38097.5 5372.5 38162.5 ;
      RECT  5537.5 38085.0 5602.5 38150.0 ;
      RECT  5537.5 38097.5 5602.5 38162.5 ;
      RECT  5537.5 38117.5 5602.5 38162.5 ;
      RECT  5570.0 38085.0 5867.5 38150.0 ;
      RECT  5867.5 38085.0 6002.5 38150.0 ;
      RECT  6572.5 38085.0 6637.5 38150.0 ;
      RECT  6572.5 38097.5 6637.5 38162.5 ;
      RECT  6355.0 38085.0 6605.0 38150.0 ;
      RECT  6572.5 38117.5 6637.5 38130.0 ;
      RECT  6605.0 38097.5 6852.5 38162.5 ;
      RECT  5022.5 39352.5 5372.5 39417.5 ;
      RECT  5537.5 39365.0 5602.5 39430.0 ;
      RECT  5537.5 39352.5 5602.5 39417.5 ;
      RECT  5537.5 39397.5 5602.5 39417.5 ;
      RECT  5570.0 39365.0 5867.5 39430.0 ;
      RECT  5867.5 39365.0 6002.5 39430.0 ;
      RECT  6572.5 39365.0 6637.5 39430.0 ;
      RECT  6572.5 39352.5 6637.5 39417.5 ;
      RECT  6355.0 39365.0 6605.0 39430.0 ;
      RECT  6572.5 39385.0 6637.5 39397.5 ;
      RECT  6605.0 39352.5 6852.5 39417.5 ;
      RECT  5022.5 40787.5 5372.5 40852.5 ;
      RECT  5537.5 40775.0 5602.5 40840.0 ;
      RECT  5537.5 40787.5 5602.5 40852.5 ;
      RECT  5537.5 40807.5 5602.5 40852.5 ;
      RECT  5570.0 40775.0 5867.5 40840.0 ;
      RECT  5867.5 40775.0 6002.5 40840.0 ;
      RECT  6572.5 40775.0 6637.5 40840.0 ;
      RECT  6572.5 40787.5 6637.5 40852.5 ;
      RECT  6355.0 40775.0 6605.0 40840.0 ;
      RECT  6572.5 40807.5 6637.5 40820.0 ;
      RECT  6605.0 40787.5 6852.5 40852.5 ;
      RECT  5675.0 21087.5 5740.0 21272.5 ;
      RECT  5675.0 19927.5 5740.0 20112.5 ;
      RECT  5315.0 20045.0 5380.0 19895.0 ;
      RECT  5315.0 20930.0 5380.0 21305.0 ;
      RECT  5505.0 20045.0 5570.0 20930.0 ;
      RECT  5315.0 20930.0 5380.0 21065.0 ;
      RECT  5505.0 20930.0 5570.0 21065.0 ;
      RECT  5505.0 20930.0 5570.0 21065.0 ;
      RECT  5315.0 20930.0 5380.0 21065.0 ;
      RECT  5315.0 20045.0 5380.0 20180.0 ;
      RECT  5505.0 20045.0 5570.0 20180.0 ;
      RECT  5505.0 20045.0 5570.0 20180.0 ;
      RECT  5315.0 20045.0 5380.0 20180.0 ;
      RECT  5675.0 21020.0 5740.0 21155.0 ;
      RECT  5675.0 20045.0 5740.0 20180.0 ;
      RECT  5372.5 20487.5 5437.5 20622.5 ;
      RECT  5372.5 20487.5 5437.5 20622.5 ;
      RECT  5537.5 20522.5 5602.5 20587.5 ;
      RECT  5247.5 21240.0 5807.5 21305.0 ;
      RECT  5247.5 19895.0 5807.5 19960.0 ;
      RECT  5875.0 20090.0 5940.0 19895.0 ;
      RECT  5875.0 20930.0 5940.0 21305.0 ;
      RECT  6255.0 20930.0 6320.0 21305.0 ;
      RECT  6425.0 21087.5 6490.0 21272.5 ;
      RECT  6425.0 19927.5 6490.0 20112.5 ;
      RECT  5875.0 20930.0 5940.0 21065.0 ;
      RECT  6065.0 20930.0 6130.0 21065.0 ;
      RECT  6065.0 20930.0 6130.0 21065.0 ;
      RECT  5875.0 20930.0 5940.0 21065.0 ;
      RECT  6065.0 20930.0 6130.0 21065.0 ;
      RECT  6255.0 20930.0 6320.0 21065.0 ;
      RECT  6255.0 20930.0 6320.0 21065.0 ;
      RECT  6065.0 20930.0 6130.0 21065.0 ;
      RECT  5875.0 20090.0 5940.0 20225.0 ;
      RECT  6065.0 20090.0 6130.0 20225.0 ;
      RECT  6065.0 20090.0 6130.0 20225.0 ;
      RECT  5875.0 20090.0 5940.0 20225.0 ;
      RECT  6065.0 20090.0 6130.0 20225.0 ;
      RECT  6255.0 20090.0 6320.0 20225.0 ;
      RECT  6255.0 20090.0 6320.0 20225.0 ;
      RECT  6065.0 20090.0 6130.0 20225.0 ;
      RECT  6425.0 21020.0 6490.0 21155.0 ;
      RECT  6425.0 20045.0 6490.0 20180.0 ;
      RECT  6260.0 20320.0 6125.0 20385.0 ;
      RECT  6002.5 20535.0 5867.5 20600.0 ;
      RECT  6065.0 20930.0 6130.0 21065.0 ;
      RECT  6255.0 20090.0 6320.0 20225.0 ;
      RECT  6355.0 20535.0 6220.0 20600.0 ;
      RECT  5867.5 20535.0 6002.5 20600.0 ;
      RECT  6125.0 20320.0 6260.0 20385.0 ;
      RECT  6220.0 20535.0 6355.0 20600.0 ;
      RECT  5807.5 21240.0 6727.5 21305.0 ;
      RECT  5807.5 19895.0 6727.5 19960.0 ;
      RECT  7155.0 21087.5 7220.0 21272.5 ;
      RECT  7155.0 19927.5 7220.0 20112.5 ;
      RECT  6795.0 20045.0 6860.0 19895.0 ;
      RECT  6795.0 20930.0 6860.0 21305.0 ;
      RECT  6985.0 20045.0 7050.0 20930.0 ;
      RECT  6795.0 20930.0 6860.0 21065.0 ;
      RECT  6985.0 20930.0 7050.0 21065.0 ;
      RECT  6985.0 20930.0 7050.0 21065.0 ;
      RECT  6795.0 20930.0 6860.0 21065.0 ;
      RECT  6795.0 20045.0 6860.0 20180.0 ;
      RECT  6985.0 20045.0 7050.0 20180.0 ;
      RECT  6985.0 20045.0 7050.0 20180.0 ;
      RECT  6795.0 20045.0 6860.0 20180.0 ;
      RECT  7155.0 21020.0 7220.0 21155.0 ;
      RECT  7155.0 20045.0 7220.0 20180.0 ;
      RECT  6852.5 20487.5 6917.5 20622.5 ;
      RECT  6852.5 20487.5 6917.5 20622.5 ;
      RECT  7017.5 20522.5 7082.5 20587.5 ;
      RECT  6727.5 21240.0 7287.5 21305.0 ;
      RECT  6727.5 19895.0 7287.5 19960.0 ;
      RECT  4990.0 20487.5 5055.0 20622.5 ;
      RECT  5130.0 20215.0 5195.0 20350.0 ;
      RECT  6125.0 20320.0 5990.0 20385.0 ;
      RECT  5675.0 21457.5 5740.0 21272.5 ;
      RECT  5675.0 22617.5 5740.0 22432.5 ;
      RECT  5315.0 22500.0 5380.0 22650.0 ;
      RECT  5315.0 21615.0 5380.0 21240.0 ;
      RECT  5505.0 22500.0 5570.0 21615.0 ;
      RECT  5315.0 21615.0 5380.0 21480.0 ;
      RECT  5505.0 21615.0 5570.0 21480.0 ;
      RECT  5505.0 21615.0 5570.0 21480.0 ;
      RECT  5315.0 21615.0 5380.0 21480.0 ;
      RECT  5315.0 22500.0 5380.0 22365.0 ;
      RECT  5505.0 22500.0 5570.0 22365.0 ;
      RECT  5505.0 22500.0 5570.0 22365.0 ;
      RECT  5315.0 22500.0 5380.0 22365.0 ;
      RECT  5675.0 21525.0 5740.0 21390.0 ;
      RECT  5675.0 22500.0 5740.0 22365.0 ;
      RECT  5372.5 22057.5 5437.5 21922.5 ;
      RECT  5372.5 22057.5 5437.5 21922.5 ;
      RECT  5537.5 22022.5 5602.5 21957.5 ;
      RECT  5247.5 21305.0 5807.5 21240.0 ;
      RECT  5247.5 22650.0 5807.5 22585.0 ;
      RECT  5875.0 22455.0 5940.0 22650.0 ;
      RECT  5875.0 21615.0 5940.0 21240.0 ;
      RECT  6255.0 21615.0 6320.0 21240.0 ;
      RECT  6425.0 21457.5 6490.0 21272.5 ;
      RECT  6425.0 22617.5 6490.0 22432.5 ;
      RECT  5875.0 21615.0 5940.0 21480.0 ;
      RECT  6065.0 21615.0 6130.0 21480.0 ;
      RECT  6065.0 21615.0 6130.0 21480.0 ;
      RECT  5875.0 21615.0 5940.0 21480.0 ;
      RECT  6065.0 21615.0 6130.0 21480.0 ;
      RECT  6255.0 21615.0 6320.0 21480.0 ;
      RECT  6255.0 21615.0 6320.0 21480.0 ;
      RECT  6065.0 21615.0 6130.0 21480.0 ;
      RECT  5875.0 22455.0 5940.0 22320.0 ;
      RECT  6065.0 22455.0 6130.0 22320.0 ;
      RECT  6065.0 22455.0 6130.0 22320.0 ;
      RECT  5875.0 22455.0 5940.0 22320.0 ;
      RECT  6065.0 22455.0 6130.0 22320.0 ;
      RECT  6255.0 22455.0 6320.0 22320.0 ;
      RECT  6255.0 22455.0 6320.0 22320.0 ;
      RECT  6065.0 22455.0 6130.0 22320.0 ;
      RECT  6425.0 21525.0 6490.0 21390.0 ;
      RECT  6425.0 22500.0 6490.0 22365.0 ;
      RECT  6260.0 22225.0 6125.0 22160.0 ;
      RECT  6002.5 22010.0 5867.5 21945.0 ;
      RECT  6065.0 21615.0 6130.0 21480.0 ;
      RECT  6255.0 22455.0 6320.0 22320.0 ;
      RECT  6355.0 22010.0 6220.0 21945.0 ;
      RECT  5867.5 22010.0 6002.5 21945.0 ;
      RECT  6125.0 22225.0 6260.0 22160.0 ;
      RECT  6220.0 22010.0 6355.0 21945.0 ;
      RECT  5807.5 21305.0 6727.5 21240.0 ;
      RECT  5807.5 22650.0 6727.5 22585.0 ;
      RECT  7155.0 21457.5 7220.0 21272.5 ;
      RECT  7155.0 22617.5 7220.0 22432.5 ;
      RECT  6795.0 22500.0 6860.0 22650.0 ;
      RECT  6795.0 21615.0 6860.0 21240.0 ;
      RECT  6985.0 22500.0 7050.0 21615.0 ;
      RECT  6795.0 21615.0 6860.0 21480.0 ;
      RECT  6985.0 21615.0 7050.0 21480.0 ;
      RECT  6985.0 21615.0 7050.0 21480.0 ;
      RECT  6795.0 21615.0 6860.0 21480.0 ;
      RECT  6795.0 22500.0 6860.0 22365.0 ;
      RECT  6985.0 22500.0 7050.0 22365.0 ;
      RECT  6985.0 22500.0 7050.0 22365.0 ;
      RECT  6795.0 22500.0 6860.0 22365.0 ;
      RECT  7155.0 21525.0 7220.0 21390.0 ;
      RECT  7155.0 22500.0 7220.0 22365.0 ;
      RECT  6852.5 22057.5 6917.5 21922.5 ;
      RECT  6852.5 22057.5 6917.5 21922.5 ;
      RECT  7017.5 22022.5 7082.5 21957.5 ;
      RECT  6727.5 21305.0 7287.5 21240.0 ;
      RECT  6727.5 22650.0 7287.5 22585.0 ;
      RECT  4990.0 21922.5 5055.0 22057.5 ;
      RECT  5130.0 22195.0 5195.0 22330.0 ;
      RECT  6125.0 22160.0 5990.0 22225.0 ;
      RECT  5675.0 23777.5 5740.0 23962.5 ;
      RECT  5675.0 22617.5 5740.0 22802.5 ;
      RECT  5315.0 22735.0 5380.0 22585.0 ;
      RECT  5315.0 23620.0 5380.0 23995.0 ;
      RECT  5505.0 22735.0 5570.0 23620.0 ;
      RECT  5315.0 23620.0 5380.0 23755.0 ;
      RECT  5505.0 23620.0 5570.0 23755.0 ;
      RECT  5505.0 23620.0 5570.0 23755.0 ;
      RECT  5315.0 23620.0 5380.0 23755.0 ;
      RECT  5315.0 22735.0 5380.0 22870.0 ;
      RECT  5505.0 22735.0 5570.0 22870.0 ;
      RECT  5505.0 22735.0 5570.0 22870.0 ;
      RECT  5315.0 22735.0 5380.0 22870.0 ;
      RECT  5675.0 23710.0 5740.0 23845.0 ;
      RECT  5675.0 22735.0 5740.0 22870.0 ;
      RECT  5372.5 23177.5 5437.5 23312.5 ;
      RECT  5372.5 23177.5 5437.5 23312.5 ;
      RECT  5537.5 23212.5 5602.5 23277.5 ;
      RECT  5247.5 23930.0 5807.5 23995.0 ;
      RECT  5247.5 22585.0 5807.5 22650.0 ;
      RECT  5875.0 22780.0 5940.0 22585.0 ;
      RECT  5875.0 23620.0 5940.0 23995.0 ;
      RECT  6255.0 23620.0 6320.0 23995.0 ;
      RECT  6425.0 23777.5 6490.0 23962.5 ;
      RECT  6425.0 22617.5 6490.0 22802.5 ;
      RECT  5875.0 23620.0 5940.0 23755.0 ;
      RECT  6065.0 23620.0 6130.0 23755.0 ;
      RECT  6065.0 23620.0 6130.0 23755.0 ;
      RECT  5875.0 23620.0 5940.0 23755.0 ;
      RECT  6065.0 23620.0 6130.0 23755.0 ;
      RECT  6255.0 23620.0 6320.0 23755.0 ;
      RECT  6255.0 23620.0 6320.0 23755.0 ;
      RECT  6065.0 23620.0 6130.0 23755.0 ;
      RECT  5875.0 22780.0 5940.0 22915.0 ;
      RECT  6065.0 22780.0 6130.0 22915.0 ;
      RECT  6065.0 22780.0 6130.0 22915.0 ;
      RECT  5875.0 22780.0 5940.0 22915.0 ;
      RECT  6065.0 22780.0 6130.0 22915.0 ;
      RECT  6255.0 22780.0 6320.0 22915.0 ;
      RECT  6255.0 22780.0 6320.0 22915.0 ;
      RECT  6065.0 22780.0 6130.0 22915.0 ;
      RECT  6425.0 23710.0 6490.0 23845.0 ;
      RECT  6425.0 22735.0 6490.0 22870.0 ;
      RECT  6260.0 23010.0 6125.0 23075.0 ;
      RECT  6002.5 23225.0 5867.5 23290.0 ;
      RECT  6065.0 23620.0 6130.0 23755.0 ;
      RECT  6255.0 22780.0 6320.0 22915.0 ;
      RECT  6355.0 23225.0 6220.0 23290.0 ;
      RECT  5867.5 23225.0 6002.5 23290.0 ;
      RECT  6125.0 23010.0 6260.0 23075.0 ;
      RECT  6220.0 23225.0 6355.0 23290.0 ;
      RECT  5807.5 23930.0 6727.5 23995.0 ;
      RECT  5807.5 22585.0 6727.5 22650.0 ;
      RECT  7155.0 23777.5 7220.0 23962.5 ;
      RECT  7155.0 22617.5 7220.0 22802.5 ;
      RECT  6795.0 22735.0 6860.0 22585.0 ;
      RECT  6795.0 23620.0 6860.0 23995.0 ;
      RECT  6985.0 22735.0 7050.0 23620.0 ;
      RECT  6795.0 23620.0 6860.0 23755.0 ;
      RECT  6985.0 23620.0 7050.0 23755.0 ;
      RECT  6985.0 23620.0 7050.0 23755.0 ;
      RECT  6795.0 23620.0 6860.0 23755.0 ;
      RECT  6795.0 22735.0 6860.0 22870.0 ;
      RECT  6985.0 22735.0 7050.0 22870.0 ;
      RECT  6985.0 22735.0 7050.0 22870.0 ;
      RECT  6795.0 22735.0 6860.0 22870.0 ;
      RECT  7155.0 23710.0 7220.0 23845.0 ;
      RECT  7155.0 22735.0 7220.0 22870.0 ;
      RECT  6852.5 23177.5 6917.5 23312.5 ;
      RECT  6852.5 23177.5 6917.5 23312.5 ;
      RECT  7017.5 23212.5 7082.5 23277.5 ;
      RECT  6727.5 23930.0 7287.5 23995.0 ;
      RECT  6727.5 22585.0 7287.5 22650.0 ;
      RECT  4990.0 23177.5 5055.0 23312.5 ;
      RECT  5130.0 22905.0 5195.0 23040.0 ;
      RECT  6125.0 23010.0 5990.0 23075.0 ;
      RECT  5675.0 24147.5 5740.0 23962.5 ;
      RECT  5675.0 25307.5 5740.0 25122.5 ;
      RECT  5315.0 25190.0 5380.0 25340.0 ;
      RECT  5315.0 24305.0 5380.0 23930.0 ;
      RECT  5505.0 25190.0 5570.0 24305.0 ;
      RECT  5315.0 24305.0 5380.0 24170.0 ;
      RECT  5505.0 24305.0 5570.0 24170.0 ;
      RECT  5505.0 24305.0 5570.0 24170.0 ;
      RECT  5315.0 24305.0 5380.0 24170.0 ;
      RECT  5315.0 25190.0 5380.0 25055.0 ;
      RECT  5505.0 25190.0 5570.0 25055.0 ;
      RECT  5505.0 25190.0 5570.0 25055.0 ;
      RECT  5315.0 25190.0 5380.0 25055.0 ;
      RECT  5675.0 24215.0 5740.0 24080.0 ;
      RECT  5675.0 25190.0 5740.0 25055.0 ;
      RECT  5372.5 24747.5 5437.5 24612.5 ;
      RECT  5372.5 24747.5 5437.5 24612.5 ;
      RECT  5537.5 24712.5 5602.5 24647.5 ;
      RECT  5247.5 23995.0 5807.5 23930.0 ;
      RECT  5247.5 25340.0 5807.5 25275.0 ;
      RECT  5875.0 25145.0 5940.0 25340.0 ;
      RECT  5875.0 24305.0 5940.0 23930.0 ;
      RECT  6255.0 24305.0 6320.0 23930.0 ;
      RECT  6425.0 24147.5 6490.0 23962.5 ;
      RECT  6425.0 25307.5 6490.0 25122.5 ;
      RECT  5875.0 24305.0 5940.0 24170.0 ;
      RECT  6065.0 24305.0 6130.0 24170.0 ;
      RECT  6065.0 24305.0 6130.0 24170.0 ;
      RECT  5875.0 24305.0 5940.0 24170.0 ;
      RECT  6065.0 24305.0 6130.0 24170.0 ;
      RECT  6255.0 24305.0 6320.0 24170.0 ;
      RECT  6255.0 24305.0 6320.0 24170.0 ;
      RECT  6065.0 24305.0 6130.0 24170.0 ;
      RECT  5875.0 25145.0 5940.0 25010.0 ;
      RECT  6065.0 25145.0 6130.0 25010.0 ;
      RECT  6065.0 25145.0 6130.0 25010.0 ;
      RECT  5875.0 25145.0 5940.0 25010.0 ;
      RECT  6065.0 25145.0 6130.0 25010.0 ;
      RECT  6255.0 25145.0 6320.0 25010.0 ;
      RECT  6255.0 25145.0 6320.0 25010.0 ;
      RECT  6065.0 25145.0 6130.0 25010.0 ;
      RECT  6425.0 24215.0 6490.0 24080.0 ;
      RECT  6425.0 25190.0 6490.0 25055.0 ;
      RECT  6260.0 24915.0 6125.0 24850.0 ;
      RECT  6002.5 24700.0 5867.5 24635.0 ;
      RECT  6065.0 24305.0 6130.0 24170.0 ;
      RECT  6255.0 25145.0 6320.0 25010.0 ;
      RECT  6355.0 24700.0 6220.0 24635.0 ;
      RECT  5867.5 24700.0 6002.5 24635.0 ;
      RECT  6125.0 24915.0 6260.0 24850.0 ;
      RECT  6220.0 24700.0 6355.0 24635.0 ;
      RECT  5807.5 23995.0 6727.5 23930.0 ;
      RECT  5807.5 25340.0 6727.5 25275.0 ;
      RECT  7155.0 24147.5 7220.0 23962.5 ;
      RECT  7155.0 25307.5 7220.0 25122.5 ;
      RECT  6795.0 25190.0 6860.0 25340.0 ;
      RECT  6795.0 24305.0 6860.0 23930.0 ;
      RECT  6985.0 25190.0 7050.0 24305.0 ;
      RECT  6795.0 24305.0 6860.0 24170.0 ;
      RECT  6985.0 24305.0 7050.0 24170.0 ;
      RECT  6985.0 24305.0 7050.0 24170.0 ;
      RECT  6795.0 24305.0 6860.0 24170.0 ;
      RECT  6795.0 25190.0 6860.0 25055.0 ;
      RECT  6985.0 25190.0 7050.0 25055.0 ;
      RECT  6985.0 25190.0 7050.0 25055.0 ;
      RECT  6795.0 25190.0 6860.0 25055.0 ;
      RECT  7155.0 24215.0 7220.0 24080.0 ;
      RECT  7155.0 25190.0 7220.0 25055.0 ;
      RECT  6852.5 24747.5 6917.5 24612.5 ;
      RECT  6852.5 24747.5 6917.5 24612.5 ;
      RECT  7017.5 24712.5 7082.5 24647.5 ;
      RECT  6727.5 23995.0 7287.5 23930.0 ;
      RECT  6727.5 25340.0 7287.5 25275.0 ;
      RECT  4990.0 24612.5 5055.0 24747.5 ;
      RECT  5130.0 24885.0 5195.0 25020.0 ;
      RECT  6125.0 24850.0 5990.0 24915.0 ;
      RECT  5675.0 26467.5 5740.0 26652.5 ;
      RECT  5675.0 25307.5 5740.0 25492.5 ;
      RECT  5315.0 25425.0 5380.0 25275.0 ;
      RECT  5315.0 26310.0 5380.0 26685.0 ;
      RECT  5505.0 25425.0 5570.0 26310.0 ;
      RECT  5315.0 26310.0 5380.0 26445.0 ;
      RECT  5505.0 26310.0 5570.0 26445.0 ;
      RECT  5505.0 26310.0 5570.0 26445.0 ;
      RECT  5315.0 26310.0 5380.0 26445.0 ;
      RECT  5315.0 25425.0 5380.0 25560.0 ;
      RECT  5505.0 25425.0 5570.0 25560.0 ;
      RECT  5505.0 25425.0 5570.0 25560.0 ;
      RECT  5315.0 25425.0 5380.0 25560.0 ;
      RECT  5675.0 26400.0 5740.0 26535.0 ;
      RECT  5675.0 25425.0 5740.0 25560.0 ;
      RECT  5372.5 25867.5 5437.5 26002.5 ;
      RECT  5372.5 25867.5 5437.5 26002.5 ;
      RECT  5537.5 25902.5 5602.5 25967.5 ;
      RECT  5247.5 26620.0 5807.5 26685.0 ;
      RECT  5247.5 25275.0 5807.5 25340.0 ;
      RECT  5875.0 25470.0 5940.0 25275.0 ;
      RECT  5875.0 26310.0 5940.0 26685.0 ;
      RECT  6255.0 26310.0 6320.0 26685.0 ;
      RECT  6425.0 26467.5 6490.0 26652.5 ;
      RECT  6425.0 25307.5 6490.0 25492.5 ;
      RECT  5875.0 26310.0 5940.0 26445.0 ;
      RECT  6065.0 26310.0 6130.0 26445.0 ;
      RECT  6065.0 26310.0 6130.0 26445.0 ;
      RECT  5875.0 26310.0 5940.0 26445.0 ;
      RECT  6065.0 26310.0 6130.0 26445.0 ;
      RECT  6255.0 26310.0 6320.0 26445.0 ;
      RECT  6255.0 26310.0 6320.0 26445.0 ;
      RECT  6065.0 26310.0 6130.0 26445.0 ;
      RECT  5875.0 25470.0 5940.0 25605.0 ;
      RECT  6065.0 25470.0 6130.0 25605.0 ;
      RECT  6065.0 25470.0 6130.0 25605.0 ;
      RECT  5875.0 25470.0 5940.0 25605.0 ;
      RECT  6065.0 25470.0 6130.0 25605.0 ;
      RECT  6255.0 25470.0 6320.0 25605.0 ;
      RECT  6255.0 25470.0 6320.0 25605.0 ;
      RECT  6065.0 25470.0 6130.0 25605.0 ;
      RECT  6425.0 26400.0 6490.0 26535.0 ;
      RECT  6425.0 25425.0 6490.0 25560.0 ;
      RECT  6260.0 25700.0 6125.0 25765.0 ;
      RECT  6002.5 25915.0 5867.5 25980.0 ;
      RECT  6065.0 26310.0 6130.0 26445.0 ;
      RECT  6255.0 25470.0 6320.0 25605.0 ;
      RECT  6355.0 25915.0 6220.0 25980.0 ;
      RECT  5867.5 25915.0 6002.5 25980.0 ;
      RECT  6125.0 25700.0 6260.0 25765.0 ;
      RECT  6220.0 25915.0 6355.0 25980.0 ;
      RECT  5807.5 26620.0 6727.5 26685.0 ;
      RECT  5807.5 25275.0 6727.5 25340.0 ;
      RECT  7155.0 26467.5 7220.0 26652.5 ;
      RECT  7155.0 25307.5 7220.0 25492.5 ;
      RECT  6795.0 25425.0 6860.0 25275.0 ;
      RECT  6795.0 26310.0 6860.0 26685.0 ;
      RECT  6985.0 25425.0 7050.0 26310.0 ;
      RECT  6795.0 26310.0 6860.0 26445.0 ;
      RECT  6985.0 26310.0 7050.0 26445.0 ;
      RECT  6985.0 26310.0 7050.0 26445.0 ;
      RECT  6795.0 26310.0 6860.0 26445.0 ;
      RECT  6795.0 25425.0 6860.0 25560.0 ;
      RECT  6985.0 25425.0 7050.0 25560.0 ;
      RECT  6985.0 25425.0 7050.0 25560.0 ;
      RECT  6795.0 25425.0 6860.0 25560.0 ;
      RECT  7155.0 26400.0 7220.0 26535.0 ;
      RECT  7155.0 25425.0 7220.0 25560.0 ;
      RECT  6852.5 25867.5 6917.5 26002.5 ;
      RECT  6852.5 25867.5 6917.5 26002.5 ;
      RECT  7017.5 25902.5 7082.5 25967.5 ;
      RECT  6727.5 26620.0 7287.5 26685.0 ;
      RECT  6727.5 25275.0 7287.5 25340.0 ;
      RECT  4990.0 25867.5 5055.0 26002.5 ;
      RECT  5130.0 25595.0 5195.0 25730.0 ;
      RECT  6125.0 25700.0 5990.0 25765.0 ;
      RECT  5675.0 26837.5 5740.0 26652.5 ;
      RECT  5675.0 27997.5 5740.0 27812.5 ;
      RECT  5315.0 27880.0 5380.0 28030.0 ;
      RECT  5315.0 26995.0 5380.0 26620.0 ;
      RECT  5505.0 27880.0 5570.0 26995.0 ;
      RECT  5315.0 26995.0 5380.0 26860.0 ;
      RECT  5505.0 26995.0 5570.0 26860.0 ;
      RECT  5505.0 26995.0 5570.0 26860.0 ;
      RECT  5315.0 26995.0 5380.0 26860.0 ;
      RECT  5315.0 27880.0 5380.0 27745.0 ;
      RECT  5505.0 27880.0 5570.0 27745.0 ;
      RECT  5505.0 27880.0 5570.0 27745.0 ;
      RECT  5315.0 27880.0 5380.0 27745.0 ;
      RECT  5675.0 26905.0 5740.0 26770.0 ;
      RECT  5675.0 27880.0 5740.0 27745.0 ;
      RECT  5372.5 27437.5 5437.5 27302.5 ;
      RECT  5372.5 27437.5 5437.5 27302.5 ;
      RECT  5537.5 27402.5 5602.5 27337.5 ;
      RECT  5247.5 26685.0 5807.5 26620.0 ;
      RECT  5247.5 28030.0 5807.5 27965.0 ;
      RECT  5875.0 27835.0 5940.0 28030.0 ;
      RECT  5875.0 26995.0 5940.0 26620.0 ;
      RECT  6255.0 26995.0 6320.0 26620.0 ;
      RECT  6425.0 26837.5 6490.0 26652.5 ;
      RECT  6425.0 27997.5 6490.0 27812.5 ;
      RECT  5875.0 26995.0 5940.0 26860.0 ;
      RECT  6065.0 26995.0 6130.0 26860.0 ;
      RECT  6065.0 26995.0 6130.0 26860.0 ;
      RECT  5875.0 26995.0 5940.0 26860.0 ;
      RECT  6065.0 26995.0 6130.0 26860.0 ;
      RECT  6255.0 26995.0 6320.0 26860.0 ;
      RECT  6255.0 26995.0 6320.0 26860.0 ;
      RECT  6065.0 26995.0 6130.0 26860.0 ;
      RECT  5875.0 27835.0 5940.0 27700.0 ;
      RECT  6065.0 27835.0 6130.0 27700.0 ;
      RECT  6065.0 27835.0 6130.0 27700.0 ;
      RECT  5875.0 27835.0 5940.0 27700.0 ;
      RECT  6065.0 27835.0 6130.0 27700.0 ;
      RECT  6255.0 27835.0 6320.0 27700.0 ;
      RECT  6255.0 27835.0 6320.0 27700.0 ;
      RECT  6065.0 27835.0 6130.0 27700.0 ;
      RECT  6425.0 26905.0 6490.0 26770.0 ;
      RECT  6425.0 27880.0 6490.0 27745.0 ;
      RECT  6260.0 27605.0 6125.0 27540.0 ;
      RECT  6002.5 27390.0 5867.5 27325.0 ;
      RECT  6065.0 26995.0 6130.0 26860.0 ;
      RECT  6255.0 27835.0 6320.0 27700.0 ;
      RECT  6355.0 27390.0 6220.0 27325.0 ;
      RECT  5867.5 27390.0 6002.5 27325.0 ;
      RECT  6125.0 27605.0 6260.0 27540.0 ;
      RECT  6220.0 27390.0 6355.0 27325.0 ;
      RECT  5807.5 26685.0 6727.5 26620.0 ;
      RECT  5807.5 28030.0 6727.5 27965.0 ;
      RECT  7155.0 26837.5 7220.0 26652.5 ;
      RECT  7155.0 27997.5 7220.0 27812.5 ;
      RECT  6795.0 27880.0 6860.0 28030.0 ;
      RECT  6795.0 26995.0 6860.0 26620.0 ;
      RECT  6985.0 27880.0 7050.0 26995.0 ;
      RECT  6795.0 26995.0 6860.0 26860.0 ;
      RECT  6985.0 26995.0 7050.0 26860.0 ;
      RECT  6985.0 26995.0 7050.0 26860.0 ;
      RECT  6795.0 26995.0 6860.0 26860.0 ;
      RECT  6795.0 27880.0 6860.0 27745.0 ;
      RECT  6985.0 27880.0 7050.0 27745.0 ;
      RECT  6985.0 27880.0 7050.0 27745.0 ;
      RECT  6795.0 27880.0 6860.0 27745.0 ;
      RECT  7155.0 26905.0 7220.0 26770.0 ;
      RECT  7155.0 27880.0 7220.0 27745.0 ;
      RECT  6852.5 27437.5 6917.5 27302.5 ;
      RECT  6852.5 27437.5 6917.5 27302.5 ;
      RECT  7017.5 27402.5 7082.5 27337.5 ;
      RECT  6727.5 26685.0 7287.5 26620.0 ;
      RECT  6727.5 28030.0 7287.5 27965.0 ;
      RECT  4990.0 27302.5 5055.0 27437.5 ;
      RECT  5130.0 27575.0 5195.0 27710.0 ;
      RECT  6125.0 27540.0 5990.0 27605.0 ;
      RECT  5675.0 29157.5 5740.0 29342.5 ;
      RECT  5675.0 27997.5 5740.0 28182.5 ;
      RECT  5315.0 28115.0 5380.0 27965.0 ;
      RECT  5315.0 29000.0 5380.0 29375.0 ;
      RECT  5505.0 28115.0 5570.0 29000.0 ;
      RECT  5315.0 29000.0 5380.0 29135.0 ;
      RECT  5505.0 29000.0 5570.0 29135.0 ;
      RECT  5505.0 29000.0 5570.0 29135.0 ;
      RECT  5315.0 29000.0 5380.0 29135.0 ;
      RECT  5315.0 28115.0 5380.0 28250.0 ;
      RECT  5505.0 28115.0 5570.0 28250.0 ;
      RECT  5505.0 28115.0 5570.0 28250.0 ;
      RECT  5315.0 28115.0 5380.0 28250.0 ;
      RECT  5675.0 29090.0 5740.0 29225.0 ;
      RECT  5675.0 28115.0 5740.0 28250.0 ;
      RECT  5372.5 28557.5 5437.5 28692.5 ;
      RECT  5372.5 28557.5 5437.5 28692.5 ;
      RECT  5537.5 28592.5 5602.5 28657.5 ;
      RECT  5247.5 29310.0 5807.5 29375.0 ;
      RECT  5247.5 27965.0 5807.5 28030.0 ;
      RECT  5875.0 28160.0 5940.0 27965.0 ;
      RECT  5875.0 29000.0 5940.0 29375.0 ;
      RECT  6255.0 29000.0 6320.0 29375.0 ;
      RECT  6425.0 29157.5 6490.0 29342.5 ;
      RECT  6425.0 27997.5 6490.0 28182.5 ;
      RECT  5875.0 29000.0 5940.0 29135.0 ;
      RECT  6065.0 29000.0 6130.0 29135.0 ;
      RECT  6065.0 29000.0 6130.0 29135.0 ;
      RECT  5875.0 29000.0 5940.0 29135.0 ;
      RECT  6065.0 29000.0 6130.0 29135.0 ;
      RECT  6255.0 29000.0 6320.0 29135.0 ;
      RECT  6255.0 29000.0 6320.0 29135.0 ;
      RECT  6065.0 29000.0 6130.0 29135.0 ;
      RECT  5875.0 28160.0 5940.0 28295.0 ;
      RECT  6065.0 28160.0 6130.0 28295.0 ;
      RECT  6065.0 28160.0 6130.0 28295.0 ;
      RECT  5875.0 28160.0 5940.0 28295.0 ;
      RECT  6065.0 28160.0 6130.0 28295.0 ;
      RECT  6255.0 28160.0 6320.0 28295.0 ;
      RECT  6255.0 28160.0 6320.0 28295.0 ;
      RECT  6065.0 28160.0 6130.0 28295.0 ;
      RECT  6425.0 29090.0 6490.0 29225.0 ;
      RECT  6425.0 28115.0 6490.0 28250.0 ;
      RECT  6260.0 28390.0 6125.0 28455.0 ;
      RECT  6002.5 28605.0 5867.5 28670.0 ;
      RECT  6065.0 29000.0 6130.0 29135.0 ;
      RECT  6255.0 28160.0 6320.0 28295.0 ;
      RECT  6355.0 28605.0 6220.0 28670.0 ;
      RECT  5867.5 28605.0 6002.5 28670.0 ;
      RECT  6125.0 28390.0 6260.0 28455.0 ;
      RECT  6220.0 28605.0 6355.0 28670.0 ;
      RECT  5807.5 29310.0 6727.5 29375.0 ;
      RECT  5807.5 27965.0 6727.5 28030.0 ;
      RECT  7155.0 29157.5 7220.0 29342.5 ;
      RECT  7155.0 27997.5 7220.0 28182.5 ;
      RECT  6795.0 28115.0 6860.0 27965.0 ;
      RECT  6795.0 29000.0 6860.0 29375.0 ;
      RECT  6985.0 28115.0 7050.0 29000.0 ;
      RECT  6795.0 29000.0 6860.0 29135.0 ;
      RECT  6985.0 29000.0 7050.0 29135.0 ;
      RECT  6985.0 29000.0 7050.0 29135.0 ;
      RECT  6795.0 29000.0 6860.0 29135.0 ;
      RECT  6795.0 28115.0 6860.0 28250.0 ;
      RECT  6985.0 28115.0 7050.0 28250.0 ;
      RECT  6985.0 28115.0 7050.0 28250.0 ;
      RECT  6795.0 28115.0 6860.0 28250.0 ;
      RECT  7155.0 29090.0 7220.0 29225.0 ;
      RECT  7155.0 28115.0 7220.0 28250.0 ;
      RECT  6852.5 28557.5 6917.5 28692.5 ;
      RECT  6852.5 28557.5 6917.5 28692.5 ;
      RECT  7017.5 28592.5 7082.5 28657.5 ;
      RECT  6727.5 29310.0 7287.5 29375.0 ;
      RECT  6727.5 27965.0 7287.5 28030.0 ;
      RECT  4990.0 28557.5 5055.0 28692.5 ;
      RECT  5130.0 28285.0 5195.0 28420.0 ;
      RECT  6125.0 28390.0 5990.0 28455.0 ;
      RECT  5675.0 29527.5 5740.0 29342.5 ;
      RECT  5675.0 30687.5 5740.0 30502.5 ;
      RECT  5315.0 30570.0 5380.0 30720.0 ;
      RECT  5315.0 29685.0 5380.0 29310.0 ;
      RECT  5505.0 30570.0 5570.0 29685.0 ;
      RECT  5315.0 29685.0 5380.0 29550.0 ;
      RECT  5505.0 29685.0 5570.0 29550.0 ;
      RECT  5505.0 29685.0 5570.0 29550.0 ;
      RECT  5315.0 29685.0 5380.0 29550.0 ;
      RECT  5315.0 30570.0 5380.0 30435.0 ;
      RECT  5505.0 30570.0 5570.0 30435.0 ;
      RECT  5505.0 30570.0 5570.0 30435.0 ;
      RECT  5315.0 30570.0 5380.0 30435.0 ;
      RECT  5675.0 29595.0 5740.0 29460.0 ;
      RECT  5675.0 30570.0 5740.0 30435.0 ;
      RECT  5372.5 30127.5 5437.5 29992.5 ;
      RECT  5372.5 30127.5 5437.5 29992.5 ;
      RECT  5537.5 30092.5 5602.5 30027.5 ;
      RECT  5247.5 29375.0 5807.5 29310.0 ;
      RECT  5247.5 30720.0 5807.5 30655.0 ;
      RECT  5875.0 30525.0 5940.0 30720.0 ;
      RECT  5875.0 29685.0 5940.0 29310.0 ;
      RECT  6255.0 29685.0 6320.0 29310.0 ;
      RECT  6425.0 29527.5 6490.0 29342.5 ;
      RECT  6425.0 30687.5 6490.0 30502.5 ;
      RECT  5875.0 29685.0 5940.0 29550.0 ;
      RECT  6065.0 29685.0 6130.0 29550.0 ;
      RECT  6065.0 29685.0 6130.0 29550.0 ;
      RECT  5875.0 29685.0 5940.0 29550.0 ;
      RECT  6065.0 29685.0 6130.0 29550.0 ;
      RECT  6255.0 29685.0 6320.0 29550.0 ;
      RECT  6255.0 29685.0 6320.0 29550.0 ;
      RECT  6065.0 29685.0 6130.0 29550.0 ;
      RECT  5875.0 30525.0 5940.0 30390.0 ;
      RECT  6065.0 30525.0 6130.0 30390.0 ;
      RECT  6065.0 30525.0 6130.0 30390.0 ;
      RECT  5875.0 30525.0 5940.0 30390.0 ;
      RECT  6065.0 30525.0 6130.0 30390.0 ;
      RECT  6255.0 30525.0 6320.0 30390.0 ;
      RECT  6255.0 30525.0 6320.0 30390.0 ;
      RECT  6065.0 30525.0 6130.0 30390.0 ;
      RECT  6425.0 29595.0 6490.0 29460.0 ;
      RECT  6425.0 30570.0 6490.0 30435.0 ;
      RECT  6260.0 30295.0 6125.0 30230.0 ;
      RECT  6002.5 30080.0 5867.5 30015.0 ;
      RECT  6065.0 29685.0 6130.0 29550.0 ;
      RECT  6255.0 30525.0 6320.0 30390.0 ;
      RECT  6355.0 30080.0 6220.0 30015.0 ;
      RECT  5867.5 30080.0 6002.5 30015.0 ;
      RECT  6125.0 30295.0 6260.0 30230.0 ;
      RECT  6220.0 30080.0 6355.0 30015.0 ;
      RECT  5807.5 29375.0 6727.5 29310.0 ;
      RECT  5807.5 30720.0 6727.5 30655.0 ;
      RECT  7155.0 29527.5 7220.0 29342.5 ;
      RECT  7155.0 30687.5 7220.0 30502.5 ;
      RECT  6795.0 30570.0 6860.0 30720.0 ;
      RECT  6795.0 29685.0 6860.0 29310.0 ;
      RECT  6985.0 30570.0 7050.0 29685.0 ;
      RECT  6795.0 29685.0 6860.0 29550.0 ;
      RECT  6985.0 29685.0 7050.0 29550.0 ;
      RECT  6985.0 29685.0 7050.0 29550.0 ;
      RECT  6795.0 29685.0 6860.0 29550.0 ;
      RECT  6795.0 30570.0 6860.0 30435.0 ;
      RECT  6985.0 30570.0 7050.0 30435.0 ;
      RECT  6985.0 30570.0 7050.0 30435.0 ;
      RECT  6795.0 30570.0 6860.0 30435.0 ;
      RECT  7155.0 29595.0 7220.0 29460.0 ;
      RECT  7155.0 30570.0 7220.0 30435.0 ;
      RECT  6852.5 30127.5 6917.5 29992.5 ;
      RECT  6852.5 30127.5 6917.5 29992.5 ;
      RECT  7017.5 30092.5 7082.5 30027.5 ;
      RECT  6727.5 29375.0 7287.5 29310.0 ;
      RECT  6727.5 30720.0 7287.5 30655.0 ;
      RECT  4990.0 29992.5 5055.0 30127.5 ;
      RECT  5130.0 30265.0 5195.0 30400.0 ;
      RECT  6125.0 30230.0 5990.0 30295.0 ;
      RECT  5675.0 31847.5 5740.0 32032.5 ;
      RECT  5675.0 30687.5 5740.0 30872.5 ;
      RECT  5315.0 30805.0 5380.0 30655.0 ;
      RECT  5315.0 31690.0 5380.0 32065.0 ;
      RECT  5505.0 30805.0 5570.0 31690.0 ;
      RECT  5315.0 31690.0 5380.0 31825.0 ;
      RECT  5505.0 31690.0 5570.0 31825.0 ;
      RECT  5505.0 31690.0 5570.0 31825.0 ;
      RECT  5315.0 31690.0 5380.0 31825.0 ;
      RECT  5315.0 30805.0 5380.0 30940.0 ;
      RECT  5505.0 30805.0 5570.0 30940.0 ;
      RECT  5505.0 30805.0 5570.0 30940.0 ;
      RECT  5315.0 30805.0 5380.0 30940.0 ;
      RECT  5675.0 31780.0 5740.0 31915.0 ;
      RECT  5675.0 30805.0 5740.0 30940.0 ;
      RECT  5372.5 31247.5 5437.5 31382.5 ;
      RECT  5372.5 31247.5 5437.5 31382.5 ;
      RECT  5537.5 31282.5 5602.5 31347.5 ;
      RECT  5247.5 32000.0 5807.5 32065.0 ;
      RECT  5247.5 30655.0 5807.5 30720.0 ;
      RECT  5875.0 30850.0 5940.0 30655.0 ;
      RECT  5875.0 31690.0 5940.0 32065.0 ;
      RECT  6255.0 31690.0 6320.0 32065.0 ;
      RECT  6425.0 31847.5 6490.0 32032.5 ;
      RECT  6425.0 30687.5 6490.0 30872.5 ;
      RECT  5875.0 31690.0 5940.0 31825.0 ;
      RECT  6065.0 31690.0 6130.0 31825.0 ;
      RECT  6065.0 31690.0 6130.0 31825.0 ;
      RECT  5875.0 31690.0 5940.0 31825.0 ;
      RECT  6065.0 31690.0 6130.0 31825.0 ;
      RECT  6255.0 31690.0 6320.0 31825.0 ;
      RECT  6255.0 31690.0 6320.0 31825.0 ;
      RECT  6065.0 31690.0 6130.0 31825.0 ;
      RECT  5875.0 30850.0 5940.0 30985.0 ;
      RECT  6065.0 30850.0 6130.0 30985.0 ;
      RECT  6065.0 30850.0 6130.0 30985.0 ;
      RECT  5875.0 30850.0 5940.0 30985.0 ;
      RECT  6065.0 30850.0 6130.0 30985.0 ;
      RECT  6255.0 30850.0 6320.0 30985.0 ;
      RECT  6255.0 30850.0 6320.0 30985.0 ;
      RECT  6065.0 30850.0 6130.0 30985.0 ;
      RECT  6425.0 31780.0 6490.0 31915.0 ;
      RECT  6425.0 30805.0 6490.0 30940.0 ;
      RECT  6260.0 31080.0 6125.0 31145.0 ;
      RECT  6002.5 31295.0 5867.5 31360.0 ;
      RECT  6065.0 31690.0 6130.0 31825.0 ;
      RECT  6255.0 30850.0 6320.0 30985.0 ;
      RECT  6355.0 31295.0 6220.0 31360.0 ;
      RECT  5867.5 31295.0 6002.5 31360.0 ;
      RECT  6125.0 31080.0 6260.0 31145.0 ;
      RECT  6220.0 31295.0 6355.0 31360.0 ;
      RECT  5807.5 32000.0 6727.5 32065.0 ;
      RECT  5807.5 30655.0 6727.5 30720.0 ;
      RECT  7155.0 31847.5 7220.0 32032.5 ;
      RECT  7155.0 30687.5 7220.0 30872.5 ;
      RECT  6795.0 30805.0 6860.0 30655.0 ;
      RECT  6795.0 31690.0 6860.0 32065.0 ;
      RECT  6985.0 30805.0 7050.0 31690.0 ;
      RECT  6795.0 31690.0 6860.0 31825.0 ;
      RECT  6985.0 31690.0 7050.0 31825.0 ;
      RECT  6985.0 31690.0 7050.0 31825.0 ;
      RECT  6795.0 31690.0 6860.0 31825.0 ;
      RECT  6795.0 30805.0 6860.0 30940.0 ;
      RECT  6985.0 30805.0 7050.0 30940.0 ;
      RECT  6985.0 30805.0 7050.0 30940.0 ;
      RECT  6795.0 30805.0 6860.0 30940.0 ;
      RECT  7155.0 31780.0 7220.0 31915.0 ;
      RECT  7155.0 30805.0 7220.0 30940.0 ;
      RECT  6852.5 31247.5 6917.5 31382.5 ;
      RECT  6852.5 31247.5 6917.5 31382.5 ;
      RECT  7017.5 31282.5 7082.5 31347.5 ;
      RECT  6727.5 32000.0 7287.5 32065.0 ;
      RECT  6727.5 30655.0 7287.5 30720.0 ;
      RECT  4990.0 31247.5 5055.0 31382.5 ;
      RECT  5130.0 30975.0 5195.0 31110.0 ;
      RECT  6125.0 31080.0 5990.0 31145.0 ;
      RECT  5675.0 32217.5 5740.0 32032.5 ;
      RECT  5675.0 33377.5 5740.0 33192.5 ;
      RECT  5315.0 33260.0 5380.0 33410.0 ;
      RECT  5315.0 32375.0 5380.0 32000.0 ;
      RECT  5505.0 33260.0 5570.0 32375.0 ;
      RECT  5315.0 32375.0 5380.0 32240.0 ;
      RECT  5505.0 32375.0 5570.0 32240.0 ;
      RECT  5505.0 32375.0 5570.0 32240.0 ;
      RECT  5315.0 32375.0 5380.0 32240.0 ;
      RECT  5315.0 33260.0 5380.0 33125.0 ;
      RECT  5505.0 33260.0 5570.0 33125.0 ;
      RECT  5505.0 33260.0 5570.0 33125.0 ;
      RECT  5315.0 33260.0 5380.0 33125.0 ;
      RECT  5675.0 32285.0 5740.0 32150.0 ;
      RECT  5675.0 33260.0 5740.0 33125.0 ;
      RECT  5372.5 32817.5 5437.5 32682.5 ;
      RECT  5372.5 32817.5 5437.5 32682.5 ;
      RECT  5537.5 32782.5 5602.5 32717.5 ;
      RECT  5247.5 32065.0 5807.5 32000.0 ;
      RECT  5247.5 33410.0 5807.5 33345.0 ;
      RECT  5875.0 33215.0 5940.0 33410.0 ;
      RECT  5875.0 32375.0 5940.0 32000.0 ;
      RECT  6255.0 32375.0 6320.0 32000.0 ;
      RECT  6425.0 32217.5 6490.0 32032.5 ;
      RECT  6425.0 33377.5 6490.0 33192.5 ;
      RECT  5875.0 32375.0 5940.0 32240.0 ;
      RECT  6065.0 32375.0 6130.0 32240.0 ;
      RECT  6065.0 32375.0 6130.0 32240.0 ;
      RECT  5875.0 32375.0 5940.0 32240.0 ;
      RECT  6065.0 32375.0 6130.0 32240.0 ;
      RECT  6255.0 32375.0 6320.0 32240.0 ;
      RECT  6255.0 32375.0 6320.0 32240.0 ;
      RECT  6065.0 32375.0 6130.0 32240.0 ;
      RECT  5875.0 33215.0 5940.0 33080.0 ;
      RECT  6065.0 33215.0 6130.0 33080.0 ;
      RECT  6065.0 33215.0 6130.0 33080.0 ;
      RECT  5875.0 33215.0 5940.0 33080.0 ;
      RECT  6065.0 33215.0 6130.0 33080.0 ;
      RECT  6255.0 33215.0 6320.0 33080.0 ;
      RECT  6255.0 33215.0 6320.0 33080.0 ;
      RECT  6065.0 33215.0 6130.0 33080.0 ;
      RECT  6425.0 32285.0 6490.0 32150.0 ;
      RECT  6425.0 33260.0 6490.0 33125.0 ;
      RECT  6260.0 32985.0 6125.0 32920.0 ;
      RECT  6002.5 32770.0 5867.5 32705.0 ;
      RECT  6065.0 32375.0 6130.0 32240.0 ;
      RECT  6255.0 33215.0 6320.0 33080.0 ;
      RECT  6355.0 32770.0 6220.0 32705.0 ;
      RECT  5867.5 32770.0 6002.5 32705.0 ;
      RECT  6125.0 32985.0 6260.0 32920.0 ;
      RECT  6220.0 32770.0 6355.0 32705.0 ;
      RECT  5807.5 32065.0 6727.5 32000.0 ;
      RECT  5807.5 33410.0 6727.5 33345.0 ;
      RECT  7155.0 32217.5 7220.0 32032.5 ;
      RECT  7155.0 33377.5 7220.0 33192.5 ;
      RECT  6795.0 33260.0 6860.0 33410.0 ;
      RECT  6795.0 32375.0 6860.0 32000.0 ;
      RECT  6985.0 33260.0 7050.0 32375.0 ;
      RECT  6795.0 32375.0 6860.0 32240.0 ;
      RECT  6985.0 32375.0 7050.0 32240.0 ;
      RECT  6985.0 32375.0 7050.0 32240.0 ;
      RECT  6795.0 32375.0 6860.0 32240.0 ;
      RECT  6795.0 33260.0 6860.0 33125.0 ;
      RECT  6985.0 33260.0 7050.0 33125.0 ;
      RECT  6985.0 33260.0 7050.0 33125.0 ;
      RECT  6795.0 33260.0 6860.0 33125.0 ;
      RECT  7155.0 32285.0 7220.0 32150.0 ;
      RECT  7155.0 33260.0 7220.0 33125.0 ;
      RECT  6852.5 32817.5 6917.5 32682.5 ;
      RECT  6852.5 32817.5 6917.5 32682.5 ;
      RECT  7017.5 32782.5 7082.5 32717.5 ;
      RECT  6727.5 32065.0 7287.5 32000.0 ;
      RECT  6727.5 33410.0 7287.5 33345.0 ;
      RECT  4990.0 32682.5 5055.0 32817.5 ;
      RECT  5130.0 32955.0 5195.0 33090.0 ;
      RECT  6125.0 32920.0 5990.0 32985.0 ;
      RECT  5675.0 34537.5 5740.0 34722.5 ;
      RECT  5675.0 33377.5 5740.0 33562.5 ;
      RECT  5315.0 33495.0 5380.0 33345.0 ;
      RECT  5315.0 34380.0 5380.0 34755.0 ;
      RECT  5505.0 33495.0 5570.0 34380.0 ;
      RECT  5315.0 34380.0 5380.0 34515.0 ;
      RECT  5505.0 34380.0 5570.0 34515.0 ;
      RECT  5505.0 34380.0 5570.0 34515.0 ;
      RECT  5315.0 34380.0 5380.0 34515.0 ;
      RECT  5315.0 33495.0 5380.0 33630.0 ;
      RECT  5505.0 33495.0 5570.0 33630.0 ;
      RECT  5505.0 33495.0 5570.0 33630.0 ;
      RECT  5315.0 33495.0 5380.0 33630.0 ;
      RECT  5675.0 34470.0 5740.0 34605.0 ;
      RECT  5675.0 33495.0 5740.0 33630.0 ;
      RECT  5372.5 33937.5 5437.5 34072.5 ;
      RECT  5372.5 33937.5 5437.5 34072.5 ;
      RECT  5537.5 33972.5 5602.5 34037.5 ;
      RECT  5247.5 34690.0 5807.5 34755.0 ;
      RECT  5247.5 33345.0 5807.5 33410.0 ;
      RECT  5875.0 33540.0 5940.0 33345.0 ;
      RECT  5875.0 34380.0 5940.0 34755.0 ;
      RECT  6255.0 34380.0 6320.0 34755.0 ;
      RECT  6425.0 34537.5 6490.0 34722.5 ;
      RECT  6425.0 33377.5 6490.0 33562.5 ;
      RECT  5875.0 34380.0 5940.0 34515.0 ;
      RECT  6065.0 34380.0 6130.0 34515.0 ;
      RECT  6065.0 34380.0 6130.0 34515.0 ;
      RECT  5875.0 34380.0 5940.0 34515.0 ;
      RECT  6065.0 34380.0 6130.0 34515.0 ;
      RECT  6255.0 34380.0 6320.0 34515.0 ;
      RECT  6255.0 34380.0 6320.0 34515.0 ;
      RECT  6065.0 34380.0 6130.0 34515.0 ;
      RECT  5875.0 33540.0 5940.0 33675.0 ;
      RECT  6065.0 33540.0 6130.0 33675.0 ;
      RECT  6065.0 33540.0 6130.0 33675.0 ;
      RECT  5875.0 33540.0 5940.0 33675.0 ;
      RECT  6065.0 33540.0 6130.0 33675.0 ;
      RECT  6255.0 33540.0 6320.0 33675.0 ;
      RECT  6255.0 33540.0 6320.0 33675.0 ;
      RECT  6065.0 33540.0 6130.0 33675.0 ;
      RECT  6425.0 34470.0 6490.0 34605.0 ;
      RECT  6425.0 33495.0 6490.0 33630.0 ;
      RECT  6260.0 33770.0 6125.0 33835.0 ;
      RECT  6002.5 33985.0 5867.5 34050.0 ;
      RECT  6065.0 34380.0 6130.0 34515.0 ;
      RECT  6255.0 33540.0 6320.0 33675.0 ;
      RECT  6355.0 33985.0 6220.0 34050.0 ;
      RECT  5867.5 33985.0 6002.5 34050.0 ;
      RECT  6125.0 33770.0 6260.0 33835.0 ;
      RECT  6220.0 33985.0 6355.0 34050.0 ;
      RECT  5807.5 34690.0 6727.5 34755.0 ;
      RECT  5807.5 33345.0 6727.5 33410.0 ;
      RECT  7155.0 34537.5 7220.0 34722.5 ;
      RECT  7155.0 33377.5 7220.0 33562.5 ;
      RECT  6795.0 33495.0 6860.0 33345.0 ;
      RECT  6795.0 34380.0 6860.0 34755.0 ;
      RECT  6985.0 33495.0 7050.0 34380.0 ;
      RECT  6795.0 34380.0 6860.0 34515.0 ;
      RECT  6985.0 34380.0 7050.0 34515.0 ;
      RECT  6985.0 34380.0 7050.0 34515.0 ;
      RECT  6795.0 34380.0 6860.0 34515.0 ;
      RECT  6795.0 33495.0 6860.0 33630.0 ;
      RECT  6985.0 33495.0 7050.0 33630.0 ;
      RECT  6985.0 33495.0 7050.0 33630.0 ;
      RECT  6795.0 33495.0 6860.0 33630.0 ;
      RECT  7155.0 34470.0 7220.0 34605.0 ;
      RECT  7155.0 33495.0 7220.0 33630.0 ;
      RECT  6852.5 33937.5 6917.5 34072.5 ;
      RECT  6852.5 33937.5 6917.5 34072.5 ;
      RECT  7017.5 33972.5 7082.5 34037.5 ;
      RECT  6727.5 34690.0 7287.5 34755.0 ;
      RECT  6727.5 33345.0 7287.5 33410.0 ;
      RECT  4990.0 33937.5 5055.0 34072.5 ;
      RECT  5130.0 33665.0 5195.0 33800.0 ;
      RECT  6125.0 33770.0 5990.0 33835.0 ;
      RECT  5675.0 34907.5 5740.0 34722.5 ;
      RECT  5675.0 36067.5 5740.0 35882.5 ;
      RECT  5315.0 35950.0 5380.0 36100.0 ;
      RECT  5315.0 35065.0 5380.0 34690.0 ;
      RECT  5505.0 35950.0 5570.0 35065.0 ;
      RECT  5315.0 35065.0 5380.0 34930.0 ;
      RECT  5505.0 35065.0 5570.0 34930.0 ;
      RECT  5505.0 35065.0 5570.0 34930.0 ;
      RECT  5315.0 35065.0 5380.0 34930.0 ;
      RECT  5315.0 35950.0 5380.0 35815.0 ;
      RECT  5505.0 35950.0 5570.0 35815.0 ;
      RECT  5505.0 35950.0 5570.0 35815.0 ;
      RECT  5315.0 35950.0 5380.0 35815.0 ;
      RECT  5675.0 34975.0 5740.0 34840.0 ;
      RECT  5675.0 35950.0 5740.0 35815.0 ;
      RECT  5372.5 35507.5 5437.5 35372.5 ;
      RECT  5372.5 35507.5 5437.5 35372.5 ;
      RECT  5537.5 35472.5 5602.5 35407.5 ;
      RECT  5247.5 34755.0 5807.5 34690.0 ;
      RECT  5247.5 36100.0 5807.5 36035.0 ;
      RECT  5875.0 35905.0 5940.0 36100.0 ;
      RECT  5875.0 35065.0 5940.0 34690.0 ;
      RECT  6255.0 35065.0 6320.0 34690.0 ;
      RECT  6425.0 34907.5 6490.0 34722.5 ;
      RECT  6425.0 36067.5 6490.0 35882.5 ;
      RECT  5875.0 35065.0 5940.0 34930.0 ;
      RECT  6065.0 35065.0 6130.0 34930.0 ;
      RECT  6065.0 35065.0 6130.0 34930.0 ;
      RECT  5875.0 35065.0 5940.0 34930.0 ;
      RECT  6065.0 35065.0 6130.0 34930.0 ;
      RECT  6255.0 35065.0 6320.0 34930.0 ;
      RECT  6255.0 35065.0 6320.0 34930.0 ;
      RECT  6065.0 35065.0 6130.0 34930.0 ;
      RECT  5875.0 35905.0 5940.0 35770.0 ;
      RECT  6065.0 35905.0 6130.0 35770.0 ;
      RECT  6065.0 35905.0 6130.0 35770.0 ;
      RECT  5875.0 35905.0 5940.0 35770.0 ;
      RECT  6065.0 35905.0 6130.0 35770.0 ;
      RECT  6255.0 35905.0 6320.0 35770.0 ;
      RECT  6255.0 35905.0 6320.0 35770.0 ;
      RECT  6065.0 35905.0 6130.0 35770.0 ;
      RECT  6425.0 34975.0 6490.0 34840.0 ;
      RECT  6425.0 35950.0 6490.0 35815.0 ;
      RECT  6260.0 35675.0 6125.0 35610.0 ;
      RECT  6002.5 35460.0 5867.5 35395.0 ;
      RECT  6065.0 35065.0 6130.0 34930.0 ;
      RECT  6255.0 35905.0 6320.0 35770.0 ;
      RECT  6355.0 35460.0 6220.0 35395.0 ;
      RECT  5867.5 35460.0 6002.5 35395.0 ;
      RECT  6125.0 35675.0 6260.0 35610.0 ;
      RECT  6220.0 35460.0 6355.0 35395.0 ;
      RECT  5807.5 34755.0 6727.5 34690.0 ;
      RECT  5807.5 36100.0 6727.5 36035.0 ;
      RECT  7155.0 34907.5 7220.0 34722.5 ;
      RECT  7155.0 36067.5 7220.0 35882.5 ;
      RECT  6795.0 35950.0 6860.0 36100.0 ;
      RECT  6795.0 35065.0 6860.0 34690.0 ;
      RECT  6985.0 35950.0 7050.0 35065.0 ;
      RECT  6795.0 35065.0 6860.0 34930.0 ;
      RECT  6985.0 35065.0 7050.0 34930.0 ;
      RECT  6985.0 35065.0 7050.0 34930.0 ;
      RECT  6795.0 35065.0 6860.0 34930.0 ;
      RECT  6795.0 35950.0 6860.0 35815.0 ;
      RECT  6985.0 35950.0 7050.0 35815.0 ;
      RECT  6985.0 35950.0 7050.0 35815.0 ;
      RECT  6795.0 35950.0 6860.0 35815.0 ;
      RECT  7155.0 34975.0 7220.0 34840.0 ;
      RECT  7155.0 35950.0 7220.0 35815.0 ;
      RECT  6852.5 35507.5 6917.5 35372.5 ;
      RECT  6852.5 35507.5 6917.5 35372.5 ;
      RECT  7017.5 35472.5 7082.5 35407.5 ;
      RECT  6727.5 34755.0 7287.5 34690.0 ;
      RECT  6727.5 36100.0 7287.5 36035.0 ;
      RECT  4990.0 35372.5 5055.0 35507.5 ;
      RECT  5130.0 35645.0 5195.0 35780.0 ;
      RECT  6125.0 35610.0 5990.0 35675.0 ;
      RECT  5675.0 37227.5 5740.0 37412.5 ;
      RECT  5675.0 36067.5 5740.0 36252.5 ;
      RECT  5315.0 36185.0 5380.0 36035.0 ;
      RECT  5315.0 37070.0 5380.0 37445.0 ;
      RECT  5505.0 36185.0 5570.0 37070.0 ;
      RECT  5315.0 37070.0 5380.0 37205.0 ;
      RECT  5505.0 37070.0 5570.0 37205.0 ;
      RECT  5505.0 37070.0 5570.0 37205.0 ;
      RECT  5315.0 37070.0 5380.0 37205.0 ;
      RECT  5315.0 36185.0 5380.0 36320.0 ;
      RECT  5505.0 36185.0 5570.0 36320.0 ;
      RECT  5505.0 36185.0 5570.0 36320.0 ;
      RECT  5315.0 36185.0 5380.0 36320.0 ;
      RECT  5675.0 37160.0 5740.0 37295.0 ;
      RECT  5675.0 36185.0 5740.0 36320.0 ;
      RECT  5372.5 36627.5 5437.5 36762.5 ;
      RECT  5372.5 36627.5 5437.5 36762.5 ;
      RECT  5537.5 36662.5 5602.5 36727.5 ;
      RECT  5247.5 37380.0 5807.5 37445.0 ;
      RECT  5247.5 36035.0 5807.5 36100.0 ;
      RECT  5875.0 36230.0 5940.0 36035.0 ;
      RECT  5875.0 37070.0 5940.0 37445.0 ;
      RECT  6255.0 37070.0 6320.0 37445.0 ;
      RECT  6425.0 37227.5 6490.0 37412.5 ;
      RECT  6425.0 36067.5 6490.0 36252.5 ;
      RECT  5875.0 37070.0 5940.0 37205.0 ;
      RECT  6065.0 37070.0 6130.0 37205.0 ;
      RECT  6065.0 37070.0 6130.0 37205.0 ;
      RECT  5875.0 37070.0 5940.0 37205.0 ;
      RECT  6065.0 37070.0 6130.0 37205.0 ;
      RECT  6255.0 37070.0 6320.0 37205.0 ;
      RECT  6255.0 37070.0 6320.0 37205.0 ;
      RECT  6065.0 37070.0 6130.0 37205.0 ;
      RECT  5875.0 36230.0 5940.0 36365.0 ;
      RECT  6065.0 36230.0 6130.0 36365.0 ;
      RECT  6065.0 36230.0 6130.0 36365.0 ;
      RECT  5875.0 36230.0 5940.0 36365.0 ;
      RECT  6065.0 36230.0 6130.0 36365.0 ;
      RECT  6255.0 36230.0 6320.0 36365.0 ;
      RECT  6255.0 36230.0 6320.0 36365.0 ;
      RECT  6065.0 36230.0 6130.0 36365.0 ;
      RECT  6425.0 37160.0 6490.0 37295.0 ;
      RECT  6425.0 36185.0 6490.0 36320.0 ;
      RECT  6260.0 36460.0 6125.0 36525.0 ;
      RECT  6002.5 36675.0 5867.5 36740.0 ;
      RECT  6065.0 37070.0 6130.0 37205.0 ;
      RECT  6255.0 36230.0 6320.0 36365.0 ;
      RECT  6355.0 36675.0 6220.0 36740.0 ;
      RECT  5867.5 36675.0 6002.5 36740.0 ;
      RECT  6125.0 36460.0 6260.0 36525.0 ;
      RECT  6220.0 36675.0 6355.0 36740.0 ;
      RECT  5807.5 37380.0 6727.5 37445.0 ;
      RECT  5807.5 36035.0 6727.5 36100.0 ;
      RECT  7155.0 37227.5 7220.0 37412.5 ;
      RECT  7155.0 36067.5 7220.0 36252.5 ;
      RECT  6795.0 36185.0 6860.0 36035.0 ;
      RECT  6795.0 37070.0 6860.0 37445.0 ;
      RECT  6985.0 36185.0 7050.0 37070.0 ;
      RECT  6795.0 37070.0 6860.0 37205.0 ;
      RECT  6985.0 37070.0 7050.0 37205.0 ;
      RECT  6985.0 37070.0 7050.0 37205.0 ;
      RECT  6795.0 37070.0 6860.0 37205.0 ;
      RECT  6795.0 36185.0 6860.0 36320.0 ;
      RECT  6985.0 36185.0 7050.0 36320.0 ;
      RECT  6985.0 36185.0 7050.0 36320.0 ;
      RECT  6795.0 36185.0 6860.0 36320.0 ;
      RECT  7155.0 37160.0 7220.0 37295.0 ;
      RECT  7155.0 36185.0 7220.0 36320.0 ;
      RECT  6852.5 36627.5 6917.5 36762.5 ;
      RECT  6852.5 36627.5 6917.5 36762.5 ;
      RECT  7017.5 36662.5 7082.5 36727.5 ;
      RECT  6727.5 37380.0 7287.5 37445.0 ;
      RECT  6727.5 36035.0 7287.5 36100.0 ;
      RECT  4990.0 36627.5 5055.0 36762.5 ;
      RECT  5130.0 36355.0 5195.0 36490.0 ;
      RECT  6125.0 36460.0 5990.0 36525.0 ;
      RECT  5675.0 37597.5 5740.0 37412.5 ;
      RECT  5675.0 38757.5 5740.0 38572.5 ;
      RECT  5315.0 38640.0 5380.0 38790.0 ;
      RECT  5315.0 37755.0 5380.0 37380.0 ;
      RECT  5505.0 38640.0 5570.0 37755.0 ;
      RECT  5315.0 37755.0 5380.0 37620.0 ;
      RECT  5505.0 37755.0 5570.0 37620.0 ;
      RECT  5505.0 37755.0 5570.0 37620.0 ;
      RECT  5315.0 37755.0 5380.0 37620.0 ;
      RECT  5315.0 38640.0 5380.0 38505.0 ;
      RECT  5505.0 38640.0 5570.0 38505.0 ;
      RECT  5505.0 38640.0 5570.0 38505.0 ;
      RECT  5315.0 38640.0 5380.0 38505.0 ;
      RECT  5675.0 37665.0 5740.0 37530.0 ;
      RECT  5675.0 38640.0 5740.0 38505.0 ;
      RECT  5372.5 38197.5 5437.5 38062.5 ;
      RECT  5372.5 38197.5 5437.5 38062.5 ;
      RECT  5537.5 38162.5 5602.5 38097.5 ;
      RECT  5247.5 37445.0 5807.5 37380.0 ;
      RECT  5247.5 38790.0 5807.5 38725.0 ;
      RECT  5875.0 38595.0 5940.0 38790.0 ;
      RECT  5875.0 37755.0 5940.0 37380.0 ;
      RECT  6255.0 37755.0 6320.0 37380.0 ;
      RECT  6425.0 37597.5 6490.0 37412.5 ;
      RECT  6425.0 38757.5 6490.0 38572.5 ;
      RECT  5875.0 37755.0 5940.0 37620.0 ;
      RECT  6065.0 37755.0 6130.0 37620.0 ;
      RECT  6065.0 37755.0 6130.0 37620.0 ;
      RECT  5875.0 37755.0 5940.0 37620.0 ;
      RECT  6065.0 37755.0 6130.0 37620.0 ;
      RECT  6255.0 37755.0 6320.0 37620.0 ;
      RECT  6255.0 37755.0 6320.0 37620.0 ;
      RECT  6065.0 37755.0 6130.0 37620.0 ;
      RECT  5875.0 38595.0 5940.0 38460.0 ;
      RECT  6065.0 38595.0 6130.0 38460.0 ;
      RECT  6065.0 38595.0 6130.0 38460.0 ;
      RECT  5875.0 38595.0 5940.0 38460.0 ;
      RECT  6065.0 38595.0 6130.0 38460.0 ;
      RECT  6255.0 38595.0 6320.0 38460.0 ;
      RECT  6255.0 38595.0 6320.0 38460.0 ;
      RECT  6065.0 38595.0 6130.0 38460.0 ;
      RECT  6425.0 37665.0 6490.0 37530.0 ;
      RECT  6425.0 38640.0 6490.0 38505.0 ;
      RECT  6260.0 38365.0 6125.0 38300.0 ;
      RECT  6002.5 38150.0 5867.5 38085.0 ;
      RECT  6065.0 37755.0 6130.0 37620.0 ;
      RECT  6255.0 38595.0 6320.0 38460.0 ;
      RECT  6355.0 38150.0 6220.0 38085.0 ;
      RECT  5867.5 38150.0 6002.5 38085.0 ;
      RECT  6125.0 38365.0 6260.0 38300.0 ;
      RECT  6220.0 38150.0 6355.0 38085.0 ;
      RECT  5807.5 37445.0 6727.5 37380.0 ;
      RECT  5807.5 38790.0 6727.5 38725.0 ;
      RECT  7155.0 37597.5 7220.0 37412.5 ;
      RECT  7155.0 38757.5 7220.0 38572.5 ;
      RECT  6795.0 38640.0 6860.0 38790.0 ;
      RECT  6795.0 37755.0 6860.0 37380.0 ;
      RECT  6985.0 38640.0 7050.0 37755.0 ;
      RECT  6795.0 37755.0 6860.0 37620.0 ;
      RECT  6985.0 37755.0 7050.0 37620.0 ;
      RECT  6985.0 37755.0 7050.0 37620.0 ;
      RECT  6795.0 37755.0 6860.0 37620.0 ;
      RECT  6795.0 38640.0 6860.0 38505.0 ;
      RECT  6985.0 38640.0 7050.0 38505.0 ;
      RECT  6985.0 38640.0 7050.0 38505.0 ;
      RECT  6795.0 38640.0 6860.0 38505.0 ;
      RECT  7155.0 37665.0 7220.0 37530.0 ;
      RECT  7155.0 38640.0 7220.0 38505.0 ;
      RECT  6852.5 38197.5 6917.5 38062.5 ;
      RECT  6852.5 38197.5 6917.5 38062.5 ;
      RECT  7017.5 38162.5 7082.5 38097.5 ;
      RECT  6727.5 37445.0 7287.5 37380.0 ;
      RECT  6727.5 38790.0 7287.5 38725.0 ;
      RECT  4990.0 38062.5 5055.0 38197.5 ;
      RECT  5130.0 38335.0 5195.0 38470.0 ;
      RECT  6125.0 38300.0 5990.0 38365.0 ;
      RECT  5675.0 39917.5 5740.0 40102.5 ;
      RECT  5675.0 38757.5 5740.0 38942.5 ;
      RECT  5315.0 38875.0 5380.0 38725.0 ;
      RECT  5315.0 39760.0 5380.0 40135.0 ;
      RECT  5505.0 38875.0 5570.0 39760.0 ;
      RECT  5315.0 39760.0 5380.0 39895.0 ;
      RECT  5505.0 39760.0 5570.0 39895.0 ;
      RECT  5505.0 39760.0 5570.0 39895.0 ;
      RECT  5315.0 39760.0 5380.0 39895.0 ;
      RECT  5315.0 38875.0 5380.0 39010.0 ;
      RECT  5505.0 38875.0 5570.0 39010.0 ;
      RECT  5505.0 38875.0 5570.0 39010.0 ;
      RECT  5315.0 38875.0 5380.0 39010.0 ;
      RECT  5675.0 39850.0 5740.0 39985.0 ;
      RECT  5675.0 38875.0 5740.0 39010.0 ;
      RECT  5372.5 39317.5 5437.5 39452.5 ;
      RECT  5372.5 39317.5 5437.5 39452.5 ;
      RECT  5537.5 39352.5 5602.5 39417.5 ;
      RECT  5247.5 40070.0 5807.5 40135.0 ;
      RECT  5247.5 38725.0 5807.5 38790.0 ;
      RECT  5875.0 38920.0 5940.0 38725.0 ;
      RECT  5875.0 39760.0 5940.0 40135.0 ;
      RECT  6255.0 39760.0 6320.0 40135.0 ;
      RECT  6425.0 39917.5 6490.0 40102.5 ;
      RECT  6425.0 38757.5 6490.0 38942.5 ;
      RECT  5875.0 39760.0 5940.0 39895.0 ;
      RECT  6065.0 39760.0 6130.0 39895.0 ;
      RECT  6065.0 39760.0 6130.0 39895.0 ;
      RECT  5875.0 39760.0 5940.0 39895.0 ;
      RECT  6065.0 39760.0 6130.0 39895.0 ;
      RECT  6255.0 39760.0 6320.0 39895.0 ;
      RECT  6255.0 39760.0 6320.0 39895.0 ;
      RECT  6065.0 39760.0 6130.0 39895.0 ;
      RECT  5875.0 38920.0 5940.0 39055.0 ;
      RECT  6065.0 38920.0 6130.0 39055.0 ;
      RECT  6065.0 38920.0 6130.0 39055.0 ;
      RECT  5875.0 38920.0 5940.0 39055.0 ;
      RECT  6065.0 38920.0 6130.0 39055.0 ;
      RECT  6255.0 38920.0 6320.0 39055.0 ;
      RECT  6255.0 38920.0 6320.0 39055.0 ;
      RECT  6065.0 38920.0 6130.0 39055.0 ;
      RECT  6425.0 39850.0 6490.0 39985.0 ;
      RECT  6425.0 38875.0 6490.0 39010.0 ;
      RECT  6260.0 39150.0 6125.0 39215.0 ;
      RECT  6002.5 39365.0 5867.5 39430.0 ;
      RECT  6065.0 39760.0 6130.0 39895.0 ;
      RECT  6255.0 38920.0 6320.0 39055.0 ;
      RECT  6355.0 39365.0 6220.0 39430.0 ;
      RECT  5867.5 39365.0 6002.5 39430.0 ;
      RECT  6125.0 39150.0 6260.0 39215.0 ;
      RECT  6220.0 39365.0 6355.0 39430.0 ;
      RECT  5807.5 40070.0 6727.5 40135.0 ;
      RECT  5807.5 38725.0 6727.5 38790.0 ;
      RECT  7155.0 39917.5 7220.0 40102.5 ;
      RECT  7155.0 38757.5 7220.0 38942.5 ;
      RECT  6795.0 38875.0 6860.0 38725.0 ;
      RECT  6795.0 39760.0 6860.0 40135.0 ;
      RECT  6985.0 38875.0 7050.0 39760.0 ;
      RECT  6795.0 39760.0 6860.0 39895.0 ;
      RECT  6985.0 39760.0 7050.0 39895.0 ;
      RECT  6985.0 39760.0 7050.0 39895.0 ;
      RECT  6795.0 39760.0 6860.0 39895.0 ;
      RECT  6795.0 38875.0 6860.0 39010.0 ;
      RECT  6985.0 38875.0 7050.0 39010.0 ;
      RECT  6985.0 38875.0 7050.0 39010.0 ;
      RECT  6795.0 38875.0 6860.0 39010.0 ;
      RECT  7155.0 39850.0 7220.0 39985.0 ;
      RECT  7155.0 38875.0 7220.0 39010.0 ;
      RECT  6852.5 39317.5 6917.5 39452.5 ;
      RECT  6852.5 39317.5 6917.5 39452.5 ;
      RECT  7017.5 39352.5 7082.5 39417.5 ;
      RECT  6727.5 40070.0 7287.5 40135.0 ;
      RECT  6727.5 38725.0 7287.5 38790.0 ;
      RECT  4990.0 39317.5 5055.0 39452.5 ;
      RECT  5130.0 39045.0 5195.0 39180.0 ;
      RECT  6125.0 39150.0 5990.0 39215.0 ;
      RECT  5675.0 40287.5 5740.0 40102.5 ;
      RECT  5675.0 41447.5 5740.0 41262.5 ;
      RECT  5315.0 41330.0 5380.0 41480.0 ;
      RECT  5315.0 40445.0 5380.0 40070.0 ;
      RECT  5505.0 41330.0 5570.0 40445.0 ;
      RECT  5315.0 40445.0 5380.0 40310.0 ;
      RECT  5505.0 40445.0 5570.0 40310.0 ;
      RECT  5505.0 40445.0 5570.0 40310.0 ;
      RECT  5315.0 40445.0 5380.0 40310.0 ;
      RECT  5315.0 41330.0 5380.0 41195.0 ;
      RECT  5505.0 41330.0 5570.0 41195.0 ;
      RECT  5505.0 41330.0 5570.0 41195.0 ;
      RECT  5315.0 41330.0 5380.0 41195.0 ;
      RECT  5675.0 40355.0 5740.0 40220.0 ;
      RECT  5675.0 41330.0 5740.0 41195.0 ;
      RECT  5372.5 40887.5 5437.5 40752.5 ;
      RECT  5372.5 40887.5 5437.5 40752.5 ;
      RECT  5537.5 40852.5 5602.5 40787.5 ;
      RECT  5247.5 40135.0 5807.5 40070.0 ;
      RECT  5247.5 41480.0 5807.5 41415.0 ;
      RECT  5875.0 41285.0 5940.0 41480.0 ;
      RECT  5875.0 40445.0 5940.0 40070.0 ;
      RECT  6255.0 40445.0 6320.0 40070.0 ;
      RECT  6425.0 40287.5 6490.0 40102.5 ;
      RECT  6425.0 41447.5 6490.0 41262.5 ;
      RECT  5875.0 40445.0 5940.0 40310.0 ;
      RECT  6065.0 40445.0 6130.0 40310.0 ;
      RECT  6065.0 40445.0 6130.0 40310.0 ;
      RECT  5875.0 40445.0 5940.0 40310.0 ;
      RECT  6065.0 40445.0 6130.0 40310.0 ;
      RECT  6255.0 40445.0 6320.0 40310.0 ;
      RECT  6255.0 40445.0 6320.0 40310.0 ;
      RECT  6065.0 40445.0 6130.0 40310.0 ;
      RECT  5875.0 41285.0 5940.0 41150.0 ;
      RECT  6065.0 41285.0 6130.0 41150.0 ;
      RECT  6065.0 41285.0 6130.0 41150.0 ;
      RECT  5875.0 41285.0 5940.0 41150.0 ;
      RECT  6065.0 41285.0 6130.0 41150.0 ;
      RECT  6255.0 41285.0 6320.0 41150.0 ;
      RECT  6255.0 41285.0 6320.0 41150.0 ;
      RECT  6065.0 41285.0 6130.0 41150.0 ;
      RECT  6425.0 40355.0 6490.0 40220.0 ;
      RECT  6425.0 41330.0 6490.0 41195.0 ;
      RECT  6260.0 41055.0 6125.0 40990.0 ;
      RECT  6002.5 40840.0 5867.5 40775.0 ;
      RECT  6065.0 40445.0 6130.0 40310.0 ;
      RECT  6255.0 41285.0 6320.0 41150.0 ;
      RECT  6355.0 40840.0 6220.0 40775.0 ;
      RECT  5867.5 40840.0 6002.5 40775.0 ;
      RECT  6125.0 41055.0 6260.0 40990.0 ;
      RECT  6220.0 40840.0 6355.0 40775.0 ;
      RECT  5807.5 40135.0 6727.5 40070.0 ;
      RECT  5807.5 41480.0 6727.5 41415.0 ;
      RECT  7155.0 40287.5 7220.0 40102.5 ;
      RECT  7155.0 41447.5 7220.0 41262.5 ;
      RECT  6795.0 41330.0 6860.0 41480.0 ;
      RECT  6795.0 40445.0 6860.0 40070.0 ;
      RECT  6985.0 41330.0 7050.0 40445.0 ;
      RECT  6795.0 40445.0 6860.0 40310.0 ;
      RECT  6985.0 40445.0 7050.0 40310.0 ;
      RECT  6985.0 40445.0 7050.0 40310.0 ;
      RECT  6795.0 40445.0 6860.0 40310.0 ;
      RECT  6795.0 41330.0 6860.0 41195.0 ;
      RECT  6985.0 41330.0 7050.0 41195.0 ;
      RECT  6985.0 41330.0 7050.0 41195.0 ;
      RECT  6795.0 41330.0 6860.0 41195.0 ;
      RECT  7155.0 40355.0 7220.0 40220.0 ;
      RECT  7155.0 41330.0 7220.0 41195.0 ;
      RECT  6852.5 40887.5 6917.5 40752.5 ;
      RECT  6852.5 40887.5 6917.5 40752.5 ;
      RECT  7017.5 40852.5 7082.5 40787.5 ;
      RECT  6727.5 40135.0 7287.5 40070.0 ;
      RECT  6727.5 41480.0 7287.5 41415.0 ;
      RECT  4990.0 40752.5 5055.0 40887.5 ;
      RECT  5130.0 41025.0 5195.0 41160.0 ;
      RECT  6125.0 40990.0 5990.0 41055.0 ;
      RECT  4792.5 20250.0 5162.5 20315.0 ;
      RECT  4792.5 22230.0 5162.5 22295.0 ;
      RECT  4792.5 22940.0 5162.5 23005.0 ;
      RECT  4792.5 24920.0 5162.5 24985.0 ;
      RECT  4792.5 25630.0 5162.5 25695.0 ;
      RECT  4792.5 27610.0 5162.5 27675.0 ;
      RECT  4792.5 28320.0 5162.5 28385.0 ;
      RECT  4792.5 30300.0 5162.5 30365.0 ;
      RECT  4792.5 31010.0 5162.5 31075.0 ;
      RECT  4792.5 32990.0 5162.5 33055.0 ;
      RECT  4792.5 33700.0 5162.5 33765.0 ;
      RECT  4792.5 35680.0 5162.5 35745.0 ;
      RECT  4792.5 36390.0 5162.5 36455.0 ;
      RECT  4792.5 38370.0 5162.5 38435.0 ;
      RECT  4792.5 39080.0 5162.5 39145.0 ;
      RECT  4792.5 41060.0 5162.5 41125.0 ;
      RECT  7017.5 20522.5 7082.5 20587.5 ;
      RECT  7017.5 21957.5 7082.5 22022.5 ;
      RECT  7017.5 23212.5 7082.5 23277.5 ;
      RECT  7017.5 24647.5 7082.5 24712.5 ;
      RECT  7017.5 25902.5 7082.5 25967.5 ;
      RECT  7017.5 27337.5 7082.5 27402.5 ;
      RECT  7017.5 28592.5 7082.5 28657.5 ;
      RECT  7017.5 30027.5 7082.5 30092.5 ;
      RECT  7017.5 31282.5 7082.5 31347.5 ;
      RECT  7017.5 32717.5 7082.5 32782.5 ;
      RECT  7017.5 33972.5 7082.5 34037.5 ;
      RECT  7017.5 35407.5 7082.5 35472.5 ;
      RECT  7017.5 36662.5 7082.5 36727.5 ;
      RECT  7017.5 38097.5 7082.5 38162.5 ;
      RECT  7017.5 39352.5 7082.5 39417.5 ;
      RECT  7017.5 40787.5 7082.5 40852.5 ;
      RECT  4792.5 21240.0 5247.5 21305.0 ;
      RECT  4792.5 23930.0 5247.5 23995.0 ;
      RECT  4792.5 26620.0 5247.5 26685.0 ;
      RECT  4792.5 29310.0 5247.5 29375.0 ;
      RECT  4792.5 32000.0 5247.5 32065.0 ;
      RECT  4792.5 34690.0 5247.5 34755.0 ;
      RECT  4792.5 37380.0 5247.5 37445.0 ;
      RECT  4792.5 40070.0 5247.5 40135.0 ;
      RECT  4792.5 19895.0 5247.5 19960.0 ;
      RECT  4792.5 22585.0 5247.5 22650.0 ;
      RECT  4792.5 25275.0 5247.5 25340.0 ;
      RECT  4792.5 27965.0 5247.5 28030.0 ;
      RECT  4792.5 30655.0 5247.5 30720.0 ;
      RECT  4792.5 33345.0 5247.5 33410.0 ;
      RECT  4792.5 36035.0 5247.5 36100.0 ;
      RECT  4792.5 38725.0 5247.5 38790.0 ;
      RECT  4792.5 41415.0 5247.5 41480.0 ;
      RECT  837.5 8757.5 7277.5 8052.5 ;
      RECT  837.5 7347.5 7277.5 8052.5 ;
      RECT  837.5 7347.5 7277.5 6642.5 ;
      RECT  837.5 5937.5 7277.5 6642.5 ;
      RECT  1042.5 8757.5 1107.5 5937.5 ;
      RECT  4047.5 8757.5 4112.5 5937.5 ;
      RECT  7007.5 8757.5 7072.5 5937.5 ;
      RECT  2057.5 8757.5 2122.5 5937.5 ;
      RECT  5017.5 8757.5 5082.5 5937.5 ;
      RECT  1202.5 8757.5 1267.5 5937.5 ;
      RECT  35.0 -3.5527136788e-12 380.0 415.0 ;
      RECT  35.0 43302.5 380.0 43717.5 ;
      RECT  11515.0 -3.5527136788e-12 11860.0 415.0 ;
      RECT  11515.0 43302.5 11860.0 43717.5 ;
      RECT  420.0 385.0 765.0 800.0 ;
      RECT  420.0 43687.5 765.0 44102.5 ;
      RECT  11900.0 385.0 12245.0 800.0 ;
      RECT  11900.0 43687.5 12245.0 44102.5 ;
      RECT  7277.5 9340.0 7142.5 9405.0 ;
      RECT  7687.5 9340.0 7552.5 9405.0 ;
      RECT  7002.5 10685.0 6867.5 10750.0 ;
      RECT  7892.5 10685.0 7757.5 10750.0 ;
      RECT  7277.5 14720.0 7142.5 14785.0 ;
      RECT  8097.5 14720.0 7962.5 14785.0 ;
      RECT  7002.5 16065.0 6867.5 16130.0 ;
      RECT  8302.5 16065.0 8167.5 16130.0 ;
      RECT  415.0 9135.0 -8.881784197e-13 9200.0 ;
      RECT  415.0 11825.0 -8.881784197e-13 11890.0 ;
      RECT  415.0 14515.0 -8.881784197e-13 14580.0 ;
      RECT  415.0 17205.0 -8.881784197e-13 17270.0 ;
      RECT  800.0 10480.0 385.0 10545.0 ;
      RECT  800.0 13170.0 385.0 13235.0 ;
      RECT  800.0 15860.0 385.0 15925.0 ;
      RECT  800.0 18550.0 385.0 18615.0 ;
      RECT  7345.0 8372.5 7210.0 8437.5 ;
      RECT  7687.5 8372.5 7552.5 8437.5 ;
      RECT  7345.0 7667.5 7210.0 7732.5 ;
      RECT  7892.5 7667.5 7757.5 7732.5 ;
      RECT  7345.0 6962.5 7210.0 7027.5 ;
      RECT  8097.5 6962.5 7962.5 7027.5 ;
      RECT  7345.0 6257.5 7210.0 6322.5 ;
      RECT  8302.5 6257.5 8167.5 6322.5 ;
      RECT  972.5 8725.0 837.5 8790.0 ;
      RECT  415.0 8725.0 -8.881784197e-13 8790.0 ;
      RECT  972.5 8020.0 837.5 8085.0 ;
      RECT  415.0 8020.0 -8.881784197e-13 8085.0 ;
      RECT  972.5 7315.0 837.5 7380.0 ;
      RECT  415.0 7315.0 -8.881784197e-13 7380.0 ;
      RECT  972.5 6610.0 837.5 6675.0 ;
      RECT  415.0 6610.0 -8.881784197e-13 6675.0 ;
      RECT  972.5 5905.0 837.5 5970.0 ;
      RECT  415.0 5905.0 -8.881784197e-13 5970.0 ;
      RECT  800.0 5700.0 385.0 5765.0 ;
      RECT  800.0 5700.0 385.0 5765.0 ;
      RECT  800.0 5700.0 385.0 5765.0 ;
      RECT  800.0 5700.0 385.0 5765.0 ;
      RECT  9122.5 4632.5 8987.5 4697.5 ;
      RECT  8712.5 2447.5 8577.5 2512.5 ;
      RECT  8917.5 3995.0 8782.5 4060.0 ;
      RECT  9122.5 42425.0 8987.5 42490.0 ;
      RECT  9327.5 11135.0 9192.5 11200.0 ;
      RECT  9532.5 15160.0 9397.5 15225.0 ;
      RECT  8507.5 8930.0 8372.5 8995.0 ;
      RECT  5090.0 41620.0 4955.0 41685.0 ;
      RECT  8507.5 41620.0 8372.5 41685.0 ;
      RECT  12280.0 43110.0 11865.0 43175.0 ;
      RECT  12280.0 19732.5 11865.0 19797.5 ;
      RECT  12280.0 11265.0 11865.0 11330.0 ;
      RECT  12280.0 7637.5 11865.0 7702.5 ;
      RECT  12280.0 10597.5 11865.0 10662.5 ;
      RECT  12280.0 5647.5 11865.0 5712.5 ;
      RECT  12280.0 8607.5 11865.0 8672.5 ;
      RECT  12280.0 2577.5 11865.0 2642.5 ;
      RECT  800.0 21240.0 385.0 21305.0 ;
      RECT  12280.0 21240.0 11865.0 21305.0 ;
      RECT  800.0 23930.0 385.0 23995.0 ;
      RECT  12280.0 23930.0 11865.0 23995.0 ;
      RECT  800.0 26620.0 385.0 26685.0 ;
      RECT  12280.0 26620.0 11865.0 26685.0 ;
      RECT  800.0 29310.0 385.0 29375.0 ;
      RECT  12280.0 29310.0 11865.0 29375.0 ;
      RECT  800.0 32000.0 385.0 32065.0 ;
      RECT  12280.0 32000.0 11865.0 32065.0 ;
      RECT  800.0 34690.0 385.0 34755.0 ;
      RECT  12280.0 34690.0 11865.0 34755.0 ;
      RECT  800.0 37380.0 385.0 37445.0 ;
      RECT  12280.0 37380.0 11865.0 37445.0 ;
      RECT  800.0 40070.0 385.0 40135.0 ;
      RECT  12280.0 40070.0 11865.0 40135.0 ;
      RECT  11895.0 3865.0 11480.0 3930.0 ;
      RECT  11895.0 15290.0 11480.0 15355.0 ;
      RECT  11895.0 4792.5 11480.0 4857.5 ;
      RECT  11895.0 12067.5 11480.0 12132.5 ;
      RECT  415.0 19895.0 -8.881784197e-13 19960.0 ;
      RECT  415.0 22585.0 -8.881784197e-13 22650.0 ;
      RECT  415.0 25275.0 -8.881784197e-13 25340.0 ;
      RECT  415.0 27965.0 -8.881784197e-13 28030.0 ;
      RECT  415.0 30655.0 -8.881784197e-13 30720.0 ;
      RECT  415.0 33345.0 -8.881784197e-13 33410.0 ;
      RECT  415.0 36035.0 -8.881784197e-13 36100.0 ;
      RECT  415.0 38725.0 -8.881784197e-13 38790.0 ;
      RECT  415.0 41415.0 -8.881784197e-13 41480.0 ;
      RECT  67.5 452.5 12212.5 732.5 ;
      RECT  67.5 43755.0 12212.5 44035.0 ;
      RECT  67.5 67.5 12212.5 347.5 ;
      RECT  67.5 43370.0 12212.5 43650.0 ;
      RECT  -720.0 24047.5 -785.0 24112.5 ;
      RECT  -752.5 24047.5 -767.5 24112.5 ;
      RECT  -720.0 24080.0 -785.0 24665.0 ;
      RECT  -720.0 25210.0 -785.0 25605.0 ;
      RECT  -720.0 26530.0 -785.0 27115.0 ;
      RECT  -1517.5 26967.5 -1895.0 27032.5 ;
      RECT  -1517.5 29927.5 -1895.0 29992.5 ;
      RECT  -1517.5 24977.5 -1895.0 25042.5 ;
      RECT  -1517.5 27937.5 -1895.0 28002.5 ;
      RECT  -735.0 24047.5 -800.0 24112.5 ;
      RECT  -720.0 25177.5 -785.0 25242.5 ;
      RECT  -2170.0 35862.5 -2235.0 36627.5 ;
      RECT  -720.0 29212.5 -785.0 30642.5 ;
      RECT  -1690.0 23962.5 -1895.0 24027.5 ;
      RECT  -2212.5 30642.5 -2277.5 32580.0 ;
      RECT  -2427.5 31052.5 -2492.5 32837.5 ;
      RECT  -795.0 32077.5 -860.0 32647.5 ;
      RECT  -655.0 31872.5 -720.0 32837.5 ;
      RECT  -515.0 31257.5 -580.0 33027.5 ;
      RECT  -795.0 33587.5 -860.0 33652.5 ;
      RECT  -795.0 33122.5 -860.0 33620.0 ;
      RECT  -767.5 33587.5 -827.5 33652.5 ;
      RECT  -700.0 33752.5 -765.0 33817.5 ;
      RECT  -732.5 33752.5 -767.5 33817.5 ;
      RECT  -700.0 33785.0 -765.0 37325.0 ;
      RECT  -3485.0 32077.5 -3550.0 33207.5 ;
      RECT  -3345.0 31257.5 -3410.0 33397.5 ;
      RECT  -3205.0 31462.5 -3270.0 33587.5 ;
      RECT  -3485.0 34147.5 -3550.0 34212.5 ;
      RECT  -3485.0 33682.5 -3550.0 34180.0 ;
      RECT  -3457.5 34147.5 -3517.5 34212.5 ;
      RECT  -3425.0 34345.0 -3490.0 34740.0 ;
      RECT  -3425.0 34905.0 -3490.0 35300.0 ;
      RECT  -2170.0 35830.0 -2235.0 35895.0 ;
      RECT  -2202.5 35830.0 -2235.0 35895.0 ;
      RECT  -2170.0 35737.5 -2235.0 35862.5 ;
      RECT  -2170.0 35145.0 -2235.0 35540.0 ;
      RECT  -2212.5 33002.5 -2277.5 33372.5 ;
      RECT  -2157.5 34077.5 -2222.5 34517.5 ;
      RECT  -3425.0 35465.0 -3490.0 35702.5 ;
      RECT  -2170.0 34742.5 -2235.0 34980.0 ;
      RECT  -107.5 23757.5 -172.5 35862.5 ;
      RECT  -107.5 30847.5 -172.5 32452.5 ;
      RECT  -1452.5 23757.5 -1517.5 35862.5 ;
      RECT  -1452.5 31667.5 -1517.5 32452.5 ;
      RECT  -2797.5 32452.5 -2862.5 35862.5 ;
      RECT  -2797.5 30847.5 -2862.5 32452.5 ;
      RECT  -4142.5 32452.5 -4207.5 35862.5 ;
      RECT  -4142.5 31667.5 -4207.5 32452.5 ;
      RECT  -4142.5 35830.0 -4207.5 35895.0 ;
      RECT  -4142.5 35657.5 -4207.5 35862.5 ;
      RECT  -4175.0 35830.0 -4220.0 35895.0 ;
      RECT  -4010.0 23757.5 -3305.0 30197.5 ;
      RECT  -2600.0 23757.5 -3305.0 30197.5 ;
      RECT  -2600.0 23757.5 -1895.0 30197.5 ;
      RECT  -4010.0 23962.5 -1895.0 24027.5 ;
      RECT  -4010.0 26967.5 -1895.0 27032.5 ;
      RECT  -4010.0 29927.5 -1895.0 29992.5 ;
      RECT  -4010.0 24977.5 -1895.0 25042.5 ;
      RECT  -4010.0 27937.5 -1895.0 28002.5 ;
      RECT  -4010.0 24122.5 -1895.0 24187.5 ;
      RECT  -1300.0 24375.0 -1485.0 24440.0 ;
      RECT  -140.0 24375.0 -325.0 24440.0 ;
      RECT  -1342.5 23825.0 -1517.5 24270.0 ;
      RECT  -257.5 24015.0 -1142.5 24080.0 ;
      RECT  -1210.0 23825.0 -1375.0 23890.0 ;
      RECT  -1210.0 24205.0 -1375.0 24270.0 ;
      RECT  -1142.5 23825.0 -1277.5 23890.0 ;
      RECT  -1142.5 24205.0 -1277.5 24270.0 ;
      RECT  -1142.5 24015.0 -1277.5 24080.0 ;
      RECT  -1142.5 24015.0 -1277.5 24080.0 ;
      RECT  -1342.5 23825.0 -1407.5 24270.0 ;
      RECT  -160.0 23825.0 -325.0 23890.0 ;
      RECT  -160.0 24205.0 -325.0 24270.0 ;
      RECT  -257.5 23825.0 -392.5 23890.0 ;
      RECT  -257.5 24205.0 -392.5 24270.0 ;
      RECT  -257.5 24015.0 -392.5 24080.0 ;
      RECT  -257.5 24015.0 -392.5 24080.0 ;
      RECT  -127.5 23825.0 -192.5 24270.0 ;
      RECT  -1232.5 24375.0 -1367.5 24440.0 ;
      RECT  -257.5 24375.0 -392.5 24440.0 ;
      RECT  -700.0 23882.5 -835.0 23947.5 ;
      RECT  -700.0 23882.5 -835.0 23947.5 ;
      RECT  -735.0 24047.5 -800.0 24112.5 ;
      RECT  -1452.5 23757.5 -1517.5 24507.5 ;
      RECT  -107.5 23757.5 -172.5 24507.5 ;
      RECT  -1300.0 25315.0 -1485.0 25380.0 ;
      RECT  -140.0 25315.0 -325.0 25380.0 ;
      RECT  -1297.5 24575.0 -1517.5 25020.0 ;
      RECT  -472.5 25145.0 -967.5 25210.0 ;
      RECT  -1165.0 24575.0 -1330.0 24640.0 ;
      RECT  -1165.0 24955.0 -1330.0 25020.0 ;
      RECT  -1000.0 24765.0 -1165.0 24830.0 ;
      RECT  -1000.0 25145.0 -1165.0 25210.0 ;
      RECT  -1097.5 24575.0 -1232.5 24640.0 ;
      RECT  -1097.5 24955.0 -1232.5 25020.0 ;
      RECT  -1097.5 24765.0 -1232.5 24830.0 ;
      RECT  -1097.5 25145.0 -1232.5 25210.0 ;
      RECT  -967.5 24765.0 -1032.5 25210.0 ;
      RECT  -1297.5 24575.0 -1362.5 25020.0 ;
      RECT  -175.0 24575.0 -340.0 24640.0 ;
      RECT  -175.0 24955.0 -340.0 25020.0 ;
      RECT  -340.0 24765.0 -505.0 24830.0 ;
      RECT  -340.0 25145.0 -505.0 25210.0 ;
      RECT  -272.5 24575.0 -407.5 24640.0 ;
      RECT  -272.5 24955.0 -407.5 25020.0 ;
      RECT  -272.5 24765.0 -407.5 24830.0 ;
      RECT  -272.5 25145.0 -407.5 25210.0 ;
      RECT  -472.5 24765.0 -537.5 25210.0 ;
      RECT  -142.5 24575.0 -207.5 25020.0 ;
      RECT  -1232.5 25315.0 -1367.5 25380.0 ;
      RECT  -257.5 25315.0 -392.5 25380.0 ;
      RECT  -685.0 24632.5 -820.0 24697.5 ;
      RECT  -685.0 24632.5 -820.0 24697.5 ;
      RECT  -720.0 25177.5 -785.0 25242.5 ;
      RECT  -1452.5 24507.5 -1517.5 25447.5 ;
      RECT  -107.5 24507.5 -172.5 25447.5 ;
      RECT  -1300.0 26825.0 -1485.0 26890.0 ;
      RECT  -140.0 26825.0 -325.0 26890.0 ;
      RECT  -1297.5 25515.0 -1517.5 26720.0 ;
      RECT  -472.5 26465.0 -967.5 26530.0 ;
      RECT  -1165.0 25515.0 -1330.0 25580.0 ;
      RECT  -1165.0 25895.0 -1330.0 25960.0 ;
      RECT  -1165.0 26275.0 -1330.0 26340.0 ;
      RECT  -1165.0 26655.0 -1330.0 26720.0 ;
      RECT  -1000.0 25705.0 -1165.0 25770.0 ;
      RECT  -1000.0 26085.0 -1165.0 26150.0 ;
      RECT  -1000.0 26465.0 -1165.0 26530.0 ;
      RECT  -1097.5 25515.0 -1232.5 25580.0 ;
      RECT  -1097.5 25895.0 -1232.5 25960.0 ;
      RECT  -1097.5 26275.0 -1232.5 26340.0 ;
      RECT  -1097.5 26655.0 -1232.5 26720.0 ;
      RECT  -1097.5 25705.0 -1232.5 25770.0 ;
      RECT  -1097.5 26085.0 -1232.5 26150.0 ;
      RECT  -1097.5 26465.0 -1232.5 26530.0 ;
      RECT  -967.5 25705.0 -1032.5 26530.0 ;
      RECT  -1297.5 25515.0 -1362.5 26720.0 ;
      RECT  -175.0 25515.0 -340.0 25580.0 ;
      RECT  -175.0 25895.0 -340.0 25960.0 ;
      RECT  -175.0 26275.0 -340.0 26340.0 ;
      RECT  -175.0 26655.0 -340.0 26720.0 ;
      RECT  -340.0 25705.0 -505.0 25770.0 ;
      RECT  -340.0 26085.0 -505.0 26150.0 ;
      RECT  -340.0 26465.0 -505.0 26530.0 ;
      RECT  -272.5 25515.0 -407.5 25580.0 ;
      RECT  -272.5 25895.0 -407.5 25960.0 ;
      RECT  -272.5 26275.0 -407.5 26340.0 ;
      RECT  -272.5 26655.0 -407.5 26720.0 ;
      RECT  -272.5 25705.0 -407.5 25770.0 ;
      RECT  -272.5 26085.0 -407.5 26150.0 ;
      RECT  -272.5 26465.0 -407.5 26530.0 ;
      RECT  -472.5 25705.0 -537.5 26530.0 ;
      RECT  -142.5 25515.0 -207.5 26720.0 ;
      RECT  -1232.5 26825.0 -1367.5 26890.0 ;
      RECT  -257.5 26825.0 -392.5 26890.0 ;
      RECT  -685.0 25572.5 -820.0 25637.5 ;
      RECT  -685.0 25572.5 -820.0 25637.5 ;
      RECT  -720.0 26497.5 -785.0 26562.5 ;
      RECT  -1452.5 25447.5 -1517.5 26957.5 ;
      RECT  -107.5 25447.5 -172.5 26957.5 ;
      RECT  -1300.0 29475.0 -1485.0 29540.0 ;
      RECT  -140.0 29475.0 -325.0 29540.0 ;
      RECT  -1297.5 27025.0 -1517.5 29370.0 ;
      RECT  -472.5 29115.0 -967.5 29180.0 ;
      RECT  -1165.0 27025.0 -1330.0 27090.0 ;
      RECT  -1165.0 27405.0 -1330.0 27470.0 ;
      RECT  -1165.0 27785.0 -1330.0 27850.0 ;
      RECT  -1165.0 28165.0 -1330.0 28230.0 ;
      RECT  -1165.0 28545.0 -1330.0 28610.0 ;
      RECT  -1165.0 28925.0 -1330.0 28990.0 ;
      RECT  -1165.0 29305.0 -1330.0 29370.0 ;
      RECT  -1000.0 27215.0 -1165.0 27280.0 ;
      RECT  -1000.0 27595.0 -1165.0 27660.0 ;
      RECT  -1000.0 27975.0 -1165.0 28040.0 ;
      RECT  -1000.0 28355.0 -1165.0 28420.0 ;
      RECT  -1000.0 28735.0 -1165.0 28800.0 ;
      RECT  -1000.0 29115.0 -1165.0 29180.0 ;
      RECT  -1097.5 27025.0 -1232.5 27090.0 ;
      RECT  -1097.5 27405.0 -1232.5 27470.0 ;
      RECT  -1097.5 27785.0 -1232.5 27850.0 ;
      RECT  -1097.5 28165.0 -1232.5 28230.0 ;
      RECT  -1097.5 28545.0 -1232.5 28610.0 ;
      RECT  -1097.5 28925.0 -1232.5 28990.0 ;
      RECT  -1097.5 29305.0 -1232.5 29370.0 ;
      RECT  -1097.5 27215.0 -1232.5 27280.0 ;
      RECT  -1097.5 27595.0 -1232.5 27660.0 ;
      RECT  -1097.5 27975.0 -1232.5 28040.0 ;
      RECT  -1097.5 28355.0 -1232.5 28420.0 ;
      RECT  -1097.5 28735.0 -1232.5 28800.0 ;
      RECT  -1097.5 29115.0 -1232.5 29180.0 ;
      RECT  -967.5 27215.0 -1032.5 29180.0 ;
      RECT  -1297.5 27025.0 -1362.5 29370.0 ;
      RECT  -175.0 27025.0 -340.0 27090.0 ;
      RECT  -175.0 27405.0 -340.0 27470.0 ;
      RECT  -175.0 27785.0 -340.0 27850.0 ;
      RECT  -175.0 28165.0 -340.0 28230.0 ;
      RECT  -175.0 28545.0 -340.0 28610.0 ;
      RECT  -175.0 28925.0 -340.0 28990.0 ;
      RECT  -175.0 29305.0 -340.0 29370.0 ;
      RECT  -340.0 27215.0 -505.0 27280.0 ;
      RECT  -340.0 27595.0 -505.0 27660.0 ;
      RECT  -340.0 27975.0 -505.0 28040.0 ;
      RECT  -340.0 28355.0 -505.0 28420.0 ;
      RECT  -340.0 28735.0 -505.0 28800.0 ;
      RECT  -340.0 29115.0 -505.0 29180.0 ;
      RECT  -272.5 27025.0 -407.5 27090.0 ;
      RECT  -272.5 27405.0 -407.5 27470.0 ;
      RECT  -272.5 27785.0 -407.5 27850.0 ;
      RECT  -272.5 28165.0 -407.5 28230.0 ;
      RECT  -272.5 28545.0 -407.5 28610.0 ;
      RECT  -272.5 28925.0 -407.5 28990.0 ;
      RECT  -272.5 29305.0 -407.5 29370.0 ;
      RECT  -272.5 27215.0 -407.5 27280.0 ;
      RECT  -272.5 27595.0 -407.5 27660.0 ;
      RECT  -272.5 27975.0 -407.5 28040.0 ;
      RECT  -272.5 28355.0 -407.5 28420.0 ;
      RECT  -272.5 28735.0 -407.5 28800.0 ;
      RECT  -272.5 29115.0 -407.5 29180.0 ;
      RECT  -472.5 27215.0 -537.5 29180.0 ;
      RECT  -142.5 27025.0 -207.5 29370.0 ;
      RECT  -1232.5 29475.0 -1367.5 29540.0 ;
      RECT  -257.5 29475.0 -392.5 29540.0 ;
      RECT  -685.0 27082.5 -820.0 27147.5 ;
      RECT  -685.0 27082.5 -820.0 27147.5 ;
      RECT  -720.0 29147.5 -785.0 29212.5 ;
      RECT  -1452.5 26957.5 -1517.5 29607.5 ;
      RECT  -107.5 26957.5 -172.5 29607.5 ;
      RECT  -302.5 32520.0 -107.5 32585.0 ;
      RECT  -1142.5 32520.0 -1517.5 32585.0 ;
      RECT  -1142.5 32900.0 -1517.5 32965.0 ;
      RECT  -1300.0 33260.0 -1485.0 33325.0 ;
      RECT  -140.0 33260.0 -325.0 33325.0 ;
      RECT  -1142.5 32520.0 -1277.5 32585.0 ;
      RECT  -1142.5 32710.0 -1277.5 32775.0 ;
      RECT  -1142.5 32710.0 -1277.5 32775.0 ;
      RECT  -1142.5 32520.0 -1277.5 32585.0 ;
      RECT  -1142.5 32710.0 -1277.5 32775.0 ;
      RECT  -1142.5 32900.0 -1277.5 32965.0 ;
      RECT  -1142.5 32900.0 -1277.5 32965.0 ;
      RECT  -1142.5 32710.0 -1277.5 32775.0 ;
      RECT  -1142.5 32900.0 -1277.5 32965.0 ;
      RECT  -1142.5 33090.0 -1277.5 33155.0 ;
      RECT  -1142.5 33090.0 -1277.5 33155.0 ;
      RECT  -1142.5 32900.0 -1277.5 32965.0 ;
      RECT  -302.5 32520.0 -437.5 32585.0 ;
      RECT  -302.5 32710.0 -437.5 32775.0 ;
      RECT  -302.5 32710.0 -437.5 32775.0 ;
      RECT  -302.5 32520.0 -437.5 32585.0 ;
      RECT  -302.5 32710.0 -437.5 32775.0 ;
      RECT  -302.5 32900.0 -437.5 32965.0 ;
      RECT  -302.5 32900.0 -437.5 32965.0 ;
      RECT  -302.5 32710.0 -437.5 32775.0 ;
      RECT  -302.5 32900.0 -437.5 32965.0 ;
      RECT  -302.5 33090.0 -437.5 33155.0 ;
      RECT  -302.5 33090.0 -437.5 33155.0 ;
      RECT  -302.5 32900.0 -437.5 32965.0 ;
      RECT  -1232.5 33260.0 -1367.5 33325.0 ;
      RECT  -257.5 33260.0 -392.5 33325.0 ;
      RECT  -515.0 33095.0 -580.0 32960.0 ;
      RECT  -655.0 32905.0 -720.0 32770.0 ;
      RECT  -795.0 32715.0 -860.0 32580.0 ;
      RECT  -1142.5 32710.0 -1277.5 32775.0 ;
      RECT  -1142.5 33090.0 -1277.5 33155.0 ;
      RECT  -302.5 33090.0 -437.5 33155.0 ;
      RECT  -760.0 33090.0 -895.0 33155.0 ;
      RECT  -795.0 32580.0 -860.0 32715.0 ;
      RECT  -655.0 32770.0 -720.0 32905.0 ;
      RECT  -515.0 32960.0 -580.0 33095.0 ;
      RECT  -760.0 33090.0 -895.0 33155.0 ;
      RECT  -1452.5 32452.5 -1517.5 33462.5 ;
      RECT  -107.5 32452.5 -172.5 33462.5 ;
      RECT  -1300.0 33890.0 -1485.0 33955.0 ;
      RECT  -140.0 33890.0 -325.0 33955.0 ;
      RECT  -257.5 33530.0 -107.5 33595.0 ;
      RECT  -1142.5 33530.0 -1517.5 33595.0 ;
      RECT  -257.5 33720.0 -1142.5 33785.0 ;
      RECT  -1142.5 33530.0 -1277.5 33595.0 ;
      RECT  -1142.5 33720.0 -1277.5 33785.0 ;
      RECT  -1142.5 33720.0 -1277.5 33785.0 ;
      RECT  -1142.5 33530.0 -1277.5 33595.0 ;
      RECT  -257.5 33530.0 -392.5 33595.0 ;
      RECT  -257.5 33720.0 -392.5 33785.0 ;
      RECT  -257.5 33720.0 -392.5 33785.0 ;
      RECT  -257.5 33530.0 -392.5 33595.0 ;
      RECT  -1232.5 33890.0 -1367.5 33955.0 ;
      RECT  -257.5 33890.0 -392.5 33955.0 ;
      RECT  -700.0 33587.5 -835.0 33652.5 ;
      RECT  -700.0 33587.5 -835.0 33652.5 ;
      RECT  -735.0 33752.5 -800.0 33817.5 ;
      RECT  -1452.5 33462.5 -1517.5 34022.5 ;
      RECT  -107.5 33462.5 -172.5 34022.5 ;
      RECT  -2712.5 32520.0 -2862.5 32585.0 ;
      RECT  -2712.5 32900.0 -2862.5 32965.0 ;
      RECT  -1895.0 32520.0 -1452.5 32585.0 ;
      RECT  -1670.0 33070.0 -1485.0 33135.0 ;
      RECT  -2830.0 33070.0 -2645.0 33135.0 ;
      RECT  -1895.0 32520.0 -1760.0 32585.0 ;
      RECT  -1895.0 32710.0 -1760.0 32775.0 ;
      RECT  -1895.0 32710.0 -1760.0 32775.0 ;
      RECT  -1895.0 32520.0 -1760.0 32585.0 ;
      RECT  -1895.0 32710.0 -1760.0 32775.0 ;
      RECT  -1895.0 32900.0 -1760.0 32965.0 ;
      RECT  -1895.0 32900.0 -1760.0 32965.0 ;
      RECT  -1895.0 32710.0 -1760.0 32775.0 ;
      RECT  -2712.5 32520.0 -2577.5 32585.0 ;
      RECT  -2712.5 32710.0 -2577.5 32775.0 ;
      RECT  -2712.5 32710.0 -2577.5 32775.0 ;
      RECT  -2712.5 32520.0 -2577.5 32585.0 ;
      RECT  -2712.5 32710.0 -2577.5 32775.0 ;
      RECT  -2712.5 32900.0 -2577.5 32965.0 ;
      RECT  -2712.5 32900.0 -2577.5 32965.0 ;
      RECT  -2712.5 32710.0 -2577.5 32775.0 ;
      RECT  -1737.5 33070.0 -1602.5 33135.0 ;
      RECT  -2712.5 33070.0 -2577.5 33135.0 ;
      RECT  -2492.5 32905.0 -2427.5 32770.0 ;
      RECT  -2277.5 32647.5 -2212.5 32512.5 ;
      RECT  -1895.0 32900.0 -1760.0 32965.0 ;
      RECT  -2677.5 32810.0 -2612.5 32675.0 ;
      RECT  -2277.5 33070.0 -2212.5 32935.0 ;
      RECT  -2277.5 32512.5 -2212.5 32647.5 ;
      RECT  -2492.5 32770.0 -2427.5 32905.0 ;
      RECT  -2277.5 32935.0 -2212.5 33070.0 ;
      RECT  -1517.5 32452.5 -1452.5 33372.5 ;
      RECT  -2862.5 32452.5 -2797.5 33372.5 ;
      RECT  -2667.5 33665.0 -2862.5 33730.0 ;
      RECT  -1827.5 33665.0 -1452.5 33730.0 ;
      RECT  -1827.5 34045.0 -1452.5 34110.0 ;
      RECT  -1670.0 34215.0 -1485.0 34280.0 ;
      RECT  -2830.0 34215.0 -2645.0 34280.0 ;
      RECT  -1827.5 33665.0 -1692.5 33730.0 ;
      RECT  -1827.5 33855.0 -1692.5 33920.0 ;
      RECT  -1827.5 33855.0 -1692.5 33920.0 ;
      RECT  -1827.5 33665.0 -1692.5 33730.0 ;
      RECT  -1827.5 33855.0 -1692.5 33920.0 ;
      RECT  -1827.5 34045.0 -1692.5 34110.0 ;
      RECT  -1827.5 34045.0 -1692.5 34110.0 ;
      RECT  -1827.5 33855.0 -1692.5 33920.0 ;
      RECT  -2667.5 33665.0 -2532.5 33730.0 ;
      RECT  -2667.5 33855.0 -2532.5 33920.0 ;
      RECT  -2667.5 33855.0 -2532.5 33920.0 ;
      RECT  -2667.5 33665.0 -2532.5 33730.0 ;
      RECT  -2667.5 33855.0 -2532.5 33920.0 ;
      RECT  -2667.5 34045.0 -2532.5 34110.0 ;
      RECT  -2667.5 34045.0 -2532.5 34110.0 ;
      RECT  -2667.5 33855.0 -2532.5 33920.0 ;
      RECT  -1737.5 34215.0 -1602.5 34280.0 ;
      RECT  -2712.5 34215.0 -2577.5 34280.0 ;
      RECT  -2437.5 34050.0 -2372.5 33915.0 ;
      RECT  -2222.5 33792.5 -2157.5 33657.5 ;
      RECT  -1827.5 33855.0 -1692.5 33920.0 ;
      RECT  -2667.5 34045.0 -2532.5 34110.0 ;
      RECT  -2222.5 34145.0 -2157.5 34010.0 ;
      RECT  -2222.5 33657.5 -2157.5 33792.5 ;
      RECT  -2437.5 33915.0 -2372.5 34050.0 ;
      RECT  -2222.5 34010.0 -2157.5 34145.0 ;
      RECT  -1517.5 33597.5 -1452.5 34517.5 ;
      RECT  -2862.5 33597.5 -2797.5 34517.5 ;
      RECT  -1670.0 34875.0 -1485.0 34810.0 ;
      RECT  -2830.0 34875.0 -2645.0 34810.0 ;
      RECT  -2712.5 35235.0 -2862.5 35170.0 ;
      RECT  -1827.5 35235.0 -1452.5 35170.0 ;
      RECT  -2712.5 35045.0 -1827.5 34980.0 ;
      RECT  -1827.5 35235.0 -1692.5 35170.0 ;
      RECT  -1827.5 35045.0 -1692.5 34980.0 ;
      RECT  -1827.5 35045.0 -1692.5 34980.0 ;
      RECT  -1827.5 35235.0 -1692.5 35170.0 ;
      RECT  -2712.5 35235.0 -2577.5 35170.0 ;
      RECT  -2712.5 35045.0 -2577.5 34980.0 ;
      RECT  -2712.5 35045.0 -2577.5 34980.0 ;
      RECT  -2712.5 35235.0 -2577.5 35170.0 ;
      RECT  -1737.5 34875.0 -1602.5 34810.0 ;
      RECT  -2712.5 34875.0 -2577.5 34810.0 ;
      RECT  -2270.0 35177.5 -2135.0 35112.5 ;
      RECT  -2270.0 35177.5 -2135.0 35112.5 ;
      RECT  -2235.0 35012.5 -2170.0 34947.5 ;
      RECT  -1517.5 35302.5 -1452.5 34742.5 ;
      RECT  -2862.5 35302.5 -2797.5 34742.5 ;
      RECT  -1670.0 35435.0 -1485.0 35370.0 ;
      RECT  -2830.0 35435.0 -2645.0 35370.0 ;
      RECT  -2712.5 35795.0 -2862.5 35730.0 ;
      RECT  -1827.5 35795.0 -1452.5 35730.0 ;
      RECT  -2712.5 35605.0 -1827.5 35540.0 ;
      RECT  -1827.5 35795.0 -1692.5 35730.0 ;
      RECT  -1827.5 35605.0 -1692.5 35540.0 ;
      RECT  -1827.5 35605.0 -1692.5 35540.0 ;
      RECT  -1827.5 35795.0 -1692.5 35730.0 ;
      RECT  -2712.5 35795.0 -2577.5 35730.0 ;
      RECT  -2712.5 35605.0 -2577.5 35540.0 ;
      RECT  -2712.5 35605.0 -2577.5 35540.0 ;
      RECT  -2712.5 35795.0 -2577.5 35730.0 ;
      RECT  -1737.5 35435.0 -1602.5 35370.0 ;
      RECT  -2712.5 35435.0 -2577.5 35370.0 ;
      RECT  -2270.0 35737.5 -2135.0 35672.5 ;
      RECT  -2270.0 35737.5 -2135.0 35672.5 ;
      RECT  -2235.0 35572.5 -2170.0 35507.5 ;
      RECT  -1517.5 35862.5 -1452.5 35302.5 ;
      RECT  -2862.5 35862.5 -2797.5 35302.5 ;
      RECT  -2992.5 33080.0 -2797.5 33145.0 ;
      RECT  -3832.5 33080.0 -4207.5 33145.0 ;
      RECT  -3832.5 33460.0 -4207.5 33525.0 ;
      RECT  -3990.0 33820.0 -4175.0 33885.0 ;
      RECT  -2830.0 33820.0 -3015.0 33885.0 ;
      RECT  -3832.5 33080.0 -3967.5 33145.0 ;
      RECT  -3832.5 33270.0 -3967.5 33335.0 ;
      RECT  -3832.5 33270.0 -3967.5 33335.0 ;
      RECT  -3832.5 33080.0 -3967.5 33145.0 ;
      RECT  -3832.5 33270.0 -3967.5 33335.0 ;
      RECT  -3832.5 33460.0 -3967.5 33525.0 ;
      RECT  -3832.5 33460.0 -3967.5 33525.0 ;
      RECT  -3832.5 33270.0 -3967.5 33335.0 ;
      RECT  -3832.5 33460.0 -3967.5 33525.0 ;
      RECT  -3832.5 33650.0 -3967.5 33715.0 ;
      RECT  -3832.5 33650.0 -3967.5 33715.0 ;
      RECT  -3832.5 33460.0 -3967.5 33525.0 ;
      RECT  -2992.5 33080.0 -3127.5 33145.0 ;
      RECT  -2992.5 33270.0 -3127.5 33335.0 ;
      RECT  -2992.5 33270.0 -3127.5 33335.0 ;
      RECT  -2992.5 33080.0 -3127.5 33145.0 ;
      RECT  -2992.5 33270.0 -3127.5 33335.0 ;
      RECT  -2992.5 33460.0 -3127.5 33525.0 ;
      RECT  -2992.5 33460.0 -3127.5 33525.0 ;
      RECT  -2992.5 33270.0 -3127.5 33335.0 ;
      RECT  -2992.5 33460.0 -3127.5 33525.0 ;
      RECT  -2992.5 33650.0 -3127.5 33715.0 ;
      RECT  -2992.5 33650.0 -3127.5 33715.0 ;
      RECT  -2992.5 33460.0 -3127.5 33525.0 ;
      RECT  -3922.5 33820.0 -4057.5 33885.0 ;
      RECT  -2947.5 33820.0 -3082.5 33885.0 ;
      RECT  -3205.0 33655.0 -3270.0 33520.0 ;
      RECT  -3345.0 33465.0 -3410.0 33330.0 ;
      RECT  -3485.0 33275.0 -3550.0 33140.0 ;
      RECT  -3832.5 33270.0 -3967.5 33335.0 ;
      RECT  -3832.5 33650.0 -3967.5 33715.0 ;
      RECT  -2992.5 33650.0 -3127.5 33715.0 ;
      RECT  -3450.0 33650.0 -3585.0 33715.0 ;
      RECT  -3485.0 33140.0 -3550.0 33275.0 ;
      RECT  -3345.0 33330.0 -3410.0 33465.0 ;
      RECT  -3205.0 33520.0 -3270.0 33655.0 ;
      RECT  -3450.0 33650.0 -3585.0 33715.0 ;
      RECT  -4142.5 33012.5 -4207.5 34022.5 ;
      RECT  -2797.5 33012.5 -2862.5 34022.5 ;
      RECT  -3990.0 34450.0 -4175.0 34515.0 ;
      RECT  -2830.0 34450.0 -3015.0 34515.0 ;
      RECT  -2947.5 34090.0 -2797.5 34155.0 ;
      RECT  -3832.5 34090.0 -4207.5 34155.0 ;
      RECT  -2947.5 34280.0 -3832.5 34345.0 ;
      RECT  -3832.5 34090.0 -3967.5 34155.0 ;
      RECT  -3832.5 34280.0 -3967.5 34345.0 ;
      RECT  -3832.5 34280.0 -3967.5 34345.0 ;
      RECT  -3832.5 34090.0 -3967.5 34155.0 ;
      RECT  -2947.5 34090.0 -3082.5 34155.0 ;
      RECT  -2947.5 34280.0 -3082.5 34345.0 ;
      RECT  -2947.5 34280.0 -3082.5 34345.0 ;
      RECT  -2947.5 34090.0 -3082.5 34155.0 ;
      RECT  -3922.5 34450.0 -4057.5 34515.0 ;
      RECT  -2947.5 34450.0 -3082.5 34515.0 ;
      RECT  -3390.0 34147.5 -3525.0 34212.5 ;
      RECT  -3390.0 34147.5 -3525.0 34212.5 ;
      RECT  -3425.0 34312.5 -3490.0 34377.5 ;
      RECT  -4142.5 34022.5 -4207.5 34582.5 ;
      RECT  -2797.5 34022.5 -2862.5 34582.5 ;
      RECT  -3990.0 35010.0 -4175.0 35075.0 ;
      RECT  -2830.0 35010.0 -3015.0 35075.0 ;
      RECT  -2947.5 34650.0 -2797.5 34715.0 ;
      RECT  -3832.5 34650.0 -4207.5 34715.0 ;
      RECT  -2947.5 34840.0 -3832.5 34905.0 ;
      RECT  -3832.5 34650.0 -3967.5 34715.0 ;
      RECT  -3832.5 34840.0 -3967.5 34905.0 ;
      RECT  -3832.5 34840.0 -3967.5 34905.0 ;
      RECT  -3832.5 34650.0 -3967.5 34715.0 ;
      RECT  -2947.5 34650.0 -3082.5 34715.0 ;
      RECT  -2947.5 34840.0 -3082.5 34905.0 ;
      RECT  -2947.5 34840.0 -3082.5 34905.0 ;
      RECT  -2947.5 34650.0 -3082.5 34715.0 ;
      RECT  -3922.5 35010.0 -4057.5 35075.0 ;
      RECT  -2947.5 35010.0 -3082.5 35075.0 ;
      RECT  -3390.0 34707.5 -3525.0 34772.5 ;
      RECT  -3390.0 34707.5 -3525.0 34772.5 ;
      RECT  -3425.0 34872.5 -3490.0 34937.5 ;
      RECT  -4142.5 34582.5 -4207.5 35142.5 ;
      RECT  -2797.5 34582.5 -2862.5 35142.5 ;
      RECT  -3990.0 35570.0 -4175.0 35635.0 ;
      RECT  -2830.0 35570.0 -3015.0 35635.0 ;
      RECT  -2947.5 35210.0 -2797.5 35275.0 ;
      RECT  -3832.5 35210.0 -4207.5 35275.0 ;
      RECT  -2947.5 35400.0 -3832.5 35465.0 ;
      RECT  -3832.5 35210.0 -3967.5 35275.0 ;
      RECT  -3832.5 35400.0 -3967.5 35465.0 ;
      RECT  -3832.5 35400.0 -3967.5 35465.0 ;
      RECT  -3832.5 35210.0 -3967.5 35275.0 ;
      RECT  -2947.5 35210.0 -3082.5 35275.0 ;
      RECT  -2947.5 35400.0 -3082.5 35465.0 ;
      RECT  -2947.5 35400.0 -3082.5 35465.0 ;
      RECT  -2947.5 35210.0 -3082.5 35275.0 ;
      RECT  -3922.5 35570.0 -4057.5 35635.0 ;
      RECT  -2947.5 35570.0 -3082.5 35635.0 ;
      RECT  -3390.0 35267.5 -3525.0 35332.5 ;
      RECT  -3390.0 35267.5 -3525.0 35332.5 ;
      RECT  -3425.0 35432.5 -3490.0 35497.5 ;
      RECT  -4142.5 35142.5 -4207.5 35702.5 ;
      RECT  -2797.5 35142.5 -2862.5 35702.5 ;
      RECT  -2797.5 42745.0 -2862.5 44172.5 ;
      RECT  -2862.5 38435.0 -3150.0 38500.0 ;
      RECT  -2862.5 40845.0 -3150.0 40910.0 ;
      RECT  -2862.5 41125.0 -3150.0 41190.0 ;
      RECT  -2862.5 43535.0 -3150.0 43600.0 ;
      RECT  -2797.5 36390.0 -3240.0 36455.0 ;
      RECT  -3240.0 36390.0 -3945.0 36455.0 ;
      RECT  -4155.0 39640.0 -3240.0 39705.0 ;
      RECT  -4155.0 42330.0 -3240.0 42395.0 ;
      RECT  -4155.0 36950.0 -3240.0 37015.0 ;
      RECT  -2170.0 37962.5 -2235.0 38662.5 ;
      RECT  -2170.0 38155.0 -2235.0 38220.0 ;
      RECT  -2170.0 37962.5 -2235.0 38187.5 ;
      RECT  -2202.5 38155.0 -3150.0 38220.0 ;
      RECT  -1485.0 38025.0 -1710.0 38090.0 ;
      RECT  -1745.0 37155.0 -1810.0 37220.0 ;
      RECT  -2170.0 37155.0 -2235.0 37220.0 ;
      RECT  -1745.0 37187.5 -1810.0 37835.0 ;
      RECT  -1777.5 37155.0 -2202.5 37220.0 ;
      RECT  -2170.0 36857.5 -2235.0 37187.5 ;
      RECT  -2202.5 37155.0 -3002.5 37220.0 ;
      RECT  -3002.5 36557.5 -3425.0 36622.5 ;
      RECT  -2135.0 36792.5 -2270.0 36857.5 ;
      RECT  -2170.0 38662.5 -2235.0 38867.5 ;
      RECT  -1670.0 36555.0 -1485.0 36490.0 ;
      RECT  -2830.0 36555.0 -2645.0 36490.0 ;
      RECT  -2712.5 36915.0 -2862.5 36850.0 ;
      RECT  -1827.5 36915.0 -1452.5 36850.0 ;
      RECT  -2712.5 36725.0 -1827.5 36660.0 ;
      RECT  -1827.5 36915.0 -1692.5 36850.0 ;
      RECT  -1827.5 36725.0 -1692.5 36660.0 ;
      RECT  -1827.5 36725.0 -1692.5 36660.0 ;
      RECT  -1827.5 36915.0 -1692.5 36850.0 ;
      RECT  -2712.5 36915.0 -2577.5 36850.0 ;
      RECT  -2712.5 36725.0 -2577.5 36660.0 ;
      RECT  -2712.5 36725.0 -2577.5 36660.0 ;
      RECT  -2712.5 36915.0 -2577.5 36850.0 ;
      RECT  -1737.5 36555.0 -1602.5 36490.0 ;
      RECT  -2712.5 36555.0 -2577.5 36490.0 ;
      RECT  -2270.0 36857.5 -2135.0 36792.5 ;
      RECT  -2270.0 36857.5 -2135.0 36792.5 ;
      RECT  -2235.0 36692.5 -2170.0 36627.5 ;
      RECT  -1517.5 36982.5 -1452.5 36422.5 ;
      RECT  -2862.5 36982.5 -2797.5 36422.5 ;
      RECT  -1845.0 37835.0 -1710.0 37900.0 ;
      RECT  -1845.0 38025.0 -1710.0 38090.0 ;
      RECT  -1845.0 38025.0 -1710.0 38090.0 ;
      RECT  -1845.0 37835.0 -1710.0 37900.0 ;
      RECT  -2862.5 42680.0 -2797.5 42745.0 ;
      RECT  -172.5 42680.0 -107.5 42745.0 ;
      RECT  -2862.5 42582.5 -2797.5 42712.5 ;
      RECT  -2830.0 42680.0 -140.0 42745.0 ;
      RECT  -172.5 42582.5 -107.5 42712.5 ;
      RECT  -1300.0 39090.0 -1485.0 39155.0 ;
      RECT  -140.0 39090.0 -325.0 39155.0 ;
      RECT  -257.5 38730.0 -107.5 38795.0 ;
      RECT  -1142.5 38730.0 -1517.5 38795.0 ;
      RECT  -257.5 38920.0 -1142.5 38985.0 ;
      RECT  -1142.5 38730.0 -1277.5 38795.0 ;
      RECT  -1142.5 38920.0 -1277.5 38985.0 ;
      RECT  -1142.5 38920.0 -1277.5 38985.0 ;
      RECT  -1142.5 38730.0 -1277.5 38795.0 ;
      RECT  -257.5 38730.0 -392.5 38795.0 ;
      RECT  -257.5 38920.0 -392.5 38985.0 ;
      RECT  -257.5 38920.0 -392.5 38985.0 ;
      RECT  -257.5 38730.0 -392.5 38795.0 ;
      RECT  -1232.5 39090.0 -1367.5 39155.0 ;
      RECT  -257.5 39090.0 -392.5 39155.0 ;
      RECT  -700.0 38787.5 -835.0 38852.5 ;
      RECT  -700.0 38787.5 -835.0 38852.5 ;
      RECT  -735.0 38952.5 -800.0 39017.5 ;
      RECT  -1452.5 38662.5 -1517.5 39222.5 ;
      RECT  -107.5 38662.5 -172.5 39222.5 ;
      RECT  -1300.0 39650.0 -1485.0 39715.0 ;
      RECT  -140.0 39650.0 -325.0 39715.0 ;
      RECT  -257.5 39290.0 -107.5 39355.0 ;
      RECT  -1142.5 39290.0 -1517.5 39355.0 ;
      RECT  -257.5 39480.0 -1142.5 39545.0 ;
      RECT  -1142.5 39290.0 -1277.5 39355.0 ;
      RECT  -1142.5 39480.0 -1277.5 39545.0 ;
      RECT  -1142.5 39480.0 -1277.5 39545.0 ;
      RECT  -1142.5 39290.0 -1277.5 39355.0 ;
      RECT  -257.5 39290.0 -392.5 39355.0 ;
      RECT  -257.5 39480.0 -392.5 39545.0 ;
      RECT  -257.5 39480.0 -392.5 39545.0 ;
      RECT  -257.5 39290.0 -392.5 39355.0 ;
      RECT  -1232.5 39650.0 -1367.5 39715.0 ;
      RECT  -257.5 39650.0 -392.5 39715.0 ;
      RECT  -700.0 39347.5 -835.0 39412.5 ;
      RECT  -700.0 39347.5 -835.0 39412.5 ;
      RECT  -735.0 39512.5 -800.0 39577.5 ;
      RECT  -1452.5 39222.5 -1517.5 39782.5 ;
      RECT  -107.5 39222.5 -172.5 39782.5 ;
      RECT  -835.0 39347.5 -700.0 39412.5 ;
      RECT  -1300.0 40210.0 -1485.0 40275.0 ;
      RECT  -140.0 40210.0 -325.0 40275.0 ;
      RECT  -257.5 39850.0 -107.5 39915.0 ;
      RECT  -1142.5 39850.0 -1517.5 39915.0 ;
      RECT  -257.5 40040.0 -1142.5 40105.0 ;
      RECT  -1142.5 39850.0 -1277.5 39915.0 ;
      RECT  -1142.5 40040.0 -1277.5 40105.0 ;
      RECT  -1142.5 40040.0 -1277.5 40105.0 ;
      RECT  -1142.5 39850.0 -1277.5 39915.0 ;
      RECT  -257.5 39850.0 -392.5 39915.0 ;
      RECT  -257.5 40040.0 -392.5 40105.0 ;
      RECT  -257.5 40040.0 -392.5 40105.0 ;
      RECT  -257.5 39850.0 -392.5 39915.0 ;
      RECT  -1232.5 40210.0 -1367.5 40275.0 ;
      RECT  -257.5 40210.0 -392.5 40275.0 ;
      RECT  -700.0 39907.5 -835.0 39972.5 ;
      RECT  -700.0 39907.5 -835.0 39972.5 ;
      RECT  -735.0 40072.5 -800.0 40137.5 ;
      RECT  -1452.5 39782.5 -1517.5 40342.5 ;
      RECT  -107.5 39782.5 -172.5 40342.5 ;
      RECT  -835.0 39907.5 -700.0 39972.5 ;
      RECT  -1300.0 40770.0 -1485.0 40835.0 ;
      RECT  -140.0 40770.0 -325.0 40835.0 ;
      RECT  -257.5 40410.0 -107.5 40475.0 ;
      RECT  -1142.5 40410.0 -1517.5 40475.0 ;
      RECT  -257.5 40600.0 -1142.5 40665.0 ;
      RECT  -1142.5 40410.0 -1277.5 40475.0 ;
      RECT  -1142.5 40600.0 -1277.5 40665.0 ;
      RECT  -1142.5 40600.0 -1277.5 40665.0 ;
      RECT  -1142.5 40410.0 -1277.5 40475.0 ;
      RECT  -257.5 40410.0 -392.5 40475.0 ;
      RECT  -257.5 40600.0 -392.5 40665.0 ;
      RECT  -257.5 40600.0 -392.5 40665.0 ;
      RECT  -257.5 40410.0 -392.5 40475.0 ;
      RECT  -1232.5 40770.0 -1367.5 40835.0 ;
      RECT  -257.5 40770.0 -392.5 40835.0 ;
      RECT  -700.0 40467.5 -835.0 40532.5 ;
      RECT  -700.0 40467.5 -835.0 40532.5 ;
      RECT  -735.0 40632.5 -800.0 40697.5 ;
      RECT  -1452.5 40342.5 -1517.5 40902.5 ;
      RECT  -107.5 40342.5 -172.5 40902.5 ;
      RECT  -835.0 40467.5 -700.0 40532.5 ;
      RECT  -1300.0 41330.0 -1485.0 41395.0 ;
      RECT  -140.0 41330.0 -325.0 41395.0 ;
      RECT  -257.5 40970.0 -107.5 41035.0 ;
      RECT  -1142.5 40970.0 -1517.5 41035.0 ;
      RECT  -257.5 41160.0 -1142.5 41225.0 ;
      RECT  -1142.5 40970.0 -1277.5 41035.0 ;
      RECT  -1142.5 41160.0 -1277.5 41225.0 ;
      RECT  -1142.5 41160.0 -1277.5 41225.0 ;
      RECT  -1142.5 40970.0 -1277.5 41035.0 ;
      RECT  -257.5 40970.0 -392.5 41035.0 ;
      RECT  -257.5 41160.0 -392.5 41225.0 ;
      RECT  -257.5 41160.0 -392.5 41225.0 ;
      RECT  -257.5 40970.0 -392.5 41035.0 ;
      RECT  -1232.5 41330.0 -1367.5 41395.0 ;
      RECT  -257.5 41330.0 -392.5 41395.0 ;
      RECT  -700.0 41027.5 -835.0 41092.5 ;
      RECT  -700.0 41027.5 -835.0 41092.5 ;
      RECT  -735.0 41192.5 -800.0 41257.5 ;
      RECT  -1452.5 40902.5 -1517.5 41462.5 ;
      RECT  -107.5 40902.5 -172.5 41462.5 ;
      RECT  -835.0 41027.5 -700.0 41092.5 ;
      RECT  -1300.0 41890.0 -1485.0 41955.0 ;
      RECT  -140.0 41890.0 -325.0 41955.0 ;
      RECT  -257.5 41530.0 -107.5 41595.0 ;
      RECT  -1142.5 41530.0 -1517.5 41595.0 ;
      RECT  -257.5 41720.0 -1142.5 41785.0 ;
      RECT  -1142.5 41530.0 -1277.5 41595.0 ;
      RECT  -1142.5 41720.0 -1277.5 41785.0 ;
      RECT  -1142.5 41720.0 -1277.5 41785.0 ;
      RECT  -1142.5 41530.0 -1277.5 41595.0 ;
      RECT  -257.5 41530.0 -392.5 41595.0 ;
      RECT  -257.5 41720.0 -392.5 41785.0 ;
      RECT  -257.5 41720.0 -392.5 41785.0 ;
      RECT  -257.5 41530.0 -392.5 41595.0 ;
      RECT  -1232.5 41890.0 -1367.5 41955.0 ;
      RECT  -257.5 41890.0 -392.5 41955.0 ;
      RECT  -700.0 41587.5 -835.0 41652.5 ;
      RECT  -700.0 41587.5 -835.0 41652.5 ;
      RECT  -735.0 41752.5 -800.0 41817.5 ;
      RECT  -1452.5 41462.5 -1517.5 42022.5 ;
      RECT  -107.5 41462.5 -172.5 42022.5 ;
      RECT  -835.0 41587.5 -700.0 41652.5 ;
      RECT  -1300.0 42450.0 -1485.0 42515.0 ;
      RECT  -140.0 42450.0 -325.0 42515.0 ;
      RECT  -257.5 42090.0 -107.5 42155.0 ;
      RECT  -1142.5 42090.0 -1517.5 42155.0 ;
      RECT  -257.5 42280.0 -1142.5 42345.0 ;
      RECT  -1142.5 42090.0 -1277.5 42155.0 ;
      RECT  -1142.5 42280.0 -1277.5 42345.0 ;
      RECT  -1142.5 42280.0 -1277.5 42345.0 ;
      RECT  -1142.5 42090.0 -1277.5 42155.0 ;
      RECT  -257.5 42090.0 -392.5 42155.0 ;
      RECT  -257.5 42280.0 -392.5 42345.0 ;
      RECT  -257.5 42280.0 -392.5 42345.0 ;
      RECT  -257.5 42090.0 -392.5 42155.0 ;
      RECT  -1232.5 42450.0 -1367.5 42515.0 ;
      RECT  -257.5 42450.0 -392.5 42515.0 ;
      RECT  -700.0 42147.5 -835.0 42212.5 ;
      RECT  -700.0 42147.5 -835.0 42212.5 ;
      RECT  -735.0 42312.5 -800.0 42377.5 ;
      RECT  -1452.5 42022.5 -1517.5 42582.5 ;
      RECT  -107.5 42022.5 -172.5 42582.5 ;
      RECT  -835.0 42147.5 -700.0 42212.5 ;
      RECT  -1670.0 41595.0 -1485.0 41530.0 ;
      RECT  -2830.0 41595.0 -2645.0 41530.0 ;
      RECT  -2712.5 41955.0 -2862.5 41890.0 ;
      RECT  -1827.5 41955.0 -1452.5 41890.0 ;
      RECT  -2712.5 41765.0 -1827.5 41700.0 ;
      RECT  -1827.5 41955.0 -1692.5 41890.0 ;
      RECT  -1827.5 41765.0 -1692.5 41700.0 ;
      RECT  -1827.5 41765.0 -1692.5 41700.0 ;
      RECT  -1827.5 41955.0 -1692.5 41890.0 ;
      RECT  -2712.5 41955.0 -2577.5 41890.0 ;
      RECT  -2712.5 41765.0 -2577.5 41700.0 ;
      RECT  -2712.5 41765.0 -2577.5 41700.0 ;
      RECT  -2712.5 41955.0 -2577.5 41890.0 ;
      RECT  -1737.5 41595.0 -1602.5 41530.0 ;
      RECT  -2712.5 41595.0 -2577.5 41530.0 ;
      RECT  -2270.0 41897.5 -2135.0 41832.5 ;
      RECT  -2270.0 41897.5 -2135.0 41832.5 ;
      RECT  -2235.0 41732.5 -2170.0 41667.5 ;
      RECT  -1517.5 42022.5 -1452.5 41462.5 ;
      RECT  -2862.5 42022.5 -2797.5 41462.5 ;
      RECT  -2270.0 41832.5 -2135.0 41897.5 ;
      RECT  -1670.0 41035.0 -1485.0 40970.0 ;
      RECT  -2830.0 41035.0 -2645.0 40970.0 ;
      RECT  -2712.5 41395.0 -2862.5 41330.0 ;
      RECT  -1827.5 41395.0 -1452.5 41330.0 ;
      RECT  -2712.5 41205.0 -1827.5 41140.0 ;
      RECT  -1827.5 41395.0 -1692.5 41330.0 ;
      RECT  -1827.5 41205.0 -1692.5 41140.0 ;
      RECT  -1827.5 41205.0 -1692.5 41140.0 ;
      RECT  -1827.5 41395.0 -1692.5 41330.0 ;
      RECT  -2712.5 41395.0 -2577.5 41330.0 ;
      RECT  -2712.5 41205.0 -2577.5 41140.0 ;
      RECT  -2712.5 41205.0 -2577.5 41140.0 ;
      RECT  -2712.5 41395.0 -2577.5 41330.0 ;
      RECT  -1737.5 41035.0 -1602.5 40970.0 ;
      RECT  -2712.5 41035.0 -2577.5 40970.0 ;
      RECT  -2270.0 41337.5 -2135.0 41272.5 ;
      RECT  -2270.0 41337.5 -2135.0 41272.5 ;
      RECT  -2235.0 41172.5 -2170.0 41107.5 ;
      RECT  -1517.5 41462.5 -1452.5 40902.5 ;
      RECT  -2862.5 41462.5 -2797.5 40902.5 ;
      RECT  -2270.0 41272.5 -2135.0 41337.5 ;
      RECT  -1670.0 40475.0 -1485.0 40410.0 ;
      RECT  -2830.0 40475.0 -2645.0 40410.0 ;
      RECT  -2712.5 40835.0 -2862.5 40770.0 ;
      RECT  -1827.5 40835.0 -1452.5 40770.0 ;
      RECT  -2712.5 40645.0 -1827.5 40580.0 ;
      RECT  -1827.5 40835.0 -1692.5 40770.0 ;
      RECT  -1827.5 40645.0 -1692.5 40580.0 ;
      RECT  -1827.5 40645.0 -1692.5 40580.0 ;
      RECT  -1827.5 40835.0 -1692.5 40770.0 ;
      RECT  -2712.5 40835.0 -2577.5 40770.0 ;
      RECT  -2712.5 40645.0 -2577.5 40580.0 ;
      RECT  -2712.5 40645.0 -2577.5 40580.0 ;
      RECT  -2712.5 40835.0 -2577.5 40770.0 ;
      RECT  -1737.5 40475.0 -1602.5 40410.0 ;
      RECT  -2712.5 40475.0 -2577.5 40410.0 ;
      RECT  -2270.0 40777.5 -2135.0 40712.5 ;
      RECT  -2270.0 40777.5 -2135.0 40712.5 ;
      RECT  -2235.0 40612.5 -2170.0 40547.5 ;
      RECT  -1517.5 40902.5 -1452.5 40342.5 ;
      RECT  -2862.5 40902.5 -2797.5 40342.5 ;
      RECT  -2270.0 40712.5 -2135.0 40777.5 ;
      RECT  -1670.0 39915.0 -1485.0 39850.0 ;
      RECT  -2830.0 39915.0 -2645.0 39850.0 ;
      RECT  -2712.5 40275.0 -2862.5 40210.0 ;
      RECT  -1827.5 40275.0 -1452.5 40210.0 ;
      RECT  -2712.5 40085.0 -1827.5 40020.0 ;
      RECT  -1827.5 40275.0 -1692.5 40210.0 ;
      RECT  -1827.5 40085.0 -1692.5 40020.0 ;
      RECT  -1827.5 40085.0 -1692.5 40020.0 ;
      RECT  -1827.5 40275.0 -1692.5 40210.0 ;
      RECT  -2712.5 40275.0 -2577.5 40210.0 ;
      RECT  -2712.5 40085.0 -2577.5 40020.0 ;
      RECT  -2712.5 40085.0 -2577.5 40020.0 ;
      RECT  -2712.5 40275.0 -2577.5 40210.0 ;
      RECT  -1737.5 39915.0 -1602.5 39850.0 ;
      RECT  -2712.5 39915.0 -2577.5 39850.0 ;
      RECT  -2270.0 40217.5 -2135.0 40152.5 ;
      RECT  -2270.0 40217.5 -2135.0 40152.5 ;
      RECT  -2235.0 40052.5 -2170.0 39987.5 ;
      RECT  -1517.5 40342.5 -1452.5 39782.5 ;
      RECT  -2862.5 40342.5 -2797.5 39782.5 ;
      RECT  -2270.0 40152.5 -2135.0 40217.5 ;
      RECT  -1670.0 39355.0 -1485.0 39290.0 ;
      RECT  -2830.0 39355.0 -2645.0 39290.0 ;
      RECT  -2712.5 39715.0 -2862.5 39650.0 ;
      RECT  -1827.5 39715.0 -1452.5 39650.0 ;
      RECT  -2712.5 39525.0 -1827.5 39460.0 ;
      RECT  -1827.5 39715.0 -1692.5 39650.0 ;
      RECT  -1827.5 39525.0 -1692.5 39460.0 ;
      RECT  -1827.5 39525.0 -1692.5 39460.0 ;
      RECT  -1827.5 39715.0 -1692.5 39650.0 ;
      RECT  -2712.5 39715.0 -2577.5 39650.0 ;
      RECT  -2712.5 39525.0 -2577.5 39460.0 ;
      RECT  -2712.5 39525.0 -2577.5 39460.0 ;
      RECT  -2712.5 39715.0 -2577.5 39650.0 ;
      RECT  -1737.5 39355.0 -1602.5 39290.0 ;
      RECT  -2712.5 39355.0 -2577.5 39290.0 ;
      RECT  -2270.0 39657.5 -2135.0 39592.5 ;
      RECT  -2270.0 39657.5 -2135.0 39592.5 ;
      RECT  -2235.0 39492.5 -2170.0 39427.5 ;
      RECT  -1517.5 39782.5 -1452.5 39222.5 ;
      RECT  -2862.5 39782.5 -2797.5 39222.5 ;
      RECT  -2270.0 39592.5 -2135.0 39657.5 ;
      RECT  -1670.0 38795.0 -1485.0 38730.0 ;
      RECT  -2830.0 38795.0 -2645.0 38730.0 ;
      RECT  -2712.5 39155.0 -2862.5 39090.0 ;
      RECT  -1827.5 39155.0 -1452.5 39090.0 ;
      RECT  -2712.5 38965.0 -1827.5 38900.0 ;
      RECT  -1827.5 39155.0 -1692.5 39090.0 ;
      RECT  -1827.5 38965.0 -1692.5 38900.0 ;
      RECT  -1827.5 38965.0 -1692.5 38900.0 ;
      RECT  -1827.5 39155.0 -1692.5 39090.0 ;
      RECT  -2712.5 39155.0 -2577.5 39090.0 ;
      RECT  -2712.5 38965.0 -2577.5 38900.0 ;
      RECT  -2712.5 38965.0 -2577.5 38900.0 ;
      RECT  -2712.5 39155.0 -2577.5 39090.0 ;
      RECT  -1737.5 38795.0 -1602.5 38730.0 ;
      RECT  -2712.5 38795.0 -2577.5 38730.0 ;
      RECT  -2270.0 39097.5 -2135.0 39032.5 ;
      RECT  -2270.0 39097.5 -2135.0 39032.5 ;
      RECT  -2235.0 38932.5 -2170.0 38867.5 ;
      RECT  -1517.5 39222.5 -1452.5 38662.5 ;
      RECT  -2862.5 39222.5 -2797.5 38662.5 ;
      RECT  -2270.0 39032.5 -2135.0 39097.5 ;
      RECT  -835.0 38952.5 -700.0 39017.5 ;
      RECT  -835.0 40632.5 -700.0 40697.5 ;
      RECT  -835.0 42312.5 -700.0 42377.5 ;
      RECT  -2270.0 40547.5 -2135.0 40612.5 ;
      RECT  -835.0 38787.5 -700.0 38852.5 ;
      RECT  -2235.0 38662.5 -2170.0 38867.5 ;
      RECT  -1517.5 38662.5 -1452.5 42582.5 ;
      RECT  -2862.5 38662.5 -2797.5 42582.5 ;
      RECT  -172.5 38662.5 -107.5 42582.5 ;
      RECT  -3240.0 38327.5 -3950.0 36982.5 ;
      RECT  -3240.0 38327.5 -3945.0 39672.5 ;
      RECT  -3240.0 41017.5 -3945.0 39672.5 ;
      RECT  -3240.0 41017.5 -3945.0 42362.5 ;
      RECT  -3240.0 43707.5 -3945.0 42362.5 ;
      RECT  -3150.0 38435.0 -4035.0 38500.0 ;
      RECT  -3150.0 40845.0 -4035.0 40910.0 ;
      RECT  -3150.0 41125.0 -4035.0 41190.0 ;
      RECT  -3150.0 43535.0 -4035.0 43600.0 ;
      RECT  -3150.0 39640.0 -4035.0 39705.0 ;
      RECT  -3150.0 42330.0 -4035.0 42395.0 ;
      RECT  -3150.0 38295.0 -4035.0 38360.0 ;
      RECT  -3150.0 40985.0 -4035.0 41050.0 ;
      RECT  -3150.0 43675.0 -4035.0 43740.0 ;
      RECT  -2830.0 38400.0 -2895.0 38535.0 ;
      RECT  -2830.0 40810.0 -2895.0 40945.0 ;
      RECT  -2830.0 41090.0 -2895.0 41225.0 ;
      RECT  -2830.0 43500.0 -2895.0 43635.0 ;
      RECT  -2832.5 38662.5 -2897.5 38797.5 ;
      RECT  -2797.5 36287.5 -2862.5 36422.5 ;
      RECT  -3307.5 36390.0 -3172.5 36455.0 ;
      RECT  -4012.5 36390.0 -3877.5 36455.0 ;
      RECT  -2170.0 37895.0 -2235.0 38030.0 ;
      RECT  -3070.0 37155.0 -2935.0 37220.0 ;
      RECT  -3070.0 36557.5 -2935.0 36622.5 ;
      RECT  -3492.5 36557.5 -3357.5 36622.5 ;
      RECT  -700.0 35862.5 -765.0 38787.5 ;
      RECT  -2170.0 35862.5 -2235.0 36627.5 ;
      RECT  -4155.0 35862.5 -4220.0 43795.0 ;
      RECT  -1452.5 35862.5 -1517.5 38662.5 ;
      RECT  -2797.5 35862.5 -2862.5 36422.5 ;
      RECT  -107.5 35862.5 -172.5 38662.5 ;
      RECT  -720.0 30710.0 -785.0 30575.0 ;
      RECT  -720.0 26630.0 -785.0 26495.0 ;
      RECT  -1657.5 24062.5 -1722.5 23927.5 ;
      RECT  -2212.5 30710.0 -2277.5 30575.0 ;
      RECT  -2427.5 31120.0 -2492.5 30985.0 ;
      RECT  -2157.5 33657.5 -2222.5 33522.5 ;
      RECT  -2372.5 33915.0 -2437.5 33780.0 ;
      RECT  -795.0 32145.0 -860.0 32010.0 ;
      RECT  -655.0 31940.0 -720.0 31805.0 ;
      RECT  -515.0 31325.0 -580.0 31190.0 ;
      RECT  -3485.0 32145.0 -3550.0 32010.0 ;
      RECT  -3345.0 31325.0 -3410.0 31190.0 ;
      RECT  -3205.0 31530.0 -3270.0 31395.0 ;
      RECT  -2177.5 33340.0 -2312.5 33405.0 ;
      RECT  -2122.5 34485.0 -2257.5 34550.0 ;
      RECT  -3390.0 35670.0 -3525.0 35735.0 ;
      RECT  -2135.0 34710.0 -2270.0 34775.0 ;
      RECT  -107.5 30915.0 -172.5 30780.0 ;
      RECT  -1452.5 31735.0 -1517.5 31600.0 ;
      RECT  -2797.5 30915.0 -2862.5 30780.0 ;
      RECT  -4142.5 31735.0 -4207.5 31600.0 ;
      RECT  -700.0 23757.5 -835.0 23947.5 ;
      RECT  -1452.5 23757.5 -1517.5 23822.5 ;
      RECT  -107.5 23757.5 -172.5 23822.5 ;
   LAYER  metal2 ;
      RECT  9430.0 34537.5 9500.0 34742.5 ;
      RECT  9225.0 35497.5 9295.0 35702.5 ;
      RECT  8815.0 33167.5 8885.0 33372.5 ;
      RECT  8610.0 34312.5 8680.0 34517.5 ;
      RECT  9020.0 31872.5 9090.0 32077.5 ;
      RECT  8405.0 30437.5 8475.0 30642.5 ;
      RECT  557.5 31462.5 627.5 31667.5 ;
      RECT  -140.0 30812.5 207.5 30882.5 ;
      RECT  8405.0 67.5 8475.0 44035.0 ;
      RECT  8610.0 67.5 8680.0 44035.0 ;
      RECT  8815.0 67.5 8885.0 44035.0 ;
      RECT  9020.0 67.5 9090.0 44035.0 ;
      RECT  9225.0 67.5 9295.0 44035.0 ;
      RECT  9430.0 67.5 9500.0 44035.0 ;
      RECT  7585.0 5527.5 7655.0 19927.5 ;
      RECT  7790.0 5527.5 7860.0 19927.5 ;
      RECT  7995.0 5527.5 8065.0 19927.5 ;
      RECT  8200.0 5527.5 8270.0 19927.5 ;
      RECT  10092.5 41602.5 10162.5 42007.5 ;
      RECT  10427.5 41602.5 10497.5 42007.5 ;
      RECT  10797.5 41602.5 10867.5 42007.5 ;
      RECT  11132.5 41602.5 11202.5 42007.5 ;
      RECT  10260.0 1277.5 10330.0 1347.5 ;
      RECT  10085.0 1277.5 10295.0 1347.5 ;
      RECT  10260.0 1312.5 10330.0 1452.5 ;
      RECT  10965.0 1277.5 11035.0 1347.5 ;
      RECT  10790.0 1277.5 11000.0 1347.5 ;
      RECT  10965.0 1312.5 11035.0 1452.5 ;
      RECT  4987.5 41447.5 5057.5 41652.5 ;
      RECT  9942.5 19927.5 10647.5 21272.5 ;
      RECT  9942.5 22617.5 10647.5 21272.5 ;
      RECT  9942.5 22617.5 10647.5 23962.5 ;
      RECT  9942.5 25307.5 10647.5 23962.5 ;
      RECT  9942.5 25307.5 10647.5 26652.5 ;
      RECT  9942.5 27997.5 10647.5 26652.5 ;
      RECT  9942.5 27997.5 10647.5 29342.5 ;
      RECT  9942.5 30687.5 10647.5 29342.5 ;
      RECT  9942.5 30687.5 10647.5 32032.5 ;
      RECT  9942.5 33377.5 10647.5 32032.5 ;
      RECT  9942.5 33377.5 10647.5 34722.5 ;
      RECT  9942.5 36067.5 10647.5 34722.5 ;
      RECT  9942.5 36067.5 10647.5 37412.5 ;
      RECT  9942.5 38757.5 10647.5 37412.5 ;
      RECT  9942.5 38757.5 10647.5 40102.5 ;
      RECT  9942.5 41447.5 10647.5 40102.5 ;
      RECT  10647.5 19927.5 11352.5 21272.5 ;
      RECT  10647.5 22617.5 11352.5 21272.5 ;
      RECT  10647.5 22617.5 11352.5 23962.5 ;
      RECT  10647.5 25307.5 11352.5 23962.5 ;
      RECT  10647.5 25307.5 11352.5 26652.5 ;
      RECT  10647.5 27997.5 11352.5 26652.5 ;
      RECT  10647.5 27997.5 11352.5 29342.5 ;
      RECT  10647.5 30687.5 11352.5 29342.5 ;
      RECT  10647.5 30687.5 11352.5 32032.5 ;
      RECT  10647.5 33377.5 11352.5 32032.5 ;
      RECT  10647.5 33377.5 11352.5 34722.5 ;
      RECT  10647.5 36067.5 11352.5 34722.5 ;
      RECT  10647.5 36067.5 11352.5 37412.5 ;
      RECT  10647.5 38757.5 11352.5 37412.5 ;
      RECT  10647.5 38757.5 11352.5 40102.5 ;
      RECT  10647.5 41447.5 11352.5 40102.5 ;
      RECT  10092.5 19827.5 10162.5 41602.5 ;
      RECT  10427.5 19827.5 10497.5 41602.5 ;
      RECT  10797.5 19827.5 10867.5 41602.5 ;
      RECT  11132.5 19827.5 11202.5 41602.5 ;
      RECT  9907.5 19827.5 9977.5 41602.5 ;
      RECT  10612.5 19827.5 10682.5 41602.5 ;
      RECT  11317.5 19827.5 11387.5 41602.5 ;
      RECT  10092.5 42130.0 10170.0 42265.0 ;
      RECT  10295.0 42130.0 10497.5 42265.0 ;
      RECT  10092.5 42660.0 10170.0 42795.0 ;
      RECT  10427.5 42660.0 10550.0 42795.0 ;
      RECT  10102.5 42130.0 10172.5 42265.0 ;
      RECT  10292.5 42130.0 10362.5 42265.0 ;
      RECT  10102.5 42660.0 10172.5 42795.0 ;
      RECT  10482.5 42660.0 10552.5 42795.0 ;
      RECT  10092.5 42007.5 10162.5 43175.0 ;
      RECT  10427.5 42007.5 10497.5 43175.0 ;
      RECT  10797.5 42130.0 10875.0 42265.0 ;
      RECT  11000.0 42130.0 11202.5 42265.0 ;
      RECT  10797.5 42660.0 10875.0 42795.0 ;
      RECT  11132.5 42660.0 11255.0 42795.0 ;
      RECT  10807.5 42130.0 10877.5 42265.0 ;
      RECT  10997.5 42130.0 11067.5 42265.0 ;
      RECT  10807.5 42660.0 10877.5 42795.0 ;
      RECT  11187.5 42660.0 11257.5 42795.0 ;
      RECT  10797.5 42007.5 10867.5 43175.0 ;
      RECT  11132.5 42007.5 11202.5 43175.0 ;
      RECT  10092.5 42007.5 10162.5 43175.0 ;
      RECT  10427.5 42007.5 10497.5 43175.0 ;
      RECT  10797.5 42007.5 10867.5 43175.0 ;
      RECT  11132.5 42007.5 11202.5 43175.0 ;
      RECT  9942.5 15042.5 10647.5 19927.5 ;
      RECT  10647.5 15042.5 11352.5 19927.5 ;
      RECT  10092.5 15042.5 10162.5 19927.5 ;
      RECT  10427.5 15042.5 10497.5 19127.5 ;
      RECT  10797.5 15042.5 10867.5 19927.5 ;
      RECT  11132.5 15042.5 11202.5 19127.5 ;
      RECT  9942.5 10867.5 10647.5 15042.5 ;
      RECT  10647.5 10867.5 11352.5 15042.5 ;
      RECT  10260.0 10867.5 10330.0 11007.5 ;
      RECT  10965.0 10867.5 11035.0 11007.5 ;
      RECT  10092.5 14742.5 10162.5 15042.5 ;
      RECT  10427.5 12602.5 10497.5 15042.5 ;
      RECT  10797.5 14742.5 10867.5 15042.5 ;
      RECT  11132.5 12602.5 11202.5 15042.5 ;
      RECT  9942.5 4427.5 10647.5 10867.5 ;
      RECT  11352.5 4427.5 10647.5 10867.5 ;
      RECT  10260.0 4427.5 10330.0 4572.5 ;
      RECT  10965.0 4427.5 11035.0 4572.5 ;
      RECT  10260.0 10597.5 10330.0 10867.5 ;
      RECT  10105.0 10180.0 10175.0 10867.5 ;
      RECT  10965.0 10597.5 11035.0 10867.5 ;
      RECT  11120.0 10180.0 11190.0 10867.5 ;
      RECT  9907.5 4427.5 9977.5 10867.5 ;
      RECT  10612.5 4427.5 10682.5 10867.5 ;
      RECT  11317.5 4427.5 11387.5 10867.5 ;
      RECT  9942.5 4427.5 10647.5 1452.5 ;
      RECT  10647.5 4427.5 11352.5 1452.5 ;
      RECT  10260.0 1692.5 10330.0 1452.5 ;
      RECT  10965.0 1692.5 11035.0 1452.5 ;
      RECT  10260.0 4427.5 10330.0 4077.5 ;
      RECT  10965.0 4427.5 11035.0 4077.5 ;
      RECT  1912.5 9167.5 1982.5 41447.5 ;
      RECT  2087.5 9167.5 2157.5 41447.5 ;
      RECT  2262.5 9167.5 2332.5 41447.5 ;
      RECT  2437.5 9167.5 2507.5 41447.5 ;
      RECT  2612.5 9167.5 2682.5 41447.5 ;
      RECT  2787.5 9167.5 2857.5 41447.5 ;
      RECT  2962.5 9167.5 3032.5 41447.5 ;
      RECT  3137.5 9167.5 3207.5 41447.5 ;
      RECT  5342.5 9167.5 5272.5 14407.5 ;
      RECT  5067.5 9167.5 4997.5 14407.5 ;
      RECT  5892.5 9167.5 5822.5 14407.5 ;
      RECT  5617.5 9167.5 5547.5 14407.5 ;
      RECT  4537.5 9772.5 4467.5 9842.5 ;
      RECT  4347.5 9772.5 4277.5 9842.5 ;
      RECT  4537.5 9807.5 4467.5 10170.0 ;
      RECT  4502.5 9772.5 4312.5 9842.5 ;
      RECT  4347.5 9465.0 4277.5 9807.5 ;
      RECT  4537.5 10170.0 4467.5 10305.0 ;
      RECT  4347.5 9330.0 4277.5 9465.0 ;
      RECT  4245.0 9772.5 4380.0 9842.5 ;
      RECT  4537.5 11252.5 4467.5 11182.5 ;
      RECT  4347.5 11252.5 4277.5 11182.5 ;
      RECT  4537.5 11217.5 4467.5 10855.0 ;
      RECT  4502.5 11252.5 4312.5 11182.5 ;
      RECT  4347.5 11560.0 4277.5 11217.5 ;
      RECT  4537.5 10855.0 4467.5 10720.0 ;
      RECT  4347.5 11695.0 4277.5 11560.0 ;
      RECT  4245.0 11252.5 4380.0 11182.5 ;
      RECT  4537.5 12462.5 4467.5 12532.5 ;
      RECT  4347.5 12462.5 4277.5 12532.5 ;
      RECT  4537.5 12497.5 4467.5 12860.0 ;
      RECT  4502.5 12462.5 4312.5 12532.5 ;
      RECT  4347.5 12155.0 4277.5 12497.5 ;
      RECT  4537.5 12860.0 4467.5 12995.0 ;
      RECT  4347.5 12020.0 4277.5 12155.0 ;
      RECT  4245.0 12462.5 4380.0 12532.5 ;
      RECT  4537.5 13942.5 4467.5 13872.5 ;
      RECT  4347.5 13942.5 4277.5 13872.5 ;
      RECT  4537.5 13907.5 4467.5 13545.0 ;
      RECT  4502.5 13942.5 4312.5 13872.5 ;
      RECT  4347.5 14250.0 4277.5 13907.5 ;
      RECT  4537.5 13545.0 4467.5 13410.0 ;
      RECT  4347.5 14385.0 4277.5 14250.0 ;
      RECT  4245.0 13942.5 4380.0 13872.5 ;
      RECT  5790.0 10282.5 5925.0 10352.5 ;
      RECT  7175.0 9760.0 7310.0 9830.0 ;
      RECT  5515.0 11627.5 5650.0 11697.5 ;
      RECT  6900.0 11195.0 7035.0 11265.0 ;
      RECT  7175.0 11957.5 7310.0 12027.5 ;
      RECT  5240.0 11957.5 5375.0 12027.5 ;
      RECT  6900.0 13302.5 7035.0 13372.5 ;
      RECT  4965.0 13302.5 5100.0 13372.5 ;
      RECT  5790.0 9772.5 5925.0 9842.5 ;
      RECT  5515.0 9557.5 5650.0 9627.5 ;
      RECT  5240.0 11182.5 5375.0 11252.5 ;
      RECT  5515.0 11397.5 5650.0 11467.5 ;
      RECT  5790.0 12462.5 5925.0 12532.5 ;
      RECT  4965.0 12247.5 5100.0 12317.5 ;
      RECT  5240.0 13872.5 5375.0 13942.5 ;
      RECT  4965.0 14087.5 5100.0 14157.5 ;
      RECT  7277.5 9167.5 7207.5 14407.5 ;
      RECT  7002.5 9167.5 6932.5 14407.5 ;
      RECT  5342.5 14547.5 5272.5 19787.5 ;
      RECT  5067.5 14547.5 4997.5 19787.5 ;
      RECT  5892.5 14547.5 5822.5 19787.5 ;
      RECT  5617.5 14547.5 5547.5 19787.5 ;
      RECT  4537.5 15152.5 4467.5 15222.5 ;
      RECT  4347.5 15152.5 4277.5 15222.5 ;
      RECT  4537.5 15187.5 4467.5 15550.0 ;
      RECT  4502.5 15152.5 4312.5 15222.5 ;
      RECT  4347.5 14845.0 4277.5 15187.5 ;
      RECT  4537.5 15550.0 4467.5 15685.0 ;
      RECT  4347.5 14710.0 4277.5 14845.0 ;
      RECT  4245.0 15152.5 4380.0 15222.5 ;
      RECT  4537.5 16632.5 4467.5 16562.5 ;
      RECT  4347.5 16632.5 4277.5 16562.5 ;
      RECT  4537.5 16597.5 4467.5 16235.0 ;
      RECT  4502.5 16632.5 4312.5 16562.5 ;
      RECT  4347.5 16940.0 4277.5 16597.5 ;
      RECT  4537.5 16235.0 4467.5 16100.0 ;
      RECT  4347.5 17075.0 4277.5 16940.0 ;
      RECT  4245.0 16632.5 4380.0 16562.5 ;
      RECT  4537.5 17842.5 4467.5 17912.5 ;
      RECT  4347.5 17842.5 4277.5 17912.5 ;
      RECT  4537.5 17877.5 4467.5 18240.0 ;
      RECT  4502.5 17842.5 4312.5 17912.5 ;
      RECT  4347.5 17535.0 4277.5 17877.5 ;
      RECT  4537.5 18240.0 4467.5 18375.0 ;
      RECT  4347.5 17400.0 4277.5 17535.0 ;
      RECT  4245.0 17842.5 4380.0 17912.5 ;
      RECT  4537.5 19322.5 4467.5 19252.5 ;
      RECT  4347.5 19322.5 4277.5 19252.5 ;
      RECT  4537.5 19287.5 4467.5 18925.0 ;
      RECT  4502.5 19322.5 4312.5 19252.5 ;
      RECT  4347.5 19630.0 4277.5 19287.5 ;
      RECT  4537.5 18925.0 4467.5 18790.0 ;
      RECT  4347.5 19765.0 4277.5 19630.0 ;
      RECT  4245.0 19322.5 4380.0 19252.5 ;
      RECT  5790.0 15662.5 5925.0 15732.5 ;
      RECT  7175.0 15140.0 7310.0 15210.0 ;
      RECT  5515.0 17007.5 5650.0 17077.5 ;
      RECT  6900.0 16575.0 7035.0 16645.0 ;
      RECT  7175.0 17337.5 7310.0 17407.5 ;
      RECT  5240.0 17337.5 5375.0 17407.5 ;
      RECT  6900.0 18682.5 7035.0 18752.5 ;
      RECT  4965.0 18682.5 5100.0 18752.5 ;
      RECT  5790.0 15152.5 5925.0 15222.5 ;
      RECT  5515.0 14937.5 5650.0 15007.5 ;
      RECT  5240.0 16562.5 5375.0 16632.5 ;
      RECT  5515.0 16777.5 5650.0 16847.5 ;
      RECT  5790.0 17842.5 5925.0 17912.5 ;
      RECT  4965.0 17627.5 5100.0 17697.5 ;
      RECT  5240.0 19252.5 5375.0 19322.5 ;
      RECT  4965.0 19467.5 5100.0 19537.5 ;
      RECT  7277.5 14547.5 7207.5 19787.5 ;
      RECT  7002.5 14547.5 6932.5 19787.5 ;
      RECT  3567.5 20532.5 3637.5 20602.5 ;
      RECT  3757.5 20532.5 3827.5 20602.5 ;
      RECT  3567.5 20567.5 3637.5 20930.0 ;
      RECT  3602.5 20532.5 3792.5 20602.5 ;
      RECT  3757.5 20225.0 3827.5 20567.5 ;
      RECT  3567.5 20930.0 3637.5 21065.0 ;
      RECT  3757.5 20090.0 3827.5 20225.0 ;
      RECT  3860.0 20532.5 3725.0 20602.5 ;
      RECT  3567.5 22012.5 3637.5 21942.5 ;
      RECT  3757.5 22012.5 3827.5 21942.5 ;
      RECT  3567.5 21977.5 3637.5 21615.0 ;
      RECT  3602.5 22012.5 3792.5 21942.5 ;
      RECT  3757.5 22320.0 3827.5 21977.5 ;
      RECT  3567.5 21615.0 3637.5 21480.0 ;
      RECT  3757.5 22455.0 3827.5 22320.0 ;
      RECT  3860.0 22012.5 3725.0 21942.5 ;
      RECT  3567.5 23222.5 3637.5 23292.5 ;
      RECT  3757.5 23222.5 3827.5 23292.5 ;
      RECT  3567.5 23257.5 3637.5 23620.0 ;
      RECT  3602.5 23222.5 3792.5 23292.5 ;
      RECT  3757.5 22915.0 3827.5 23257.5 ;
      RECT  3567.5 23620.0 3637.5 23755.0 ;
      RECT  3757.5 22780.0 3827.5 22915.0 ;
      RECT  3860.0 23222.5 3725.0 23292.5 ;
      RECT  3567.5 24702.5 3637.5 24632.5 ;
      RECT  3757.5 24702.5 3827.5 24632.5 ;
      RECT  3567.5 24667.5 3637.5 24305.0 ;
      RECT  3602.5 24702.5 3792.5 24632.5 ;
      RECT  3757.5 25010.0 3827.5 24667.5 ;
      RECT  3567.5 24305.0 3637.5 24170.0 ;
      RECT  3757.5 25145.0 3827.5 25010.0 ;
      RECT  3860.0 24702.5 3725.0 24632.5 ;
      RECT  3567.5 25912.5 3637.5 25982.5 ;
      RECT  3757.5 25912.5 3827.5 25982.5 ;
      RECT  3567.5 25947.5 3637.5 26310.0 ;
      RECT  3602.5 25912.5 3792.5 25982.5 ;
      RECT  3757.5 25605.0 3827.5 25947.5 ;
      RECT  3567.5 26310.0 3637.5 26445.0 ;
      RECT  3757.5 25470.0 3827.5 25605.0 ;
      RECT  3860.0 25912.5 3725.0 25982.5 ;
      RECT  3567.5 27392.5 3637.5 27322.5 ;
      RECT  3757.5 27392.5 3827.5 27322.5 ;
      RECT  3567.5 27357.5 3637.5 26995.0 ;
      RECT  3602.5 27392.5 3792.5 27322.5 ;
      RECT  3757.5 27700.0 3827.5 27357.5 ;
      RECT  3567.5 26995.0 3637.5 26860.0 ;
      RECT  3757.5 27835.0 3827.5 27700.0 ;
      RECT  3860.0 27392.5 3725.0 27322.5 ;
      RECT  3567.5 28602.5 3637.5 28672.5 ;
      RECT  3757.5 28602.5 3827.5 28672.5 ;
      RECT  3567.5 28637.5 3637.5 29000.0 ;
      RECT  3602.5 28602.5 3792.5 28672.5 ;
      RECT  3757.5 28295.0 3827.5 28637.5 ;
      RECT  3567.5 29000.0 3637.5 29135.0 ;
      RECT  3757.5 28160.0 3827.5 28295.0 ;
      RECT  3860.0 28602.5 3725.0 28672.5 ;
      RECT  3567.5 30082.5 3637.5 30012.5 ;
      RECT  3757.5 30082.5 3827.5 30012.5 ;
      RECT  3567.5 30047.5 3637.5 29685.0 ;
      RECT  3602.5 30082.5 3792.5 30012.5 ;
      RECT  3757.5 30390.0 3827.5 30047.5 ;
      RECT  3567.5 29685.0 3637.5 29550.0 ;
      RECT  3757.5 30525.0 3827.5 30390.0 ;
      RECT  3860.0 30082.5 3725.0 30012.5 ;
      RECT  3567.5 31292.5 3637.5 31362.5 ;
      RECT  3757.5 31292.5 3827.5 31362.5 ;
      RECT  3567.5 31327.5 3637.5 31690.0 ;
      RECT  3602.5 31292.5 3792.5 31362.5 ;
      RECT  3757.5 30985.0 3827.5 31327.5 ;
      RECT  3567.5 31690.0 3637.5 31825.0 ;
      RECT  3757.5 30850.0 3827.5 30985.0 ;
      RECT  3860.0 31292.5 3725.0 31362.5 ;
      RECT  3567.5 32772.5 3637.5 32702.5 ;
      RECT  3757.5 32772.5 3827.5 32702.5 ;
      RECT  3567.5 32737.5 3637.5 32375.0 ;
      RECT  3602.5 32772.5 3792.5 32702.5 ;
      RECT  3757.5 33080.0 3827.5 32737.5 ;
      RECT  3567.5 32375.0 3637.5 32240.0 ;
      RECT  3757.5 33215.0 3827.5 33080.0 ;
      RECT  3860.0 32772.5 3725.0 32702.5 ;
      RECT  3567.5 33982.5 3637.5 34052.5 ;
      RECT  3757.5 33982.5 3827.5 34052.5 ;
      RECT  3567.5 34017.5 3637.5 34380.0 ;
      RECT  3602.5 33982.5 3792.5 34052.5 ;
      RECT  3757.5 33675.0 3827.5 34017.5 ;
      RECT  3567.5 34380.0 3637.5 34515.0 ;
      RECT  3757.5 33540.0 3827.5 33675.0 ;
      RECT  3860.0 33982.5 3725.0 34052.5 ;
      RECT  3567.5 35462.5 3637.5 35392.5 ;
      RECT  3757.5 35462.5 3827.5 35392.5 ;
      RECT  3567.5 35427.5 3637.5 35065.0 ;
      RECT  3602.5 35462.5 3792.5 35392.5 ;
      RECT  3757.5 35770.0 3827.5 35427.5 ;
      RECT  3567.5 35065.0 3637.5 34930.0 ;
      RECT  3757.5 35905.0 3827.5 35770.0 ;
      RECT  3860.0 35462.5 3725.0 35392.5 ;
      RECT  3567.5 36672.5 3637.5 36742.5 ;
      RECT  3757.5 36672.5 3827.5 36742.5 ;
      RECT  3567.5 36707.5 3637.5 37070.0 ;
      RECT  3602.5 36672.5 3792.5 36742.5 ;
      RECT  3757.5 36365.0 3827.5 36707.5 ;
      RECT  3567.5 37070.0 3637.5 37205.0 ;
      RECT  3757.5 36230.0 3827.5 36365.0 ;
      RECT  3860.0 36672.5 3725.0 36742.5 ;
      RECT  3567.5 38152.5 3637.5 38082.5 ;
      RECT  3757.5 38152.5 3827.5 38082.5 ;
      RECT  3567.5 38117.5 3637.5 37755.0 ;
      RECT  3602.5 38152.5 3792.5 38082.5 ;
      RECT  3757.5 38460.0 3827.5 38117.5 ;
      RECT  3567.5 37755.0 3637.5 37620.0 ;
      RECT  3757.5 38595.0 3827.5 38460.0 ;
      RECT  3860.0 38152.5 3725.0 38082.5 ;
      RECT  3567.5 39362.5 3637.5 39432.5 ;
      RECT  3757.5 39362.5 3827.5 39432.5 ;
      RECT  3567.5 39397.5 3637.5 39760.0 ;
      RECT  3602.5 39362.5 3792.5 39432.5 ;
      RECT  3757.5 39055.0 3827.5 39397.5 ;
      RECT  3567.5 39760.0 3637.5 39895.0 ;
      RECT  3757.5 38920.0 3827.5 39055.0 ;
      RECT  3860.0 39362.5 3725.0 39432.5 ;
      RECT  3567.5 40842.5 3637.5 40772.5 ;
      RECT  3757.5 40842.5 3827.5 40772.5 ;
      RECT  3567.5 40807.5 3637.5 40445.0 ;
      RECT  3602.5 40842.5 3792.5 40772.5 ;
      RECT  3757.5 41150.0 3827.5 40807.5 ;
      RECT  3567.5 40445.0 3637.5 40310.0 ;
      RECT  3757.5 41285.0 3827.5 41150.0 ;
      RECT  3860.0 40842.5 3725.0 40772.5 ;
      RECT  2015.0 9760.0 1880.0 9830.0 ;
      RECT  2190.0 11195.0 2055.0 11265.0 ;
      RECT  2365.0 12450.0 2230.0 12520.0 ;
      RECT  2540.0 13885.0 2405.0 13955.0 ;
      RECT  2715.0 15140.0 2580.0 15210.0 ;
      RECT  2890.0 16575.0 2755.0 16645.0 ;
      RECT  3065.0 17830.0 2930.0 17900.0 ;
      RECT  3240.0 19265.0 3105.0 19335.0 ;
      RECT  2015.0 20532.5 1880.0 20602.5 ;
      RECT  2715.0 20317.5 2580.0 20387.5 ;
      RECT  2015.0 21942.5 1880.0 22012.5 ;
      RECT  2890.0 22157.5 2755.0 22227.5 ;
      RECT  2015.0 23222.5 1880.0 23292.5 ;
      RECT  3065.0 23007.5 2930.0 23077.5 ;
      RECT  2015.0 24632.5 1880.0 24702.5 ;
      RECT  3240.0 24847.5 3105.0 24917.5 ;
      RECT  2190.0 25912.5 2055.0 25982.5 ;
      RECT  2715.0 25697.5 2580.0 25767.5 ;
      RECT  2190.0 27322.5 2055.0 27392.5 ;
      RECT  2890.0 27537.5 2755.0 27607.5 ;
      RECT  2190.0 28602.5 2055.0 28672.5 ;
      RECT  3065.0 28387.5 2930.0 28457.5 ;
      RECT  2190.0 30012.5 2055.0 30082.5 ;
      RECT  3240.0 30227.5 3105.0 30297.5 ;
      RECT  2365.0 31292.5 2230.0 31362.5 ;
      RECT  2715.0 31077.5 2580.0 31147.5 ;
      RECT  2365.0 32702.5 2230.0 32772.5 ;
      RECT  2890.0 32917.5 2755.0 32987.5 ;
      RECT  2365.0 33982.5 2230.0 34052.5 ;
      RECT  3065.0 33767.5 2930.0 33837.5 ;
      RECT  2365.0 35392.5 2230.0 35462.5 ;
      RECT  3240.0 35607.5 3105.0 35677.5 ;
      RECT  2540.0 36672.5 2405.0 36742.5 ;
      RECT  2715.0 36457.5 2580.0 36527.5 ;
      RECT  2540.0 38082.5 2405.0 38152.5 ;
      RECT  2890.0 38297.5 2755.0 38367.5 ;
      RECT  2540.0 39362.5 2405.0 39432.5 ;
      RECT  3065.0 39147.5 2930.0 39217.5 ;
      RECT  2540.0 40772.5 2405.0 40842.5 ;
      RECT  3240.0 40987.5 3105.0 41057.5 ;
      RECT  7207.5 9167.5 7277.5 14407.5 ;
      RECT  6932.5 9167.5 7002.5 14407.5 ;
      RECT  7207.5 14547.5 7277.5 19787.5 ;
      RECT  6932.5 14547.5 7002.5 19787.5 ;
      RECT  5127.5 20317.5 5197.5 20387.5 ;
      RECT  5127.5 20282.5 5197.5 20352.5 ;
      RECT  5162.5 20317.5 6125.0 20387.5 ;
      RECT  5127.5 22157.5 5197.5 22227.5 ;
      RECT  5127.5 22192.5 5197.5 22262.5 ;
      RECT  5162.5 22157.5 6125.0 22227.5 ;
      RECT  5127.5 23007.5 5197.5 23077.5 ;
      RECT  5127.5 22972.5 5197.5 23042.5 ;
      RECT  5162.5 23007.5 6125.0 23077.5 ;
      RECT  5127.5 24847.5 5197.5 24917.5 ;
      RECT  5127.5 24882.5 5197.5 24952.5 ;
      RECT  5162.5 24847.5 6125.0 24917.5 ;
      RECT  5127.5 25697.5 5197.5 25767.5 ;
      RECT  5127.5 25662.5 5197.5 25732.5 ;
      RECT  5162.5 25697.5 6125.0 25767.5 ;
      RECT  5127.5 27537.5 5197.5 27607.5 ;
      RECT  5127.5 27572.5 5197.5 27642.5 ;
      RECT  5162.5 27537.5 6125.0 27607.5 ;
      RECT  5127.5 28387.5 5197.5 28457.5 ;
      RECT  5127.5 28352.5 5197.5 28422.5 ;
      RECT  5162.5 28387.5 6125.0 28457.5 ;
      RECT  5127.5 30227.5 5197.5 30297.5 ;
      RECT  5127.5 30262.5 5197.5 30332.5 ;
      RECT  5162.5 30227.5 6125.0 30297.5 ;
      RECT  5127.5 31077.5 5197.5 31147.5 ;
      RECT  5127.5 31042.5 5197.5 31112.5 ;
      RECT  5162.5 31077.5 6125.0 31147.5 ;
      RECT  5127.5 32917.5 5197.5 32987.5 ;
      RECT  5127.5 32952.5 5197.5 33022.5 ;
      RECT  5162.5 32917.5 6125.0 32987.5 ;
      RECT  5127.5 33767.5 5197.5 33837.5 ;
      RECT  5127.5 33732.5 5197.5 33802.5 ;
      RECT  5162.5 33767.5 6125.0 33837.5 ;
      RECT  5127.5 35607.5 5197.5 35677.5 ;
      RECT  5127.5 35642.5 5197.5 35712.5 ;
      RECT  5162.5 35607.5 6125.0 35677.5 ;
      RECT  5127.5 36457.5 5197.5 36527.5 ;
      RECT  5127.5 36422.5 5197.5 36492.5 ;
      RECT  5162.5 36457.5 6125.0 36527.5 ;
      RECT  5127.5 38297.5 5197.5 38367.5 ;
      RECT  5127.5 38332.5 5197.5 38402.5 ;
      RECT  5162.5 38297.5 6125.0 38367.5 ;
      RECT  5127.5 39147.5 5197.5 39217.5 ;
      RECT  5127.5 39112.5 5197.5 39182.5 ;
      RECT  5162.5 39147.5 6125.0 39217.5 ;
      RECT  5127.5 40987.5 5197.5 41057.5 ;
      RECT  5127.5 41022.5 5197.5 41092.5 ;
      RECT  5162.5 40987.5 6125.0 41057.5 ;
      RECT  6062.5 20532.5 6132.5 20602.5 ;
      RECT  6252.5 20532.5 6322.5 20602.5 ;
      RECT  6062.5 20567.5 6132.5 20930.0 ;
      RECT  6097.5 20532.5 6287.5 20602.5 ;
      RECT  6252.5 20225.0 6322.5 20567.5 ;
      RECT  6062.5 20930.0 6132.5 21065.0 ;
      RECT  6252.5 20090.0 6322.5 20225.0 ;
      RECT  6355.0 20532.5 6220.0 20602.5 ;
      RECT  4987.5 20487.5 5057.5 20622.5 ;
      RECT  5127.5 20215.0 5197.5 20350.0 ;
      RECT  6125.0 20317.5 5990.0 20387.5 ;
      RECT  6062.5 22012.5 6132.5 21942.5 ;
      RECT  6252.5 22012.5 6322.5 21942.5 ;
      RECT  6062.5 21977.5 6132.5 21615.0 ;
      RECT  6097.5 22012.5 6287.5 21942.5 ;
      RECT  6252.5 22320.0 6322.5 21977.5 ;
      RECT  6062.5 21615.0 6132.5 21480.0 ;
      RECT  6252.5 22455.0 6322.5 22320.0 ;
      RECT  6355.0 22012.5 6220.0 21942.5 ;
      RECT  4987.5 21922.5 5057.5 22057.5 ;
      RECT  5127.5 22195.0 5197.5 22330.0 ;
      RECT  6125.0 22157.5 5990.0 22227.5 ;
      RECT  6062.5 23222.5 6132.5 23292.5 ;
      RECT  6252.5 23222.5 6322.5 23292.5 ;
      RECT  6062.5 23257.5 6132.5 23620.0 ;
      RECT  6097.5 23222.5 6287.5 23292.5 ;
      RECT  6252.5 22915.0 6322.5 23257.5 ;
      RECT  6062.5 23620.0 6132.5 23755.0 ;
      RECT  6252.5 22780.0 6322.5 22915.0 ;
      RECT  6355.0 23222.5 6220.0 23292.5 ;
      RECT  4987.5 23177.5 5057.5 23312.5 ;
      RECT  5127.5 22905.0 5197.5 23040.0 ;
      RECT  6125.0 23007.5 5990.0 23077.5 ;
      RECT  6062.5 24702.5 6132.5 24632.5 ;
      RECT  6252.5 24702.5 6322.5 24632.5 ;
      RECT  6062.5 24667.5 6132.5 24305.0 ;
      RECT  6097.5 24702.5 6287.5 24632.5 ;
      RECT  6252.5 25010.0 6322.5 24667.5 ;
      RECT  6062.5 24305.0 6132.5 24170.0 ;
      RECT  6252.5 25145.0 6322.5 25010.0 ;
      RECT  6355.0 24702.5 6220.0 24632.5 ;
      RECT  4987.5 24612.5 5057.5 24747.5 ;
      RECT  5127.5 24885.0 5197.5 25020.0 ;
      RECT  6125.0 24847.5 5990.0 24917.5 ;
      RECT  6062.5 25912.5 6132.5 25982.5 ;
      RECT  6252.5 25912.5 6322.5 25982.5 ;
      RECT  6062.5 25947.5 6132.5 26310.0 ;
      RECT  6097.5 25912.5 6287.5 25982.5 ;
      RECT  6252.5 25605.0 6322.5 25947.5 ;
      RECT  6062.5 26310.0 6132.5 26445.0 ;
      RECT  6252.5 25470.0 6322.5 25605.0 ;
      RECT  6355.0 25912.5 6220.0 25982.5 ;
      RECT  4987.5 25867.5 5057.5 26002.5 ;
      RECT  5127.5 25595.0 5197.5 25730.0 ;
      RECT  6125.0 25697.5 5990.0 25767.5 ;
      RECT  6062.5 27392.5 6132.5 27322.5 ;
      RECT  6252.5 27392.5 6322.5 27322.5 ;
      RECT  6062.5 27357.5 6132.5 26995.0 ;
      RECT  6097.5 27392.5 6287.5 27322.5 ;
      RECT  6252.5 27700.0 6322.5 27357.5 ;
      RECT  6062.5 26995.0 6132.5 26860.0 ;
      RECT  6252.5 27835.0 6322.5 27700.0 ;
      RECT  6355.0 27392.5 6220.0 27322.5 ;
      RECT  4987.5 27302.5 5057.5 27437.5 ;
      RECT  5127.5 27575.0 5197.5 27710.0 ;
      RECT  6125.0 27537.5 5990.0 27607.5 ;
      RECT  6062.5 28602.5 6132.5 28672.5 ;
      RECT  6252.5 28602.5 6322.5 28672.5 ;
      RECT  6062.5 28637.5 6132.5 29000.0 ;
      RECT  6097.5 28602.5 6287.5 28672.5 ;
      RECT  6252.5 28295.0 6322.5 28637.5 ;
      RECT  6062.5 29000.0 6132.5 29135.0 ;
      RECT  6252.5 28160.0 6322.5 28295.0 ;
      RECT  6355.0 28602.5 6220.0 28672.5 ;
      RECT  4987.5 28557.5 5057.5 28692.5 ;
      RECT  5127.5 28285.0 5197.5 28420.0 ;
      RECT  6125.0 28387.5 5990.0 28457.5 ;
      RECT  6062.5 30082.5 6132.5 30012.5 ;
      RECT  6252.5 30082.5 6322.5 30012.5 ;
      RECT  6062.5 30047.5 6132.5 29685.0 ;
      RECT  6097.5 30082.5 6287.5 30012.5 ;
      RECT  6252.5 30390.0 6322.5 30047.5 ;
      RECT  6062.5 29685.0 6132.5 29550.0 ;
      RECT  6252.5 30525.0 6322.5 30390.0 ;
      RECT  6355.0 30082.5 6220.0 30012.5 ;
      RECT  4987.5 29992.5 5057.5 30127.5 ;
      RECT  5127.5 30265.0 5197.5 30400.0 ;
      RECT  6125.0 30227.5 5990.0 30297.5 ;
      RECT  6062.5 31292.5 6132.5 31362.5 ;
      RECT  6252.5 31292.5 6322.5 31362.5 ;
      RECT  6062.5 31327.5 6132.5 31690.0 ;
      RECT  6097.5 31292.5 6287.5 31362.5 ;
      RECT  6252.5 30985.0 6322.5 31327.5 ;
      RECT  6062.5 31690.0 6132.5 31825.0 ;
      RECT  6252.5 30850.0 6322.5 30985.0 ;
      RECT  6355.0 31292.5 6220.0 31362.5 ;
      RECT  4987.5 31247.5 5057.5 31382.5 ;
      RECT  5127.5 30975.0 5197.5 31110.0 ;
      RECT  6125.0 31077.5 5990.0 31147.5 ;
      RECT  6062.5 32772.5 6132.5 32702.5 ;
      RECT  6252.5 32772.5 6322.5 32702.5 ;
      RECT  6062.5 32737.5 6132.5 32375.0 ;
      RECT  6097.5 32772.5 6287.5 32702.5 ;
      RECT  6252.5 33080.0 6322.5 32737.5 ;
      RECT  6062.5 32375.0 6132.5 32240.0 ;
      RECT  6252.5 33215.0 6322.5 33080.0 ;
      RECT  6355.0 32772.5 6220.0 32702.5 ;
      RECT  4987.5 32682.5 5057.5 32817.5 ;
      RECT  5127.5 32955.0 5197.5 33090.0 ;
      RECT  6125.0 32917.5 5990.0 32987.5 ;
      RECT  6062.5 33982.5 6132.5 34052.5 ;
      RECT  6252.5 33982.5 6322.5 34052.5 ;
      RECT  6062.5 34017.5 6132.5 34380.0 ;
      RECT  6097.5 33982.5 6287.5 34052.5 ;
      RECT  6252.5 33675.0 6322.5 34017.5 ;
      RECT  6062.5 34380.0 6132.5 34515.0 ;
      RECT  6252.5 33540.0 6322.5 33675.0 ;
      RECT  6355.0 33982.5 6220.0 34052.5 ;
      RECT  4987.5 33937.5 5057.5 34072.5 ;
      RECT  5127.5 33665.0 5197.5 33800.0 ;
      RECT  6125.0 33767.5 5990.0 33837.5 ;
      RECT  6062.5 35462.5 6132.5 35392.5 ;
      RECT  6252.5 35462.5 6322.5 35392.5 ;
      RECT  6062.5 35427.5 6132.5 35065.0 ;
      RECT  6097.5 35462.5 6287.5 35392.5 ;
      RECT  6252.5 35770.0 6322.5 35427.5 ;
      RECT  6062.5 35065.0 6132.5 34930.0 ;
      RECT  6252.5 35905.0 6322.5 35770.0 ;
      RECT  6355.0 35462.5 6220.0 35392.5 ;
      RECT  4987.5 35372.5 5057.5 35507.5 ;
      RECT  5127.5 35645.0 5197.5 35780.0 ;
      RECT  6125.0 35607.5 5990.0 35677.5 ;
      RECT  6062.5 36672.5 6132.5 36742.5 ;
      RECT  6252.5 36672.5 6322.5 36742.5 ;
      RECT  6062.5 36707.5 6132.5 37070.0 ;
      RECT  6097.5 36672.5 6287.5 36742.5 ;
      RECT  6252.5 36365.0 6322.5 36707.5 ;
      RECT  6062.5 37070.0 6132.5 37205.0 ;
      RECT  6252.5 36230.0 6322.5 36365.0 ;
      RECT  6355.0 36672.5 6220.0 36742.5 ;
      RECT  4987.5 36627.5 5057.5 36762.5 ;
      RECT  5127.5 36355.0 5197.5 36490.0 ;
      RECT  6125.0 36457.5 5990.0 36527.5 ;
      RECT  6062.5 38152.5 6132.5 38082.5 ;
      RECT  6252.5 38152.5 6322.5 38082.5 ;
      RECT  6062.5 38117.5 6132.5 37755.0 ;
      RECT  6097.5 38152.5 6287.5 38082.5 ;
      RECT  6252.5 38460.0 6322.5 38117.5 ;
      RECT  6062.5 37755.0 6132.5 37620.0 ;
      RECT  6252.5 38595.0 6322.5 38460.0 ;
      RECT  6355.0 38152.5 6220.0 38082.5 ;
      RECT  4987.5 38062.5 5057.5 38197.5 ;
      RECT  5127.5 38335.0 5197.5 38470.0 ;
      RECT  6125.0 38297.5 5990.0 38367.5 ;
      RECT  6062.5 39362.5 6132.5 39432.5 ;
      RECT  6252.5 39362.5 6322.5 39432.5 ;
      RECT  6062.5 39397.5 6132.5 39760.0 ;
      RECT  6097.5 39362.5 6287.5 39432.5 ;
      RECT  6252.5 39055.0 6322.5 39397.5 ;
      RECT  6062.5 39760.0 6132.5 39895.0 ;
      RECT  6252.5 38920.0 6322.5 39055.0 ;
      RECT  6355.0 39362.5 6220.0 39432.5 ;
      RECT  4987.5 39317.5 5057.5 39452.5 ;
      RECT  5127.5 39045.0 5197.5 39180.0 ;
      RECT  6125.0 39147.5 5990.0 39217.5 ;
      RECT  6062.5 40842.5 6132.5 40772.5 ;
      RECT  6252.5 40842.5 6322.5 40772.5 ;
      RECT  6062.5 40807.5 6132.5 40445.0 ;
      RECT  6097.5 40842.5 6287.5 40772.5 ;
      RECT  6252.5 41150.0 6322.5 40807.5 ;
      RECT  6062.5 40445.0 6132.5 40310.0 ;
      RECT  6252.5 41285.0 6322.5 41150.0 ;
      RECT  6355.0 40842.5 6220.0 40772.5 ;
      RECT  4987.5 40752.5 5057.5 40887.5 ;
      RECT  5127.5 41025.0 5197.5 41160.0 ;
      RECT  6125.0 40987.5 5990.0 41057.5 ;
      RECT  4987.5 19927.5 5057.5 41447.5 ;
      RECT  837.5 8757.5 7277.5 8052.5 ;
      RECT  837.5 7347.5 7277.5 8052.5 ;
      RECT  837.5 7347.5 7277.5 6642.5 ;
      RECT  837.5 5937.5 7277.5 6642.5 ;
      RECT  837.5 8440.0 982.5 8370.0 ;
      RECT  837.5 7735.0 982.5 7665.0 ;
      RECT  837.5 7030.0 982.5 6960.0 ;
      RECT  837.5 6325.0 982.5 6255.0 ;
      RECT  7007.5 8440.0 7277.5 8370.0 ;
      RECT  6590.0 8595.0 7277.5 8525.0 ;
      RECT  7007.5 7735.0 7277.5 7665.0 ;
      RECT  6590.0 7580.0 7277.5 7510.0 ;
      RECT  7007.5 7030.0 7277.5 6960.0 ;
      RECT  6590.0 7185.0 7277.5 7115.0 ;
      RECT  7007.5 6325.0 7277.5 6255.0 ;
      RECT  6590.0 6170.0 7277.5 6100.0 ;
      RECT  837.5 8792.5 7277.5 8722.5 ;
      RECT  837.5 8087.5 7277.5 8017.5 ;
      RECT  837.5 7382.5 7277.5 7312.5 ;
      RECT  837.5 6677.5 7277.5 6607.5 ;
      RECT  837.5 5972.5 7277.5 5902.5 ;
      RECT  35.0 -3.5527136788e-12 380.0 415.0 ;
      RECT  35.0 43302.5 380.0 43717.5 ;
      RECT  11515.0 -3.5527136788e-12 11860.0 415.0 ;
      RECT  11515.0 43302.5 11860.0 43717.5 ;
      RECT  420.0 385.0 765.0 800.0 ;
      RECT  420.0 43687.5 765.0 44102.5 ;
      RECT  11900.0 385.0 12245.0 800.0 ;
      RECT  11900.0 43687.5 12245.0 44102.5 ;
      RECT  10050.0 1277.5 10120.0 1412.5 ;
      RECT  10755.0 1277.5 10825.0 1412.5 ;
      RECT  10260.0 67.5 10330.0 202.5 ;
      RECT  10965.0 67.5 11035.0 202.5 ;
      RECT  7277.5 9337.5 7142.5 9407.5 ;
      RECT  7687.5 9337.5 7552.5 9407.5 ;
      RECT  7002.5 10682.5 6867.5 10752.5 ;
      RECT  7892.5 10682.5 7757.5 10752.5 ;
      RECT  7277.5 14717.5 7142.5 14787.5 ;
      RECT  8097.5 14717.5 7962.5 14787.5 ;
      RECT  7002.5 16062.5 6867.5 16132.5 ;
      RECT  8302.5 16062.5 8167.5 16132.5 ;
      RECT  415.0 9132.5 -8.881784197e-13 9202.5 ;
      RECT  415.0 11822.5 -8.881784197e-13 11892.5 ;
      RECT  415.0 14512.5 -8.881784197e-13 14582.5 ;
      RECT  415.0 17202.5 -8.881784197e-13 17272.5 ;
      RECT  800.0 10477.5 385.0 10547.5 ;
      RECT  800.0 13167.5 385.0 13237.5 ;
      RECT  800.0 15857.5 385.0 15927.5 ;
      RECT  800.0 18547.5 385.0 18617.5 ;
      RECT  7345.0 8370.0 7210.0 8440.0 ;
      RECT  7687.5 8370.0 7552.5 8440.0 ;
      RECT  7345.0 7665.0 7210.0 7735.0 ;
      RECT  7892.5 7665.0 7757.5 7735.0 ;
      RECT  7345.0 6960.0 7210.0 7030.0 ;
      RECT  8097.5 6960.0 7962.5 7030.0 ;
      RECT  7345.0 6255.0 7210.0 6325.0 ;
      RECT  8302.5 6255.0 8167.5 6325.0 ;
      RECT  972.5 8722.5 837.5 8792.5 ;
      RECT  415.0 8722.5 -8.881784197e-13 8792.5 ;
      RECT  972.5 8017.5 837.5 8087.5 ;
      RECT  415.0 8017.5 -8.881784197e-13 8087.5 ;
      RECT  972.5 7312.5 837.5 7382.5 ;
      RECT  415.0 7312.5 -8.881784197e-13 7382.5 ;
      RECT  972.5 6607.5 837.5 6677.5 ;
      RECT  415.0 6607.5 -8.881784197e-13 6677.5 ;
      RECT  972.5 5902.5 837.5 5972.5 ;
      RECT  415.0 5902.5 -8.881784197e-13 5972.5 ;
      RECT  800.0 5697.5 385.0 5767.5 ;
      RECT  800.0 5697.5 385.0 5767.5 ;
      RECT  800.0 5697.5 385.0 5767.5 ;
      RECT  800.0 5697.5 385.0 5767.5 ;
      RECT  9122.5 4630.0 8987.5 4700.0 ;
      RECT  8712.5 2445.0 8577.5 2515.0 ;
      RECT  8917.5 3992.5 8782.5 4062.5 ;
      RECT  9122.5 42422.5 8987.5 42492.5 ;
      RECT  9327.5 11132.5 9192.5 11202.5 ;
      RECT  9532.5 15157.5 9397.5 15227.5 ;
      RECT  8507.5 8927.5 8372.5 8997.5 ;
      RECT  5090.0 41617.5 4955.0 41687.5 ;
      RECT  8507.5 41617.5 8372.5 41687.5 ;
      RECT  12280.0 43107.5 11865.0 43177.5 ;
      RECT  12280.0 19730.0 11865.0 19800.0 ;
      RECT  12280.0 11262.5 11865.0 11332.5 ;
      RECT  12280.0 7635.0 11865.0 7705.0 ;
      RECT  12280.0 10595.0 11865.0 10665.0 ;
      RECT  12280.0 5645.0 11865.0 5715.0 ;
      RECT  12280.0 8605.0 11865.0 8675.0 ;
      RECT  12280.0 2575.0 11865.0 2645.0 ;
      RECT  800.0 21237.5 385.0 21307.5 ;
      RECT  12280.0 21237.5 11865.0 21307.5 ;
      RECT  800.0 23927.5 385.0 23997.5 ;
      RECT  12280.0 23927.5 11865.0 23997.5 ;
      RECT  800.0 26617.5 385.0 26687.5 ;
      RECT  12280.0 26617.5 11865.0 26687.5 ;
      RECT  800.0 29307.5 385.0 29377.5 ;
      RECT  12280.0 29307.5 11865.0 29377.5 ;
      RECT  800.0 31997.5 385.0 32067.5 ;
      RECT  12280.0 31997.5 11865.0 32067.5 ;
      RECT  800.0 34687.5 385.0 34757.5 ;
      RECT  12280.0 34687.5 11865.0 34757.5 ;
      RECT  800.0 37377.5 385.0 37447.5 ;
      RECT  12280.0 37377.5 11865.0 37447.5 ;
      RECT  800.0 40067.5 385.0 40137.5 ;
      RECT  12280.0 40067.5 11865.0 40137.5 ;
      RECT  11895.0 3862.5 11480.0 3932.5 ;
      RECT  11895.0 15287.5 11480.0 15357.5 ;
      RECT  11895.0 4790.0 11480.0 4860.0 ;
      RECT  11895.0 12065.0 11480.0 12135.0 ;
      RECT  415.0 19892.5 -8.881784197e-13 19962.5 ;
      RECT  415.0 22582.5 -8.881784197e-13 22652.5 ;
      RECT  415.0 25272.5 -8.881784197e-13 25342.5 ;
      RECT  415.0 27962.5 -8.881784197e-13 28032.5 ;
      RECT  415.0 30652.5 -8.881784197e-13 30722.5 ;
      RECT  415.0 33342.5 -8.881784197e-13 33412.5 ;
      RECT  415.0 36032.5 -8.881784197e-13 36102.5 ;
      RECT  415.0 38722.5 -8.881784197e-13 38792.5 ;
      RECT  415.0 41412.5 -8.881784197e-13 41482.5 ;
      RECT  10260.0 67.5 10330.0 207.5 ;
      RECT  10965.0 67.5 11035.0 207.5 ;
      RECT  9430.0 67.5 9500.0 44035.0 ;
      RECT  9225.0 67.5 9295.0 44035.0 ;
      RECT  8610.0 67.5 8680.0 44035.0 ;
      RECT  8815.0 67.5 8885.0 44035.0 ;
      RECT  9020.0 67.5 9090.0 44035.0 ;
      RECT  8405.0 67.5 8475.0 44035.0 ;
      RECT  452.5 67.5 732.5 44035.0 ;
      RECT  11932.5 67.5 12212.5 44035.0 ;
      RECT  67.5 67.5 347.5 44035.0 ;
      RECT  11547.5 67.5 11827.5 44035.0 ;
      RECT  -140.0 31017.5 -4175.0 31087.5 ;
      RECT  -140.0 31222.5 -4175.0 31292.5 ;
      RECT  -140.0 31427.5 -4175.0 31497.5 ;
      RECT  -140.0 31837.5 -4175.0 31907.5 ;
      RECT  -752.5 26527.5 -1485.0 26597.5 ;
      RECT  -1655.0 23995.0 -1725.0 30642.5 ;
      RECT  -140.0 30812.5 -345.0 30882.5 ;
      RECT  -1280.0 31632.5 -1485.0 31702.5 ;
      RECT  -2625.0 30812.5 -2830.0 30882.5 ;
      RECT  -3970.0 31632.5 -4175.0 31702.5 ;
      RECT  -4010.0 23757.5 -3305.0 30197.5 ;
      RECT  -2600.0 23757.5 -3305.0 30197.5 ;
      RECT  -2600.0 23757.5 -1895.0 30197.5 ;
      RECT  -3692.5 23757.5 -3622.5 23902.5 ;
      RECT  -2987.5 23757.5 -2917.5 23902.5 ;
      RECT  -2282.5 23757.5 -2212.5 23902.5 ;
      RECT  -3692.5 29927.5 -3622.5 30197.5 ;
      RECT  -3847.5 29510.0 -3777.5 30197.5 ;
      RECT  -2987.5 29927.5 -2917.5 30197.5 ;
      RECT  -2832.5 29510.0 -2762.5 30197.5 ;
      RECT  -2282.5 29927.5 -2212.5 30197.5 ;
      RECT  -2437.5 29510.0 -2367.5 30197.5 ;
      RECT  -4045.0 23757.5 -3975.0 30197.5 ;
      RECT  -3340.0 23757.5 -3270.0 30197.5 ;
      RECT  -2635.0 23757.5 -2565.0 30197.5 ;
      RECT  -1930.0 23757.5 -1860.0 30197.5 ;
      RECT  -437.5 33087.5 -1142.5 33157.5 ;
      RECT  -792.5 32707.5 -862.5 32777.5 ;
      RECT  -792.5 33087.5 -862.5 33157.5 ;
      RECT  -827.5 32707.5 -1142.5 32777.5 ;
      RECT  -792.5 32742.5 -862.5 33122.5 ;
      RECT  -437.5 33087.5 -827.5 33157.5 ;
      RECT  -1142.5 32707.5 -1277.5 32777.5 ;
      RECT  -1142.5 33087.5 -1277.5 33157.5 ;
      RECT  -302.5 33087.5 -437.5 33157.5 ;
      RECT  -760.0 33087.5 -895.0 33157.5 ;
      RECT  -2280.0 32897.5 -2210.0 32967.5 ;
      RECT  -2245.0 32897.5 -1895.0 32967.5 ;
      RECT  -2280.0 32932.5 -2210.0 33002.5 ;
      RECT  -2680.0 32897.5 -2610.0 32967.5 ;
      RECT  -2680.0 32775.0 -2610.0 32932.5 ;
      RECT  -2645.0 32897.5 -2245.0 32967.5 ;
      RECT  -1895.0 32897.5 -1760.0 32967.5 ;
      RECT  -2680.0 32810.0 -2610.0 32675.0 ;
      RECT  -2280.0 33070.0 -2210.0 32935.0 ;
      RECT  -2225.0 33852.5 -2155.0 33922.5 ;
      RECT  -2225.0 34042.5 -2155.0 34112.5 ;
      RECT  -2190.0 33852.5 -1827.5 33922.5 ;
      RECT  -2225.0 33887.5 -2155.0 34077.5 ;
      RECT  -2532.5 34042.5 -2190.0 34112.5 ;
      RECT  -1827.5 33852.5 -1692.5 33922.5 ;
      RECT  -2667.5 34042.5 -2532.5 34112.5 ;
      RECT  -2225.0 34145.0 -2155.0 34010.0 ;
      RECT  -3127.5 33647.5 -3832.5 33717.5 ;
      RECT  -3482.5 33267.5 -3552.5 33337.5 ;
      RECT  -3482.5 33647.5 -3552.5 33717.5 ;
      RECT  -3517.5 33267.5 -3832.5 33337.5 ;
      RECT  -3482.5 33302.5 -3552.5 33682.5 ;
      RECT  -3127.5 33647.5 -3517.5 33717.5 ;
      RECT  -3832.5 33267.5 -3967.5 33337.5 ;
      RECT  -3832.5 33647.5 -3967.5 33717.5 ;
      RECT  -2992.5 33647.5 -3127.5 33717.5 ;
      RECT  -3450.0 33647.5 -3585.0 33717.5 ;
      RECT  -3777.5 30265.0 -3847.5 30130.0 ;
      RECT  -3777.5 31940.0 -3847.5 31805.0 ;
      RECT  -3622.5 30265.0 -3692.5 30130.0 ;
      RECT  -3622.5 31120.0 -3692.5 30985.0 ;
      RECT  -2762.5 30265.0 -2832.5 30130.0 ;
      RECT  -2762.5 31325.0 -2832.5 31190.0 ;
      RECT  -2367.5 30265.0 -2437.5 30130.0 ;
      RECT  -2367.5 31530.0 -2437.5 31395.0 ;
      RECT  -3975.0 30265.0 -4045.0 30130.0 ;
      RECT  -3975.0 30915.0 -4045.0 30780.0 ;
      RECT  -3270.0 30265.0 -3340.0 30130.0 ;
      RECT  -3270.0 30915.0 -3340.0 30780.0 ;
      RECT  -2565.0 30265.0 -2635.0 30130.0 ;
      RECT  -2565.0 30915.0 -2635.0 30780.0 ;
      RECT  -1860.0 30265.0 -1930.0 30130.0 ;
      RECT  -1860.0 30915.0 -1930.0 30780.0 ;
      RECT  -2795.0 36422.5 -2865.0 44172.5 ;
      RECT  -3205.0 36422.5 -3275.0 43862.5 ;
      RECT  -3910.0 36422.5 -3980.0 43862.5 ;
      RECT  -2967.5 36590.0 -3037.5 37187.5 ;
      RECT  -3390.0 36590.0 -3460.0 36870.0 ;
      RECT  -802.5 38985.0 -732.5 39380.0 ;
      RECT  -802.5 39380.0 -732.5 39940.0 ;
      RECT  -802.5 39940.0 -732.5 40500.0 ;
      RECT  -802.5 40665.0 -732.5 41060.0 ;
      RECT  -802.5 41060.0 -732.5 41620.0 ;
      RECT  -802.5 41620.0 -732.5 42180.0 ;
      RECT  -1520.0 42310.0 -1450.0 42380.0 ;
      RECT  -1520.0 41830.0 -1450.0 41900.0 ;
      RECT  -1485.0 42310.0 -767.5 42380.0 ;
      RECT  -1520.0 41865.0 -1450.0 42345.0 ;
      RECT  -2202.5 41830.0 -1485.0 41900.0 ;
      RECT  -2237.5 41305.0 -2167.5 41865.0 ;
      RECT  -2237.5 40745.0 -2167.5 41305.0 ;
      RECT  -2237.5 40185.0 -2167.5 40580.0 ;
      RECT  -2237.5 39625.0 -2167.5 40185.0 ;
      RECT  -2237.5 39065.0 -2167.5 39625.0 ;
      RECT  -835.0 39345.0 -700.0 39415.0 ;
      RECT  -835.0 39905.0 -700.0 39975.0 ;
      RECT  -835.0 40465.0 -700.0 40535.0 ;
      RECT  -835.0 41025.0 -700.0 41095.0 ;
      RECT  -835.0 41585.0 -700.0 41655.0 ;
      RECT  -835.0 42145.0 -700.0 42215.0 ;
      RECT  -2270.0 41830.0 -2135.0 41900.0 ;
      RECT  -2270.0 41270.0 -2135.0 41340.0 ;
      RECT  -2270.0 40710.0 -2135.0 40780.0 ;
      RECT  -2270.0 40150.0 -2135.0 40220.0 ;
      RECT  -2270.0 39590.0 -2135.0 39660.0 ;
      RECT  -2270.0 39030.0 -2135.0 39100.0 ;
      RECT  -835.0 38950.0 -700.0 39020.0 ;
      RECT  -835.0 40630.0 -700.0 40700.0 ;
      RECT  -835.0 42310.0 -700.0 42380.0 ;
      RECT  -2270.0 40545.0 -2135.0 40615.0 ;
      RECT  -3240.0 38327.5 -3950.0 36982.5 ;
      RECT  -3240.0 38327.5 -3945.0 39672.5 ;
      RECT  -3240.0 41017.5 -3945.0 39672.5 ;
      RECT  -3240.0 41017.5 -3945.0 42362.5 ;
      RECT  -3240.0 43707.5 -3945.0 42362.5 ;
      RECT  -3390.0 38227.5 -3460.0 43862.5 ;
      RECT  -3725.0 38227.5 -3795.0 43862.5 ;
      RECT  -3205.0 38227.5 -3275.0 43862.5 ;
      RECT  -3910.0 38227.5 -3980.0 43862.5 ;
      RECT  -2827.5 38400.0 -2897.5 38535.0 ;
      RECT  -2827.5 40810.0 -2897.5 40945.0 ;
      RECT  -2827.5 41090.0 -2897.5 41225.0 ;
      RECT  -2827.5 43500.0 -2897.5 43635.0 ;
      RECT  -2830.0 38662.5 -2900.0 38797.5 ;
      RECT  -2795.0 36287.5 -2865.0 36422.5 ;
      RECT  -3307.5 36387.5 -3172.5 36457.5 ;
      RECT  -4012.5 36387.5 -3877.5 36457.5 ;
      RECT  -3070.0 37152.5 -2935.0 37222.5 ;
      RECT  -3070.0 36555.0 -2935.0 36625.0 ;
      RECT  -3492.5 36555.0 -3357.5 36625.0 ;
      RECT  -717.5 30710.0 -787.5 30575.0 ;
      RECT  -717.5 26630.0 -787.5 26495.0 ;
      RECT  -1450.0 26630.0 -1520.0 26495.0 ;
      RECT  -1450.0 32145.0 -1520.0 32010.0 ;
      RECT  -1655.0 24062.5 -1725.0 23927.5 ;
      RECT  -2210.0 30710.0 -2280.0 30575.0 ;
      RECT  -2425.0 31120.0 -2495.0 30985.0 ;
      RECT  -2155.0 33657.5 -2225.0 33522.5 ;
      RECT  -2155.0 33657.5 -2225.0 33522.5 ;
      RECT  -2155.0 32145.0 -2225.0 32010.0 ;
      RECT  -2370.0 33915.0 -2440.0 33780.0 ;
      RECT  -2370.0 33915.0 -2440.0 33780.0 ;
      RECT  -2370.0 31940.0 -2440.0 31805.0 ;
      RECT  -792.5 32145.0 -862.5 32010.0 ;
      RECT  -652.5 31940.0 -722.5 31805.0 ;
      RECT  -512.5 31325.0 -582.5 31190.0 ;
      RECT  -3482.5 32145.0 -3552.5 32010.0 ;
      RECT  -3342.5 31325.0 -3412.5 31190.0 ;
      RECT  -3202.5 31530.0 -3272.5 31395.0 ;
      RECT  -2177.5 33337.5 -2312.5 33407.5 ;
      RECT  -2122.5 34482.5 -2257.5 34552.5 ;
      RECT  -3390.0 35667.5 -3525.0 35737.5 ;
      RECT  -2135.0 34707.5 -2270.0 34777.5 ;
      RECT  -105.0 30915.0 -175.0 30780.0 ;
      RECT  -1450.0 31735.0 -1520.0 31600.0 ;
      RECT  -2795.0 30915.0 -2865.0 30780.0 ;
      RECT  -4140.0 31735.0 -4210.0 31600.0 ;
      RECT  -140.0 34707.5 -2202.5 34777.5 ;
      RECT  -140.0 35667.5 -3457.5 35737.5 ;
      RECT  -140.0 33337.5 -2245.0 33407.5 ;
      RECT  -140.0 34482.5 -2190.0 34552.5 ;
      RECT  -140.0 32042.5 -4175.0 32112.5 ;
      RECT  -140.0 30607.5 -4175.0 30677.5 ;
      RECT  -140.0 31632.5 -4175.0 31702.5 ;
      RECT  -140.0 30812.5 -4175.0 30882.5 ;
      RECT  9532.5 34707.5 9397.5 34777.5 ;
      RECT  -140.0 34707.5 -275.0 34777.5 ;
      RECT  9327.5 35667.5 9192.5 35737.5 ;
      RECT  -140.0 35667.5 -275.0 35737.5 ;
      RECT  8917.5 33337.5 8782.5 33407.5 ;
      RECT  -140.0 33337.5 -275.0 33407.5 ;
      RECT  8712.5 34482.5 8577.5 34552.5 ;
      RECT  -140.0 34482.5 -275.0 34552.5 ;
      RECT  9122.5 32042.5 8987.5 32112.5 ;
      RECT  -140.0 32042.5 -275.0 32112.5 ;
      RECT  8507.5 30607.5 8372.5 30677.5 ;
      RECT  -140.0 30607.5 -275.0 30677.5 ;
      RECT  660.0 31632.5 525.0 31702.5 ;
      RECT  -140.0 31632.5 -275.0 31702.5 ;
   LAYER  metal3 ;
      RECT  -140.0 34707.5 9465.0 34777.5 ;
      RECT  -140.0 35667.5 9260.0 35737.5 ;
      RECT  -140.0 33337.5 8850.0 33407.5 ;
      RECT  -140.0 34482.5 8645.0 34552.5 ;
      RECT  -140.0 32042.5 9055.0 32112.5 ;
      RECT  -140.0 30607.5 8440.0 30677.5 ;
      RECT  -140.0 31632.5 592.5 31702.5 ;
      RECT  10050.0 19822.5 10120.0 19892.5 ;
      RECT  10050.0 1312.5 10120.0 19857.5 ;
      RECT  10085.0 19822.5 10255.0 19892.5 ;
      RECT  10755.0 19822.5 10825.0 19892.5 ;
      RECT  10755.0 1312.5 10825.0 19857.5 ;
      RECT  10790.0 19822.5 10960.0 19892.5 ;
      RECT  10260.0 67.5 10330.0 4427.5 ;
      RECT  10965.0 67.5 11035.0 4427.5 ;
      RECT  10255.0 19787.5 10325.0 19927.5 ;
      RECT  10960.0 19787.5 11030.0 19927.5 ;
      RECT  10260.0 4427.5 10330.0 4567.5 ;
      RECT  10965.0 4427.5 11035.0 4567.5 ;
      RECT  837.5 8440.0 977.5 8370.0 ;
      RECT  837.5 7735.0 977.5 7665.0 ;
      RECT  837.5 7030.0 977.5 6960.0 ;
      RECT  837.5 6325.0 977.5 6255.0 ;
      RECT  10050.0 1277.5 10120.0 1412.5 ;
      RECT  10755.0 1277.5 10825.0 1412.5 ;
      RECT  10260.0 67.5 10330.0 202.5 ;
      RECT  10965.0 67.5 11035.0 202.5 ;
      RECT  67.5 8370.0 837.5 8440.0 ;
      RECT  67.5 7665.0 837.5 7735.0 ;
      RECT  67.5 6960.0 837.5 7030.0 ;
      RECT  67.5 6255.0 837.5 6325.0 ;
      RECT  -3777.5 30197.5 -3847.5 31872.5 ;
      RECT  -3622.5 30197.5 -3692.5 31052.5 ;
      RECT  -2762.5 30197.5 -2832.5 31257.5 ;
      RECT  -2367.5 30197.5 -2437.5 31462.5 ;
      RECT  -3975.0 30197.5 -4045.0 30847.5 ;
      RECT  -3270.0 30197.5 -3340.0 30847.5 ;
      RECT  -2565.0 30197.5 -2635.0 30847.5 ;
      RECT  -1860.0 30197.5 -1930.0 30847.5 ;
      RECT  -1450.0 26562.5 -1520.0 32077.5 ;
      RECT  -2155.0 32077.5 -2225.0 33590.0 ;
      RECT  -2370.0 31872.5 -2440.0 33847.5 ;
      RECT  -3692.5 23757.5 -3622.5 23897.5 ;
      RECT  -2987.5 23757.5 -2917.5 23897.5 ;
      RECT  -2282.5 23757.5 -2212.5 23897.5 ;
      RECT  -3777.5 30265.0 -3847.5 30130.0 ;
      RECT  -3777.5 31940.0 -3847.5 31805.0 ;
      RECT  -3622.5 30265.0 -3692.5 30130.0 ;
      RECT  -3622.5 31120.0 -3692.5 30985.0 ;
      RECT  -2762.5 30265.0 -2832.5 30130.0 ;
      RECT  -2762.5 31325.0 -2832.5 31190.0 ;
      RECT  -2367.5 30265.0 -2437.5 30130.0 ;
      RECT  -2367.5 31530.0 -2437.5 31395.0 ;
      RECT  -3975.0 30265.0 -4045.0 30130.0 ;
      RECT  -3975.0 30915.0 -4045.0 30780.0 ;
      RECT  -3270.0 30265.0 -3340.0 30130.0 ;
      RECT  -3270.0 30915.0 -3340.0 30780.0 ;
      RECT  -2565.0 30265.0 -2635.0 30130.0 ;
      RECT  -2565.0 30915.0 -2635.0 30780.0 ;
      RECT  -1860.0 30265.0 -1930.0 30130.0 ;
      RECT  -1860.0 30915.0 -1930.0 30780.0 ;
      RECT  -1450.0 26630.0 -1520.0 26495.0 ;
      RECT  -1450.0 32145.0 -1520.0 32010.0 ;
      RECT  -2155.0 33657.5 -2225.0 33522.5 ;
      RECT  -2155.0 32145.0 -2225.0 32010.0 ;
      RECT  -2370.0 33915.0 -2440.0 33780.0 ;
      RECT  -2370.0 31940.0 -2440.0 31805.0 ;
      RECT  -2917.5 23757.5 -2987.5 23897.5 ;
      RECT  -2212.5 23757.5 -2282.5 23897.5 ;
      RECT  -3622.5 23757.5 -3692.5 23897.5 ;
      RECT  9532.5 34707.5 9397.5 34777.5 ;
      RECT  -140.0 34707.5 -275.0 34777.5 ;
      RECT  9327.5 35667.5 9192.5 35737.5 ;
      RECT  -140.0 35667.5 -275.0 35737.5 ;
      RECT  8917.5 33337.5 8782.5 33407.5 ;
      RECT  -140.0 33337.5 -275.0 33407.5 ;
      RECT  8712.5 34482.5 8577.5 34552.5 ;
      RECT  -140.0 34482.5 -275.0 34552.5 ;
      RECT  9122.5 32042.5 8987.5 32112.5 ;
      RECT  -140.0 32042.5 -275.0 32112.5 ;
      RECT  8507.5 30607.5 8372.5 30677.5 ;
      RECT  -140.0 30607.5 -275.0 30677.5 ;
      RECT  660.0 31632.5 525.0 31702.5 ;
      RECT  -140.0 31632.5 -275.0 31702.5 ;
   END
   END    sram_2_16_1_freepdk45
END    LIBRARY
