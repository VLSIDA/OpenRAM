magic
tech sky130A
magscale 1 2
timestamp 1595931502
<< checkpaint >>
rect -1319 -1316 1577 1566
<< nwell >>
rect -54 -54 312 306
<< scpmos >>
rect 60 0 90 252
rect 168 0 198 252
<< pdiff >>
rect 0 0 60 252
rect 90 0 168 252
rect 198 0 258 252
<< poly >>
rect 60 252 90 278
rect 168 252 198 278
rect 60 -26 90 0
rect 168 -26 198 0
rect 60 -56 198 -26
<< locali >>
rect 8 93 42 159
rect 112 93 146 159
rect 216 93 250 159
use contact_11  contact_11_2
timestamp 1595931502
transform 1 0 0 0 1 93
box -59 -51 109 117
use contact_11  contact_11_1
timestamp 1595931502
transform 1 0 104 0 1 93
box -59 -51 109 117
use contact_11  contact_11_0
timestamp 1595931502
transform 1 0 208 0 1 93
box -59 -51 109 117
<< labels >>
rlabel poly s 129 -41 129 -41 4 G
rlabel corelocali s 233 126 233 126 4 S
rlabel corelocali s 25 126 25 126 4 S
rlabel corelocali s 129 126 129 126 4 D
<< properties >>
string FIXED_BBOX -54 -54 312 306
<< end >>
