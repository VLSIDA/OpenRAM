magic
tech sky130A
magscale 1 2
timestamp 1595931502
<< checkpaint >>
rect -1309 -1311 31567 29327
<< metal1 >>
rect 5632 14266 5660 22347
rect 5712 14266 5740 23905
rect 5792 14266 5820 25175
rect 5872 14266 5900 26733
rect 14720 22632 14766 22886
rect 15590 22632 15636 22886
rect 14720 7958 14766 8212
rect 15590 7958 15636 8212
rect 24580 4111 24608 14266
rect 24660 5669 24688 14266
rect 24740 6939 24768 14266
rect 24820 8497 24848 14266
<< metal2 >>
rect 30055 27426 30121 27478
rect 25020 27311 25118 27339
rect 27227 27333 27255 27361
rect 4415 26778 4481 26830
rect 5858 26709 5914 26757
rect 5778 25151 5834 25199
rect 4415 25078 4481 25130
rect 4415 23950 4481 24002
rect 5698 23881 5754 23929
rect 17236 22956 17264 23067
rect 5618 22323 5674 22371
rect 4415 22250 4481 22302
rect 1748 10342 1776 11994
rect 5516 2881 5544 22020
rect 17360 21691 17388 22984
rect 17484 18728 17512 20213
rect 12748 10631 12776 12116
rect 25020 8824 25048 27311
rect 28482 18850 28510 20502
rect 26083 8542 26149 8594
rect 24806 8473 24862 8521
rect 12872 5681 12900 6363
rect 12996 5681 13024 7815
rect 24726 6915 24782 6963
rect 26083 6842 26149 6894
rect 26083 5714 26149 5766
rect 13120 4949 13148 5709
rect 24646 5645 24702 5693
rect 24566 4087 24622 4135
rect 26083 4014 26149 4066
rect 6751 3111 6817 3163
rect 7919 3111 7985 3163
rect 137 2238 203 2290
rect 5493 721 5567 2881
rect 5446 707 5567 721
rect 5446 693 5544 707
rect 3087 655 3115 683
rect 137 538 203 590
<< metal3 >>
rect 25153 27967 25251 28065
rect 30209 27969 30307 28067
rect 4813 27319 4911 27417
rect 5393 26703 5886 26763
rect 25153 26553 25251 26651
rect 30209 26553 30307 26651
rect 4813 25905 4911 26003
rect 5393 25145 5806 25205
rect 25153 25139 25251 25237
rect 4813 24491 4911 24589
rect 5393 23875 5726 23935
rect 25153 23725 25251 23823
rect 4813 23077 4911 23175
rect 17250 23037 25118 23097
rect 14948 22729 15046 22827
rect 15310 22729 15408 22827
rect 14948 22407 15046 22505
rect 15310 22407 15408 22505
rect 5393 22317 5646 22377
rect 25153 22311 25251 22409
rect 5446 21983 5530 22057
rect 4813 21663 4911 21761
rect 399 21503 497 21601
rect 1135 21503 1233 21601
rect 14936 21569 15034 21667
rect 15322 21569 15420 21667
rect 17374 21661 25118 21721
rect 25153 20897 25251 20995
rect 15018 20795 15116 20893
rect 15240 20795 15338 20893
rect 399 20383 497 20481
rect 1135 20383 1233 20481
rect 24950 20472 28496 20532
rect 17498 20183 25118 20243
rect 14760 19685 14858 19783
rect 15622 19685 15720 19783
rect 16008 19685 16106 19783
rect 25153 19483 25251 19581
rect 399 19263 497 19361
rect 1135 19263 1233 19361
rect 29025 19323 29123 19421
rect 29761 19323 29859 19421
rect 14255 19094 14353 19192
rect 14898 19113 14958 19173
rect 15522 19113 15582 19173
rect 16127 19094 16225 19192
rect 13578 18789 13638 18849
rect 16842 18789 16902 18849
rect 13578 18552 13638 18612
rect 16842 18552 16902 18612
rect 13578 18315 13638 18375
rect 16842 18315 16902 18375
rect 399 18143 497 18241
rect 1135 18143 1233 18241
rect 9833 18174 9931 18272
rect 10258 18174 10356 18272
rect 10637 18167 10735 18265
rect 10909 18167 11007 18265
rect 19473 18167 19571 18265
rect 19745 18167 19843 18265
rect 20124 18174 20222 18272
rect 20549 18174 20647 18272
rect 29025 18203 29123 18301
rect 29761 18203 29859 18301
rect 13578 17999 13638 18059
rect 16842 17999 16902 18059
rect 9833 17802 9931 17900
rect 10258 17804 10356 17902
rect 10637 17772 10735 17870
rect 10909 17772 11007 17870
rect 13578 17762 13638 17822
rect 16842 17762 16902 17822
rect 19473 17772 19571 17870
rect 19745 17772 19843 17870
rect 20124 17804 20222 17902
rect 20549 17802 20647 17900
rect 13578 17525 13638 17585
rect 16842 17525 16902 17585
rect 9833 17384 9931 17482
rect 10258 17384 10356 17482
rect 10637 17377 10735 17475
rect 10909 17377 11007 17475
rect 19473 17377 19571 17475
rect 19745 17377 19843 17475
rect 20124 17384 20222 17482
rect 20549 17384 20647 17482
rect 13578 17209 13638 17269
rect 16842 17209 16902 17269
rect 399 17023 497 17121
rect 1135 17023 1233 17121
rect 9833 17012 9931 17110
rect 10258 17014 10356 17112
rect 10637 16982 10735 17080
rect 10909 16982 11007 17080
rect 13578 16972 13638 17032
rect 16842 16972 16902 17032
rect 19473 16982 19571 17080
rect 19745 16982 19843 17080
rect 20124 17014 20222 17112
rect 20549 17012 20647 17110
rect 29025 17083 29123 17181
rect 29761 17083 29859 17181
rect 13578 16735 13638 16795
rect 16842 16735 16902 16795
rect 9833 16594 9931 16692
rect 10258 16594 10356 16692
rect 10637 16587 10735 16685
rect 10909 16587 11007 16685
rect 19473 16587 19571 16685
rect 19745 16587 19843 16685
rect 20124 16594 20222 16692
rect 20549 16594 20647 16692
rect 13578 16419 13638 16479
rect 16842 16419 16902 16479
rect 9833 16222 9931 16320
rect 10258 16224 10356 16322
rect 10637 16192 10735 16290
rect 10909 16192 11007 16290
rect 13578 16182 13638 16242
rect 16842 16182 16902 16242
rect 19473 16192 19571 16290
rect 19745 16192 19843 16290
rect 20124 16224 20222 16322
rect 20549 16222 20647 16320
rect 399 15903 497 16001
rect 1135 15903 1233 16001
rect 13578 15945 13638 16005
rect 16842 15945 16902 16005
rect 29025 15963 29123 16061
rect 29761 15963 29859 16061
rect 7619 15804 7717 15902
rect 8044 15804 8142 15902
rect 8423 15797 8521 15895
rect 8695 15797 8793 15895
rect 9833 15804 9931 15902
rect 10258 15804 10356 15902
rect 10637 15797 10735 15895
rect 10909 15797 11007 15895
rect 19473 15797 19571 15895
rect 19745 15797 19843 15895
rect 20124 15804 20222 15902
rect 20549 15804 20647 15902
rect 21687 15797 21785 15895
rect 21959 15797 22057 15895
rect 22338 15804 22436 15902
rect 22763 15804 22861 15902
rect 13578 15629 13638 15689
rect 16842 15629 16902 15689
rect 9833 15432 9931 15530
rect 10258 15434 10356 15532
rect 10637 15402 10735 15500
rect 10909 15402 11007 15500
rect 11355 15358 11453 15456
rect 11780 15357 11878 15455
rect 12197 15373 12295 15471
rect 12695 15373 12793 15471
rect 13578 15392 13638 15452
rect 16842 15392 16902 15452
rect 17687 15373 17785 15471
rect 18185 15373 18283 15471
rect 18602 15357 18700 15455
rect 19027 15358 19125 15456
rect 19473 15402 19571 15500
rect 19745 15402 19843 15500
rect 20124 15434 20222 15532
rect 20549 15432 20647 15530
rect 13578 15155 13638 15215
rect 16842 15155 16902 15215
rect 6449 15007 6547 15105
rect 6721 15007 6819 15105
rect 7619 15014 7717 15112
rect 8044 15014 8142 15112
rect 8423 15007 8521 15105
rect 8695 15007 8793 15105
rect 9833 15014 9931 15112
rect 10258 15014 10356 15112
rect 10637 15007 10735 15105
rect 10909 15007 11007 15105
rect 19473 15007 19571 15105
rect 19745 15007 19843 15105
rect 20124 15014 20222 15112
rect 20549 15014 20647 15112
rect 21687 15007 21785 15105
rect 21959 15007 22057 15105
rect 22338 15014 22436 15112
rect 22763 15014 22861 15112
rect 23661 15007 23759 15105
rect 23933 15007 24031 15105
rect 399 14783 497 14881
rect 1135 14783 1233 14881
rect 13578 14839 13638 14899
rect 16842 14839 16902 14899
rect 29025 14843 29123 14941
rect 29761 14843 29859 14941
rect 9833 14642 9931 14740
rect 10258 14644 10356 14742
rect 10637 14612 10735 14710
rect 10909 14612 11007 14710
rect 13578 14602 13638 14662
rect 16842 14602 16902 14662
rect 19473 14612 19571 14710
rect 19745 14612 19843 14710
rect 20124 14644 20222 14742
rect 20549 14642 20647 14740
rect 13578 14365 13638 14425
rect 16842 14365 16902 14425
rect 9833 14224 9931 14322
rect 10258 14224 10356 14322
rect 10637 14217 10735 14315
rect 10909 14217 11007 14315
rect 19473 14217 19571 14315
rect 19745 14217 19843 14315
rect 20124 14224 20222 14322
rect 20549 14224 20647 14322
rect 13578 14049 13638 14109
rect 16842 14049 16902 14109
rect 9833 13852 9931 13950
rect 10258 13854 10356 13952
rect 10637 13822 10735 13920
rect 10909 13822 11007 13920
rect 13578 13812 13638 13872
rect 16842 13812 16902 13872
rect 19473 13822 19571 13920
rect 19745 13822 19843 13920
rect 20124 13854 20222 13952
rect 20549 13852 20647 13950
rect 399 13663 497 13761
rect 1135 13663 1233 13761
rect 29025 13723 29123 13821
rect 29761 13723 29859 13821
rect 13578 13575 13638 13635
rect 16842 13575 16902 13635
rect 7619 13434 7717 13532
rect 8044 13434 8142 13532
rect 8423 13427 8521 13525
rect 8695 13427 8793 13525
rect 9833 13434 9931 13532
rect 10258 13434 10356 13532
rect 10637 13427 10735 13525
rect 10909 13427 11007 13525
rect 19473 13427 19571 13525
rect 19745 13427 19843 13525
rect 20124 13434 20222 13532
rect 20549 13434 20647 13532
rect 21687 13427 21785 13525
rect 21959 13427 22057 13525
rect 22338 13434 22436 13532
rect 22763 13434 22861 13532
rect 13578 13259 13638 13319
rect 16842 13259 16902 13319
rect 9833 13062 9931 13160
rect 10258 13064 10356 13162
rect 10637 13032 10735 13130
rect 10909 13032 11007 13130
rect 13578 13022 13638 13082
rect 16842 13022 16902 13082
rect 19473 13032 19571 13130
rect 19745 13032 19843 13130
rect 20124 13064 20222 13162
rect 20549 13062 20647 13160
rect 13578 12785 13638 12845
rect 16842 12785 16902 12845
rect 399 12543 497 12641
rect 1135 12543 1233 12641
rect 6449 12637 6547 12735
rect 6721 12637 6819 12735
rect 7619 12644 7717 12742
rect 8044 12644 8142 12742
rect 8423 12637 8521 12735
rect 8695 12637 8793 12735
rect 9833 12644 9931 12742
rect 10258 12644 10356 12742
rect 10637 12637 10735 12735
rect 10909 12637 11007 12735
rect 19473 12637 19571 12735
rect 19745 12637 19843 12735
rect 20124 12644 20222 12742
rect 20549 12644 20647 12742
rect 21687 12637 21785 12735
rect 21959 12637 22057 12735
rect 22338 12644 22436 12742
rect 22763 12644 22861 12742
rect 23661 12637 23759 12735
rect 23933 12637 24031 12735
rect 29025 12603 29123 12701
rect 29761 12603 29859 12701
rect 13578 12469 13638 12529
rect 16842 12469 16902 12529
rect 13578 12232 13638 12292
rect 16842 12232 16902 12292
rect 13578 11995 13638 12055
rect 16842 11995 16902 12055
rect 14255 11652 14353 11750
rect 14898 11671 14958 11731
rect 15522 11671 15582 11731
rect 16127 11652 16225 11750
rect 399 11423 497 11521
rect 1135 11423 1233 11521
rect 29025 11483 29123 11581
rect 29761 11483 29859 11581
rect 5313 11263 5411 11361
rect 14374 11061 14472 11159
rect 14760 11061 14858 11159
rect 15622 11061 15720 11159
rect 5446 10601 12762 10661
rect 1762 10312 14536 10372
rect 29025 10363 29123 10461
rect 29761 10363 29859 10461
rect 15018 9951 15116 10049
rect 15240 9951 15338 10049
rect 5313 9849 5411 9947
rect 14936 9177 15034 9275
rect 15322 9177 15420 9275
rect 29025 9243 29123 9341
rect 29761 9243 29859 9341
rect 25653 9083 25751 9181
rect 25034 8787 25118 8861
rect 5313 8435 5411 8533
rect 24834 8467 25171 8527
rect 14948 8339 15046 8437
rect 15310 8339 15408 8437
rect 14948 8017 15046 8115
rect 15310 8017 15408 8115
rect 5446 7785 13010 7845
rect 25653 7669 25751 7767
rect 14834 7224 14932 7322
rect 15424 7224 15522 7322
rect 5313 7021 5411 7119
rect 24754 6909 25171 6969
rect 14823 6787 14921 6885
rect 15435 6787 15533 6885
rect 14944 6455 15042 6553
rect 15314 6455 15412 6553
rect 5446 6333 12886 6393
rect 14829 6253 14927 6351
rect 15429 6253 15527 6351
rect 25653 6255 25751 6353
rect 14843 5837 14941 5935
rect 15415 5837 15513 5935
rect 5313 5607 5411 5705
rect 24674 5639 25171 5699
rect 5446 4919 13134 4979
rect 25653 4841 25751 4939
rect 5313 4193 5411 4291
rect 24594 4081 25171 4141
rect 7149 3938 7247 4036
rect 8317 3938 8415 4036
rect 25653 3427 25751 3525
rect -49 2781 49 2879
rect 5313 2779 5411 2877
rect 5530 2851 7782 2911
rect 7149 2524 7247 2622
rect 8317 2524 8415 2622
rect -49 1365 49 1463
rect 5313 1365 5411 1463
rect -49 -51 49 47
rect 5313 -49 5411 49
use contact_9  contact_9_31
timestamp 1595931502
transform 1 0 5413 0 1 10594
box 0 0 66 74
use contact_9  contact_9_30
timestamp 1595931502
transform 1 0 12729 0 1 10594
box 0 0 66 74
use contact_9  contact_9_29
timestamp 1595931502
transform 1 0 5413 0 1 6326
box 0 0 66 74
use contact_9  contact_9_28
timestamp 1595931502
transform 1 0 12853 0 1 6326
box 0 0 66 74
use contact_9  contact_9_27
timestamp 1595931502
transform 1 0 5413 0 1 7778
box 0 0 66 74
use contact_9  contact_9_26
timestamp 1595931502
transform 1 0 12977 0 1 7778
box 0 0 66 74
use contact_9  contact_9_25
timestamp 1595931502
transform 1 0 5413 0 1 4912
box 0 0 66 74
use contact_9  contact_9_24
timestamp 1595931502
transform 1 0 13101 0 1 4912
box 0 0 66 74
use contact_9  contact_9_23
timestamp 1595931502
transform 1 0 25085 0 1 20176
box 0 0 66 74
use contact_9  contact_9_22
timestamp 1595931502
transform 1 0 17465 0 1 20176
box 0 0 66 74
use contact_9  contact_9_21
timestamp 1595931502
transform 1 0 25085 0 1 21654
box 0 0 66 74
use contact_9  contact_9_20
timestamp 1595931502
transform 1 0 17341 0 1 21654
box 0 0 66 74
use contact_9  contact_9_19
timestamp 1595931502
transform 1 0 25085 0 1 23030
box 0 0 66 74
use contact_9  contact_9_18
timestamp 1595931502
transform 1 0 17217 0 1 23030
box 0 0 66 74
use contact_9  contact_9_17
timestamp 1595931502
transform 1 0 10042 0 1 10305
box 0 0 66 74
use contact_9  contact_9_16
timestamp 1595931502
transform 1 0 20414 0 1 20465
box 0 0 66 74
use contact_9  contact_9_15
timestamp 1595931502
transform 1 0 5360 0 1 22310
box 0 0 66 74
use contact_9  contact_9_14
timestamp 1595931502
transform 1 0 5613 0 1 22310
box 0 0 66 74
use contact_9  contact_9_13
timestamp 1595931502
transform 1 0 5360 0 1 23868
box 0 0 66 74
use contact_9  contact_9_12
timestamp 1595931502
transform 1 0 5693 0 1 23868
box 0 0 66 74
use contact_9  contact_9_11
timestamp 1595931502
transform 1 0 5360 0 1 25138
box 0 0 66 74
use contact_9  contact_9_10
timestamp 1595931502
transform 1 0 5773 0 1 25138
box 0 0 66 74
use contact_9  contact_9_9
timestamp 1595931502
transform 1 0 5360 0 1 26696
box 0 0 66 74
use contact_9  contact_9_8
timestamp 1595931502
transform 1 0 5853 0 1 26696
box 0 0 66 74
use contact_9  contact_9_7
timestamp 1595931502
transform 1 0 25138 0 1 8460
box 0 0 66 74
use contact_9  contact_9_6
timestamp 1595931502
transform 1 0 24801 0 1 8460
box 0 0 66 74
use contact_9  contact_9_5
timestamp 1595931502
transform 1 0 25138 0 1 6902
box 0 0 66 74
use contact_9  contact_9_4
timestamp 1595931502
transform 1 0 24721 0 1 6902
box 0 0 66 74
use contact_9  contact_9_3
timestamp 1595931502
transform 1 0 25138 0 1 5632
box 0 0 66 74
use contact_9  contact_9_2
timestamp 1595931502
transform 1 0 24641 0 1 5632
box 0 0 66 74
use contact_9  contact_9_1
timestamp 1595931502
transform 1 0 25138 0 1 4074
box 0 0 66 74
use contact_9  contact_9_0
timestamp 1595931502
transform 1 0 24561 0 1 4074
box 0 0 66 74
use cr_0  cr_0_0
timestamp 1595931502
transform 1 0 5614 0 1 5695
box 2083 -2475 9873 36
use control_logic_r  control_logic_r_0
timestamp 1595931502
transform -1 0 30258 0 -1 28016
box -49 -51 5140 18781
use control_logic_rw  control_logic_rw_0
timestamp 1595931502
transform 1 0 0 0 1 0
box -49 -51 5446 21609
use row_addr_dff  row_addr_dff_1
timestamp 1595931502
transform 1 0 4278 0 1 21712
box -8 -49 1176 5705
use row_addr_dff  row_addr_dff_0
timestamp 1595931502
transform -1 0 26286 0 -1 9132
box -8 -49 1176 5705
use contact_8  contact_8_7
timestamp 1595931502
transform 1 0 5614 0 1 22315
box 0 0 64 64
use contact_8  contact_8_6
timestamp 1595931502
transform 1 0 5694 0 1 23873
box 0 0 64 64
use contact_8  contact_8_5
timestamp 1595931502
transform 1 0 5774 0 1 25143
box 0 0 64 64
use contact_8  contact_8_4
timestamp 1595931502
transform 1 0 5854 0 1 26701
box 0 0 64 64
use contact_8  contact_8_3
timestamp 1595931502
transform 1 0 24802 0 1 8465
box 0 0 64 64
use contact_8  contact_8_2
timestamp 1595931502
transform 1 0 24722 0 1 6907
box 0 0 64 64
use contact_8  contact_8_1
timestamp 1595931502
transform 1 0 24642 0 1 5637
box 0 0 64 64
use contact_8  contact_8_0
timestamp 1595931502
transform 1 0 24562 0 1 4079
box 0 0 64 64
use bank  bank_0
timestamp 1595931502
transform 1 0 5614 0 1 5695
box 0 0 19336 17275
use contact_27  contact_27_4
timestamp 1595931502
transform 1 0 5497 0 1 21983
box 0 0 66 74
use contact_27  contact_27_3
timestamp 1595931502
transform 1 0 5497 0 1 2844
box 0 0 66 74
use contact_27  contact_27_2
timestamp 1595931502
transform 1 0 25001 0 1 8787
box 0 0 66 74
use contact_27  contact_27_1
timestamp 1595931502
transform 1 0 1729 0 1 10305
box 0 0 66 74
use contact_27  contact_27_0
timestamp 1595931502
transform 1 0 28463 0 1 20465
box 0 0 66 74
use data_dff  data_dff_0
timestamp 1595931502
transform 1 0 6614 0 1 2573
box -8 -49 2344 1467
<< labels >>
rlabel metal2 s 4572 10631 4572 10631 4 s_en
rlabel metal2 s 4680 6363 4680 6363 4 w_en
rlabel metal2 s 4749 7815 4749 7815 4 p_en_bar
rlabel metal2 s 4882 4949 4882 4949 4 wl_en
rlabel metal2 s 5155 707 5155 707 4 clk_buf
rlabel metal2 s 7952 3137 7952 3137 4 din0[1]
rlabel metal2 s 4448 25104 4448 25104 4 addr0[2]
rlabel metal1 s 15613 8085 15613 8085 4 dout0[1]
rlabel metal1 s 14743 22759 14743 22759 4 dout1[0]
rlabel metal2 s 3101 669 3101 669 4 clk0
rlabel metal2 s 4448 22276 4448 22276 4 addr0[0]
rlabel metal1 s 14743 8085 14743 8085 4 dout0[0]
rlabel metal2 s 1762 11733 1762 11733 4 rbl_bl0
rlabel metal2 s 170 564 170 564 4 csb0
rlabel metal2 s 6784 3137 6784 3137 4 din0[0]
rlabel metal3 s 16872 16765 16872 16765 4 gnd
rlabel metal3 s 19794 15451 19794 15451 4 gnd
rlabel metal3 s 23982 12686 23982 12686 4 gnd
rlabel metal3 s 10686 13871 10686 13871 4 gnd
rlabel metal3 s 9882 17851 9882 17851 4 gnd
rlabel metal3 s 23982 15056 23982 15056 4 gnd
rlabel metal3 s 22812 15853 22812 15853 4 gnd
rlabel metal3 s 14997 22778 14997 22778 4 gnd
rlabel metal3 s 22812 15063 22812 15063 4 gnd
rlabel metal3 s 20598 17061 20598 17061 4 gnd
rlabel metal3 s 15363 6504 15363 6504 4 gnd
rlabel metal3 s 16872 13289 16872 13289 4 gnd
rlabel metal3 s 10686 14661 10686 14661 4 gnd
rlabel metal3 s 16872 17002 16872 17002 4 gnd
rlabel metal3 s 22812 13483 22812 13483 4 gnd
rlabel metal3 s 5362 0 5362 0 4 gnd
rlabel metal3 s 19794 17821 19794 17821 4 gnd
rlabel metal3 s 25202 19532 25202 19532 4 gnd
rlabel metal3 s 9882 18223 9882 18223 4 gnd
rlabel metal3 s 10686 15846 10686 15846 4 gnd
rlabel metal3 s 8472 15846 8472 15846 4 gnd
rlabel metal3 s 9882 14273 9882 14273 4 gnd
rlabel metal3 s 20598 15853 20598 15853 4 gnd
rlabel metal3 s 9882 17433 9882 17433 4 gnd
rlabel metal3 s 22008 15846 22008 15846 4 gnd
rlabel metal3 s 12246 15422 12246 15422 4 gnd
rlabel metal3 s 448 15952 448 15952 4 gnd
rlabel metal3 s 16872 14395 16872 14395 4 gnd
rlabel metal3 s 20598 13901 20598 13901 4 gnd
rlabel metal3 s 16872 15659 16872 15659 4 gnd
rlabel metal3 s 19794 13476 19794 13476 4 gnd
rlabel metal3 s 16872 12815 16872 12815 4 gnd
rlabel metal3 s 6498 12686 6498 12686 4 gnd
rlabel metal3 s 25202 25188 25202 25188 4 gnd
rlabel metal3 s 15067 10000 15067 10000 4 gnd
rlabel metal3 s 20598 13111 20598 13111 4 gnd
rlabel metal3 s 19794 15056 19794 15056 4 gnd
rlabel metal3 s 16872 12499 16872 12499 4 gnd
rlabel metal3 s 9882 17061 9882 17061 4 gnd
rlabel metal3 s 10686 12686 10686 12686 4 gnd
rlabel metal3 s 14878 6302 14878 6302 4 gnd
rlabel metal3 s 7668 13483 7668 13483 4 gnd
rlabel metal3 s 448 13712 448 13712 4 gnd
rlabel metal3 s 20598 15481 20598 15481 4 gnd
rlabel metal3 s 11404 15407 11404 15407 4 gnd
rlabel metal3 s 19794 12686 19794 12686 4 gnd
rlabel metal3 s 10686 17031 10686 17031 4 gnd
rlabel metal3 s 15289 10000 15289 10000 4 gnd
rlabel metal3 s 30258 28018 30258 28018 4 gnd
rlabel metal3 s 9882 12693 9882 12693 4 gnd
rlabel metal3 s 20598 17433 20598 17433 4 gnd
rlabel metal3 s 29074 17132 29074 17132 4 gnd
rlabel metal3 s 19794 17031 19794 17031 4 gnd
rlabel metal3 s 29810 17132 29810 17132 4 gnd
rlabel metal3 s 16872 16212 16872 16212 4 gnd
rlabel metal3 s 13608 13842 13608 13842 4 gnd
rlabel metal3 s 13608 18582 13608 18582 4 gnd
rlabel metal3 s 9882 15853 9882 15853 4 gnd
rlabel metal3 s 29074 14892 29074 14892 4 gnd
rlabel metal3 s 29074 12652 29074 12652 4 gnd
rlabel metal3 s 1184 18192 1184 18192 4 gnd
rlabel metal3 s 16872 17239 16872 17239 4 gnd
rlabel metal3 s 16872 15422 16872 15422 4 gnd
rlabel metal3 s 13608 15659 13608 15659 4 gnd
rlabel metal3 s 13608 14632 13608 14632 4 gnd
rlabel metal3 s 14883 7273 14883 7273 4 gnd
rlabel metal3 s 5362 11312 5362 11312 4 gnd
rlabel metal3 s 9882 13901 9882 13901 4 gnd
rlabel metal3 s 16872 16449 16872 16449 4 gnd
rlabel metal3 s 7668 15063 7668 15063 4 gnd
rlabel metal3 s 16872 13052 16872 13052 4 gnd
rlabel metal3 s 9882 15481 9882 15481 4 gnd
rlabel metal3 s 448 11472 448 11472 4 gnd
rlabel metal3 s 29074 19372 29074 19372 4 gnd
rlabel metal3 s 19076 15407 19076 15407 4 gnd
rlabel metal3 s 13608 12262 13608 12262 4 gnd
rlabel metal3 s 4862 24540 4862 24540 4 gnd
rlabel metal3 s 19794 14661 19794 14661 4 gnd
rlabel metal3 s 13608 18819 13608 18819 4 gnd
rlabel metal3 s 13608 16449 13608 16449 4 gnd
rlabel metal3 s 16872 14632 16872 14632 4 gnd
rlabel metal3 s 20598 15063 20598 15063 4 gnd
rlabel metal3 s 16872 14079 16872 14079 4 gnd
rlabel metal3 s 25702 3476 25702 3476 4 gnd
rlabel metal3 s 13608 16765 13608 16765 4 gnd
rlabel metal3 s 13608 16212 13608 16212 4 gnd
rlabel metal3 s 13608 13289 13608 13289 4 gnd
rlabel metal3 s 8472 12686 8472 12686 4 gnd
rlabel metal3 s 8366 2573 8366 2573 4 gnd
rlabel metal3 s 22008 15056 22008 15056 4 gnd
rlabel metal3 s 19794 16636 19794 16636 4 gnd
rlabel metal3 s 16872 18819 16872 18819 4 gnd
rlabel metal3 s 13608 17792 13608 17792 4 gnd
rlabel metal3 s 18234 15422 18234 15422 4 gnd
rlabel metal3 s 4862 21712 4862 21712 4 gnd
rlabel metal3 s 10686 18216 10686 18216 4 gnd
rlabel metal3 s 1184 15952 1184 15952 4 gnd
rlabel metal3 s 10686 17821 10686 17821 4 gnd
rlabel metal3 s 19794 14266 19794 14266 4 gnd
rlabel metal3 s 5362 5656 5362 5656 4 gnd
rlabel metal3 s 16872 18029 16872 18029 4 gnd
rlabel metal3 s 19794 16241 19794 16241 4 gnd
rlabel metal3 s 16872 18345 16872 18345 4 gnd
rlabel metal3 s 13608 15422 13608 15422 4 gnd
rlabel metal3 s 15473 7273 15473 7273 4 gnd
rlabel metal3 s 13608 12025 13608 12025 4 gnd
rlabel metal3 s 19794 18216 19794 18216 4 gnd
rlabel metal3 s 13608 13605 13608 13605 4 gnd
rlabel metal3 s 22812 12693 22812 12693 4 gnd
rlabel metal3 s 13608 14869 13608 14869 4 gnd
rlabel metal3 s 13608 17002 13608 17002 4 gnd
rlabel metal3 s 1184 20432 1184 20432 4 gnd
rlabel metal3 s 9882 13111 9882 13111 4 gnd
rlabel metal3 s 13608 14079 13608 14079 4 gnd
rlabel metal3 s 25702 9132 25702 9132 4 gnd
rlabel metal3 s 16872 14869 16872 14869 4 gnd
rlabel metal3 s 20598 14273 20598 14273 4 gnd
rlabel metal3 s 16872 12262 16872 12262 4 gnd
rlabel metal3 s 20598 13483 20598 13483 4 gnd
rlabel metal3 s 15359 8066 15359 8066 4 gnd
rlabel metal3 s 8472 15056 8472 15056 4 gnd
rlabel metal3 s 13608 12815 13608 12815 4 gnd
rlabel metal3 s 29810 12652 29810 12652 4 gnd
rlabel metal3 s 15289 20844 15289 20844 4 gnd
rlabel metal3 s 25702 6304 25702 6304 4 gnd
rlabel metal3 s 9882 14691 9882 14691 4 gnd
rlabel metal3 s 20598 16643 20598 16643 4 gnd
rlabel metal3 s 20598 12693 20598 12693 4 gnd
rlabel metal3 s 10686 13081 10686 13081 4 gnd
rlabel metal3 s 14993 6504 14993 6504 4 gnd
rlabel metal3 s 13608 15185 13608 15185 4 gnd
rlabel metal3 s 15478 6302 15478 6302 4 gnd
rlabel metal3 s 9882 16271 9882 16271 4 gnd
rlabel metal3 s 19794 13081 19794 13081 4 gnd
rlabel metal3 s 13608 18029 13608 18029 4 gnd
rlabel metal3 s 20598 17851 20598 17851 4 gnd
rlabel metal3 s 10686 16241 10686 16241 4 gnd
rlabel metal3 s 20598 18223 20598 18223 4 gnd
rlabel metal3 s 16872 17555 16872 17555 4 gnd
rlabel metal3 s 7198 2573 7198 2573 4 gnd
rlabel metal3 s 19794 15846 19794 15846 4 gnd
rlabel metal3 s 16872 13842 16872 13842 4 gnd
rlabel metal3 s 7668 15853 7668 15853 4 gnd
rlabel metal3 s 29074 10412 29074 10412 4 gnd
rlabel metal3 s 10686 13476 10686 13476 4 gnd
rlabel metal3 s 9882 15063 9882 15063 4 gnd
rlabel metal3 s 9882 16643 9882 16643 4 gnd
rlabel metal3 s 448 20432 448 20432 4 gnd
rlabel metal3 s 25202 22360 25202 22360 4 gnd
rlabel metal3 s 4862 27368 4862 27368 4 gnd
rlabel metal3 s 0 2830 0 2830 4 gnd
rlabel metal3 s 448 18192 448 18192 4 gnd
rlabel metal3 s 10686 16636 10686 16636 4 gnd
rlabel metal3 s 8472 13476 8472 13476 4 gnd
rlabel metal3 s 13608 18345 13608 18345 4 gnd
rlabel metal3 s 14997 8066 14997 8066 4 gnd
rlabel metal3 s 13608 15975 13608 15975 4 gnd
rlabel metal3 s 29810 10412 29810 10412 4 gnd
rlabel metal3 s 0 -2 0 -2 4 gnd
rlabel metal3 s 13608 17239 13608 17239 4 gnd
rlabel metal3 s 19794 13871 19794 13871 4 gnd
rlabel metal3 s 16872 17792 16872 17792 4 gnd
rlabel metal3 s 16872 18582 16872 18582 4 gnd
rlabel metal3 s 6498 15056 6498 15056 4 gnd
rlabel metal3 s 9882 13483 9882 13483 4 gnd
rlabel metal3 s 10686 17426 10686 17426 4 gnd
rlabel metal3 s 29810 14892 29810 14892 4 gnd
rlabel metal3 s 16872 12025 16872 12025 4 gnd
rlabel metal3 s 13608 12499 13608 12499 4 gnd
rlabel metal3 s 29810 19372 29810 19372 4 gnd
rlabel metal3 s 16872 15975 16872 15975 4 gnd
rlabel metal3 s 15359 22778 15359 22778 4 gnd
rlabel metal3 s 1184 11472 1184 11472 4 gnd
rlabel metal3 s 22008 12686 22008 12686 4 gnd
rlabel metal3 s 20598 14691 20598 14691 4 gnd
rlabel metal3 s 1184 13712 1184 13712 4 gnd
rlabel metal3 s 19794 17426 19794 17426 4 gnd
rlabel metal3 s 5362 2828 5362 2828 4 gnd
rlabel metal3 s 16872 13605 16872 13605 4 gnd
rlabel metal3 s 5362 8484 5362 8484 4 gnd
rlabel metal3 s 10686 14266 10686 14266 4 gnd
rlabel metal3 s 10686 15451 10686 15451 4 gnd
rlabel metal3 s 22008 13476 22008 13476 4 gnd
rlabel metal3 s 13608 17555 13608 17555 4 gnd
rlabel metal3 s 7668 12693 7668 12693 4 gnd
rlabel metal3 s 13608 13052 13608 13052 4 gnd
rlabel metal3 s 10686 15056 10686 15056 4 gnd
rlabel metal3 s 25202 28016 25202 28016 4 gnd
rlabel metal3 s 16872 15185 16872 15185 4 gnd
rlabel metal3 s 13608 14395 13608 14395 4 gnd
rlabel metal3 s 20598 16271 20598 16271 4 gnd
rlabel metal3 s 15067 20844 15067 20844 4 gnd
rlabel metal2 s 26116 5740 26116 5740 4 addr1[2]
rlabel metal2 s 26116 6868 26116 6868 4 addr1[1]
rlabel metal2 s 4448 26804 4448 26804 4 addr0[3]
rlabel metal2 s 30088 27452 30088 27452 4 csb1
rlabel metal2 s 26116 4040 26116 4040 4 addr1[3]
rlabel metal2 s 28496 19111 28496 19111 4 rbl_bl1
rlabel metal2 s 26116 8568 26116 8568 4 addr1[0]
rlabel metal2 s 27241 27347 27241 27347 4 clk1
rlabel metal2 s 4448 23976 4448 23976 4 addr0[1]
rlabel metal2 s 170 2264 170 2264 4 web0
rlabel metal3 s 25702 4890 25702 4890 4 vdd
rlabel metal3 s 10958 12686 10958 12686 4 vdd
rlabel metal3 s 10958 17821 10958 17821 4 vdd
rlabel metal3 s 10958 18216 10958 18216 4 vdd
rlabel metal3 s 29810 16012 29810 16012 4 vdd
rlabel metal3 s 5362 4242 5362 4242 4 vdd
rlabel metal3 s 18651 15406 18651 15406 4 vdd
rlabel metal3 s 25202 20946 25202 20946 4 vdd
rlabel metal3 s 8366 3987 8366 3987 4 vdd
rlabel metal3 s 15552 19143 15552 19143 4 vdd
rlabel metal3 s 8744 15846 8744 15846 4 vdd
rlabel metal3 s 448 17072 448 17072 4 vdd
rlabel metal3 s 17736 15422 17736 15422 4 vdd
rlabel metal3 s 10958 13081 10958 13081 4 vdd
rlabel metal3 s 16057 19734 16057 19734 4 vdd
rlabel metal3 s 19522 17821 19522 17821 4 vdd
rlabel metal3 s 14809 11110 14809 11110 4 vdd
rlabel metal3 s 19522 14661 19522 14661 4 vdd
rlabel metal3 s 29074 18252 29074 18252 4 vdd
rlabel metal3 s 10958 15846 10958 15846 4 vdd
rlabel metal3 s 14997 22456 14997 22456 4 vdd
rlabel metal3 s 14985 21618 14985 21618 4 vdd
rlabel metal3 s 10307 17433 10307 17433 4 vdd
rlabel metal3 s 14304 19143 14304 19143 4 vdd
rlabel metal3 s 5362 7070 5362 7070 4 vdd
rlabel metal3 s 8744 12686 8744 12686 4 vdd
rlabel metal3 s 15359 8388 15359 8388 4 vdd
rlabel metal3 s 8093 12693 8093 12693 4 vdd
rlabel metal3 s 8093 15853 8093 15853 4 vdd
rlabel metal3 s 19522 14266 19522 14266 4 vdd
rlabel metal3 s 10307 16643 10307 16643 4 vdd
rlabel metal3 s 19522 16241 19522 16241 4 vdd
rlabel metal3 s 29074 11532 29074 11532 4 vdd
rlabel metal3 s 10958 17031 10958 17031 4 vdd
rlabel metal3 s 20173 13903 20173 13903 4 vdd
rlabel metal3 s 10958 17426 10958 17426 4 vdd
rlabel metal3 s 14985 9226 14985 9226 4 vdd
rlabel metal3 s 21736 15846 21736 15846 4 vdd
rlabel metal3 s 448 14832 448 14832 4 vdd
rlabel metal3 s 10958 15056 10958 15056 4 vdd
rlabel metal3 s 20173 16643 20173 16643 4 vdd
rlabel metal3 s 29810 13772 29810 13772 4 vdd
rlabel metal3 s 14423 11110 14423 11110 4 vdd
rlabel metal3 s 21736 15056 21736 15056 4 vdd
rlabel metal3 s 29810 11532 29810 11532 4 vdd
rlabel metal3 s 19522 16636 19522 16636 4 vdd
rlabel metal3 s 6770 12686 6770 12686 4 vdd
rlabel metal3 s 19522 18216 19522 18216 4 vdd
rlabel metal3 s 448 12592 448 12592 4 vdd
rlabel metal3 s 20173 13113 20173 13113 4 vdd
rlabel metal3 s 20173 14693 20173 14693 4 vdd
rlabel metal3 s 10958 13476 10958 13476 4 vdd
rlabel metal3 s 0 1414 0 1414 4 vdd
rlabel metal3 s 5362 1414 5362 1414 4 vdd
rlabel metal3 s 15484 6836 15484 6836 4 vdd
rlabel metal3 s 1184 14832 1184 14832 4 vdd
rlabel metal3 s 15464 5886 15464 5886 4 vdd
rlabel metal3 s 20173 17063 20173 17063 4 vdd
rlabel metal3 s 20173 15483 20173 15483 4 vdd
rlabel metal3 s 25702 7718 25702 7718 4 vdd
rlabel metal3 s 20173 16273 20173 16273 4 vdd
rlabel metal3 s 1184 21552 1184 21552 4 vdd
rlabel metal3 s 23710 12686 23710 12686 4 vdd
rlabel metal3 s 448 19312 448 19312 4 vdd
rlabel metal3 s 1184 12592 1184 12592 4 vdd
rlabel metal3 s 5362 9898 5362 9898 4 vdd
rlabel metal3 s 25202 26602 25202 26602 4 vdd
rlabel metal3 s 29074 9292 29074 9292 4 vdd
rlabel metal3 s 8093 15063 8093 15063 4 vdd
rlabel metal3 s 14928 19143 14928 19143 4 vdd
rlabel metal3 s 1184 17072 1184 17072 4 vdd
rlabel metal3 s 22387 15853 22387 15853 4 vdd
rlabel metal3 s 14928 11701 14928 11701 4 vdd
rlabel metal3 s 448 21552 448 21552 4 vdd
rlabel metal3 s 8744 15056 8744 15056 4 vdd
rlabel metal3 s 6770 15056 6770 15056 4 vdd
rlabel metal3 s 10307 15483 10307 15483 4 vdd
rlabel metal3 s 20173 17433 20173 17433 4 vdd
rlabel metal3 s 20173 15853 20173 15853 4 vdd
rlabel metal3 s 14892 5886 14892 5886 4 vdd
rlabel metal3 s 20173 14273 20173 14273 4 vdd
rlabel metal3 s 19522 15056 19522 15056 4 vdd
rlabel metal3 s 10958 16241 10958 16241 4 vdd
rlabel metal3 s 10307 14693 10307 14693 4 vdd
rlabel metal3 s 20173 12693 20173 12693 4 vdd
rlabel metal3 s 10958 16636 10958 16636 4 vdd
rlabel metal3 s 19522 13081 19522 13081 4 vdd
rlabel metal3 s 23710 15056 23710 15056 4 vdd
rlabel metal3 s 20173 17853 20173 17853 4 vdd
rlabel metal3 s 21736 12686 21736 12686 4 vdd
rlabel metal3 s 22387 13483 22387 13483 4 vdd
rlabel metal3 s 10307 18223 10307 18223 4 vdd
rlabel metal3 s 1184 19312 1184 19312 4 vdd
rlabel metal3 s 19522 15451 19522 15451 4 vdd
rlabel metal3 s 10307 13483 10307 13483 4 vdd
rlabel metal3 s 29074 13772 29074 13772 4 vdd
rlabel metal3 s 21736 13476 21736 13476 4 vdd
rlabel metal3 s 19522 13476 19522 13476 4 vdd
rlabel metal3 s 10307 14273 10307 14273 4 vdd
rlabel metal3 s 11829 15406 11829 15406 4 vdd
rlabel metal3 s 22387 12693 22387 12693 4 vdd
rlabel metal3 s 10958 13871 10958 13871 4 vdd
rlabel metal3 s 20173 18223 20173 18223 4 vdd
rlabel metal3 s 10307 15853 10307 15853 4 vdd
rlabel metal3 s 19522 13871 19522 13871 4 vdd
rlabel metal3 s 29810 9292 29810 9292 4 vdd
rlabel metal3 s 12744 15422 12744 15422 4 vdd
rlabel metal3 s 10958 14661 10958 14661 4 vdd
rlabel metal3 s 8093 13483 8093 13483 4 vdd
rlabel metal3 s 10958 15451 10958 15451 4 vdd
rlabel metal3 s 19522 15846 19522 15846 4 vdd
rlabel metal3 s 22387 15063 22387 15063 4 vdd
rlabel metal3 s 29810 18252 29810 18252 4 vdd
rlabel metal3 s 4862 23126 4862 23126 4 vdd
rlabel metal3 s 10307 13903 10307 13903 4 vdd
rlabel metal3 s 10307 12693 10307 12693 4 vdd
rlabel metal3 s 19522 17426 19522 17426 4 vdd
rlabel metal3 s 10307 16273 10307 16273 4 vdd
rlabel metal3 s 15671 11110 15671 11110 4 vdd
rlabel metal3 s 10307 15063 10307 15063 4 vdd
rlabel metal3 s 20173 15063 20173 15063 4 vdd
rlabel metal3 s 15552 11701 15552 11701 4 vdd
rlabel metal3 s 10307 17853 10307 17853 4 vdd
rlabel metal3 s 14997 8388 14997 8388 4 vdd
rlabel metal3 s 14304 11701 14304 11701 4 vdd
rlabel metal3 s 14809 19734 14809 19734 4 vdd
rlabel metal3 s 10958 14266 10958 14266 4 vdd
rlabel metal3 s 7198 3987 7198 3987 4 vdd
rlabel metal3 s 14872 6836 14872 6836 4 vdd
rlabel metal3 s 16176 19143 16176 19143 4 vdd
rlabel metal3 s 4862 25954 4862 25954 4 vdd
rlabel metal3 s 15671 19734 15671 19734 4 vdd
rlabel metal3 s 8744 13476 8744 13476 4 vdd
rlabel metal3 s 19522 12686 19522 12686 4 vdd
rlabel metal3 s 10307 13113 10307 13113 4 vdd
rlabel metal3 s 30258 26602 30258 26602 4 vdd
rlabel metal3 s 16176 11701 16176 11701 4 vdd
rlabel metal3 s 15359 22456 15359 22456 4 vdd
rlabel metal3 s 15371 9226 15371 9226 4 vdd
rlabel metal3 s 19522 17031 19522 17031 4 vdd
rlabel metal3 s 10307 17063 10307 17063 4 vdd
rlabel metal3 s 15371 21618 15371 21618 4 vdd
rlabel metal3 s 29074 16012 29074 16012 4 vdd
rlabel metal3 s 25202 23774 25202 23774 4 vdd
rlabel metal3 s 20173 13483 20173 13483 4 vdd
rlabel metal1 s 15613 22759 15613 22759 4 dout1[1]
<< properties >>
string FIXED_BBOX 0 0 30258 28016
<< end >>
