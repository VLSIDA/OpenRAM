magic
tech gf180mcuD
magscale 1 10
timestamp 1694492161
<< nwell >>
rect 625 -40 1305 640
<< nmos >>
rect 161 300 331 360
rect 161 190 331 250
<< pmos >>
rect 715 330 1056 390
rect 715 160 1056 220
<< ndiff >>
rect 161 438 331 460
rect 161 392 223 438
rect 269 392 331 438
rect 161 360 331 392
rect 161 250 331 300
rect 161 158 331 190
rect 161 112 223 158
rect 269 112 331 158
rect 161 90 331 112
<< pdiff >>
rect 715 468 1056 490
rect 715 422 768 468
rect 1002 422 1056 468
rect 715 390 1056 422
rect 715 298 1056 330
rect 715 252 768 298
rect 1002 252 1056 298
rect 715 220 1056 252
rect 715 128 1056 160
rect 715 82 768 128
rect 1002 82 1056 128
rect 715 60 1056 82
<< ndiffc >>
rect 223 392 269 438
rect 223 112 269 158
<< pdiffc >>
rect 768 422 1002 468
rect 768 252 1002 298
rect 768 82 1002 128
<< psubdiff >>
rect 24 23 131 40
rect 24 -23 64 23
rect 110 -23 131 23
rect 24 -40 131 -23
<< nsubdiff >>
rect 1122 107 1202 144
rect 1122 61 1139 107
rect 1185 61 1202 107
rect 1122 37 1202 61
<< psubdiffcont >>
rect 64 -23 110 23
<< nsubdiffcont >>
rect 1139 61 1185 107
<< polysilicon >>
rect 38 373 121 400
rect 38 327 54 373
rect 100 360 121 373
rect 381 360 715 390
rect 100 327 161 360
rect 38 300 161 327
rect 331 330 715 360
rect 1056 330 1106 390
rect 331 300 421 330
rect 38 234 161 250
rect 38 188 54 234
rect 100 190 161 234
rect 331 220 421 250
rect 331 190 715 220
rect 100 188 121 190
rect 38 150 121 188
rect 381 160 715 190
rect 1056 160 1106 220
<< polycontact >>
rect 54 327 100 373
rect 54 188 100 234
<< metal1 >>
rect 161 438 401 440
rect 51 373 103 425
rect 161 392 223 438
rect 269 392 401 438
rect 757 422 768 468
rect 1002 422 1014 468
rect 853 416 865 422
rect 917 416 929 422
rect 161 390 401 392
rect 51 327 54 373
rect 100 327 103 373
rect 51 313 103 327
rect 351 300 401 390
rect 1080 300 1132 463
rect 351 298 1132 300
rect 351 252 768 298
rect 1002 252 1132 298
rect 351 250 1132 252
rect 51 234 103 248
rect 51 188 54 234
rect 100 188 103 234
rect 51 129 103 188
rect 191 106 223 158
rect 275 106 298 158
rect 853 128 865 134
rect 917 128 929 134
rect 191 100 298 106
rect 757 82 768 128
rect 1002 82 1014 128
rect 1089 58 1136 110
rect 1188 58 1200 110
rect 30 26 129 36
rect 30 -26 61 26
rect 113 -26 129 26
rect 30 -34 129 -26
<< via1 >>
rect 865 422 917 468
rect 865 416 917 422
rect 223 112 269 158
rect 269 112 275 158
rect 223 106 275 112
rect 865 128 917 134
rect 865 82 917 128
rect 1136 107 1188 110
rect 1136 61 1139 107
rect 1139 61 1185 107
rect 1185 61 1188 107
rect 1136 58 1188 61
rect 61 23 113 26
rect 61 -23 64 23
rect 64 -23 110 23
rect 110 -23 113 23
rect 61 -26 113 -23
<< metal2 >>
rect 221 158 277 520
rect 221 106 223 158
rect 275 106 277 158
rect 221 28 277 106
rect 39 26 277 28
rect 39 -26 61 26
rect 113 -26 277 26
rect 863 468 919 520
rect 863 416 865 468
rect 917 416 919 468
rect 863 134 919 416
rect 863 82 865 134
rect 917 112 919 134
rect 917 110 1200 112
rect 917 82 1136 110
rect 863 58 1136 82
rect 1188 58 1200 110
rect 863 56 1200 58
rect 863 8 919 56
rect 39 -28 277 -26
<< labels >>
rlabel metal1 s 1106 439 1106 439 4 Y
rlabel metal1 s 77 211 77 211 4 B
rlabel metal1 s 77 350 77 350 4 A
rlabel metal2 s 891 33 891 33 4 VDD
rlabel metal2 s 250 56 250 56 4 GND
<< properties >>
string FIXED_BBOX 0 0 1305 522
<< end >>
