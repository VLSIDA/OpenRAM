magic
tech sky130A
magscale 1 2
timestamp 1595931502
<< checkpaint >>
rect -1260 -1260 20596 18535
<< locali >>
rect 11498 12757 11641 12777
rect 7466 12723 7645 12757
rect 11498 12743 11786 12757
rect 11607 12723 11786 12743
rect 7611 12557 7645 12723
rect 7611 12523 7754 12557
rect 7611 12427 7754 12461
rect 7611 12261 7645 12427
rect 7466 12227 7645 12261
rect 11607 12241 11786 12261
rect 11498 12227 11786 12241
rect 11498 12207 11641 12227
rect 11498 11967 11641 11987
rect 7466 11933 7645 11967
rect 11498 11953 11786 11967
rect 11607 11933 11786 11953
rect 7611 11767 7645 11933
rect 7611 11733 7754 11767
rect 7611 11637 7754 11671
rect 7611 11471 7645 11637
rect 7466 11437 7645 11471
rect 11607 11451 11786 11471
rect 11498 11437 11786 11451
rect 11498 11417 11641 11437
rect 11498 11177 11641 11197
rect 7466 11143 7645 11177
rect 11498 11163 11786 11177
rect 11607 11143 11786 11163
rect 7611 10977 7645 11143
rect 7611 10943 7754 10977
rect 7611 10847 7754 10881
rect 7611 10681 7645 10847
rect 7466 10647 7645 10681
rect 11607 10661 11786 10681
rect 11498 10647 11786 10661
rect 11498 10627 11641 10647
rect 11498 10387 11641 10407
rect 7466 10353 7645 10387
rect 11498 10373 11786 10387
rect 11607 10353 11786 10373
rect 7611 10187 7645 10353
rect 7611 10153 7754 10187
rect 7611 10057 7754 10091
rect 7611 9891 7645 10057
rect 7466 9857 7645 9891
rect 11607 9871 11786 9891
rect 11498 9857 11786 9871
rect 11498 9837 11641 9857
rect 11498 9597 11641 9617
rect 7466 9563 7645 9597
rect 11498 9583 11786 9597
rect 11607 9563 11786 9583
rect 7611 9397 7645 9563
rect 7611 9363 7754 9397
rect 7611 9267 7754 9301
rect 7611 9101 7645 9267
rect 7466 9067 7645 9101
rect 11607 9081 11786 9101
rect 11498 9067 11786 9081
rect 11498 9047 11641 9067
rect 11498 8807 11641 8827
rect 7466 8773 7645 8807
rect 11498 8793 11786 8807
rect 11607 8773 11786 8793
rect 7611 8607 7645 8773
rect 7611 8573 7754 8607
rect 7611 8477 7754 8511
rect 7611 8311 7645 8477
rect 7466 8277 7645 8311
rect 11607 8291 11786 8311
rect 11498 8277 11786 8291
rect 11498 8257 11641 8277
rect 11498 8017 11641 8037
rect 7466 7983 7645 8017
rect 11498 8003 11786 8017
rect 11607 7983 11786 8003
rect 7611 7817 7645 7983
rect 7611 7783 7754 7817
rect 7611 7687 7754 7721
rect 7611 7521 7645 7687
rect 7466 7487 7645 7521
rect 11607 7501 11786 7521
rect 11498 7487 11786 7501
rect 11498 7467 11641 7487
rect 11498 7227 11641 7247
rect 7466 7193 7645 7227
rect 11498 7213 11786 7227
rect 11607 7193 11786 7213
rect 7611 7027 7645 7193
rect 7611 6993 7754 7027
rect 7611 6897 7754 6931
rect 7611 6731 7645 6897
rect 7466 6697 7645 6731
rect 11607 6711 11786 6731
rect 11498 6697 11786 6711
rect 11498 6677 11641 6697
<< metal1 >>
rect 9106 16937 9152 17191
rect 9976 16937 10022 17191
rect 10316 14683 10344 14807
rect 9068 13817 9096 13929
rect 9532 13817 9560 13929
rect 9068 13789 9328 13817
rect 9300 13677 9328 13789
rect 9372 13789 9560 13817
rect 9692 13817 9720 13929
rect 10156 13817 10184 13929
rect 9692 13789 9880 13817
rect 9372 13677 9400 13789
rect 9852 13677 9880 13789
rect 9924 13789 10184 13817
rect 10316 13817 10344 13929
rect 10780 13817 10808 13929
rect 10316 13789 10576 13817
rect 9924 13677 9952 13789
rect 10548 13677 10576 13789
rect 10620 13789 10808 13817
rect 10620 13677 10648 13789
rect 11636 13377 13648 13405
rect 11466 12734 11530 12786
rect 7722 12514 7786 12566
rect 7722 12418 7786 12470
rect 11466 12198 11530 12250
rect 11466 11944 11530 11996
rect 7722 11724 7786 11776
rect 7722 11628 7786 11680
rect 11466 11408 11530 11460
rect 11466 11154 11530 11206
rect 7722 10934 7786 10986
rect 7722 10838 7786 10890
rect 11466 10618 11530 10670
rect 18 6596 46 10546
rect 98 6596 126 10546
rect 178 6596 206 10546
rect 258 6596 286 10546
rect 11466 10364 11530 10416
rect 7722 10144 7786 10196
rect 7722 10048 7786 10100
rect 11466 9828 11530 9880
rect 11466 9574 11530 9626
rect 7722 9354 7786 9406
rect 7722 9258 7786 9310
rect 11466 9038 11530 9090
rect 11466 8784 11530 8836
rect 7722 8564 7786 8616
rect 7722 8468 7786 8520
rect 11466 8248 11530 8300
rect 11466 7994 11530 8046
rect 7722 7774 7786 7826
rect 7722 7678 7786 7730
rect 11466 7458 11530 7510
rect 11466 7204 11530 7256
rect 7722 6984 7786 7036
rect 7722 6888 7786 6940
rect 11466 6668 11530 6720
rect 18966 6596 18994 10546
rect 19046 6596 19074 10546
rect 19126 6596 19154 10546
rect 19206 6596 19234 10546
rect 5604 6049 7520 6077
rect 8820 5665 8848 5777
rect 8444 5637 8848 5665
rect 8892 5665 8920 5777
rect 9084 5665 9112 5777
rect 8892 5637 8936 5665
rect 8444 5525 8472 5637
rect 8908 5525 8936 5637
rect 9068 5637 9112 5665
rect 9156 5665 9184 5777
rect 10068 5665 10096 5777
rect 9156 5637 9560 5665
rect 9068 5525 9096 5637
rect 9532 5525 9560 5637
rect 9692 5637 10096 5665
rect 10140 5665 10168 5777
rect 10140 5637 10184 5665
rect 9692 5525 9720 5637
rect 10156 5525 10184 5637
rect 8908 4647 8936 4771
rect 9106 2263 9152 2517
rect 9976 2263 10022 2517
rect 7272 94 9626 122
rect 9257 4 9317 60
rect 9811 4 9871 60
<< metal2 >>
rect 10302 14783 10358 14831
rect 11622 13028 11650 17275
rect 11746 13047 11774 17275
rect 11870 13047 11898 17275
rect 9626 13000 11650 13028
rect 13634 12887 13662 13391
rect 5590 6063 5618 6567
rect 7134 0 7162 6407
rect 7258 0 7286 6407
rect 7382 0 7410 6407
rect 7506 6234 7534 6407
rect 7506 6206 9626 6234
rect 7506 0 7534 6206
rect 8894 4623 8950 4671
<< metal3 >>
rect 9334 17034 9432 17132
rect 9696 17034 9794 17132
rect 9334 16712 9432 16810
rect 9696 16712 9794 16810
rect 9322 15874 9420 15972
rect 9708 15874 9806 15972
rect 9404 15100 9502 15198
rect 9626 15100 9724 15198
rect 9626 14967 11884 15027
rect 10330 14777 19336 14837
rect 9938 14628 11760 14688
rect 9146 13990 9244 14088
rect 10008 13990 10106 14088
rect 10394 13990 10492 14088
rect 8641 13399 8739 13497
rect 9284 13418 9344 13478
rect 9908 13418 9968 13478
rect 10513 13399 10611 13497
rect 7964 13094 8024 13154
rect 11228 13094 11288 13154
rect 7964 12857 8024 12917
rect 11228 12857 11288 12917
rect 7964 12620 8024 12680
rect 11228 12620 11288 12680
rect 4219 12479 4317 12577
rect 4644 12479 4742 12577
rect 5023 12472 5121 12570
rect 5295 12472 5393 12570
rect 13859 12472 13957 12570
rect 14131 12472 14229 12570
rect 14510 12479 14608 12577
rect 14935 12479 15033 12577
rect 7964 12304 8024 12364
rect 11228 12304 11288 12364
rect 4219 12107 4317 12205
rect 4644 12109 4742 12207
rect 5023 12077 5121 12175
rect 5295 12077 5393 12175
rect 7964 12067 8024 12127
rect 11228 12067 11288 12127
rect 13859 12077 13957 12175
rect 14131 12077 14229 12175
rect 14510 12109 14608 12207
rect 14935 12107 15033 12205
rect 7964 11830 8024 11890
rect 11228 11830 11288 11890
rect 4219 11689 4317 11787
rect 4644 11689 4742 11787
rect 5023 11682 5121 11780
rect 5295 11682 5393 11780
rect 13859 11682 13957 11780
rect 14131 11682 14229 11780
rect 14510 11689 14608 11787
rect 14935 11689 15033 11787
rect 7964 11514 8024 11574
rect 11228 11514 11288 11574
rect 4219 11317 4317 11415
rect 4644 11319 4742 11417
rect 5023 11287 5121 11385
rect 5295 11287 5393 11385
rect 7964 11277 8024 11337
rect 11228 11277 11288 11337
rect 13859 11287 13957 11385
rect 14131 11287 14229 11385
rect 14510 11319 14608 11417
rect 14935 11317 15033 11415
rect 7964 11040 8024 11100
rect 11228 11040 11288 11100
rect 4219 10899 4317 10997
rect 4644 10899 4742 10997
rect 5023 10892 5121 10990
rect 5295 10892 5393 10990
rect 13859 10892 13957 10990
rect 14131 10892 14229 10990
rect 14510 10899 14608 10997
rect 14935 10899 15033 10997
rect 7964 10724 8024 10784
rect 11228 10724 11288 10784
rect 4219 10527 4317 10625
rect 4644 10529 4742 10627
rect 5023 10497 5121 10595
rect 5295 10497 5393 10595
rect 7964 10487 8024 10547
rect 11228 10487 11288 10547
rect 13859 10497 13957 10595
rect 14131 10497 14229 10595
rect 14510 10529 14608 10627
rect 14935 10527 15033 10625
rect 7964 10250 8024 10310
rect 11228 10250 11288 10310
rect 2005 10109 2103 10207
rect 2430 10109 2528 10207
rect 2809 10102 2907 10200
rect 3081 10102 3179 10200
rect 4219 10109 4317 10207
rect 4644 10109 4742 10207
rect 5023 10102 5121 10200
rect 5295 10102 5393 10200
rect 13859 10102 13957 10200
rect 14131 10102 14229 10200
rect 14510 10109 14608 10207
rect 14935 10109 15033 10207
rect 16073 10102 16171 10200
rect 16345 10102 16443 10200
rect 16724 10109 16822 10207
rect 17149 10109 17247 10207
rect 7964 9934 8024 9994
rect 11228 9934 11288 9994
rect 4219 9737 4317 9835
rect 4644 9739 4742 9837
rect 5023 9707 5121 9805
rect 5295 9707 5393 9805
rect 5741 9663 5839 9761
rect 6166 9662 6264 9760
rect 6583 9678 6681 9776
rect 7081 9678 7179 9776
rect 7964 9697 8024 9757
rect 11228 9697 11288 9757
rect 12073 9678 12171 9776
rect 12571 9678 12669 9776
rect 12988 9662 13086 9760
rect 13413 9663 13511 9761
rect 13859 9707 13957 9805
rect 14131 9707 14229 9805
rect 14510 9739 14608 9837
rect 14935 9737 15033 9835
rect 7964 9460 8024 9520
rect 11228 9460 11288 9520
rect 835 9312 933 9410
rect 1107 9312 1205 9410
rect 2005 9319 2103 9417
rect 2430 9319 2528 9417
rect 2809 9312 2907 9410
rect 3081 9312 3179 9410
rect 4219 9319 4317 9417
rect 4644 9319 4742 9417
rect 5023 9312 5121 9410
rect 5295 9312 5393 9410
rect 13859 9312 13957 9410
rect 14131 9312 14229 9410
rect 14510 9319 14608 9417
rect 14935 9319 15033 9417
rect 16073 9312 16171 9410
rect 16345 9312 16443 9410
rect 16724 9319 16822 9417
rect 17149 9319 17247 9417
rect 18047 9312 18145 9410
rect 18319 9312 18417 9410
rect 7964 9144 8024 9204
rect 11228 9144 11288 9204
rect 4219 8947 4317 9045
rect 4644 8949 4742 9047
rect 5023 8917 5121 9015
rect 5295 8917 5393 9015
rect 7964 8907 8024 8967
rect 11228 8907 11288 8967
rect 13859 8917 13957 9015
rect 14131 8917 14229 9015
rect 14510 8949 14608 9047
rect 14935 8947 15033 9045
rect 7964 8670 8024 8730
rect 11228 8670 11288 8730
rect 4219 8529 4317 8627
rect 4644 8529 4742 8627
rect 5023 8522 5121 8620
rect 5295 8522 5393 8620
rect 13859 8522 13957 8620
rect 14131 8522 14229 8620
rect 14510 8529 14608 8627
rect 14935 8529 15033 8627
rect 7964 8354 8024 8414
rect 11228 8354 11288 8414
rect 4219 8157 4317 8255
rect 4644 8159 4742 8257
rect 5023 8127 5121 8225
rect 5295 8127 5393 8225
rect 7964 8117 8024 8177
rect 11228 8117 11288 8177
rect 13859 8127 13957 8225
rect 14131 8127 14229 8225
rect 14510 8159 14608 8257
rect 14935 8157 15033 8255
rect 7964 7880 8024 7940
rect 11228 7880 11288 7940
rect 2005 7739 2103 7837
rect 2430 7739 2528 7837
rect 2809 7732 2907 7830
rect 3081 7732 3179 7830
rect 4219 7739 4317 7837
rect 4644 7739 4742 7837
rect 5023 7732 5121 7830
rect 5295 7732 5393 7830
rect 13859 7732 13957 7830
rect 14131 7732 14229 7830
rect 14510 7739 14608 7837
rect 14935 7739 15033 7837
rect 16073 7732 16171 7830
rect 16345 7732 16443 7830
rect 16724 7739 16822 7837
rect 17149 7739 17247 7837
rect 7964 7564 8024 7624
rect 11228 7564 11288 7624
rect 4219 7367 4317 7465
rect 4644 7369 4742 7467
rect 5023 7337 5121 7435
rect 5295 7337 5393 7435
rect 7964 7327 8024 7387
rect 11228 7327 11288 7387
rect 13859 7337 13957 7435
rect 14131 7337 14229 7435
rect 14510 7369 14608 7467
rect 14935 7367 15033 7465
rect 7964 7090 8024 7150
rect 11228 7090 11288 7150
rect 835 6942 933 7040
rect 1107 6942 1205 7040
rect 2005 6949 2103 7047
rect 2430 6949 2528 7047
rect 2809 6942 2907 7040
rect 3081 6942 3179 7040
rect 4219 6949 4317 7047
rect 4644 6949 4742 7047
rect 5023 6942 5121 7040
rect 5295 6942 5393 7040
rect 13859 6942 13957 7040
rect 14131 6942 14229 7040
rect 14510 6949 14608 7047
rect 14935 6949 15033 7047
rect 16073 6942 16171 7040
rect 16345 6942 16443 7040
rect 16724 6949 16822 7047
rect 17149 6949 17247 7047
rect 18047 6942 18145 7040
rect 18319 6942 18417 7040
rect 7964 6774 8024 6834
rect 11228 6774 11288 6834
rect 7964 6537 8024 6597
rect 11228 6537 11288 6597
rect 7964 6300 8024 6360
rect 11228 6300 11288 6360
rect 8641 5957 8739 6055
rect 9284 5976 9344 6036
rect 9908 5976 9968 6036
rect 10513 5957 10611 6055
rect 8760 5366 8858 5464
rect 9146 5366 9244 5464
rect 10008 5366 10106 5464
rect 7396 4766 9314 4826
rect 0 4617 8922 4677
rect 7148 4427 9626 4487
rect 9404 4256 9502 4354
rect 9626 4256 9724 4354
rect 9322 3482 9420 3580
rect 9708 3482 9806 3580
rect 9334 2644 9432 2742
rect 9696 2644 9794 2742
rect 9334 2322 9432 2420
rect 9696 2322 9794 2420
rect 9220 1529 9318 1627
rect 9810 1529 9908 1627
rect 9209 1092 9307 1190
rect 9821 1092 9919 1190
rect 9330 760 9428 858
rect 9700 760 9798 858
rect 9215 558 9313 656
rect 9815 558 9913 656
rect 9229 142 9327 240
rect 9801 142 9899 240
use port_address  port_address_1
timestamp 1595931502
transform 1 0 0 0 1 6567
box 0 -56 7484 6405
use port_address  port_address_0
timestamp 1595931502
transform -1 0 19252 0 1 6567
box 0 -56 7484 6405
use contact_9  contact_9_5
timestamp 1595931502
transform 1 0 8889 0 1 4610
box 0 0 66 74
use contact_9  contact_9_4
timestamp 1595931502
transform 1 0 7363 0 1 4759
box 0 0 66 74
use contact_9  contact_9_3
timestamp 1595931502
transform 1 0 7115 0 1 4420
box 0 0 66 74
use contact_9  contact_9_2
timestamp 1595931502
transform 1 0 10297 0 1 14770
box 0 0 66 74
use contact_9  contact_9_1
timestamp 1595931502
transform 1 0 11727 0 1 14621
box 0 0 66 74
use contact_9  contact_9_0
timestamp 1595931502
transform 1 0 11851 0 1 14960
box 0 0 66 74
use replica_bitcell_array  replica_bitcell_array_0
timestamp 1595931502
transform 1 0 7754 0 1 5777
box -42 0 3786 7900
use port_data_0  port_data_0_0
timestamp 1595931502
transform 1 0 9002 0 1 13677
box -160 238 1872 3514
use port_data  port_data_0
timestamp 1595931502
transform 1 0 8378 0 -1 5777
box 0 238 1908 5773
use contact_8  contact_8_6
timestamp 1595931502
transform 1 0 8890 0 1 4615
box 0 0 64 64
use contact_8  contact_8_5
timestamp 1595931502
transform 1 0 7240 0 1 76
box 0 0 64 64
use contact_8  contact_8_4
timestamp 1595931502
transform 1 0 5572 0 1 6031
box 0 0 64 64
use contact_8  contact_8_3
timestamp 1595931502
transform 1 0 7488 0 1 6031
box 0 0 64 64
use contact_8  contact_8_2
timestamp 1595931502
transform 1 0 10298 0 1 14775
box 0 0 64 64
use contact_8  contact_8_1
timestamp 1595931502
transform 1 0 13616 0 1 13359
box 0 0 64 64
use contact_8  contact_8_0
timestamp 1595931502
transform 1 0 11604 0 1 13359
box 0 0 64 64
use contact_22  contact_22_31
timestamp 1595931502
transform 1 0 7722 0 1 6888
box 0 0 64 52
use contact_22  contact_22_30
timestamp 1595931502
transform 1 0 7722 0 1 6984
box 0 0 64 52
use contact_22  contact_22_29
timestamp 1595931502
transform 1 0 7722 0 1 7678
box 0 0 64 52
use contact_22  contact_22_28
timestamp 1595931502
transform 1 0 7722 0 1 7774
box 0 0 64 52
use contact_22  contact_22_27
timestamp 1595931502
transform 1 0 7722 0 1 8468
box 0 0 64 52
use contact_22  contact_22_26
timestamp 1595931502
transform 1 0 7722 0 1 8564
box 0 0 64 52
use contact_22  contact_22_25
timestamp 1595931502
transform 1 0 7722 0 1 9258
box 0 0 64 52
use contact_22  contact_22_24
timestamp 1595931502
transform 1 0 7722 0 1 9354
box 0 0 64 52
use contact_22  contact_22_23
timestamp 1595931502
transform 1 0 7722 0 1 10048
box 0 0 64 52
use contact_22  contact_22_22
timestamp 1595931502
transform 1 0 7722 0 1 10144
box 0 0 64 52
use contact_22  contact_22_21
timestamp 1595931502
transform 1 0 7722 0 1 10838
box 0 0 64 52
use contact_22  contact_22_20
timestamp 1595931502
transform 1 0 7722 0 1 10934
box 0 0 64 52
use contact_22  contact_22_19
timestamp 1595931502
transform 1 0 7722 0 1 11628
box 0 0 64 52
use contact_22  contact_22_18
timestamp 1595931502
transform 1 0 7722 0 1 11724
box 0 0 64 52
use contact_22  contact_22_17
timestamp 1595931502
transform 1 0 7722 0 1 12418
box 0 0 64 52
use contact_22  contact_22_16
timestamp 1595931502
transform 1 0 7722 0 1 12514
box 0 0 64 52
use contact_22  contact_22_15
timestamp 1595931502
transform 1 0 11466 0 1 6668
box 0 0 64 52
use contact_22  contact_22_14
timestamp 1595931502
transform 1 0 11466 0 1 7204
box 0 0 64 52
use contact_22  contact_22_13
timestamp 1595931502
transform 1 0 11466 0 1 7458
box 0 0 64 52
use contact_22  contact_22_12
timestamp 1595931502
transform 1 0 11466 0 1 7994
box 0 0 64 52
use contact_22  contact_22_11
timestamp 1595931502
transform 1 0 11466 0 1 8248
box 0 0 64 52
use contact_22  contact_22_10
timestamp 1595931502
transform 1 0 11466 0 1 8784
box 0 0 64 52
use contact_22  contact_22_9
timestamp 1595931502
transform 1 0 11466 0 1 9038
box 0 0 64 52
use contact_22  contact_22_8
timestamp 1595931502
transform 1 0 11466 0 1 9574
box 0 0 64 52
use contact_22  contact_22_7
timestamp 1595931502
transform 1 0 11466 0 1 9828
box 0 0 64 52
use contact_22  contact_22_6
timestamp 1595931502
transform 1 0 11466 0 1 10364
box 0 0 64 52
use contact_22  contact_22_5
timestamp 1595931502
transform 1 0 11466 0 1 10618
box 0 0 64 52
use contact_22  contact_22_4
timestamp 1595931502
transform 1 0 11466 0 1 11154
box 0 0 64 52
use contact_22  contact_22_3
timestamp 1595931502
transform 1 0 11466 0 1 11408
box 0 0 64 52
use contact_22  contact_22_2
timestamp 1595931502
transform 1 0 11466 0 1 11944
box 0 0 64 52
use contact_22  contact_22_1
timestamp 1595931502
transform 1 0 11466 0 1 12198
box 0 0 64 52
use contact_22  contact_22_0
timestamp 1595931502
transform 1 0 11466 0 1 12734
box 0 0 64 52
use contact_21  contact_21_31
timestamp 1595931502
transform 1 0 7721 0 1 6891
box 0 0 66 46
use contact_21  contact_21_30
timestamp 1595931502
transform 1 0 7721 0 1 6987
box 0 0 66 46
use contact_21  contact_21_29
timestamp 1595931502
transform 1 0 7721 0 1 7681
box 0 0 66 46
use contact_21  contact_21_28
timestamp 1595931502
transform 1 0 7721 0 1 7777
box 0 0 66 46
use contact_21  contact_21_27
timestamp 1595931502
transform 1 0 7721 0 1 8471
box 0 0 66 46
use contact_21  contact_21_26
timestamp 1595931502
transform 1 0 7721 0 1 8567
box 0 0 66 46
use contact_21  contact_21_25
timestamp 1595931502
transform 1 0 7721 0 1 9261
box 0 0 66 46
use contact_21  contact_21_24
timestamp 1595931502
transform 1 0 7721 0 1 9357
box 0 0 66 46
use contact_21  contact_21_23
timestamp 1595931502
transform 1 0 7721 0 1 10051
box 0 0 66 46
use contact_21  contact_21_22
timestamp 1595931502
transform 1 0 7721 0 1 10147
box 0 0 66 46
use contact_21  contact_21_21
timestamp 1595931502
transform 1 0 7721 0 1 10841
box 0 0 66 46
use contact_21  contact_21_20
timestamp 1595931502
transform 1 0 7721 0 1 10937
box 0 0 66 46
use contact_21  contact_21_19
timestamp 1595931502
transform 1 0 7721 0 1 11631
box 0 0 66 46
use contact_21  contact_21_18
timestamp 1595931502
transform 1 0 7721 0 1 11727
box 0 0 66 46
use contact_21  contact_21_17
timestamp 1595931502
transform 1 0 7721 0 1 12421
box 0 0 66 46
use contact_21  contact_21_16
timestamp 1595931502
transform 1 0 7721 0 1 12517
box 0 0 66 46
use contact_21  contact_21_15
timestamp 1595931502
transform 1 0 11465 0 1 6671
box 0 0 66 46
use contact_21  contact_21_14
timestamp 1595931502
transform 1 0 11465 0 1 7207
box 0 0 66 46
use contact_21  contact_21_13
timestamp 1595931502
transform 1 0 11465 0 1 7461
box 0 0 66 46
use contact_21  contact_21_12
timestamp 1595931502
transform 1 0 11465 0 1 7997
box 0 0 66 46
use contact_21  contact_21_11
timestamp 1595931502
transform 1 0 11465 0 1 8251
box 0 0 66 46
use contact_21  contact_21_10
timestamp 1595931502
transform 1 0 11465 0 1 8787
box 0 0 66 46
use contact_21  contact_21_9
timestamp 1595931502
transform 1 0 11465 0 1 9041
box 0 0 66 46
use contact_21  contact_21_8
timestamp 1595931502
transform 1 0 11465 0 1 9577
box 0 0 66 46
use contact_21  contact_21_7
timestamp 1595931502
transform 1 0 11465 0 1 9831
box 0 0 66 46
use contact_21  contact_21_6
timestamp 1595931502
transform 1 0 11465 0 1 10367
box 0 0 66 46
use contact_21  contact_21_5
timestamp 1595931502
transform 1 0 11465 0 1 10621
box 0 0 66 46
use contact_21  contact_21_4
timestamp 1595931502
transform 1 0 11465 0 1 11157
box 0 0 66 46
use contact_21  contact_21_3
timestamp 1595931502
transform 1 0 11465 0 1 11411
box 0 0 66 46
use contact_21  contact_21_2
timestamp 1595931502
transform 1 0 11465 0 1 11947
box 0 0 66 46
use contact_21  contact_21_1
timestamp 1595931502
transform 1 0 11465 0 1 12201
box 0 0 66 46
use contact_21  contact_21_0
timestamp 1595931502
transform 1 0 11465 0 1 12737
box 0 0 66 46
<< labels >>
rlabel metal1 s 9999 17064 9999 17064 4 dout1_1
rlabel metal1 s 19220 8571 19220 8571 4 addr1_0
rlabel metal2 s 11884 15161 11884 15161 4 s_en1
rlabel metal1 s 272 8571 272 8571 4 addr0_3
rlabel metal2 s 11760 15161 11760 15161 4 p_en_bar1
rlabel metal1 s 18980 8571 18980 8571 4 addr1_3
rlabel metal1 s 9129 17064 9129 17064 4 dout1_0
rlabel metal1 s 9999 2390 9999 2390 4 dout0_1
rlabel metal1 s 192 8571 192 8571 4 addr0_2
rlabel metal3 s 4461 4647 4461 4647 4 rbl_bl0
rlabel metal1 s 9841 32 9841 32 4 din0_1
rlabel metal3 s 7994 12097 7994 12097 4 gnd
rlabel metal3 s 9383 17083 9383 17083 4 gnd
rlabel metal3 s 9745 2371 9745 2371 4 gnd
rlabel metal3 s 11258 7120 11258 7120 4 gnd
rlabel metal3 s 5072 6991 5072 6991 4 gnd
rlabel metal3 s 4268 10158 4268 10158 4 gnd
rlabel metal3 s 17198 9368 17198 9368 4 gnd
rlabel metal3 s 7994 11544 7994 11544 4 gnd
rlabel metal3 s 14984 12156 14984 12156 4 gnd
rlabel metal3 s 11258 8147 11258 8147 4 gnd
rlabel metal3 s 14984 9786 14984 9786 4 gnd
rlabel metal3 s 18368 6991 18368 6991 4 gnd
rlabel metal3 s 4268 7788 4268 7788 4 gnd
rlabel metal3 s 14180 12521 14180 12521 4 gnd
rlabel metal3 s 11258 7910 11258 7910 4 gnd
rlabel metal3 s 2054 7788 2054 7788 4 gnd
rlabel metal3 s 5072 10151 5072 10151 4 gnd
rlabel metal3 s 14180 11336 14180 11336 4 gnd
rlabel metal3 s 4268 6998 4268 6998 4 gnd
rlabel metal3 s 4268 8996 4268 8996 4 gnd
rlabel metal3 s 11258 7594 11258 7594 4 gnd
rlabel metal3 s 7994 12887 7994 12887 4 gnd
rlabel metal3 s 4268 9786 4268 9786 4 gnd
rlabel metal3 s 9269 1578 9269 1578 4 gnd
rlabel metal3 s 16394 6991 16394 6991 4 gnd
rlabel metal3 s 7994 8384 7994 8384 4 gnd
rlabel metal3 s 11258 11070 11258 11070 4 gnd
rlabel metal3 s 9264 607 9264 607 4 gnd
rlabel metal3 s 2858 10151 2858 10151 4 gnd
rlabel metal3 s 7994 8147 7994 8147 4 gnd
rlabel metal3 s 11258 10517 11258 10517 4 gnd
rlabel metal3 s 11258 12887 11258 12887 4 gnd
rlabel metal3 s 4268 10948 4268 10948 4 gnd
rlabel metal3 s 11258 12334 11258 12334 4 gnd
rlabel metal3 s 11258 9727 11258 9727 4 gnd
rlabel metal3 s 14984 8206 14984 8206 4 gnd
rlabel metal3 s 14180 8571 14180 8571 4 gnd
rlabel metal3 s 11258 8700 11258 8700 4 gnd
rlabel metal3 s 7994 7357 7994 7357 4 gnd
rlabel metal3 s 5072 9361 5072 9361 4 gnd
rlabel metal3 s 11258 10280 11258 10280 4 gnd
rlabel metal3 s 2858 9361 2858 9361 4 gnd
rlabel metal3 s 14984 7416 14984 7416 4 gnd
rlabel metal3 s 7994 6567 7994 6567 4 gnd
rlabel metal3 s 4268 8206 4268 8206 4 gnd
rlabel metal3 s 14984 11738 14984 11738 4 gnd
rlabel metal3 s 9749 809 9749 809 4 gnd
rlabel metal3 s 14984 9368 14984 9368 4 gnd
rlabel metal3 s 14180 10151 14180 10151 4 gnd
rlabel metal3 s 7994 9174 7994 9174 4 gnd
rlabel metal3 s 7994 11070 7994 11070 4 gnd
rlabel metal3 s 7994 9490 7994 9490 4 gnd
rlabel metal3 s 7994 7910 7994 7910 4 gnd
rlabel metal3 s 17198 6998 17198 6998 4 gnd
rlabel metal3 s 5072 11336 5072 11336 4 gnd
rlabel metal3 s 7994 7120 7994 7120 4 gnd
rlabel metal3 s 14984 6998 14984 6998 4 gnd
rlabel metal3 s 11258 8937 11258 8937 4 gnd
rlabel metal3 s 4268 8578 4268 8578 4 gnd
rlabel metal3 s 12620 9727 12620 9727 4 gnd
rlabel metal3 s 7994 9727 7994 9727 4 gnd
rlabel metal3 s 4268 12528 4268 12528 4 gnd
rlabel metal3 s 4268 11738 4268 11738 4 gnd
rlabel metal3 s 2858 7781 2858 7781 4 gnd
rlabel metal3 s 7994 10754 7994 10754 4 gnd
rlabel metal3 s 2054 10158 2054 10158 4 gnd
rlabel metal3 s 14984 8996 14984 8996 4 gnd
rlabel metal3 s 9859 1578 9859 1578 4 gnd
rlabel metal3 s 4268 7416 4268 7416 4 gnd
rlabel metal3 s 9745 17083 9745 17083 4 gnd
rlabel metal3 s 5072 8571 5072 8571 4 gnd
rlabel metal3 s 884 6991 884 6991 4 gnd
rlabel metal3 s 5072 10546 5072 10546 4 gnd
rlabel metal3 s 11258 6567 11258 6567 4 gnd
rlabel metal3 s 11258 7357 11258 7357 4 gnd
rlabel metal3 s 14984 11366 14984 11366 4 gnd
rlabel metal3 s 11258 12650 11258 12650 4 gnd
rlabel metal3 s 14180 11731 14180 11731 4 gnd
rlabel metal3 s 7994 13124 7994 13124 4 gnd
rlabel metal3 s 11258 8384 11258 8384 4 gnd
rlabel metal3 s 14180 10546 14180 10546 4 gnd
rlabel metal3 s 5072 8966 5072 8966 4 gnd
rlabel metal3 s 5790 9712 5790 9712 4 gnd
rlabel metal3 s 9453 15149 9453 15149 4 gnd
rlabel metal3 s 17198 7788 17198 7788 4 gnd
rlabel metal3 s 7994 11860 7994 11860 4 gnd
rlabel metal3 s 7994 9964 7994 9964 4 gnd
rlabel metal3 s 2054 9368 2054 9368 4 gnd
rlabel metal3 s 7994 12650 7994 12650 4 gnd
rlabel metal3 s 2858 6991 2858 6991 4 gnd
rlabel metal3 s 14180 7781 14180 7781 4 gnd
rlabel metal3 s 18368 9361 18368 9361 4 gnd
rlabel metal3 s 5072 9756 5072 9756 4 gnd
rlabel metal3 s 7994 8937 7994 8937 4 gnd
rlabel metal3 s 5072 10941 5072 10941 4 gnd
rlabel metal3 s 11258 11860 11258 11860 4 gnd
rlabel metal3 s 7994 10517 7994 10517 4 gnd
rlabel metal3 s 11258 12097 11258 12097 4 gnd
rlabel metal3 s 9383 2371 9383 2371 4 gnd
rlabel metal3 s 9379 809 9379 809 4 gnd
rlabel metal3 s 4268 12156 4268 12156 4 gnd
rlabel metal3 s 14984 10948 14984 10948 4 gnd
rlabel metal3 s 6632 9727 6632 9727 4 gnd
rlabel metal3 s 14180 10941 14180 10941 4 gnd
rlabel metal3 s 16394 10151 16394 10151 4 gnd
rlabel metal3 s 14180 6991 14180 6991 4 gnd
rlabel metal3 s 11258 9964 11258 9964 4 gnd
rlabel metal3 s 11258 13124 11258 13124 4 gnd
rlabel metal3 s 7994 8700 7994 8700 4 gnd
rlabel metal3 s 7994 12334 7994 12334 4 gnd
rlabel metal3 s 5072 8176 5072 8176 4 gnd
rlabel metal3 s 11258 9174 11258 9174 4 gnd
rlabel metal3 s 11258 6330 11258 6330 4 gnd
rlabel metal3 s 11258 9490 11258 9490 4 gnd
rlabel metal3 s 5072 12521 5072 12521 4 gnd
rlabel metal3 s 13462 9712 13462 9712 4 gnd
rlabel metal3 s 7994 11307 7994 11307 4 gnd
rlabel metal3 s 14984 7788 14984 7788 4 gnd
rlabel metal3 s 5072 11731 5072 11731 4 gnd
rlabel metal3 s 4268 10576 4268 10576 4 gnd
rlabel metal3 s 11258 11544 11258 11544 4 gnd
rlabel metal3 s 14180 9361 14180 9361 4 gnd
rlabel metal3 s 5072 7781 5072 7781 4 gnd
rlabel metal3 s 9864 607 9864 607 4 gnd
rlabel metal3 s 14984 8578 14984 8578 4 gnd
rlabel metal3 s 14984 10158 14984 10158 4 gnd
rlabel metal3 s 17198 10158 17198 10158 4 gnd
rlabel metal3 s 9675 4305 9675 4305 4 gnd
rlabel metal3 s 11258 10754 11258 10754 4 gnd
rlabel metal3 s 4268 11366 4268 11366 4 gnd
rlabel metal3 s 11258 11307 11258 11307 4 gnd
rlabel metal3 s 9675 15149 9675 15149 4 gnd
rlabel metal3 s 14984 12528 14984 12528 4 gnd
rlabel metal3 s 7994 6804 7994 6804 4 gnd
rlabel metal3 s 884 9361 884 9361 4 gnd
rlabel metal3 s 5072 12126 5072 12126 4 gnd
rlabel metal3 s 14984 10576 14984 10576 4 gnd
rlabel metal3 s 14180 7386 14180 7386 4 gnd
rlabel metal3 s 11258 6804 11258 6804 4 gnd
rlabel metal3 s 14180 8176 14180 8176 4 gnd
rlabel metal3 s 5072 7386 5072 7386 4 gnd
rlabel metal3 s 2054 6998 2054 6998 4 gnd
rlabel metal3 s 7994 10280 7994 10280 4 gnd
rlabel metal3 s 9453 4305 9453 4305 4 gnd
rlabel metal3 s 14180 8966 14180 8966 4 gnd
rlabel metal3 s 4268 9368 4268 9368 4 gnd
rlabel metal3 s 14180 12126 14180 12126 4 gnd
rlabel metal3 s 14180 9756 14180 9756 4 gnd
rlabel metal3 s 7994 6330 7994 6330 4 gnd
rlabel metal3 s 16394 9361 16394 9361 4 gnd
rlabel metal3 s 7994 7594 7994 7594 4 gnd
rlabel metal3 s 16394 7781 16394 7781 4 gnd
rlabel metal2 s 11636 15161 11636 15161 4 wl_en1
rlabel metal2 s 7520 3203 7520 3203 4 wl_en0
rlabel metal1 s 9129 2390 9129 2390 4 dout0_0
rlabel metal1 s 32 8571 32 8571 4 addr0_0
rlabel metal2 s 7396 3203 7396 3203 4 p_en_bar0
rlabel metal1 s 112 8571 112 8571 4 addr0_1
rlabel metal3 s 14833 14807 14833 14807 4 rbl_bl1
rlabel metal2 s 7272 3203 7272 3203 4 w_en0
rlabel metal1 s 9287 32 9287 32 4 din0_0
rlabel metal1 s 19060 8571 19060 8571 4 addr1_2
rlabel metal1 s 19140 8571 19140 8571 4 addr1_1
rlabel metal2 s 7148 3203 7148 3203 4 s_en0
rlabel metal3 s 4693 10158 4693 10158 4 vdd
rlabel metal3 s 18096 6991 18096 6991 4 vdd
rlabel metal3 s 9314 13448 9314 13448 4 vdd
rlabel metal3 s 9195 5415 9195 5415 4 vdd
rlabel metal3 s 14559 7418 14559 7418 4 vdd
rlabel metal3 s 9870 1141 9870 1141 4 vdd
rlabel metal3 s 9745 16761 9745 16761 4 vdd
rlabel metal3 s 13908 11731 13908 11731 4 vdd
rlabel metal3 s 16773 10158 16773 10158 4 vdd
rlabel metal3 s 5344 11336 5344 11336 4 vdd
rlabel metal3 s 4693 7788 4693 7788 4 vdd
rlabel metal3 s 5344 8966 5344 8966 4 vdd
rlabel metal3 s 13908 6991 13908 6991 4 vdd
rlabel metal3 s 14559 10948 14559 10948 4 vdd
rlabel metal3 s 13908 8571 13908 8571 4 vdd
rlabel metal3 s 1156 9361 1156 9361 4 vdd
rlabel metal3 s 8809 5415 8809 5415 4 vdd
rlabel metal3 s 5344 11731 5344 11731 4 vdd
rlabel metal3 s 14559 10158 14559 10158 4 vdd
rlabel metal3 s 10562 13448 10562 13448 4 vdd
rlabel metal3 s 5344 9756 5344 9756 4 vdd
rlabel metal3 s 9314 6006 9314 6006 4 vdd
rlabel metal3 s 14559 8578 14559 8578 4 vdd
rlabel metal3 s 3130 9361 3130 9361 4 vdd
rlabel metal3 s 14559 11738 14559 11738 4 vdd
rlabel metal3 s 1156 6991 1156 6991 4 vdd
rlabel metal3 s 9278 191 9278 191 4 vdd
rlabel metal3 s 4693 11368 4693 11368 4 vdd
rlabel metal3 s 5344 10941 5344 10941 4 vdd
rlabel metal3 s 14559 7788 14559 7788 4 vdd
rlabel metal3 s 9371 15923 9371 15923 4 vdd
rlabel metal3 s 5344 8571 5344 8571 4 vdd
rlabel metal3 s 13037 9711 13037 9711 4 vdd
rlabel metal3 s 9383 16761 9383 16761 4 vdd
rlabel metal3 s 13908 10151 13908 10151 4 vdd
rlabel metal3 s 4693 9788 4693 9788 4 vdd
rlabel metal3 s 13908 8966 13908 8966 4 vdd
rlabel metal3 s 10057 5415 10057 5415 4 vdd
rlabel metal3 s 16773 6998 16773 6998 4 vdd
rlabel metal3 s 2479 10158 2479 10158 4 vdd
rlabel metal3 s 5344 8176 5344 8176 4 vdd
rlabel metal3 s 4693 12158 4693 12158 4 vdd
rlabel metal3 s 4693 12528 4693 12528 4 vdd
rlabel metal3 s 14559 12158 14559 12158 4 vdd
rlabel metal3 s 14559 8208 14559 8208 4 vdd
rlabel metal3 s 9938 6006 9938 6006 4 vdd
rlabel metal3 s 9757 3531 9757 3531 4 vdd
rlabel metal3 s 4693 8578 4693 8578 4 vdd
rlabel metal3 s 14559 9368 14559 9368 4 vdd
rlabel metal3 s 9757 15923 9757 15923 4 vdd
rlabel metal3 s 2479 7788 2479 7788 4 vdd
rlabel metal3 s 16122 7781 16122 7781 4 vdd
rlabel metal3 s 5344 7781 5344 7781 4 vdd
rlabel metal3 s 18096 9361 18096 9361 4 vdd
rlabel metal3 s 9850 191 9850 191 4 vdd
rlabel metal3 s 4693 9368 4693 9368 4 vdd
rlabel metal3 s 14559 6998 14559 6998 4 vdd
rlabel metal3 s 8690 6006 8690 6006 4 vdd
rlabel metal3 s 14559 9788 14559 9788 4 vdd
rlabel metal3 s 9195 14039 9195 14039 4 vdd
rlabel metal3 s 9745 2693 9745 2693 4 vdd
rlabel metal3 s 5344 10546 5344 10546 4 vdd
rlabel metal3 s 4693 10578 4693 10578 4 vdd
rlabel metal3 s 16122 6991 16122 6991 4 vdd
rlabel metal3 s 8690 13448 8690 13448 4 vdd
rlabel metal3 s 9258 1141 9258 1141 4 vdd
rlabel metal3 s 13908 9756 13908 9756 4 vdd
rlabel metal3 s 4693 11738 4693 11738 4 vdd
rlabel metal3 s 3130 10151 3130 10151 4 vdd
rlabel metal3 s 5344 10151 5344 10151 4 vdd
rlabel metal3 s 5344 12521 5344 12521 4 vdd
rlabel metal3 s 6215 9711 6215 9711 4 vdd
rlabel metal3 s 9938 13448 9938 13448 4 vdd
rlabel metal3 s 16122 9361 16122 9361 4 vdd
rlabel metal3 s 9371 3531 9371 3531 4 vdd
rlabel metal3 s 13908 9361 13908 9361 4 vdd
rlabel metal3 s 12122 9727 12122 9727 4 vdd
rlabel metal3 s 4693 6998 4693 6998 4 vdd
rlabel metal3 s 4693 7418 4693 7418 4 vdd
rlabel metal3 s 16122 10151 16122 10151 4 vdd
rlabel metal3 s 4693 8998 4693 8998 4 vdd
rlabel metal3 s 4693 10948 4693 10948 4 vdd
rlabel metal3 s 13908 10546 13908 10546 4 vdd
rlabel metal3 s 5344 12126 5344 12126 4 vdd
rlabel metal3 s 3130 7781 3130 7781 4 vdd
rlabel metal3 s 4693 8208 4693 8208 4 vdd
rlabel metal3 s 10443 14039 10443 14039 4 vdd
rlabel metal3 s 13908 7781 13908 7781 4 vdd
rlabel metal3 s 14559 10578 14559 10578 4 vdd
rlabel metal3 s 13908 12126 13908 12126 4 vdd
rlabel metal3 s 13908 12521 13908 12521 4 vdd
rlabel metal3 s 10562 6006 10562 6006 4 vdd
rlabel metal3 s 3130 6991 3130 6991 4 vdd
rlabel metal3 s 5344 7386 5344 7386 4 vdd
rlabel metal3 s 13908 11336 13908 11336 4 vdd
rlabel metal3 s 14559 8998 14559 8998 4 vdd
rlabel metal3 s 16773 7788 16773 7788 4 vdd
rlabel metal3 s 13908 10941 13908 10941 4 vdd
rlabel metal3 s 13908 7386 13908 7386 4 vdd
rlabel metal3 s 14559 12528 14559 12528 4 vdd
rlabel metal3 s 13908 8176 13908 8176 4 vdd
rlabel metal3 s 10057 14039 10057 14039 4 vdd
rlabel metal3 s 7130 9727 7130 9727 4 vdd
rlabel metal3 s 14559 11368 14559 11368 4 vdd
rlabel metal3 s 9383 2693 9383 2693 4 vdd
rlabel metal3 s 2479 9368 2479 9368 4 vdd
rlabel metal3 s 16773 9368 16773 9368 4 vdd
rlabel metal3 s 2479 6998 2479 6998 4 vdd
rlabel metal3 s 5344 9361 5344 9361 4 vdd
rlabel metal3 s 5344 6991 5344 6991 4 vdd
<< properties >>
string FIXED_BBOX 0 0 19336 17275
<< end >>
