* SPICE3 file created from replica_cell_6t.ext - technology: scmos

M1000 a_36_40# vdd vdd vdd pfet w=0.6u l=0.8u
+  ad=0.76p pd=3.6u as=2.76p ps=12.4u
** SOURCE/DRAIN TIED
M1001 vdd a_36_40# vdd vdd pfet w=0.8u l=0.6u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_36_40# vdd gnd gnd nfet w=1.6u l=0.4u
+  ad=2.4p pd=7.2u as=4.48p ps=12u
M1003 gnd a_36_40# vdd gnd nfet w=1.6u l=0.4u
+  ad=0p pd=0u as=3.04p ps=10.4u
M1004 a_36_40# wl bl gnd nfet w=0.8u l=0.4u
+  ad=0p pd=0u as=0.8p ps=3.6u
M1005 vdd wl br gnd nfet w=0.8u l=0.4u
+  ad=0p pd=0u as=0.8p ps=3.6u
C0 vdd 0 2.60fF
