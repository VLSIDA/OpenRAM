magic
tech sky130A
magscale 1 2
timestamp 1595931502
<< checkpaint >>
rect -1302 -1364 2550 1680
<< ndiffc >>
rect 404 378 438 380
rect 810 378 844 380
rect 596 221 599 253
rect 649 221 652 253
rect 42 94 76 96
rect 1172 94 1206 96
rect 42 62 76 64
rect 1172 62 1206 64
<< locali >>
rect 42 395 76 412
rect 404 395 438 410
rect 810 395 844 410
rect 1172 395 1206 412
rect -14 253 17 254
rect -14 221 0 253
rect -14 220 17 221
rect 107 213 109 241
rect 139 207 141 241
rect 339 233 341 267
rect 371 233 373 261
rect 463 253 497 254
rect 565 253 596 254
rect 652 253 683 254
rect 751 253 785 254
rect 875 233 877 261
rect 907 233 909 267
rect 1231 253 1262 254
rect 463 220 497 221
rect 565 220 596 221
rect 652 220 683 221
rect 751 220 785 221
rect 1107 207 1109 241
rect 1139 213 1141 241
rect 1248 221 1262 253
rect 1231 220 1262 221
<< metal1 >>
rect 78 0 114 395
rect 150 0 186 395
rect 222 79 258 420
rect 294 0 330 395
rect 366 0 402 395
rect 846 0 882 395
rect 918 0 954 395
rect 990 79 1026 420
rect 1062 0 1098 395
rect 1134 0 1170 395
<< metal2 >>
rect 0 323 1248 371
rect 186 199 294 275
rect 954 199 1062 275
rect 0 103 1248 151
rect 186 -55 294 55
rect 954 -55 1062 55
use dummy_cell_1rw_1r  dummy_cell_1rw_1r_0
timestamp 1595931502
transform -1 0 1248 0 1 0
box -42 -104 624 420
use dummy_cell_1rw_1r  dummy_cell_1rw_1r_1
timestamp 1595931502
transform 1 0 0 0 1 0
box -42 -104 624 420
<< labels >>
rlabel metal2 s 1008 237 1008 237 4 gnd
rlabel metal2 s 1008 0 1008 0 4 gnd
rlabel metal2 s 240 237 240 237 4 gnd
rlabel metal2 s 240 0 240 0 4 gnd
rlabel metal1 s 168 197 168 197 4 br0_0
rlabel metal1 s 1080 197 1080 197 4 br0_1
rlabel metal2 s 624 127 624 127 4 wl1_0
rlabel metal1 s 384 197 384 197 4 br1_0
rlabel metal1 s 936 197 936 197 4 bl1_1
rlabel metal2 s 624 347 624 347 4 wl0_0
rlabel metal1 s 96 197 96 197 4 bl0_0
rlabel metal1 s 312 197 312 197 4 bl1_0
rlabel metal1 s 864 197 864 197 4 br1_1
rlabel metal1 s 1152 197 1152 197 4 bl0_1
rlabel metal1 s 1008 249 1008 249 4 vdd
rlabel metal1 s 240 249 240 249 4 vdd
<< properties >>
string FIXED_BBOX 0 0 1248 395
<< end >>
