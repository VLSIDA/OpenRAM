
*********************** "cell_6t" ******************************
.SUBCKT cell_6t bl br wl vdd gnd
* SPICE3 file created from cell_6t.ext - technology: scmos

M1000 a_36_40# a_28_32# vdd vdd p w=0.6u l=0.8u
M1001 vdd a_36_40# a_28_32# vdd p w=0.6u l=0.8u
M1002 a_36_40# a_28_32# gnd gnd n w=1.6u l=0.4u
M1003 gnd a_36_40# a_28_32# gnd n w=1.6u l=0.4u
M1004 a_36_40# wl bl gnd n w=0.8u l=0.4u
M1005 a_28_32# wl br gnd n w=0.8u l=0.4u

.ENDS
