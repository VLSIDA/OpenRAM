VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO sram_2_16_scn4m_subm
   CLASS BLOCK ;
   SIZE 216.9 BY 423.6 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  180.9 56.6 181.7 57.4 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  202.7 56.6 203.5 57.4 ;
      END
   END din0[1]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  65.2 352.2 66.0 353.0 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  65.2 374.2 66.0 375.0 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  65.2 392.2 66.0 393.0 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  65.2 414.2 66.0 415.0 ;
      END
   END addr0[3]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  10.0 10.2 10.8 11.0 ;
      END
   END csb0
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  10.0 32.2 10.8 33.0 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  54.1 1.6 54.7 11.4 ;
      END
   END clk0
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER m2 ;
         RECT  187.5 119.8 188.3 122.8 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER m2 ;
         RECT  194.3 119.8 195.1 122.8 ;
      END
   END dout0[1]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER m3 ;
         RECT  196.8 307.7 197.4 308.3 ;
         LAYER m3 ;
         RECT  93.1 276.8 93.9 277.6 ;
         LAYER m3 ;
         RECT  176.4 203.7 177.0 204.3 ;
         LAYER m3 ;
         RECT  152.0 245.6 152.8 246.4 ;
         LAYER m3 ;
         RECT  0.0 60.0 214.8 61.2 ;
         LAYER m3 ;
         RECT  172.8 213.6 214.8 214.8 ;
         LAYER m3 ;
         RECT  69.6 343.2 169.2 344.4 ;
         LAYER m3 ;
         RECT  0.0 170.4 214.8 171.6 ;
         LAYER m3 ;
         RECT  2.7 262.0 3.5 262.8 ;
         LAYER m3 ;
         RECT  79.2 160.8 214.8 162.0 ;
         LAYER m4 ;
         RECT  55.2 0.0 56.4 421.2 ;
         LAYER m3 ;
         RECT  136.8 247.2 214.8 248.4 ;
         LAYER m3 ;
         RECT  23.2 340.4 24.0 341.2 ;
         LAYER m3 ;
         RECT  93.1 224.8 93.9 225.6 ;
         LAYER m4 ;
         RECT  108.0 0.0 109.2 421.2 ;
         LAYER m4 ;
         RECT  213.6 0.0 214.8 421.2 ;
         LAYER m3 ;
         RECT  203.6 349.3 204.2 349.9 ;
         LAYER m3 ;
         RECT  0.0 122.4 34.8 123.6 ;
         LAYER m4 ;
         RECT  194.4 0.0 195.6 421.2 ;
         LAYER m3 ;
         RECT  129.6 280.8 169.2 282.0 ;
         LAYER m3 ;
         RECT  0.0 160.8 73.2 162.0 ;
         LAYER m3 ;
         RECT  176.4 182.9 177.0 183.5 ;
         LAYER m3 ;
         RECT  197.2 166.8 198.0 167.6 ;
         LAYER m3 ;
         RECT  190.4 166.8 191.2 167.6 ;
         LAYER m3 ;
         RECT  203.6 307.7 204.2 308.3 ;
         LAYER m4 ;
         RECT  165.6 0.0 166.8 421.2 ;
         LAYER m3 ;
         RECT  196.8 349.3 197.4 349.9 ;
         LAYER m3 ;
         RECT  172.8 319.2 214.8 320.4 ;
         LAYER m4 ;
         RECT  36.0 0.0 37.2 421.2 ;
         LAYER m4 ;
         RECT  160.8 0.0 162.0 421.2 ;
         LAYER m3 ;
         RECT  0.0 21.6 214.8 22.8 ;
         LAYER m3 ;
         RECT  0.0 348.0 54.0 349.2 ;
         LAYER m3 ;
         RECT  0.0 132.0 214.8 133.2 ;
         LAYER m3 ;
         RECT  134.4 223.2 214.8 224.4 ;
         LAYER m3 ;
         RECT  2.7 183.6 3.5 184.4 ;
         LAYER m3 ;
         RECT  2.7 340.4 3.5 341.2 ;
         LAYER m3 ;
         RECT  0.0 88.8 75.6 90.0 ;
         LAYER m3 ;
         RECT  0.0 314.4 169.2 315.6 ;
         LAYER m3 ;
         RECT  203.6 266.1 204.2 266.7 ;
         LAYER m3 ;
         RECT  108.1 256.0 108.9 256.8 ;
         LAYER m3 ;
         RECT  196.8 224.5 197.4 225.1 ;
         LAYER m3 ;
         RECT  172.8 194.4 214.8 195.6 ;
         LAYER m3 ;
         RECT  129.6 252.0 169.2 253.2 ;
         LAYER m3 ;
         RECT  86.4 352.8 169.2 354.0 ;
         LAYER m3 ;
         RECT  176.4 224.5 177.0 225.1 ;
         LAYER m3 ;
         RECT  0.0 184.8 214.8 186.0 ;
         LAYER m3 ;
         RECT  0.0 93.6 188.4 94.8 ;
         LAYER m3 ;
         RECT  108.1 276.8 108.9 277.6 ;
         LAYER m3 ;
         RECT  132.0 204.0 214.8 205.2 ;
         LAYER m3 ;
         RECT  33.6 213.6 87.6 214.8 ;
         LAYER m3 ;
         RECT  0.0 218.4 116.4 219.6 ;
         LAYER m3 ;
         RECT  33.6 271.2 116.4 272.4 ;
         LAYER m3 ;
         RECT  176.4 328.5 177.0 329.1 ;
         LAYER m3 ;
         RECT  0.0 112.8 75.6 114.0 ;
         LAYER m3 ;
         RECT  190.1 98.6 190.9 99.4 ;
         LAYER m3 ;
         RECT  0.0 391.2 70.8 392.4 ;
         LAYER m4 ;
         RECT  84.0 0.0 85.2 421.2 ;
         LAYER m3 ;
         RECT  203.6 182.9 204.2 183.5 ;
         LAYER m3 ;
         RECT  77.6 141.2 78.4 142.0 ;
         LAYER m3 ;
         RECT  0.0 45.6 178.8 46.8 ;
         LAYER m3 ;
         RECT  33.6 290.4 169.2 291.6 ;
         LAYER m3 ;
         RECT  0.0 103.2 214.8 104.4 ;
         LAYER m4 ;
         RECT  199.2 0.0 200.4 421.2 ;
         LAYER m4 ;
         RECT  45.6 0.0 46.8 421.2 ;
         LAYER m3 ;
         RECT  0.0 386.4 214.8 387.6 ;
         LAYER m3 ;
         RECT  172.8 357.6 214.8 358.8 ;
         LAYER m3 ;
         RECT  176.4 245.3 177.0 245.9 ;
         LAYER m3 ;
         RECT  112.8 232.8 147.6 234.0 ;
         LAYER m3 ;
         RECT  52.8 12.0 214.8 13.2 ;
         LAYER m3 ;
         RECT  203.6 245.3 204.2 245.9 ;
         LAYER m4 ;
         RECT  112.8 0.0 114.0 421.2 ;
         LAYER m3 ;
         RECT  203.6 328.5 204.2 329.1 ;
         LAYER m3 ;
         RECT  0.0 180.0 214.8 181.2 ;
         LAYER m3 ;
         RECT  33.6 252.0 116.4 253.2 ;
         LAYER m3 ;
         RECT  0.0 146.4 188.4 147.6 ;
         LAYER m3 ;
         RECT  2.0 21.2 2.8 22.0 ;
         LAYER m3 ;
         RECT  0.0 295.2 147.6 296.4 ;
         LAYER m3 ;
         RECT  88.8 372.0 214.8 373.2 ;
         LAYER m3 ;
         RECT  93.1 256.0 93.9 256.8 ;
         LAYER m3 ;
         RECT  196.8 203.7 197.4 204.3 ;
         LAYER m3 ;
         RECT  190.0 370.1 190.6 370.7 ;
         LAYER m3 ;
         RECT  190.0 286.9 190.6 287.5 ;
         LAYER m3 ;
         RECT  183.1 224.4 183.9 225.2 ;
         LAYER m3 ;
         RECT  0.0 396.0 214.8 397.2 ;
         LAYER m3 ;
         RECT  0.0 16.8 214.8 18.0 ;
         LAYER m3 ;
         RECT  33.6 175.2 214.8 176.4 ;
         LAYER m3 ;
         RECT  190.0 307.7 190.6 308.3 ;
         LAYER m3 ;
         RECT  0.0 208.8 116.4 210.0 ;
         LAYER m3 ;
         RECT  26.4 242.4 214.8 243.6 ;
         LAYER m3 ;
         RECT  0.0 98.4 214.8 99.6 ;
         LAYER m3 ;
         RECT  33.6 194.4 87.6 195.6 ;
         LAYER m3 ;
         RECT  93.1 204.0 93.9 204.8 ;
         LAYER m3 ;
         RECT  0.0 237.6 214.8 238.8 ;
         LAYER m3 ;
         RECT  172.8 295.2 214.8 296.4 ;
         LAYER m3 ;
         RECT  190.0 266.1 190.6 266.7 ;
         LAYER m3 ;
         RECT  183.1 182.8 183.9 183.6 ;
         LAYER m3 ;
         RECT  0.0 420.0 214.8 421.2 ;
         LAYER m4 ;
         RECT  180.0 0.0 181.2 421.2 ;
         LAYER m3 ;
         RECT  0.0 247.2 87.6 248.4 ;
         LAYER m3 ;
         RECT  79.2 40.8 214.8 42.0 ;
         LAYER m3 ;
         RECT  0.0 400.8 214.8 402.0 ;
         LAYER m3 ;
         RECT  2.7 301.2 3.5 302.0 ;
         LAYER m3 ;
         RECT  152.0 328.8 152.8 329.6 ;
         LAYER m3 ;
         RECT  23.2 183.6 24.0 184.4 ;
         LAYER m3 ;
         RECT  0.0 333.6 169.2 334.8 ;
         LAYER m3 ;
         RECT  167.5 245.6 168.3 246.4 ;
         LAYER m3 ;
         RECT  129.6 271.2 169.2 272.4 ;
         LAYER m3 ;
         RECT  167.5 287.2 168.3 288.0 ;
         LAYER m3 ;
         RECT  68.1 363.2 68.9 364.0 ;
         LAYER m3 ;
         RECT  205.6 67.6 206.4 68.4 ;
         LAYER m4 ;
         RECT  12.0 0.0 13.2 421.2 ;
         LAYER m4 ;
         RECT  127.2 0.0 128.4 421.2 ;
         LAYER m3 ;
         RECT  167.5 349.6 168.3 350.4 ;
         LAYER m4 ;
         RECT  16.8 0.0 18.0 421.2 ;
         LAYER m3 ;
         RECT  0.0 31.2 214.8 32.4 ;
         LAYER m4 ;
         RECT  88.8 0.0 90.0 421.2 ;
         LAYER m3 ;
         RECT  199.1 132.6 199.9 133.4 ;
         LAYER m3 ;
         RECT  190.0 328.5 190.6 329.1 ;
         LAYER m4 ;
         RECT  136.8 0.0 138.0 421.2 ;
         LAYER m4 ;
         RECT  175.2 0.0 176.4 421.2 ;
         LAYER m3 ;
         RECT  4.8 40.8 73.2 42.0 ;
         LAYER m3 ;
         RECT  129.6 228.0 169.2 229.2 ;
         LAYER m3 ;
         RECT  112.8 285.6 214.8 286.8 ;
         LAYER m3 ;
         RECT  190.0 182.9 190.6 183.5 ;
         LAYER m3 ;
         RECT  23.2 222.8 24.0 223.6 ;
         LAYER m3 ;
         RECT  0.0 36.0 34.8 37.2 ;
         LAYER m3 ;
         RECT  172.8 232.8 214.8 234.0 ;
         LAYER m4 ;
         RECT  146.4 0.0 147.6 421.2 ;
         LAYER m3 ;
         RECT  196.8 370.1 197.4 370.7 ;
         LAYER m4 ;
         RECT  21.6 0.0 22.8 421.2 ;
         LAYER m3 ;
         RECT  0.0 108.0 183.6 109.2 ;
         LAYER m3 ;
         RECT  33.6 232.8 87.6 234.0 ;
         LAYER m3 ;
         RECT  129.6 261.6 169.2 262.8 ;
         LAYER m4 ;
         RECT  79.2 0.0 80.4 421.2 ;
         LAYER m3 ;
         RECT  203.6 203.7 204.2 204.3 ;
         LAYER m3 ;
         RECT  183.1 286.8 183.9 287.6 ;
         LAYER m3 ;
         RECT  196.8 182.9 197.4 183.5 ;
         LAYER m3 ;
         RECT  183.1 203.6 183.9 204.4 ;
         LAYER m3 ;
         RECT  23.2 301.2 24.0 302.0 ;
         LAYER m3 ;
         RECT  0.0 300.0 214.8 301.2 ;
         LAYER m3 ;
         RECT  203.6 370.1 204.2 370.7 ;
         LAYER m3 ;
         RECT  0.0 285.6 87.6 286.8 ;
         LAYER m4 ;
         RECT  60.0 0.0 61.2 421.2 ;
         LAYER m3 ;
         RECT  86.4 348.0 214.8 349.2 ;
         LAYER m3 ;
         RECT  0.0 372.0 70.8 373.2 ;
         LAYER m4 ;
         RECT  40.8 0.0 42.0 421.2 ;
         LAYER m3 ;
         RECT  33.6 328.8 214.8 330.0 ;
         LAYER m3 ;
         RECT  196.8 245.3 197.4 245.9 ;
         LAYER m3 ;
         RECT  0.0 74.4 214.8 75.6 ;
         LAYER m3 ;
         RECT  0.0 228.0 121.2 229.2 ;
         LAYER m4 ;
         RECT  122.4 0.0 123.6 421.2 ;
         LAYER m4 ;
         RECT  170.4 0.0 171.6 421.2 ;
         LAYER m4 ;
         RECT  2.4 0.0 3.6 421.2 ;
         LAYER m3 ;
         RECT  108.1 224.8 108.9 225.6 ;
         LAYER m3 ;
         RECT  33.6 309.6 214.8 310.8 ;
         LAYER m3 ;
         RECT  81.6 122.4 214.8 123.6 ;
         LAYER m3 ;
         RECT  196.8 266.1 197.4 266.7 ;
         LAYER m4 ;
         RECT  93.6 0.0 94.8 421.2 ;
         LAYER m3 ;
         RECT  77.6 61.2 78.4 62.0 ;
         LAYER m3 ;
         RECT  0.0 50.4 39.6 51.6 ;
         LAYER m3 ;
         RECT  26.4 319.2 147.6 320.4 ;
         LAYER m3 ;
         RECT  203.6 286.9 204.2 287.5 ;
         LAYER m3 ;
         RECT  196.8 286.9 197.4 287.5 ;
         LAYER m3 ;
         RECT  0.0 156.0 27.6 157.2 ;
         LAYER m4 ;
         RECT  50.4 0.0 51.6 421.2 ;
         LAYER m3 ;
         RECT  0.0 362.4 214.8 363.6 ;
         LAYER m3 ;
         RECT  167.5 204.0 168.3 204.8 ;
         LAYER m3 ;
         RECT  152.0 349.6 152.8 350.4 ;
         LAYER m3 ;
         RECT  0.0 199.2 116.4 200.4 ;
         LAYER m3 ;
         RECT  176.4 370.1 177.0 370.7 ;
         LAYER m3 ;
         RECT  0.0 117.6 214.8 118.8 ;
         LAYER m3 ;
         RECT  172.8 276.0 214.8 277.2 ;
         LAYER m3 ;
         RECT  190.0 349.3 190.6 349.9 ;
         LAYER m4 ;
         RECT  26.4 0.0 27.6 421.2 ;
         LAYER m4 ;
         RECT  208.8 0.0 210.0 421.2 ;
         LAYER m3 ;
         RECT  2.7 222.8 3.5 223.6 ;
         LAYER m3 ;
         RECT  172.8 151.2 214.8 152.4 ;
         LAYER m3 ;
         RECT  152.0 308.0 152.8 308.8 ;
         LAYER m3 ;
         RECT  192.3 132.6 193.1 133.4 ;
         LAYER m3 ;
         RECT  0.0 367.2 214.8 368.4 ;
         LAYER m3 ;
         RECT  0.0 141.6 214.8 142.8 ;
         LAYER m3 ;
         RECT  0.0 343.2 63.6 344.4 ;
         LAYER m3 ;
         RECT  72.0 381.6 214.8 382.8 ;
         LAYER m3 ;
         RECT  0.0 256.8 121.2 258.0 ;
         LAYER m3 ;
         RECT  0.0 7.2 214.8 8.4 ;
         LAYER m3 ;
         RECT  0.0 69.6 214.8 70.8 ;
         LAYER m4 ;
         RECT  132.0 0.0 133.2 421.2 ;
         LAYER m4 ;
         RECT  184.8 0.0 186.0 421.2 ;
         LAYER m4 ;
         RECT  64.8 0.0 66.0 421.2 ;
         LAYER m3 ;
         RECT  196.8 328.5 197.4 329.1 ;
         LAYER m3 ;
         RECT  0.0 151.2 75.6 152.4 ;
         LAYER m3 ;
         RECT  0.0 376.8 214.8 378.0 ;
         LAYER m3 ;
         RECT  183.1 328.4 183.9 329.2 ;
         LAYER m3 ;
         RECT  152.0 266.4 152.8 267.2 ;
         LAYER m3 ;
         RECT  190.0 245.3 190.6 245.9 ;
         LAYER m3 ;
         RECT  0.0 84.0 214.8 85.2 ;
         LAYER m3 ;
         RECT  0.0 189.6 169.2 190.8 ;
         LAYER m3 ;
         RECT  129.6 218.4 169.2 219.6 ;
         LAYER m4 ;
         RECT  69.6 0.0 70.8 421.2 ;
         LAYER m3 ;
         RECT  190.7 81.2 191.5 82.0 ;
         LAYER m3 ;
         RECT  0.0 338.4 147.6 339.6 ;
         LAYER m3 ;
         RECT  0.0 352.8 70.8 354.0 ;
         LAYER m3 ;
         RECT  0.0 415.2 214.8 416.4 ;
         LAYER m3 ;
         RECT  183.1 245.2 183.9 246.0 ;
         LAYER m3 ;
         RECT  0.0 26.4 214.8 27.6 ;
         LAYER m3 ;
         RECT  81.6 79.2 214.8 80.4 ;
         LAYER m3 ;
         RECT  0.0 410.4 214.8 411.6 ;
         LAYER m3 ;
         RECT  152.0 204.0 152.8 204.8 ;
         LAYER m3 ;
         RECT  183.8 67.6 184.6 68.4 ;
         LAYER m3 ;
         RECT  175.2 112.8 214.8 114.0 ;
         LAYER m3 ;
         RECT  176.4 307.7 177.0 308.3 ;
         LAYER m3 ;
         RECT  0.0 261.6 116.4 262.8 ;
         LAYER m3 ;
         RECT  0.0 276.0 121.2 277.2 ;
         LAYER m3 ;
         RECT  23.2 262.0 24.0 262.8 ;
         LAYER m3 ;
         RECT  91.2 391.2 214.8 392.4 ;
         LAYER m3 ;
         RECT  0.0 12.0 27.6 13.2 ;
         LAYER m3 ;
         RECT  0.0 127.2 214.8 128.4 ;
         LAYER m3 ;
         RECT  183.1 370.0 183.9 370.8 ;
         LAYER m3 ;
         RECT  81.6 2.4 214.8 3.6 ;
         LAYER m3 ;
         RECT  190.0 224.5 190.6 225.1 ;
         LAYER m3 ;
         RECT  196.9 98.6 197.7 99.4 ;
         LAYER m3 ;
         RECT  0.0 55.2 214.8 56.4 ;
         LAYER m3 ;
         RECT  0.0 79.2 73.2 80.4 ;
         LAYER m4 ;
         RECT  7.2 0.0 8.4 421.2 ;
         LAYER m4 ;
         RECT  151.2 0.0 152.4 421.2 ;
         LAYER m3 ;
         RECT  176.4 286.9 177.0 287.5 ;
         LAYER m3 ;
         RECT  77.6 101.2 78.4 102.0 ;
         LAYER m3 ;
         RECT  187.2 156.0 214.8 157.2 ;
         LAYER m3 ;
         RECT  129.6 199.2 169.2 200.4 ;
         LAYER m3 ;
         RECT  0.0 266.4 90.0 267.6 ;
         LAYER m3 ;
         RECT  68.1 403.2 68.9 404.0 ;
         LAYER m3 ;
         RECT  4.8 2.4 44.4 3.6 ;
         LAYER m4 ;
         RECT  117.6 0.0 118.8 421.2 ;
         LAYER m3 ;
         RECT  0.0 324.0 169.2 325.2 ;
         LAYER m3 ;
         RECT  0.0 304.8 214.8 306.0 ;
         LAYER m3 ;
         RECT  176.4 349.3 177.0 349.9 ;
         LAYER m3 ;
         RECT  167.5 266.4 168.3 267.2 ;
         LAYER m3 ;
         RECT  190.0 203.7 190.6 204.3 ;
         LAYER m3 ;
         RECT  172.8 338.4 214.8 339.6 ;
         LAYER m3 ;
         RECT  0.0 357.6 147.6 358.8 ;
         LAYER m4 ;
         RECT  31.2 0.0 32.4 421.2 ;
         LAYER m3 ;
         RECT  167.5 328.8 168.3 329.6 ;
         LAYER m4 ;
         RECT  74.4 0.0 75.6 421.2 ;
         LAYER m3 ;
         RECT  108.1 204.0 108.9 204.8 ;
         LAYER m4 ;
         RECT  98.4 0.0 99.6 421.2 ;
         LAYER m3 ;
         RECT  77.6 21.2 78.4 22.0 ;
         LAYER m3 ;
         RECT  197.5 81.2 198.3 82.0 ;
         LAYER m3 ;
         RECT  152.0 287.2 152.8 288.0 ;
         LAYER m3 ;
         RECT  0.0 64.8 214.8 66.0 ;
         LAYER m3 ;
         RECT  172.8 256.8 214.8 258.0 ;
         LAYER m3 ;
         RECT  0.0 381.6 63.6 382.8 ;
         LAYER m3 ;
         RECT  183.1 266.0 183.9 266.8 ;
         LAYER m3 ;
         RECT  183.1 307.6 183.9 308.4 ;
         LAYER m3 ;
         RECT  183.1 349.2 183.9 350.0 ;
         LAYER m3 ;
         RECT  26.4 165.6 214.8 166.8 ;
         LAYER m3 ;
         RECT  0.0 223.2 121.2 224.4 ;
         LAYER m4 ;
         RECT  204.0 0.0 205.2 421.2 ;
         LAYER m4 ;
         RECT  141.6 0.0 142.8 421.2 ;
         LAYER m4 ;
         RECT  156.0 0.0 157.2 421.2 ;
         LAYER m3 ;
         RECT  0.0 405.6 214.8 406.8 ;
         LAYER m3 ;
         RECT  139.2 266.4 214.8 267.6 ;
         LAYER m3 ;
         RECT  26.4 280.8 116.4 282.0 ;
         LAYER m3 ;
         RECT  203.6 224.5 204.2 225.1 ;
         LAYER m3 ;
         RECT  183.6 166.8 184.4 167.6 ;
         LAYER m3 ;
         RECT  0.0 136.8 214.8 138.0 ;
         LAYER m3 ;
         RECT  67.2 36.0 214.8 37.2 ;
         LAYER m4 ;
         RECT  103.2 0.0 104.4 421.2 ;
         LAYER m3 ;
         RECT  26.4 204.0 121.2 205.2 ;
         LAYER m3 ;
         RECT  167.5 224.8 168.3 225.6 ;
         LAYER m3 ;
         RECT  152.0 224.8 152.8 225.6 ;
         LAYER m3 ;
         RECT  129.6 208.8 169.2 210.0 ;
         LAYER m4 ;
         RECT  189.6 0.0 190.8 421.2 ;
         LAYER m3 ;
         RECT  176.4 266.1 177.0 266.7 ;
         LAYER m3 ;
         RECT  167.5 308.0 168.3 308.8 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER m3 ;
         RECT  179.8 333.5 180.4 334.1 ;
         LAYER m4 ;
         RECT  19.2 0.0 20.4 421.2 ;
         LAYER m3 ;
         RECT  200.2 219.5 200.8 220.1 ;
         LAYER m3 ;
         RECT  200.2 177.9 200.8 178.5 ;
         LAYER m3 ;
         RECT  200.2 312.7 200.8 313.3 ;
         LAYER m3 ;
         RECT  132.0 192.0 214.8 193.2 ;
         LAYER m3 ;
         RECT  0.0 91.2 75.6 92.4 ;
         LAYER m3 ;
         RECT  72.0 364.8 214.8 366.0 ;
         LAYER m3 ;
         RECT  186.5 229.4 187.3 230.2 ;
         LAYER m3 ;
         RECT  93.1 245.6 93.9 246.4 ;
         LAYER m3 ;
         RECT  200.2 187.9 200.8 188.5 ;
         LAYER m3 ;
         RECT  179.8 302.7 180.4 303.3 ;
         LAYER m3 ;
         RECT  0.0 388.8 214.8 390.0 ;
         LAYER m3 ;
         RECT  186.6 291.9 187.2 292.5 ;
         LAYER m3 ;
         RECT  141.6 278.4 214.8 279.6 ;
         LAYER m3 ;
         RECT  186.5 302.6 187.3 303.4 ;
         LAYER m3 ;
         RECT  0.0 345.6 54.0 346.8 ;
         LAYER m3 ;
         RECT  48.0 28.8 214.8 30.0 ;
         LAYER m3 ;
         RECT  0.0 393.6 70.8 394.8 ;
         LAYER m3 ;
         RECT  179.7 261.0 180.5 261.8 ;
         LAYER m4 ;
         RECT  129.6 0.0 130.8 421.2 ;
         LAYER m4 ;
         RECT  168.0 0.0 169.2 421.2 ;
         LAYER m4 ;
         RECT  134.4 0.0 135.6 421.2 ;
         LAYER m3 ;
         RECT  207.0 187.9 207.6 188.5 ;
         LAYER m3 ;
         RECT  68.1 423.2 68.9 424.0 ;
         LAYER m3 ;
         RECT  186.5 177.8 187.3 178.6 ;
         LAYER m3 ;
         RECT  186.5 250.2 187.3 251.0 ;
         LAYER m3 ;
         RECT  0.0 283.2 116.4 284.4 ;
         LAYER m3 ;
         RECT  179.8 177.9 180.4 178.5 ;
         LAYER m3 ;
         RECT  186.6 177.9 187.2 178.5 ;
         LAYER m3 ;
         RECT  200.1 146.0 200.9 146.8 ;
         LAYER m3 ;
         RECT  193.4 198.7 194.0 199.3 ;
         LAYER m3 ;
         RECT  173.0 177.9 173.6 178.5 ;
         LAYER m3 ;
         RECT  198.9 92.2 199.7 93.0 ;
         LAYER m4 ;
         RECT  187.2 0.0 188.4 421.2 ;
         LAYER m3 ;
         RECT  0.0 177.6 214.8 178.8 ;
         LAYER m4 ;
         RECT  62.4 0.0 63.6 421.2 ;
         LAYER m3 ;
         RECT  186.6 312.7 187.2 313.3 ;
         LAYER m3 ;
         RECT  167.5 297.6 168.3 298.4 ;
         LAYER m3 ;
         RECT  0.0 24.0 37.2 25.2 ;
         LAYER m3 ;
         RECT  207.0 302.7 207.6 303.3 ;
         LAYER m3 ;
         RECT  129.6 283.2 214.8 284.4 ;
         LAYER m3 ;
         RECT  207.0 198.7 207.6 199.3 ;
         LAYER m3 ;
         RECT  0.0 57.6 214.8 58.8 ;
         LAYER m4 ;
         RECT  192.0 0.0 193.2 421.2 ;
         LAYER m3 ;
         RECT  193.4 187.9 194.0 188.5 ;
         LAYER m3 ;
         RECT  179.7 333.4 180.5 334.2 ;
         LAYER m3 ;
         RECT  193.4 177.9 194.0 178.5 ;
         LAYER m3 ;
         RECT  179.7 240.2 180.5 241.0 ;
         LAYER m3 ;
         RECT  207.0 219.5 207.6 220.1 ;
         LAYER m3 ;
         RECT  2.7 164.0 3.5 164.8 ;
         LAYER m3 ;
         RECT  200.2 229.5 200.8 230.1 ;
         LAYER m3 ;
         RECT  112.8 201.6 147.6 202.8 ;
         LAYER m4 ;
         RECT  211.2 0.0 212.4 421.2 ;
         LAYER m3 ;
         RECT  200.2 261.1 200.8 261.7 ;
         LAYER m3 ;
         RECT  186.5 291.8 187.3 292.6 ;
         LAYER m3 ;
         RECT  108.1 266.4 108.9 267.2 ;
         LAYER m3 ;
         RECT  179.8 187.9 180.4 188.5 ;
         LAYER m3 ;
         RECT  152.0 339.2 152.8 340.0 ;
         LAYER m3 ;
         RECT  179.8 240.3 180.4 240.9 ;
         LAYER m3 ;
         RECT  0.0 76.8 214.8 78.0 ;
         LAYER m3 ;
         RECT  167.5 318.4 168.3 319.2 ;
         LAYER m3 ;
         RECT  0.0 14.4 27.6 15.6 ;
         LAYER m4 ;
         RECT  206.4 0.0 207.6 421.2 ;
         LAYER m3 ;
         RECT  167.5 193.6 168.3 194.4 ;
         LAYER m3 ;
         RECT  108.1 245.6 108.9 246.4 ;
         LAYER m3 ;
         RECT  179.7 229.4 180.5 230.2 ;
         LAYER m3 ;
         RECT  179.7 344.2 180.5 345.0 ;
         LAYER m3 ;
         RECT  179.8 271.1 180.4 271.7 ;
         LAYER m3 ;
         RECT  0.0 321.6 214.8 322.8 ;
         LAYER m3 ;
         RECT  207.0 261.1 207.6 261.7 ;
         LAYER m3 ;
         RECT  152.0 193.6 152.8 194.4 ;
         LAYER m3 ;
         RECT  0.0 129.6 214.8 130.8 ;
         LAYER m3 ;
         RECT  0.0 216.0 121.2 217.2 ;
         LAYER m3 ;
         RECT  91.2 412.8 214.8 414.0 ;
         LAYER m3 ;
         RECT  186.5 333.4 187.3 334.2 ;
         LAYER m3 ;
         RECT  152.0 256.0 152.8 256.8 ;
         LAYER m3 ;
         RECT  179.7 323.4 180.5 324.2 ;
         LAYER m3 ;
         RECT  0.0 403.2 63.6 404.4 ;
         LAYER m4 ;
         RECT  148.8 0.0 150.0 421.2 ;
         LAYER m4 ;
         RECT  76.8 0.0 78.0 421.2 ;
         LAYER m3 ;
         RECT  189.3 106.8 190.1 107.6 ;
         LAYER m3 ;
         RECT  0.0 43.2 214.8 44.4 ;
         LAYER m3 ;
         RECT  186.5 281.8 187.3 282.6 ;
         LAYER m4 ;
         RECT  201.6 0.0 202.8 421.2 ;
         LAYER m3 ;
         RECT  186.6 354.3 187.2 354.9 ;
         LAYER m3 ;
         RECT  200.2 281.9 200.8 282.5 ;
         LAYER m3 ;
         RECT  0.0 235.2 214.8 236.4 ;
         LAYER m3 ;
         RECT  69.6 403.2 214.8 404.4 ;
         LAYER m3 ;
         RECT  0.0 168.0 178.8 169.2 ;
         LAYER m3 ;
         RECT  26.4 264.0 147.6 265.2 ;
         LAYER m3 ;
         RECT  91.2 393.6 214.8 394.8 ;
         LAYER m3 ;
         RECT  179.8 208.7 180.4 209.3 ;
         LAYER m4 ;
         RECT  4.8 0.0 6.0 421.2 ;
         LAYER m4 ;
         RECT  120.0 0.0 121.2 421.2 ;
         LAYER m3 ;
         RECT  167.5 235.2 168.3 236.0 ;
         LAYER m3 ;
         RECT  23.2 281.6 24.0 282.4 ;
         LAYER m3 ;
         RECT  0.0 244.8 121.2 246.0 ;
         LAYER m4 ;
         RECT  14.4 0.0 15.6 421.2 ;
         LAYER m3 ;
         RECT  68.1 343.2 68.9 344.0 ;
         LAYER m3 ;
         RECT  33.6 292.8 214.8 294.0 ;
         LAYER m4 ;
         RECT  158.4 0.0 159.6 421.2 ;
         LAYER m3 ;
         RECT  179.7 219.4 180.5 220.2 ;
         LAYER m3 ;
         RECT  200.2 354.3 200.8 354.9 ;
         LAYER m3 ;
         RECT  193.4 354.3 194.0 354.9 ;
         LAYER m3 ;
         RECT  26.4 220.8 116.4 222.0 ;
         LAYER m3 ;
         RECT  179.8 250.3 180.4 250.9 ;
         LAYER m3 ;
         RECT  2.7 203.2 3.5 204.0 ;
         LAYER m3 ;
         RECT  2.7 320.8 3.5 321.6 ;
         LAYER m3 ;
         RECT  152.0 360.0 152.8 360.8 ;
         LAYER m3 ;
         RECT  179.8 198.7 180.4 199.3 ;
         LAYER m3 ;
         RECT  193.4 229.5 194.0 230.1 ;
         LAYER m3 ;
         RECT  183.8 47.6 184.6 48.4 ;
         LAYER m3 ;
         RECT  152.0 214.4 152.8 215.2 ;
         LAYER m3 ;
         RECT  33.6 312.0 214.8 313.2 ;
         LAYER m3 ;
         RECT  129.6 268.8 214.8 270.0 ;
         LAYER m3 ;
         RECT  193.4 312.7 194.0 313.3 ;
         LAYER m3 ;
         RECT  93.1 266.4 93.9 267.2 ;
         LAYER m3 ;
         RECT  173.0 208.7 173.6 209.3 ;
         LAYER m3 ;
         RECT  186.6 281.9 187.2 282.5 ;
         LAYER m3 ;
         RECT  179.7 302.6 180.5 303.4 ;
         LAYER m3 ;
         RECT  173.0 271.1 173.6 271.7 ;
         LAYER m3 ;
         RECT  0.0 417.6 214.8 418.8 ;
         LAYER m3 ;
         RECT  77.6 41.2 78.4 42.0 ;
         LAYER m3 ;
         RECT  0.0 86.4 214.8 87.6 ;
         LAYER m3 ;
         RECT  200.2 323.5 200.8 324.1 ;
         LAYER m3 ;
         RECT  108.1 287.2 108.9 288.0 ;
         LAYER m3 ;
         RECT  179.8 291.9 180.4 292.5 ;
         LAYER m3 ;
         RECT  0.0 67.2 178.8 68.4 ;
         LAYER m3 ;
         RECT  193.4 291.9 194.0 292.5 ;
         LAYER m3 ;
         RECT  26.4 340.8 214.8 342.0 ;
         LAYER m3 ;
         RECT  0.0 148.8 214.8 150.0 ;
         LAYER m3 ;
         RECT  0.0 153.6 214.8 154.8 ;
         LAYER m4 ;
         RECT  9.6 0.0 10.8 421.2 ;
         LAYER m3 ;
         RECT  0.0 72.0 75.6 73.2 ;
         LAYER m3 ;
         RECT  33.6 331.2 214.8 332.4 ;
         LAYER m3 ;
         RECT  179.8 344.3 180.4 344.9 ;
         LAYER m3 ;
         RECT  0.0 364.8 63.6 366.0 ;
         LAYER m3 ;
         RECT  23.2 164.0 24.0 164.8 ;
         LAYER m3 ;
         RECT  33.6 192.0 121.2 193.2 ;
         LAYER m3 ;
         RECT  129.6 206.4 214.8 207.6 ;
         LAYER m3 ;
         RECT  0.0 240.0 214.8 241.2 ;
         LAYER m3 ;
         RECT  0.0 360.0 214.8 361.2 ;
         LAYER m3 ;
         RECT  0.0 4.8 214.8 6.0 ;
         LAYER m4 ;
         RECT  110.4 0.0 111.6 421.2 ;
         LAYER m3 ;
         RECT  186.5 312.6 187.3 313.4 ;
         LAYER m3 ;
         RECT  186.5 208.6 187.3 209.4 ;
         LAYER m3 ;
         RECT  170.4 91.2 214.8 92.4 ;
         LAYER m3 ;
         RECT  173.0 323.5 173.6 324.1 ;
         LAYER m3 ;
         RECT  179.7 250.2 180.5 251.0 ;
         LAYER m3 ;
         RECT  186.6 229.5 187.2 230.1 ;
         LAYER m3 ;
         RECT  167.5 256.0 168.3 256.8 ;
         LAYER m3 ;
         RECT  0.0 307.2 147.6 308.4 ;
         LAYER m3 ;
         RECT  0.0 144.0 214.8 145.2 ;
         LAYER m4 ;
         RECT  172.8 0.0 174.0 421.2 ;
         LAYER m3 ;
         RECT  207.0 177.9 207.6 178.5 ;
         LAYER m3 ;
         RECT  179.8 323.5 180.4 324.1 ;
         LAYER m3 ;
         RECT  186.5 271.0 187.3 271.8 ;
         LAYER m3 ;
         RECT  179.7 365.0 180.5 365.8 ;
         LAYER m4 ;
         RECT  86.4 0.0 87.6 421.2 ;
         LAYER m3 ;
         RECT  200.2 302.7 200.8 303.3 ;
         LAYER m3 ;
         RECT  193.4 240.3 194.0 240.9 ;
         LAYER m3 ;
         RECT  81.6 19.2 214.8 20.4 ;
         LAYER m3 ;
         RECT  129.6 249.6 214.8 250.8 ;
         LAYER m3 ;
         RECT  200.2 271.1 200.8 271.7 ;
         LAYER m3 ;
         RECT  200.2 365.1 200.8 365.7 ;
         LAYER m3 ;
         RECT  179.7 208.6 180.5 209.4 ;
         LAYER m3 ;
         RECT  0.0 201.6 87.6 202.8 ;
         LAYER m3 ;
         RECT  179.7 312.6 180.5 313.4 ;
         LAYER m3 ;
         RECT  179.7 187.8 180.5 188.6 ;
         LAYER m3 ;
         RECT  77.6 81.2 78.4 82.0 ;
         LAYER m4 ;
         RECT  24.0 0.0 25.2 421.2 ;
         LAYER m3 ;
         RECT  193.4 323.5 194.0 324.1 ;
         LAYER m3 ;
         RECT  33.6 172.8 214.8 174.0 ;
         LAYER m3 ;
         RECT  0.0 268.8 121.2 270.0 ;
         LAYER m3 ;
         RECT  192.1 92.2 192.9 93.0 ;
         LAYER m3 ;
         RECT  0.0 412.8 70.8 414.0 ;
         LAYER m3 ;
         RECT  197.5 87.8 198.3 88.6 ;
         LAYER m3 ;
         RECT  179.7 281.8 180.5 282.6 ;
         LAYER m3 ;
         RECT  207.0 323.5 207.6 324.1 ;
         LAYER m3 ;
         RECT  86.4 345.6 214.8 346.8 ;
         LAYER m3 ;
         RECT  4.8 19.2 73.2 20.4 ;
         LAYER m3 ;
         RECT  193.4 208.7 194.0 209.3 ;
         LAYER m3 ;
         RECT  207.0 229.5 207.6 230.1 ;
         LAYER m4 ;
         RECT  153.6 0.0 154.8 421.2 ;
         LAYER m4 ;
         RECT  91.2 0.0 92.4 421.2 ;
         LAYER m3 ;
         RECT  0.0 316.8 214.8 318.0 ;
         LAYER m3 ;
         RECT  167.5 339.2 168.3 340.0 ;
         LAYER m3 ;
         RECT  190.7 87.8 191.5 88.6 ;
         LAYER m3 ;
         RECT  108.1 214.4 108.9 215.2 ;
         LAYER m3 ;
         RECT  0.0 206.4 121.2 207.6 ;
         LAYER m3 ;
         RECT  0.0 52.8 214.8 54.0 ;
         LAYER m3 ;
         RECT  0.0 369.6 171.6 370.8 ;
         LAYER m3 ;
         RECT  179.8 281.9 180.4 282.5 ;
         LAYER m3 ;
         RECT  108.1 235.2 108.9 236.0 ;
         LAYER m3 ;
         RECT  207.0 240.3 207.6 240.9 ;
         LAYER m3 ;
         RECT  77.6 121.2 78.4 122.0 ;
         LAYER m3 ;
         RECT  186.5 219.4 187.3 220.2 ;
         LAYER m4 ;
         RECT  38.4 0.0 39.6 421.2 ;
         LAYER m3 ;
         RECT  207.0 365.1 207.6 365.7 ;
         LAYER m3 ;
         RECT  129.6 230.4 214.8 231.6 ;
         LAYER m3 ;
         RECT  93.1 193.6 93.9 194.4 ;
         LAYER m3 ;
         RECT  173.0 250.3 173.6 250.9 ;
         LAYER m3 ;
         RECT  207.0 333.5 207.6 334.1 ;
         LAYER m3 ;
         RECT  0.0 249.6 116.4 250.8 ;
         LAYER m3 ;
         RECT  207.0 281.9 207.6 282.5 ;
         LAYER m3 ;
         RECT  81.6 139.2 214.8 140.4 ;
         LAYER m4 ;
         RECT  196.8 0.0 198.0 421.2 ;
         LAYER m3 ;
         RECT  0.0 124.8 214.8 126.0 ;
         LAYER m3 ;
         RECT  186.6 219.5 187.2 220.1 ;
         LAYER m3 ;
         RECT  152.0 235.2 152.8 236.0 ;
         LAYER m3 ;
         RECT  207.0 291.9 207.6 292.5 ;
         LAYER m3 ;
         RECT  23.2 320.8 24.0 321.6 ;
         LAYER m3 ;
         RECT  179.7 271.0 180.5 271.8 ;
         LAYER m3 ;
         RECT  26.4 182.4 171.6 183.6 ;
         LAYER m4 ;
         RECT  52.8 0.0 54.0 421.2 ;
         LAYER m3 ;
         RECT  207.0 312.7 207.6 313.3 ;
         LAYER m3 ;
         RECT  186.6 365.1 187.2 365.7 ;
         LAYER m3 ;
         RECT  193.4 219.5 194.0 220.1 ;
         LAYER m3 ;
         RECT  193.4 281.9 194.0 282.5 ;
         LAYER m4 ;
         RECT  0.0 0.0 1.2 421.2 ;
         LAYER m3 ;
         RECT  173.0 240.3 173.6 240.9 ;
         LAYER m3 ;
         RECT  136.8 254.4 214.8 255.6 ;
         LAYER m3 ;
         RECT  0.0 297.6 214.8 298.8 ;
         LAYER m3 ;
         RECT  179.8 229.5 180.4 230.1 ;
         LAYER m3 ;
         RECT  193.4 250.3 194.0 250.9 ;
         LAYER m3 ;
         RECT  52.8 14.4 214.8 15.6 ;
         LAYER m3 ;
         RECT  0.0 187.2 214.8 188.4 ;
         LAYER m3 ;
         RECT  179.7 177.8 180.5 178.6 ;
         LAYER m3 ;
         RECT  74.4 24.0 214.8 25.2 ;
         LAYER m3 ;
         RECT  0.0 48.0 214.8 49.2 ;
         LAYER m3 ;
         RECT  173.0 261.1 173.6 261.7 ;
         LAYER m3 ;
         RECT  77.6 161.2 78.4 162.0 ;
         LAYER m4 ;
         RECT  81.6 0.0 82.8 421.2 ;
         LAYER m3 ;
         RECT  93.1 214.4 93.9 215.2 ;
         LAYER m3 ;
         RECT  186.5 365.0 187.3 365.8 ;
         LAYER m3 ;
         RECT  0.0 196.8 116.4 198.0 ;
         LAYER m4 ;
         RECT  67.2 0.0 68.4 421.2 ;
         LAYER m3 ;
         RECT  0.0 9.6 214.8 10.8 ;
         LAYER m3 ;
         RECT  186.5 354.2 187.3 355.0 ;
         LAYER m3 ;
         RECT  2.0 41.2 2.8 42.0 ;
         LAYER m3 ;
         RECT  200.2 208.7 200.8 209.3 ;
         LAYER m3 ;
         RECT  193.4 261.1 194.0 261.7 ;
         LAYER m3 ;
         RECT  186.6 333.5 187.2 334.1 ;
         LAYER m3 ;
         RECT  0.0 379.2 214.8 380.4 ;
         LAYER m3 ;
         RECT  2.0 1.2 2.8 2.0 ;
         LAYER m3 ;
         RECT  0.0 96.0 214.8 97.2 ;
         LAYER m3 ;
         RECT  167.5 276.8 168.3 277.6 ;
         LAYER m3 ;
         RECT  193.4 271.1 194.0 271.7 ;
         LAYER m4 ;
         RECT  43.2 0.0 44.4 421.2 ;
         LAYER m3 ;
         RECT  193.3 146.0 194.1 146.8 ;
         LAYER m3 ;
         RECT  186.6 208.7 187.2 209.3 ;
         LAYER m3 ;
         RECT  186.5 198.6 187.3 199.4 ;
         LAYER m3 ;
         RECT  108.1 193.6 108.9 194.4 ;
         LAYER m3 ;
         RECT  23.2 242.4 24.0 243.2 ;
         LAYER m3 ;
         RECT  2.7 242.4 3.5 243.2 ;
         LAYER m3 ;
         RECT  186.6 344.3 187.2 344.9 ;
         LAYER m3 ;
         RECT  0.0 288.0 147.6 289.2 ;
         LAYER m3 ;
         RECT  179.7 198.6 180.5 199.4 ;
         LAYER m3 ;
         RECT  0.0 230.4 116.4 231.6 ;
         LAYER m3 ;
         RECT  0.0 384.0 214.8 385.2 ;
         LAYER m3 ;
         RECT  179.8 312.7 180.4 313.3 ;
         LAYER m3 ;
         RECT  0.0 115.2 214.8 116.4 ;
         LAYER m3 ;
         RECT  173.0 229.5 173.6 230.1 ;
         LAYER m4 ;
         RECT  100.8 0.0 102.0 421.2 ;
         LAYER m3 ;
         RECT  200.2 344.3 200.8 344.9 ;
         LAYER m3 ;
         RECT  173.0 187.9 173.6 188.5 ;
         LAYER m3 ;
         RECT  67.2 33.6 214.8 34.8 ;
         LAYER m3 ;
         RECT  186.6 187.9 187.2 188.5 ;
         LAYER m3 ;
         RECT  186.6 198.7 187.2 199.3 ;
         LAYER m3 ;
         RECT  93.1 287.2 93.9 288.0 ;
         LAYER m3 ;
         RECT  129.6 220.8 214.8 222.0 ;
         LAYER m3 ;
         RECT  173.0 344.3 173.6 344.9 ;
         LAYER m3 ;
         RECT  173.0 198.7 173.6 199.3 ;
         LAYER m4 ;
         RECT  163.2 0.0 164.4 421.2 ;
         LAYER m3 ;
         RECT  0.0 139.2 73.2 140.4 ;
         LAYER m3 ;
         RECT  200.2 291.9 200.8 292.5 ;
         LAYER m3 ;
         RECT  173.0 365.1 173.6 365.7 ;
         LAYER m4 ;
         RECT  33.6 0.0 34.8 421.2 ;
         LAYER m3 ;
         RECT  152.0 297.6 152.8 298.4 ;
         LAYER m3 ;
         RECT  0.0 28.8 27.6 30.0 ;
         LAYER m3 ;
         RECT  186.6 302.7 187.2 303.3 ;
         LAYER m3 ;
         RECT  196.1 106.8 196.9 107.6 ;
         LAYER m3 ;
         RECT  193.4 302.7 194.0 303.3 ;
         LAYER m3 ;
         RECT  0.0 398.4 214.8 399.6 ;
         LAYER m3 ;
         RECT  0.0 254.4 87.6 255.6 ;
         LAYER m3 ;
         RECT  186.6 261.1 187.2 261.7 ;
         LAYER m4 ;
         RECT  28.8 0.0 30.0 421.2 ;
         LAYER m3 ;
         RECT  186.5 344.2 187.3 345.0 ;
         LAYER m3 ;
         RECT  0.0 350.4 147.6 351.6 ;
         LAYER m3 ;
         RECT  93.1 235.2 93.9 236.0 ;
         LAYER m3 ;
         RECT  173.0 333.5 173.6 334.1 ;
         LAYER m3 ;
         RECT  134.4 216.0 214.8 217.2 ;
         LAYER m4 ;
         RECT  48.0 0.0 49.2 421.2 ;
         LAYER m4 ;
         RECT  144.0 0.0 145.2 421.2 ;
         LAYER m3 ;
         RECT  0.0 0.0 214.8 1.2 ;
         LAYER m3 ;
         RECT  0.0 158.4 214.8 159.6 ;
         LAYER m4 ;
         RECT  105.6 0.0 106.8 421.2 ;
         LAYER m3 ;
         RECT  129.6 259.2 214.8 260.4 ;
         LAYER m3 ;
         RECT  167.5 214.4 168.3 215.2 ;
         LAYER m3 ;
         RECT  186.5 323.4 187.3 324.2 ;
         LAYER m4 ;
         RECT  115.2 0.0 116.4 421.2 ;
         LAYER m3 ;
         RECT  179.7 354.2 180.5 355.0 ;
         LAYER m3 ;
         RECT  33.6 273.6 214.8 274.8 ;
         LAYER m3 ;
         RECT  186.6 250.3 187.2 250.9 ;
         LAYER m3 ;
         RECT  0.0 100.8 73.2 102.0 ;
         LAYER m3 ;
         RECT  0.0 120.0 214.8 121.2 ;
         LAYER m3 ;
         RECT  79.2 100.8 214.8 102.0 ;
         LAYER m3 ;
         RECT  0.0 134.4 188.4 135.6 ;
         LAYER m3 ;
         RECT  175.2 72.0 214.8 73.2 ;
         LAYER m3 ;
         RECT  186.5 240.2 187.3 241.0 ;
         LAYER m3 ;
         RECT  0.0 374.4 70.8 375.6 ;
         LAYER m3 ;
         RECT  173.0 281.9 173.6 282.5 ;
         LAYER m3 ;
         RECT  173.0 302.7 173.6 303.3 ;
         LAYER m3 ;
         RECT  200.2 250.3 200.8 250.9 ;
         LAYER m3 ;
         RECT  173.0 219.5 173.6 220.1 ;
         LAYER m3 ;
         RECT  152.0 276.8 152.8 277.6 ;
         LAYER m3 ;
         RECT  81.6 62.4 214.8 63.6 ;
         LAYER m4 ;
         RECT  57.6 0.0 58.8 421.2 ;
         LAYER m3 ;
         RECT  77.6 1.2 78.4 2.0 ;
         LAYER m3 ;
         RECT  175.2 110.4 214.8 111.6 ;
         LAYER m3 ;
         RECT  193.4 365.1 194.0 365.7 ;
         LAYER m3 ;
         RECT  23.2 203.2 24.0 204.0 ;
         LAYER m3 ;
         RECT  186.5 187.8 187.3 188.6 ;
         LAYER m3 ;
         RECT  179.8 261.1 180.4 261.7 ;
         LAYER m3 ;
         RECT  179.7 291.8 180.5 292.6 ;
         LAYER m3 ;
         RECT  186.6 323.5 187.2 324.1 ;
         LAYER m3 ;
         RECT  179.8 354.3 180.4 354.9 ;
         LAYER m3 ;
         RECT  0.0 62.4 73.2 63.6 ;
         LAYER m3 ;
         RECT  167.5 360.0 168.3 360.8 ;
         LAYER m3 ;
         RECT  0.0 278.4 87.6 279.6 ;
         LAYER m3 ;
         RECT  186.6 271.1 187.2 271.7 ;
         LAYER m3 ;
         RECT  179.8 219.5 180.4 220.1 ;
         LAYER m3 ;
         RECT  205.6 47.6 206.4 48.4 ;
         LAYER m3 ;
         RECT  173.0 354.3 173.6 354.9 ;
         LAYER m3 ;
         RECT  2.7 281.6 3.5 282.4 ;
         LAYER m4 ;
         RECT  177.6 0.0 178.8 421.2 ;
         LAYER m4 ;
         RECT  96.0 0.0 97.2 421.2 ;
         LAYER m3 ;
         RECT  173.0 291.9 173.6 292.5 ;
         LAYER m3 ;
         RECT  200.2 198.7 200.8 199.3 ;
         LAYER m3 ;
         RECT  207.0 344.3 207.6 344.9 ;
         LAYER m3 ;
         RECT  88.8 374.4 214.8 375.6 ;
         LAYER m3 ;
         RECT  207.0 250.3 207.6 250.9 ;
         LAYER m3 ;
         RECT  26.4 302.4 214.8 303.6 ;
         LAYER m4 ;
         RECT  182.4 0.0 183.6 421.2 ;
         LAYER m3 ;
         RECT  0.0 225.6 87.6 226.8 ;
         LAYER m3 ;
         RECT  0.0 259.2 121.2 260.4 ;
         LAYER m3 ;
         RECT  0.0 110.4 75.6 111.6 ;
         LAYER m4 ;
         RECT  139.2 0.0 140.4 421.2 ;
         LAYER m3 ;
         RECT  0.0 105.6 214.8 106.8 ;
         LAYER m3 ;
         RECT  200.2 240.3 200.8 240.9 ;
         LAYER m3 ;
         RECT  0.0 408.0 214.8 409.2 ;
         LAYER m3 ;
         RECT  0.0 33.6 34.8 34.8 ;
         LAYER m3 ;
         RECT  207.0 354.3 207.6 354.9 ;
         LAYER m3 ;
         RECT  186.5 261.0 187.3 261.8 ;
         LAYER m3 ;
         RECT  173.0 312.7 173.6 313.3 ;
         LAYER m3 ;
         RECT  207.0 208.7 207.6 209.3 ;
         LAYER m3 ;
         RECT  193.4 344.3 194.0 344.9 ;
         LAYER m3 ;
         RECT  129.6 196.8 214.8 198.0 ;
         LAYER m4 ;
         RECT  72.0 0.0 73.2 421.2 ;
         LAYER m3 ;
         RECT  200.2 333.5 200.8 334.1 ;
         LAYER m3 ;
         RECT  0.0 355.2 214.8 356.4 ;
         LAYER m3 ;
         RECT  207.0 271.1 207.6 271.7 ;
         LAYER m3 ;
         RECT  33.6 211.2 214.8 212.4 ;
         LAYER m3 ;
         RECT  0.0 336.0 214.8 337.2 ;
         LAYER m3 ;
         RECT  179.8 365.1 180.4 365.7 ;
         LAYER m3 ;
         RECT  0.0 81.6 186.0 82.8 ;
         LAYER m4 ;
         RECT  124.8 0.0 126.0 421.2 ;
         LAYER m3 ;
         RECT  193.4 333.5 194.0 334.1 ;
         LAYER m3 ;
         RECT  0.0 163.2 214.8 164.4 ;
         LAYER m3 ;
         RECT  186.6 240.3 187.2 240.9 ;
         LAYER m3 ;
         RECT  0.0 326.4 147.6 327.6 ;
         LAYER m3 ;
         RECT  68.1 383.2 68.9 384.0 ;
         LAYER m3 ;
         RECT  152.0 318.4 152.8 319.2 ;
         LAYER m3 ;
         RECT  0.0 38.4 214.8 39.6 ;
      END
   END gnd
   OBS
   LAYER  m1 ;
      RECT  188.9 197.6 189.9 198.4 ;
      RECT  191.3 202.0 192.3 202.8 ;
      RECT  191.5 198.4 192.3 198.8 ;
      RECT  190.3 196.6 191.1 196.8 ;
      RECT  193.3 197.2 194.1 201.4 ;
      RECT  189.1 200.6 190.7 201.4 ;
      RECT  191.5 197.6 192.5 198.4 ;
      RECT  186.5 203.6 194.1 204.4 ;
      RECT  186.5 202.0 187.3 203.6 ;
      RECT  189.1 202.0 190.1 202.8 ;
      RECT  189.1 201.4 189.9 202.0 ;
      RECT  191.5 199.6 192.3 202.0 ;
      RECT  191.1 198.8 192.3 199.6 ;
      RECT  186.5 195.8 194.1 196.6 ;
      RECT  186.5 197.2 187.3 201.4 ;
      RECT  189.1 198.4 189.9 200.6 ;
      RECT  190.9 194.4 192.5 195.2 ;
      RECT  193.3 202.0 194.1 203.6 ;
      RECT  188.1 194.4 189.7 195.2 ;
      RECT  188.9 210.4 189.9 209.6 ;
      RECT  191.3 206.0 192.3 205.2 ;
      RECT  191.5 209.6 192.3 209.2 ;
      RECT  190.3 211.4 191.1 211.2 ;
      RECT  193.3 210.8 194.1 206.6 ;
      RECT  189.1 207.4 190.7 206.6 ;
      RECT  191.5 210.4 192.5 209.6 ;
      RECT  186.5 204.4 194.1 203.6 ;
      RECT  186.5 206.0 187.3 204.4 ;
      RECT  189.1 206.0 190.1 205.2 ;
      RECT  189.1 206.6 189.9 206.0 ;
      RECT  191.5 208.4 192.3 206.0 ;
      RECT  191.1 209.2 192.3 208.4 ;
      RECT  186.5 212.2 194.1 211.4 ;
      RECT  186.5 210.8 187.3 206.6 ;
      RECT  189.1 209.6 189.9 207.4 ;
      RECT  190.9 213.6 192.5 212.8 ;
      RECT  193.3 206.0 194.1 204.4 ;
      RECT  188.1 213.6 189.7 212.8 ;
      RECT  188.9 218.4 189.9 219.2 ;
      RECT  191.3 222.8 192.3 223.6 ;
      RECT  191.5 219.2 192.3 219.6 ;
      RECT  190.3 217.4 191.1 217.6 ;
      RECT  193.3 218.0 194.1 222.2 ;
      RECT  189.1 221.4 190.7 222.2 ;
      RECT  191.5 218.4 192.5 219.2 ;
      RECT  186.5 224.4 194.1 225.2 ;
      RECT  186.5 222.8 187.3 224.4 ;
      RECT  189.1 222.8 190.1 223.6 ;
      RECT  189.1 222.2 189.9 222.8 ;
      RECT  191.5 220.4 192.3 222.8 ;
      RECT  191.1 219.6 192.3 220.4 ;
      RECT  186.5 216.6 194.1 217.4 ;
      RECT  186.5 218.0 187.3 222.2 ;
      RECT  189.1 219.2 189.9 221.4 ;
      RECT  190.9 215.2 192.5 216.0 ;
      RECT  193.3 222.8 194.1 224.4 ;
      RECT  188.1 215.2 189.7 216.0 ;
      RECT  188.9 231.2 189.9 230.4 ;
      RECT  191.3 226.8 192.3 226.0 ;
      RECT  191.5 230.4 192.3 230.0 ;
      RECT  190.3 232.2 191.1 232.0 ;
      RECT  193.3 231.6 194.1 227.4 ;
      RECT  189.1 228.2 190.7 227.4 ;
      RECT  191.5 231.2 192.5 230.4 ;
      RECT  186.5 225.2 194.1 224.4 ;
      RECT  186.5 226.8 187.3 225.2 ;
      RECT  189.1 226.8 190.1 226.0 ;
      RECT  189.1 227.4 189.9 226.8 ;
      RECT  191.5 229.2 192.3 226.8 ;
      RECT  191.1 230.0 192.3 229.2 ;
      RECT  186.5 233.0 194.1 232.2 ;
      RECT  186.5 231.6 187.3 227.4 ;
      RECT  189.1 230.4 189.9 228.2 ;
      RECT  190.9 234.4 192.5 233.6 ;
      RECT  193.3 226.8 194.1 225.2 ;
      RECT  188.1 234.4 189.7 233.6 ;
      RECT  188.9 239.2 189.9 240.0 ;
      RECT  191.3 243.6 192.3 244.4 ;
      RECT  191.5 240.0 192.3 240.4 ;
      RECT  190.3 238.2 191.1 238.4 ;
      RECT  193.3 238.8 194.1 243.0 ;
      RECT  189.1 242.2 190.7 243.0 ;
      RECT  191.5 239.2 192.5 240.0 ;
      RECT  186.5 245.2 194.1 246.0 ;
      RECT  186.5 243.6 187.3 245.2 ;
      RECT  189.1 243.6 190.1 244.4 ;
      RECT  189.1 243.0 189.9 243.6 ;
      RECT  191.5 241.2 192.3 243.6 ;
      RECT  191.1 240.4 192.3 241.2 ;
      RECT  186.5 237.4 194.1 238.2 ;
      RECT  186.5 238.8 187.3 243.0 ;
      RECT  189.1 240.0 189.9 242.2 ;
      RECT  190.9 236.0 192.5 236.8 ;
      RECT  193.3 243.6 194.1 245.2 ;
      RECT  188.1 236.0 189.7 236.8 ;
      RECT  188.9 252.0 189.9 251.2 ;
      RECT  191.3 247.6 192.3 246.8 ;
      RECT  191.5 251.2 192.3 250.8 ;
      RECT  190.3 253.0 191.1 252.8 ;
      RECT  193.3 252.4 194.1 248.2 ;
      RECT  189.1 249.0 190.7 248.2 ;
      RECT  191.5 252.0 192.5 251.2 ;
      RECT  186.5 246.0 194.1 245.2 ;
      RECT  186.5 247.6 187.3 246.0 ;
      RECT  189.1 247.6 190.1 246.8 ;
      RECT  189.1 248.2 189.9 247.6 ;
      RECT  191.5 250.0 192.3 247.6 ;
      RECT  191.1 250.8 192.3 250.0 ;
      RECT  186.5 253.8 194.1 253.0 ;
      RECT  186.5 252.4 187.3 248.2 ;
      RECT  189.1 251.2 189.9 249.0 ;
      RECT  190.9 255.2 192.5 254.4 ;
      RECT  193.3 247.6 194.1 246.0 ;
      RECT  188.1 255.2 189.7 254.4 ;
      RECT  188.9 260.0 189.9 260.8 ;
      RECT  191.3 264.4 192.3 265.2 ;
      RECT  191.5 260.8 192.3 261.2 ;
      RECT  190.3 259.0 191.1 259.2 ;
      RECT  193.3 259.6 194.1 263.8 ;
      RECT  189.1 263.0 190.7 263.8 ;
      RECT  191.5 260.0 192.5 260.8 ;
      RECT  186.5 266.0 194.1 266.8 ;
      RECT  186.5 264.4 187.3 266.0 ;
      RECT  189.1 264.4 190.1 265.2 ;
      RECT  189.1 263.8 189.9 264.4 ;
      RECT  191.5 262.0 192.3 264.4 ;
      RECT  191.1 261.2 192.3 262.0 ;
      RECT  186.5 258.2 194.1 259.0 ;
      RECT  186.5 259.6 187.3 263.8 ;
      RECT  189.1 260.8 189.9 263.0 ;
      RECT  190.9 256.8 192.5 257.6 ;
      RECT  193.3 264.4 194.1 266.0 ;
      RECT  188.1 256.8 189.7 257.6 ;
      RECT  188.9 272.8 189.9 272.0 ;
      RECT  191.3 268.4 192.3 267.6 ;
      RECT  191.5 272.0 192.3 271.6 ;
      RECT  190.3 273.8 191.1 273.6 ;
      RECT  193.3 273.2 194.1 269.0 ;
      RECT  189.1 269.8 190.7 269.0 ;
      RECT  191.5 272.8 192.5 272.0 ;
      RECT  186.5 266.8 194.1 266.0 ;
      RECT  186.5 268.4 187.3 266.8 ;
      RECT  189.1 268.4 190.1 267.6 ;
      RECT  189.1 269.0 189.9 268.4 ;
      RECT  191.5 270.8 192.3 268.4 ;
      RECT  191.1 271.6 192.3 270.8 ;
      RECT  186.5 274.6 194.1 273.8 ;
      RECT  186.5 273.2 187.3 269.0 ;
      RECT  189.1 272.0 189.9 269.8 ;
      RECT  190.9 276.0 192.5 275.2 ;
      RECT  193.3 268.4 194.1 266.8 ;
      RECT  188.1 276.0 189.7 275.2 ;
      RECT  188.9 280.8 189.9 281.6 ;
      RECT  191.3 285.2 192.3 286.0 ;
      RECT  191.5 281.6 192.3 282.0 ;
      RECT  190.3 279.8 191.1 280.0 ;
      RECT  193.3 280.4 194.1 284.6 ;
      RECT  189.1 283.8 190.7 284.6 ;
      RECT  191.5 280.8 192.5 281.6 ;
      RECT  186.5 286.8 194.1 287.6 ;
      RECT  186.5 285.2 187.3 286.8 ;
      RECT  189.1 285.2 190.1 286.0 ;
      RECT  189.1 284.6 189.9 285.2 ;
      RECT  191.5 282.8 192.3 285.2 ;
      RECT  191.1 282.0 192.3 282.8 ;
      RECT  186.5 279.0 194.1 279.8 ;
      RECT  186.5 280.4 187.3 284.6 ;
      RECT  189.1 281.6 189.9 283.8 ;
      RECT  190.9 277.6 192.5 278.4 ;
      RECT  193.3 285.2 194.1 286.8 ;
      RECT  188.1 277.6 189.7 278.4 ;
      RECT  188.9 293.6 189.9 292.8 ;
      RECT  191.3 289.2 192.3 288.4 ;
      RECT  191.5 292.8 192.3 292.4 ;
      RECT  190.3 294.6 191.1 294.4 ;
      RECT  193.3 294.0 194.1 289.8 ;
      RECT  189.1 290.6 190.7 289.8 ;
      RECT  191.5 293.6 192.5 292.8 ;
      RECT  186.5 287.6 194.1 286.8 ;
      RECT  186.5 289.2 187.3 287.6 ;
      RECT  189.1 289.2 190.1 288.4 ;
      RECT  189.1 289.8 189.9 289.2 ;
      RECT  191.5 291.6 192.3 289.2 ;
      RECT  191.1 292.4 192.3 291.6 ;
      RECT  186.5 295.4 194.1 294.6 ;
      RECT  186.5 294.0 187.3 289.8 ;
      RECT  189.1 292.8 189.9 290.6 ;
      RECT  190.9 296.8 192.5 296.0 ;
      RECT  193.3 289.2 194.1 287.6 ;
      RECT  188.1 296.8 189.7 296.0 ;
      RECT  188.9 301.6 189.9 302.4 ;
      RECT  191.3 306.0 192.3 306.8 ;
      RECT  191.5 302.4 192.3 302.8 ;
      RECT  190.3 300.6 191.1 300.8 ;
      RECT  193.3 301.2 194.1 305.4 ;
      RECT  189.1 304.6 190.7 305.4 ;
      RECT  191.5 301.6 192.5 302.4 ;
      RECT  186.5 307.6 194.1 308.4 ;
      RECT  186.5 306.0 187.3 307.6 ;
      RECT  189.1 306.0 190.1 306.8 ;
      RECT  189.1 305.4 189.9 306.0 ;
      RECT  191.5 303.6 192.3 306.0 ;
      RECT  191.1 302.8 192.3 303.6 ;
      RECT  186.5 299.8 194.1 300.6 ;
      RECT  186.5 301.2 187.3 305.4 ;
      RECT  189.1 302.4 189.9 304.6 ;
      RECT  190.9 298.4 192.5 299.2 ;
      RECT  193.3 306.0 194.1 307.6 ;
      RECT  188.1 298.4 189.7 299.2 ;
      RECT  188.9 314.4 189.9 313.6 ;
      RECT  191.3 310.0 192.3 309.2 ;
      RECT  191.5 313.6 192.3 313.2 ;
      RECT  190.3 315.4 191.1 315.2 ;
      RECT  193.3 314.8 194.1 310.6 ;
      RECT  189.1 311.4 190.7 310.6 ;
      RECT  191.5 314.4 192.5 313.6 ;
      RECT  186.5 308.4 194.1 307.6 ;
      RECT  186.5 310.0 187.3 308.4 ;
      RECT  189.1 310.0 190.1 309.2 ;
      RECT  189.1 310.6 189.9 310.0 ;
      RECT  191.5 312.4 192.3 310.0 ;
      RECT  191.1 313.2 192.3 312.4 ;
      RECT  186.5 316.2 194.1 315.4 ;
      RECT  186.5 314.8 187.3 310.6 ;
      RECT  189.1 313.6 189.9 311.4 ;
      RECT  190.9 317.6 192.5 316.8 ;
      RECT  193.3 310.0 194.1 308.4 ;
      RECT  188.1 317.6 189.7 316.8 ;
      RECT  188.9 322.4 189.9 323.2 ;
      RECT  191.3 326.8 192.3 327.6 ;
      RECT  191.5 323.2 192.3 323.6 ;
      RECT  190.3 321.4 191.1 321.6 ;
      RECT  193.3 322.0 194.1 326.2 ;
      RECT  189.1 325.4 190.7 326.2 ;
      RECT  191.5 322.4 192.5 323.2 ;
      RECT  186.5 328.4 194.1 329.2 ;
      RECT  186.5 326.8 187.3 328.4 ;
      RECT  189.1 326.8 190.1 327.6 ;
      RECT  189.1 326.2 189.9 326.8 ;
      RECT  191.5 324.4 192.3 326.8 ;
      RECT  191.1 323.6 192.3 324.4 ;
      RECT  186.5 320.6 194.1 321.4 ;
      RECT  186.5 322.0 187.3 326.2 ;
      RECT  189.1 323.2 189.9 325.4 ;
      RECT  190.9 319.2 192.5 320.0 ;
      RECT  193.3 326.8 194.1 328.4 ;
      RECT  188.1 319.2 189.7 320.0 ;
      RECT  188.9 335.2 189.9 334.4 ;
      RECT  191.3 330.8 192.3 330.0 ;
      RECT  191.5 334.4 192.3 334.0 ;
      RECT  190.3 336.2 191.1 336.0 ;
      RECT  193.3 335.6 194.1 331.4 ;
      RECT  189.1 332.2 190.7 331.4 ;
      RECT  191.5 335.2 192.5 334.4 ;
      RECT  186.5 329.2 194.1 328.4 ;
      RECT  186.5 330.8 187.3 329.2 ;
      RECT  189.1 330.8 190.1 330.0 ;
      RECT  189.1 331.4 189.9 330.8 ;
      RECT  191.5 333.2 192.3 330.8 ;
      RECT  191.1 334.0 192.3 333.2 ;
      RECT  186.5 337.0 194.1 336.2 ;
      RECT  186.5 335.6 187.3 331.4 ;
      RECT  189.1 334.4 189.9 332.2 ;
      RECT  190.9 338.4 192.5 337.6 ;
      RECT  193.3 330.8 194.1 329.2 ;
      RECT  188.1 338.4 189.7 337.6 ;
      RECT  188.9 343.2 189.9 344.0 ;
      RECT  191.3 347.6 192.3 348.4 ;
      RECT  191.5 344.0 192.3 344.4 ;
      RECT  190.3 342.2 191.1 342.4 ;
      RECT  193.3 342.8 194.1 347.0 ;
      RECT  189.1 346.2 190.7 347.0 ;
      RECT  191.5 343.2 192.5 344.0 ;
      RECT  186.5 349.2 194.1 350.0 ;
      RECT  186.5 347.6 187.3 349.2 ;
      RECT  189.1 347.6 190.1 348.4 ;
      RECT  189.1 347.0 189.9 347.6 ;
      RECT  191.5 345.2 192.3 347.6 ;
      RECT  191.1 344.4 192.3 345.2 ;
      RECT  186.5 341.4 194.1 342.2 ;
      RECT  186.5 342.8 187.3 347.0 ;
      RECT  189.1 344.0 189.9 346.2 ;
      RECT  190.9 340.0 192.5 340.8 ;
      RECT  193.3 347.6 194.1 349.2 ;
      RECT  188.1 340.0 189.7 340.8 ;
      RECT  188.9 356.0 189.9 355.2 ;
      RECT  191.3 351.6 192.3 350.8 ;
      RECT  191.5 355.2 192.3 354.8 ;
      RECT  190.3 357.0 191.1 356.8 ;
      RECT  193.3 356.4 194.1 352.2 ;
      RECT  189.1 353.0 190.7 352.2 ;
      RECT  191.5 356.0 192.5 355.2 ;
      RECT  186.5 350.0 194.1 349.2 ;
      RECT  186.5 351.6 187.3 350.0 ;
      RECT  189.1 351.6 190.1 350.8 ;
      RECT  189.1 352.2 189.9 351.6 ;
      RECT  191.5 354.0 192.3 351.6 ;
      RECT  191.1 354.8 192.3 354.0 ;
      RECT  186.5 357.8 194.1 357.0 ;
      RECT  186.5 356.4 187.3 352.2 ;
      RECT  189.1 355.2 189.9 353.0 ;
      RECT  190.9 359.2 192.5 358.4 ;
      RECT  193.3 351.6 194.1 350.0 ;
      RECT  188.1 359.2 189.7 358.4 ;
      RECT  195.7 197.6 196.7 198.4 ;
      RECT  198.1 202.0 199.1 202.8 ;
      RECT  198.3 198.4 199.1 198.8 ;
      RECT  197.1 196.6 197.9 196.8 ;
      RECT  200.1 197.2 200.9 201.4 ;
      RECT  195.9 200.6 197.5 201.4 ;
      RECT  198.3 197.6 199.3 198.4 ;
      RECT  193.3 203.6 200.9 204.4 ;
      RECT  193.3 202.0 194.1 203.6 ;
      RECT  195.9 202.0 196.9 202.8 ;
      RECT  195.9 201.4 196.7 202.0 ;
      RECT  198.3 199.6 199.1 202.0 ;
      RECT  197.9 198.8 199.1 199.6 ;
      RECT  193.3 195.8 200.9 196.6 ;
      RECT  193.3 197.2 194.1 201.4 ;
      RECT  195.9 198.4 196.7 200.6 ;
      RECT  197.7 194.4 199.3 195.2 ;
      RECT  200.1 202.0 200.9 203.6 ;
      RECT  194.9 194.4 196.5 195.2 ;
      RECT  195.7 210.4 196.7 209.6 ;
      RECT  198.1 206.0 199.1 205.2 ;
      RECT  198.3 209.6 199.1 209.2 ;
      RECT  197.1 211.4 197.9 211.2 ;
      RECT  200.1 210.8 200.9 206.6 ;
      RECT  195.9 207.4 197.5 206.6 ;
      RECT  198.3 210.4 199.3 209.6 ;
      RECT  193.3 204.4 200.9 203.6 ;
      RECT  193.3 206.0 194.1 204.4 ;
      RECT  195.9 206.0 196.9 205.2 ;
      RECT  195.9 206.6 196.7 206.0 ;
      RECT  198.3 208.4 199.1 206.0 ;
      RECT  197.9 209.2 199.1 208.4 ;
      RECT  193.3 212.2 200.9 211.4 ;
      RECT  193.3 210.8 194.1 206.6 ;
      RECT  195.9 209.6 196.7 207.4 ;
      RECT  197.7 213.6 199.3 212.8 ;
      RECT  200.1 206.0 200.9 204.4 ;
      RECT  194.9 213.6 196.5 212.8 ;
      RECT  195.7 218.4 196.7 219.2 ;
      RECT  198.1 222.8 199.1 223.6 ;
      RECT  198.3 219.2 199.1 219.6 ;
      RECT  197.1 217.4 197.9 217.6 ;
      RECT  200.1 218.0 200.9 222.2 ;
      RECT  195.9 221.4 197.5 222.2 ;
      RECT  198.3 218.4 199.3 219.2 ;
      RECT  193.3 224.4 200.9 225.2 ;
      RECT  193.3 222.8 194.1 224.4 ;
      RECT  195.9 222.8 196.9 223.6 ;
      RECT  195.9 222.2 196.7 222.8 ;
      RECT  198.3 220.4 199.1 222.8 ;
      RECT  197.9 219.6 199.1 220.4 ;
      RECT  193.3 216.6 200.9 217.4 ;
      RECT  193.3 218.0 194.1 222.2 ;
      RECT  195.9 219.2 196.7 221.4 ;
      RECT  197.7 215.2 199.3 216.0 ;
      RECT  200.1 222.8 200.9 224.4 ;
      RECT  194.9 215.2 196.5 216.0 ;
      RECT  195.7 231.2 196.7 230.4 ;
      RECT  198.1 226.8 199.1 226.0 ;
      RECT  198.3 230.4 199.1 230.0 ;
      RECT  197.1 232.2 197.9 232.0 ;
      RECT  200.1 231.6 200.9 227.4 ;
      RECT  195.9 228.2 197.5 227.4 ;
      RECT  198.3 231.2 199.3 230.4 ;
      RECT  193.3 225.2 200.9 224.4 ;
      RECT  193.3 226.8 194.1 225.2 ;
      RECT  195.9 226.8 196.9 226.0 ;
      RECT  195.9 227.4 196.7 226.8 ;
      RECT  198.3 229.2 199.1 226.8 ;
      RECT  197.9 230.0 199.1 229.2 ;
      RECT  193.3 233.0 200.9 232.2 ;
      RECT  193.3 231.6 194.1 227.4 ;
      RECT  195.9 230.4 196.7 228.2 ;
      RECT  197.7 234.4 199.3 233.6 ;
      RECT  200.1 226.8 200.9 225.2 ;
      RECT  194.9 234.4 196.5 233.6 ;
      RECT  195.7 239.2 196.7 240.0 ;
      RECT  198.1 243.6 199.1 244.4 ;
      RECT  198.3 240.0 199.1 240.4 ;
      RECT  197.1 238.2 197.9 238.4 ;
      RECT  200.1 238.8 200.9 243.0 ;
      RECT  195.9 242.2 197.5 243.0 ;
      RECT  198.3 239.2 199.3 240.0 ;
      RECT  193.3 245.2 200.9 246.0 ;
      RECT  193.3 243.6 194.1 245.2 ;
      RECT  195.9 243.6 196.9 244.4 ;
      RECT  195.9 243.0 196.7 243.6 ;
      RECT  198.3 241.2 199.1 243.6 ;
      RECT  197.9 240.4 199.1 241.2 ;
      RECT  193.3 237.4 200.9 238.2 ;
      RECT  193.3 238.8 194.1 243.0 ;
      RECT  195.9 240.0 196.7 242.2 ;
      RECT  197.7 236.0 199.3 236.8 ;
      RECT  200.1 243.6 200.9 245.2 ;
      RECT  194.9 236.0 196.5 236.8 ;
      RECT  195.7 252.0 196.7 251.2 ;
      RECT  198.1 247.6 199.1 246.8 ;
      RECT  198.3 251.2 199.1 250.8 ;
      RECT  197.1 253.0 197.9 252.8 ;
      RECT  200.1 252.4 200.9 248.2 ;
      RECT  195.9 249.0 197.5 248.2 ;
      RECT  198.3 252.0 199.3 251.2 ;
      RECT  193.3 246.0 200.9 245.2 ;
      RECT  193.3 247.6 194.1 246.0 ;
      RECT  195.9 247.6 196.9 246.8 ;
      RECT  195.9 248.2 196.7 247.6 ;
      RECT  198.3 250.0 199.1 247.6 ;
      RECT  197.9 250.8 199.1 250.0 ;
      RECT  193.3 253.8 200.9 253.0 ;
      RECT  193.3 252.4 194.1 248.2 ;
      RECT  195.9 251.2 196.7 249.0 ;
      RECT  197.7 255.2 199.3 254.4 ;
      RECT  200.1 247.6 200.9 246.0 ;
      RECT  194.9 255.2 196.5 254.4 ;
      RECT  195.7 260.0 196.7 260.8 ;
      RECT  198.1 264.4 199.1 265.2 ;
      RECT  198.3 260.8 199.1 261.2 ;
      RECT  197.1 259.0 197.9 259.2 ;
      RECT  200.1 259.6 200.9 263.8 ;
      RECT  195.9 263.0 197.5 263.8 ;
      RECT  198.3 260.0 199.3 260.8 ;
      RECT  193.3 266.0 200.9 266.8 ;
      RECT  193.3 264.4 194.1 266.0 ;
      RECT  195.9 264.4 196.9 265.2 ;
      RECT  195.9 263.8 196.7 264.4 ;
      RECT  198.3 262.0 199.1 264.4 ;
      RECT  197.9 261.2 199.1 262.0 ;
      RECT  193.3 258.2 200.9 259.0 ;
      RECT  193.3 259.6 194.1 263.8 ;
      RECT  195.9 260.8 196.7 263.0 ;
      RECT  197.7 256.8 199.3 257.6 ;
      RECT  200.1 264.4 200.9 266.0 ;
      RECT  194.9 256.8 196.5 257.6 ;
      RECT  195.7 272.8 196.7 272.0 ;
      RECT  198.1 268.4 199.1 267.6 ;
      RECT  198.3 272.0 199.1 271.6 ;
      RECT  197.1 273.8 197.9 273.6 ;
      RECT  200.1 273.2 200.9 269.0 ;
      RECT  195.9 269.8 197.5 269.0 ;
      RECT  198.3 272.8 199.3 272.0 ;
      RECT  193.3 266.8 200.9 266.0 ;
      RECT  193.3 268.4 194.1 266.8 ;
      RECT  195.9 268.4 196.9 267.6 ;
      RECT  195.9 269.0 196.7 268.4 ;
      RECT  198.3 270.8 199.1 268.4 ;
      RECT  197.9 271.6 199.1 270.8 ;
      RECT  193.3 274.6 200.9 273.8 ;
      RECT  193.3 273.2 194.1 269.0 ;
      RECT  195.9 272.0 196.7 269.8 ;
      RECT  197.7 276.0 199.3 275.2 ;
      RECT  200.1 268.4 200.9 266.8 ;
      RECT  194.9 276.0 196.5 275.2 ;
      RECT  195.7 280.8 196.7 281.6 ;
      RECT  198.1 285.2 199.1 286.0 ;
      RECT  198.3 281.6 199.1 282.0 ;
      RECT  197.1 279.8 197.9 280.0 ;
      RECT  200.1 280.4 200.9 284.6 ;
      RECT  195.9 283.8 197.5 284.6 ;
      RECT  198.3 280.8 199.3 281.6 ;
      RECT  193.3 286.8 200.9 287.6 ;
      RECT  193.3 285.2 194.1 286.8 ;
      RECT  195.9 285.2 196.9 286.0 ;
      RECT  195.9 284.6 196.7 285.2 ;
      RECT  198.3 282.8 199.1 285.2 ;
      RECT  197.9 282.0 199.1 282.8 ;
      RECT  193.3 279.0 200.9 279.8 ;
      RECT  193.3 280.4 194.1 284.6 ;
      RECT  195.9 281.6 196.7 283.8 ;
      RECT  197.7 277.6 199.3 278.4 ;
      RECT  200.1 285.2 200.9 286.8 ;
      RECT  194.9 277.6 196.5 278.4 ;
      RECT  195.7 293.6 196.7 292.8 ;
      RECT  198.1 289.2 199.1 288.4 ;
      RECT  198.3 292.8 199.1 292.4 ;
      RECT  197.1 294.6 197.9 294.4 ;
      RECT  200.1 294.0 200.9 289.8 ;
      RECT  195.9 290.6 197.5 289.8 ;
      RECT  198.3 293.6 199.3 292.8 ;
      RECT  193.3 287.6 200.9 286.8 ;
      RECT  193.3 289.2 194.1 287.6 ;
      RECT  195.9 289.2 196.9 288.4 ;
      RECT  195.9 289.8 196.7 289.2 ;
      RECT  198.3 291.6 199.1 289.2 ;
      RECT  197.9 292.4 199.1 291.6 ;
      RECT  193.3 295.4 200.9 294.6 ;
      RECT  193.3 294.0 194.1 289.8 ;
      RECT  195.9 292.8 196.7 290.6 ;
      RECT  197.7 296.8 199.3 296.0 ;
      RECT  200.1 289.2 200.9 287.6 ;
      RECT  194.9 296.8 196.5 296.0 ;
      RECT  195.7 301.6 196.7 302.4 ;
      RECT  198.1 306.0 199.1 306.8 ;
      RECT  198.3 302.4 199.1 302.8 ;
      RECT  197.1 300.6 197.9 300.8 ;
      RECT  200.1 301.2 200.9 305.4 ;
      RECT  195.9 304.6 197.5 305.4 ;
      RECT  198.3 301.6 199.3 302.4 ;
      RECT  193.3 307.6 200.9 308.4 ;
      RECT  193.3 306.0 194.1 307.6 ;
      RECT  195.9 306.0 196.9 306.8 ;
      RECT  195.9 305.4 196.7 306.0 ;
      RECT  198.3 303.6 199.1 306.0 ;
      RECT  197.9 302.8 199.1 303.6 ;
      RECT  193.3 299.8 200.9 300.6 ;
      RECT  193.3 301.2 194.1 305.4 ;
      RECT  195.9 302.4 196.7 304.6 ;
      RECT  197.7 298.4 199.3 299.2 ;
      RECT  200.1 306.0 200.9 307.6 ;
      RECT  194.9 298.4 196.5 299.2 ;
      RECT  195.7 314.4 196.7 313.6 ;
      RECT  198.1 310.0 199.1 309.2 ;
      RECT  198.3 313.6 199.1 313.2 ;
      RECT  197.1 315.4 197.9 315.2 ;
      RECT  200.1 314.8 200.9 310.6 ;
      RECT  195.9 311.4 197.5 310.6 ;
      RECT  198.3 314.4 199.3 313.6 ;
      RECT  193.3 308.4 200.9 307.6 ;
      RECT  193.3 310.0 194.1 308.4 ;
      RECT  195.9 310.0 196.9 309.2 ;
      RECT  195.9 310.6 196.7 310.0 ;
      RECT  198.3 312.4 199.1 310.0 ;
      RECT  197.9 313.2 199.1 312.4 ;
      RECT  193.3 316.2 200.9 315.4 ;
      RECT  193.3 314.8 194.1 310.6 ;
      RECT  195.9 313.6 196.7 311.4 ;
      RECT  197.7 317.6 199.3 316.8 ;
      RECT  200.1 310.0 200.9 308.4 ;
      RECT  194.9 317.6 196.5 316.8 ;
      RECT  195.7 322.4 196.7 323.2 ;
      RECT  198.1 326.8 199.1 327.6 ;
      RECT  198.3 323.2 199.1 323.6 ;
      RECT  197.1 321.4 197.9 321.6 ;
      RECT  200.1 322.0 200.9 326.2 ;
      RECT  195.9 325.4 197.5 326.2 ;
      RECT  198.3 322.4 199.3 323.2 ;
      RECT  193.3 328.4 200.9 329.2 ;
      RECT  193.3 326.8 194.1 328.4 ;
      RECT  195.9 326.8 196.9 327.6 ;
      RECT  195.9 326.2 196.7 326.8 ;
      RECT  198.3 324.4 199.1 326.8 ;
      RECT  197.9 323.6 199.1 324.4 ;
      RECT  193.3 320.6 200.9 321.4 ;
      RECT  193.3 322.0 194.1 326.2 ;
      RECT  195.9 323.2 196.7 325.4 ;
      RECT  197.7 319.2 199.3 320.0 ;
      RECT  200.1 326.8 200.9 328.4 ;
      RECT  194.9 319.2 196.5 320.0 ;
      RECT  195.7 335.2 196.7 334.4 ;
      RECT  198.1 330.8 199.1 330.0 ;
      RECT  198.3 334.4 199.1 334.0 ;
      RECT  197.1 336.2 197.9 336.0 ;
      RECT  200.1 335.6 200.9 331.4 ;
      RECT  195.9 332.2 197.5 331.4 ;
      RECT  198.3 335.2 199.3 334.4 ;
      RECT  193.3 329.2 200.9 328.4 ;
      RECT  193.3 330.8 194.1 329.2 ;
      RECT  195.9 330.8 196.9 330.0 ;
      RECT  195.9 331.4 196.7 330.8 ;
      RECT  198.3 333.2 199.1 330.8 ;
      RECT  197.9 334.0 199.1 333.2 ;
      RECT  193.3 337.0 200.9 336.2 ;
      RECT  193.3 335.6 194.1 331.4 ;
      RECT  195.9 334.4 196.7 332.2 ;
      RECT  197.7 338.4 199.3 337.6 ;
      RECT  200.1 330.8 200.9 329.2 ;
      RECT  194.9 338.4 196.5 337.6 ;
      RECT  195.7 343.2 196.7 344.0 ;
      RECT  198.1 347.6 199.1 348.4 ;
      RECT  198.3 344.0 199.1 344.4 ;
      RECT  197.1 342.2 197.9 342.4 ;
      RECT  200.1 342.8 200.9 347.0 ;
      RECT  195.9 346.2 197.5 347.0 ;
      RECT  198.3 343.2 199.3 344.0 ;
      RECT  193.3 349.2 200.9 350.0 ;
      RECT  193.3 347.6 194.1 349.2 ;
      RECT  195.9 347.6 196.9 348.4 ;
      RECT  195.9 347.0 196.7 347.6 ;
      RECT  198.3 345.2 199.1 347.6 ;
      RECT  197.9 344.4 199.1 345.2 ;
      RECT  193.3 341.4 200.9 342.2 ;
      RECT  193.3 342.8 194.1 347.0 ;
      RECT  195.9 344.0 196.7 346.2 ;
      RECT  197.7 340.0 199.3 340.8 ;
      RECT  200.1 347.6 200.9 349.2 ;
      RECT  194.9 340.0 196.5 340.8 ;
      RECT  195.7 356.0 196.7 355.2 ;
      RECT  198.1 351.6 199.1 350.8 ;
      RECT  198.3 355.2 199.1 354.8 ;
      RECT  197.1 357.0 197.9 356.8 ;
      RECT  200.1 356.4 200.9 352.2 ;
      RECT  195.9 353.0 197.5 352.2 ;
      RECT  198.3 356.0 199.3 355.2 ;
      RECT  193.3 350.0 200.9 349.2 ;
      RECT  193.3 351.6 194.1 350.0 ;
      RECT  195.9 351.6 196.9 350.8 ;
      RECT  195.9 352.2 196.7 351.6 ;
      RECT  198.3 354.0 199.1 351.6 ;
      RECT  197.9 354.8 199.1 354.0 ;
      RECT  193.3 357.8 200.9 357.0 ;
      RECT  193.3 356.4 194.1 352.2 ;
      RECT  195.9 355.2 196.7 353.0 ;
      RECT  197.7 359.2 199.3 358.4 ;
      RECT  200.1 351.6 200.9 350.0 ;
      RECT  194.9 359.2 196.5 358.4 ;
      RECT  186.9 195.8 200.5 196.6 ;
      RECT  186.9 211.4 200.5 212.2 ;
      RECT  186.9 216.6 200.5 217.4 ;
      RECT  186.9 232.2 200.5 233.0 ;
      RECT  186.9 237.4 200.5 238.2 ;
      RECT  186.9 253.0 200.5 253.8 ;
      RECT  186.9 258.2 200.5 259.0 ;
      RECT  186.9 273.8 200.5 274.6 ;
      RECT  186.9 279.0 200.5 279.8 ;
      RECT  186.9 294.6 200.5 295.4 ;
      RECT  186.9 299.8 200.5 300.6 ;
      RECT  186.9 315.4 200.5 316.2 ;
      RECT  186.9 320.6 200.5 321.4 ;
      RECT  186.9 336.2 200.5 337.0 ;
      RECT  186.9 341.4 200.5 342.2 ;
      RECT  186.9 357.0 200.5 357.8 ;
      RECT  182.1 176.8 183.1 177.6 ;
      RECT  184.5 181.2 185.5 182.0 ;
      RECT  184.7 177.6 185.5 178.0 ;
      RECT  183.5 175.8 184.3 176.0 ;
      RECT  186.5 176.4 187.3 180.6 ;
      RECT  182.3 179.8 183.9 180.6 ;
      RECT  184.7 176.8 185.7 177.6 ;
      RECT  182.1 173.6 182.9 174.4 ;
      RECT  179.7 182.8 187.3 183.6 ;
      RECT  179.7 181.2 180.5 182.8 ;
      RECT  182.3 181.2 183.3 182.0 ;
      RECT  182.3 180.6 183.1 181.2 ;
      RECT  184.7 178.8 185.5 181.2 ;
      RECT  184.3 178.0 185.5 178.8 ;
      RECT  179.7 175.0 187.3 175.8 ;
      RECT  184.9 173.6 185.7 174.4 ;
      RECT  179.7 176.4 180.5 180.6 ;
      RECT  182.3 177.6 183.1 179.8 ;
      RECT  186.5 181.2 187.3 182.8 ;
      RECT  182.1 189.6 183.1 188.8 ;
      RECT  184.5 185.2 185.5 184.4 ;
      RECT  184.7 188.8 185.5 188.4 ;
      RECT  183.5 190.6 184.3 190.4 ;
      RECT  186.5 190.0 187.3 185.8 ;
      RECT  182.3 186.6 183.9 185.8 ;
      RECT  184.5 184.4 185.3 183.6 ;
      RECT  184.7 189.6 185.7 188.8 ;
      RECT  179.7 183.6 187.3 182.8 ;
      RECT  179.7 185.2 180.5 183.6 ;
      RECT  182.3 185.2 183.3 184.4 ;
      RECT  182.3 185.8 183.1 185.2 ;
      RECT  184.7 187.6 185.5 185.2 ;
      RECT  184.3 188.4 185.5 187.6 ;
      RECT  179.7 191.4 187.3 190.6 ;
      RECT  179.7 190.0 180.5 185.8 ;
      RECT  182.3 188.8 183.1 186.6 ;
      RECT  184.1 192.8 185.7 192.0 ;
      RECT  186.5 185.2 187.3 183.6 ;
      RECT  181.3 192.8 182.9 192.0 ;
      RECT  182.1 197.6 183.1 198.4 ;
      RECT  184.5 202.0 185.5 202.8 ;
      RECT  184.7 198.4 185.5 198.8 ;
      RECT  183.5 196.6 184.3 196.8 ;
      RECT  186.5 197.2 187.3 201.4 ;
      RECT  182.3 200.6 183.9 201.4 ;
      RECT  184.5 202.8 185.3 203.6 ;
      RECT  184.7 197.6 185.7 198.4 ;
      RECT  179.7 203.6 187.3 204.4 ;
      RECT  179.7 202.0 180.5 203.6 ;
      RECT  182.3 202.0 183.3 202.8 ;
      RECT  182.3 201.4 183.1 202.0 ;
      RECT  184.7 199.6 185.5 202.0 ;
      RECT  184.3 198.8 185.5 199.6 ;
      RECT  179.7 195.8 187.3 196.6 ;
      RECT  179.7 197.2 180.5 201.4 ;
      RECT  182.3 198.4 183.1 200.6 ;
      RECT  184.1 194.4 185.7 195.2 ;
      RECT  186.5 202.0 187.3 203.6 ;
      RECT  181.3 194.4 182.9 195.2 ;
      RECT  182.1 210.4 183.1 209.6 ;
      RECT  184.5 206.0 185.5 205.2 ;
      RECT  184.7 209.6 185.5 209.2 ;
      RECT  183.5 211.4 184.3 211.2 ;
      RECT  186.5 210.8 187.3 206.6 ;
      RECT  182.3 207.4 183.9 206.6 ;
      RECT  184.5 205.2 185.3 204.4 ;
      RECT  184.7 210.4 185.7 209.6 ;
      RECT  179.7 204.4 187.3 203.6 ;
      RECT  179.7 206.0 180.5 204.4 ;
      RECT  182.3 206.0 183.3 205.2 ;
      RECT  182.3 206.6 183.1 206.0 ;
      RECT  184.7 208.4 185.5 206.0 ;
      RECT  184.3 209.2 185.5 208.4 ;
      RECT  179.7 212.2 187.3 211.4 ;
      RECT  179.7 210.8 180.5 206.6 ;
      RECT  182.3 209.6 183.1 207.4 ;
      RECT  184.1 213.6 185.7 212.8 ;
      RECT  186.5 206.0 187.3 204.4 ;
      RECT  181.3 213.6 182.9 212.8 ;
      RECT  182.1 218.4 183.1 219.2 ;
      RECT  184.5 222.8 185.5 223.6 ;
      RECT  184.7 219.2 185.5 219.6 ;
      RECT  183.5 217.4 184.3 217.6 ;
      RECT  186.5 218.0 187.3 222.2 ;
      RECT  182.3 221.4 183.9 222.2 ;
      RECT  184.5 223.6 185.3 224.4 ;
      RECT  184.7 218.4 185.7 219.2 ;
      RECT  179.7 224.4 187.3 225.2 ;
      RECT  179.7 222.8 180.5 224.4 ;
      RECT  182.3 222.8 183.3 223.6 ;
      RECT  182.3 222.2 183.1 222.8 ;
      RECT  184.7 220.4 185.5 222.8 ;
      RECT  184.3 219.6 185.5 220.4 ;
      RECT  179.7 216.6 187.3 217.4 ;
      RECT  179.7 218.0 180.5 222.2 ;
      RECT  182.3 219.2 183.1 221.4 ;
      RECT  184.1 215.2 185.7 216.0 ;
      RECT  186.5 222.8 187.3 224.4 ;
      RECT  181.3 215.2 182.9 216.0 ;
      RECT  182.1 231.2 183.1 230.4 ;
      RECT  184.5 226.8 185.5 226.0 ;
      RECT  184.7 230.4 185.5 230.0 ;
      RECT  183.5 232.2 184.3 232.0 ;
      RECT  186.5 231.6 187.3 227.4 ;
      RECT  182.3 228.2 183.9 227.4 ;
      RECT  184.5 226.0 185.3 225.2 ;
      RECT  184.7 231.2 185.7 230.4 ;
      RECT  179.7 225.2 187.3 224.4 ;
      RECT  179.7 226.8 180.5 225.2 ;
      RECT  182.3 226.8 183.3 226.0 ;
      RECT  182.3 227.4 183.1 226.8 ;
      RECT  184.7 229.2 185.5 226.8 ;
      RECT  184.3 230.0 185.5 229.2 ;
      RECT  179.7 233.0 187.3 232.2 ;
      RECT  179.7 231.6 180.5 227.4 ;
      RECT  182.3 230.4 183.1 228.2 ;
      RECT  184.1 234.4 185.7 233.6 ;
      RECT  186.5 226.8 187.3 225.2 ;
      RECT  181.3 234.4 182.9 233.6 ;
      RECT  182.1 239.2 183.1 240.0 ;
      RECT  184.5 243.6 185.5 244.4 ;
      RECT  184.7 240.0 185.5 240.4 ;
      RECT  183.5 238.2 184.3 238.4 ;
      RECT  186.5 238.8 187.3 243.0 ;
      RECT  182.3 242.2 183.9 243.0 ;
      RECT  184.5 244.4 185.3 245.2 ;
      RECT  184.7 239.2 185.7 240.0 ;
      RECT  179.7 245.2 187.3 246.0 ;
      RECT  179.7 243.6 180.5 245.2 ;
      RECT  182.3 243.6 183.3 244.4 ;
      RECT  182.3 243.0 183.1 243.6 ;
      RECT  184.7 241.2 185.5 243.6 ;
      RECT  184.3 240.4 185.5 241.2 ;
      RECT  179.7 237.4 187.3 238.2 ;
      RECT  179.7 238.8 180.5 243.0 ;
      RECT  182.3 240.0 183.1 242.2 ;
      RECT  184.1 236.0 185.7 236.8 ;
      RECT  186.5 243.6 187.3 245.2 ;
      RECT  181.3 236.0 182.9 236.8 ;
      RECT  182.1 252.0 183.1 251.2 ;
      RECT  184.5 247.6 185.5 246.8 ;
      RECT  184.7 251.2 185.5 250.8 ;
      RECT  183.5 253.0 184.3 252.8 ;
      RECT  186.5 252.4 187.3 248.2 ;
      RECT  182.3 249.0 183.9 248.2 ;
      RECT  184.5 246.8 185.3 246.0 ;
      RECT  184.7 252.0 185.7 251.2 ;
      RECT  179.7 246.0 187.3 245.2 ;
      RECT  179.7 247.6 180.5 246.0 ;
      RECT  182.3 247.6 183.3 246.8 ;
      RECT  182.3 248.2 183.1 247.6 ;
      RECT  184.7 250.0 185.5 247.6 ;
      RECT  184.3 250.8 185.5 250.0 ;
      RECT  179.7 253.8 187.3 253.0 ;
      RECT  179.7 252.4 180.5 248.2 ;
      RECT  182.3 251.2 183.1 249.0 ;
      RECT  184.1 255.2 185.7 254.4 ;
      RECT  186.5 247.6 187.3 246.0 ;
      RECT  181.3 255.2 182.9 254.4 ;
      RECT  182.1 260.0 183.1 260.8 ;
      RECT  184.5 264.4 185.5 265.2 ;
      RECT  184.7 260.8 185.5 261.2 ;
      RECT  183.5 259.0 184.3 259.2 ;
      RECT  186.5 259.6 187.3 263.8 ;
      RECT  182.3 263.0 183.9 263.8 ;
      RECT  184.5 265.2 185.3 266.0 ;
      RECT  184.7 260.0 185.7 260.8 ;
      RECT  179.7 266.0 187.3 266.8 ;
      RECT  179.7 264.4 180.5 266.0 ;
      RECT  182.3 264.4 183.3 265.2 ;
      RECT  182.3 263.8 183.1 264.4 ;
      RECT  184.7 262.0 185.5 264.4 ;
      RECT  184.3 261.2 185.5 262.0 ;
      RECT  179.7 258.2 187.3 259.0 ;
      RECT  179.7 259.6 180.5 263.8 ;
      RECT  182.3 260.8 183.1 263.0 ;
      RECT  184.1 256.8 185.7 257.6 ;
      RECT  186.5 264.4 187.3 266.0 ;
      RECT  181.3 256.8 182.9 257.6 ;
      RECT  182.1 272.8 183.1 272.0 ;
      RECT  184.5 268.4 185.5 267.6 ;
      RECT  184.7 272.0 185.5 271.6 ;
      RECT  183.5 273.8 184.3 273.6 ;
      RECT  186.5 273.2 187.3 269.0 ;
      RECT  182.3 269.8 183.9 269.0 ;
      RECT  184.5 267.6 185.3 266.8 ;
      RECT  184.7 272.8 185.7 272.0 ;
      RECT  179.7 266.8 187.3 266.0 ;
      RECT  179.7 268.4 180.5 266.8 ;
      RECT  182.3 268.4 183.3 267.6 ;
      RECT  182.3 269.0 183.1 268.4 ;
      RECT  184.7 270.8 185.5 268.4 ;
      RECT  184.3 271.6 185.5 270.8 ;
      RECT  179.7 274.6 187.3 273.8 ;
      RECT  179.7 273.2 180.5 269.0 ;
      RECT  182.3 272.0 183.1 269.8 ;
      RECT  184.1 276.0 185.7 275.2 ;
      RECT  186.5 268.4 187.3 266.8 ;
      RECT  181.3 276.0 182.9 275.2 ;
      RECT  182.1 280.8 183.1 281.6 ;
      RECT  184.5 285.2 185.5 286.0 ;
      RECT  184.7 281.6 185.5 282.0 ;
      RECT  183.5 279.8 184.3 280.0 ;
      RECT  186.5 280.4 187.3 284.6 ;
      RECT  182.3 283.8 183.9 284.6 ;
      RECT  184.5 286.0 185.3 286.8 ;
      RECT  184.7 280.8 185.7 281.6 ;
      RECT  179.7 286.8 187.3 287.6 ;
      RECT  179.7 285.2 180.5 286.8 ;
      RECT  182.3 285.2 183.3 286.0 ;
      RECT  182.3 284.6 183.1 285.2 ;
      RECT  184.7 282.8 185.5 285.2 ;
      RECT  184.3 282.0 185.5 282.8 ;
      RECT  179.7 279.0 187.3 279.8 ;
      RECT  179.7 280.4 180.5 284.6 ;
      RECT  182.3 281.6 183.1 283.8 ;
      RECT  184.1 277.6 185.7 278.4 ;
      RECT  186.5 285.2 187.3 286.8 ;
      RECT  181.3 277.6 182.9 278.4 ;
      RECT  182.1 293.6 183.1 292.8 ;
      RECT  184.5 289.2 185.5 288.4 ;
      RECT  184.7 292.8 185.5 292.4 ;
      RECT  183.5 294.6 184.3 294.4 ;
      RECT  186.5 294.0 187.3 289.8 ;
      RECT  182.3 290.6 183.9 289.8 ;
      RECT  184.5 288.4 185.3 287.6 ;
      RECT  184.7 293.6 185.7 292.8 ;
      RECT  179.7 287.6 187.3 286.8 ;
      RECT  179.7 289.2 180.5 287.6 ;
      RECT  182.3 289.2 183.3 288.4 ;
      RECT  182.3 289.8 183.1 289.2 ;
      RECT  184.7 291.6 185.5 289.2 ;
      RECT  184.3 292.4 185.5 291.6 ;
      RECT  179.7 295.4 187.3 294.6 ;
      RECT  179.7 294.0 180.5 289.8 ;
      RECT  182.3 292.8 183.1 290.6 ;
      RECT  184.1 296.8 185.7 296.0 ;
      RECT  186.5 289.2 187.3 287.6 ;
      RECT  181.3 296.8 182.9 296.0 ;
      RECT  182.1 301.6 183.1 302.4 ;
      RECT  184.5 306.0 185.5 306.8 ;
      RECT  184.7 302.4 185.5 302.8 ;
      RECT  183.5 300.6 184.3 300.8 ;
      RECT  186.5 301.2 187.3 305.4 ;
      RECT  182.3 304.6 183.9 305.4 ;
      RECT  184.5 306.8 185.3 307.6 ;
      RECT  184.7 301.6 185.7 302.4 ;
      RECT  179.7 307.6 187.3 308.4 ;
      RECT  179.7 306.0 180.5 307.6 ;
      RECT  182.3 306.0 183.3 306.8 ;
      RECT  182.3 305.4 183.1 306.0 ;
      RECT  184.7 303.6 185.5 306.0 ;
      RECT  184.3 302.8 185.5 303.6 ;
      RECT  179.7 299.8 187.3 300.6 ;
      RECT  179.7 301.2 180.5 305.4 ;
      RECT  182.3 302.4 183.1 304.6 ;
      RECT  184.1 298.4 185.7 299.2 ;
      RECT  186.5 306.0 187.3 307.6 ;
      RECT  181.3 298.4 182.9 299.2 ;
      RECT  182.1 314.4 183.1 313.6 ;
      RECT  184.5 310.0 185.5 309.2 ;
      RECT  184.7 313.6 185.5 313.2 ;
      RECT  183.5 315.4 184.3 315.2 ;
      RECT  186.5 314.8 187.3 310.6 ;
      RECT  182.3 311.4 183.9 310.6 ;
      RECT  184.5 309.2 185.3 308.4 ;
      RECT  184.7 314.4 185.7 313.6 ;
      RECT  179.7 308.4 187.3 307.6 ;
      RECT  179.7 310.0 180.5 308.4 ;
      RECT  182.3 310.0 183.3 309.2 ;
      RECT  182.3 310.6 183.1 310.0 ;
      RECT  184.7 312.4 185.5 310.0 ;
      RECT  184.3 313.2 185.5 312.4 ;
      RECT  179.7 316.2 187.3 315.4 ;
      RECT  179.7 314.8 180.5 310.6 ;
      RECT  182.3 313.6 183.1 311.4 ;
      RECT  184.1 317.6 185.7 316.8 ;
      RECT  186.5 310.0 187.3 308.4 ;
      RECT  181.3 317.6 182.9 316.8 ;
      RECT  182.1 322.4 183.1 323.2 ;
      RECT  184.5 326.8 185.5 327.6 ;
      RECT  184.7 323.2 185.5 323.6 ;
      RECT  183.5 321.4 184.3 321.6 ;
      RECT  186.5 322.0 187.3 326.2 ;
      RECT  182.3 325.4 183.9 326.2 ;
      RECT  184.5 327.6 185.3 328.4 ;
      RECT  184.7 322.4 185.7 323.2 ;
      RECT  179.7 328.4 187.3 329.2 ;
      RECT  179.7 326.8 180.5 328.4 ;
      RECT  182.3 326.8 183.3 327.6 ;
      RECT  182.3 326.2 183.1 326.8 ;
      RECT  184.7 324.4 185.5 326.8 ;
      RECT  184.3 323.6 185.5 324.4 ;
      RECT  179.7 320.6 187.3 321.4 ;
      RECT  179.7 322.0 180.5 326.2 ;
      RECT  182.3 323.2 183.1 325.4 ;
      RECT  184.1 319.2 185.7 320.0 ;
      RECT  186.5 326.8 187.3 328.4 ;
      RECT  181.3 319.2 182.9 320.0 ;
      RECT  182.1 335.2 183.1 334.4 ;
      RECT  184.5 330.8 185.5 330.0 ;
      RECT  184.7 334.4 185.5 334.0 ;
      RECT  183.5 336.2 184.3 336.0 ;
      RECT  186.5 335.6 187.3 331.4 ;
      RECT  182.3 332.2 183.9 331.4 ;
      RECT  184.5 330.0 185.3 329.2 ;
      RECT  184.7 335.2 185.7 334.4 ;
      RECT  179.7 329.2 187.3 328.4 ;
      RECT  179.7 330.8 180.5 329.2 ;
      RECT  182.3 330.8 183.3 330.0 ;
      RECT  182.3 331.4 183.1 330.8 ;
      RECT  184.7 333.2 185.5 330.8 ;
      RECT  184.3 334.0 185.5 333.2 ;
      RECT  179.7 337.0 187.3 336.2 ;
      RECT  179.7 335.6 180.5 331.4 ;
      RECT  182.3 334.4 183.1 332.2 ;
      RECT  184.1 338.4 185.7 337.6 ;
      RECT  186.5 330.8 187.3 329.2 ;
      RECT  181.3 338.4 182.9 337.6 ;
      RECT  182.1 343.2 183.1 344.0 ;
      RECT  184.5 347.6 185.5 348.4 ;
      RECT  184.7 344.0 185.5 344.4 ;
      RECT  183.5 342.2 184.3 342.4 ;
      RECT  186.5 342.8 187.3 347.0 ;
      RECT  182.3 346.2 183.9 347.0 ;
      RECT  184.5 348.4 185.3 349.2 ;
      RECT  184.7 343.2 185.7 344.0 ;
      RECT  179.7 349.2 187.3 350.0 ;
      RECT  179.7 347.6 180.5 349.2 ;
      RECT  182.3 347.6 183.3 348.4 ;
      RECT  182.3 347.0 183.1 347.6 ;
      RECT  184.7 345.2 185.5 347.6 ;
      RECT  184.3 344.4 185.5 345.2 ;
      RECT  179.7 341.4 187.3 342.2 ;
      RECT  179.7 342.8 180.5 347.0 ;
      RECT  182.3 344.0 183.1 346.2 ;
      RECT  184.1 340.0 185.7 340.8 ;
      RECT  186.5 347.6 187.3 349.2 ;
      RECT  181.3 340.0 182.9 340.8 ;
      RECT  182.1 356.0 183.1 355.2 ;
      RECT  184.5 351.6 185.5 350.8 ;
      RECT  184.7 355.2 185.5 354.8 ;
      RECT  183.5 357.0 184.3 356.8 ;
      RECT  186.5 356.4 187.3 352.2 ;
      RECT  182.3 353.0 183.9 352.2 ;
      RECT  184.5 350.8 185.3 350.0 ;
      RECT  184.7 356.0 185.7 355.2 ;
      RECT  179.7 350.0 187.3 349.2 ;
      RECT  179.7 351.6 180.5 350.0 ;
      RECT  182.3 351.6 183.3 350.8 ;
      RECT  182.3 352.2 183.1 351.6 ;
      RECT  184.7 354.0 185.5 351.6 ;
      RECT  184.3 354.8 185.5 354.0 ;
      RECT  179.7 357.8 187.3 357.0 ;
      RECT  179.7 356.4 180.5 352.2 ;
      RECT  182.3 355.2 183.1 353.0 ;
      RECT  184.1 359.2 185.7 358.4 ;
      RECT  186.5 351.6 187.3 350.0 ;
      RECT  181.3 359.2 182.9 358.4 ;
      RECT  182.1 364.0 183.1 364.8 ;
      RECT  184.5 368.4 185.5 369.2 ;
      RECT  184.7 364.8 185.5 365.2 ;
      RECT  183.5 363.0 184.3 363.2 ;
      RECT  186.5 363.6 187.3 367.8 ;
      RECT  182.3 367.0 183.9 367.8 ;
      RECT  184.7 364.0 185.7 364.8 ;
      RECT  182.1 360.8 182.9 361.6 ;
      RECT  179.7 370.0 187.3 370.8 ;
      RECT  179.7 368.4 180.5 370.0 ;
      RECT  182.3 368.4 183.3 369.2 ;
      RECT  182.3 367.8 183.1 368.4 ;
      RECT  184.7 366.0 185.5 368.4 ;
      RECT  184.3 365.2 185.5 366.0 ;
      RECT  179.7 362.2 187.3 363.0 ;
      RECT  184.9 360.8 185.7 361.6 ;
      RECT  179.7 363.6 180.5 367.8 ;
      RECT  182.3 364.8 183.1 367.0 ;
      RECT  186.5 368.4 187.3 370.0 ;
      RECT  180.1 175.0 186.9 175.8 ;
      RECT  180.1 190.6 186.9 191.4 ;
      RECT  180.1 195.8 186.9 196.6 ;
      RECT  180.1 211.4 186.9 212.2 ;
      RECT  180.1 216.6 186.9 217.4 ;
      RECT  180.1 232.2 186.9 233.0 ;
      RECT  180.1 237.4 186.9 238.2 ;
      RECT  180.1 253.0 186.9 253.8 ;
      RECT  180.1 258.2 186.9 259.0 ;
      RECT  180.1 273.8 186.9 274.6 ;
      RECT  180.1 279.0 186.9 279.8 ;
      RECT  180.1 294.6 186.9 295.4 ;
      RECT  180.1 299.8 186.9 300.6 ;
      RECT  180.1 315.4 186.9 316.2 ;
      RECT  180.1 320.6 186.9 321.4 ;
      RECT  180.1 336.2 186.9 337.0 ;
      RECT  180.1 341.4 186.9 342.2 ;
      RECT  180.1 357.0 186.9 357.8 ;
      RECT  180.1 362.2 186.9 363.0 ;
      RECT  188.9 189.6 189.9 188.8 ;
      RECT  191.3 185.2 192.3 184.4 ;
      RECT  191.5 188.8 192.3 188.4 ;
      RECT  190.3 190.6 191.1 190.4 ;
      RECT  193.3 190.0 194.1 185.8 ;
      RECT  189.1 186.6 190.7 185.8 ;
      RECT  191.5 189.6 192.5 188.8 ;
      RECT  188.9 192.8 189.7 192.0 ;
      RECT  186.5 183.6 194.1 182.8 ;
      RECT  186.5 185.2 187.3 183.6 ;
      RECT  189.1 185.2 190.1 184.4 ;
      RECT  189.1 185.8 189.9 185.2 ;
      RECT  191.5 187.6 192.3 185.2 ;
      RECT  191.1 188.4 192.3 187.6 ;
      RECT  186.5 191.4 194.1 190.6 ;
      RECT  191.7 192.8 192.5 192.0 ;
      RECT  186.5 190.0 187.3 185.8 ;
      RECT  189.1 188.8 189.9 186.6 ;
      RECT  193.3 185.2 194.1 183.6 ;
      RECT  195.7 189.6 196.7 188.8 ;
      RECT  198.1 185.2 199.1 184.4 ;
      RECT  198.3 188.8 199.1 188.4 ;
      RECT  197.1 190.6 197.9 190.4 ;
      RECT  200.1 190.0 200.9 185.8 ;
      RECT  195.9 186.6 197.5 185.8 ;
      RECT  198.3 189.6 199.3 188.8 ;
      RECT  195.7 192.8 196.5 192.0 ;
      RECT  193.3 183.6 200.9 182.8 ;
      RECT  193.3 185.2 194.1 183.6 ;
      RECT  195.9 185.2 196.9 184.4 ;
      RECT  195.9 185.8 196.7 185.2 ;
      RECT  198.3 187.6 199.1 185.2 ;
      RECT  197.9 188.4 199.1 187.6 ;
      RECT  193.3 191.4 200.9 190.6 ;
      RECT  198.5 192.8 199.3 192.0 ;
      RECT  193.3 190.0 194.1 185.8 ;
      RECT  195.9 188.8 196.7 186.6 ;
      RECT  200.1 185.2 200.9 183.6 ;
      RECT  186.9 191.4 200.5 190.6 ;
      RECT  188.9 176.8 189.9 177.6 ;
      RECT  191.3 181.2 192.3 182.0 ;
      RECT  191.5 177.6 192.3 178.0 ;
      RECT  190.3 175.8 191.1 176.0 ;
      RECT  193.3 176.4 194.1 180.6 ;
      RECT  189.1 179.8 190.7 180.6 ;
      RECT  191.5 176.8 192.5 177.6 ;
      RECT  188.9 173.6 189.7 174.4 ;
      RECT  186.5 182.8 194.1 183.6 ;
      RECT  186.5 181.2 187.3 182.8 ;
      RECT  189.1 181.2 190.1 182.0 ;
      RECT  189.1 180.6 189.9 181.2 ;
      RECT  191.5 178.8 192.3 181.2 ;
      RECT  191.1 178.0 192.3 178.8 ;
      RECT  186.5 175.0 194.1 175.8 ;
      RECT  191.7 173.6 192.5 174.4 ;
      RECT  186.5 176.4 187.3 180.6 ;
      RECT  189.1 177.6 189.9 179.8 ;
      RECT  193.3 181.2 194.1 182.8 ;
      RECT  195.7 176.8 196.7 177.6 ;
      RECT  198.1 181.2 199.1 182.0 ;
      RECT  198.3 177.6 199.1 178.0 ;
      RECT  197.1 175.8 197.9 176.0 ;
      RECT  200.1 176.4 200.9 180.6 ;
      RECT  195.9 179.8 197.5 180.6 ;
      RECT  198.3 176.8 199.3 177.6 ;
      RECT  195.7 173.6 196.5 174.4 ;
      RECT  193.3 182.8 200.9 183.6 ;
      RECT  193.3 181.2 194.1 182.8 ;
      RECT  195.9 181.2 196.9 182.0 ;
      RECT  195.9 180.6 196.7 181.2 ;
      RECT  198.3 178.8 199.1 181.2 ;
      RECT  197.9 178.0 199.1 178.8 ;
      RECT  193.3 175.0 200.9 175.8 ;
      RECT  198.5 173.6 199.3 174.4 ;
      RECT  193.3 176.4 194.1 180.6 ;
      RECT  195.9 177.6 196.7 179.8 ;
      RECT  200.1 181.2 200.9 182.8 ;
      RECT  186.9 175.0 200.5 175.8 ;
      RECT  188.9 364.0 189.9 364.8 ;
      RECT  191.3 368.4 192.3 369.2 ;
      RECT  191.5 364.8 192.3 365.2 ;
      RECT  190.3 363.0 191.1 363.2 ;
      RECT  193.3 363.6 194.1 367.8 ;
      RECT  189.1 367.0 190.7 367.8 ;
      RECT  191.5 364.0 192.5 364.8 ;
      RECT  188.9 360.8 189.7 361.6 ;
      RECT  186.5 370.0 194.1 370.8 ;
      RECT  186.5 368.4 187.3 370.0 ;
      RECT  189.1 368.4 190.1 369.2 ;
      RECT  189.1 367.8 189.9 368.4 ;
      RECT  191.5 366.0 192.3 368.4 ;
      RECT  191.1 365.2 192.3 366.0 ;
      RECT  186.5 362.2 194.1 363.0 ;
      RECT  191.7 360.8 192.5 361.6 ;
      RECT  186.5 363.6 187.3 367.8 ;
      RECT  189.1 364.8 189.9 367.0 ;
      RECT  193.3 368.4 194.1 370.0 ;
      RECT  195.7 364.0 196.7 364.8 ;
      RECT  198.1 368.4 199.1 369.2 ;
      RECT  198.3 364.8 199.1 365.2 ;
      RECT  197.1 363.0 197.9 363.2 ;
      RECT  200.1 363.6 200.9 367.8 ;
      RECT  195.9 367.0 197.5 367.8 ;
      RECT  198.3 364.0 199.3 364.8 ;
      RECT  195.7 360.8 196.5 361.6 ;
      RECT  193.3 370.0 200.9 370.8 ;
      RECT  193.3 368.4 194.1 370.0 ;
      RECT  195.9 368.4 196.9 369.2 ;
      RECT  195.9 367.8 196.7 368.4 ;
      RECT  198.3 366.0 199.1 368.4 ;
      RECT  197.9 365.2 199.1 366.0 ;
      RECT  193.3 362.2 200.9 363.0 ;
      RECT  198.5 360.8 199.3 361.6 ;
      RECT  193.3 363.6 194.1 367.8 ;
      RECT  195.9 364.8 196.7 367.0 ;
      RECT  200.1 368.4 200.9 370.0 ;
      RECT  186.9 362.2 200.5 363.0 ;
      RECT  175.3 176.8 176.3 177.6 ;
      RECT  177.7 181.2 178.7 182.0 ;
      RECT  177.9 177.6 178.7 178.0 ;
      RECT  176.7 175.8 177.5 176.0 ;
      RECT  179.7 176.4 180.5 180.6 ;
      RECT  175.5 179.8 177.1 180.6 ;
      RECT  177.9 176.8 178.9 177.6 ;
      RECT  175.3 173.6 176.1 174.4 ;
      RECT  172.9 182.8 180.5 183.6 ;
      RECT  172.9 181.2 173.7 182.8 ;
      RECT  175.5 181.2 176.5 182.0 ;
      RECT  175.5 180.6 176.3 181.2 ;
      RECT  177.9 178.8 178.7 181.2 ;
      RECT  177.5 178.0 178.7 178.8 ;
      RECT  172.9 175.0 180.5 175.8 ;
      RECT  178.1 173.6 178.9 174.4 ;
      RECT  172.9 176.4 173.7 180.6 ;
      RECT  175.5 177.6 176.3 179.8 ;
      RECT  179.7 181.2 180.5 182.8 ;
      RECT  175.3 189.6 176.3 188.8 ;
      RECT  177.7 185.2 178.7 184.4 ;
      RECT  177.9 188.8 178.7 188.4 ;
      RECT  176.7 190.6 177.5 190.4 ;
      RECT  179.7 190.0 180.5 185.8 ;
      RECT  175.5 186.6 177.1 185.8 ;
      RECT  177.9 189.6 178.9 188.8 ;
      RECT  175.3 192.8 176.1 192.0 ;
      RECT  172.9 183.6 180.5 182.8 ;
      RECT  172.9 185.2 173.7 183.6 ;
      RECT  175.5 185.2 176.5 184.4 ;
      RECT  175.5 185.8 176.3 185.2 ;
      RECT  177.9 187.6 178.7 185.2 ;
      RECT  177.5 188.4 178.7 187.6 ;
      RECT  172.9 191.4 180.5 190.6 ;
      RECT  178.1 192.8 178.9 192.0 ;
      RECT  172.9 190.0 173.7 185.8 ;
      RECT  175.5 188.8 176.3 186.6 ;
      RECT  179.7 185.2 180.5 183.6 ;
      RECT  175.3 197.6 176.3 198.4 ;
      RECT  177.7 202.0 178.7 202.8 ;
      RECT  177.9 198.4 178.7 198.8 ;
      RECT  176.7 196.6 177.5 196.8 ;
      RECT  179.7 197.2 180.5 201.4 ;
      RECT  175.5 200.6 177.1 201.4 ;
      RECT  177.9 197.6 178.9 198.4 ;
      RECT  175.3 194.4 176.1 195.2 ;
      RECT  172.9 203.6 180.5 204.4 ;
      RECT  172.9 202.0 173.7 203.6 ;
      RECT  175.5 202.0 176.5 202.8 ;
      RECT  175.5 201.4 176.3 202.0 ;
      RECT  177.9 199.6 178.7 202.0 ;
      RECT  177.5 198.8 178.7 199.6 ;
      RECT  172.9 195.8 180.5 196.6 ;
      RECT  178.1 194.4 178.9 195.2 ;
      RECT  172.9 197.2 173.7 201.4 ;
      RECT  175.5 198.4 176.3 200.6 ;
      RECT  179.7 202.0 180.5 203.6 ;
      RECT  175.3 210.4 176.3 209.6 ;
      RECT  177.7 206.0 178.7 205.2 ;
      RECT  177.9 209.6 178.7 209.2 ;
      RECT  176.7 211.4 177.5 211.2 ;
      RECT  179.7 210.8 180.5 206.6 ;
      RECT  175.5 207.4 177.1 206.6 ;
      RECT  177.9 210.4 178.9 209.6 ;
      RECT  175.3 213.6 176.1 212.8 ;
      RECT  172.9 204.4 180.5 203.6 ;
      RECT  172.9 206.0 173.7 204.4 ;
      RECT  175.5 206.0 176.5 205.2 ;
      RECT  175.5 206.6 176.3 206.0 ;
      RECT  177.9 208.4 178.7 206.0 ;
      RECT  177.5 209.2 178.7 208.4 ;
      RECT  172.9 212.2 180.5 211.4 ;
      RECT  178.1 213.6 178.9 212.8 ;
      RECT  172.9 210.8 173.7 206.6 ;
      RECT  175.5 209.6 176.3 207.4 ;
      RECT  179.7 206.0 180.5 204.4 ;
      RECT  175.3 218.4 176.3 219.2 ;
      RECT  177.7 222.8 178.7 223.6 ;
      RECT  177.9 219.2 178.7 219.6 ;
      RECT  176.7 217.4 177.5 217.6 ;
      RECT  179.7 218.0 180.5 222.2 ;
      RECT  175.5 221.4 177.1 222.2 ;
      RECT  177.9 218.4 178.9 219.2 ;
      RECT  175.3 215.2 176.1 216.0 ;
      RECT  172.9 224.4 180.5 225.2 ;
      RECT  172.9 222.8 173.7 224.4 ;
      RECT  175.5 222.8 176.5 223.6 ;
      RECT  175.5 222.2 176.3 222.8 ;
      RECT  177.9 220.4 178.7 222.8 ;
      RECT  177.5 219.6 178.7 220.4 ;
      RECT  172.9 216.6 180.5 217.4 ;
      RECT  178.1 215.2 178.9 216.0 ;
      RECT  172.9 218.0 173.7 222.2 ;
      RECT  175.5 219.2 176.3 221.4 ;
      RECT  179.7 222.8 180.5 224.4 ;
      RECT  175.3 231.2 176.3 230.4 ;
      RECT  177.7 226.8 178.7 226.0 ;
      RECT  177.9 230.4 178.7 230.0 ;
      RECT  176.7 232.2 177.5 232.0 ;
      RECT  179.7 231.6 180.5 227.4 ;
      RECT  175.5 228.2 177.1 227.4 ;
      RECT  177.9 231.2 178.9 230.4 ;
      RECT  175.3 234.4 176.1 233.6 ;
      RECT  172.9 225.2 180.5 224.4 ;
      RECT  172.9 226.8 173.7 225.2 ;
      RECT  175.5 226.8 176.5 226.0 ;
      RECT  175.5 227.4 176.3 226.8 ;
      RECT  177.9 229.2 178.7 226.8 ;
      RECT  177.5 230.0 178.7 229.2 ;
      RECT  172.9 233.0 180.5 232.2 ;
      RECT  178.1 234.4 178.9 233.6 ;
      RECT  172.9 231.6 173.7 227.4 ;
      RECT  175.5 230.4 176.3 228.2 ;
      RECT  179.7 226.8 180.5 225.2 ;
      RECT  175.3 239.2 176.3 240.0 ;
      RECT  177.7 243.6 178.7 244.4 ;
      RECT  177.9 240.0 178.7 240.4 ;
      RECT  176.7 238.2 177.5 238.4 ;
      RECT  179.7 238.8 180.5 243.0 ;
      RECT  175.5 242.2 177.1 243.0 ;
      RECT  177.9 239.2 178.9 240.0 ;
      RECT  175.3 236.0 176.1 236.8 ;
      RECT  172.9 245.2 180.5 246.0 ;
      RECT  172.9 243.6 173.7 245.2 ;
      RECT  175.5 243.6 176.5 244.4 ;
      RECT  175.5 243.0 176.3 243.6 ;
      RECT  177.9 241.2 178.7 243.6 ;
      RECT  177.5 240.4 178.7 241.2 ;
      RECT  172.9 237.4 180.5 238.2 ;
      RECT  178.1 236.0 178.9 236.8 ;
      RECT  172.9 238.8 173.7 243.0 ;
      RECT  175.5 240.0 176.3 242.2 ;
      RECT  179.7 243.6 180.5 245.2 ;
      RECT  175.3 252.0 176.3 251.2 ;
      RECT  177.7 247.6 178.7 246.8 ;
      RECT  177.9 251.2 178.7 250.8 ;
      RECT  176.7 253.0 177.5 252.8 ;
      RECT  179.7 252.4 180.5 248.2 ;
      RECT  175.5 249.0 177.1 248.2 ;
      RECT  177.9 252.0 178.9 251.2 ;
      RECT  175.3 255.2 176.1 254.4 ;
      RECT  172.9 246.0 180.5 245.2 ;
      RECT  172.9 247.6 173.7 246.0 ;
      RECT  175.5 247.6 176.5 246.8 ;
      RECT  175.5 248.2 176.3 247.6 ;
      RECT  177.9 250.0 178.7 247.6 ;
      RECT  177.5 250.8 178.7 250.0 ;
      RECT  172.9 253.8 180.5 253.0 ;
      RECT  178.1 255.2 178.9 254.4 ;
      RECT  172.9 252.4 173.7 248.2 ;
      RECT  175.5 251.2 176.3 249.0 ;
      RECT  179.7 247.6 180.5 246.0 ;
      RECT  175.3 260.0 176.3 260.8 ;
      RECT  177.7 264.4 178.7 265.2 ;
      RECT  177.9 260.8 178.7 261.2 ;
      RECT  176.7 259.0 177.5 259.2 ;
      RECT  179.7 259.6 180.5 263.8 ;
      RECT  175.5 263.0 177.1 263.8 ;
      RECT  177.9 260.0 178.9 260.8 ;
      RECT  175.3 256.8 176.1 257.6 ;
      RECT  172.9 266.0 180.5 266.8 ;
      RECT  172.9 264.4 173.7 266.0 ;
      RECT  175.5 264.4 176.5 265.2 ;
      RECT  175.5 263.8 176.3 264.4 ;
      RECT  177.9 262.0 178.7 264.4 ;
      RECT  177.5 261.2 178.7 262.0 ;
      RECT  172.9 258.2 180.5 259.0 ;
      RECT  178.1 256.8 178.9 257.6 ;
      RECT  172.9 259.6 173.7 263.8 ;
      RECT  175.5 260.8 176.3 263.0 ;
      RECT  179.7 264.4 180.5 266.0 ;
      RECT  175.3 272.8 176.3 272.0 ;
      RECT  177.7 268.4 178.7 267.6 ;
      RECT  177.9 272.0 178.7 271.6 ;
      RECT  176.7 273.8 177.5 273.6 ;
      RECT  179.7 273.2 180.5 269.0 ;
      RECT  175.5 269.8 177.1 269.0 ;
      RECT  177.9 272.8 178.9 272.0 ;
      RECT  175.3 276.0 176.1 275.2 ;
      RECT  172.9 266.8 180.5 266.0 ;
      RECT  172.9 268.4 173.7 266.8 ;
      RECT  175.5 268.4 176.5 267.6 ;
      RECT  175.5 269.0 176.3 268.4 ;
      RECT  177.9 270.8 178.7 268.4 ;
      RECT  177.5 271.6 178.7 270.8 ;
      RECT  172.9 274.6 180.5 273.8 ;
      RECT  178.1 276.0 178.9 275.2 ;
      RECT  172.9 273.2 173.7 269.0 ;
      RECT  175.5 272.0 176.3 269.8 ;
      RECT  179.7 268.4 180.5 266.8 ;
      RECT  175.3 280.8 176.3 281.6 ;
      RECT  177.7 285.2 178.7 286.0 ;
      RECT  177.9 281.6 178.7 282.0 ;
      RECT  176.7 279.8 177.5 280.0 ;
      RECT  179.7 280.4 180.5 284.6 ;
      RECT  175.5 283.8 177.1 284.6 ;
      RECT  177.9 280.8 178.9 281.6 ;
      RECT  175.3 277.6 176.1 278.4 ;
      RECT  172.9 286.8 180.5 287.6 ;
      RECT  172.9 285.2 173.7 286.8 ;
      RECT  175.5 285.2 176.5 286.0 ;
      RECT  175.5 284.6 176.3 285.2 ;
      RECT  177.9 282.8 178.7 285.2 ;
      RECT  177.5 282.0 178.7 282.8 ;
      RECT  172.9 279.0 180.5 279.8 ;
      RECT  178.1 277.6 178.9 278.4 ;
      RECT  172.9 280.4 173.7 284.6 ;
      RECT  175.5 281.6 176.3 283.8 ;
      RECT  179.7 285.2 180.5 286.8 ;
      RECT  175.3 293.6 176.3 292.8 ;
      RECT  177.7 289.2 178.7 288.4 ;
      RECT  177.9 292.8 178.7 292.4 ;
      RECT  176.7 294.6 177.5 294.4 ;
      RECT  179.7 294.0 180.5 289.8 ;
      RECT  175.5 290.6 177.1 289.8 ;
      RECT  177.9 293.6 178.9 292.8 ;
      RECT  175.3 296.8 176.1 296.0 ;
      RECT  172.9 287.6 180.5 286.8 ;
      RECT  172.9 289.2 173.7 287.6 ;
      RECT  175.5 289.2 176.5 288.4 ;
      RECT  175.5 289.8 176.3 289.2 ;
      RECT  177.9 291.6 178.7 289.2 ;
      RECT  177.5 292.4 178.7 291.6 ;
      RECT  172.9 295.4 180.5 294.6 ;
      RECT  178.1 296.8 178.9 296.0 ;
      RECT  172.9 294.0 173.7 289.8 ;
      RECT  175.5 292.8 176.3 290.6 ;
      RECT  179.7 289.2 180.5 287.6 ;
      RECT  175.3 301.6 176.3 302.4 ;
      RECT  177.7 306.0 178.7 306.8 ;
      RECT  177.9 302.4 178.7 302.8 ;
      RECT  176.7 300.6 177.5 300.8 ;
      RECT  179.7 301.2 180.5 305.4 ;
      RECT  175.5 304.6 177.1 305.4 ;
      RECT  177.9 301.6 178.9 302.4 ;
      RECT  175.3 298.4 176.1 299.2 ;
      RECT  172.9 307.6 180.5 308.4 ;
      RECT  172.9 306.0 173.7 307.6 ;
      RECT  175.5 306.0 176.5 306.8 ;
      RECT  175.5 305.4 176.3 306.0 ;
      RECT  177.9 303.6 178.7 306.0 ;
      RECT  177.5 302.8 178.7 303.6 ;
      RECT  172.9 299.8 180.5 300.6 ;
      RECT  178.1 298.4 178.9 299.2 ;
      RECT  172.9 301.2 173.7 305.4 ;
      RECT  175.5 302.4 176.3 304.6 ;
      RECT  179.7 306.0 180.5 307.6 ;
      RECT  175.3 314.4 176.3 313.6 ;
      RECT  177.7 310.0 178.7 309.2 ;
      RECT  177.9 313.6 178.7 313.2 ;
      RECT  176.7 315.4 177.5 315.2 ;
      RECT  179.7 314.8 180.5 310.6 ;
      RECT  175.5 311.4 177.1 310.6 ;
      RECT  177.9 314.4 178.9 313.6 ;
      RECT  175.3 317.6 176.1 316.8 ;
      RECT  172.9 308.4 180.5 307.6 ;
      RECT  172.9 310.0 173.7 308.4 ;
      RECT  175.5 310.0 176.5 309.2 ;
      RECT  175.5 310.6 176.3 310.0 ;
      RECT  177.9 312.4 178.7 310.0 ;
      RECT  177.5 313.2 178.7 312.4 ;
      RECT  172.9 316.2 180.5 315.4 ;
      RECT  178.1 317.6 178.9 316.8 ;
      RECT  172.9 314.8 173.7 310.6 ;
      RECT  175.5 313.6 176.3 311.4 ;
      RECT  179.7 310.0 180.5 308.4 ;
      RECT  175.3 322.4 176.3 323.2 ;
      RECT  177.7 326.8 178.7 327.6 ;
      RECT  177.9 323.2 178.7 323.6 ;
      RECT  176.7 321.4 177.5 321.6 ;
      RECT  179.7 322.0 180.5 326.2 ;
      RECT  175.5 325.4 177.1 326.2 ;
      RECT  177.9 322.4 178.9 323.2 ;
      RECT  175.3 319.2 176.1 320.0 ;
      RECT  172.9 328.4 180.5 329.2 ;
      RECT  172.9 326.8 173.7 328.4 ;
      RECT  175.5 326.8 176.5 327.6 ;
      RECT  175.5 326.2 176.3 326.8 ;
      RECT  177.9 324.4 178.7 326.8 ;
      RECT  177.5 323.6 178.7 324.4 ;
      RECT  172.9 320.6 180.5 321.4 ;
      RECT  178.1 319.2 178.9 320.0 ;
      RECT  172.9 322.0 173.7 326.2 ;
      RECT  175.5 323.2 176.3 325.4 ;
      RECT  179.7 326.8 180.5 328.4 ;
      RECT  175.3 335.2 176.3 334.4 ;
      RECT  177.7 330.8 178.7 330.0 ;
      RECT  177.9 334.4 178.7 334.0 ;
      RECT  176.7 336.2 177.5 336.0 ;
      RECT  179.7 335.6 180.5 331.4 ;
      RECT  175.5 332.2 177.1 331.4 ;
      RECT  177.9 335.2 178.9 334.4 ;
      RECT  175.3 338.4 176.1 337.6 ;
      RECT  172.9 329.2 180.5 328.4 ;
      RECT  172.9 330.8 173.7 329.2 ;
      RECT  175.5 330.8 176.5 330.0 ;
      RECT  175.5 331.4 176.3 330.8 ;
      RECT  177.9 333.2 178.7 330.8 ;
      RECT  177.5 334.0 178.7 333.2 ;
      RECT  172.9 337.0 180.5 336.2 ;
      RECT  178.1 338.4 178.9 337.6 ;
      RECT  172.9 335.6 173.7 331.4 ;
      RECT  175.5 334.4 176.3 332.2 ;
      RECT  179.7 330.8 180.5 329.2 ;
      RECT  175.3 343.2 176.3 344.0 ;
      RECT  177.7 347.6 178.7 348.4 ;
      RECT  177.9 344.0 178.7 344.4 ;
      RECT  176.7 342.2 177.5 342.4 ;
      RECT  179.7 342.8 180.5 347.0 ;
      RECT  175.5 346.2 177.1 347.0 ;
      RECT  177.9 343.2 178.9 344.0 ;
      RECT  175.3 340.0 176.1 340.8 ;
      RECT  172.9 349.2 180.5 350.0 ;
      RECT  172.9 347.6 173.7 349.2 ;
      RECT  175.5 347.6 176.5 348.4 ;
      RECT  175.5 347.0 176.3 347.6 ;
      RECT  177.9 345.2 178.7 347.6 ;
      RECT  177.5 344.4 178.7 345.2 ;
      RECT  172.9 341.4 180.5 342.2 ;
      RECT  178.1 340.0 178.9 340.8 ;
      RECT  172.9 342.8 173.7 347.0 ;
      RECT  175.5 344.0 176.3 346.2 ;
      RECT  179.7 347.6 180.5 349.2 ;
      RECT  175.3 356.0 176.3 355.2 ;
      RECT  177.7 351.6 178.7 350.8 ;
      RECT  177.9 355.2 178.7 354.8 ;
      RECT  176.7 357.0 177.5 356.8 ;
      RECT  179.7 356.4 180.5 352.2 ;
      RECT  175.5 353.0 177.1 352.2 ;
      RECT  177.9 356.0 178.9 355.2 ;
      RECT  175.3 359.2 176.1 358.4 ;
      RECT  172.9 350.0 180.5 349.2 ;
      RECT  172.9 351.6 173.7 350.0 ;
      RECT  175.5 351.6 176.5 350.8 ;
      RECT  175.5 352.2 176.3 351.6 ;
      RECT  177.9 354.0 178.7 351.6 ;
      RECT  177.5 354.8 178.7 354.0 ;
      RECT  172.9 357.8 180.5 357.0 ;
      RECT  178.1 359.2 178.9 358.4 ;
      RECT  172.9 356.4 173.7 352.2 ;
      RECT  175.5 355.2 176.3 353.0 ;
      RECT  179.7 351.6 180.5 350.0 ;
      RECT  175.3 364.0 176.3 364.8 ;
      RECT  177.7 368.4 178.7 369.2 ;
      RECT  177.9 364.8 178.7 365.2 ;
      RECT  176.7 363.0 177.5 363.2 ;
      RECT  179.7 363.6 180.5 367.8 ;
      RECT  175.5 367.0 177.1 367.8 ;
      RECT  177.9 364.0 178.9 364.8 ;
      RECT  175.3 360.8 176.1 361.6 ;
      RECT  172.9 370.0 180.5 370.8 ;
      RECT  172.9 368.4 173.7 370.0 ;
      RECT  175.5 368.4 176.5 369.2 ;
      RECT  175.5 367.8 176.3 368.4 ;
      RECT  177.9 366.0 178.7 368.4 ;
      RECT  177.5 365.2 178.7 366.0 ;
      RECT  172.9 362.2 180.5 363.0 ;
      RECT  178.1 360.8 178.9 361.6 ;
      RECT  172.9 363.6 173.7 367.8 ;
      RECT  175.5 364.8 176.3 367.0 ;
      RECT  179.7 368.4 180.5 370.0 ;
      RECT  173.3 175.0 180.1 175.8 ;
      RECT  173.3 190.6 180.1 191.4 ;
      RECT  173.3 195.8 180.1 196.6 ;
      RECT  173.3 211.4 180.1 212.2 ;
      RECT  173.3 216.6 180.1 217.4 ;
      RECT  173.3 232.2 180.1 233.0 ;
      RECT  173.3 237.4 180.1 238.2 ;
      RECT  173.3 253.0 180.1 253.8 ;
      RECT  173.3 258.2 180.1 259.0 ;
      RECT  173.3 273.8 180.1 274.6 ;
      RECT  173.3 279.0 180.1 279.8 ;
      RECT  173.3 294.6 180.1 295.4 ;
      RECT  173.3 299.8 180.1 300.6 ;
      RECT  173.3 315.4 180.1 316.2 ;
      RECT  173.3 320.6 180.1 321.4 ;
      RECT  173.3 336.2 180.1 337.0 ;
      RECT  173.3 341.4 180.1 342.2 ;
      RECT  173.3 357.0 180.1 357.8 ;
      RECT  173.3 362.2 180.1 363.0 ;
      RECT  202.5 176.8 203.5 177.6 ;
      RECT  204.9 181.2 205.9 182.0 ;
      RECT  205.1 177.6 205.9 178.0 ;
      RECT  203.9 175.8 204.7 176.0 ;
      RECT  206.9 176.4 207.7 180.6 ;
      RECT  202.7 179.8 204.3 180.6 ;
      RECT  205.1 176.8 206.1 177.6 ;
      RECT  202.5 173.6 203.3 174.4 ;
      RECT  200.1 182.8 207.7 183.6 ;
      RECT  200.1 181.2 200.9 182.8 ;
      RECT  202.7 181.2 203.7 182.0 ;
      RECT  202.7 180.6 203.5 181.2 ;
      RECT  205.1 178.8 205.9 181.2 ;
      RECT  204.7 178.0 205.9 178.8 ;
      RECT  200.1 175.0 207.7 175.8 ;
      RECT  205.3 173.6 206.1 174.4 ;
      RECT  200.1 176.4 200.9 180.6 ;
      RECT  202.7 177.6 203.5 179.8 ;
      RECT  206.9 181.2 207.7 182.8 ;
      RECT  202.5 189.6 203.5 188.8 ;
      RECT  204.9 185.2 205.9 184.4 ;
      RECT  205.1 188.8 205.9 188.4 ;
      RECT  203.9 190.6 204.7 190.4 ;
      RECT  206.9 190.0 207.7 185.8 ;
      RECT  202.7 186.6 204.3 185.8 ;
      RECT  205.1 189.6 206.1 188.8 ;
      RECT  202.5 192.8 203.3 192.0 ;
      RECT  200.1 183.6 207.7 182.8 ;
      RECT  200.1 185.2 200.9 183.6 ;
      RECT  202.7 185.2 203.7 184.4 ;
      RECT  202.7 185.8 203.5 185.2 ;
      RECT  205.1 187.6 205.9 185.2 ;
      RECT  204.7 188.4 205.9 187.6 ;
      RECT  200.1 191.4 207.7 190.6 ;
      RECT  205.3 192.8 206.1 192.0 ;
      RECT  200.1 190.0 200.9 185.8 ;
      RECT  202.7 188.8 203.5 186.6 ;
      RECT  206.9 185.2 207.7 183.6 ;
      RECT  202.5 197.6 203.5 198.4 ;
      RECT  204.9 202.0 205.9 202.8 ;
      RECT  205.1 198.4 205.9 198.8 ;
      RECT  203.9 196.6 204.7 196.8 ;
      RECT  206.9 197.2 207.7 201.4 ;
      RECT  202.7 200.6 204.3 201.4 ;
      RECT  205.1 197.6 206.1 198.4 ;
      RECT  202.5 194.4 203.3 195.2 ;
      RECT  200.1 203.6 207.7 204.4 ;
      RECT  200.1 202.0 200.9 203.6 ;
      RECT  202.7 202.0 203.7 202.8 ;
      RECT  202.7 201.4 203.5 202.0 ;
      RECT  205.1 199.6 205.9 202.0 ;
      RECT  204.7 198.8 205.9 199.6 ;
      RECT  200.1 195.8 207.7 196.6 ;
      RECT  205.3 194.4 206.1 195.2 ;
      RECT  200.1 197.2 200.9 201.4 ;
      RECT  202.7 198.4 203.5 200.6 ;
      RECT  206.9 202.0 207.7 203.6 ;
      RECT  202.5 210.4 203.5 209.6 ;
      RECT  204.9 206.0 205.9 205.2 ;
      RECT  205.1 209.6 205.9 209.2 ;
      RECT  203.9 211.4 204.7 211.2 ;
      RECT  206.9 210.8 207.7 206.6 ;
      RECT  202.7 207.4 204.3 206.6 ;
      RECT  205.1 210.4 206.1 209.6 ;
      RECT  202.5 213.6 203.3 212.8 ;
      RECT  200.1 204.4 207.7 203.6 ;
      RECT  200.1 206.0 200.9 204.4 ;
      RECT  202.7 206.0 203.7 205.2 ;
      RECT  202.7 206.6 203.5 206.0 ;
      RECT  205.1 208.4 205.9 206.0 ;
      RECT  204.7 209.2 205.9 208.4 ;
      RECT  200.1 212.2 207.7 211.4 ;
      RECT  205.3 213.6 206.1 212.8 ;
      RECT  200.1 210.8 200.9 206.6 ;
      RECT  202.7 209.6 203.5 207.4 ;
      RECT  206.9 206.0 207.7 204.4 ;
      RECT  202.5 218.4 203.5 219.2 ;
      RECT  204.9 222.8 205.9 223.6 ;
      RECT  205.1 219.2 205.9 219.6 ;
      RECT  203.9 217.4 204.7 217.6 ;
      RECT  206.9 218.0 207.7 222.2 ;
      RECT  202.7 221.4 204.3 222.2 ;
      RECT  205.1 218.4 206.1 219.2 ;
      RECT  202.5 215.2 203.3 216.0 ;
      RECT  200.1 224.4 207.7 225.2 ;
      RECT  200.1 222.8 200.9 224.4 ;
      RECT  202.7 222.8 203.7 223.6 ;
      RECT  202.7 222.2 203.5 222.8 ;
      RECT  205.1 220.4 205.9 222.8 ;
      RECT  204.7 219.6 205.9 220.4 ;
      RECT  200.1 216.6 207.7 217.4 ;
      RECT  205.3 215.2 206.1 216.0 ;
      RECT  200.1 218.0 200.9 222.2 ;
      RECT  202.7 219.2 203.5 221.4 ;
      RECT  206.9 222.8 207.7 224.4 ;
      RECT  202.5 231.2 203.5 230.4 ;
      RECT  204.9 226.8 205.9 226.0 ;
      RECT  205.1 230.4 205.9 230.0 ;
      RECT  203.9 232.2 204.7 232.0 ;
      RECT  206.9 231.6 207.7 227.4 ;
      RECT  202.7 228.2 204.3 227.4 ;
      RECT  205.1 231.2 206.1 230.4 ;
      RECT  202.5 234.4 203.3 233.6 ;
      RECT  200.1 225.2 207.7 224.4 ;
      RECT  200.1 226.8 200.9 225.2 ;
      RECT  202.7 226.8 203.7 226.0 ;
      RECT  202.7 227.4 203.5 226.8 ;
      RECT  205.1 229.2 205.9 226.8 ;
      RECT  204.7 230.0 205.9 229.2 ;
      RECT  200.1 233.0 207.7 232.2 ;
      RECT  205.3 234.4 206.1 233.6 ;
      RECT  200.1 231.6 200.9 227.4 ;
      RECT  202.7 230.4 203.5 228.2 ;
      RECT  206.9 226.8 207.7 225.2 ;
      RECT  202.5 239.2 203.5 240.0 ;
      RECT  204.9 243.6 205.9 244.4 ;
      RECT  205.1 240.0 205.9 240.4 ;
      RECT  203.9 238.2 204.7 238.4 ;
      RECT  206.9 238.8 207.7 243.0 ;
      RECT  202.7 242.2 204.3 243.0 ;
      RECT  205.1 239.2 206.1 240.0 ;
      RECT  202.5 236.0 203.3 236.8 ;
      RECT  200.1 245.2 207.7 246.0 ;
      RECT  200.1 243.6 200.9 245.2 ;
      RECT  202.7 243.6 203.7 244.4 ;
      RECT  202.7 243.0 203.5 243.6 ;
      RECT  205.1 241.2 205.9 243.6 ;
      RECT  204.7 240.4 205.9 241.2 ;
      RECT  200.1 237.4 207.7 238.2 ;
      RECT  205.3 236.0 206.1 236.8 ;
      RECT  200.1 238.8 200.9 243.0 ;
      RECT  202.7 240.0 203.5 242.2 ;
      RECT  206.9 243.6 207.7 245.2 ;
      RECT  202.5 252.0 203.5 251.2 ;
      RECT  204.9 247.6 205.9 246.8 ;
      RECT  205.1 251.2 205.9 250.8 ;
      RECT  203.9 253.0 204.7 252.8 ;
      RECT  206.9 252.4 207.7 248.2 ;
      RECT  202.7 249.0 204.3 248.2 ;
      RECT  205.1 252.0 206.1 251.2 ;
      RECT  202.5 255.2 203.3 254.4 ;
      RECT  200.1 246.0 207.7 245.2 ;
      RECT  200.1 247.6 200.9 246.0 ;
      RECT  202.7 247.6 203.7 246.8 ;
      RECT  202.7 248.2 203.5 247.6 ;
      RECT  205.1 250.0 205.9 247.6 ;
      RECT  204.7 250.8 205.9 250.0 ;
      RECT  200.1 253.8 207.7 253.0 ;
      RECT  205.3 255.2 206.1 254.4 ;
      RECT  200.1 252.4 200.9 248.2 ;
      RECT  202.7 251.2 203.5 249.0 ;
      RECT  206.9 247.6 207.7 246.0 ;
      RECT  202.5 260.0 203.5 260.8 ;
      RECT  204.9 264.4 205.9 265.2 ;
      RECT  205.1 260.8 205.9 261.2 ;
      RECT  203.9 259.0 204.7 259.2 ;
      RECT  206.9 259.6 207.7 263.8 ;
      RECT  202.7 263.0 204.3 263.8 ;
      RECT  205.1 260.0 206.1 260.8 ;
      RECT  202.5 256.8 203.3 257.6 ;
      RECT  200.1 266.0 207.7 266.8 ;
      RECT  200.1 264.4 200.9 266.0 ;
      RECT  202.7 264.4 203.7 265.2 ;
      RECT  202.7 263.8 203.5 264.4 ;
      RECT  205.1 262.0 205.9 264.4 ;
      RECT  204.7 261.2 205.9 262.0 ;
      RECT  200.1 258.2 207.7 259.0 ;
      RECT  205.3 256.8 206.1 257.6 ;
      RECT  200.1 259.6 200.9 263.8 ;
      RECT  202.7 260.8 203.5 263.0 ;
      RECT  206.9 264.4 207.7 266.0 ;
      RECT  202.5 272.8 203.5 272.0 ;
      RECT  204.9 268.4 205.9 267.6 ;
      RECT  205.1 272.0 205.9 271.6 ;
      RECT  203.9 273.8 204.7 273.6 ;
      RECT  206.9 273.2 207.7 269.0 ;
      RECT  202.7 269.8 204.3 269.0 ;
      RECT  205.1 272.8 206.1 272.0 ;
      RECT  202.5 276.0 203.3 275.2 ;
      RECT  200.1 266.8 207.7 266.0 ;
      RECT  200.1 268.4 200.9 266.8 ;
      RECT  202.7 268.4 203.7 267.6 ;
      RECT  202.7 269.0 203.5 268.4 ;
      RECT  205.1 270.8 205.9 268.4 ;
      RECT  204.7 271.6 205.9 270.8 ;
      RECT  200.1 274.6 207.7 273.8 ;
      RECT  205.3 276.0 206.1 275.2 ;
      RECT  200.1 273.2 200.9 269.0 ;
      RECT  202.7 272.0 203.5 269.8 ;
      RECT  206.9 268.4 207.7 266.8 ;
      RECT  202.5 280.8 203.5 281.6 ;
      RECT  204.9 285.2 205.9 286.0 ;
      RECT  205.1 281.6 205.9 282.0 ;
      RECT  203.9 279.8 204.7 280.0 ;
      RECT  206.9 280.4 207.7 284.6 ;
      RECT  202.7 283.8 204.3 284.6 ;
      RECT  205.1 280.8 206.1 281.6 ;
      RECT  202.5 277.6 203.3 278.4 ;
      RECT  200.1 286.8 207.7 287.6 ;
      RECT  200.1 285.2 200.9 286.8 ;
      RECT  202.7 285.2 203.7 286.0 ;
      RECT  202.7 284.6 203.5 285.2 ;
      RECT  205.1 282.8 205.9 285.2 ;
      RECT  204.7 282.0 205.9 282.8 ;
      RECT  200.1 279.0 207.7 279.8 ;
      RECT  205.3 277.6 206.1 278.4 ;
      RECT  200.1 280.4 200.9 284.6 ;
      RECT  202.7 281.6 203.5 283.8 ;
      RECT  206.9 285.2 207.7 286.8 ;
      RECT  202.5 293.6 203.5 292.8 ;
      RECT  204.9 289.2 205.9 288.4 ;
      RECT  205.1 292.8 205.9 292.4 ;
      RECT  203.9 294.6 204.7 294.4 ;
      RECT  206.9 294.0 207.7 289.8 ;
      RECT  202.7 290.6 204.3 289.8 ;
      RECT  205.1 293.6 206.1 292.8 ;
      RECT  202.5 296.8 203.3 296.0 ;
      RECT  200.1 287.6 207.7 286.8 ;
      RECT  200.1 289.2 200.9 287.6 ;
      RECT  202.7 289.2 203.7 288.4 ;
      RECT  202.7 289.8 203.5 289.2 ;
      RECT  205.1 291.6 205.9 289.2 ;
      RECT  204.7 292.4 205.9 291.6 ;
      RECT  200.1 295.4 207.7 294.6 ;
      RECT  205.3 296.8 206.1 296.0 ;
      RECT  200.1 294.0 200.9 289.8 ;
      RECT  202.7 292.8 203.5 290.6 ;
      RECT  206.9 289.2 207.7 287.6 ;
      RECT  202.5 301.6 203.5 302.4 ;
      RECT  204.9 306.0 205.9 306.8 ;
      RECT  205.1 302.4 205.9 302.8 ;
      RECT  203.9 300.6 204.7 300.8 ;
      RECT  206.9 301.2 207.7 305.4 ;
      RECT  202.7 304.6 204.3 305.4 ;
      RECT  205.1 301.6 206.1 302.4 ;
      RECT  202.5 298.4 203.3 299.2 ;
      RECT  200.1 307.6 207.7 308.4 ;
      RECT  200.1 306.0 200.9 307.6 ;
      RECT  202.7 306.0 203.7 306.8 ;
      RECT  202.7 305.4 203.5 306.0 ;
      RECT  205.1 303.6 205.9 306.0 ;
      RECT  204.7 302.8 205.9 303.6 ;
      RECT  200.1 299.8 207.7 300.6 ;
      RECT  205.3 298.4 206.1 299.2 ;
      RECT  200.1 301.2 200.9 305.4 ;
      RECT  202.7 302.4 203.5 304.6 ;
      RECT  206.9 306.0 207.7 307.6 ;
      RECT  202.5 314.4 203.5 313.6 ;
      RECT  204.9 310.0 205.9 309.2 ;
      RECT  205.1 313.6 205.9 313.2 ;
      RECT  203.9 315.4 204.7 315.2 ;
      RECT  206.9 314.8 207.7 310.6 ;
      RECT  202.7 311.4 204.3 310.6 ;
      RECT  205.1 314.4 206.1 313.6 ;
      RECT  202.5 317.6 203.3 316.8 ;
      RECT  200.1 308.4 207.7 307.6 ;
      RECT  200.1 310.0 200.9 308.4 ;
      RECT  202.7 310.0 203.7 309.2 ;
      RECT  202.7 310.6 203.5 310.0 ;
      RECT  205.1 312.4 205.9 310.0 ;
      RECT  204.7 313.2 205.9 312.4 ;
      RECT  200.1 316.2 207.7 315.4 ;
      RECT  205.3 317.6 206.1 316.8 ;
      RECT  200.1 314.8 200.9 310.6 ;
      RECT  202.7 313.6 203.5 311.4 ;
      RECT  206.9 310.0 207.7 308.4 ;
      RECT  202.5 322.4 203.5 323.2 ;
      RECT  204.9 326.8 205.9 327.6 ;
      RECT  205.1 323.2 205.9 323.6 ;
      RECT  203.9 321.4 204.7 321.6 ;
      RECT  206.9 322.0 207.7 326.2 ;
      RECT  202.7 325.4 204.3 326.2 ;
      RECT  205.1 322.4 206.1 323.2 ;
      RECT  202.5 319.2 203.3 320.0 ;
      RECT  200.1 328.4 207.7 329.2 ;
      RECT  200.1 326.8 200.9 328.4 ;
      RECT  202.7 326.8 203.7 327.6 ;
      RECT  202.7 326.2 203.5 326.8 ;
      RECT  205.1 324.4 205.9 326.8 ;
      RECT  204.7 323.6 205.9 324.4 ;
      RECT  200.1 320.6 207.7 321.4 ;
      RECT  205.3 319.2 206.1 320.0 ;
      RECT  200.1 322.0 200.9 326.2 ;
      RECT  202.7 323.2 203.5 325.4 ;
      RECT  206.9 326.8 207.7 328.4 ;
      RECT  202.5 335.2 203.5 334.4 ;
      RECT  204.9 330.8 205.9 330.0 ;
      RECT  205.1 334.4 205.9 334.0 ;
      RECT  203.9 336.2 204.7 336.0 ;
      RECT  206.9 335.6 207.7 331.4 ;
      RECT  202.7 332.2 204.3 331.4 ;
      RECT  205.1 335.2 206.1 334.4 ;
      RECT  202.5 338.4 203.3 337.6 ;
      RECT  200.1 329.2 207.7 328.4 ;
      RECT  200.1 330.8 200.9 329.2 ;
      RECT  202.7 330.8 203.7 330.0 ;
      RECT  202.7 331.4 203.5 330.8 ;
      RECT  205.1 333.2 205.9 330.8 ;
      RECT  204.7 334.0 205.9 333.2 ;
      RECT  200.1 337.0 207.7 336.2 ;
      RECT  205.3 338.4 206.1 337.6 ;
      RECT  200.1 335.6 200.9 331.4 ;
      RECT  202.7 334.4 203.5 332.2 ;
      RECT  206.9 330.8 207.7 329.2 ;
      RECT  202.5 343.2 203.5 344.0 ;
      RECT  204.9 347.6 205.9 348.4 ;
      RECT  205.1 344.0 205.9 344.4 ;
      RECT  203.9 342.2 204.7 342.4 ;
      RECT  206.9 342.8 207.7 347.0 ;
      RECT  202.7 346.2 204.3 347.0 ;
      RECT  205.1 343.2 206.1 344.0 ;
      RECT  202.5 340.0 203.3 340.8 ;
      RECT  200.1 349.2 207.7 350.0 ;
      RECT  200.1 347.6 200.9 349.2 ;
      RECT  202.7 347.6 203.7 348.4 ;
      RECT  202.7 347.0 203.5 347.6 ;
      RECT  205.1 345.2 205.9 347.6 ;
      RECT  204.7 344.4 205.9 345.2 ;
      RECT  200.1 341.4 207.7 342.2 ;
      RECT  205.3 340.0 206.1 340.8 ;
      RECT  200.1 342.8 200.9 347.0 ;
      RECT  202.7 344.0 203.5 346.2 ;
      RECT  206.9 347.6 207.7 349.2 ;
      RECT  202.5 356.0 203.5 355.2 ;
      RECT  204.9 351.6 205.9 350.8 ;
      RECT  205.1 355.2 205.9 354.8 ;
      RECT  203.9 357.0 204.7 356.8 ;
      RECT  206.9 356.4 207.7 352.2 ;
      RECT  202.7 353.0 204.3 352.2 ;
      RECT  205.1 356.0 206.1 355.2 ;
      RECT  202.5 359.2 203.3 358.4 ;
      RECT  200.1 350.0 207.7 349.2 ;
      RECT  200.1 351.6 200.9 350.0 ;
      RECT  202.7 351.6 203.7 350.8 ;
      RECT  202.7 352.2 203.5 351.6 ;
      RECT  205.1 354.0 205.9 351.6 ;
      RECT  204.7 354.8 205.9 354.0 ;
      RECT  200.1 357.8 207.7 357.0 ;
      RECT  205.3 359.2 206.1 358.4 ;
      RECT  200.1 356.4 200.9 352.2 ;
      RECT  202.7 355.2 203.5 353.0 ;
      RECT  206.9 351.6 207.7 350.0 ;
      RECT  202.5 364.0 203.5 364.8 ;
      RECT  204.9 368.4 205.9 369.2 ;
      RECT  205.1 364.8 205.9 365.2 ;
      RECT  203.9 363.0 204.7 363.2 ;
      RECT  206.9 363.6 207.7 367.8 ;
      RECT  202.7 367.0 204.3 367.8 ;
      RECT  205.1 364.0 206.1 364.8 ;
      RECT  202.5 360.8 203.3 361.6 ;
      RECT  200.1 370.0 207.7 370.8 ;
      RECT  200.1 368.4 200.9 370.0 ;
      RECT  202.7 368.4 203.7 369.2 ;
      RECT  202.7 367.8 203.5 368.4 ;
      RECT  205.1 366.0 205.9 368.4 ;
      RECT  204.7 365.2 205.9 366.0 ;
      RECT  200.1 362.2 207.7 363.0 ;
      RECT  205.3 360.8 206.1 361.6 ;
      RECT  200.1 363.6 200.9 367.8 ;
      RECT  202.7 364.8 203.5 367.0 ;
      RECT  206.9 368.4 207.7 370.0 ;
      RECT  200.5 175.0 207.3 175.8 ;
      RECT  200.5 190.6 207.3 191.4 ;
      RECT  200.5 195.8 207.3 196.6 ;
      RECT  200.5 211.4 207.3 212.2 ;
      RECT  200.5 216.6 207.3 217.4 ;
      RECT  200.5 232.2 207.3 233.0 ;
      RECT  200.5 237.4 207.3 238.2 ;
      RECT  200.5 253.0 207.3 253.8 ;
      RECT  200.5 258.2 207.3 259.0 ;
      RECT  200.5 273.8 207.3 274.6 ;
      RECT  200.5 279.0 207.3 279.8 ;
      RECT  200.5 294.6 207.3 295.4 ;
      RECT  200.5 299.8 207.3 300.6 ;
      RECT  200.5 315.4 207.3 316.2 ;
      RECT  200.5 320.6 207.3 321.4 ;
      RECT  200.5 336.2 207.3 337.0 ;
      RECT  200.5 341.4 207.3 342.2 ;
      RECT  200.5 357.0 207.3 357.8 ;
      RECT  200.5 362.2 207.3 363.0 ;
      RECT  173.3 195.8 207.3 196.6 ;
      RECT  173.3 211.4 207.3 212.2 ;
      RECT  173.3 216.6 207.3 217.4 ;
      RECT  173.3 232.2 207.3 233.0 ;
      RECT  173.3 237.4 207.3 238.2 ;
      RECT  173.3 253.0 207.3 253.8 ;
      RECT  173.3 258.2 207.3 259.0 ;
      RECT  173.3 273.8 207.3 274.6 ;
      RECT  173.3 279.0 207.3 279.8 ;
      RECT  173.3 294.6 207.3 295.4 ;
      RECT  173.3 299.8 207.3 300.6 ;
      RECT  173.3 315.4 207.3 316.2 ;
      RECT  173.3 320.6 207.3 321.4 ;
      RECT  173.3 336.2 207.3 337.0 ;
      RECT  173.3 341.4 207.3 342.2 ;
      RECT  173.3 357.0 207.3 357.8 ;
      RECT  173.3 190.6 207.3 191.4 ;
      RECT  183.6 159.6 184.4 160.4 ;
      RECT  181.6 159.6 182.4 160.4 ;
      RECT  183.6 164.0 184.4 164.8 ;
      RECT  181.6 164.0 182.4 164.8 ;
      RECT  185.6 164.0 186.4 164.8 ;
      RECT  183.6 164.0 184.4 164.8 ;
      RECT  180.1 157.5 186.9 158.1 ;
      RECT  190.4 159.6 191.2 160.4 ;
      RECT  188.4 159.6 189.2 160.4 ;
      RECT  190.4 164.0 191.2 164.8 ;
      RECT  188.4 164.0 189.2 164.8 ;
      RECT  192.4 164.0 193.2 164.8 ;
      RECT  190.4 164.0 191.2 164.8 ;
      RECT  186.9 157.5 193.7 158.1 ;
      RECT  197.2 159.6 198.0 160.4 ;
      RECT  195.2 159.6 196.0 160.4 ;
      RECT  197.2 164.0 198.0 164.8 ;
      RECT  195.2 164.0 196.0 164.8 ;
      RECT  199.2 164.0 200.0 164.8 ;
      RECT  197.2 164.0 198.0 164.8 ;
      RECT  193.7 157.5 200.5 158.1 ;
      RECT  180.1 157.5 200.5 158.1 ;
      RECT  189.7 123.8 190.5 128.6 ;
      RECT  192.3 133.0 193.1 134.2 ;
      RECT  191.5 140.8 192.3 143.2 ;
      RECT  189.9 141.4 190.7 143.2 ;
      RECT  193.3 147.2 194.1 148.0 ;
      RECT  188.1 124.4 188.9 128.6 ;
      RECT  189.9 134.2 193.1 134.8 ;
      RECT  188.3 133.6 189.1 143.2 ;
      RECT  193.1 128.6 193.7 130.0 ;
      RECT  186.5 149.6 194.1 150.4 ;
      RECT  188.3 132.8 189.5 133.6 ;
      RECT  188.1 130.0 189.5 130.6 ;
      RECT  188.7 130.6 189.5 130.8 ;
      RECT  191.7 147.2 192.5 147.6 ;
      RECT  191.3 123.8 192.1 129.4 ;
      RECT  189.5 128.6 190.3 129.4 ;
      RECT  188.1 128.6 188.7 130.0 ;
      RECT  190.1 143.2 190.7 145.8 ;
      RECT  192.9 123.8 193.7 128.6 ;
      RECT  190.1 145.8 190.9 147.6 ;
      RECT  187.5 122.0 188.3 123.8 ;
      RECT  191.5 135.4 192.3 140.0 ;
      RECT  187.5 123.8 188.9 124.4 ;
      RECT  192.7 130.0 193.7 130.8 ;
      RECT  189.9 135.4 190.7 139.0 ;
      RECT  191.7 146.4 194.1 147.2 ;
      RECT  189.9 134.8 190.5 135.4 ;
      RECT  191.5 140.0 192.9 140.8 ;
      RECT  191.7 145.8 192.5 146.4 ;
      RECT  196.5 123.8 197.3 128.6 ;
      RECT  199.1 133.0 199.9 134.2 ;
      RECT  198.3 140.8 199.1 143.2 ;
      RECT  196.7 141.4 197.5 143.2 ;
      RECT  200.1 147.2 200.9 148.0 ;
      RECT  194.9 124.4 195.7 128.6 ;
      RECT  196.7 134.2 199.9 134.8 ;
      RECT  195.1 133.6 195.9 143.2 ;
      RECT  199.9 128.6 200.5 130.0 ;
      RECT  193.3 149.6 200.9 150.4 ;
      RECT  195.1 132.8 196.3 133.6 ;
      RECT  194.9 130.0 196.3 130.6 ;
      RECT  195.5 130.6 196.3 130.8 ;
      RECT  198.5 147.2 199.3 147.6 ;
      RECT  198.1 123.8 198.9 129.4 ;
      RECT  196.3 128.6 197.1 129.4 ;
      RECT  194.9 128.6 195.5 130.0 ;
      RECT  196.9 143.2 197.5 145.8 ;
      RECT  199.7 123.8 200.5 128.6 ;
      RECT  196.9 145.8 197.7 147.6 ;
      RECT  194.3 122.0 195.1 123.8 ;
      RECT  198.3 135.4 199.1 140.0 ;
      RECT  194.3 123.8 195.7 124.4 ;
      RECT  199.5 130.0 200.5 130.8 ;
      RECT  196.7 135.4 197.5 139.0 ;
      RECT  198.5 146.4 200.9 147.2 ;
      RECT  196.7 134.8 197.3 135.4 ;
      RECT  198.3 140.0 199.7 140.8 ;
      RECT  198.5 145.8 199.3 146.4 ;
      RECT  186.9 149.6 200.5 150.2 ;
      RECT  187.9 91.4 188.7 95.2 ;
      RECT  191.1 94.2 192.3 95.0 ;
      RECT  187.5 79.8 193.1 80.6 ;
      RECT  187.9 113.6 189.7 114.4 ;
      RECT  187.5 82.0 188.3 84.0 ;
      RECT  190.9 100.0 191.7 102.6 ;
      RECT  189.5 96.4 190.3 98.6 ;
      RECT  187.5 81.2 191.5 82.0 ;
      RECT  189.5 91.4 190.3 92.8 ;
      RECT  187.9 95.8 188.7 97.8 ;
      RECT  189.1 82.6 189.9 84.6 ;
      RECT  187.5 85.2 188.3 87.8 ;
      RECT  190.9 103.4 191.7 104.6 ;
      RECT  187.7 100.0 188.5 108.6 ;
      RECT  187.9 95.2 191.9 95.8 ;
      RECT  189.3 98.6 190.9 99.4 ;
      RECT  190.7 82.0 191.5 84.0 ;
      RECT  191.1 95.8 191.9 97.8 ;
      RECT  189.1 86.4 189.9 87.8 ;
      RECT  191.1 95.0 191.9 95.2 ;
      RECT  190.9 110.6 191.7 113.8 ;
      RECT  189.3 99.4 190.1 101.4 ;
      RECT  190.9 102.6 193.5 103.4 ;
      RECT  187.5 89.2 188.3 90.0 ;
      RECT  191.9 92.8 192.9 93.0 ;
      RECT  187.9 113.0 188.5 113.6 ;
      RECT  189.3 103.8 190.1 113.0 ;
      RECT  187.7 110.6 188.5 113.0 ;
      RECT  187.5 84.6 189.9 85.2 ;
      RECT  192.5 111.4 193.5 112.2 ;
      RECT  187.7 87.8 188.3 89.2 ;
      RECT  189.9 76.2 190.7 77.8 ;
      RECT  190.7 86.4 191.5 88.6 ;
      RECT  192.9 103.4 193.5 111.4 ;
      RECT  191.5 90.0 193.1 90.8 ;
      RECT  191.1 91.4 192.9 92.8 ;
      RECT  192.3 82.6 193.1 90.0 ;
      RECT  194.7 91.4 195.5 95.2 ;
      RECT  197.9 94.2 199.1 95.0 ;
      RECT  194.3 79.8 199.9 80.6 ;
      RECT  194.7 113.6 196.5 114.4 ;
      RECT  194.3 82.0 195.1 84.0 ;
      RECT  197.7 100.0 198.5 102.6 ;
      RECT  196.3 96.4 197.1 98.6 ;
      RECT  194.3 81.2 198.3 82.0 ;
      RECT  196.3 91.4 197.1 92.8 ;
      RECT  194.7 95.8 195.5 97.8 ;
      RECT  195.9 82.6 196.7 84.6 ;
      RECT  194.3 85.2 195.1 87.8 ;
      RECT  197.7 103.4 198.5 104.6 ;
      RECT  194.5 100.0 195.3 108.6 ;
      RECT  194.7 95.2 198.7 95.8 ;
      RECT  196.1 98.6 197.7 99.4 ;
      RECT  197.5 82.0 198.3 84.0 ;
      RECT  197.9 95.8 198.7 97.8 ;
      RECT  195.9 86.4 196.7 87.8 ;
      RECT  197.9 95.0 198.7 95.2 ;
      RECT  197.7 110.6 198.5 113.8 ;
      RECT  196.1 99.4 196.9 101.4 ;
      RECT  197.7 102.6 200.3 103.4 ;
      RECT  194.3 89.2 195.1 90.0 ;
      RECT  198.7 92.8 199.7 93.0 ;
      RECT  194.7 113.0 195.3 113.6 ;
      RECT  196.1 103.8 196.9 113.0 ;
      RECT  194.5 110.6 195.3 113.0 ;
      RECT  194.3 84.6 196.7 85.2 ;
      RECT  199.3 111.4 200.3 112.2 ;
      RECT  194.5 87.8 195.1 89.2 ;
      RECT  196.7 76.2 197.5 77.8 ;
      RECT  197.5 86.4 198.3 88.6 ;
      RECT  199.7 103.4 200.3 111.4 ;
      RECT  198.3 90.0 199.9 90.8 ;
      RECT  197.9 91.4 199.7 92.8 ;
      RECT  199.1 82.6 199.9 90.0 ;
      RECT  186.9 79.8 200.5 80.4 ;
      RECT  186.9 150.2 200.5 149.6 ;
      RECT  180.1 158.1 200.5 157.5 ;
      RECT  186.9 80.4 200.5 79.8 ;
      RECT  97.3 202.3 98.1 203.1 ;
      RECT  95.3 202.3 96.1 203.1 ;
      RECT  97.3 194.9 98.1 195.7 ;
      RECT  95.3 194.9 96.1 195.7 ;
      RECT  95.7 198.6 96.5 199.4 ;
      RECT  97.7 198.7 98.3 199.3 ;
      RECT  94.1 204.1 100.7 204.7 ;
      RECT  94.1 193.7 100.7 194.3 ;
      RECT  97.3 206.5 98.1 205.7 ;
      RECT  95.3 206.5 96.1 205.7 ;
      RECT  97.3 213.9 98.1 213.1 ;
      RECT  95.3 213.9 96.1 213.1 ;
      RECT  95.7 210.2 96.5 209.4 ;
      RECT  97.7 210.1 98.3 209.5 ;
      RECT  94.1 204.7 100.7 204.1 ;
      RECT  94.1 215.1 100.7 214.5 ;
      RECT  112.3 202.3 113.1 203.1 ;
      RECT  110.3 202.3 111.1 203.1 ;
      RECT  114.3 202.3 115.1 203.1 ;
      RECT  112.3 202.3 113.1 203.1 ;
      RECT  110.3 195.3 111.1 196.1 ;
      RECT  114.3 195.3 115.1 196.1 ;
      RECT  111.3 196.8 112.1 197.6 ;
      RECT  113.3 199.6 114.1 200.4 ;
      RECT  115.8 201.0 116.4 201.6 ;
      RECT  109.1 204.1 117.7 204.7 ;
      RECT  109.1 193.7 117.7 194.3 ;
      RECT  120.9 202.3 121.7 203.1 ;
      RECT  118.9 202.3 119.7 203.1 ;
      RECT  120.9 194.9 121.7 195.7 ;
      RECT  118.9 194.9 119.7 195.7 ;
      RECT  119.3 198.6 120.1 199.4 ;
      RECT  121.3 198.7 121.9 199.3 ;
      RECT  117.7 204.1 124.3 204.7 ;
      RECT  117.7 193.7 124.3 194.3 ;
      RECT  111.3 196.8 112.1 197.6 ;
      RECT  113.3 199.6 114.1 200.4 ;
      RECT  121.3 198.7 121.9 199.3 ;
      RECT  109.1 204.1 124.3 204.7 ;
      RECT  109.1 193.7 124.3 194.3 ;
      RECT  112.3 206.5 113.1 205.7 ;
      RECT  110.3 206.5 111.1 205.7 ;
      RECT  114.3 206.5 115.1 205.7 ;
      RECT  112.3 206.5 113.1 205.7 ;
      RECT  110.3 213.5 111.1 212.7 ;
      RECT  114.3 213.5 115.1 212.7 ;
      RECT  111.3 212.0 112.1 211.2 ;
      RECT  113.3 209.2 114.1 208.4 ;
      RECT  115.8 207.8 116.4 207.2 ;
      RECT  109.1 204.7 117.7 204.1 ;
      RECT  109.1 215.1 117.7 214.5 ;
      RECT  120.9 206.5 121.7 205.7 ;
      RECT  118.9 206.5 119.7 205.7 ;
      RECT  120.9 213.9 121.7 213.1 ;
      RECT  118.9 213.9 119.7 213.1 ;
      RECT  119.3 210.2 120.1 209.4 ;
      RECT  121.3 210.1 121.9 209.5 ;
      RECT  117.7 204.7 124.3 204.1 ;
      RECT  117.7 215.1 124.3 214.5 ;
      RECT  111.3 212.0 112.1 211.2 ;
      RECT  113.3 209.2 114.1 208.4 ;
      RECT  121.3 210.1 121.9 209.5 ;
      RECT  109.1 204.7 124.3 204.1 ;
      RECT  109.1 215.1 124.3 214.5 ;
      RECT  112.3 223.1 113.1 223.9 ;
      RECT  110.3 223.1 111.1 223.9 ;
      RECT  114.3 223.1 115.1 223.9 ;
      RECT  112.3 223.1 113.1 223.9 ;
      RECT  110.3 216.1 111.1 216.9 ;
      RECT  114.3 216.1 115.1 216.9 ;
      RECT  111.3 217.6 112.1 218.4 ;
      RECT  113.3 220.4 114.1 221.2 ;
      RECT  115.8 221.8 116.4 222.4 ;
      RECT  109.1 224.9 117.7 225.5 ;
      RECT  109.1 214.5 117.7 215.1 ;
      RECT  120.9 223.1 121.7 223.9 ;
      RECT  118.9 223.1 119.7 223.9 ;
      RECT  120.9 215.7 121.7 216.5 ;
      RECT  118.9 215.7 119.7 216.5 ;
      RECT  119.3 219.4 120.1 220.2 ;
      RECT  121.3 219.5 121.9 220.1 ;
      RECT  117.7 224.9 124.3 225.5 ;
      RECT  117.7 214.5 124.3 215.1 ;
      RECT  111.3 217.6 112.1 218.4 ;
      RECT  113.3 220.4 114.1 221.2 ;
      RECT  121.3 219.5 121.9 220.1 ;
      RECT  109.1 224.9 124.3 225.5 ;
      RECT  109.1 214.5 124.3 215.1 ;
      RECT  112.3 227.3 113.1 226.5 ;
      RECT  110.3 227.3 111.1 226.5 ;
      RECT  114.3 227.3 115.1 226.5 ;
      RECT  112.3 227.3 113.1 226.5 ;
      RECT  110.3 234.3 111.1 233.5 ;
      RECT  114.3 234.3 115.1 233.5 ;
      RECT  111.3 232.8 112.1 232.0 ;
      RECT  113.3 230.0 114.1 229.2 ;
      RECT  115.8 228.6 116.4 228.0 ;
      RECT  109.1 225.5 117.7 224.9 ;
      RECT  109.1 235.9 117.7 235.3 ;
      RECT  120.9 227.3 121.7 226.5 ;
      RECT  118.9 227.3 119.7 226.5 ;
      RECT  120.9 234.7 121.7 233.9 ;
      RECT  118.9 234.7 119.7 233.9 ;
      RECT  119.3 231.0 120.1 230.2 ;
      RECT  121.3 230.9 121.9 230.3 ;
      RECT  117.7 225.5 124.3 224.9 ;
      RECT  117.7 235.9 124.3 235.3 ;
      RECT  111.3 232.8 112.1 232.0 ;
      RECT  113.3 230.0 114.1 229.2 ;
      RECT  121.3 230.9 121.9 230.3 ;
      RECT  109.1 225.5 124.3 224.9 ;
      RECT  109.1 235.9 124.3 235.3 ;
      RECT  121.3 198.7 121.9 199.3 ;
      RECT  121.3 209.5 121.9 210.1 ;
      RECT  121.3 219.5 121.9 220.1 ;
      RECT  121.3 230.3 121.9 230.9 ;
      RECT  97.3 254.3 98.1 255.1 ;
      RECT  95.3 254.3 96.1 255.1 ;
      RECT  97.3 246.9 98.1 247.7 ;
      RECT  95.3 246.9 96.1 247.7 ;
      RECT  95.7 250.6 96.5 251.4 ;
      RECT  97.7 250.7 98.3 251.3 ;
      RECT  94.1 256.1 100.7 256.7 ;
      RECT  94.1 245.7 100.7 246.3 ;
      RECT  97.3 258.5 98.1 257.7 ;
      RECT  95.3 258.5 96.1 257.7 ;
      RECT  97.3 265.9 98.1 265.1 ;
      RECT  95.3 265.9 96.1 265.1 ;
      RECT  95.7 262.2 96.5 261.4 ;
      RECT  97.7 262.1 98.3 261.5 ;
      RECT  94.1 256.7 100.7 256.1 ;
      RECT  94.1 267.1 100.7 266.5 ;
      RECT  112.3 254.3 113.1 255.1 ;
      RECT  110.3 254.3 111.1 255.1 ;
      RECT  114.3 254.3 115.1 255.1 ;
      RECT  112.3 254.3 113.1 255.1 ;
      RECT  110.3 247.3 111.1 248.1 ;
      RECT  114.3 247.3 115.1 248.1 ;
      RECT  111.3 248.8 112.1 249.6 ;
      RECT  113.3 251.6 114.1 252.4 ;
      RECT  115.8 253.0 116.4 253.6 ;
      RECT  109.1 256.1 117.7 256.7 ;
      RECT  109.1 245.7 117.7 246.3 ;
      RECT  120.9 254.3 121.7 255.1 ;
      RECT  118.9 254.3 119.7 255.1 ;
      RECT  120.9 246.9 121.7 247.7 ;
      RECT  118.9 246.9 119.7 247.7 ;
      RECT  119.3 250.6 120.1 251.4 ;
      RECT  121.3 250.7 121.9 251.3 ;
      RECT  117.7 256.1 124.3 256.7 ;
      RECT  117.7 245.7 124.3 246.3 ;
      RECT  111.3 248.8 112.1 249.6 ;
      RECT  113.3 251.6 114.1 252.4 ;
      RECT  121.3 250.7 121.9 251.3 ;
      RECT  109.1 256.1 124.3 256.7 ;
      RECT  109.1 245.7 124.3 246.3 ;
      RECT  112.3 258.5 113.1 257.7 ;
      RECT  110.3 258.5 111.1 257.7 ;
      RECT  114.3 258.5 115.1 257.7 ;
      RECT  112.3 258.5 113.1 257.7 ;
      RECT  110.3 265.5 111.1 264.7 ;
      RECT  114.3 265.5 115.1 264.7 ;
      RECT  111.3 264.0 112.1 263.2 ;
      RECT  113.3 261.2 114.1 260.4 ;
      RECT  115.8 259.8 116.4 259.2 ;
      RECT  109.1 256.7 117.7 256.1 ;
      RECT  109.1 267.1 117.7 266.5 ;
      RECT  120.9 258.5 121.7 257.7 ;
      RECT  118.9 258.5 119.7 257.7 ;
      RECT  120.9 265.9 121.7 265.1 ;
      RECT  118.9 265.9 119.7 265.1 ;
      RECT  119.3 262.2 120.1 261.4 ;
      RECT  121.3 262.1 121.9 261.5 ;
      RECT  117.7 256.7 124.3 256.1 ;
      RECT  117.7 267.1 124.3 266.5 ;
      RECT  111.3 264.0 112.1 263.2 ;
      RECT  113.3 261.2 114.1 260.4 ;
      RECT  121.3 262.1 121.9 261.5 ;
      RECT  109.1 256.7 124.3 256.1 ;
      RECT  109.1 267.1 124.3 266.5 ;
      RECT  112.3 275.1 113.1 275.9 ;
      RECT  110.3 275.1 111.1 275.9 ;
      RECT  114.3 275.1 115.1 275.9 ;
      RECT  112.3 275.1 113.1 275.9 ;
      RECT  110.3 268.1 111.1 268.9 ;
      RECT  114.3 268.1 115.1 268.9 ;
      RECT  111.3 269.6 112.1 270.4 ;
      RECT  113.3 272.4 114.1 273.2 ;
      RECT  115.8 273.8 116.4 274.4 ;
      RECT  109.1 276.9 117.7 277.5 ;
      RECT  109.1 266.5 117.7 267.1 ;
      RECT  120.9 275.1 121.7 275.9 ;
      RECT  118.9 275.1 119.7 275.9 ;
      RECT  120.9 267.7 121.7 268.5 ;
      RECT  118.9 267.7 119.7 268.5 ;
      RECT  119.3 271.4 120.1 272.2 ;
      RECT  121.3 271.5 121.9 272.1 ;
      RECT  117.7 276.9 124.3 277.5 ;
      RECT  117.7 266.5 124.3 267.1 ;
      RECT  111.3 269.6 112.1 270.4 ;
      RECT  113.3 272.4 114.1 273.2 ;
      RECT  121.3 271.5 121.9 272.1 ;
      RECT  109.1 276.9 124.3 277.5 ;
      RECT  109.1 266.5 124.3 267.1 ;
      RECT  112.3 279.3 113.1 278.5 ;
      RECT  110.3 279.3 111.1 278.5 ;
      RECT  114.3 279.3 115.1 278.5 ;
      RECT  112.3 279.3 113.1 278.5 ;
      RECT  110.3 286.3 111.1 285.5 ;
      RECT  114.3 286.3 115.1 285.5 ;
      RECT  111.3 284.8 112.1 284.0 ;
      RECT  113.3 282.0 114.1 281.2 ;
      RECT  115.8 280.6 116.4 280.0 ;
      RECT  109.1 277.5 117.7 276.9 ;
      RECT  109.1 287.9 117.7 287.3 ;
      RECT  120.9 279.3 121.7 278.5 ;
      RECT  118.9 279.3 119.7 278.5 ;
      RECT  120.9 286.7 121.7 285.9 ;
      RECT  118.9 286.7 119.7 285.9 ;
      RECT  119.3 283.0 120.1 282.2 ;
      RECT  121.3 282.9 121.9 282.3 ;
      RECT  117.7 277.5 124.3 276.9 ;
      RECT  117.7 287.9 124.3 287.3 ;
      RECT  111.3 284.8 112.1 284.0 ;
      RECT  113.3 282.0 114.1 281.2 ;
      RECT  121.3 282.9 121.9 282.3 ;
      RECT  109.1 277.5 124.3 276.9 ;
      RECT  109.1 287.9 124.3 287.3 ;
      RECT  121.3 250.7 121.9 251.3 ;
      RECT  121.3 261.5 121.9 262.1 ;
      RECT  121.3 271.5 121.9 272.1 ;
      RECT  121.3 282.3 121.9 282.9 ;
      RECT  140.1 202.3 140.9 203.1 ;
      RECT  138.1 202.3 138.9 203.1 ;
      RECT  142.1 202.3 142.9 203.1 ;
      RECT  140.1 202.3 140.9 203.1 ;
      RECT  138.1 195.3 138.9 196.1 ;
      RECT  142.1 195.3 142.9 196.1 ;
      RECT  139.1 196.8 139.9 197.6 ;
      RECT  141.1 199.6 141.9 200.4 ;
      RECT  143.6 201.0 144.2 201.6 ;
      RECT  136.9 204.1 145.5 204.7 ;
      RECT  136.9 193.7 145.5 194.3 ;
      RECT  148.7 202.3 149.5 203.1 ;
      RECT  146.7 202.3 147.5 203.1 ;
      RECT  148.7 194.9 149.5 195.7 ;
      RECT  146.7 194.9 147.5 195.7 ;
      RECT  147.1 198.6 147.9 199.4 ;
      RECT  149.1 198.7 149.7 199.3 ;
      RECT  145.5 204.1 152.1 204.7 ;
      RECT  145.5 193.7 152.1 194.3 ;
      RECT  139.1 196.8 139.9 197.6 ;
      RECT  141.1 199.6 141.9 200.4 ;
      RECT  149.1 198.7 149.7 199.3 ;
      RECT  136.9 204.1 152.1 204.7 ;
      RECT  136.9 193.7 152.1 194.3 ;
      RECT  140.1 206.5 140.9 205.7 ;
      RECT  138.1 206.5 138.9 205.7 ;
      RECT  142.1 206.5 142.9 205.7 ;
      RECT  140.1 206.5 140.9 205.7 ;
      RECT  138.1 213.5 138.9 212.7 ;
      RECT  142.1 213.5 142.9 212.7 ;
      RECT  139.1 212.0 139.9 211.2 ;
      RECT  141.1 209.2 141.9 208.4 ;
      RECT  143.6 207.8 144.2 207.2 ;
      RECT  136.9 204.7 145.5 204.1 ;
      RECT  136.9 215.1 145.5 214.5 ;
      RECT  148.7 206.5 149.5 205.7 ;
      RECT  146.7 206.5 147.5 205.7 ;
      RECT  148.7 213.9 149.5 213.1 ;
      RECT  146.7 213.9 147.5 213.1 ;
      RECT  147.1 210.2 147.9 209.4 ;
      RECT  149.1 210.1 149.7 209.5 ;
      RECT  145.5 204.7 152.1 204.1 ;
      RECT  145.5 215.1 152.1 214.5 ;
      RECT  139.1 212.0 139.9 211.2 ;
      RECT  141.1 209.2 141.9 208.4 ;
      RECT  149.1 210.1 149.7 209.5 ;
      RECT  136.9 204.7 152.1 204.1 ;
      RECT  136.9 215.1 152.1 214.5 ;
      RECT  140.1 223.1 140.9 223.9 ;
      RECT  138.1 223.1 138.9 223.9 ;
      RECT  142.1 223.1 142.9 223.9 ;
      RECT  140.1 223.1 140.9 223.9 ;
      RECT  138.1 216.1 138.9 216.9 ;
      RECT  142.1 216.1 142.9 216.9 ;
      RECT  139.1 217.6 139.9 218.4 ;
      RECT  141.1 220.4 141.9 221.2 ;
      RECT  143.6 221.8 144.2 222.4 ;
      RECT  136.9 224.9 145.5 225.5 ;
      RECT  136.9 214.5 145.5 215.1 ;
      RECT  148.7 223.1 149.5 223.9 ;
      RECT  146.7 223.1 147.5 223.9 ;
      RECT  148.7 215.7 149.5 216.5 ;
      RECT  146.7 215.7 147.5 216.5 ;
      RECT  147.1 219.4 147.9 220.2 ;
      RECT  149.1 219.5 149.7 220.1 ;
      RECT  145.5 224.9 152.1 225.5 ;
      RECT  145.5 214.5 152.1 215.1 ;
      RECT  139.1 217.6 139.9 218.4 ;
      RECT  141.1 220.4 141.9 221.2 ;
      RECT  149.1 219.5 149.7 220.1 ;
      RECT  136.9 224.9 152.1 225.5 ;
      RECT  136.9 214.5 152.1 215.1 ;
      RECT  140.1 227.3 140.9 226.5 ;
      RECT  138.1 227.3 138.9 226.5 ;
      RECT  142.1 227.3 142.9 226.5 ;
      RECT  140.1 227.3 140.9 226.5 ;
      RECT  138.1 234.3 138.9 233.5 ;
      RECT  142.1 234.3 142.9 233.5 ;
      RECT  139.1 232.8 139.9 232.0 ;
      RECT  141.1 230.0 141.9 229.2 ;
      RECT  143.6 228.6 144.2 228.0 ;
      RECT  136.9 225.5 145.5 224.9 ;
      RECT  136.9 235.9 145.5 235.3 ;
      RECT  148.7 227.3 149.5 226.5 ;
      RECT  146.7 227.3 147.5 226.5 ;
      RECT  148.7 234.7 149.5 233.9 ;
      RECT  146.7 234.7 147.5 233.9 ;
      RECT  147.1 231.0 147.9 230.2 ;
      RECT  149.1 230.9 149.7 230.3 ;
      RECT  145.5 225.5 152.1 224.9 ;
      RECT  145.5 235.9 152.1 235.3 ;
      RECT  139.1 232.8 139.9 232.0 ;
      RECT  141.1 230.0 141.9 229.2 ;
      RECT  149.1 230.9 149.7 230.3 ;
      RECT  136.9 225.5 152.1 224.9 ;
      RECT  136.9 235.9 152.1 235.3 ;
      RECT  140.1 243.9 140.9 244.7 ;
      RECT  138.1 243.9 138.9 244.7 ;
      RECT  142.1 243.9 142.9 244.7 ;
      RECT  140.1 243.9 140.9 244.7 ;
      RECT  138.1 236.9 138.9 237.7 ;
      RECT  142.1 236.9 142.9 237.7 ;
      RECT  139.1 238.4 139.9 239.2 ;
      RECT  141.1 241.2 141.9 242.0 ;
      RECT  143.6 242.6 144.2 243.2 ;
      RECT  136.9 245.7 145.5 246.3 ;
      RECT  136.9 235.3 145.5 235.9 ;
      RECT  148.7 243.9 149.5 244.7 ;
      RECT  146.7 243.9 147.5 244.7 ;
      RECT  148.7 236.5 149.5 237.3 ;
      RECT  146.7 236.5 147.5 237.3 ;
      RECT  147.1 240.2 147.9 241.0 ;
      RECT  149.1 240.3 149.7 240.9 ;
      RECT  145.5 245.7 152.1 246.3 ;
      RECT  145.5 235.3 152.1 235.9 ;
      RECT  139.1 238.4 139.9 239.2 ;
      RECT  141.1 241.2 141.9 242.0 ;
      RECT  149.1 240.3 149.7 240.9 ;
      RECT  136.9 245.7 152.1 246.3 ;
      RECT  136.9 235.3 152.1 235.9 ;
      RECT  140.1 248.1 140.9 247.3 ;
      RECT  138.1 248.1 138.9 247.3 ;
      RECT  142.1 248.1 142.9 247.3 ;
      RECT  140.1 248.1 140.9 247.3 ;
      RECT  138.1 255.1 138.9 254.3 ;
      RECT  142.1 255.1 142.9 254.3 ;
      RECT  139.1 253.6 139.9 252.8 ;
      RECT  141.1 250.8 141.9 250.0 ;
      RECT  143.6 249.4 144.2 248.8 ;
      RECT  136.9 246.3 145.5 245.7 ;
      RECT  136.9 256.7 145.5 256.1 ;
      RECT  148.7 248.1 149.5 247.3 ;
      RECT  146.7 248.1 147.5 247.3 ;
      RECT  148.7 255.5 149.5 254.7 ;
      RECT  146.7 255.5 147.5 254.7 ;
      RECT  147.1 251.8 147.9 251.0 ;
      RECT  149.1 251.7 149.7 251.1 ;
      RECT  145.5 246.3 152.1 245.7 ;
      RECT  145.5 256.7 152.1 256.1 ;
      RECT  139.1 253.6 139.9 252.8 ;
      RECT  141.1 250.8 141.9 250.0 ;
      RECT  149.1 251.7 149.7 251.1 ;
      RECT  136.9 246.3 152.1 245.7 ;
      RECT  136.9 256.7 152.1 256.1 ;
      RECT  140.1 264.7 140.9 265.5 ;
      RECT  138.1 264.7 138.9 265.5 ;
      RECT  142.1 264.7 142.9 265.5 ;
      RECT  140.1 264.7 140.9 265.5 ;
      RECT  138.1 257.7 138.9 258.5 ;
      RECT  142.1 257.7 142.9 258.5 ;
      RECT  139.1 259.2 139.9 260.0 ;
      RECT  141.1 262.0 141.9 262.8 ;
      RECT  143.6 263.4 144.2 264.0 ;
      RECT  136.9 266.5 145.5 267.1 ;
      RECT  136.9 256.1 145.5 256.7 ;
      RECT  148.7 264.7 149.5 265.5 ;
      RECT  146.7 264.7 147.5 265.5 ;
      RECT  148.7 257.3 149.5 258.1 ;
      RECT  146.7 257.3 147.5 258.1 ;
      RECT  147.1 261.0 147.9 261.8 ;
      RECT  149.1 261.1 149.7 261.7 ;
      RECT  145.5 266.5 152.1 267.1 ;
      RECT  145.5 256.1 152.1 256.7 ;
      RECT  139.1 259.2 139.9 260.0 ;
      RECT  141.1 262.0 141.9 262.8 ;
      RECT  149.1 261.1 149.7 261.7 ;
      RECT  136.9 266.5 152.1 267.1 ;
      RECT  136.9 256.1 152.1 256.7 ;
      RECT  140.1 268.9 140.9 268.1 ;
      RECT  138.1 268.9 138.9 268.1 ;
      RECT  142.1 268.9 142.9 268.1 ;
      RECT  140.1 268.9 140.9 268.1 ;
      RECT  138.1 275.9 138.9 275.1 ;
      RECT  142.1 275.9 142.9 275.1 ;
      RECT  139.1 274.4 139.9 273.6 ;
      RECT  141.1 271.6 141.9 270.8 ;
      RECT  143.6 270.2 144.2 269.6 ;
      RECT  136.9 267.1 145.5 266.5 ;
      RECT  136.9 277.5 145.5 276.9 ;
      RECT  148.7 268.9 149.5 268.1 ;
      RECT  146.7 268.9 147.5 268.1 ;
      RECT  148.7 276.3 149.5 275.5 ;
      RECT  146.7 276.3 147.5 275.5 ;
      RECT  147.1 272.6 147.9 271.8 ;
      RECT  149.1 272.5 149.7 271.9 ;
      RECT  145.5 267.1 152.1 266.5 ;
      RECT  145.5 277.5 152.1 276.9 ;
      RECT  139.1 274.4 139.9 273.6 ;
      RECT  141.1 271.6 141.9 270.8 ;
      RECT  149.1 272.5 149.7 271.9 ;
      RECT  136.9 267.1 152.1 266.5 ;
      RECT  136.9 277.5 152.1 276.9 ;
      RECT  140.1 285.5 140.9 286.3 ;
      RECT  138.1 285.5 138.9 286.3 ;
      RECT  142.1 285.5 142.9 286.3 ;
      RECT  140.1 285.5 140.9 286.3 ;
      RECT  138.1 278.5 138.9 279.3 ;
      RECT  142.1 278.5 142.9 279.3 ;
      RECT  139.1 280.0 139.9 280.8 ;
      RECT  141.1 282.8 141.9 283.6 ;
      RECT  143.6 284.2 144.2 284.8 ;
      RECT  136.9 287.3 145.5 287.9 ;
      RECT  136.9 276.9 145.5 277.5 ;
      RECT  148.7 285.5 149.5 286.3 ;
      RECT  146.7 285.5 147.5 286.3 ;
      RECT  148.7 278.1 149.5 278.9 ;
      RECT  146.7 278.1 147.5 278.9 ;
      RECT  147.1 281.8 147.9 282.6 ;
      RECT  149.1 281.9 149.7 282.5 ;
      RECT  145.5 287.3 152.1 287.9 ;
      RECT  145.5 276.9 152.1 277.5 ;
      RECT  139.1 280.0 139.9 280.8 ;
      RECT  141.1 282.8 141.9 283.6 ;
      RECT  149.1 281.9 149.7 282.5 ;
      RECT  136.9 287.3 152.1 287.9 ;
      RECT  136.9 276.9 152.1 277.5 ;
      RECT  140.1 289.7 140.9 288.9 ;
      RECT  138.1 289.7 138.9 288.9 ;
      RECT  142.1 289.7 142.9 288.9 ;
      RECT  140.1 289.7 140.9 288.9 ;
      RECT  138.1 296.7 138.9 295.9 ;
      RECT  142.1 296.7 142.9 295.9 ;
      RECT  139.1 295.2 139.9 294.4 ;
      RECT  141.1 292.4 141.9 291.6 ;
      RECT  143.6 291.0 144.2 290.4 ;
      RECT  136.9 287.9 145.5 287.3 ;
      RECT  136.9 298.3 145.5 297.7 ;
      RECT  148.7 289.7 149.5 288.9 ;
      RECT  146.7 289.7 147.5 288.9 ;
      RECT  148.7 297.1 149.5 296.3 ;
      RECT  146.7 297.1 147.5 296.3 ;
      RECT  147.1 293.4 147.9 292.6 ;
      RECT  149.1 293.3 149.7 292.7 ;
      RECT  145.5 287.9 152.1 287.3 ;
      RECT  145.5 298.3 152.1 297.7 ;
      RECT  139.1 295.2 139.9 294.4 ;
      RECT  141.1 292.4 141.9 291.6 ;
      RECT  149.1 293.3 149.7 292.7 ;
      RECT  136.9 287.9 152.1 287.3 ;
      RECT  136.9 298.3 152.1 297.7 ;
      RECT  140.1 306.3 140.9 307.1 ;
      RECT  138.1 306.3 138.9 307.1 ;
      RECT  142.1 306.3 142.9 307.1 ;
      RECT  140.1 306.3 140.9 307.1 ;
      RECT  138.1 299.3 138.9 300.1 ;
      RECT  142.1 299.3 142.9 300.1 ;
      RECT  139.1 300.8 139.9 301.6 ;
      RECT  141.1 303.6 141.9 304.4 ;
      RECT  143.6 305.0 144.2 305.6 ;
      RECT  136.9 308.1 145.5 308.7 ;
      RECT  136.9 297.7 145.5 298.3 ;
      RECT  148.7 306.3 149.5 307.1 ;
      RECT  146.7 306.3 147.5 307.1 ;
      RECT  148.7 298.9 149.5 299.7 ;
      RECT  146.7 298.9 147.5 299.7 ;
      RECT  147.1 302.6 147.9 303.4 ;
      RECT  149.1 302.7 149.7 303.3 ;
      RECT  145.5 308.1 152.1 308.7 ;
      RECT  145.5 297.7 152.1 298.3 ;
      RECT  139.1 300.8 139.9 301.6 ;
      RECT  141.1 303.6 141.9 304.4 ;
      RECT  149.1 302.7 149.7 303.3 ;
      RECT  136.9 308.1 152.1 308.7 ;
      RECT  136.9 297.7 152.1 298.3 ;
      RECT  140.1 310.5 140.9 309.7 ;
      RECT  138.1 310.5 138.9 309.7 ;
      RECT  142.1 310.5 142.9 309.7 ;
      RECT  140.1 310.5 140.9 309.7 ;
      RECT  138.1 317.5 138.9 316.7 ;
      RECT  142.1 317.5 142.9 316.7 ;
      RECT  139.1 316.0 139.9 315.2 ;
      RECT  141.1 313.2 141.9 312.4 ;
      RECT  143.6 311.8 144.2 311.2 ;
      RECT  136.9 308.7 145.5 308.1 ;
      RECT  136.9 319.1 145.5 318.5 ;
      RECT  148.7 310.5 149.5 309.7 ;
      RECT  146.7 310.5 147.5 309.7 ;
      RECT  148.7 317.9 149.5 317.1 ;
      RECT  146.7 317.9 147.5 317.1 ;
      RECT  147.1 314.2 147.9 313.4 ;
      RECT  149.1 314.1 149.7 313.5 ;
      RECT  145.5 308.7 152.1 308.1 ;
      RECT  145.5 319.1 152.1 318.5 ;
      RECT  139.1 316.0 139.9 315.2 ;
      RECT  141.1 313.2 141.9 312.4 ;
      RECT  149.1 314.1 149.7 313.5 ;
      RECT  136.9 308.7 152.1 308.1 ;
      RECT  136.9 319.1 152.1 318.5 ;
      RECT  140.1 327.1 140.9 327.9 ;
      RECT  138.1 327.1 138.9 327.9 ;
      RECT  142.1 327.1 142.9 327.9 ;
      RECT  140.1 327.1 140.9 327.9 ;
      RECT  138.1 320.1 138.9 320.9 ;
      RECT  142.1 320.1 142.9 320.9 ;
      RECT  139.1 321.6 139.9 322.4 ;
      RECT  141.1 324.4 141.9 325.2 ;
      RECT  143.6 325.8 144.2 326.4 ;
      RECT  136.9 328.9 145.5 329.5 ;
      RECT  136.9 318.5 145.5 319.1 ;
      RECT  148.7 327.1 149.5 327.9 ;
      RECT  146.7 327.1 147.5 327.9 ;
      RECT  148.7 319.7 149.5 320.5 ;
      RECT  146.7 319.7 147.5 320.5 ;
      RECT  147.1 323.4 147.9 324.2 ;
      RECT  149.1 323.5 149.7 324.1 ;
      RECT  145.5 328.9 152.1 329.5 ;
      RECT  145.5 318.5 152.1 319.1 ;
      RECT  139.1 321.6 139.9 322.4 ;
      RECT  141.1 324.4 141.9 325.2 ;
      RECT  149.1 323.5 149.7 324.1 ;
      RECT  136.9 328.9 152.1 329.5 ;
      RECT  136.9 318.5 152.1 319.1 ;
      RECT  140.1 331.3 140.9 330.5 ;
      RECT  138.1 331.3 138.9 330.5 ;
      RECT  142.1 331.3 142.9 330.5 ;
      RECT  140.1 331.3 140.9 330.5 ;
      RECT  138.1 338.3 138.9 337.5 ;
      RECT  142.1 338.3 142.9 337.5 ;
      RECT  139.1 336.8 139.9 336.0 ;
      RECT  141.1 334.0 141.9 333.2 ;
      RECT  143.6 332.6 144.2 332.0 ;
      RECT  136.9 329.5 145.5 328.9 ;
      RECT  136.9 339.9 145.5 339.3 ;
      RECT  148.7 331.3 149.5 330.5 ;
      RECT  146.7 331.3 147.5 330.5 ;
      RECT  148.7 338.7 149.5 337.9 ;
      RECT  146.7 338.7 147.5 337.9 ;
      RECT  147.1 335.0 147.9 334.2 ;
      RECT  149.1 334.9 149.7 334.3 ;
      RECT  145.5 329.5 152.1 328.9 ;
      RECT  145.5 339.9 152.1 339.3 ;
      RECT  139.1 336.8 139.9 336.0 ;
      RECT  141.1 334.0 141.9 333.2 ;
      RECT  149.1 334.9 149.7 334.3 ;
      RECT  136.9 329.5 152.1 328.9 ;
      RECT  136.9 339.9 152.1 339.3 ;
      RECT  140.1 347.9 140.9 348.7 ;
      RECT  138.1 347.9 138.9 348.7 ;
      RECT  142.1 347.9 142.9 348.7 ;
      RECT  140.1 347.9 140.9 348.7 ;
      RECT  138.1 340.9 138.9 341.7 ;
      RECT  142.1 340.9 142.9 341.7 ;
      RECT  139.1 342.4 139.9 343.2 ;
      RECT  141.1 345.2 141.9 346.0 ;
      RECT  143.6 346.6 144.2 347.2 ;
      RECT  136.9 349.7 145.5 350.3 ;
      RECT  136.9 339.3 145.5 339.9 ;
      RECT  148.7 347.9 149.5 348.7 ;
      RECT  146.7 347.9 147.5 348.7 ;
      RECT  148.7 340.5 149.5 341.3 ;
      RECT  146.7 340.5 147.5 341.3 ;
      RECT  147.1 344.2 147.9 345.0 ;
      RECT  149.1 344.3 149.7 344.9 ;
      RECT  145.5 349.7 152.1 350.3 ;
      RECT  145.5 339.3 152.1 339.9 ;
      RECT  139.1 342.4 139.9 343.2 ;
      RECT  141.1 345.2 141.9 346.0 ;
      RECT  149.1 344.3 149.7 344.9 ;
      RECT  136.9 349.7 152.1 350.3 ;
      RECT  136.9 339.3 152.1 339.9 ;
      RECT  140.1 352.1 140.9 351.3 ;
      RECT  138.1 352.1 138.9 351.3 ;
      RECT  142.1 352.1 142.9 351.3 ;
      RECT  140.1 352.1 140.9 351.3 ;
      RECT  138.1 359.1 138.9 358.3 ;
      RECT  142.1 359.1 142.9 358.3 ;
      RECT  139.1 357.6 139.9 356.8 ;
      RECT  141.1 354.8 141.9 354.0 ;
      RECT  143.6 353.4 144.2 352.8 ;
      RECT  136.9 350.3 145.5 349.7 ;
      RECT  136.9 360.7 145.5 360.1 ;
      RECT  148.7 352.1 149.5 351.3 ;
      RECT  146.7 352.1 147.5 351.3 ;
      RECT  148.7 359.5 149.5 358.7 ;
      RECT  146.7 359.5 147.5 358.7 ;
      RECT  147.1 355.8 147.9 355.0 ;
      RECT  149.1 355.7 149.7 355.1 ;
      RECT  145.5 350.3 152.1 349.7 ;
      RECT  145.5 360.7 152.1 360.1 ;
      RECT  139.1 357.6 139.9 356.8 ;
      RECT  141.1 354.8 141.9 354.0 ;
      RECT  149.1 355.7 149.7 355.1 ;
      RECT  136.9 350.3 152.1 349.7 ;
      RECT  136.9 360.7 152.1 360.1 ;
      RECT  149.1 198.7 149.7 199.3 ;
      RECT  149.1 209.5 149.7 210.1 ;
      RECT  149.1 219.5 149.7 220.1 ;
      RECT  149.1 230.3 149.7 230.9 ;
      RECT  149.1 240.3 149.7 240.9 ;
      RECT  149.1 251.1 149.7 251.7 ;
      RECT  149.1 261.1 149.7 261.7 ;
      RECT  149.1 271.9 149.7 272.5 ;
      RECT  149.1 281.9 149.7 282.5 ;
      RECT  149.1 292.7 149.7 293.3 ;
      RECT  149.1 302.7 149.7 303.3 ;
      RECT  149.1 313.5 149.7 314.1 ;
      RECT  149.1 323.5 149.7 324.1 ;
      RECT  149.1 334.3 149.7 334.9 ;
      RECT  149.1 344.3 149.7 344.9 ;
      RECT  149.1 355.1 149.7 355.7 ;
      RECT  155.9 202.3 156.7 203.1 ;
      RECT  153.9 202.3 154.7 203.1 ;
      RECT  157.9 202.3 158.7 203.1 ;
      RECT  155.9 202.3 156.7 203.1 ;
      RECT  153.9 195.3 154.7 196.1 ;
      RECT  157.9 195.3 158.7 196.1 ;
      RECT  154.9 196.8 155.7 197.6 ;
      RECT  156.9 199.6 157.7 200.4 ;
      RECT  159.4 201.0 160.0 201.6 ;
      RECT  152.7 204.1 161.3 204.7 ;
      RECT  152.7 193.7 161.3 194.3 ;
      RECT  164.5 201.5 165.3 202.3 ;
      RECT  162.5 201.5 163.3 202.3 ;
      RECT  164.5 195.3 165.3 196.1 ;
      RECT  162.5 195.3 163.3 196.1 ;
      RECT  162.9 198.4 163.7 199.2 ;
      RECT  164.9 198.5 165.5 199.1 ;
      RECT  161.3 204.1 167.9 204.7 ;
      RECT  161.3 193.7 167.9 194.3 ;
      RECT  154.9 196.8 155.7 197.6 ;
      RECT  156.9 199.6 157.7 200.4 ;
      RECT  164.9 198.5 165.5 199.1 ;
      RECT  152.7 204.1 167.9 204.7 ;
      RECT  152.7 193.7 167.9 194.3 ;
      RECT  155.9 206.5 156.7 205.7 ;
      RECT  153.9 206.5 154.7 205.7 ;
      RECT  157.9 206.5 158.7 205.7 ;
      RECT  155.9 206.5 156.7 205.7 ;
      RECT  153.9 213.5 154.7 212.7 ;
      RECT  157.9 213.5 158.7 212.7 ;
      RECT  154.9 212.0 155.7 211.2 ;
      RECT  156.9 209.2 157.7 208.4 ;
      RECT  159.4 207.8 160.0 207.2 ;
      RECT  152.7 204.7 161.3 204.1 ;
      RECT  152.7 215.1 161.3 214.5 ;
      RECT  164.5 207.3 165.3 206.5 ;
      RECT  162.5 207.3 163.3 206.5 ;
      RECT  164.5 213.5 165.3 212.7 ;
      RECT  162.5 213.5 163.3 212.7 ;
      RECT  162.9 210.4 163.7 209.6 ;
      RECT  164.9 210.3 165.5 209.7 ;
      RECT  161.3 204.7 167.9 204.1 ;
      RECT  161.3 215.1 167.9 214.5 ;
      RECT  154.9 212.0 155.7 211.2 ;
      RECT  156.9 209.2 157.7 208.4 ;
      RECT  164.9 210.3 165.5 209.7 ;
      RECT  152.7 204.7 167.9 204.1 ;
      RECT  152.7 215.1 167.9 214.5 ;
      RECT  155.9 223.1 156.7 223.9 ;
      RECT  153.9 223.1 154.7 223.9 ;
      RECT  157.9 223.1 158.7 223.9 ;
      RECT  155.9 223.1 156.7 223.9 ;
      RECT  153.9 216.1 154.7 216.9 ;
      RECT  157.9 216.1 158.7 216.9 ;
      RECT  154.9 217.6 155.7 218.4 ;
      RECT  156.9 220.4 157.7 221.2 ;
      RECT  159.4 221.8 160.0 222.4 ;
      RECT  152.7 224.9 161.3 225.5 ;
      RECT  152.7 214.5 161.3 215.1 ;
      RECT  164.5 222.3 165.3 223.1 ;
      RECT  162.5 222.3 163.3 223.1 ;
      RECT  164.5 216.1 165.3 216.9 ;
      RECT  162.5 216.1 163.3 216.9 ;
      RECT  162.9 219.2 163.7 220.0 ;
      RECT  164.9 219.3 165.5 219.9 ;
      RECT  161.3 224.9 167.9 225.5 ;
      RECT  161.3 214.5 167.9 215.1 ;
      RECT  154.9 217.6 155.7 218.4 ;
      RECT  156.9 220.4 157.7 221.2 ;
      RECT  164.9 219.3 165.5 219.9 ;
      RECT  152.7 224.9 167.9 225.5 ;
      RECT  152.7 214.5 167.9 215.1 ;
      RECT  155.9 227.3 156.7 226.5 ;
      RECT  153.9 227.3 154.7 226.5 ;
      RECT  157.9 227.3 158.7 226.5 ;
      RECT  155.9 227.3 156.7 226.5 ;
      RECT  153.9 234.3 154.7 233.5 ;
      RECT  157.9 234.3 158.7 233.5 ;
      RECT  154.9 232.8 155.7 232.0 ;
      RECT  156.9 230.0 157.7 229.2 ;
      RECT  159.4 228.6 160.0 228.0 ;
      RECT  152.7 225.5 161.3 224.9 ;
      RECT  152.7 235.9 161.3 235.3 ;
      RECT  164.5 228.1 165.3 227.3 ;
      RECT  162.5 228.1 163.3 227.3 ;
      RECT  164.5 234.3 165.3 233.5 ;
      RECT  162.5 234.3 163.3 233.5 ;
      RECT  162.9 231.2 163.7 230.4 ;
      RECT  164.9 231.1 165.5 230.5 ;
      RECT  161.3 225.5 167.9 224.9 ;
      RECT  161.3 235.9 167.9 235.3 ;
      RECT  154.9 232.8 155.7 232.0 ;
      RECT  156.9 230.0 157.7 229.2 ;
      RECT  164.9 231.1 165.5 230.5 ;
      RECT  152.7 225.5 167.9 224.9 ;
      RECT  152.7 235.9 167.9 235.3 ;
      RECT  155.9 243.9 156.7 244.7 ;
      RECT  153.9 243.9 154.7 244.7 ;
      RECT  157.9 243.9 158.7 244.7 ;
      RECT  155.9 243.9 156.7 244.7 ;
      RECT  153.9 236.9 154.7 237.7 ;
      RECT  157.9 236.9 158.7 237.7 ;
      RECT  154.9 238.4 155.7 239.2 ;
      RECT  156.9 241.2 157.7 242.0 ;
      RECT  159.4 242.6 160.0 243.2 ;
      RECT  152.7 245.7 161.3 246.3 ;
      RECT  152.7 235.3 161.3 235.9 ;
      RECT  164.5 243.1 165.3 243.9 ;
      RECT  162.5 243.1 163.3 243.9 ;
      RECT  164.5 236.9 165.3 237.7 ;
      RECT  162.5 236.9 163.3 237.7 ;
      RECT  162.9 240.0 163.7 240.8 ;
      RECT  164.9 240.1 165.5 240.7 ;
      RECT  161.3 245.7 167.9 246.3 ;
      RECT  161.3 235.3 167.9 235.9 ;
      RECT  154.9 238.4 155.7 239.2 ;
      RECT  156.9 241.2 157.7 242.0 ;
      RECT  164.9 240.1 165.5 240.7 ;
      RECT  152.7 245.7 167.9 246.3 ;
      RECT  152.7 235.3 167.9 235.9 ;
      RECT  155.9 248.1 156.7 247.3 ;
      RECT  153.9 248.1 154.7 247.3 ;
      RECT  157.9 248.1 158.7 247.3 ;
      RECT  155.9 248.1 156.7 247.3 ;
      RECT  153.9 255.1 154.7 254.3 ;
      RECT  157.9 255.1 158.7 254.3 ;
      RECT  154.9 253.6 155.7 252.8 ;
      RECT  156.9 250.8 157.7 250.0 ;
      RECT  159.4 249.4 160.0 248.8 ;
      RECT  152.7 246.3 161.3 245.7 ;
      RECT  152.7 256.7 161.3 256.1 ;
      RECT  164.5 248.9 165.3 248.1 ;
      RECT  162.5 248.9 163.3 248.1 ;
      RECT  164.5 255.1 165.3 254.3 ;
      RECT  162.5 255.1 163.3 254.3 ;
      RECT  162.9 252.0 163.7 251.2 ;
      RECT  164.9 251.9 165.5 251.3 ;
      RECT  161.3 246.3 167.9 245.7 ;
      RECT  161.3 256.7 167.9 256.1 ;
      RECT  154.9 253.6 155.7 252.8 ;
      RECT  156.9 250.8 157.7 250.0 ;
      RECT  164.9 251.9 165.5 251.3 ;
      RECT  152.7 246.3 167.9 245.7 ;
      RECT  152.7 256.7 167.9 256.1 ;
      RECT  155.9 264.7 156.7 265.5 ;
      RECT  153.9 264.7 154.7 265.5 ;
      RECT  157.9 264.7 158.7 265.5 ;
      RECT  155.9 264.7 156.7 265.5 ;
      RECT  153.9 257.7 154.7 258.5 ;
      RECT  157.9 257.7 158.7 258.5 ;
      RECT  154.9 259.2 155.7 260.0 ;
      RECT  156.9 262.0 157.7 262.8 ;
      RECT  159.4 263.4 160.0 264.0 ;
      RECT  152.7 266.5 161.3 267.1 ;
      RECT  152.7 256.1 161.3 256.7 ;
      RECT  164.5 263.9 165.3 264.7 ;
      RECT  162.5 263.9 163.3 264.7 ;
      RECT  164.5 257.7 165.3 258.5 ;
      RECT  162.5 257.7 163.3 258.5 ;
      RECT  162.9 260.8 163.7 261.6 ;
      RECT  164.9 260.9 165.5 261.5 ;
      RECT  161.3 266.5 167.9 267.1 ;
      RECT  161.3 256.1 167.9 256.7 ;
      RECT  154.9 259.2 155.7 260.0 ;
      RECT  156.9 262.0 157.7 262.8 ;
      RECT  164.9 260.9 165.5 261.5 ;
      RECT  152.7 266.5 167.9 267.1 ;
      RECT  152.7 256.1 167.9 256.7 ;
      RECT  155.9 268.9 156.7 268.1 ;
      RECT  153.9 268.9 154.7 268.1 ;
      RECT  157.9 268.9 158.7 268.1 ;
      RECT  155.9 268.9 156.7 268.1 ;
      RECT  153.9 275.9 154.7 275.1 ;
      RECT  157.9 275.9 158.7 275.1 ;
      RECT  154.9 274.4 155.7 273.6 ;
      RECT  156.9 271.6 157.7 270.8 ;
      RECT  159.4 270.2 160.0 269.6 ;
      RECT  152.7 267.1 161.3 266.5 ;
      RECT  152.7 277.5 161.3 276.9 ;
      RECT  164.5 269.7 165.3 268.9 ;
      RECT  162.5 269.7 163.3 268.9 ;
      RECT  164.5 275.9 165.3 275.1 ;
      RECT  162.5 275.9 163.3 275.1 ;
      RECT  162.9 272.8 163.7 272.0 ;
      RECT  164.9 272.7 165.5 272.1 ;
      RECT  161.3 267.1 167.9 266.5 ;
      RECT  161.3 277.5 167.9 276.9 ;
      RECT  154.9 274.4 155.7 273.6 ;
      RECT  156.9 271.6 157.7 270.8 ;
      RECT  164.9 272.7 165.5 272.1 ;
      RECT  152.7 267.1 167.9 266.5 ;
      RECT  152.7 277.5 167.9 276.9 ;
      RECT  155.9 285.5 156.7 286.3 ;
      RECT  153.9 285.5 154.7 286.3 ;
      RECT  157.9 285.5 158.7 286.3 ;
      RECT  155.9 285.5 156.7 286.3 ;
      RECT  153.9 278.5 154.7 279.3 ;
      RECT  157.9 278.5 158.7 279.3 ;
      RECT  154.9 280.0 155.7 280.8 ;
      RECT  156.9 282.8 157.7 283.6 ;
      RECT  159.4 284.2 160.0 284.8 ;
      RECT  152.7 287.3 161.3 287.9 ;
      RECT  152.7 276.9 161.3 277.5 ;
      RECT  164.5 284.7 165.3 285.5 ;
      RECT  162.5 284.7 163.3 285.5 ;
      RECT  164.5 278.5 165.3 279.3 ;
      RECT  162.5 278.5 163.3 279.3 ;
      RECT  162.9 281.6 163.7 282.4 ;
      RECT  164.9 281.7 165.5 282.3 ;
      RECT  161.3 287.3 167.9 287.9 ;
      RECT  161.3 276.9 167.9 277.5 ;
      RECT  154.9 280.0 155.7 280.8 ;
      RECT  156.9 282.8 157.7 283.6 ;
      RECT  164.9 281.7 165.5 282.3 ;
      RECT  152.7 287.3 167.9 287.9 ;
      RECT  152.7 276.9 167.9 277.5 ;
      RECT  155.9 289.7 156.7 288.9 ;
      RECT  153.9 289.7 154.7 288.9 ;
      RECT  157.9 289.7 158.7 288.9 ;
      RECT  155.9 289.7 156.7 288.9 ;
      RECT  153.9 296.7 154.7 295.9 ;
      RECT  157.9 296.7 158.7 295.9 ;
      RECT  154.9 295.2 155.7 294.4 ;
      RECT  156.9 292.4 157.7 291.6 ;
      RECT  159.4 291.0 160.0 290.4 ;
      RECT  152.7 287.9 161.3 287.3 ;
      RECT  152.7 298.3 161.3 297.7 ;
      RECT  164.5 290.5 165.3 289.7 ;
      RECT  162.5 290.5 163.3 289.7 ;
      RECT  164.5 296.7 165.3 295.9 ;
      RECT  162.5 296.7 163.3 295.9 ;
      RECT  162.9 293.6 163.7 292.8 ;
      RECT  164.9 293.5 165.5 292.9 ;
      RECT  161.3 287.9 167.9 287.3 ;
      RECT  161.3 298.3 167.9 297.7 ;
      RECT  154.9 295.2 155.7 294.4 ;
      RECT  156.9 292.4 157.7 291.6 ;
      RECT  164.9 293.5 165.5 292.9 ;
      RECT  152.7 287.9 167.9 287.3 ;
      RECT  152.7 298.3 167.9 297.7 ;
      RECT  155.9 306.3 156.7 307.1 ;
      RECT  153.9 306.3 154.7 307.1 ;
      RECT  157.9 306.3 158.7 307.1 ;
      RECT  155.9 306.3 156.7 307.1 ;
      RECT  153.9 299.3 154.7 300.1 ;
      RECT  157.9 299.3 158.7 300.1 ;
      RECT  154.9 300.8 155.7 301.6 ;
      RECT  156.9 303.6 157.7 304.4 ;
      RECT  159.4 305.0 160.0 305.6 ;
      RECT  152.7 308.1 161.3 308.7 ;
      RECT  152.7 297.7 161.3 298.3 ;
      RECT  164.5 305.5 165.3 306.3 ;
      RECT  162.5 305.5 163.3 306.3 ;
      RECT  164.5 299.3 165.3 300.1 ;
      RECT  162.5 299.3 163.3 300.1 ;
      RECT  162.9 302.4 163.7 303.2 ;
      RECT  164.9 302.5 165.5 303.1 ;
      RECT  161.3 308.1 167.9 308.7 ;
      RECT  161.3 297.7 167.9 298.3 ;
      RECT  154.9 300.8 155.7 301.6 ;
      RECT  156.9 303.6 157.7 304.4 ;
      RECT  164.9 302.5 165.5 303.1 ;
      RECT  152.7 308.1 167.9 308.7 ;
      RECT  152.7 297.7 167.9 298.3 ;
      RECT  155.9 310.5 156.7 309.7 ;
      RECT  153.9 310.5 154.7 309.7 ;
      RECT  157.9 310.5 158.7 309.7 ;
      RECT  155.9 310.5 156.7 309.7 ;
      RECT  153.9 317.5 154.7 316.7 ;
      RECT  157.9 317.5 158.7 316.7 ;
      RECT  154.9 316.0 155.7 315.2 ;
      RECT  156.9 313.2 157.7 312.4 ;
      RECT  159.4 311.8 160.0 311.2 ;
      RECT  152.7 308.7 161.3 308.1 ;
      RECT  152.7 319.1 161.3 318.5 ;
      RECT  164.5 311.3 165.3 310.5 ;
      RECT  162.5 311.3 163.3 310.5 ;
      RECT  164.5 317.5 165.3 316.7 ;
      RECT  162.5 317.5 163.3 316.7 ;
      RECT  162.9 314.4 163.7 313.6 ;
      RECT  164.9 314.3 165.5 313.7 ;
      RECT  161.3 308.7 167.9 308.1 ;
      RECT  161.3 319.1 167.9 318.5 ;
      RECT  154.9 316.0 155.7 315.2 ;
      RECT  156.9 313.2 157.7 312.4 ;
      RECT  164.9 314.3 165.5 313.7 ;
      RECT  152.7 308.7 167.9 308.1 ;
      RECT  152.7 319.1 167.9 318.5 ;
      RECT  155.9 327.1 156.7 327.9 ;
      RECT  153.9 327.1 154.7 327.9 ;
      RECT  157.9 327.1 158.7 327.9 ;
      RECT  155.9 327.1 156.7 327.9 ;
      RECT  153.9 320.1 154.7 320.9 ;
      RECT  157.9 320.1 158.7 320.9 ;
      RECT  154.9 321.6 155.7 322.4 ;
      RECT  156.9 324.4 157.7 325.2 ;
      RECT  159.4 325.8 160.0 326.4 ;
      RECT  152.7 328.9 161.3 329.5 ;
      RECT  152.7 318.5 161.3 319.1 ;
      RECT  164.5 326.3 165.3 327.1 ;
      RECT  162.5 326.3 163.3 327.1 ;
      RECT  164.5 320.1 165.3 320.9 ;
      RECT  162.5 320.1 163.3 320.9 ;
      RECT  162.9 323.2 163.7 324.0 ;
      RECT  164.9 323.3 165.5 323.9 ;
      RECT  161.3 328.9 167.9 329.5 ;
      RECT  161.3 318.5 167.9 319.1 ;
      RECT  154.9 321.6 155.7 322.4 ;
      RECT  156.9 324.4 157.7 325.2 ;
      RECT  164.9 323.3 165.5 323.9 ;
      RECT  152.7 328.9 167.9 329.5 ;
      RECT  152.7 318.5 167.9 319.1 ;
      RECT  155.9 331.3 156.7 330.5 ;
      RECT  153.9 331.3 154.7 330.5 ;
      RECT  157.9 331.3 158.7 330.5 ;
      RECT  155.9 331.3 156.7 330.5 ;
      RECT  153.9 338.3 154.7 337.5 ;
      RECT  157.9 338.3 158.7 337.5 ;
      RECT  154.9 336.8 155.7 336.0 ;
      RECT  156.9 334.0 157.7 333.2 ;
      RECT  159.4 332.6 160.0 332.0 ;
      RECT  152.7 329.5 161.3 328.9 ;
      RECT  152.7 339.9 161.3 339.3 ;
      RECT  164.5 332.1 165.3 331.3 ;
      RECT  162.5 332.1 163.3 331.3 ;
      RECT  164.5 338.3 165.3 337.5 ;
      RECT  162.5 338.3 163.3 337.5 ;
      RECT  162.9 335.2 163.7 334.4 ;
      RECT  164.9 335.1 165.5 334.5 ;
      RECT  161.3 329.5 167.9 328.9 ;
      RECT  161.3 339.9 167.9 339.3 ;
      RECT  154.9 336.8 155.7 336.0 ;
      RECT  156.9 334.0 157.7 333.2 ;
      RECT  164.9 335.1 165.5 334.5 ;
      RECT  152.7 329.5 167.9 328.9 ;
      RECT  152.7 339.9 167.9 339.3 ;
      RECT  155.9 347.9 156.7 348.7 ;
      RECT  153.9 347.9 154.7 348.7 ;
      RECT  157.9 347.9 158.7 348.7 ;
      RECT  155.9 347.9 156.7 348.7 ;
      RECT  153.9 340.9 154.7 341.7 ;
      RECT  157.9 340.9 158.7 341.7 ;
      RECT  154.9 342.4 155.7 343.2 ;
      RECT  156.9 345.2 157.7 346.0 ;
      RECT  159.4 346.6 160.0 347.2 ;
      RECT  152.7 349.7 161.3 350.3 ;
      RECT  152.7 339.3 161.3 339.9 ;
      RECT  164.5 347.1 165.3 347.9 ;
      RECT  162.5 347.1 163.3 347.9 ;
      RECT  164.5 340.9 165.3 341.7 ;
      RECT  162.5 340.9 163.3 341.7 ;
      RECT  162.9 344.0 163.7 344.8 ;
      RECT  164.9 344.1 165.5 344.7 ;
      RECT  161.3 349.7 167.9 350.3 ;
      RECT  161.3 339.3 167.9 339.9 ;
      RECT  154.9 342.4 155.7 343.2 ;
      RECT  156.9 345.2 157.7 346.0 ;
      RECT  164.9 344.1 165.5 344.7 ;
      RECT  152.7 349.7 167.9 350.3 ;
      RECT  152.7 339.3 167.9 339.9 ;
      RECT  155.9 352.1 156.7 351.3 ;
      RECT  153.9 352.1 154.7 351.3 ;
      RECT  157.9 352.1 158.7 351.3 ;
      RECT  155.9 352.1 156.7 351.3 ;
      RECT  153.9 359.1 154.7 358.3 ;
      RECT  157.9 359.1 158.7 358.3 ;
      RECT  154.9 357.6 155.7 356.8 ;
      RECT  156.9 354.8 157.7 354.0 ;
      RECT  159.4 353.4 160.0 352.8 ;
      RECT  152.7 350.3 161.3 349.7 ;
      RECT  152.7 360.7 161.3 360.1 ;
      RECT  164.5 352.9 165.3 352.1 ;
      RECT  162.5 352.9 163.3 352.1 ;
      RECT  164.5 359.1 165.3 358.3 ;
      RECT  162.5 359.1 163.3 358.3 ;
      RECT  162.9 356.0 163.7 355.2 ;
      RECT  164.9 355.9 165.5 355.3 ;
      RECT  161.3 350.3 167.9 349.7 ;
      RECT  161.3 360.7 167.9 360.1 ;
      RECT  154.9 357.6 155.7 356.8 ;
      RECT  156.9 354.8 157.7 354.0 ;
      RECT  164.9 355.9 165.5 355.3 ;
      RECT  152.7 350.3 167.9 349.7 ;
      RECT  152.7 360.7 167.9 360.1 ;
      RECT  154.9 196.8 155.7 197.6 ;
      RECT  154.9 211.2 155.7 212.0 ;
      RECT  154.9 217.6 155.7 218.4 ;
      RECT  154.9 232.0 155.7 232.8 ;
      RECT  154.9 238.4 155.7 239.2 ;
      RECT  154.9 252.8 155.7 253.6 ;
      RECT  154.9 259.2 155.7 260.0 ;
      RECT  154.9 273.6 155.7 274.4 ;
      RECT  154.9 280.0 155.7 280.8 ;
      RECT  154.9 294.4 155.7 295.2 ;
      RECT  154.9 300.8 155.7 301.6 ;
      RECT  154.9 315.2 155.7 316.0 ;
      RECT  154.9 321.6 155.7 322.4 ;
      RECT  154.9 336.0 155.7 336.8 ;
      RECT  154.9 342.4 155.7 343.2 ;
      RECT  154.9 356.8 155.7 357.6 ;
      RECT  164.9 198.5 165.5 199.1 ;
      RECT  164.9 209.7 165.5 210.3 ;
      RECT  164.9 219.3 165.5 219.9 ;
      RECT  164.9 230.5 165.5 231.1 ;
      RECT  164.9 240.1 165.5 240.7 ;
      RECT  164.9 251.3 165.5 251.9 ;
      RECT  164.9 260.9 165.5 261.5 ;
      RECT  164.9 272.1 165.5 272.7 ;
      RECT  164.9 281.7 165.5 282.3 ;
      RECT  164.9 292.9 165.5 293.5 ;
      RECT  164.9 302.5 165.5 303.1 ;
      RECT  164.9 313.7 165.5 314.3 ;
      RECT  164.9 323.3 165.5 323.9 ;
      RECT  164.9 334.5 165.5 335.1 ;
      RECT  164.9 344.1 165.5 344.7 ;
      RECT  164.9 355.3 165.5 355.9 ;
      RECT  164.9 198.5 165.5 199.1 ;
      RECT  164.9 209.7 165.5 210.3 ;
      RECT  164.9 219.3 165.5 219.9 ;
      RECT  164.9 230.5 165.5 231.1 ;
      RECT  164.9 240.1 165.5 240.7 ;
      RECT  164.9 251.3 165.5 251.9 ;
      RECT  164.9 260.9 165.5 261.5 ;
      RECT  164.9 272.1 165.5 272.7 ;
      RECT  164.9 281.7 165.5 282.3 ;
      RECT  164.9 292.9 165.5 293.5 ;
      RECT  164.9 302.5 165.5 303.1 ;
      RECT  164.9 313.7 165.5 314.3 ;
      RECT  164.9 323.3 165.5 323.9 ;
      RECT  164.9 334.5 165.5 335.1 ;
      RECT  164.9 344.1 165.5 344.7 ;
      RECT  164.9 355.3 165.5 355.9 ;
      RECT  16.4 9.6 17.2 9.8 ;
      RECT  3.6 2.8 4.4 7.6 ;
      RECT  12.4 15.8 13.0 16.4 ;
      RECT  10.2 15.2 13.8 15.8 ;
      RECT  3.6 11.4 9.2 11.6 ;
      RECT  4.4 8.4 15.4 9.0 ;
      RECT  21.2 11.8 22.0 20.4 ;
      RECT  12.4 4.8 13.0 5.4 ;
      RECT  8.0 2.8 8.8 4.2 ;
      RECT  10.2 15.0 11.0 15.2 ;
      RECT  16.4 15.6 17.2 16.4 ;
      RECT  12.8 12.4 13.4 13.6 ;
      RECT  6.8 16.4 8.8 17.0 ;
      RECT  14.0 2.2 14.8 4.8 ;
      RECT  10.2 5.4 13.0 6.0 ;
      RECT  6.8 4.2 8.8 4.8 ;
      RECT  21.2 7.8 22.0 11.2 ;
      RECT  16.6 16.4 17.8 20.4 ;
      RECT  5.2 12.6 6.0 21.0 ;
      RECT  6.8 13.0 12.2 13.6 ;
      RECT  14.8 9.0 15.4 12.2 ;
      RECT  2.4 21.0 24.2 22.2 ;
      RECT  17.8 11.2 22.0 11.8 ;
      RECT  19.6 12.4 20.4 21.0 ;
      RECT  22.8 2.2 23.6 3.6 ;
      RECT  16.6 12.8 17.2 13.8 ;
      RECT  14.8 12.2 17.2 12.8 ;
      RECT  3.6 12.0 4.4 20.4 ;
      RECT  16.4 4.2 17.8 4.8 ;
      RECT  12.8 13.6 15.0 14.2 ;
      RECT  8.0 17.0 8.8 20.4 ;
      RECT  5.8 10.2 10.8 10.8 ;
      RECT  22.8 19.4 23.6 21.0 ;
      RECT  16.4 9.8 20.2 10.4 ;
      RECT  16.4 4.8 17.2 5.6 ;
      RECT  2.4 1.0 24.2 2.2 ;
      RECT  10.0 10.8 10.8 11.0 ;
      RECT  7.4 9.0 8.2 9.2 ;
      RECT  13.0 15.0 13.8 15.2 ;
      RECT  21.2 2.8 22.0 7.2 ;
      RECT  4.4 8.2 6.0 8.4 ;
      RECT  6.8 15.6 7.6 16.4 ;
      RECT  12.4 2.8 13.2 4.8 ;
      RECT  5.8 10.0 6.6 10.2 ;
      RECT  6.8 13.6 7.6 13.8 ;
      RECT  18.2 7.0 19.0 7.2 ;
      RECT  8.4 5.4 9.2 6.2 ;
      RECT  19.6 2.2 20.4 6.6 ;
      RECT  14.2 13.4 15.0 13.6 ;
      RECT  10.6 2.2 11.6 4.8 ;
      RECT  8.6 6.2 9.2 8.4 ;
      RECT  14.0 16.4 14.8 21.0 ;
      RECT  10.8 16.4 11.6 21.0 ;
      RECT  14.2 8.2 15.0 8.4 ;
      RECT  8.6 12.0 13.4 12.4 ;
      RECT  3.6 11.6 9.4 11.8 ;
      RECT  12.4 16.4 13.2 20.4 ;
      RECT  19.4 10.4 20.2 10.6 ;
      RECT  3.6 11.8 13.4 12.0 ;
      RECT  11.4 13.6 12.2 13.8 ;
      RECT  16.6 2.8 17.8 4.2 ;
      RECT  10.2 6.0 11.0 6.2 ;
      RECT  16.6 13.8 18.0 14.6 ;
      RECT  17.8 11.0 18.6 11.2 ;
      RECT  6.8 4.8 7.6 5.6 ;
      RECT  5.2 2.2 6.0 6.8 ;
      RECT  18.2 7.2 22.0 7.8 ;
      RECT  29.8 18.7 30.6 19.5 ;
      RECT  27.8 18.7 28.6 19.5 ;
      RECT  29.8 2.9 30.6 3.7 ;
      RECT  27.8 2.9 28.6 3.7 ;
      RECT  28.2 10.8 29.0 11.6 ;
      RECT  30.2 10.9 30.8 11.5 ;
      RECT  26.6 21.3 33.2 21.9 ;
      RECT  26.6 1.3 33.2 1.9 ;
      RECT  36.4 17.1 37.2 17.9 ;
      RECT  34.4 17.1 35.2 17.9 ;
      RECT  36.4 3.7 37.2 4.5 ;
      RECT  34.4 3.7 35.2 4.5 ;
      RECT  34.8 10.4 35.6 11.2 ;
      RECT  36.8 10.5 37.4 11.1 ;
      RECT  33.2 21.3 39.8 21.9 ;
      RECT  33.2 1.3 39.8 1.9 ;
      RECT  2.4 21.0 39.8 22.2 ;
      RECT  2.4 1.0 39.8 2.2 ;
      RECT  16.4 33.6 17.2 33.4 ;
      RECT  3.6 40.4 4.4 35.6 ;
      RECT  12.4 27.4 13.0 26.8 ;
      RECT  10.2 28.0 13.8 27.4 ;
      RECT  3.6 31.8 9.2 31.6 ;
      RECT  4.4 34.8 15.4 34.2 ;
      RECT  21.2 31.4 22.0 22.8 ;
      RECT  12.4 38.4 13.0 37.8 ;
      RECT  8.0 40.4 8.8 39.0 ;
      RECT  10.2 28.2 11.0 28.0 ;
      RECT  16.4 27.6 17.2 26.8 ;
      RECT  12.8 30.8 13.4 29.6 ;
      RECT  6.8 26.8 8.8 26.2 ;
      RECT  14.0 41.0 14.8 38.4 ;
      RECT  10.2 37.8 13.0 37.2 ;
      RECT  6.8 39.0 8.8 38.4 ;
      RECT  21.2 35.4 22.0 32.0 ;
      RECT  16.6 26.8 17.8 22.8 ;
      RECT  5.2 30.6 6.0 22.2 ;
      RECT  6.8 30.2 12.2 29.6 ;
      RECT  14.8 34.2 15.4 31.0 ;
      RECT  2.4 22.2 24.2 21.0 ;
      RECT  17.8 32.0 22.0 31.4 ;
      RECT  19.6 30.8 20.4 22.2 ;
      RECT  22.8 41.0 23.6 39.6 ;
      RECT  16.6 30.4 17.2 29.4 ;
      RECT  14.8 31.0 17.2 30.4 ;
      RECT  3.6 31.2 4.4 22.8 ;
      RECT  16.4 39.0 17.8 38.4 ;
      RECT  12.8 29.6 15.0 29.0 ;
      RECT  8.0 26.2 8.8 22.8 ;
      RECT  5.8 33.0 10.8 32.4 ;
      RECT  22.8 23.8 23.6 22.2 ;
      RECT  16.4 33.4 20.2 32.8 ;
      RECT  16.4 38.4 17.2 37.6 ;
      RECT  2.4 42.2 24.2 41.0 ;
      RECT  10.0 32.4 10.8 32.2 ;
      RECT  7.4 34.2 8.2 34.0 ;
      RECT  13.0 28.2 13.8 28.0 ;
      RECT  21.2 40.4 22.0 36.0 ;
      RECT  4.4 35.0 6.0 34.8 ;
      RECT  6.8 27.6 7.6 26.8 ;
      RECT  12.4 40.4 13.2 38.4 ;
      RECT  5.8 33.2 6.6 33.0 ;
      RECT  6.8 29.6 7.6 29.4 ;
      RECT  18.2 36.2 19.0 36.0 ;
      RECT  8.4 37.8 9.2 37.0 ;
      RECT  19.6 41.0 20.4 36.6 ;
      RECT  14.2 29.8 15.0 29.6 ;
      RECT  10.6 41.0 11.6 38.4 ;
      RECT  8.6 37.0 9.2 34.8 ;
      RECT  14.0 26.8 14.8 22.2 ;
      RECT  10.8 26.8 11.6 22.2 ;
      RECT  14.2 35.0 15.0 34.8 ;
      RECT  8.6 31.2 13.4 30.8 ;
      RECT  3.6 31.6 9.4 31.4 ;
      RECT  12.4 26.8 13.2 22.8 ;
      RECT  19.4 32.8 20.2 32.6 ;
      RECT  3.6 31.4 13.4 31.2 ;
      RECT  11.4 29.6 12.2 29.4 ;
      RECT  16.6 40.4 17.8 39.0 ;
      RECT  10.2 37.2 11.0 37.0 ;
      RECT  16.6 29.4 18.0 28.6 ;
      RECT  17.8 32.2 18.6 32.0 ;
      RECT  6.8 38.4 7.6 37.6 ;
      RECT  5.2 41.0 6.0 36.4 ;
      RECT  18.2 36.0 22.0 35.4 ;
      RECT  29.8 24.5 30.6 23.7 ;
      RECT  27.8 24.5 28.6 23.7 ;
      RECT  29.8 40.3 30.6 39.5 ;
      RECT  27.8 40.3 28.6 39.5 ;
      RECT  28.2 32.4 29.0 31.6 ;
      RECT  30.2 32.3 30.8 31.7 ;
      RECT  26.6 21.9 33.2 21.3 ;
      RECT  26.6 41.9 33.2 41.3 ;
      RECT  36.4 26.1 37.2 25.3 ;
      RECT  34.4 26.1 35.2 25.3 ;
      RECT  36.4 39.5 37.2 38.7 ;
      RECT  34.4 39.5 35.2 38.7 ;
      RECT  34.8 32.8 35.6 32.0 ;
      RECT  36.8 32.7 37.4 32.1 ;
      RECT  33.2 21.9 39.8 21.3 ;
      RECT  33.2 41.9 39.8 41.3 ;
      RECT  2.4 22.2 39.8 21.0 ;
      RECT  2.4 42.2 39.8 41.0 ;
      RECT  55.6 19.5 56.4 20.3 ;
      RECT  53.6 19.5 54.4 20.3 ;
      RECT  55.6 2.5 56.4 3.3 ;
      RECT  53.6 2.5 54.4 3.3 ;
      RECT  54.0 11.0 54.8 11.8 ;
      RECT  56.0 11.1 56.6 11.7 ;
      RECT  52.4 21.3 59.0 21.9 ;
      RECT  52.4 1.3 59.0 1.9 ;
      RECT  62.2 18.7 63.0 19.5 ;
      RECT  60.2 18.7 61.0 19.5 ;
      RECT  62.2 2.9 63.0 3.7 ;
      RECT  60.2 2.9 61.0 3.7 ;
      RECT  60.6 10.8 61.4 11.6 ;
      RECT  62.6 10.9 63.2 11.5 ;
      RECT  59.0 21.3 64.2 21.9 ;
      RECT  59.0 1.3 64.2 1.9 ;
      RECT  67.4 16.3 68.2 17.1 ;
      RECT  65.4 16.3 66.2 17.1 ;
      RECT  67.4 4.1 68.2 4.9 ;
      RECT  65.4 4.1 66.2 4.9 ;
      RECT  65.8 10.2 66.6 11.0 ;
      RECT  67.8 10.3 68.4 10.9 ;
      RECT  64.2 21.3 69.4 21.9 ;
      RECT  64.2 1.3 69.4 1.9 ;
      RECT  72.5 15.1 76.5 15.7 ;
      RECT  70.6 16.3 71.4 17.1 ;
      RECT  74.0 16.3 74.8 17.1 ;
      RECT  72.5 5.5 76.5 6.1 ;
      RECT  74.0 4.1 74.8 4.9 ;
      RECT  70.6 4.1 71.4 4.9 ;
      RECT  71.0 10.2 71.8 11.0 ;
      RECT  74.5 10.3 75.1 10.9 ;
      RECT  69.4 21.3 78.0 21.9 ;
      RECT  69.4 1.3 78.0 1.9 ;
      RECT  54.0 11.0 54.8 11.8 ;
      RECT  74.5 10.3 75.1 10.9 ;
      RECT  52.4 21.3 78.0 21.9 ;
      RECT  52.4 1.3 78.0 1.9 ;
      RECT  55.6 23.7 56.4 22.9 ;
      RECT  53.6 23.7 54.4 22.9 ;
      RECT  55.6 40.7 56.4 39.9 ;
      RECT  53.6 40.7 54.4 39.9 ;
      RECT  54.0 32.2 54.8 31.4 ;
      RECT  56.0 32.1 56.6 31.5 ;
      RECT  52.4 21.9 59.0 21.3 ;
      RECT  52.4 41.9 59.0 41.3 ;
      RECT  62.2 23.7 63.0 22.9 ;
      RECT  60.2 23.7 61.0 22.9 ;
      RECT  64.2 23.7 65.0 22.9 ;
      RECT  62.2 23.7 63.0 22.9 ;
      RECT  60.2 40.3 61.0 39.5 ;
      RECT  64.2 40.3 65.0 39.5 ;
      RECT  61.2 38.8 62.0 38.0 ;
      RECT  63.2 36.0 64.0 35.2 ;
      RECT  65.7 25.0 66.3 24.4 ;
      RECT  59.0 21.9 66.6 21.3 ;
      RECT  59.0 41.9 66.6 41.3 ;
      RECT  69.7 27.3 73.7 26.7 ;
      RECT  71.2 26.1 72.0 25.3 ;
      RECT  67.8 26.1 68.6 25.3 ;
      RECT  69.7 38.1 73.7 37.5 ;
      RECT  71.2 39.5 72.0 38.7 ;
      RECT  67.8 39.5 68.6 38.7 ;
      RECT  68.2 32.8 69.0 32.0 ;
      RECT  71.7 32.7 72.3 32.1 ;
      RECT  66.6 21.9 76.4 21.3 ;
      RECT  66.6 41.9 76.4 41.3 ;
      RECT  68.2 32.8 69.0 32.0 ;
      RECT  71.7 32.7 72.3 32.1 ;
      RECT  66.6 21.9 76.4 21.3 ;
      RECT  66.6 41.9 76.4 41.3 ;
      RECT  61.2 38.8 62.0 38.0 ;
      RECT  63.2 36.0 64.0 35.2 ;
      RECT  71.7 32.7 72.3 32.1 ;
      RECT  59.0 21.9 76.4 21.3 ;
      RECT  59.0 41.9 76.4 41.3 ;
      RECT  55.6 59.5 56.4 60.3 ;
      RECT  53.6 59.5 54.4 60.3 ;
      RECT  57.6 59.5 58.4 60.3 ;
      RECT  55.6 59.5 56.4 60.3 ;
      RECT  53.6 42.9 54.4 43.7 ;
      RECT  57.6 42.9 58.4 43.7 ;
      RECT  54.6 44.4 55.4 45.2 ;
      RECT  56.6 47.2 57.4 48.0 ;
      RECT  59.1 58.2 59.7 58.8 ;
      RECT  52.4 61.3 60.0 61.9 ;
      RECT  52.4 41.3 60.0 41.9 ;
      RECT  63.1 55.9 67.1 56.5 ;
      RECT  64.6 57.1 65.4 57.9 ;
      RECT  61.2 57.1 62.0 57.9 ;
      RECT  63.1 45.1 67.1 45.7 ;
      RECT  64.6 43.7 65.4 44.5 ;
      RECT  61.2 43.7 62.0 44.5 ;
      RECT  61.6 50.4 62.4 51.2 ;
      RECT  65.1 50.5 65.7 51.1 ;
      RECT  60.0 61.3 69.8 61.9 ;
      RECT  60.0 41.3 69.8 41.9 ;
      RECT  61.6 50.4 62.4 51.2 ;
      RECT  65.1 50.5 65.7 51.1 ;
      RECT  60.0 61.3 69.8 61.9 ;
      RECT  60.0 41.3 69.8 41.9 ;
      RECT  54.6 44.4 55.4 45.2 ;
      RECT  56.6 47.2 57.4 48.0 ;
      RECT  65.1 50.5 65.7 51.1 ;
      RECT  52.4 61.3 69.8 61.9 ;
      RECT  52.4 41.3 69.8 41.9 ;
      RECT  55.6 63.7 56.4 62.9 ;
      RECT  53.6 63.7 54.4 62.9 ;
      RECT  55.6 80.7 56.4 79.9 ;
      RECT  53.6 80.7 54.4 79.9 ;
      RECT  54.0 72.2 54.8 71.4 ;
      RECT  56.0 72.1 56.6 71.5 ;
      RECT  52.4 61.9 59.0 61.3 ;
      RECT  52.4 81.9 59.0 81.3 ;
      RECT  62.2 63.7 63.0 62.9 ;
      RECT  60.2 63.7 61.0 62.9 ;
      RECT  62.2 80.7 63.0 79.9 ;
      RECT  60.2 80.7 61.0 79.9 ;
      RECT  60.6 72.2 61.4 71.4 ;
      RECT  62.6 72.1 63.2 71.5 ;
      RECT  59.0 61.9 64.2 61.3 ;
      RECT  59.0 81.9 64.2 81.3 ;
      RECT  67.4 64.5 68.2 63.7 ;
      RECT  65.4 64.5 66.2 63.7 ;
      RECT  67.4 80.3 68.2 79.5 ;
      RECT  65.4 80.3 66.2 79.5 ;
      RECT  65.8 72.4 66.6 71.6 ;
      RECT  67.8 72.3 68.4 71.7 ;
      RECT  64.2 61.9 69.4 61.3 ;
      RECT  64.2 81.9 69.4 81.3 ;
      RECT  72.6 66.9 73.4 66.1 ;
      RECT  70.6 66.9 71.4 66.1 ;
      RECT  72.6 79.1 73.4 78.3 ;
      RECT  70.6 79.1 71.4 78.3 ;
      RECT  71.0 73.0 71.8 72.2 ;
      RECT  73.0 72.9 73.6 72.3 ;
      RECT  69.4 61.9 74.6 61.3 ;
      RECT  69.4 81.9 74.6 81.3 ;
      RECT  54.0 72.2 54.8 71.4 ;
      RECT  73.0 72.9 73.6 72.3 ;
      RECT  52.4 61.9 74.6 61.3 ;
      RECT  52.4 81.9 74.6 81.3 ;
      RECT  55.6 139.5 56.4 140.3 ;
      RECT  53.6 139.5 54.4 140.3 ;
      RECT  55.6 122.5 56.4 123.3 ;
      RECT  53.6 122.5 54.4 123.3 ;
      RECT  54.0 131.0 54.8 131.8 ;
      RECT  56.0 131.1 56.6 131.7 ;
      RECT  52.4 141.3 59.0 141.9 ;
      RECT  52.4 121.3 59.0 121.9 ;
      RECT  55.6 99.5 56.4 100.3 ;
      RECT  53.6 99.5 54.4 100.3 ;
      RECT  57.6 99.5 58.4 100.3 ;
      RECT  55.6 99.5 56.4 100.3 ;
      RECT  59.6 99.5 60.4 100.3 ;
      RECT  57.6 99.5 58.4 100.3 ;
      RECT  53.6 82.9 54.4 83.7 ;
      RECT  59.6 82.9 60.4 83.7 ;
      RECT  54.2 84.4 55.0 85.2 ;
      RECT  56.6 85.7 57.4 86.5 ;
      RECT  59.0 87.0 59.8 87.8 ;
      RECT  61.1 98.3 61.7 98.9 ;
      RECT  52.4 101.3 62.0 101.9 ;
      RECT  52.4 81.3 62.0 81.9 ;
      RECT  65.0 96.3 65.8 97.1 ;
      RECT  63.2 96.3 64.0 97.1 ;
      RECT  66.8 96.3 67.6 97.1 ;
      RECT  65.0 84.1 65.8 84.9 ;
      RECT  66.8 84.1 67.6 84.9 ;
      RECT  63.2 84.1 64.0 84.9 ;
      RECT  63.6 90.2 64.4 91.0 ;
      RECT  65.4 90.3 66.0 90.9 ;
      RECT  62.0 101.3 70.2 101.9 ;
      RECT  62.0 81.3 70.2 81.9 ;
      RECT  63.6 90.2 64.4 91.0 ;
      RECT  65.4 90.3 66.0 90.9 ;
      RECT  62.0 101.3 70.2 101.9 ;
      RECT  62.0 81.3 70.2 81.9 ;
      RECT  54.2 84.4 55.0 85.2 ;
      RECT  56.6 85.7 57.4 86.5 ;
      RECT  59.0 87.0 59.8 87.8 ;
      RECT  65.4 90.3 66.0 90.9 ;
      RECT  52.4 101.3 70.2 101.9 ;
      RECT  52.4 81.3 70.2 81.9 ;
      RECT  55.6 143.7 56.4 142.9 ;
      RECT  53.6 143.7 54.4 142.9 ;
      RECT  57.6 143.7 58.4 142.9 ;
      RECT  55.6 143.7 56.4 142.9 ;
      RECT  59.6 143.7 60.4 142.9 ;
      RECT  57.6 143.7 58.4 142.9 ;
      RECT  53.6 160.3 54.4 159.5 ;
      RECT  59.6 160.3 60.4 159.5 ;
      RECT  54.2 158.8 55.0 158.0 ;
      RECT  56.6 157.5 57.4 156.7 ;
      RECT  59.0 156.2 59.8 155.4 ;
      RECT  61.1 144.9 61.7 144.3 ;
      RECT  52.4 141.9 62.0 141.3 ;
      RECT  52.4 161.9 62.0 161.3 ;
      RECT  65.2 144.5 66.0 143.7 ;
      RECT  63.2 144.5 64.0 143.7 ;
      RECT  65.2 160.3 66.0 159.5 ;
      RECT  63.2 160.3 64.0 159.5 ;
      RECT  63.6 152.4 64.4 151.6 ;
      RECT  65.6 152.3 66.2 151.7 ;
      RECT  62.0 141.9 68.6 141.3 ;
      RECT  62.0 161.9 68.6 161.3 ;
      RECT  63.6 152.4 64.4 151.6 ;
      RECT  65.6 152.3 66.2 151.7 ;
      RECT  62.0 141.9 68.6 141.3 ;
      RECT  62.0 161.9 68.6 161.3 ;
      RECT  54.2 158.8 55.0 158.0 ;
      RECT  56.6 157.5 57.4 156.7 ;
      RECT  59.0 156.2 59.8 155.4 ;
      RECT  65.6 152.3 66.2 151.7 ;
      RECT  52.4 141.9 68.6 141.3 ;
      RECT  52.4 161.9 68.6 161.3 ;
      RECT  32.2 181.9 31.4 182.7 ;
      RECT  34.2 181.9 33.4 182.7 ;
      RECT  32.2 165.3 31.4 166.1 ;
      RECT  34.2 165.3 33.4 166.1 ;
      RECT  33.8 173.6 33.0 174.4 ;
      RECT  31.8 173.7 31.2 174.3 ;
      RECT  35.4 183.7 28.8 184.3 ;
      RECT  35.4 164.1 28.8 164.7 ;
      RECT  25.6 181.9 24.8 182.7 ;
      RECT  27.6 181.9 26.8 182.7 ;
      RECT  25.6 165.3 24.8 166.1 ;
      RECT  27.6 165.3 26.8 166.1 ;
      RECT  27.2 173.6 26.4 174.4 ;
      RECT  25.2 173.7 24.6 174.3 ;
      RECT  28.8 183.7 22.2 184.3 ;
      RECT  28.8 164.1 22.2 164.7 ;
      RECT  19.0 181.9 18.2 182.7 ;
      RECT  21.0 181.9 20.2 182.7 ;
      RECT  19.0 165.3 18.2 166.1 ;
      RECT  21.0 165.3 20.2 166.1 ;
      RECT  20.6 173.6 19.8 174.4 ;
      RECT  18.6 173.7 18.0 174.3 ;
      RECT  22.2 183.7 15.6 184.3 ;
      RECT  22.2 164.1 15.6 164.7 ;
      RECT  12.4 181.9 11.6 182.7 ;
      RECT  14.4 181.9 13.6 182.7 ;
      RECT  12.4 165.3 11.6 166.1 ;
      RECT  14.4 165.3 13.6 166.1 ;
      RECT  14.0 173.6 13.2 174.4 ;
      RECT  12.0 173.7 11.4 174.3 ;
      RECT  15.6 183.7 9.0 184.3 ;
      RECT  15.6 164.1 9.0 164.7 ;
      RECT  5.8 181.9 5.0 182.7 ;
      RECT  7.8 181.9 7.0 182.7 ;
      RECT  5.8 165.3 5.0 166.1 ;
      RECT  7.8 165.3 7.0 166.1 ;
      RECT  7.4 173.6 6.6 174.4 ;
      RECT  5.4 173.7 4.8 174.3 ;
      RECT  9.0 183.7 2.4 184.3 ;
      RECT  9.0 164.1 2.4 164.7 ;
      RECT  32.2 186.1 31.4 185.3 ;
      RECT  34.2 186.1 33.4 185.3 ;
      RECT  32.2 202.7 31.4 201.9 ;
      RECT  34.2 202.7 33.4 201.9 ;
      RECT  33.8 194.4 33.0 193.6 ;
      RECT  31.8 194.3 31.2 193.7 ;
      RECT  35.4 184.3 28.8 183.7 ;
      RECT  35.4 203.9 28.8 203.3 ;
      RECT  25.6 186.1 24.8 185.3 ;
      RECT  27.6 186.1 26.8 185.3 ;
      RECT  25.6 202.7 24.8 201.9 ;
      RECT  27.6 202.7 26.8 201.9 ;
      RECT  27.2 194.4 26.4 193.6 ;
      RECT  25.2 194.3 24.6 193.7 ;
      RECT  28.8 184.3 22.2 183.7 ;
      RECT  28.8 203.9 22.2 203.3 ;
      RECT  19.0 186.1 18.2 185.3 ;
      RECT  21.0 186.1 20.2 185.3 ;
      RECT  19.0 202.7 18.2 201.9 ;
      RECT  21.0 202.7 20.2 201.9 ;
      RECT  20.6 194.4 19.8 193.6 ;
      RECT  18.6 194.3 18.0 193.7 ;
      RECT  22.2 184.3 15.6 183.7 ;
      RECT  22.2 203.9 15.6 203.3 ;
      RECT  12.4 186.1 11.6 185.3 ;
      RECT  14.4 186.1 13.6 185.3 ;
      RECT  12.4 202.7 11.6 201.9 ;
      RECT  14.4 202.7 13.6 201.9 ;
      RECT  14.0 194.4 13.2 193.6 ;
      RECT  12.0 194.3 11.4 193.7 ;
      RECT  15.6 184.3 9.0 183.7 ;
      RECT  15.6 203.9 9.0 203.3 ;
      RECT  5.8 186.1 5.0 185.3 ;
      RECT  7.8 186.1 7.0 185.3 ;
      RECT  5.8 202.7 5.0 201.9 ;
      RECT  7.8 202.7 7.0 201.9 ;
      RECT  7.4 194.4 6.6 193.6 ;
      RECT  5.4 194.3 4.8 193.7 ;
      RECT  9.0 184.3 2.4 183.7 ;
      RECT  9.0 203.9 2.4 203.3 ;
      RECT  32.2 221.1 31.4 221.9 ;
      RECT  34.2 221.1 33.4 221.9 ;
      RECT  32.2 204.5 31.4 205.3 ;
      RECT  34.2 204.5 33.4 205.3 ;
      RECT  33.8 212.8 33.0 213.6 ;
      RECT  31.8 212.9 31.2 213.5 ;
      RECT  35.4 222.9 28.8 223.5 ;
      RECT  35.4 203.3 28.8 203.9 ;
      RECT  25.6 221.1 24.8 221.9 ;
      RECT  27.6 221.1 26.8 221.9 ;
      RECT  25.6 204.5 24.8 205.3 ;
      RECT  27.6 204.5 26.8 205.3 ;
      RECT  27.2 212.8 26.4 213.6 ;
      RECT  25.2 212.9 24.6 213.5 ;
      RECT  28.8 222.9 22.2 223.5 ;
      RECT  28.8 203.3 22.2 203.9 ;
      RECT  19.0 221.1 18.2 221.9 ;
      RECT  21.0 221.1 20.2 221.9 ;
      RECT  19.0 204.5 18.2 205.3 ;
      RECT  21.0 204.5 20.2 205.3 ;
      RECT  20.6 212.8 19.8 213.6 ;
      RECT  18.6 212.9 18.0 213.5 ;
      RECT  22.2 222.9 15.6 223.5 ;
      RECT  22.2 203.3 15.6 203.9 ;
      RECT  12.4 221.1 11.6 221.9 ;
      RECT  14.4 221.1 13.6 221.9 ;
      RECT  12.4 204.5 11.6 205.3 ;
      RECT  14.4 204.5 13.6 205.3 ;
      RECT  14.0 212.8 13.2 213.6 ;
      RECT  12.0 212.9 11.4 213.5 ;
      RECT  15.6 222.9 9.0 223.5 ;
      RECT  15.6 203.3 9.0 203.9 ;
      RECT  5.8 221.1 5.0 221.9 ;
      RECT  7.8 221.1 7.0 221.9 ;
      RECT  5.8 204.5 5.0 205.3 ;
      RECT  7.8 204.5 7.0 205.3 ;
      RECT  7.4 212.8 6.6 213.6 ;
      RECT  5.4 212.9 4.8 213.5 ;
      RECT  9.0 222.9 2.4 223.5 ;
      RECT  9.0 203.3 2.4 203.9 ;
      RECT  32.2 225.3 31.4 224.5 ;
      RECT  34.2 225.3 33.4 224.5 ;
      RECT  32.2 241.9 31.4 241.1 ;
      RECT  34.2 241.9 33.4 241.1 ;
      RECT  33.8 233.6 33.0 232.8 ;
      RECT  31.8 233.5 31.2 232.9 ;
      RECT  35.4 223.5 28.8 222.9 ;
      RECT  35.4 243.1 28.8 242.5 ;
      RECT  25.6 225.3 24.8 224.5 ;
      RECT  27.6 225.3 26.8 224.5 ;
      RECT  25.6 241.9 24.8 241.1 ;
      RECT  27.6 241.9 26.8 241.1 ;
      RECT  27.2 233.6 26.4 232.8 ;
      RECT  25.2 233.5 24.6 232.9 ;
      RECT  28.8 223.5 22.2 222.9 ;
      RECT  28.8 243.1 22.2 242.5 ;
      RECT  19.0 225.3 18.2 224.5 ;
      RECT  21.0 225.3 20.2 224.5 ;
      RECT  19.0 241.9 18.2 241.1 ;
      RECT  21.0 241.9 20.2 241.1 ;
      RECT  20.6 233.6 19.8 232.8 ;
      RECT  18.6 233.5 18.0 232.9 ;
      RECT  22.2 223.5 15.6 222.9 ;
      RECT  22.2 243.1 15.6 242.5 ;
      RECT  12.4 225.3 11.6 224.5 ;
      RECT  14.4 225.3 13.6 224.5 ;
      RECT  12.4 241.9 11.6 241.1 ;
      RECT  14.4 241.9 13.6 241.1 ;
      RECT  14.0 233.6 13.2 232.8 ;
      RECT  12.0 233.5 11.4 232.9 ;
      RECT  15.6 223.5 9.0 222.9 ;
      RECT  15.6 243.1 9.0 242.5 ;
      RECT  5.8 225.3 5.0 224.5 ;
      RECT  7.8 225.3 7.0 224.5 ;
      RECT  5.8 241.9 5.0 241.1 ;
      RECT  7.8 241.9 7.0 241.1 ;
      RECT  7.4 233.6 6.6 232.8 ;
      RECT  5.4 233.5 4.8 232.9 ;
      RECT  9.0 223.5 2.4 222.9 ;
      RECT  9.0 243.1 2.4 242.5 ;
      RECT  32.2 260.3 31.4 261.1 ;
      RECT  34.2 260.3 33.4 261.1 ;
      RECT  32.2 243.7 31.4 244.5 ;
      RECT  34.2 243.7 33.4 244.5 ;
      RECT  33.8 252.0 33.0 252.8 ;
      RECT  31.8 252.1 31.2 252.7 ;
      RECT  35.4 262.1 28.8 262.7 ;
      RECT  35.4 242.5 28.8 243.1 ;
      RECT  25.6 260.3 24.8 261.1 ;
      RECT  27.6 260.3 26.8 261.1 ;
      RECT  25.6 243.7 24.8 244.5 ;
      RECT  27.6 243.7 26.8 244.5 ;
      RECT  27.2 252.0 26.4 252.8 ;
      RECT  25.2 252.1 24.6 252.7 ;
      RECT  28.8 262.1 22.2 262.7 ;
      RECT  28.8 242.5 22.2 243.1 ;
      RECT  19.0 260.3 18.2 261.1 ;
      RECT  21.0 260.3 20.2 261.1 ;
      RECT  19.0 243.7 18.2 244.5 ;
      RECT  21.0 243.7 20.2 244.5 ;
      RECT  20.6 252.0 19.8 252.8 ;
      RECT  18.6 252.1 18.0 252.7 ;
      RECT  22.2 262.1 15.6 262.7 ;
      RECT  22.2 242.5 15.6 243.1 ;
      RECT  12.4 260.3 11.6 261.1 ;
      RECT  14.4 260.3 13.6 261.1 ;
      RECT  12.4 243.7 11.6 244.5 ;
      RECT  14.4 243.7 13.6 244.5 ;
      RECT  14.0 252.0 13.2 252.8 ;
      RECT  12.0 252.1 11.4 252.7 ;
      RECT  15.6 262.1 9.0 262.7 ;
      RECT  15.6 242.5 9.0 243.1 ;
      RECT  5.8 260.3 5.0 261.1 ;
      RECT  7.8 260.3 7.0 261.1 ;
      RECT  5.8 243.7 5.0 244.5 ;
      RECT  7.8 243.7 7.0 244.5 ;
      RECT  7.4 252.0 6.6 252.8 ;
      RECT  5.4 252.1 4.8 252.7 ;
      RECT  9.0 262.1 2.4 262.7 ;
      RECT  9.0 242.5 2.4 243.1 ;
      RECT  32.2 264.5 31.4 263.7 ;
      RECT  34.2 264.5 33.4 263.7 ;
      RECT  32.2 281.1 31.4 280.3 ;
      RECT  34.2 281.1 33.4 280.3 ;
      RECT  33.8 272.8 33.0 272.0 ;
      RECT  31.8 272.7 31.2 272.1 ;
      RECT  35.4 262.7 28.8 262.1 ;
      RECT  35.4 282.3 28.8 281.7 ;
      RECT  25.6 264.5 24.8 263.7 ;
      RECT  27.6 264.5 26.8 263.7 ;
      RECT  25.6 281.1 24.8 280.3 ;
      RECT  27.6 281.1 26.8 280.3 ;
      RECT  27.2 272.8 26.4 272.0 ;
      RECT  25.2 272.7 24.6 272.1 ;
      RECT  28.8 262.7 22.2 262.1 ;
      RECT  28.8 282.3 22.2 281.7 ;
      RECT  19.0 264.5 18.2 263.7 ;
      RECT  21.0 264.5 20.2 263.7 ;
      RECT  19.0 281.1 18.2 280.3 ;
      RECT  21.0 281.1 20.2 280.3 ;
      RECT  20.6 272.8 19.8 272.0 ;
      RECT  18.6 272.7 18.0 272.1 ;
      RECT  22.2 262.7 15.6 262.1 ;
      RECT  22.2 282.3 15.6 281.7 ;
      RECT  12.4 264.5 11.6 263.7 ;
      RECT  14.4 264.5 13.6 263.7 ;
      RECT  12.4 281.1 11.6 280.3 ;
      RECT  14.4 281.1 13.6 280.3 ;
      RECT  14.0 272.8 13.2 272.0 ;
      RECT  12.0 272.7 11.4 272.1 ;
      RECT  15.6 262.7 9.0 262.1 ;
      RECT  15.6 282.3 9.0 281.7 ;
      RECT  5.8 264.5 5.0 263.7 ;
      RECT  7.8 264.5 7.0 263.7 ;
      RECT  5.8 281.1 5.0 280.3 ;
      RECT  7.8 281.1 7.0 280.3 ;
      RECT  7.4 272.8 6.6 272.0 ;
      RECT  5.4 272.7 4.8 272.1 ;
      RECT  9.0 262.7 2.4 262.1 ;
      RECT  9.0 282.3 2.4 281.7 ;
      RECT  32.2 299.5 31.4 300.3 ;
      RECT  34.2 299.5 33.4 300.3 ;
      RECT  32.2 282.9 31.4 283.7 ;
      RECT  34.2 282.9 33.4 283.7 ;
      RECT  33.8 291.2 33.0 292.0 ;
      RECT  31.8 291.3 31.2 291.9 ;
      RECT  35.4 301.3 28.8 301.9 ;
      RECT  35.4 281.7 28.8 282.3 ;
      RECT  25.6 299.5 24.8 300.3 ;
      RECT  27.6 299.5 26.8 300.3 ;
      RECT  25.6 282.9 24.8 283.7 ;
      RECT  27.6 282.9 26.8 283.7 ;
      RECT  27.2 291.2 26.4 292.0 ;
      RECT  25.2 291.3 24.6 291.9 ;
      RECT  28.8 301.3 22.2 301.9 ;
      RECT  28.8 281.7 22.2 282.3 ;
      RECT  19.0 299.5 18.2 300.3 ;
      RECT  21.0 299.5 20.2 300.3 ;
      RECT  19.0 282.9 18.2 283.7 ;
      RECT  21.0 282.9 20.2 283.7 ;
      RECT  20.6 291.2 19.8 292.0 ;
      RECT  18.6 291.3 18.0 291.9 ;
      RECT  22.2 301.3 15.6 301.9 ;
      RECT  22.2 281.7 15.6 282.3 ;
      RECT  12.4 299.5 11.6 300.3 ;
      RECT  14.4 299.5 13.6 300.3 ;
      RECT  12.4 282.9 11.6 283.7 ;
      RECT  14.4 282.9 13.6 283.7 ;
      RECT  14.0 291.2 13.2 292.0 ;
      RECT  12.0 291.3 11.4 291.9 ;
      RECT  15.6 301.3 9.0 301.9 ;
      RECT  15.6 281.7 9.0 282.3 ;
      RECT  5.8 299.5 5.0 300.3 ;
      RECT  7.8 299.5 7.0 300.3 ;
      RECT  5.8 282.9 5.0 283.7 ;
      RECT  7.8 282.9 7.0 283.7 ;
      RECT  7.4 291.2 6.6 292.0 ;
      RECT  5.4 291.3 4.8 291.9 ;
      RECT  9.0 301.3 2.4 301.9 ;
      RECT  9.0 281.7 2.4 282.3 ;
      RECT  32.2 303.7 31.4 302.9 ;
      RECT  34.2 303.7 33.4 302.9 ;
      RECT  32.2 320.3 31.4 319.5 ;
      RECT  34.2 320.3 33.4 319.5 ;
      RECT  33.8 312.0 33.0 311.2 ;
      RECT  31.8 311.9 31.2 311.3 ;
      RECT  35.4 301.9 28.8 301.3 ;
      RECT  35.4 321.5 28.8 320.9 ;
      RECT  25.6 303.7 24.8 302.9 ;
      RECT  27.6 303.7 26.8 302.9 ;
      RECT  25.6 320.3 24.8 319.5 ;
      RECT  27.6 320.3 26.8 319.5 ;
      RECT  27.2 312.0 26.4 311.2 ;
      RECT  25.2 311.9 24.6 311.3 ;
      RECT  28.8 301.9 22.2 301.3 ;
      RECT  28.8 321.5 22.2 320.9 ;
      RECT  19.0 303.7 18.2 302.9 ;
      RECT  21.0 303.7 20.2 302.9 ;
      RECT  19.0 320.3 18.2 319.5 ;
      RECT  21.0 320.3 20.2 319.5 ;
      RECT  20.6 312.0 19.8 311.2 ;
      RECT  18.6 311.9 18.0 311.3 ;
      RECT  22.2 301.9 15.6 301.3 ;
      RECT  22.2 321.5 15.6 320.9 ;
      RECT  12.4 303.7 11.6 302.9 ;
      RECT  14.4 303.7 13.6 302.9 ;
      RECT  12.4 320.3 11.6 319.5 ;
      RECT  14.4 320.3 13.6 319.5 ;
      RECT  14.0 312.0 13.2 311.2 ;
      RECT  12.0 311.9 11.4 311.3 ;
      RECT  15.6 301.9 9.0 301.3 ;
      RECT  15.6 321.5 9.0 320.9 ;
      RECT  5.8 303.7 5.0 302.9 ;
      RECT  7.8 303.7 7.0 302.9 ;
      RECT  5.8 320.3 5.0 319.5 ;
      RECT  7.8 320.3 7.0 319.5 ;
      RECT  7.4 312.0 6.6 311.2 ;
      RECT  5.4 311.9 4.8 311.3 ;
      RECT  9.0 301.9 2.4 301.3 ;
      RECT  9.0 321.5 2.4 320.9 ;
      RECT  32.2 338.7 31.4 339.5 ;
      RECT  34.2 338.7 33.4 339.5 ;
      RECT  32.2 322.1 31.4 322.9 ;
      RECT  34.2 322.1 33.4 322.9 ;
      RECT  33.8 330.4 33.0 331.2 ;
      RECT  31.8 330.5 31.2 331.1 ;
      RECT  35.4 340.5 28.8 341.1 ;
      RECT  35.4 320.9 28.8 321.5 ;
      RECT  25.6 338.7 24.8 339.5 ;
      RECT  27.6 338.7 26.8 339.5 ;
      RECT  25.6 322.1 24.8 322.9 ;
      RECT  27.6 322.1 26.8 322.9 ;
      RECT  27.2 330.4 26.4 331.2 ;
      RECT  25.2 330.5 24.6 331.1 ;
      RECT  28.8 340.5 22.2 341.1 ;
      RECT  28.8 320.9 22.2 321.5 ;
      RECT  19.0 338.7 18.2 339.5 ;
      RECT  21.0 338.7 20.2 339.5 ;
      RECT  19.0 322.1 18.2 322.9 ;
      RECT  21.0 322.1 20.2 322.9 ;
      RECT  20.6 330.4 19.8 331.2 ;
      RECT  18.6 330.5 18.0 331.1 ;
      RECT  22.2 340.5 15.6 341.1 ;
      RECT  22.2 320.9 15.6 321.5 ;
      RECT  12.4 338.7 11.6 339.5 ;
      RECT  14.4 338.7 13.6 339.5 ;
      RECT  12.4 322.1 11.6 322.9 ;
      RECT  14.4 322.1 13.6 322.9 ;
      RECT  14.0 330.4 13.2 331.2 ;
      RECT  12.0 330.5 11.4 331.1 ;
      RECT  15.6 340.5 9.0 341.1 ;
      RECT  15.6 320.9 9.0 321.5 ;
      RECT  5.8 338.7 5.0 339.5 ;
      RECT  7.8 338.7 7.0 339.5 ;
      RECT  5.8 322.1 5.0 322.9 ;
      RECT  7.8 322.1 7.0 322.9 ;
      RECT  7.4 330.4 6.6 331.2 ;
      RECT  5.4 330.5 4.8 331.1 ;
      RECT  9.0 340.5 2.4 341.1 ;
      RECT  9.0 320.9 2.4 321.5 ;
      RECT  55.6 103.7 56.4 102.9 ;
      RECT  53.6 103.7 54.4 102.9 ;
      RECT  57.6 103.7 58.4 102.9 ;
      RECT  55.6 103.7 56.4 102.9 ;
      RECT  53.6 120.3 54.4 119.5 ;
      RECT  57.6 120.3 58.4 119.5 ;
      RECT  54.6 118.8 55.4 118.0 ;
      RECT  56.6 116.0 57.4 115.2 ;
      RECT  59.1 105.0 59.7 104.4 ;
      RECT  52.4 101.9 61.0 101.3 ;
      RECT  52.4 121.9 61.0 121.3 ;
      RECT  64.2 103.7 65.0 102.9 ;
      RECT  62.2 103.7 63.0 102.9 ;
      RECT  64.2 120.7 65.0 119.9 ;
      RECT  62.2 120.7 63.0 119.9 ;
      RECT  62.6 112.2 63.4 111.4 ;
      RECT  64.6 112.1 65.2 111.5 ;
      RECT  61.0 101.9 67.6 101.3 ;
      RECT  61.0 121.9 67.6 121.3 ;
      RECT  70.8 103.7 71.6 102.9 ;
      RECT  68.8 103.7 69.6 102.9 ;
      RECT  70.8 120.7 71.6 119.9 ;
      RECT  68.8 120.7 69.6 119.9 ;
      RECT  69.2 112.2 70.0 111.4 ;
      RECT  71.2 112.1 71.8 111.5 ;
      RECT  67.6 101.9 72.8 101.3 ;
      RECT  67.6 121.9 72.8 121.3 ;
      RECT  62.6 112.2 63.4 111.4 ;
      RECT  71.2 112.1 71.8 111.5 ;
      RECT  61.0 101.9 72.8 101.3 ;
      RECT  61.0 121.9 72.8 121.3 ;
      RECT  65.9 151.7 79.4 152.3 ;
      RECT  65.7 90.3 79.4 90.9 ;
      RECT  71.5 111.5 79.4 112.1 ;
      RECT  73.3 72.3 79.4 72.9 ;
      RECT  74.8 10.3 79.4 10.9 ;
      RECT  71.6 351.6 72.4 351.8 ;
      RECT  58.8 344.8 59.6 349.6 ;
      RECT  67.6 357.8 68.2 358.4 ;
      RECT  65.4 357.2 69.0 357.8 ;
      RECT  58.8 353.4 64.4 353.6 ;
      RECT  59.6 350.4 70.6 351.0 ;
      RECT  76.4 353.8 77.2 362.4 ;
      RECT  67.6 346.8 68.2 347.4 ;
      RECT  63.2 344.8 64.0 346.2 ;
      RECT  65.4 357.0 66.2 357.2 ;
      RECT  71.6 357.6 72.4 358.4 ;
      RECT  68.0 354.4 68.6 355.6 ;
      RECT  62.0 358.4 64.0 359.0 ;
      RECT  69.2 344.2 70.0 346.8 ;
      RECT  65.4 347.4 68.2 348.0 ;
      RECT  62.0 346.2 64.0 346.8 ;
      RECT  76.4 349.8 77.2 353.2 ;
      RECT  71.8 358.4 73.0 362.4 ;
      RECT  60.4 354.6 61.2 363.0 ;
      RECT  62.0 355.0 67.4 355.6 ;
      RECT  70.0 351.0 70.6 354.2 ;
      RECT  57.6 363.0 79.4 364.2 ;
      RECT  73.0 353.2 77.2 353.8 ;
      RECT  74.8 354.4 75.6 363.0 ;
      RECT  78.0 344.2 78.8 345.6 ;
      RECT  71.8 354.8 72.4 355.8 ;
      RECT  70.0 354.2 72.4 354.8 ;
      RECT  58.8 354.0 59.6 362.4 ;
      RECT  71.6 346.2 73.0 346.8 ;
      RECT  68.0 355.6 70.2 356.2 ;
      RECT  63.2 359.0 64.0 362.4 ;
      RECT  61.0 352.2 66.0 352.8 ;
      RECT  78.0 361.4 78.8 363.0 ;
      RECT  71.6 351.8 75.4 352.4 ;
      RECT  71.6 346.8 72.4 347.6 ;
      RECT  57.6 343.0 79.4 344.2 ;
      RECT  65.2 352.8 66.0 353.0 ;
      RECT  62.6 351.0 63.4 351.2 ;
      RECT  68.2 357.0 69.0 357.2 ;
      RECT  76.4 344.8 77.2 349.2 ;
      RECT  59.6 350.2 61.2 350.4 ;
      RECT  62.0 357.6 62.8 358.4 ;
      RECT  67.6 344.8 68.4 346.8 ;
      RECT  61.0 352.0 61.8 352.2 ;
      RECT  62.0 355.6 62.8 355.8 ;
      RECT  73.4 349.0 74.2 349.2 ;
      RECT  63.6 347.4 64.4 348.2 ;
      RECT  74.8 344.2 75.6 348.6 ;
      RECT  69.4 355.4 70.2 355.6 ;
      RECT  65.8 344.2 66.8 346.8 ;
      RECT  63.8 348.2 64.4 350.4 ;
      RECT  69.2 358.4 70.0 363.0 ;
      RECT  66.0 358.4 66.8 363.0 ;
      RECT  69.4 350.2 70.2 350.4 ;
      RECT  63.8 354.0 68.6 354.4 ;
      RECT  58.8 353.6 64.6 353.8 ;
      RECT  67.6 358.4 68.4 362.4 ;
      RECT  74.6 352.4 75.4 352.6 ;
      RECT  58.8 353.8 68.6 354.0 ;
      RECT  66.6 355.6 67.4 355.8 ;
      RECT  71.8 344.8 73.0 346.2 ;
      RECT  65.4 348.0 66.2 348.2 ;
      RECT  71.8 355.8 73.2 356.6 ;
      RECT  73.0 353.0 73.8 353.2 ;
      RECT  62.0 346.8 62.8 347.6 ;
      RECT  60.4 344.2 61.2 348.8 ;
      RECT  73.4 349.2 77.2 349.8 ;
      RECT  71.6 375.6 72.4 375.4 ;
      RECT  58.8 382.4 59.6 377.6 ;
      RECT  67.6 369.4 68.2 368.8 ;
      RECT  65.4 370.0 69.0 369.4 ;
      RECT  58.8 373.8 64.4 373.6 ;
      RECT  59.6 376.8 70.6 376.2 ;
      RECT  76.4 373.4 77.2 364.8 ;
      RECT  67.6 380.4 68.2 379.8 ;
      RECT  63.2 382.4 64.0 381.0 ;
      RECT  65.4 370.2 66.2 370.0 ;
      RECT  71.6 369.6 72.4 368.8 ;
      RECT  68.0 372.8 68.6 371.6 ;
      RECT  62.0 368.8 64.0 368.2 ;
      RECT  69.2 383.0 70.0 380.4 ;
      RECT  65.4 379.8 68.2 379.2 ;
      RECT  62.0 381.0 64.0 380.4 ;
      RECT  76.4 377.4 77.2 374.0 ;
      RECT  71.8 368.8 73.0 364.8 ;
      RECT  60.4 372.6 61.2 364.2 ;
      RECT  62.0 372.2 67.4 371.6 ;
      RECT  70.0 376.2 70.6 373.0 ;
      RECT  57.6 364.2 79.4 363.0 ;
      RECT  73.0 374.0 77.2 373.4 ;
      RECT  74.8 372.8 75.6 364.2 ;
      RECT  78.0 383.0 78.8 381.6 ;
      RECT  71.8 372.4 72.4 371.4 ;
      RECT  70.0 373.0 72.4 372.4 ;
      RECT  58.8 373.2 59.6 364.8 ;
      RECT  71.6 381.0 73.0 380.4 ;
      RECT  68.0 371.6 70.2 371.0 ;
      RECT  63.2 368.2 64.0 364.8 ;
      RECT  61.0 375.0 66.0 374.4 ;
      RECT  78.0 365.8 78.8 364.2 ;
      RECT  71.6 375.4 75.4 374.8 ;
      RECT  71.6 380.4 72.4 379.6 ;
      RECT  57.6 384.2 79.4 383.0 ;
      RECT  65.2 374.4 66.0 374.2 ;
      RECT  62.6 376.2 63.4 376.0 ;
      RECT  68.2 370.2 69.0 370.0 ;
      RECT  76.4 382.4 77.2 378.0 ;
      RECT  59.6 377.0 61.2 376.8 ;
      RECT  62.0 369.6 62.8 368.8 ;
      RECT  67.6 382.4 68.4 380.4 ;
      RECT  61.0 375.2 61.8 375.0 ;
      RECT  62.0 371.6 62.8 371.4 ;
      RECT  73.4 378.2 74.2 378.0 ;
      RECT  63.6 379.8 64.4 379.0 ;
      RECT  74.8 383.0 75.6 378.6 ;
      RECT  69.4 371.8 70.2 371.6 ;
      RECT  65.8 383.0 66.8 380.4 ;
      RECT  63.8 379.0 64.4 376.8 ;
      RECT  69.2 368.8 70.0 364.2 ;
      RECT  66.0 368.8 66.8 364.2 ;
      RECT  69.4 377.0 70.2 376.8 ;
      RECT  63.8 373.2 68.6 372.8 ;
      RECT  58.8 373.6 64.6 373.4 ;
      RECT  67.6 368.8 68.4 364.8 ;
      RECT  74.6 374.8 75.4 374.6 ;
      RECT  58.8 373.4 68.6 373.2 ;
      RECT  66.6 371.6 67.4 371.4 ;
      RECT  71.8 382.4 73.0 381.0 ;
      RECT  65.4 379.2 66.2 379.0 ;
      RECT  71.8 371.4 73.2 370.6 ;
      RECT  73.0 374.2 73.8 374.0 ;
      RECT  62.0 380.4 62.8 379.6 ;
      RECT  60.4 383.0 61.2 378.4 ;
      RECT  73.4 378.0 77.2 377.4 ;
      RECT  71.6 391.6 72.4 391.8 ;
      RECT  58.8 384.8 59.6 389.6 ;
      RECT  67.6 397.8 68.2 398.4 ;
      RECT  65.4 397.2 69.0 397.8 ;
      RECT  58.8 393.4 64.4 393.6 ;
      RECT  59.6 390.4 70.6 391.0 ;
      RECT  76.4 393.8 77.2 402.4 ;
      RECT  67.6 386.8 68.2 387.4 ;
      RECT  63.2 384.8 64.0 386.2 ;
      RECT  65.4 397.0 66.2 397.2 ;
      RECT  71.6 397.6 72.4 398.4 ;
      RECT  68.0 394.4 68.6 395.6 ;
      RECT  62.0 398.4 64.0 399.0 ;
      RECT  69.2 384.2 70.0 386.8 ;
      RECT  65.4 387.4 68.2 388.0 ;
      RECT  62.0 386.2 64.0 386.8 ;
      RECT  76.4 389.8 77.2 393.2 ;
      RECT  71.8 398.4 73.0 402.4 ;
      RECT  60.4 394.6 61.2 403.0 ;
      RECT  62.0 395.0 67.4 395.6 ;
      RECT  70.0 391.0 70.6 394.2 ;
      RECT  57.6 403.0 79.4 404.2 ;
      RECT  73.0 393.2 77.2 393.8 ;
      RECT  74.8 394.4 75.6 403.0 ;
      RECT  78.0 384.2 78.8 385.6 ;
      RECT  71.8 394.8 72.4 395.8 ;
      RECT  70.0 394.2 72.4 394.8 ;
      RECT  58.8 394.0 59.6 402.4 ;
      RECT  71.6 386.2 73.0 386.8 ;
      RECT  68.0 395.6 70.2 396.2 ;
      RECT  63.2 399.0 64.0 402.4 ;
      RECT  61.0 392.2 66.0 392.8 ;
      RECT  78.0 401.4 78.8 403.0 ;
      RECT  71.6 391.8 75.4 392.4 ;
      RECT  71.6 386.8 72.4 387.6 ;
      RECT  57.6 383.0 79.4 384.2 ;
      RECT  65.2 392.8 66.0 393.0 ;
      RECT  62.6 391.0 63.4 391.2 ;
      RECT  68.2 397.0 69.0 397.2 ;
      RECT  76.4 384.8 77.2 389.2 ;
      RECT  59.6 390.2 61.2 390.4 ;
      RECT  62.0 397.6 62.8 398.4 ;
      RECT  67.6 384.8 68.4 386.8 ;
      RECT  61.0 392.0 61.8 392.2 ;
      RECT  62.0 395.6 62.8 395.8 ;
      RECT  73.4 389.0 74.2 389.2 ;
      RECT  63.6 387.4 64.4 388.2 ;
      RECT  74.8 384.2 75.6 388.6 ;
      RECT  69.4 395.4 70.2 395.6 ;
      RECT  65.8 384.2 66.8 386.8 ;
      RECT  63.8 388.2 64.4 390.4 ;
      RECT  69.2 398.4 70.0 403.0 ;
      RECT  66.0 398.4 66.8 403.0 ;
      RECT  69.4 390.2 70.2 390.4 ;
      RECT  63.8 394.0 68.6 394.4 ;
      RECT  58.8 393.6 64.6 393.8 ;
      RECT  67.6 398.4 68.4 402.4 ;
      RECT  74.6 392.4 75.4 392.6 ;
      RECT  58.8 393.8 68.6 394.0 ;
      RECT  66.6 395.6 67.4 395.8 ;
      RECT  71.8 384.8 73.0 386.2 ;
      RECT  65.4 388.0 66.2 388.2 ;
      RECT  71.8 395.8 73.2 396.6 ;
      RECT  73.0 393.0 73.8 393.2 ;
      RECT  62.0 386.8 62.8 387.6 ;
      RECT  60.4 384.2 61.2 388.8 ;
      RECT  73.4 389.2 77.2 389.8 ;
      RECT  71.6 415.6 72.4 415.4 ;
      RECT  58.8 422.4 59.6 417.6 ;
      RECT  67.6 409.4 68.2 408.8 ;
      RECT  65.4 410.0 69.0 409.4 ;
      RECT  58.8 413.8 64.4 413.6 ;
      RECT  59.6 416.8 70.6 416.2 ;
      RECT  76.4 413.4 77.2 404.8 ;
      RECT  67.6 420.4 68.2 419.8 ;
      RECT  63.2 422.4 64.0 421.0 ;
      RECT  65.4 410.2 66.2 410.0 ;
      RECT  71.6 409.6 72.4 408.8 ;
      RECT  68.0 412.8 68.6 411.6 ;
      RECT  62.0 408.8 64.0 408.2 ;
      RECT  69.2 423.0 70.0 420.4 ;
      RECT  65.4 419.8 68.2 419.2 ;
      RECT  62.0 421.0 64.0 420.4 ;
      RECT  76.4 417.4 77.2 414.0 ;
      RECT  71.8 408.8 73.0 404.8 ;
      RECT  60.4 412.6 61.2 404.2 ;
      RECT  62.0 412.2 67.4 411.6 ;
      RECT  70.0 416.2 70.6 413.0 ;
      RECT  57.6 404.2 79.4 403.0 ;
      RECT  73.0 414.0 77.2 413.4 ;
      RECT  74.8 412.8 75.6 404.2 ;
      RECT  78.0 423.0 78.8 421.6 ;
      RECT  71.8 412.4 72.4 411.4 ;
      RECT  70.0 413.0 72.4 412.4 ;
      RECT  58.8 413.2 59.6 404.8 ;
      RECT  71.6 421.0 73.0 420.4 ;
      RECT  68.0 411.6 70.2 411.0 ;
      RECT  63.2 408.2 64.0 404.8 ;
      RECT  61.0 415.0 66.0 414.4 ;
      RECT  78.0 405.8 78.8 404.2 ;
      RECT  71.6 415.4 75.4 414.8 ;
      RECT  71.6 420.4 72.4 419.6 ;
      RECT  57.6 424.2 79.4 423.0 ;
      RECT  65.2 414.4 66.0 414.2 ;
      RECT  62.6 416.2 63.4 416.0 ;
      RECT  68.2 410.2 69.0 410.0 ;
      RECT  76.4 422.4 77.2 418.0 ;
      RECT  59.6 417.0 61.2 416.8 ;
      RECT  62.0 409.6 62.8 408.8 ;
      RECT  67.6 422.4 68.4 420.4 ;
      RECT  61.0 415.2 61.8 415.0 ;
      RECT  62.0 411.6 62.8 411.4 ;
      RECT  73.4 418.2 74.2 418.0 ;
      RECT  63.6 419.8 64.4 419.0 ;
      RECT  74.8 423.0 75.6 418.6 ;
      RECT  69.4 411.8 70.2 411.6 ;
      RECT  65.8 423.0 66.8 420.4 ;
      RECT  63.8 419.0 64.4 416.8 ;
      RECT  69.2 408.8 70.0 404.2 ;
      RECT  66.0 408.8 66.8 404.2 ;
      RECT  69.4 417.0 70.2 416.8 ;
      RECT  63.8 413.2 68.6 412.8 ;
      RECT  58.8 413.6 64.6 413.4 ;
      RECT  67.6 408.8 68.4 404.8 ;
      RECT  74.6 414.8 75.4 414.6 ;
      RECT  58.8 413.4 68.6 413.2 ;
      RECT  66.6 411.6 67.4 411.4 ;
      RECT  71.8 422.4 73.0 421.0 ;
      RECT  65.4 419.2 66.2 419.0 ;
      RECT  71.8 411.4 73.2 410.6 ;
      RECT  73.0 414.2 73.8 414.0 ;
      RECT  62.0 420.4 62.8 419.6 ;
      RECT  60.4 423.0 61.2 418.4 ;
      RECT  73.4 418.0 77.2 417.4 ;
      RECT  187.3 56.0 188.1 56.2 ;
      RECT  174.5 49.2 175.3 54.0 ;
      RECT  183.3 62.2 183.9 62.8 ;
      RECT  181.1 61.6 184.7 62.2 ;
      RECT  174.5 57.8 180.1 58.0 ;
      RECT  175.3 54.8 186.3 55.4 ;
      RECT  192.1 58.2 192.9 66.8 ;
      RECT  183.3 51.2 183.9 51.8 ;
      RECT  178.9 49.2 179.7 50.6 ;
      RECT  181.1 61.4 181.9 61.6 ;
      RECT  187.3 62.0 188.1 62.8 ;
      RECT  183.7 58.8 184.3 60.0 ;
      RECT  177.7 62.8 179.7 63.4 ;
      RECT  184.9 48.6 185.7 51.2 ;
      RECT  181.1 51.8 183.9 52.4 ;
      RECT  177.7 50.6 179.7 51.2 ;
      RECT  192.1 54.2 192.9 57.6 ;
      RECT  187.5 62.8 188.7 66.8 ;
      RECT  176.1 59.0 176.9 67.4 ;
      RECT  177.7 59.4 183.1 60.0 ;
      RECT  185.7 55.4 186.3 58.6 ;
      RECT  173.3 67.4 195.1 68.6 ;
      RECT  188.7 57.6 192.9 58.2 ;
      RECT  190.5 58.8 191.3 67.4 ;
      RECT  193.7 48.6 194.5 50.0 ;
      RECT  187.5 59.2 188.1 60.2 ;
      RECT  185.7 58.6 188.1 59.2 ;
      RECT  174.5 58.4 175.3 66.8 ;
      RECT  187.3 50.6 188.7 51.2 ;
      RECT  183.7 60.0 185.9 60.6 ;
      RECT  178.9 63.4 179.7 66.8 ;
      RECT  176.7 56.6 181.7 57.2 ;
      RECT  193.7 65.8 194.5 67.4 ;
      RECT  187.3 56.2 191.1 56.8 ;
      RECT  187.3 51.2 188.1 52.0 ;
      RECT  173.3 47.4 195.1 48.6 ;
      RECT  180.9 57.2 181.7 57.4 ;
      RECT  178.3 55.4 179.1 55.6 ;
      RECT  183.9 61.4 184.7 61.6 ;
      RECT  192.1 49.2 192.9 53.6 ;
      RECT  175.3 54.6 176.9 54.8 ;
      RECT  177.7 62.0 178.5 62.8 ;
      RECT  183.3 49.2 184.1 51.2 ;
      RECT  176.7 56.4 177.5 56.6 ;
      RECT  177.7 60.0 178.5 60.2 ;
      RECT  189.1 53.4 189.9 53.6 ;
      RECT  179.3 51.8 180.1 52.6 ;
      RECT  190.5 48.6 191.3 53.0 ;
      RECT  185.1 59.8 185.9 60.0 ;
      RECT  181.5 48.6 182.5 51.2 ;
      RECT  179.5 52.6 180.1 54.8 ;
      RECT  184.9 62.8 185.7 67.4 ;
      RECT  181.7 62.8 182.5 67.4 ;
      RECT  185.1 54.6 185.9 54.8 ;
      RECT  179.5 58.4 184.3 58.8 ;
      RECT  174.5 58.0 180.3 58.2 ;
      RECT  183.3 62.8 184.1 66.8 ;
      RECT  190.3 56.8 191.1 57.0 ;
      RECT  174.5 58.2 184.3 58.4 ;
      RECT  182.3 60.0 183.1 60.2 ;
      RECT  187.5 49.2 188.7 50.6 ;
      RECT  181.1 52.4 181.9 52.6 ;
      RECT  187.5 60.2 188.9 61.0 ;
      RECT  188.7 57.4 189.5 57.6 ;
      RECT  177.7 51.2 178.5 52.0 ;
      RECT  176.1 48.6 176.9 53.2 ;
      RECT  189.1 53.6 192.9 54.2 ;
      RECT  209.1 56.0 209.9 56.2 ;
      RECT  196.3 49.2 197.1 54.0 ;
      RECT  205.1 62.2 205.7 62.8 ;
      RECT  202.9 61.6 206.5 62.2 ;
      RECT  196.3 57.8 201.9 58.0 ;
      RECT  197.1 54.8 208.1 55.4 ;
      RECT  213.9 58.2 214.7 66.8 ;
      RECT  205.1 51.2 205.7 51.8 ;
      RECT  200.7 49.2 201.5 50.6 ;
      RECT  202.9 61.4 203.7 61.6 ;
      RECT  209.1 62.0 209.9 62.8 ;
      RECT  205.5 58.8 206.1 60.0 ;
      RECT  199.5 62.8 201.5 63.4 ;
      RECT  206.7 48.6 207.5 51.2 ;
      RECT  202.9 51.8 205.7 52.4 ;
      RECT  199.5 50.6 201.5 51.2 ;
      RECT  213.9 54.2 214.7 57.6 ;
      RECT  209.3 62.8 210.5 66.8 ;
      RECT  197.9 59.0 198.7 67.4 ;
      RECT  199.5 59.4 204.9 60.0 ;
      RECT  207.5 55.4 208.1 58.6 ;
      RECT  195.1 67.4 216.9 68.6 ;
      RECT  210.5 57.6 214.7 58.2 ;
      RECT  212.3 58.8 213.1 67.4 ;
      RECT  215.5 48.6 216.3 50.0 ;
      RECT  209.3 59.2 209.9 60.2 ;
      RECT  207.5 58.6 209.9 59.2 ;
      RECT  196.3 58.4 197.1 66.8 ;
      RECT  209.1 50.6 210.5 51.2 ;
      RECT  205.5 60.0 207.7 60.6 ;
      RECT  200.7 63.4 201.5 66.8 ;
      RECT  198.5 56.6 203.5 57.2 ;
      RECT  215.5 65.8 216.3 67.4 ;
      RECT  209.1 56.2 212.9 56.8 ;
      RECT  209.1 51.2 209.9 52.0 ;
      RECT  195.1 47.4 216.9 48.6 ;
      RECT  202.7 57.2 203.5 57.4 ;
      RECT  200.1 55.4 200.9 55.6 ;
      RECT  205.7 61.4 206.5 61.6 ;
      RECT  213.9 49.2 214.7 53.6 ;
      RECT  197.1 54.6 198.7 54.8 ;
      RECT  199.5 62.0 200.3 62.8 ;
      RECT  205.1 49.2 205.9 51.2 ;
      RECT  198.5 56.4 199.3 56.6 ;
      RECT  199.5 60.0 200.3 60.2 ;
      RECT  210.9 53.4 211.7 53.6 ;
      RECT  201.1 51.8 201.9 52.6 ;
      RECT  212.3 48.6 213.1 53.0 ;
      RECT  206.9 59.8 207.7 60.0 ;
      RECT  203.3 48.6 204.3 51.2 ;
      RECT  201.3 52.6 201.9 54.8 ;
      RECT  206.7 62.8 207.5 67.4 ;
      RECT  203.5 62.8 204.3 67.4 ;
      RECT  206.9 54.6 207.7 54.8 ;
      RECT  201.3 58.4 206.1 58.8 ;
      RECT  196.3 58.0 202.1 58.2 ;
      RECT  205.1 62.8 205.9 66.8 ;
      RECT  212.1 56.8 212.9 57.0 ;
      RECT  196.3 58.2 206.1 58.4 ;
      RECT  204.1 60.0 204.9 60.2 ;
      RECT  209.3 49.2 210.5 50.6 ;
      RECT  202.9 52.4 203.7 52.6 ;
      RECT  209.3 60.2 210.7 61.0 ;
      RECT  210.5 57.4 211.3 57.6 ;
      RECT  199.5 51.2 200.3 52.0 ;
      RECT  197.9 48.6 198.7 53.2 ;
      RECT  210.9 53.6 214.7 54.2 ;
   LAYER  m2 ;
      RECT  189.9 203.6 190.7 204.4 ;
      RECT  186.5 193.6 187.3 204.4 ;
      RECT  191.7 195.2 192.5 204.4 ;
      RECT  188.1 193.6 188.9 204.4 ;
      RECT  190.9 194.4 192.5 195.2 ;
      RECT  193.3 193.6 194.1 204.4 ;
      RECT  191.7 193.6 192.5 194.4 ;
      RECT  189.9 204.4 190.7 203.6 ;
      RECT  186.5 214.4 187.3 203.6 ;
      RECT  191.7 212.8 192.5 203.6 ;
      RECT  188.1 214.4 188.9 203.6 ;
      RECT  190.9 213.6 192.5 212.8 ;
      RECT  193.3 214.4 194.1 203.6 ;
      RECT  191.7 214.4 192.5 213.6 ;
      RECT  189.9 224.4 190.7 225.2 ;
      RECT  186.5 214.4 187.3 225.2 ;
      RECT  191.7 216.0 192.5 225.2 ;
      RECT  188.1 214.4 188.9 225.2 ;
      RECT  190.9 215.2 192.5 216.0 ;
      RECT  193.3 214.4 194.1 225.2 ;
      RECT  191.7 214.4 192.5 215.2 ;
      RECT  189.9 225.2 190.7 224.4 ;
      RECT  186.5 235.2 187.3 224.4 ;
      RECT  191.7 233.6 192.5 224.4 ;
      RECT  188.1 235.2 188.9 224.4 ;
      RECT  190.9 234.4 192.5 233.6 ;
      RECT  193.3 235.2 194.1 224.4 ;
      RECT  191.7 235.2 192.5 234.4 ;
      RECT  189.9 245.2 190.7 246.0 ;
      RECT  186.5 235.2 187.3 246.0 ;
      RECT  191.7 236.8 192.5 246.0 ;
      RECT  188.1 235.2 188.9 246.0 ;
      RECT  190.9 236.0 192.5 236.8 ;
      RECT  193.3 235.2 194.1 246.0 ;
      RECT  191.7 235.2 192.5 236.0 ;
      RECT  189.9 246.0 190.7 245.2 ;
      RECT  186.5 256.0 187.3 245.2 ;
      RECT  191.7 254.4 192.5 245.2 ;
      RECT  188.1 256.0 188.9 245.2 ;
      RECT  190.9 255.2 192.5 254.4 ;
      RECT  193.3 256.0 194.1 245.2 ;
      RECT  191.7 256.0 192.5 255.2 ;
      RECT  189.9 266.0 190.7 266.8 ;
      RECT  186.5 256.0 187.3 266.8 ;
      RECT  191.7 257.6 192.5 266.8 ;
      RECT  188.1 256.0 188.9 266.8 ;
      RECT  190.9 256.8 192.5 257.6 ;
      RECT  193.3 256.0 194.1 266.8 ;
      RECT  191.7 256.0 192.5 256.8 ;
      RECT  189.9 266.8 190.7 266.0 ;
      RECT  186.5 276.8 187.3 266.0 ;
      RECT  191.7 275.2 192.5 266.0 ;
      RECT  188.1 276.8 188.9 266.0 ;
      RECT  190.9 276.0 192.5 275.2 ;
      RECT  193.3 276.8 194.1 266.0 ;
      RECT  191.7 276.8 192.5 276.0 ;
      RECT  189.9 286.8 190.7 287.6 ;
      RECT  186.5 276.8 187.3 287.6 ;
      RECT  191.7 278.4 192.5 287.6 ;
      RECT  188.1 276.8 188.9 287.6 ;
      RECT  190.9 277.6 192.5 278.4 ;
      RECT  193.3 276.8 194.1 287.6 ;
      RECT  191.7 276.8 192.5 277.6 ;
      RECT  189.9 287.6 190.7 286.8 ;
      RECT  186.5 297.6 187.3 286.8 ;
      RECT  191.7 296.0 192.5 286.8 ;
      RECT  188.1 297.6 188.9 286.8 ;
      RECT  190.9 296.8 192.5 296.0 ;
      RECT  193.3 297.6 194.1 286.8 ;
      RECT  191.7 297.6 192.5 296.8 ;
      RECT  189.9 307.6 190.7 308.4 ;
      RECT  186.5 297.6 187.3 308.4 ;
      RECT  191.7 299.2 192.5 308.4 ;
      RECT  188.1 297.6 188.9 308.4 ;
      RECT  190.9 298.4 192.5 299.2 ;
      RECT  193.3 297.6 194.1 308.4 ;
      RECT  191.7 297.6 192.5 298.4 ;
      RECT  189.9 308.4 190.7 307.6 ;
      RECT  186.5 318.4 187.3 307.6 ;
      RECT  191.7 316.8 192.5 307.6 ;
      RECT  188.1 318.4 188.9 307.6 ;
      RECT  190.9 317.6 192.5 316.8 ;
      RECT  193.3 318.4 194.1 307.6 ;
      RECT  191.7 318.4 192.5 317.6 ;
      RECT  189.9 328.4 190.7 329.2 ;
      RECT  186.5 318.4 187.3 329.2 ;
      RECT  191.7 320.0 192.5 329.2 ;
      RECT  188.1 318.4 188.9 329.2 ;
      RECT  190.9 319.2 192.5 320.0 ;
      RECT  193.3 318.4 194.1 329.2 ;
      RECT  191.7 318.4 192.5 319.2 ;
      RECT  189.9 329.2 190.7 328.4 ;
      RECT  186.5 339.2 187.3 328.4 ;
      RECT  191.7 337.6 192.5 328.4 ;
      RECT  188.1 339.2 188.9 328.4 ;
      RECT  190.9 338.4 192.5 337.6 ;
      RECT  193.3 339.2 194.1 328.4 ;
      RECT  191.7 339.2 192.5 338.4 ;
      RECT  189.9 349.2 190.7 350.0 ;
      RECT  186.5 339.2 187.3 350.0 ;
      RECT  191.7 340.8 192.5 350.0 ;
      RECT  188.1 339.2 188.9 350.0 ;
      RECT  190.9 340.0 192.5 340.8 ;
      RECT  193.3 339.2 194.1 350.0 ;
      RECT  191.7 339.2 192.5 340.0 ;
      RECT  189.9 350.0 190.7 349.2 ;
      RECT  186.5 360.0 187.3 349.2 ;
      RECT  191.7 358.4 192.5 349.2 ;
      RECT  188.1 360.0 188.9 349.2 ;
      RECT  190.9 359.2 192.5 358.4 ;
      RECT  193.3 360.0 194.1 349.2 ;
      RECT  191.7 360.0 192.5 359.2 ;
      RECT  196.7 203.6 197.5 204.4 ;
      RECT  193.3 193.6 194.1 204.4 ;
      RECT  198.5 195.2 199.3 204.4 ;
      RECT  194.9 193.6 195.7 204.4 ;
      RECT  197.7 194.4 199.3 195.2 ;
      RECT  200.1 193.6 200.9 204.4 ;
      RECT  198.5 193.6 199.3 194.4 ;
      RECT  196.7 204.4 197.5 203.6 ;
      RECT  193.3 214.4 194.1 203.6 ;
      RECT  198.5 212.8 199.3 203.6 ;
      RECT  194.9 214.4 195.7 203.6 ;
      RECT  197.7 213.6 199.3 212.8 ;
      RECT  200.1 214.4 200.9 203.6 ;
      RECT  198.5 214.4 199.3 213.6 ;
      RECT  196.7 224.4 197.5 225.2 ;
      RECT  193.3 214.4 194.1 225.2 ;
      RECT  198.5 216.0 199.3 225.2 ;
      RECT  194.9 214.4 195.7 225.2 ;
      RECT  197.7 215.2 199.3 216.0 ;
      RECT  200.1 214.4 200.9 225.2 ;
      RECT  198.5 214.4 199.3 215.2 ;
      RECT  196.7 225.2 197.5 224.4 ;
      RECT  193.3 235.2 194.1 224.4 ;
      RECT  198.5 233.6 199.3 224.4 ;
      RECT  194.9 235.2 195.7 224.4 ;
      RECT  197.7 234.4 199.3 233.6 ;
      RECT  200.1 235.2 200.9 224.4 ;
      RECT  198.5 235.2 199.3 234.4 ;
      RECT  196.7 245.2 197.5 246.0 ;
      RECT  193.3 235.2 194.1 246.0 ;
      RECT  198.5 236.8 199.3 246.0 ;
      RECT  194.9 235.2 195.7 246.0 ;
      RECT  197.7 236.0 199.3 236.8 ;
      RECT  200.1 235.2 200.9 246.0 ;
      RECT  198.5 235.2 199.3 236.0 ;
      RECT  196.7 246.0 197.5 245.2 ;
      RECT  193.3 256.0 194.1 245.2 ;
      RECT  198.5 254.4 199.3 245.2 ;
      RECT  194.9 256.0 195.7 245.2 ;
      RECT  197.7 255.2 199.3 254.4 ;
      RECT  200.1 256.0 200.9 245.2 ;
      RECT  198.5 256.0 199.3 255.2 ;
      RECT  196.7 266.0 197.5 266.8 ;
      RECT  193.3 256.0 194.1 266.8 ;
      RECT  198.5 257.6 199.3 266.8 ;
      RECT  194.9 256.0 195.7 266.8 ;
      RECT  197.7 256.8 199.3 257.6 ;
      RECT  200.1 256.0 200.9 266.8 ;
      RECT  198.5 256.0 199.3 256.8 ;
      RECT  196.7 266.8 197.5 266.0 ;
      RECT  193.3 276.8 194.1 266.0 ;
      RECT  198.5 275.2 199.3 266.0 ;
      RECT  194.9 276.8 195.7 266.0 ;
      RECT  197.7 276.0 199.3 275.2 ;
      RECT  200.1 276.8 200.9 266.0 ;
      RECT  198.5 276.8 199.3 276.0 ;
      RECT  196.7 286.8 197.5 287.6 ;
      RECT  193.3 276.8 194.1 287.6 ;
      RECT  198.5 278.4 199.3 287.6 ;
      RECT  194.9 276.8 195.7 287.6 ;
      RECT  197.7 277.6 199.3 278.4 ;
      RECT  200.1 276.8 200.9 287.6 ;
      RECT  198.5 276.8 199.3 277.6 ;
      RECT  196.7 287.6 197.5 286.8 ;
      RECT  193.3 297.6 194.1 286.8 ;
      RECT  198.5 296.0 199.3 286.8 ;
      RECT  194.9 297.6 195.7 286.8 ;
      RECT  197.7 296.8 199.3 296.0 ;
      RECT  200.1 297.6 200.9 286.8 ;
      RECT  198.5 297.6 199.3 296.8 ;
      RECT  196.7 307.6 197.5 308.4 ;
      RECT  193.3 297.6 194.1 308.4 ;
      RECT  198.5 299.2 199.3 308.4 ;
      RECT  194.9 297.6 195.7 308.4 ;
      RECT  197.7 298.4 199.3 299.2 ;
      RECT  200.1 297.6 200.9 308.4 ;
      RECT  198.5 297.6 199.3 298.4 ;
      RECT  196.7 308.4 197.5 307.6 ;
      RECT  193.3 318.4 194.1 307.6 ;
      RECT  198.5 316.8 199.3 307.6 ;
      RECT  194.9 318.4 195.7 307.6 ;
      RECT  197.7 317.6 199.3 316.8 ;
      RECT  200.1 318.4 200.9 307.6 ;
      RECT  198.5 318.4 199.3 317.6 ;
      RECT  196.7 328.4 197.5 329.2 ;
      RECT  193.3 318.4 194.1 329.2 ;
      RECT  198.5 320.0 199.3 329.2 ;
      RECT  194.9 318.4 195.7 329.2 ;
      RECT  197.7 319.2 199.3 320.0 ;
      RECT  200.1 318.4 200.9 329.2 ;
      RECT  198.5 318.4 199.3 319.2 ;
      RECT  196.7 329.2 197.5 328.4 ;
      RECT  193.3 339.2 194.1 328.4 ;
      RECT  198.5 337.6 199.3 328.4 ;
      RECT  194.9 339.2 195.7 328.4 ;
      RECT  197.7 338.4 199.3 337.6 ;
      RECT  200.1 339.2 200.9 328.4 ;
      RECT  198.5 339.2 199.3 338.4 ;
      RECT  196.7 349.2 197.5 350.0 ;
      RECT  193.3 339.2 194.1 350.0 ;
      RECT  198.5 340.8 199.3 350.0 ;
      RECT  194.9 339.2 195.7 350.0 ;
      RECT  197.7 340.0 199.3 340.8 ;
      RECT  200.1 339.2 200.9 350.0 ;
      RECT  198.5 339.2 199.3 340.0 ;
      RECT  196.7 350.0 197.5 349.2 ;
      RECT  193.3 360.0 194.1 349.2 ;
      RECT  198.5 358.4 199.3 349.2 ;
      RECT  194.9 360.0 195.7 349.2 ;
      RECT  197.7 359.2 199.3 358.4 ;
      RECT  200.1 360.0 200.9 349.2 ;
      RECT  198.5 360.0 199.3 359.2 ;
      RECT  188.1 193.6 188.9 360.0 ;
      RECT  191.7 193.6 192.5 360.0 ;
      RECT  194.9 193.6 195.7 360.0 ;
      RECT  198.5 193.6 199.3 360.0 ;
      RECT  183.1 182.8 183.9 183.6 ;
      RECT  179.7 172.8 180.5 183.6 ;
      RECT  181.3 172.8 182.1 183.6 ;
      RECT  184.9 172.8 185.7 183.6 ;
      RECT  186.5 172.8 187.3 183.6 ;
      RECT  183.1 183.6 183.9 182.8 ;
      RECT  179.7 193.6 180.5 182.8 ;
      RECT  184.9 192.0 185.7 182.8 ;
      RECT  181.3 193.6 182.1 182.8 ;
      RECT  184.1 192.8 185.7 192.0 ;
      RECT  186.5 193.6 187.3 182.8 ;
      RECT  184.9 193.6 185.7 192.8 ;
      RECT  183.1 203.6 183.9 204.4 ;
      RECT  179.7 193.6 180.5 204.4 ;
      RECT  184.9 195.2 185.7 204.4 ;
      RECT  181.3 193.6 182.1 204.4 ;
      RECT  184.1 194.4 185.7 195.2 ;
      RECT  186.5 193.6 187.3 204.4 ;
      RECT  184.9 193.6 185.7 194.4 ;
      RECT  183.1 204.4 183.9 203.6 ;
      RECT  179.7 214.4 180.5 203.6 ;
      RECT  184.9 212.8 185.7 203.6 ;
      RECT  181.3 214.4 182.1 203.6 ;
      RECT  184.1 213.6 185.7 212.8 ;
      RECT  186.5 214.4 187.3 203.6 ;
      RECT  184.9 214.4 185.7 213.6 ;
      RECT  183.1 224.4 183.9 225.2 ;
      RECT  179.7 214.4 180.5 225.2 ;
      RECT  184.9 216.0 185.7 225.2 ;
      RECT  181.3 214.4 182.1 225.2 ;
      RECT  184.1 215.2 185.7 216.0 ;
      RECT  186.5 214.4 187.3 225.2 ;
      RECT  184.9 214.4 185.7 215.2 ;
      RECT  183.1 225.2 183.9 224.4 ;
      RECT  179.7 235.2 180.5 224.4 ;
      RECT  184.9 233.6 185.7 224.4 ;
      RECT  181.3 235.2 182.1 224.4 ;
      RECT  184.1 234.4 185.7 233.6 ;
      RECT  186.5 235.2 187.3 224.4 ;
      RECT  184.9 235.2 185.7 234.4 ;
      RECT  183.1 245.2 183.9 246.0 ;
      RECT  179.7 235.2 180.5 246.0 ;
      RECT  184.9 236.8 185.7 246.0 ;
      RECT  181.3 235.2 182.1 246.0 ;
      RECT  184.1 236.0 185.7 236.8 ;
      RECT  186.5 235.2 187.3 246.0 ;
      RECT  184.9 235.2 185.7 236.0 ;
      RECT  183.1 246.0 183.9 245.2 ;
      RECT  179.7 256.0 180.5 245.2 ;
      RECT  184.9 254.4 185.7 245.2 ;
      RECT  181.3 256.0 182.1 245.2 ;
      RECT  184.1 255.2 185.7 254.4 ;
      RECT  186.5 256.0 187.3 245.2 ;
      RECT  184.9 256.0 185.7 255.2 ;
      RECT  183.1 266.0 183.9 266.8 ;
      RECT  179.7 256.0 180.5 266.8 ;
      RECT  184.9 257.6 185.7 266.8 ;
      RECT  181.3 256.0 182.1 266.8 ;
      RECT  184.1 256.8 185.7 257.6 ;
      RECT  186.5 256.0 187.3 266.8 ;
      RECT  184.9 256.0 185.7 256.8 ;
      RECT  183.1 266.8 183.9 266.0 ;
      RECT  179.7 276.8 180.5 266.0 ;
      RECT  184.9 275.2 185.7 266.0 ;
      RECT  181.3 276.8 182.1 266.0 ;
      RECT  184.1 276.0 185.7 275.2 ;
      RECT  186.5 276.8 187.3 266.0 ;
      RECT  184.9 276.8 185.7 276.0 ;
      RECT  183.1 286.8 183.9 287.6 ;
      RECT  179.7 276.8 180.5 287.6 ;
      RECT  184.9 278.4 185.7 287.6 ;
      RECT  181.3 276.8 182.1 287.6 ;
      RECT  184.1 277.6 185.7 278.4 ;
      RECT  186.5 276.8 187.3 287.6 ;
      RECT  184.9 276.8 185.7 277.6 ;
      RECT  183.1 287.6 183.9 286.8 ;
      RECT  179.7 297.6 180.5 286.8 ;
      RECT  184.9 296.0 185.7 286.8 ;
      RECT  181.3 297.6 182.1 286.8 ;
      RECT  184.1 296.8 185.7 296.0 ;
      RECT  186.5 297.6 187.3 286.8 ;
      RECT  184.9 297.6 185.7 296.8 ;
      RECT  183.1 307.6 183.9 308.4 ;
      RECT  179.7 297.6 180.5 308.4 ;
      RECT  184.9 299.2 185.7 308.4 ;
      RECT  181.3 297.6 182.1 308.4 ;
      RECT  184.1 298.4 185.7 299.2 ;
      RECT  186.5 297.6 187.3 308.4 ;
      RECT  184.9 297.6 185.7 298.4 ;
      RECT  183.1 308.4 183.9 307.6 ;
      RECT  179.7 318.4 180.5 307.6 ;
      RECT  184.9 316.8 185.7 307.6 ;
      RECT  181.3 318.4 182.1 307.6 ;
      RECT  184.1 317.6 185.7 316.8 ;
      RECT  186.5 318.4 187.3 307.6 ;
      RECT  184.9 318.4 185.7 317.6 ;
      RECT  183.1 328.4 183.9 329.2 ;
      RECT  179.7 318.4 180.5 329.2 ;
      RECT  184.9 320.0 185.7 329.2 ;
      RECT  181.3 318.4 182.1 329.2 ;
      RECT  184.1 319.2 185.7 320.0 ;
      RECT  186.5 318.4 187.3 329.2 ;
      RECT  184.9 318.4 185.7 319.2 ;
      RECT  183.1 329.2 183.9 328.4 ;
      RECT  179.7 339.2 180.5 328.4 ;
      RECT  184.9 337.6 185.7 328.4 ;
      RECT  181.3 339.2 182.1 328.4 ;
      RECT  184.1 338.4 185.7 337.6 ;
      RECT  186.5 339.2 187.3 328.4 ;
      RECT  184.9 339.2 185.7 338.4 ;
      RECT  183.1 349.2 183.9 350.0 ;
      RECT  179.7 339.2 180.5 350.0 ;
      RECT  184.9 340.8 185.7 350.0 ;
      RECT  181.3 339.2 182.1 350.0 ;
      RECT  184.1 340.0 185.7 340.8 ;
      RECT  186.5 339.2 187.3 350.0 ;
      RECT  184.9 339.2 185.7 340.0 ;
      RECT  183.1 350.0 183.9 349.2 ;
      RECT  179.7 360.0 180.5 349.2 ;
      RECT  184.9 358.4 185.7 349.2 ;
      RECT  181.3 360.0 182.1 349.2 ;
      RECT  184.1 359.2 185.7 358.4 ;
      RECT  186.5 360.0 187.3 349.2 ;
      RECT  184.9 360.0 185.7 359.2 ;
      RECT  183.1 370.0 183.9 370.8 ;
      RECT  179.7 360.0 180.5 370.8 ;
      RECT  181.3 360.0 182.1 370.8 ;
      RECT  184.9 360.0 185.7 370.8 ;
      RECT  186.5 360.0 187.3 370.8 ;
      RECT  183.1 349.2 183.9 350.0 ;
      RECT  183.1 224.4 183.9 225.2 ;
      RECT  183.1 224.4 183.9 225.2 ;
      RECT  183.1 370.0 183.9 370.8 ;
      RECT  183.1 203.6 183.9 204.4 ;
      RECT  183.1 266.0 183.9 266.8 ;
      RECT  183.1 245.2 183.9 246.0 ;
      RECT  183.1 307.6 183.9 308.4 ;
      RECT  183.1 286.8 183.9 287.6 ;
      RECT  183.1 286.8 183.9 287.6 ;
      RECT  183.1 307.6 183.9 308.4 ;
      RECT  183.1 328.4 183.9 329.2 ;
      RECT  183.1 182.8 183.9 183.6 ;
      RECT  186.5 224.4 187.3 235.2 ;
      RECT  179.7 328.4 180.5 339.2 ;
      RECT  186.5 328.4 187.3 339.2 ;
      RECT  186.5 349.2 187.3 360.0 ;
      RECT  186.5 256.0 187.3 266.8 ;
      RECT  186.5 266.0 187.3 276.8 ;
      RECT  186.5 339.2 187.3 350.0 ;
      RECT  186.5 360.0 187.3 370.8 ;
      RECT  179.7 235.2 180.5 246.0 ;
      RECT  179.7 256.0 180.5 266.8 ;
      RECT  179.7 318.4 180.5 329.2 ;
      RECT  179.7 193.6 180.5 204.4 ;
      RECT  179.7 182.8 180.5 193.6 ;
      RECT  179.7 266.0 180.5 276.8 ;
      RECT  179.7 203.6 180.5 214.4 ;
      RECT  179.7 349.2 180.5 360.0 ;
      RECT  186.5 245.2 187.3 256.0 ;
      RECT  179.7 214.4 180.5 225.2 ;
      RECT  186.5 286.8 187.3 297.6 ;
      RECT  186.5 203.6 187.3 214.4 ;
      RECT  186.5 214.4 187.3 225.2 ;
      RECT  186.5 182.8 187.3 193.6 ;
      RECT  179.7 172.8 180.5 183.6 ;
      RECT  179.7 339.2 180.5 350.0 ;
      RECT  179.7 286.8 180.5 297.6 ;
      RECT  179.7 276.8 180.5 287.6 ;
      RECT  186.5 193.6 187.3 204.4 ;
      RECT  186.5 307.6 187.3 318.4 ;
      RECT  179.7 224.4 180.5 235.2 ;
      RECT  186.5 235.2 187.3 246.0 ;
      RECT  186.5 297.6 187.3 308.4 ;
      RECT  186.5 276.8 187.3 287.6 ;
      RECT  179.7 360.0 180.5 370.8 ;
      RECT  179.7 245.2 180.5 256.0 ;
      RECT  186.5 318.4 187.3 329.2 ;
      RECT  179.7 297.6 180.5 308.4 ;
      RECT  186.5 172.8 187.3 183.6 ;
      RECT  179.7 307.6 180.5 318.4 ;
      RECT  189.9 183.6 190.7 182.8 ;
      RECT  186.5 193.6 187.3 182.8 ;
      RECT  188.1 193.6 188.9 182.8 ;
      RECT  191.7 193.6 192.5 182.8 ;
      RECT  193.3 193.6 194.1 182.8 ;
      RECT  196.7 183.6 197.5 182.8 ;
      RECT  193.3 193.6 194.1 182.8 ;
      RECT  194.9 193.6 195.7 182.8 ;
      RECT  198.5 193.6 199.3 182.8 ;
      RECT  200.1 193.6 200.9 182.8 ;
      RECT  188.1 193.6 188.9 183.2 ;
      RECT  191.7 193.6 192.5 183.2 ;
      RECT  194.9 193.6 195.7 183.2 ;
      RECT  198.5 193.6 199.3 183.2 ;
      RECT  189.9 182.8 190.7 183.6 ;
      RECT  186.5 172.8 187.3 183.6 ;
      RECT  188.1 172.8 188.9 183.6 ;
      RECT  191.7 172.8 192.5 183.6 ;
      RECT  193.3 172.8 194.1 183.6 ;
      RECT  196.7 182.8 197.5 183.6 ;
      RECT  193.3 172.8 194.1 183.6 ;
      RECT  194.9 172.8 195.7 183.6 ;
      RECT  198.5 172.8 199.3 183.6 ;
      RECT  200.1 172.8 200.9 183.6 ;
      RECT  188.1 172.8 188.9 183.2 ;
      RECT  191.7 172.8 192.5 183.2 ;
      RECT  194.9 172.8 195.7 183.2 ;
      RECT  198.5 172.8 199.3 183.2 ;
      RECT  189.9 370.0 190.7 370.8 ;
      RECT  186.5 360.0 187.3 370.8 ;
      RECT  188.1 360.0 188.9 370.8 ;
      RECT  191.7 360.0 192.5 370.8 ;
      RECT  193.3 360.0 194.1 370.8 ;
      RECT  196.7 370.0 197.5 370.8 ;
      RECT  193.3 360.0 194.1 370.8 ;
      RECT  194.9 360.0 195.7 370.8 ;
      RECT  198.5 360.0 199.3 370.8 ;
      RECT  200.1 360.0 200.9 370.8 ;
      RECT  188.1 360.0 188.9 370.4 ;
      RECT  191.7 360.0 192.5 370.4 ;
      RECT  194.9 360.0 195.7 370.4 ;
      RECT  198.5 360.0 199.3 370.4 ;
      RECT  176.3 182.8 177.1 183.6 ;
      RECT  172.9 172.8 173.7 183.6 ;
      RECT  174.5 172.8 175.3 183.6 ;
      RECT  178.1 172.8 178.9 183.6 ;
      RECT  179.7 172.8 180.5 183.6 ;
      RECT  176.3 183.6 177.1 182.8 ;
      RECT  172.9 193.6 173.7 182.8 ;
      RECT  174.5 193.6 175.3 182.8 ;
      RECT  178.1 193.6 178.9 182.8 ;
      RECT  179.7 193.6 180.5 182.8 ;
      RECT  176.3 203.6 177.1 204.4 ;
      RECT  172.9 193.6 173.7 204.4 ;
      RECT  174.5 193.6 175.3 204.4 ;
      RECT  178.1 193.6 178.9 204.4 ;
      RECT  179.7 193.6 180.5 204.4 ;
      RECT  176.3 204.4 177.1 203.6 ;
      RECT  172.9 214.4 173.7 203.6 ;
      RECT  174.5 214.4 175.3 203.6 ;
      RECT  178.1 214.4 178.9 203.6 ;
      RECT  179.7 214.4 180.5 203.6 ;
      RECT  176.3 224.4 177.1 225.2 ;
      RECT  172.9 214.4 173.7 225.2 ;
      RECT  174.5 214.4 175.3 225.2 ;
      RECT  178.1 214.4 178.9 225.2 ;
      RECT  179.7 214.4 180.5 225.2 ;
      RECT  176.3 225.2 177.1 224.4 ;
      RECT  172.9 235.2 173.7 224.4 ;
      RECT  174.5 235.2 175.3 224.4 ;
      RECT  178.1 235.2 178.9 224.4 ;
      RECT  179.7 235.2 180.5 224.4 ;
      RECT  176.3 245.2 177.1 246.0 ;
      RECT  172.9 235.2 173.7 246.0 ;
      RECT  174.5 235.2 175.3 246.0 ;
      RECT  178.1 235.2 178.9 246.0 ;
      RECT  179.7 235.2 180.5 246.0 ;
      RECT  176.3 246.0 177.1 245.2 ;
      RECT  172.9 256.0 173.7 245.2 ;
      RECT  174.5 256.0 175.3 245.2 ;
      RECT  178.1 256.0 178.9 245.2 ;
      RECT  179.7 256.0 180.5 245.2 ;
      RECT  176.3 266.0 177.1 266.8 ;
      RECT  172.9 256.0 173.7 266.8 ;
      RECT  174.5 256.0 175.3 266.8 ;
      RECT  178.1 256.0 178.9 266.8 ;
      RECT  179.7 256.0 180.5 266.8 ;
      RECT  176.3 266.8 177.1 266.0 ;
      RECT  172.9 276.8 173.7 266.0 ;
      RECT  174.5 276.8 175.3 266.0 ;
      RECT  178.1 276.8 178.9 266.0 ;
      RECT  179.7 276.8 180.5 266.0 ;
      RECT  176.3 286.8 177.1 287.6 ;
      RECT  172.9 276.8 173.7 287.6 ;
      RECT  174.5 276.8 175.3 287.6 ;
      RECT  178.1 276.8 178.9 287.6 ;
      RECT  179.7 276.8 180.5 287.6 ;
      RECT  176.3 287.6 177.1 286.8 ;
      RECT  172.9 297.6 173.7 286.8 ;
      RECT  174.5 297.6 175.3 286.8 ;
      RECT  178.1 297.6 178.9 286.8 ;
      RECT  179.7 297.6 180.5 286.8 ;
      RECT  176.3 307.6 177.1 308.4 ;
      RECT  172.9 297.6 173.7 308.4 ;
      RECT  174.5 297.6 175.3 308.4 ;
      RECT  178.1 297.6 178.9 308.4 ;
      RECT  179.7 297.6 180.5 308.4 ;
      RECT  176.3 308.4 177.1 307.6 ;
      RECT  172.9 318.4 173.7 307.6 ;
      RECT  174.5 318.4 175.3 307.6 ;
      RECT  178.1 318.4 178.9 307.6 ;
      RECT  179.7 318.4 180.5 307.6 ;
      RECT  176.3 328.4 177.1 329.2 ;
      RECT  172.9 318.4 173.7 329.2 ;
      RECT  174.5 318.4 175.3 329.2 ;
      RECT  178.1 318.4 178.9 329.2 ;
      RECT  179.7 318.4 180.5 329.2 ;
      RECT  176.3 329.2 177.1 328.4 ;
      RECT  172.9 339.2 173.7 328.4 ;
      RECT  174.5 339.2 175.3 328.4 ;
      RECT  178.1 339.2 178.9 328.4 ;
      RECT  179.7 339.2 180.5 328.4 ;
      RECT  176.3 349.2 177.1 350.0 ;
      RECT  172.9 339.2 173.7 350.0 ;
      RECT  174.5 339.2 175.3 350.0 ;
      RECT  178.1 339.2 178.9 350.0 ;
      RECT  179.7 339.2 180.5 350.0 ;
      RECT  176.3 350.0 177.1 349.2 ;
      RECT  172.9 360.0 173.7 349.2 ;
      RECT  174.5 360.0 175.3 349.2 ;
      RECT  178.1 360.0 178.9 349.2 ;
      RECT  179.7 360.0 180.5 349.2 ;
      RECT  176.3 370.0 177.1 370.8 ;
      RECT  172.9 360.0 173.7 370.8 ;
      RECT  174.5 360.0 175.3 370.8 ;
      RECT  178.1 360.0 178.9 370.8 ;
      RECT  179.7 360.0 180.5 370.8 ;
      RECT  174.5 172.8 175.3 370.4 ;
      RECT  178.1 172.8 178.9 370.4 ;
      RECT  203.5 182.8 204.3 183.6 ;
      RECT  200.1 172.8 200.9 183.6 ;
      RECT  201.7 172.8 202.5 183.6 ;
      RECT  205.3 172.8 206.1 183.6 ;
      RECT  206.9 172.8 207.7 183.6 ;
      RECT  203.5 183.6 204.3 182.8 ;
      RECT  200.1 193.6 200.9 182.8 ;
      RECT  201.7 193.6 202.5 182.8 ;
      RECT  205.3 193.6 206.1 182.8 ;
      RECT  206.9 193.6 207.7 182.8 ;
      RECT  203.5 203.6 204.3 204.4 ;
      RECT  200.1 193.6 200.9 204.4 ;
      RECT  201.7 193.6 202.5 204.4 ;
      RECT  205.3 193.6 206.1 204.4 ;
      RECT  206.9 193.6 207.7 204.4 ;
      RECT  203.5 204.4 204.3 203.6 ;
      RECT  200.1 214.4 200.9 203.6 ;
      RECT  201.7 214.4 202.5 203.6 ;
      RECT  205.3 214.4 206.1 203.6 ;
      RECT  206.9 214.4 207.7 203.6 ;
      RECT  203.5 224.4 204.3 225.2 ;
      RECT  200.1 214.4 200.9 225.2 ;
      RECT  201.7 214.4 202.5 225.2 ;
      RECT  205.3 214.4 206.1 225.2 ;
      RECT  206.9 214.4 207.7 225.2 ;
      RECT  203.5 225.2 204.3 224.4 ;
      RECT  200.1 235.2 200.9 224.4 ;
      RECT  201.7 235.2 202.5 224.4 ;
      RECT  205.3 235.2 206.1 224.4 ;
      RECT  206.9 235.2 207.7 224.4 ;
      RECT  203.5 245.2 204.3 246.0 ;
      RECT  200.1 235.2 200.9 246.0 ;
      RECT  201.7 235.2 202.5 246.0 ;
      RECT  205.3 235.2 206.1 246.0 ;
      RECT  206.9 235.2 207.7 246.0 ;
      RECT  203.5 246.0 204.3 245.2 ;
      RECT  200.1 256.0 200.9 245.2 ;
      RECT  201.7 256.0 202.5 245.2 ;
      RECT  205.3 256.0 206.1 245.2 ;
      RECT  206.9 256.0 207.7 245.2 ;
      RECT  203.5 266.0 204.3 266.8 ;
      RECT  200.1 256.0 200.9 266.8 ;
      RECT  201.7 256.0 202.5 266.8 ;
      RECT  205.3 256.0 206.1 266.8 ;
      RECT  206.9 256.0 207.7 266.8 ;
      RECT  203.5 266.8 204.3 266.0 ;
      RECT  200.1 276.8 200.9 266.0 ;
      RECT  201.7 276.8 202.5 266.0 ;
      RECT  205.3 276.8 206.1 266.0 ;
      RECT  206.9 276.8 207.7 266.0 ;
      RECT  203.5 286.8 204.3 287.6 ;
      RECT  200.1 276.8 200.9 287.6 ;
      RECT  201.7 276.8 202.5 287.6 ;
      RECT  205.3 276.8 206.1 287.6 ;
      RECT  206.9 276.8 207.7 287.6 ;
      RECT  203.5 287.6 204.3 286.8 ;
      RECT  200.1 297.6 200.9 286.8 ;
      RECT  201.7 297.6 202.5 286.8 ;
      RECT  205.3 297.6 206.1 286.8 ;
      RECT  206.9 297.6 207.7 286.8 ;
      RECT  203.5 307.6 204.3 308.4 ;
      RECT  200.1 297.6 200.9 308.4 ;
      RECT  201.7 297.6 202.5 308.4 ;
      RECT  205.3 297.6 206.1 308.4 ;
      RECT  206.9 297.6 207.7 308.4 ;
      RECT  203.5 308.4 204.3 307.6 ;
      RECT  200.1 318.4 200.9 307.6 ;
      RECT  201.7 318.4 202.5 307.6 ;
      RECT  205.3 318.4 206.1 307.6 ;
      RECT  206.9 318.4 207.7 307.6 ;
      RECT  203.5 328.4 204.3 329.2 ;
      RECT  200.1 318.4 200.9 329.2 ;
      RECT  201.7 318.4 202.5 329.2 ;
      RECT  205.3 318.4 206.1 329.2 ;
      RECT  206.9 318.4 207.7 329.2 ;
      RECT  203.5 329.2 204.3 328.4 ;
      RECT  200.1 339.2 200.9 328.4 ;
      RECT  201.7 339.2 202.5 328.4 ;
      RECT  205.3 339.2 206.1 328.4 ;
      RECT  206.9 339.2 207.7 328.4 ;
      RECT  203.5 349.2 204.3 350.0 ;
      RECT  200.1 339.2 200.9 350.0 ;
      RECT  201.7 339.2 202.5 350.0 ;
      RECT  205.3 339.2 206.1 350.0 ;
      RECT  206.9 339.2 207.7 350.0 ;
      RECT  203.5 350.0 204.3 349.2 ;
      RECT  200.1 360.0 200.9 349.2 ;
      RECT  201.7 360.0 202.5 349.2 ;
      RECT  205.3 360.0 206.1 349.2 ;
      RECT  206.9 360.0 207.7 349.2 ;
      RECT  203.5 370.0 204.3 370.8 ;
      RECT  200.1 360.0 200.9 370.8 ;
      RECT  201.7 360.0 202.5 370.8 ;
      RECT  205.3 360.0 206.1 370.8 ;
      RECT  206.9 360.0 207.7 370.8 ;
      RECT  201.7 172.8 202.5 370.4 ;
      RECT  205.3 172.8 206.1 370.4 ;
      RECT  188.1 172.8 188.9 370.4 ;
      RECT  191.7 172.8 192.5 370.4 ;
      RECT  194.9 172.8 195.7 370.4 ;
      RECT  198.5 172.8 199.3 370.4 ;
      RECT  181.3 172.8 182.1 370.4 ;
      RECT  184.9 172.8 185.7 370.4 ;
      RECT  181.2 156.6 181.8 168.6 ;
      RECT  185.2 156.6 185.8 168.6 ;
      RECT  188.0 156.6 188.6 168.6 ;
      RECT  192.0 156.6 192.6 168.6 ;
      RECT  194.8 156.6 195.4 168.6 ;
      RECT  198.8 156.6 199.4 168.6 ;
      RECT  181.2 156.6 181.8 168.6 ;
      RECT  185.2 156.6 185.8 168.6 ;
      RECT  188.0 156.6 188.6 168.6 ;
      RECT  192.0 156.6 192.6 168.6 ;
      RECT  194.8 156.6 195.4 168.6 ;
      RECT  198.8 156.6 199.4 168.6 ;
      RECT  188.9 129.4 189.7 152.4 ;
      RECT  190.9 129.4 191.7 152.4 ;
      RECT  190.9 119.8 191.7 128.6 ;
      RECT  187.5 119.8 188.3 122.8 ;
      RECT  193.3 145.6 194.1 147.2 ;
      RECT  190.9 128.6 192.1 129.4 ;
      RECT  188.9 119.8 189.7 128.6 ;
      RECT  192.3 132.2 193.1 133.8 ;
      RECT  188.9 128.6 190.3 129.4 ;
      RECT  195.7 129.4 196.5 152.4 ;
      RECT  197.7 129.4 198.5 152.4 ;
      RECT  197.7 119.8 198.5 128.6 ;
      RECT  194.3 119.8 195.1 122.8 ;
      RECT  200.1 145.6 200.9 147.2 ;
      RECT  197.7 128.6 198.9 129.4 ;
      RECT  195.7 119.8 196.5 128.6 ;
      RECT  199.1 132.2 199.9 133.8 ;
      RECT  195.7 128.6 197.1 129.4 ;
      RECT  187.5 119.8 188.3 122.8 ;
      RECT  188.9 129.4 189.7 152.4 ;
      RECT  190.9 129.4 191.7 152.4 ;
      RECT  194.3 119.8 195.1 122.8 ;
      RECT  195.7 129.4 196.5 152.4 ;
      RECT  197.7 129.4 198.5 152.4 ;
      RECT  190.9 110.6 191.7 115.6 ;
      RECT  192.1 92.2 192.9 93.0 ;
      RECT  190.7 87.8 191.5 88.6 ;
      RECT  188.9 113.6 189.7 115.6 ;
      RECT  189.3 106.8 190.1 107.6 ;
      RECT  190.1 98.6 190.9 99.4 ;
      RECT  189.9 75.0 190.7 77.0 ;
      RECT  190.7 81.2 191.5 82.0 ;
      RECT  197.7 110.6 198.5 115.6 ;
      RECT  198.9 92.2 199.7 93.0 ;
      RECT  197.5 87.8 198.3 88.6 ;
      RECT  195.7 113.6 196.5 115.6 ;
      RECT  196.1 106.8 196.9 107.6 ;
      RECT  196.9 98.6 197.7 99.4 ;
      RECT  196.7 75.0 197.5 77.0 ;
      RECT  197.5 81.2 198.3 82.0 ;
      RECT  189.9 75.0 190.7 77.0 ;
      RECT  196.7 75.0 197.5 77.0 ;
      RECT  188.9 113.6 189.7 115.6 ;
      RECT  190.9 110.6 191.7 115.6 ;
      RECT  195.7 113.6 196.5 115.6 ;
      RECT  197.7 110.6 198.5 115.6 ;
      RECT  181.2 168.6 181.8 156.6 ;
      RECT  185.2 168.6 185.8 156.6 ;
      RECT  188.0 168.6 188.6 156.6 ;
      RECT  192.0 168.6 192.6 156.6 ;
      RECT  194.8 168.6 195.4 156.6 ;
      RECT  198.8 168.6 199.4 156.6 ;
      RECT  187.5 122.8 188.3 119.8 ;
      RECT  194.3 122.8 195.1 119.8 ;
      RECT  189.9 77.0 190.7 75.0 ;
      RECT  196.7 77.0 197.5 75.0 ;
      RECT  89.8 198.6 90.6 199.4 ;
      RECT  91.2 209.4 92.0 210.2 ;
      RECT  89.8 250.6 90.6 251.4 ;
      RECT  91.2 261.4 92.0 262.2 ;
      RECT  82.3 194.0 82.9 287.6 ;
      RECT  83.7 194.0 84.3 287.6 ;
      RECT  85.1 194.0 85.7 287.6 ;
      RECT  86.5 194.0 87.1 287.6 ;
      RECT  156.9 194.0 157.5 360.4 ;
      RECT  82.3 194.0 82.9 287.6 ;
      RECT  83.7 194.0 84.3 287.6 ;
      RECT  85.1 194.0 85.7 287.6 ;
      RECT  86.5 194.0 87.1 287.6 ;
      RECT  156.9 194.0 157.5 360.4 ;
      RECT  187.5 119.8 188.3 122.8 ;
      RECT  194.3 119.8 195.1 122.8 ;
      RECT  189.9 75.0 190.7 77.0 ;
      RECT  196.7 75.0 197.5 77.0 ;
      RECT  82.3 194.0 82.9 287.6 ;
      RECT  83.7 194.0 84.3 287.6 ;
      RECT  85.1 194.0 85.7 287.6 ;
      RECT  86.5 194.0 87.1 287.6 ;
      RECT  167.7 75.0 168.3 190.8 ;
      RECT  169.1 75.0 169.7 190.8 ;
      RECT  166.3 75.0 166.9 190.8 ;
      RECT  170.5 75.0 171.1 190.8 ;
      RECT  10.0 10.2 10.8 11.0 ;
      RECT  21.2 11.0 22.0 11.8 ;
      RECT  5.2 8.2 6.0 9.0 ;
      RECT  3.6 6.8 4.4 12.4 ;
      RECT  6.8 4.8 7.6 16.4 ;
      RECT  16.4 4.8 17.2 16.4 ;
      RECT  10.0 10.2 10.8 11.0 ;
      RECT  38.2 7.7 38.8 8.3 ;
      RECT  32.6 13.7 33.2 14.3 ;
      RECT  5.2 8.2 6.0 9.0 ;
      RECT  10.0 33.0 10.8 32.2 ;
      RECT  21.2 32.2 22.0 31.4 ;
      RECT  5.2 35.0 6.0 34.2 ;
      RECT  3.6 36.4 4.4 30.8 ;
      RECT  6.8 38.4 7.6 26.8 ;
      RECT  16.4 38.4 17.2 26.8 ;
      RECT  10.0 33.0 10.8 32.2 ;
      RECT  38.2 35.5 38.8 34.9 ;
      RECT  32.6 29.5 33.2 28.9 ;
      RECT  5.2 35.0 6.0 34.2 ;
      RECT  10.0 10.2 10.8 11.0 ;
      RECT  10.0 32.2 10.8 33.0 ;
      RECT  38.2 7.7 38.8 8.3 ;
      RECT  32.6 13.7 33.2 14.3 ;
      RECT  38.2 34.9 38.8 35.5 ;
      RECT  32.6 28.9 33.2 29.5 ;
      RECT  5.2 1.6 5.8 41.6 ;
      RECT  33.8 164.4 33.2 174.0 ;
      RECT  5.5 164.4 4.9 330.8 ;
      RECT  10.0 10.2 10.8 11.0 ;
      RECT  10.0 32.2 10.8 33.0 ;
      RECT  54.1 1.6 54.7 11.4 ;
      RECT  33.2 164.4 33.8 174.0 ;
      RECT  65.2 352.2 66.0 353.0 ;
      RECT  76.4 353.0 77.2 353.8 ;
      RECT  60.4 350.2 61.2 351.0 ;
      RECT  58.8 348.8 59.6 354.4 ;
      RECT  62.0 346.8 62.8 358.4 ;
      RECT  71.6 346.8 72.4 358.4 ;
      RECT  65.2 375.0 66.0 374.2 ;
      RECT  76.4 374.2 77.2 373.4 ;
      RECT  60.4 377.0 61.2 376.2 ;
      RECT  58.8 378.4 59.6 372.8 ;
      RECT  62.0 380.4 62.8 368.8 ;
      RECT  71.6 380.4 72.4 368.8 ;
      RECT  65.2 392.2 66.0 393.0 ;
      RECT  76.4 393.0 77.2 393.8 ;
      RECT  60.4 390.2 61.2 391.0 ;
      RECT  58.8 388.8 59.6 394.4 ;
      RECT  62.0 386.8 62.8 398.4 ;
      RECT  71.6 386.8 72.4 398.4 ;
      RECT  65.2 415.0 66.0 414.2 ;
      RECT  76.4 414.2 77.2 413.4 ;
      RECT  60.4 417.0 61.2 416.2 ;
      RECT  58.8 418.4 59.6 412.8 ;
      RECT  62.0 420.4 62.8 408.8 ;
      RECT  71.6 420.4 72.4 408.8 ;
      RECT  65.2 352.2 66.0 353.0 ;
      RECT  65.2 374.2 66.0 375.0 ;
      RECT  65.2 392.2 66.0 393.0 ;
      RECT  65.2 414.2 66.0 415.0 ;
      RECT  76.4 353.0 77.2 353.8 ;
      RECT  76.4 373.4 77.2 374.2 ;
      RECT  76.4 393.0 77.2 393.8 ;
      RECT  76.4 413.4 77.2 414.2 ;
      RECT  180.9 56.6 181.7 57.4 ;
      RECT  192.1 57.4 192.9 58.2 ;
      RECT  176.1 54.6 176.9 55.4 ;
      RECT  174.5 53.2 175.3 58.8 ;
      RECT  177.7 51.2 178.5 62.8 ;
      RECT  187.3 51.2 188.1 62.8 ;
      RECT  202.7 56.6 203.5 57.4 ;
      RECT  213.9 57.4 214.7 58.2 ;
      RECT  197.9 54.6 198.7 55.4 ;
      RECT  196.3 53.2 197.1 58.8 ;
      RECT  199.5 51.2 200.3 62.8 ;
      RECT  209.1 51.2 209.9 62.8 ;
      RECT  180.9 56.6 181.7 57.4 ;
      RECT  202.7 56.6 203.5 57.4 ;
      RECT  192.1 57.4 192.9 58.2 ;
      RECT  213.9 57.4 214.7 58.2 ;
   LAYER  m3 ;
      RECT  189.9 286.8 190.7 287.6 ;
      RECT  196.7 307.6 197.5 308.4 ;
      RECT  189.9 203.6 190.7 204.4 ;
      RECT  189.9 307.6 190.7 308.4 ;
      RECT  196.7 224.4 197.5 225.2 ;
      RECT  196.7 286.8 197.5 287.6 ;
      RECT  189.9 349.2 190.7 350.0 ;
      RECT  196.7 245.2 197.5 246.0 ;
      RECT  196.7 245.2 197.5 246.0 ;
      RECT  196.7 349.2 197.5 350.0 ;
      RECT  189.9 266.0 190.7 266.8 ;
      RECT  189.9 245.2 190.7 246.0 ;
      RECT  189.9 245.2 190.7 246.0 ;
      RECT  189.9 224.4 190.7 225.2 ;
      RECT  189.9 328.4 190.7 329.2 ;
      RECT  189.9 328.4 190.7 329.2 ;
      RECT  196.7 203.6 197.5 204.4 ;
      RECT  196.7 266.0 197.5 266.8 ;
      RECT  196.7 328.4 197.5 329.2 ;
      RECT  196.7 328.4 197.5 329.2 ;
      RECT  193.3 323.4 194.1 324.2 ;
      RECT  186.5 281.8 187.3 282.6 ;
      RECT  200.1 219.4 200.9 220.2 ;
      RECT  186.5 208.6 187.3 209.4 ;
      RECT  186.5 219.4 187.3 220.2 ;
      RECT  200.1 333.4 200.9 334.2 ;
      RECT  200.1 312.6 200.9 313.4 ;
      RECT  186.5 312.6 187.3 313.4 ;
      RECT  193.3 354.2 194.1 355.0 ;
      RECT  193.3 229.4 194.1 230.2 ;
      RECT  193.3 291.8 194.1 292.6 ;
      RECT  200.1 302.6 200.9 303.4 ;
      RECT  200.1 344.2 200.9 345.0 ;
      RECT  200.1 354.2 200.9 355.0 ;
      RECT  200.1 229.4 200.9 230.2 ;
      RECT  200.1 261.0 200.9 261.8 ;
      RECT  186.5 229.4 187.3 230.2 ;
      RECT  200.1 250.2 200.9 251.0 ;
      RECT  186.5 302.6 187.3 303.4 ;
      RECT  186.5 333.4 187.3 334.2 ;
      RECT  193.3 333.4 194.1 334.2 ;
      RECT  186.5 344.2 187.3 345.0 ;
      RECT  193.3 344.2 194.1 345.0 ;
      RECT  193.3 219.4 194.1 220.2 ;
      RECT  200.1 281.8 200.9 282.6 ;
      RECT  186.5 198.6 187.3 199.4 ;
      RECT  200.1 271.0 200.9 271.8 ;
      RECT  193.3 208.6 194.1 209.4 ;
      RECT  193.3 250.2 194.1 251.0 ;
      RECT  186.5 250.2 187.3 251.0 ;
      RECT  193.3 261.0 194.1 261.8 ;
      RECT  186.5 354.2 187.3 355.0 ;
      RECT  186.5 240.2 187.3 241.0 ;
      RECT  193.3 302.6 194.1 303.4 ;
      RECT  200.1 208.6 200.9 209.4 ;
      RECT  186.5 323.4 187.3 324.2 ;
      RECT  186.5 261.0 187.3 261.8 ;
      RECT  193.3 240.2 194.1 241.0 ;
      RECT  193.3 281.8 194.1 282.6 ;
      RECT  186.5 271.0 187.3 271.8 ;
      RECT  200.1 291.8 200.9 292.6 ;
      RECT  200.1 240.2 200.9 241.0 ;
      RECT  200.1 323.4 200.9 324.2 ;
      RECT  193.3 271.0 194.1 271.8 ;
      RECT  200.1 198.6 200.9 199.4 ;
      RECT  186.5 291.8 187.3 292.6 ;
      RECT  193.3 312.6 194.1 313.4 ;
      RECT  193.3 198.6 194.1 199.4 ;
      RECT  196.7 183.6 197.5 182.8 ;
      RECT  189.9 183.6 190.7 182.8 ;
      RECT  186.5 188.6 187.3 187.8 ;
      RECT  193.3 188.6 194.1 187.8 ;
      RECT  200.1 188.6 200.9 187.8 ;
      RECT  196.7 182.8 197.5 183.6 ;
      RECT  189.9 182.8 190.7 183.6 ;
      RECT  186.5 177.8 187.3 178.6 ;
      RECT  193.3 177.8 194.1 178.6 ;
      RECT  200.1 177.8 200.9 178.6 ;
      RECT  196.7 370.0 197.5 370.8 ;
      RECT  189.9 370.0 190.7 370.8 ;
      RECT  186.5 365.0 187.3 365.8 ;
      RECT  193.3 365.0 194.1 365.8 ;
      RECT  200.1 365.0 200.9 365.8 ;
      RECT  176.3 266.0 177.1 266.8 ;
      RECT  176.3 245.2 177.1 246.0 ;
      RECT  176.3 307.6 177.1 308.4 ;
      RECT  176.3 307.6 177.1 308.4 ;
      RECT  176.3 224.4 177.1 225.2 ;
      RECT  176.3 224.4 177.1 225.2 ;
      RECT  176.3 370.0 177.1 370.8 ;
      RECT  176.3 328.4 177.1 329.2 ;
      RECT  176.3 349.2 177.1 350.0 ;
      RECT  176.3 203.6 177.1 204.4 ;
      RECT  176.3 182.8 177.1 183.6 ;
      RECT  176.3 286.8 177.1 287.6 ;
      RECT  179.7 302.6 180.5 303.4 ;
      RECT  172.9 261.0 173.7 261.8 ;
      RECT  179.7 344.2 180.5 345.0 ;
      RECT  172.9 187.8 173.7 188.6 ;
      RECT  172.9 198.6 173.7 199.4 ;
      RECT  172.9 354.2 173.7 355.0 ;
      RECT  179.7 354.2 180.5 355.0 ;
      RECT  172.9 291.8 173.7 292.6 ;
      RECT  179.7 333.4 180.5 334.2 ;
      RECT  179.7 208.6 180.5 209.4 ;
      RECT  179.7 271.0 180.5 271.8 ;
      RECT  172.9 344.2 173.7 345.0 ;
      RECT  172.9 365.0 173.7 365.8 ;
      RECT  172.9 323.4 173.7 324.2 ;
      RECT  172.9 208.6 173.7 209.4 ;
      RECT  179.7 312.6 180.5 313.4 ;
      RECT  172.9 281.8 173.7 282.6 ;
      RECT  172.9 312.6 173.7 313.4 ;
      RECT  179.7 323.4 180.5 324.2 ;
      RECT  179.7 198.6 180.5 199.4 ;
      RECT  172.9 177.8 173.7 178.6 ;
      RECT  179.7 187.8 180.5 188.6 ;
      RECT  179.7 229.4 180.5 230.2 ;
      RECT  172.9 229.4 173.7 230.2 ;
      RECT  179.7 240.2 180.5 241.0 ;
      RECT  172.9 333.4 173.7 334.2 ;
      RECT  172.9 219.4 173.7 220.2 ;
      RECT  179.7 281.8 180.5 282.6 ;
      RECT  179.7 365.0 180.5 365.8 ;
      RECT  172.9 302.6 173.7 303.4 ;
      RECT  172.9 240.2 173.7 241.0 ;
      RECT  179.7 219.4 180.5 220.2 ;
      RECT  179.7 261.0 180.5 261.8 ;
      RECT  172.9 250.2 173.7 251.0 ;
      RECT  179.7 250.2 180.5 251.0 ;
      RECT  172.9 271.0 173.7 271.8 ;
      RECT  179.7 291.8 180.5 292.6 ;
      RECT  179.7 177.8 180.5 178.6 ;
      RECT  203.5 266.0 204.3 266.8 ;
      RECT  203.5 245.2 204.3 246.0 ;
      RECT  203.5 307.6 204.3 308.4 ;
      RECT  203.5 307.6 204.3 308.4 ;
      RECT  203.5 224.4 204.3 225.2 ;
      RECT  203.5 224.4 204.3 225.2 ;
      RECT  203.5 370.0 204.3 370.8 ;
      RECT  203.5 328.4 204.3 329.2 ;
      RECT  203.5 349.2 204.3 350.0 ;
      RECT  203.5 203.6 204.3 204.4 ;
      RECT  203.5 182.8 204.3 183.6 ;
      RECT  203.5 286.8 204.3 287.6 ;
      RECT  206.9 302.6 207.7 303.4 ;
      RECT  200.1 261.0 200.9 261.8 ;
      RECT  206.9 344.2 207.7 345.0 ;
      RECT  200.1 187.8 200.9 188.6 ;
      RECT  200.1 198.6 200.9 199.4 ;
      RECT  200.1 354.2 200.9 355.0 ;
      RECT  206.9 354.2 207.7 355.0 ;
      RECT  200.1 291.8 200.9 292.6 ;
      RECT  206.9 333.4 207.7 334.2 ;
      RECT  206.9 208.6 207.7 209.4 ;
      RECT  206.9 271.0 207.7 271.8 ;
      RECT  200.1 344.2 200.9 345.0 ;
      RECT  200.1 365.0 200.9 365.8 ;
      RECT  200.1 323.4 200.9 324.2 ;
      RECT  200.1 208.6 200.9 209.4 ;
      RECT  206.9 312.6 207.7 313.4 ;
      RECT  200.1 281.8 200.9 282.6 ;
      RECT  200.1 312.6 200.9 313.4 ;
      RECT  206.9 323.4 207.7 324.2 ;
      RECT  206.9 198.6 207.7 199.4 ;
      RECT  200.1 177.8 200.9 178.6 ;
      RECT  206.9 187.8 207.7 188.6 ;
      RECT  206.9 229.4 207.7 230.2 ;
      RECT  200.1 229.4 200.9 230.2 ;
      RECT  206.9 240.2 207.7 241.0 ;
      RECT  200.1 333.4 200.9 334.2 ;
      RECT  200.1 219.4 200.9 220.2 ;
      RECT  206.9 281.8 207.7 282.6 ;
      RECT  206.9 365.0 207.7 365.8 ;
      RECT  200.1 302.6 200.9 303.4 ;
      RECT  200.1 240.2 200.9 241.0 ;
      RECT  206.9 219.4 207.7 220.2 ;
      RECT  206.9 261.0 207.7 261.8 ;
      RECT  200.1 250.2 200.9 251.0 ;
      RECT  206.9 250.2 207.7 251.0 ;
      RECT  200.1 271.0 200.9 271.8 ;
      RECT  206.9 291.8 207.7 292.6 ;
      RECT  206.9 177.8 207.7 178.6 ;
      RECT  190.0 182.9 190.6 183.5 ;
      RECT  190.0 286.9 190.6 287.5 ;
      RECT  176.4 370.1 177.0 370.7 ;
      RECT  183.1 286.8 183.9 287.6 ;
      RECT  203.6 286.9 204.2 287.5 ;
      RECT  196.8 182.9 197.4 183.5 ;
      RECT  196.8 286.9 197.4 287.5 ;
      RECT  176.4 182.9 177.0 183.5 ;
      RECT  203.6 370.1 204.2 370.7 ;
      RECT  183.1 370.0 183.9 370.8 ;
      RECT  176.4 203.7 177.0 204.3 ;
      RECT  203.6 307.7 204.2 308.3 ;
      RECT  203.6 224.5 204.2 225.1 ;
      RECT  203.6 328.5 204.2 329.1 ;
      RECT  190.0 203.7 190.6 204.3 ;
      RECT  183.1 203.6 183.9 204.4 ;
      RECT  183.1 266.0 183.9 266.8 ;
      RECT  183.1 328.4 183.9 329.2 ;
      RECT  183.1 224.4 183.9 225.2 ;
      RECT  190.0 328.5 190.6 329.1 ;
      RECT  196.8 266.1 197.4 266.7 ;
      RECT  190.0 266.1 190.6 266.7 ;
      RECT  203.6 182.9 204.2 183.5 ;
      RECT  190.0 224.5 190.6 225.1 ;
      RECT  190.0 245.3 190.6 245.9 ;
      RECT  190.0 370.1 190.6 370.7 ;
      RECT  183.1 349.2 183.9 350.0 ;
      RECT  176.4 245.3 177.0 245.9 ;
      RECT  196.8 307.7 197.4 308.3 ;
      RECT  176.4 349.3 177.0 349.9 ;
      RECT  176.4 224.5 177.0 225.1 ;
      RECT  190.0 307.7 190.6 308.3 ;
      RECT  196.8 349.3 197.4 349.9 ;
      RECT  196.8 224.5 197.4 225.1 ;
      RECT  196.8 370.1 197.4 370.7 ;
      RECT  176.4 307.7 177.0 308.3 ;
      RECT  203.6 349.3 204.2 349.9 ;
      RECT  203.6 245.3 204.2 245.9 ;
      RECT  203.6 203.7 204.2 204.3 ;
      RECT  196.8 245.3 197.4 245.9 ;
      RECT  176.4 286.9 177.0 287.5 ;
      RECT  203.6 266.1 204.2 266.7 ;
      RECT  183.1 182.8 183.9 183.6 ;
      RECT  176.4 328.5 177.0 329.1 ;
      RECT  183.1 245.2 183.9 246.0 ;
      RECT  196.8 203.7 197.4 204.3 ;
      RECT  183.1 307.6 183.9 308.4 ;
      RECT  176.4 266.1 177.0 266.7 ;
      RECT  190.0 349.3 190.6 349.9 ;
      RECT  196.8 328.5 197.4 329.1 ;
      RECT  200.2 333.5 200.8 334.1 ;
      RECT  179.8 291.9 180.4 292.5 ;
      RECT  179.7 333.4 180.5 334.2 ;
      RECT  179.7 208.6 180.5 209.4 ;
      RECT  186.5 281.8 187.3 282.6 ;
      RECT  207.0 344.3 207.6 344.9 ;
      RECT  200.2 250.3 200.8 250.9 ;
      RECT  193.4 261.1 194.0 261.7 ;
      RECT  173.0 354.3 173.6 354.9 ;
      RECT  207.0 177.9 207.6 178.5 ;
      RECT  173.0 240.3 173.6 240.9 ;
      RECT  179.8 302.7 180.4 303.3 ;
      RECT  179.8 312.7 180.4 313.3 ;
      RECT  173.0 229.5 173.6 230.1 ;
      RECT  179.8 271.1 180.4 271.7 ;
      RECT  200.2 344.3 200.8 344.9 ;
      RECT  207.0 312.7 207.6 313.3 ;
      RECT  179.8 177.9 180.4 178.5 ;
      RECT  186.6 250.3 187.2 250.9 ;
      RECT  179.7 187.8 180.5 188.6 ;
      RECT  179.7 229.4 180.5 230.2 ;
      RECT  179.7 240.2 180.5 241.0 ;
      RECT  200.2 261.1 200.8 261.7 ;
      RECT  186.5 365.0 187.3 365.8 ;
      RECT  179.7 281.8 180.5 282.6 ;
      RECT  179.8 281.9 180.4 282.5 ;
      RECT  207.0 198.7 207.6 199.3 ;
      RECT  193.4 344.3 194.0 344.9 ;
      RECT  179.7 261.0 180.5 261.8 ;
      RECT  200.2 302.7 200.8 303.3 ;
      RECT  200.2 302.7 200.8 303.3 ;
      RECT  173.0 333.5 173.6 334.1 ;
      RECT  193.4 208.7 194.0 209.3 ;
      RECT  173.0 344.3 173.6 344.9 ;
      RECT  186.5 177.8 187.3 178.6 ;
      RECT  186.6 291.9 187.2 292.5 ;
      RECT  193.4 365.1 194.0 365.7 ;
      RECT  179.7 177.8 180.5 178.6 ;
      RECT  193.4 354.3 194.0 354.9 ;
      RECT  193.4 177.9 194.0 178.5 ;
      RECT  179.8 208.7 180.4 209.3 ;
      RECT  179.7 302.6 180.5 303.4 ;
      RECT  179.8 261.1 180.4 261.7 ;
      RECT  193.4 323.5 194.0 324.1 ;
      RECT  179.7 344.2 180.5 345.0 ;
      RECT  200.2 281.9 200.8 282.5 ;
      RECT  200.2 229.5 200.8 230.1 ;
      RECT  173.0 198.7 173.6 199.3 ;
      RECT  200.2 229.5 200.8 230.1 ;
      RECT  186.5 291.8 187.3 292.6 ;
      RECT  207.0 229.5 207.6 230.1 ;
      RECT  186.6 240.3 187.2 240.9 ;
      RECT  179.7 271.0 180.5 271.8 ;
      RECT  186.5 323.4 187.3 324.2 ;
      RECT  173.0 281.9 173.6 282.5 ;
      RECT  186.6 261.1 187.2 261.7 ;
      RECT  179.8 323.5 180.4 324.1 ;
      RECT  173.0 323.5 173.6 324.1 ;
      RECT  179.7 323.4 180.5 324.2 ;
      RECT  179.7 312.6 180.5 313.4 ;
      RECT  207.0 208.7 207.6 209.3 ;
      RECT  200.2 312.7 200.8 313.3 ;
      RECT  200.2 312.7 200.8 313.3 ;
      RECT  193.4 291.9 194.0 292.5 ;
      RECT  207.0 354.3 207.6 354.9 ;
      RECT  186.6 177.9 187.2 178.5 ;
      RECT  193.4 187.9 194.0 188.5 ;
      RECT  186.5 261.0 187.3 261.8 ;
      RECT  179.8 354.3 180.4 354.9 ;
      RECT  186.5 344.2 187.3 345.0 ;
      RECT  173.0 208.7 173.6 209.3 ;
      RECT  186.5 354.2 187.3 355.0 ;
      RECT  207.0 365.1 207.6 365.7 ;
      RECT  179.8 333.5 180.4 334.1 ;
      RECT  179.8 229.5 180.4 230.1 ;
      RECT  193.4 312.7 194.0 313.3 ;
      RECT  186.6 365.1 187.2 365.7 ;
      RECT  186.6 312.7 187.2 313.3 ;
      RECT  186.5 271.0 187.3 271.8 ;
      RECT  200.2 291.9 200.8 292.5 ;
      RECT  173.0 187.9 173.6 188.5 ;
      RECT  186.6 271.1 187.2 271.7 ;
      RECT  186.5 219.4 187.3 220.2 ;
      RECT  186.5 302.6 187.3 303.4 ;
      RECT  179.7 291.8 180.5 292.6 ;
      RECT  200.2 365.1 200.8 365.7 ;
      RECT  207.0 302.7 207.6 303.3 ;
      RECT  207.0 261.1 207.6 261.7 ;
      RECT  179.8 250.3 180.4 250.9 ;
      RECT  200.2 271.1 200.8 271.7 ;
      RECT  173.0 261.1 173.6 261.7 ;
      RECT  186.6 281.9 187.2 282.5 ;
      RECT  186.5 312.6 187.3 313.4 ;
      RECT  193.4 229.5 194.0 230.1 ;
      RECT  179.8 365.1 180.4 365.7 ;
      RECT  179.8 344.3 180.4 344.9 ;
      RECT  207.0 333.5 207.6 334.1 ;
      RECT  186.6 344.3 187.2 344.9 ;
      RECT  207.0 250.3 207.6 250.9 ;
      RECT  186.5 208.6 187.3 209.4 ;
      RECT  186.5 240.2 187.3 241.0 ;
      RECT  207.0 240.3 207.6 240.9 ;
      RECT  173.0 312.7 173.6 313.3 ;
      RECT  193.4 198.7 194.0 199.3 ;
      RECT  179.7 198.6 180.5 199.4 ;
      RECT  207.0 187.9 207.6 188.5 ;
      RECT  186.5 250.2 187.3 251.0 ;
      RECT  200.2 219.5 200.8 220.1 ;
      RECT  200.2 354.3 200.8 354.9 ;
      RECT  200.2 323.5 200.8 324.1 ;
      RECT  186.5 187.8 187.3 188.6 ;
      RECT  186.6 219.5 187.2 220.1 ;
      RECT  193.4 281.9 194.0 282.5 ;
      RECT  179.8 187.9 180.4 188.5 ;
      RECT  179.7 250.2 180.5 251.0 ;
      RECT  186.6 323.5 187.2 324.1 ;
      RECT  179.8 219.5 180.4 220.1 ;
      RECT  200.2 177.9 200.8 178.5 ;
      RECT  207.0 219.5 207.6 220.1 ;
      RECT  186.6 208.7 187.2 209.3 ;
      RECT  186.5 198.6 187.3 199.4 ;
      RECT  179.7 354.2 180.5 355.0 ;
      RECT  207.0 271.1 207.6 271.7 ;
      RECT  173.0 291.9 173.6 292.5 ;
      RECT  173.0 271.1 173.6 271.7 ;
      RECT  193.4 219.5 194.0 220.1 ;
      RECT  193.4 240.3 194.0 240.9 ;
      RECT  186.5 333.4 187.3 334.2 ;
      RECT  193.4 271.1 194.0 271.7 ;
      RECT  173.0 177.9 173.6 178.5 ;
      RECT  186.5 229.4 187.3 230.2 ;
      RECT  200.2 187.9 200.8 188.5 ;
      RECT  186.6 229.5 187.2 230.1 ;
      RECT  173.0 302.7 173.6 303.3 ;
      RECT  179.8 240.3 180.4 240.9 ;
      RECT  207.0 291.9 207.6 292.5 ;
      RECT  193.4 333.5 194.0 334.1 ;
      RECT  207.0 323.5 207.6 324.1 ;
      RECT  186.6 187.9 187.2 188.5 ;
      RECT  179.8 198.7 180.4 199.3 ;
      RECT  186.6 333.5 187.2 334.1 ;
      RECT  200.2 208.7 200.8 209.3 ;
      RECT  173.0 365.1 173.6 365.7 ;
      RECT  173.0 219.5 173.6 220.1 ;
      RECT  193.4 302.7 194.0 303.3 ;
      RECT  179.7 365.0 180.5 365.8 ;
      RECT  200.2 198.7 200.8 199.3 ;
      RECT  207.0 281.9 207.6 282.5 ;
      RECT  179.7 219.4 180.5 220.2 ;
      RECT  193.4 250.3 194.0 250.9 ;
      RECT  173.0 250.3 173.6 250.9 ;
      RECT  200.2 240.3 200.8 240.9 ;
      RECT  186.6 354.3 187.2 354.9 ;
      RECT  186.6 302.7 187.2 303.3 ;
      RECT  186.6 198.7 187.2 199.3 ;
      RECT  183.6 166.8 184.4 167.6 ;
      RECT  190.4 166.8 191.2 167.6 ;
      RECT  197.2 166.8 198.0 167.6 ;
      RECT  183.6 166.8 184.4 167.6 ;
      RECT  197.2 166.8 198.0 167.6 ;
      RECT  190.4 166.8 191.2 167.6 ;
      RECT  192.3 132.6 193.1 133.4 ;
      RECT  199.1 132.6 199.9 133.4 ;
      RECT  193.3 146.0 194.1 146.8 ;
      RECT  200.1 146.0 200.9 146.8 ;
      RECT  197.5 81.2 198.3 82.0 ;
      RECT  190.1 98.6 190.9 99.4 ;
      RECT  196.9 98.6 197.7 99.4 ;
      RECT  190.7 81.2 191.5 82.0 ;
      RECT  190.7 87.8 191.5 88.6 ;
      RECT  198.9 92.2 199.7 93.0 ;
      RECT  192.1 92.2 192.9 93.0 ;
      RECT  196.1 106.8 196.9 107.6 ;
      RECT  189.3 106.8 190.1 107.6 ;
      RECT  197.5 87.8 198.3 88.6 ;
      RECT  190.7 82.0 191.5 81.2 ;
      RECT  190.1 99.4 190.9 98.6 ;
      RECT  196.9 99.4 197.7 98.6 ;
      RECT  199.1 133.4 199.9 132.6 ;
      RECT  183.6 167.6 184.4 166.8 ;
      RECT  197.2 167.6 198.0 166.8 ;
      RECT  197.5 82.0 198.3 81.2 ;
      RECT  190.4 167.6 191.2 166.8 ;
      RECT  192.3 133.4 193.1 132.6 ;
      RECT  198.9 93.0 199.7 92.2 ;
      RECT  200.1 146.8 200.9 146.0 ;
      RECT  196.1 107.6 196.9 106.8 ;
      RECT  192.1 93.0 192.9 92.2 ;
      RECT  197.5 88.6 198.3 87.8 ;
      RECT  193.3 146.8 194.1 146.0 ;
      RECT  189.3 107.6 190.1 106.8 ;
      RECT  190.7 88.6 191.5 87.8 ;
      RECT  93.1 224.8 93.9 225.6 ;
      RECT  93.1 204.0 93.9 204.8 ;
      RECT  93.1 204.0 93.9 204.8 ;
      RECT  93.1 224.8 93.9 225.6 ;
      RECT  108.1 204.0 108.9 204.8 ;
      RECT  108.1 204.0 108.9 204.8 ;
      RECT  108.1 224.8 108.9 225.6 ;
      RECT  108.1 224.8 108.9 225.6 ;
      RECT  108.1 193.6 108.9 194.4 ;
      RECT  93.1 193.6 93.9 194.4 ;
      RECT  108.1 214.4 108.9 215.2 ;
      RECT  108.1 235.2 108.9 236.0 ;
      RECT  93.1 235.2 93.9 236.0 ;
      RECT  93.1 214.4 93.9 215.2 ;
      RECT  93.1 276.8 93.9 277.6 ;
      RECT  93.1 256.0 93.9 256.8 ;
      RECT  93.1 256.0 93.9 256.8 ;
      RECT  93.1 276.8 93.9 277.6 ;
      RECT  108.1 256.0 108.9 256.8 ;
      RECT  108.1 256.0 108.9 256.8 ;
      RECT  108.1 276.8 108.9 277.6 ;
      RECT  108.1 276.8 108.9 277.6 ;
      RECT  108.1 245.6 108.9 246.4 ;
      RECT  93.1 245.6 93.9 246.4 ;
      RECT  108.1 266.4 108.9 267.2 ;
      RECT  108.1 287.2 108.9 288.0 ;
      RECT  93.1 287.2 93.9 288.0 ;
      RECT  93.1 266.4 93.9 267.2 ;
      RECT  152.0 204.0 152.8 204.8 ;
      RECT  152.0 204.0 152.8 204.8 ;
      RECT  152.0 308.0 152.8 308.8 ;
      RECT  108.1 224.8 108.9 225.6 ;
      RECT  108.1 204.0 108.9 204.8 ;
      RECT  108.1 256.0 108.9 256.8 ;
      RECT  152.0 266.4 152.8 267.2 ;
      RECT  152.0 266.4 152.8 267.2 ;
      RECT  93.1 204.0 93.9 204.8 ;
      RECT  152.0 224.8 152.8 225.6 ;
      RECT  152.0 224.8 152.8 225.6 ;
      RECT  108.1 276.8 108.9 277.6 ;
      RECT  152.0 349.6 152.8 350.4 ;
      RECT  152.0 287.2 152.8 288.0 ;
      RECT  152.0 287.2 152.8 288.0 ;
      RECT  93.1 224.8 93.9 225.6 ;
      RECT  93.1 256.0 93.9 256.8 ;
      RECT  152.0 328.8 152.8 329.6 ;
      RECT  93.1 276.8 93.9 277.6 ;
      RECT  152.0 245.6 152.8 246.4 ;
      RECT  108.1 193.6 108.9 194.4 ;
      RECT  108.1 266.4 108.9 267.2 ;
      RECT  152.0 339.2 152.8 340.0 ;
      RECT  108.1 235.2 108.9 236.0 ;
      RECT  93.1 235.2 93.9 236.0 ;
      RECT  93.1 287.2 93.9 288.0 ;
      RECT  152.0 276.8 152.8 277.6 ;
      RECT  108.1 287.2 108.9 288.0 ;
      RECT  152.0 256.0 152.8 256.8 ;
      RECT  152.0 360.0 152.8 360.8 ;
      RECT  152.0 193.6 152.8 194.4 ;
      RECT  93.1 266.4 93.9 267.2 ;
      RECT  108.1 214.4 108.9 215.2 ;
      RECT  152.0 297.6 152.8 298.4 ;
      RECT  152.0 235.2 152.8 236.0 ;
      RECT  93.1 245.6 93.9 246.4 ;
      RECT  93.1 214.4 93.9 215.2 ;
      RECT  152.0 318.4 152.8 319.2 ;
      RECT  152.0 214.4 152.8 215.2 ;
      RECT  93.1 193.6 93.9 194.4 ;
      RECT  108.1 245.6 108.9 246.4 ;
      RECT  167.5 245.6 168.3 246.4 ;
      RECT  167.5 349.6 168.3 350.4 ;
      RECT  167.5 224.8 168.3 225.6 ;
      RECT  167.5 224.8 168.3 225.6 ;
      RECT  167.5 204.0 168.3 204.8 ;
      RECT  167.5 204.0 168.3 204.8 ;
      RECT  167.5 266.4 168.3 267.2 ;
      RECT  167.5 266.4 168.3 267.2 ;
      RECT  167.5 287.2 168.3 288.0 ;
      RECT  167.5 287.2 168.3 288.0 ;
      RECT  167.5 308.0 168.3 308.8 ;
      RECT  167.5 328.8 168.3 329.6 ;
      RECT  167.5 214.4 168.3 215.2 ;
      RECT  167.5 318.4 168.3 319.2 ;
      RECT  167.5 256.0 168.3 256.8 ;
      RECT  167.5 193.6 168.3 194.4 ;
      RECT  167.5 339.2 168.3 340.0 ;
      RECT  167.5 297.6 168.3 298.4 ;
      RECT  167.5 276.8 168.3 277.6 ;
      RECT  167.5 235.2 168.3 236.0 ;
      RECT  167.5 360.0 168.3 360.8 ;
      RECT  93.1 204.0 93.9 204.8 ;
      RECT  152.0 287.2 152.8 288.0 ;
      RECT  167.5 245.6 168.3 246.4 ;
      RECT  167.5 287.2 168.3 288.0 ;
      RECT  152.0 328.8 152.8 329.6 ;
      RECT  152.0 245.6 152.8 246.4 ;
      RECT  108.1 224.8 108.9 225.6 ;
      RECT  108.1 256.0 108.9 256.8 ;
      RECT  167.5 266.4 168.3 267.2 ;
      RECT  152.0 266.4 152.8 267.2 ;
      RECT  93.1 256.0 93.9 256.8 ;
      RECT  152.0 224.8 152.8 225.6 ;
      RECT  152.0 308.0 152.8 308.8 ;
      RECT  108.1 276.8 108.9 277.6 ;
      RECT  93.1 224.8 93.9 225.6 ;
      RECT  167.5 224.8 168.3 225.6 ;
      RECT  152.0 204.0 152.8 204.8 ;
      RECT  152.0 349.6 152.8 350.4 ;
      RECT  167.5 204.0 168.3 204.8 ;
      RECT  167.5 349.6 168.3 350.4 ;
      RECT  167.5 308.0 168.3 308.8 ;
      RECT  93.1 276.8 93.9 277.6 ;
      RECT  108.1 204.0 108.9 204.8 ;
      RECT  167.5 328.8 168.3 329.6 ;
      RECT  167.5 297.6 168.3 298.4 ;
      RECT  167.5 339.2 168.3 340.0 ;
      RECT  93.1 235.2 93.9 236.0 ;
      RECT  108.1 193.6 108.9 194.4 ;
      RECT  167.5 256.0 168.3 256.8 ;
      RECT  167.5 193.6 168.3 194.4 ;
      RECT  93.1 266.4 93.9 267.2 ;
      RECT  152.0 276.8 152.8 277.6 ;
      RECT  167.5 318.4 168.3 319.2 ;
      RECT  152.0 193.6 152.8 194.4 ;
      RECT  93.1 287.2 93.9 288.0 ;
      RECT  152.0 214.4 152.8 215.2 ;
      RECT  152.0 256.0 152.8 256.8 ;
      RECT  167.5 235.2 168.3 236.0 ;
      RECT  108.1 235.2 108.9 236.0 ;
      RECT  167.5 214.4 168.3 215.2 ;
      RECT  108.1 214.4 108.9 215.2 ;
      RECT  93.1 193.6 93.9 194.4 ;
      RECT  108.1 245.6 108.9 246.4 ;
      RECT  152.0 339.2 152.8 340.0 ;
      RECT  108.1 266.4 108.9 267.2 ;
      RECT  167.5 360.0 168.3 360.8 ;
      RECT  152.0 360.0 152.8 360.8 ;
      RECT  93.1 214.4 93.9 215.2 ;
      RECT  152.0 297.6 152.8 298.4 ;
      RECT  93.1 245.6 93.9 246.4 ;
      RECT  108.1 287.2 108.9 288.0 ;
      RECT  152.0 235.2 152.8 236.0 ;
      RECT  152.0 318.4 152.8 319.2 ;
      RECT  167.5 276.8 168.3 277.6 ;
      RECT  108.1 224.8 108.9 225.6 ;
      RECT  183.6 166.8 184.4 167.6 ;
      RECT  203.6 224.5 204.2 225.1 ;
      RECT  203.6 328.5 204.2 329.1 ;
      RECT  190.0 203.7 190.6 204.3 ;
      RECT  183.1 266.0 183.9 266.8 ;
      RECT  190.0 328.5 190.6 329.1 ;
      RECT  108.1 256.0 108.9 256.8 ;
      RECT  190.0 224.5 190.6 225.1 ;
      RECT  167.5 266.4 168.3 267.2 ;
      RECT  196.8 307.7 197.4 308.3 ;
      RECT  93.1 256.0 93.9 256.8 ;
      RECT  196.8 349.3 197.4 349.9 ;
      RECT  167.5 328.8 168.3 329.6 ;
      RECT  196.8 370.1 197.4 370.7 ;
      RECT  167.5 349.6 168.3 350.4 ;
      RECT  183.1 182.8 183.9 183.6 ;
      RECT  183.1 245.2 183.9 246.0 ;
      RECT  190.0 349.3 190.6 349.9 ;
      RECT  108.1 276.8 108.9 277.6 ;
      RECT  93.1 204.0 93.9 204.8 ;
      RECT  203.6 307.7 204.2 308.3 ;
      RECT  152.0 349.6 152.8 350.4 ;
      RECT  183.1 328.4 183.9 329.2 ;
      RECT  183.1 224.4 183.9 225.2 ;
      RECT  190.4 166.8 191.2 167.6 ;
      RECT  196.8 266.1 197.4 266.7 ;
      RECT  190.0 245.3 190.6 245.9 ;
      RECT  176.4 245.3 177.0 245.9 ;
      RECT  176.4 349.3 177.0 349.9 ;
      RECT  199.1 132.6 199.9 133.4 ;
      RECT  197.5 81.2 198.3 82.0 ;
      RECT  176.4 224.5 177.0 225.1 ;
      RECT  190.0 307.7 190.6 308.3 ;
      RECT  196.8 224.5 197.4 225.1 ;
      RECT  203.6 349.3 204.2 349.9 ;
      RECT  93.1 276.8 93.9 277.6 ;
      RECT  196.8 245.3 197.4 245.9 ;
      RECT  176.4 286.9 177.0 287.5 ;
      RECT  196.8 203.7 197.4 204.3 ;
      RECT  197.2 166.8 198.0 167.6 ;
      RECT  93.1 224.8 93.9 225.6 ;
      RECT  152.0 266.4 152.8 267.2 ;
      RECT  152.0 204.0 152.8 204.8 ;
      RECT  167.5 204.0 168.3 204.8 ;
      RECT  152.0 328.8 152.8 329.6 ;
      RECT  196.8 182.9 197.4 183.5 ;
      RECT  196.8 286.9 197.4 287.5 ;
      RECT  176.4 182.9 177.0 183.5 ;
      RECT  203.6 370.1 204.2 370.7 ;
      RECT  108.1 204.0 108.9 204.8 ;
      RECT  196.9 98.6 197.7 99.4 ;
      RECT  183.1 203.6 183.9 204.4 ;
      RECT  203.6 182.9 204.2 183.5 ;
      RECT  152.0 245.6 152.8 246.4 ;
      RECT  190.1 98.6 190.9 99.4 ;
      RECT  190.0 370.1 190.6 370.7 ;
      RECT  176.4 307.7 177.0 308.3 ;
      RECT  203.6 203.7 204.2 204.3 ;
      RECT  203.6 266.1 204.2 266.7 ;
      RECT  176.4 328.5 177.0 329.1 ;
      RECT  152.0 287.2 152.8 288.0 ;
      RECT  152.0 308.0 152.8 308.8 ;
      RECT  176.4 266.1 177.0 266.7 ;
      RECT  190.0 182.9 190.6 183.5 ;
      RECT  167.5 287.2 168.3 288.0 ;
      RECT  190.0 286.9 190.6 287.5 ;
      RECT  176.4 370.1 177.0 370.7 ;
      RECT  183.1 286.8 183.9 287.6 ;
      RECT  203.6 286.9 204.2 287.5 ;
      RECT  167.5 308.0 168.3 308.8 ;
      RECT  183.1 370.0 183.9 370.8 ;
      RECT  176.4 203.7 177.0 204.3 ;
      RECT  167.5 224.8 168.3 225.6 ;
      RECT  190.0 266.1 190.6 266.7 ;
      RECT  167.5 245.6 168.3 246.4 ;
      RECT  183.1 349.2 183.9 350.0 ;
      RECT  190.7 81.2 191.5 82.0 ;
      RECT  192.3 132.6 193.1 133.4 ;
      RECT  152.0 224.8 152.8 225.6 ;
      RECT  203.6 245.3 204.2 245.9 ;
      RECT  183.1 307.6 183.9 308.4 ;
      RECT  196.8 328.5 197.4 329.1 ;
      RECT  200.2 333.5 200.8 334.1 ;
      RECT  167.5 276.8 168.3 277.6 ;
      RECT  179.8 291.9 180.4 292.5 ;
      RECT  179.7 333.4 180.5 334.2 ;
      RECT  179.7 208.6 180.5 209.4 ;
      RECT  186.5 281.8 187.3 282.6 ;
      RECT  93.1 266.4 93.9 267.2 ;
      RECT  207.0 344.3 207.6 344.9 ;
      RECT  152.0 339.2 152.8 340.0 ;
      RECT  200.2 250.3 200.8 250.9 ;
      RECT  193.4 261.1 194.0 261.7 ;
      RECT  173.0 354.3 173.6 354.9 ;
      RECT  207.0 177.9 207.6 178.5 ;
      RECT  173.0 240.3 173.6 240.9 ;
      RECT  190.7 87.8 191.5 88.6 ;
      RECT  152.0 256.0 152.8 256.8 ;
      RECT  179.8 302.7 180.4 303.3 ;
      RECT  179.8 312.7 180.4 313.3 ;
      RECT  173.0 229.5 173.6 230.1 ;
      RECT  179.8 271.1 180.4 271.7 ;
      RECT  200.2 344.3 200.8 344.9 ;
      RECT  207.0 312.7 207.6 313.3 ;
      RECT  179.8 177.9 180.4 178.5 ;
      RECT  186.6 250.3 187.2 250.9 ;
      RECT  179.7 187.8 180.5 188.6 ;
      RECT  179.7 229.4 180.5 230.2 ;
      RECT  167.5 235.2 168.3 236.0 ;
      RECT  179.7 240.2 180.5 241.0 ;
      RECT  200.2 261.1 200.8 261.7 ;
      RECT  186.5 365.0 187.3 365.8 ;
      RECT  179.7 281.8 180.5 282.6 ;
      RECT  179.8 281.9 180.4 282.5 ;
      RECT  207.0 198.7 207.6 199.3 ;
      RECT  193.4 344.3 194.0 344.9 ;
      RECT  179.7 261.0 180.5 261.8 ;
      RECT  200.2 302.7 200.8 303.3 ;
      RECT  152.0 360.0 152.8 360.8 ;
      RECT  173.0 333.5 173.6 334.1 ;
      RECT  189.3 106.8 190.1 107.6 ;
      RECT  193.4 208.7 194.0 209.3 ;
      RECT  173.0 344.3 173.6 344.9 ;
      RECT  93.1 193.6 93.9 194.4 ;
      RECT  186.5 177.8 187.3 178.6 ;
      RECT  186.6 291.9 187.2 292.5 ;
      RECT  193.4 365.1 194.0 365.7 ;
      RECT  179.7 177.8 180.5 178.6 ;
      RECT  193.4 354.3 194.0 354.9 ;
      RECT  193.4 177.9 194.0 178.5 ;
      RECT  179.8 208.7 180.4 209.3 ;
      RECT  179.7 302.6 180.5 303.4 ;
      RECT  152.0 193.6 152.8 194.4 ;
      RECT  179.8 261.1 180.4 261.7 ;
      RECT  108.1 287.2 108.9 288.0 ;
      RECT  193.4 323.5 194.0 324.1 ;
      RECT  179.7 344.2 180.5 345.0 ;
      RECT  200.2 281.9 200.8 282.5 ;
      RECT  200.2 229.5 200.8 230.1 ;
      RECT  173.0 198.7 173.6 199.3 ;
      RECT  186.5 291.8 187.3 292.6 ;
      RECT  207.0 229.5 207.6 230.1 ;
      RECT  108.1 193.6 108.9 194.4 ;
      RECT  186.6 240.3 187.2 240.9 ;
      RECT  179.7 271.0 180.5 271.8 ;
      RECT  186.5 323.4 187.3 324.2 ;
      RECT  173.0 281.9 173.6 282.5 ;
      RECT  186.6 261.1 187.2 261.7 ;
      RECT  179.8 323.5 180.4 324.1 ;
      RECT  173.0 323.5 173.6 324.1 ;
      RECT  152.0 235.2 152.8 236.0 ;
      RECT  179.7 323.4 180.5 324.2 ;
      RECT  179.7 312.6 180.5 313.4 ;
      RECT  207.0 208.7 207.6 209.3 ;
      RECT  200.2 312.7 200.8 313.3 ;
      RECT  152.0 214.4 152.8 215.2 ;
      RECT  108.1 235.2 108.9 236.0 ;
      RECT  193.4 291.9 194.0 292.5 ;
      RECT  207.0 354.3 207.6 354.9 ;
      RECT  186.6 177.9 187.2 178.5 ;
      RECT  193.4 187.9 194.0 188.5 ;
      RECT  186.5 261.0 187.3 261.8 ;
      RECT  179.8 354.3 180.4 354.9 ;
      RECT  200.1 146.0 200.9 146.8 ;
      RECT  186.5 344.2 187.3 345.0 ;
      RECT  173.0 208.7 173.6 209.3 ;
      RECT  167.5 297.6 168.3 298.4 ;
      RECT  186.5 354.2 187.3 355.0 ;
      RECT  207.0 365.1 207.6 365.7 ;
      RECT  179.8 333.5 180.4 334.1 ;
      RECT  179.8 229.5 180.4 230.1 ;
      RECT  152.0 297.6 152.8 298.4 ;
      RECT  193.4 312.7 194.0 313.3 ;
      RECT  108.1 245.6 108.9 246.4 ;
      RECT  186.6 365.1 187.2 365.7 ;
      RECT  93.1 235.2 93.9 236.0 ;
      RECT  186.6 312.7 187.2 313.3 ;
      RECT  186.5 271.0 187.3 271.8 ;
      RECT  200.2 291.9 200.8 292.5 ;
      RECT  173.0 187.9 173.6 188.5 ;
      RECT  186.6 271.1 187.2 271.7 ;
      RECT  186.5 219.4 187.3 220.2 ;
      RECT  186.5 302.6 187.3 303.4 ;
      RECT  179.7 291.8 180.5 292.6 ;
      RECT  200.2 365.1 200.8 365.7 ;
      RECT  207.0 302.7 207.6 303.3 ;
      RECT  207.0 261.1 207.6 261.7 ;
      RECT  179.8 250.3 180.4 250.9 ;
      RECT  200.2 271.1 200.8 271.7 ;
      RECT  173.0 261.1 173.6 261.7 ;
      RECT  186.6 281.9 187.2 282.5 ;
      RECT  186.5 312.6 187.3 313.4 ;
      RECT  93.1 245.6 93.9 246.4 ;
      RECT  193.4 229.5 194.0 230.1 ;
      RECT  179.8 365.1 180.4 365.7 ;
      RECT  179.8 344.3 180.4 344.9 ;
      RECT  207.0 333.5 207.6 334.1 ;
      RECT  186.6 344.3 187.2 344.9 ;
      RECT  207.0 250.3 207.6 250.9 ;
      RECT  186.5 208.6 187.3 209.4 ;
      RECT  186.5 240.2 187.3 241.0 ;
      RECT  207.0 240.3 207.6 240.9 ;
      RECT  167.5 318.4 168.3 319.2 ;
      RECT  173.0 312.7 173.6 313.3 ;
      RECT  193.4 198.7 194.0 199.3 ;
      RECT  196.1 106.8 196.9 107.6 ;
      RECT  179.7 198.6 180.5 199.4 ;
      RECT  207.0 187.9 207.6 188.5 ;
      RECT  192.1 92.2 192.9 93.0 ;
      RECT  186.5 250.2 187.3 251.0 ;
      RECT  200.2 219.5 200.8 220.1 ;
      RECT  152.0 276.8 152.8 277.6 ;
      RECT  200.2 354.3 200.8 354.9 ;
      RECT  200.2 323.5 200.8 324.1 ;
      RECT  186.5 187.8 187.3 188.6 ;
      RECT  186.6 219.5 187.2 220.1 ;
      RECT  108.1 214.4 108.9 215.2 ;
      RECT  193.4 281.9 194.0 282.5 ;
      RECT  179.8 187.9 180.4 188.5 ;
      RECT  179.7 250.2 180.5 251.0 ;
      RECT  167.5 214.4 168.3 215.2 ;
      RECT  186.6 323.5 187.2 324.1 ;
      RECT  179.8 219.5 180.4 220.1 ;
      RECT  167.5 339.2 168.3 340.0 ;
      RECT  200.2 177.9 200.8 178.5 ;
      RECT  152.0 318.4 152.8 319.2 ;
      RECT  207.0 219.5 207.6 220.1 ;
      RECT  186.6 208.7 187.2 209.3 ;
      RECT  193.3 146.0 194.1 146.8 ;
      RECT  186.5 198.6 187.3 199.4 ;
      RECT  179.7 354.2 180.5 355.0 ;
      RECT  207.0 271.1 207.6 271.7 ;
      RECT  173.0 291.9 173.6 292.5 ;
      RECT  173.0 271.1 173.6 271.7 ;
      RECT  193.4 219.5 194.0 220.1 ;
      RECT  197.5 87.8 198.3 88.6 ;
      RECT  193.4 240.3 194.0 240.9 ;
      RECT  186.5 333.4 187.3 334.2 ;
      RECT  193.4 271.1 194.0 271.7 ;
      RECT  173.0 177.9 173.6 178.5 ;
      RECT  186.5 229.4 187.3 230.2 ;
      RECT  200.2 187.9 200.8 188.5 ;
      RECT  186.6 229.5 187.2 230.1 ;
      RECT  173.0 302.7 173.6 303.3 ;
      RECT  179.8 240.3 180.4 240.9 ;
      RECT  207.0 291.9 207.6 292.5 ;
      RECT  193.4 333.5 194.0 334.1 ;
      RECT  207.0 323.5 207.6 324.1 ;
      RECT  167.5 256.0 168.3 256.8 ;
      RECT  186.6 187.9 187.2 188.5 ;
      RECT  179.8 198.7 180.4 199.3 ;
      RECT  167.5 360.0 168.3 360.8 ;
      RECT  93.1 214.4 93.9 215.2 ;
      RECT  186.6 333.5 187.2 334.1 ;
      RECT  200.2 208.7 200.8 209.3 ;
      RECT  173.0 365.1 173.6 365.7 ;
      RECT  173.0 219.5 173.6 220.1 ;
      RECT  193.4 302.7 194.0 303.3 ;
      RECT  179.7 365.0 180.5 365.8 ;
      RECT  198.9 92.2 199.7 93.0 ;
      RECT  200.2 198.7 200.8 199.3 ;
      RECT  207.0 281.9 207.6 282.5 ;
      RECT  179.7 219.4 180.5 220.2 ;
      RECT  167.5 193.6 168.3 194.4 ;
      RECT  193.4 250.3 194.0 250.9 ;
      RECT  173.0 250.3 173.6 250.9 ;
      RECT  200.2 240.3 200.8 240.9 ;
      RECT  93.1 287.2 93.9 288.0 ;
      RECT  108.1 266.4 108.9 267.2 ;
      RECT  186.6 354.3 187.2 354.9 ;
      RECT  186.6 302.7 187.2 303.3 ;
      RECT  186.6 198.7 187.2 199.3 ;
      RECT  2.0 21.2 2.8 22.0 ;
      RECT  2.0 1.2 2.8 2.0 ;
      RECT  2.0 41.2 2.8 42.0 ;
      RECT  3.5 340.4 2.7 341.2 ;
      RECT  24.0 262.0 23.2 262.8 ;
      RECT  24.0 222.8 23.2 223.6 ;
      RECT  3.5 183.6 2.7 184.4 ;
      RECT  24.0 301.2 23.2 302.0 ;
      RECT  3.5 222.8 2.7 223.6 ;
      RECT  3.5 262.0 2.7 262.8 ;
      RECT  24.0 340.4 23.2 341.2 ;
      RECT  24.0 183.6 23.2 184.4 ;
      RECT  3.5 301.2 2.7 302.0 ;
      RECT  24.0 320.8 23.2 321.6 ;
      RECT  24.0 203.2 23.2 204.0 ;
      RECT  24.0 242.4 23.2 243.2 ;
      RECT  24.0 164.0 23.2 164.8 ;
      RECT  3.5 242.4 2.7 243.2 ;
      RECT  24.0 281.6 23.2 282.4 ;
      RECT  3.5 281.6 2.7 282.4 ;
      RECT  3.5 164.0 2.7 164.8 ;
      RECT  3.5 320.8 2.7 321.6 ;
      RECT  3.5 203.2 2.7 204.0 ;
      RECT  23.2 183.6 24.0 184.4 ;
      RECT  23.2 262.0 24.0 262.8 ;
      RECT  2.7 222.8 3.5 223.6 ;
      RECT  77.6 61.2 78.4 62.0 ;
      RECT  77.6 141.2 78.4 142.0 ;
      RECT  77.6 21.2 78.4 22.0 ;
      RECT  2.7 340.4 3.5 341.2 ;
      RECT  23.2 301.2 24.0 302.0 ;
      RECT  2.0 21.2 2.8 22.0 ;
      RECT  23.2 222.8 24.0 223.6 ;
      RECT  2.7 301.2 3.5 302.0 ;
      RECT  2.7 262.0 3.5 262.8 ;
      RECT  2.7 183.6 3.5 184.4 ;
      RECT  23.2 340.4 24.0 341.2 ;
      RECT  77.6 101.2 78.4 102.0 ;
      RECT  23.2 320.8 24.0 321.6 ;
      RECT  23.2 281.6 24.0 282.4 ;
      RECT  2.7 203.2 3.5 204.0 ;
      RECT  77.6 81.2 78.4 82.0 ;
      RECT  2.7 281.6 3.5 282.4 ;
      RECT  2.0 41.2 2.8 42.0 ;
      RECT  23.2 203.2 24.0 204.0 ;
      RECT  2.7 164.0 3.5 164.8 ;
      RECT  77.6 1.2 78.4 2.0 ;
      RECT  2.7 320.8 3.5 321.6 ;
      RECT  2.7 242.4 3.5 243.2 ;
      RECT  77.6 121.2 78.4 122.0 ;
      RECT  23.2 164.0 24.0 164.8 ;
      RECT  23.2 242.4 24.0 243.2 ;
      RECT  2.0 1.2 2.8 2.0 ;
      RECT  77.6 161.2 78.4 162.0 ;
      RECT  77.6 41.2 78.4 42.0 ;
      RECT  57.6 346.7 79.4 347.3 ;
      RECT  68.1 403.2 68.9 404.0 ;
      RECT  68.1 363.2 68.9 364.0 ;
      RECT  68.1 383.2 68.9 384.0 ;
      RECT  68.1 343.2 68.9 344.0 ;
      RECT  68.1 423.2 68.9 424.0 ;
      RECT  173.3 51.1 216.9 51.7 ;
      RECT  205.6 67.6 206.4 68.4 ;
      RECT  183.8 67.6 184.6 68.4 ;
      RECT  205.6 47.6 206.4 48.4 ;
      RECT  183.8 47.6 184.6 48.4 ;
   LAYER  m4 ;
   END
   END    sram_2_16_scn4m_subm
END    LIBRARY
