
.SUBCKT col_cap_cell_1rw_1r bl0 br0 bl1 br1 vdd

.ENDS
