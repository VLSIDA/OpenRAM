magic
tech scmos
timestamp 1577067400
<< nwell >>
rect 0 46 54 75
<< pwell >>
rect 0 0 54 46
<< ntransistor >>
rect 14 33 16 37
rect 22 29 24 37
rect 30 29 32 37
rect 38 33 40 37
rect 14 17 16 23
rect 22 17 24 23
rect 30 17 32 23
rect 38 17 40 23
<< ptransistor >>
rect 22 54 24 57
rect 30 54 32 57
<< ndiffusion >>
rect 13 33 14 37
rect 16 33 17 37
rect 21 33 22 37
rect 17 29 22 33
rect 24 29 25 37
rect 29 29 30 37
rect 32 33 33 37
rect 37 33 38 37
rect 40 33 41 37
rect 32 29 37 33
rect 9 21 14 23
rect 13 17 14 21
rect 16 17 22 23
rect 24 17 25 23
rect 29 17 30 23
rect 32 17 38 23
rect 40 21 45 23
rect 40 17 41 21
<< pdiffusion >>
rect 21 54 22 57
rect 24 54 25 57
rect 29 54 30 57
rect 32 54 33 57
<< ndcontact >>
rect 9 33 13 37
rect 17 33 21 37
rect 25 29 29 37
rect 33 33 37 37
rect 41 33 45 37
rect 9 17 13 21
rect 25 17 29 23
rect 41 17 45 21
<< pdcontact >>
rect 17 54 21 58
rect 25 54 29 58
rect 33 54 37 58
<< psubstratepcontact >>
rect 25 9 29 13
<< nsubstratencontact >>
rect 25 68 29 72
<< polysilicon >>
rect 22 57 24 60
rect 30 57 32 60
rect 22 44 24 54
rect 30 51 32 54
rect 31 47 32 51
rect 14 37 16 44
rect 22 40 23 44
rect 22 37 24 40
rect 30 37 32 47
rect 38 37 40 44
rect 14 31 16 33
rect 38 31 40 33
rect 14 23 16 24
rect 22 23 24 29
rect 30 23 32 29
rect 38 23 40 24
rect 14 15 16 17
rect 22 15 24 17
rect 30 15 32 17
rect 38 15 40 17
<< polycontact >>
rect 27 47 31 51
rect 10 40 14 44
rect 23 40 27 44
rect 40 40 44 44
rect 12 24 16 28
rect 38 24 42 28
<< metal1 >>
rect 0 68 25 72
rect 29 68 54 72
rect 0 61 54 65
rect 10 44 14 61
rect 17 51 20 54
rect 17 47 27 51
rect 17 37 20 47
rect 34 44 37 54
rect 27 40 37 44
rect 40 44 44 61
rect 34 37 37 40
rect 2 33 9 37
rect 45 33 52 37
rect 25 23 29 29
rect 25 13 29 17
rect 0 9 25 13
rect 29 9 54 13
rect 0 2 16 6
rect 20 2 34 6
rect 38 2 54 6
<< m2contact >>
rect 25 68 29 72
rect 25 54 29 58
rect 16 24 20 28
rect 34 24 38 28
rect 16 2 20 6
rect 34 2 38 6
<< metal2 >>
rect 2 0 6 72
rect 9 0 13 72
rect 25 58 29 68
rect 16 6 20 24
rect 34 6 38 24
rect 41 0 45 72
rect 48 0 52 72
<< comment >>
rect 0 0 54 70
<< labels >>
rlabel metal1 19 63 19 63 1 wl0
rlabel metal1 19 70 19 70 5 vdd
rlabel metal1 27 4 27 4 1 wl1
rlabel psubstratepcontact 27 11 27 11 1 gnd
rlabel metal2 4 7 4 7 2 bl0
rlabel metal2 11 7 11 7 1 bl1
rlabel metal2 43 7 43 7 1 br1
rlabel metal2 50 7 50 7 8 br0
rlabel polycontact 29 49 29 49 1 Q
rlabel polycontact 25 42 25 42 1 Q_bar
<< end >>
