VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 1000 ;
END UNITS
SITE  MacroSite
   CLASS Core ;
   SIZE 106535.0 by 115787.5 ;
END  MacroSite
MACRO sram_1rw_32b_256w_1bank_freepdk45
   CLASS BLOCK ;
   SIZE 106535.0 BY 115787.5 ;
   SYMMETRY X Y R90 ;
   SITE MacroSite ;
   PIN DATA[0]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  16067.5 35.0 16137.5 175.0 ;
      END
   END DATA[0]
   PIN DATA[1]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  18887.5 35.0 18957.5 175.0 ;
      END
   END DATA[1]
   PIN DATA[2]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  21707.5 35.0 21777.5 175.0 ;
      END
   END DATA[2]
   PIN DATA[3]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  24527.5 35.0 24597.5 175.0 ;
      END
   END DATA[3]
   PIN DATA[4]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  27347.5 35.0 27417.5 175.0 ;
      END
   END DATA[4]
   PIN DATA[5]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  30167.5 35.0 30237.5 175.0 ;
      END
   END DATA[5]
   PIN DATA[6]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  32987.5 35.0 33057.5 175.0 ;
      END
   END DATA[6]
   PIN DATA[7]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  35807.5 35.0 35877.5 175.0 ;
      END
   END DATA[7]
   PIN DATA[8]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  38627.5 35.0 38697.5 175.0 ;
      END
   END DATA[8]
   PIN DATA[9]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  41447.5 35.0 41517.5 175.0 ;
      END
   END DATA[9]
   PIN DATA[10]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  44267.5 35.0 44337.5 175.0 ;
      END
   END DATA[10]
   PIN DATA[11]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  47087.5 35.0 47157.5 175.0 ;
      END
   END DATA[11]
   PIN DATA[12]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  49907.5 35.0 49977.5 175.0 ;
      END
   END DATA[12]
   PIN DATA[13]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  52727.5 35.0 52797.5 175.0 ;
      END
   END DATA[13]
   PIN DATA[14]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  55547.5 35.0 55617.5 175.0 ;
      END
   END DATA[14]
   PIN DATA[15]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  58367.5 35.0 58437.5 175.0 ;
      END
   END DATA[15]
   PIN DATA[16]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  61187.5 35.0 61257.5 175.0 ;
      END
   END DATA[16]
   PIN DATA[17]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  64007.5 35.0 64077.5 175.0 ;
      END
   END DATA[17]
   PIN DATA[18]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  66827.5 35.0 66897.5 175.0 ;
      END
   END DATA[18]
   PIN DATA[19]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  69647.5 35.0 69717.5 175.0 ;
      END
   END DATA[19]
   PIN DATA[20]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  72467.5 35.0 72537.5 175.0 ;
      END
   END DATA[20]
   PIN DATA[21]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  75287.5 35.0 75357.5 175.0 ;
      END
   END DATA[21]
   PIN DATA[22]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  78107.5 35.0 78177.5 175.0 ;
      END
   END DATA[22]
   PIN DATA[23]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  80927.5 35.0 80997.5 175.0 ;
      END
   END DATA[23]
   PIN DATA[24]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  83747.5 35.0 83817.5 175.0 ;
      END
   END DATA[24]
   PIN DATA[25]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  86567.5 35.0 86637.5 175.0 ;
      END
   END DATA[25]
   PIN DATA[26]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  89387.5 35.0 89457.5 175.0 ;
      END
   END DATA[26]
   PIN DATA[27]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  92207.5 35.0 92277.5 175.0 ;
      END
   END DATA[27]
   PIN DATA[28]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  95027.5 35.0 95097.5 175.0 ;
      END
   END DATA[28]
   PIN DATA[29]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  97847.5 35.0 97917.5 175.0 ;
      END
   END DATA[29]
   PIN DATA[30]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  100667.5 35.0 100737.5 175.0 ;
      END
   END DATA[30]
   PIN DATA[31]
      DIRECTION INOUT ;
      PORT
         LAYER metal2 ;
         RECT  103487.5 35.0 103557.5 175.0 ;
      END
   END DATA[31]
   PIN ADDR[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  4175.0 11077.5 4655.0 11147.5 ;
      END
   END ADDR[0]
   PIN ADDR[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  4175.0 10372.5 4655.0 10442.5 ;
      END
   END ADDR[1]
   PIN ADDR[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  4175.0 9667.5 4655.0 9737.5 ;
      END
   END ADDR[2]
   PIN ADDR[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  4175.0 8962.5 4655.0 9032.5 ;
      END
   END ADDR[3]
   PIN ADDR[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  4175.0 8257.5 4655.0 8327.5 ;
      END
   END ADDR[4]
   PIN ADDR[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  4175.0 7552.5 4655.0 7622.5 ;
      END
   END ADDR[5]
   PIN ADDR[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  4175.0 6847.5 4655.0 6917.5 ;
      END
   END ADDR[6]
   PIN ADDR[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  4175.0 6142.5 4655.0 6212.5 ;
      END
   END ADDR[7]
   PIN CSb
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1187.5 28155.0 1257.5 28295.0 ;
      END
   END CSb
   PIN WEb
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  1892.5 28155.0 1962.5 28295.0 ;
      END
   END WEb
   PIN OEb
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  482.5 28155.0 552.5 28295.0 ;
      END
   END OEb
   PIN clk
      DIRECTION INPUT ;
      PORT
         LAYER metal1 ;
         RECT  3340.0 28155.0 3475.0 28345.0 ;
      END
   END clk
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal1 ;
         RECT  106185.0 35.0 106535.0 115822.5 ;
         LAYER metal1 ;
         RECT  4175.0 35.0 4525.0 115822.5 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal2 ;
         RECT  13657.5 35.0 14007.5 115822.5 ;
      END
   END gnd
   OBS
   LAYER  metal1 ;
      RECT  4317.5 35860.0 4382.5 36065.0 ;
      RECT  8565.0 28610.0 8630.0 28675.0 ;
      RECT  8565.0 28337.5 8630.0 28402.5 ;
      RECT  8495.0 28610.0 8597.5 28675.0 ;
      RECT  8565.0 28370.0 8630.0 28642.5 ;
      RECT  8597.5 28337.5 8700.0 28402.5 ;
      RECT  13292.5 28610.0 13357.5 28675.0 ;
      RECT  13292.5 28122.5 13357.5 28187.5 ;
      RECT  10990.0 28610.0 13325.0 28675.0 ;
      RECT  13292.5 28155.0 13357.5 28642.5 ;
      RECT  13325.0 28122.5 15660.0 28187.5 ;
      RECT  8565.0 30045.0 8630.0 30110.0 ;
      RECT  8565.0 30317.5 8630.0 30382.5 ;
      RECT  8495.0 30045.0 8597.5 30110.0 ;
      RECT  8565.0 30077.5 8630.0 30350.0 ;
      RECT  8597.5 30317.5 8700.0 30382.5 ;
      RECT  13292.5 30045.0 13357.5 30110.0 ;
      RECT  13292.5 30532.5 13357.5 30597.5 ;
      RECT  10990.0 30045.0 13325.0 30110.0 ;
      RECT  13292.5 30077.5 13357.5 30565.0 ;
      RECT  13325.0 30532.5 15660.0 30597.5 ;
      RECT  8565.0 31300.0 8630.0 31365.0 ;
      RECT  8565.0 31027.5 8630.0 31092.5 ;
      RECT  8495.0 31300.0 8597.5 31365.0 ;
      RECT  8565.0 31060.0 8630.0 31332.5 ;
      RECT  8597.5 31027.5 8700.0 31092.5 ;
      RECT  13292.5 31300.0 13357.5 31365.0 ;
      RECT  13292.5 30812.5 13357.5 30877.5 ;
      RECT  10990.0 31300.0 13325.0 31365.0 ;
      RECT  13292.5 30845.0 13357.5 31332.5 ;
      RECT  13325.0 30812.5 15660.0 30877.5 ;
      RECT  8565.0 32735.0 8630.0 32800.0 ;
      RECT  8565.0 33007.5 8630.0 33072.5 ;
      RECT  8495.0 32735.0 8597.5 32800.0 ;
      RECT  8565.0 32767.5 8630.0 33040.0 ;
      RECT  8597.5 33007.5 8700.0 33072.5 ;
      RECT  13292.5 32735.0 13357.5 32800.0 ;
      RECT  13292.5 33222.5 13357.5 33287.5 ;
      RECT  10990.0 32735.0 13325.0 32800.0 ;
      RECT  13292.5 32767.5 13357.5 33255.0 ;
      RECT  13325.0 33222.5 15660.0 33287.5 ;
      RECT  8565.0 33990.0 8630.0 34055.0 ;
      RECT  8565.0 33717.5 8630.0 33782.5 ;
      RECT  8495.0 33990.0 8597.5 34055.0 ;
      RECT  8565.0 33750.0 8630.0 34022.5 ;
      RECT  8597.5 33717.5 8700.0 33782.5 ;
      RECT  13292.5 33990.0 13357.5 34055.0 ;
      RECT  13292.5 33502.5 13357.5 33567.5 ;
      RECT  10990.0 33990.0 13325.0 34055.0 ;
      RECT  13292.5 33535.0 13357.5 34022.5 ;
      RECT  13325.0 33502.5 15660.0 33567.5 ;
      RECT  8565.0 35425.0 8630.0 35490.0 ;
      RECT  8565.0 35697.5 8630.0 35762.5 ;
      RECT  8495.0 35425.0 8597.5 35490.0 ;
      RECT  8565.0 35457.5 8630.0 35730.0 ;
      RECT  8597.5 35697.5 8700.0 35762.5 ;
      RECT  13292.5 35425.0 13357.5 35490.0 ;
      RECT  13292.5 35912.5 13357.5 35977.5 ;
      RECT  10990.0 35425.0 13325.0 35490.0 ;
      RECT  13292.5 35457.5 13357.5 35945.0 ;
      RECT  13325.0 35912.5 15660.0 35977.5 ;
      RECT  8565.0 36680.0 8630.0 36745.0 ;
      RECT  8565.0 36407.5 8630.0 36472.5 ;
      RECT  8495.0 36680.0 8597.5 36745.0 ;
      RECT  8565.0 36440.0 8630.0 36712.5 ;
      RECT  8597.5 36407.5 8700.0 36472.5 ;
      RECT  13292.5 36680.0 13357.5 36745.0 ;
      RECT  13292.5 36192.5 13357.5 36257.5 ;
      RECT  10990.0 36680.0 13325.0 36745.0 ;
      RECT  13292.5 36225.0 13357.5 36712.5 ;
      RECT  13325.0 36192.5 15660.0 36257.5 ;
      RECT  8565.0 38115.0 8630.0 38180.0 ;
      RECT  8565.0 38387.5 8630.0 38452.5 ;
      RECT  8495.0 38115.0 8597.5 38180.0 ;
      RECT  8565.0 38147.5 8630.0 38420.0 ;
      RECT  8597.5 38387.5 8700.0 38452.5 ;
      RECT  13292.5 38115.0 13357.5 38180.0 ;
      RECT  13292.5 38602.5 13357.5 38667.5 ;
      RECT  10990.0 38115.0 13325.0 38180.0 ;
      RECT  13292.5 38147.5 13357.5 38635.0 ;
      RECT  13325.0 38602.5 15660.0 38667.5 ;
      RECT  8565.0 39370.0 8630.0 39435.0 ;
      RECT  8565.0 39097.5 8630.0 39162.5 ;
      RECT  8495.0 39370.0 8597.5 39435.0 ;
      RECT  8565.0 39130.0 8630.0 39402.5 ;
      RECT  8597.5 39097.5 8700.0 39162.5 ;
      RECT  13292.5 39370.0 13357.5 39435.0 ;
      RECT  13292.5 38882.5 13357.5 38947.5 ;
      RECT  10990.0 39370.0 13325.0 39435.0 ;
      RECT  13292.5 38915.0 13357.5 39402.5 ;
      RECT  13325.0 38882.5 15660.0 38947.5 ;
      RECT  8565.0 40805.0 8630.0 40870.0 ;
      RECT  8565.0 41077.5 8630.0 41142.5 ;
      RECT  8495.0 40805.0 8597.5 40870.0 ;
      RECT  8565.0 40837.5 8630.0 41110.0 ;
      RECT  8597.5 41077.5 8700.0 41142.5 ;
      RECT  13292.5 40805.0 13357.5 40870.0 ;
      RECT  13292.5 41292.5 13357.5 41357.5 ;
      RECT  10990.0 40805.0 13325.0 40870.0 ;
      RECT  13292.5 40837.5 13357.5 41325.0 ;
      RECT  13325.0 41292.5 15660.0 41357.5 ;
      RECT  8565.0 42060.0 8630.0 42125.0 ;
      RECT  8565.0 41787.5 8630.0 41852.5 ;
      RECT  8495.0 42060.0 8597.5 42125.0 ;
      RECT  8565.0 41820.0 8630.0 42092.5 ;
      RECT  8597.5 41787.5 8700.0 41852.5 ;
      RECT  13292.5 42060.0 13357.5 42125.0 ;
      RECT  13292.5 41572.5 13357.5 41637.5 ;
      RECT  10990.0 42060.0 13325.0 42125.0 ;
      RECT  13292.5 41605.0 13357.5 42092.5 ;
      RECT  13325.0 41572.5 15660.0 41637.5 ;
      RECT  8565.0 43495.0 8630.0 43560.0 ;
      RECT  8565.0 43767.5 8630.0 43832.5 ;
      RECT  8495.0 43495.0 8597.5 43560.0 ;
      RECT  8565.0 43527.5 8630.0 43800.0 ;
      RECT  8597.5 43767.5 8700.0 43832.5 ;
      RECT  13292.5 43495.0 13357.5 43560.0 ;
      RECT  13292.5 43982.5 13357.5 44047.5 ;
      RECT  10990.0 43495.0 13325.0 43560.0 ;
      RECT  13292.5 43527.5 13357.5 44015.0 ;
      RECT  13325.0 43982.5 15660.0 44047.5 ;
      RECT  8565.0 44750.0 8630.0 44815.0 ;
      RECT  8565.0 44477.5 8630.0 44542.5 ;
      RECT  8495.0 44750.0 8597.5 44815.0 ;
      RECT  8565.0 44510.0 8630.0 44782.5 ;
      RECT  8597.5 44477.5 8700.0 44542.5 ;
      RECT  13292.5 44750.0 13357.5 44815.0 ;
      RECT  13292.5 44262.5 13357.5 44327.5 ;
      RECT  10990.0 44750.0 13325.0 44815.0 ;
      RECT  13292.5 44295.0 13357.5 44782.5 ;
      RECT  13325.0 44262.5 15660.0 44327.5 ;
      RECT  8565.0 46185.0 8630.0 46250.0 ;
      RECT  8565.0 46457.5 8630.0 46522.5 ;
      RECT  8495.0 46185.0 8597.5 46250.0 ;
      RECT  8565.0 46217.5 8630.0 46490.0 ;
      RECT  8597.5 46457.5 8700.0 46522.5 ;
      RECT  13292.5 46185.0 13357.5 46250.0 ;
      RECT  13292.5 46672.5 13357.5 46737.5 ;
      RECT  10990.0 46185.0 13325.0 46250.0 ;
      RECT  13292.5 46217.5 13357.5 46705.0 ;
      RECT  13325.0 46672.5 15660.0 46737.5 ;
      RECT  8565.0 47440.0 8630.0 47505.0 ;
      RECT  8565.0 47167.5 8630.0 47232.5 ;
      RECT  8495.0 47440.0 8597.5 47505.0 ;
      RECT  8565.0 47200.0 8630.0 47472.5 ;
      RECT  8597.5 47167.5 8700.0 47232.5 ;
      RECT  13292.5 47440.0 13357.5 47505.0 ;
      RECT  13292.5 46952.5 13357.5 47017.5 ;
      RECT  10990.0 47440.0 13325.0 47505.0 ;
      RECT  13292.5 46985.0 13357.5 47472.5 ;
      RECT  13325.0 46952.5 15660.0 47017.5 ;
      RECT  8565.0 48875.0 8630.0 48940.0 ;
      RECT  8565.0 49147.5 8630.0 49212.5 ;
      RECT  8495.0 48875.0 8597.5 48940.0 ;
      RECT  8565.0 48907.5 8630.0 49180.0 ;
      RECT  8597.5 49147.5 8700.0 49212.5 ;
      RECT  13292.5 48875.0 13357.5 48940.0 ;
      RECT  13292.5 49362.5 13357.5 49427.5 ;
      RECT  10990.0 48875.0 13325.0 48940.0 ;
      RECT  13292.5 48907.5 13357.5 49395.0 ;
      RECT  13325.0 49362.5 15660.0 49427.5 ;
      RECT  8565.0 50130.0 8630.0 50195.0 ;
      RECT  8565.0 49857.5 8630.0 49922.5 ;
      RECT  8495.0 50130.0 8597.5 50195.0 ;
      RECT  8565.0 49890.0 8630.0 50162.5 ;
      RECT  8597.5 49857.5 8700.0 49922.5 ;
      RECT  13292.5 50130.0 13357.5 50195.0 ;
      RECT  13292.5 49642.5 13357.5 49707.5 ;
      RECT  10990.0 50130.0 13325.0 50195.0 ;
      RECT  13292.5 49675.0 13357.5 50162.5 ;
      RECT  13325.0 49642.5 15660.0 49707.5 ;
      RECT  8565.0 51565.0 8630.0 51630.0 ;
      RECT  8565.0 51837.5 8630.0 51902.5 ;
      RECT  8495.0 51565.0 8597.5 51630.0 ;
      RECT  8565.0 51597.5 8630.0 51870.0 ;
      RECT  8597.5 51837.5 8700.0 51902.5 ;
      RECT  13292.5 51565.0 13357.5 51630.0 ;
      RECT  13292.5 52052.5 13357.5 52117.5 ;
      RECT  10990.0 51565.0 13325.0 51630.0 ;
      RECT  13292.5 51597.5 13357.5 52085.0 ;
      RECT  13325.0 52052.5 15660.0 52117.5 ;
      RECT  8565.0 52820.0 8630.0 52885.0 ;
      RECT  8565.0 52547.5 8630.0 52612.5 ;
      RECT  8495.0 52820.0 8597.5 52885.0 ;
      RECT  8565.0 52580.0 8630.0 52852.5 ;
      RECT  8597.5 52547.5 8700.0 52612.5 ;
      RECT  13292.5 52820.0 13357.5 52885.0 ;
      RECT  13292.5 52332.5 13357.5 52397.5 ;
      RECT  10990.0 52820.0 13325.0 52885.0 ;
      RECT  13292.5 52365.0 13357.5 52852.5 ;
      RECT  13325.0 52332.5 15660.0 52397.5 ;
      RECT  8565.0 54255.0 8630.0 54320.0 ;
      RECT  8565.0 54527.5 8630.0 54592.5 ;
      RECT  8495.0 54255.0 8597.5 54320.0 ;
      RECT  8565.0 54287.5 8630.0 54560.0 ;
      RECT  8597.5 54527.5 8700.0 54592.5 ;
      RECT  13292.5 54255.0 13357.5 54320.0 ;
      RECT  13292.5 54742.5 13357.5 54807.5 ;
      RECT  10990.0 54255.0 13325.0 54320.0 ;
      RECT  13292.5 54287.5 13357.5 54775.0 ;
      RECT  13325.0 54742.5 15660.0 54807.5 ;
      RECT  8565.0 55510.0 8630.0 55575.0 ;
      RECT  8565.0 55237.5 8630.0 55302.5 ;
      RECT  8495.0 55510.0 8597.5 55575.0 ;
      RECT  8565.0 55270.0 8630.0 55542.5 ;
      RECT  8597.5 55237.5 8700.0 55302.5 ;
      RECT  13292.5 55510.0 13357.5 55575.0 ;
      RECT  13292.5 55022.5 13357.5 55087.5 ;
      RECT  10990.0 55510.0 13325.0 55575.0 ;
      RECT  13292.5 55055.0 13357.5 55542.5 ;
      RECT  13325.0 55022.5 15660.0 55087.5 ;
      RECT  8565.0 56945.0 8630.0 57010.0 ;
      RECT  8565.0 57217.5 8630.0 57282.5 ;
      RECT  8495.0 56945.0 8597.5 57010.0 ;
      RECT  8565.0 56977.5 8630.0 57250.0 ;
      RECT  8597.5 57217.5 8700.0 57282.5 ;
      RECT  13292.5 56945.0 13357.5 57010.0 ;
      RECT  13292.5 57432.5 13357.5 57497.5 ;
      RECT  10990.0 56945.0 13325.0 57010.0 ;
      RECT  13292.5 56977.5 13357.5 57465.0 ;
      RECT  13325.0 57432.5 15660.0 57497.5 ;
      RECT  8565.0 58200.0 8630.0 58265.0 ;
      RECT  8565.0 57927.5 8630.0 57992.5 ;
      RECT  8495.0 58200.0 8597.5 58265.0 ;
      RECT  8565.0 57960.0 8630.0 58232.5 ;
      RECT  8597.5 57927.5 8700.0 57992.5 ;
      RECT  13292.5 58200.0 13357.5 58265.0 ;
      RECT  13292.5 57712.5 13357.5 57777.5 ;
      RECT  10990.0 58200.0 13325.0 58265.0 ;
      RECT  13292.5 57745.0 13357.5 58232.5 ;
      RECT  13325.0 57712.5 15660.0 57777.5 ;
      RECT  8565.0 59635.0 8630.0 59700.0 ;
      RECT  8565.0 59907.5 8630.0 59972.5 ;
      RECT  8495.0 59635.0 8597.5 59700.0 ;
      RECT  8565.0 59667.5 8630.0 59940.0 ;
      RECT  8597.5 59907.5 8700.0 59972.5 ;
      RECT  13292.5 59635.0 13357.5 59700.0 ;
      RECT  13292.5 60122.5 13357.5 60187.5 ;
      RECT  10990.0 59635.0 13325.0 59700.0 ;
      RECT  13292.5 59667.5 13357.5 60155.0 ;
      RECT  13325.0 60122.5 15660.0 60187.5 ;
      RECT  8565.0 60890.0 8630.0 60955.0 ;
      RECT  8565.0 60617.5 8630.0 60682.5 ;
      RECT  8495.0 60890.0 8597.5 60955.0 ;
      RECT  8565.0 60650.0 8630.0 60922.5 ;
      RECT  8597.5 60617.5 8700.0 60682.5 ;
      RECT  13292.5 60890.0 13357.5 60955.0 ;
      RECT  13292.5 60402.5 13357.5 60467.5 ;
      RECT  10990.0 60890.0 13325.0 60955.0 ;
      RECT  13292.5 60435.0 13357.5 60922.5 ;
      RECT  13325.0 60402.5 15660.0 60467.5 ;
      RECT  8565.0 62325.0 8630.0 62390.0 ;
      RECT  8565.0 62597.5 8630.0 62662.5 ;
      RECT  8495.0 62325.0 8597.5 62390.0 ;
      RECT  8565.0 62357.5 8630.0 62630.0 ;
      RECT  8597.5 62597.5 8700.0 62662.5 ;
      RECT  13292.5 62325.0 13357.5 62390.0 ;
      RECT  13292.5 62812.5 13357.5 62877.5 ;
      RECT  10990.0 62325.0 13325.0 62390.0 ;
      RECT  13292.5 62357.5 13357.5 62845.0 ;
      RECT  13325.0 62812.5 15660.0 62877.5 ;
      RECT  8565.0 63580.0 8630.0 63645.0 ;
      RECT  8565.0 63307.5 8630.0 63372.5 ;
      RECT  8495.0 63580.0 8597.5 63645.0 ;
      RECT  8565.0 63340.0 8630.0 63612.5 ;
      RECT  8597.5 63307.5 8700.0 63372.5 ;
      RECT  13292.5 63580.0 13357.5 63645.0 ;
      RECT  13292.5 63092.5 13357.5 63157.5 ;
      RECT  10990.0 63580.0 13325.0 63645.0 ;
      RECT  13292.5 63125.0 13357.5 63612.5 ;
      RECT  13325.0 63092.5 15660.0 63157.5 ;
      RECT  8565.0 65015.0 8630.0 65080.0 ;
      RECT  8565.0 65287.5 8630.0 65352.5 ;
      RECT  8495.0 65015.0 8597.5 65080.0 ;
      RECT  8565.0 65047.5 8630.0 65320.0 ;
      RECT  8597.5 65287.5 8700.0 65352.5 ;
      RECT  13292.5 65015.0 13357.5 65080.0 ;
      RECT  13292.5 65502.5 13357.5 65567.5 ;
      RECT  10990.0 65015.0 13325.0 65080.0 ;
      RECT  13292.5 65047.5 13357.5 65535.0 ;
      RECT  13325.0 65502.5 15660.0 65567.5 ;
      RECT  8565.0 66270.0 8630.0 66335.0 ;
      RECT  8565.0 65997.5 8630.0 66062.5 ;
      RECT  8495.0 66270.0 8597.5 66335.0 ;
      RECT  8565.0 66030.0 8630.0 66302.5 ;
      RECT  8597.5 65997.5 8700.0 66062.5 ;
      RECT  13292.5 66270.0 13357.5 66335.0 ;
      RECT  13292.5 65782.5 13357.5 65847.5 ;
      RECT  10990.0 66270.0 13325.0 66335.0 ;
      RECT  13292.5 65815.0 13357.5 66302.5 ;
      RECT  13325.0 65782.5 15660.0 65847.5 ;
      RECT  8565.0 67705.0 8630.0 67770.0 ;
      RECT  8565.0 67977.5 8630.0 68042.5 ;
      RECT  8495.0 67705.0 8597.5 67770.0 ;
      RECT  8565.0 67737.5 8630.0 68010.0 ;
      RECT  8597.5 67977.5 8700.0 68042.5 ;
      RECT  13292.5 67705.0 13357.5 67770.0 ;
      RECT  13292.5 68192.5 13357.5 68257.5 ;
      RECT  10990.0 67705.0 13325.0 67770.0 ;
      RECT  13292.5 67737.5 13357.5 68225.0 ;
      RECT  13325.0 68192.5 15660.0 68257.5 ;
      RECT  8565.0 68960.0 8630.0 69025.0 ;
      RECT  8565.0 68687.5 8630.0 68752.5 ;
      RECT  8495.0 68960.0 8597.5 69025.0 ;
      RECT  8565.0 68720.0 8630.0 68992.5 ;
      RECT  8597.5 68687.5 8700.0 68752.5 ;
      RECT  13292.5 68960.0 13357.5 69025.0 ;
      RECT  13292.5 68472.5 13357.5 68537.5 ;
      RECT  10990.0 68960.0 13325.0 69025.0 ;
      RECT  13292.5 68505.0 13357.5 68992.5 ;
      RECT  13325.0 68472.5 15660.0 68537.5 ;
      RECT  8565.0 70395.0 8630.0 70460.0 ;
      RECT  8565.0 70667.5 8630.0 70732.5 ;
      RECT  8495.0 70395.0 8597.5 70460.0 ;
      RECT  8565.0 70427.5 8630.0 70700.0 ;
      RECT  8597.5 70667.5 8700.0 70732.5 ;
      RECT  13292.5 70395.0 13357.5 70460.0 ;
      RECT  13292.5 70882.5 13357.5 70947.5 ;
      RECT  10990.0 70395.0 13325.0 70460.0 ;
      RECT  13292.5 70427.5 13357.5 70915.0 ;
      RECT  13325.0 70882.5 15660.0 70947.5 ;
      RECT  8565.0 71650.0 8630.0 71715.0 ;
      RECT  8565.0 71377.5 8630.0 71442.5 ;
      RECT  8495.0 71650.0 8597.5 71715.0 ;
      RECT  8565.0 71410.0 8630.0 71682.5 ;
      RECT  8597.5 71377.5 8700.0 71442.5 ;
      RECT  13292.5 71650.0 13357.5 71715.0 ;
      RECT  13292.5 71162.5 13357.5 71227.5 ;
      RECT  10990.0 71650.0 13325.0 71715.0 ;
      RECT  13292.5 71195.0 13357.5 71682.5 ;
      RECT  13325.0 71162.5 15660.0 71227.5 ;
      RECT  8565.0 73085.0 8630.0 73150.0 ;
      RECT  8565.0 73357.5 8630.0 73422.5 ;
      RECT  8495.0 73085.0 8597.5 73150.0 ;
      RECT  8565.0 73117.5 8630.0 73390.0 ;
      RECT  8597.5 73357.5 8700.0 73422.5 ;
      RECT  13292.5 73085.0 13357.5 73150.0 ;
      RECT  13292.5 73572.5 13357.5 73637.5 ;
      RECT  10990.0 73085.0 13325.0 73150.0 ;
      RECT  13292.5 73117.5 13357.5 73605.0 ;
      RECT  13325.0 73572.5 15660.0 73637.5 ;
      RECT  8565.0 74340.0 8630.0 74405.0 ;
      RECT  8565.0 74067.5 8630.0 74132.5 ;
      RECT  8495.0 74340.0 8597.5 74405.0 ;
      RECT  8565.0 74100.0 8630.0 74372.5 ;
      RECT  8597.5 74067.5 8700.0 74132.5 ;
      RECT  13292.5 74340.0 13357.5 74405.0 ;
      RECT  13292.5 73852.5 13357.5 73917.5 ;
      RECT  10990.0 74340.0 13325.0 74405.0 ;
      RECT  13292.5 73885.0 13357.5 74372.5 ;
      RECT  13325.0 73852.5 15660.0 73917.5 ;
      RECT  8565.0 75775.0 8630.0 75840.0 ;
      RECT  8565.0 76047.5 8630.0 76112.5 ;
      RECT  8495.0 75775.0 8597.5 75840.0 ;
      RECT  8565.0 75807.5 8630.0 76080.0 ;
      RECT  8597.5 76047.5 8700.0 76112.5 ;
      RECT  13292.5 75775.0 13357.5 75840.0 ;
      RECT  13292.5 76262.5 13357.5 76327.5 ;
      RECT  10990.0 75775.0 13325.0 75840.0 ;
      RECT  13292.5 75807.5 13357.5 76295.0 ;
      RECT  13325.0 76262.5 15660.0 76327.5 ;
      RECT  8565.0 77030.0 8630.0 77095.0 ;
      RECT  8565.0 76757.5 8630.0 76822.5 ;
      RECT  8495.0 77030.0 8597.5 77095.0 ;
      RECT  8565.0 76790.0 8630.0 77062.5 ;
      RECT  8597.5 76757.5 8700.0 76822.5 ;
      RECT  13292.5 77030.0 13357.5 77095.0 ;
      RECT  13292.5 76542.5 13357.5 76607.5 ;
      RECT  10990.0 77030.0 13325.0 77095.0 ;
      RECT  13292.5 76575.0 13357.5 77062.5 ;
      RECT  13325.0 76542.5 15660.0 76607.5 ;
      RECT  8565.0 78465.0 8630.0 78530.0 ;
      RECT  8565.0 78737.5 8630.0 78802.5 ;
      RECT  8495.0 78465.0 8597.5 78530.0 ;
      RECT  8565.0 78497.5 8630.0 78770.0 ;
      RECT  8597.5 78737.5 8700.0 78802.5 ;
      RECT  13292.5 78465.0 13357.5 78530.0 ;
      RECT  13292.5 78952.5 13357.5 79017.5 ;
      RECT  10990.0 78465.0 13325.0 78530.0 ;
      RECT  13292.5 78497.5 13357.5 78985.0 ;
      RECT  13325.0 78952.5 15660.0 79017.5 ;
      RECT  8565.0 79720.0 8630.0 79785.0 ;
      RECT  8565.0 79447.5 8630.0 79512.5 ;
      RECT  8495.0 79720.0 8597.5 79785.0 ;
      RECT  8565.0 79480.0 8630.0 79752.5 ;
      RECT  8597.5 79447.5 8700.0 79512.5 ;
      RECT  13292.5 79720.0 13357.5 79785.0 ;
      RECT  13292.5 79232.5 13357.5 79297.5 ;
      RECT  10990.0 79720.0 13325.0 79785.0 ;
      RECT  13292.5 79265.0 13357.5 79752.5 ;
      RECT  13325.0 79232.5 15660.0 79297.5 ;
      RECT  8565.0 81155.0 8630.0 81220.0 ;
      RECT  8565.0 81427.5 8630.0 81492.5 ;
      RECT  8495.0 81155.0 8597.5 81220.0 ;
      RECT  8565.0 81187.5 8630.0 81460.0 ;
      RECT  8597.5 81427.5 8700.0 81492.5 ;
      RECT  13292.5 81155.0 13357.5 81220.0 ;
      RECT  13292.5 81642.5 13357.5 81707.5 ;
      RECT  10990.0 81155.0 13325.0 81220.0 ;
      RECT  13292.5 81187.5 13357.5 81675.0 ;
      RECT  13325.0 81642.5 15660.0 81707.5 ;
      RECT  8565.0 82410.0 8630.0 82475.0 ;
      RECT  8565.0 82137.5 8630.0 82202.5 ;
      RECT  8495.0 82410.0 8597.5 82475.0 ;
      RECT  8565.0 82170.0 8630.0 82442.5 ;
      RECT  8597.5 82137.5 8700.0 82202.5 ;
      RECT  13292.5 82410.0 13357.5 82475.0 ;
      RECT  13292.5 81922.5 13357.5 81987.5 ;
      RECT  10990.0 82410.0 13325.0 82475.0 ;
      RECT  13292.5 81955.0 13357.5 82442.5 ;
      RECT  13325.0 81922.5 15660.0 81987.5 ;
      RECT  8565.0 83845.0 8630.0 83910.0 ;
      RECT  8565.0 84117.5 8630.0 84182.5 ;
      RECT  8495.0 83845.0 8597.5 83910.0 ;
      RECT  8565.0 83877.5 8630.0 84150.0 ;
      RECT  8597.5 84117.5 8700.0 84182.5 ;
      RECT  13292.5 83845.0 13357.5 83910.0 ;
      RECT  13292.5 84332.5 13357.5 84397.5 ;
      RECT  10990.0 83845.0 13325.0 83910.0 ;
      RECT  13292.5 83877.5 13357.5 84365.0 ;
      RECT  13325.0 84332.5 15660.0 84397.5 ;
      RECT  8565.0 85100.0 8630.0 85165.0 ;
      RECT  8565.0 84827.5 8630.0 84892.5 ;
      RECT  8495.0 85100.0 8597.5 85165.0 ;
      RECT  8565.0 84860.0 8630.0 85132.5 ;
      RECT  8597.5 84827.5 8700.0 84892.5 ;
      RECT  13292.5 85100.0 13357.5 85165.0 ;
      RECT  13292.5 84612.5 13357.5 84677.5 ;
      RECT  10990.0 85100.0 13325.0 85165.0 ;
      RECT  13292.5 84645.0 13357.5 85132.5 ;
      RECT  13325.0 84612.5 15660.0 84677.5 ;
      RECT  8565.0 86535.0 8630.0 86600.0 ;
      RECT  8565.0 86807.5 8630.0 86872.5 ;
      RECT  8495.0 86535.0 8597.5 86600.0 ;
      RECT  8565.0 86567.5 8630.0 86840.0 ;
      RECT  8597.5 86807.5 8700.0 86872.5 ;
      RECT  13292.5 86535.0 13357.5 86600.0 ;
      RECT  13292.5 87022.5 13357.5 87087.5 ;
      RECT  10990.0 86535.0 13325.0 86600.0 ;
      RECT  13292.5 86567.5 13357.5 87055.0 ;
      RECT  13325.0 87022.5 15660.0 87087.5 ;
      RECT  8565.0 87790.0 8630.0 87855.0 ;
      RECT  8565.0 87517.5 8630.0 87582.5 ;
      RECT  8495.0 87790.0 8597.5 87855.0 ;
      RECT  8565.0 87550.0 8630.0 87822.5 ;
      RECT  8597.5 87517.5 8700.0 87582.5 ;
      RECT  13292.5 87790.0 13357.5 87855.0 ;
      RECT  13292.5 87302.5 13357.5 87367.5 ;
      RECT  10990.0 87790.0 13325.0 87855.0 ;
      RECT  13292.5 87335.0 13357.5 87822.5 ;
      RECT  13325.0 87302.5 15660.0 87367.5 ;
      RECT  8565.0 89225.0 8630.0 89290.0 ;
      RECT  8565.0 89497.5 8630.0 89562.5 ;
      RECT  8495.0 89225.0 8597.5 89290.0 ;
      RECT  8565.0 89257.5 8630.0 89530.0 ;
      RECT  8597.5 89497.5 8700.0 89562.5 ;
      RECT  13292.5 89225.0 13357.5 89290.0 ;
      RECT  13292.5 89712.5 13357.5 89777.5 ;
      RECT  10990.0 89225.0 13325.0 89290.0 ;
      RECT  13292.5 89257.5 13357.5 89745.0 ;
      RECT  13325.0 89712.5 15660.0 89777.5 ;
      RECT  8565.0 90480.0 8630.0 90545.0 ;
      RECT  8565.0 90207.5 8630.0 90272.5 ;
      RECT  8495.0 90480.0 8597.5 90545.0 ;
      RECT  8565.0 90240.0 8630.0 90512.5 ;
      RECT  8597.5 90207.5 8700.0 90272.5 ;
      RECT  13292.5 90480.0 13357.5 90545.0 ;
      RECT  13292.5 89992.5 13357.5 90057.5 ;
      RECT  10990.0 90480.0 13325.0 90545.0 ;
      RECT  13292.5 90025.0 13357.5 90512.5 ;
      RECT  13325.0 89992.5 15660.0 90057.5 ;
      RECT  8565.0 91915.0 8630.0 91980.0 ;
      RECT  8565.0 92187.5 8630.0 92252.5 ;
      RECT  8495.0 91915.0 8597.5 91980.0 ;
      RECT  8565.0 91947.5 8630.0 92220.0 ;
      RECT  8597.5 92187.5 8700.0 92252.5 ;
      RECT  13292.5 91915.0 13357.5 91980.0 ;
      RECT  13292.5 92402.5 13357.5 92467.5 ;
      RECT  10990.0 91915.0 13325.0 91980.0 ;
      RECT  13292.5 91947.5 13357.5 92435.0 ;
      RECT  13325.0 92402.5 15660.0 92467.5 ;
      RECT  8565.0 93170.0 8630.0 93235.0 ;
      RECT  8565.0 92897.5 8630.0 92962.5 ;
      RECT  8495.0 93170.0 8597.5 93235.0 ;
      RECT  8565.0 92930.0 8630.0 93202.5 ;
      RECT  8597.5 92897.5 8700.0 92962.5 ;
      RECT  13292.5 93170.0 13357.5 93235.0 ;
      RECT  13292.5 92682.5 13357.5 92747.5 ;
      RECT  10990.0 93170.0 13325.0 93235.0 ;
      RECT  13292.5 92715.0 13357.5 93202.5 ;
      RECT  13325.0 92682.5 15660.0 92747.5 ;
      RECT  8565.0 94605.0 8630.0 94670.0 ;
      RECT  8565.0 94877.5 8630.0 94942.5 ;
      RECT  8495.0 94605.0 8597.5 94670.0 ;
      RECT  8565.0 94637.5 8630.0 94910.0 ;
      RECT  8597.5 94877.5 8700.0 94942.5 ;
      RECT  13292.5 94605.0 13357.5 94670.0 ;
      RECT  13292.5 95092.5 13357.5 95157.5 ;
      RECT  10990.0 94605.0 13325.0 94670.0 ;
      RECT  13292.5 94637.5 13357.5 95125.0 ;
      RECT  13325.0 95092.5 15660.0 95157.5 ;
      RECT  8565.0 95860.0 8630.0 95925.0 ;
      RECT  8565.0 95587.5 8630.0 95652.5 ;
      RECT  8495.0 95860.0 8597.5 95925.0 ;
      RECT  8565.0 95620.0 8630.0 95892.5 ;
      RECT  8597.5 95587.5 8700.0 95652.5 ;
      RECT  13292.5 95860.0 13357.5 95925.0 ;
      RECT  13292.5 95372.5 13357.5 95437.5 ;
      RECT  10990.0 95860.0 13325.0 95925.0 ;
      RECT  13292.5 95405.0 13357.5 95892.5 ;
      RECT  13325.0 95372.5 15660.0 95437.5 ;
      RECT  8565.0 97295.0 8630.0 97360.0 ;
      RECT  8565.0 97567.5 8630.0 97632.5 ;
      RECT  8495.0 97295.0 8597.5 97360.0 ;
      RECT  8565.0 97327.5 8630.0 97600.0 ;
      RECT  8597.5 97567.5 8700.0 97632.5 ;
      RECT  13292.5 97295.0 13357.5 97360.0 ;
      RECT  13292.5 97782.5 13357.5 97847.5 ;
      RECT  10990.0 97295.0 13325.0 97360.0 ;
      RECT  13292.5 97327.5 13357.5 97815.0 ;
      RECT  13325.0 97782.5 15660.0 97847.5 ;
      RECT  8565.0 98550.0 8630.0 98615.0 ;
      RECT  8565.0 98277.5 8630.0 98342.5 ;
      RECT  8495.0 98550.0 8597.5 98615.0 ;
      RECT  8565.0 98310.0 8630.0 98582.5 ;
      RECT  8597.5 98277.5 8700.0 98342.5 ;
      RECT  13292.5 98550.0 13357.5 98615.0 ;
      RECT  13292.5 98062.5 13357.5 98127.5 ;
      RECT  10990.0 98550.0 13325.0 98615.0 ;
      RECT  13292.5 98095.0 13357.5 98582.5 ;
      RECT  13325.0 98062.5 15660.0 98127.5 ;
      RECT  8565.0 99985.0 8630.0 100050.0 ;
      RECT  8565.0 100257.5 8630.0 100322.5 ;
      RECT  8495.0 99985.0 8597.5 100050.0 ;
      RECT  8565.0 100017.5 8630.0 100290.0 ;
      RECT  8597.5 100257.5 8700.0 100322.5 ;
      RECT  13292.5 99985.0 13357.5 100050.0 ;
      RECT  13292.5 100472.5 13357.5 100537.5 ;
      RECT  10990.0 99985.0 13325.0 100050.0 ;
      RECT  13292.5 100017.5 13357.5 100505.0 ;
      RECT  13325.0 100472.5 15660.0 100537.5 ;
      RECT  8565.0 101240.0 8630.0 101305.0 ;
      RECT  8565.0 100967.5 8630.0 101032.5 ;
      RECT  8495.0 101240.0 8597.5 101305.0 ;
      RECT  8565.0 101000.0 8630.0 101272.5 ;
      RECT  8597.5 100967.5 8700.0 101032.5 ;
      RECT  13292.5 101240.0 13357.5 101305.0 ;
      RECT  13292.5 100752.5 13357.5 100817.5 ;
      RECT  10990.0 101240.0 13325.0 101305.0 ;
      RECT  13292.5 100785.0 13357.5 101272.5 ;
      RECT  13325.0 100752.5 15660.0 100817.5 ;
      RECT  8565.0 102675.0 8630.0 102740.0 ;
      RECT  8565.0 102947.5 8630.0 103012.5 ;
      RECT  8495.0 102675.0 8597.5 102740.0 ;
      RECT  8565.0 102707.5 8630.0 102980.0 ;
      RECT  8597.5 102947.5 8700.0 103012.5 ;
      RECT  13292.5 102675.0 13357.5 102740.0 ;
      RECT  13292.5 103162.5 13357.5 103227.5 ;
      RECT  10990.0 102675.0 13325.0 102740.0 ;
      RECT  13292.5 102707.5 13357.5 103195.0 ;
      RECT  13325.0 103162.5 15660.0 103227.5 ;
      RECT  8565.0 103930.0 8630.0 103995.0 ;
      RECT  8565.0 103657.5 8630.0 103722.5 ;
      RECT  8495.0 103930.0 8597.5 103995.0 ;
      RECT  8565.0 103690.0 8630.0 103962.5 ;
      RECT  8597.5 103657.5 8700.0 103722.5 ;
      RECT  13292.5 103930.0 13357.5 103995.0 ;
      RECT  13292.5 103442.5 13357.5 103507.5 ;
      RECT  10990.0 103930.0 13325.0 103995.0 ;
      RECT  13292.5 103475.0 13357.5 103962.5 ;
      RECT  13325.0 103442.5 15660.0 103507.5 ;
      RECT  8565.0 105365.0 8630.0 105430.0 ;
      RECT  8565.0 105637.5 8630.0 105702.5 ;
      RECT  8495.0 105365.0 8597.5 105430.0 ;
      RECT  8565.0 105397.5 8630.0 105670.0 ;
      RECT  8597.5 105637.5 8700.0 105702.5 ;
      RECT  13292.5 105365.0 13357.5 105430.0 ;
      RECT  13292.5 105852.5 13357.5 105917.5 ;
      RECT  10990.0 105365.0 13325.0 105430.0 ;
      RECT  13292.5 105397.5 13357.5 105885.0 ;
      RECT  13325.0 105852.5 15660.0 105917.5 ;
      RECT  8565.0 106620.0 8630.0 106685.0 ;
      RECT  8565.0 106347.5 8630.0 106412.5 ;
      RECT  8495.0 106620.0 8597.5 106685.0 ;
      RECT  8565.0 106380.0 8630.0 106652.5 ;
      RECT  8597.5 106347.5 8700.0 106412.5 ;
      RECT  13292.5 106620.0 13357.5 106685.0 ;
      RECT  13292.5 106132.5 13357.5 106197.5 ;
      RECT  10990.0 106620.0 13325.0 106685.0 ;
      RECT  13292.5 106165.0 13357.5 106652.5 ;
      RECT  13325.0 106132.5 15660.0 106197.5 ;
      RECT  8565.0 108055.0 8630.0 108120.0 ;
      RECT  8565.0 108327.5 8630.0 108392.5 ;
      RECT  8495.0 108055.0 8597.5 108120.0 ;
      RECT  8565.0 108087.5 8630.0 108360.0 ;
      RECT  8597.5 108327.5 8700.0 108392.5 ;
      RECT  13292.5 108055.0 13357.5 108120.0 ;
      RECT  13292.5 108542.5 13357.5 108607.5 ;
      RECT  10990.0 108055.0 13325.0 108120.0 ;
      RECT  13292.5 108087.5 13357.5 108575.0 ;
      RECT  13325.0 108542.5 15660.0 108607.5 ;
      RECT  8565.0 109310.0 8630.0 109375.0 ;
      RECT  8565.0 109037.5 8630.0 109102.5 ;
      RECT  8495.0 109310.0 8597.5 109375.0 ;
      RECT  8565.0 109070.0 8630.0 109342.5 ;
      RECT  8597.5 109037.5 8700.0 109102.5 ;
      RECT  13292.5 109310.0 13357.5 109375.0 ;
      RECT  13292.5 108822.5 13357.5 108887.5 ;
      RECT  10990.0 109310.0 13325.0 109375.0 ;
      RECT  13292.5 108855.0 13357.5 109342.5 ;
      RECT  13325.0 108822.5 15660.0 108887.5 ;
      RECT  8565.0 110745.0 8630.0 110810.0 ;
      RECT  8565.0 111017.5 8630.0 111082.5 ;
      RECT  8495.0 110745.0 8597.5 110810.0 ;
      RECT  8565.0 110777.5 8630.0 111050.0 ;
      RECT  8597.5 111017.5 8700.0 111082.5 ;
      RECT  13292.5 110745.0 13357.5 110810.0 ;
      RECT  13292.5 111232.5 13357.5 111297.5 ;
      RECT  10990.0 110745.0 13325.0 110810.0 ;
      RECT  13292.5 110777.5 13357.5 111265.0 ;
      RECT  13325.0 111232.5 15660.0 111297.5 ;
      RECT  8565.0 112000.0 8630.0 112065.0 ;
      RECT  8565.0 111727.5 8630.0 111792.5 ;
      RECT  8495.0 112000.0 8597.5 112065.0 ;
      RECT  8565.0 111760.0 8630.0 112032.5 ;
      RECT  8597.5 111727.5 8700.0 111792.5 ;
      RECT  13292.5 112000.0 13357.5 112065.0 ;
      RECT  13292.5 111512.5 13357.5 111577.5 ;
      RECT  10990.0 112000.0 13325.0 112065.0 ;
      RECT  13292.5 111545.0 13357.5 112032.5 ;
      RECT  13325.0 111512.5 15660.0 111577.5 ;
      RECT  8565.0 113435.0 8630.0 113500.0 ;
      RECT  8565.0 113707.5 8630.0 113772.5 ;
      RECT  8495.0 113435.0 8597.5 113500.0 ;
      RECT  8565.0 113467.5 8630.0 113740.0 ;
      RECT  8597.5 113707.5 8700.0 113772.5 ;
      RECT  13292.5 113435.0 13357.5 113500.0 ;
      RECT  13292.5 113922.5 13357.5 113987.5 ;
      RECT  10990.0 113435.0 13325.0 113500.0 ;
      RECT  13292.5 113467.5 13357.5 113955.0 ;
      RECT  13325.0 113922.5 15660.0 113987.5 ;
      RECT  9155.0 27982.5 15750.0 28047.5 ;
      RECT  9155.0 30672.5 15750.0 30737.5 ;
      RECT  9155.0 33362.5 15750.0 33427.5 ;
      RECT  9155.0 36052.5 15750.0 36117.5 ;
      RECT  9155.0 38742.5 15750.0 38807.5 ;
      RECT  9155.0 41432.5 15750.0 41497.5 ;
      RECT  9155.0 44122.5 15750.0 44187.5 ;
      RECT  9155.0 46812.5 15750.0 46877.5 ;
      RECT  9155.0 49502.5 15750.0 49567.5 ;
      RECT  9155.0 52192.5 15750.0 52257.5 ;
      RECT  9155.0 54882.5 15750.0 54947.5 ;
      RECT  9155.0 57572.5 15750.0 57637.5 ;
      RECT  9155.0 60262.5 15750.0 60327.5 ;
      RECT  9155.0 62952.5 15750.0 63017.5 ;
      RECT  9155.0 65642.5 15750.0 65707.5 ;
      RECT  9155.0 68332.5 15750.0 68397.5 ;
      RECT  9155.0 71022.5 15750.0 71087.5 ;
      RECT  9155.0 73712.5 15750.0 73777.5 ;
      RECT  9155.0 76402.5 15750.0 76467.5 ;
      RECT  9155.0 79092.5 15750.0 79157.5 ;
      RECT  9155.0 81782.5 15750.0 81847.5 ;
      RECT  9155.0 84472.5 15750.0 84537.5 ;
      RECT  9155.0 87162.5 15750.0 87227.5 ;
      RECT  9155.0 89852.5 15750.0 89917.5 ;
      RECT  9155.0 92542.5 15750.0 92607.5 ;
      RECT  9155.0 95232.5 15750.0 95297.5 ;
      RECT  9155.0 97922.5 15750.0 97987.5 ;
      RECT  9155.0 100612.5 15750.0 100677.5 ;
      RECT  9155.0 103302.5 15750.0 103367.5 ;
      RECT  9155.0 105992.5 15750.0 106057.5 ;
      RECT  9155.0 108682.5 15750.0 108747.5 ;
      RECT  9155.0 111372.5 15750.0 111437.5 ;
      RECT  9155.0 114062.5 15750.0 114127.5 ;
      RECT  4175.0 29327.5 106535.0 29392.5 ;
      RECT  4175.0 32017.5 106535.0 32082.5 ;
      RECT  4175.0 34707.5 106535.0 34772.5 ;
      RECT  4175.0 37397.5 106535.0 37462.5 ;
      RECT  4175.0 40087.5 106535.0 40152.5 ;
      RECT  4175.0 42777.5 106535.0 42842.5 ;
      RECT  4175.0 45467.5 106535.0 45532.5 ;
      RECT  4175.0 48157.5 106535.0 48222.5 ;
      RECT  4175.0 50847.5 106535.0 50912.5 ;
      RECT  4175.0 53537.5 106535.0 53602.5 ;
      RECT  4175.0 56227.5 106535.0 56292.5 ;
      RECT  4175.0 58917.5 106535.0 58982.5 ;
      RECT  4175.0 61607.5 106535.0 61672.5 ;
      RECT  4175.0 64297.5 106535.0 64362.5 ;
      RECT  4175.0 66987.5 106535.0 67052.5 ;
      RECT  4175.0 69677.5 106535.0 69742.5 ;
      RECT  4175.0 72367.5 106535.0 72432.5 ;
      RECT  4175.0 75057.5 106535.0 75122.5 ;
      RECT  4175.0 77747.5 106535.0 77812.5 ;
      RECT  4175.0 80437.5 106535.0 80502.5 ;
      RECT  4175.0 83127.5 106535.0 83192.5 ;
      RECT  4175.0 85817.5 106535.0 85882.5 ;
      RECT  4175.0 88507.5 106535.0 88572.5 ;
      RECT  4175.0 91197.5 106535.0 91262.5 ;
      RECT  4175.0 93887.5 106535.0 93952.5 ;
      RECT  4175.0 96577.5 106535.0 96642.5 ;
      RECT  4175.0 99267.5 106535.0 99332.5 ;
      RECT  4175.0 101957.5 106535.0 102022.5 ;
      RECT  4175.0 104647.5 106535.0 104712.5 ;
      RECT  4175.0 107337.5 106535.0 107402.5 ;
      RECT  4175.0 110027.5 106535.0 110092.5 ;
      RECT  4175.0 112717.5 106535.0 112782.5 ;
      RECT  11095.0 12047.5 11437.5 12112.5 ;
      RECT  10820.0 13392.5 11642.5 13457.5 ;
      RECT  11095.0 17427.5 11847.5 17492.5 ;
      RECT  10820.0 18772.5 12052.5 18837.5 ;
      RECT  11095.0 22807.5 12257.5 22872.5 ;
      RECT  10820.0 24152.5 12462.5 24217.5 ;
      RECT  11095.0 11842.5 11232.5 11907.5 ;
      RECT  11095.0 14532.5 11232.5 14597.5 ;
      RECT  11095.0 17222.5 11232.5 17287.5 ;
      RECT  11095.0 19912.5 11232.5 19977.5 ;
      RECT  11095.0 22602.5 11232.5 22667.5 ;
      RECT  11095.0 25292.5 11232.5 25357.5 ;
      RECT  4175.0 13187.5 11095.0 13252.5 ;
      RECT  4175.0 15877.5 11095.0 15942.5 ;
      RECT  4175.0 18567.5 11095.0 18632.5 ;
      RECT  4175.0 21257.5 11095.0 21322.5 ;
      RECT  4175.0 23947.5 11095.0 24012.5 ;
      RECT  4175.0 26637.5 11095.0 26702.5 ;
      RECT  12667.5 26012.5 15750.0 26077.5 ;
      RECT  12872.5 25872.5 15750.0 25937.5 ;
      RECT  13077.5 25732.5 15750.0 25797.5 ;
      RECT  13282.5 25592.5 15750.0 25657.5 ;
      RECT  10685.0 630.0 12667.5 695.0 ;
      RECT  10685.0 2065.0 12872.5 2130.0 ;
      RECT  10685.0 3320.0 13077.5 3385.0 ;
      RECT  10685.0 4755.0 13282.5 4820.0 ;
      RECT  10685.0 2.5 13657.5 67.5 ;
      RECT  10685.0 2692.5 13657.5 2757.5 ;
      RECT  10685.0 5382.5 13657.5 5447.5 ;
      RECT  4175.0 1347.5 13657.5 1412.5 ;
      RECT  4175.0 4037.5 13657.5 4102.5 ;
      RECT  11095.0 11080.0 11437.5 11145.0 ;
      RECT  11095.0 10375.0 11642.5 10440.0 ;
      RECT  11095.0 9670.0 11847.5 9735.0 ;
      RECT  11095.0 8965.0 12052.5 9030.0 ;
      RECT  11095.0 8260.0 12257.5 8325.0 ;
      RECT  11095.0 7555.0 12462.5 7620.0 ;
      RECT  11095.0 11432.5 13792.5 11497.5 ;
      RECT  11095.0 10727.5 13792.5 10792.5 ;
      RECT  11095.0 10022.5 13792.5 10087.5 ;
      RECT  11095.0 9317.5 13792.5 9382.5 ;
      RECT  11095.0 8612.5 13792.5 8677.5 ;
      RECT  11095.0 7907.5 13792.5 7972.5 ;
      RECT  11095.0 7202.5 13792.5 7267.5 ;
      RECT  11095.0 6497.5 13792.5 6562.5 ;
      RECT  11095.0 5792.5 13792.5 5857.5 ;
      RECT  7865.0 5587.5 7930.0 5652.5 ;
      RECT  7865.0 5620.0 7930.0 5825.0 ;
      RECT  4175.0 5587.5 7897.5 5652.5 ;
      RECT  10825.0 5587.5 10890.0 5652.5 ;
      RECT  10825.0 5620.0 10890.0 5825.0 ;
      RECT  4175.0 5587.5 10857.5 5652.5 ;
      RECT  5875.0 5587.5 5940.0 5652.5 ;
      RECT  5875.0 5620.0 5940.0 5825.0 ;
      RECT  4175.0 5587.5 5907.5 5652.5 ;
      RECT  8835.0 5587.5 8900.0 5652.5 ;
      RECT  8835.0 5620.0 8900.0 5825.0 ;
      RECT  4175.0 5587.5 8867.5 5652.5 ;
      RECT  14862.5 9875.0 15750.0 9940.0 ;
      RECT  14452.5 7690.0 15750.0 7755.0 ;
      RECT  14657.5 9237.5 15750.0 9302.5 ;
      RECT  14862.5 115072.5 15750.0 115137.5 ;
      RECT  15067.5 16377.5 15750.0 16442.5 ;
      RECT  15272.5 20402.5 15750.0 20467.5 ;
      RECT  4860.0 11637.5 4925.0 11702.5 ;
      RECT  4860.0 11465.0 4925.0 11670.0 ;
      RECT  4892.5 11637.5 14247.5 11702.5 ;
      RECT  8930.0 114267.5 14312.5 114332.5 ;
      RECT  15750.0 115757.5 106185.0 115822.5 ;
      RECT  15750.0 24975.0 106185.0 25040.0 ;
      RECT  15750.0 16507.5 106185.0 16572.5 ;
      RECT  15750.0 12880.0 106185.0 12945.0 ;
      RECT  15750.0 15840.0 106185.0 15905.0 ;
      RECT  15750.0 10890.0 106185.0 10955.0 ;
      RECT  15750.0 13850.0 106185.0 13915.0 ;
      RECT  15750.0 7820.0 106185.0 7885.0 ;
      RECT  14007.5 9107.5 15750.0 9172.5 ;
      RECT  14007.5 20532.5 15750.0 20597.5 ;
      RECT  14007.5 10035.0 15750.0 10100.0 ;
      RECT  14007.5 17310.0 15750.0 17375.0 ;
      RECT  15750.0 28015.0 16455.0 29360.0 ;
      RECT  15750.0 30705.0 16455.0 29360.0 ;
      RECT  15750.0 30705.0 16455.0 32050.0 ;
      RECT  15750.0 33395.0 16455.0 32050.0 ;
      RECT  15750.0 33395.0 16455.0 34740.0 ;
      RECT  15750.0 36085.0 16455.0 34740.0 ;
      RECT  15750.0 36085.0 16455.0 37430.0 ;
      RECT  15750.0 38775.0 16455.0 37430.0 ;
      RECT  15750.0 38775.0 16455.0 40120.0 ;
      RECT  15750.0 41465.0 16455.0 40120.0 ;
      RECT  15750.0 41465.0 16455.0 42810.0 ;
      RECT  15750.0 44155.0 16455.0 42810.0 ;
      RECT  15750.0 44155.0 16455.0 45500.0 ;
      RECT  15750.0 46845.0 16455.0 45500.0 ;
      RECT  15750.0 46845.0 16455.0 48190.0 ;
      RECT  15750.0 49535.0 16455.0 48190.0 ;
      RECT  15750.0 49535.0 16455.0 50880.0 ;
      RECT  15750.0 52225.0 16455.0 50880.0 ;
      RECT  15750.0 52225.0 16455.0 53570.0 ;
      RECT  15750.0 54915.0 16455.0 53570.0 ;
      RECT  15750.0 54915.0 16455.0 56260.0 ;
      RECT  15750.0 57605.0 16455.0 56260.0 ;
      RECT  15750.0 57605.0 16455.0 58950.0 ;
      RECT  15750.0 60295.0 16455.0 58950.0 ;
      RECT  15750.0 60295.0 16455.0 61640.0 ;
      RECT  15750.0 62985.0 16455.0 61640.0 ;
      RECT  15750.0 62985.0 16455.0 64330.0 ;
      RECT  15750.0 65675.0 16455.0 64330.0 ;
      RECT  15750.0 65675.0 16455.0 67020.0 ;
      RECT  15750.0 68365.0 16455.0 67020.0 ;
      RECT  15750.0 68365.0 16455.0 69710.0 ;
      RECT  15750.0 71055.0 16455.0 69710.0 ;
      RECT  15750.0 71055.0 16455.0 72400.0 ;
      RECT  15750.0 73745.0 16455.0 72400.0 ;
      RECT  15750.0 73745.0 16455.0 75090.0 ;
      RECT  15750.0 76435.0 16455.0 75090.0 ;
      RECT  15750.0 76435.0 16455.0 77780.0 ;
      RECT  15750.0 79125.0 16455.0 77780.0 ;
      RECT  15750.0 79125.0 16455.0 80470.0 ;
      RECT  15750.0 81815.0 16455.0 80470.0 ;
      RECT  15750.0 81815.0 16455.0 83160.0 ;
      RECT  15750.0 84505.0 16455.0 83160.0 ;
      RECT  15750.0 84505.0 16455.0 85850.0 ;
      RECT  15750.0 87195.0 16455.0 85850.0 ;
      RECT  15750.0 87195.0 16455.0 88540.0 ;
      RECT  15750.0 89885.0 16455.0 88540.0 ;
      RECT  15750.0 89885.0 16455.0 91230.0 ;
      RECT  15750.0 92575.0 16455.0 91230.0 ;
      RECT  15750.0 92575.0 16455.0 93920.0 ;
      RECT  15750.0 95265.0 16455.0 93920.0 ;
      RECT  15750.0 95265.0 16455.0 96610.0 ;
      RECT  15750.0 97955.0 16455.0 96610.0 ;
      RECT  15750.0 97955.0 16455.0 99300.0 ;
      RECT  15750.0 100645.0 16455.0 99300.0 ;
      RECT  15750.0 100645.0 16455.0 101990.0 ;
      RECT  15750.0 103335.0 16455.0 101990.0 ;
      RECT  15750.0 103335.0 16455.0 104680.0 ;
      RECT  15750.0 106025.0 16455.0 104680.0 ;
      RECT  15750.0 106025.0 16455.0 107370.0 ;
      RECT  15750.0 108715.0 16455.0 107370.0 ;
      RECT  15750.0 108715.0 16455.0 110060.0 ;
      RECT  15750.0 111405.0 16455.0 110060.0 ;
      RECT  15750.0 111405.0 16455.0 112750.0 ;
      RECT  15750.0 114095.0 16455.0 112750.0 ;
      RECT  16455.0 28015.0 17160.0 29360.0 ;
      RECT  16455.0 30705.0 17160.0 29360.0 ;
      RECT  16455.0 30705.0 17160.0 32050.0 ;
      RECT  16455.0 33395.0 17160.0 32050.0 ;
      RECT  16455.0 33395.0 17160.0 34740.0 ;
      RECT  16455.0 36085.0 17160.0 34740.0 ;
      RECT  16455.0 36085.0 17160.0 37430.0 ;
      RECT  16455.0 38775.0 17160.0 37430.0 ;
      RECT  16455.0 38775.0 17160.0 40120.0 ;
      RECT  16455.0 41465.0 17160.0 40120.0 ;
      RECT  16455.0 41465.0 17160.0 42810.0 ;
      RECT  16455.0 44155.0 17160.0 42810.0 ;
      RECT  16455.0 44155.0 17160.0 45500.0 ;
      RECT  16455.0 46845.0 17160.0 45500.0 ;
      RECT  16455.0 46845.0 17160.0 48190.0 ;
      RECT  16455.0 49535.0 17160.0 48190.0 ;
      RECT  16455.0 49535.0 17160.0 50880.0 ;
      RECT  16455.0 52225.0 17160.0 50880.0 ;
      RECT  16455.0 52225.0 17160.0 53570.0 ;
      RECT  16455.0 54915.0 17160.0 53570.0 ;
      RECT  16455.0 54915.0 17160.0 56260.0 ;
      RECT  16455.0 57605.0 17160.0 56260.0 ;
      RECT  16455.0 57605.0 17160.0 58950.0 ;
      RECT  16455.0 60295.0 17160.0 58950.0 ;
      RECT  16455.0 60295.0 17160.0 61640.0 ;
      RECT  16455.0 62985.0 17160.0 61640.0 ;
      RECT  16455.0 62985.0 17160.0 64330.0 ;
      RECT  16455.0 65675.0 17160.0 64330.0 ;
      RECT  16455.0 65675.0 17160.0 67020.0 ;
      RECT  16455.0 68365.0 17160.0 67020.0 ;
      RECT  16455.0 68365.0 17160.0 69710.0 ;
      RECT  16455.0 71055.0 17160.0 69710.0 ;
      RECT  16455.0 71055.0 17160.0 72400.0 ;
      RECT  16455.0 73745.0 17160.0 72400.0 ;
      RECT  16455.0 73745.0 17160.0 75090.0 ;
      RECT  16455.0 76435.0 17160.0 75090.0 ;
      RECT  16455.0 76435.0 17160.0 77780.0 ;
      RECT  16455.0 79125.0 17160.0 77780.0 ;
      RECT  16455.0 79125.0 17160.0 80470.0 ;
      RECT  16455.0 81815.0 17160.0 80470.0 ;
      RECT  16455.0 81815.0 17160.0 83160.0 ;
      RECT  16455.0 84505.0 17160.0 83160.0 ;
      RECT  16455.0 84505.0 17160.0 85850.0 ;
      RECT  16455.0 87195.0 17160.0 85850.0 ;
      RECT  16455.0 87195.0 17160.0 88540.0 ;
      RECT  16455.0 89885.0 17160.0 88540.0 ;
      RECT  16455.0 89885.0 17160.0 91230.0 ;
      RECT  16455.0 92575.0 17160.0 91230.0 ;
      RECT  16455.0 92575.0 17160.0 93920.0 ;
      RECT  16455.0 95265.0 17160.0 93920.0 ;
      RECT  16455.0 95265.0 17160.0 96610.0 ;
      RECT  16455.0 97955.0 17160.0 96610.0 ;
      RECT  16455.0 97955.0 17160.0 99300.0 ;
      RECT  16455.0 100645.0 17160.0 99300.0 ;
      RECT  16455.0 100645.0 17160.0 101990.0 ;
      RECT  16455.0 103335.0 17160.0 101990.0 ;
      RECT  16455.0 103335.0 17160.0 104680.0 ;
      RECT  16455.0 106025.0 17160.0 104680.0 ;
      RECT  16455.0 106025.0 17160.0 107370.0 ;
      RECT  16455.0 108715.0 17160.0 107370.0 ;
      RECT  16455.0 108715.0 17160.0 110060.0 ;
      RECT  16455.0 111405.0 17160.0 110060.0 ;
      RECT  16455.0 111405.0 17160.0 112750.0 ;
      RECT  16455.0 114095.0 17160.0 112750.0 ;
      RECT  17160.0 28015.0 17865.0 29360.0 ;
      RECT  17160.0 30705.0 17865.0 29360.0 ;
      RECT  17160.0 30705.0 17865.0 32050.0 ;
      RECT  17160.0 33395.0 17865.0 32050.0 ;
      RECT  17160.0 33395.0 17865.0 34740.0 ;
      RECT  17160.0 36085.0 17865.0 34740.0 ;
      RECT  17160.0 36085.0 17865.0 37430.0 ;
      RECT  17160.0 38775.0 17865.0 37430.0 ;
      RECT  17160.0 38775.0 17865.0 40120.0 ;
      RECT  17160.0 41465.0 17865.0 40120.0 ;
      RECT  17160.0 41465.0 17865.0 42810.0 ;
      RECT  17160.0 44155.0 17865.0 42810.0 ;
      RECT  17160.0 44155.0 17865.0 45500.0 ;
      RECT  17160.0 46845.0 17865.0 45500.0 ;
      RECT  17160.0 46845.0 17865.0 48190.0 ;
      RECT  17160.0 49535.0 17865.0 48190.0 ;
      RECT  17160.0 49535.0 17865.0 50880.0 ;
      RECT  17160.0 52225.0 17865.0 50880.0 ;
      RECT  17160.0 52225.0 17865.0 53570.0 ;
      RECT  17160.0 54915.0 17865.0 53570.0 ;
      RECT  17160.0 54915.0 17865.0 56260.0 ;
      RECT  17160.0 57605.0 17865.0 56260.0 ;
      RECT  17160.0 57605.0 17865.0 58950.0 ;
      RECT  17160.0 60295.0 17865.0 58950.0 ;
      RECT  17160.0 60295.0 17865.0 61640.0 ;
      RECT  17160.0 62985.0 17865.0 61640.0 ;
      RECT  17160.0 62985.0 17865.0 64330.0 ;
      RECT  17160.0 65675.0 17865.0 64330.0 ;
      RECT  17160.0 65675.0 17865.0 67020.0 ;
      RECT  17160.0 68365.0 17865.0 67020.0 ;
      RECT  17160.0 68365.0 17865.0 69710.0 ;
      RECT  17160.0 71055.0 17865.0 69710.0 ;
      RECT  17160.0 71055.0 17865.0 72400.0 ;
      RECT  17160.0 73745.0 17865.0 72400.0 ;
      RECT  17160.0 73745.0 17865.0 75090.0 ;
      RECT  17160.0 76435.0 17865.0 75090.0 ;
      RECT  17160.0 76435.0 17865.0 77780.0 ;
      RECT  17160.0 79125.0 17865.0 77780.0 ;
      RECT  17160.0 79125.0 17865.0 80470.0 ;
      RECT  17160.0 81815.0 17865.0 80470.0 ;
      RECT  17160.0 81815.0 17865.0 83160.0 ;
      RECT  17160.0 84505.0 17865.0 83160.0 ;
      RECT  17160.0 84505.0 17865.0 85850.0 ;
      RECT  17160.0 87195.0 17865.0 85850.0 ;
      RECT  17160.0 87195.0 17865.0 88540.0 ;
      RECT  17160.0 89885.0 17865.0 88540.0 ;
      RECT  17160.0 89885.0 17865.0 91230.0 ;
      RECT  17160.0 92575.0 17865.0 91230.0 ;
      RECT  17160.0 92575.0 17865.0 93920.0 ;
      RECT  17160.0 95265.0 17865.0 93920.0 ;
      RECT  17160.0 95265.0 17865.0 96610.0 ;
      RECT  17160.0 97955.0 17865.0 96610.0 ;
      RECT  17160.0 97955.0 17865.0 99300.0 ;
      RECT  17160.0 100645.0 17865.0 99300.0 ;
      RECT  17160.0 100645.0 17865.0 101990.0 ;
      RECT  17160.0 103335.0 17865.0 101990.0 ;
      RECT  17160.0 103335.0 17865.0 104680.0 ;
      RECT  17160.0 106025.0 17865.0 104680.0 ;
      RECT  17160.0 106025.0 17865.0 107370.0 ;
      RECT  17160.0 108715.0 17865.0 107370.0 ;
      RECT  17160.0 108715.0 17865.0 110060.0 ;
      RECT  17160.0 111405.0 17865.0 110060.0 ;
      RECT  17160.0 111405.0 17865.0 112750.0 ;
      RECT  17160.0 114095.0 17865.0 112750.0 ;
      RECT  17865.0 28015.0 18570.0 29360.0 ;
      RECT  17865.0 30705.0 18570.0 29360.0 ;
      RECT  17865.0 30705.0 18570.0 32050.0 ;
      RECT  17865.0 33395.0 18570.0 32050.0 ;
      RECT  17865.0 33395.0 18570.0 34740.0 ;
      RECT  17865.0 36085.0 18570.0 34740.0 ;
      RECT  17865.0 36085.0 18570.0 37430.0 ;
      RECT  17865.0 38775.0 18570.0 37430.0 ;
      RECT  17865.0 38775.0 18570.0 40120.0 ;
      RECT  17865.0 41465.0 18570.0 40120.0 ;
      RECT  17865.0 41465.0 18570.0 42810.0 ;
      RECT  17865.0 44155.0 18570.0 42810.0 ;
      RECT  17865.0 44155.0 18570.0 45500.0 ;
      RECT  17865.0 46845.0 18570.0 45500.0 ;
      RECT  17865.0 46845.0 18570.0 48190.0 ;
      RECT  17865.0 49535.0 18570.0 48190.0 ;
      RECT  17865.0 49535.0 18570.0 50880.0 ;
      RECT  17865.0 52225.0 18570.0 50880.0 ;
      RECT  17865.0 52225.0 18570.0 53570.0 ;
      RECT  17865.0 54915.0 18570.0 53570.0 ;
      RECT  17865.0 54915.0 18570.0 56260.0 ;
      RECT  17865.0 57605.0 18570.0 56260.0 ;
      RECT  17865.0 57605.0 18570.0 58950.0 ;
      RECT  17865.0 60295.0 18570.0 58950.0 ;
      RECT  17865.0 60295.0 18570.0 61640.0 ;
      RECT  17865.0 62985.0 18570.0 61640.0 ;
      RECT  17865.0 62985.0 18570.0 64330.0 ;
      RECT  17865.0 65675.0 18570.0 64330.0 ;
      RECT  17865.0 65675.0 18570.0 67020.0 ;
      RECT  17865.0 68365.0 18570.0 67020.0 ;
      RECT  17865.0 68365.0 18570.0 69710.0 ;
      RECT  17865.0 71055.0 18570.0 69710.0 ;
      RECT  17865.0 71055.0 18570.0 72400.0 ;
      RECT  17865.0 73745.0 18570.0 72400.0 ;
      RECT  17865.0 73745.0 18570.0 75090.0 ;
      RECT  17865.0 76435.0 18570.0 75090.0 ;
      RECT  17865.0 76435.0 18570.0 77780.0 ;
      RECT  17865.0 79125.0 18570.0 77780.0 ;
      RECT  17865.0 79125.0 18570.0 80470.0 ;
      RECT  17865.0 81815.0 18570.0 80470.0 ;
      RECT  17865.0 81815.0 18570.0 83160.0 ;
      RECT  17865.0 84505.0 18570.0 83160.0 ;
      RECT  17865.0 84505.0 18570.0 85850.0 ;
      RECT  17865.0 87195.0 18570.0 85850.0 ;
      RECT  17865.0 87195.0 18570.0 88540.0 ;
      RECT  17865.0 89885.0 18570.0 88540.0 ;
      RECT  17865.0 89885.0 18570.0 91230.0 ;
      RECT  17865.0 92575.0 18570.0 91230.0 ;
      RECT  17865.0 92575.0 18570.0 93920.0 ;
      RECT  17865.0 95265.0 18570.0 93920.0 ;
      RECT  17865.0 95265.0 18570.0 96610.0 ;
      RECT  17865.0 97955.0 18570.0 96610.0 ;
      RECT  17865.0 97955.0 18570.0 99300.0 ;
      RECT  17865.0 100645.0 18570.0 99300.0 ;
      RECT  17865.0 100645.0 18570.0 101990.0 ;
      RECT  17865.0 103335.0 18570.0 101990.0 ;
      RECT  17865.0 103335.0 18570.0 104680.0 ;
      RECT  17865.0 106025.0 18570.0 104680.0 ;
      RECT  17865.0 106025.0 18570.0 107370.0 ;
      RECT  17865.0 108715.0 18570.0 107370.0 ;
      RECT  17865.0 108715.0 18570.0 110060.0 ;
      RECT  17865.0 111405.0 18570.0 110060.0 ;
      RECT  17865.0 111405.0 18570.0 112750.0 ;
      RECT  17865.0 114095.0 18570.0 112750.0 ;
      RECT  18570.0 28015.0 19275.0 29360.0 ;
      RECT  18570.0 30705.0 19275.0 29360.0 ;
      RECT  18570.0 30705.0 19275.0 32050.0 ;
      RECT  18570.0 33395.0 19275.0 32050.0 ;
      RECT  18570.0 33395.0 19275.0 34740.0 ;
      RECT  18570.0 36085.0 19275.0 34740.0 ;
      RECT  18570.0 36085.0 19275.0 37430.0 ;
      RECT  18570.0 38775.0 19275.0 37430.0 ;
      RECT  18570.0 38775.0 19275.0 40120.0 ;
      RECT  18570.0 41465.0 19275.0 40120.0 ;
      RECT  18570.0 41465.0 19275.0 42810.0 ;
      RECT  18570.0 44155.0 19275.0 42810.0 ;
      RECT  18570.0 44155.0 19275.0 45500.0 ;
      RECT  18570.0 46845.0 19275.0 45500.0 ;
      RECT  18570.0 46845.0 19275.0 48190.0 ;
      RECT  18570.0 49535.0 19275.0 48190.0 ;
      RECT  18570.0 49535.0 19275.0 50880.0 ;
      RECT  18570.0 52225.0 19275.0 50880.0 ;
      RECT  18570.0 52225.0 19275.0 53570.0 ;
      RECT  18570.0 54915.0 19275.0 53570.0 ;
      RECT  18570.0 54915.0 19275.0 56260.0 ;
      RECT  18570.0 57605.0 19275.0 56260.0 ;
      RECT  18570.0 57605.0 19275.0 58950.0 ;
      RECT  18570.0 60295.0 19275.0 58950.0 ;
      RECT  18570.0 60295.0 19275.0 61640.0 ;
      RECT  18570.0 62985.0 19275.0 61640.0 ;
      RECT  18570.0 62985.0 19275.0 64330.0 ;
      RECT  18570.0 65675.0 19275.0 64330.0 ;
      RECT  18570.0 65675.0 19275.0 67020.0 ;
      RECT  18570.0 68365.0 19275.0 67020.0 ;
      RECT  18570.0 68365.0 19275.0 69710.0 ;
      RECT  18570.0 71055.0 19275.0 69710.0 ;
      RECT  18570.0 71055.0 19275.0 72400.0 ;
      RECT  18570.0 73745.0 19275.0 72400.0 ;
      RECT  18570.0 73745.0 19275.0 75090.0 ;
      RECT  18570.0 76435.0 19275.0 75090.0 ;
      RECT  18570.0 76435.0 19275.0 77780.0 ;
      RECT  18570.0 79125.0 19275.0 77780.0 ;
      RECT  18570.0 79125.0 19275.0 80470.0 ;
      RECT  18570.0 81815.0 19275.0 80470.0 ;
      RECT  18570.0 81815.0 19275.0 83160.0 ;
      RECT  18570.0 84505.0 19275.0 83160.0 ;
      RECT  18570.0 84505.0 19275.0 85850.0 ;
      RECT  18570.0 87195.0 19275.0 85850.0 ;
      RECT  18570.0 87195.0 19275.0 88540.0 ;
      RECT  18570.0 89885.0 19275.0 88540.0 ;
      RECT  18570.0 89885.0 19275.0 91230.0 ;
      RECT  18570.0 92575.0 19275.0 91230.0 ;
      RECT  18570.0 92575.0 19275.0 93920.0 ;
      RECT  18570.0 95265.0 19275.0 93920.0 ;
      RECT  18570.0 95265.0 19275.0 96610.0 ;
      RECT  18570.0 97955.0 19275.0 96610.0 ;
      RECT  18570.0 97955.0 19275.0 99300.0 ;
      RECT  18570.0 100645.0 19275.0 99300.0 ;
      RECT  18570.0 100645.0 19275.0 101990.0 ;
      RECT  18570.0 103335.0 19275.0 101990.0 ;
      RECT  18570.0 103335.0 19275.0 104680.0 ;
      RECT  18570.0 106025.0 19275.0 104680.0 ;
      RECT  18570.0 106025.0 19275.0 107370.0 ;
      RECT  18570.0 108715.0 19275.0 107370.0 ;
      RECT  18570.0 108715.0 19275.0 110060.0 ;
      RECT  18570.0 111405.0 19275.0 110060.0 ;
      RECT  18570.0 111405.0 19275.0 112750.0 ;
      RECT  18570.0 114095.0 19275.0 112750.0 ;
      RECT  19275.0 28015.0 19980.0 29360.0 ;
      RECT  19275.0 30705.0 19980.0 29360.0 ;
      RECT  19275.0 30705.0 19980.0 32050.0 ;
      RECT  19275.0 33395.0 19980.0 32050.0 ;
      RECT  19275.0 33395.0 19980.0 34740.0 ;
      RECT  19275.0 36085.0 19980.0 34740.0 ;
      RECT  19275.0 36085.0 19980.0 37430.0 ;
      RECT  19275.0 38775.0 19980.0 37430.0 ;
      RECT  19275.0 38775.0 19980.0 40120.0 ;
      RECT  19275.0 41465.0 19980.0 40120.0 ;
      RECT  19275.0 41465.0 19980.0 42810.0 ;
      RECT  19275.0 44155.0 19980.0 42810.0 ;
      RECT  19275.0 44155.0 19980.0 45500.0 ;
      RECT  19275.0 46845.0 19980.0 45500.0 ;
      RECT  19275.0 46845.0 19980.0 48190.0 ;
      RECT  19275.0 49535.0 19980.0 48190.0 ;
      RECT  19275.0 49535.0 19980.0 50880.0 ;
      RECT  19275.0 52225.0 19980.0 50880.0 ;
      RECT  19275.0 52225.0 19980.0 53570.0 ;
      RECT  19275.0 54915.0 19980.0 53570.0 ;
      RECT  19275.0 54915.0 19980.0 56260.0 ;
      RECT  19275.0 57605.0 19980.0 56260.0 ;
      RECT  19275.0 57605.0 19980.0 58950.0 ;
      RECT  19275.0 60295.0 19980.0 58950.0 ;
      RECT  19275.0 60295.0 19980.0 61640.0 ;
      RECT  19275.0 62985.0 19980.0 61640.0 ;
      RECT  19275.0 62985.0 19980.0 64330.0 ;
      RECT  19275.0 65675.0 19980.0 64330.0 ;
      RECT  19275.0 65675.0 19980.0 67020.0 ;
      RECT  19275.0 68365.0 19980.0 67020.0 ;
      RECT  19275.0 68365.0 19980.0 69710.0 ;
      RECT  19275.0 71055.0 19980.0 69710.0 ;
      RECT  19275.0 71055.0 19980.0 72400.0 ;
      RECT  19275.0 73745.0 19980.0 72400.0 ;
      RECT  19275.0 73745.0 19980.0 75090.0 ;
      RECT  19275.0 76435.0 19980.0 75090.0 ;
      RECT  19275.0 76435.0 19980.0 77780.0 ;
      RECT  19275.0 79125.0 19980.0 77780.0 ;
      RECT  19275.0 79125.0 19980.0 80470.0 ;
      RECT  19275.0 81815.0 19980.0 80470.0 ;
      RECT  19275.0 81815.0 19980.0 83160.0 ;
      RECT  19275.0 84505.0 19980.0 83160.0 ;
      RECT  19275.0 84505.0 19980.0 85850.0 ;
      RECT  19275.0 87195.0 19980.0 85850.0 ;
      RECT  19275.0 87195.0 19980.0 88540.0 ;
      RECT  19275.0 89885.0 19980.0 88540.0 ;
      RECT  19275.0 89885.0 19980.0 91230.0 ;
      RECT  19275.0 92575.0 19980.0 91230.0 ;
      RECT  19275.0 92575.0 19980.0 93920.0 ;
      RECT  19275.0 95265.0 19980.0 93920.0 ;
      RECT  19275.0 95265.0 19980.0 96610.0 ;
      RECT  19275.0 97955.0 19980.0 96610.0 ;
      RECT  19275.0 97955.0 19980.0 99300.0 ;
      RECT  19275.0 100645.0 19980.0 99300.0 ;
      RECT  19275.0 100645.0 19980.0 101990.0 ;
      RECT  19275.0 103335.0 19980.0 101990.0 ;
      RECT  19275.0 103335.0 19980.0 104680.0 ;
      RECT  19275.0 106025.0 19980.0 104680.0 ;
      RECT  19275.0 106025.0 19980.0 107370.0 ;
      RECT  19275.0 108715.0 19980.0 107370.0 ;
      RECT  19275.0 108715.0 19980.0 110060.0 ;
      RECT  19275.0 111405.0 19980.0 110060.0 ;
      RECT  19275.0 111405.0 19980.0 112750.0 ;
      RECT  19275.0 114095.0 19980.0 112750.0 ;
      RECT  19980.0 28015.0 20685.0 29360.0 ;
      RECT  19980.0 30705.0 20685.0 29360.0 ;
      RECT  19980.0 30705.0 20685.0 32050.0 ;
      RECT  19980.0 33395.0 20685.0 32050.0 ;
      RECT  19980.0 33395.0 20685.0 34740.0 ;
      RECT  19980.0 36085.0 20685.0 34740.0 ;
      RECT  19980.0 36085.0 20685.0 37430.0 ;
      RECT  19980.0 38775.0 20685.0 37430.0 ;
      RECT  19980.0 38775.0 20685.0 40120.0 ;
      RECT  19980.0 41465.0 20685.0 40120.0 ;
      RECT  19980.0 41465.0 20685.0 42810.0 ;
      RECT  19980.0 44155.0 20685.0 42810.0 ;
      RECT  19980.0 44155.0 20685.0 45500.0 ;
      RECT  19980.0 46845.0 20685.0 45500.0 ;
      RECT  19980.0 46845.0 20685.0 48190.0 ;
      RECT  19980.0 49535.0 20685.0 48190.0 ;
      RECT  19980.0 49535.0 20685.0 50880.0 ;
      RECT  19980.0 52225.0 20685.0 50880.0 ;
      RECT  19980.0 52225.0 20685.0 53570.0 ;
      RECT  19980.0 54915.0 20685.0 53570.0 ;
      RECT  19980.0 54915.0 20685.0 56260.0 ;
      RECT  19980.0 57605.0 20685.0 56260.0 ;
      RECT  19980.0 57605.0 20685.0 58950.0 ;
      RECT  19980.0 60295.0 20685.0 58950.0 ;
      RECT  19980.0 60295.0 20685.0 61640.0 ;
      RECT  19980.0 62985.0 20685.0 61640.0 ;
      RECT  19980.0 62985.0 20685.0 64330.0 ;
      RECT  19980.0 65675.0 20685.0 64330.0 ;
      RECT  19980.0 65675.0 20685.0 67020.0 ;
      RECT  19980.0 68365.0 20685.0 67020.0 ;
      RECT  19980.0 68365.0 20685.0 69710.0 ;
      RECT  19980.0 71055.0 20685.0 69710.0 ;
      RECT  19980.0 71055.0 20685.0 72400.0 ;
      RECT  19980.0 73745.0 20685.0 72400.0 ;
      RECT  19980.0 73745.0 20685.0 75090.0 ;
      RECT  19980.0 76435.0 20685.0 75090.0 ;
      RECT  19980.0 76435.0 20685.0 77780.0 ;
      RECT  19980.0 79125.0 20685.0 77780.0 ;
      RECT  19980.0 79125.0 20685.0 80470.0 ;
      RECT  19980.0 81815.0 20685.0 80470.0 ;
      RECT  19980.0 81815.0 20685.0 83160.0 ;
      RECT  19980.0 84505.0 20685.0 83160.0 ;
      RECT  19980.0 84505.0 20685.0 85850.0 ;
      RECT  19980.0 87195.0 20685.0 85850.0 ;
      RECT  19980.0 87195.0 20685.0 88540.0 ;
      RECT  19980.0 89885.0 20685.0 88540.0 ;
      RECT  19980.0 89885.0 20685.0 91230.0 ;
      RECT  19980.0 92575.0 20685.0 91230.0 ;
      RECT  19980.0 92575.0 20685.0 93920.0 ;
      RECT  19980.0 95265.0 20685.0 93920.0 ;
      RECT  19980.0 95265.0 20685.0 96610.0 ;
      RECT  19980.0 97955.0 20685.0 96610.0 ;
      RECT  19980.0 97955.0 20685.0 99300.0 ;
      RECT  19980.0 100645.0 20685.0 99300.0 ;
      RECT  19980.0 100645.0 20685.0 101990.0 ;
      RECT  19980.0 103335.0 20685.0 101990.0 ;
      RECT  19980.0 103335.0 20685.0 104680.0 ;
      RECT  19980.0 106025.0 20685.0 104680.0 ;
      RECT  19980.0 106025.0 20685.0 107370.0 ;
      RECT  19980.0 108715.0 20685.0 107370.0 ;
      RECT  19980.0 108715.0 20685.0 110060.0 ;
      RECT  19980.0 111405.0 20685.0 110060.0 ;
      RECT  19980.0 111405.0 20685.0 112750.0 ;
      RECT  19980.0 114095.0 20685.0 112750.0 ;
      RECT  20685.0 28015.0 21390.0 29360.0 ;
      RECT  20685.0 30705.0 21390.0 29360.0 ;
      RECT  20685.0 30705.0 21390.0 32050.0 ;
      RECT  20685.0 33395.0 21390.0 32050.0 ;
      RECT  20685.0 33395.0 21390.0 34740.0 ;
      RECT  20685.0 36085.0 21390.0 34740.0 ;
      RECT  20685.0 36085.0 21390.0 37430.0 ;
      RECT  20685.0 38775.0 21390.0 37430.0 ;
      RECT  20685.0 38775.0 21390.0 40120.0 ;
      RECT  20685.0 41465.0 21390.0 40120.0 ;
      RECT  20685.0 41465.0 21390.0 42810.0 ;
      RECT  20685.0 44155.0 21390.0 42810.0 ;
      RECT  20685.0 44155.0 21390.0 45500.0 ;
      RECT  20685.0 46845.0 21390.0 45500.0 ;
      RECT  20685.0 46845.0 21390.0 48190.0 ;
      RECT  20685.0 49535.0 21390.0 48190.0 ;
      RECT  20685.0 49535.0 21390.0 50880.0 ;
      RECT  20685.0 52225.0 21390.0 50880.0 ;
      RECT  20685.0 52225.0 21390.0 53570.0 ;
      RECT  20685.0 54915.0 21390.0 53570.0 ;
      RECT  20685.0 54915.0 21390.0 56260.0 ;
      RECT  20685.0 57605.0 21390.0 56260.0 ;
      RECT  20685.0 57605.0 21390.0 58950.0 ;
      RECT  20685.0 60295.0 21390.0 58950.0 ;
      RECT  20685.0 60295.0 21390.0 61640.0 ;
      RECT  20685.0 62985.0 21390.0 61640.0 ;
      RECT  20685.0 62985.0 21390.0 64330.0 ;
      RECT  20685.0 65675.0 21390.0 64330.0 ;
      RECT  20685.0 65675.0 21390.0 67020.0 ;
      RECT  20685.0 68365.0 21390.0 67020.0 ;
      RECT  20685.0 68365.0 21390.0 69710.0 ;
      RECT  20685.0 71055.0 21390.0 69710.0 ;
      RECT  20685.0 71055.0 21390.0 72400.0 ;
      RECT  20685.0 73745.0 21390.0 72400.0 ;
      RECT  20685.0 73745.0 21390.0 75090.0 ;
      RECT  20685.0 76435.0 21390.0 75090.0 ;
      RECT  20685.0 76435.0 21390.0 77780.0 ;
      RECT  20685.0 79125.0 21390.0 77780.0 ;
      RECT  20685.0 79125.0 21390.0 80470.0 ;
      RECT  20685.0 81815.0 21390.0 80470.0 ;
      RECT  20685.0 81815.0 21390.0 83160.0 ;
      RECT  20685.0 84505.0 21390.0 83160.0 ;
      RECT  20685.0 84505.0 21390.0 85850.0 ;
      RECT  20685.0 87195.0 21390.0 85850.0 ;
      RECT  20685.0 87195.0 21390.0 88540.0 ;
      RECT  20685.0 89885.0 21390.0 88540.0 ;
      RECT  20685.0 89885.0 21390.0 91230.0 ;
      RECT  20685.0 92575.0 21390.0 91230.0 ;
      RECT  20685.0 92575.0 21390.0 93920.0 ;
      RECT  20685.0 95265.0 21390.0 93920.0 ;
      RECT  20685.0 95265.0 21390.0 96610.0 ;
      RECT  20685.0 97955.0 21390.0 96610.0 ;
      RECT  20685.0 97955.0 21390.0 99300.0 ;
      RECT  20685.0 100645.0 21390.0 99300.0 ;
      RECT  20685.0 100645.0 21390.0 101990.0 ;
      RECT  20685.0 103335.0 21390.0 101990.0 ;
      RECT  20685.0 103335.0 21390.0 104680.0 ;
      RECT  20685.0 106025.0 21390.0 104680.0 ;
      RECT  20685.0 106025.0 21390.0 107370.0 ;
      RECT  20685.0 108715.0 21390.0 107370.0 ;
      RECT  20685.0 108715.0 21390.0 110060.0 ;
      RECT  20685.0 111405.0 21390.0 110060.0 ;
      RECT  20685.0 111405.0 21390.0 112750.0 ;
      RECT  20685.0 114095.0 21390.0 112750.0 ;
      RECT  21390.0 28015.0 22095.0 29360.0 ;
      RECT  21390.0 30705.0 22095.0 29360.0 ;
      RECT  21390.0 30705.0 22095.0 32050.0 ;
      RECT  21390.0 33395.0 22095.0 32050.0 ;
      RECT  21390.0 33395.0 22095.0 34740.0 ;
      RECT  21390.0 36085.0 22095.0 34740.0 ;
      RECT  21390.0 36085.0 22095.0 37430.0 ;
      RECT  21390.0 38775.0 22095.0 37430.0 ;
      RECT  21390.0 38775.0 22095.0 40120.0 ;
      RECT  21390.0 41465.0 22095.0 40120.0 ;
      RECT  21390.0 41465.0 22095.0 42810.0 ;
      RECT  21390.0 44155.0 22095.0 42810.0 ;
      RECT  21390.0 44155.0 22095.0 45500.0 ;
      RECT  21390.0 46845.0 22095.0 45500.0 ;
      RECT  21390.0 46845.0 22095.0 48190.0 ;
      RECT  21390.0 49535.0 22095.0 48190.0 ;
      RECT  21390.0 49535.0 22095.0 50880.0 ;
      RECT  21390.0 52225.0 22095.0 50880.0 ;
      RECT  21390.0 52225.0 22095.0 53570.0 ;
      RECT  21390.0 54915.0 22095.0 53570.0 ;
      RECT  21390.0 54915.0 22095.0 56260.0 ;
      RECT  21390.0 57605.0 22095.0 56260.0 ;
      RECT  21390.0 57605.0 22095.0 58950.0 ;
      RECT  21390.0 60295.0 22095.0 58950.0 ;
      RECT  21390.0 60295.0 22095.0 61640.0 ;
      RECT  21390.0 62985.0 22095.0 61640.0 ;
      RECT  21390.0 62985.0 22095.0 64330.0 ;
      RECT  21390.0 65675.0 22095.0 64330.0 ;
      RECT  21390.0 65675.0 22095.0 67020.0 ;
      RECT  21390.0 68365.0 22095.0 67020.0 ;
      RECT  21390.0 68365.0 22095.0 69710.0 ;
      RECT  21390.0 71055.0 22095.0 69710.0 ;
      RECT  21390.0 71055.0 22095.0 72400.0 ;
      RECT  21390.0 73745.0 22095.0 72400.0 ;
      RECT  21390.0 73745.0 22095.0 75090.0 ;
      RECT  21390.0 76435.0 22095.0 75090.0 ;
      RECT  21390.0 76435.0 22095.0 77780.0 ;
      RECT  21390.0 79125.0 22095.0 77780.0 ;
      RECT  21390.0 79125.0 22095.0 80470.0 ;
      RECT  21390.0 81815.0 22095.0 80470.0 ;
      RECT  21390.0 81815.0 22095.0 83160.0 ;
      RECT  21390.0 84505.0 22095.0 83160.0 ;
      RECT  21390.0 84505.0 22095.0 85850.0 ;
      RECT  21390.0 87195.0 22095.0 85850.0 ;
      RECT  21390.0 87195.0 22095.0 88540.0 ;
      RECT  21390.0 89885.0 22095.0 88540.0 ;
      RECT  21390.0 89885.0 22095.0 91230.0 ;
      RECT  21390.0 92575.0 22095.0 91230.0 ;
      RECT  21390.0 92575.0 22095.0 93920.0 ;
      RECT  21390.0 95265.0 22095.0 93920.0 ;
      RECT  21390.0 95265.0 22095.0 96610.0 ;
      RECT  21390.0 97955.0 22095.0 96610.0 ;
      RECT  21390.0 97955.0 22095.0 99300.0 ;
      RECT  21390.0 100645.0 22095.0 99300.0 ;
      RECT  21390.0 100645.0 22095.0 101990.0 ;
      RECT  21390.0 103335.0 22095.0 101990.0 ;
      RECT  21390.0 103335.0 22095.0 104680.0 ;
      RECT  21390.0 106025.0 22095.0 104680.0 ;
      RECT  21390.0 106025.0 22095.0 107370.0 ;
      RECT  21390.0 108715.0 22095.0 107370.0 ;
      RECT  21390.0 108715.0 22095.0 110060.0 ;
      RECT  21390.0 111405.0 22095.0 110060.0 ;
      RECT  21390.0 111405.0 22095.0 112750.0 ;
      RECT  21390.0 114095.0 22095.0 112750.0 ;
      RECT  22095.0 28015.0 22800.0 29360.0 ;
      RECT  22095.0 30705.0 22800.0 29360.0 ;
      RECT  22095.0 30705.0 22800.0 32050.0 ;
      RECT  22095.0 33395.0 22800.0 32050.0 ;
      RECT  22095.0 33395.0 22800.0 34740.0 ;
      RECT  22095.0 36085.0 22800.0 34740.0 ;
      RECT  22095.0 36085.0 22800.0 37430.0 ;
      RECT  22095.0 38775.0 22800.0 37430.0 ;
      RECT  22095.0 38775.0 22800.0 40120.0 ;
      RECT  22095.0 41465.0 22800.0 40120.0 ;
      RECT  22095.0 41465.0 22800.0 42810.0 ;
      RECT  22095.0 44155.0 22800.0 42810.0 ;
      RECT  22095.0 44155.0 22800.0 45500.0 ;
      RECT  22095.0 46845.0 22800.0 45500.0 ;
      RECT  22095.0 46845.0 22800.0 48190.0 ;
      RECT  22095.0 49535.0 22800.0 48190.0 ;
      RECT  22095.0 49535.0 22800.0 50880.0 ;
      RECT  22095.0 52225.0 22800.0 50880.0 ;
      RECT  22095.0 52225.0 22800.0 53570.0 ;
      RECT  22095.0 54915.0 22800.0 53570.0 ;
      RECT  22095.0 54915.0 22800.0 56260.0 ;
      RECT  22095.0 57605.0 22800.0 56260.0 ;
      RECT  22095.0 57605.0 22800.0 58950.0 ;
      RECT  22095.0 60295.0 22800.0 58950.0 ;
      RECT  22095.0 60295.0 22800.0 61640.0 ;
      RECT  22095.0 62985.0 22800.0 61640.0 ;
      RECT  22095.0 62985.0 22800.0 64330.0 ;
      RECT  22095.0 65675.0 22800.0 64330.0 ;
      RECT  22095.0 65675.0 22800.0 67020.0 ;
      RECT  22095.0 68365.0 22800.0 67020.0 ;
      RECT  22095.0 68365.0 22800.0 69710.0 ;
      RECT  22095.0 71055.0 22800.0 69710.0 ;
      RECT  22095.0 71055.0 22800.0 72400.0 ;
      RECT  22095.0 73745.0 22800.0 72400.0 ;
      RECT  22095.0 73745.0 22800.0 75090.0 ;
      RECT  22095.0 76435.0 22800.0 75090.0 ;
      RECT  22095.0 76435.0 22800.0 77780.0 ;
      RECT  22095.0 79125.0 22800.0 77780.0 ;
      RECT  22095.0 79125.0 22800.0 80470.0 ;
      RECT  22095.0 81815.0 22800.0 80470.0 ;
      RECT  22095.0 81815.0 22800.0 83160.0 ;
      RECT  22095.0 84505.0 22800.0 83160.0 ;
      RECT  22095.0 84505.0 22800.0 85850.0 ;
      RECT  22095.0 87195.0 22800.0 85850.0 ;
      RECT  22095.0 87195.0 22800.0 88540.0 ;
      RECT  22095.0 89885.0 22800.0 88540.0 ;
      RECT  22095.0 89885.0 22800.0 91230.0 ;
      RECT  22095.0 92575.0 22800.0 91230.0 ;
      RECT  22095.0 92575.0 22800.0 93920.0 ;
      RECT  22095.0 95265.0 22800.0 93920.0 ;
      RECT  22095.0 95265.0 22800.0 96610.0 ;
      RECT  22095.0 97955.0 22800.0 96610.0 ;
      RECT  22095.0 97955.0 22800.0 99300.0 ;
      RECT  22095.0 100645.0 22800.0 99300.0 ;
      RECT  22095.0 100645.0 22800.0 101990.0 ;
      RECT  22095.0 103335.0 22800.0 101990.0 ;
      RECT  22095.0 103335.0 22800.0 104680.0 ;
      RECT  22095.0 106025.0 22800.0 104680.0 ;
      RECT  22095.0 106025.0 22800.0 107370.0 ;
      RECT  22095.0 108715.0 22800.0 107370.0 ;
      RECT  22095.0 108715.0 22800.0 110060.0 ;
      RECT  22095.0 111405.0 22800.0 110060.0 ;
      RECT  22095.0 111405.0 22800.0 112750.0 ;
      RECT  22095.0 114095.0 22800.0 112750.0 ;
      RECT  22800.0 28015.0 23505.0 29360.0 ;
      RECT  22800.0 30705.0 23505.0 29360.0 ;
      RECT  22800.0 30705.0 23505.0 32050.0 ;
      RECT  22800.0 33395.0 23505.0 32050.0 ;
      RECT  22800.0 33395.0 23505.0 34740.0 ;
      RECT  22800.0 36085.0 23505.0 34740.0 ;
      RECT  22800.0 36085.0 23505.0 37430.0 ;
      RECT  22800.0 38775.0 23505.0 37430.0 ;
      RECT  22800.0 38775.0 23505.0 40120.0 ;
      RECT  22800.0 41465.0 23505.0 40120.0 ;
      RECT  22800.0 41465.0 23505.0 42810.0 ;
      RECT  22800.0 44155.0 23505.0 42810.0 ;
      RECT  22800.0 44155.0 23505.0 45500.0 ;
      RECT  22800.0 46845.0 23505.0 45500.0 ;
      RECT  22800.0 46845.0 23505.0 48190.0 ;
      RECT  22800.0 49535.0 23505.0 48190.0 ;
      RECT  22800.0 49535.0 23505.0 50880.0 ;
      RECT  22800.0 52225.0 23505.0 50880.0 ;
      RECT  22800.0 52225.0 23505.0 53570.0 ;
      RECT  22800.0 54915.0 23505.0 53570.0 ;
      RECT  22800.0 54915.0 23505.0 56260.0 ;
      RECT  22800.0 57605.0 23505.0 56260.0 ;
      RECT  22800.0 57605.0 23505.0 58950.0 ;
      RECT  22800.0 60295.0 23505.0 58950.0 ;
      RECT  22800.0 60295.0 23505.0 61640.0 ;
      RECT  22800.0 62985.0 23505.0 61640.0 ;
      RECT  22800.0 62985.0 23505.0 64330.0 ;
      RECT  22800.0 65675.0 23505.0 64330.0 ;
      RECT  22800.0 65675.0 23505.0 67020.0 ;
      RECT  22800.0 68365.0 23505.0 67020.0 ;
      RECT  22800.0 68365.0 23505.0 69710.0 ;
      RECT  22800.0 71055.0 23505.0 69710.0 ;
      RECT  22800.0 71055.0 23505.0 72400.0 ;
      RECT  22800.0 73745.0 23505.0 72400.0 ;
      RECT  22800.0 73745.0 23505.0 75090.0 ;
      RECT  22800.0 76435.0 23505.0 75090.0 ;
      RECT  22800.0 76435.0 23505.0 77780.0 ;
      RECT  22800.0 79125.0 23505.0 77780.0 ;
      RECT  22800.0 79125.0 23505.0 80470.0 ;
      RECT  22800.0 81815.0 23505.0 80470.0 ;
      RECT  22800.0 81815.0 23505.0 83160.0 ;
      RECT  22800.0 84505.0 23505.0 83160.0 ;
      RECT  22800.0 84505.0 23505.0 85850.0 ;
      RECT  22800.0 87195.0 23505.0 85850.0 ;
      RECT  22800.0 87195.0 23505.0 88540.0 ;
      RECT  22800.0 89885.0 23505.0 88540.0 ;
      RECT  22800.0 89885.0 23505.0 91230.0 ;
      RECT  22800.0 92575.0 23505.0 91230.0 ;
      RECT  22800.0 92575.0 23505.0 93920.0 ;
      RECT  22800.0 95265.0 23505.0 93920.0 ;
      RECT  22800.0 95265.0 23505.0 96610.0 ;
      RECT  22800.0 97955.0 23505.0 96610.0 ;
      RECT  22800.0 97955.0 23505.0 99300.0 ;
      RECT  22800.0 100645.0 23505.0 99300.0 ;
      RECT  22800.0 100645.0 23505.0 101990.0 ;
      RECT  22800.0 103335.0 23505.0 101990.0 ;
      RECT  22800.0 103335.0 23505.0 104680.0 ;
      RECT  22800.0 106025.0 23505.0 104680.0 ;
      RECT  22800.0 106025.0 23505.0 107370.0 ;
      RECT  22800.0 108715.0 23505.0 107370.0 ;
      RECT  22800.0 108715.0 23505.0 110060.0 ;
      RECT  22800.0 111405.0 23505.0 110060.0 ;
      RECT  22800.0 111405.0 23505.0 112750.0 ;
      RECT  22800.0 114095.0 23505.0 112750.0 ;
      RECT  23505.0 28015.0 24210.0 29360.0 ;
      RECT  23505.0 30705.0 24210.0 29360.0 ;
      RECT  23505.0 30705.0 24210.0 32050.0 ;
      RECT  23505.0 33395.0 24210.0 32050.0 ;
      RECT  23505.0 33395.0 24210.0 34740.0 ;
      RECT  23505.0 36085.0 24210.0 34740.0 ;
      RECT  23505.0 36085.0 24210.0 37430.0 ;
      RECT  23505.0 38775.0 24210.0 37430.0 ;
      RECT  23505.0 38775.0 24210.0 40120.0 ;
      RECT  23505.0 41465.0 24210.0 40120.0 ;
      RECT  23505.0 41465.0 24210.0 42810.0 ;
      RECT  23505.0 44155.0 24210.0 42810.0 ;
      RECT  23505.0 44155.0 24210.0 45500.0 ;
      RECT  23505.0 46845.0 24210.0 45500.0 ;
      RECT  23505.0 46845.0 24210.0 48190.0 ;
      RECT  23505.0 49535.0 24210.0 48190.0 ;
      RECT  23505.0 49535.0 24210.0 50880.0 ;
      RECT  23505.0 52225.0 24210.0 50880.0 ;
      RECT  23505.0 52225.0 24210.0 53570.0 ;
      RECT  23505.0 54915.0 24210.0 53570.0 ;
      RECT  23505.0 54915.0 24210.0 56260.0 ;
      RECT  23505.0 57605.0 24210.0 56260.0 ;
      RECT  23505.0 57605.0 24210.0 58950.0 ;
      RECT  23505.0 60295.0 24210.0 58950.0 ;
      RECT  23505.0 60295.0 24210.0 61640.0 ;
      RECT  23505.0 62985.0 24210.0 61640.0 ;
      RECT  23505.0 62985.0 24210.0 64330.0 ;
      RECT  23505.0 65675.0 24210.0 64330.0 ;
      RECT  23505.0 65675.0 24210.0 67020.0 ;
      RECT  23505.0 68365.0 24210.0 67020.0 ;
      RECT  23505.0 68365.0 24210.0 69710.0 ;
      RECT  23505.0 71055.0 24210.0 69710.0 ;
      RECT  23505.0 71055.0 24210.0 72400.0 ;
      RECT  23505.0 73745.0 24210.0 72400.0 ;
      RECT  23505.0 73745.0 24210.0 75090.0 ;
      RECT  23505.0 76435.0 24210.0 75090.0 ;
      RECT  23505.0 76435.0 24210.0 77780.0 ;
      RECT  23505.0 79125.0 24210.0 77780.0 ;
      RECT  23505.0 79125.0 24210.0 80470.0 ;
      RECT  23505.0 81815.0 24210.0 80470.0 ;
      RECT  23505.0 81815.0 24210.0 83160.0 ;
      RECT  23505.0 84505.0 24210.0 83160.0 ;
      RECT  23505.0 84505.0 24210.0 85850.0 ;
      RECT  23505.0 87195.0 24210.0 85850.0 ;
      RECT  23505.0 87195.0 24210.0 88540.0 ;
      RECT  23505.0 89885.0 24210.0 88540.0 ;
      RECT  23505.0 89885.0 24210.0 91230.0 ;
      RECT  23505.0 92575.0 24210.0 91230.0 ;
      RECT  23505.0 92575.0 24210.0 93920.0 ;
      RECT  23505.0 95265.0 24210.0 93920.0 ;
      RECT  23505.0 95265.0 24210.0 96610.0 ;
      RECT  23505.0 97955.0 24210.0 96610.0 ;
      RECT  23505.0 97955.0 24210.0 99300.0 ;
      RECT  23505.0 100645.0 24210.0 99300.0 ;
      RECT  23505.0 100645.0 24210.0 101990.0 ;
      RECT  23505.0 103335.0 24210.0 101990.0 ;
      RECT  23505.0 103335.0 24210.0 104680.0 ;
      RECT  23505.0 106025.0 24210.0 104680.0 ;
      RECT  23505.0 106025.0 24210.0 107370.0 ;
      RECT  23505.0 108715.0 24210.0 107370.0 ;
      RECT  23505.0 108715.0 24210.0 110060.0 ;
      RECT  23505.0 111405.0 24210.0 110060.0 ;
      RECT  23505.0 111405.0 24210.0 112750.0 ;
      RECT  23505.0 114095.0 24210.0 112750.0 ;
      RECT  24210.0 28015.0 24915.0 29360.0 ;
      RECT  24210.0 30705.0 24915.0 29360.0 ;
      RECT  24210.0 30705.0 24915.0 32050.0 ;
      RECT  24210.0 33395.0 24915.0 32050.0 ;
      RECT  24210.0 33395.0 24915.0 34740.0 ;
      RECT  24210.0 36085.0 24915.0 34740.0 ;
      RECT  24210.0 36085.0 24915.0 37430.0 ;
      RECT  24210.0 38775.0 24915.0 37430.0 ;
      RECT  24210.0 38775.0 24915.0 40120.0 ;
      RECT  24210.0 41465.0 24915.0 40120.0 ;
      RECT  24210.0 41465.0 24915.0 42810.0 ;
      RECT  24210.0 44155.0 24915.0 42810.0 ;
      RECT  24210.0 44155.0 24915.0 45500.0 ;
      RECT  24210.0 46845.0 24915.0 45500.0 ;
      RECT  24210.0 46845.0 24915.0 48190.0 ;
      RECT  24210.0 49535.0 24915.0 48190.0 ;
      RECT  24210.0 49535.0 24915.0 50880.0 ;
      RECT  24210.0 52225.0 24915.0 50880.0 ;
      RECT  24210.0 52225.0 24915.0 53570.0 ;
      RECT  24210.0 54915.0 24915.0 53570.0 ;
      RECT  24210.0 54915.0 24915.0 56260.0 ;
      RECT  24210.0 57605.0 24915.0 56260.0 ;
      RECT  24210.0 57605.0 24915.0 58950.0 ;
      RECT  24210.0 60295.0 24915.0 58950.0 ;
      RECT  24210.0 60295.0 24915.0 61640.0 ;
      RECT  24210.0 62985.0 24915.0 61640.0 ;
      RECT  24210.0 62985.0 24915.0 64330.0 ;
      RECT  24210.0 65675.0 24915.0 64330.0 ;
      RECT  24210.0 65675.0 24915.0 67020.0 ;
      RECT  24210.0 68365.0 24915.0 67020.0 ;
      RECT  24210.0 68365.0 24915.0 69710.0 ;
      RECT  24210.0 71055.0 24915.0 69710.0 ;
      RECT  24210.0 71055.0 24915.0 72400.0 ;
      RECT  24210.0 73745.0 24915.0 72400.0 ;
      RECT  24210.0 73745.0 24915.0 75090.0 ;
      RECT  24210.0 76435.0 24915.0 75090.0 ;
      RECT  24210.0 76435.0 24915.0 77780.0 ;
      RECT  24210.0 79125.0 24915.0 77780.0 ;
      RECT  24210.0 79125.0 24915.0 80470.0 ;
      RECT  24210.0 81815.0 24915.0 80470.0 ;
      RECT  24210.0 81815.0 24915.0 83160.0 ;
      RECT  24210.0 84505.0 24915.0 83160.0 ;
      RECT  24210.0 84505.0 24915.0 85850.0 ;
      RECT  24210.0 87195.0 24915.0 85850.0 ;
      RECT  24210.0 87195.0 24915.0 88540.0 ;
      RECT  24210.0 89885.0 24915.0 88540.0 ;
      RECT  24210.0 89885.0 24915.0 91230.0 ;
      RECT  24210.0 92575.0 24915.0 91230.0 ;
      RECT  24210.0 92575.0 24915.0 93920.0 ;
      RECT  24210.0 95265.0 24915.0 93920.0 ;
      RECT  24210.0 95265.0 24915.0 96610.0 ;
      RECT  24210.0 97955.0 24915.0 96610.0 ;
      RECT  24210.0 97955.0 24915.0 99300.0 ;
      RECT  24210.0 100645.0 24915.0 99300.0 ;
      RECT  24210.0 100645.0 24915.0 101990.0 ;
      RECT  24210.0 103335.0 24915.0 101990.0 ;
      RECT  24210.0 103335.0 24915.0 104680.0 ;
      RECT  24210.0 106025.0 24915.0 104680.0 ;
      RECT  24210.0 106025.0 24915.0 107370.0 ;
      RECT  24210.0 108715.0 24915.0 107370.0 ;
      RECT  24210.0 108715.0 24915.0 110060.0 ;
      RECT  24210.0 111405.0 24915.0 110060.0 ;
      RECT  24210.0 111405.0 24915.0 112750.0 ;
      RECT  24210.0 114095.0 24915.0 112750.0 ;
      RECT  24915.0 28015.0 25620.0 29360.0 ;
      RECT  24915.0 30705.0 25620.0 29360.0 ;
      RECT  24915.0 30705.0 25620.0 32050.0 ;
      RECT  24915.0 33395.0 25620.0 32050.0 ;
      RECT  24915.0 33395.0 25620.0 34740.0 ;
      RECT  24915.0 36085.0 25620.0 34740.0 ;
      RECT  24915.0 36085.0 25620.0 37430.0 ;
      RECT  24915.0 38775.0 25620.0 37430.0 ;
      RECT  24915.0 38775.0 25620.0 40120.0 ;
      RECT  24915.0 41465.0 25620.0 40120.0 ;
      RECT  24915.0 41465.0 25620.0 42810.0 ;
      RECT  24915.0 44155.0 25620.0 42810.0 ;
      RECT  24915.0 44155.0 25620.0 45500.0 ;
      RECT  24915.0 46845.0 25620.0 45500.0 ;
      RECT  24915.0 46845.0 25620.0 48190.0 ;
      RECT  24915.0 49535.0 25620.0 48190.0 ;
      RECT  24915.0 49535.0 25620.0 50880.0 ;
      RECT  24915.0 52225.0 25620.0 50880.0 ;
      RECT  24915.0 52225.0 25620.0 53570.0 ;
      RECT  24915.0 54915.0 25620.0 53570.0 ;
      RECT  24915.0 54915.0 25620.0 56260.0 ;
      RECT  24915.0 57605.0 25620.0 56260.0 ;
      RECT  24915.0 57605.0 25620.0 58950.0 ;
      RECT  24915.0 60295.0 25620.0 58950.0 ;
      RECT  24915.0 60295.0 25620.0 61640.0 ;
      RECT  24915.0 62985.0 25620.0 61640.0 ;
      RECT  24915.0 62985.0 25620.0 64330.0 ;
      RECT  24915.0 65675.0 25620.0 64330.0 ;
      RECT  24915.0 65675.0 25620.0 67020.0 ;
      RECT  24915.0 68365.0 25620.0 67020.0 ;
      RECT  24915.0 68365.0 25620.0 69710.0 ;
      RECT  24915.0 71055.0 25620.0 69710.0 ;
      RECT  24915.0 71055.0 25620.0 72400.0 ;
      RECT  24915.0 73745.0 25620.0 72400.0 ;
      RECT  24915.0 73745.0 25620.0 75090.0 ;
      RECT  24915.0 76435.0 25620.0 75090.0 ;
      RECT  24915.0 76435.0 25620.0 77780.0 ;
      RECT  24915.0 79125.0 25620.0 77780.0 ;
      RECT  24915.0 79125.0 25620.0 80470.0 ;
      RECT  24915.0 81815.0 25620.0 80470.0 ;
      RECT  24915.0 81815.0 25620.0 83160.0 ;
      RECT  24915.0 84505.0 25620.0 83160.0 ;
      RECT  24915.0 84505.0 25620.0 85850.0 ;
      RECT  24915.0 87195.0 25620.0 85850.0 ;
      RECT  24915.0 87195.0 25620.0 88540.0 ;
      RECT  24915.0 89885.0 25620.0 88540.0 ;
      RECT  24915.0 89885.0 25620.0 91230.0 ;
      RECT  24915.0 92575.0 25620.0 91230.0 ;
      RECT  24915.0 92575.0 25620.0 93920.0 ;
      RECT  24915.0 95265.0 25620.0 93920.0 ;
      RECT  24915.0 95265.0 25620.0 96610.0 ;
      RECT  24915.0 97955.0 25620.0 96610.0 ;
      RECT  24915.0 97955.0 25620.0 99300.0 ;
      RECT  24915.0 100645.0 25620.0 99300.0 ;
      RECT  24915.0 100645.0 25620.0 101990.0 ;
      RECT  24915.0 103335.0 25620.0 101990.0 ;
      RECT  24915.0 103335.0 25620.0 104680.0 ;
      RECT  24915.0 106025.0 25620.0 104680.0 ;
      RECT  24915.0 106025.0 25620.0 107370.0 ;
      RECT  24915.0 108715.0 25620.0 107370.0 ;
      RECT  24915.0 108715.0 25620.0 110060.0 ;
      RECT  24915.0 111405.0 25620.0 110060.0 ;
      RECT  24915.0 111405.0 25620.0 112750.0 ;
      RECT  24915.0 114095.0 25620.0 112750.0 ;
      RECT  25620.0 28015.0 26325.0 29360.0 ;
      RECT  25620.0 30705.0 26325.0 29360.0 ;
      RECT  25620.0 30705.0 26325.0 32050.0 ;
      RECT  25620.0 33395.0 26325.0 32050.0 ;
      RECT  25620.0 33395.0 26325.0 34740.0 ;
      RECT  25620.0 36085.0 26325.0 34740.0 ;
      RECT  25620.0 36085.0 26325.0 37430.0 ;
      RECT  25620.0 38775.0 26325.0 37430.0 ;
      RECT  25620.0 38775.0 26325.0 40120.0 ;
      RECT  25620.0 41465.0 26325.0 40120.0 ;
      RECT  25620.0 41465.0 26325.0 42810.0 ;
      RECT  25620.0 44155.0 26325.0 42810.0 ;
      RECT  25620.0 44155.0 26325.0 45500.0 ;
      RECT  25620.0 46845.0 26325.0 45500.0 ;
      RECT  25620.0 46845.0 26325.0 48190.0 ;
      RECT  25620.0 49535.0 26325.0 48190.0 ;
      RECT  25620.0 49535.0 26325.0 50880.0 ;
      RECT  25620.0 52225.0 26325.0 50880.0 ;
      RECT  25620.0 52225.0 26325.0 53570.0 ;
      RECT  25620.0 54915.0 26325.0 53570.0 ;
      RECT  25620.0 54915.0 26325.0 56260.0 ;
      RECT  25620.0 57605.0 26325.0 56260.0 ;
      RECT  25620.0 57605.0 26325.0 58950.0 ;
      RECT  25620.0 60295.0 26325.0 58950.0 ;
      RECT  25620.0 60295.0 26325.0 61640.0 ;
      RECT  25620.0 62985.0 26325.0 61640.0 ;
      RECT  25620.0 62985.0 26325.0 64330.0 ;
      RECT  25620.0 65675.0 26325.0 64330.0 ;
      RECT  25620.0 65675.0 26325.0 67020.0 ;
      RECT  25620.0 68365.0 26325.0 67020.0 ;
      RECT  25620.0 68365.0 26325.0 69710.0 ;
      RECT  25620.0 71055.0 26325.0 69710.0 ;
      RECT  25620.0 71055.0 26325.0 72400.0 ;
      RECT  25620.0 73745.0 26325.0 72400.0 ;
      RECT  25620.0 73745.0 26325.0 75090.0 ;
      RECT  25620.0 76435.0 26325.0 75090.0 ;
      RECT  25620.0 76435.0 26325.0 77780.0 ;
      RECT  25620.0 79125.0 26325.0 77780.0 ;
      RECT  25620.0 79125.0 26325.0 80470.0 ;
      RECT  25620.0 81815.0 26325.0 80470.0 ;
      RECT  25620.0 81815.0 26325.0 83160.0 ;
      RECT  25620.0 84505.0 26325.0 83160.0 ;
      RECT  25620.0 84505.0 26325.0 85850.0 ;
      RECT  25620.0 87195.0 26325.0 85850.0 ;
      RECT  25620.0 87195.0 26325.0 88540.0 ;
      RECT  25620.0 89885.0 26325.0 88540.0 ;
      RECT  25620.0 89885.0 26325.0 91230.0 ;
      RECT  25620.0 92575.0 26325.0 91230.0 ;
      RECT  25620.0 92575.0 26325.0 93920.0 ;
      RECT  25620.0 95265.0 26325.0 93920.0 ;
      RECT  25620.0 95265.0 26325.0 96610.0 ;
      RECT  25620.0 97955.0 26325.0 96610.0 ;
      RECT  25620.0 97955.0 26325.0 99300.0 ;
      RECT  25620.0 100645.0 26325.0 99300.0 ;
      RECT  25620.0 100645.0 26325.0 101990.0 ;
      RECT  25620.0 103335.0 26325.0 101990.0 ;
      RECT  25620.0 103335.0 26325.0 104680.0 ;
      RECT  25620.0 106025.0 26325.0 104680.0 ;
      RECT  25620.0 106025.0 26325.0 107370.0 ;
      RECT  25620.0 108715.0 26325.0 107370.0 ;
      RECT  25620.0 108715.0 26325.0 110060.0 ;
      RECT  25620.0 111405.0 26325.0 110060.0 ;
      RECT  25620.0 111405.0 26325.0 112750.0 ;
      RECT  25620.0 114095.0 26325.0 112750.0 ;
      RECT  26325.0 28015.0 27030.0 29360.0 ;
      RECT  26325.0 30705.0 27030.0 29360.0 ;
      RECT  26325.0 30705.0 27030.0 32050.0 ;
      RECT  26325.0 33395.0 27030.0 32050.0 ;
      RECT  26325.0 33395.0 27030.0 34740.0 ;
      RECT  26325.0 36085.0 27030.0 34740.0 ;
      RECT  26325.0 36085.0 27030.0 37430.0 ;
      RECT  26325.0 38775.0 27030.0 37430.0 ;
      RECT  26325.0 38775.0 27030.0 40120.0 ;
      RECT  26325.0 41465.0 27030.0 40120.0 ;
      RECT  26325.0 41465.0 27030.0 42810.0 ;
      RECT  26325.0 44155.0 27030.0 42810.0 ;
      RECT  26325.0 44155.0 27030.0 45500.0 ;
      RECT  26325.0 46845.0 27030.0 45500.0 ;
      RECT  26325.0 46845.0 27030.0 48190.0 ;
      RECT  26325.0 49535.0 27030.0 48190.0 ;
      RECT  26325.0 49535.0 27030.0 50880.0 ;
      RECT  26325.0 52225.0 27030.0 50880.0 ;
      RECT  26325.0 52225.0 27030.0 53570.0 ;
      RECT  26325.0 54915.0 27030.0 53570.0 ;
      RECT  26325.0 54915.0 27030.0 56260.0 ;
      RECT  26325.0 57605.0 27030.0 56260.0 ;
      RECT  26325.0 57605.0 27030.0 58950.0 ;
      RECT  26325.0 60295.0 27030.0 58950.0 ;
      RECT  26325.0 60295.0 27030.0 61640.0 ;
      RECT  26325.0 62985.0 27030.0 61640.0 ;
      RECT  26325.0 62985.0 27030.0 64330.0 ;
      RECT  26325.0 65675.0 27030.0 64330.0 ;
      RECT  26325.0 65675.0 27030.0 67020.0 ;
      RECT  26325.0 68365.0 27030.0 67020.0 ;
      RECT  26325.0 68365.0 27030.0 69710.0 ;
      RECT  26325.0 71055.0 27030.0 69710.0 ;
      RECT  26325.0 71055.0 27030.0 72400.0 ;
      RECT  26325.0 73745.0 27030.0 72400.0 ;
      RECT  26325.0 73745.0 27030.0 75090.0 ;
      RECT  26325.0 76435.0 27030.0 75090.0 ;
      RECT  26325.0 76435.0 27030.0 77780.0 ;
      RECT  26325.0 79125.0 27030.0 77780.0 ;
      RECT  26325.0 79125.0 27030.0 80470.0 ;
      RECT  26325.0 81815.0 27030.0 80470.0 ;
      RECT  26325.0 81815.0 27030.0 83160.0 ;
      RECT  26325.0 84505.0 27030.0 83160.0 ;
      RECT  26325.0 84505.0 27030.0 85850.0 ;
      RECT  26325.0 87195.0 27030.0 85850.0 ;
      RECT  26325.0 87195.0 27030.0 88540.0 ;
      RECT  26325.0 89885.0 27030.0 88540.0 ;
      RECT  26325.0 89885.0 27030.0 91230.0 ;
      RECT  26325.0 92575.0 27030.0 91230.0 ;
      RECT  26325.0 92575.0 27030.0 93920.0 ;
      RECT  26325.0 95265.0 27030.0 93920.0 ;
      RECT  26325.0 95265.0 27030.0 96610.0 ;
      RECT  26325.0 97955.0 27030.0 96610.0 ;
      RECT  26325.0 97955.0 27030.0 99300.0 ;
      RECT  26325.0 100645.0 27030.0 99300.0 ;
      RECT  26325.0 100645.0 27030.0 101990.0 ;
      RECT  26325.0 103335.0 27030.0 101990.0 ;
      RECT  26325.0 103335.0 27030.0 104680.0 ;
      RECT  26325.0 106025.0 27030.0 104680.0 ;
      RECT  26325.0 106025.0 27030.0 107370.0 ;
      RECT  26325.0 108715.0 27030.0 107370.0 ;
      RECT  26325.0 108715.0 27030.0 110060.0 ;
      RECT  26325.0 111405.0 27030.0 110060.0 ;
      RECT  26325.0 111405.0 27030.0 112750.0 ;
      RECT  26325.0 114095.0 27030.0 112750.0 ;
      RECT  27030.0 28015.0 27735.0 29360.0 ;
      RECT  27030.0 30705.0 27735.0 29360.0 ;
      RECT  27030.0 30705.0 27735.0 32050.0 ;
      RECT  27030.0 33395.0 27735.0 32050.0 ;
      RECT  27030.0 33395.0 27735.0 34740.0 ;
      RECT  27030.0 36085.0 27735.0 34740.0 ;
      RECT  27030.0 36085.0 27735.0 37430.0 ;
      RECT  27030.0 38775.0 27735.0 37430.0 ;
      RECT  27030.0 38775.0 27735.0 40120.0 ;
      RECT  27030.0 41465.0 27735.0 40120.0 ;
      RECT  27030.0 41465.0 27735.0 42810.0 ;
      RECT  27030.0 44155.0 27735.0 42810.0 ;
      RECT  27030.0 44155.0 27735.0 45500.0 ;
      RECT  27030.0 46845.0 27735.0 45500.0 ;
      RECT  27030.0 46845.0 27735.0 48190.0 ;
      RECT  27030.0 49535.0 27735.0 48190.0 ;
      RECT  27030.0 49535.0 27735.0 50880.0 ;
      RECT  27030.0 52225.0 27735.0 50880.0 ;
      RECT  27030.0 52225.0 27735.0 53570.0 ;
      RECT  27030.0 54915.0 27735.0 53570.0 ;
      RECT  27030.0 54915.0 27735.0 56260.0 ;
      RECT  27030.0 57605.0 27735.0 56260.0 ;
      RECT  27030.0 57605.0 27735.0 58950.0 ;
      RECT  27030.0 60295.0 27735.0 58950.0 ;
      RECT  27030.0 60295.0 27735.0 61640.0 ;
      RECT  27030.0 62985.0 27735.0 61640.0 ;
      RECT  27030.0 62985.0 27735.0 64330.0 ;
      RECT  27030.0 65675.0 27735.0 64330.0 ;
      RECT  27030.0 65675.0 27735.0 67020.0 ;
      RECT  27030.0 68365.0 27735.0 67020.0 ;
      RECT  27030.0 68365.0 27735.0 69710.0 ;
      RECT  27030.0 71055.0 27735.0 69710.0 ;
      RECT  27030.0 71055.0 27735.0 72400.0 ;
      RECT  27030.0 73745.0 27735.0 72400.0 ;
      RECT  27030.0 73745.0 27735.0 75090.0 ;
      RECT  27030.0 76435.0 27735.0 75090.0 ;
      RECT  27030.0 76435.0 27735.0 77780.0 ;
      RECT  27030.0 79125.0 27735.0 77780.0 ;
      RECT  27030.0 79125.0 27735.0 80470.0 ;
      RECT  27030.0 81815.0 27735.0 80470.0 ;
      RECT  27030.0 81815.0 27735.0 83160.0 ;
      RECT  27030.0 84505.0 27735.0 83160.0 ;
      RECT  27030.0 84505.0 27735.0 85850.0 ;
      RECT  27030.0 87195.0 27735.0 85850.0 ;
      RECT  27030.0 87195.0 27735.0 88540.0 ;
      RECT  27030.0 89885.0 27735.0 88540.0 ;
      RECT  27030.0 89885.0 27735.0 91230.0 ;
      RECT  27030.0 92575.0 27735.0 91230.0 ;
      RECT  27030.0 92575.0 27735.0 93920.0 ;
      RECT  27030.0 95265.0 27735.0 93920.0 ;
      RECT  27030.0 95265.0 27735.0 96610.0 ;
      RECT  27030.0 97955.0 27735.0 96610.0 ;
      RECT  27030.0 97955.0 27735.0 99300.0 ;
      RECT  27030.0 100645.0 27735.0 99300.0 ;
      RECT  27030.0 100645.0 27735.0 101990.0 ;
      RECT  27030.0 103335.0 27735.0 101990.0 ;
      RECT  27030.0 103335.0 27735.0 104680.0 ;
      RECT  27030.0 106025.0 27735.0 104680.0 ;
      RECT  27030.0 106025.0 27735.0 107370.0 ;
      RECT  27030.0 108715.0 27735.0 107370.0 ;
      RECT  27030.0 108715.0 27735.0 110060.0 ;
      RECT  27030.0 111405.0 27735.0 110060.0 ;
      RECT  27030.0 111405.0 27735.0 112750.0 ;
      RECT  27030.0 114095.0 27735.0 112750.0 ;
      RECT  27735.0 28015.0 28440.0 29360.0 ;
      RECT  27735.0 30705.0 28440.0 29360.0 ;
      RECT  27735.0 30705.0 28440.0 32050.0 ;
      RECT  27735.0 33395.0 28440.0 32050.0 ;
      RECT  27735.0 33395.0 28440.0 34740.0 ;
      RECT  27735.0 36085.0 28440.0 34740.0 ;
      RECT  27735.0 36085.0 28440.0 37430.0 ;
      RECT  27735.0 38775.0 28440.0 37430.0 ;
      RECT  27735.0 38775.0 28440.0 40120.0 ;
      RECT  27735.0 41465.0 28440.0 40120.0 ;
      RECT  27735.0 41465.0 28440.0 42810.0 ;
      RECT  27735.0 44155.0 28440.0 42810.0 ;
      RECT  27735.0 44155.0 28440.0 45500.0 ;
      RECT  27735.0 46845.0 28440.0 45500.0 ;
      RECT  27735.0 46845.0 28440.0 48190.0 ;
      RECT  27735.0 49535.0 28440.0 48190.0 ;
      RECT  27735.0 49535.0 28440.0 50880.0 ;
      RECT  27735.0 52225.0 28440.0 50880.0 ;
      RECT  27735.0 52225.0 28440.0 53570.0 ;
      RECT  27735.0 54915.0 28440.0 53570.0 ;
      RECT  27735.0 54915.0 28440.0 56260.0 ;
      RECT  27735.0 57605.0 28440.0 56260.0 ;
      RECT  27735.0 57605.0 28440.0 58950.0 ;
      RECT  27735.0 60295.0 28440.0 58950.0 ;
      RECT  27735.0 60295.0 28440.0 61640.0 ;
      RECT  27735.0 62985.0 28440.0 61640.0 ;
      RECT  27735.0 62985.0 28440.0 64330.0 ;
      RECT  27735.0 65675.0 28440.0 64330.0 ;
      RECT  27735.0 65675.0 28440.0 67020.0 ;
      RECT  27735.0 68365.0 28440.0 67020.0 ;
      RECT  27735.0 68365.0 28440.0 69710.0 ;
      RECT  27735.0 71055.0 28440.0 69710.0 ;
      RECT  27735.0 71055.0 28440.0 72400.0 ;
      RECT  27735.0 73745.0 28440.0 72400.0 ;
      RECT  27735.0 73745.0 28440.0 75090.0 ;
      RECT  27735.0 76435.0 28440.0 75090.0 ;
      RECT  27735.0 76435.0 28440.0 77780.0 ;
      RECT  27735.0 79125.0 28440.0 77780.0 ;
      RECT  27735.0 79125.0 28440.0 80470.0 ;
      RECT  27735.0 81815.0 28440.0 80470.0 ;
      RECT  27735.0 81815.0 28440.0 83160.0 ;
      RECT  27735.0 84505.0 28440.0 83160.0 ;
      RECT  27735.0 84505.0 28440.0 85850.0 ;
      RECT  27735.0 87195.0 28440.0 85850.0 ;
      RECT  27735.0 87195.0 28440.0 88540.0 ;
      RECT  27735.0 89885.0 28440.0 88540.0 ;
      RECT  27735.0 89885.0 28440.0 91230.0 ;
      RECT  27735.0 92575.0 28440.0 91230.0 ;
      RECT  27735.0 92575.0 28440.0 93920.0 ;
      RECT  27735.0 95265.0 28440.0 93920.0 ;
      RECT  27735.0 95265.0 28440.0 96610.0 ;
      RECT  27735.0 97955.0 28440.0 96610.0 ;
      RECT  27735.0 97955.0 28440.0 99300.0 ;
      RECT  27735.0 100645.0 28440.0 99300.0 ;
      RECT  27735.0 100645.0 28440.0 101990.0 ;
      RECT  27735.0 103335.0 28440.0 101990.0 ;
      RECT  27735.0 103335.0 28440.0 104680.0 ;
      RECT  27735.0 106025.0 28440.0 104680.0 ;
      RECT  27735.0 106025.0 28440.0 107370.0 ;
      RECT  27735.0 108715.0 28440.0 107370.0 ;
      RECT  27735.0 108715.0 28440.0 110060.0 ;
      RECT  27735.0 111405.0 28440.0 110060.0 ;
      RECT  27735.0 111405.0 28440.0 112750.0 ;
      RECT  27735.0 114095.0 28440.0 112750.0 ;
      RECT  28440.0 28015.0 29145.0 29360.0 ;
      RECT  28440.0 30705.0 29145.0 29360.0 ;
      RECT  28440.0 30705.0 29145.0 32050.0 ;
      RECT  28440.0 33395.0 29145.0 32050.0 ;
      RECT  28440.0 33395.0 29145.0 34740.0 ;
      RECT  28440.0 36085.0 29145.0 34740.0 ;
      RECT  28440.0 36085.0 29145.0 37430.0 ;
      RECT  28440.0 38775.0 29145.0 37430.0 ;
      RECT  28440.0 38775.0 29145.0 40120.0 ;
      RECT  28440.0 41465.0 29145.0 40120.0 ;
      RECT  28440.0 41465.0 29145.0 42810.0 ;
      RECT  28440.0 44155.0 29145.0 42810.0 ;
      RECT  28440.0 44155.0 29145.0 45500.0 ;
      RECT  28440.0 46845.0 29145.0 45500.0 ;
      RECT  28440.0 46845.0 29145.0 48190.0 ;
      RECT  28440.0 49535.0 29145.0 48190.0 ;
      RECT  28440.0 49535.0 29145.0 50880.0 ;
      RECT  28440.0 52225.0 29145.0 50880.0 ;
      RECT  28440.0 52225.0 29145.0 53570.0 ;
      RECT  28440.0 54915.0 29145.0 53570.0 ;
      RECT  28440.0 54915.0 29145.0 56260.0 ;
      RECT  28440.0 57605.0 29145.0 56260.0 ;
      RECT  28440.0 57605.0 29145.0 58950.0 ;
      RECT  28440.0 60295.0 29145.0 58950.0 ;
      RECT  28440.0 60295.0 29145.0 61640.0 ;
      RECT  28440.0 62985.0 29145.0 61640.0 ;
      RECT  28440.0 62985.0 29145.0 64330.0 ;
      RECT  28440.0 65675.0 29145.0 64330.0 ;
      RECT  28440.0 65675.0 29145.0 67020.0 ;
      RECT  28440.0 68365.0 29145.0 67020.0 ;
      RECT  28440.0 68365.0 29145.0 69710.0 ;
      RECT  28440.0 71055.0 29145.0 69710.0 ;
      RECT  28440.0 71055.0 29145.0 72400.0 ;
      RECT  28440.0 73745.0 29145.0 72400.0 ;
      RECT  28440.0 73745.0 29145.0 75090.0 ;
      RECT  28440.0 76435.0 29145.0 75090.0 ;
      RECT  28440.0 76435.0 29145.0 77780.0 ;
      RECT  28440.0 79125.0 29145.0 77780.0 ;
      RECT  28440.0 79125.0 29145.0 80470.0 ;
      RECT  28440.0 81815.0 29145.0 80470.0 ;
      RECT  28440.0 81815.0 29145.0 83160.0 ;
      RECT  28440.0 84505.0 29145.0 83160.0 ;
      RECT  28440.0 84505.0 29145.0 85850.0 ;
      RECT  28440.0 87195.0 29145.0 85850.0 ;
      RECT  28440.0 87195.0 29145.0 88540.0 ;
      RECT  28440.0 89885.0 29145.0 88540.0 ;
      RECT  28440.0 89885.0 29145.0 91230.0 ;
      RECT  28440.0 92575.0 29145.0 91230.0 ;
      RECT  28440.0 92575.0 29145.0 93920.0 ;
      RECT  28440.0 95265.0 29145.0 93920.0 ;
      RECT  28440.0 95265.0 29145.0 96610.0 ;
      RECT  28440.0 97955.0 29145.0 96610.0 ;
      RECT  28440.0 97955.0 29145.0 99300.0 ;
      RECT  28440.0 100645.0 29145.0 99300.0 ;
      RECT  28440.0 100645.0 29145.0 101990.0 ;
      RECT  28440.0 103335.0 29145.0 101990.0 ;
      RECT  28440.0 103335.0 29145.0 104680.0 ;
      RECT  28440.0 106025.0 29145.0 104680.0 ;
      RECT  28440.0 106025.0 29145.0 107370.0 ;
      RECT  28440.0 108715.0 29145.0 107370.0 ;
      RECT  28440.0 108715.0 29145.0 110060.0 ;
      RECT  28440.0 111405.0 29145.0 110060.0 ;
      RECT  28440.0 111405.0 29145.0 112750.0 ;
      RECT  28440.0 114095.0 29145.0 112750.0 ;
      RECT  29145.0 28015.0 29850.0 29360.0 ;
      RECT  29145.0 30705.0 29850.0 29360.0 ;
      RECT  29145.0 30705.0 29850.0 32050.0 ;
      RECT  29145.0 33395.0 29850.0 32050.0 ;
      RECT  29145.0 33395.0 29850.0 34740.0 ;
      RECT  29145.0 36085.0 29850.0 34740.0 ;
      RECT  29145.0 36085.0 29850.0 37430.0 ;
      RECT  29145.0 38775.0 29850.0 37430.0 ;
      RECT  29145.0 38775.0 29850.0 40120.0 ;
      RECT  29145.0 41465.0 29850.0 40120.0 ;
      RECT  29145.0 41465.0 29850.0 42810.0 ;
      RECT  29145.0 44155.0 29850.0 42810.0 ;
      RECT  29145.0 44155.0 29850.0 45500.0 ;
      RECT  29145.0 46845.0 29850.0 45500.0 ;
      RECT  29145.0 46845.0 29850.0 48190.0 ;
      RECT  29145.0 49535.0 29850.0 48190.0 ;
      RECT  29145.0 49535.0 29850.0 50880.0 ;
      RECT  29145.0 52225.0 29850.0 50880.0 ;
      RECT  29145.0 52225.0 29850.0 53570.0 ;
      RECT  29145.0 54915.0 29850.0 53570.0 ;
      RECT  29145.0 54915.0 29850.0 56260.0 ;
      RECT  29145.0 57605.0 29850.0 56260.0 ;
      RECT  29145.0 57605.0 29850.0 58950.0 ;
      RECT  29145.0 60295.0 29850.0 58950.0 ;
      RECT  29145.0 60295.0 29850.0 61640.0 ;
      RECT  29145.0 62985.0 29850.0 61640.0 ;
      RECT  29145.0 62985.0 29850.0 64330.0 ;
      RECT  29145.0 65675.0 29850.0 64330.0 ;
      RECT  29145.0 65675.0 29850.0 67020.0 ;
      RECT  29145.0 68365.0 29850.0 67020.0 ;
      RECT  29145.0 68365.0 29850.0 69710.0 ;
      RECT  29145.0 71055.0 29850.0 69710.0 ;
      RECT  29145.0 71055.0 29850.0 72400.0 ;
      RECT  29145.0 73745.0 29850.0 72400.0 ;
      RECT  29145.0 73745.0 29850.0 75090.0 ;
      RECT  29145.0 76435.0 29850.0 75090.0 ;
      RECT  29145.0 76435.0 29850.0 77780.0 ;
      RECT  29145.0 79125.0 29850.0 77780.0 ;
      RECT  29145.0 79125.0 29850.0 80470.0 ;
      RECT  29145.0 81815.0 29850.0 80470.0 ;
      RECT  29145.0 81815.0 29850.0 83160.0 ;
      RECT  29145.0 84505.0 29850.0 83160.0 ;
      RECT  29145.0 84505.0 29850.0 85850.0 ;
      RECT  29145.0 87195.0 29850.0 85850.0 ;
      RECT  29145.0 87195.0 29850.0 88540.0 ;
      RECT  29145.0 89885.0 29850.0 88540.0 ;
      RECT  29145.0 89885.0 29850.0 91230.0 ;
      RECT  29145.0 92575.0 29850.0 91230.0 ;
      RECT  29145.0 92575.0 29850.0 93920.0 ;
      RECT  29145.0 95265.0 29850.0 93920.0 ;
      RECT  29145.0 95265.0 29850.0 96610.0 ;
      RECT  29145.0 97955.0 29850.0 96610.0 ;
      RECT  29145.0 97955.0 29850.0 99300.0 ;
      RECT  29145.0 100645.0 29850.0 99300.0 ;
      RECT  29145.0 100645.0 29850.0 101990.0 ;
      RECT  29145.0 103335.0 29850.0 101990.0 ;
      RECT  29145.0 103335.0 29850.0 104680.0 ;
      RECT  29145.0 106025.0 29850.0 104680.0 ;
      RECT  29145.0 106025.0 29850.0 107370.0 ;
      RECT  29145.0 108715.0 29850.0 107370.0 ;
      RECT  29145.0 108715.0 29850.0 110060.0 ;
      RECT  29145.0 111405.0 29850.0 110060.0 ;
      RECT  29145.0 111405.0 29850.0 112750.0 ;
      RECT  29145.0 114095.0 29850.0 112750.0 ;
      RECT  29850.0 28015.0 30555.0 29360.0 ;
      RECT  29850.0 30705.0 30555.0 29360.0 ;
      RECT  29850.0 30705.0 30555.0 32050.0 ;
      RECT  29850.0 33395.0 30555.0 32050.0 ;
      RECT  29850.0 33395.0 30555.0 34740.0 ;
      RECT  29850.0 36085.0 30555.0 34740.0 ;
      RECT  29850.0 36085.0 30555.0 37430.0 ;
      RECT  29850.0 38775.0 30555.0 37430.0 ;
      RECT  29850.0 38775.0 30555.0 40120.0 ;
      RECT  29850.0 41465.0 30555.0 40120.0 ;
      RECT  29850.0 41465.0 30555.0 42810.0 ;
      RECT  29850.0 44155.0 30555.0 42810.0 ;
      RECT  29850.0 44155.0 30555.0 45500.0 ;
      RECT  29850.0 46845.0 30555.0 45500.0 ;
      RECT  29850.0 46845.0 30555.0 48190.0 ;
      RECT  29850.0 49535.0 30555.0 48190.0 ;
      RECT  29850.0 49535.0 30555.0 50880.0 ;
      RECT  29850.0 52225.0 30555.0 50880.0 ;
      RECT  29850.0 52225.0 30555.0 53570.0 ;
      RECT  29850.0 54915.0 30555.0 53570.0 ;
      RECT  29850.0 54915.0 30555.0 56260.0 ;
      RECT  29850.0 57605.0 30555.0 56260.0 ;
      RECT  29850.0 57605.0 30555.0 58950.0 ;
      RECT  29850.0 60295.0 30555.0 58950.0 ;
      RECT  29850.0 60295.0 30555.0 61640.0 ;
      RECT  29850.0 62985.0 30555.0 61640.0 ;
      RECT  29850.0 62985.0 30555.0 64330.0 ;
      RECT  29850.0 65675.0 30555.0 64330.0 ;
      RECT  29850.0 65675.0 30555.0 67020.0 ;
      RECT  29850.0 68365.0 30555.0 67020.0 ;
      RECT  29850.0 68365.0 30555.0 69710.0 ;
      RECT  29850.0 71055.0 30555.0 69710.0 ;
      RECT  29850.0 71055.0 30555.0 72400.0 ;
      RECT  29850.0 73745.0 30555.0 72400.0 ;
      RECT  29850.0 73745.0 30555.0 75090.0 ;
      RECT  29850.0 76435.0 30555.0 75090.0 ;
      RECT  29850.0 76435.0 30555.0 77780.0 ;
      RECT  29850.0 79125.0 30555.0 77780.0 ;
      RECT  29850.0 79125.0 30555.0 80470.0 ;
      RECT  29850.0 81815.0 30555.0 80470.0 ;
      RECT  29850.0 81815.0 30555.0 83160.0 ;
      RECT  29850.0 84505.0 30555.0 83160.0 ;
      RECT  29850.0 84505.0 30555.0 85850.0 ;
      RECT  29850.0 87195.0 30555.0 85850.0 ;
      RECT  29850.0 87195.0 30555.0 88540.0 ;
      RECT  29850.0 89885.0 30555.0 88540.0 ;
      RECT  29850.0 89885.0 30555.0 91230.0 ;
      RECT  29850.0 92575.0 30555.0 91230.0 ;
      RECT  29850.0 92575.0 30555.0 93920.0 ;
      RECT  29850.0 95265.0 30555.0 93920.0 ;
      RECT  29850.0 95265.0 30555.0 96610.0 ;
      RECT  29850.0 97955.0 30555.0 96610.0 ;
      RECT  29850.0 97955.0 30555.0 99300.0 ;
      RECT  29850.0 100645.0 30555.0 99300.0 ;
      RECT  29850.0 100645.0 30555.0 101990.0 ;
      RECT  29850.0 103335.0 30555.0 101990.0 ;
      RECT  29850.0 103335.0 30555.0 104680.0 ;
      RECT  29850.0 106025.0 30555.0 104680.0 ;
      RECT  29850.0 106025.0 30555.0 107370.0 ;
      RECT  29850.0 108715.0 30555.0 107370.0 ;
      RECT  29850.0 108715.0 30555.0 110060.0 ;
      RECT  29850.0 111405.0 30555.0 110060.0 ;
      RECT  29850.0 111405.0 30555.0 112750.0 ;
      RECT  29850.0 114095.0 30555.0 112750.0 ;
      RECT  30555.0 28015.0 31260.0 29360.0 ;
      RECT  30555.0 30705.0 31260.0 29360.0 ;
      RECT  30555.0 30705.0 31260.0 32050.0 ;
      RECT  30555.0 33395.0 31260.0 32050.0 ;
      RECT  30555.0 33395.0 31260.0 34740.0 ;
      RECT  30555.0 36085.0 31260.0 34740.0 ;
      RECT  30555.0 36085.0 31260.0 37430.0 ;
      RECT  30555.0 38775.0 31260.0 37430.0 ;
      RECT  30555.0 38775.0 31260.0 40120.0 ;
      RECT  30555.0 41465.0 31260.0 40120.0 ;
      RECT  30555.0 41465.0 31260.0 42810.0 ;
      RECT  30555.0 44155.0 31260.0 42810.0 ;
      RECT  30555.0 44155.0 31260.0 45500.0 ;
      RECT  30555.0 46845.0 31260.0 45500.0 ;
      RECT  30555.0 46845.0 31260.0 48190.0 ;
      RECT  30555.0 49535.0 31260.0 48190.0 ;
      RECT  30555.0 49535.0 31260.0 50880.0 ;
      RECT  30555.0 52225.0 31260.0 50880.0 ;
      RECT  30555.0 52225.0 31260.0 53570.0 ;
      RECT  30555.0 54915.0 31260.0 53570.0 ;
      RECT  30555.0 54915.0 31260.0 56260.0 ;
      RECT  30555.0 57605.0 31260.0 56260.0 ;
      RECT  30555.0 57605.0 31260.0 58950.0 ;
      RECT  30555.0 60295.0 31260.0 58950.0 ;
      RECT  30555.0 60295.0 31260.0 61640.0 ;
      RECT  30555.0 62985.0 31260.0 61640.0 ;
      RECT  30555.0 62985.0 31260.0 64330.0 ;
      RECT  30555.0 65675.0 31260.0 64330.0 ;
      RECT  30555.0 65675.0 31260.0 67020.0 ;
      RECT  30555.0 68365.0 31260.0 67020.0 ;
      RECT  30555.0 68365.0 31260.0 69710.0 ;
      RECT  30555.0 71055.0 31260.0 69710.0 ;
      RECT  30555.0 71055.0 31260.0 72400.0 ;
      RECT  30555.0 73745.0 31260.0 72400.0 ;
      RECT  30555.0 73745.0 31260.0 75090.0 ;
      RECT  30555.0 76435.0 31260.0 75090.0 ;
      RECT  30555.0 76435.0 31260.0 77780.0 ;
      RECT  30555.0 79125.0 31260.0 77780.0 ;
      RECT  30555.0 79125.0 31260.0 80470.0 ;
      RECT  30555.0 81815.0 31260.0 80470.0 ;
      RECT  30555.0 81815.0 31260.0 83160.0 ;
      RECT  30555.0 84505.0 31260.0 83160.0 ;
      RECT  30555.0 84505.0 31260.0 85850.0 ;
      RECT  30555.0 87195.0 31260.0 85850.0 ;
      RECT  30555.0 87195.0 31260.0 88540.0 ;
      RECT  30555.0 89885.0 31260.0 88540.0 ;
      RECT  30555.0 89885.0 31260.0 91230.0 ;
      RECT  30555.0 92575.0 31260.0 91230.0 ;
      RECT  30555.0 92575.0 31260.0 93920.0 ;
      RECT  30555.0 95265.0 31260.0 93920.0 ;
      RECT  30555.0 95265.0 31260.0 96610.0 ;
      RECT  30555.0 97955.0 31260.0 96610.0 ;
      RECT  30555.0 97955.0 31260.0 99300.0 ;
      RECT  30555.0 100645.0 31260.0 99300.0 ;
      RECT  30555.0 100645.0 31260.0 101990.0 ;
      RECT  30555.0 103335.0 31260.0 101990.0 ;
      RECT  30555.0 103335.0 31260.0 104680.0 ;
      RECT  30555.0 106025.0 31260.0 104680.0 ;
      RECT  30555.0 106025.0 31260.0 107370.0 ;
      RECT  30555.0 108715.0 31260.0 107370.0 ;
      RECT  30555.0 108715.0 31260.0 110060.0 ;
      RECT  30555.0 111405.0 31260.0 110060.0 ;
      RECT  30555.0 111405.0 31260.0 112750.0 ;
      RECT  30555.0 114095.0 31260.0 112750.0 ;
      RECT  31260.0 28015.0 31965.0 29360.0 ;
      RECT  31260.0 30705.0 31965.0 29360.0 ;
      RECT  31260.0 30705.0 31965.0 32050.0 ;
      RECT  31260.0 33395.0 31965.0 32050.0 ;
      RECT  31260.0 33395.0 31965.0 34740.0 ;
      RECT  31260.0 36085.0 31965.0 34740.0 ;
      RECT  31260.0 36085.0 31965.0 37430.0 ;
      RECT  31260.0 38775.0 31965.0 37430.0 ;
      RECT  31260.0 38775.0 31965.0 40120.0 ;
      RECT  31260.0 41465.0 31965.0 40120.0 ;
      RECT  31260.0 41465.0 31965.0 42810.0 ;
      RECT  31260.0 44155.0 31965.0 42810.0 ;
      RECT  31260.0 44155.0 31965.0 45500.0 ;
      RECT  31260.0 46845.0 31965.0 45500.0 ;
      RECT  31260.0 46845.0 31965.0 48190.0 ;
      RECT  31260.0 49535.0 31965.0 48190.0 ;
      RECT  31260.0 49535.0 31965.0 50880.0 ;
      RECT  31260.0 52225.0 31965.0 50880.0 ;
      RECT  31260.0 52225.0 31965.0 53570.0 ;
      RECT  31260.0 54915.0 31965.0 53570.0 ;
      RECT  31260.0 54915.0 31965.0 56260.0 ;
      RECT  31260.0 57605.0 31965.0 56260.0 ;
      RECT  31260.0 57605.0 31965.0 58950.0 ;
      RECT  31260.0 60295.0 31965.0 58950.0 ;
      RECT  31260.0 60295.0 31965.0 61640.0 ;
      RECT  31260.0 62985.0 31965.0 61640.0 ;
      RECT  31260.0 62985.0 31965.0 64330.0 ;
      RECT  31260.0 65675.0 31965.0 64330.0 ;
      RECT  31260.0 65675.0 31965.0 67020.0 ;
      RECT  31260.0 68365.0 31965.0 67020.0 ;
      RECT  31260.0 68365.0 31965.0 69710.0 ;
      RECT  31260.0 71055.0 31965.0 69710.0 ;
      RECT  31260.0 71055.0 31965.0 72400.0 ;
      RECT  31260.0 73745.0 31965.0 72400.0 ;
      RECT  31260.0 73745.0 31965.0 75090.0 ;
      RECT  31260.0 76435.0 31965.0 75090.0 ;
      RECT  31260.0 76435.0 31965.0 77780.0 ;
      RECT  31260.0 79125.0 31965.0 77780.0 ;
      RECT  31260.0 79125.0 31965.0 80470.0 ;
      RECT  31260.0 81815.0 31965.0 80470.0 ;
      RECT  31260.0 81815.0 31965.0 83160.0 ;
      RECT  31260.0 84505.0 31965.0 83160.0 ;
      RECT  31260.0 84505.0 31965.0 85850.0 ;
      RECT  31260.0 87195.0 31965.0 85850.0 ;
      RECT  31260.0 87195.0 31965.0 88540.0 ;
      RECT  31260.0 89885.0 31965.0 88540.0 ;
      RECT  31260.0 89885.0 31965.0 91230.0 ;
      RECT  31260.0 92575.0 31965.0 91230.0 ;
      RECT  31260.0 92575.0 31965.0 93920.0 ;
      RECT  31260.0 95265.0 31965.0 93920.0 ;
      RECT  31260.0 95265.0 31965.0 96610.0 ;
      RECT  31260.0 97955.0 31965.0 96610.0 ;
      RECT  31260.0 97955.0 31965.0 99300.0 ;
      RECT  31260.0 100645.0 31965.0 99300.0 ;
      RECT  31260.0 100645.0 31965.0 101990.0 ;
      RECT  31260.0 103335.0 31965.0 101990.0 ;
      RECT  31260.0 103335.0 31965.0 104680.0 ;
      RECT  31260.0 106025.0 31965.0 104680.0 ;
      RECT  31260.0 106025.0 31965.0 107370.0 ;
      RECT  31260.0 108715.0 31965.0 107370.0 ;
      RECT  31260.0 108715.0 31965.0 110060.0 ;
      RECT  31260.0 111405.0 31965.0 110060.0 ;
      RECT  31260.0 111405.0 31965.0 112750.0 ;
      RECT  31260.0 114095.0 31965.0 112750.0 ;
      RECT  31965.0 28015.0 32670.0 29360.0 ;
      RECT  31965.0 30705.0 32670.0 29360.0 ;
      RECT  31965.0 30705.0 32670.0 32050.0 ;
      RECT  31965.0 33395.0 32670.0 32050.0 ;
      RECT  31965.0 33395.0 32670.0 34740.0 ;
      RECT  31965.0 36085.0 32670.0 34740.0 ;
      RECT  31965.0 36085.0 32670.0 37430.0 ;
      RECT  31965.0 38775.0 32670.0 37430.0 ;
      RECT  31965.0 38775.0 32670.0 40120.0 ;
      RECT  31965.0 41465.0 32670.0 40120.0 ;
      RECT  31965.0 41465.0 32670.0 42810.0 ;
      RECT  31965.0 44155.0 32670.0 42810.0 ;
      RECT  31965.0 44155.0 32670.0 45500.0 ;
      RECT  31965.0 46845.0 32670.0 45500.0 ;
      RECT  31965.0 46845.0 32670.0 48190.0 ;
      RECT  31965.0 49535.0 32670.0 48190.0 ;
      RECT  31965.0 49535.0 32670.0 50880.0 ;
      RECT  31965.0 52225.0 32670.0 50880.0 ;
      RECT  31965.0 52225.0 32670.0 53570.0 ;
      RECT  31965.0 54915.0 32670.0 53570.0 ;
      RECT  31965.0 54915.0 32670.0 56260.0 ;
      RECT  31965.0 57605.0 32670.0 56260.0 ;
      RECT  31965.0 57605.0 32670.0 58950.0 ;
      RECT  31965.0 60295.0 32670.0 58950.0 ;
      RECT  31965.0 60295.0 32670.0 61640.0 ;
      RECT  31965.0 62985.0 32670.0 61640.0 ;
      RECT  31965.0 62985.0 32670.0 64330.0 ;
      RECT  31965.0 65675.0 32670.0 64330.0 ;
      RECT  31965.0 65675.0 32670.0 67020.0 ;
      RECT  31965.0 68365.0 32670.0 67020.0 ;
      RECT  31965.0 68365.0 32670.0 69710.0 ;
      RECT  31965.0 71055.0 32670.0 69710.0 ;
      RECT  31965.0 71055.0 32670.0 72400.0 ;
      RECT  31965.0 73745.0 32670.0 72400.0 ;
      RECT  31965.0 73745.0 32670.0 75090.0 ;
      RECT  31965.0 76435.0 32670.0 75090.0 ;
      RECT  31965.0 76435.0 32670.0 77780.0 ;
      RECT  31965.0 79125.0 32670.0 77780.0 ;
      RECT  31965.0 79125.0 32670.0 80470.0 ;
      RECT  31965.0 81815.0 32670.0 80470.0 ;
      RECT  31965.0 81815.0 32670.0 83160.0 ;
      RECT  31965.0 84505.0 32670.0 83160.0 ;
      RECT  31965.0 84505.0 32670.0 85850.0 ;
      RECT  31965.0 87195.0 32670.0 85850.0 ;
      RECT  31965.0 87195.0 32670.0 88540.0 ;
      RECT  31965.0 89885.0 32670.0 88540.0 ;
      RECT  31965.0 89885.0 32670.0 91230.0 ;
      RECT  31965.0 92575.0 32670.0 91230.0 ;
      RECT  31965.0 92575.0 32670.0 93920.0 ;
      RECT  31965.0 95265.0 32670.0 93920.0 ;
      RECT  31965.0 95265.0 32670.0 96610.0 ;
      RECT  31965.0 97955.0 32670.0 96610.0 ;
      RECT  31965.0 97955.0 32670.0 99300.0 ;
      RECT  31965.0 100645.0 32670.0 99300.0 ;
      RECT  31965.0 100645.0 32670.0 101990.0 ;
      RECT  31965.0 103335.0 32670.0 101990.0 ;
      RECT  31965.0 103335.0 32670.0 104680.0 ;
      RECT  31965.0 106025.0 32670.0 104680.0 ;
      RECT  31965.0 106025.0 32670.0 107370.0 ;
      RECT  31965.0 108715.0 32670.0 107370.0 ;
      RECT  31965.0 108715.0 32670.0 110060.0 ;
      RECT  31965.0 111405.0 32670.0 110060.0 ;
      RECT  31965.0 111405.0 32670.0 112750.0 ;
      RECT  31965.0 114095.0 32670.0 112750.0 ;
      RECT  32670.0 28015.0 33375.0 29360.0 ;
      RECT  32670.0 30705.0 33375.0 29360.0 ;
      RECT  32670.0 30705.0 33375.0 32050.0 ;
      RECT  32670.0 33395.0 33375.0 32050.0 ;
      RECT  32670.0 33395.0 33375.0 34740.0 ;
      RECT  32670.0 36085.0 33375.0 34740.0 ;
      RECT  32670.0 36085.0 33375.0 37430.0 ;
      RECT  32670.0 38775.0 33375.0 37430.0 ;
      RECT  32670.0 38775.0 33375.0 40120.0 ;
      RECT  32670.0 41465.0 33375.0 40120.0 ;
      RECT  32670.0 41465.0 33375.0 42810.0 ;
      RECT  32670.0 44155.0 33375.0 42810.0 ;
      RECT  32670.0 44155.0 33375.0 45500.0 ;
      RECT  32670.0 46845.0 33375.0 45500.0 ;
      RECT  32670.0 46845.0 33375.0 48190.0 ;
      RECT  32670.0 49535.0 33375.0 48190.0 ;
      RECT  32670.0 49535.0 33375.0 50880.0 ;
      RECT  32670.0 52225.0 33375.0 50880.0 ;
      RECT  32670.0 52225.0 33375.0 53570.0 ;
      RECT  32670.0 54915.0 33375.0 53570.0 ;
      RECT  32670.0 54915.0 33375.0 56260.0 ;
      RECT  32670.0 57605.0 33375.0 56260.0 ;
      RECT  32670.0 57605.0 33375.0 58950.0 ;
      RECT  32670.0 60295.0 33375.0 58950.0 ;
      RECT  32670.0 60295.0 33375.0 61640.0 ;
      RECT  32670.0 62985.0 33375.0 61640.0 ;
      RECT  32670.0 62985.0 33375.0 64330.0 ;
      RECT  32670.0 65675.0 33375.0 64330.0 ;
      RECT  32670.0 65675.0 33375.0 67020.0 ;
      RECT  32670.0 68365.0 33375.0 67020.0 ;
      RECT  32670.0 68365.0 33375.0 69710.0 ;
      RECT  32670.0 71055.0 33375.0 69710.0 ;
      RECT  32670.0 71055.0 33375.0 72400.0 ;
      RECT  32670.0 73745.0 33375.0 72400.0 ;
      RECT  32670.0 73745.0 33375.0 75090.0 ;
      RECT  32670.0 76435.0 33375.0 75090.0 ;
      RECT  32670.0 76435.0 33375.0 77780.0 ;
      RECT  32670.0 79125.0 33375.0 77780.0 ;
      RECT  32670.0 79125.0 33375.0 80470.0 ;
      RECT  32670.0 81815.0 33375.0 80470.0 ;
      RECT  32670.0 81815.0 33375.0 83160.0 ;
      RECT  32670.0 84505.0 33375.0 83160.0 ;
      RECT  32670.0 84505.0 33375.0 85850.0 ;
      RECT  32670.0 87195.0 33375.0 85850.0 ;
      RECT  32670.0 87195.0 33375.0 88540.0 ;
      RECT  32670.0 89885.0 33375.0 88540.0 ;
      RECT  32670.0 89885.0 33375.0 91230.0 ;
      RECT  32670.0 92575.0 33375.0 91230.0 ;
      RECT  32670.0 92575.0 33375.0 93920.0 ;
      RECT  32670.0 95265.0 33375.0 93920.0 ;
      RECT  32670.0 95265.0 33375.0 96610.0 ;
      RECT  32670.0 97955.0 33375.0 96610.0 ;
      RECT  32670.0 97955.0 33375.0 99300.0 ;
      RECT  32670.0 100645.0 33375.0 99300.0 ;
      RECT  32670.0 100645.0 33375.0 101990.0 ;
      RECT  32670.0 103335.0 33375.0 101990.0 ;
      RECT  32670.0 103335.0 33375.0 104680.0 ;
      RECT  32670.0 106025.0 33375.0 104680.0 ;
      RECT  32670.0 106025.0 33375.0 107370.0 ;
      RECT  32670.0 108715.0 33375.0 107370.0 ;
      RECT  32670.0 108715.0 33375.0 110060.0 ;
      RECT  32670.0 111405.0 33375.0 110060.0 ;
      RECT  32670.0 111405.0 33375.0 112750.0 ;
      RECT  32670.0 114095.0 33375.0 112750.0 ;
      RECT  33375.0 28015.0 34080.0 29360.0 ;
      RECT  33375.0 30705.0 34080.0 29360.0 ;
      RECT  33375.0 30705.0 34080.0 32050.0 ;
      RECT  33375.0 33395.0 34080.0 32050.0 ;
      RECT  33375.0 33395.0 34080.0 34740.0 ;
      RECT  33375.0 36085.0 34080.0 34740.0 ;
      RECT  33375.0 36085.0 34080.0 37430.0 ;
      RECT  33375.0 38775.0 34080.0 37430.0 ;
      RECT  33375.0 38775.0 34080.0 40120.0 ;
      RECT  33375.0 41465.0 34080.0 40120.0 ;
      RECT  33375.0 41465.0 34080.0 42810.0 ;
      RECT  33375.0 44155.0 34080.0 42810.0 ;
      RECT  33375.0 44155.0 34080.0 45500.0 ;
      RECT  33375.0 46845.0 34080.0 45500.0 ;
      RECT  33375.0 46845.0 34080.0 48190.0 ;
      RECT  33375.0 49535.0 34080.0 48190.0 ;
      RECT  33375.0 49535.0 34080.0 50880.0 ;
      RECT  33375.0 52225.0 34080.0 50880.0 ;
      RECT  33375.0 52225.0 34080.0 53570.0 ;
      RECT  33375.0 54915.0 34080.0 53570.0 ;
      RECT  33375.0 54915.0 34080.0 56260.0 ;
      RECT  33375.0 57605.0 34080.0 56260.0 ;
      RECT  33375.0 57605.0 34080.0 58950.0 ;
      RECT  33375.0 60295.0 34080.0 58950.0 ;
      RECT  33375.0 60295.0 34080.0 61640.0 ;
      RECT  33375.0 62985.0 34080.0 61640.0 ;
      RECT  33375.0 62985.0 34080.0 64330.0 ;
      RECT  33375.0 65675.0 34080.0 64330.0 ;
      RECT  33375.0 65675.0 34080.0 67020.0 ;
      RECT  33375.0 68365.0 34080.0 67020.0 ;
      RECT  33375.0 68365.0 34080.0 69710.0 ;
      RECT  33375.0 71055.0 34080.0 69710.0 ;
      RECT  33375.0 71055.0 34080.0 72400.0 ;
      RECT  33375.0 73745.0 34080.0 72400.0 ;
      RECT  33375.0 73745.0 34080.0 75090.0 ;
      RECT  33375.0 76435.0 34080.0 75090.0 ;
      RECT  33375.0 76435.0 34080.0 77780.0 ;
      RECT  33375.0 79125.0 34080.0 77780.0 ;
      RECT  33375.0 79125.0 34080.0 80470.0 ;
      RECT  33375.0 81815.0 34080.0 80470.0 ;
      RECT  33375.0 81815.0 34080.0 83160.0 ;
      RECT  33375.0 84505.0 34080.0 83160.0 ;
      RECT  33375.0 84505.0 34080.0 85850.0 ;
      RECT  33375.0 87195.0 34080.0 85850.0 ;
      RECT  33375.0 87195.0 34080.0 88540.0 ;
      RECT  33375.0 89885.0 34080.0 88540.0 ;
      RECT  33375.0 89885.0 34080.0 91230.0 ;
      RECT  33375.0 92575.0 34080.0 91230.0 ;
      RECT  33375.0 92575.0 34080.0 93920.0 ;
      RECT  33375.0 95265.0 34080.0 93920.0 ;
      RECT  33375.0 95265.0 34080.0 96610.0 ;
      RECT  33375.0 97955.0 34080.0 96610.0 ;
      RECT  33375.0 97955.0 34080.0 99300.0 ;
      RECT  33375.0 100645.0 34080.0 99300.0 ;
      RECT  33375.0 100645.0 34080.0 101990.0 ;
      RECT  33375.0 103335.0 34080.0 101990.0 ;
      RECT  33375.0 103335.0 34080.0 104680.0 ;
      RECT  33375.0 106025.0 34080.0 104680.0 ;
      RECT  33375.0 106025.0 34080.0 107370.0 ;
      RECT  33375.0 108715.0 34080.0 107370.0 ;
      RECT  33375.0 108715.0 34080.0 110060.0 ;
      RECT  33375.0 111405.0 34080.0 110060.0 ;
      RECT  33375.0 111405.0 34080.0 112750.0 ;
      RECT  33375.0 114095.0 34080.0 112750.0 ;
      RECT  34080.0 28015.0 34785.0 29360.0 ;
      RECT  34080.0 30705.0 34785.0 29360.0 ;
      RECT  34080.0 30705.0 34785.0 32050.0 ;
      RECT  34080.0 33395.0 34785.0 32050.0 ;
      RECT  34080.0 33395.0 34785.0 34740.0 ;
      RECT  34080.0 36085.0 34785.0 34740.0 ;
      RECT  34080.0 36085.0 34785.0 37430.0 ;
      RECT  34080.0 38775.0 34785.0 37430.0 ;
      RECT  34080.0 38775.0 34785.0 40120.0 ;
      RECT  34080.0 41465.0 34785.0 40120.0 ;
      RECT  34080.0 41465.0 34785.0 42810.0 ;
      RECT  34080.0 44155.0 34785.0 42810.0 ;
      RECT  34080.0 44155.0 34785.0 45500.0 ;
      RECT  34080.0 46845.0 34785.0 45500.0 ;
      RECT  34080.0 46845.0 34785.0 48190.0 ;
      RECT  34080.0 49535.0 34785.0 48190.0 ;
      RECT  34080.0 49535.0 34785.0 50880.0 ;
      RECT  34080.0 52225.0 34785.0 50880.0 ;
      RECT  34080.0 52225.0 34785.0 53570.0 ;
      RECT  34080.0 54915.0 34785.0 53570.0 ;
      RECT  34080.0 54915.0 34785.0 56260.0 ;
      RECT  34080.0 57605.0 34785.0 56260.0 ;
      RECT  34080.0 57605.0 34785.0 58950.0 ;
      RECT  34080.0 60295.0 34785.0 58950.0 ;
      RECT  34080.0 60295.0 34785.0 61640.0 ;
      RECT  34080.0 62985.0 34785.0 61640.0 ;
      RECT  34080.0 62985.0 34785.0 64330.0 ;
      RECT  34080.0 65675.0 34785.0 64330.0 ;
      RECT  34080.0 65675.0 34785.0 67020.0 ;
      RECT  34080.0 68365.0 34785.0 67020.0 ;
      RECT  34080.0 68365.0 34785.0 69710.0 ;
      RECT  34080.0 71055.0 34785.0 69710.0 ;
      RECT  34080.0 71055.0 34785.0 72400.0 ;
      RECT  34080.0 73745.0 34785.0 72400.0 ;
      RECT  34080.0 73745.0 34785.0 75090.0 ;
      RECT  34080.0 76435.0 34785.0 75090.0 ;
      RECT  34080.0 76435.0 34785.0 77780.0 ;
      RECT  34080.0 79125.0 34785.0 77780.0 ;
      RECT  34080.0 79125.0 34785.0 80470.0 ;
      RECT  34080.0 81815.0 34785.0 80470.0 ;
      RECT  34080.0 81815.0 34785.0 83160.0 ;
      RECT  34080.0 84505.0 34785.0 83160.0 ;
      RECT  34080.0 84505.0 34785.0 85850.0 ;
      RECT  34080.0 87195.0 34785.0 85850.0 ;
      RECT  34080.0 87195.0 34785.0 88540.0 ;
      RECT  34080.0 89885.0 34785.0 88540.0 ;
      RECT  34080.0 89885.0 34785.0 91230.0 ;
      RECT  34080.0 92575.0 34785.0 91230.0 ;
      RECT  34080.0 92575.0 34785.0 93920.0 ;
      RECT  34080.0 95265.0 34785.0 93920.0 ;
      RECT  34080.0 95265.0 34785.0 96610.0 ;
      RECT  34080.0 97955.0 34785.0 96610.0 ;
      RECT  34080.0 97955.0 34785.0 99300.0 ;
      RECT  34080.0 100645.0 34785.0 99300.0 ;
      RECT  34080.0 100645.0 34785.0 101990.0 ;
      RECT  34080.0 103335.0 34785.0 101990.0 ;
      RECT  34080.0 103335.0 34785.0 104680.0 ;
      RECT  34080.0 106025.0 34785.0 104680.0 ;
      RECT  34080.0 106025.0 34785.0 107370.0 ;
      RECT  34080.0 108715.0 34785.0 107370.0 ;
      RECT  34080.0 108715.0 34785.0 110060.0 ;
      RECT  34080.0 111405.0 34785.0 110060.0 ;
      RECT  34080.0 111405.0 34785.0 112750.0 ;
      RECT  34080.0 114095.0 34785.0 112750.0 ;
      RECT  34785.0 28015.0 35490.0 29360.0 ;
      RECT  34785.0 30705.0 35490.0 29360.0 ;
      RECT  34785.0 30705.0 35490.0 32050.0 ;
      RECT  34785.0 33395.0 35490.0 32050.0 ;
      RECT  34785.0 33395.0 35490.0 34740.0 ;
      RECT  34785.0 36085.0 35490.0 34740.0 ;
      RECT  34785.0 36085.0 35490.0 37430.0 ;
      RECT  34785.0 38775.0 35490.0 37430.0 ;
      RECT  34785.0 38775.0 35490.0 40120.0 ;
      RECT  34785.0 41465.0 35490.0 40120.0 ;
      RECT  34785.0 41465.0 35490.0 42810.0 ;
      RECT  34785.0 44155.0 35490.0 42810.0 ;
      RECT  34785.0 44155.0 35490.0 45500.0 ;
      RECT  34785.0 46845.0 35490.0 45500.0 ;
      RECT  34785.0 46845.0 35490.0 48190.0 ;
      RECT  34785.0 49535.0 35490.0 48190.0 ;
      RECT  34785.0 49535.0 35490.0 50880.0 ;
      RECT  34785.0 52225.0 35490.0 50880.0 ;
      RECT  34785.0 52225.0 35490.0 53570.0 ;
      RECT  34785.0 54915.0 35490.0 53570.0 ;
      RECT  34785.0 54915.0 35490.0 56260.0 ;
      RECT  34785.0 57605.0 35490.0 56260.0 ;
      RECT  34785.0 57605.0 35490.0 58950.0 ;
      RECT  34785.0 60295.0 35490.0 58950.0 ;
      RECT  34785.0 60295.0 35490.0 61640.0 ;
      RECT  34785.0 62985.0 35490.0 61640.0 ;
      RECT  34785.0 62985.0 35490.0 64330.0 ;
      RECT  34785.0 65675.0 35490.0 64330.0 ;
      RECT  34785.0 65675.0 35490.0 67020.0 ;
      RECT  34785.0 68365.0 35490.0 67020.0 ;
      RECT  34785.0 68365.0 35490.0 69710.0 ;
      RECT  34785.0 71055.0 35490.0 69710.0 ;
      RECT  34785.0 71055.0 35490.0 72400.0 ;
      RECT  34785.0 73745.0 35490.0 72400.0 ;
      RECT  34785.0 73745.0 35490.0 75090.0 ;
      RECT  34785.0 76435.0 35490.0 75090.0 ;
      RECT  34785.0 76435.0 35490.0 77780.0 ;
      RECT  34785.0 79125.0 35490.0 77780.0 ;
      RECT  34785.0 79125.0 35490.0 80470.0 ;
      RECT  34785.0 81815.0 35490.0 80470.0 ;
      RECT  34785.0 81815.0 35490.0 83160.0 ;
      RECT  34785.0 84505.0 35490.0 83160.0 ;
      RECT  34785.0 84505.0 35490.0 85850.0 ;
      RECT  34785.0 87195.0 35490.0 85850.0 ;
      RECT  34785.0 87195.0 35490.0 88540.0 ;
      RECT  34785.0 89885.0 35490.0 88540.0 ;
      RECT  34785.0 89885.0 35490.0 91230.0 ;
      RECT  34785.0 92575.0 35490.0 91230.0 ;
      RECT  34785.0 92575.0 35490.0 93920.0 ;
      RECT  34785.0 95265.0 35490.0 93920.0 ;
      RECT  34785.0 95265.0 35490.0 96610.0 ;
      RECT  34785.0 97955.0 35490.0 96610.0 ;
      RECT  34785.0 97955.0 35490.0 99300.0 ;
      RECT  34785.0 100645.0 35490.0 99300.0 ;
      RECT  34785.0 100645.0 35490.0 101990.0 ;
      RECT  34785.0 103335.0 35490.0 101990.0 ;
      RECT  34785.0 103335.0 35490.0 104680.0 ;
      RECT  34785.0 106025.0 35490.0 104680.0 ;
      RECT  34785.0 106025.0 35490.0 107370.0 ;
      RECT  34785.0 108715.0 35490.0 107370.0 ;
      RECT  34785.0 108715.0 35490.0 110060.0 ;
      RECT  34785.0 111405.0 35490.0 110060.0 ;
      RECT  34785.0 111405.0 35490.0 112750.0 ;
      RECT  34785.0 114095.0 35490.0 112750.0 ;
      RECT  35490.0 28015.0 36195.0 29360.0 ;
      RECT  35490.0 30705.0 36195.0 29360.0 ;
      RECT  35490.0 30705.0 36195.0 32050.0 ;
      RECT  35490.0 33395.0 36195.0 32050.0 ;
      RECT  35490.0 33395.0 36195.0 34740.0 ;
      RECT  35490.0 36085.0 36195.0 34740.0 ;
      RECT  35490.0 36085.0 36195.0 37430.0 ;
      RECT  35490.0 38775.0 36195.0 37430.0 ;
      RECT  35490.0 38775.0 36195.0 40120.0 ;
      RECT  35490.0 41465.0 36195.0 40120.0 ;
      RECT  35490.0 41465.0 36195.0 42810.0 ;
      RECT  35490.0 44155.0 36195.0 42810.0 ;
      RECT  35490.0 44155.0 36195.0 45500.0 ;
      RECT  35490.0 46845.0 36195.0 45500.0 ;
      RECT  35490.0 46845.0 36195.0 48190.0 ;
      RECT  35490.0 49535.0 36195.0 48190.0 ;
      RECT  35490.0 49535.0 36195.0 50880.0 ;
      RECT  35490.0 52225.0 36195.0 50880.0 ;
      RECT  35490.0 52225.0 36195.0 53570.0 ;
      RECT  35490.0 54915.0 36195.0 53570.0 ;
      RECT  35490.0 54915.0 36195.0 56260.0 ;
      RECT  35490.0 57605.0 36195.0 56260.0 ;
      RECT  35490.0 57605.0 36195.0 58950.0 ;
      RECT  35490.0 60295.0 36195.0 58950.0 ;
      RECT  35490.0 60295.0 36195.0 61640.0 ;
      RECT  35490.0 62985.0 36195.0 61640.0 ;
      RECT  35490.0 62985.0 36195.0 64330.0 ;
      RECT  35490.0 65675.0 36195.0 64330.0 ;
      RECT  35490.0 65675.0 36195.0 67020.0 ;
      RECT  35490.0 68365.0 36195.0 67020.0 ;
      RECT  35490.0 68365.0 36195.0 69710.0 ;
      RECT  35490.0 71055.0 36195.0 69710.0 ;
      RECT  35490.0 71055.0 36195.0 72400.0 ;
      RECT  35490.0 73745.0 36195.0 72400.0 ;
      RECT  35490.0 73745.0 36195.0 75090.0 ;
      RECT  35490.0 76435.0 36195.0 75090.0 ;
      RECT  35490.0 76435.0 36195.0 77780.0 ;
      RECT  35490.0 79125.0 36195.0 77780.0 ;
      RECT  35490.0 79125.0 36195.0 80470.0 ;
      RECT  35490.0 81815.0 36195.0 80470.0 ;
      RECT  35490.0 81815.0 36195.0 83160.0 ;
      RECT  35490.0 84505.0 36195.0 83160.0 ;
      RECT  35490.0 84505.0 36195.0 85850.0 ;
      RECT  35490.0 87195.0 36195.0 85850.0 ;
      RECT  35490.0 87195.0 36195.0 88540.0 ;
      RECT  35490.0 89885.0 36195.0 88540.0 ;
      RECT  35490.0 89885.0 36195.0 91230.0 ;
      RECT  35490.0 92575.0 36195.0 91230.0 ;
      RECT  35490.0 92575.0 36195.0 93920.0 ;
      RECT  35490.0 95265.0 36195.0 93920.0 ;
      RECT  35490.0 95265.0 36195.0 96610.0 ;
      RECT  35490.0 97955.0 36195.0 96610.0 ;
      RECT  35490.0 97955.0 36195.0 99300.0 ;
      RECT  35490.0 100645.0 36195.0 99300.0 ;
      RECT  35490.0 100645.0 36195.0 101990.0 ;
      RECT  35490.0 103335.0 36195.0 101990.0 ;
      RECT  35490.0 103335.0 36195.0 104680.0 ;
      RECT  35490.0 106025.0 36195.0 104680.0 ;
      RECT  35490.0 106025.0 36195.0 107370.0 ;
      RECT  35490.0 108715.0 36195.0 107370.0 ;
      RECT  35490.0 108715.0 36195.0 110060.0 ;
      RECT  35490.0 111405.0 36195.0 110060.0 ;
      RECT  35490.0 111405.0 36195.0 112750.0 ;
      RECT  35490.0 114095.0 36195.0 112750.0 ;
      RECT  36195.0 28015.0 36900.0 29360.0 ;
      RECT  36195.0 30705.0 36900.0 29360.0 ;
      RECT  36195.0 30705.0 36900.0 32050.0 ;
      RECT  36195.0 33395.0 36900.0 32050.0 ;
      RECT  36195.0 33395.0 36900.0 34740.0 ;
      RECT  36195.0 36085.0 36900.0 34740.0 ;
      RECT  36195.0 36085.0 36900.0 37430.0 ;
      RECT  36195.0 38775.0 36900.0 37430.0 ;
      RECT  36195.0 38775.0 36900.0 40120.0 ;
      RECT  36195.0 41465.0 36900.0 40120.0 ;
      RECT  36195.0 41465.0 36900.0 42810.0 ;
      RECT  36195.0 44155.0 36900.0 42810.0 ;
      RECT  36195.0 44155.0 36900.0 45500.0 ;
      RECT  36195.0 46845.0 36900.0 45500.0 ;
      RECT  36195.0 46845.0 36900.0 48190.0 ;
      RECT  36195.0 49535.0 36900.0 48190.0 ;
      RECT  36195.0 49535.0 36900.0 50880.0 ;
      RECT  36195.0 52225.0 36900.0 50880.0 ;
      RECT  36195.0 52225.0 36900.0 53570.0 ;
      RECT  36195.0 54915.0 36900.0 53570.0 ;
      RECT  36195.0 54915.0 36900.0 56260.0 ;
      RECT  36195.0 57605.0 36900.0 56260.0 ;
      RECT  36195.0 57605.0 36900.0 58950.0 ;
      RECT  36195.0 60295.0 36900.0 58950.0 ;
      RECT  36195.0 60295.0 36900.0 61640.0 ;
      RECT  36195.0 62985.0 36900.0 61640.0 ;
      RECT  36195.0 62985.0 36900.0 64330.0 ;
      RECT  36195.0 65675.0 36900.0 64330.0 ;
      RECT  36195.0 65675.0 36900.0 67020.0 ;
      RECT  36195.0 68365.0 36900.0 67020.0 ;
      RECT  36195.0 68365.0 36900.0 69710.0 ;
      RECT  36195.0 71055.0 36900.0 69710.0 ;
      RECT  36195.0 71055.0 36900.0 72400.0 ;
      RECT  36195.0 73745.0 36900.0 72400.0 ;
      RECT  36195.0 73745.0 36900.0 75090.0 ;
      RECT  36195.0 76435.0 36900.0 75090.0 ;
      RECT  36195.0 76435.0 36900.0 77780.0 ;
      RECT  36195.0 79125.0 36900.0 77780.0 ;
      RECT  36195.0 79125.0 36900.0 80470.0 ;
      RECT  36195.0 81815.0 36900.0 80470.0 ;
      RECT  36195.0 81815.0 36900.0 83160.0 ;
      RECT  36195.0 84505.0 36900.0 83160.0 ;
      RECT  36195.0 84505.0 36900.0 85850.0 ;
      RECT  36195.0 87195.0 36900.0 85850.0 ;
      RECT  36195.0 87195.0 36900.0 88540.0 ;
      RECT  36195.0 89885.0 36900.0 88540.0 ;
      RECT  36195.0 89885.0 36900.0 91230.0 ;
      RECT  36195.0 92575.0 36900.0 91230.0 ;
      RECT  36195.0 92575.0 36900.0 93920.0 ;
      RECT  36195.0 95265.0 36900.0 93920.0 ;
      RECT  36195.0 95265.0 36900.0 96610.0 ;
      RECT  36195.0 97955.0 36900.0 96610.0 ;
      RECT  36195.0 97955.0 36900.0 99300.0 ;
      RECT  36195.0 100645.0 36900.0 99300.0 ;
      RECT  36195.0 100645.0 36900.0 101990.0 ;
      RECT  36195.0 103335.0 36900.0 101990.0 ;
      RECT  36195.0 103335.0 36900.0 104680.0 ;
      RECT  36195.0 106025.0 36900.0 104680.0 ;
      RECT  36195.0 106025.0 36900.0 107370.0 ;
      RECT  36195.0 108715.0 36900.0 107370.0 ;
      RECT  36195.0 108715.0 36900.0 110060.0 ;
      RECT  36195.0 111405.0 36900.0 110060.0 ;
      RECT  36195.0 111405.0 36900.0 112750.0 ;
      RECT  36195.0 114095.0 36900.0 112750.0 ;
      RECT  36900.0 28015.0 37605.0 29360.0 ;
      RECT  36900.0 30705.0 37605.0 29360.0 ;
      RECT  36900.0 30705.0 37605.0 32050.0 ;
      RECT  36900.0 33395.0 37605.0 32050.0 ;
      RECT  36900.0 33395.0 37605.0 34740.0 ;
      RECT  36900.0 36085.0 37605.0 34740.0 ;
      RECT  36900.0 36085.0 37605.0 37430.0 ;
      RECT  36900.0 38775.0 37605.0 37430.0 ;
      RECT  36900.0 38775.0 37605.0 40120.0 ;
      RECT  36900.0 41465.0 37605.0 40120.0 ;
      RECT  36900.0 41465.0 37605.0 42810.0 ;
      RECT  36900.0 44155.0 37605.0 42810.0 ;
      RECT  36900.0 44155.0 37605.0 45500.0 ;
      RECT  36900.0 46845.0 37605.0 45500.0 ;
      RECT  36900.0 46845.0 37605.0 48190.0 ;
      RECT  36900.0 49535.0 37605.0 48190.0 ;
      RECT  36900.0 49535.0 37605.0 50880.0 ;
      RECT  36900.0 52225.0 37605.0 50880.0 ;
      RECT  36900.0 52225.0 37605.0 53570.0 ;
      RECT  36900.0 54915.0 37605.0 53570.0 ;
      RECT  36900.0 54915.0 37605.0 56260.0 ;
      RECT  36900.0 57605.0 37605.0 56260.0 ;
      RECT  36900.0 57605.0 37605.0 58950.0 ;
      RECT  36900.0 60295.0 37605.0 58950.0 ;
      RECT  36900.0 60295.0 37605.0 61640.0 ;
      RECT  36900.0 62985.0 37605.0 61640.0 ;
      RECT  36900.0 62985.0 37605.0 64330.0 ;
      RECT  36900.0 65675.0 37605.0 64330.0 ;
      RECT  36900.0 65675.0 37605.0 67020.0 ;
      RECT  36900.0 68365.0 37605.0 67020.0 ;
      RECT  36900.0 68365.0 37605.0 69710.0 ;
      RECT  36900.0 71055.0 37605.0 69710.0 ;
      RECT  36900.0 71055.0 37605.0 72400.0 ;
      RECT  36900.0 73745.0 37605.0 72400.0 ;
      RECT  36900.0 73745.0 37605.0 75090.0 ;
      RECT  36900.0 76435.0 37605.0 75090.0 ;
      RECT  36900.0 76435.0 37605.0 77780.0 ;
      RECT  36900.0 79125.0 37605.0 77780.0 ;
      RECT  36900.0 79125.0 37605.0 80470.0 ;
      RECT  36900.0 81815.0 37605.0 80470.0 ;
      RECT  36900.0 81815.0 37605.0 83160.0 ;
      RECT  36900.0 84505.0 37605.0 83160.0 ;
      RECT  36900.0 84505.0 37605.0 85850.0 ;
      RECT  36900.0 87195.0 37605.0 85850.0 ;
      RECT  36900.0 87195.0 37605.0 88540.0 ;
      RECT  36900.0 89885.0 37605.0 88540.0 ;
      RECT  36900.0 89885.0 37605.0 91230.0 ;
      RECT  36900.0 92575.0 37605.0 91230.0 ;
      RECT  36900.0 92575.0 37605.0 93920.0 ;
      RECT  36900.0 95265.0 37605.0 93920.0 ;
      RECT  36900.0 95265.0 37605.0 96610.0 ;
      RECT  36900.0 97955.0 37605.0 96610.0 ;
      RECT  36900.0 97955.0 37605.0 99300.0 ;
      RECT  36900.0 100645.0 37605.0 99300.0 ;
      RECT  36900.0 100645.0 37605.0 101990.0 ;
      RECT  36900.0 103335.0 37605.0 101990.0 ;
      RECT  36900.0 103335.0 37605.0 104680.0 ;
      RECT  36900.0 106025.0 37605.0 104680.0 ;
      RECT  36900.0 106025.0 37605.0 107370.0 ;
      RECT  36900.0 108715.0 37605.0 107370.0 ;
      RECT  36900.0 108715.0 37605.0 110060.0 ;
      RECT  36900.0 111405.0 37605.0 110060.0 ;
      RECT  36900.0 111405.0 37605.0 112750.0 ;
      RECT  36900.0 114095.0 37605.0 112750.0 ;
      RECT  37605.0 28015.0 38310.0 29360.0 ;
      RECT  37605.0 30705.0 38310.0 29360.0 ;
      RECT  37605.0 30705.0 38310.0 32050.0 ;
      RECT  37605.0 33395.0 38310.0 32050.0 ;
      RECT  37605.0 33395.0 38310.0 34740.0 ;
      RECT  37605.0 36085.0 38310.0 34740.0 ;
      RECT  37605.0 36085.0 38310.0 37430.0 ;
      RECT  37605.0 38775.0 38310.0 37430.0 ;
      RECT  37605.0 38775.0 38310.0 40120.0 ;
      RECT  37605.0 41465.0 38310.0 40120.0 ;
      RECT  37605.0 41465.0 38310.0 42810.0 ;
      RECT  37605.0 44155.0 38310.0 42810.0 ;
      RECT  37605.0 44155.0 38310.0 45500.0 ;
      RECT  37605.0 46845.0 38310.0 45500.0 ;
      RECT  37605.0 46845.0 38310.0 48190.0 ;
      RECT  37605.0 49535.0 38310.0 48190.0 ;
      RECT  37605.0 49535.0 38310.0 50880.0 ;
      RECT  37605.0 52225.0 38310.0 50880.0 ;
      RECT  37605.0 52225.0 38310.0 53570.0 ;
      RECT  37605.0 54915.0 38310.0 53570.0 ;
      RECT  37605.0 54915.0 38310.0 56260.0 ;
      RECT  37605.0 57605.0 38310.0 56260.0 ;
      RECT  37605.0 57605.0 38310.0 58950.0 ;
      RECT  37605.0 60295.0 38310.0 58950.0 ;
      RECT  37605.0 60295.0 38310.0 61640.0 ;
      RECT  37605.0 62985.0 38310.0 61640.0 ;
      RECT  37605.0 62985.0 38310.0 64330.0 ;
      RECT  37605.0 65675.0 38310.0 64330.0 ;
      RECT  37605.0 65675.0 38310.0 67020.0 ;
      RECT  37605.0 68365.0 38310.0 67020.0 ;
      RECT  37605.0 68365.0 38310.0 69710.0 ;
      RECT  37605.0 71055.0 38310.0 69710.0 ;
      RECT  37605.0 71055.0 38310.0 72400.0 ;
      RECT  37605.0 73745.0 38310.0 72400.0 ;
      RECT  37605.0 73745.0 38310.0 75090.0 ;
      RECT  37605.0 76435.0 38310.0 75090.0 ;
      RECT  37605.0 76435.0 38310.0 77780.0 ;
      RECT  37605.0 79125.0 38310.0 77780.0 ;
      RECT  37605.0 79125.0 38310.0 80470.0 ;
      RECT  37605.0 81815.0 38310.0 80470.0 ;
      RECT  37605.0 81815.0 38310.0 83160.0 ;
      RECT  37605.0 84505.0 38310.0 83160.0 ;
      RECT  37605.0 84505.0 38310.0 85850.0 ;
      RECT  37605.0 87195.0 38310.0 85850.0 ;
      RECT  37605.0 87195.0 38310.0 88540.0 ;
      RECT  37605.0 89885.0 38310.0 88540.0 ;
      RECT  37605.0 89885.0 38310.0 91230.0 ;
      RECT  37605.0 92575.0 38310.0 91230.0 ;
      RECT  37605.0 92575.0 38310.0 93920.0 ;
      RECT  37605.0 95265.0 38310.0 93920.0 ;
      RECT  37605.0 95265.0 38310.0 96610.0 ;
      RECT  37605.0 97955.0 38310.0 96610.0 ;
      RECT  37605.0 97955.0 38310.0 99300.0 ;
      RECT  37605.0 100645.0 38310.0 99300.0 ;
      RECT  37605.0 100645.0 38310.0 101990.0 ;
      RECT  37605.0 103335.0 38310.0 101990.0 ;
      RECT  37605.0 103335.0 38310.0 104680.0 ;
      RECT  37605.0 106025.0 38310.0 104680.0 ;
      RECT  37605.0 106025.0 38310.0 107370.0 ;
      RECT  37605.0 108715.0 38310.0 107370.0 ;
      RECT  37605.0 108715.0 38310.0 110060.0 ;
      RECT  37605.0 111405.0 38310.0 110060.0 ;
      RECT  37605.0 111405.0 38310.0 112750.0 ;
      RECT  37605.0 114095.0 38310.0 112750.0 ;
      RECT  38310.0 28015.0 39015.0 29360.0 ;
      RECT  38310.0 30705.0 39015.0 29360.0 ;
      RECT  38310.0 30705.0 39015.0 32050.0 ;
      RECT  38310.0 33395.0 39015.0 32050.0 ;
      RECT  38310.0 33395.0 39015.0 34740.0 ;
      RECT  38310.0 36085.0 39015.0 34740.0 ;
      RECT  38310.0 36085.0 39015.0 37430.0 ;
      RECT  38310.0 38775.0 39015.0 37430.0 ;
      RECT  38310.0 38775.0 39015.0 40120.0 ;
      RECT  38310.0 41465.0 39015.0 40120.0 ;
      RECT  38310.0 41465.0 39015.0 42810.0 ;
      RECT  38310.0 44155.0 39015.0 42810.0 ;
      RECT  38310.0 44155.0 39015.0 45500.0 ;
      RECT  38310.0 46845.0 39015.0 45500.0 ;
      RECT  38310.0 46845.0 39015.0 48190.0 ;
      RECT  38310.0 49535.0 39015.0 48190.0 ;
      RECT  38310.0 49535.0 39015.0 50880.0 ;
      RECT  38310.0 52225.0 39015.0 50880.0 ;
      RECT  38310.0 52225.0 39015.0 53570.0 ;
      RECT  38310.0 54915.0 39015.0 53570.0 ;
      RECT  38310.0 54915.0 39015.0 56260.0 ;
      RECT  38310.0 57605.0 39015.0 56260.0 ;
      RECT  38310.0 57605.0 39015.0 58950.0 ;
      RECT  38310.0 60295.0 39015.0 58950.0 ;
      RECT  38310.0 60295.0 39015.0 61640.0 ;
      RECT  38310.0 62985.0 39015.0 61640.0 ;
      RECT  38310.0 62985.0 39015.0 64330.0 ;
      RECT  38310.0 65675.0 39015.0 64330.0 ;
      RECT  38310.0 65675.0 39015.0 67020.0 ;
      RECT  38310.0 68365.0 39015.0 67020.0 ;
      RECT  38310.0 68365.0 39015.0 69710.0 ;
      RECT  38310.0 71055.0 39015.0 69710.0 ;
      RECT  38310.0 71055.0 39015.0 72400.0 ;
      RECT  38310.0 73745.0 39015.0 72400.0 ;
      RECT  38310.0 73745.0 39015.0 75090.0 ;
      RECT  38310.0 76435.0 39015.0 75090.0 ;
      RECT  38310.0 76435.0 39015.0 77780.0 ;
      RECT  38310.0 79125.0 39015.0 77780.0 ;
      RECT  38310.0 79125.0 39015.0 80470.0 ;
      RECT  38310.0 81815.0 39015.0 80470.0 ;
      RECT  38310.0 81815.0 39015.0 83160.0 ;
      RECT  38310.0 84505.0 39015.0 83160.0 ;
      RECT  38310.0 84505.0 39015.0 85850.0 ;
      RECT  38310.0 87195.0 39015.0 85850.0 ;
      RECT  38310.0 87195.0 39015.0 88540.0 ;
      RECT  38310.0 89885.0 39015.0 88540.0 ;
      RECT  38310.0 89885.0 39015.0 91230.0 ;
      RECT  38310.0 92575.0 39015.0 91230.0 ;
      RECT  38310.0 92575.0 39015.0 93920.0 ;
      RECT  38310.0 95265.0 39015.0 93920.0 ;
      RECT  38310.0 95265.0 39015.0 96610.0 ;
      RECT  38310.0 97955.0 39015.0 96610.0 ;
      RECT  38310.0 97955.0 39015.0 99300.0 ;
      RECT  38310.0 100645.0 39015.0 99300.0 ;
      RECT  38310.0 100645.0 39015.0 101990.0 ;
      RECT  38310.0 103335.0 39015.0 101990.0 ;
      RECT  38310.0 103335.0 39015.0 104680.0 ;
      RECT  38310.0 106025.0 39015.0 104680.0 ;
      RECT  38310.0 106025.0 39015.0 107370.0 ;
      RECT  38310.0 108715.0 39015.0 107370.0 ;
      RECT  38310.0 108715.0 39015.0 110060.0 ;
      RECT  38310.0 111405.0 39015.0 110060.0 ;
      RECT  38310.0 111405.0 39015.0 112750.0 ;
      RECT  38310.0 114095.0 39015.0 112750.0 ;
      RECT  39015.0 28015.0 39720.0 29360.0 ;
      RECT  39015.0 30705.0 39720.0 29360.0 ;
      RECT  39015.0 30705.0 39720.0 32050.0 ;
      RECT  39015.0 33395.0 39720.0 32050.0 ;
      RECT  39015.0 33395.0 39720.0 34740.0 ;
      RECT  39015.0 36085.0 39720.0 34740.0 ;
      RECT  39015.0 36085.0 39720.0 37430.0 ;
      RECT  39015.0 38775.0 39720.0 37430.0 ;
      RECT  39015.0 38775.0 39720.0 40120.0 ;
      RECT  39015.0 41465.0 39720.0 40120.0 ;
      RECT  39015.0 41465.0 39720.0 42810.0 ;
      RECT  39015.0 44155.0 39720.0 42810.0 ;
      RECT  39015.0 44155.0 39720.0 45500.0 ;
      RECT  39015.0 46845.0 39720.0 45500.0 ;
      RECT  39015.0 46845.0 39720.0 48190.0 ;
      RECT  39015.0 49535.0 39720.0 48190.0 ;
      RECT  39015.0 49535.0 39720.0 50880.0 ;
      RECT  39015.0 52225.0 39720.0 50880.0 ;
      RECT  39015.0 52225.0 39720.0 53570.0 ;
      RECT  39015.0 54915.0 39720.0 53570.0 ;
      RECT  39015.0 54915.0 39720.0 56260.0 ;
      RECT  39015.0 57605.0 39720.0 56260.0 ;
      RECT  39015.0 57605.0 39720.0 58950.0 ;
      RECT  39015.0 60295.0 39720.0 58950.0 ;
      RECT  39015.0 60295.0 39720.0 61640.0 ;
      RECT  39015.0 62985.0 39720.0 61640.0 ;
      RECT  39015.0 62985.0 39720.0 64330.0 ;
      RECT  39015.0 65675.0 39720.0 64330.0 ;
      RECT  39015.0 65675.0 39720.0 67020.0 ;
      RECT  39015.0 68365.0 39720.0 67020.0 ;
      RECT  39015.0 68365.0 39720.0 69710.0 ;
      RECT  39015.0 71055.0 39720.0 69710.0 ;
      RECT  39015.0 71055.0 39720.0 72400.0 ;
      RECT  39015.0 73745.0 39720.0 72400.0 ;
      RECT  39015.0 73745.0 39720.0 75090.0 ;
      RECT  39015.0 76435.0 39720.0 75090.0 ;
      RECT  39015.0 76435.0 39720.0 77780.0 ;
      RECT  39015.0 79125.0 39720.0 77780.0 ;
      RECT  39015.0 79125.0 39720.0 80470.0 ;
      RECT  39015.0 81815.0 39720.0 80470.0 ;
      RECT  39015.0 81815.0 39720.0 83160.0 ;
      RECT  39015.0 84505.0 39720.0 83160.0 ;
      RECT  39015.0 84505.0 39720.0 85850.0 ;
      RECT  39015.0 87195.0 39720.0 85850.0 ;
      RECT  39015.0 87195.0 39720.0 88540.0 ;
      RECT  39015.0 89885.0 39720.0 88540.0 ;
      RECT  39015.0 89885.0 39720.0 91230.0 ;
      RECT  39015.0 92575.0 39720.0 91230.0 ;
      RECT  39015.0 92575.0 39720.0 93920.0 ;
      RECT  39015.0 95265.0 39720.0 93920.0 ;
      RECT  39015.0 95265.0 39720.0 96610.0 ;
      RECT  39015.0 97955.0 39720.0 96610.0 ;
      RECT  39015.0 97955.0 39720.0 99300.0 ;
      RECT  39015.0 100645.0 39720.0 99300.0 ;
      RECT  39015.0 100645.0 39720.0 101990.0 ;
      RECT  39015.0 103335.0 39720.0 101990.0 ;
      RECT  39015.0 103335.0 39720.0 104680.0 ;
      RECT  39015.0 106025.0 39720.0 104680.0 ;
      RECT  39015.0 106025.0 39720.0 107370.0 ;
      RECT  39015.0 108715.0 39720.0 107370.0 ;
      RECT  39015.0 108715.0 39720.0 110060.0 ;
      RECT  39015.0 111405.0 39720.0 110060.0 ;
      RECT  39015.0 111405.0 39720.0 112750.0 ;
      RECT  39015.0 114095.0 39720.0 112750.0 ;
      RECT  39720.0 28015.0 40425.0 29360.0 ;
      RECT  39720.0 30705.0 40425.0 29360.0 ;
      RECT  39720.0 30705.0 40425.0 32050.0 ;
      RECT  39720.0 33395.0 40425.0 32050.0 ;
      RECT  39720.0 33395.0 40425.0 34740.0 ;
      RECT  39720.0 36085.0 40425.0 34740.0 ;
      RECT  39720.0 36085.0 40425.0 37430.0 ;
      RECT  39720.0 38775.0 40425.0 37430.0 ;
      RECT  39720.0 38775.0 40425.0 40120.0 ;
      RECT  39720.0 41465.0 40425.0 40120.0 ;
      RECT  39720.0 41465.0 40425.0 42810.0 ;
      RECT  39720.0 44155.0 40425.0 42810.0 ;
      RECT  39720.0 44155.0 40425.0 45500.0 ;
      RECT  39720.0 46845.0 40425.0 45500.0 ;
      RECT  39720.0 46845.0 40425.0 48190.0 ;
      RECT  39720.0 49535.0 40425.0 48190.0 ;
      RECT  39720.0 49535.0 40425.0 50880.0 ;
      RECT  39720.0 52225.0 40425.0 50880.0 ;
      RECT  39720.0 52225.0 40425.0 53570.0 ;
      RECT  39720.0 54915.0 40425.0 53570.0 ;
      RECT  39720.0 54915.0 40425.0 56260.0 ;
      RECT  39720.0 57605.0 40425.0 56260.0 ;
      RECT  39720.0 57605.0 40425.0 58950.0 ;
      RECT  39720.0 60295.0 40425.0 58950.0 ;
      RECT  39720.0 60295.0 40425.0 61640.0 ;
      RECT  39720.0 62985.0 40425.0 61640.0 ;
      RECT  39720.0 62985.0 40425.0 64330.0 ;
      RECT  39720.0 65675.0 40425.0 64330.0 ;
      RECT  39720.0 65675.0 40425.0 67020.0 ;
      RECT  39720.0 68365.0 40425.0 67020.0 ;
      RECT  39720.0 68365.0 40425.0 69710.0 ;
      RECT  39720.0 71055.0 40425.0 69710.0 ;
      RECT  39720.0 71055.0 40425.0 72400.0 ;
      RECT  39720.0 73745.0 40425.0 72400.0 ;
      RECT  39720.0 73745.0 40425.0 75090.0 ;
      RECT  39720.0 76435.0 40425.0 75090.0 ;
      RECT  39720.0 76435.0 40425.0 77780.0 ;
      RECT  39720.0 79125.0 40425.0 77780.0 ;
      RECT  39720.0 79125.0 40425.0 80470.0 ;
      RECT  39720.0 81815.0 40425.0 80470.0 ;
      RECT  39720.0 81815.0 40425.0 83160.0 ;
      RECT  39720.0 84505.0 40425.0 83160.0 ;
      RECT  39720.0 84505.0 40425.0 85850.0 ;
      RECT  39720.0 87195.0 40425.0 85850.0 ;
      RECT  39720.0 87195.0 40425.0 88540.0 ;
      RECT  39720.0 89885.0 40425.0 88540.0 ;
      RECT  39720.0 89885.0 40425.0 91230.0 ;
      RECT  39720.0 92575.0 40425.0 91230.0 ;
      RECT  39720.0 92575.0 40425.0 93920.0 ;
      RECT  39720.0 95265.0 40425.0 93920.0 ;
      RECT  39720.0 95265.0 40425.0 96610.0 ;
      RECT  39720.0 97955.0 40425.0 96610.0 ;
      RECT  39720.0 97955.0 40425.0 99300.0 ;
      RECT  39720.0 100645.0 40425.0 99300.0 ;
      RECT  39720.0 100645.0 40425.0 101990.0 ;
      RECT  39720.0 103335.0 40425.0 101990.0 ;
      RECT  39720.0 103335.0 40425.0 104680.0 ;
      RECT  39720.0 106025.0 40425.0 104680.0 ;
      RECT  39720.0 106025.0 40425.0 107370.0 ;
      RECT  39720.0 108715.0 40425.0 107370.0 ;
      RECT  39720.0 108715.0 40425.0 110060.0 ;
      RECT  39720.0 111405.0 40425.0 110060.0 ;
      RECT  39720.0 111405.0 40425.0 112750.0 ;
      RECT  39720.0 114095.0 40425.0 112750.0 ;
      RECT  40425.0 28015.0 41130.0 29360.0 ;
      RECT  40425.0 30705.0 41130.0 29360.0 ;
      RECT  40425.0 30705.0 41130.0 32050.0 ;
      RECT  40425.0 33395.0 41130.0 32050.0 ;
      RECT  40425.0 33395.0 41130.0 34740.0 ;
      RECT  40425.0 36085.0 41130.0 34740.0 ;
      RECT  40425.0 36085.0 41130.0 37430.0 ;
      RECT  40425.0 38775.0 41130.0 37430.0 ;
      RECT  40425.0 38775.0 41130.0 40120.0 ;
      RECT  40425.0 41465.0 41130.0 40120.0 ;
      RECT  40425.0 41465.0 41130.0 42810.0 ;
      RECT  40425.0 44155.0 41130.0 42810.0 ;
      RECT  40425.0 44155.0 41130.0 45500.0 ;
      RECT  40425.0 46845.0 41130.0 45500.0 ;
      RECT  40425.0 46845.0 41130.0 48190.0 ;
      RECT  40425.0 49535.0 41130.0 48190.0 ;
      RECT  40425.0 49535.0 41130.0 50880.0 ;
      RECT  40425.0 52225.0 41130.0 50880.0 ;
      RECT  40425.0 52225.0 41130.0 53570.0 ;
      RECT  40425.0 54915.0 41130.0 53570.0 ;
      RECT  40425.0 54915.0 41130.0 56260.0 ;
      RECT  40425.0 57605.0 41130.0 56260.0 ;
      RECT  40425.0 57605.0 41130.0 58950.0 ;
      RECT  40425.0 60295.0 41130.0 58950.0 ;
      RECT  40425.0 60295.0 41130.0 61640.0 ;
      RECT  40425.0 62985.0 41130.0 61640.0 ;
      RECT  40425.0 62985.0 41130.0 64330.0 ;
      RECT  40425.0 65675.0 41130.0 64330.0 ;
      RECT  40425.0 65675.0 41130.0 67020.0 ;
      RECT  40425.0 68365.0 41130.0 67020.0 ;
      RECT  40425.0 68365.0 41130.0 69710.0 ;
      RECT  40425.0 71055.0 41130.0 69710.0 ;
      RECT  40425.0 71055.0 41130.0 72400.0 ;
      RECT  40425.0 73745.0 41130.0 72400.0 ;
      RECT  40425.0 73745.0 41130.0 75090.0 ;
      RECT  40425.0 76435.0 41130.0 75090.0 ;
      RECT  40425.0 76435.0 41130.0 77780.0 ;
      RECT  40425.0 79125.0 41130.0 77780.0 ;
      RECT  40425.0 79125.0 41130.0 80470.0 ;
      RECT  40425.0 81815.0 41130.0 80470.0 ;
      RECT  40425.0 81815.0 41130.0 83160.0 ;
      RECT  40425.0 84505.0 41130.0 83160.0 ;
      RECT  40425.0 84505.0 41130.0 85850.0 ;
      RECT  40425.0 87195.0 41130.0 85850.0 ;
      RECT  40425.0 87195.0 41130.0 88540.0 ;
      RECT  40425.0 89885.0 41130.0 88540.0 ;
      RECT  40425.0 89885.0 41130.0 91230.0 ;
      RECT  40425.0 92575.0 41130.0 91230.0 ;
      RECT  40425.0 92575.0 41130.0 93920.0 ;
      RECT  40425.0 95265.0 41130.0 93920.0 ;
      RECT  40425.0 95265.0 41130.0 96610.0 ;
      RECT  40425.0 97955.0 41130.0 96610.0 ;
      RECT  40425.0 97955.0 41130.0 99300.0 ;
      RECT  40425.0 100645.0 41130.0 99300.0 ;
      RECT  40425.0 100645.0 41130.0 101990.0 ;
      RECT  40425.0 103335.0 41130.0 101990.0 ;
      RECT  40425.0 103335.0 41130.0 104680.0 ;
      RECT  40425.0 106025.0 41130.0 104680.0 ;
      RECT  40425.0 106025.0 41130.0 107370.0 ;
      RECT  40425.0 108715.0 41130.0 107370.0 ;
      RECT  40425.0 108715.0 41130.0 110060.0 ;
      RECT  40425.0 111405.0 41130.0 110060.0 ;
      RECT  40425.0 111405.0 41130.0 112750.0 ;
      RECT  40425.0 114095.0 41130.0 112750.0 ;
      RECT  41130.0 28015.0 41835.0 29360.0 ;
      RECT  41130.0 30705.0 41835.0 29360.0 ;
      RECT  41130.0 30705.0 41835.0 32050.0 ;
      RECT  41130.0 33395.0 41835.0 32050.0 ;
      RECT  41130.0 33395.0 41835.0 34740.0 ;
      RECT  41130.0 36085.0 41835.0 34740.0 ;
      RECT  41130.0 36085.0 41835.0 37430.0 ;
      RECT  41130.0 38775.0 41835.0 37430.0 ;
      RECT  41130.0 38775.0 41835.0 40120.0 ;
      RECT  41130.0 41465.0 41835.0 40120.0 ;
      RECT  41130.0 41465.0 41835.0 42810.0 ;
      RECT  41130.0 44155.0 41835.0 42810.0 ;
      RECT  41130.0 44155.0 41835.0 45500.0 ;
      RECT  41130.0 46845.0 41835.0 45500.0 ;
      RECT  41130.0 46845.0 41835.0 48190.0 ;
      RECT  41130.0 49535.0 41835.0 48190.0 ;
      RECT  41130.0 49535.0 41835.0 50880.0 ;
      RECT  41130.0 52225.0 41835.0 50880.0 ;
      RECT  41130.0 52225.0 41835.0 53570.0 ;
      RECT  41130.0 54915.0 41835.0 53570.0 ;
      RECT  41130.0 54915.0 41835.0 56260.0 ;
      RECT  41130.0 57605.0 41835.0 56260.0 ;
      RECT  41130.0 57605.0 41835.0 58950.0 ;
      RECT  41130.0 60295.0 41835.0 58950.0 ;
      RECT  41130.0 60295.0 41835.0 61640.0 ;
      RECT  41130.0 62985.0 41835.0 61640.0 ;
      RECT  41130.0 62985.0 41835.0 64330.0 ;
      RECT  41130.0 65675.0 41835.0 64330.0 ;
      RECT  41130.0 65675.0 41835.0 67020.0 ;
      RECT  41130.0 68365.0 41835.0 67020.0 ;
      RECT  41130.0 68365.0 41835.0 69710.0 ;
      RECT  41130.0 71055.0 41835.0 69710.0 ;
      RECT  41130.0 71055.0 41835.0 72400.0 ;
      RECT  41130.0 73745.0 41835.0 72400.0 ;
      RECT  41130.0 73745.0 41835.0 75090.0 ;
      RECT  41130.0 76435.0 41835.0 75090.0 ;
      RECT  41130.0 76435.0 41835.0 77780.0 ;
      RECT  41130.0 79125.0 41835.0 77780.0 ;
      RECT  41130.0 79125.0 41835.0 80470.0 ;
      RECT  41130.0 81815.0 41835.0 80470.0 ;
      RECT  41130.0 81815.0 41835.0 83160.0 ;
      RECT  41130.0 84505.0 41835.0 83160.0 ;
      RECT  41130.0 84505.0 41835.0 85850.0 ;
      RECT  41130.0 87195.0 41835.0 85850.0 ;
      RECT  41130.0 87195.0 41835.0 88540.0 ;
      RECT  41130.0 89885.0 41835.0 88540.0 ;
      RECT  41130.0 89885.0 41835.0 91230.0 ;
      RECT  41130.0 92575.0 41835.0 91230.0 ;
      RECT  41130.0 92575.0 41835.0 93920.0 ;
      RECT  41130.0 95265.0 41835.0 93920.0 ;
      RECT  41130.0 95265.0 41835.0 96610.0 ;
      RECT  41130.0 97955.0 41835.0 96610.0 ;
      RECT  41130.0 97955.0 41835.0 99300.0 ;
      RECT  41130.0 100645.0 41835.0 99300.0 ;
      RECT  41130.0 100645.0 41835.0 101990.0 ;
      RECT  41130.0 103335.0 41835.0 101990.0 ;
      RECT  41130.0 103335.0 41835.0 104680.0 ;
      RECT  41130.0 106025.0 41835.0 104680.0 ;
      RECT  41130.0 106025.0 41835.0 107370.0 ;
      RECT  41130.0 108715.0 41835.0 107370.0 ;
      RECT  41130.0 108715.0 41835.0 110060.0 ;
      RECT  41130.0 111405.0 41835.0 110060.0 ;
      RECT  41130.0 111405.0 41835.0 112750.0 ;
      RECT  41130.0 114095.0 41835.0 112750.0 ;
      RECT  41835.0 28015.0 42540.0 29360.0 ;
      RECT  41835.0 30705.0 42540.0 29360.0 ;
      RECT  41835.0 30705.0 42540.0 32050.0 ;
      RECT  41835.0 33395.0 42540.0 32050.0 ;
      RECT  41835.0 33395.0 42540.0 34740.0 ;
      RECT  41835.0 36085.0 42540.0 34740.0 ;
      RECT  41835.0 36085.0 42540.0 37430.0 ;
      RECT  41835.0 38775.0 42540.0 37430.0 ;
      RECT  41835.0 38775.0 42540.0 40120.0 ;
      RECT  41835.0 41465.0 42540.0 40120.0 ;
      RECT  41835.0 41465.0 42540.0 42810.0 ;
      RECT  41835.0 44155.0 42540.0 42810.0 ;
      RECT  41835.0 44155.0 42540.0 45500.0 ;
      RECT  41835.0 46845.0 42540.0 45500.0 ;
      RECT  41835.0 46845.0 42540.0 48190.0 ;
      RECT  41835.0 49535.0 42540.0 48190.0 ;
      RECT  41835.0 49535.0 42540.0 50880.0 ;
      RECT  41835.0 52225.0 42540.0 50880.0 ;
      RECT  41835.0 52225.0 42540.0 53570.0 ;
      RECT  41835.0 54915.0 42540.0 53570.0 ;
      RECT  41835.0 54915.0 42540.0 56260.0 ;
      RECT  41835.0 57605.0 42540.0 56260.0 ;
      RECT  41835.0 57605.0 42540.0 58950.0 ;
      RECT  41835.0 60295.0 42540.0 58950.0 ;
      RECT  41835.0 60295.0 42540.0 61640.0 ;
      RECT  41835.0 62985.0 42540.0 61640.0 ;
      RECT  41835.0 62985.0 42540.0 64330.0 ;
      RECT  41835.0 65675.0 42540.0 64330.0 ;
      RECT  41835.0 65675.0 42540.0 67020.0 ;
      RECT  41835.0 68365.0 42540.0 67020.0 ;
      RECT  41835.0 68365.0 42540.0 69710.0 ;
      RECT  41835.0 71055.0 42540.0 69710.0 ;
      RECT  41835.0 71055.0 42540.0 72400.0 ;
      RECT  41835.0 73745.0 42540.0 72400.0 ;
      RECT  41835.0 73745.0 42540.0 75090.0 ;
      RECT  41835.0 76435.0 42540.0 75090.0 ;
      RECT  41835.0 76435.0 42540.0 77780.0 ;
      RECT  41835.0 79125.0 42540.0 77780.0 ;
      RECT  41835.0 79125.0 42540.0 80470.0 ;
      RECT  41835.0 81815.0 42540.0 80470.0 ;
      RECT  41835.0 81815.0 42540.0 83160.0 ;
      RECT  41835.0 84505.0 42540.0 83160.0 ;
      RECT  41835.0 84505.0 42540.0 85850.0 ;
      RECT  41835.0 87195.0 42540.0 85850.0 ;
      RECT  41835.0 87195.0 42540.0 88540.0 ;
      RECT  41835.0 89885.0 42540.0 88540.0 ;
      RECT  41835.0 89885.0 42540.0 91230.0 ;
      RECT  41835.0 92575.0 42540.0 91230.0 ;
      RECT  41835.0 92575.0 42540.0 93920.0 ;
      RECT  41835.0 95265.0 42540.0 93920.0 ;
      RECT  41835.0 95265.0 42540.0 96610.0 ;
      RECT  41835.0 97955.0 42540.0 96610.0 ;
      RECT  41835.0 97955.0 42540.0 99300.0 ;
      RECT  41835.0 100645.0 42540.0 99300.0 ;
      RECT  41835.0 100645.0 42540.0 101990.0 ;
      RECT  41835.0 103335.0 42540.0 101990.0 ;
      RECT  41835.0 103335.0 42540.0 104680.0 ;
      RECT  41835.0 106025.0 42540.0 104680.0 ;
      RECT  41835.0 106025.0 42540.0 107370.0 ;
      RECT  41835.0 108715.0 42540.0 107370.0 ;
      RECT  41835.0 108715.0 42540.0 110060.0 ;
      RECT  41835.0 111405.0 42540.0 110060.0 ;
      RECT  41835.0 111405.0 42540.0 112750.0 ;
      RECT  41835.0 114095.0 42540.0 112750.0 ;
      RECT  42540.0 28015.0 43245.0 29360.0 ;
      RECT  42540.0 30705.0 43245.0 29360.0 ;
      RECT  42540.0 30705.0 43245.0 32050.0 ;
      RECT  42540.0 33395.0 43245.0 32050.0 ;
      RECT  42540.0 33395.0 43245.0 34740.0 ;
      RECT  42540.0 36085.0 43245.0 34740.0 ;
      RECT  42540.0 36085.0 43245.0 37430.0 ;
      RECT  42540.0 38775.0 43245.0 37430.0 ;
      RECT  42540.0 38775.0 43245.0 40120.0 ;
      RECT  42540.0 41465.0 43245.0 40120.0 ;
      RECT  42540.0 41465.0 43245.0 42810.0 ;
      RECT  42540.0 44155.0 43245.0 42810.0 ;
      RECT  42540.0 44155.0 43245.0 45500.0 ;
      RECT  42540.0 46845.0 43245.0 45500.0 ;
      RECT  42540.0 46845.0 43245.0 48190.0 ;
      RECT  42540.0 49535.0 43245.0 48190.0 ;
      RECT  42540.0 49535.0 43245.0 50880.0 ;
      RECT  42540.0 52225.0 43245.0 50880.0 ;
      RECT  42540.0 52225.0 43245.0 53570.0 ;
      RECT  42540.0 54915.0 43245.0 53570.0 ;
      RECT  42540.0 54915.0 43245.0 56260.0 ;
      RECT  42540.0 57605.0 43245.0 56260.0 ;
      RECT  42540.0 57605.0 43245.0 58950.0 ;
      RECT  42540.0 60295.0 43245.0 58950.0 ;
      RECT  42540.0 60295.0 43245.0 61640.0 ;
      RECT  42540.0 62985.0 43245.0 61640.0 ;
      RECT  42540.0 62985.0 43245.0 64330.0 ;
      RECT  42540.0 65675.0 43245.0 64330.0 ;
      RECT  42540.0 65675.0 43245.0 67020.0 ;
      RECT  42540.0 68365.0 43245.0 67020.0 ;
      RECT  42540.0 68365.0 43245.0 69710.0 ;
      RECT  42540.0 71055.0 43245.0 69710.0 ;
      RECT  42540.0 71055.0 43245.0 72400.0 ;
      RECT  42540.0 73745.0 43245.0 72400.0 ;
      RECT  42540.0 73745.0 43245.0 75090.0 ;
      RECT  42540.0 76435.0 43245.0 75090.0 ;
      RECT  42540.0 76435.0 43245.0 77780.0 ;
      RECT  42540.0 79125.0 43245.0 77780.0 ;
      RECT  42540.0 79125.0 43245.0 80470.0 ;
      RECT  42540.0 81815.0 43245.0 80470.0 ;
      RECT  42540.0 81815.0 43245.0 83160.0 ;
      RECT  42540.0 84505.0 43245.0 83160.0 ;
      RECT  42540.0 84505.0 43245.0 85850.0 ;
      RECT  42540.0 87195.0 43245.0 85850.0 ;
      RECT  42540.0 87195.0 43245.0 88540.0 ;
      RECT  42540.0 89885.0 43245.0 88540.0 ;
      RECT  42540.0 89885.0 43245.0 91230.0 ;
      RECT  42540.0 92575.0 43245.0 91230.0 ;
      RECT  42540.0 92575.0 43245.0 93920.0 ;
      RECT  42540.0 95265.0 43245.0 93920.0 ;
      RECT  42540.0 95265.0 43245.0 96610.0 ;
      RECT  42540.0 97955.0 43245.0 96610.0 ;
      RECT  42540.0 97955.0 43245.0 99300.0 ;
      RECT  42540.0 100645.0 43245.0 99300.0 ;
      RECT  42540.0 100645.0 43245.0 101990.0 ;
      RECT  42540.0 103335.0 43245.0 101990.0 ;
      RECT  42540.0 103335.0 43245.0 104680.0 ;
      RECT  42540.0 106025.0 43245.0 104680.0 ;
      RECT  42540.0 106025.0 43245.0 107370.0 ;
      RECT  42540.0 108715.0 43245.0 107370.0 ;
      RECT  42540.0 108715.0 43245.0 110060.0 ;
      RECT  42540.0 111405.0 43245.0 110060.0 ;
      RECT  42540.0 111405.0 43245.0 112750.0 ;
      RECT  42540.0 114095.0 43245.0 112750.0 ;
      RECT  43245.0 28015.0 43950.0 29360.0 ;
      RECT  43245.0 30705.0 43950.0 29360.0 ;
      RECT  43245.0 30705.0 43950.0 32050.0 ;
      RECT  43245.0 33395.0 43950.0 32050.0 ;
      RECT  43245.0 33395.0 43950.0 34740.0 ;
      RECT  43245.0 36085.0 43950.0 34740.0 ;
      RECT  43245.0 36085.0 43950.0 37430.0 ;
      RECT  43245.0 38775.0 43950.0 37430.0 ;
      RECT  43245.0 38775.0 43950.0 40120.0 ;
      RECT  43245.0 41465.0 43950.0 40120.0 ;
      RECT  43245.0 41465.0 43950.0 42810.0 ;
      RECT  43245.0 44155.0 43950.0 42810.0 ;
      RECT  43245.0 44155.0 43950.0 45500.0 ;
      RECT  43245.0 46845.0 43950.0 45500.0 ;
      RECT  43245.0 46845.0 43950.0 48190.0 ;
      RECT  43245.0 49535.0 43950.0 48190.0 ;
      RECT  43245.0 49535.0 43950.0 50880.0 ;
      RECT  43245.0 52225.0 43950.0 50880.0 ;
      RECT  43245.0 52225.0 43950.0 53570.0 ;
      RECT  43245.0 54915.0 43950.0 53570.0 ;
      RECT  43245.0 54915.0 43950.0 56260.0 ;
      RECT  43245.0 57605.0 43950.0 56260.0 ;
      RECT  43245.0 57605.0 43950.0 58950.0 ;
      RECT  43245.0 60295.0 43950.0 58950.0 ;
      RECT  43245.0 60295.0 43950.0 61640.0 ;
      RECT  43245.0 62985.0 43950.0 61640.0 ;
      RECT  43245.0 62985.0 43950.0 64330.0 ;
      RECT  43245.0 65675.0 43950.0 64330.0 ;
      RECT  43245.0 65675.0 43950.0 67020.0 ;
      RECT  43245.0 68365.0 43950.0 67020.0 ;
      RECT  43245.0 68365.0 43950.0 69710.0 ;
      RECT  43245.0 71055.0 43950.0 69710.0 ;
      RECT  43245.0 71055.0 43950.0 72400.0 ;
      RECT  43245.0 73745.0 43950.0 72400.0 ;
      RECT  43245.0 73745.0 43950.0 75090.0 ;
      RECT  43245.0 76435.0 43950.0 75090.0 ;
      RECT  43245.0 76435.0 43950.0 77780.0 ;
      RECT  43245.0 79125.0 43950.0 77780.0 ;
      RECT  43245.0 79125.0 43950.0 80470.0 ;
      RECT  43245.0 81815.0 43950.0 80470.0 ;
      RECT  43245.0 81815.0 43950.0 83160.0 ;
      RECT  43245.0 84505.0 43950.0 83160.0 ;
      RECT  43245.0 84505.0 43950.0 85850.0 ;
      RECT  43245.0 87195.0 43950.0 85850.0 ;
      RECT  43245.0 87195.0 43950.0 88540.0 ;
      RECT  43245.0 89885.0 43950.0 88540.0 ;
      RECT  43245.0 89885.0 43950.0 91230.0 ;
      RECT  43245.0 92575.0 43950.0 91230.0 ;
      RECT  43245.0 92575.0 43950.0 93920.0 ;
      RECT  43245.0 95265.0 43950.0 93920.0 ;
      RECT  43245.0 95265.0 43950.0 96610.0 ;
      RECT  43245.0 97955.0 43950.0 96610.0 ;
      RECT  43245.0 97955.0 43950.0 99300.0 ;
      RECT  43245.0 100645.0 43950.0 99300.0 ;
      RECT  43245.0 100645.0 43950.0 101990.0 ;
      RECT  43245.0 103335.0 43950.0 101990.0 ;
      RECT  43245.0 103335.0 43950.0 104680.0 ;
      RECT  43245.0 106025.0 43950.0 104680.0 ;
      RECT  43245.0 106025.0 43950.0 107370.0 ;
      RECT  43245.0 108715.0 43950.0 107370.0 ;
      RECT  43245.0 108715.0 43950.0 110060.0 ;
      RECT  43245.0 111405.0 43950.0 110060.0 ;
      RECT  43245.0 111405.0 43950.0 112750.0 ;
      RECT  43245.0 114095.0 43950.0 112750.0 ;
      RECT  43950.0 28015.0 44655.0 29360.0 ;
      RECT  43950.0 30705.0 44655.0 29360.0 ;
      RECT  43950.0 30705.0 44655.0 32050.0 ;
      RECT  43950.0 33395.0 44655.0 32050.0 ;
      RECT  43950.0 33395.0 44655.0 34740.0 ;
      RECT  43950.0 36085.0 44655.0 34740.0 ;
      RECT  43950.0 36085.0 44655.0 37430.0 ;
      RECT  43950.0 38775.0 44655.0 37430.0 ;
      RECT  43950.0 38775.0 44655.0 40120.0 ;
      RECT  43950.0 41465.0 44655.0 40120.0 ;
      RECT  43950.0 41465.0 44655.0 42810.0 ;
      RECT  43950.0 44155.0 44655.0 42810.0 ;
      RECT  43950.0 44155.0 44655.0 45500.0 ;
      RECT  43950.0 46845.0 44655.0 45500.0 ;
      RECT  43950.0 46845.0 44655.0 48190.0 ;
      RECT  43950.0 49535.0 44655.0 48190.0 ;
      RECT  43950.0 49535.0 44655.0 50880.0 ;
      RECT  43950.0 52225.0 44655.0 50880.0 ;
      RECT  43950.0 52225.0 44655.0 53570.0 ;
      RECT  43950.0 54915.0 44655.0 53570.0 ;
      RECT  43950.0 54915.0 44655.0 56260.0 ;
      RECT  43950.0 57605.0 44655.0 56260.0 ;
      RECT  43950.0 57605.0 44655.0 58950.0 ;
      RECT  43950.0 60295.0 44655.0 58950.0 ;
      RECT  43950.0 60295.0 44655.0 61640.0 ;
      RECT  43950.0 62985.0 44655.0 61640.0 ;
      RECT  43950.0 62985.0 44655.0 64330.0 ;
      RECT  43950.0 65675.0 44655.0 64330.0 ;
      RECT  43950.0 65675.0 44655.0 67020.0 ;
      RECT  43950.0 68365.0 44655.0 67020.0 ;
      RECT  43950.0 68365.0 44655.0 69710.0 ;
      RECT  43950.0 71055.0 44655.0 69710.0 ;
      RECT  43950.0 71055.0 44655.0 72400.0 ;
      RECT  43950.0 73745.0 44655.0 72400.0 ;
      RECT  43950.0 73745.0 44655.0 75090.0 ;
      RECT  43950.0 76435.0 44655.0 75090.0 ;
      RECT  43950.0 76435.0 44655.0 77780.0 ;
      RECT  43950.0 79125.0 44655.0 77780.0 ;
      RECT  43950.0 79125.0 44655.0 80470.0 ;
      RECT  43950.0 81815.0 44655.0 80470.0 ;
      RECT  43950.0 81815.0 44655.0 83160.0 ;
      RECT  43950.0 84505.0 44655.0 83160.0 ;
      RECT  43950.0 84505.0 44655.0 85850.0 ;
      RECT  43950.0 87195.0 44655.0 85850.0 ;
      RECT  43950.0 87195.0 44655.0 88540.0 ;
      RECT  43950.0 89885.0 44655.0 88540.0 ;
      RECT  43950.0 89885.0 44655.0 91230.0 ;
      RECT  43950.0 92575.0 44655.0 91230.0 ;
      RECT  43950.0 92575.0 44655.0 93920.0 ;
      RECT  43950.0 95265.0 44655.0 93920.0 ;
      RECT  43950.0 95265.0 44655.0 96610.0 ;
      RECT  43950.0 97955.0 44655.0 96610.0 ;
      RECT  43950.0 97955.0 44655.0 99300.0 ;
      RECT  43950.0 100645.0 44655.0 99300.0 ;
      RECT  43950.0 100645.0 44655.0 101990.0 ;
      RECT  43950.0 103335.0 44655.0 101990.0 ;
      RECT  43950.0 103335.0 44655.0 104680.0 ;
      RECT  43950.0 106025.0 44655.0 104680.0 ;
      RECT  43950.0 106025.0 44655.0 107370.0 ;
      RECT  43950.0 108715.0 44655.0 107370.0 ;
      RECT  43950.0 108715.0 44655.0 110060.0 ;
      RECT  43950.0 111405.0 44655.0 110060.0 ;
      RECT  43950.0 111405.0 44655.0 112750.0 ;
      RECT  43950.0 114095.0 44655.0 112750.0 ;
      RECT  44655.0 28015.0 45360.0 29360.0 ;
      RECT  44655.0 30705.0 45360.0 29360.0 ;
      RECT  44655.0 30705.0 45360.0 32050.0 ;
      RECT  44655.0 33395.0 45360.0 32050.0 ;
      RECT  44655.0 33395.0 45360.0 34740.0 ;
      RECT  44655.0 36085.0 45360.0 34740.0 ;
      RECT  44655.0 36085.0 45360.0 37430.0 ;
      RECT  44655.0 38775.0 45360.0 37430.0 ;
      RECT  44655.0 38775.0 45360.0 40120.0 ;
      RECT  44655.0 41465.0 45360.0 40120.0 ;
      RECT  44655.0 41465.0 45360.0 42810.0 ;
      RECT  44655.0 44155.0 45360.0 42810.0 ;
      RECT  44655.0 44155.0 45360.0 45500.0 ;
      RECT  44655.0 46845.0 45360.0 45500.0 ;
      RECT  44655.0 46845.0 45360.0 48190.0 ;
      RECT  44655.0 49535.0 45360.0 48190.0 ;
      RECT  44655.0 49535.0 45360.0 50880.0 ;
      RECT  44655.0 52225.0 45360.0 50880.0 ;
      RECT  44655.0 52225.0 45360.0 53570.0 ;
      RECT  44655.0 54915.0 45360.0 53570.0 ;
      RECT  44655.0 54915.0 45360.0 56260.0 ;
      RECT  44655.0 57605.0 45360.0 56260.0 ;
      RECT  44655.0 57605.0 45360.0 58950.0 ;
      RECT  44655.0 60295.0 45360.0 58950.0 ;
      RECT  44655.0 60295.0 45360.0 61640.0 ;
      RECT  44655.0 62985.0 45360.0 61640.0 ;
      RECT  44655.0 62985.0 45360.0 64330.0 ;
      RECT  44655.0 65675.0 45360.0 64330.0 ;
      RECT  44655.0 65675.0 45360.0 67020.0 ;
      RECT  44655.0 68365.0 45360.0 67020.0 ;
      RECT  44655.0 68365.0 45360.0 69710.0 ;
      RECT  44655.0 71055.0 45360.0 69710.0 ;
      RECT  44655.0 71055.0 45360.0 72400.0 ;
      RECT  44655.0 73745.0 45360.0 72400.0 ;
      RECT  44655.0 73745.0 45360.0 75090.0 ;
      RECT  44655.0 76435.0 45360.0 75090.0 ;
      RECT  44655.0 76435.0 45360.0 77780.0 ;
      RECT  44655.0 79125.0 45360.0 77780.0 ;
      RECT  44655.0 79125.0 45360.0 80470.0 ;
      RECT  44655.0 81815.0 45360.0 80470.0 ;
      RECT  44655.0 81815.0 45360.0 83160.0 ;
      RECT  44655.0 84505.0 45360.0 83160.0 ;
      RECT  44655.0 84505.0 45360.0 85850.0 ;
      RECT  44655.0 87195.0 45360.0 85850.0 ;
      RECT  44655.0 87195.0 45360.0 88540.0 ;
      RECT  44655.0 89885.0 45360.0 88540.0 ;
      RECT  44655.0 89885.0 45360.0 91230.0 ;
      RECT  44655.0 92575.0 45360.0 91230.0 ;
      RECT  44655.0 92575.0 45360.0 93920.0 ;
      RECT  44655.0 95265.0 45360.0 93920.0 ;
      RECT  44655.0 95265.0 45360.0 96610.0 ;
      RECT  44655.0 97955.0 45360.0 96610.0 ;
      RECT  44655.0 97955.0 45360.0 99300.0 ;
      RECT  44655.0 100645.0 45360.0 99300.0 ;
      RECT  44655.0 100645.0 45360.0 101990.0 ;
      RECT  44655.0 103335.0 45360.0 101990.0 ;
      RECT  44655.0 103335.0 45360.0 104680.0 ;
      RECT  44655.0 106025.0 45360.0 104680.0 ;
      RECT  44655.0 106025.0 45360.0 107370.0 ;
      RECT  44655.0 108715.0 45360.0 107370.0 ;
      RECT  44655.0 108715.0 45360.0 110060.0 ;
      RECT  44655.0 111405.0 45360.0 110060.0 ;
      RECT  44655.0 111405.0 45360.0 112750.0 ;
      RECT  44655.0 114095.0 45360.0 112750.0 ;
      RECT  45360.0 28015.0 46065.0 29360.0 ;
      RECT  45360.0 30705.0 46065.0 29360.0 ;
      RECT  45360.0 30705.0 46065.0 32050.0 ;
      RECT  45360.0 33395.0 46065.0 32050.0 ;
      RECT  45360.0 33395.0 46065.0 34740.0 ;
      RECT  45360.0 36085.0 46065.0 34740.0 ;
      RECT  45360.0 36085.0 46065.0 37430.0 ;
      RECT  45360.0 38775.0 46065.0 37430.0 ;
      RECT  45360.0 38775.0 46065.0 40120.0 ;
      RECT  45360.0 41465.0 46065.0 40120.0 ;
      RECT  45360.0 41465.0 46065.0 42810.0 ;
      RECT  45360.0 44155.0 46065.0 42810.0 ;
      RECT  45360.0 44155.0 46065.0 45500.0 ;
      RECT  45360.0 46845.0 46065.0 45500.0 ;
      RECT  45360.0 46845.0 46065.0 48190.0 ;
      RECT  45360.0 49535.0 46065.0 48190.0 ;
      RECT  45360.0 49535.0 46065.0 50880.0 ;
      RECT  45360.0 52225.0 46065.0 50880.0 ;
      RECT  45360.0 52225.0 46065.0 53570.0 ;
      RECT  45360.0 54915.0 46065.0 53570.0 ;
      RECT  45360.0 54915.0 46065.0 56260.0 ;
      RECT  45360.0 57605.0 46065.0 56260.0 ;
      RECT  45360.0 57605.0 46065.0 58950.0 ;
      RECT  45360.0 60295.0 46065.0 58950.0 ;
      RECT  45360.0 60295.0 46065.0 61640.0 ;
      RECT  45360.0 62985.0 46065.0 61640.0 ;
      RECT  45360.0 62985.0 46065.0 64330.0 ;
      RECT  45360.0 65675.0 46065.0 64330.0 ;
      RECT  45360.0 65675.0 46065.0 67020.0 ;
      RECT  45360.0 68365.0 46065.0 67020.0 ;
      RECT  45360.0 68365.0 46065.0 69710.0 ;
      RECT  45360.0 71055.0 46065.0 69710.0 ;
      RECT  45360.0 71055.0 46065.0 72400.0 ;
      RECT  45360.0 73745.0 46065.0 72400.0 ;
      RECT  45360.0 73745.0 46065.0 75090.0 ;
      RECT  45360.0 76435.0 46065.0 75090.0 ;
      RECT  45360.0 76435.0 46065.0 77780.0 ;
      RECT  45360.0 79125.0 46065.0 77780.0 ;
      RECT  45360.0 79125.0 46065.0 80470.0 ;
      RECT  45360.0 81815.0 46065.0 80470.0 ;
      RECT  45360.0 81815.0 46065.0 83160.0 ;
      RECT  45360.0 84505.0 46065.0 83160.0 ;
      RECT  45360.0 84505.0 46065.0 85850.0 ;
      RECT  45360.0 87195.0 46065.0 85850.0 ;
      RECT  45360.0 87195.0 46065.0 88540.0 ;
      RECT  45360.0 89885.0 46065.0 88540.0 ;
      RECT  45360.0 89885.0 46065.0 91230.0 ;
      RECT  45360.0 92575.0 46065.0 91230.0 ;
      RECT  45360.0 92575.0 46065.0 93920.0 ;
      RECT  45360.0 95265.0 46065.0 93920.0 ;
      RECT  45360.0 95265.0 46065.0 96610.0 ;
      RECT  45360.0 97955.0 46065.0 96610.0 ;
      RECT  45360.0 97955.0 46065.0 99300.0 ;
      RECT  45360.0 100645.0 46065.0 99300.0 ;
      RECT  45360.0 100645.0 46065.0 101990.0 ;
      RECT  45360.0 103335.0 46065.0 101990.0 ;
      RECT  45360.0 103335.0 46065.0 104680.0 ;
      RECT  45360.0 106025.0 46065.0 104680.0 ;
      RECT  45360.0 106025.0 46065.0 107370.0 ;
      RECT  45360.0 108715.0 46065.0 107370.0 ;
      RECT  45360.0 108715.0 46065.0 110060.0 ;
      RECT  45360.0 111405.0 46065.0 110060.0 ;
      RECT  45360.0 111405.0 46065.0 112750.0 ;
      RECT  45360.0 114095.0 46065.0 112750.0 ;
      RECT  46065.0 28015.0 46770.0 29360.0 ;
      RECT  46065.0 30705.0 46770.0 29360.0 ;
      RECT  46065.0 30705.0 46770.0 32050.0 ;
      RECT  46065.0 33395.0 46770.0 32050.0 ;
      RECT  46065.0 33395.0 46770.0 34740.0 ;
      RECT  46065.0 36085.0 46770.0 34740.0 ;
      RECT  46065.0 36085.0 46770.0 37430.0 ;
      RECT  46065.0 38775.0 46770.0 37430.0 ;
      RECT  46065.0 38775.0 46770.0 40120.0 ;
      RECT  46065.0 41465.0 46770.0 40120.0 ;
      RECT  46065.0 41465.0 46770.0 42810.0 ;
      RECT  46065.0 44155.0 46770.0 42810.0 ;
      RECT  46065.0 44155.0 46770.0 45500.0 ;
      RECT  46065.0 46845.0 46770.0 45500.0 ;
      RECT  46065.0 46845.0 46770.0 48190.0 ;
      RECT  46065.0 49535.0 46770.0 48190.0 ;
      RECT  46065.0 49535.0 46770.0 50880.0 ;
      RECT  46065.0 52225.0 46770.0 50880.0 ;
      RECT  46065.0 52225.0 46770.0 53570.0 ;
      RECT  46065.0 54915.0 46770.0 53570.0 ;
      RECT  46065.0 54915.0 46770.0 56260.0 ;
      RECT  46065.0 57605.0 46770.0 56260.0 ;
      RECT  46065.0 57605.0 46770.0 58950.0 ;
      RECT  46065.0 60295.0 46770.0 58950.0 ;
      RECT  46065.0 60295.0 46770.0 61640.0 ;
      RECT  46065.0 62985.0 46770.0 61640.0 ;
      RECT  46065.0 62985.0 46770.0 64330.0 ;
      RECT  46065.0 65675.0 46770.0 64330.0 ;
      RECT  46065.0 65675.0 46770.0 67020.0 ;
      RECT  46065.0 68365.0 46770.0 67020.0 ;
      RECT  46065.0 68365.0 46770.0 69710.0 ;
      RECT  46065.0 71055.0 46770.0 69710.0 ;
      RECT  46065.0 71055.0 46770.0 72400.0 ;
      RECT  46065.0 73745.0 46770.0 72400.0 ;
      RECT  46065.0 73745.0 46770.0 75090.0 ;
      RECT  46065.0 76435.0 46770.0 75090.0 ;
      RECT  46065.0 76435.0 46770.0 77780.0 ;
      RECT  46065.0 79125.0 46770.0 77780.0 ;
      RECT  46065.0 79125.0 46770.0 80470.0 ;
      RECT  46065.0 81815.0 46770.0 80470.0 ;
      RECT  46065.0 81815.0 46770.0 83160.0 ;
      RECT  46065.0 84505.0 46770.0 83160.0 ;
      RECT  46065.0 84505.0 46770.0 85850.0 ;
      RECT  46065.0 87195.0 46770.0 85850.0 ;
      RECT  46065.0 87195.0 46770.0 88540.0 ;
      RECT  46065.0 89885.0 46770.0 88540.0 ;
      RECT  46065.0 89885.0 46770.0 91230.0 ;
      RECT  46065.0 92575.0 46770.0 91230.0 ;
      RECT  46065.0 92575.0 46770.0 93920.0 ;
      RECT  46065.0 95265.0 46770.0 93920.0 ;
      RECT  46065.0 95265.0 46770.0 96610.0 ;
      RECT  46065.0 97955.0 46770.0 96610.0 ;
      RECT  46065.0 97955.0 46770.0 99300.0 ;
      RECT  46065.0 100645.0 46770.0 99300.0 ;
      RECT  46065.0 100645.0 46770.0 101990.0 ;
      RECT  46065.0 103335.0 46770.0 101990.0 ;
      RECT  46065.0 103335.0 46770.0 104680.0 ;
      RECT  46065.0 106025.0 46770.0 104680.0 ;
      RECT  46065.0 106025.0 46770.0 107370.0 ;
      RECT  46065.0 108715.0 46770.0 107370.0 ;
      RECT  46065.0 108715.0 46770.0 110060.0 ;
      RECT  46065.0 111405.0 46770.0 110060.0 ;
      RECT  46065.0 111405.0 46770.0 112750.0 ;
      RECT  46065.0 114095.0 46770.0 112750.0 ;
      RECT  46770.0 28015.0 47475.0 29360.0 ;
      RECT  46770.0 30705.0 47475.0 29360.0 ;
      RECT  46770.0 30705.0 47475.0 32050.0 ;
      RECT  46770.0 33395.0 47475.0 32050.0 ;
      RECT  46770.0 33395.0 47475.0 34740.0 ;
      RECT  46770.0 36085.0 47475.0 34740.0 ;
      RECT  46770.0 36085.0 47475.0 37430.0 ;
      RECT  46770.0 38775.0 47475.0 37430.0 ;
      RECT  46770.0 38775.0 47475.0 40120.0 ;
      RECT  46770.0 41465.0 47475.0 40120.0 ;
      RECT  46770.0 41465.0 47475.0 42810.0 ;
      RECT  46770.0 44155.0 47475.0 42810.0 ;
      RECT  46770.0 44155.0 47475.0 45500.0 ;
      RECT  46770.0 46845.0 47475.0 45500.0 ;
      RECT  46770.0 46845.0 47475.0 48190.0 ;
      RECT  46770.0 49535.0 47475.0 48190.0 ;
      RECT  46770.0 49535.0 47475.0 50880.0 ;
      RECT  46770.0 52225.0 47475.0 50880.0 ;
      RECT  46770.0 52225.0 47475.0 53570.0 ;
      RECT  46770.0 54915.0 47475.0 53570.0 ;
      RECT  46770.0 54915.0 47475.0 56260.0 ;
      RECT  46770.0 57605.0 47475.0 56260.0 ;
      RECT  46770.0 57605.0 47475.0 58950.0 ;
      RECT  46770.0 60295.0 47475.0 58950.0 ;
      RECT  46770.0 60295.0 47475.0 61640.0 ;
      RECT  46770.0 62985.0 47475.0 61640.0 ;
      RECT  46770.0 62985.0 47475.0 64330.0 ;
      RECT  46770.0 65675.0 47475.0 64330.0 ;
      RECT  46770.0 65675.0 47475.0 67020.0 ;
      RECT  46770.0 68365.0 47475.0 67020.0 ;
      RECT  46770.0 68365.0 47475.0 69710.0 ;
      RECT  46770.0 71055.0 47475.0 69710.0 ;
      RECT  46770.0 71055.0 47475.0 72400.0 ;
      RECT  46770.0 73745.0 47475.0 72400.0 ;
      RECT  46770.0 73745.0 47475.0 75090.0 ;
      RECT  46770.0 76435.0 47475.0 75090.0 ;
      RECT  46770.0 76435.0 47475.0 77780.0 ;
      RECT  46770.0 79125.0 47475.0 77780.0 ;
      RECT  46770.0 79125.0 47475.0 80470.0 ;
      RECT  46770.0 81815.0 47475.0 80470.0 ;
      RECT  46770.0 81815.0 47475.0 83160.0 ;
      RECT  46770.0 84505.0 47475.0 83160.0 ;
      RECT  46770.0 84505.0 47475.0 85850.0 ;
      RECT  46770.0 87195.0 47475.0 85850.0 ;
      RECT  46770.0 87195.0 47475.0 88540.0 ;
      RECT  46770.0 89885.0 47475.0 88540.0 ;
      RECT  46770.0 89885.0 47475.0 91230.0 ;
      RECT  46770.0 92575.0 47475.0 91230.0 ;
      RECT  46770.0 92575.0 47475.0 93920.0 ;
      RECT  46770.0 95265.0 47475.0 93920.0 ;
      RECT  46770.0 95265.0 47475.0 96610.0 ;
      RECT  46770.0 97955.0 47475.0 96610.0 ;
      RECT  46770.0 97955.0 47475.0 99300.0 ;
      RECT  46770.0 100645.0 47475.0 99300.0 ;
      RECT  46770.0 100645.0 47475.0 101990.0 ;
      RECT  46770.0 103335.0 47475.0 101990.0 ;
      RECT  46770.0 103335.0 47475.0 104680.0 ;
      RECT  46770.0 106025.0 47475.0 104680.0 ;
      RECT  46770.0 106025.0 47475.0 107370.0 ;
      RECT  46770.0 108715.0 47475.0 107370.0 ;
      RECT  46770.0 108715.0 47475.0 110060.0 ;
      RECT  46770.0 111405.0 47475.0 110060.0 ;
      RECT  46770.0 111405.0 47475.0 112750.0 ;
      RECT  46770.0 114095.0 47475.0 112750.0 ;
      RECT  47475.0 28015.0 48180.0 29360.0 ;
      RECT  47475.0 30705.0 48180.0 29360.0 ;
      RECT  47475.0 30705.0 48180.0 32050.0 ;
      RECT  47475.0 33395.0 48180.0 32050.0 ;
      RECT  47475.0 33395.0 48180.0 34740.0 ;
      RECT  47475.0 36085.0 48180.0 34740.0 ;
      RECT  47475.0 36085.0 48180.0 37430.0 ;
      RECT  47475.0 38775.0 48180.0 37430.0 ;
      RECT  47475.0 38775.0 48180.0 40120.0 ;
      RECT  47475.0 41465.0 48180.0 40120.0 ;
      RECT  47475.0 41465.0 48180.0 42810.0 ;
      RECT  47475.0 44155.0 48180.0 42810.0 ;
      RECT  47475.0 44155.0 48180.0 45500.0 ;
      RECT  47475.0 46845.0 48180.0 45500.0 ;
      RECT  47475.0 46845.0 48180.0 48190.0 ;
      RECT  47475.0 49535.0 48180.0 48190.0 ;
      RECT  47475.0 49535.0 48180.0 50880.0 ;
      RECT  47475.0 52225.0 48180.0 50880.0 ;
      RECT  47475.0 52225.0 48180.0 53570.0 ;
      RECT  47475.0 54915.0 48180.0 53570.0 ;
      RECT  47475.0 54915.0 48180.0 56260.0 ;
      RECT  47475.0 57605.0 48180.0 56260.0 ;
      RECT  47475.0 57605.0 48180.0 58950.0 ;
      RECT  47475.0 60295.0 48180.0 58950.0 ;
      RECT  47475.0 60295.0 48180.0 61640.0 ;
      RECT  47475.0 62985.0 48180.0 61640.0 ;
      RECT  47475.0 62985.0 48180.0 64330.0 ;
      RECT  47475.0 65675.0 48180.0 64330.0 ;
      RECT  47475.0 65675.0 48180.0 67020.0 ;
      RECT  47475.0 68365.0 48180.0 67020.0 ;
      RECT  47475.0 68365.0 48180.0 69710.0 ;
      RECT  47475.0 71055.0 48180.0 69710.0 ;
      RECT  47475.0 71055.0 48180.0 72400.0 ;
      RECT  47475.0 73745.0 48180.0 72400.0 ;
      RECT  47475.0 73745.0 48180.0 75090.0 ;
      RECT  47475.0 76435.0 48180.0 75090.0 ;
      RECT  47475.0 76435.0 48180.0 77780.0 ;
      RECT  47475.0 79125.0 48180.0 77780.0 ;
      RECT  47475.0 79125.0 48180.0 80470.0 ;
      RECT  47475.0 81815.0 48180.0 80470.0 ;
      RECT  47475.0 81815.0 48180.0 83160.0 ;
      RECT  47475.0 84505.0 48180.0 83160.0 ;
      RECT  47475.0 84505.0 48180.0 85850.0 ;
      RECT  47475.0 87195.0 48180.0 85850.0 ;
      RECT  47475.0 87195.0 48180.0 88540.0 ;
      RECT  47475.0 89885.0 48180.0 88540.0 ;
      RECT  47475.0 89885.0 48180.0 91230.0 ;
      RECT  47475.0 92575.0 48180.0 91230.0 ;
      RECT  47475.0 92575.0 48180.0 93920.0 ;
      RECT  47475.0 95265.0 48180.0 93920.0 ;
      RECT  47475.0 95265.0 48180.0 96610.0 ;
      RECT  47475.0 97955.0 48180.0 96610.0 ;
      RECT  47475.0 97955.0 48180.0 99300.0 ;
      RECT  47475.0 100645.0 48180.0 99300.0 ;
      RECT  47475.0 100645.0 48180.0 101990.0 ;
      RECT  47475.0 103335.0 48180.0 101990.0 ;
      RECT  47475.0 103335.0 48180.0 104680.0 ;
      RECT  47475.0 106025.0 48180.0 104680.0 ;
      RECT  47475.0 106025.0 48180.0 107370.0 ;
      RECT  47475.0 108715.0 48180.0 107370.0 ;
      RECT  47475.0 108715.0 48180.0 110060.0 ;
      RECT  47475.0 111405.0 48180.0 110060.0 ;
      RECT  47475.0 111405.0 48180.0 112750.0 ;
      RECT  47475.0 114095.0 48180.0 112750.0 ;
      RECT  48180.0 28015.0 48885.0 29360.0 ;
      RECT  48180.0 30705.0 48885.0 29360.0 ;
      RECT  48180.0 30705.0 48885.0 32050.0 ;
      RECT  48180.0 33395.0 48885.0 32050.0 ;
      RECT  48180.0 33395.0 48885.0 34740.0 ;
      RECT  48180.0 36085.0 48885.0 34740.0 ;
      RECT  48180.0 36085.0 48885.0 37430.0 ;
      RECT  48180.0 38775.0 48885.0 37430.0 ;
      RECT  48180.0 38775.0 48885.0 40120.0 ;
      RECT  48180.0 41465.0 48885.0 40120.0 ;
      RECT  48180.0 41465.0 48885.0 42810.0 ;
      RECT  48180.0 44155.0 48885.0 42810.0 ;
      RECT  48180.0 44155.0 48885.0 45500.0 ;
      RECT  48180.0 46845.0 48885.0 45500.0 ;
      RECT  48180.0 46845.0 48885.0 48190.0 ;
      RECT  48180.0 49535.0 48885.0 48190.0 ;
      RECT  48180.0 49535.0 48885.0 50880.0 ;
      RECT  48180.0 52225.0 48885.0 50880.0 ;
      RECT  48180.0 52225.0 48885.0 53570.0 ;
      RECT  48180.0 54915.0 48885.0 53570.0 ;
      RECT  48180.0 54915.0 48885.0 56260.0 ;
      RECT  48180.0 57605.0 48885.0 56260.0 ;
      RECT  48180.0 57605.0 48885.0 58950.0 ;
      RECT  48180.0 60295.0 48885.0 58950.0 ;
      RECT  48180.0 60295.0 48885.0 61640.0 ;
      RECT  48180.0 62985.0 48885.0 61640.0 ;
      RECT  48180.0 62985.0 48885.0 64330.0 ;
      RECT  48180.0 65675.0 48885.0 64330.0 ;
      RECT  48180.0 65675.0 48885.0 67020.0 ;
      RECT  48180.0 68365.0 48885.0 67020.0 ;
      RECT  48180.0 68365.0 48885.0 69710.0 ;
      RECT  48180.0 71055.0 48885.0 69710.0 ;
      RECT  48180.0 71055.0 48885.0 72400.0 ;
      RECT  48180.0 73745.0 48885.0 72400.0 ;
      RECT  48180.0 73745.0 48885.0 75090.0 ;
      RECT  48180.0 76435.0 48885.0 75090.0 ;
      RECT  48180.0 76435.0 48885.0 77780.0 ;
      RECT  48180.0 79125.0 48885.0 77780.0 ;
      RECT  48180.0 79125.0 48885.0 80470.0 ;
      RECT  48180.0 81815.0 48885.0 80470.0 ;
      RECT  48180.0 81815.0 48885.0 83160.0 ;
      RECT  48180.0 84505.0 48885.0 83160.0 ;
      RECT  48180.0 84505.0 48885.0 85850.0 ;
      RECT  48180.0 87195.0 48885.0 85850.0 ;
      RECT  48180.0 87195.0 48885.0 88540.0 ;
      RECT  48180.0 89885.0 48885.0 88540.0 ;
      RECT  48180.0 89885.0 48885.0 91230.0 ;
      RECT  48180.0 92575.0 48885.0 91230.0 ;
      RECT  48180.0 92575.0 48885.0 93920.0 ;
      RECT  48180.0 95265.0 48885.0 93920.0 ;
      RECT  48180.0 95265.0 48885.0 96610.0 ;
      RECT  48180.0 97955.0 48885.0 96610.0 ;
      RECT  48180.0 97955.0 48885.0 99300.0 ;
      RECT  48180.0 100645.0 48885.0 99300.0 ;
      RECT  48180.0 100645.0 48885.0 101990.0 ;
      RECT  48180.0 103335.0 48885.0 101990.0 ;
      RECT  48180.0 103335.0 48885.0 104680.0 ;
      RECT  48180.0 106025.0 48885.0 104680.0 ;
      RECT  48180.0 106025.0 48885.0 107370.0 ;
      RECT  48180.0 108715.0 48885.0 107370.0 ;
      RECT  48180.0 108715.0 48885.0 110060.0 ;
      RECT  48180.0 111405.0 48885.0 110060.0 ;
      RECT  48180.0 111405.0 48885.0 112750.0 ;
      RECT  48180.0 114095.0 48885.0 112750.0 ;
      RECT  48885.0 28015.0 49590.0 29360.0 ;
      RECT  48885.0 30705.0 49590.0 29360.0 ;
      RECT  48885.0 30705.0 49590.0 32050.0 ;
      RECT  48885.0 33395.0 49590.0 32050.0 ;
      RECT  48885.0 33395.0 49590.0 34740.0 ;
      RECT  48885.0 36085.0 49590.0 34740.0 ;
      RECT  48885.0 36085.0 49590.0 37430.0 ;
      RECT  48885.0 38775.0 49590.0 37430.0 ;
      RECT  48885.0 38775.0 49590.0 40120.0 ;
      RECT  48885.0 41465.0 49590.0 40120.0 ;
      RECT  48885.0 41465.0 49590.0 42810.0 ;
      RECT  48885.0 44155.0 49590.0 42810.0 ;
      RECT  48885.0 44155.0 49590.0 45500.0 ;
      RECT  48885.0 46845.0 49590.0 45500.0 ;
      RECT  48885.0 46845.0 49590.0 48190.0 ;
      RECT  48885.0 49535.0 49590.0 48190.0 ;
      RECT  48885.0 49535.0 49590.0 50880.0 ;
      RECT  48885.0 52225.0 49590.0 50880.0 ;
      RECT  48885.0 52225.0 49590.0 53570.0 ;
      RECT  48885.0 54915.0 49590.0 53570.0 ;
      RECT  48885.0 54915.0 49590.0 56260.0 ;
      RECT  48885.0 57605.0 49590.0 56260.0 ;
      RECT  48885.0 57605.0 49590.0 58950.0 ;
      RECT  48885.0 60295.0 49590.0 58950.0 ;
      RECT  48885.0 60295.0 49590.0 61640.0 ;
      RECT  48885.0 62985.0 49590.0 61640.0 ;
      RECT  48885.0 62985.0 49590.0 64330.0 ;
      RECT  48885.0 65675.0 49590.0 64330.0 ;
      RECT  48885.0 65675.0 49590.0 67020.0 ;
      RECT  48885.0 68365.0 49590.0 67020.0 ;
      RECT  48885.0 68365.0 49590.0 69710.0 ;
      RECT  48885.0 71055.0 49590.0 69710.0 ;
      RECT  48885.0 71055.0 49590.0 72400.0 ;
      RECT  48885.0 73745.0 49590.0 72400.0 ;
      RECT  48885.0 73745.0 49590.0 75090.0 ;
      RECT  48885.0 76435.0 49590.0 75090.0 ;
      RECT  48885.0 76435.0 49590.0 77780.0 ;
      RECT  48885.0 79125.0 49590.0 77780.0 ;
      RECT  48885.0 79125.0 49590.0 80470.0 ;
      RECT  48885.0 81815.0 49590.0 80470.0 ;
      RECT  48885.0 81815.0 49590.0 83160.0 ;
      RECT  48885.0 84505.0 49590.0 83160.0 ;
      RECT  48885.0 84505.0 49590.0 85850.0 ;
      RECT  48885.0 87195.0 49590.0 85850.0 ;
      RECT  48885.0 87195.0 49590.0 88540.0 ;
      RECT  48885.0 89885.0 49590.0 88540.0 ;
      RECT  48885.0 89885.0 49590.0 91230.0 ;
      RECT  48885.0 92575.0 49590.0 91230.0 ;
      RECT  48885.0 92575.0 49590.0 93920.0 ;
      RECT  48885.0 95265.0 49590.0 93920.0 ;
      RECT  48885.0 95265.0 49590.0 96610.0 ;
      RECT  48885.0 97955.0 49590.0 96610.0 ;
      RECT  48885.0 97955.0 49590.0 99300.0 ;
      RECT  48885.0 100645.0 49590.0 99300.0 ;
      RECT  48885.0 100645.0 49590.0 101990.0 ;
      RECT  48885.0 103335.0 49590.0 101990.0 ;
      RECT  48885.0 103335.0 49590.0 104680.0 ;
      RECT  48885.0 106025.0 49590.0 104680.0 ;
      RECT  48885.0 106025.0 49590.0 107370.0 ;
      RECT  48885.0 108715.0 49590.0 107370.0 ;
      RECT  48885.0 108715.0 49590.0 110060.0 ;
      RECT  48885.0 111405.0 49590.0 110060.0 ;
      RECT  48885.0 111405.0 49590.0 112750.0 ;
      RECT  48885.0 114095.0 49590.0 112750.0 ;
      RECT  49590.0 28015.0 50295.0 29360.0 ;
      RECT  49590.0 30705.0 50295.0 29360.0 ;
      RECT  49590.0 30705.0 50295.0 32050.0 ;
      RECT  49590.0 33395.0 50295.0 32050.0 ;
      RECT  49590.0 33395.0 50295.0 34740.0 ;
      RECT  49590.0 36085.0 50295.0 34740.0 ;
      RECT  49590.0 36085.0 50295.0 37430.0 ;
      RECT  49590.0 38775.0 50295.0 37430.0 ;
      RECT  49590.0 38775.0 50295.0 40120.0 ;
      RECT  49590.0 41465.0 50295.0 40120.0 ;
      RECT  49590.0 41465.0 50295.0 42810.0 ;
      RECT  49590.0 44155.0 50295.0 42810.0 ;
      RECT  49590.0 44155.0 50295.0 45500.0 ;
      RECT  49590.0 46845.0 50295.0 45500.0 ;
      RECT  49590.0 46845.0 50295.0 48190.0 ;
      RECT  49590.0 49535.0 50295.0 48190.0 ;
      RECT  49590.0 49535.0 50295.0 50880.0 ;
      RECT  49590.0 52225.0 50295.0 50880.0 ;
      RECT  49590.0 52225.0 50295.0 53570.0 ;
      RECT  49590.0 54915.0 50295.0 53570.0 ;
      RECT  49590.0 54915.0 50295.0 56260.0 ;
      RECT  49590.0 57605.0 50295.0 56260.0 ;
      RECT  49590.0 57605.0 50295.0 58950.0 ;
      RECT  49590.0 60295.0 50295.0 58950.0 ;
      RECT  49590.0 60295.0 50295.0 61640.0 ;
      RECT  49590.0 62985.0 50295.0 61640.0 ;
      RECT  49590.0 62985.0 50295.0 64330.0 ;
      RECT  49590.0 65675.0 50295.0 64330.0 ;
      RECT  49590.0 65675.0 50295.0 67020.0 ;
      RECT  49590.0 68365.0 50295.0 67020.0 ;
      RECT  49590.0 68365.0 50295.0 69710.0 ;
      RECT  49590.0 71055.0 50295.0 69710.0 ;
      RECT  49590.0 71055.0 50295.0 72400.0 ;
      RECT  49590.0 73745.0 50295.0 72400.0 ;
      RECT  49590.0 73745.0 50295.0 75090.0 ;
      RECT  49590.0 76435.0 50295.0 75090.0 ;
      RECT  49590.0 76435.0 50295.0 77780.0 ;
      RECT  49590.0 79125.0 50295.0 77780.0 ;
      RECT  49590.0 79125.0 50295.0 80470.0 ;
      RECT  49590.0 81815.0 50295.0 80470.0 ;
      RECT  49590.0 81815.0 50295.0 83160.0 ;
      RECT  49590.0 84505.0 50295.0 83160.0 ;
      RECT  49590.0 84505.0 50295.0 85850.0 ;
      RECT  49590.0 87195.0 50295.0 85850.0 ;
      RECT  49590.0 87195.0 50295.0 88540.0 ;
      RECT  49590.0 89885.0 50295.0 88540.0 ;
      RECT  49590.0 89885.0 50295.0 91230.0 ;
      RECT  49590.0 92575.0 50295.0 91230.0 ;
      RECT  49590.0 92575.0 50295.0 93920.0 ;
      RECT  49590.0 95265.0 50295.0 93920.0 ;
      RECT  49590.0 95265.0 50295.0 96610.0 ;
      RECT  49590.0 97955.0 50295.0 96610.0 ;
      RECT  49590.0 97955.0 50295.0 99300.0 ;
      RECT  49590.0 100645.0 50295.0 99300.0 ;
      RECT  49590.0 100645.0 50295.0 101990.0 ;
      RECT  49590.0 103335.0 50295.0 101990.0 ;
      RECT  49590.0 103335.0 50295.0 104680.0 ;
      RECT  49590.0 106025.0 50295.0 104680.0 ;
      RECT  49590.0 106025.0 50295.0 107370.0 ;
      RECT  49590.0 108715.0 50295.0 107370.0 ;
      RECT  49590.0 108715.0 50295.0 110060.0 ;
      RECT  49590.0 111405.0 50295.0 110060.0 ;
      RECT  49590.0 111405.0 50295.0 112750.0 ;
      RECT  49590.0 114095.0 50295.0 112750.0 ;
      RECT  50295.0 28015.0 51000.0 29360.0 ;
      RECT  50295.0 30705.0 51000.0 29360.0 ;
      RECT  50295.0 30705.0 51000.0 32050.0 ;
      RECT  50295.0 33395.0 51000.0 32050.0 ;
      RECT  50295.0 33395.0 51000.0 34740.0 ;
      RECT  50295.0 36085.0 51000.0 34740.0 ;
      RECT  50295.0 36085.0 51000.0 37430.0 ;
      RECT  50295.0 38775.0 51000.0 37430.0 ;
      RECT  50295.0 38775.0 51000.0 40120.0 ;
      RECT  50295.0 41465.0 51000.0 40120.0 ;
      RECT  50295.0 41465.0 51000.0 42810.0 ;
      RECT  50295.0 44155.0 51000.0 42810.0 ;
      RECT  50295.0 44155.0 51000.0 45500.0 ;
      RECT  50295.0 46845.0 51000.0 45500.0 ;
      RECT  50295.0 46845.0 51000.0 48190.0 ;
      RECT  50295.0 49535.0 51000.0 48190.0 ;
      RECT  50295.0 49535.0 51000.0 50880.0 ;
      RECT  50295.0 52225.0 51000.0 50880.0 ;
      RECT  50295.0 52225.0 51000.0 53570.0 ;
      RECT  50295.0 54915.0 51000.0 53570.0 ;
      RECT  50295.0 54915.0 51000.0 56260.0 ;
      RECT  50295.0 57605.0 51000.0 56260.0 ;
      RECT  50295.0 57605.0 51000.0 58950.0 ;
      RECT  50295.0 60295.0 51000.0 58950.0 ;
      RECT  50295.0 60295.0 51000.0 61640.0 ;
      RECT  50295.0 62985.0 51000.0 61640.0 ;
      RECT  50295.0 62985.0 51000.0 64330.0 ;
      RECT  50295.0 65675.0 51000.0 64330.0 ;
      RECT  50295.0 65675.0 51000.0 67020.0 ;
      RECT  50295.0 68365.0 51000.0 67020.0 ;
      RECT  50295.0 68365.0 51000.0 69710.0 ;
      RECT  50295.0 71055.0 51000.0 69710.0 ;
      RECT  50295.0 71055.0 51000.0 72400.0 ;
      RECT  50295.0 73745.0 51000.0 72400.0 ;
      RECT  50295.0 73745.0 51000.0 75090.0 ;
      RECT  50295.0 76435.0 51000.0 75090.0 ;
      RECT  50295.0 76435.0 51000.0 77780.0 ;
      RECT  50295.0 79125.0 51000.0 77780.0 ;
      RECT  50295.0 79125.0 51000.0 80470.0 ;
      RECT  50295.0 81815.0 51000.0 80470.0 ;
      RECT  50295.0 81815.0 51000.0 83160.0 ;
      RECT  50295.0 84505.0 51000.0 83160.0 ;
      RECT  50295.0 84505.0 51000.0 85850.0 ;
      RECT  50295.0 87195.0 51000.0 85850.0 ;
      RECT  50295.0 87195.0 51000.0 88540.0 ;
      RECT  50295.0 89885.0 51000.0 88540.0 ;
      RECT  50295.0 89885.0 51000.0 91230.0 ;
      RECT  50295.0 92575.0 51000.0 91230.0 ;
      RECT  50295.0 92575.0 51000.0 93920.0 ;
      RECT  50295.0 95265.0 51000.0 93920.0 ;
      RECT  50295.0 95265.0 51000.0 96610.0 ;
      RECT  50295.0 97955.0 51000.0 96610.0 ;
      RECT  50295.0 97955.0 51000.0 99300.0 ;
      RECT  50295.0 100645.0 51000.0 99300.0 ;
      RECT  50295.0 100645.0 51000.0 101990.0 ;
      RECT  50295.0 103335.0 51000.0 101990.0 ;
      RECT  50295.0 103335.0 51000.0 104680.0 ;
      RECT  50295.0 106025.0 51000.0 104680.0 ;
      RECT  50295.0 106025.0 51000.0 107370.0 ;
      RECT  50295.0 108715.0 51000.0 107370.0 ;
      RECT  50295.0 108715.0 51000.0 110060.0 ;
      RECT  50295.0 111405.0 51000.0 110060.0 ;
      RECT  50295.0 111405.0 51000.0 112750.0 ;
      RECT  50295.0 114095.0 51000.0 112750.0 ;
      RECT  51000.0 28015.0 51705.0 29360.0 ;
      RECT  51000.0 30705.0 51705.0 29360.0 ;
      RECT  51000.0 30705.0 51705.0 32050.0 ;
      RECT  51000.0 33395.0 51705.0 32050.0 ;
      RECT  51000.0 33395.0 51705.0 34740.0 ;
      RECT  51000.0 36085.0 51705.0 34740.0 ;
      RECT  51000.0 36085.0 51705.0 37430.0 ;
      RECT  51000.0 38775.0 51705.0 37430.0 ;
      RECT  51000.0 38775.0 51705.0 40120.0 ;
      RECT  51000.0 41465.0 51705.0 40120.0 ;
      RECT  51000.0 41465.0 51705.0 42810.0 ;
      RECT  51000.0 44155.0 51705.0 42810.0 ;
      RECT  51000.0 44155.0 51705.0 45500.0 ;
      RECT  51000.0 46845.0 51705.0 45500.0 ;
      RECT  51000.0 46845.0 51705.0 48190.0 ;
      RECT  51000.0 49535.0 51705.0 48190.0 ;
      RECT  51000.0 49535.0 51705.0 50880.0 ;
      RECT  51000.0 52225.0 51705.0 50880.0 ;
      RECT  51000.0 52225.0 51705.0 53570.0 ;
      RECT  51000.0 54915.0 51705.0 53570.0 ;
      RECT  51000.0 54915.0 51705.0 56260.0 ;
      RECT  51000.0 57605.0 51705.0 56260.0 ;
      RECT  51000.0 57605.0 51705.0 58950.0 ;
      RECT  51000.0 60295.0 51705.0 58950.0 ;
      RECT  51000.0 60295.0 51705.0 61640.0 ;
      RECT  51000.0 62985.0 51705.0 61640.0 ;
      RECT  51000.0 62985.0 51705.0 64330.0 ;
      RECT  51000.0 65675.0 51705.0 64330.0 ;
      RECT  51000.0 65675.0 51705.0 67020.0 ;
      RECT  51000.0 68365.0 51705.0 67020.0 ;
      RECT  51000.0 68365.0 51705.0 69710.0 ;
      RECT  51000.0 71055.0 51705.0 69710.0 ;
      RECT  51000.0 71055.0 51705.0 72400.0 ;
      RECT  51000.0 73745.0 51705.0 72400.0 ;
      RECT  51000.0 73745.0 51705.0 75090.0 ;
      RECT  51000.0 76435.0 51705.0 75090.0 ;
      RECT  51000.0 76435.0 51705.0 77780.0 ;
      RECT  51000.0 79125.0 51705.0 77780.0 ;
      RECT  51000.0 79125.0 51705.0 80470.0 ;
      RECT  51000.0 81815.0 51705.0 80470.0 ;
      RECT  51000.0 81815.0 51705.0 83160.0 ;
      RECT  51000.0 84505.0 51705.0 83160.0 ;
      RECT  51000.0 84505.0 51705.0 85850.0 ;
      RECT  51000.0 87195.0 51705.0 85850.0 ;
      RECT  51000.0 87195.0 51705.0 88540.0 ;
      RECT  51000.0 89885.0 51705.0 88540.0 ;
      RECT  51000.0 89885.0 51705.0 91230.0 ;
      RECT  51000.0 92575.0 51705.0 91230.0 ;
      RECT  51000.0 92575.0 51705.0 93920.0 ;
      RECT  51000.0 95265.0 51705.0 93920.0 ;
      RECT  51000.0 95265.0 51705.0 96610.0 ;
      RECT  51000.0 97955.0 51705.0 96610.0 ;
      RECT  51000.0 97955.0 51705.0 99300.0 ;
      RECT  51000.0 100645.0 51705.0 99300.0 ;
      RECT  51000.0 100645.0 51705.0 101990.0 ;
      RECT  51000.0 103335.0 51705.0 101990.0 ;
      RECT  51000.0 103335.0 51705.0 104680.0 ;
      RECT  51000.0 106025.0 51705.0 104680.0 ;
      RECT  51000.0 106025.0 51705.0 107370.0 ;
      RECT  51000.0 108715.0 51705.0 107370.0 ;
      RECT  51000.0 108715.0 51705.0 110060.0 ;
      RECT  51000.0 111405.0 51705.0 110060.0 ;
      RECT  51000.0 111405.0 51705.0 112750.0 ;
      RECT  51000.0 114095.0 51705.0 112750.0 ;
      RECT  51705.0 28015.0 52410.0 29360.0 ;
      RECT  51705.0 30705.0 52410.0 29360.0 ;
      RECT  51705.0 30705.0 52410.0 32050.0 ;
      RECT  51705.0 33395.0 52410.0 32050.0 ;
      RECT  51705.0 33395.0 52410.0 34740.0 ;
      RECT  51705.0 36085.0 52410.0 34740.0 ;
      RECT  51705.0 36085.0 52410.0 37430.0 ;
      RECT  51705.0 38775.0 52410.0 37430.0 ;
      RECT  51705.0 38775.0 52410.0 40120.0 ;
      RECT  51705.0 41465.0 52410.0 40120.0 ;
      RECT  51705.0 41465.0 52410.0 42810.0 ;
      RECT  51705.0 44155.0 52410.0 42810.0 ;
      RECT  51705.0 44155.0 52410.0 45500.0 ;
      RECT  51705.0 46845.0 52410.0 45500.0 ;
      RECT  51705.0 46845.0 52410.0 48190.0 ;
      RECT  51705.0 49535.0 52410.0 48190.0 ;
      RECT  51705.0 49535.0 52410.0 50880.0 ;
      RECT  51705.0 52225.0 52410.0 50880.0 ;
      RECT  51705.0 52225.0 52410.0 53570.0 ;
      RECT  51705.0 54915.0 52410.0 53570.0 ;
      RECT  51705.0 54915.0 52410.0 56260.0 ;
      RECT  51705.0 57605.0 52410.0 56260.0 ;
      RECT  51705.0 57605.0 52410.0 58950.0 ;
      RECT  51705.0 60295.0 52410.0 58950.0 ;
      RECT  51705.0 60295.0 52410.0 61640.0 ;
      RECT  51705.0 62985.0 52410.0 61640.0 ;
      RECT  51705.0 62985.0 52410.0 64330.0 ;
      RECT  51705.0 65675.0 52410.0 64330.0 ;
      RECT  51705.0 65675.0 52410.0 67020.0 ;
      RECT  51705.0 68365.0 52410.0 67020.0 ;
      RECT  51705.0 68365.0 52410.0 69710.0 ;
      RECT  51705.0 71055.0 52410.0 69710.0 ;
      RECT  51705.0 71055.0 52410.0 72400.0 ;
      RECT  51705.0 73745.0 52410.0 72400.0 ;
      RECT  51705.0 73745.0 52410.0 75090.0 ;
      RECT  51705.0 76435.0 52410.0 75090.0 ;
      RECT  51705.0 76435.0 52410.0 77780.0 ;
      RECT  51705.0 79125.0 52410.0 77780.0 ;
      RECT  51705.0 79125.0 52410.0 80470.0 ;
      RECT  51705.0 81815.0 52410.0 80470.0 ;
      RECT  51705.0 81815.0 52410.0 83160.0 ;
      RECT  51705.0 84505.0 52410.0 83160.0 ;
      RECT  51705.0 84505.0 52410.0 85850.0 ;
      RECT  51705.0 87195.0 52410.0 85850.0 ;
      RECT  51705.0 87195.0 52410.0 88540.0 ;
      RECT  51705.0 89885.0 52410.0 88540.0 ;
      RECT  51705.0 89885.0 52410.0 91230.0 ;
      RECT  51705.0 92575.0 52410.0 91230.0 ;
      RECT  51705.0 92575.0 52410.0 93920.0 ;
      RECT  51705.0 95265.0 52410.0 93920.0 ;
      RECT  51705.0 95265.0 52410.0 96610.0 ;
      RECT  51705.0 97955.0 52410.0 96610.0 ;
      RECT  51705.0 97955.0 52410.0 99300.0 ;
      RECT  51705.0 100645.0 52410.0 99300.0 ;
      RECT  51705.0 100645.0 52410.0 101990.0 ;
      RECT  51705.0 103335.0 52410.0 101990.0 ;
      RECT  51705.0 103335.0 52410.0 104680.0 ;
      RECT  51705.0 106025.0 52410.0 104680.0 ;
      RECT  51705.0 106025.0 52410.0 107370.0 ;
      RECT  51705.0 108715.0 52410.0 107370.0 ;
      RECT  51705.0 108715.0 52410.0 110060.0 ;
      RECT  51705.0 111405.0 52410.0 110060.0 ;
      RECT  51705.0 111405.0 52410.0 112750.0 ;
      RECT  51705.0 114095.0 52410.0 112750.0 ;
      RECT  52410.0 28015.0 53115.0 29360.0 ;
      RECT  52410.0 30705.0 53115.0 29360.0 ;
      RECT  52410.0 30705.0 53115.0 32050.0 ;
      RECT  52410.0 33395.0 53115.0 32050.0 ;
      RECT  52410.0 33395.0 53115.0 34740.0 ;
      RECT  52410.0 36085.0 53115.0 34740.0 ;
      RECT  52410.0 36085.0 53115.0 37430.0 ;
      RECT  52410.0 38775.0 53115.0 37430.0 ;
      RECT  52410.0 38775.0 53115.0 40120.0 ;
      RECT  52410.0 41465.0 53115.0 40120.0 ;
      RECT  52410.0 41465.0 53115.0 42810.0 ;
      RECT  52410.0 44155.0 53115.0 42810.0 ;
      RECT  52410.0 44155.0 53115.0 45500.0 ;
      RECT  52410.0 46845.0 53115.0 45500.0 ;
      RECT  52410.0 46845.0 53115.0 48190.0 ;
      RECT  52410.0 49535.0 53115.0 48190.0 ;
      RECT  52410.0 49535.0 53115.0 50880.0 ;
      RECT  52410.0 52225.0 53115.0 50880.0 ;
      RECT  52410.0 52225.0 53115.0 53570.0 ;
      RECT  52410.0 54915.0 53115.0 53570.0 ;
      RECT  52410.0 54915.0 53115.0 56260.0 ;
      RECT  52410.0 57605.0 53115.0 56260.0 ;
      RECT  52410.0 57605.0 53115.0 58950.0 ;
      RECT  52410.0 60295.0 53115.0 58950.0 ;
      RECT  52410.0 60295.0 53115.0 61640.0 ;
      RECT  52410.0 62985.0 53115.0 61640.0 ;
      RECT  52410.0 62985.0 53115.0 64330.0 ;
      RECT  52410.0 65675.0 53115.0 64330.0 ;
      RECT  52410.0 65675.0 53115.0 67020.0 ;
      RECT  52410.0 68365.0 53115.0 67020.0 ;
      RECT  52410.0 68365.0 53115.0 69710.0 ;
      RECT  52410.0 71055.0 53115.0 69710.0 ;
      RECT  52410.0 71055.0 53115.0 72400.0 ;
      RECT  52410.0 73745.0 53115.0 72400.0 ;
      RECT  52410.0 73745.0 53115.0 75090.0 ;
      RECT  52410.0 76435.0 53115.0 75090.0 ;
      RECT  52410.0 76435.0 53115.0 77780.0 ;
      RECT  52410.0 79125.0 53115.0 77780.0 ;
      RECT  52410.0 79125.0 53115.0 80470.0 ;
      RECT  52410.0 81815.0 53115.0 80470.0 ;
      RECT  52410.0 81815.0 53115.0 83160.0 ;
      RECT  52410.0 84505.0 53115.0 83160.0 ;
      RECT  52410.0 84505.0 53115.0 85850.0 ;
      RECT  52410.0 87195.0 53115.0 85850.0 ;
      RECT  52410.0 87195.0 53115.0 88540.0 ;
      RECT  52410.0 89885.0 53115.0 88540.0 ;
      RECT  52410.0 89885.0 53115.0 91230.0 ;
      RECT  52410.0 92575.0 53115.0 91230.0 ;
      RECT  52410.0 92575.0 53115.0 93920.0 ;
      RECT  52410.0 95265.0 53115.0 93920.0 ;
      RECT  52410.0 95265.0 53115.0 96610.0 ;
      RECT  52410.0 97955.0 53115.0 96610.0 ;
      RECT  52410.0 97955.0 53115.0 99300.0 ;
      RECT  52410.0 100645.0 53115.0 99300.0 ;
      RECT  52410.0 100645.0 53115.0 101990.0 ;
      RECT  52410.0 103335.0 53115.0 101990.0 ;
      RECT  52410.0 103335.0 53115.0 104680.0 ;
      RECT  52410.0 106025.0 53115.0 104680.0 ;
      RECT  52410.0 106025.0 53115.0 107370.0 ;
      RECT  52410.0 108715.0 53115.0 107370.0 ;
      RECT  52410.0 108715.0 53115.0 110060.0 ;
      RECT  52410.0 111405.0 53115.0 110060.0 ;
      RECT  52410.0 111405.0 53115.0 112750.0 ;
      RECT  52410.0 114095.0 53115.0 112750.0 ;
      RECT  53115.0 28015.0 53820.0 29360.0 ;
      RECT  53115.0 30705.0 53820.0 29360.0 ;
      RECT  53115.0 30705.0 53820.0 32050.0 ;
      RECT  53115.0 33395.0 53820.0 32050.0 ;
      RECT  53115.0 33395.0 53820.0 34740.0 ;
      RECT  53115.0 36085.0 53820.0 34740.0 ;
      RECT  53115.0 36085.0 53820.0 37430.0 ;
      RECT  53115.0 38775.0 53820.0 37430.0 ;
      RECT  53115.0 38775.0 53820.0 40120.0 ;
      RECT  53115.0 41465.0 53820.0 40120.0 ;
      RECT  53115.0 41465.0 53820.0 42810.0 ;
      RECT  53115.0 44155.0 53820.0 42810.0 ;
      RECT  53115.0 44155.0 53820.0 45500.0 ;
      RECT  53115.0 46845.0 53820.0 45500.0 ;
      RECT  53115.0 46845.0 53820.0 48190.0 ;
      RECT  53115.0 49535.0 53820.0 48190.0 ;
      RECT  53115.0 49535.0 53820.0 50880.0 ;
      RECT  53115.0 52225.0 53820.0 50880.0 ;
      RECT  53115.0 52225.0 53820.0 53570.0 ;
      RECT  53115.0 54915.0 53820.0 53570.0 ;
      RECT  53115.0 54915.0 53820.0 56260.0 ;
      RECT  53115.0 57605.0 53820.0 56260.0 ;
      RECT  53115.0 57605.0 53820.0 58950.0 ;
      RECT  53115.0 60295.0 53820.0 58950.0 ;
      RECT  53115.0 60295.0 53820.0 61640.0 ;
      RECT  53115.0 62985.0 53820.0 61640.0 ;
      RECT  53115.0 62985.0 53820.0 64330.0 ;
      RECT  53115.0 65675.0 53820.0 64330.0 ;
      RECT  53115.0 65675.0 53820.0 67020.0 ;
      RECT  53115.0 68365.0 53820.0 67020.0 ;
      RECT  53115.0 68365.0 53820.0 69710.0 ;
      RECT  53115.0 71055.0 53820.0 69710.0 ;
      RECT  53115.0 71055.0 53820.0 72400.0 ;
      RECT  53115.0 73745.0 53820.0 72400.0 ;
      RECT  53115.0 73745.0 53820.0 75090.0 ;
      RECT  53115.0 76435.0 53820.0 75090.0 ;
      RECT  53115.0 76435.0 53820.0 77780.0 ;
      RECT  53115.0 79125.0 53820.0 77780.0 ;
      RECT  53115.0 79125.0 53820.0 80470.0 ;
      RECT  53115.0 81815.0 53820.0 80470.0 ;
      RECT  53115.0 81815.0 53820.0 83160.0 ;
      RECT  53115.0 84505.0 53820.0 83160.0 ;
      RECT  53115.0 84505.0 53820.0 85850.0 ;
      RECT  53115.0 87195.0 53820.0 85850.0 ;
      RECT  53115.0 87195.0 53820.0 88540.0 ;
      RECT  53115.0 89885.0 53820.0 88540.0 ;
      RECT  53115.0 89885.0 53820.0 91230.0 ;
      RECT  53115.0 92575.0 53820.0 91230.0 ;
      RECT  53115.0 92575.0 53820.0 93920.0 ;
      RECT  53115.0 95265.0 53820.0 93920.0 ;
      RECT  53115.0 95265.0 53820.0 96610.0 ;
      RECT  53115.0 97955.0 53820.0 96610.0 ;
      RECT  53115.0 97955.0 53820.0 99300.0 ;
      RECT  53115.0 100645.0 53820.0 99300.0 ;
      RECT  53115.0 100645.0 53820.0 101990.0 ;
      RECT  53115.0 103335.0 53820.0 101990.0 ;
      RECT  53115.0 103335.0 53820.0 104680.0 ;
      RECT  53115.0 106025.0 53820.0 104680.0 ;
      RECT  53115.0 106025.0 53820.0 107370.0 ;
      RECT  53115.0 108715.0 53820.0 107370.0 ;
      RECT  53115.0 108715.0 53820.0 110060.0 ;
      RECT  53115.0 111405.0 53820.0 110060.0 ;
      RECT  53115.0 111405.0 53820.0 112750.0 ;
      RECT  53115.0 114095.0 53820.0 112750.0 ;
      RECT  53820.0 28015.0 54525.0 29360.0 ;
      RECT  53820.0 30705.0 54525.0 29360.0 ;
      RECT  53820.0 30705.0 54525.0 32050.0 ;
      RECT  53820.0 33395.0 54525.0 32050.0 ;
      RECT  53820.0 33395.0 54525.0 34740.0 ;
      RECT  53820.0 36085.0 54525.0 34740.0 ;
      RECT  53820.0 36085.0 54525.0 37430.0 ;
      RECT  53820.0 38775.0 54525.0 37430.0 ;
      RECT  53820.0 38775.0 54525.0 40120.0 ;
      RECT  53820.0 41465.0 54525.0 40120.0 ;
      RECT  53820.0 41465.0 54525.0 42810.0 ;
      RECT  53820.0 44155.0 54525.0 42810.0 ;
      RECT  53820.0 44155.0 54525.0 45500.0 ;
      RECT  53820.0 46845.0 54525.0 45500.0 ;
      RECT  53820.0 46845.0 54525.0 48190.0 ;
      RECT  53820.0 49535.0 54525.0 48190.0 ;
      RECT  53820.0 49535.0 54525.0 50880.0 ;
      RECT  53820.0 52225.0 54525.0 50880.0 ;
      RECT  53820.0 52225.0 54525.0 53570.0 ;
      RECT  53820.0 54915.0 54525.0 53570.0 ;
      RECT  53820.0 54915.0 54525.0 56260.0 ;
      RECT  53820.0 57605.0 54525.0 56260.0 ;
      RECT  53820.0 57605.0 54525.0 58950.0 ;
      RECT  53820.0 60295.0 54525.0 58950.0 ;
      RECT  53820.0 60295.0 54525.0 61640.0 ;
      RECT  53820.0 62985.0 54525.0 61640.0 ;
      RECT  53820.0 62985.0 54525.0 64330.0 ;
      RECT  53820.0 65675.0 54525.0 64330.0 ;
      RECT  53820.0 65675.0 54525.0 67020.0 ;
      RECT  53820.0 68365.0 54525.0 67020.0 ;
      RECT  53820.0 68365.0 54525.0 69710.0 ;
      RECT  53820.0 71055.0 54525.0 69710.0 ;
      RECT  53820.0 71055.0 54525.0 72400.0 ;
      RECT  53820.0 73745.0 54525.0 72400.0 ;
      RECT  53820.0 73745.0 54525.0 75090.0 ;
      RECT  53820.0 76435.0 54525.0 75090.0 ;
      RECT  53820.0 76435.0 54525.0 77780.0 ;
      RECT  53820.0 79125.0 54525.0 77780.0 ;
      RECT  53820.0 79125.0 54525.0 80470.0 ;
      RECT  53820.0 81815.0 54525.0 80470.0 ;
      RECT  53820.0 81815.0 54525.0 83160.0 ;
      RECT  53820.0 84505.0 54525.0 83160.0 ;
      RECT  53820.0 84505.0 54525.0 85850.0 ;
      RECT  53820.0 87195.0 54525.0 85850.0 ;
      RECT  53820.0 87195.0 54525.0 88540.0 ;
      RECT  53820.0 89885.0 54525.0 88540.0 ;
      RECT  53820.0 89885.0 54525.0 91230.0 ;
      RECT  53820.0 92575.0 54525.0 91230.0 ;
      RECT  53820.0 92575.0 54525.0 93920.0 ;
      RECT  53820.0 95265.0 54525.0 93920.0 ;
      RECT  53820.0 95265.0 54525.0 96610.0 ;
      RECT  53820.0 97955.0 54525.0 96610.0 ;
      RECT  53820.0 97955.0 54525.0 99300.0 ;
      RECT  53820.0 100645.0 54525.0 99300.0 ;
      RECT  53820.0 100645.0 54525.0 101990.0 ;
      RECT  53820.0 103335.0 54525.0 101990.0 ;
      RECT  53820.0 103335.0 54525.0 104680.0 ;
      RECT  53820.0 106025.0 54525.0 104680.0 ;
      RECT  53820.0 106025.0 54525.0 107370.0 ;
      RECT  53820.0 108715.0 54525.0 107370.0 ;
      RECT  53820.0 108715.0 54525.0 110060.0 ;
      RECT  53820.0 111405.0 54525.0 110060.0 ;
      RECT  53820.0 111405.0 54525.0 112750.0 ;
      RECT  53820.0 114095.0 54525.0 112750.0 ;
      RECT  54525.0 28015.0 55230.0 29360.0 ;
      RECT  54525.0 30705.0 55230.0 29360.0 ;
      RECT  54525.0 30705.0 55230.0 32050.0 ;
      RECT  54525.0 33395.0 55230.0 32050.0 ;
      RECT  54525.0 33395.0 55230.0 34740.0 ;
      RECT  54525.0 36085.0 55230.0 34740.0 ;
      RECT  54525.0 36085.0 55230.0 37430.0 ;
      RECT  54525.0 38775.0 55230.0 37430.0 ;
      RECT  54525.0 38775.0 55230.0 40120.0 ;
      RECT  54525.0 41465.0 55230.0 40120.0 ;
      RECT  54525.0 41465.0 55230.0 42810.0 ;
      RECT  54525.0 44155.0 55230.0 42810.0 ;
      RECT  54525.0 44155.0 55230.0 45500.0 ;
      RECT  54525.0 46845.0 55230.0 45500.0 ;
      RECT  54525.0 46845.0 55230.0 48190.0 ;
      RECT  54525.0 49535.0 55230.0 48190.0 ;
      RECT  54525.0 49535.0 55230.0 50880.0 ;
      RECT  54525.0 52225.0 55230.0 50880.0 ;
      RECT  54525.0 52225.0 55230.0 53570.0 ;
      RECT  54525.0 54915.0 55230.0 53570.0 ;
      RECT  54525.0 54915.0 55230.0 56260.0 ;
      RECT  54525.0 57605.0 55230.0 56260.0 ;
      RECT  54525.0 57605.0 55230.0 58950.0 ;
      RECT  54525.0 60295.0 55230.0 58950.0 ;
      RECT  54525.0 60295.0 55230.0 61640.0 ;
      RECT  54525.0 62985.0 55230.0 61640.0 ;
      RECT  54525.0 62985.0 55230.0 64330.0 ;
      RECT  54525.0 65675.0 55230.0 64330.0 ;
      RECT  54525.0 65675.0 55230.0 67020.0 ;
      RECT  54525.0 68365.0 55230.0 67020.0 ;
      RECT  54525.0 68365.0 55230.0 69710.0 ;
      RECT  54525.0 71055.0 55230.0 69710.0 ;
      RECT  54525.0 71055.0 55230.0 72400.0 ;
      RECT  54525.0 73745.0 55230.0 72400.0 ;
      RECT  54525.0 73745.0 55230.0 75090.0 ;
      RECT  54525.0 76435.0 55230.0 75090.0 ;
      RECT  54525.0 76435.0 55230.0 77780.0 ;
      RECT  54525.0 79125.0 55230.0 77780.0 ;
      RECT  54525.0 79125.0 55230.0 80470.0 ;
      RECT  54525.0 81815.0 55230.0 80470.0 ;
      RECT  54525.0 81815.0 55230.0 83160.0 ;
      RECT  54525.0 84505.0 55230.0 83160.0 ;
      RECT  54525.0 84505.0 55230.0 85850.0 ;
      RECT  54525.0 87195.0 55230.0 85850.0 ;
      RECT  54525.0 87195.0 55230.0 88540.0 ;
      RECT  54525.0 89885.0 55230.0 88540.0 ;
      RECT  54525.0 89885.0 55230.0 91230.0 ;
      RECT  54525.0 92575.0 55230.0 91230.0 ;
      RECT  54525.0 92575.0 55230.0 93920.0 ;
      RECT  54525.0 95265.0 55230.0 93920.0 ;
      RECT  54525.0 95265.0 55230.0 96610.0 ;
      RECT  54525.0 97955.0 55230.0 96610.0 ;
      RECT  54525.0 97955.0 55230.0 99300.0 ;
      RECT  54525.0 100645.0 55230.0 99300.0 ;
      RECT  54525.0 100645.0 55230.0 101990.0 ;
      RECT  54525.0 103335.0 55230.0 101990.0 ;
      RECT  54525.0 103335.0 55230.0 104680.0 ;
      RECT  54525.0 106025.0 55230.0 104680.0 ;
      RECT  54525.0 106025.0 55230.0 107370.0 ;
      RECT  54525.0 108715.0 55230.0 107370.0 ;
      RECT  54525.0 108715.0 55230.0 110060.0 ;
      RECT  54525.0 111405.0 55230.0 110060.0 ;
      RECT  54525.0 111405.0 55230.0 112750.0 ;
      RECT  54525.0 114095.0 55230.0 112750.0 ;
      RECT  55230.0 28015.0 55935.0 29360.0 ;
      RECT  55230.0 30705.0 55935.0 29360.0 ;
      RECT  55230.0 30705.0 55935.0 32050.0 ;
      RECT  55230.0 33395.0 55935.0 32050.0 ;
      RECT  55230.0 33395.0 55935.0 34740.0 ;
      RECT  55230.0 36085.0 55935.0 34740.0 ;
      RECT  55230.0 36085.0 55935.0 37430.0 ;
      RECT  55230.0 38775.0 55935.0 37430.0 ;
      RECT  55230.0 38775.0 55935.0 40120.0 ;
      RECT  55230.0 41465.0 55935.0 40120.0 ;
      RECT  55230.0 41465.0 55935.0 42810.0 ;
      RECT  55230.0 44155.0 55935.0 42810.0 ;
      RECT  55230.0 44155.0 55935.0 45500.0 ;
      RECT  55230.0 46845.0 55935.0 45500.0 ;
      RECT  55230.0 46845.0 55935.0 48190.0 ;
      RECT  55230.0 49535.0 55935.0 48190.0 ;
      RECT  55230.0 49535.0 55935.0 50880.0 ;
      RECT  55230.0 52225.0 55935.0 50880.0 ;
      RECT  55230.0 52225.0 55935.0 53570.0 ;
      RECT  55230.0 54915.0 55935.0 53570.0 ;
      RECT  55230.0 54915.0 55935.0 56260.0 ;
      RECT  55230.0 57605.0 55935.0 56260.0 ;
      RECT  55230.0 57605.0 55935.0 58950.0 ;
      RECT  55230.0 60295.0 55935.0 58950.0 ;
      RECT  55230.0 60295.0 55935.0 61640.0 ;
      RECT  55230.0 62985.0 55935.0 61640.0 ;
      RECT  55230.0 62985.0 55935.0 64330.0 ;
      RECT  55230.0 65675.0 55935.0 64330.0 ;
      RECT  55230.0 65675.0 55935.0 67020.0 ;
      RECT  55230.0 68365.0 55935.0 67020.0 ;
      RECT  55230.0 68365.0 55935.0 69710.0 ;
      RECT  55230.0 71055.0 55935.0 69710.0 ;
      RECT  55230.0 71055.0 55935.0 72400.0 ;
      RECT  55230.0 73745.0 55935.0 72400.0 ;
      RECT  55230.0 73745.0 55935.0 75090.0 ;
      RECT  55230.0 76435.0 55935.0 75090.0 ;
      RECT  55230.0 76435.0 55935.0 77780.0 ;
      RECT  55230.0 79125.0 55935.0 77780.0 ;
      RECT  55230.0 79125.0 55935.0 80470.0 ;
      RECT  55230.0 81815.0 55935.0 80470.0 ;
      RECT  55230.0 81815.0 55935.0 83160.0 ;
      RECT  55230.0 84505.0 55935.0 83160.0 ;
      RECT  55230.0 84505.0 55935.0 85850.0 ;
      RECT  55230.0 87195.0 55935.0 85850.0 ;
      RECT  55230.0 87195.0 55935.0 88540.0 ;
      RECT  55230.0 89885.0 55935.0 88540.0 ;
      RECT  55230.0 89885.0 55935.0 91230.0 ;
      RECT  55230.0 92575.0 55935.0 91230.0 ;
      RECT  55230.0 92575.0 55935.0 93920.0 ;
      RECT  55230.0 95265.0 55935.0 93920.0 ;
      RECT  55230.0 95265.0 55935.0 96610.0 ;
      RECT  55230.0 97955.0 55935.0 96610.0 ;
      RECT  55230.0 97955.0 55935.0 99300.0 ;
      RECT  55230.0 100645.0 55935.0 99300.0 ;
      RECT  55230.0 100645.0 55935.0 101990.0 ;
      RECT  55230.0 103335.0 55935.0 101990.0 ;
      RECT  55230.0 103335.0 55935.0 104680.0 ;
      RECT  55230.0 106025.0 55935.0 104680.0 ;
      RECT  55230.0 106025.0 55935.0 107370.0 ;
      RECT  55230.0 108715.0 55935.0 107370.0 ;
      RECT  55230.0 108715.0 55935.0 110060.0 ;
      RECT  55230.0 111405.0 55935.0 110060.0 ;
      RECT  55230.0 111405.0 55935.0 112750.0 ;
      RECT  55230.0 114095.0 55935.0 112750.0 ;
      RECT  55935.0 28015.0 56640.0 29360.0 ;
      RECT  55935.0 30705.0 56640.0 29360.0 ;
      RECT  55935.0 30705.0 56640.0 32050.0 ;
      RECT  55935.0 33395.0 56640.0 32050.0 ;
      RECT  55935.0 33395.0 56640.0 34740.0 ;
      RECT  55935.0 36085.0 56640.0 34740.0 ;
      RECT  55935.0 36085.0 56640.0 37430.0 ;
      RECT  55935.0 38775.0 56640.0 37430.0 ;
      RECT  55935.0 38775.0 56640.0 40120.0 ;
      RECT  55935.0 41465.0 56640.0 40120.0 ;
      RECT  55935.0 41465.0 56640.0 42810.0 ;
      RECT  55935.0 44155.0 56640.0 42810.0 ;
      RECT  55935.0 44155.0 56640.0 45500.0 ;
      RECT  55935.0 46845.0 56640.0 45500.0 ;
      RECT  55935.0 46845.0 56640.0 48190.0 ;
      RECT  55935.0 49535.0 56640.0 48190.0 ;
      RECT  55935.0 49535.0 56640.0 50880.0 ;
      RECT  55935.0 52225.0 56640.0 50880.0 ;
      RECT  55935.0 52225.0 56640.0 53570.0 ;
      RECT  55935.0 54915.0 56640.0 53570.0 ;
      RECT  55935.0 54915.0 56640.0 56260.0 ;
      RECT  55935.0 57605.0 56640.0 56260.0 ;
      RECT  55935.0 57605.0 56640.0 58950.0 ;
      RECT  55935.0 60295.0 56640.0 58950.0 ;
      RECT  55935.0 60295.0 56640.0 61640.0 ;
      RECT  55935.0 62985.0 56640.0 61640.0 ;
      RECT  55935.0 62985.0 56640.0 64330.0 ;
      RECT  55935.0 65675.0 56640.0 64330.0 ;
      RECT  55935.0 65675.0 56640.0 67020.0 ;
      RECT  55935.0 68365.0 56640.0 67020.0 ;
      RECT  55935.0 68365.0 56640.0 69710.0 ;
      RECT  55935.0 71055.0 56640.0 69710.0 ;
      RECT  55935.0 71055.0 56640.0 72400.0 ;
      RECT  55935.0 73745.0 56640.0 72400.0 ;
      RECT  55935.0 73745.0 56640.0 75090.0 ;
      RECT  55935.0 76435.0 56640.0 75090.0 ;
      RECT  55935.0 76435.0 56640.0 77780.0 ;
      RECT  55935.0 79125.0 56640.0 77780.0 ;
      RECT  55935.0 79125.0 56640.0 80470.0 ;
      RECT  55935.0 81815.0 56640.0 80470.0 ;
      RECT  55935.0 81815.0 56640.0 83160.0 ;
      RECT  55935.0 84505.0 56640.0 83160.0 ;
      RECT  55935.0 84505.0 56640.0 85850.0 ;
      RECT  55935.0 87195.0 56640.0 85850.0 ;
      RECT  55935.0 87195.0 56640.0 88540.0 ;
      RECT  55935.0 89885.0 56640.0 88540.0 ;
      RECT  55935.0 89885.0 56640.0 91230.0 ;
      RECT  55935.0 92575.0 56640.0 91230.0 ;
      RECT  55935.0 92575.0 56640.0 93920.0 ;
      RECT  55935.0 95265.0 56640.0 93920.0 ;
      RECT  55935.0 95265.0 56640.0 96610.0 ;
      RECT  55935.0 97955.0 56640.0 96610.0 ;
      RECT  55935.0 97955.0 56640.0 99300.0 ;
      RECT  55935.0 100645.0 56640.0 99300.0 ;
      RECT  55935.0 100645.0 56640.0 101990.0 ;
      RECT  55935.0 103335.0 56640.0 101990.0 ;
      RECT  55935.0 103335.0 56640.0 104680.0 ;
      RECT  55935.0 106025.0 56640.0 104680.0 ;
      RECT  55935.0 106025.0 56640.0 107370.0 ;
      RECT  55935.0 108715.0 56640.0 107370.0 ;
      RECT  55935.0 108715.0 56640.0 110060.0 ;
      RECT  55935.0 111405.0 56640.0 110060.0 ;
      RECT  55935.0 111405.0 56640.0 112750.0 ;
      RECT  55935.0 114095.0 56640.0 112750.0 ;
      RECT  56640.0 28015.0 57345.0 29360.0 ;
      RECT  56640.0 30705.0 57345.0 29360.0 ;
      RECT  56640.0 30705.0 57345.0 32050.0 ;
      RECT  56640.0 33395.0 57345.0 32050.0 ;
      RECT  56640.0 33395.0 57345.0 34740.0 ;
      RECT  56640.0 36085.0 57345.0 34740.0 ;
      RECT  56640.0 36085.0 57345.0 37430.0 ;
      RECT  56640.0 38775.0 57345.0 37430.0 ;
      RECT  56640.0 38775.0 57345.0 40120.0 ;
      RECT  56640.0 41465.0 57345.0 40120.0 ;
      RECT  56640.0 41465.0 57345.0 42810.0 ;
      RECT  56640.0 44155.0 57345.0 42810.0 ;
      RECT  56640.0 44155.0 57345.0 45500.0 ;
      RECT  56640.0 46845.0 57345.0 45500.0 ;
      RECT  56640.0 46845.0 57345.0 48190.0 ;
      RECT  56640.0 49535.0 57345.0 48190.0 ;
      RECT  56640.0 49535.0 57345.0 50880.0 ;
      RECT  56640.0 52225.0 57345.0 50880.0 ;
      RECT  56640.0 52225.0 57345.0 53570.0 ;
      RECT  56640.0 54915.0 57345.0 53570.0 ;
      RECT  56640.0 54915.0 57345.0 56260.0 ;
      RECT  56640.0 57605.0 57345.0 56260.0 ;
      RECT  56640.0 57605.0 57345.0 58950.0 ;
      RECT  56640.0 60295.0 57345.0 58950.0 ;
      RECT  56640.0 60295.0 57345.0 61640.0 ;
      RECT  56640.0 62985.0 57345.0 61640.0 ;
      RECT  56640.0 62985.0 57345.0 64330.0 ;
      RECT  56640.0 65675.0 57345.0 64330.0 ;
      RECT  56640.0 65675.0 57345.0 67020.0 ;
      RECT  56640.0 68365.0 57345.0 67020.0 ;
      RECT  56640.0 68365.0 57345.0 69710.0 ;
      RECT  56640.0 71055.0 57345.0 69710.0 ;
      RECT  56640.0 71055.0 57345.0 72400.0 ;
      RECT  56640.0 73745.0 57345.0 72400.0 ;
      RECT  56640.0 73745.0 57345.0 75090.0 ;
      RECT  56640.0 76435.0 57345.0 75090.0 ;
      RECT  56640.0 76435.0 57345.0 77780.0 ;
      RECT  56640.0 79125.0 57345.0 77780.0 ;
      RECT  56640.0 79125.0 57345.0 80470.0 ;
      RECT  56640.0 81815.0 57345.0 80470.0 ;
      RECT  56640.0 81815.0 57345.0 83160.0 ;
      RECT  56640.0 84505.0 57345.0 83160.0 ;
      RECT  56640.0 84505.0 57345.0 85850.0 ;
      RECT  56640.0 87195.0 57345.0 85850.0 ;
      RECT  56640.0 87195.0 57345.0 88540.0 ;
      RECT  56640.0 89885.0 57345.0 88540.0 ;
      RECT  56640.0 89885.0 57345.0 91230.0 ;
      RECT  56640.0 92575.0 57345.0 91230.0 ;
      RECT  56640.0 92575.0 57345.0 93920.0 ;
      RECT  56640.0 95265.0 57345.0 93920.0 ;
      RECT  56640.0 95265.0 57345.0 96610.0 ;
      RECT  56640.0 97955.0 57345.0 96610.0 ;
      RECT  56640.0 97955.0 57345.0 99300.0 ;
      RECT  56640.0 100645.0 57345.0 99300.0 ;
      RECT  56640.0 100645.0 57345.0 101990.0 ;
      RECT  56640.0 103335.0 57345.0 101990.0 ;
      RECT  56640.0 103335.0 57345.0 104680.0 ;
      RECT  56640.0 106025.0 57345.0 104680.0 ;
      RECT  56640.0 106025.0 57345.0 107370.0 ;
      RECT  56640.0 108715.0 57345.0 107370.0 ;
      RECT  56640.0 108715.0 57345.0 110060.0 ;
      RECT  56640.0 111405.0 57345.0 110060.0 ;
      RECT  56640.0 111405.0 57345.0 112750.0 ;
      RECT  56640.0 114095.0 57345.0 112750.0 ;
      RECT  57345.0 28015.0 58050.0 29360.0 ;
      RECT  57345.0 30705.0 58050.0 29360.0 ;
      RECT  57345.0 30705.0 58050.0 32050.0 ;
      RECT  57345.0 33395.0 58050.0 32050.0 ;
      RECT  57345.0 33395.0 58050.0 34740.0 ;
      RECT  57345.0 36085.0 58050.0 34740.0 ;
      RECT  57345.0 36085.0 58050.0 37430.0 ;
      RECT  57345.0 38775.0 58050.0 37430.0 ;
      RECT  57345.0 38775.0 58050.0 40120.0 ;
      RECT  57345.0 41465.0 58050.0 40120.0 ;
      RECT  57345.0 41465.0 58050.0 42810.0 ;
      RECT  57345.0 44155.0 58050.0 42810.0 ;
      RECT  57345.0 44155.0 58050.0 45500.0 ;
      RECT  57345.0 46845.0 58050.0 45500.0 ;
      RECT  57345.0 46845.0 58050.0 48190.0 ;
      RECT  57345.0 49535.0 58050.0 48190.0 ;
      RECT  57345.0 49535.0 58050.0 50880.0 ;
      RECT  57345.0 52225.0 58050.0 50880.0 ;
      RECT  57345.0 52225.0 58050.0 53570.0 ;
      RECT  57345.0 54915.0 58050.0 53570.0 ;
      RECT  57345.0 54915.0 58050.0 56260.0 ;
      RECT  57345.0 57605.0 58050.0 56260.0 ;
      RECT  57345.0 57605.0 58050.0 58950.0 ;
      RECT  57345.0 60295.0 58050.0 58950.0 ;
      RECT  57345.0 60295.0 58050.0 61640.0 ;
      RECT  57345.0 62985.0 58050.0 61640.0 ;
      RECT  57345.0 62985.0 58050.0 64330.0 ;
      RECT  57345.0 65675.0 58050.0 64330.0 ;
      RECT  57345.0 65675.0 58050.0 67020.0 ;
      RECT  57345.0 68365.0 58050.0 67020.0 ;
      RECT  57345.0 68365.0 58050.0 69710.0 ;
      RECT  57345.0 71055.0 58050.0 69710.0 ;
      RECT  57345.0 71055.0 58050.0 72400.0 ;
      RECT  57345.0 73745.0 58050.0 72400.0 ;
      RECT  57345.0 73745.0 58050.0 75090.0 ;
      RECT  57345.0 76435.0 58050.0 75090.0 ;
      RECT  57345.0 76435.0 58050.0 77780.0 ;
      RECT  57345.0 79125.0 58050.0 77780.0 ;
      RECT  57345.0 79125.0 58050.0 80470.0 ;
      RECT  57345.0 81815.0 58050.0 80470.0 ;
      RECT  57345.0 81815.0 58050.0 83160.0 ;
      RECT  57345.0 84505.0 58050.0 83160.0 ;
      RECT  57345.0 84505.0 58050.0 85850.0 ;
      RECT  57345.0 87195.0 58050.0 85850.0 ;
      RECT  57345.0 87195.0 58050.0 88540.0 ;
      RECT  57345.0 89885.0 58050.0 88540.0 ;
      RECT  57345.0 89885.0 58050.0 91230.0 ;
      RECT  57345.0 92575.0 58050.0 91230.0 ;
      RECT  57345.0 92575.0 58050.0 93920.0 ;
      RECT  57345.0 95265.0 58050.0 93920.0 ;
      RECT  57345.0 95265.0 58050.0 96610.0 ;
      RECT  57345.0 97955.0 58050.0 96610.0 ;
      RECT  57345.0 97955.0 58050.0 99300.0 ;
      RECT  57345.0 100645.0 58050.0 99300.0 ;
      RECT  57345.0 100645.0 58050.0 101990.0 ;
      RECT  57345.0 103335.0 58050.0 101990.0 ;
      RECT  57345.0 103335.0 58050.0 104680.0 ;
      RECT  57345.0 106025.0 58050.0 104680.0 ;
      RECT  57345.0 106025.0 58050.0 107370.0 ;
      RECT  57345.0 108715.0 58050.0 107370.0 ;
      RECT  57345.0 108715.0 58050.0 110060.0 ;
      RECT  57345.0 111405.0 58050.0 110060.0 ;
      RECT  57345.0 111405.0 58050.0 112750.0 ;
      RECT  57345.0 114095.0 58050.0 112750.0 ;
      RECT  58050.0 28015.0 58755.0 29360.0 ;
      RECT  58050.0 30705.0 58755.0 29360.0 ;
      RECT  58050.0 30705.0 58755.0 32050.0 ;
      RECT  58050.0 33395.0 58755.0 32050.0 ;
      RECT  58050.0 33395.0 58755.0 34740.0 ;
      RECT  58050.0 36085.0 58755.0 34740.0 ;
      RECT  58050.0 36085.0 58755.0 37430.0 ;
      RECT  58050.0 38775.0 58755.0 37430.0 ;
      RECT  58050.0 38775.0 58755.0 40120.0 ;
      RECT  58050.0 41465.0 58755.0 40120.0 ;
      RECT  58050.0 41465.0 58755.0 42810.0 ;
      RECT  58050.0 44155.0 58755.0 42810.0 ;
      RECT  58050.0 44155.0 58755.0 45500.0 ;
      RECT  58050.0 46845.0 58755.0 45500.0 ;
      RECT  58050.0 46845.0 58755.0 48190.0 ;
      RECT  58050.0 49535.0 58755.0 48190.0 ;
      RECT  58050.0 49535.0 58755.0 50880.0 ;
      RECT  58050.0 52225.0 58755.0 50880.0 ;
      RECT  58050.0 52225.0 58755.0 53570.0 ;
      RECT  58050.0 54915.0 58755.0 53570.0 ;
      RECT  58050.0 54915.0 58755.0 56260.0 ;
      RECT  58050.0 57605.0 58755.0 56260.0 ;
      RECT  58050.0 57605.0 58755.0 58950.0 ;
      RECT  58050.0 60295.0 58755.0 58950.0 ;
      RECT  58050.0 60295.0 58755.0 61640.0 ;
      RECT  58050.0 62985.0 58755.0 61640.0 ;
      RECT  58050.0 62985.0 58755.0 64330.0 ;
      RECT  58050.0 65675.0 58755.0 64330.0 ;
      RECT  58050.0 65675.0 58755.0 67020.0 ;
      RECT  58050.0 68365.0 58755.0 67020.0 ;
      RECT  58050.0 68365.0 58755.0 69710.0 ;
      RECT  58050.0 71055.0 58755.0 69710.0 ;
      RECT  58050.0 71055.0 58755.0 72400.0 ;
      RECT  58050.0 73745.0 58755.0 72400.0 ;
      RECT  58050.0 73745.0 58755.0 75090.0 ;
      RECT  58050.0 76435.0 58755.0 75090.0 ;
      RECT  58050.0 76435.0 58755.0 77780.0 ;
      RECT  58050.0 79125.0 58755.0 77780.0 ;
      RECT  58050.0 79125.0 58755.0 80470.0 ;
      RECT  58050.0 81815.0 58755.0 80470.0 ;
      RECT  58050.0 81815.0 58755.0 83160.0 ;
      RECT  58050.0 84505.0 58755.0 83160.0 ;
      RECT  58050.0 84505.0 58755.0 85850.0 ;
      RECT  58050.0 87195.0 58755.0 85850.0 ;
      RECT  58050.0 87195.0 58755.0 88540.0 ;
      RECT  58050.0 89885.0 58755.0 88540.0 ;
      RECT  58050.0 89885.0 58755.0 91230.0 ;
      RECT  58050.0 92575.0 58755.0 91230.0 ;
      RECT  58050.0 92575.0 58755.0 93920.0 ;
      RECT  58050.0 95265.0 58755.0 93920.0 ;
      RECT  58050.0 95265.0 58755.0 96610.0 ;
      RECT  58050.0 97955.0 58755.0 96610.0 ;
      RECT  58050.0 97955.0 58755.0 99300.0 ;
      RECT  58050.0 100645.0 58755.0 99300.0 ;
      RECT  58050.0 100645.0 58755.0 101990.0 ;
      RECT  58050.0 103335.0 58755.0 101990.0 ;
      RECT  58050.0 103335.0 58755.0 104680.0 ;
      RECT  58050.0 106025.0 58755.0 104680.0 ;
      RECT  58050.0 106025.0 58755.0 107370.0 ;
      RECT  58050.0 108715.0 58755.0 107370.0 ;
      RECT  58050.0 108715.0 58755.0 110060.0 ;
      RECT  58050.0 111405.0 58755.0 110060.0 ;
      RECT  58050.0 111405.0 58755.0 112750.0 ;
      RECT  58050.0 114095.0 58755.0 112750.0 ;
      RECT  58755.0 28015.0 59460.0 29360.0 ;
      RECT  58755.0 30705.0 59460.0 29360.0 ;
      RECT  58755.0 30705.0 59460.0 32050.0 ;
      RECT  58755.0 33395.0 59460.0 32050.0 ;
      RECT  58755.0 33395.0 59460.0 34740.0 ;
      RECT  58755.0 36085.0 59460.0 34740.0 ;
      RECT  58755.0 36085.0 59460.0 37430.0 ;
      RECT  58755.0 38775.0 59460.0 37430.0 ;
      RECT  58755.0 38775.0 59460.0 40120.0 ;
      RECT  58755.0 41465.0 59460.0 40120.0 ;
      RECT  58755.0 41465.0 59460.0 42810.0 ;
      RECT  58755.0 44155.0 59460.0 42810.0 ;
      RECT  58755.0 44155.0 59460.0 45500.0 ;
      RECT  58755.0 46845.0 59460.0 45500.0 ;
      RECT  58755.0 46845.0 59460.0 48190.0 ;
      RECT  58755.0 49535.0 59460.0 48190.0 ;
      RECT  58755.0 49535.0 59460.0 50880.0 ;
      RECT  58755.0 52225.0 59460.0 50880.0 ;
      RECT  58755.0 52225.0 59460.0 53570.0 ;
      RECT  58755.0 54915.0 59460.0 53570.0 ;
      RECT  58755.0 54915.0 59460.0 56260.0 ;
      RECT  58755.0 57605.0 59460.0 56260.0 ;
      RECT  58755.0 57605.0 59460.0 58950.0 ;
      RECT  58755.0 60295.0 59460.0 58950.0 ;
      RECT  58755.0 60295.0 59460.0 61640.0 ;
      RECT  58755.0 62985.0 59460.0 61640.0 ;
      RECT  58755.0 62985.0 59460.0 64330.0 ;
      RECT  58755.0 65675.0 59460.0 64330.0 ;
      RECT  58755.0 65675.0 59460.0 67020.0 ;
      RECT  58755.0 68365.0 59460.0 67020.0 ;
      RECT  58755.0 68365.0 59460.0 69710.0 ;
      RECT  58755.0 71055.0 59460.0 69710.0 ;
      RECT  58755.0 71055.0 59460.0 72400.0 ;
      RECT  58755.0 73745.0 59460.0 72400.0 ;
      RECT  58755.0 73745.0 59460.0 75090.0 ;
      RECT  58755.0 76435.0 59460.0 75090.0 ;
      RECT  58755.0 76435.0 59460.0 77780.0 ;
      RECT  58755.0 79125.0 59460.0 77780.0 ;
      RECT  58755.0 79125.0 59460.0 80470.0 ;
      RECT  58755.0 81815.0 59460.0 80470.0 ;
      RECT  58755.0 81815.0 59460.0 83160.0 ;
      RECT  58755.0 84505.0 59460.0 83160.0 ;
      RECT  58755.0 84505.0 59460.0 85850.0 ;
      RECT  58755.0 87195.0 59460.0 85850.0 ;
      RECT  58755.0 87195.0 59460.0 88540.0 ;
      RECT  58755.0 89885.0 59460.0 88540.0 ;
      RECT  58755.0 89885.0 59460.0 91230.0 ;
      RECT  58755.0 92575.0 59460.0 91230.0 ;
      RECT  58755.0 92575.0 59460.0 93920.0 ;
      RECT  58755.0 95265.0 59460.0 93920.0 ;
      RECT  58755.0 95265.0 59460.0 96610.0 ;
      RECT  58755.0 97955.0 59460.0 96610.0 ;
      RECT  58755.0 97955.0 59460.0 99300.0 ;
      RECT  58755.0 100645.0 59460.0 99300.0 ;
      RECT  58755.0 100645.0 59460.0 101990.0 ;
      RECT  58755.0 103335.0 59460.0 101990.0 ;
      RECT  58755.0 103335.0 59460.0 104680.0 ;
      RECT  58755.0 106025.0 59460.0 104680.0 ;
      RECT  58755.0 106025.0 59460.0 107370.0 ;
      RECT  58755.0 108715.0 59460.0 107370.0 ;
      RECT  58755.0 108715.0 59460.0 110060.0 ;
      RECT  58755.0 111405.0 59460.0 110060.0 ;
      RECT  58755.0 111405.0 59460.0 112750.0 ;
      RECT  58755.0 114095.0 59460.0 112750.0 ;
      RECT  59460.0 28015.0 60165.0 29360.0 ;
      RECT  59460.0 30705.0 60165.0 29360.0 ;
      RECT  59460.0 30705.0 60165.0 32050.0 ;
      RECT  59460.0 33395.0 60165.0 32050.0 ;
      RECT  59460.0 33395.0 60165.0 34740.0 ;
      RECT  59460.0 36085.0 60165.0 34740.0 ;
      RECT  59460.0 36085.0 60165.0 37430.0 ;
      RECT  59460.0 38775.0 60165.0 37430.0 ;
      RECT  59460.0 38775.0 60165.0 40120.0 ;
      RECT  59460.0 41465.0 60165.0 40120.0 ;
      RECT  59460.0 41465.0 60165.0 42810.0 ;
      RECT  59460.0 44155.0 60165.0 42810.0 ;
      RECT  59460.0 44155.0 60165.0 45500.0 ;
      RECT  59460.0 46845.0 60165.0 45500.0 ;
      RECT  59460.0 46845.0 60165.0 48190.0 ;
      RECT  59460.0 49535.0 60165.0 48190.0 ;
      RECT  59460.0 49535.0 60165.0 50880.0 ;
      RECT  59460.0 52225.0 60165.0 50880.0 ;
      RECT  59460.0 52225.0 60165.0 53570.0 ;
      RECT  59460.0 54915.0 60165.0 53570.0 ;
      RECT  59460.0 54915.0 60165.0 56260.0 ;
      RECT  59460.0 57605.0 60165.0 56260.0 ;
      RECT  59460.0 57605.0 60165.0 58950.0 ;
      RECT  59460.0 60295.0 60165.0 58950.0 ;
      RECT  59460.0 60295.0 60165.0 61640.0 ;
      RECT  59460.0 62985.0 60165.0 61640.0 ;
      RECT  59460.0 62985.0 60165.0 64330.0 ;
      RECT  59460.0 65675.0 60165.0 64330.0 ;
      RECT  59460.0 65675.0 60165.0 67020.0 ;
      RECT  59460.0 68365.0 60165.0 67020.0 ;
      RECT  59460.0 68365.0 60165.0 69710.0 ;
      RECT  59460.0 71055.0 60165.0 69710.0 ;
      RECT  59460.0 71055.0 60165.0 72400.0 ;
      RECT  59460.0 73745.0 60165.0 72400.0 ;
      RECT  59460.0 73745.0 60165.0 75090.0 ;
      RECT  59460.0 76435.0 60165.0 75090.0 ;
      RECT  59460.0 76435.0 60165.0 77780.0 ;
      RECT  59460.0 79125.0 60165.0 77780.0 ;
      RECT  59460.0 79125.0 60165.0 80470.0 ;
      RECT  59460.0 81815.0 60165.0 80470.0 ;
      RECT  59460.0 81815.0 60165.0 83160.0 ;
      RECT  59460.0 84505.0 60165.0 83160.0 ;
      RECT  59460.0 84505.0 60165.0 85850.0 ;
      RECT  59460.0 87195.0 60165.0 85850.0 ;
      RECT  59460.0 87195.0 60165.0 88540.0 ;
      RECT  59460.0 89885.0 60165.0 88540.0 ;
      RECT  59460.0 89885.0 60165.0 91230.0 ;
      RECT  59460.0 92575.0 60165.0 91230.0 ;
      RECT  59460.0 92575.0 60165.0 93920.0 ;
      RECT  59460.0 95265.0 60165.0 93920.0 ;
      RECT  59460.0 95265.0 60165.0 96610.0 ;
      RECT  59460.0 97955.0 60165.0 96610.0 ;
      RECT  59460.0 97955.0 60165.0 99300.0 ;
      RECT  59460.0 100645.0 60165.0 99300.0 ;
      RECT  59460.0 100645.0 60165.0 101990.0 ;
      RECT  59460.0 103335.0 60165.0 101990.0 ;
      RECT  59460.0 103335.0 60165.0 104680.0 ;
      RECT  59460.0 106025.0 60165.0 104680.0 ;
      RECT  59460.0 106025.0 60165.0 107370.0 ;
      RECT  59460.0 108715.0 60165.0 107370.0 ;
      RECT  59460.0 108715.0 60165.0 110060.0 ;
      RECT  59460.0 111405.0 60165.0 110060.0 ;
      RECT  59460.0 111405.0 60165.0 112750.0 ;
      RECT  59460.0 114095.0 60165.0 112750.0 ;
      RECT  60165.0 28015.0 60870.0 29360.0 ;
      RECT  60165.0 30705.0 60870.0 29360.0 ;
      RECT  60165.0 30705.0 60870.0 32050.0 ;
      RECT  60165.0 33395.0 60870.0 32050.0 ;
      RECT  60165.0 33395.0 60870.0 34740.0 ;
      RECT  60165.0 36085.0 60870.0 34740.0 ;
      RECT  60165.0 36085.0 60870.0 37430.0 ;
      RECT  60165.0 38775.0 60870.0 37430.0 ;
      RECT  60165.0 38775.0 60870.0 40120.0 ;
      RECT  60165.0 41465.0 60870.0 40120.0 ;
      RECT  60165.0 41465.0 60870.0 42810.0 ;
      RECT  60165.0 44155.0 60870.0 42810.0 ;
      RECT  60165.0 44155.0 60870.0 45500.0 ;
      RECT  60165.0 46845.0 60870.0 45500.0 ;
      RECT  60165.0 46845.0 60870.0 48190.0 ;
      RECT  60165.0 49535.0 60870.0 48190.0 ;
      RECT  60165.0 49535.0 60870.0 50880.0 ;
      RECT  60165.0 52225.0 60870.0 50880.0 ;
      RECT  60165.0 52225.0 60870.0 53570.0 ;
      RECT  60165.0 54915.0 60870.0 53570.0 ;
      RECT  60165.0 54915.0 60870.0 56260.0 ;
      RECT  60165.0 57605.0 60870.0 56260.0 ;
      RECT  60165.0 57605.0 60870.0 58950.0 ;
      RECT  60165.0 60295.0 60870.0 58950.0 ;
      RECT  60165.0 60295.0 60870.0 61640.0 ;
      RECT  60165.0 62985.0 60870.0 61640.0 ;
      RECT  60165.0 62985.0 60870.0 64330.0 ;
      RECT  60165.0 65675.0 60870.0 64330.0 ;
      RECT  60165.0 65675.0 60870.0 67020.0 ;
      RECT  60165.0 68365.0 60870.0 67020.0 ;
      RECT  60165.0 68365.0 60870.0 69710.0 ;
      RECT  60165.0 71055.0 60870.0 69710.0 ;
      RECT  60165.0 71055.0 60870.0 72400.0 ;
      RECT  60165.0 73745.0 60870.0 72400.0 ;
      RECT  60165.0 73745.0 60870.0 75090.0 ;
      RECT  60165.0 76435.0 60870.0 75090.0 ;
      RECT  60165.0 76435.0 60870.0 77780.0 ;
      RECT  60165.0 79125.0 60870.0 77780.0 ;
      RECT  60165.0 79125.0 60870.0 80470.0 ;
      RECT  60165.0 81815.0 60870.0 80470.0 ;
      RECT  60165.0 81815.0 60870.0 83160.0 ;
      RECT  60165.0 84505.0 60870.0 83160.0 ;
      RECT  60165.0 84505.0 60870.0 85850.0 ;
      RECT  60165.0 87195.0 60870.0 85850.0 ;
      RECT  60165.0 87195.0 60870.0 88540.0 ;
      RECT  60165.0 89885.0 60870.0 88540.0 ;
      RECT  60165.0 89885.0 60870.0 91230.0 ;
      RECT  60165.0 92575.0 60870.0 91230.0 ;
      RECT  60165.0 92575.0 60870.0 93920.0 ;
      RECT  60165.0 95265.0 60870.0 93920.0 ;
      RECT  60165.0 95265.0 60870.0 96610.0 ;
      RECT  60165.0 97955.0 60870.0 96610.0 ;
      RECT  60165.0 97955.0 60870.0 99300.0 ;
      RECT  60165.0 100645.0 60870.0 99300.0 ;
      RECT  60165.0 100645.0 60870.0 101990.0 ;
      RECT  60165.0 103335.0 60870.0 101990.0 ;
      RECT  60165.0 103335.0 60870.0 104680.0 ;
      RECT  60165.0 106025.0 60870.0 104680.0 ;
      RECT  60165.0 106025.0 60870.0 107370.0 ;
      RECT  60165.0 108715.0 60870.0 107370.0 ;
      RECT  60165.0 108715.0 60870.0 110060.0 ;
      RECT  60165.0 111405.0 60870.0 110060.0 ;
      RECT  60165.0 111405.0 60870.0 112750.0 ;
      RECT  60165.0 114095.0 60870.0 112750.0 ;
      RECT  60870.0 28015.0 61575.0 29360.0 ;
      RECT  60870.0 30705.0 61575.0 29360.0 ;
      RECT  60870.0 30705.0 61575.0 32050.0 ;
      RECT  60870.0 33395.0 61575.0 32050.0 ;
      RECT  60870.0 33395.0 61575.0 34740.0 ;
      RECT  60870.0 36085.0 61575.0 34740.0 ;
      RECT  60870.0 36085.0 61575.0 37430.0 ;
      RECT  60870.0 38775.0 61575.0 37430.0 ;
      RECT  60870.0 38775.0 61575.0 40120.0 ;
      RECT  60870.0 41465.0 61575.0 40120.0 ;
      RECT  60870.0 41465.0 61575.0 42810.0 ;
      RECT  60870.0 44155.0 61575.0 42810.0 ;
      RECT  60870.0 44155.0 61575.0 45500.0 ;
      RECT  60870.0 46845.0 61575.0 45500.0 ;
      RECT  60870.0 46845.0 61575.0 48190.0 ;
      RECT  60870.0 49535.0 61575.0 48190.0 ;
      RECT  60870.0 49535.0 61575.0 50880.0 ;
      RECT  60870.0 52225.0 61575.0 50880.0 ;
      RECT  60870.0 52225.0 61575.0 53570.0 ;
      RECT  60870.0 54915.0 61575.0 53570.0 ;
      RECT  60870.0 54915.0 61575.0 56260.0 ;
      RECT  60870.0 57605.0 61575.0 56260.0 ;
      RECT  60870.0 57605.0 61575.0 58950.0 ;
      RECT  60870.0 60295.0 61575.0 58950.0 ;
      RECT  60870.0 60295.0 61575.0 61640.0 ;
      RECT  60870.0 62985.0 61575.0 61640.0 ;
      RECT  60870.0 62985.0 61575.0 64330.0 ;
      RECT  60870.0 65675.0 61575.0 64330.0 ;
      RECT  60870.0 65675.0 61575.0 67020.0 ;
      RECT  60870.0 68365.0 61575.0 67020.0 ;
      RECT  60870.0 68365.0 61575.0 69710.0 ;
      RECT  60870.0 71055.0 61575.0 69710.0 ;
      RECT  60870.0 71055.0 61575.0 72400.0 ;
      RECT  60870.0 73745.0 61575.0 72400.0 ;
      RECT  60870.0 73745.0 61575.0 75090.0 ;
      RECT  60870.0 76435.0 61575.0 75090.0 ;
      RECT  60870.0 76435.0 61575.0 77780.0 ;
      RECT  60870.0 79125.0 61575.0 77780.0 ;
      RECT  60870.0 79125.0 61575.0 80470.0 ;
      RECT  60870.0 81815.0 61575.0 80470.0 ;
      RECT  60870.0 81815.0 61575.0 83160.0 ;
      RECT  60870.0 84505.0 61575.0 83160.0 ;
      RECT  60870.0 84505.0 61575.0 85850.0 ;
      RECT  60870.0 87195.0 61575.0 85850.0 ;
      RECT  60870.0 87195.0 61575.0 88540.0 ;
      RECT  60870.0 89885.0 61575.0 88540.0 ;
      RECT  60870.0 89885.0 61575.0 91230.0 ;
      RECT  60870.0 92575.0 61575.0 91230.0 ;
      RECT  60870.0 92575.0 61575.0 93920.0 ;
      RECT  60870.0 95265.0 61575.0 93920.0 ;
      RECT  60870.0 95265.0 61575.0 96610.0 ;
      RECT  60870.0 97955.0 61575.0 96610.0 ;
      RECT  60870.0 97955.0 61575.0 99300.0 ;
      RECT  60870.0 100645.0 61575.0 99300.0 ;
      RECT  60870.0 100645.0 61575.0 101990.0 ;
      RECT  60870.0 103335.0 61575.0 101990.0 ;
      RECT  60870.0 103335.0 61575.0 104680.0 ;
      RECT  60870.0 106025.0 61575.0 104680.0 ;
      RECT  60870.0 106025.0 61575.0 107370.0 ;
      RECT  60870.0 108715.0 61575.0 107370.0 ;
      RECT  60870.0 108715.0 61575.0 110060.0 ;
      RECT  60870.0 111405.0 61575.0 110060.0 ;
      RECT  60870.0 111405.0 61575.0 112750.0 ;
      RECT  60870.0 114095.0 61575.0 112750.0 ;
      RECT  61575.0 28015.0 62280.0 29360.0 ;
      RECT  61575.0 30705.0 62280.0 29360.0 ;
      RECT  61575.0 30705.0 62280.0 32050.0 ;
      RECT  61575.0 33395.0 62280.0 32050.0 ;
      RECT  61575.0 33395.0 62280.0 34740.0 ;
      RECT  61575.0 36085.0 62280.0 34740.0 ;
      RECT  61575.0 36085.0 62280.0 37430.0 ;
      RECT  61575.0 38775.0 62280.0 37430.0 ;
      RECT  61575.0 38775.0 62280.0 40120.0 ;
      RECT  61575.0 41465.0 62280.0 40120.0 ;
      RECT  61575.0 41465.0 62280.0 42810.0 ;
      RECT  61575.0 44155.0 62280.0 42810.0 ;
      RECT  61575.0 44155.0 62280.0 45500.0 ;
      RECT  61575.0 46845.0 62280.0 45500.0 ;
      RECT  61575.0 46845.0 62280.0 48190.0 ;
      RECT  61575.0 49535.0 62280.0 48190.0 ;
      RECT  61575.0 49535.0 62280.0 50880.0 ;
      RECT  61575.0 52225.0 62280.0 50880.0 ;
      RECT  61575.0 52225.0 62280.0 53570.0 ;
      RECT  61575.0 54915.0 62280.0 53570.0 ;
      RECT  61575.0 54915.0 62280.0 56260.0 ;
      RECT  61575.0 57605.0 62280.0 56260.0 ;
      RECT  61575.0 57605.0 62280.0 58950.0 ;
      RECT  61575.0 60295.0 62280.0 58950.0 ;
      RECT  61575.0 60295.0 62280.0 61640.0 ;
      RECT  61575.0 62985.0 62280.0 61640.0 ;
      RECT  61575.0 62985.0 62280.0 64330.0 ;
      RECT  61575.0 65675.0 62280.0 64330.0 ;
      RECT  61575.0 65675.0 62280.0 67020.0 ;
      RECT  61575.0 68365.0 62280.0 67020.0 ;
      RECT  61575.0 68365.0 62280.0 69710.0 ;
      RECT  61575.0 71055.0 62280.0 69710.0 ;
      RECT  61575.0 71055.0 62280.0 72400.0 ;
      RECT  61575.0 73745.0 62280.0 72400.0 ;
      RECT  61575.0 73745.0 62280.0 75090.0 ;
      RECT  61575.0 76435.0 62280.0 75090.0 ;
      RECT  61575.0 76435.0 62280.0 77780.0 ;
      RECT  61575.0 79125.0 62280.0 77780.0 ;
      RECT  61575.0 79125.0 62280.0 80470.0 ;
      RECT  61575.0 81815.0 62280.0 80470.0 ;
      RECT  61575.0 81815.0 62280.0 83160.0 ;
      RECT  61575.0 84505.0 62280.0 83160.0 ;
      RECT  61575.0 84505.0 62280.0 85850.0 ;
      RECT  61575.0 87195.0 62280.0 85850.0 ;
      RECT  61575.0 87195.0 62280.0 88540.0 ;
      RECT  61575.0 89885.0 62280.0 88540.0 ;
      RECT  61575.0 89885.0 62280.0 91230.0 ;
      RECT  61575.0 92575.0 62280.0 91230.0 ;
      RECT  61575.0 92575.0 62280.0 93920.0 ;
      RECT  61575.0 95265.0 62280.0 93920.0 ;
      RECT  61575.0 95265.0 62280.0 96610.0 ;
      RECT  61575.0 97955.0 62280.0 96610.0 ;
      RECT  61575.0 97955.0 62280.0 99300.0 ;
      RECT  61575.0 100645.0 62280.0 99300.0 ;
      RECT  61575.0 100645.0 62280.0 101990.0 ;
      RECT  61575.0 103335.0 62280.0 101990.0 ;
      RECT  61575.0 103335.0 62280.0 104680.0 ;
      RECT  61575.0 106025.0 62280.0 104680.0 ;
      RECT  61575.0 106025.0 62280.0 107370.0 ;
      RECT  61575.0 108715.0 62280.0 107370.0 ;
      RECT  61575.0 108715.0 62280.0 110060.0 ;
      RECT  61575.0 111405.0 62280.0 110060.0 ;
      RECT  61575.0 111405.0 62280.0 112750.0 ;
      RECT  61575.0 114095.0 62280.0 112750.0 ;
      RECT  62280.0 28015.0 62985.0 29360.0 ;
      RECT  62280.0 30705.0 62985.0 29360.0 ;
      RECT  62280.0 30705.0 62985.0 32050.0 ;
      RECT  62280.0 33395.0 62985.0 32050.0 ;
      RECT  62280.0 33395.0 62985.0 34740.0 ;
      RECT  62280.0 36085.0 62985.0 34740.0 ;
      RECT  62280.0 36085.0 62985.0 37430.0 ;
      RECT  62280.0 38775.0 62985.0 37430.0 ;
      RECT  62280.0 38775.0 62985.0 40120.0 ;
      RECT  62280.0 41465.0 62985.0 40120.0 ;
      RECT  62280.0 41465.0 62985.0 42810.0 ;
      RECT  62280.0 44155.0 62985.0 42810.0 ;
      RECT  62280.0 44155.0 62985.0 45500.0 ;
      RECT  62280.0 46845.0 62985.0 45500.0 ;
      RECT  62280.0 46845.0 62985.0 48190.0 ;
      RECT  62280.0 49535.0 62985.0 48190.0 ;
      RECT  62280.0 49535.0 62985.0 50880.0 ;
      RECT  62280.0 52225.0 62985.0 50880.0 ;
      RECT  62280.0 52225.0 62985.0 53570.0 ;
      RECT  62280.0 54915.0 62985.0 53570.0 ;
      RECT  62280.0 54915.0 62985.0 56260.0 ;
      RECT  62280.0 57605.0 62985.0 56260.0 ;
      RECT  62280.0 57605.0 62985.0 58950.0 ;
      RECT  62280.0 60295.0 62985.0 58950.0 ;
      RECT  62280.0 60295.0 62985.0 61640.0 ;
      RECT  62280.0 62985.0 62985.0 61640.0 ;
      RECT  62280.0 62985.0 62985.0 64330.0 ;
      RECT  62280.0 65675.0 62985.0 64330.0 ;
      RECT  62280.0 65675.0 62985.0 67020.0 ;
      RECT  62280.0 68365.0 62985.0 67020.0 ;
      RECT  62280.0 68365.0 62985.0 69710.0 ;
      RECT  62280.0 71055.0 62985.0 69710.0 ;
      RECT  62280.0 71055.0 62985.0 72400.0 ;
      RECT  62280.0 73745.0 62985.0 72400.0 ;
      RECT  62280.0 73745.0 62985.0 75090.0 ;
      RECT  62280.0 76435.0 62985.0 75090.0 ;
      RECT  62280.0 76435.0 62985.0 77780.0 ;
      RECT  62280.0 79125.0 62985.0 77780.0 ;
      RECT  62280.0 79125.0 62985.0 80470.0 ;
      RECT  62280.0 81815.0 62985.0 80470.0 ;
      RECT  62280.0 81815.0 62985.0 83160.0 ;
      RECT  62280.0 84505.0 62985.0 83160.0 ;
      RECT  62280.0 84505.0 62985.0 85850.0 ;
      RECT  62280.0 87195.0 62985.0 85850.0 ;
      RECT  62280.0 87195.0 62985.0 88540.0 ;
      RECT  62280.0 89885.0 62985.0 88540.0 ;
      RECT  62280.0 89885.0 62985.0 91230.0 ;
      RECT  62280.0 92575.0 62985.0 91230.0 ;
      RECT  62280.0 92575.0 62985.0 93920.0 ;
      RECT  62280.0 95265.0 62985.0 93920.0 ;
      RECT  62280.0 95265.0 62985.0 96610.0 ;
      RECT  62280.0 97955.0 62985.0 96610.0 ;
      RECT  62280.0 97955.0 62985.0 99300.0 ;
      RECT  62280.0 100645.0 62985.0 99300.0 ;
      RECT  62280.0 100645.0 62985.0 101990.0 ;
      RECT  62280.0 103335.0 62985.0 101990.0 ;
      RECT  62280.0 103335.0 62985.0 104680.0 ;
      RECT  62280.0 106025.0 62985.0 104680.0 ;
      RECT  62280.0 106025.0 62985.0 107370.0 ;
      RECT  62280.0 108715.0 62985.0 107370.0 ;
      RECT  62280.0 108715.0 62985.0 110060.0 ;
      RECT  62280.0 111405.0 62985.0 110060.0 ;
      RECT  62280.0 111405.0 62985.0 112750.0 ;
      RECT  62280.0 114095.0 62985.0 112750.0 ;
      RECT  62985.0 28015.0 63690.0 29360.0 ;
      RECT  62985.0 30705.0 63690.0 29360.0 ;
      RECT  62985.0 30705.0 63690.0 32050.0 ;
      RECT  62985.0 33395.0 63690.0 32050.0 ;
      RECT  62985.0 33395.0 63690.0 34740.0 ;
      RECT  62985.0 36085.0 63690.0 34740.0 ;
      RECT  62985.0 36085.0 63690.0 37430.0 ;
      RECT  62985.0 38775.0 63690.0 37430.0 ;
      RECT  62985.0 38775.0 63690.0 40120.0 ;
      RECT  62985.0 41465.0 63690.0 40120.0 ;
      RECT  62985.0 41465.0 63690.0 42810.0 ;
      RECT  62985.0 44155.0 63690.0 42810.0 ;
      RECT  62985.0 44155.0 63690.0 45500.0 ;
      RECT  62985.0 46845.0 63690.0 45500.0 ;
      RECT  62985.0 46845.0 63690.0 48190.0 ;
      RECT  62985.0 49535.0 63690.0 48190.0 ;
      RECT  62985.0 49535.0 63690.0 50880.0 ;
      RECT  62985.0 52225.0 63690.0 50880.0 ;
      RECT  62985.0 52225.0 63690.0 53570.0 ;
      RECT  62985.0 54915.0 63690.0 53570.0 ;
      RECT  62985.0 54915.0 63690.0 56260.0 ;
      RECT  62985.0 57605.0 63690.0 56260.0 ;
      RECT  62985.0 57605.0 63690.0 58950.0 ;
      RECT  62985.0 60295.0 63690.0 58950.0 ;
      RECT  62985.0 60295.0 63690.0 61640.0 ;
      RECT  62985.0 62985.0 63690.0 61640.0 ;
      RECT  62985.0 62985.0 63690.0 64330.0 ;
      RECT  62985.0 65675.0 63690.0 64330.0 ;
      RECT  62985.0 65675.0 63690.0 67020.0 ;
      RECT  62985.0 68365.0 63690.0 67020.0 ;
      RECT  62985.0 68365.0 63690.0 69710.0 ;
      RECT  62985.0 71055.0 63690.0 69710.0 ;
      RECT  62985.0 71055.0 63690.0 72400.0 ;
      RECT  62985.0 73745.0 63690.0 72400.0 ;
      RECT  62985.0 73745.0 63690.0 75090.0 ;
      RECT  62985.0 76435.0 63690.0 75090.0 ;
      RECT  62985.0 76435.0 63690.0 77780.0 ;
      RECT  62985.0 79125.0 63690.0 77780.0 ;
      RECT  62985.0 79125.0 63690.0 80470.0 ;
      RECT  62985.0 81815.0 63690.0 80470.0 ;
      RECT  62985.0 81815.0 63690.0 83160.0 ;
      RECT  62985.0 84505.0 63690.0 83160.0 ;
      RECT  62985.0 84505.0 63690.0 85850.0 ;
      RECT  62985.0 87195.0 63690.0 85850.0 ;
      RECT  62985.0 87195.0 63690.0 88540.0 ;
      RECT  62985.0 89885.0 63690.0 88540.0 ;
      RECT  62985.0 89885.0 63690.0 91230.0 ;
      RECT  62985.0 92575.0 63690.0 91230.0 ;
      RECT  62985.0 92575.0 63690.0 93920.0 ;
      RECT  62985.0 95265.0 63690.0 93920.0 ;
      RECT  62985.0 95265.0 63690.0 96610.0 ;
      RECT  62985.0 97955.0 63690.0 96610.0 ;
      RECT  62985.0 97955.0 63690.0 99300.0 ;
      RECT  62985.0 100645.0 63690.0 99300.0 ;
      RECT  62985.0 100645.0 63690.0 101990.0 ;
      RECT  62985.0 103335.0 63690.0 101990.0 ;
      RECT  62985.0 103335.0 63690.0 104680.0 ;
      RECT  62985.0 106025.0 63690.0 104680.0 ;
      RECT  62985.0 106025.0 63690.0 107370.0 ;
      RECT  62985.0 108715.0 63690.0 107370.0 ;
      RECT  62985.0 108715.0 63690.0 110060.0 ;
      RECT  62985.0 111405.0 63690.0 110060.0 ;
      RECT  62985.0 111405.0 63690.0 112750.0 ;
      RECT  62985.0 114095.0 63690.0 112750.0 ;
      RECT  63690.0 28015.0 64395.0 29360.0 ;
      RECT  63690.0 30705.0 64395.0 29360.0 ;
      RECT  63690.0 30705.0 64395.0 32050.0 ;
      RECT  63690.0 33395.0 64395.0 32050.0 ;
      RECT  63690.0 33395.0 64395.0 34740.0 ;
      RECT  63690.0 36085.0 64395.0 34740.0 ;
      RECT  63690.0 36085.0 64395.0 37430.0 ;
      RECT  63690.0 38775.0 64395.0 37430.0 ;
      RECT  63690.0 38775.0 64395.0 40120.0 ;
      RECT  63690.0 41465.0 64395.0 40120.0 ;
      RECT  63690.0 41465.0 64395.0 42810.0 ;
      RECT  63690.0 44155.0 64395.0 42810.0 ;
      RECT  63690.0 44155.0 64395.0 45500.0 ;
      RECT  63690.0 46845.0 64395.0 45500.0 ;
      RECT  63690.0 46845.0 64395.0 48190.0 ;
      RECT  63690.0 49535.0 64395.0 48190.0 ;
      RECT  63690.0 49535.0 64395.0 50880.0 ;
      RECT  63690.0 52225.0 64395.0 50880.0 ;
      RECT  63690.0 52225.0 64395.0 53570.0 ;
      RECT  63690.0 54915.0 64395.0 53570.0 ;
      RECT  63690.0 54915.0 64395.0 56260.0 ;
      RECT  63690.0 57605.0 64395.0 56260.0 ;
      RECT  63690.0 57605.0 64395.0 58950.0 ;
      RECT  63690.0 60295.0 64395.0 58950.0 ;
      RECT  63690.0 60295.0 64395.0 61640.0 ;
      RECT  63690.0 62985.0 64395.0 61640.0 ;
      RECT  63690.0 62985.0 64395.0 64330.0 ;
      RECT  63690.0 65675.0 64395.0 64330.0 ;
      RECT  63690.0 65675.0 64395.0 67020.0 ;
      RECT  63690.0 68365.0 64395.0 67020.0 ;
      RECT  63690.0 68365.0 64395.0 69710.0 ;
      RECT  63690.0 71055.0 64395.0 69710.0 ;
      RECT  63690.0 71055.0 64395.0 72400.0 ;
      RECT  63690.0 73745.0 64395.0 72400.0 ;
      RECT  63690.0 73745.0 64395.0 75090.0 ;
      RECT  63690.0 76435.0 64395.0 75090.0 ;
      RECT  63690.0 76435.0 64395.0 77780.0 ;
      RECT  63690.0 79125.0 64395.0 77780.0 ;
      RECT  63690.0 79125.0 64395.0 80470.0 ;
      RECT  63690.0 81815.0 64395.0 80470.0 ;
      RECT  63690.0 81815.0 64395.0 83160.0 ;
      RECT  63690.0 84505.0 64395.0 83160.0 ;
      RECT  63690.0 84505.0 64395.0 85850.0 ;
      RECT  63690.0 87195.0 64395.0 85850.0 ;
      RECT  63690.0 87195.0 64395.0 88540.0 ;
      RECT  63690.0 89885.0 64395.0 88540.0 ;
      RECT  63690.0 89885.0 64395.0 91230.0 ;
      RECT  63690.0 92575.0 64395.0 91230.0 ;
      RECT  63690.0 92575.0 64395.0 93920.0 ;
      RECT  63690.0 95265.0 64395.0 93920.0 ;
      RECT  63690.0 95265.0 64395.0 96610.0 ;
      RECT  63690.0 97955.0 64395.0 96610.0 ;
      RECT  63690.0 97955.0 64395.0 99300.0 ;
      RECT  63690.0 100645.0 64395.0 99300.0 ;
      RECT  63690.0 100645.0 64395.0 101990.0 ;
      RECT  63690.0 103335.0 64395.0 101990.0 ;
      RECT  63690.0 103335.0 64395.0 104680.0 ;
      RECT  63690.0 106025.0 64395.0 104680.0 ;
      RECT  63690.0 106025.0 64395.0 107370.0 ;
      RECT  63690.0 108715.0 64395.0 107370.0 ;
      RECT  63690.0 108715.0 64395.0 110060.0 ;
      RECT  63690.0 111405.0 64395.0 110060.0 ;
      RECT  63690.0 111405.0 64395.0 112750.0 ;
      RECT  63690.0 114095.0 64395.0 112750.0 ;
      RECT  64395.0 28015.0 65100.0 29360.0 ;
      RECT  64395.0 30705.0 65100.0 29360.0 ;
      RECT  64395.0 30705.0 65100.0 32050.0 ;
      RECT  64395.0 33395.0 65100.0 32050.0 ;
      RECT  64395.0 33395.0 65100.0 34740.0 ;
      RECT  64395.0 36085.0 65100.0 34740.0 ;
      RECT  64395.0 36085.0 65100.0 37430.0 ;
      RECT  64395.0 38775.0 65100.0 37430.0 ;
      RECT  64395.0 38775.0 65100.0 40120.0 ;
      RECT  64395.0 41465.0 65100.0 40120.0 ;
      RECT  64395.0 41465.0 65100.0 42810.0 ;
      RECT  64395.0 44155.0 65100.0 42810.0 ;
      RECT  64395.0 44155.0 65100.0 45500.0 ;
      RECT  64395.0 46845.0 65100.0 45500.0 ;
      RECT  64395.0 46845.0 65100.0 48190.0 ;
      RECT  64395.0 49535.0 65100.0 48190.0 ;
      RECT  64395.0 49535.0 65100.0 50880.0 ;
      RECT  64395.0 52225.0 65100.0 50880.0 ;
      RECT  64395.0 52225.0 65100.0 53570.0 ;
      RECT  64395.0 54915.0 65100.0 53570.0 ;
      RECT  64395.0 54915.0 65100.0 56260.0 ;
      RECT  64395.0 57605.0 65100.0 56260.0 ;
      RECT  64395.0 57605.0 65100.0 58950.0 ;
      RECT  64395.0 60295.0 65100.0 58950.0 ;
      RECT  64395.0 60295.0 65100.0 61640.0 ;
      RECT  64395.0 62985.0 65100.0 61640.0 ;
      RECT  64395.0 62985.0 65100.0 64330.0 ;
      RECT  64395.0 65675.0 65100.0 64330.0 ;
      RECT  64395.0 65675.0 65100.0 67020.0 ;
      RECT  64395.0 68365.0 65100.0 67020.0 ;
      RECT  64395.0 68365.0 65100.0 69710.0 ;
      RECT  64395.0 71055.0 65100.0 69710.0 ;
      RECT  64395.0 71055.0 65100.0 72400.0 ;
      RECT  64395.0 73745.0 65100.0 72400.0 ;
      RECT  64395.0 73745.0 65100.0 75090.0 ;
      RECT  64395.0 76435.0 65100.0 75090.0 ;
      RECT  64395.0 76435.0 65100.0 77780.0 ;
      RECT  64395.0 79125.0 65100.0 77780.0 ;
      RECT  64395.0 79125.0 65100.0 80470.0 ;
      RECT  64395.0 81815.0 65100.0 80470.0 ;
      RECT  64395.0 81815.0 65100.0 83160.0 ;
      RECT  64395.0 84505.0 65100.0 83160.0 ;
      RECT  64395.0 84505.0 65100.0 85850.0 ;
      RECT  64395.0 87195.0 65100.0 85850.0 ;
      RECT  64395.0 87195.0 65100.0 88540.0 ;
      RECT  64395.0 89885.0 65100.0 88540.0 ;
      RECT  64395.0 89885.0 65100.0 91230.0 ;
      RECT  64395.0 92575.0 65100.0 91230.0 ;
      RECT  64395.0 92575.0 65100.0 93920.0 ;
      RECT  64395.0 95265.0 65100.0 93920.0 ;
      RECT  64395.0 95265.0 65100.0 96610.0 ;
      RECT  64395.0 97955.0 65100.0 96610.0 ;
      RECT  64395.0 97955.0 65100.0 99300.0 ;
      RECT  64395.0 100645.0 65100.0 99300.0 ;
      RECT  64395.0 100645.0 65100.0 101990.0 ;
      RECT  64395.0 103335.0 65100.0 101990.0 ;
      RECT  64395.0 103335.0 65100.0 104680.0 ;
      RECT  64395.0 106025.0 65100.0 104680.0 ;
      RECT  64395.0 106025.0 65100.0 107370.0 ;
      RECT  64395.0 108715.0 65100.0 107370.0 ;
      RECT  64395.0 108715.0 65100.0 110060.0 ;
      RECT  64395.0 111405.0 65100.0 110060.0 ;
      RECT  64395.0 111405.0 65100.0 112750.0 ;
      RECT  64395.0 114095.0 65100.0 112750.0 ;
      RECT  65100.0 28015.0 65805.0 29360.0 ;
      RECT  65100.0 30705.0 65805.0 29360.0 ;
      RECT  65100.0 30705.0 65805.0 32050.0 ;
      RECT  65100.0 33395.0 65805.0 32050.0 ;
      RECT  65100.0 33395.0 65805.0 34740.0 ;
      RECT  65100.0 36085.0 65805.0 34740.0 ;
      RECT  65100.0 36085.0 65805.0 37430.0 ;
      RECT  65100.0 38775.0 65805.0 37430.0 ;
      RECT  65100.0 38775.0 65805.0 40120.0 ;
      RECT  65100.0 41465.0 65805.0 40120.0 ;
      RECT  65100.0 41465.0 65805.0 42810.0 ;
      RECT  65100.0 44155.0 65805.0 42810.0 ;
      RECT  65100.0 44155.0 65805.0 45500.0 ;
      RECT  65100.0 46845.0 65805.0 45500.0 ;
      RECT  65100.0 46845.0 65805.0 48190.0 ;
      RECT  65100.0 49535.0 65805.0 48190.0 ;
      RECT  65100.0 49535.0 65805.0 50880.0 ;
      RECT  65100.0 52225.0 65805.0 50880.0 ;
      RECT  65100.0 52225.0 65805.0 53570.0 ;
      RECT  65100.0 54915.0 65805.0 53570.0 ;
      RECT  65100.0 54915.0 65805.0 56260.0 ;
      RECT  65100.0 57605.0 65805.0 56260.0 ;
      RECT  65100.0 57605.0 65805.0 58950.0 ;
      RECT  65100.0 60295.0 65805.0 58950.0 ;
      RECT  65100.0 60295.0 65805.0 61640.0 ;
      RECT  65100.0 62985.0 65805.0 61640.0 ;
      RECT  65100.0 62985.0 65805.0 64330.0 ;
      RECT  65100.0 65675.0 65805.0 64330.0 ;
      RECT  65100.0 65675.0 65805.0 67020.0 ;
      RECT  65100.0 68365.0 65805.0 67020.0 ;
      RECT  65100.0 68365.0 65805.0 69710.0 ;
      RECT  65100.0 71055.0 65805.0 69710.0 ;
      RECT  65100.0 71055.0 65805.0 72400.0 ;
      RECT  65100.0 73745.0 65805.0 72400.0 ;
      RECT  65100.0 73745.0 65805.0 75090.0 ;
      RECT  65100.0 76435.0 65805.0 75090.0 ;
      RECT  65100.0 76435.0 65805.0 77780.0 ;
      RECT  65100.0 79125.0 65805.0 77780.0 ;
      RECT  65100.0 79125.0 65805.0 80470.0 ;
      RECT  65100.0 81815.0 65805.0 80470.0 ;
      RECT  65100.0 81815.0 65805.0 83160.0 ;
      RECT  65100.0 84505.0 65805.0 83160.0 ;
      RECT  65100.0 84505.0 65805.0 85850.0 ;
      RECT  65100.0 87195.0 65805.0 85850.0 ;
      RECT  65100.0 87195.0 65805.0 88540.0 ;
      RECT  65100.0 89885.0 65805.0 88540.0 ;
      RECT  65100.0 89885.0 65805.0 91230.0 ;
      RECT  65100.0 92575.0 65805.0 91230.0 ;
      RECT  65100.0 92575.0 65805.0 93920.0 ;
      RECT  65100.0 95265.0 65805.0 93920.0 ;
      RECT  65100.0 95265.0 65805.0 96610.0 ;
      RECT  65100.0 97955.0 65805.0 96610.0 ;
      RECT  65100.0 97955.0 65805.0 99300.0 ;
      RECT  65100.0 100645.0 65805.0 99300.0 ;
      RECT  65100.0 100645.0 65805.0 101990.0 ;
      RECT  65100.0 103335.0 65805.0 101990.0 ;
      RECT  65100.0 103335.0 65805.0 104680.0 ;
      RECT  65100.0 106025.0 65805.0 104680.0 ;
      RECT  65100.0 106025.0 65805.0 107370.0 ;
      RECT  65100.0 108715.0 65805.0 107370.0 ;
      RECT  65100.0 108715.0 65805.0 110060.0 ;
      RECT  65100.0 111405.0 65805.0 110060.0 ;
      RECT  65100.0 111405.0 65805.0 112750.0 ;
      RECT  65100.0 114095.0 65805.0 112750.0 ;
      RECT  65805.0 28015.0 66510.0 29360.0 ;
      RECT  65805.0 30705.0 66510.0 29360.0 ;
      RECT  65805.0 30705.0 66510.0 32050.0 ;
      RECT  65805.0 33395.0 66510.0 32050.0 ;
      RECT  65805.0 33395.0 66510.0 34740.0 ;
      RECT  65805.0 36085.0 66510.0 34740.0 ;
      RECT  65805.0 36085.0 66510.0 37430.0 ;
      RECT  65805.0 38775.0 66510.0 37430.0 ;
      RECT  65805.0 38775.0 66510.0 40120.0 ;
      RECT  65805.0 41465.0 66510.0 40120.0 ;
      RECT  65805.0 41465.0 66510.0 42810.0 ;
      RECT  65805.0 44155.0 66510.0 42810.0 ;
      RECT  65805.0 44155.0 66510.0 45500.0 ;
      RECT  65805.0 46845.0 66510.0 45500.0 ;
      RECT  65805.0 46845.0 66510.0 48190.0 ;
      RECT  65805.0 49535.0 66510.0 48190.0 ;
      RECT  65805.0 49535.0 66510.0 50880.0 ;
      RECT  65805.0 52225.0 66510.0 50880.0 ;
      RECT  65805.0 52225.0 66510.0 53570.0 ;
      RECT  65805.0 54915.0 66510.0 53570.0 ;
      RECT  65805.0 54915.0 66510.0 56260.0 ;
      RECT  65805.0 57605.0 66510.0 56260.0 ;
      RECT  65805.0 57605.0 66510.0 58950.0 ;
      RECT  65805.0 60295.0 66510.0 58950.0 ;
      RECT  65805.0 60295.0 66510.0 61640.0 ;
      RECT  65805.0 62985.0 66510.0 61640.0 ;
      RECT  65805.0 62985.0 66510.0 64330.0 ;
      RECT  65805.0 65675.0 66510.0 64330.0 ;
      RECT  65805.0 65675.0 66510.0 67020.0 ;
      RECT  65805.0 68365.0 66510.0 67020.0 ;
      RECT  65805.0 68365.0 66510.0 69710.0 ;
      RECT  65805.0 71055.0 66510.0 69710.0 ;
      RECT  65805.0 71055.0 66510.0 72400.0 ;
      RECT  65805.0 73745.0 66510.0 72400.0 ;
      RECT  65805.0 73745.0 66510.0 75090.0 ;
      RECT  65805.0 76435.0 66510.0 75090.0 ;
      RECT  65805.0 76435.0 66510.0 77780.0 ;
      RECT  65805.0 79125.0 66510.0 77780.0 ;
      RECT  65805.0 79125.0 66510.0 80470.0 ;
      RECT  65805.0 81815.0 66510.0 80470.0 ;
      RECT  65805.0 81815.0 66510.0 83160.0 ;
      RECT  65805.0 84505.0 66510.0 83160.0 ;
      RECT  65805.0 84505.0 66510.0 85850.0 ;
      RECT  65805.0 87195.0 66510.0 85850.0 ;
      RECT  65805.0 87195.0 66510.0 88540.0 ;
      RECT  65805.0 89885.0 66510.0 88540.0 ;
      RECT  65805.0 89885.0 66510.0 91230.0 ;
      RECT  65805.0 92575.0 66510.0 91230.0 ;
      RECT  65805.0 92575.0 66510.0 93920.0 ;
      RECT  65805.0 95265.0 66510.0 93920.0 ;
      RECT  65805.0 95265.0 66510.0 96610.0 ;
      RECT  65805.0 97955.0 66510.0 96610.0 ;
      RECT  65805.0 97955.0 66510.0 99300.0 ;
      RECT  65805.0 100645.0 66510.0 99300.0 ;
      RECT  65805.0 100645.0 66510.0 101990.0 ;
      RECT  65805.0 103335.0 66510.0 101990.0 ;
      RECT  65805.0 103335.0 66510.0 104680.0 ;
      RECT  65805.0 106025.0 66510.0 104680.0 ;
      RECT  65805.0 106025.0 66510.0 107370.0 ;
      RECT  65805.0 108715.0 66510.0 107370.0 ;
      RECT  65805.0 108715.0 66510.0 110060.0 ;
      RECT  65805.0 111405.0 66510.0 110060.0 ;
      RECT  65805.0 111405.0 66510.0 112750.0 ;
      RECT  65805.0 114095.0 66510.0 112750.0 ;
      RECT  66510.0 28015.0 67215.0 29360.0 ;
      RECT  66510.0 30705.0 67215.0 29360.0 ;
      RECT  66510.0 30705.0 67215.0 32050.0 ;
      RECT  66510.0 33395.0 67215.0 32050.0 ;
      RECT  66510.0 33395.0 67215.0 34740.0 ;
      RECT  66510.0 36085.0 67215.0 34740.0 ;
      RECT  66510.0 36085.0 67215.0 37430.0 ;
      RECT  66510.0 38775.0 67215.0 37430.0 ;
      RECT  66510.0 38775.0 67215.0 40120.0 ;
      RECT  66510.0 41465.0 67215.0 40120.0 ;
      RECT  66510.0 41465.0 67215.0 42810.0 ;
      RECT  66510.0 44155.0 67215.0 42810.0 ;
      RECT  66510.0 44155.0 67215.0 45500.0 ;
      RECT  66510.0 46845.0 67215.0 45500.0 ;
      RECT  66510.0 46845.0 67215.0 48190.0 ;
      RECT  66510.0 49535.0 67215.0 48190.0 ;
      RECT  66510.0 49535.0 67215.0 50880.0 ;
      RECT  66510.0 52225.0 67215.0 50880.0 ;
      RECT  66510.0 52225.0 67215.0 53570.0 ;
      RECT  66510.0 54915.0 67215.0 53570.0 ;
      RECT  66510.0 54915.0 67215.0 56260.0 ;
      RECT  66510.0 57605.0 67215.0 56260.0 ;
      RECT  66510.0 57605.0 67215.0 58950.0 ;
      RECT  66510.0 60295.0 67215.0 58950.0 ;
      RECT  66510.0 60295.0 67215.0 61640.0 ;
      RECT  66510.0 62985.0 67215.0 61640.0 ;
      RECT  66510.0 62985.0 67215.0 64330.0 ;
      RECT  66510.0 65675.0 67215.0 64330.0 ;
      RECT  66510.0 65675.0 67215.0 67020.0 ;
      RECT  66510.0 68365.0 67215.0 67020.0 ;
      RECT  66510.0 68365.0 67215.0 69710.0 ;
      RECT  66510.0 71055.0 67215.0 69710.0 ;
      RECT  66510.0 71055.0 67215.0 72400.0 ;
      RECT  66510.0 73745.0 67215.0 72400.0 ;
      RECT  66510.0 73745.0 67215.0 75090.0 ;
      RECT  66510.0 76435.0 67215.0 75090.0 ;
      RECT  66510.0 76435.0 67215.0 77780.0 ;
      RECT  66510.0 79125.0 67215.0 77780.0 ;
      RECT  66510.0 79125.0 67215.0 80470.0 ;
      RECT  66510.0 81815.0 67215.0 80470.0 ;
      RECT  66510.0 81815.0 67215.0 83160.0 ;
      RECT  66510.0 84505.0 67215.0 83160.0 ;
      RECT  66510.0 84505.0 67215.0 85850.0 ;
      RECT  66510.0 87195.0 67215.0 85850.0 ;
      RECT  66510.0 87195.0 67215.0 88540.0 ;
      RECT  66510.0 89885.0 67215.0 88540.0 ;
      RECT  66510.0 89885.0 67215.0 91230.0 ;
      RECT  66510.0 92575.0 67215.0 91230.0 ;
      RECT  66510.0 92575.0 67215.0 93920.0 ;
      RECT  66510.0 95265.0 67215.0 93920.0 ;
      RECT  66510.0 95265.0 67215.0 96610.0 ;
      RECT  66510.0 97955.0 67215.0 96610.0 ;
      RECT  66510.0 97955.0 67215.0 99300.0 ;
      RECT  66510.0 100645.0 67215.0 99300.0 ;
      RECT  66510.0 100645.0 67215.0 101990.0 ;
      RECT  66510.0 103335.0 67215.0 101990.0 ;
      RECT  66510.0 103335.0 67215.0 104680.0 ;
      RECT  66510.0 106025.0 67215.0 104680.0 ;
      RECT  66510.0 106025.0 67215.0 107370.0 ;
      RECT  66510.0 108715.0 67215.0 107370.0 ;
      RECT  66510.0 108715.0 67215.0 110060.0 ;
      RECT  66510.0 111405.0 67215.0 110060.0 ;
      RECT  66510.0 111405.0 67215.0 112750.0 ;
      RECT  66510.0 114095.0 67215.0 112750.0 ;
      RECT  67215.0 28015.0 67920.0 29360.0 ;
      RECT  67215.0 30705.0 67920.0 29360.0 ;
      RECT  67215.0 30705.0 67920.0 32050.0 ;
      RECT  67215.0 33395.0 67920.0 32050.0 ;
      RECT  67215.0 33395.0 67920.0 34740.0 ;
      RECT  67215.0 36085.0 67920.0 34740.0 ;
      RECT  67215.0 36085.0 67920.0 37430.0 ;
      RECT  67215.0 38775.0 67920.0 37430.0 ;
      RECT  67215.0 38775.0 67920.0 40120.0 ;
      RECT  67215.0 41465.0 67920.0 40120.0 ;
      RECT  67215.0 41465.0 67920.0 42810.0 ;
      RECT  67215.0 44155.0 67920.0 42810.0 ;
      RECT  67215.0 44155.0 67920.0 45500.0 ;
      RECT  67215.0 46845.0 67920.0 45500.0 ;
      RECT  67215.0 46845.0 67920.0 48190.0 ;
      RECT  67215.0 49535.0 67920.0 48190.0 ;
      RECT  67215.0 49535.0 67920.0 50880.0 ;
      RECT  67215.0 52225.0 67920.0 50880.0 ;
      RECT  67215.0 52225.0 67920.0 53570.0 ;
      RECT  67215.0 54915.0 67920.0 53570.0 ;
      RECT  67215.0 54915.0 67920.0 56260.0 ;
      RECT  67215.0 57605.0 67920.0 56260.0 ;
      RECT  67215.0 57605.0 67920.0 58950.0 ;
      RECT  67215.0 60295.0 67920.0 58950.0 ;
      RECT  67215.0 60295.0 67920.0 61640.0 ;
      RECT  67215.0 62985.0 67920.0 61640.0 ;
      RECT  67215.0 62985.0 67920.0 64330.0 ;
      RECT  67215.0 65675.0 67920.0 64330.0 ;
      RECT  67215.0 65675.0 67920.0 67020.0 ;
      RECT  67215.0 68365.0 67920.0 67020.0 ;
      RECT  67215.0 68365.0 67920.0 69710.0 ;
      RECT  67215.0 71055.0 67920.0 69710.0 ;
      RECT  67215.0 71055.0 67920.0 72400.0 ;
      RECT  67215.0 73745.0 67920.0 72400.0 ;
      RECT  67215.0 73745.0 67920.0 75090.0 ;
      RECT  67215.0 76435.0 67920.0 75090.0 ;
      RECT  67215.0 76435.0 67920.0 77780.0 ;
      RECT  67215.0 79125.0 67920.0 77780.0 ;
      RECT  67215.0 79125.0 67920.0 80470.0 ;
      RECT  67215.0 81815.0 67920.0 80470.0 ;
      RECT  67215.0 81815.0 67920.0 83160.0 ;
      RECT  67215.0 84505.0 67920.0 83160.0 ;
      RECT  67215.0 84505.0 67920.0 85850.0 ;
      RECT  67215.0 87195.0 67920.0 85850.0 ;
      RECT  67215.0 87195.0 67920.0 88540.0 ;
      RECT  67215.0 89885.0 67920.0 88540.0 ;
      RECT  67215.0 89885.0 67920.0 91230.0 ;
      RECT  67215.0 92575.0 67920.0 91230.0 ;
      RECT  67215.0 92575.0 67920.0 93920.0 ;
      RECT  67215.0 95265.0 67920.0 93920.0 ;
      RECT  67215.0 95265.0 67920.0 96610.0 ;
      RECT  67215.0 97955.0 67920.0 96610.0 ;
      RECT  67215.0 97955.0 67920.0 99300.0 ;
      RECT  67215.0 100645.0 67920.0 99300.0 ;
      RECT  67215.0 100645.0 67920.0 101990.0 ;
      RECT  67215.0 103335.0 67920.0 101990.0 ;
      RECT  67215.0 103335.0 67920.0 104680.0 ;
      RECT  67215.0 106025.0 67920.0 104680.0 ;
      RECT  67215.0 106025.0 67920.0 107370.0 ;
      RECT  67215.0 108715.0 67920.0 107370.0 ;
      RECT  67215.0 108715.0 67920.0 110060.0 ;
      RECT  67215.0 111405.0 67920.0 110060.0 ;
      RECT  67215.0 111405.0 67920.0 112750.0 ;
      RECT  67215.0 114095.0 67920.0 112750.0 ;
      RECT  67920.0 28015.0 68625.0 29360.0 ;
      RECT  67920.0 30705.0 68625.0 29360.0 ;
      RECT  67920.0 30705.0 68625.0 32050.0 ;
      RECT  67920.0 33395.0 68625.0 32050.0 ;
      RECT  67920.0 33395.0 68625.0 34740.0 ;
      RECT  67920.0 36085.0 68625.0 34740.0 ;
      RECT  67920.0 36085.0 68625.0 37430.0 ;
      RECT  67920.0 38775.0 68625.0 37430.0 ;
      RECT  67920.0 38775.0 68625.0 40120.0 ;
      RECT  67920.0 41465.0 68625.0 40120.0 ;
      RECT  67920.0 41465.0 68625.0 42810.0 ;
      RECT  67920.0 44155.0 68625.0 42810.0 ;
      RECT  67920.0 44155.0 68625.0 45500.0 ;
      RECT  67920.0 46845.0 68625.0 45500.0 ;
      RECT  67920.0 46845.0 68625.0 48190.0 ;
      RECT  67920.0 49535.0 68625.0 48190.0 ;
      RECT  67920.0 49535.0 68625.0 50880.0 ;
      RECT  67920.0 52225.0 68625.0 50880.0 ;
      RECT  67920.0 52225.0 68625.0 53570.0 ;
      RECT  67920.0 54915.0 68625.0 53570.0 ;
      RECT  67920.0 54915.0 68625.0 56260.0 ;
      RECT  67920.0 57605.0 68625.0 56260.0 ;
      RECT  67920.0 57605.0 68625.0 58950.0 ;
      RECT  67920.0 60295.0 68625.0 58950.0 ;
      RECT  67920.0 60295.0 68625.0 61640.0 ;
      RECT  67920.0 62985.0 68625.0 61640.0 ;
      RECT  67920.0 62985.0 68625.0 64330.0 ;
      RECT  67920.0 65675.0 68625.0 64330.0 ;
      RECT  67920.0 65675.0 68625.0 67020.0 ;
      RECT  67920.0 68365.0 68625.0 67020.0 ;
      RECT  67920.0 68365.0 68625.0 69710.0 ;
      RECT  67920.0 71055.0 68625.0 69710.0 ;
      RECT  67920.0 71055.0 68625.0 72400.0 ;
      RECT  67920.0 73745.0 68625.0 72400.0 ;
      RECT  67920.0 73745.0 68625.0 75090.0 ;
      RECT  67920.0 76435.0 68625.0 75090.0 ;
      RECT  67920.0 76435.0 68625.0 77780.0 ;
      RECT  67920.0 79125.0 68625.0 77780.0 ;
      RECT  67920.0 79125.0 68625.0 80470.0 ;
      RECT  67920.0 81815.0 68625.0 80470.0 ;
      RECT  67920.0 81815.0 68625.0 83160.0 ;
      RECT  67920.0 84505.0 68625.0 83160.0 ;
      RECT  67920.0 84505.0 68625.0 85850.0 ;
      RECT  67920.0 87195.0 68625.0 85850.0 ;
      RECT  67920.0 87195.0 68625.0 88540.0 ;
      RECT  67920.0 89885.0 68625.0 88540.0 ;
      RECT  67920.0 89885.0 68625.0 91230.0 ;
      RECT  67920.0 92575.0 68625.0 91230.0 ;
      RECT  67920.0 92575.0 68625.0 93920.0 ;
      RECT  67920.0 95265.0 68625.0 93920.0 ;
      RECT  67920.0 95265.0 68625.0 96610.0 ;
      RECT  67920.0 97955.0 68625.0 96610.0 ;
      RECT  67920.0 97955.0 68625.0 99300.0 ;
      RECT  67920.0 100645.0 68625.0 99300.0 ;
      RECT  67920.0 100645.0 68625.0 101990.0 ;
      RECT  67920.0 103335.0 68625.0 101990.0 ;
      RECT  67920.0 103335.0 68625.0 104680.0 ;
      RECT  67920.0 106025.0 68625.0 104680.0 ;
      RECT  67920.0 106025.0 68625.0 107370.0 ;
      RECT  67920.0 108715.0 68625.0 107370.0 ;
      RECT  67920.0 108715.0 68625.0 110060.0 ;
      RECT  67920.0 111405.0 68625.0 110060.0 ;
      RECT  67920.0 111405.0 68625.0 112750.0 ;
      RECT  67920.0 114095.0 68625.0 112750.0 ;
      RECT  68625.0 28015.0 69330.0 29360.0 ;
      RECT  68625.0 30705.0 69330.0 29360.0 ;
      RECT  68625.0 30705.0 69330.0 32050.0 ;
      RECT  68625.0 33395.0 69330.0 32050.0 ;
      RECT  68625.0 33395.0 69330.0 34740.0 ;
      RECT  68625.0 36085.0 69330.0 34740.0 ;
      RECT  68625.0 36085.0 69330.0 37430.0 ;
      RECT  68625.0 38775.0 69330.0 37430.0 ;
      RECT  68625.0 38775.0 69330.0 40120.0 ;
      RECT  68625.0 41465.0 69330.0 40120.0 ;
      RECT  68625.0 41465.0 69330.0 42810.0 ;
      RECT  68625.0 44155.0 69330.0 42810.0 ;
      RECT  68625.0 44155.0 69330.0 45500.0 ;
      RECT  68625.0 46845.0 69330.0 45500.0 ;
      RECT  68625.0 46845.0 69330.0 48190.0 ;
      RECT  68625.0 49535.0 69330.0 48190.0 ;
      RECT  68625.0 49535.0 69330.0 50880.0 ;
      RECT  68625.0 52225.0 69330.0 50880.0 ;
      RECT  68625.0 52225.0 69330.0 53570.0 ;
      RECT  68625.0 54915.0 69330.0 53570.0 ;
      RECT  68625.0 54915.0 69330.0 56260.0 ;
      RECT  68625.0 57605.0 69330.0 56260.0 ;
      RECT  68625.0 57605.0 69330.0 58950.0 ;
      RECT  68625.0 60295.0 69330.0 58950.0 ;
      RECT  68625.0 60295.0 69330.0 61640.0 ;
      RECT  68625.0 62985.0 69330.0 61640.0 ;
      RECT  68625.0 62985.0 69330.0 64330.0 ;
      RECT  68625.0 65675.0 69330.0 64330.0 ;
      RECT  68625.0 65675.0 69330.0 67020.0 ;
      RECT  68625.0 68365.0 69330.0 67020.0 ;
      RECT  68625.0 68365.0 69330.0 69710.0 ;
      RECT  68625.0 71055.0 69330.0 69710.0 ;
      RECT  68625.0 71055.0 69330.0 72400.0 ;
      RECT  68625.0 73745.0 69330.0 72400.0 ;
      RECT  68625.0 73745.0 69330.0 75090.0 ;
      RECT  68625.0 76435.0 69330.0 75090.0 ;
      RECT  68625.0 76435.0 69330.0 77780.0 ;
      RECT  68625.0 79125.0 69330.0 77780.0 ;
      RECT  68625.0 79125.0 69330.0 80470.0 ;
      RECT  68625.0 81815.0 69330.0 80470.0 ;
      RECT  68625.0 81815.0 69330.0 83160.0 ;
      RECT  68625.0 84505.0 69330.0 83160.0 ;
      RECT  68625.0 84505.0 69330.0 85850.0 ;
      RECT  68625.0 87195.0 69330.0 85850.0 ;
      RECT  68625.0 87195.0 69330.0 88540.0 ;
      RECT  68625.0 89885.0 69330.0 88540.0 ;
      RECT  68625.0 89885.0 69330.0 91230.0 ;
      RECT  68625.0 92575.0 69330.0 91230.0 ;
      RECT  68625.0 92575.0 69330.0 93920.0 ;
      RECT  68625.0 95265.0 69330.0 93920.0 ;
      RECT  68625.0 95265.0 69330.0 96610.0 ;
      RECT  68625.0 97955.0 69330.0 96610.0 ;
      RECT  68625.0 97955.0 69330.0 99300.0 ;
      RECT  68625.0 100645.0 69330.0 99300.0 ;
      RECT  68625.0 100645.0 69330.0 101990.0 ;
      RECT  68625.0 103335.0 69330.0 101990.0 ;
      RECT  68625.0 103335.0 69330.0 104680.0 ;
      RECT  68625.0 106025.0 69330.0 104680.0 ;
      RECT  68625.0 106025.0 69330.0 107370.0 ;
      RECT  68625.0 108715.0 69330.0 107370.0 ;
      RECT  68625.0 108715.0 69330.0 110060.0 ;
      RECT  68625.0 111405.0 69330.0 110060.0 ;
      RECT  68625.0 111405.0 69330.0 112750.0 ;
      RECT  68625.0 114095.0 69330.0 112750.0 ;
      RECT  69330.0 28015.0 70035.0 29360.0 ;
      RECT  69330.0 30705.0 70035.0 29360.0 ;
      RECT  69330.0 30705.0 70035.0 32050.0 ;
      RECT  69330.0 33395.0 70035.0 32050.0 ;
      RECT  69330.0 33395.0 70035.0 34740.0 ;
      RECT  69330.0 36085.0 70035.0 34740.0 ;
      RECT  69330.0 36085.0 70035.0 37430.0 ;
      RECT  69330.0 38775.0 70035.0 37430.0 ;
      RECT  69330.0 38775.0 70035.0 40120.0 ;
      RECT  69330.0 41465.0 70035.0 40120.0 ;
      RECT  69330.0 41465.0 70035.0 42810.0 ;
      RECT  69330.0 44155.0 70035.0 42810.0 ;
      RECT  69330.0 44155.0 70035.0 45500.0 ;
      RECT  69330.0 46845.0 70035.0 45500.0 ;
      RECT  69330.0 46845.0 70035.0 48190.0 ;
      RECT  69330.0 49535.0 70035.0 48190.0 ;
      RECT  69330.0 49535.0 70035.0 50880.0 ;
      RECT  69330.0 52225.0 70035.0 50880.0 ;
      RECT  69330.0 52225.0 70035.0 53570.0 ;
      RECT  69330.0 54915.0 70035.0 53570.0 ;
      RECT  69330.0 54915.0 70035.0 56260.0 ;
      RECT  69330.0 57605.0 70035.0 56260.0 ;
      RECT  69330.0 57605.0 70035.0 58950.0 ;
      RECT  69330.0 60295.0 70035.0 58950.0 ;
      RECT  69330.0 60295.0 70035.0 61640.0 ;
      RECT  69330.0 62985.0 70035.0 61640.0 ;
      RECT  69330.0 62985.0 70035.0 64330.0 ;
      RECT  69330.0 65675.0 70035.0 64330.0 ;
      RECT  69330.0 65675.0 70035.0 67020.0 ;
      RECT  69330.0 68365.0 70035.0 67020.0 ;
      RECT  69330.0 68365.0 70035.0 69710.0 ;
      RECT  69330.0 71055.0 70035.0 69710.0 ;
      RECT  69330.0 71055.0 70035.0 72400.0 ;
      RECT  69330.0 73745.0 70035.0 72400.0 ;
      RECT  69330.0 73745.0 70035.0 75090.0 ;
      RECT  69330.0 76435.0 70035.0 75090.0 ;
      RECT  69330.0 76435.0 70035.0 77780.0 ;
      RECT  69330.0 79125.0 70035.0 77780.0 ;
      RECT  69330.0 79125.0 70035.0 80470.0 ;
      RECT  69330.0 81815.0 70035.0 80470.0 ;
      RECT  69330.0 81815.0 70035.0 83160.0 ;
      RECT  69330.0 84505.0 70035.0 83160.0 ;
      RECT  69330.0 84505.0 70035.0 85850.0 ;
      RECT  69330.0 87195.0 70035.0 85850.0 ;
      RECT  69330.0 87195.0 70035.0 88540.0 ;
      RECT  69330.0 89885.0 70035.0 88540.0 ;
      RECT  69330.0 89885.0 70035.0 91230.0 ;
      RECT  69330.0 92575.0 70035.0 91230.0 ;
      RECT  69330.0 92575.0 70035.0 93920.0 ;
      RECT  69330.0 95265.0 70035.0 93920.0 ;
      RECT  69330.0 95265.0 70035.0 96610.0 ;
      RECT  69330.0 97955.0 70035.0 96610.0 ;
      RECT  69330.0 97955.0 70035.0 99300.0 ;
      RECT  69330.0 100645.0 70035.0 99300.0 ;
      RECT  69330.0 100645.0 70035.0 101990.0 ;
      RECT  69330.0 103335.0 70035.0 101990.0 ;
      RECT  69330.0 103335.0 70035.0 104680.0 ;
      RECT  69330.0 106025.0 70035.0 104680.0 ;
      RECT  69330.0 106025.0 70035.0 107370.0 ;
      RECT  69330.0 108715.0 70035.0 107370.0 ;
      RECT  69330.0 108715.0 70035.0 110060.0 ;
      RECT  69330.0 111405.0 70035.0 110060.0 ;
      RECT  69330.0 111405.0 70035.0 112750.0 ;
      RECT  69330.0 114095.0 70035.0 112750.0 ;
      RECT  70035.0 28015.0 70740.0 29360.0 ;
      RECT  70035.0 30705.0 70740.0 29360.0 ;
      RECT  70035.0 30705.0 70740.0 32050.0 ;
      RECT  70035.0 33395.0 70740.0 32050.0 ;
      RECT  70035.0 33395.0 70740.0 34740.0 ;
      RECT  70035.0 36085.0 70740.0 34740.0 ;
      RECT  70035.0 36085.0 70740.0 37430.0 ;
      RECT  70035.0 38775.0 70740.0 37430.0 ;
      RECT  70035.0 38775.0 70740.0 40120.0 ;
      RECT  70035.0 41465.0 70740.0 40120.0 ;
      RECT  70035.0 41465.0 70740.0 42810.0 ;
      RECT  70035.0 44155.0 70740.0 42810.0 ;
      RECT  70035.0 44155.0 70740.0 45500.0 ;
      RECT  70035.0 46845.0 70740.0 45500.0 ;
      RECT  70035.0 46845.0 70740.0 48190.0 ;
      RECT  70035.0 49535.0 70740.0 48190.0 ;
      RECT  70035.0 49535.0 70740.0 50880.0 ;
      RECT  70035.0 52225.0 70740.0 50880.0 ;
      RECT  70035.0 52225.0 70740.0 53570.0 ;
      RECT  70035.0 54915.0 70740.0 53570.0 ;
      RECT  70035.0 54915.0 70740.0 56260.0 ;
      RECT  70035.0 57605.0 70740.0 56260.0 ;
      RECT  70035.0 57605.0 70740.0 58950.0 ;
      RECT  70035.0 60295.0 70740.0 58950.0 ;
      RECT  70035.0 60295.0 70740.0 61640.0 ;
      RECT  70035.0 62985.0 70740.0 61640.0 ;
      RECT  70035.0 62985.0 70740.0 64330.0 ;
      RECT  70035.0 65675.0 70740.0 64330.0 ;
      RECT  70035.0 65675.0 70740.0 67020.0 ;
      RECT  70035.0 68365.0 70740.0 67020.0 ;
      RECT  70035.0 68365.0 70740.0 69710.0 ;
      RECT  70035.0 71055.0 70740.0 69710.0 ;
      RECT  70035.0 71055.0 70740.0 72400.0 ;
      RECT  70035.0 73745.0 70740.0 72400.0 ;
      RECT  70035.0 73745.0 70740.0 75090.0 ;
      RECT  70035.0 76435.0 70740.0 75090.0 ;
      RECT  70035.0 76435.0 70740.0 77780.0 ;
      RECT  70035.0 79125.0 70740.0 77780.0 ;
      RECT  70035.0 79125.0 70740.0 80470.0 ;
      RECT  70035.0 81815.0 70740.0 80470.0 ;
      RECT  70035.0 81815.0 70740.0 83160.0 ;
      RECT  70035.0 84505.0 70740.0 83160.0 ;
      RECT  70035.0 84505.0 70740.0 85850.0 ;
      RECT  70035.0 87195.0 70740.0 85850.0 ;
      RECT  70035.0 87195.0 70740.0 88540.0 ;
      RECT  70035.0 89885.0 70740.0 88540.0 ;
      RECT  70035.0 89885.0 70740.0 91230.0 ;
      RECT  70035.0 92575.0 70740.0 91230.0 ;
      RECT  70035.0 92575.0 70740.0 93920.0 ;
      RECT  70035.0 95265.0 70740.0 93920.0 ;
      RECT  70035.0 95265.0 70740.0 96610.0 ;
      RECT  70035.0 97955.0 70740.0 96610.0 ;
      RECT  70035.0 97955.0 70740.0 99300.0 ;
      RECT  70035.0 100645.0 70740.0 99300.0 ;
      RECT  70035.0 100645.0 70740.0 101990.0 ;
      RECT  70035.0 103335.0 70740.0 101990.0 ;
      RECT  70035.0 103335.0 70740.0 104680.0 ;
      RECT  70035.0 106025.0 70740.0 104680.0 ;
      RECT  70035.0 106025.0 70740.0 107370.0 ;
      RECT  70035.0 108715.0 70740.0 107370.0 ;
      RECT  70035.0 108715.0 70740.0 110060.0 ;
      RECT  70035.0 111405.0 70740.0 110060.0 ;
      RECT  70035.0 111405.0 70740.0 112750.0 ;
      RECT  70035.0 114095.0 70740.0 112750.0 ;
      RECT  70740.0 28015.0 71445.0 29360.0 ;
      RECT  70740.0 30705.0 71445.0 29360.0 ;
      RECT  70740.0 30705.0 71445.0 32050.0 ;
      RECT  70740.0 33395.0 71445.0 32050.0 ;
      RECT  70740.0 33395.0 71445.0 34740.0 ;
      RECT  70740.0 36085.0 71445.0 34740.0 ;
      RECT  70740.0 36085.0 71445.0 37430.0 ;
      RECT  70740.0 38775.0 71445.0 37430.0 ;
      RECT  70740.0 38775.0 71445.0 40120.0 ;
      RECT  70740.0 41465.0 71445.0 40120.0 ;
      RECT  70740.0 41465.0 71445.0 42810.0 ;
      RECT  70740.0 44155.0 71445.0 42810.0 ;
      RECT  70740.0 44155.0 71445.0 45500.0 ;
      RECT  70740.0 46845.0 71445.0 45500.0 ;
      RECT  70740.0 46845.0 71445.0 48190.0 ;
      RECT  70740.0 49535.0 71445.0 48190.0 ;
      RECT  70740.0 49535.0 71445.0 50880.0 ;
      RECT  70740.0 52225.0 71445.0 50880.0 ;
      RECT  70740.0 52225.0 71445.0 53570.0 ;
      RECT  70740.0 54915.0 71445.0 53570.0 ;
      RECT  70740.0 54915.0 71445.0 56260.0 ;
      RECT  70740.0 57605.0 71445.0 56260.0 ;
      RECT  70740.0 57605.0 71445.0 58950.0 ;
      RECT  70740.0 60295.0 71445.0 58950.0 ;
      RECT  70740.0 60295.0 71445.0 61640.0 ;
      RECT  70740.0 62985.0 71445.0 61640.0 ;
      RECT  70740.0 62985.0 71445.0 64330.0 ;
      RECT  70740.0 65675.0 71445.0 64330.0 ;
      RECT  70740.0 65675.0 71445.0 67020.0 ;
      RECT  70740.0 68365.0 71445.0 67020.0 ;
      RECT  70740.0 68365.0 71445.0 69710.0 ;
      RECT  70740.0 71055.0 71445.0 69710.0 ;
      RECT  70740.0 71055.0 71445.0 72400.0 ;
      RECT  70740.0 73745.0 71445.0 72400.0 ;
      RECT  70740.0 73745.0 71445.0 75090.0 ;
      RECT  70740.0 76435.0 71445.0 75090.0 ;
      RECT  70740.0 76435.0 71445.0 77780.0 ;
      RECT  70740.0 79125.0 71445.0 77780.0 ;
      RECT  70740.0 79125.0 71445.0 80470.0 ;
      RECT  70740.0 81815.0 71445.0 80470.0 ;
      RECT  70740.0 81815.0 71445.0 83160.0 ;
      RECT  70740.0 84505.0 71445.0 83160.0 ;
      RECT  70740.0 84505.0 71445.0 85850.0 ;
      RECT  70740.0 87195.0 71445.0 85850.0 ;
      RECT  70740.0 87195.0 71445.0 88540.0 ;
      RECT  70740.0 89885.0 71445.0 88540.0 ;
      RECT  70740.0 89885.0 71445.0 91230.0 ;
      RECT  70740.0 92575.0 71445.0 91230.0 ;
      RECT  70740.0 92575.0 71445.0 93920.0 ;
      RECT  70740.0 95265.0 71445.0 93920.0 ;
      RECT  70740.0 95265.0 71445.0 96610.0 ;
      RECT  70740.0 97955.0 71445.0 96610.0 ;
      RECT  70740.0 97955.0 71445.0 99300.0 ;
      RECT  70740.0 100645.0 71445.0 99300.0 ;
      RECT  70740.0 100645.0 71445.0 101990.0 ;
      RECT  70740.0 103335.0 71445.0 101990.0 ;
      RECT  70740.0 103335.0 71445.0 104680.0 ;
      RECT  70740.0 106025.0 71445.0 104680.0 ;
      RECT  70740.0 106025.0 71445.0 107370.0 ;
      RECT  70740.0 108715.0 71445.0 107370.0 ;
      RECT  70740.0 108715.0 71445.0 110060.0 ;
      RECT  70740.0 111405.0 71445.0 110060.0 ;
      RECT  70740.0 111405.0 71445.0 112750.0 ;
      RECT  70740.0 114095.0 71445.0 112750.0 ;
      RECT  71445.0 28015.0 72150.0 29360.0 ;
      RECT  71445.0 30705.0 72150.0 29360.0 ;
      RECT  71445.0 30705.0 72150.0 32050.0 ;
      RECT  71445.0 33395.0 72150.0 32050.0 ;
      RECT  71445.0 33395.0 72150.0 34740.0 ;
      RECT  71445.0 36085.0 72150.0 34740.0 ;
      RECT  71445.0 36085.0 72150.0 37430.0 ;
      RECT  71445.0 38775.0 72150.0 37430.0 ;
      RECT  71445.0 38775.0 72150.0 40120.0 ;
      RECT  71445.0 41465.0 72150.0 40120.0 ;
      RECT  71445.0 41465.0 72150.0 42810.0 ;
      RECT  71445.0 44155.0 72150.0 42810.0 ;
      RECT  71445.0 44155.0 72150.0 45500.0 ;
      RECT  71445.0 46845.0 72150.0 45500.0 ;
      RECT  71445.0 46845.0 72150.0 48190.0 ;
      RECT  71445.0 49535.0 72150.0 48190.0 ;
      RECT  71445.0 49535.0 72150.0 50880.0 ;
      RECT  71445.0 52225.0 72150.0 50880.0 ;
      RECT  71445.0 52225.0 72150.0 53570.0 ;
      RECT  71445.0 54915.0 72150.0 53570.0 ;
      RECT  71445.0 54915.0 72150.0 56260.0 ;
      RECT  71445.0 57605.0 72150.0 56260.0 ;
      RECT  71445.0 57605.0 72150.0 58950.0 ;
      RECT  71445.0 60295.0 72150.0 58950.0 ;
      RECT  71445.0 60295.0 72150.0 61640.0 ;
      RECT  71445.0 62985.0 72150.0 61640.0 ;
      RECT  71445.0 62985.0 72150.0 64330.0 ;
      RECT  71445.0 65675.0 72150.0 64330.0 ;
      RECT  71445.0 65675.0 72150.0 67020.0 ;
      RECT  71445.0 68365.0 72150.0 67020.0 ;
      RECT  71445.0 68365.0 72150.0 69710.0 ;
      RECT  71445.0 71055.0 72150.0 69710.0 ;
      RECT  71445.0 71055.0 72150.0 72400.0 ;
      RECT  71445.0 73745.0 72150.0 72400.0 ;
      RECT  71445.0 73745.0 72150.0 75090.0 ;
      RECT  71445.0 76435.0 72150.0 75090.0 ;
      RECT  71445.0 76435.0 72150.0 77780.0 ;
      RECT  71445.0 79125.0 72150.0 77780.0 ;
      RECT  71445.0 79125.0 72150.0 80470.0 ;
      RECT  71445.0 81815.0 72150.0 80470.0 ;
      RECT  71445.0 81815.0 72150.0 83160.0 ;
      RECT  71445.0 84505.0 72150.0 83160.0 ;
      RECT  71445.0 84505.0 72150.0 85850.0 ;
      RECT  71445.0 87195.0 72150.0 85850.0 ;
      RECT  71445.0 87195.0 72150.0 88540.0 ;
      RECT  71445.0 89885.0 72150.0 88540.0 ;
      RECT  71445.0 89885.0 72150.0 91230.0 ;
      RECT  71445.0 92575.0 72150.0 91230.0 ;
      RECT  71445.0 92575.0 72150.0 93920.0 ;
      RECT  71445.0 95265.0 72150.0 93920.0 ;
      RECT  71445.0 95265.0 72150.0 96610.0 ;
      RECT  71445.0 97955.0 72150.0 96610.0 ;
      RECT  71445.0 97955.0 72150.0 99300.0 ;
      RECT  71445.0 100645.0 72150.0 99300.0 ;
      RECT  71445.0 100645.0 72150.0 101990.0 ;
      RECT  71445.0 103335.0 72150.0 101990.0 ;
      RECT  71445.0 103335.0 72150.0 104680.0 ;
      RECT  71445.0 106025.0 72150.0 104680.0 ;
      RECT  71445.0 106025.0 72150.0 107370.0 ;
      RECT  71445.0 108715.0 72150.0 107370.0 ;
      RECT  71445.0 108715.0 72150.0 110060.0 ;
      RECT  71445.0 111405.0 72150.0 110060.0 ;
      RECT  71445.0 111405.0 72150.0 112750.0 ;
      RECT  71445.0 114095.0 72150.0 112750.0 ;
      RECT  72150.0 28015.0 72855.0 29360.0 ;
      RECT  72150.0 30705.0 72855.0 29360.0 ;
      RECT  72150.0 30705.0 72855.0 32050.0 ;
      RECT  72150.0 33395.0 72855.0 32050.0 ;
      RECT  72150.0 33395.0 72855.0 34740.0 ;
      RECT  72150.0 36085.0 72855.0 34740.0 ;
      RECT  72150.0 36085.0 72855.0 37430.0 ;
      RECT  72150.0 38775.0 72855.0 37430.0 ;
      RECT  72150.0 38775.0 72855.0 40120.0 ;
      RECT  72150.0 41465.0 72855.0 40120.0 ;
      RECT  72150.0 41465.0 72855.0 42810.0 ;
      RECT  72150.0 44155.0 72855.0 42810.0 ;
      RECT  72150.0 44155.0 72855.0 45500.0 ;
      RECT  72150.0 46845.0 72855.0 45500.0 ;
      RECT  72150.0 46845.0 72855.0 48190.0 ;
      RECT  72150.0 49535.0 72855.0 48190.0 ;
      RECT  72150.0 49535.0 72855.0 50880.0 ;
      RECT  72150.0 52225.0 72855.0 50880.0 ;
      RECT  72150.0 52225.0 72855.0 53570.0 ;
      RECT  72150.0 54915.0 72855.0 53570.0 ;
      RECT  72150.0 54915.0 72855.0 56260.0 ;
      RECT  72150.0 57605.0 72855.0 56260.0 ;
      RECT  72150.0 57605.0 72855.0 58950.0 ;
      RECT  72150.0 60295.0 72855.0 58950.0 ;
      RECT  72150.0 60295.0 72855.0 61640.0 ;
      RECT  72150.0 62985.0 72855.0 61640.0 ;
      RECT  72150.0 62985.0 72855.0 64330.0 ;
      RECT  72150.0 65675.0 72855.0 64330.0 ;
      RECT  72150.0 65675.0 72855.0 67020.0 ;
      RECT  72150.0 68365.0 72855.0 67020.0 ;
      RECT  72150.0 68365.0 72855.0 69710.0 ;
      RECT  72150.0 71055.0 72855.0 69710.0 ;
      RECT  72150.0 71055.0 72855.0 72400.0 ;
      RECT  72150.0 73745.0 72855.0 72400.0 ;
      RECT  72150.0 73745.0 72855.0 75090.0 ;
      RECT  72150.0 76435.0 72855.0 75090.0 ;
      RECT  72150.0 76435.0 72855.0 77780.0 ;
      RECT  72150.0 79125.0 72855.0 77780.0 ;
      RECT  72150.0 79125.0 72855.0 80470.0 ;
      RECT  72150.0 81815.0 72855.0 80470.0 ;
      RECT  72150.0 81815.0 72855.0 83160.0 ;
      RECT  72150.0 84505.0 72855.0 83160.0 ;
      RECT  72150.0 84505.0 72855.0 85850.0 ;
      RECT  72150.0 87195.0 72855.0 85850.0 ;
      RECT  72150.0 87195.0 72855.0 88540.0 ;
      RECT  72150.0 89885.0 72855.0 88540.0 ;
      RECT  72150.0 89885.0 72855.0 91230.0 ;
      RECT  72150.0 92575.0 72855.0 91230.0 ;
      RECT  72150.0 92575.0 72855.0 93920.0 ;
      RECT  72150.0 95265.0 72855.0 93920.0 ;
      RECT  72150.0 95265.0 72855.0 96610.0 ;
      RECT  72150.0 97955.0 72855.0 96610.0 ;
      RECT  72150.0 97955.0 72855.0 99300.0 ;
      RECT  72150.0 100645.0 72855.0 99300.0 ;
      RECT  72150.0 100645.0 72855.0 101990.0 ;
      RECT  72150.0 103335.0 72855.0 101990.0 ;
      RECT  72150.0 103335.0 72855.0 104680.0 ;
      RECT  72150.0 106025.0 72855.0 104680.0 ;
      RECT  72150.0 106025.0 72855.0 107370.0 ;
      RECT  72150.0 108715.0 72855.0 107370.0 ;
      RECT  72150.0 108715.0 72855.0 110060.0 ;
      RECT  72150.0 111405.0 72855.0 110060.0 ;
      RECT  72150.0 111405.0 72855.0 112750.0 ;
      RECT  72150.0 114095.0 72855.0 112750.0 ;
      RECT  72855.0 28015.0 73560.0 29360.0 ;
      RECT  72855.0 30705.0 73560.0 29360.0 ;
      RECT  72855.0 30705.0 73560.0 32050.0 ;
      RECT  72855.0 33395.0 73560.0 32050.0 ;
      RECT  72855.0 33395.0 73560.0 34740.0 ;
      RECT  72855.0 36085.0 73560.0 34740.0 ;
      RECT  72855.0 36085.0 73560.0 37430.0 ;
      RECT  72855.0 38775.0 73560.0 37430.0 ;
      RECT  72855.0 38775.0 73560.0 40120.0 ;
      RECT  72855.0 41465.0 73560.0 40120.0 ;
      RECT  72855.0 41465.0 73560.0 42810.0 ;
      RECT  72855.0 44155.0 73560.0 42810.0 ;
      RECT  72855.0 44155.0 73560.0 45500.0 ;
      RECT  72855.0 46845.0 73560.0 45500.0 ;
      RECT  72855.0 46845.0 73560.0 48190.0 ;
      RECT  72855.0 49535.0 73560.0 48190.0 ;
      RECT  72855.0 49535.0 73560.0 50880.0 ;
      RECT  72855.0 52225.0 73560.0 50880.0 ;
      RECT  72855.0 52225.0 73560.0 53570.0 ;
      RECT  72855.0 54915.0 73560.0 53570.0 ;
      RECT  72855.0 54915.0 73560.0 56260.0 ;
      RECT  72855.0 57605.0 73560.0 56260.0 ;
      RECT  72855.0 57605.0 73560.0 58950.0 ;
      RECT  72855.0 60295.0 73560.0 58950.0 ;
      RECT  72855.0 60295.0 73560.0 61640.0 ;
      RECT  72855.0 62985.0 73560.0 61640.0 ;
      RECT  72855.0 62985.0 73560.0 64330.0 ;
      RECT  72855.0 65675.0 73560.0 64330.0 ;
      RECT  72855.0 65675.0 73560.0 67020.0 ;
      RECT  72855.0 68365.0 73560.0 67020.0 ;
      RECT  72855.0 68365.0 73560.0 69710.0 ;
      RECT  72855.0 71055.0 73560.0 69710.0 ;
      RECT  72855.0 71055.0 73560.0 72400.0 ;
      RECT  72855.0 73745.0 73560.0 72400.0 ;
      RECT  72855.0 73745.0 73560.0 75090.0 ;
      RECT  72855.0 76435.0 73560.0 75090.0 ;
      RECT  72855.0 76435.0 73560.0 77780.0 ;
      RECT  72855.0 79125.0 73560.0 77780.0 ;
      RECT  72855.0 79125.0 73560.0 80470.0 ;
      RECT  72855.0 81815.0 73560.0 80470.0 ;
      RECT  72855.0 81815.0 73560.0 83160.0 ;
      RECT  72855.0 84505.0 73560.0 83160.0 ;
      RECT  72855.0 84505.0 73560.0 85850.0 ;
      RECT  72855.0 87195.0 73560.0 85850.0 ;
      RECT  72855.0 87195.0 73560.0 88540.0 ;
      RECT  72855.0 89885.0 73560.0 88540.0 ;
      RECT  72855.0 89885.0 73560.0 91230.0 ;
      RECT  72855.0 92575.0 73560.0 91230.0 ;
      RECT  72855.0 92575.0 73560.0 93920.0 ;
      RECT  72855.0 95265.0 73560.0 93920.0 ;
      RECT  72855.0 95265.0 73560.0 96610.0 ;
      RECT  72855.0 97955.0 73560.0 96610.0 ;
      RECT  72855.0 97955.0 73560.0 99300.0 ;
      RECT  72855.0 100645.0 73560.0 99300.0 ;
      RECT  72855.0 100645.0 73560.0 101990.0 ;
      RECT  72855.0 103335.0 73560.0 101990.0 ;
      RECT  72855.0 103335.0 73560.0 104680.0 ;
      RECT  72855.0 106025.0 73560.0 104680.0 ;
      RECT  72855.0 106025.0 73560.0 107370.0 ;
      RECT  72855.0 108715.0 73560.0 107370.0 ;
      RECT  72855.0 108715.0 73560.0 110060.0 ;
      RECT  72855.0 111405.0 73560.0 110060.0 ;
      RECT  72855.0 111405.0 73560.0 112750.0 ;
      RECT  72855.0 114095.0 73560.0 112750.0 ;
      RECT  73560.0 28015.0 74265.0 29360.0 ;
      RECT  73560.0 30705.0 74265.0 29360.0 ;
      RECT  73560.0 30705.0 74265.0 32050.0 ;
      RECT  73560.0 33395.0 74265.0 32050.0 ;
      RECT  73560.0 33395.0 74265.0 34740.0 ;
      RECT  73560.0 36085.0 74265.0 34740.0 ;
      RECT  73560.0 36085.0 74265.0 37430.0 ;
      RECT  73560.0 38775.0 74265.0 37430.0 ;
      RECT  73560.0 38775.0 74265.0 40120.0 ;
      RECT  73560.0 41465.0 74265.0 40120.0 ;
      RECT  73560.0 41465.0 74265.0 42810.0 ;
      RECT  73560.0 44155.0 74265.0 42810.0 ;
      RECT  73560.0 44155.0 74265.0 45500.0 ;
      RECT  73560.0 46845.0 74265.0 45500.0 ;
      RECT  73560.0 46845.0 74265.0 48190.0 ;
      RECT  73560.0 49535.0 74265.0 48190.0 ;
      RECT  73560.0 49535.0 74265.0 50880.0 ;
      RECT  73560.0 52225.0 74265.0 50880.0 ;
      RECT  73560.0 52225.0 74265.0 53570.0 ;
      RECT  73560.0 54915.0 74265.0 53570.0 ;
      RECT  73560.0 54915.0 74265.0 56260.0 ;
      RECT  73560.0 57605.0 74265.0 56260.0 ;
      RECT  73560.0 57605.0 74265.0 58950.0 ;
      RECT  73560.0 60295.0 74265.0 58950.0 ;
      RECT  73560.0 60295.0 74265.0 61640.0 ;
      RECT  73560.0 62985.0 74265.0 61640.0 ;
      RECT  73560.0 62985.0 74265.0 64330.0 ;
      RECT  73560.0 65675.0 74265.0 64330.0 ;
      RECT  73560.0 65675.0 74265.0 67020.0 ;
      RECT  73560.0 68365.0 74265.0 67020.0 ;
      RECT  73560.0 68365.0 74265.0 69710.0 ;
      RECT  73560.0 71055.0 74265.0 69710.0 ;
      RECT  73560.0 71055.0 74265.0 72400.0 ;
      RECT  73560.0 73745.0 74265.0 72400.0 ;
      RECT  73560.0 73745.0 74265.0 75090.0 ;
      RECT  73560.0 76435.0 74265.0 75090.0 ;
      RECT  73560.0 76435.0 74265.0 77780.0 ;
      RECT  73560.0 79125.0 74265.0 77780.0 ;
      RECT  73560.0 79125.0 74265.0 80470.0 ;
      RECT  73560.0 81815.0 74265.0 80470.0 ;
      RECT  73560.0 81815.0 74265.0 83160.0 ;
      RECT  73560.0 84505.0 74265.0 83160.0 ;
      RECT  73560.0 84505.0 74265.0 85850.0 ;
      RECT  73560.0 87195.0 74265.0 85850.0 ;
      RECT  73560.0 87195.0 74265.0 88540.0 ;
      RECT  73560.0 89885.0 74265.0 88540.0 ;
      RECT  73560.0 89885.0 74265.0 91230.0 ;
      RECT  73560.0 92575.0 74265.0 91230.0 ;
      RECT  73560.0 92575.0 74265.0 93920.0 ;
      RECT  73560.0 95265.0 74265.0 93920.0 ;
      RECT  73560.0 95265.0 74265.0 96610.0 ;
      RECT  73560.0 97955.0 74265.0 96610.0 ;
      RECT  73560.0 97955.0 74265.0 99300.0 ;
      RECT  73560.0 100645.0 74265.0 99300.0 ;
      RECT  73560.0 100645.0 74265.0 101990.0 ;
      RECT  73560.0 103335.0 74265.0 101990.0 ;
      RECT  73560.0 103335.0 74265.0 104680.0 ;
      RECT  73560.0 106025.0 74265.0 104680.0 ;
      RECT  73560.0 106025.0 74265.0 107370.0 ;
      RECT  73560.0 108715.0 74265.0 107370.0 ;
      RECT  73560.0 108715.0 74265.0 110060.0 ;
      RECT  73560.0 111405.0 74265.0 110060.0 ;
      RECT  73560.0 111405.0 74265.0 112750.0 ;
      RECT  73560.0 114095.0 74265.0 112750.0 ;
      RECT  74265.0 28015.0 74970.0 29360.0 ;
      RECT  74265.0 30705.0 74970.0 29360.0 ;
      RECT  74265.0 30705.0 74970.0 32050.0 ;
      RECT  74265.0 33395.0 74970.0 32050.0 ;
      RECT  74265.0 33395.0 74970.0 34740.0 ;
      RECT  74265.0 36085.0 74970.0 34740.0 ;
      RECT  74265.0 36085.0 74970.0 37430.0 ;
      RECT  74265.0 38775.0 74970.0 37430.0 ;
      RECT  74265.0 38775.0 74970.0 40120.0 ;
      RECT  74265.0 41465.0 74970.0 40120.0 ;
      RECT  74265.0 41465.0 74970.0 42810.0 ;
      RECT  74265.0 44155.0 74970.0 42810.0 ;
      RECT  74265.0 44155.0 74970.0 45500.0 ;
      RECT  74265.0 46845.0 74970.0 45500.0 ;
      RECT  74265.0 46845.0 74970.0 48190.0 ;
      RECT  74265.0 49535.0 74970.0 48190.0 ;
      RECT  74265.0 49535.0 74970.0 50880.0 ;
      RECT  74265.0 52225.0 74970.0 50880.0 ;
      RECT  74265.0 52225.0 74970.0 53570.0 ;
      RECT  74265.0 54915.0 74970.0 53570.0 ;
      RECT  74265.0 54915.0 74970.0 56260.0 ;
      RECT  74265.0 57605.0 74970.0 56260.0 ;
      RECT  74265.0 57605.0 74970.0 58950.0 ;
      RECT  74265.0 60295.0 74970.0 58950.0 ;
      RECT  74265.0 60295.0 74970.0 61640.0 ;
      RECT  74265.0 62985.0 74970.0 61640.0 ;
      RECT  74265.0 62985.0 74970.0 64330.0 ;
      RECT  74265.0 65675.0 74970.0 64330.0 ;
      RECT  74265.0 65675.0 74970.0 67020.0 ;
      RECT  74265.0 68365.0 74970.0 67020.0 ;
      RECT  74265.0 68365.0 74970.0 69710.0 ;
      RECT  74265.0 71055.0 74970.0 69710.0 ;
      RECT  74265.0 71055.0 74970.0 72400.0 ;
      RECT  74265.0 73745.0 74970.0 72400.0 ;
      RECT  74265.0 73745.0 74970.0 75090.0 ;
      RECT  74265.0 76435.0 74970.0 75090.0 ;
      RECT  74265.0 76435.0 74970.0 77780.0 ;
      RECT  74265.0 79125.0 74970.0 77780.0 ;
      RECT  74265.0 79125.0 74970.0 80470.0 ;
      RECT  74265.0 81815.0 74970.0 80470.0 ;
      RECT  74265.0 81815.0 74970.0 83160.0 ;
      RECT  74265.0 84505.0 74970.0 83160.0 ;
      RECT  74265.0 84505.0 74970.0 85850.0 ;
      RECT  74265.0 87195.0 74970.0 85850.0 ;
      RECT  74265.0 87195.0 74970.0 88540.0 ;
      RECT  74265.0 89885.0 74970.0 88540.0 ;
      RECT  74265.0 89885.0 74970.0 91230.0 ;
      RECT  74265.0 92575.0 74970.0 91230.0 ;
      RECT  74265.0 92575.0 74970.0 93920.0 ;
      RECT  74265.0 95265.0 74970.0 93920.0 ;
      RECT  74265.0 95265.0 74970.0 96610.0 ;
      RECT  74265.0 97955.0 74970.0 96610.0 ;
      RECT  74265.0 97955.0 74970.0 99300.0 ;
      RECT  74265.0 100645.0 74970.0 99300.0 ;
      RECT  74265.0 100645.0 74970.0 101990.0 ;
      RECT  74265.0 103335.0 74970.0 101990.0 ;
      RECT  74265.0 103335.0 74970.0 104680.0 ;
      RECT  74265.0 106025.0 74970.0 104680.0 ;
      RECT  74265.0 106025.0 74970.0 107370.0 ;
      RECT  74265.0 108715.0 74970.0 107370.0 ;
      RECT  74265.0 108715.0 74970.0 110060.0 ;
      RECT  74265.0 111405.0 74970.0 110060.0 ;
      RECT  74265.0 111405.0 74970.0 112750.0 ;
      RECT  74265.0 114095.0 74970.0 112750.0 ;
      RECT  74970.0 28015.0 75675.0 29360.0 ;
      RECT  74970.0 30705.0 75675.0 29360.0 ;
      RECT  74970.0 30705.0 75675.0 32050.0 ;
      RECT  74970.0 33395.0 75675.0 32050.0 ;
      RECT  74970.0 33395.0 75675.0 34740.0 ;
      RECT  74970.0 36085.0 75675.0 34740.0 ;
      RECT  74970.0 36085.0 75675.0 37430.0 ;
      RECT  74970.0 38775.0 75675.0 37430.0 ;
      RECT  74970.0 38775.0 75675.0 40120.0 ;
      RECT  74970.0 41465.0 75675.0 40120.0 ;
      RECT  74970.0 41465.0 75675.0 42810.0 ;
      RECT  74970.0 44155.0 75675.0 42810.0 ;
      RECT  74970.0 44155.0 75675.0 45500.0 ;
      RECT  74970.0 46845.0 75675.0 45500.0 ;
      RECT  74970.0 46845.0 75675.0 48190.0 ;
      RECT  74970.0 49535.0 75675.0 48190.0 ;
      RECT  74970.0 49535.0 75675.0 50880.0 ;
      RECT  74970.0 52225.0 75675.0 50880.0 ;
      RECT  74970.0 52225.0 75675.0 53570.0 ;
      RECT  74970.0 54915.0 75675.0 53570.0 ;
      RECT  74970.0 54915.0 75675.0 56260.0 ;
      RECT  74970.0 57605.0 75675.0 56260.0 ;
      RECT  74970.0 57605.0 75675.0 58950.0 ;
      RECT  74970.0 60295.0 75675.0 58950.0 ;
      RECT  74970.0 60295.0 75675.0 61640.0 ;
      RECT  74970.0 62985.0 75675.0 61640.0 ;
      RECT  74970.0 62985.0 75675.0 64330.0 ;
      RECT  74970.0 65675.0 75675.0 64330.0 ;
      RECT  74970.0 65675.0 75675.0 67020.0 ;
      RECT  74970.0 68365.0 75675.0 67020.0 ;
      RECT  74970.0 68365.0 75675.0 69710.0 ;
      RECT  74970.0 71055.0 75675.0 69710.0 ;
      RECT  74970.0 71055.0 75675.0 72400.0 ;
      RECT  74970.0 73745.0 75675.0 72400.0 ;
      RECT  74970.0 73745.0 75675.0 75090.0 ;
      RECT  74970.0 76435.0 75675.0 75090.0 ;
      RECT  74970.0 76435.0 75675.0 77780.0 ;
      RECT  74970.0 79125.0 75675.0 77780.0 ;
      RECT  74970.0 79125.0 75675.0 80470.0 ;
      RECT  74970.0 81815.0 75675.0 80470.0 ;
      RECT  74970.0 81815.0 75675.0 83160.0 ;
      RECT  74970.0 84505.0 75675.0 83160.0 ;
      RECT  74970.0 84505.0 75675.0 85850.0 ;
      RECT  74970.0 87195.0 75675.0 85850.0 ;
      RECT  74970.0 87195.0 75675.0 88540.0 ;
      RECT  74970.0 89885.0 75675.0 88540.0 ;
      RECT  74970.0 89885.0 75675.0 91230.0 ;
      RECT  74970.0 92575.0 75675.0 91230.0 ;
      RECT  74970.0 92575.0 75675.0 93920.0 ;
      RECT  74970.0 95265.0 75675.0 93920.0 ;
      RECT  74970.0 95265.0 75675.0 96610.0 ;
      RECT  74970.0 97955.0 75675.0 96610.0 ;
      RECT  74970.0 97955.0 75675.0 99300.0 ;
      RECT  74970.0 100645.0 75675.0 99300.0 ;
      RECT  74970.0 100645.0 75675.0 101990.0 ;
      RECT  74970.0 103335.0 75675.0 101990.0 ;
      RECT  74970.0 103335.0 75675.0 104680.0 ;
      RECT  74970.0 106025.0 75675.0 104680.0 ;
      RECT  74970.0 106025.0 75675.0 107370.0 ;
      RECT  74970.0 108715.0 75675.0 107370.0 ;
      RECT  74970.0 108715.0 75675.0 110060.0 ;
      RECT  74970.0 111405.0 75675.0 110060.0 ;
      RECT  74970.0 111405.0 75675.0 112750.0 ;
      RECT  74970.0 114095.0 75675.0 112750.0 ;
      RECT  75675.0 28015.0 76380.0 29360.0 ;
      RECT  75675.0 30705.0 76380.0 29360.0 ;
      RECT  75675.0 30705.0 76380.0 32050.0 ;
      RECT  75675.0 33395.0 76380.0 32050.0 ;
      RECT  75675.0 33395.0 76380.0 34740.0 ;
      RECT  75675.0 36085.0 76380.0 34740.0 ;
      RECT  75675.0 36085.0 76380.0 37430.0 ;
      RECT  75675.0 38775.0 76380.0 37430.0 ;
      RECT  75675.0 38775.0 76380.0 40120.0 ;
      RECT  75675.0 41465.0 76380.0 40120.0 ;
      RECT  75675.0 41465.0 76380.0 42810.0 ;
      RECT  75675.0 44155.0 76380.0 42810.0 ;
      RECT  75675.0 44155.0 76380.0 45500.0 ;
      RECT  75675.0 46845.0 76380.0 45500.0 ;
      RECT  75675.0 46845.0 76380.0 48190.0 ;
      RECT  75675.0 49535.0 76380.0 48190.0 ;
      RECT  75675.0 49535.0 76380.0 50880.0 ;
      RECT  75675.0 52225.0 76380.0 50880.0 ;
      RECT  75675.0 52225.0 76380.0 53570.0 ;
      RECT  75675.0 54915.0 76380.0 53570.0 ;
      RECT  75675.0 54915.0 76380.0 56260.0 ;
      RECT  75675.0 57605.0 76380.0 56260.0 ;
      RECT  75675.0 57605.0 76380.0 58950.0 ;
      RECT  75675.0 60295.0 76380.0 58950.0 ;
      RECT  75675.0 60295.0 76380.0 61640.0 ;
      RECT  75675.0 62985.0 76380.0 61640.0 ;
      RECT  75675.0 62985.0 76380.0 64330.0 ;
      RECT  75675.0 65675.0 76380.0 64330.0 ;
      RECT  75675.0 65675.0 76380.0 67020.0 ;
      RECT  75675.0 68365.0 76380.0 67020.0 ;
      RECT  75675.0 68365.0 76380.0 69710.0 ;
      RECT  75675.0 71055.0 76380.0 69710.0 ;
      RECT  75675.0 71055.0 76380.0 72400.0 ;
      RECT  75675.0 73745.0 76380.0 72400.0 ;
      RECT  75675.0 73745.0 76380.0 75090.0 ;
      RECT  75675.0 76435.0 76380.0 75090.0 ;
      RECT  75675.0 76435.0 76380.0 77780.0 ;
      RECT  75675.0 79125.0 76380.0 77780.0 ;
      RECT  75675.0 79125.0 76380.0 80470.0 ;
      RECT  75675.0 81815.0 76380.0 80470.0 ;
      RECT  75675.0 81815.0 76380.0 83160.0 ;
      RECT  75675.0 84505.0 76380.0 83160.0 ;
      RECT  75675.0 84505.0 76380.0 85850.0 ;
      RECT  75675.0 87195.0 76380.0 85850.0 ;
      RECT  75675.0 87195.0 76380.0 88540.0 ;
      RECT  75675.0 89885.0 76380.0 88540.0 ;
      RECT  75675.0 89885.0 76380.0 91230.0 ;
      RECT  75675.0 92575.0 76380.0 91230.0 ;
      RECT  75675.0 92575.0 76380.0 93920.0 ;
      RECT  75675.0 95265.0 76380.0 93920.0 ;
      RECT  75675.0 95265.0 76380.0 96610.0 ;
      RECT  75675.0 97955.0 76380.0 96610.0 ;
      RECT  75675.0 97955.0 76380.0 99300.0 ;
      RECT  75675.0 100645.0 76380.0 99300.0 ;
      RECT  75675.0 100645.0 76380.0 101990.0 ;
      RECT  75675.0 103335.0 76380.0 101990.0 ;
      RECT  75675.0 103335.0 76380.0 104680.0 ;
      RECT  75675.0 106025.0 76380.0 104680.0 ;
      RECT  75675.0 106025.0 76380.0 107370.0 ;
      RECT  75675.0 108715.0 76380.0 107370.0 ;
      RECT  75675.0 108715.0 76380.0 110060.0 ;
      RECT  75675.0 111405.0 76380.0 110060.0 ;
      RECT  75675.0 111405.0 76380.0 112750.0 ;
      RECT  75675.0 114095.0 76380.0 112750.0 ;
      RECT  76380.0 28015.0 77085.0 29360.0 ;
      RECT  76380.0 30705.0 77085.0 29360.0 ;
      RECT  76380.0 30705.0 77085.0 32050.0 ;
      RECT  76380.0 33395.0 77085.0 32050.0 ;
      RECT  76380.0 33395.0 77085.0 34740.0 ;
      RECT  76380.0 36085.0 77085.0 34740.0 ;
      RECT  76380.0 36085.0 77085.0 37430.0 ;
      RECT  76380.0 38775.0 77085.0 37430.0 ;
      RECT  76380.0 38775.0 77085.0 40120.0 ;
      RECT  76380.0 41465.0 77085.0 40120.0 ;
      RECT  76380.0 41465.0 77085.0 42810.0 ;
      RECT  76380.0 44155.0 77085.0 42810.0 ;
      RECT  76380.0 44155.0 77085.0 45500.0 ;
      RECT  76380.0 46845.0 77085.0 45500.0 ;
      RECT  76380.0 46845.0 77085.0 48190.0 ;
      RECT  76380.0 49535.0 77085.0 48190.0 ;
      RECT  76380.0 49535.0 77085.0 50880.0 ;
      RECT  76380.0 52225.0 77085.0 50880.0 ;
      RECT  76380.0 52225.0 77085.0 53570.0 ;
      RECT  76380.0 54915.0 77085.0 53570.0 ;
      RECT  76380.0 54915.0 77085.0 56260.0 ;
      RECT  76380.0 57605.0 77085.0 56260.0 ;
      RECT  76380.0 57605.0 77085.0 58950.0 ;
      RECT  76380.0 60295.0 77085.0 58950.0 ;
      RECT  76380.0 60295.0 77085.0 61640.0 ;
      RECT  76380.0 62985.0 77085.0 61640.0 ;
      RECT  76380.0 62985.0 77085.0 64330.0 ;
      RECT  76380.0 65675.0 77085.0 64330.0 ;
      RECT  76380.0 65675.0 77085.0 67020.0 ;
      RECT  76380.0 68365.0 77085.0 67020.0 ;
      RECT  76380.0 68365.0 77085.0 69710.0 ;
      RECT  76380.0 71055.0 77085.0 69710.0 ;
      RECT  76380.0 71055.0 77085.0 72400.0 ;
      RECT  76380.0 73745.0 77085.0 72400.0 ;
      RECT  76380.0 73745.0 77085.0 75090.0 ;
      RECT  76380.0 76435.0 77085.0 75090.0 ;
      RECT  76380.0 76435.0 77085.0 77780.0 ;
      RECT  76380.0 79125.0 77085.0 77780.0 ;
      RECT  76380.0 79125.0 77085.0 80470.0 ;
      RECT  76380.0 81815.0 77085.0 80470.0 ;
      RECT  76380.0 81815.0 77085.0 83160.0 ;
      RECT  76380.0 84505.0 77085.0 83160.0 ;
      RECT  76380.0 84505.0 77085.0 85850.0 ;
      RECT  76380.0 87195.0 77085.0 85850.0 ;
      RECT  76380.0 87195.0 77085.0 88540.0 ;
      RECT  76380.0 89885.0 77085.0 88540.0 ;
      RECT  76380.0 89885.0 77085.0 91230.0 ;
      RECT  76380.0 92575.0 77085.0 91230.0 ;
      RECT  76380.0 92575.0 77085.0 93920.0 ;
      RECT  76380.0 95265.0 77085.0 93920.0 ;
      RECT  76380.0 95265.0 77085.0 96610.0 ;
      RECT  76380.0 97955.0 77085.0 96610.0 ;
      RECT  76380.0 97955.0 77085.0 99300.0 ;
      RECT  76380.0 100645.0 77085.0 99300.0 ;
      RECT  76380.0 100645.0 77085.0 101990.0 ;
      RECT  76380.0 103335.0 77085.0 101990.0 ;
      RECT  76380.0 103335.0 77085.0 104680.0 ;
      RECT  76380.0 106025.0 77085.0 104680.0 ;
      RECT  76380.0 106025.0 77085.0 107370.0 ;
      RECT  76380.0 108715.0 77085.0 107370.0 ;
      RECT  76380.0 108715.0 77085.0 110060.0 ;
      RECT  76380.0 111405.0 77085.0 110060.0 ;
      RECT  76380.0 111405.0 77085.0 112750.0 ;
      RECT  76380.0 114095.0 77085.0 112750.0 ;
      RECT  77085.0 28015.0 77790.0 29360.0 ;
      RECT  77085.0 30705.0 77790.0 29360.0 ;
      RECT  77085.0 30705.0 77790.0 32050.0 ;
      RECT  77085.0 33395.0 77790.0 32050.0 ;
      RECT  77085.0 33395.0 77790.0 34740.0 ;
      RECT  77085.0 36085.0 77790.0 34740.0 ;
      RECT  77085.0 36085.0 77790.0 37430.0 ;
      RECT  77085.0 38775.0 77790.0 37430.0 ;
      RECT  77085.0 38775.0 77790.0 40120.0 ;
      RECT  77085.0 41465.0 77790.0 40120.0 ;
      RECT  77085.0 41465.0 77790.0 42810.0 ;
      RECT  77085.0 44155.0 77790.0 42810.0 ;
      RECT  77085.0 44155.0 77790.0 45500.0 ;
      RECT  77085.0 46845.0 77790.0 45500.0 ;
      RECT  77085.0 46845.0 77790.0 48190.0 ;
      RECT  77085.0 49535.0 77790.0 48190.0 ;
      RECT  77085.0 49535.0 77790.0 50880.0 ;
      RECT  77085.0 52225.0 77790.0 50880.0 ;
      RECT  77085.0 52225.0 77790.0 53570.0 ;
      RECT  77085.0 54915.0 77790.0 53570.0 ;
      RECT  77085.0 54915.0 77790.0 56260.0 ;
      RECT  77085.0 57605.0 77790.0 56260.0 ;
      RECT  77085.0 57605.0 77790.0 58950.0 ;
      RECT  77085.0 60295.0 77790.0 58950.0 ;
      RECT  77085.0 60295.0 77790.0 61640.0 ;
      RECT  77085.0 62985.0 77790.0 61640.0 ;
      RECT  77085.0 62985.0 77790.0 64330.0 ;
      RECT  77085.0 65675.0 77790.0 64330.0 ;
      RECT  77085.0 65675.0 77790.0 67020.0 ;
      RECT  77085.0 68365.0 77790.0 67020.0 ;
      RECT  77085.0 68365.0 77790.0 69710.0 ;
      RECT  77085.0 71055.0 77790.0 69710.0 ;
      RECT  77085.0 71055.0 77790.0 72400.0 ;
      RECT  77085.0 73745.0 77790.0 72400.0 ;
      RECT  77085.0 73745.0 77790.0 75090.0 ;
      RECT  77085.0 76435.0 77790.0 75090.0 ;
      RECT  77085.0 76435.0 77790.0 77780.0 ;
      RECT  77085.0 79125.0 77790.0 77780.0 ;
      RECT  77085.0 79125.0 77790.0 80470.0 ;
      RECT  77085.0 81815.0 77790.0 80470.0 ;
      RECT  77085.0 81815.0 77790.0 83160.0 ;
      RECT  77085.0 84505.0 77790.0 83160.0 ;
      RECT  77085.0 84505.0 77790.0 85850.0 ;
      RECT  77085.0 87195.0 77790.0 85850.0 ;
      RECT  77085.0 87195.0 77790.0 88540.0 ;
      RECT  77085.0 89885.0 77790.0 88540.0 ;
      RECT  77085.0 89885.0 77790.0 91230.0 ;
      RECT  77085.0 92575.0 77790.0 91230.0 ;
      RECT  77085.0 92575.0 77790.0 93920.0 ;
      RECT  77085.0 95265.0 77790.0 93920.0 ;
      RECT  77085.0 95265.0 77790.0 96610.0 ;
      RECT  77085.0 97955.0 77790.0 96610.0 ;
      RECT  77085.0 97955.0 77790.0 99300.0 ;
      RECT  77085.0 100645.0 77790.0 99300.0 ;
      RECT  77085.0 100645.0 77790.0 101990.0 ;
      RECT  77085.0 103335.0 77790.0 101990.0 ;
      RECT  77085.0 103335.0 77790.0 104680.0 ;
      RECT  77085.0 106025.0 77790.0 104680.0 ;
      RECT  77085.0 106025.0 77790.0 107370.0 ;
      RECT  77085.0 108715.0 77790.0 107370.0 ;
      RECT  77085.0 108715.0 77790.0 110060.0 ;
      RECT  77085.0 111405.0 77790.0 110060.0 ;
      RECT  77085.0 111405.0 77790.0 112750.0 ;
      RECT  77085.0 114095.0 77790.0 112750.0 ;
      RECT  77790.0 28015.0 78495.0 29360.0 ;
      RECT  77790.0 30705.0 78495.0 29360.0 ;
      RECT  77790.0 30705.0 78495.0 32050.0 ;
      RECT  77790.0 33395.0 78495.0 32050.0 ;
      RECT  77790.0 33395.0 78495.0 34740.0 ;
      RECT  77790.0 36085.0 78495.0 34740.0 ;
      RECT  77790.0 36085.0 78495.0 37430.0 ;
      RECT  77790.0 38775.0 78495.0 37430.0 ;
      RECT  77790.0 38775.0 78495.0 40120.0 ;
      RECT  77790.0 41465.0 78495.0 40120.0 ;
      RECT  77790.0 41465.0 78495.0 42810.0 ;
      RECT  77790.0 44155.0 78495.0 42810.0 ;
      RECT  77790.0 44155.0 78495.0 45500.0 ;
      RECT  77790.0 46845.0 78495.0 45500.0 ;
      RECT  77790.0 46845.0 78495.0 48190.0 ;
      RECT  77790.0 49535.0 78495.0 48190.0 ;
      RECT  77790.0 49535.0 78495.0 50880.0 ;
      RECT  77790.0 52225.0 78495.0 50880.0 ;
      RECT  77790.0 52225.0 78495.0 53570.0 ;
      RECT  77790.0 54915.0 78495.0 53570.0 ;
      RECT  77790.0 54915.0 78495.0 56260.0 ;
      RECT  77790.0 57605.0 78495.0 56260.0 ;
      RECT  77790.0 57605.0 78495.0 58950.0 ;
      RECT  77790.0 60295.0 78495.0 58950.0 ;
      RECT  77790.0 60295.0 78495.0 61640.0 ;
      RECT  77790.0 62985.0 78495.0 61640.0 ;
      RECT  77790.0 62985.0 78495.0 64330.0 ;
      RECT  77790.0 65675.0 78495.0 64330.0 ;
      RECT  77790.0 65675.0 78495.0 67020.0 ;
      RECT  77790.0 68365.0 78495.0 67020.0 ;
      RECT  77790.0 68365.0 78495.0 69710.0 ;
      RECT  77790.0 71055.0 78495.0 69710.0 ;
      RECT  77790.0 71055.0 78495.0 72400.0 ;
      RECT  77790.0 73745.0 78495.0 72400.0 ;
      RECT  77790.0 73745.0 78495.0 75090.0 ;
      RECT  77790.0 76435.0 78495.0 75090.0 ;
      RECT  77790.0 76435.0 78495.0 77780.0 ;
      RECT  77790.0 79125.0 78495.0 77780.0 ;
      RECT  77790.0 79125.0 78495.0 80470.0 ;
      RECT  77790.0 81815.0 78495.0 80470.0 ;
      RECT  77790.0 81815.0 78495.0 83160.0 ;
      RECT  77790.0 84505.0 78495.0 83160.0 ;
      RECT  77790.0 84505.0 78495.0 85850.0 ;
      RECT  77790.0 87195.0 78495.0 85850.0 ;
      RECT  77790.0 87195.0 78495.0 88540.0 ;
      RECT  77790.0 89885.0 78495.0 88540.0 ;
      RECT  77790.0 89885.0 78495.0 91230.0 ;
      RECT  77790.0 92575.0 78495.0 91230.0 ;
      RECT  77790.0 92575.0 78495.0 93920.0 ;
      RECT  77790.0 95265.0 78495.0 93920.0 ;
      RECT  77790.0 95265.0 78495.0 96610.0 ;
      RECT  77790.0 97955.0 78495.0 96610.0 ;
      RECT  77790.0 97955.0 78495.0 99300.0 ;
      RECT  77790.0 100645.0 78495.0 99300.0 ;
      RECT  77790.0 100645.0 78495.0 101990.0 ;
      RECT  77790.0 103335.0 78495.0 101990.0 ;
      RECT  77790.0 103335.0 78495.0 104680.0 ;
      RECT  77790.0 106025.0 78495.0 104680.0 ;
      RECT  77790.0 106025.0 78495.0 107370.0 ;
      RECT  77790.0 108715.0 78495.0 107370.0 ;
      RECT  77790.0 108715.0 78495.0 110060.0 ;
      RECT  77790.0 111405.0 78495.0 110060.0 ;
      RECT  77790.0 111405.0 78495.0 112750.0 ;
      RECT  77790.0 114095.0 78495.0 112750.0 ;
      RECT  78495.0 28015.0 79200.0 29360.0 ;
      RECT  78495.0 30705.0 79200.0 29360.0 ;
      RECT  78495.0 30705.0 79200.0 32050.0 ;
      RECT  78495.0 33395.0 79200.0 32050.0 ;
      RECT  78495.0 33395.0 79200.0 34740.0 ;
      RECT  78495.0 36085.0 79200.0 34740.0 ;
      RECT  78495.0 36085.0 79200.0 37430.0 ;
      RECT  78495.0 38775.0 79200.0 37430.0 ;
      RECT  78495.0 38775.0 79200.0 40120.0 ;
      RECT  78495.0 41465.0 79200.0 40120.0 ;
      RECT  78495.0 41465.0 79200.0 42810.0 ;
      RECT  78495.0 44155.0 79200.0 42810.0 ;
      RECT  78495.0 44155.0 79200.0 45500.0 ;
      RECT  78495.0 46845.0 79200.0 45500.0 ;
      RECT  78495.0 46845.0 79200.0 48190.0 ;
      RECT  78495.0 49535.0 79200.0 48190.0 ;
      RECT  78495.0 49535.0 79200.0 50880.0 ;
      RECT  78495.0 52225.0 79200.0 50880.0 ;
      RECT  78495.0 52225.0 79200.0 53570.0 ;
      RECT  78495.0 54915.0 79200.0 53570.0 ;
      RECT  78495.0 54915.0 79200.0 56260.0 ;
      RECT  78495.0 57605.0 79200.0 56260.0 ;
      RECT  78495.0 57605.0 79200.0 58950.0 ;
      RECT  78495.0 60295.0 79200.0 58950.0 ;
      RECT  78495.0 60295.0 79200.0 61640.0 ;
      RECT  78495.0 62985.0 79200.0 61640.0 ;
      RECT  78495.0 62985.0 79200.0 64330.0 ;
      RECT  78495.0 65675.0 79200.0 64330.0 ;
      RECT  78495.0 65675.0 79200.0 67020.0 ;
      RECT  78495.0 68365.0 79200.0 67020.0 ;
      RECT  78495.0 68365.0 79200.0 69710.0 ;
      RECT  78495.0 71055.0 79200.0 69710.0 ;
      RECT  78495.0 71055.0 79200.0 72400.0 ;
      RECT  78495.0 73745.0 79200.0 72400.0 ;
      RECT  78495.0 73745.0 79200.0 75090.0 ;
      RECT  78495.0 76435.0 79200.0 75090.0 ;
      RECT  78495.0 76435.0 79200.0 77780.0 ;
      RECT  78495.0 79125.0 79200.0 77780.0 ;
      RECT  78495.0 79125.0 79200.0 80470.0 ;
      RECT  78495.0 81815.0 79200.0 80470.0 ;
      RECT  78495.0 81815.0 79200.0 83160.0 ;
      RECT  78495.0 84505.0 79200.0 83160.0 ;
      RECT  78495.0 84505.0 79200.0 85850.0 ;
      RECT  78495.0 87195.0 79200.0 85850.0 ;
      RECT  78495.0 87195.0 79200.0 88540.0 ;
      RECT  78495.0 89885.0 79200.0 88540.0 ;
      RECT  78495.0 89885.0 79200.0 91230.0 ;
      RECT  78495.0 92575.0 79200.0 91230.0 ;
      RECT  78495.0 92575.0 79200.0 93920.0 ;
      RECT  78495.0 95265.0 79200.0 93920.0 ;
      RECT  78495.0 95265.0 79200.0 96610.0 ;
      RECT  78495.0 97955.0 79200.0 96610.0 ;
      RECT  78495.0 97955.0 79200.0 99300.0 ;
      RECT  78495.0 100645.0 79200.0 99300.0 ;
      RECT  78495.0 100645.0 79200.0 101990.0 ;
      RECT  78495.0 103335.0 79200.0 101990.0 ;
      RECT  78495.0 103335.0 79200.0 104680.0 ;
      RECT  78495.0 106025.0 79200.0 104680.0 ;
      RECT  78495.0 106025.0 79200.0 107370.0 ;
      RECT  78495.0 108715.0 79200.0 107370.0 ;
      RECT  78495.0 108715.0 79200.0 110060.0 ;
      RECT  78495.0 111405.0 79200.0 110060.0 ;
      RECT  78495.0 111405.0 79200.0 112750.0 ;
      RECT  78495.0 114095.0 79200.0 112750.0 ;
      RECT  79200.0 28015.0 79905.0 29360.0 ;
      RECT  79200.0 30705.0 79905.0 29360.0 ;
      RECT  79200.0 30705.0 79905.0 32050.0 ;
      RECT  79200.0 33395.0 79905.0 32050.0 ;
      RECT  79200.0 33395.0 79905.0 34740.0 ;
      RECT  79200.0 36085.0 79905.0 34740.0 ;
      RECT  79200.0 36085.0 79905.0 37430.0 ;
      RECT  79200.0 38775.0 79905.0 37430.0 ;
      RECT  79200.0 38775.0 79905.0 40120.0 ;
      RECT  79200.0 41465.0 79905.0 40120.0 ;
      RECT  79200.0 41465.0 79905.0 42810.0 ;
      RECT  79200.0 44155.0 79905.0 42810.0 ;
      RECT  79200.0 44155.0 79905.0 45500.0 ;
      RECT  79200.0 46845.0 79905.0 45500.0 ;
      RECT  79200.0 46845.0 79905.0 48190.0 ;
      RECT  79200.0 49535.0 79905.0 48190.0 ;
      RECT  79200.0 49535.0 79905.0 50880.0 ;
      RECT  79200.0 52225.0 79905.0 50880.0 ;
      RECT  79200.0 52225.0 79905.0 53570.0 ;
      RECT  79200.0 54915.0 79905.0 53570.0 ;
      RECT  79200.0 54915.0 79905.0 56260.0 ;
      RECT  79200.0 57605.0 79905.0 56260.0 ;
      RECT  79200.0 57605.0 79905.0 58950.0 ;
      RECT  79200.0 60295.0 79905.0 58950.0 ;
      RECT  79200.0 60295.0 79905.0 61640.0 ;
      RECT  79200.0 62985.0 79905.0 61640.0 ;
      RECT  79200.0 62985.0 79905.0 64330.0 ;
      RECT  79200.0 65675.0 79905.0 64330.0 ;
      RECT  79200.0 65675.0 79905.0 67020.0 ;
      RECT  79200.0 68365.0 79905.0 67020.0 ;
      RECT  79200.0 68365.0 79905.0 69710.0 ;
      RECT  79200.0 71055.0 79905.0 69710.0 ;
      RECT  79200.0 71055.0 79905.0 72400.0 ;
      RECT  79200.0 73745.0 79905.0 72400.0 ;
      RECT  79200.0 73745.0 79905.0 75090.0 ;
      RECT  79200.0 76435.0 79905.0 75090.0 ;
      RECT  79200.0 76435.0 79905.0 77780.0 ;
      RECT  79200.0 79125.0 79905.0 77780.0 ;
      RECT  79200.0 79125.0 79905.0 80470.0 ;
      RECT  79200.0 81815.0 79905.0 80470.0 ;
      RECT  79200.0 81815.0 79905.0 83160.0 ;
      RECT  79200.0 84505.0 79905.0 83160.0 ;
      RECT  79200.0 84505.0 79905.0 85850.0 ;
      RECT  79200.0 87195.0 79905.0 85850.0 ;
      RECT  79200.0 87195.0 79905.0 88540.0 ;
      RECT  79200.0 89885.0 79905.0 88540.0 ;
      RECT  79200.0 89885.0 79905.0 91230.0 ;
      RECT  79200.0 92575.0 79905.0 91230.0 ;
      RECT  79200.0 92575.0 79905.0 93920.0 ;
      RECT  79200.0 95265.0 79905.0 93920.0 ;
      RECT  79200.0 95265.0 79905.0 96610.0 ;
      RECT  79200.0 97955.0 79905.0 96610.0 ;
      RECT  79200.0 97955.0 79905.0 99300.0 ;
      RECT  79200.0 100645.0 79905.0 99300.0 ;
      RECT  79200.0 100645.0 79905.0 101990.0 ;
      RECT  79200.0 103335.0 79905.0 101990.0 ;
      RECT  79200.0 103335.0 79905.0 104680.0 ;
      RECT  79200.0 106025.0 79905.0 104680.0 ;
      RECT  79200.0 106025.0 79905.0 107370.0 ;
      RECT  79200.0 108715.0 79905.0 107370.0 ;
      RECT  79200.0 108715.0 79905.0 110060.0 ;
      RECT  79200.0 111405.0 79905.0 110060.0 ;
      RECT  79200.0 111405.0 79905.0 112750.0 ;
      RECT  79200.0 114095.0 79905.0 112750.0 ;
      RECT  79905.0 28015.0 80610.0 29360.0 ;
      RECT  79905.0 30705.0 80610.0 29360.0 ;
      RECT  79905.0 30705.0 80610.0 32050.0 ;
      RECT  79905.0 33395.0 80610.0 32050.0 ;
      RECT  79905.0 33395.0 80610.0 34740.0 ;
      RECT  79905.0 36085.0 80610.0 34740.0 ;
      RECT  79905.0 36085.0 80610.0 37430.0 ;
      RECT  79905.0 38775.0 80610.0 37430.0 ;
      RECT  79905.0 38775.0 80610.0 40120.0 ;
      RECT  79905.0 41465.0 80610.0 40120.0 ;
      RECT  79905.0 41465.0 80610.0 42810.0 ;
      RECT  79905.0 44155.0 80610.0 42810.0 ;
      RECT  79905.0 44155.0 80610.0 45500.0 ;
      RECT  79905.0 46845.0 80610.0 45500.0 ;
      RECT  79905.0 46845.0 80610.0 48190.0 ;
      RECT  79905.0 49535.0 80610.0 48190.0 ;
      RECT  79905.0 49535.0 80610.0 50880.0 ;
      RECT  79905.0 52225.0 80610.0 50880.0 ;
      RECT  79905.0 52225.0 80610.0 53570.0 ;
      RECT  79905.0 54915.0 80610.0 53570.0 ;
      RECT  79905.0 54915.0 80610.0 56260.0 ;
      RECT  79905.0 57605.0 80610.0 56260.0 ;
      RECT  79905.0 57605.0 80610.0 58950.0 ;
      RECT  79905.0 60295.0 80610.0 58950.0 ;
      RECT  79905.0 60295.0 80610.0 61640.0 ;
      RECT  79905.0 62985.0 80610.0 61640.0 ;
      RECT  79905.0 62985.0 80610.0 64330.0 ;
      RECT  79905.0 65675.0 80610.0 64330.0 ;
      RECT  79905.0 65675.0 80610.0 67020.0 ;
      RECT  79905.0 68365.0 80610.0 67020.0 ;
      RECT  79905.0 68365.0 80610.0 69710.0 ;
      RECT  79905.0 71055.0 80610.0 69710.0 ;
      RECT  79905.0 71055.0 80610.0 72400.0 ;
      RECT  79905.0 73745.0 80610.0 72400.0 ;
      RECT  79905.0 73745.0 80610.0 75090.0 ;
      RECT  79905.0 76435.0 80610.0 75090.0 ;
      RECT  79905.0 76435.0 80610.0 77780.0 ;
      RECT  79905.0 79125.0 80610.0 77780.0 ;
      RECT  79905.0 79125.0 80610.0 80470.0 ;
      RECT  79905.0 81815.0 80610.0 80470.0 ;
      RECT  79905.0 81815.0 80610.0 83160.0 ;
      RECT  79905.0 84505.0 80610.0 83160.0 ;
      RECT  79905.0 84505.0 80610.0 85850.0 ;
      RECT  79905.0 87195.0 80610.0 85850.0 ;
      RECT  79905.0 87195.0 80610.0 88540.0 ;
      RECT  79905.0 89885.0 80610.0 88540.0 ;
      RECT  79905.0 89885.0 80610.0 91230.0 ;
      RECT  79905.0 92575.0 80610.0 91230.0 ;
      RECT  79905.0 92575.0 80610.0 93920.0 ;
      RECT  79905.0 95265.0 80610.0 93920.0 ;
      RECT  79905.0 95265.0 80610.0 96610.0 ;
      RECT  79905.0 97955.0 80610.0 96610.0 ;
      RECT  79905.0 97955.0 80610.0 99300.0 ;
      RECT  79905.0 100645.0 80610.0 99300.0 ;
      RECT  79905.0 100645.0 80610.0 101990.0 ;
      RECT  79905.0 103335.0 80610.0 101990.0 ;
      RECT  79905.0 103335.0 80610.0 104680.0 ;
      RECT  79905.0 106025.0 80610.0 104680.0 ;
      RECT  79905.0 106025.0 80610.0 107370.0 ;
      RECT  79905.0 108715.0 80610.0 107370.0 ;
      RECT  79905.0 108715.0 80610.0 110060.0 ;
      RECT  79905.0 111405.0 80610.0 110060.0 ;
      RECT  79905.0 111405.0 80610.0 112750.0 ;
      RECT  79905.0 114095.0 80610.0 112750.0 ;
      RECT  80610.0 28015.0 81315.0 29360.0 ;
      RECT  80610.0 30705.0 81315.0 29360.0 ;
      RECT  80610.0 30705.0 81315.0 32050.0 ;
      RECT  80610.0 33395.0 81315.0 32050.0 ;
      RECT  80610.0 33395.0 81315.0 34740.0 ;
      RECT  80610.0 36085.0 81315.0 34740.0 ;
      RECT  80610.0 36085.0 81315.0 37430.0 ;
      RECT  80610.0 38775.0 81315.0 37430.0 ;
      RECT  80610.0 38775.0 81315.0 40120.0 ;
      RECT  80610.0 41465.0 81315.0 40120.0 ;
      RECT  80610.0 41465.0 81315.0 42810.0 ;
      RECT  80610.0 44155.0 81315.0 42810.0 ;
      RECT  80610.0 44155.0 81315.0 45500.0 ;
      RECT  80610.0 46845.0 81315.0 45500.0 ;
      RECT  80610.0 46845.0 81315.0 48190.0 ;
      RECT  80610.0 49535.0 81315.0 48190.0 ;
      RECT  80610.0 49535.0 81315.0 50880.0 ;
      RECT  80610.0 52225.0 81315.0 50880.0 ;
      RECT  80610.0 52225.0 81315.0 53570.0 ;
      RECT  80610.0 54915.0 81315.0 53570.0 ;
      RECT  80610.0 54915.0 81315.0 56260.0 ;
      RECT  80610.0 57605.0 81315.0 56260.0 ;
      RECT  80610.0 57605.0 81315.0 58950.0 ;
      RECT  80610.0 60295.0 81315.0 58950.0 ;
      RECT  80610.0 60295.0 81315.0 61640.0 ;
      RECT  80610.0 62985.0 81315.0 61640.0 ;
      RECT  80610.0 62985.0 81315.0 64330.0 ;
      RECT  80610.0 65675.0 81315.0 64330.0 ;
      RECT  80610.0 65675.0 81315.0 67020.0 ;
      RECT  80610.0 68365.0 81315.0 67020.0 ;
      RECT  80610.0 68365.0 81315.0 69710.0 ;
      RECT  80610.0 71055.0 81315.0 69710.0 ;
      RECT  80610.0 71055.0 81315.0 72400.0 ;
      RECT  80610.0 73745.0 81315.0 72400.0 ;
      RECT  80610.0 73745.0 81315.0 75090.0 ;
      RECT  80610.0 76435.0 81315.0 75090.0 ;
      RECT  80610.0 76435.0 81315.0 77780.0 ;
      RECT  80610.0 79125.0 81315.0 77780.0 ;
      RECT  80610.0 79125.0 81315.0 80470.0 ;
      RECT  80610.0 81815.0 81315.0 80470.0 ;
      RECT  80610.0 81815.0 81315.0 83160.0 ;
      RECT  80610.0 84505.0 81315.0 83160.0 ;
      RECT  80610.0 84505.0 81315.0 85850.0 ;
      RECT  80610.0 87195.0 81315.0 85850.0 ;
      RECT  80610.0 87195.0 81315.0 88540.0 ;
      RECT  80610.0 89885.0 81315.0 88540.0 ;
      RECT  80610.0 89885.0 81315.0 91230.0 ;
      RECT  80610.0 92575.0 81315.0 91230.0 ;
      RECT  80610.0 92575.0 81315.0 93920.0 ;
      RECT  80610.0 95265.0 81315.0 93920.0 ;
      RECT  80610.0 95265.0 81315.0 96610.0 ;
      RECT  80610.0 97955.0 81315.0 96610.0 ;
      RECT  80610.0 97955.0 81315.0 99300.0 ;
      RECT  80610.0 100645.0 81315.0 99300.0 ;
      RECT  80610.0 100645.0 81315.0 101990.0 ;
      RECT  80610.0 103335.0 81315.0 101990.0 ;
      RECT  80610.0 103335.0 81315.0 104680.0 ;
      RECT  80610.0 106025.0 81315.0 104680.0 ;
      RECT  80610.0 106025.0 81315.0 107370.0 ;
      RECT  80610.0 108715.0 81315.0 107370.0 ;
      RECT  80610.0 108715.0 81315.0 110060.0 ;
      RECT  80610.0 111405.0 81315.0 110060.0 ;
      RECT  80610.0 111405.0 81315.0 112750.0 ;
      RECT  80610.0 114095.0 81315.0 112750.0 ;
      RECT  81315.0 28015.0 82020.0 29360.0 ;
      RECT  81315.0 30705.0 82020.0 29360.0 ;
      RECT  81315.0 30705.0 82020.0 32050.0 ;
      RECT  81315.0 33395.0 82020.0 32050.0 ;
      RECT  81315.0 33395.0 82020.0 34740.0 ;
      RECT  81315.0 36085.0 82020.0 34740.0 ;
      RECT  81315.0 36085.0 82020.0 37430.0 ;
      RECT  81315.0 38775.0 82020.0 37430.0 ;
      RECT  81315.0 38775.0 82020.0 40120.0 ;
      RECT  81315.0 41465.0 82020.0 40120.0 ;
      RECT  81315.0 41465.0 82020.0 42810.0 ;
      RECT  81315.0 44155.0 82020.0 42810.0 ;
      RECT  81315.0 44155.0 82020.0 45500.0 ;
      RECT  81315.0 46845.0 82020.0 45500.0 ;
      RECT  81315.0 46845.0 82020.0 48190.0 ;
      RECT  81315.0 49535.0 82020.0 48190.0 ;
      RECT  81315.0 49535.0 82020.0 50880.0 ;
      RECT  81315.0 52225.0 82020.0 50880.0 ;
      RECT  81315.0 52225.0 82020.0 53570.0 ;
      RECT  81315.0 54915.0 82020.0 53570.0 ;
      RECT  81315.0 54915.0 82020.0 56260.0 ;
      RECT  81315.0 57605.0 82020.0 56260.0 ;
      RECT  81315.0 57605.0 82020.0 58950.0 ;
      RECT  81315.0 60295.0 82020.0 58950.0 ;
      RECT  81315.0 60295.0 82020.0 61640.0 ;
      RECT  81315.0 62985.0 82020.0 61640.0 ;
      RECT  81315.0 62985.0 82020.0 64330.0 ;
      RECT  81315.0 65675.0 82020.0 64330.0 ;
      RECT  81315.0 65675.0 82020.0 67020.0 ;
      RECT  81315.0 68365.0 82020.0 67020.0 ;
      RECT  81315.0 68365.0 82020.0 69710.0 ;
      RECT  81315.0 71055.0 82020.0 69710.0 ;
      RECT  81315.0 71055.0 82020.0 72400.0 ;
      RECT  81315.0 73745.0 82020.0 72400.0 ;
      RECT  81315.0 73745.0 82020.0 75090.0 ;
      RECT  81315.0 76435.0 82020.0 75090.0 ;
      RECT  81315.0 76435.0 82020.0 77780.0 ;
      RECT  81315.0 79125.0 82020.0 77780.0 ;
      RECT  81315.0 79125.0 82020.0 80470.0 ;
      RECT  81315.0 81815.0 82020.0 80470.0 ;
      RECT  81315.0 81815.0 82020.0 83160.0 ;
      RECT  81315.0 84505.0 82020.0 83160.0 ;
      RECT  81315.0 84505.0 82020.0 85850.0 ;
      RECT  81315.0 87195.0 82020.0 85850.0 ;
      RECT  81315.0 87195.0 82020.0 88540.0 ;
      RECT  81315.0 89885.0 82020.0 88540.0 ;
      RECT  81315.0 89885.0 82020.0 91230.0 ;
      RECT  81315.0 92575.0 82020.0 91230.0 ;
      RECT  81315.0 92575.0 82020.0 93920.0 ;
      RECT  81315.0 95265.0 82020.0 93920.0 ;
      RECT  81315.0 95265.0 82020.0 96610.0 ;
      RECT  81315.0 97955.0 82020.0 96610.0 ;
      RECT  81315.0 97955.0 82020.0 99300.0 ;
      RECT  81315.0 100645.0 82020.0 99300.0 ;
      RECT  81315.0 100645.0 82020.0 101990.0 ;
      RECT  81315.0 103335.0 82020.0 101990.0 ;
      RECT  81315.0 103335.0 82020.0 104680.0 ;
      RECT  81315.0 106025.0 82020.0 104680.0 ;
      RECT  81315.0 106025.0 82020.0 107370.0 ;
      RECT  81315.0 108715.0 82020.0 107370.0 ;
      RECT  81315.0 108715.0 82020.0 110060.0 ;
      RECT  81315.0 111405.0 82020.0 110060.0 ;
      RECT  81315.0 111405.0 82020.0 112750.0 ;
      RECT  81315.0 114095.0 82020.0 112750.0 ;
      RECT  82020.0 28015.0 82725.0 29360.0 ;
      RECT  82020.0 30705.0 82725.0 29360.0 ;
      RECT  82020.0 30705.0 82725.0 32050.0 ;
      RECT  82020.0 33395.0 82725.0 32050.0 ;
      RECT  82020.0 33395.0 82725.0 34740.0 ;
      RECT  82020.0 36085.0 82725.0 34740.0 ;
      RECT  82020.0 36085.0 82725.0 37430.0 ;
      RECT  82020.0 38775.0 82725.0 37430.0 ;
      RECT  82020.0 38775.0 82725.0 40120.0 ;
      RECT  82020.0 41465.0 82725.0 40120.0 ;
      RECT  82020.0 41465.0 82725.0 42810.0 ;
      RECT  82020.0 44155.0 82725.0 42810.0 ;
      RECT  82020.0 44155.0 82725.0 45500.0 ;
      RECT  82020.0 46845.0 82725.0 45500.0 ;
      RECT  82020.0 46845.0 82725.0 48190.0 ;
      RECT  82020.0 49535.0 82725.0 48190.0 ;
      RECT  82020.0 49535.0 82725.0 50880.0 ;
      RECT  82020.0 52225.0 82725.0 50880.0 ;
      RECT  82020.0 52225.0 82725.0 53570.0 ;
      RECT  82020.0 54915.0 82725.0 53570.0 ;
      RECT  82020.0 54915.0 82725.0 56260.0 ;
      RECT  82020.0 57605.0 82725.0 56260.0 ;
      RECT  82020.0 57605.0 82725.0 58950.0 ;
      RECT  82020.0 60295.0 82725.0 58950.0 ;
      RECT  82020.0 60295.0 82725.0 61640.0 ;
      RECT  82020.0 62985.0 82725.0 61640.0 ;
      RECT  82020.0 62985.0 82725.0 64330.0 ;
      RECT  82020.0 65675.0 82725.0 64330.0 ;
      RECT  82020.0 65675.0 82725.0 67020.0 ;
      RECT  82020.0 68365.0 82725.0 67020.0 ;
      RECT  82020.0 68365.0 82725.0 69710.0 ;
      RECT  82020.0 71055.0 82725.0 69710.0 ;
      RECT  82020.0 71055.0 82725.0 72400.0 ;
      RECT  82020.0 73745.0 82725.0 72400.0 ;
      RECT  82020.0 73745.0 82725.0 75090.0 ;
      RECT  82020.0 76435.0 82725.0 75090.0 ;
      RECT  82020.0 76435.0 82725.0 77780.0 ;
      RECT  82020.0 79125.0 82725.0 77780.0 ;
      RECT  82020.0 79125.0 82725.0 80470.0 ;
      RECT  82020.0 81815.0 82725.0 80470.0 ;
      RECT  82020.0 81815.0 82725.0 83160.0 ;
      RECT  82020.0 84505.0 82725.0 83160.0 ;
      RECT  82020.0 84505.0 82725.0 85850.0 ;
      RECT  82020.0 87195.0 82725.0 85850.0 ;
      RECT  82020.0 87195.0 82725.0 88540.0 ;
      RECT  82020.0 89885.0 82725.0 88540.0 ;
      RECT  82020.0 89885.0 82725.0 91230.0 ;
      RECT  82020.0 92575.0 82725.0 91230.0 ;
      RECT  82020.0 92575.0 82725.0 93920.0 ;
      RECT  82020.0 95265.0 82725.0 93920.0 ;
      RECT  82020.0 95265.0 82725.0 96610.0 ;
      RECT  82020.0 97955.0 82725.0 96610.0 ;
      RECT  82020.0 97955.0 82725.0 99300.0 ;
      RECT  82020.0 100645.0 82725.0 99300.0 ;
      RECT  82020.0 100645.0 82725.0 101990.0 ;
      RECT  82020.0 103335.0 82725.0 101990.0 ;
      RECT  82020.0 103335.0 82725.0 104680.0 ;
      RECT  82020.0 106025.0 82725.0 104680.0 ;
      RECT  82020.0 106025.0 82725.0 107370.0 ;
      RECT  82020.0 108715.0 82725.0 107370.0 ;
      RECT  82020.0 108715.0 82725.0 110060.0 ;
      RECT  82020.0 111405.0 82725.0 110060.0 ;
      RECT  82020.0 111405.0 82725.0 112750.0 ;
      RECT  82020.0 114095.0 82725.0 112750.0 ;
      RECT  82725.0 28015.0 83430.0 29360.0 ;
      RECT  82725.0 30705.0 83430.0 29360.0 ;
      RECT  82725.0 30705.0 83430.0 32050.0 ;
      RECT  82725.0 33395.0 83430.0 32050.0 ;
      RECT  82725.0 33395.0 83430.0 34740.0 ;
      RECT  82725.0 36085.0 83430.0 34740.0 ;
      RECT  82725.0 36085.0 83430.0 37430.0 ;
      RECT  82725.0 38775.0 83430.0 37430.0 ;
      RECT  82725.0 38775.0 83430.0 40120.0 ;
      RECT  82725.0 41465.0 83430.0 40120.0 ;
      RECT  82725.0 41465.0 83430.0 42810.0 ;
      RECT  82725.0 44155.0 83430.0 42810.0 ;
      RECT  82725.0 44155.0 83430.0 45500.0 ;
      RECT  82725.0 46845.0 83430.0 45500.0 ;
      RECT  82725.0 46845.0 83430.0 48190.0 ;
      RECT  82725.0 49535.0 83430.0 48190.0 ;
      RECT  82725.0 49535.0 83430.0 50880.0 ;
      RECT  82725.0 52225.0 83430.0 50880.0 ;
      RECT  82725.0 52225.0 83430.0 53570.0 ;
      RECT  82725.0 54915.0 83430.0 53570.0 ;
      RECT  82725.0 54915.0 83430.0 56260.0 ;
      RECT  82725.0 57605.0 83430.0 56260.0 ;
      RECT  82725.0 57605.0 83430.0 58950.0 ;
      RECT  82725.0 60295.0 83430.0 58950.0 ;
      RECT  82725.0 60295.0 83430.0 61640.0 ;
      RECT  82725.0 62985.0 83430.0 61640.0 ;
      RECT  82725.0 62985.0 83430.0 64330.0 ;
      RECT  82725.0 65675.0 83430.0 64330.0 ;
      RECT  82725.0 65675.0 83430.0 67020.0 ;
      RECT  82725.0 68365.0 83430.0 67020.0 ;
      RECT  82725.0 68365.0 83430.0 69710.0 ;
      RECT  82725.0 71055.0 83430.0 69710.0 ;
      RECT  82725.0 71055.0 83430.0 72400.0 ;
      RECT  82725.0 73745.0 83430.0 72400.0 ;
      RECT  82725.0 73745.0 83430.0 75090.0 ;
      RECT  82725.0 76435.0 83430.0 75090.0 ;
      RECT  82725.0 76435.0 83430.0 77780.0 ;
      RECT  82725.0 79125.0 83430.0 77780.0 ;
      RECT  82725.0 79125.0 83430.0 80470.0 ;
      RECT  82725.0 81815.0 83430.0 80470.0 ;
      RECT  82725.0 81815.0 83430.0 83160.0 ;
      RECT  82725.0 84505.0 83430.0 83160.0 ;
      RECT  82725.0 84505.0 83430.0 85850.0 ;
      RECT  82725.0 87195.0 83430.0 85850.0 ;
      RECT  82725.0 87195.0 83430.0 88540.0 ;
      RECT  82725.0 89885.0 83430.0 88540.0 ;
      RECT  82725.0 89885.0 83430.0 91230.0 ;
      RECT  82725.0 92575.0 83430.0 91230.0 ;
      RECT  82725.0 92575.0 83430.0 93920.0 ;
      RECT  82725.0 95265.0 83430.0 93920.0 ;
      RECT  82725.0 95265.0 83430.0 96610.0 ;
      RECT  82725.0 97955.0 83430.0 96610.0 ;
      RECT  82725.0 97955.0 83430.0 99300.0 ;
      RECT  82725.0 100645.0 83430.0 99300.0 ;
      RECT  82725.0 100645.0 83430.0 101990.0 ;
      RECT  82725.0 103335.0 83430.0 101990.0 ;
      RECT  82725.0 103335.0 83430.0 104680.0 ;
      RECT  82725.0 106025.0 83430.0 104680.0 ;
      RECT  82725.0 106025.0 83430.0 107370.0 ;
      RECT  82725.0 108715.0 83430.0 107370.0 ;
      RECT  82725.0 108715.0 83430.0 110060.0 ;
      RECT  82725.0 111405.0 83430.0 110060.0 ;
      RECT  82725.0 111405.0 83430.0 112750.0 ;
      RECT  82725.0 114095.0 83430.0 112750.0 ;
      RECT  83430.0 28015.0 84135.0 29360.0 ;
      RECT  83430.0 30705.0 84135.0 29360.0 ;
      RECT  83430.0 30705.0 84135.0 32050.0 ;
      RECT  83430.0 33395.0 84135.0 32050.0 ;
      RECT  83430.0 33395.0 84135.0 34740.0 ;
      RECT  83430.0 36085.0 84135.0 34740.0 ;
      RECT  83430.0 36085.0 84135.0 37430.0 ;
      RECT  83430.0 38775.0 84135.0 37430.0 ;
      RECT  83430.0 38775.0 84135.0 40120.0 ;
      RECT  83430.0 41465.0 84135.0 40120.0 ;
      RECT  83430.0 41465.0 84135.0 42810.0 ;
      RECT  83430.0 44155.0 84135.0 42810.0 ;
      RECT  83430.0 44155.0 84135.0 45500.0 ;
      RECT  83430.0 46845.0 84135.0 45500.0 ;
      RECT  83430.0 46845.0 84135.0 48190.0 ;
      RECT  83430.0 49535.0 84135.0 48190.0 ;
      RECT  83430.0 49535.0 84135.0 50880.0 ;
      RECT  83430.0 52225.0 84135.0 50880.0 ;
      RECT  83430.0 52225.0 84135.0 53570.0 ;
      RECT  83430.0 54915.0 84135.0 53570.0 ;
      RECT  83430.0 54915.0 84135.0 56260.0 ;
      RECT  83430.0 57605.0 84135.0 56260.0 ;
      RECT  83430.0 57605.0 84135.0 58950.0 ;
      RECT  83430.0 60295.0 84135.0 58950.0 ;
      RECT  83430.0 60295.0 84135.0 61640.0 ;
      RECT  83430.0 62985.0 84135.0 61640.0 ;
      RECT  83430.0 62985.0 84135.0 64330.0 ;
      RECT  83430.0 65675.0 84135.0 64330.0 ;
      RECT  83430.0 65675.0 84135.0 67020.0 ;
      RECT  83430.0 68365.0 84135.0 67020.0 ;
      RECT  83430.0 68365.0 84135.0 69710.0 ;
      RECT  83430.0 71055.0 84135.0 69710.0 ;
      RECT  83430.0 71055.0 84135.0 72400.0 ;
      RECT  83430.0 73745.0 84135.0 72400.0 ;
      RECT  83430.0 73745.0 84135.0 75090.0 ;
      RECT  83430.0 76435.0 84135.0 75090.0 ;
      RECT  83430.0 76435.0 84135.0 77780.0 ;
      RECT  83430.0 79125.0 84135.0 77780.0 ;
      RECT  83430.0 79125.0 84135.0 80470.0 ;
      RECT  83430.0 81815.0 84135.0 80470.0 ;
      RECT  83430.0 81815.0 84135.0 83160.0 ;
      RECT  83430.0 84505.0 84135.0 83160.0 ;
      RECT  83430.0 84505.0 84135.0 85850.0 ;
      RECT  83430.0 87195.0 84135.0 85850.0 ;
      RECT  83430.0 87195.0 84135.0 88540.0 ;
      RECT  83430.0 89885.0 84135.0 88540.0 ;
      RECT  83430.0 89885.0 84135.0 91230.0 ;
      RECT  83430.0 92575.0 84135.0 91230.0 ;
      RECT  83430.0 92575.0 84135.0 93920.0 ;
      RECT  83430.0 95265.0 84135.0 93920.0 ;
      RECT  83430.0 95265.0 84135.0 96610.0 ;
      RECT  83430.0 97955.0 84135.0 96610.0 ;
      RECT  83430.0 97955.0 84135.0 99300.0 ;
      RECT  83430.0 100645.0 84135.0 99300.0 ;
      RECT  83430.0 100645.0 84135.0 101990.0 ;
      RECT  83430.0 103335.0 84135.0 101990.0 ;
      RECT  83430.0 103335.0 84135.0 104680.0 ;
      RECT  83430.0 106025.0 84135.0 104680.0 ;
      RECT  83430.0 106025.0 84135.0 107370.0 ;
      RECT  83430.0 108715.0 84135.0 107370.0 ;
      RECT  83430.0 108715.0 84135.0 110060.0 ;
      RECT  83430.0 111405.0 84135.0 110060.0 ;
      RECT  83430.0 111405.0 84135.0 112750.0 ;
      RECT  83430.0 114095.0 84135.0 112750.0 ;
      RECT  84135.0 28015.0 84840.0 29360.0 ;
      RECT  84135.0 30705.0 84840.0 29360.0 ;
      RECT  84135.0 30705.0 84840.0 32050.0 ;
      RECT  84135.0 33395.0 84840.0 32050.0 ;
      RECT  84135.0 33395.0 84840.0 34740.0 ;
      RECT  84135.0 36085.0 84840.0 34740.0 ;
      RECT  84135.0 36085.0 84840.0 37430.0 ;
      RECT  84135.0 38775.0 84840.0 37430.0 ;
      RECT  84135.0 38775.0 84840.0 40120.0 ;
      RECT  84135.0 41465.0 84840.0 40120.0 ;
      RECT  84135.0 41465.0 84840.0 42810.0 ;
      RECT  84135.0 44155.0 84840.0 42810.0 ;
      RECT  84135.0 44155.0 84840.0 45500.0 ;
      RECT  84135.0 46845.0 84840.0 45500.0 ;
      RECT  84135.0 46845.0 84840.0 48190.0 ;
      RECT  84135.0 49535.0 84840.0 48190.0 ;
      RECT  84135.0 49535.0 84840.0 50880.0 ;
      RECT  84135.0 52225.0 84840.0 50880.0 ;
      RECT  84135.0 52225.0 84840.0 53570.0 ;
      RECT  84135.0 54915.0 84840.0 53570.0 ;
      RECT  84135.0 54915.0 84840.0 56260.0 ;
      RECT  84135.0 57605.0 84840.0 56260.0 ;
      RECT  84135.0 57605.0 84840.0 58950.0 ;
      RECT  84135.0 60295.0 84840.0 58950.0 ;
      RECT  84135.0 60295.0 84840.0 61640.0 ;
      RECT  84135.0 62985.0 84840.0 61640.0 ;
      RECT  84135.0 62985.0 84840.0 64330.0 ;
      RECT  84135.0 65675.0 84840.0 64330.0 ;
      RECT  84135.0 65675.0 84840.0 67020.0 ;
      RECT  84135.0 68365.0 84840.0 67020.0 ;
      RECT  84135.0 68365.0 84840.0 69710.0 ;
      RECT  84135.0 71055.0 84840.0 69710.0 ;
      RECT  84135.0 71055.0 84840.0 72400.0 ;
      RECT  84135.0 73745.0 84840.0 72400.0 ;
      RECT  84135.0 73745.0 84840.0 75090.0 ;
      RECT  84135.0 76435.0 84840.0 75090.0 ;
      RECT  84135.0 76435.0 84840.0 77780.0 ;
      RECT  84135.0 79125.0 84840.0 77780.0 ;
      RECT  84135.0 79125.0 84840.0 80470.0 ;
      RECT  84135.0 81815.0 84840.0 80470.0 ;
      RECT  84135.0 81815.0 84840.0 83160.0 ;
      RECT  84135.0 84505.0 84840.0 83160.0 ;
      RECT  84135.0 84505.0 84840.0 85850.0 ;
      RECT  84135.0 87195.0 84840.0 85850.0 ;
      RECT  84135.0 87195.0 84840.0 88540.0 ;
      RECT  84135.0 89885.0 84840.0 88540.0 ;
      RECT  84135.0 89885.0 84840.0 91230.0 ;
      RECT  84135.0 92575.0 84840.0 91230.0 ;
      RECT  84135.0 92575.0 84840.0 93920.0 ;
      RECT  84135.0 95265.0 84840.0 93920.0 ;
      RECT  84135.0 95265.0 84840.0 96610.0 ;
      RECT  84135.0 97955.0 84840.0 96610.0 ;
      RECT  84135.0 97955.0 84840.0 99300.0 ;
      RECT  84135.0 100645.0 84840.0 99300.0 ;
      RECT  84135.0 100645.0 84840.0 101990.0 ;
      RECT  84135.0 103335.0 84840.0 101990.0 ;
      RECT  84135.0 103335.0 84840.0 104680.0 ;
      RECT  84135.0 106025.0 84840.0 104680.0 ;
      RECT  84135.0 106025.0 84840.0 107370.0 ;
      RECT  84135.0 108715.0 84840.0 107370.0 ;
      RECT  84135.0 108715.0 84840.0 110060.0 ;
      RECT  84135.0 111405.0 84840.0 110060.0 ;
      RECT  84135.0 111405.0 84840.0 112750.0 ;
      RECT  84135.0 114095.0 84840.0 112750.0 ;
      RECT  84840.0 28015.0 85545.0 29360.0 ;
      RECT  84840.0 30705.0 85545.0 29360.0 ;
      RECT  84840.0 30705.0 85545.0 32050.0 ;
      RECT  84840.0 33395.0 85545.0 32050.0 ;
      RECT  84840.0 33395.0 85545.0 34740.0 ;
      RECT  84840.0 36085.0 85545.0 34740.0 ;
      RECT  84840.0 36085.0 85545.0 37430.0 ;
      RECT  84840.0 38775.0 85545.0 37430.0 ;
      RECT  84840.0 38775.0 85545.0 40120.0 ;
      RECT  84840.0 41465.0 85545.0 40120.0 ;
      RECT  84840.0 41465.0 85545.0 42810.0 ;
      RECT  84840.0 44155.0 85545.0 42810.0 ;
      RECT  84840.0 44155.0 85545.0 45500.0 ;
      RECT  84840.0 46845.0 85545.0 45500.0 ;
      RECT  84840.0 46845.0 85545.0 48190.0 ;
      RECT  84840.0 49535.0 85545.0 48190.0 ;
      RECT  84840.0 49535.0 85545.0 50880.0 ;
      RECT  84840.0 52225.0 85545.0 50880.0 ;
      RECT  84840.0 52225.0 85545.0 53570.0 ;
      RECT  84840.0 54915.0 85545.0 53570.0 ;
      RECT  84840.0 54915.0 85545.0 56260.0 ;
      RECT  84840.0 57605.0 85545.0 56260.0 ;
      RECT  84840.0 57605.0 85545.0 58950.0 ;
      RECT  84840.0 60295.0 85545.0 58950.0 ;
      RECT  84840.0 60295.0 85545.0 61640.0 ;
      RECT  84840.0 62985.0 85545.0 61640.0 ;
      RECT  84840.0 62985.0 85545.0 64330.0 ;
      RECT  84840.0 65675.0 85545.0 64330.0 ;
      RECT  84840.0 65675.0 85545.0 67020.0 ;
      RECT  84840.0 68365.0 85545.0 67020.0 ;
      RECT  84840.0 68365.0 85545.0 69710.0 ;
      RECT  84840.0 71055.0 85545.0 69710.0 ;
      RECT  84840.0 71055.0 85545.0 72400.0 ;
      RECT  84840.0 73745.0 85545.0 72400.0 ;
      RECT  84840.0 73745.0 85545.0 75090.0 ;
      RECT  84840.0 76435.0 85545.0 75090.0 ;
      RECT  84840.0 76435.0 85545.0 77780.0 ;
      RECT  84840.0 79125.0 85545.0 77780.0 ;
      RECT  84840.0 79125.0 85545.0 80470.0 ;
      RECT  84840.0 81815.0 85545.0 80470.0 ;
      RECT  84840.0 81815.0 85545.0 83160.0 ;
      RECT  84840.0 84505.0 85545.0 83160.0 ;
      RECT  84840.0 84505.0 85545.0 85850.0 ;
      RECT  84840.0 87195.0 85545.0 85850.0 ;
      RECT  84840.0 87195.0 85545.0 88540.0 ;
      RECT  84840.0 89885.0 85545.0 88540.0 ;
      RECT  84840.0 89885.0 85545.0 91230.0 ;
      RECT  84840.0 92575.0 85545.0 91230.0 ;
      RECT  84840.0 92575.0 85545.0 93920.0 ;
      RECT  84840.0 95265.0 85545.0 93920.0 ;
      RECT  84840.0 95265.0 85545.0 96610.0 ;
      RECT  84840.0 97955.0 85545.0 96610.0 ;
      RECT  84840.0 97955.0 85545.0 99300.0 ;
      RECT  84840.0 100645.0 85545.0 99300.0 ;
      RECT  84840.0 100645.0 85545.0 101990.0 ;
      RECT  84840.0 103335.0 85545.0 101990.0 ;
      RECT  84840.0 103335.0 85545.0 104680.0 ;
      RECT  84840.0 106025.0 85545.0 104680.0 ;
      RECT  84840.0 106025.0 85545.0 107370.0 ;
      RECT  84840.0 108715.0 85545.0 107370.0 ;
      RECT  84840.0 108715.0 85545.0 110060.0 ;
      RECT  84840.0 111405.0 85545.0 110060.0 ;
      RECT  84840.0 111405.0 85545.0 112750.0 ;
      RECT  84840.0 114095.0 85545.0 112750.0 ;
      RECT  85545.0 28015.0 86250.0 29360.0 ;
      RECT  85545.0 30705.0 86250.0 29360.0 ;
      RECT  85545.0 30705.0 86250.0 32050.0 ;
      RECT  85545.0 33395.0 86250.0 32050.0 ;
      RECT  85545.0 33395.0 86250.0 34740.0 ;
      RECT  85545.0 36085.0 86250.0 34740.0 ;
      RECT  85545.0 36085.0 86250.0 37430.0 ;
      RECT  85545.0 38775.0 86250.0 37430.0 ;
      RECT  85545.0 38775.0 86250.0 40120.0 ;
      RECT  85545.0 41465.0 86250.0 40120.0 ;
      RECT  85545.0 41465.0 86250.0 42810.0 ;
      RECT  85545.0 44155.0 86250.0 42810.0 ;
      RECT  85545.0 44155.0 86250.0 45500.0 ;
      RECT  85545.0 46845.0 86250.0 45500.0 ;
      RECT  85545.0 46845.0 86250.0 48190.0 ;
      RECT  85545.0 49535.0 86250.0 48190.0 ;
      RECT  85545.0 49535.0 86250.0 50880.0 ;
      RECT  85545.0 52225.0 86250.0 50880.0 ;
      RECT  85545.0 52225.0 86250.0 53570.0 ;
      RECT  85545.0 54915.0 86250.0 53570.0 ;
      RECT  85545.0 54915.0 86250.0 56260.0 ;
      RECT  85545.0 57605.0 86250.0 56260.0 ;
      RECT  85545.0 57605.0 86250.0 58950.0 ;
      RECT  85545.0 60295.0 86250.0 58950.0 ;
      RECT  85545.0 60295.0 86250.0 61640.0 ;
      RECT  85545.0 62985.0 86250.0 61640.0 ;
      RECT  85545.0 62985.0 86250.0 64330.0 ;
      RECT  85545.0 65675.0 86250.0 64330.0 ;
      RECT  85545.0 65675.0 86250.0 67020.0 ;
      RECT  85545.0 68365.0 86250.0 67020.0 ;
      RECT  85545.0 68365.0 86250.0 69710.0 ;
      RECT  85545.0 71055.0 86250.0 69710.0 ;
      RECT  85545.0 71055.0 86250.0 72400.0 ;
      RECT  85545.0 73745.0 86250.0 72400.0 ;
      RECT  85545.0 73745.0 86250.0 75090.0 ;
      RECT  85545.0 76435.0 86250.0 75090.0 ;
      RECT  85545.0 76435.0 86250.0 77780.0 ;
      RECT  85545.0 79125.0 86250.0 77780.0 ;
      RECT  85545.0 79125.0 86250.0 80470.0 ;
      RECT  85545.0 81815.0 86250.0 80470.0 ;
      RECT  85545.0 81815.0 86250.0 83160.0 ;
      RECT  85545.0 84505.0 86250.0 83160.0 ;
      RECT  85545.0 84505.0 86250.0 85850.0 ;
      RECT  85545.0 87195.0 86250.0 85850.0 ;
      RECT  85545.0 87195.0 86250.0 88540.0 ;
      RECT  85545.0 89885.0 86250.0 88540.0 ;
      RECT  85545.0 89885.0 86250.0 91230.0 ;
      RECT  85545.0 92575.0 86250.0 91230.0 ;
      RECT  85545.0 92575.0 86250.0 93920.0 ;
      RECT  85545.0 95265.0 86250.0 93920.0 ;
      RECT  85545.0 95265.0 86250.0 96610.0 ;
      RECT  85545.0 97955.0 86250.0 96610.0 ;
      RECT  85545.0 97955.0 86250.0 99300.0 ;
      RECT  85545.0 100645.0 86250.0 99300.0 ;
      RECT  85545.0 100645.0 86250.0 101990.0 ;
      RECT  85545.0 103335.0 86250.0 101990.0 ;
      RECT  85545.0 103335.0 86250.0 104680.0 ;
      RECT  85545.0 106025.0 86250.0 104680.0 ;
      RECT  85545.0 106025.0 86250.0 107370.0 ;
      RECT  85545.0 108715.0 86250.0 107370.0 ;
      RECT  85545.0 108715.0 86250.0 110060.0 ;
      RECT  85545.0 111405.0 86250.0 110060.0 ;
      RECT  85545.0 111405.0 86250.0 112750.0 ;
      RECT  85545.0 114095.0 86250.0 112750.0 ;
      RECT  86250.0 28015.0 86955.0 29360.0 ;
      RECT  86250.0 30705.0 86955.0 29360.0 ;
      RECT  86250.0 30705.0 86955.0 32050.0 ;
      RECT  86250.0 33395.0 86955.0 32050.0 ;
      RECT  86250.0 33395.0 86955.0 34740.0 ;
      RECT  86250.0 36085.0 86955.0 34740.0 ;
      RECT  86250.0 36085.0 86955.0 37430.0 ;
      RECT  86250.0 38775.0 86955.0 37430.0 ;
      RECT  86250.0 38775.0 86955.0 40120.0 ;
      RECT  86250.0 41465.0 86955.0 40120.0 ;
      RECT  86250.0 41465.0 86955.0 42810.0 ;
      RECT  86250.0 44155.0 86955.0 42810.0 ;
      RECT  86250.0 44155.0 86955.0 45500.0 ;
      RECT  86250.0 46845.0 86955.0 45500.0 ;
      RECT  86250.0 46845.0 86955.0 48190.0 ;
      RECT  86250.0 49535.0 86955.0 48190.0 ;
      RECT  86250.0 49535.0 86955.0 50880.0 ;
      RECT  86250.0 52225.0 86955.0 50880.0 ;
      RECT  86250.0 52225.0 86955.0 53570.0 ;
      RECT  86250.0 54915.0 86955.0 53570.0 ;
      RECT  86250.0 54915.0 86955.0 56260.0 ;
      RECT  86250.0 57605.0 86955.0 56260.0 ;
      RECT  86250.0 57605.0 86955.0 58950.0 ;
      RECT  86250.0 60295.0 86955.0 58950.0 ;
      RECT  86250.0 60295.0 86955.0 61640.0 ;
      RECT  86250.0 62985.0 86955.0 61640.0 ;
      RECT  86250.0 62985.0 86955.0 64330.0 ;
      RECT  86250.0 65675.0 86955.0 64330.0 ;
      RECT  86250.0 65675.0 86955.0 67020.0 ;
      RECT  86250.0 68365.0 86955.0 67020.0 ;
      RECT  86250.0 68365.0 86955.0 69710.0 ;
      RECT  86250.0 71055.0 86955.0 69710.0 ;
      RECT  86250.0 71055.0 86955.0 72400.0 ;
      RECT  86250.0 73745.0 86955.0 72400.0 ;
      RECT  86250.0 73745.0 86955.0 75090.0 ;
      RECT  86250.0 76435.0 86955.0 75090.0 ;
      RECT  86250.0 76435.0 86955.0 77780.0 ;
      RECT  86250.0 79125.0 86955.0 77780.0 ;
      RECT  86250.0 79125.0 86955.0 80470.0 ;
      RECT  86250.0 81815.0 86955.0 80470.0 ;
      RECT  86250.0 81815.0 86955.0 83160.0 ;
      RECT  86250.0 84505.0 86955.0 83160.0 ;
      RECT  86250.0 84505.0 86955.0 85850.0 ;
      RECT  86250.0 87195.0 86955.0 85850.0 ;
      RECT  86250.0 87195.0 86955.0 88540.0 ;
      RECT  86250.0 89885.0 86955.0 88540.0 ;
      RECT  86250.0 89885.0 86955.0 91230.0 ;
      RECT  86250.0 92575.0 86955.0 91230.0 ;
      RECT  86250.0 92575.0 86955.0 93920.0 ;
      RECT  86250.0 95265.0 86955.0 93920.0 ;
      RECT  86250.0 95265.0 86955.0 96610.0 ;
      RECT  86250.0 97955.0 86955.0 96610.0 ;
      RECT  86250.0 97955.0 86955.0 99300.0 ;
      RECT  86250.0 100645.0 86955.0 99300.0 ;
      RECT  86250.0 100645.0 86955.0 101990.0 ;
      RECT  86250.0 103335.0 86955.0 101990.0 ;
      RECT  86250.0 103335.0 86955.0 104680.0 ;
      RECT  86250.0 106025.0 86955.0 104680.0 ;
      RECT  86250.0 106025.0 86955.0 107370.0 ;
      RECT  86250.0 108715.0 86955.0 107370.0 ;
      RECT  86250.0 108715.0 86955.0 110060.0 ;
      RECT  86250.0 111405.0 86955.0 110060.0 ;
      RECT  86250.0 111405.0 86955.0 112750.0 ;
      RECT  86250.0 114095.0 86955.0 112750.0 ;
      RECT  86955.0 28015.0 87660.0 29360.0 ;
      RECT  86955.0 30705.0 87660.0 29360.0 ;
      RECT  86955.0 30705.0 87660.0 32050.0 ;
      RECT  86955.0 33395.0 87660.0 32050.0 ;
      RECT  86955.0 33395.0 87660.0 34740.0 ;
      RECT  86955.0 36085.0 87660.0 34740.0 ;
      RECT  86955.0 36085.0 87660.0 37430.0 ;
      RECT  86955.0 38775.0 87660.0 37430.0 ;
      RECT  86955.0 38775.0 87660.0 40120.0 ;
      RECT  86955.0 41465.0 87660.0 40120.0 ;
      RECT  86955.0 41465.0 87660.0 42810.0 ;
      RECT  86955.0 44155.0 87660.0 42810.0 ;
      RECT  86955.0 44155.0 87660.0 45500.0 ;
      RECT  86955.0 46845.0 87660.0 45500.0 ;
      RECT  86955.0 46845.0 87660.0 48190.0 ;
      RECT  86955.0 49535.0 87660.0 48190.0 ;
      RECT  86955.0 49535.0 87660.0 50880.0 ;
      RECT  86955.0 52225.0 87660.0 50880.0 ;
      RECT  86955.0 52225.0 87660.0 53570.0 ;
      RECT  86955.0 54915.0 87660.0 53570.0 ;
      RECT  86955.0 54915.0 87660.0 56260.0 ;
      RECT  86955.0 57605.0 87660.0 56260.0 ;
      RECT  86955.0 57605.0 87660.0 58950.0 ;
      RECT  86955.0 60295.0 87660.0 58950.0 ;
      RECT  86955.0 60295.0 87660.0 61640.0 ;
      RECT  86955.0 62985.0 87660.0 61640.0 ;
      RECT  86955.0 62985.0 87660.0 64330.0 ;
      RECT  86955.0 65675.0 87660.0 64330.0 ;
      RECT  86955.0 65675.0 87660.0 67020.0 ;
      RECT  86955.0 68365.0 87660.0 67020.0 ;
      RECT  86955.0 68365.0 87660.0 69710.0 ;
      RECT  86955.0 71055.0 87660.0 69710.0 ;
      RECT  86955.0 71055.0 87660.0 72400.0 ;
      RECT  86955.0 73745.0 87660.0 72400.0 ;
      RECT  86955.0 73745.0 87660.0 75090.0 ;
      RECT  86955.0 76435.0 87660.0 75090.0 ;
      RECT  86955.0 76435.0 87660.0 77780.0 ;
      RECT  86955.0 79125.0 87660.0 77780.0 ;
      RECT  86955.0 79125.0 87660.0 80470.0 ;
      RECT  86955.0 81815.0 87660.0 80470.0 ;
      RECT  86955.0 81815.0 87660.0 83160.0 ;
      RECT  86955.0 84505.0 87660.0 83160.0 ;
      RECT  86955.0 84505.0 87660.0 85850.0 ;
      RECT  86955.0 87195.0 87660.0 85850.0 ;
      RECT  86955.0 87195.0 87660.0 88540.0 ;
      RECT  86955.0 89885.0 87660.0 88540.0 ;
      RECT  86955.0 89885.0 87660.0 91230.0 ;
      RECT  86955.0 92575.0 87660.0 91230.0 ;
      RECT  86955.0 92575.0 87660.0 93920.0 ;
      RECT  86955.0 95265.0 87660.0 93920.0 ;
      RECT  86955.0 95265.0 87660.0 96610.0 ;
      RECT  86955.0 97955.0 87660.0 96610.0 ;
      RECT  86955.0 97955.0 87660.0 99300.0 ;
      RECT  86955.0 100645.0 87660.0 99300.0 ;
      RECT  86955.0 100645.0 87660.0 101990.0 ;
      RECT  86955.0 103335.0 87660.0 101990.0 ;
      RECT  86955.0 103335.0 87660.0 104680.0 ;
      RECT  86955.0 106025.0 87660.0 104680.0 ;
      RECT  86955.0 106025.0 87660.0 107370.0 ;
      RECT  86955.0 108715.0 87660.0 107370.0 ;
      RECT  86955.0 108715.0 87660.0 110060.0 ;
      RECT  86955.0 111405.0 87660.0 110060.0 ;
      RECT  86955.0 111405.0 87660.0 112750.0 ;
      RECT  86955.0 114095.0 87660.0 112750.0 ;
      RECT  87660.0 28015.0 88365.0 29360.0 ;
      RECT  87660.0 30705.0 88365.0 29360.0 ;
      RECT  87660.0 30705.0 88365.0 32050.0 ;
      RECT  87660.0 33395.0 88365.0 32050.0 ;
      RECT  87660.0 33395.0 88365.0 34740.0 ;
      RECT  87660.0 36085.0 88365.0 34740.0 ;
      RECT  87660.0 36085.0 88365.0 37430.0 ;
      RECT  87660.0 38775.0 88365.0 37430.0 ;
      RECT  87660.0 38775.0 88365.0 40120.0 ;
      RECT  87660.0 41465.0 88365.0 40120.0 ;
      RECT  87660.0 41465.0 88365.0 42810.0 ;
      RECT  87660.0 44155.0 88365.0 42810.0 ;
      RECT  87660.0 44155.0 88365.0 45500.0 ;
      RECT  87660.0 46845.0 88365.0 45500.0 ;
      RECT  87660.0 46845.0 88365.0 48190.0 ;
      RECT  87660.0 49535.0 88365.0 48190.0 ;
      RECT  87660.0 49535.0 88365.0 50880.0 ;
      RECT  87660.0 52225.0 88365.0 50880.0 ;
      RECT  87660.0 52225.0 88365.0 53570.0 ;
      RECT  87660.0 54915.0 88365.0 53570.0 ;
      RECT  87660.0 54915.0 88365.0 56260.0 ;
      RECT  87660.0 57605.0 88365.0 56260.0 ;
      RECT  87660.0 57605.0 88365.0 58950.0 ;
      RECT  87660.0 60295.0 88365.0 58950.0 ;
      RECT  87660.0 60295.0 88365.0 61640.0 ;
      RECT  87660.0 62985.0 88365.0 61640.0 ;
      RECT  87660.0 62985.0 88365.0 64330.0 ;
      RECT  87660.0 65675.0 88365.0 64330.0 ;
      RECT  87660.0 65675.0 88365.0 67020.0 ;
      RECT  87660.0 68365.0 88365.0 67020.0 ;
      RECT  87660.0 68365.0 88365.0 69710.0 ;
      RECT  87660.0 71055.0 88365.0 69710.0 ;
      RECT  87660.0 71055.0 88365.0 72400.0 ;
      RECT  87660.0 73745.0 88365.0 72400.0 ;
      RECT  87660.0 73745.0 88365.0 75090.0 ;
      RECT  87660.0 76435.0 88365.0 75090.0 ;
      RECT  87660.0 76435.0 88365.0 77780.0 ;
      RECT  87660.0 79125.0 88365.0 77780.0 ;
      RECT  87660.0 79125.0 88365.0 80470.0 ;
      RECT  87660.0 81815.0 88365.0 80470.0 ;
      RECT  87660.0 81815.0 88365.0 83160.0 ;
      RECT  87660.0 84505.0 88365.0 83160.0 ;
      RECT  87660.0 84505.0 88365.0 85850.0 ;
      RECT  87660.0 87195.0 88365.0 85850.0 ;
      RECT  87660.0 87195.0 88365.0 88540.0 ;
      RECT  87660.0 89885.0 88365.0 88540.0 ;
      RECT  87660.0 89885.0 88365.0 91230.0 ;
      RECT  87660.0 92575.0 88365.0 91230.0 ;
      RECT  87660.0 92575.0 88365.0 93920.0 ;
      RECT  87660.0 95265.0 88365.0 93920.0 ;
      RECT  87660.0 95265.0 88365.0 96610.0 ;
      RECT  87660.0 97955.0 88365.0 96610.0 ;
      RECT  87660.0 97955.0 88365.0 99300.0 ;
      RECT  87660.0 100645.0 88365.0 99300.0 ;
      RECT  87660.0 100645.0 88365.0 101990.0 ;
      RECT  87660.0 103335.0 88365.0 101990.0 ;
      RECT  87660.0 103335.0 88365.0 104680.0 ;
      RECT  87660.0 106025.0 88365.0 104680.0 ;
      RECT  87660.0 106025.0 88365.0 107370.0 ;
      RECT  87660.0 108715.0 88365.0 107370.0 ;
      RECT  87660.0 108715.0 88365.0 110060.0 ;
      RECT  87660.0 111405.0 88365.0 110060.0 ;
      RECT  87660.0 111405.0 88365.0 112750.0 ;
      RECT  87660.0 114095.0 88365.0 112750.0 ;
      RECT  88365.0 28015.0 89070.0 29360.0 ;
      RECT  88365.0 30705.0 89070.0 29360.0 ;
      RECT  88365.0 30705.0 89070.0 32050.0 ;
      RECT  88365.0 33395.0 89070.0 32050.0 ;
      RECT  88365.0 33395.0 89070.0 34740.0 ;
      RECT  88365.0 36085.0 89070.0 34740.0 ;
      RECT  88365.0 36085.0 89070.0 37430.0 ;
      RECT  88365.0 38775.0 89070.0 37430.0 ;
      RECT  88365.0 38775.0 89070.0 40120.0 ;
      RECT  88365.0 41465.0 89070.0 40120.0 ;
      RECT  88365.0 41465.0 89070.0 42810.0 ;
      RECT  88365.0 44155.0 89070.0 42810.0 ;
      RECT  88365.0 44155.0 89070.0 45500.0 ;
      RECT  88365.0 46845.0 89070.0 45500.0 ;
      RECT  88365.0 46845.0 89070.0 48190.0 ;
      RECT  88365.0 49535.0 89070.0 48190.0 ;
      RECT  88365.0 49535.0 89070.0 50880.0 ;
      RECT  88365.0 52225.0 89070.0 50880.0 ;
      RECT  88365.0 52225.0 89070.0 53570.0 ;
      RECT  88365.0 54915.0 89070.0 53570.0 ;
      RECT  88365.0 54915.0 89070.0 56260.0 ;
      RECT  88365.0 57605.0 89070.0 56260.0 ;
      RECT  88365.0 57605.0 89070.0 58950.0 ;
      RECT  88365.0 60295.0 89070.0 58950.0 ;
      RECT  88365.0 60295.0 89070.0 61640.0 ;
      RECT  88365.0 62985.0 89070.0 61640.0 ;
      RECT  88365.0 62985.0 89070.0 64330.0 ;
      RECT  88365.0 65675.0 89070.0 64330.0 ;
      RECT  88365.0 65675.0 89070.0 67020.0 ;
      RECT  88365.0 68365.0 89070.0 67020.0 ;
      RECT  88365.0 68365.0 89070.0 69710.0 ;
      RECT  88365.0 71055.0 89070.0 69710.0 ;
      RECT  88365.0 71055.0 89070.0 72400.0 ;
      RECT  88365.0 73745.0 89070.0 72400.0 ;
      RECT  88365.0 73745.0 89070.0 75090.0 ;
      RECT  88365.0 76435.0 89070.0 75090.0 ;
      RECT  88365.0 76435.0 89070.0 77780.0 ;
      RECT  88365.0 79125.0 89070.0 77780.0 ;
      RECT  88365.0 79125.0 89070.0 80470.0 ;
      RECT  88365.0 81815.0 89070.0 80470.0 ;
      RECT  88365.0 81815.0 89070.0 83160.0 ;
      RECT  88365.0 84505.0 89070.0 83160.0 ;
      RECT  88365.0 84505.0 89070.0 85850.0 ;
      RECT  88365.0 87195.0 89070.0 85850.0 ;
      RECT  88365.0 87195.0 89070.0 88540.0 ;
      RECT  88365.0 89885.0 89070.0 88540.0 ;
      RECT  88365.0 89885.0 89070.0 91230.0 ;
      RECT  88365.0 92575.0 89070.0 91230.0 ;
      RECT  88365.0 92575.0 89070.0 93920.0 ;
      RECT  88365.0 95265.0 89070.0 93920.0 ;
      RECT  88365.0 95265.0 89070.0 96610.0 ;
      RECT  88365.0 97955.0 89070.0 96610.0 ;
      RECT  88365.0 97955.0 89070.0 99300.0 ;
      RECT  88365.0 100645.0 89070.0 99300.0 ;
      RECT  88365.0 100645.0 89070.0 101990.0 ;
      RECT  88365.0 103335.0 89070.0 101990.0 ;
      RECT  88365.0 103335.0 89070.0 104680.0 ;
      RECT  88365.0 106025.0 89070.0 104680.0 ;
      RECT  88365.0 106025.0 89070.0 107370.0 ;
      RECT  88365.0 108715.0 89070.0 107370.0 ;
      RECT  88365.0 108715.0 89070.0 110060.0 ;
      RECT  88365.0 111405.0 89070.0 110060.0 ;
      RECT  88365.0 111405.0 89070.0 112750.0 ;
      RECT  88365.0 114095.0 89070.0 112750.0 ;
      RECT  89070.0 28015.0 89775.0 29360.0 ;
      RECT  89070.0 30705.0 89775.0 29360.0 ;
      RECT  89070.0 30705.0 89775.0 32050.0 ;
      RECT  89070.0 33395.0 89775.0 32050.0 ;
      RECT  89070.0 33395.0 89775.0 34740.0 ;
      RECT  89070.0 36085.0 89775.0 34740.0 ;
      RECT  89070.0 36085.0 89775.0 37430.0 ;
      RECT  89070.0 38775.0 89775.0 37430.0 ;
      RECT  89070.0 38775.0 89775.0 40120.0 ;
      RECT  89070.0 41465.0 89775.0 40120.0 ;
      RECT  89070.0 41465.0 89775.0 42810.0 ;
      RECT  89070.0 44155.0 89775.0 42810.0 ;
      RECT  89070.0 44155.0 89775.0 45500.0 ;
      RECT  89070.0 46845.0 89775.0 45500.0 ;
      RECT  89070.0 46845.0 89775.0 48190.0 ;
      RECT  89070.0 49535.0 89775.0 48190.0 ;
      RECT  89070.0 49535.0 89775.0 50880.0 ;
      RECT  89070.0 52225.0 89775.0 50880.0 ;
      RECT  89070.0 52225.0 89775.0 53570.0 ;
      RECT  89070.0 54915.0 89775.0 53570.0 ;
      RECT  89070.0 54915.0 89775.0 56260.0 ;
      RECT  89070.0 57605.0 89775.0 56260.0 ;
      RECT  89070.0 57605.0 89775.0 58950.0 ;
      RECT  89070.0 60295.0 89775.0 58950.0 ;
      RECT  89070.0 60295.0 89775.0 61640.0 ;
      RECT  89070.0 62985.0 89775.0 61640.0 ;
      RECT  89070.0 62985.0 89775.0 64330.0 ;
      RECT  89070.0 65675.0 89775.0 64330.0 ;
      RECT  89070.0 65675.0 89775.0 67020.0 ;
      RECT  89070.0 68365.0 89775.0 67020.0 ;
      RECT  89070.0 68365.0 89775.0 69710.0 ;
      RECT  89070.0 71055.0 89775.0 69710.0 ;
      RECT  89070.0 71055.0 89775.0 72400.0 ;
      RECT  89070.0 73745.0 89775.0 72400.0 ;
      RECT  89070.0 73745.0 89775.0 75090.0 ;
      RECT  89070.0 76435.0 89775.0 75090.0 ;
      RECT  89070.0 76435.0 89775.0 77780.0 ;
      RECT  89070.0 79125.0 89775.0 77780.0 ;
      RECT  89070.0 79125.0 89775.0 80470.0 ;
      RECT  89070.0 81815.0 89775.0 80470.0 ;
      RECT  89070.0 81815.0 89775.0 83160.0 ;
      RECT  89070.0 84505.0 89775.0 83160.0 ;
      RECT  89070.0 84505.0 89775.0 85850.0 ;
      RECT  89070.0 87195.0 89775.0 85850.0 ;
      RECT  89070.0 87195.0 89775.0 88540.0 ;
      RECT  89070.0 89885.0 89775.0 88540.0 ;
      RECT  89070.0 89885.0 89775.0 91230.0 ;
      RECT  89070.0 92575.0 89775.0 91230.0 ;
      RECT  89070.0 92575.0 89775.0 93920.0 ;
      RECT  89070.0 95265.0 89775.0 93920.0 ;
      RECT  89070.0 95265.0 89775.0 96610.0 ;
      RECT  89070.0 97955.0 89775.0 96610.0 ;
      RECT  89070.0 97955.0 89775.0 99300.0 ;
      RECT  89070.0 100645.0 89775.0 99300.0 ;
      RECT  89070.0 100645.0 89775.0 101990.0 ;
      RECT  89070.0 103335.0 89775.0 101990.0 ;
      RECT  89070.0 103335.0 89775.0 104680.0 ;
      RECT  89070.0 106025.0 89775.0 104680.0 ;
      RECT  89070.0 106025.0 89775.0 107370.0 ;
      RECT  89070.0 108715.0 89775.0 107370.0 ;
      RECT  89070.0 108715.0 89775.0 110060.0 ;
      RECT  89070.0 111405.0 89775.0 110060.0 ;
      RECT  89070.0 111405.0 89775.0 112750.0 ;
      RECT  89070.0 114095.0 89775.0 112750.0 ;
      RECT  89775.0 28015.0 90480.0 29360.0 ;
      RECT  89775.0 30705.0 90480.0 29360.0 ;
      RECT  89775.0 30705.0 90480.0 32050.0 ;
      RECT  89775.0 33395.0 90480.0 32050.0 ;
      RECT  89775.0 33395.0 90480.0 34740.0 ;
      RECT  89775.0 36085.0 90480.0 34740.0 ;
      RECT  89775.0 36085.0 90480.0 37430.0 ;
      RECT  89775.0 38775.0 90480.0 37430.0 ;
      RECT  89775.0 38775.0 90480.0 40120.0 ;
      RECT  89775.0 41465.0 90480.0 40120.0 ;
      RECT  89775.0 41465.0 90480.0 42810.0 ;
      RECT  89775.0 44155.0 90480.0 42810.0 ;
      RECT  89775.0 44155.0 90480.0 45500.0 ;
      RECT  89775.0 46845.0 90480.0 45500.0 ;
      RECT  89775.0 46845.0 90480.0 48190.0 ;
      RECT  89775.0 49535.0 90480.0 48190.0 ;
      RECT  89775.0 49535.0 90480.0 50880.0 ;
      RECT  89775.0 52225.0 90480.0 50880.0 ;
      RECT  89775.0 52225.0 90480.0 53570.0 ;
      RECT  89775.0 54915.0 90480.0 53570.0 ;
      RECT  89775.0 54915.0 90480.0 56260.0 ;
      RECT  89775.0 57605.0 90480.0 56260.0 ;
      RECT  89775.0 57605.0 90480.0 58950.0 ;
      RECT  89775.0 60295.0 90480.0 58950.0 ;
      RECT  89775.0 60295.0 90480.0 61640.0 ;
      RECT  89775.0 62985.0 90480.0 61640.0 ;
      RECT  89775.0 62985.0 90480.0 64330.0 ;
      RECT  89775.0 65675.0 90480.0 64330.0 ;
      RECT  89775.0 65675.0 90480.0 67020.0 ;
      RECT  89775.0 68365.0 90480.0 67020.0 ;
      RECT  89775.0 68365.0 90480.0 69710.0 ;
      RECT  89775.0 71055.0 90480.0 69710.0 ;
      RECT  89775.0 71055.0 90480.0 72400.0 ;
      RECT  89775.0 73745.0 90480.0 72400.0 ;
      RECT  89775.0 73745.0 90480.0 75090.0 ;
      RECT  89775.0 76435.0 90480.0 75090.0 ;
      RECT  89775.0 76435.0 90480.0 77780.0 ;
      RECT  89775.0 79125.0 90480.0 77780.0 ;
      RECT  89775.0 79125.0 90480.0 80470.0 ;
      RECT  89775.0 81815.0 90480.0 80470.0 ;
      RECT  89775.0 81815.0 90480.0 83160.0 ;
      RECT  89775.0 84505.0 90480.0 83160.0 ;
      RECT  89775.0 84505.0 90480.0 85850.0 ;
      RECT  89775.0 87195.0 90480.0 85850.0 ;
      RECT  89775.0 87195.0 90480.0 88540.0 ;
      RECT  89775.0 89885.0 90480.0 88540.0 ;
      RECT  89775.0 89885.0 90480.0 91230.0 ;
      RECT  89775.0 92575.0 90480.0 91230.0 ;
      RECT  89775.0 92575.0 90480.0 93920.0 ;
      RECT  89775.0 95265.0 90480.0 93920.0 ;
      RECT  89775.0 95265.0 90480.0 96610.0 ;
      RECT  89775.0 97955.0 90480.0 96610.0 ;
      RECT  89775.0 97955.0 90480.0 99300.0 ;
      RECT  89775.0 100645.0 90480.0 99300.0 ;
      RECT  89775.0 100645.0 90480.0 101990.0 ;
      RECT  89775.0 103335.0 90480.0 101990.0 ;
      RECT  89775.0 103335.0 90480.0 104680.0 ;
      RECT  89775.0 106025.0 90480.0 104680.0 ;
      RECT  89775.0 106025.0 90480.0 107370.0 ;
      RECT  89775.0 108715.0 90480.0 107370.0 ;
      RECT  89775.0 108715.0 90480.0 110060.0 ;
      RECT  89775.0 111405.0 90480.0 110060.0 ;
      RECT  89775.0 111405.0 90480.0 112750.0 ;
      RECT  89775.0 114095.0 90480.0 112750.0 ;
      RECT  90480.0 28015.0 91185.0 29360.0 ;
      RECT  90480.0 30705.0 91185.0 29360.0 ;
      RECT  90480.0 30705.0 91185.0 32050.0 ;
      RECT  90480.0 33395.0 91185.0 32050.0 ;
      RECT  90480.0 33395.0 91185.0 34740.0 ;
      RECT  90480.0 36085.0 91185.0 34740.0 ;
      RECT  90480.0 36085.0 91185.0 37430.0 ;
      RECT  90480.0 38775.0 91185.0 37430.0 ;
      RECT  90480.0 38775.0 91185.0 40120.0 ;
      RECT  90480.0 41465.0 91185.0 40120.0 ;
      RECT  90480.0 41465.0 91185.0 42810.0 ;
      RECT  90480.0 44155.0 91185.0 42810.0 ;
      RECT  90480.0 44155.0 91185.0 45500.0 ;
      RECT  90480.0 46845.0 91185.0 45500.0 ;
      RECT  90480.0 46845.0 91185.0 48190.0 ;
      RECT  90480.0 49535.0 91185.0 48190.0 ;
      RECT  90480.0 49535.0 91185.0 50880.0 ;
      RECT  90480.0 52225.0 91185.0 50880.0 ;
      RECT  90480.0 52225.0 91185.0 53570.0 ;
      RECT  90480.0 54915.0 91185.0 53570.0 ;
      RECT  90480.0 54915.0 91185.0 56260.0 ;
      RECT  90480.0 57605.0 91185.0 56260.0 ;
      RECT  90480.0 57605.0 91185.0 58950.0 ;
      RECT  90480.0 60295.0 91185.0 58950.0 ;
      RECT  90480.0 60295.0 91185.0 61640.0 ;
      RECT  90480.0 62985.0 91185.0 61640.0 ;
      RECT  90480.0 62985.0 91185.0 64330.0 ;
      RECT  90480.0 65675.0 91185.0 64330.0 ;
      RECT  90480.0 65675.0 91185.0 67020.0 ;
      RECT  90480.0 68365.0 91185.0 67020.0 ;
      RECT  90480.0 68365.0 91185.0 69710.0 ;
      RECT  90480.0 71055.0 91185.0 69710.0 ;
      RECT  90480.0 71055.0 91185.0 72400.0 ;
      RECT  90480.0 73745.0 91185.0 72400.0 ;
      RECT  90480.0 73745.0 91185.0 75090.0 ;
      RECT  90480.0 76435.0 91185.0 75090.0 ;
      RECT  90480.0 76435.0 91185.0 77780.0 ;
      RECT  90480.0 79125.0 91185.0 77780.0 ;
      RECT  90480.0 79125.0 91185.0 80470.0 ;
      RECT  90480.0 81815.0 91185.0 80470.0 ;
      RECT  90480.0 81815.0 91185.0 83160.0 ;
      RECT  90480.0 84505.0 91185.0 83160.0 ;
      RECT  90480.0 84505.0 91185.0 85850.0 ;
      RECT  90480.0 87195.0 91185.0 85850.0 ;
      RECT  90480.0 87195.0 91185.0 88540.0 ;
      RECT  90480.0 89885.0 91185.0 88540.0 ;
      RECT  90480.0 89885.0 91185.0 91230.0 ;
      RECT  90480.0 92575.0 91185.0 91230.0 ;
      RECT  90480.0 92575.0 91185.0 93920.0 ;
      RECT  90480.0 95265.0 91185.0 93920.0 ;
      RECT  90480.0 95265.0 91185.0 96610.0 ;
      RECT  90480.0 97955.0 91185.0 96610.0 ;
      RECT  90480.0 97955.0 91185.0 99300.0 ;
      RECT  90480.0 100645.0 91185.0 99300.0 ;
      RECT  90480.0 100645.0 91185.0 101990.0 ;
      RECT  90480.0 103335.0 91185.0 101990.0 ;
      RECT  90480.0 103335.0 91185.0 104680.0 ;
      RECT  90480.0 106025.0 91185.0 104680.0 ;
      RECT  90480.0 106025.0 91185.0 107370.0 ;
      RECT  90480.0 108715.0 91185.0 107370.0 ;
      RECT  90480.0 108715.0 91185.0 110060.0 ;
      RECT  90480.0 111405.0 91185.0 110060.0 ;
      RECT  90480.0 111405.0 91185.0 112750.0 ;
      RECT  90480.0 114095.0 91185.0 112750.0 ;
      RECT  91185.0 28015.0 91890.0 29360.0 ;
      RECT  91185.0 30705.0 91890.0 29360.0 ;
      RECT  91185.0 30705.0 91890.0 32050.0 ;
      RECT  91185.0 33395.0 91890.0 32050.0 ;
      RECT  91185.0 33395.0 91890.0 34740.0 ;
      RECT  91185.0 36085.0 91890.0 34740.0 ;
      RECT  91185.0 36085.0 91890.0 37430.0 ;
      RECT  91185.0 38775.0 91890.0 37430.0 ;
      RECT  91185.0 38775.0 91890.0 40120.0 ;
      RECT  91185.0 41465.0 91890.0 40120.0 ;
      RECT  91185.0 41465.0 91890.0 42810.0 ;
      RECT  91185.0 44155.0 91890.0 42810.0 ;
      RECT  91185.0 44155.0 91890.0 45500.0 ;
      RECT  91185.0 46845.0 91890.0 45500.0 ;
      RECT  91185.0 46845.0 91890.0 48190.0 ;
      RECT  91185.0 49535.0 91890.0 48190.0 ;
      RECT  91185.0 49535.0 91890.0 50880.0 ;
      RECT  91185.0 52225.0 91890.0 50880.0 ;
      RECT  91185.0 52225.0 91890.0 53570.0 ;
      RECT  91185.0 54915.0 91890.0 53570.0 ;
      RECT  91185.0 54915.0 91890.0 56260.0 ;
      RECT  91185.0 57605.0 91890.0 56260.0 ;
      RECT  91185.0 57605.0 91890.0 58950.0 ;
      RECT  91185.0 60295.0 91890.0 58950.0 ;
      RECT  91185.0 60295.0 91890.0 61640.0 ;
      RECT  91185.0 62985.0 91890.0 61640.0 ;
      RECT  91185.0 62985.0 91890.0 64330.0 ;
      RECT  91185.0 65675.0 91890.0 64330.0 ;
      RECT  91185.0 65675.0 91890.0 67020.0 ;
      RECT  91185.0 68365.0 91890.0 67020.0 ;
      RECT  91185.0 68365.0 91890.0 69710.0 ;
      RECT  91185.0 71055.0 91890.0 69710.0 ;
      RECT  91185.0 71055.0 91890.0 72400.0 ;
      RECT  91185.0 73745.0 91890.0 72400.0 ;
      RECT  91185.0 73745.0 91890.0 75090.0 ;
      RECT  91185.0 76435.0 91890.0 75090.0 ;
      RECT  91185.0 76435.0 91890.0 77780.0 ;
      RECT  91185.0 79125.0 91890.0 77780.0 ;
      RECT  91185.0 79125.0 91890.0 80470.0 ;
      RECT  91185.0 81815.0 91890.0 80470.0 ;
      RECT  91185.0 81815.0 91890.0 83160.0 ;
      RECT  91185.0 84505.0 91890.0 83160.0 ;
      RECT  91185.0 84505.0 91890.0 85850.0 ;
      RECT  91185.0 87195.0 91890.0 85850.0 ;
      RECT  91185.0 87195.0 91890.0 88540.0 ;
      RECT  91185.0 89885.0 91890.0 88540.0 ;
      RECT  91185.0 89885.0 91890.0 91230.0 ;
      RECT  91185.0 92575.0 91890.0 91230.0 ;
      RECT  91185.0 92575.0 91890.0 93920.0 ;
      RECT  91185.0 95265.0 91890.0 93920.0 ;
      RECT  91185.0 95265.0 91890.0 96610.0 ;
      RECT  91185.0 97955.0 91890.0 96610.0 ;
      RECT  91185.0 97955.0 91890.0 99300.0 ;
      RECT  91185.0 100645.0 91890.0 99300.0 ;
      RECT  91185.0 100645.0 91890.0 101990.0 ;
      RECT  91185.0 103335.0 91890.0 101990.0 ;
      RECT  91185.0 103335.0 91890.0 104680.0 ;
      RECT  91185.0 106025.0 91890.0 104680.0 ;
      RECT  91185.0 106025.0 91890.0 107370.0 ;
      RECT  91185.0 108715.0 91890.0 107370.0 ;
      RECT  91185.0 108715.0 91890.0 110060.0 ;
      RECT  91185.0 111405.0 91890.0 110060.0 ;
      RECT  91185.0 111405.0 91890.0 112750.0 ;
      RECT  91185.0 114095.0 91890.0 112750.0 ;
      RECT  91890.0 28015.0 92595.0 29360.0 ;
      RECT  91890.0 30705.0 92595.0 29360.0 ;
      RECT  91890.0 30705.0 92595.0 32050.0 ;
      RECT  91890.0 33395.0 92595.0 32050.0 ;
      RECT  91890.0 33395.0 92595.0 34740.0 ;
      RECT  91890.0 36085.0 92595.0 34740.0 ;
      RECT  91890.0 36085.0 92595.0 37430.0 ;
      RECT  91890.0 38775.0 92595.0 37430.0 ;
      RECT  91890.0 38775.0 92595.0 40120.0 ;
      RECT  91890.0 41465.0 92595.0 40120.0 ;
      RECT  91890.0 41465.0 92595.0 42810.0 ;
      RECT  91890.0 44155.0 92595.0 42810.0 ;
      RECT  91890.0 44155.0 92595.0 45500.0 ;
      RECT  91890.0 46845.0 92595.0 45500.0 ;
      RECT  91890.0 46845.0 92595.0 48190.0 ;
      RECT  91890.0 49535.0 92595.0 48190.0 ;
      RECT  91890.0 49535.0 92595.0 50880.0 ;
      RECT  91890.0 52225.0 92595.0 50880.0 ;
      RECT  91890.0 52225.0 92595.0 53570.0 ;
      RECT  91890.0 54915.0 92595.0 53570.0 ;
      RECT  91890.0 54915.0 92595.0 56260.0 ;
      RECT  91890.0 57605.0 92595.0 56260.0 ;
      RECT  91890.0 57605.0 92595.0 58950.0 ;
      RECT  91890.0 60295.0 92595.0 58950.0 ;
      RECT  91890.0 60295.0 92595.0 61640.0 ;
      RECT  91890.0 62985.0 92595.0 61640.0 ;
      RECT  91890.0 62985.0 92595.0 64330.0 ;
      RECT  91890.0 65675.0 92595.0 64330.0 ;
      RECT  91890.0 65675.0 92595.0 67020.0 ;
      RECT  91890.0 68365.0 92595.0 67020.0 ;
      RECT  91890.0 68365.0 92595.0 69710.0 ;
      RECT  91890.0 71055.0 92595.0 69710.0 ;
      RECT  91890.0 71055.0 92595.0 72400.0 ;
      RECT  91890.0 73745.0 92595.0 72400.0 ;
      RECT  91890.0 73745.0 92595.0 75090.0 ;
      RECT  91890.0 76435.0 92595.0 75090.0 ;
      RECT  91890.0 76435.0 92595.0 77780.0 ;
      RECT  91890.0 79125.0 92595.0 77780.0 ;
      RECT  91890.0 79125.0 92595.0 80470.0 ;
      RECT  91890.0 81815.0 92595.0 80470.0 ;
      RECT  91890.0 81815.0 92595.0 83160.0 ;
      RECT  91890.0 84505.0 92595.0 83160.0 ;
      RECT  91890.0 84505.0 92595.0 85850.0 ;
      RECT  91890.0 87195.0 92595.0 85850.0 ;
      RECT  91890.0 87195.0 92595.0 88540.0 ;
      RECT  91890.0 89885.0 92595.0 88540.0 ;
      RECT  91890.0 89885.0 92595.0 91230.0 ;
      RECT  91890.0 92575.0 92595.0 91230.0 ;
      RECT  91890.0 92575.0 92595.0 93920.0 ;
      RECT  91890.0 95265.0 92595.0 93920.0 ;
      RECT  91890.0 95265.0 92595.0 96610.0 ;
      RECT  91890.0 97955.0 92595.0 96610.0 ;
      RECT  91890.0 97955.0 92595.0 99300.0 ;
      RECT  91890.0 100645.0 92595.0 99300.0 ;
      RECT  91890.0 100645.0 92595.0 101990.0 ;
      RECT  91890.0 103335.0 92595.0 101990.0 ;
      RECT  91890.0 103335.0 92595.0 104680.0 ;
      RECT  91890.0 106025.0 92595.0 104680.0 ;
      RECT  91890.0 106025.0 92595.0 107370.0 ;
      RECT  91890.0 108715.0 92595.0 107370.0 ;
      RECT  91890.0 108715.0 92595.0 110060.0 ;
      RECT  91890.0 111405.0 92595.0 110060.0 ;
      RECT  91890.0 111405.0 92595.0 112750.0 ;
      RECT  91890.0 114095.0 92595.0 112750.0 ;
      RECT  92595.0 28015.0 93300.0 29360.0 ;
      RECT  92595.0 30705.0 93300.0 29360.0 ;
      RECT  92595.0 30705.0 93300.0 32050.0 ;
      RECT  92595.0 33395.0 93300.0 32050.0 ;
      RECT  92595.0 33395.0 93300.0 34740.0 ;
      RECT  92595.0 36085.0 93300.0 34740.0 ;
      RECT  92595.0 36085.0 93300.0 37430.0 ;
      RECT  92595.0 38775.0 93300.0 37430.0 ;
      RECT  92595.0 38775.0 93300.0 40120.0 ;
      RECT  92595.0 41465.0 93300.0 40120.0 ;
      RECT  92595.0 41465.0 93300.0 42810.0 ;
      RECT  92595.0 44155.0 93300.0 42810.0 ;
      RECT  92595.0 44155.0 93300.0 45500.0 ;
      RECT  92595.0 46845.0 93300.0 45500.0 ;
      RECT  92595.0 46845.0 93300.0 48190.0 ;
      RECT  92595.0 49535.0 93300.0 48190.0 ;
      RECT  92595.0 49535.0 93300.0 50880.0 ;
      RECT  92595.0 52225.0 93300.0 50880.0 ;
      RECT  92595.0 52225.0 93300.0 53570.0 ;
      RECT  92595.0 54915.0 93300.0 53570.0 ;
      RECT  92595.0 54915.0 93300.0 56260.0 ;
      RECT  92595.0 57605.0 93300.0 56260.0 ;
      RECT  92595.0 57605.0 93300.0 58950.0 ;
      RECT  92595.0 60295.0 93300.0 58950.0 ;
      RECT  92595.0 60295.0 93300.0 61640.0 ;
      RECT  92595.0 62985.0 93300.0 61640.0 ;
      RECT  92595.0 62985.0 93300.0 64330.0 ;
      RECT  92595.0 65675.0 93300.0 64330.0 ;
      RECT  92595.0 65675.0 93300.0 67020.0 ;
      RECT  92595.0 68365.0 93300.0 67020.0 ;
      RECT  92595.0 68365.0 93300.0 69710.0 ;
      RECT  92595.0 71055.0 93300.0 69710.0 ;
      RECT  92595.0 71055.0 93300.0 72400.0 ;
      RECT  92595.0 73745.0 93300.0 72400.0 ;
      RECT  92595.0 73745.0 93300.0 75090.0 ;
      RECT  92595.0 76435.0 93300.0 75090.0 ;
      RECT  92595.0 76435.0 93300.0 77780.0 ;
      RECT  92595.0 79125.0 93300.0 77780.0 ;
      RECT  92595.0 79125.0 93300.0 80470.0 ;
      RECT  92595.0 81815.0 93300.0 80470.0 ;
      RECT  92595.0 81815.0 93300.0 83160.0 ;
      RECT  92595.0 84505.0 93300.0 83160.0 ;
      RECT  92595.0 84505.0 93300.0 85850.0 ;
      RECT  92595.0 87195.0 93300.0 85850.0 ;
      RECT  92595.0 87195.0 93300.0 88540.0 ;
      RECT  92595.0 89885.0 93300.0 88540.0 ;
      RECT  92595.0 89885.0 93300.0 91230.0 ;
      RECT  92595.0 92575.0 93300.0 91230.0 ;
      RECT  92595.0 92575.0 93300.0 93920.0 ;
      RECT  92595.0 95265.0 93300.0 93920.0 ;
      RECT  92595.0 95265.0 93300.0 96610.0 ;
      RECT  92595.0 97955.0 93300.0 96610.0 ;
      RECT  92595.0 97955.0 93300.0 99300.0 ;
      RECT  92595.0 100645.0 93300.0 99300.0 ;
      RECT  92595.0 100645.0 93300.0 101990.0 ;
      RECT  92595.0 103335.0 93300.0 101990.0 ;
      RECT  92595.0 103335.0 93300.0 104680.0 ;
      RECT  92595.0 106025.0 93300.0 104680.0 ;
      RECT  92595.0 106025.0 93300.0 107370.0 ;
      RECT  92595.0 108715.0 93300.0 107370.0 ;
      RECT  92595.0 108715.0 93300.0 110060.0 ;
      RECT  92595.0 111405.0 93300.0 110060.0 ;
      RECT  92595.0 111405.0 93300.0 112750.0 ;
      RECT  92595.0 114095.0 93300.0 112750.0 ;
      RECT  93300.0 28015.0 94005.0 29360.0 ;
      RECT  93300.0 30705.0 94005.0 29360.0 ;
      RECT  93300.0 30705.0 94005.0 32050.0 ;
      RECT  93300.0 33395.0 94005.0 32050.0 ;
      RECT  93300.0 33395.0 94005.0 34740.0 ;
      RECT  93300.0 36085.0 94005.0 34740.0 ;
      RECT  93300.0 36085.0 94005.0 37430.0 ;
      RECT  93300.0 38775.0 94005.0 37430.0 ;
      RECT  93300.0 38775.0 94005.0 40120.0 ;
      RECT  93300.0 41465.0 94005.0 40120.0 ;
      RECT  93300.0 41465.0 94005.0 42810.0 ;
      RECT  93300.0 44155.0 94005.0 42810.0 ;
      RECT  93300.0 44155.0 94005.0 45500.0 ;
      RECT  93300.0 46845.0 94005.0 45500.0 ;
      RECT  93300.0 46845.0 94005.0 48190.0 ;
      RECT  93300.0 49535.0 94005.0 48190.0 ;
      RECT  93300.0 49535.0 94005.0 50880.0 ;
      RECT  93300.0 52225.0 94005.0 50880.0 ;
      RECT  93300.0 52225.0 94005.0 53570.0 ;
      RECT  93300.0 54915.0 94005.0 53570.0 ;
      RECT  93300.0 54915.0 94005.0 56260.0 ;
      RECT  93300.0 57605.0 94005.0 56260.0 ;
      RECT  93300.0 57605.0 94005.0 58950.0 ;
      RECT  93300.0 60295.0 94005.0 58950.0 ;
      RECT  93300.0 60295.0 94005.0 61640.0 ;
      RECT  93300.0 62985.0 94005.0 61640.0 ;
      RECT  93300.0 62985.0 94005.0 64330.0 ;
      RECT  93300.0 65675.0 94005.0 64330.0 ;
      RECT  93300.0 65675.0 94005.0 67020.0 ;
      RECT  93300.0 68365.0 94005.0 67020.0 ;
      RECT  93300.0 68365.0 94005.0 69710.0 ;
      RECT  93300.0 71055.0 94005.0 69710.0 ;
      RECT  93300.0 71055.0 94005.0 72400.0 ;
      RECT  93300.0 73745.0 94005.0 72400.0 ;
      RECT  93300.0 73745.0 94005.0 75090.0 ;
      RECT  93300.0 76435.0 94005.0 75090.0 ;
      RECT  93300.0 76435.0 94005.0 77780.0 ;
      RECT  93300.0 79125.0 94005.0 77780.0 ;
      RECT  93300.0 79125.0 94005.0 80470.0 ;
      RECT  93300.0 81815.0 94005.0 80470.0 ;
      RECT  93300.0 81815.0 94005.0 83160.0 ;
      RECT  93300.0 84505.0 94005.0 83160.0 ;
      RECT  93300.0 84505.0 94005.0 85850.0 ;
      RECT  93300.0 87195.0 94005.0 85850.0 ;
      RECT  93300.0 87195.0 94005.0 88540.0 ;
      RECT  93300.0 89885.0 94005.0 88540.0 ;
      RECT  93300.0 89885.0 94005.0 91230.0 ;
      RECT  93300.0 92575.0 94005.0 91230.0 ;
      RECT  93300.0 92575.0 94005.0 93920.0 ;
      RECT  93300.0 95265.0 94005.0 93920.0 ;
      RECT  93300.0 95265.0 94005.0 96610.0 ;
      RECT  93300.0 97955.0 94005.0 96610.0 ;
      RECT  93300.0 97955.0 94005.0 99300.0 ;
      RECT  93300.0 100645.0 94005.0 99300.0 ;
      RECT  93300.0 100645.0 94005.0 101990.0 ;
      RECT  93300.0 103335.0 94005.0 101990.0 ;
      RECT  93300.0 103335.0 94005.0 104680.0 ;
      RECT  93300.0 106025.0 94005.0 104680.0 ;
      RECT  93300.0 106025.0 94005.0 107370.0 ;
      RECT  93300.0 108715.0 94005.0 107370.0 ;
      RECT  93300.0 108715.0 94005.0 110060.0 ;
      RECT  93300.0 111405.0 94005.0 110060.0 ;
      RECT  93300.0 111405.0 94005.0 112750.0 ;
      RECT  93300.0 114095.0 94005.0 112750.0 ;
      RECT  94005.0 28015.0 94710.0 29360.0 ;
      RECT  94005.0 30705.0 94710.0 29360.0 ;
      RECT  94005.0 30705.0 94710.0 32050.0 ;
      RECT  94005.0 33395.0 94710.0 32050.0 ;
      RECT  94005.0 33395.0 94710.0 34740.0 ;
      RECT  94005.0 36085.0 94710.0 34740.0 ;
      RECT  94005.0 36085.0 94710.0 37430.0 ;
      RECT  94005.0 38775.0 94710.0 37430.0 ;
      RECT  94005.0 38775.0 94710.0 40120.0 ;
      RECT  94005.0 41465.0 94710.0 40120.0 ;
      RECT  94005.0 41465.0 94710.0 42810.0 ;
      RECT  94005.0 44155.0 94710.0 42810.0 ;
      RECT  94005.0 44155.0 94710.0 45500.0 ;
      RECT  94005.0 46845.0 94710.0 45500.0 ;
      RECT  94005.0 46845.0 94710.0 48190.0 ;
      RECT  94005.0 49535.0 94710.0 48190.0 ;
      RECT  94005.0 49535.0 94710.0 50880.0 ;
      RECT  94005.0 52225.0 94710.0 50880.0 ;
      RECT  94005.0 52225.0 94710.0 53570.0 ;
      RECT  94005.0 54915.0 94710.0 53570.0 ;
      RECT  94005.0 54915.0 94710.0 56260.0 ;
      RECT  94005.0 57605.0 94710.0 56260.0 ;
      RECT  94005.0 57605.0 94710.0 58950.0 ;
      RECT  94005.0 60295.0 94710.0 58950.0 ;
      RECT  94005.0 60295.0 94710.0 61640.0 ;
      RECT  94005.0 62985.0 94710.0 61640.0 ;
      RECT  94005.0 62985.0 94710.0 64330.0 ;
      RECT  94005.0 65675.0 94710.0 64330.0 ;
      RECT  94005.0 65675.0 94710.0 67020.0 ;
      RECT  94005.0 68365.0 94710.0 67020.0 ;
      RECT  94005.0 68365.0 94710.0 69710.0 ;
      RECT  94005.0 71055.0 94710.0 69710.0 ;
      RECT  94005.0 71055.0 94710.0 72400.0 ;
      RECT  94005.0 73745.0 94710.0 72400.0 ;
      RECT  94005.0 73745.0 94710.0 75090.0 ;
      RECT  94005.0 76435.0 94710.0 75090.0 ;
      RECT  94005.0 76435.0 94710.0 77780.0 ;
      RECT  94005.0 79125.0 94710.0 77780.0 ;
      RECT  94005.0 79125.0 94710.0 80470.0 ;
      RECT  94005.0 81815.0 94710.0 80470.0 ;
      RECT  94005.0 81815.0 94710.0 83160.0 ;
      RECT  94005.0 84505.0 94710.0 83160.0 ;
      RECT  94005.0 84505.0 94710.0 85850.0 ;
      RECT  94005.0 87195.0 94710.0 85850.0 ;
      RECT  94005.0 87195.0 94710.0 88540.0 ;
      RECT  94005.0 89885.0 94710.0 88540.0 ;
      RECT  94005.0 89885.0 94710.0 91230.0 ;
      RECT  94005.0 92575.0 94710.0 91230.0 ;
      RECT  94005.0 92575.0 94710.0 93920.0 ;
      RECT  94005.0 95265.0 94710.0 93920.0 ;
      RECT  94005.0 95265.0 94710.0 96610.0 ;
      RECT  94005.0 97955.0 94710.0 96610.0 ;
      RECT  94005.0 97955.0 94710.0 99300.0 ;
      RECT  94005.0 100645.0 94710.0 99300.0 ;
      RECT  94005.0 100645.0 94710.0 101990.0 ;
      RECT  94005.0 103335.0 94710.0 101990.0 ;
      RECT  94005.0 103335.0 94710.0 104680.0 ;
      RECT  94005.0 106025.0 94710.0 104680.0 ;
      RECT  94005.0 106025.0 94710.0 107370.0 ;
      RECT  94005.0 108715.0 94710.0 107370.0 ;
      RECT  94005.0 108715.0 94710.0 110060.0 ;
      RECT  94005.0 111405.0 94710.0 110060.0 ;
      RECT  94005.0 111405.0 94710.0 112750.0 ;
      RECT  94005.0 114095.0 94710.0 112750.0 ;
      RECT  94710.0 28015.0 95415.0 29360.0 ;
      RECT  94710.0 30705.0 95415.0 29360.0 ;
      RECT  94710.0 30705.0 95415.0 32050.0 ;
      RECT  94710.0 33395.0 95415.0 32050.0 ;
      RECT  94710.0 33395.0 95415.0 34740.0 ;
      RECT  94710.0 36085.0 95415.0 34740.0 ;
      RECT  94710.0 36085.0 95415.0 37430.0 ;
      RECT  94710.0 38775.0 95415.0 37430.0 ;
      RECT  94710.0 38775.0 95415.0 40120.0 ;
      RECT  94710.0 41465.0 95415.0 40120.0 ;
      RECT  94710.0 41465.0 95415.0 42810.0 ;
      RECT  94710.0 44155.0 95415.0 42810.0 ;
      RECT  94710.0 44155.0 95415.0 45500.0 ;
      RECT  94710.0 46845.0 95415.0 45500.0 ;
      RECT  94710.0 46845.0 95415.0 48190.0 ;
      RECT  94710.0 49535.0 95415.0 48190.0 ;
      RECT  94710.0 49535.0 95415.0 50880.0 ;
      RECT  94710.0 52225.0 95415.0 50880.0 ;
      RECT  94710.0 52225.0 95415.0 53570.0 ;
      RECT  94710.0 54915.0 95415.0 53570.0 ;
      RECT  94710.0 54915.0 95415.0 56260.0 ;
      RECT  94710.0 57605.0 95415.0 56260.0 ;
      RECT  94710.0 57605.0 95415.0 58950.0 ;
      RECT  94710.0 60295.0 95415.0 58950.0 ;
      RECT  94710.0 60295.0 95415.0 61640.0 ;
      RECT  94710.0 62985.0 95415.0 61640.0 ;
      RECT  94710.0 62985.0 95415.0 64330.0 ;
      RECT  94710.0 65675.0 95415.0 64330.0 ;
      RECT  94710.0 65675.0 95415.0 67020.0 ;
      RECT  94710.0 68365.0 95415.0 67020.0 ;
      RECT  94710.0 68365.0 95415.0 69710.0 ;
      RECT  94710.0 71055.0 95415.0 69710.0 ;
      RECT  94710.0 71055.0 95415.0 72400.0 ;
      RECT  94710.0 73745.0 95415.0 72400.0 ;
      RECT  94710.0 73745.0 95415.0 75090.0 ;
      RECT  94710.0 76435.0 95415.0 75090.0 ;
      RECT  94710.0 76435.0 95415.0 77780.0 ;
      RECT  94710.0 79125.0 95415.0 77780.0 ;
      RECT  94710.0 79125.0 95415.0 80470.0 ;
      RECT  94710.0 81815.0 95415.0 80470.0 ;
      RECT  94710.0 81815.0 95415.0 83160.0 ;
      RECT  94710.0 84505.0 95415.0 83160.0 ;
      RECT  94710.0 84505.0 95415.0 85850.0 ;
      RECT  94710.0 87195.0 95415.0 85850.0 ;
      RECT  94710.0 87195.0 95415.0 88540.0 ;
      RECT  94710.0 89885.0 95415.0 88540.0 ;
      RECT  94710.0 89885.0 95415.0 91230.0 ;
      RECT  94710.0 92575.0 95415.0 91230.0 ;
      RECT  94710.0 92575.0 95415.0 93920.0 ;
      RECT  94710.0 95265.0 95415.0 93920.0 ;
      RECT  94710.0 95265.0 95415.0 96610.0 ;
      RECT  94710.0 97955.0 95415.0 96610.0 ;
      RECT  94710.0 97955.0 95415.0 99300.0 ;
      RECT  94710.0 100645.0 95415.0 99300.0 ;
      RECT  94710.0 100645.0 95415.0 101990.0 ;
      RECT  94710.0 103335.0 95415.0 101990.0 ;
      RECT  94710.0 103335.0 95415.0 104680.0 ;
      RECT  94710.0 106025.0 95415.0 104680.0 ;
      RECT  94710.0 106025.0 95415.0 107370.0 ;
      RECT  94710.0 108715.0 95415.0 107370.0 ;
      RECT  94710.0 108715.0 95415.0 110060.0 ;
      RECT  94710.0 111405.0 95415.0 110060.0 ;
      RECT  94710.0 111405.0 95415.0 112750.0 ;
      RECT  94710.0 114095.0 95415.0 112750.0 ;
      RECT  95415.0 28015.0 96120.0 29360.0 ;
      RECT  95415.0 30705.0 96120.0 29360.0 ;
      RECT  95415.0 30705.0 96120.0 32050.0 ;
      RECT  95415.0 33395.0 96120.0 32050.0 ;
      RECT  95415.0 33395.0 96120.0 34740.0 ;
      RECT  95415.0 36085.0 96120.0 34740.0 ;
      RECT  95415.0 36085.0 96120.0 37430.0 ;
      RECT  95415.0 38775.0 96120.0 37430.0 ;
      RECT  95415.0 38775.0 96120.0 40120.0 ;
      RECT  95415.0 41465.0 96120.0 40120.0 ;
      RECT  95415.0 41465.0 96120.0 42810.0 ;
      RECT  95415.0 44155.0 96120.0 42810.0 ;
      RECT  95415.0 44155.0 96120.0 45500.0 ;
      RECT  95415.0 46845.0 96120.0 45500.0 ;
      RECT  95415.0 46845.0 96120.0 48190.0 ;
      RECT  95415.0 49535.0 96120.0 48190.0 ;
      RECT  95415.0 49535.0 96120.0 50880.0 ;
      RECT  95415.0 52225.0 96120.0 50880.0 ;
      RECT  95415.0 52225.0 96120.0 53570.0 ;
      RECT  95415.0 54915.0 96120.0 53570.0 ;
      RECT  95415.0 54915.0 96120.0 56260.0 ;
      RECT  95415.0 57605.0 96120.0 56260.0 ;
      RECT  95415.0 57605.0 96120.0 58950.0 ;
      RECT  95415.0 60295.0 96120.0 58950.0 ;
      RECT  95415.0 60295.0 96120.0 61640.0 ;
      RECT  95415.0 62985.0 96120.0 61640.0 ;
      RECT  95415.0 62985.0 96120.0 64330.0 ;
      RECT  95415.0 65675.0 96120.0 64330.0 ;
      RECT  95415.0 65675.0 96120.0 67020.0 ;
      RECT  95415.0 68365.0 96120.0 67020.0 ;
      RECT  95415.0 68365.0 96120.0 69710.0 ;
      RECT  95415.0 71055.0 96120.0 69710.0 ;
      RECT  95415.0 71055.0 96120.0 72400.0 ;
      RECT  95415.0 73745.0 96120.0 72400.0 ;
      RECT  95415.0 73745.0 96120.0 75090.0 ;
      RECT  95415.0 76435.0 96120.0 75090.0 ;
      RECT  95415.0 76435.0 96120.0 77780.0 ;
      RECT  95415.0 79125.0 96120.0 77780.0 ;
      RECT  95415.0 79125.0 96120.0 80470.0 ;
      RECT  95415.0 81815.0 96120.0 80470.0 ;
      RECT  95415.0 81815.0 96120.0 83160.0 ;
      RECT  95415.0 84505.0 96120.0 83160.0 ;
      RECT  95415.0 84505.0 96120.0 85850.0 ;
      RECT  95415.0 87195.0 96120.0 85850.0 ;
      RECT  95415.0 87195.0 96120.0 88540.0 ;
      RECT  95415.0 89885.0 96120.0 88540.0 ;
      RECT  95415.0 89885.0 96120.0 91230.0 ;
      RECT  95415.0 92575.0 96120.0 91230.0 ;
      RECT  95415.0 92575.0 96120.0 93920.0 ;
      RECT  95415.0 95265.0 96120.0 93920.0 ;
      RECT  95415.0 95265.0 96120.0 96610.0 ;
      RECT  95415.0 97955.0 96120.0 96610.0 ;
      RECT  95415.0 97955.0 96120.0 99300.0 ;
      RECT  95415.0 100645.0 96120.0 99300.0 ;
      RECT  95415.0 100645.0 96120.0 101990.0 ;
      RECT  95415.0 103335.0 96120.0 101990.0 ;
      RECT  95415.0 103335.0 96120.0 104680.0 ;
      RECT  95415.0 106025.0 96120.0 104680.0 ;
      RECT  95415.0 106025.0 96120.0 107370.0 ;
      RECT  95415.0 108715.0 96120.0 107370.0 ;
      RECT  95415.0 108715.0 96120.0 110060.0 ;
      RECT  95415.0 111405.0 96120.0 110060.0 ;
      RECT  95415.0 111405.0 96120.0 112750.0 ;
      RECT  95415.0 114095.0 96120.0 112750.0 ;
      RECT  96120.0 28015.0 96825.0 29360.0 ;
      RECT  96120.0 30705.0 96825.0 29360.0 ;
      RECT  96120.0 30705.0 96825.0 32050.0 ;
      RECT  96120.0 33395.0 96825.0 32050.0 ;
      RECT  96120.0 33395.0 96825.0 34740.0 ;
      RECT  96120.0 36085.0 96825.0 34740.0 ;
      RECT  96120.0 36085.0 96825.0 37430.0 ;
      RECT  96120.0 38775.0 96825.0 37430.0 ;
      RECT  96120.0 38775.0 96825.0 40120.0 ;
      RECT  96120.0 41465.0 96825.0 40120.0 ;
      RECT  96120.0 41465.0 96825.0 42810.0 ;
      RECT  96120.0 44155.0 96825.0 42810.0 ;
      RECT  96120.0 44155.0 96825.0 45500.0 ;
      RECT  96120.0 46845.0 96825.0 45500.0 ;
      RECT  96120.0 46845.0 96825.0 48190.0 ;
      RECT  96120.0 49535.0 96825.0 48190.0 ;
      RECT  96120.0 49535.0 96825.0 50880.0 ;
      RECT  96120.0 52225.0 96825.0 50880.0 ;
      RECT  96120.0 52225.0 96825.0 53570.0 ;
      RECT  96120.0 54915.0 96825.0 53570.0 ;
      RECT  96120.0 54915.0 96825.0 56260.0 ;
      RECT  96120.0 57605.0 96825.0 56260.0 ;
      RECT  96120.0 57605.0 96825.0 58950.0 ;
      RECT  96120.0 60295.0 96825.0 58950.0 ;
      RECT  96120.0 60295.0 96825.0 61640.0 ;
      RECT  96120.0 62985.0 96825.0 61640.0 ;
      RECT  96120.0 62985.0 96825.0 64330.0 ;
      RECT  96120.0 65675.0 96825.0 64330.0 ;
      RECT  96120.0 65675.0 96825.0 67020.0 ;
      RECT  96120.0 68365.0 96825.0 67020.0 ;
      RECT  96120.0 68365.0 96825.0 69710.0 ;
      RECT  96120.0 71055.0 96825.0 69710.0 ;
      RECT  96120.0 71055.0 96825.0 72400.0 ;
      RECT  96120.0 73745.0 96825.0 72400.0 ;
      RECT  96120.0 73745.0 96825.0 75090.0 ;
      RECT  96120.0 76435.0 96825.0 75090.0 ;
      RECT  96120.0 76435.0 96825.0 77780.0 ;
      RECT  96120.0 79125.0 96825.0 77780.0 ;
      RECT  96120.0 79125.0 96825.0 80470.0 ;
      RECT  96120.0 81815.0 96825.0 80470.0 ;
      RECT  96120.0 81815.0 96825.0 83160.0 ;
      RECT  96120.0 84505.0 96825.0 83160.0 ;
      RECT  96120.0 84505.0 96825.0 85850.0 ;
      RECT  96120.0 87195.0 96825.0 85850.0 ;
      RECT  96120.0 87195.0 96825.0 88540.0 ;
      RECT  96120.0 89885.0 96825.0 88540.0 ;
      RECT  96120.0 89885.0 96825.0 91230.0 ;
      RECT  96120.0 92575.0 96825.0 91230.0 ;
      RECT  96120.0 92575.0 96825.0 93920.0 ;
      RECT  96120.0 95265.0 96825.0 93920.0 ;
      RECT  96120.0 95265.0 96825.0 96610.0 ;
      RECT  96120.0 97955.0 96825.0 96610.0 ;
      RECT  96120.0 97955.0 96825.0 99300.0 ;
      RECT  96120.0 100645.0 96825.0 99300.0 ;
      RECT  96120.0 100645.0 96825.0 101990.0 ;
      RECT  96120.0 103335.0 96825.0 101990.0 ;
      RECT  96120.0 103335.0 96825.0 104680.0 ;
      RECT  96120.0 106025.0 96825.0 104680.0 ;
      RECT  96120.0 106025.0 96825.0 107370.0 ;
      RECT  96120.0 108715.0 96825.0 107370.0 ;
      RECT  96120.0 108715.0 96825.0 110060.0 ;
      RECT  96120.0 111405.0 96825.0 110060.0 ;
      RECT  96120.0 111405.0 96825.0 112750.0 ;
      RECT  96120.0 114095.0 96825.0 112750.0 ;
      RECT  96825.0 28015.0 97530.0 29360.0 ;
      RECT  96825.0 30705.0 97530.0 29360.0 ;
      RECT  96825.0 30705.0 97530.0 32050.0 ;
      RECT  96825.0 33395.0 97530.0 32050.0 ;
      RECT  96825.0 33395.0 97530.0 34740.0 ;
      RECT  96825.0 36085.0 97530.0 34740.0 ;
      RECT  96825.0 36085.0 97530.0 37430.0 ;
      RECT  96825.0 38775.0 97530.0 37430.0 ;
      RECT  96825.0 38775.0 97530.0 40120.0 ;
      RECT  96825.0 41465.0 97530.0 40120.0 ;
      RECT  96825.0 41465.0 97530.0 42810.0 ;
      RECT  96825.0 44155.0 97530.0 42810.0 ;
      RECT  96825.0 44155.0 97530.0 45500.0 ;
      RECT  96825.0 46845.0 97530.0 45500.0 ;
      RECT  96825.0 46845.0 97530.0 48190.0 ;
      RECT  96825.0 49535.0 97530.0 48190.0 ;
      RECT  96825.0 49535.0 97530.0 50880.0 ;
      RECT  96825.0 52225.0 97530.0 50880.0 ;
      RECT  96825.0 52225.0 97530.0 53570.0 ;
      RECT  96825.0 54915.0 97530.0 53570.0 ;
      RECT  96825.0 54915.0 97530.0 56260.0 ;
      RECT  96825.0 57605.0 97530.0 56260.0 ;
      RECT  96825.0 57605.0 97530.0 58950.0 ;
      RECT  96825.0 60295.0 97530.0 58950.0 ;
      RECT  96825.0 60295.0 97530.0 61640.0 ;
      RECT  96825.0 62985.0 97530.0 61640.0 ;
      RECT  96825.0 62985.0 97530.0 64330.0 ;
      RECT  96825.0 65675.0 97530.0 64330.0 ;
      RECT  96825.0 65675.0 97530.0 67020.0 ;
      RECT  96825.0 68365.0 97530.0 67020.0 ;
      RECT  96825.0 68365.0 97530.0 69710.0 ;
      RECT  96825.0 71055.0 97530.0 69710.0 ;
      RECT  96825.0 71055.0 97530.0 72400.0 ;
      RECT  96825.0 73745.0 97530.0 72400.0 ;
      RECT  96825.0 73745.0 97530.0 75090.0 ;
      RECT  96825.0 76435.0 97530.0 75090.0 ;
      RECT  96825.0 76435.0 97530.0 77780.0 ;
      RECT  96825.0 79125.0 97530.0 77780.0 ;
      RECT  96825.0 79125.0 97530.0 80470.0 ;
      RECT  96825.0 81815.0 97530.0 80470.0 ;
      RECT  96825.0 81815.0 97530.0 83160.0 ;
      RECT  96825.0 84505.0 97530.0 83160.0 ;
      RECT  96825.0 84505.0 97530.0 85850.0 ;
      RECT  96825.0 87195.0 97530.0 85850.0 ;
      RECT  96825.0 87195.0 97530.0 88540.0 ;
      RECT  96825.0 89885.0 97530.0 88540.0 ;
      RECT  96825.0 89885.0 97530.0 91230.0 ;
      RECT  96825.0 92575.0 97530.0 91230.0 ;
      RECT  96825.0 92575.0 97530.0 93920.0 ;
      RECT  96825.0 95265.0 97530.0 93920.0 ;
      RECT  96825.0 95265.0 97530.0 96610.0 ;
      RECT  96825.0 97955.0 97530.0 96610.0 ;
      RECT  96825.0 97955.0 97530.0 99300.0 ;
      RECT  96825.0 100645.0 97530.0 99300.0 ;
      RECT  96825.0 100645.0 97530.0 101990.0 ;
      RECT  96825.0 103335.0 97530.0 101990.0 ;
      RECT  96825.0 103335.0 97530.0 104680.0 ;
      RECT  96825.0 106025.0 97530.0 104680.0 ;
      RECT  96825.0 106025.0 97530.0 107370.0 ;
      RECT  96825.0 108715.0 97530.0 107370.0 ;
      RECT  96825.0 108715.0 97530.0 110060.0 ;
      RECT  96825.0 111405.0 97530.0 110060.0 ;
      RECT  96825.0 111405.0 97530.0 112750.0 ;
      RECT  96825.0 114095.0 97530.0 112750.0 ;
      RECT  97530.0 28015.0 98235.0 29360.0 ;
      RECT  97530.0 30705.0 98235.0 29360.0 ;
      RECT  97530.0 30705.0 98235.0 32050.0 ;
      RECT  97530.0 33395.0 98235.0 32050.0 ;
      RECT  97530.0 33395.0 98235.0 34740.0 ;
      RECT  97530.0 36085.0 98235.0 34740.0 ;
      RECT  97530.0 36085.0 98235.0 37430.0 ;
      RECT  97530.0 38775.0 98235.0 37430.0 ;
      RECT  97530.0 38775.0 98235.0 40120.0 ;
      RECT  97530.0 41465.0 98235.0 40120.0 ;
      RECT  97530.0 41465.0 98235.0 42810.0 ;
      RECT  97530.0 44155.0 98235.0 42810.0 ;
      RECT  97530.0 44155.0 98235.0 45500.0 ;
      RECT  97530.0 46845.0 98235.0 45500.0 ;
      RECT  97530.0 46845.0 98235.0 48190.0 ;
      RECT  97530.0 49535.0 98235.0 48190.0 ;
      RECT  97530.0 49535.0 98235.0 50880.0 ;
      RECT  97530.0 52225.0 98235.0 50880.0 ;
      RECT  97530.0 52225.0 98235.0 53570.0 ;
      RECT  97530.0 54915.0 98235.0 53570.0 ;
      RECT  97530.0 54915.0 98235.0 56260.0 ;
      RECT  97530.0 57605.0 98235.0 56260.0 ;
      RECT  97530.0 57605.0 98235.0 58950.0 ;
      RECT  97530.0 60295.0 98235.0 58950.0 ;
      RECT  97530.0 60295.0 98235.0 61640.0 ;
      RECT  97530.0 62985.0 98235.0 61640.0 ;
      RECT  97530.0 62985.0 98235.0 64330.0 ;
      RECT  97530.0 65675.0 98235.0 64330.0 ;
      RECT  97530.0 65675.0 98235.0 67020.0 ;
      RECT  97530.0 68365.0 98235.0 67020.0 ;
      RECT  97530.0 68365.0 98235.0 69710.0 ;
      RECT  97530.0 71055.0 98235.0 69710.0 ;
      RECT  97530.0 71055.0 98235.0 72400.0 ;
      RECT  97530.0 73745.0 98235.0 72400.0 ;
      RECT  97530.0 73745.0 98235.0 75090.0 ;
      RECT  97530.0 76435.0 98235.0 75090.0 ;
      RECT  97530.0 76435.0 98235.0 77780.0 ;
      RECT  97530.0 79125.0 98235.0 77780.0 ;
      RECT  97530.0 79125.0 98235.0 80470.0 ;
      RECT  97530.0 81815.0 98235.0 80470.0 ;
      RECT  97530.0 81815.0 98235.0 83160.0 ;
      RECT  97530.0 84505.0 98235.0 83160.0 ;
      RECT  97530.0 84505.0 98235.0 85850.0 ;
      RECT  97530.0 87195.0 98235.0 85850.0 ;
      RECT  97530.0 87195.0 98235.0 88540.0 ;
      RECT  97530.0 89885.0 98235.0 88540.0 ;
      RECT  97530.0 89885.0 98235.0 91230.0 ;
      RECT  97530.0 92575.0 98235.0 91230.0 ;
      RECT  97530.0 92575.0 98235.0 93920.0 ;
      RECT  97530.0 95265.0 98235.0 93920.0 ;
      RECT  97530.0 95265.0 98235.0 96610.0 ;
      RECT  97530.0 97955.0 98235.0 96610.0 ;
      RECT  97530.0 97955.0 98235.0 99300.0 ;
      RECT  97530.0 100645.0 98235.0 99300.0 ;
      RECT  97530.0 100645.0 98235.0 101990.0 ;
      RECT  97530.0 103335.0 98235.0 101990.0 ;
      RECT  97530.0 103335.0 98235.0 104680.0 ;
      RECT  97530.0 106025.0 98235.0 104680.0 ;
      RECT  97530.0 106025.0 98235.0 107370.0 ;
      RECT  97530.0 108715.0 98235.0 107370.0 ;
      RECT  97530.0 108715.0 98235.0 110060.0 ;
      RECT  97530.0 111405.0 98235.0 110060.0 ;
      RECT  97530.0 111405.0 98235.0 112750.0 ;
      RECT  97530.0 114095.0 98235.0 112750.0 ;
      RECT  98235.0 28015.0 98940.0 29360.0 ;
      RECT  98235.0 30705.0 98940.0 29360.0 ;
      RECT  98235.0 30705.0 98940.0 32050.0 ;
      RECT  98235.0 33395.0 98940.0 32050.0 ;
      RECT  98235.0 33395.0 98940.0 34740.0 ;
      RECT  98235.0 36085.0 98940.0 34740.0 ;
      RECT  98235.0 36085.0 98940.0 37430.0 ;
      RECT  98235.0 38775.0 98940.0 37430.0 ;
      RECT  98235.0 38775.0 98940.0 40120.0 ;
      RECT  98235.0 41465.0 98940.0 40120.0 ;
      RECT  98235.0 41465.0 98940.0 42810.0 ;
      RECT  98235.0 44155.0 98940.0 42810.0 ;
      RECT  98235.0 44155.0 98940.0 45500.0 ;
      RECT  98235.0 46845.0 98940.0 45500.0 ;
      RECT  98235.0 46845.0 98940.0 48190.0 ;
      RECT  98235.0 49535.0 98940.0 48190.0 ;
      RECT  98235.0 49535.0 98940.0 50880.0 ;
      RECT  98235.0 52225.0 98940.0 50880.0 ;
      RECT  98235.0 52225.0 98940.0 53570.0 ;
      RECT  98235.0 54915.0 98940.0 53570.0 ;
      RECT  98235.0 54915.0 98940.0 56260.0 ;
      RECT  98235.0 57605.0 98940.0 56260.0 ;
      RECT  98235.0 57605.0 98940.0 58950.0 ;
      RECT  98235.0 60295.0 98940.0 58950.0 ;
      RECT  98235.0 60295.0 98940.0 61640.0 ;
      RECT  98235.0 62985.0 98940.0 61640.0 ;
      RECT  98235.0 62985.0 98940.0 64330.0 ;
      RECT  98235.0 65675.0 98940.0 64330.0 ;
      RECT  98235.0 65675.0 98940.0 67020.0 ;
      RECT  98235.0 68365.0 98940.0 67020.0 ;
      RECT  98235.0 68365.0 98940.0 69710.0 ;
      RECT  98235.0 71055.0 98940.0 69710.0 ;
      RECT  98235.0 71055.0 98940.0 72400.0 ;
      RECT  98235.0 73745.0 98940.0 72400.0 ;
      RECT  98235.0 73745.0 98940.0 75090.0 ;
      RECT  98235.0 76435.0 98940.0 75090.0 ;
      RECT  98235.0 76435.0 98940.0 77780.0 ;
      RECT  98235.0 79125.0 98940.0 77780.0 ;
      RECT  98235.0 79125.0 98940.0 80470.0 ;
      RECT  98235.0 81815.0 98940.0 80470.0 ;
      RECT  98235.0 81815.0 98940.0 83160.0 ;
      RECT  98235.0 84505.0 98940.0 83160.0 ;
      RECT  98235.0 84505.0 98940.0 85850.0 ;
      RECT  98235.0 87195.0 98940.0 85850.0 ;
      RECT  98235.0 87195.0 98940.0 88540.0 ;
      RECT  98235.0 89885.0 98940.0 88540.0 ;
      RECT  98235.0 89885.0 98940.0 91230.0 ;
      RECT  98235.0 92575.0 98940.0 91230.0 ;
      RECT  98235.0 92575.0 98940.0 93920.0 ;
      RECT  98235.0 95265.0 98940.0 93920.0 ;
      RECT  98235.0 95265.0 98940.0 96610.0 ;
      RECT  98235.0 97955.0 98940.0 96610.0 ;
      RECT  98235.0 97955.0 98940.0 99300.0 ;
      RECT  98235.0 100645.0 98940.0 99300.0 ;
      RECT  98235.0 100645.0 98940.0 101990.0 ;
      RECT  98235.0 103335.0 98940.0 101990.0 ;
      RECT  98235.0 103335.0 98940.0 104680.0 ;
      RECT  98235.0 106025.0 98940.0 104680.0 ;
      RECT  98235.0 106025.0 98940.0 107370.0 ;
      RECT  98235.0 108715.0 98940.0 107370.0 ;
      RECT  98235.0 108715.0 98940.0 110060.0 ;
      RECT  98235.0 111405.0 98940.0 110060.0 ;
      RECT  98235.0 111405.0 98940.0 112750.0 ;
      RECT  98235.0 114095.0 98940.0 112750.0 ;
      RECT  98940.0 28015.0 99645.0 29360.0 ;
      RECT  98940.0 30705.0 99645.0 29360.0 ;
      RECT  98940.0 30705.0 99645.0 32050.0 ;
      RECT  98940.0 33395.0 99645.0 32050.0 ;
      RECT  98940.0 33395.0 99645.0 34740.0 ;
      RECT  98940.0 36085.0 99645.0 34740.0 ;
      RECT  98940.0 36085.0 99645.0 37430.0 ;
      RECT  98940.0 38775.0 99645.0 37430.0 ;
      RECT  98940.0 38775.0 99645.0 40120.0 ;
      RECT  98940.0 41465.0 99645.0 40120.0 ;
      RECT  98940.0 41465.0 99645.0 42810.0 ;
      RECT  98940.0 44155.0 99645.0 42810.0 ;
      RECT  98940.0 44155.0 99645.0 45500.0 ;
      RECT  98940.0 46845.0 99645.0 45500.0 ;
      RECT  98940.0 46845.0 99645.0 48190.0 ;
      RECT  98940.0 49535.0 99645.0 48190.0 ;
      RECT  98940.0 49535.0 99645.0 50880.0 ;
      RECT  98940.0 52225.0 99645.0 50880.0 ;
      RECT  98940.0 52225.0 99645.0 53570.0 ;
      RECT  98940.0 54915.0 99645.0 53570.0 ;
      RECT  98940.0 54915.0 99645.0 56260.0 ;
      RECT  98940.0 57605.0 99645.0 56260.0 ;
      RECT  98940.0 57605.0 99645.0 58950.0 ;
      RECT  98940.0 60295.0 99645.0 58950.0 ;
      RECT  98940.0 60295.0 99645.0 61640.0 ;
      RECT  98940.0 62985.0 99645.0 61640.0 ;
      RECT  98940.0 62985.0 99645.0 64330.0 ;
      RECT  98940.0 65675.0 99645.0 64330.0 ;
      RECT  98940.0 65675.0 99645.0 67020.0 ;
      RECT  98940.0 68365.0 99645.0 67020.0 ;
      RECT  98940.0 68365.0 99645.0 69710.0 ;
      RECT  98940.0 71055.0 99645.0 69710.0 ;
      RECT  98940.0 71055.0 99645.0 72400.0 ;
      RECT  98940.0 73745.0 99645.0 72400.0 ;
      RECT  98940.0 73745.0 99645.0 75090.0 ;
      RECT  98940.0 76435.0 99645.0 75090.0 ;
      RECT  98940.0 76435.0 99645.0 77780.0 ;
      RECT  98940.0 79125.0 99645.0 77780.0 ;
      RECT  98940.0 79125.0 99645.0 80470.0 ;
      RECT  98940.0 81815.0 99645.0 80470.0 ;
      RECT  98940.0 81815.0 99645.0 83160.0 ;
      RECT  98940.0 84505.0 99645.0 83160.0 ;
      RECT  98940.0 84505.0 99645.0 85850.0 ;
      RECT  98940.0 87195.0 99645.0 85850.0 ;
      RECT  98940.0 87195.0 99645.0 88540.0 ;
      RECT  98940.0 89885.0 99645.0 88540.0 ;
      RECT  98940.0 89885.0 99645.0 91230.0 ;
      RECT  98940.0 92575.0 99645.0 91230.0 ;
      RECT  98940.0 92575.0 99645.0 93920.0 ;
      RECT  98940.0 95265.0 99645.0 93920.0 ;
      RECT  98940.0 95265.0 99645.0 96610.0 ;
      RECT  98940.0 97955.0 99645.0 96610.0 ;
      RECT  98940.0 97955.0 99645.0 99300.0 ;
      RECT  98940.0 100645.0 99645.0 99300.0 ;
      RECT  98940.0 100645.0 99645.0 101990.0 ;
      RECT  98940.0 103335.0 99645.0 101990.0 ;
      RECT  98940.0 103335.0 99645.0 104680.0 ;
      RECT  98940.0 106025.0 99645.0 104680.0 ;
      RECT  98940.0 106025.0 99645.0 107370.0 ;
      RECT  98940.0 108715.0 99645.0 107370.0 ;
      RECT  98940.0 108715.0 99645.0 110060.0 ;
      RECT  98940.0 111405.0 99645.0 110060.0 ;
      RECT  98940.0 111405.0 99645.0 112750.0 ;
      RECT  98940.0 114095.0 99645.0 112750.0 ;
      RECT  99645.0 28015.0 100350.0 29360.0 ;
      RECT  99645.0 30705.0 100350.0 29360.0 ;
      RECT  99645.0 30705.0 100350.0 32050.0 ;
      RECT  99645.0 33395.0 100350.0 32050.0 ;
      RECT  99645.0 33395.0 100350.0 34740.0 ;
      RECT  99645.0 36085.0 100350.0 34740.0 ;
      RECT  99645.0 36085.0 100350.0 37430.0 ;
      RECT  99645.0 38775.0 100350.0 37430.0 ;
      RECT  99645.0 38775.0 100350.0 40120.0 ;
      RECT  99645.0 41465.0 100350.0 40120.0 ;
      RECT  99645.0 41465.0 100350.0 42810.0 ;
      RECT  99645.0 44155.0 100350.0 42810.0 ;
      RECT  99645.0 44155.0 100350.0 45500.0 ;
      RECT  99645.0 46845.0 100350.0 45500.0 ;
      RECT  99645.0 46845.0 100350.0 48190.0 ;
      RECT  99645.0 49535.0 100350.0 48190.0 ;
      RECT  99645.0 49535.0 100350.0 50880.0 ;
      RECT  99645.0 52225.0 100350.0 50880.0 ;
      RECT  99645.0 52225.0 100350.0 53570.0 ;
      RECT  99645.0 54915.0 100350.0 53570.0 ;
      RECT  99645.0 54915.0 100350.0 56260.0 ;
      RECT  99645.0 57605.0 100350.0 56260.0 ;
      RECT  99645.0 57605.0 100350.0 58950.0 ;
      RECT  99645.0 60295.0 100350.0 58950.0 ;
      RECT  99645.0 60295.0 100350.0 61640.0 ;
      RECT  99645.0 62985.0 100350.0 61640.0 ;
      RECT  99645.0 62985.0 100350.0 64330.0 ;
      RECT  99645.0 65675.0 100350.0 64330.0 ;
      RECT  99645.0 65675.0 100350.0 67020.0 ;
      RECT  99645.0 68365.0 100350.0 67020.0 ;
      RECT  99645.0 68365.0 100350.0 69710.0 ;
      RECT  99645.0 71055.0 100350.0 69710.0 ;
      RECT  99645.0 71055.0 100350.0 72400.0 ;
      RECT  99645.0 73745.0 100350.0 72400.0 ;
      RECT  99645.0 73745.0 100350.0 75090.0 ;
      RECT  99645.0 76435.0 100350.0 75090.0 ;
      RECT  99645.0 76435.0 100350.0 77780.0 ;
      RECT  99645.0 79125.0 100350.0 77780.0 ;
      RECT  99645.0 79125.0 100350.0 80470.0 ;
      RECT  99645.0 81815.0 100350.0 80470.0 ;
      RECT  99645.0 81815.0 100350.0 83160.0 ;
      RECT  99645.0 84505.0 100350.0 83160.0 ;
      RECT  99645.0 84505.0 100350.0 85850.0 ;
      RECT  99645.0 87195.0 100350.0 85850.0 ;
      RECT  99645.0 87195.0 100350.0 88540.0 ;
      RECT  99645.0 89885.0 100350.0 88540.0 ;
      RECT  99645.0 89885.0 100350.0 91230.0 ;
      RECT  99645.0 92575.0 100350.0 91230.0 ;
      RECT  99645.0 92575.0 100350.0 93920.0 ;
      RECT  99645.0 95265.0 100350.0 93920.0 ;
      RECT  99645.0 95265.0 100350.0 96610.0 ;
      RECT  99645.0 97955.0 100350.0 96610.0 ;
      RECT  99645.0 97955.0 100350.0 99300.0 ;
      RECT  99645.0 100645.0 100350.0 99300.0 ;
      RECT  99645.0 100645.0 100350.0 101990.0 ;
      RECT  99645.0 103335.0 100350.0 101990.0 ;
      RECT  99645.0 103335.0 100350.0 104680.0 ;
      RECT  99645.0 106025.0 100350.0 104680.0 ;
      RECT  99645.0 106025.0 100350.0 107370.0 ;
      RECT  99645.0 108715.0 100350.0 107370.0 ;
      RECT  99645.0 108715.0 100350.0 110060.0 ;
      RECT  99645.0 111405.0 100350.0 110060.0 ;
      RECT  99645.0 111405.0 100350.0 112750.0 ;
      RECT  99645.0 114095.0 100350.0 112750.0 ;
      RECT  100350.0 28015.0 101055.0 29360.0 ;
      RECT  100350.0 30705.0 101055.0 29360.0 ;
      RECT  100350.0 30705.0 101055.0 32050.0 ;
      RECT  100350.0 33395.0 101055.0 32050.0 ;
      RECT  100350.0 33395.0 101055.0 34740.0 ;
      RECT  100350.0 36085.0 101055.0 34740.0 ;
      RECT  100350.0 36085.0 101055.0 37430.0 ;
      RECT  100350.0 38775.0 101055.0 37430.0 ;
      RECT  100350.0 38775.0 101055.0 40120.0 ;
      RECT  100350.0 41465.0 101055.0 40120.0 ;
      RECT  100350.0 41465.0 101055.0 42810.0 ;
      RECT  100350.0 44155.0 101055.0 42810.0 ;
      RECT  100350.0 44155.0 101055.0 45500.0 ;
      RECT  100350.0 46845.0 101055.0 45500.0 ;
      RECT  100350.0 46845.0 101055.0 48190.0 ;
      RECT  100350.0 49535.0 101055.0 48190.0 ;
      RECT  100350.0 49535.0 101055.0 50880.0 ;
      RECT  100350.0 52225.0 101055.0 50880.0 ;
      RECT  100350.0 52225.0 101055.0 53570.0 ;
      RECT  100350.0 54915.0 101055.0 53570.0 ;
      RECT  100350.0 54915.0 101055.0 56260.0 ;
      RECT  100350.0 57605.0 101055.0 56260.0 ;
      RECT  100350.0 57605.0 101055.0 58950.0 ;
      RECT  100350.0 60295.0 101055.0 58950.0 ;
      RECT  100350.0 60295.0 101055.0 61640.0 ;
      RECT  100350.0 62985.0 101055.0 61640.0 ;
      RECT  100350.0 62985.0 101055.0 64330.0 ;
      RECT  100350.0 65675.0 101055.0 64330.0 ;
      RECT  100350.0 65675.0 101055.0 67020.0 ;
      RECT  100350.0 68365.0 101055.0 67020.0 ;
      RECT  100350.0 68365.0 101055.0 69710.0 ;
      RECT  100350.0 71055.0 101055.0 69710.0 ;
      RECT  100350.0 71055.0 101055.0 72400.0 ;
      RECT  100350.0 73745.0 101055.0 72400.0 ;
      RECT  100350.0 73745.0 101055.0 75090.0 ;
      RECT  100350.0 76435.0 101055.0 75090.0 ;
      RECT  100350.0 76435.0 101055.0 77780.0 ;
      RECT  100350.0 79125.0 101055.0 77780.0 ;
      RECT  100350.0 79125.0 101055.0 80470.0 ;
      RECT  100350.0 81815.0 101055.0 80470.0 ;
      RECT  100350.0 81815.0 101055.0 83160.0 ;
      RECT  100350.0 84505.0 101055.0 83160.0 ;
      RECT  100350.0 84505.0 101055.0 85850.0 ;
      RECT  100350.0 87195.0 101055.0 85850.0 ;
      RECT  100350.0 87195.0 101055.0 88540.0 ;
      RECT  100350.0 89885.0 101055.0 88540.0 ;
      RECT  100350.0 89885.0 101055.0 91230.0 ;
      RECT  100350.0 92575.0 101055.0 91230.0 ;
      RECT  100350.0 92575.0 101055.0 93920.0 ;
      RECT  100350.0 95265.0 101055.0 93920.0 ;
      RECT  100350.0 95265.0 101055.0 96610.0 ;
      RECT  100350.0 97955.0 101055.0 96610.0 ;
      RECT  100350.0 97955.0 101055.0 99300.0 ;
      RECT  100350.0 100645.0 101055.0 99300.0 ;
      RECT  100350.0 100645.0 101055.0 101990.0 ;
      RECT  100350.0 103335.0 101055.0 101990.0 ;
      RECT  100350.0 103335.0 101055.0 104680.0 ;
      RECT  100350.0 106025.0 101055.0 104680.0 ;
      RECT  100350.0 106025.0 101055.0 107370.0 ;
      RECT  100350.0 108715.0 101055.0 107370.0 ;
      RECT  100350.0 108715.0 101055.0 110060.0 ;
      RECT  100350.0 111405.0 101055.0 110060.0 ;
      RECT  100350.0 111405.0 101055.0 112750.0 ;
      RECT  100350.0 114095.0 101055.0 112750.0 ;
      RECT  101055.0 28015.0 101760.0 29360.0 ;
      RECT  101055.0 30705.0 101760.0 29360.0 ;
      RECT  101055.0 30705.0 101760.0 32050.0 ;
      RECT  101055.0 33395.0 101760.0 32050.0 ;
      RECT  101055.0 33395.0 101760.0 34740.0 ;
      RECT  101055.0 36085.0 101760.0 34740.0 ;
      RECT  101055.0 36085.0 101760.0 37430.0 ;
      RECT  101055.0 38775.0 101760.0 37430.0 ;
      RECT  101055.0 38775.0 101760.0 40120.0 ;
      RECT  101055.0 41465.0 101760.0 40120.0 ;
      RECT  101055.0 41465.0 101760.0 42810.0 ;
      RECT  101055.0 44155.0 101760.0 42810.0 ;
      RECT  101055.0 44155.0 101760.0 45500.0 ;
      RECT  101055.0 46845.0 101760.0 45500.0 ;
      RECT  101055.0 46845.0 101760.0 48190.0 ;
      RECT  101055.0 49535.0 101760.0 48190.0 ;
      RECT  101055.0 49535.0 101760.0 50880.0 ;
      RECT  101055.0 52225.0 101760.0 50880.0 ;
      RECT  101055.0 52225.0 101760.0 53570.0 ;
      RECT  101055.0 54915.0 101760.0 53570.0 ;
      RECT  101055.0 54915.0 101760.0 56260.0 ;
      RECT  101055.0 57605.0 101760.0 56260.0 ;
      RECT  101055.0 57605.0 101760.0 58950.0 ;
      RECT  101055.0 60295.0 101760.0 58950.0 ;
      RECT  101055.0 60295.0 101760.0 61640.0 ;
      RECT  101055.0 62985.0 101760.0 61640.0 ;
      RECT  101055.0 62985.0 101760.0 64330.0 ;
      RECT  101055.0 65675.0 101760.0 64330.0 ;
      RECT  101055.0 65675.0 101760.0 67020.0 ;
      RECT  101055.0 68365.0 101760.0 67020.0 ;
      RECT  101055.0 68365.0 101760.0 69710.0 ;
      RECT  101055.0 71055.0 101760.0 69710.0 ;
      RECT  101055.0 71055.0 101760.0 72400.0 ;
      RECT  101055.0 73745.0 101760.0 72400.0 ;
      RECT  101055.0 73745.0 101760.0 75090.0 ;
      RECT  101055.0 76435.0 101760.0 75090.0 ;
      RECT  101055.0 76435.0 101760.0 77780.0 ;
      RECT  101055.0 79125.0 101760.0 77780.0 ;
      RECT  101055.0 79125.0 101760.0 80470.0 ;
      RECT  101055.0 81815.0 101760.0 80470.0 ;
      RECT  101055.0 81815.0 101760.0 83160.0 ;
      RECT  101055.0 84505.0 101760.0 83160.0 ;
      RECT  101055.0 84505.0 101760.0 85850.0 ;
      RECT  101055.0 87195.0 101760.0 85850.0 ;
      RECT  101055.0 87195.0 101760.0 88540.0 ;
      RECT  101055.0 89885.0 101760.0 88540.0 ;
      RECT  101055.0 89885.0 101760.0 91230.0 ;
      RECT  101055.0 92575.0 101760.0 91230.0 ;
      RECT  101055.0 92575.0 101760.0 93920.0 ;
      RECT  101055.0 95265.0 101760.0 93920.0 ;
      RECT  101055.0 95265.0 101760.0 96610.0 ;
      RECT  101055.0 97955.0 101760.0 96610.0 ;
      RECT  101055.0 97955.0 101760.0 99300.0 ;
      RECT  101055.0 100645.0 101760.0 99300.0 ;
      RECT  101055.0 100645.0 101760.0 101990.0 ;
      RECT  101055.0 103335.0 101760.0 101990.0 ;
      RECT  101055.0 103335.0 101760.0 104680.0 ;
      RECT  101055.0 106025.0 101760.0 104680.0 ;
      RECT  101055.0 106025.0 101760.0 107370.0 ;
      RECT  101055.0 108715.0 101760.0 107370.0 ;
      RECT  101055.0 108715.0 101760.0 110060.0 ;
      RECT  101055.0 111405.0 101760.0 110060.0 ;
      RECT  101055.0 111405.0 101760.0 112750.0 ;
      RECT  101055.0 114095.0 101760.0 112750.0 ;
      RECT  101760.0 28015.0 102465.0 29360.0 ;
      RECT  101760.0 30705.0 102465.0 29360.0 ;
      RECT  101760.0 30705.0 102465.0 32050.0 ;
      RECT  101760.0 33395.0 102465.0 32050.0 ;
      RECT  101760.0 33395.0 102465.0 34740.0 ;
      RECT  101760.0 36085.0 102465.0 34740.0 ;
      RECT  101760.0 36085.0 102465.0 37430.0 ;
      RECT  101760.0 38775.0 102465.0 37430.0 ;
      RECT  101760.0 38775.0 102465.0 40120.0 ;
      RECT  101760.0 41465.0 102465.0 40120.0 ;
      RECT  101760.0 41465.0 102465.0 42810.0 ;
      RECT  101760.0 44155.0 102465.0 42810.0 ;
      RECT  101760.0 44155.0 102465.0 45500.0 ;
      RECT  101760.0 46845.0 102465.0 45500.0 ;
      RECT  101760.0 46845.0 102465.0 48190.0 ;
      RECT  101760.0 49535.0 102465.0 48190.0 ;
      RECT  101760.0 49535.0 102465.0 50880.0 ;
      RECT  101760.0 52225.0 102465.0 50880.0 ;
      RECT  101760.0 52225.0 102465.0 53570.0 ;
      RECT  101760.0 54915.0 102465.0 53570.0 ;
      RECT  101760.0 54915.0 102465.0 56260.0 ;
      RECT  101760.0 57605.0 102465.0 56260.0 ;
      RECT  101760.0 57605.0 102465.0 58950.0 ;
      RECT  101760.0 60295.0 102465.0 58950.0 ;
      RECT  101760.0 60295.0 102465.0 61640.0 ;
      RECT  101760.0 62985.0 102465.0 61640.0 ;
      RECT  101760.0 62985.0 102465.0 64330.0 ;
      RECT  101760.0 65675.0 102465.0 64330.0 ;
      RECT  101760.0 65675.0 102465.0 67020.0 ;
      RECT  101760.0 68365.0 102465.0 67020.0 ;
      RECT  101760.0 68365.0 102465.0 69710.0 ;
      RECT  101760.0 71055.0 102465.0 69710.0 ;
      RECT  101760.0 71055.0 102465.0 72400.0 ;
      RECT  101760.0 73745.0 102465.0 72400.0 ;
      RECT  101760.0 73745.0 102465.0 75090.0 ;
      RECT  101760.0 76435.0 102465.0 75090.0 ;
      RECT  101760.0 76435.0 102465.0 77780.0 ;
      RECT  101760.0 79125.0 102465.0 77780.0 ;
      RECT  101760.0 79125.0 102465.0 80470.0 ;
      RECT  101760.0 81815.0 102465.0 80470.0 ;
      RECT  101760.0 81815.0 102465.0 83160.0 ;
      RECT  101760.0 84505.0 102465.0 83160.0 ;
      RECT  101760.0 84505.0 102465.0 85850.0 ;
      RECT  101760.0 87195.0 102465.0 85850.0 ;
      RECT  101760.0 87195.0 102465.0 88540.0 ;
      RECT  101760.0 89885.0 102465.0 88540.0 ;
      RECT  101760.0 89885.0 102465.0 91230.0 ;
      RECT  101760.0 92575.0 102465.0 91230.0 ;
      RECT  101760.0 92575.0 102465.0 93920.0 ;
      RECT  101760.0 95265.0 102465.0 93920.0 ;
      RECT  101760.0 95265.0 102465.0 96610.0 ;
      RECT  101760.0 97955.0 102465.0 96610.0 ;
      RECT  101760.0 97955.0 102465.0 99300.0 ;
      RECT  101760.0 100645.0 102465.0 99300.0 ;
      RECT  101760.0 100645.0 102465.0 101990.0 ;
      RECT  101760.0 103335.0 102465.0 101990.0 ;
      RECT  101760.0 103335.0 102465.0 104680.0 ;
      RECT  101760.0 106025.0 102465.0 104680.0 ;
      RECT  101760.0 106025.0 102465.0 107370.0 ;
      RECT  101760.0 108715.0 102465.0 107370.0 ;
      RECT  101760.0 108715.0 102465.0 110060.0 ;
      RECT  101760.0 111405.0 102465.0 110060.0 ;
      RECT  101760.0 111405.0 102465.0 112750.0 ;
      RECT  101760.0 114095.0 102465.0 112750.0 ;
      RECT  102465.0 28015.0 103170.0 29360.0 ;
      RECT  102465.0 30705.0 103170.0 29360.0 ;
      RECT  102465.0 30705.0 103170.0 32050.0 ;
      RECT  102465.0 33395.0 103170.0 32050.0 ;
      RECT  102465.0 33395.0 103170.0 34740.0 ;
      RECT  102465.0 36085.0 103170.0 34740.0 ;
      RECT  102465.0 36085.0 103170.0 37430.0 ;
      RECT  102465.0 38775.0 103170.0 37430.0 ;
      RECT  102465.0 38775.0 103170.0 40120.0 ;
      RECT  102465.0 41465.0 103170.0 40120.0 ;
      RECT  102465.0 41465.0 103170.0 42810.0 ;
      RECT  102465.0 44155.0 103170.0 42810.0 ;
      RECT  102465.0 44155.0 103170.0 45500.0 ;
      RECT  102465.0 46845.0 103170.0 45500.0 ;
      RECT  102465.0 46845.0 103170.0 48190.0 ;
      RECT  102465.0 49535.0 103170.0 48190.0 ;
      RECT  102465.0 49535.0 103170.0 50880.0 ;
      RECT  102465.0 52225.0 103170.0 50880.0 ;
      RECT  102465.0 52225.0 103170.0 53570.0 ;
      RECT  102465.0 54915.0 103170.0 53570.0 ;
      RECT  102465.0 54915.0 103170.0 56260.0 ;
      RECT  102465.0 57605.0 103170.0 56260.0 ;
      RECT  102465.0 57605.0 103170.0 58950.0 ;
      RECT  102465.0 60295.0 103170.0 58950.0 ;
      RECT  102465.0 60295.0 103170.0 61640.0 ;
      RECT  102465.0 62985.0 103170.0 61640.0 ;
      RECT  102465.0 62985.0 103170.0 64330.0 ;
      RECT  102465.0 65675.0 103170.0 64330.0 ;
      RECT  102465.0 65675.0 103170.0 67020.0 ;
      RECT  102465.0 68365.0 103170.0 67020.0 ;
      RECT  102465.0 68365.0 103170.0 69710.0 ;
      RECT  102465.0 71055.0 103170.0 69710.0 ;
      RECT  102465.0 71055.0 103170.0 72400.0 ;
      RECT  102465.0 73745.0 103170.0 72400.0 ;
      RECT  102465.0 73745.0 103170.0 75090.0 ;
      RECT  102465.0 76435.0 103170.0 75090.0 ;
      RECT  102465.0 76435.0 103170.0 77780.0 ;
      RECT  102465.0 79125.0 103170.0 77780.0 ;
      RECT  102465.0 79125.0 103170.0 80470.0 ;
      RECT  102465.0 81815.0 103170.0 80470.0 ;
      RECT  102465.0 81815.0 103170.0 83160.0 ;
      RECT  102465.0 84505.0 103170.0 83160.0 ;
      RECT  102465.0 84505.0 103170.0 85850.0 ;
      RECT  102465.0 87195.0 103170.0 85850.0 ;
      RECT  102465.0 87195.0 103170.0 88540.0 ;
      RECT  102465.0 89885.0 103170.0 88540.0 ;
      RECT  102465.0 89885.0 103170.0 91230.0 ;
      RECT  102465.0 92575.0 103170.0 91230.0 ;
      RECT  102465.0 92575.0 103170.0 93920.0 ;
      RECT  102465.0 95265.0 103170.0 93920.0 ;
      RECT  102465.0 95265.0 103170.0 96610.0 ;
      RECT  102465.0 97955.0 103170.0 96610.0 ;
      RECT  102465.0 97955.0 103170.0 99300.0 ;
      RECT  102465.0 100645.0 103170.0 99300.0 ;
      RECT  102465.0 100645.0 103170.0 101990.0 ;
      RECT  102465.0 103335.0 103170.0 101990.0 ;
      RECT  102465.0 103335.0 103170.0 104680.0 ;
      RECT  102465.0 106025.0 103170.0 104680.0 ;
      RECT  102465.0 106025.0 103170.0 107370.0 ;
      RECT  102465.0 108715.0 103170.0 107370.0 ;
      RECT  102465.0 108715.0 103170.0 110060.0 ;
      RECT  102465.0 111405.0 103170.0 110060.0 ;
      RECT  102465.0 111405.0 103170.0 112750.0 ;
      RECT  102465.0 114095.0 103170.0 112750.0 ;
      RECT  103170.0 28015.0 103875.0 29360.0 ;
      RECT  103170.0 30705.0 103875.0 29360.0 ;
      RECT  103170.0 30705.0 103875.0 32050.0 ;
      RECT  103170.0 33395.0 103875.0 32050.0 ;
      RECT  103170.0 33395.0 103875.0 34740.0 ;
      RECT  103170.0 36085.0 103875.0 34740.0 ;
      RECT  103170.0 36085.0 103875.0 37430.0 ;
      RECT  103170.0 38775.0 103875.0 37430.0 ;
      RECT  103170.0 38775.0 103875.0 40120.0 ;
      RECT  103170.0 41465.0 103875.0 40120.0 ;
      RECT  103170.0 41465.0 103875.0 42810.0 ;
      RECT  103170.0 44155.0 103875.0 42810.0 ;
      RECT  103170.0 44155.0 103875.0 45500.0 ;
      RECT  103170.0 46845.0 103875.0 45500.0 ;
      RECT  103170.0 46845.0 103875.0 48190.0 ;
      RECT  103170.0 49535.0 103875.0 48190.0 ;
      RECT  103170.0 49535.0 103875.0 50880.0 ;
      RECT  103170.0 52225.0 103875.0 50880.0 ;
      RECT  103170.0 52225.0 103875.0 53570.0 ;
      RECT  103170.0 54915.0 103875.0 53570.0 ;
      RECT  103170.0 54915.0 103875.0 56260.0 ;
      RECT  103170.0 57605.0 103875.0 56260.0 ;
      RECT  103170.0 57605.0 103875.0 58950.0 ;
      RECT  103170.0 60295.0 103875.0 58950.0 ;
      RECT  103170.0 60295.0 103875.0 61640.0 ;
      RECT  103170.0 62985.0 103875.0 61640.0 ;
      RECT  103170.0 62985.0 103875.0 64330.0 ;
      RECT  103170.0 65675.0 103875.0 64330.0 ;
      RECT  103170.0 65675.0 103875.0 67020.0 ;
      RECT  103170.0 68365.0 103875.0 67020.0 ;
      RECT  103170.0 68365.0 103875.0 69710.0 ;
      RECT  103170.0 71055.0 103875.0 69710.0 ;
      RECT  103170.0 71055.0 103875.0 72400.0 ;
      RECT  103170.0 73745.0 103875.0 72400.0 ;
      RECT  103170.0 73745.0 103875.0 75090.0 ;
      RECT  103170.0 76435.0 103875.0 75090.0 ;
      RECT  103170.0 76435.0 103875.0 77780.0 ;
      RECT  103170.0 79125.0 103875.0 77780.0 ;
      RECT  103170.0 79125.0 103875.0 80470.0 ;
      RECT  103170.0 81815.0 103875.0 80470.0 ;
      RECT  103170.0 81815.0 103875.0 83160.0 ;
      RECT  103170.0 84505.0 103875.0 83160.0 ;
      RECT  103170.0 84505.0 103875.0 85850.0 ;
      RECT  103170.0 87195.0 103875.0 85850.0 ;
      RECT  103170.0 87195.0 103875.0 88540.0 ;
      RECT  103170.0 89885.0 103875.0 88540.0 ;
      RECT  103170.0 89885.0 103875.0 91230.0 ;
      RECT  103170.0 92575.0 103875.0 91230.0 ;
      RECT  103170.0 92575.0 103875.0 93920.0 ;
      RECT  103170.0 95265.0 103875.0 93920.0 ;
      RECT  103170.0 95265.0 103875.0 96610.0 ;
      RECT  103170.0 97955.0 103875.0 96610.0 ;
      RECT  103170.0 97955.0 103875.0 99300.0 ;
      RECT  103170.0 100645.0 103875.0 99300.0 ;
      RECT  103170.0 100645.0 103875.0 101990.0 ;
      RECT  103170.0 103335.0 103875.0 101990.0 ;
      RECT  103170.0 103335.0 103875.0 104680.0 ;
      RECT  103170.0 106025.0 103875.0 104680.0 ;
      RECT  103170.0 106025.0 103875.0 107370.0 ;
      RECT  103170.0 108715.0 103875.0 107370.0 ;
      RECT  103170.0 108715.0 103875.0 110060.0 ;
      RECT  103170.0 111405.0 103875.0 110060.0 ;
      RECT  103170.0 111405.0 103875.0 112750.0 ;
      RECT  103170.0 114095.0 103875.0 112750.0 ;
      RECT  103875.0 28015.0 104580.0 29360.0 ;
      RECT  103875.0 30705.0 104580.0 29360.0 ;
      RECT  103875.0 30705.0 104580.0 32050.0 ;
      RECT  103875.0 33395.0 104580.0 32050.0 ;
      RECT  103875.0 33395.0 104580.0 34740.0 ;
      RECT  103875.0 36085.0 104580.0 34740.0 ;
      RECT  103875.0 36085.0 104580.0 37430.0 ;
      RECT  103875.0 38775.0 104580.0 37430.0 ;
      RECT  103875.0 38775.0 104580.0 40120.0 ;
      RECT  103875.0 41465.0 104580.0 40120.0 ;
      RECT  103875.0 41465.0 104580.0 42810.0 ;
      RECT  103875.0 44155.0 104580.0 42810.0 ;
      RECT  103875.0 44155.0 104580.0 45500.0 ;
      RECT  103875.0 46845.0 104580.0 45500.0 ;
      RECT  103875.0 46845.0 104580.0 48190.0 ;
      RECT  103875.0 49535.0 104580.0 48190.0 ;
      RECT  103875.0 49535.0 104580.0 50880.0 ;
      RECT  103875.0 52225.0 104580.0 50880.0 ;
      RECT  103875.0 52225.0 104580.0 53570.0 ;
      RECT  103875.0 54915.0 104580.0 53570.0 ;
      RECT  103875.0 54915.0 104580.0 56260.0 ;
      RECT  103875.0 57605.0 104580.0 56260.0 ;
      RECT  103875.0 57605.0 104580.0 58950.0 ;
      RECT  103875.0 60295.0 104580.0 58950.0 ;
      RECT  103875.0 60295.0 104580.0 61640.0 ;
      RECT  103875.0 62985.0 104580.0 61640.0 ;
      RECT  103875.0 62985.0 104580.0 64330.0 ;
      RECT  103875.0 65675.0 104580.0 64330.0 ;
      RECT  103875.0 65675.0 104580.0 67020.0 ;
      RECT  103875.0 68365.0 104580.0 67020.0 ;
      RECT  103875.0 68365.0 104580.0 69710.0 ;
      RECT  103875.0 71055.0 104580.0 69710.0 ;
      RECT  103875.0 71055.0 104580.0 72400.0 ;
      RECT  103875.0 73745.0 104580.0 72400.0 ;
      RECT  103875.0 73745.0 104580.0 75090.0 ;
      RECT  103875.0 76435.0 104580.0 75090.0 ;
      RECT  103875.0 76435.0 104580.0 77780.0 ;
      RECT  103875.0 79125.0 104580.0 77780.0 ;
      RECT  103875.0 79125.0 104580.0 80470.0 ;
      RECT  103875.0 81815.0 104580.0 80470.0 ;
      RECT  103875.0 81815.0 104580.0 83160.0 ;
      RECT  103875.0 84505.0 104580.0 83160.0 ;
      RECT  103875.0 84505.0 104580.0 85850.0 ;
      RECT  103875.0 87195.0 104580.0 85850.0 ;
      RECT  103875.0 87195.0 104580.0 88540.0 ;
      RECT  103875.0 89885.0 104580.0 88540.0 ;
      RECT  103875.0 89885.0 104580.0 91230.0 ;
      RECT  103875.0 92575.0 104580.0 91230.0 ;
      RECT  103875.0 92575.0 104580.0 93920.0 ;
      RECT  103875.0 95265.0 104580.0 93920.0 ;
      RECT  103875.0 95265.0 104580.0 96610.0 ;
      RECT  103875.0 97955.0 104580.0 96610.0 ;
      RECT  103875.0 97955.0 104580.0 99300.0 ;
      RECT  103875.0 100645.0 104580.0 99300.0 ;
      RECT  103875.0 100645.0 104580.0 101990.0 ;
      RECT  103875.0 103335.0 104580.0 101990.0 ;
      RECT  103875.0 103335.0 104580.0 104680.0 ;
      RECT  103875.0 106025.0 104580.0 104680.0 ;
      RECT  103875.0 106025.0 104580.0 107370.0 ;
      RECT  103875.0 108715.0 104580.0 107370.0 ;
      RECT  103875.0 108715.0 104580.0 110060.0 ;
      RECT  103875.0 111405.0 104580.0 110060.0 ;
      RECT  103875.0 111405.0 104580.0 112750.0 ;
      RECT  103875.0 114095.0 104580.0 112750.0 ;
      RECT  104580.0 28015.0 105285.0 29360.0 ;
      RECT  104580.0 30705.0 105285.0 29360.0 ;
      RECT  104580.0 30705.0 105285.0 32050.0 ;
      RECT  104580.0 33395.0 105285.0 32050.0 ;
      RECT  104580.0 33395.0 105285.0 34740.0 ;
      RECT  104580.0 36085.0 105285.0 34740.0 ;
      RECT  104580.0 36085.0 105285.0 37430.0 ;
      RECT  104580.0 38775.0 105285.0 37430.0 ;
      RECT  104580.0 38775.0 105285.0 40120.0 ;
      RECT  104580.0 41465.0 105285.0 40120.0 ;
      RECT  104580.0 41465.0 105285.0 42810.0 ;
      RECT  104580.0 44155.0 105285.0 42810.0 ;
      RECT  104580.0 44155.0 105285.0 45500.0 ;
      RECT  104580.0 46845.0 105285.0 45500.0 ;
      RECT  104580.0 46845.0 105285.0 48190.0 ;
      RECT  104580.0 49535.0 105285.0 48190.0 ;
      RECT  104580.0 49535.0 105285.0 50880.0 ;
      RECT  104580.0 52225.0 105285.0 50880.0 ;
      RECT  104580.0 52225.0 105285.0 53570.0 ;
      RECT  104580.0 54915.0 105285.0 53570.0 ;
      RECT  104580.0 54915.0 105285.0 56260.0 ;
      RECT  104580.0 57605.0 105285.0 56260.0 ;
      RECT  104580.0 57605.0 105285.0 58950.0 ;
      RECT  104580.0 60295.0 105285.0 58950.0 ;
      RECT  104580.0 60295.0 105285.0 61640.0 ;
      RECT  104580.0 62985.0 105285.0 61640.0 ;
      RECT  104580.0 62985.0 105285.0 64330.0 ;
      RECT  104580.0 65675.0 105285.0 64330.0 ;
      RECT  104580.0 65675.0 105285.0 67020.0 ;
      RECT  104580.0 68365.0 105285.0 67020.0 ;
      RECT  104580.0 68365.0 105285.0 69710.0 ;
      RECT  104580.0 71055.0 105285.0 69710.0 ;
      RECT  104580.0 71055.0 105285.0 72400.0 ;
      RECT  104580.0 73745.0 105285.0 72400.0 ;
      RECT  104580.0 73745.0 105285.0 75090.0 ;
      RECT  104580.0 76435.0 105285.0 75090.0 ;
      RECT  104580.0 76435.0 105285.0 77780.0 ;
      RECT  104580.0 79125.0 105285.0 77780.0 ;
      RECT  104580.0 79125.0 105285.0 80470.0 ;
      RECT  104580.0 81815.0 105285.0 80470.0 ;
      RECT  104580.0 81815.0 105285.0 83160.0 ;
      RECT  104580.0 84505.0 105285.0 83160.0 ;
      RECT  104580.0 84505.0 105285.0 85850.0 ;
      RECT  104580.0 87195.0 105285.0 85850.0 ;
      RECT  104580.0 87195.0 105285.0 88540.0 ;
      RECT  104580.0 89885.0 105285.0 88540.0 ;
      RECT  104580.0 89885.0 105285.0 91230.0 ;
      RECT  104580.0 92575.0 105285.0 91230.0 ;
      RECT  104580.0 92575.0 105285.0 93920.0 ;
      RECT  104580.0 95265.0 105285.0 93920.0 ;
      RECT  104580.0 95265.0 105285.0 96610.0 ;
      RECT  104580.0 97955.0 105285.0 96610.0 ;
      RECT  104580.0 97955.0 105285.0 99300.0 ;
      RECT  104580.0 100645.0 105285.0 99300.0 ;
      RECT  104580.0 100645.0 105285.0 101990.0 ;
      RECT  104580.0 103335.0 105285.0 101990.0 ;
      RECT  104580.0 103335.0 105285.0 104680.0 ;
      RECT  104580.0 106025.0 105285.0 104680.0 ;
      RECT  104580.0 106025.0 105285.0 107370.0 ;
      RECT  104580.0 108715.0 105285.0 107370.0 ;
      RECT  104580.0 108715.0 105285.0 110060.0 ;
      RECT  104580.0 111405.0 105285.0 110060.0 ;
      RECT  104580.0 111405.0 105285.0 112750.0 ;
      RECT  104580.0 114095.0 105285.0 112750.0 ;
      RECT  105285.0 28015.0 105990.0 29360.0 ;
      RECT  105285.0 30705.0 105990.0 29360.0 ;
      RECT  105285.0 30705.0 105990.0 32050.0 ;
      RECT  105285.0 33395.0 105990.0 32050.0 ;
      RECT  105285.0 33395.0 105990.0 34740.0 ;
      RECT  105285.0 36085.0 105990.0 34740.0 ;
      RECT  105285.0 36085.0 105990.0 37430.0 ;
      RECT  105285.0 38775.0 105990.0 37430.0 ;
      RECT  105285.0 38775.0 105990.0 40120.0 ;
      RECT  105285.0 41465.0 105990.0 40120.0 ;
      RECT  105285.0 41465.0 105990.0 42810.0 ;
      RECT  105285.0 44155.0 105990.0 42810.0 ;
      RECT  105285.0 44155.0 105990.0 45500.0 ;
      RECT  105285.0 46845.0 105990.0 45500.0 ;
      RECT  105285.0 46845.0 105990.0 48190.0 ;
      RECT  105285.0 49535.0 105990.0 48190.0 ;
      RECT  105285.0 49535.0 105990.0 50880.0 ;
      RECT  105285.0 52225.0 105990.0 50880.0 ;
      RECT  105285.0 52225.0 105990.0 53570.0 ;
      RECT  105285.0 54915.0 105990.0 53570.0 ;
      RECT  105285.0 54915.0 105990.0 56260.0 ;
      RECT  105285.0 57605.0 105990.0 56260.0 ;
      RECT  105285.0 57605.0 105990.0 58950.0 ;
      RECT  105285.0 60295.0 105990.0 58950.0 ;
      RECT  105285.0 60295.0 105990.0 61640.0 ;
      RECT  105285.0 62985.0 105990.0 61640.0 ;
      RECT  105285.0 62985.0 105990.0 64330.0 ;
      RECT  105285.0 65675.0 105990.0 64330.0 ;
      RECT  105285.0 65675.0 105990.0 67020.0 ;
      RECT  105285.0 68365.0 105990.0 67020.0 ;
      RECT  105285.0 68365.0 105990.0 69710.0 ;
      RECT  105285.0 71055.0 105990.0 69710.0 ;
      RECT  105285.0 71055.0 105990.0 72400.0 ;
      RECT  105285.0 73745.0 105990.0 72400.0 ;
      RECT  105285.0 73745.0 105990.0 75090.0 ;
      RECT  105285.0 76435.0 105990.0 75090.0 ;
      RECT  105285.0 76435.0 105990.0 77780.0 ;
      RECT  105285.0 79125.0 105990.0 77780.0 ;
      RECT  105285.0 79125.0 105990.0 80470.0 ;
      RECT  105285.0 81815.0 105990.0 80470.0 ;
      RECT  105285.0 81815.0 105990.0 83160.0 ;
      RECT  105285.0 84505.0 105990.0 83160.0 ;
      RECT  105285.0 84505.0 105990.0 85850.0 ;
      RECT  105285.0 87195.0 105990.0 85850.0 ;
      RECT  105285.0 87195.0 105990.0 88540.0 ;
      RECT  105285.0 89885.0 105990.0 88540.0 ;
      RECT  105285.0 89885.0 105990.0 91230.0 ;
      RECT  105285.0 92575.0 105990.0 91230.0 ;
      RECT  105285.0 92575.0 105990.0 93920.0 ;
      RECT  105285.0 95265.0 105990.0 93920.0 ;
      RECT  105285.0 95265.0 105990.0 96610.0 ;
      RECT  105285.0 97955.0 105990.0 96610.0 ;
      RECT  105285.0 97955.0 105990.0 99300.0 ;
      RECT  105285.0 100645.0 105990.0 99300.0 ;
      RECT  105285.0 100645.0 105990.0 101990.0 ;
      RECT  105285.0 103335.0 105990.0 101990.0 ;
      RECT  105285.0 103335.0 105990.0 104680.0 ;
      RECT  105285.0 106025.0 105990.0 104680.0 ;
      RECT  105285.0 106025.0 105990.0 107370.0 ;
      RECT  105285.0 108715.0 105990.0 107370.0 ;
      RECT  105285.0 108715.0 105990.0 110060.0 ;
      RECT  105285.0 111405.0 105990.0 110060.0 ;
      RECT  105285.0 111405.0 105990.0 112750.0 ;
      RECT  105285.0 114095.0 105990.0 112750.0 ;
      RECT  15660.0 28122.5 106080.0 28187.5 ;
      RECT  15660.0 30532.5 106080.0 30597.5 ;
      RECT  15660.0 30812.5 106080.0 30877.5 ;
      RECT  15660.0 33222.5 106080.0 33287.5 ;
      RECT  15660.0 33502.5 106080.0 33567.5 ;
      RECT  15660.0 35912.5 106080.0 35977.5 ;
      RECT  15660.0 36192.5 106080.0 36257.5 ;
      RECT  15660.0 38602.5 106080.0 38667.5 ;
      RECT  15660.0 38882.5 106080.0 38947.5 ;
      RECT  15660.0 41292.5 106080.0 41357.5 ;
      RECT  15660.0 41572.5 106080.0 41637.5 ;
      RECT  15660.0 43982.5 106080.0 44047.5 ;
      RECT  15660.0 44262.5 106080.0 44327.5 ;
      RECT  15660.0 46672.5 106080.0 46737.5 ;
      RECT  15660.0 46952.5 106080.0 47017.5 ;
      RECT  15660.0 49362.5 106080.0 49427.5 ;
      RECT  15660.0 49642.5 106080.0 49707.5 ;
      RECT  15660.0 52052.5 106080.0 52117.5 ;
      RECT  15660.0 52332.5 106080.0 52397.5 ;
      RECT  15660.0 54742.5 106080.0 54807.5 ;
      RECT  15660.0 55022.5 106080.0 55087.5 ;
      RECT  15660.0 57432.5 106080.0 57497.5 ;
      RECT  15660.0 57712.5 106080.0 57777.5 ;
      RECT  15660.0 60122.5 106080.0 60187.5 ;
      RECT  15660.0 60402.5 106080.0 60467.5 ;
      RECT  15660.0 62812.5 106080.0 62877.5 ;
      RECT  15660.0 63092.5 106080.0 63157.5 ;
      RECT  15660.0 65502.5 106080.0 65567.5 ;
      RECT  15660.0 65782.5 106080.0 65847.5 ;
      RECT  15660.0 68192.5 106080.0 68257.5 ;
      RECT  15660.0 68472.5 106080.0 68537.5 ;
      RECT  15660.0 70882.5 106080.0 70947.5 ;
      RECT  15660.0 71162.5 106080.0 71227.5 ;
      RECT  15660.0 73572.5 106080.0 73637.5 ;
      RECT  15660.0 73852.5 106080.0 73917.5 ;
      RECT  15660.0 76262.5 106080.0 76327.5 ;
      RECT  15660.0 76542.5 106080.0 76607.5 ;
      RECT  15660.0 78952.5 106080.0 79017.5 ;
      RECT  15660.0 79232.5 106080.0 79297.5 ;
      RECT  15660.0 81642.5 106080.0 81707.5 ;
      RECT  15660.0 81922.5 106080.0 81987.5 ;
      RECT  15660.0 84332.5 106080.0 84397.5 ;
      RECT  15660.0 84612.5 106080.0 84677.5 ;
      RECT  15660.0 87022.5 106080.0 87087.5 ;
      RECT  15660.0 87302.5 106080.0 87367.5 ;
      RECT  15660.0 89712.5 106080.0 89777.5 ;
      RECT  15660.0 89992.5 106080.0 90057.5 ;
      RECT  15660.0 92402.5 106080.0 92467.5 ;
      RECT  15660.0 92682.5 106080.0 92747.5 ;
      RECT  15660.0 95092.5 106080.0 95157.5 ;
      RECT  15660.0 95372.5 106080.0 95437.5 ;
      RECT  15660.0 97782.5 106080.0 97847.5 ;
      RECT  15660.0 98062.5 106080.0 98127.5 ;
      RECT  15660.0 100472.5 106080.0 100537.5 ;
      RECT  15660.0 100752.5 106080.0 100817.5 ;
      RECT  15660.0 103162.5 106080.0 103227.5 ;
      RECT  15660.0 103442.5 106080.0 103507.5 ;
      RECT  15660.0 105852.5 106080.0 105917.5 ;
      RECT  15660.0 106132.5 106080.0 106197.5 ;
      RECT  15660.0 108542.5 106080.0 108607.5 ;
      RECT  15660.0 108822.5 106080.0 108887.5 ;
      RECT  15660.0 111232.5 106080.0 111297.5 ;
      RECT  15660.0 111512.5 106080.0 111577.5 ;
      RECT  15660.0 113922.5 106080.0 113987.5 ;
      RECT  15660.0 29327.5 106080.0 29392.5 ;
      RECT  15660.0 32017.5 106080.0 32082.5 ;
      RECT  15660.0 34707.5 106080.0 34772.5 ;
      RECT  15660.0 37397.5 106080.0 37462.5 ;
      RECT  15660.0 40087.5 106080.0 40152.5 ;
      RECT  15660.0 42777.5 106080.0 42842.5 ;
      RECT  15660.0 45467.5 106080.0 45532.5 ;
      RECT  15660.0 48157.5 106080.0 48222.5 ;
      RECT  15660.0 50847.5 106080.0 50912.5 ;
      RECT  15660.0 53537.5 106080.0 53602.5 ;
      RECT  15660.0 56227.5 106080.0 56292.5 ;
      RECT  15660.0 58917.5 106080.0 58982.5 ;
      RECT  15660.0 61607.5 106080.0 61672.5 ;
      RECT  15660.0 64297.5 106080.0 64362.5 ;
      RECT  15660.0 66987.5 106080.0 67052.5 ;
      RECT  15660.0 69677.5 106080.0 69742.5 ;
      RECT  15660.0 72367.5 106080.0 72432.5 ;
      RECT  15660.0 75057.5 106080.0 75122.5 ;
      RECT  15660.0 77747.5 106080.0 77812.5 ;
      RECT  15660.0 80437.5 106080.0 80502.5 ;
      RECT  15660.0 83127.5 106080.0 83192.5 ;
      RECT  15660.0 85817.5 106080.0 85882.5 ;
      RECT  15660.0 88507.5 106080.0 88572.5 ;
      RECT  15660.0 91197.5 106080.0 91262.5 ;
      RECT  15660.0 93887.5 106080.0 93952.5 ;
      RECT  15660.0 96577.5 106080.0 96642.5 ;
      RECT  15660.0 99267.5 106080.0 99332.5 ;
      RECT  15660.0 101957.5 106080.0 102022.5 ;
      RECT  15660.0 104647.5 106080.0 104712.5 ;
      RECT  15660.0 107337.5 106080.0 107402.5 ;
      RECT  15660.0 110027.5 106080.0 110092.5 ;
      RECT  15660.0 112717.5 106080.0 112782.5 ;
      RECT  15660.0 27982.5 106080.0 28047.5 ;
      RECT  15660.0 30672.5 106080.0 30737.5 ;
      RECT  15660.0 33362.5 106080.0 33427.5 ;
      RECT  15660.0 36052.5 106080.0 36117.5 ;
      RECT  15660.0 38742.5 106080.0 38807.5 ;
      RECT  15660.0 41432.5 106080.0 41497.5 ;
      RECT  15660.0 44122.5 106080.0 44187.5 ;
      RECT  15660.0 46812.5 106080.0 46877.5 ;
      RECT  15660.0 49502.5 106080.0 49567.5 ;
      RECT  15660.0 52192.5 106080.0 52257.5 ;
      RECT  15660.0 54882.5 106080.0 54947.5 ;
      RECT  15660.0 57572.5 106080.0 57637.5 ;
      RECT  15660.0 60262.5 106080.0 60327.5 ;
      RECT  15660.0 62952.5 106080.0 63017.5 ;
      RECT  15660.0 65642.5 106080.0 65707.5 ;
      RECT  15660.0 68332.5 106080.0 68397.5 ;
      RECT  15660.0 71022.5 106080.0 71087.5 ;
      RECT  15660.0 73712.5 106080.0 73777.5 ;
      RECT  15660.0 76402.5 106080.0 76467.5 ;
      RECT  15660.0 79092.5 106080.0 79157.5 ;
      RECT  15660.0 81782.5 106080.0 81847.5 ;
      RECT  15660.0 84472.5 106080.0 84537.5 ;
      RECT  15660.0 87162.5 106080.0 87227.5 ;
      RECT  15660.0 89852.5 106080.0 89917.5 ;
      RECT  15660.0 92542.5 106080.0 92607.5 ;
      RECT  15660.0 95232.5 106080.0 95297.5 ;
      RECT  15660.0 97922.5 106080.0 97987.5 ;
      RECT  15660.0 100612.5 106080.0 100677.5 ;
      RECT  15660.0 103302.5 106080.0 103367.5 ;
      RECT  15660.0 105992.5 106080.0 106057.5 ;
      RECT  15660.0 108682.5 106080.0 108747.5 ;
      RECT  15660.0 111372.5 106080.0 111437.5 ;
      RECT  15660.0 114062.5 106080.0 114127.5 ;
      RECT  16102.5 115307.5 16167.5 115822.5 ;
      RECT  15912.5 114777.5 15977.5 114912.5 ;
      RECT  16102.5 114777.5 16167.5 114912.5 ;
      RECT  16102.5 114777.5 16167.5 114912.5 ;
      RECT  15912.5 114777.5 15977.5 114912.5 ;
      RECT  15912.5 115307.5 15977.5 115442.5 ;
      RECT  16102.5 115307.5 16167.5 115442.5 ;
      RECT  16102.5 115307.5 16167.5 115442.5 ;
      RECT  15912.5 115307.5 15977.5 115442.5 ;
      RECT  16102.5 115307.5 16167.5 115442.5 ;
      RECT  16292.5 115307.5 16357.5 115442.5 ;
      RECT  16292.5 115307.5 16357.5 115442.5 ;
      RECT  16102.5 115307.5 16167.5 115442.5 ;
      RECT  16082.5 115072.5 15947.5 115137.5 ;
      RECT  16102.5 115620.0 16167.5 115755.0 ;
      RECT  15912.5 114777.5 15977.5 114912.5 ;
      RECT  16102.5 114777.5 16167.5 114912.5 ;
      RECT  15912.5 115307.5 15977.5 115442.5 ;
      RECT  16292.5 115307.5 16357.5 115442.5 ;
      RECT  15750.0 115072.5 16455.0 115137.5 ;
      RECT  15750.0 115757.5 16455.0 115822.5 ;
      RECT  16807.5 115307.5 16872.5 115822.5 ;
      RECT  16617.5 114777.5 16682.5 114912.5 ;
      RECT  16807.5 114777.5 16872.5 114912.5 ;
      RECT  16807.5 114777.5 16872.5 114912.5 ;
      RECT  16617.5 114777.5 16682.5 114912.5 ;
      RECT  16617.5 115307.5 16682.5 115442.5 ;
      RECT  16807.5 115307.5 16872.5 115442.5 ;
      RECT  16807.5 115307.5 16872.5 115442.5 ;
      RECT  16617.5 115307.5 16682.5 115442.5 ;
      RECT  16807.5 115307.5 16872.5 115442.5 ;
      RECT  16997.5 115307.5 17062.5 115442.5 ;
      RECT  16997.5 115307.5 17062.5 115442.5 ;
      RECT  16807.5 115307.5 16872.5 115442.5 ;
      RECT  16787.5 115072.5 16652.5 115137.5 ;
      RECT  16807.5 115620.0 16872.5 115755.0 ;
      RECT  16617.5 114777.5 16682.5 114912.5 ;
      RECT  16807.5 114777.5 16872.5 114912.5 ;
      RECT  16617.5 115307.5 16682.5 115442.5 ;
      RECT  16997.5 115307.5 17062.5 115442.5 ;
      RECT  16455.0 115072.5 17160.0 115137.5 ;
      RECT  16455.0 115757.5 17160.0 115822.5 ;
      RECT  17512.5 115307.5 17577.5 115822.5 ;
      RECT  17322.5 114777.5 17387.5 114912.5 ;
      RECT  17512.5 114777.5 17577.5 114912.5 ;
      RECT  17512.5 114777.5 17577.5 114912.5 ;
      RECT  17322.5 114777.5 17387.5 114912.5 ;
      RECT  17322.5 115307.5 17387.5 115442.5 ;
      RECT  17512.5 115307.5 17577.5 115442.5 ;
      RECT  17512.5 115307.5 17577.5 115442.5 ;
      RECT  17322.5 115307.5 17387.5 115442.5 ;
      RECT  17512.5 115307.5 17577.5 115442.5 ;
      RECT  17702.5 115307.5 17767.5 115442.5 ;
      RECT  17702.5 115307.5 17767.5 115442.5 ;
      RECT  17512.5 115307.5 17577.5 115442.5 ;
      RECT  17492.5 115072.5 17357.5 115137.5 ;
      RECT  17512.5 115620.0 17577.5 115755.0 ;
      RECT  17322.5 114777.5 17387.5 114912.5 ;
      RECT  17512.5 114777.5 17577.5 114912.5 ;
      RECT  17322.5 115307.5 17387.5 115442.5 ;
      RECT  17702.5 115307.5 17767.5 115442.5 ;
      RECT  17160.0 115072.5 17865.0 115137.5 ;
      RECT  17160.0 115757.5 17865.0 115822.5 ;
      RECT  18217.5 115307.5 18282.5 115822.5 ;
      RECT  18027.5 114777.5 18092.5 114912.5 ;
      RECT  18217.5 114777.5 18282.5 114912.5 ;
      RECT  18217.5 114777.5 18282.5 114912.5 ;
      RECT  18027.5 114777.5 18092.5 114912.5 ;
      RECT  18027.5 115307.5 18092.5 115442.5 ;
      RECT  18217.5 115307.5 18282.5 115442.5 ;
      RECT  18217.5 115307.5 18282.5 115442.5 ;
      RECT  18027.5 115307.5 18092.5 115442.5 ;
      RECT  18217.5 115307.5 18282.5 115442.5 ;
      RECT  18407.5 115307.5 18472.5 115442.5 ;
      RECT  18407.5 115307.5 18472.5 115442.5 ;
      RECT  18217.5 115307.5 18282.5 115442.5 ;
      RECT  18197.5 115072.5 18062.5 115137.5 ;
      RECT  18217.5 115620.0 18282.5 115755.0 ;
      RECT  18027.5 114777.5 18092.5 114912.5 ;
      RECT  18217.5 114777.5 18282.5 114912.5 ;
      RECT  18027.5 115307.5 18092.5 115442.5 ;
      RECT  18407.5 115307.5 18472.5 115442.5 ;
      RECT  17865.0 115072.5 18570.0 115137.5 ;
      RECT  17865.0 115757.5 18570.0 115822.5 ;
      RECT  18922.5 115307.5 18987.5 115822.5 ;
      RECT  18732.5 114777.5 18797.5 114912.5 ;
      RECT  18922.5 114777.5 18987.5 114912.5 ;
      RECT  18922.5 114777.5 18987.5 114912.5 ;
      RECT  18732.5 114777.5 18797.5 114912.5 ;
      RECT  18732.5 115307.5 18797.5 115442.5 ;
      RECT  18922.5 115307.5 18987.5 115442.5 ;
      RECT  18922.5 115307.5 18987.5 115442.5 ;
      RECT  18732.5 115307.5 18797.5 115442.5 ;
      RECT  18922.5 115307.5 18987.5 115442.5 ;
      RECT  19112.5 115307.5 19177.5 115442.5 ;
      RECT  19112.5 115307.5 19177.5 115442.5 ;
      RECT  18922.5 115307.5 18987.5 115442.5 ;
      RECT  18902.5 115072.5 18767.5 115137.5 ;
      RECT  18922.5 115620.0 18987.5 115755.0 ;
      RECT  18732.5 114777.5 18797.5 114912.5 ;
      RECT  18922.5 114777.5 18987.5 114912.5 ;
      RECT  18732.5 115307.5 18797.5 115442.5 ;
      RECT  19112.5 115307.5 19177.5 115442.5 ;
      RECT  18570.0 115072.5 19275.0 115137.5 ;
      RECT  18570.0 115757.5 19275.0 115822.5 ;
      RECT  19627.5 115307.5 19692.5 115822.5 ;
      RECT  19437.5 114777.5 19502.5 114912.5 ;
      RECT  19627.5 114777.5 19692.5 114912.5 ;
      RECT  19627.5 114777.5 19692.5 114912.5 ;
      RECT  19437.5 114777.5 19502.5 114912.5 ;
      RECT  19437.5 115307.5 19502.5 115442.5 ;
      RECT  19627.5 115307.5 19692.5 115442.5 ;
      RECT  19627.5 115307.5 19692.5 115442.5 ;
      RECT  19437.5 115307.5 19502.5 115442.5 ;
      RECT  19627.5 115307.5 19692.5 115442.5 ;
      RECT  19817.5 115307.5 19882.5 115442.5 ;
      RECT  19817.5 115307.5 19882.5 115442.5 ;
      RECT  19627.5 115307.5 19692.5 115442.5 ;
      RECT  19607.5 115072.5 19472.5 115137.5 ;
      RECT  19627.5 115620.0 19692.5 115755.0 ;
      RECT  19437.5 114777.5 19502.5 114912.5 ;
      RECT  19627.5 114777.5 19692.5 114912.5 ;
      RECT  19437.5 115307.5 19502.5 115442.5 ;
      RECT  19817.5 115307.5 19882.5 115442.5 ;
      RECT  19275.0 115072.5 19980.0 115137.5 ;
      RECT  19275.0 115757.5 19980.0 115822.5 ;
      RECT  20332.5 115307.5 20397.5 115822.5 ;
      RECT  20142.5 114777.5 20207.5 114912.5 ;
      RECT  20332.5 114777.5 20397.5 114912.5 ;
      RECT  20332.5 114777.5 20397.5 114912.5 ;
      RECT  20142.5 114777.5 20207.5 114912.5 ;
      RECT  20142.5 115307.5 20207.5 115442.5 ;
      RECT  20332.5 115307.5 20397.5 115442.5 ;
      RECT  20332.5 115307.5 20397.5 115442.5 ;
      RECT  20142.5 115307.5 20207.5 115442.5 ;
      RECT  20332.5 115307.5 20397.5 115442.5 ;
      RECT  20522.5 115307.5 20587.5 115442.5 ;
      RECT  20522.5 115307.5 20587.5 115442.5 ;
      RECT  20332.5 115307.5 20397.5 115442.5 ;
      RECT  20312.5 115072.5 20177.5 115137.5 ;
      RECT  20332.5 115620.0 20397.5 115755.0 ;
      RECT  20142.5 114777.5 20207.5 114912.5 ;
      RECT  20332.5 114777.5 20397.5 114912.5 ;
      RECT  20142.5 115307.5 20207.5 115442.5 ;
      RECT  20522.5 115307.5 20587.5 115442.5 ;
      RECT  19980.0 115072.5 20685.0 115137.5 ;
      RECT  19980.0 115757.5 20685.0 115822.5 ;
      RECT  21037.5 115307.5 21102.5 115822.5 ;
      RECT  20847.5 114777.5 20912.5 114912.5 ;
      RECT  21037.5 114777.5 21102.5 114912.5 ;
      RECT  21037.5 114777.5 21102.5 114912.5 ;
      RECT  20847.5 114777.5 20912.5 114912.5 ;
      RECT  20847.5 115307.5 20912.5 115442.5 ;
      RECT  21037.5 115307.5 21102.5 115442.5 ;
      RECT  21037.5 115307.5 21102.5 115442.5 ;
      RECT  20847.5 115307.5 20912.5 115442.5 ;
      RECT  21037.5 115307.5 21102.5 115442.5 ;
      RECT  21227.5 115307.5 21292.5 115442.5 ;
      RECT  21227.5 115307.5 21292.5 115442.5 ;
      RECT  21037.5 115307.5 21102.5 115442.5 ;
      RECT  21017.5 115072.5 20882.5 115137.5 ;
      RECT  21037.5 115620.0 21102.5 115755.0 ;
      RECT  20847.5 114777.5 20912.5 114912.5 ;
      RECT  21037.5 114777.5 21102.5 114912.5 ;
      RECT  20847.5 115307.5 20912.5 115442.5 ;
      RECT  21227.5 115307.5 21292.5 115442.5 ;
      RECT  20685.0 115072.5 21390.0 115137.5 ;
      RECT  20685.0 115757.5 21390.0 115822.5 ;
      RECT  21742.5 115307.5 21807.5 115822.5 ;
      RECT  21552.5 114777.5 21617.5 114912.5 ;
      RECT  21742.5 114777.5 21807.5 114912.5 ;
      RECT  21742.5 114777.5 21807.5 114912.5 ;
      RECT  21552.5 114777.5 21617.5 114912.5 ;
      RECT  21552.5 115307.5 21617.5 115442.5 ;
      RECT  21742.5 115307.5 21807.5 115442.5 ;
      RECT  21742.5 115307.5 21807.5 115442.5 ;
      RECT  21552.5 115307.5 21617.5 115442.5 ;
      RECT  21742.5 115307.5 21807.5 115442.5 ;
      RECT  21932.5 115307.5 21997.5 115442.5 ;
      RECT  21932.5 115307.5 21997.5 115442.5 ;
      RECT  21742.5 115307.5 21807.5 115442.5 ;
      RECT  21722.5 115072.5 21587.5 115137.5 ;
      RECT  21742.5 115620.0 21807.5 115755.0 ;
      RECT  21552.5 114777.5 21617.5 114912.5 ;
      RECT  21742.5 114777.5 21807.5 114912.5 ;
      RECT  21552.5 115307.5 21617.5 115442.5 ;
      RECT  21932.5 115307.5 21997.5 115442.5 ;
      RECT  21390.0 115072.5 22095.0 115137.5 ;
      RECT  21390.0 115757.5 22095.0 115822.5 ;
      RECT  22447.5 115307.5 22512.5 115822.5 ;
      RECT  22257.5 114777.5 22322.5 114912.5 ;
      RECT  22447.5 114777.5 22512.5 114912.5 ;
      RECT  22447.5 114777.5 22512.5 114912.5 ;
      RECT  22257.5 114777.5 22322.5 114912.5 ;
      RECT  22257.5 115307.5 22322.5 115442.5 ;
      RECT  22447.5 115307.5 22512.5 115442.5 ;
      RECT  22447.5 115307.5 22512.5 115442.5 ;
      RECT  22257.5 115307.5 22322.5 115442.5 ;
      RECT  22447.5 115307.5 22512.5 115442.5 ;
      RECT  22637.5 115307.5 22702.5 115442.5 ;
      RECT  22637.5 115307.5 22702.5 115442.5 ;
      RECT  22447.5 115307.5 22512.5 115442.5 ;
      RECT  22427.5 115072.5 22292.5 115137.5 ;
      RECT  22447.5 115620.0 22512.5 115755.0 ;
      RECT  22257.5 114777.5 22322.5 114912.5 ;
      RECT  22447.5 114777.5 22512.5 114912.5 ;
      RECT  22257.5 115307.5 22322.5 115442.5 ;
      RECT  22637.5 115307.5 22702.5 115442.5 ;
      RECT  22095.0 115072.5 22800.0 115137.5 ;
      RECT  22095.0 115757.5 22800.0 115822.5 ;
      RECT  23152.5 115307.5 23217.5 115822.5 ;
      RECT  22962.5 114777.5 23027.5 114912.5 ;
      RECT  23152.5 114777.5 23217.5 114912.5 ;
      RECT  23152.5 114777.5 23217.5 114912.5 ;
      RECT  22962.5 114777.5 23027.5 114912.5 ;
      RECT  22962.5 115307.5 23027.5 115442.5 ;
      RECT  23152.5 115307.5 23217.5 115442.5 ;
      RECT  23152.5 115307.5 23217.5 115442.5 ;
      RECT  22962.5 115307.5 23027.5 115442.5 ;
      RECT  23152.5 115307.5 23217.5 115442.5 ;
      RECT  23342.5 115307.5 23407.5 115442.5 ;
      RECT  23342.5 115307.5 23407.5 115442.5 ;
      RECT  23152.5 115307.5 23217.5 115442.5 ;
      RECT  23132.5 115072.5 22997.5 115137.5 ;
      RECT  23152.5 115620.0 23217.5 115755.0 ;
      RECT  22962.5 114777.5 23027.5 114912.5 ;
      RECT  23152.5 114777.5 23217.5 114912.5 ;
      RECT  22962.5 115307.5 23027.5 115442.5 ;
      RECT  23342.5 115307.5 23407.5 115442.5 ;
      RECT  22800.0 115072.5 23505.0 115137.5 ;
      RECT  22800.0 115757.5 23505.0 115822.5 ;
      RECT  23857.5 115307.5 23922.5 115822.5 ;
      RECT  23667.5 114777.5 23732.5 114912.5 ;
      RECT  23857.5 114777.5 23922.5 114912.5 ;
      RECT  23857.5 114777.5 23922.5 114912.5 ;
      RECT  23667.5 114777.5 23732.5 114912.5 ;
      RECT  23667.5 115307.5 23732.5 115442.5 ;
      RECT  23857.5 115307.5 23922.5 115442.5 ;
      RECT  23857.5 115307.5 23922.5 115442.5 ;
      RECT  23667.5 115307.5 23732.5 115442.5 ;
      RECT  23857.5 115307.5 23922.5 115442.5 ;
      RECT  24047.5 115307.5 24112.5 115442.5 ;
      RECT  24047.5 115307.5 24112.5 115442.5 ;
      RECT  23857.5 115307.5 23922.5 115442.5 ;
      RECT  23837.5 115072.5 23702.5 115137.5 ;
      RECT  23857.5 115620.0 23922.5 115755.0 ;
      RECT  23667.5 114777.5 23732.5 114912.5 ;
      RECT  23857.5 114777.5 23922.5 114912.5 ;
      RECT  23667.5 115307.5 23732.5 115442.5 ;
      RECT  24047.5 115307.5 24112.5 115442.5 ;
      RECT  23505.0 115072.5 24210.0 115137.5 ;
      RECT  23505.0 115757.5 24210.0 115822.5 ;
      RECT  24562.5 115307.5 24627.5 115822.5 ;
      RECT  24372.5 114777.5 24437.5 114912.5 ;
      RECT  24562.5 114777.5 24627.5 114912.5 ;
      RECT  24562.5 114777.5 24627.5 114912.5 ;
      RECT  24372.5 114777.5 24437.5 114912.5 ;
      RECT  24372.5 115307.5 24437.5 115442.5 ;
      RECT  24562.5 115307.5 24627.5 115442.5 ;
      RECT  24562.5 115307.5 24627.5 115442.5 ;
      RECT  24372.5 115307.5 24437.5 115442.5 ;
      RECT  24562.5 115307.5 24627.5 115442.5 ;
      RECT  24752.5 115307.5 24817.5 115442.5 ;
      RECT  24752.5 115307.5 24817.5 115442.5 ;
      RECT  24562.5 115307.5 24627.5 115442.5 ;
      RECT  24542.5 115072.5 24407.5 115137.5 ;
      RECT  24562.5 115620.0 24627.5 115755.0 ;
      RECT  24372.5 114777.5 24437.5 114912.5 ;
      RECT  24562.5 114777.5 24627.5 114912.5 ;
      RECT  24372.5 115307.5 24437.5 115442.5 ;
      RECT  24752.5 115307.5 24817.5 115442.5 ;
      RECT  24210.0 115072.5 24915.0 115137.5 ;
      RECT  24210.0 115757.5 24915.0 115822.5 ;
      RECT  25267.5 115307.5 25332.5 115822.5 ;
      RECT  25077.5 114777.5 25142.5 114912.5 ;
      RECT  25267.5 114777.5 25332.5 114912.5 ;
      RECT  25267.5 114777.5 25332.5 114912.5 ;
      RECT  25077.5 114777.5 25142.5 114912.5 ;
      RECT  25077.5 115307.5 25142.5 115442.5 ;
      RECT  25267.5 115307.5 25332.5 115442.5 ;
      RECT  25267.5 115307.5 25332.5 115442.5 ;
      RECT  25077.5 115307.5 25142.5 115442.5 ;
      RECT  25267.5 115307.5 25332.5 115442.5 ;
      RECT  25457.5 115307.5 25522.5 115442.5 ;
      RECT  25457.5 115307.5 25522.5 115442.5 ;
      RECT  25267.5 115307.5 25332.5 115442.5 ;
      RECT  25247.5 115072.5 25112.5 115137.5 ;
      RECT  25267.5 115620.0 25332.5 115755.0 ;
      RECT  25077.5 114777.5 25142.5 114912.5 ;
      RECT  25267.5 114777.5 25332.5 114912.5 ;
      RECT  25077.5 115307.5 25142.5 115442.5 ;
      RECT  25457.5 115307.5 25522.5 115442.5 ;
      RECT  24915.0 115072.5 25620.0 115137.5 ;
      RECT  24915.0 115757.5 25620.0 115822.5 ;
      RECT  25972.5 115307.5 26037.5 115822.5 ;
      RECT  25782.5 114777.5 25847.5 114912.5 ;
      RECT  25972.5 114777.5 26037.5 114912.5 ;
      RECT  25972.5 114777.5 26037.5 114912.5 ;
      RECT  25782.5 114777.5 25847.5 114912.5 ;
      RECT  25782.5 115307.5 25847.5 115442.5 ;
      RECT  25972.5 115307.5 26037.5 115442.5 ;
      RECT  25972.5 115307.5 26037.5 115442.5 ;
      RECT  25782.5 115307.5 25847.5 115442.5 ;
      RECT  25972.5 115307.5 26037.5 115442.5 ;
      RECT  26162.5 115307.5 26227.5 115442.5 ;
      RECT  26162.5 115307.5 26227.5 115442.5 ;
      RECT  25972.5 115307.5 26037.5 115442.5 ;
      RECT  25952.5 115072.5 25817.5 115137.5 ;
      RECT  25972.5 115620.0 26037.5 115755.0 ;
      RECT  25782.5 114777.5 25847.5 114912.5 ;
      RECT  25972.5 114777.5 26037.5 114912.5 ;
      RECT  25782.5 115307.5 25847.5 115442.5 ;
      RECT  26162.5 115307.5 26227.5 115442.5 ;
      RECT  25620.0 115072.5 26325.0 115137.5 ;
      RECT  25620.0 115757.5 26325.0 115822.5 ;
      RECT  26677.5 115307.5 26742.5 115822.5 ;
      RECT  26487.5 114777.5 26552.5 114912.5 ;
      RECT  26677.5 114777.5 26742.5 114912.5 ;
      RECT  26677.5 114777.5 26742.5 114912.5 ;
      RECT  26487.5 114777.5 26552.5 114912.5 ;
      RECT  26487.5 115307.5 26552.5 115442.5 ;
      RECT  26677.5 115307.5 26742.5 115442.5 ;
      RECT  26677.5 115307.5 26742.5 115442.5 ;
      RECT  26487.5 115307.5 26552.5 115442.5 ;
      RECT  26677.5 115307.5 26742.5 115442.5 ;
      RECT  26867.5 115307.5 26932.5 115442.5 ;
      RECT  26867.5 115307.5 26932.5 115442.5 ;
      RECT  26677.5 115307.5 26742.5 115442.5 ;
      RECT  26657.5 115072.5 26522.5 115137.5 ;
      RECT  26677.5 115620.0 26742.5 115755.0 ;
      RECT  26487.5 114777.5 26552.5 114912.5 ;
      RECT  26677.5 114777.5 26742.5 114912.5 ;
      RECT  26487.5 115307.5 26552.5 115442.5 ;
      RECT  26867.5 115307.5 26932.5 115442.5 ;
      RECT  26325.0 115072.5 27030.0 115137.5 ;
      RECT  26325.0 115757.5 27030.0 115822.5 ;
      RECT  27382.5 115307.5 27447.5 115822.5 ;
      RECT  27192.5 114777.5 27257.5 114912.5 ;
      RECT  27382.5 114777.5 27447.5 114912.5 ;
      RECT  27382.5 114777.5 27447.5 114912.5 ;
      RECT  27192.5 114777.5 27257.5 114912.5 ;
      RECT  27192.5 115307.5 27257.5 115442.5 ;
      RECT  27382.5 115307.5 27447.5 115442.5 ;
      RECT  27382.5 115307.5 27447.5 115442.5 ;
      RECT  27192.5 115307.5 27257.5 115442.5 ;
      RECT  27382.5 115307.5 27447.5 115442.5 ;
      RECT  27572.5 115307.5 27637.5 115442.5 ;
      RECT  27572.5 115307.5 27637.5 115442.5 ;
      RECT  27382.5 115307.5 27447.5 115442.5 ;
      RECT  27362.5 115072.5 27227.5 115137.5 ;
      RECT  27382.5 115620.0 27447.5 115755.0 ;
      RECT  27192.5 114777.5 27257.5 114912.5 ;
      RECT  27382.5 114777.5 27447.5 114912.5 ;
      RECT  27192.5 115307.5 27257.5 115442.5 ;
      RECT  27572.5 115307.5 27637.5 115442.5 ;
      RECT  27030.0 115072.5 27735.0 115137.5 ;
      RECT  27030.0 115757.5 27735.0 115822.5 ;
      RECT  28087.5 115307.5 28152.5 115822.5 ;
      RECT  27897.5 114777.5 27962.5 114912.5 ;
      RECT  28087.5 114777.5 28152.5 114912.5 ;
      RECT  28087.5 114777.5 28152.5 114912.5 ;
      RECT  27897.5 114777.5 27962.5 114912.5 ;
      RECT  27897.5 115307.5 27962.5 115442.5 ;
      RECT  28087.5 115307.5 28152.5 115442.5 ;
      RECT  28087.5 115307.5 28152.5 115442.5 ;
      RECT  27897.5 115307.5 27962.5 115442.5 ;
      RECT  28087.5 115307.5 28152.5 115442.5 ;
      RECT  28277.5 115307.5 28342.5 115442.5 ;
      RECT  28277.5 115307.5 28342.5 115442.5 ;
      RECT  28087.5 115307.5 28152.5 115442.5 ;
      RECT  28067.5 115072.5 27932.5 115137.5 ;
      RECT  28087.5 115620.0 28152.5 115755.0 ;
      RECT  27897.5 114777.5 27962.5 114912.5 ;
      RECT  28087.5 114777.5 28152.5 114912.5 ;
      RECT  27897.5 115307.5 27962.5 115442.5 ;
      RECT  28277.5 115307.5 28342.5 115442.5 ;
      RECT  27735.0 115072.5 28440.0 115137.5 ;
      RECT  27735.0 115757.5 28440.0 115822.5 ;
      RECT  28792.5 115307.5 28857.5 115822.5 ;
      RECT  28602.5 114777.5 28667.5 114912.5 ;
      RECT  28792.5 114777.5 28857.5 114912.5 ;
      RECT  28792.5 114777.5 28857.5 114912.5 ;
      RECT  28602.5 114777.5 28667.5 114912.5 ;
      RECT  28602.5 115307.5 28667.5 115442.5 ;
      RECT  28792.5 115307.5 28857.5 115442.5 ;
      RECT  28792.5 115307.5 28857.5 115442.5 ;
      RECT  28602.5 115307.5 28667.5 115442.5 ;
      RECT  28792.5 115307.5 28857.5 115442.5 ;
      RECT  28982.5 115307.5 29047.5 115442.5 ;
      RECT  28982.5 115307.5 29047.5 115442.5 ;
      RECT  28792.5 115307.5 28857.5 115442.5 ;
      RECT  28772.5 115072.5 28637.5 115137.5 ;
      RECT  28792.5 115620.0 28857.5 115755.0 ;
      RECT  28602.5 114777.5 28667.5 114912.5 ;
      RECT  28792.5 114777.5 28857.5 114912.5 ;
      RECT  28602.5 115307.5 28667.5 115442.5 ;
      RECT  28982.5 115307.5 29047.5 115442.5 ;
      RECT  28440.0 115072.5 29145.0 115137.5 ;
      RECT  28440.0 115757.5 29145.0 115822.5 ;
      RECT  29497.5 115307.5 29562.5 115822.5 ;
      RECT  29307.5 114777.5 29372.5 114912.5 ;
      RECT  29497.5 114777.5 29562.5 114912.5 ;
      RECT  29497.5 114777.5 29562.5 114912.5 ;
      RECT  29307.5 114777.5 29372.5 114912.5 ;
      RECT  29307.5 115307.5 29372.5 115442.5 ;
      RECT  29497.5 115307.5 29562.5 115442.5 ;
      RECT  29497.5 115307.5 29562.5 115442.5 ;
      RECT  29307.5 115307.5 29372.5 115442.5 ;
      RECT  29497.5 115307.5 29562.5 115442.5 ;
      RECT  29687.5 115307.5 29752.5 115442.5 ;
      RECT  29687.5 115307.5 29752.5 115442.5 ;
      RECT  29497.5 115307.5 29562.5 115442.5 ;
      RECT  29477.5 115072.5 29342.5 115137.5 ;
      RECT  29497.5 115620.0 29562.5 115755.0 ;
      RECT  29307.5 114777.5 29372.5 114912.5 ;
      RECT  29497.5 114777.5 29562.5 114912.5 ;
      RECT  29307.5 115307.5 29372.5 115442.5 ;
      RECT  29687.5 115307.5 29752.5 115442.5 ;
      RECT  29145.0 115072.5 29850.0 115137.5 ;
      RECT  29145.0 115757.5 29850.0 115822.5 ;
      RECT  30202.5 115307.5 30267.5 115822.5 ;
      RECT  30012.5 114777.5 30077.5 114912.5 ;
      RECT  30202.5 114777.5 30267.5 114912.5 ;
      RECT  30202.5 114777.5 30267.5 114912.5 ;
      RECT  30012.5 114777.5 30077.5 114912.5 ;
      RECT  30012.5 115307.5 30077.5 115442.5 ;
      RECT  30202.5 115307.5 30267.5 115442.5 ;
      RECT  30202.5 115307.5 30267.5 115442.5 ;
      RECT  30012.5 115307.5 30077.5 115442.5 ;
      RECT  30202.5 115307.5 30267.5 115442.5 ;
      RECT  30392.5 115307.5 30457.5 115442.5 ;
      RECT  30392.5 115307.5 30457.5 115442.5 ;
      RECT  30202.5 115307.5 30267.5 115442.5 ;
      RECT  30182.5 115072.5 30047.5 115137.5 ;
      RECT  30202.5 115620.0 30267.5 115755.0 ;
      RECT  30012.5 114777.5 30077.5 114912.5 ;
      RECT  30202.5 114777.5 30267.5 114912.5 ;
      RECT  30012.5 115307.5 30077.5 115442.5 ;
      RECT  30392.5 115307.5 30457.5 115442.5 ;
      RECT  29850.0 115072.5 30555.0 115137.5 ;
      RECT  29850.0 115757.5 30555.0 115822.5 ;
      RECT  30907.5 115307.5 30972.5 115822.5 ;
      RECT  30717.5 114777.5 30782.5 114912.5 ;
      RECT  30907.5 114777.5 30972.5 114912.5 ;
      RECT  30907.5 114777.5 30972.5 114912.5 ;
      RECT  30717.5 114777.5 30782.5 114912.5 ;
      RECT  30717.5 115307.5 30782.5 115442.5 ;
      RECT  30907.5 115307.5 30972.5 115442.5 ;
      RECT  30907.5 115307.5 30972.5 115442.5 ;
      RECT  30717.5 115307.5 30782.5 115442.5 ;
      RECT  30907.5 115307.5 30972.5 115442.5 ;
      RECT  31097.5 115307.5 31162.5 115442.5 ;
      RECT  31097.5 115307.5 31162.5 115442.5 ;
      RECT  30907.5 115307.5 30972.5 115442.5 ;
      RECT  30887.5 115072.5 30752.5 115137.5 ;
      RECT  30907.5 115620.0 30972.5 115755.0 ;
      RECT  30717.5 114777.5 30782.5 114912.5 ;
      RECT  30907.5 114777.5 30972.5 114912.5 ;
      RECT  30717.5 115307.5 30782.5 115442.5 ;
      RECT  31097.5 115307.5 31162.5 115442.5 ;
      RECT  30555.0 115072.5 31260.0 115137.5 ;
      RECT  30555.0 115757.5 31260.0 115822.5 ;
      RECT  31612.5 115307.5 31677.5 115822.5 ;
      RECT  31422.5 114777.5 31487.5 114912.5 ;
      RECT  31612.5 114777.5 31677.5 114912.5 ;
      RECT  31612.5 114777.5 31677.5 114912.5 ;
      RECT  31422.5 114777.5 31487.5 114912.5 ;
      RECT  31422.5 115307.5 31487.5 115442.5 ;
      RECT  31612.5 115307.5 31677.5 115442.5 ;
      RECT  31612.5 115307.5 31677.5 115442.5 ;
      RECT  31422.5 115307.5 31487.5 115442.5 ;
      RECT  31612.5 115307.5 31677.5 115442.5 ;
      RECT  31802.5 115307.5 31867.5 115442.5 ;
      RECT  31802.5 115307.5 31867.5 115442.5 ;
      RECT  31612.5 115307.5 31677.5 115442.5 ;
      RECT  31592.5 115072.5 31457.5 115137.5 ;
      RECT  31612.5 115620.0 31677.5 115755.0 ;
      RECT  31422.5 114777.5 31487.5 114912.5 ;
      RECT  31612.5 114777.5 31677.5 114912.5 ;
      RECT  31422.5 115307.5 31487.5 115442.5 ;
      RECT  31802.5 115307.5 31867.5 115442.5 ;
      RECT  31260.0 115072.5 31965.0 115137.5 ;
      RECT  31260.0 115757.5 31965.0 115822.5 ;
      RECT  32317.5 115307.5 32382.5 115822.5 ;
      RECT  32127.5 114777.5 32192.5 114912.5 ;
      RECT  32317.5 114777.5 32382.5 114912.5 ;
      RECT  32317.5 114777.5 32382.5 114912.5 ;
      RECT  32127.5 114777.5 32192.5 114912.5 ;
      RECT  32127.5 115307.5 32192.5 115442.5 ;
      RECT  32317.5 115307.5 32382.5 115442.5 ;
      RECT  32317.5 115307.5 32382.5 115442.5 ;
      RECT  32127.5 115307.5 32192.5 115442.5 ;
      RECT  32317.5 115307.5 32382.5 115442.5 ;
      RECT  32507.5 115307.5 32572.5 115442.5 ;
      RECT  32507.5 115307.5 32572.5 115442.5 ;
      RECT  32317.5 115307.5 32382.5 115442.5 ;
      RECT  32297.5 115072.5 32162.5 115137.5 ;
      RECT  32317.5 115620.0 32382.5 115755.0 ;
      RECT  32127.5 114777.5 32192.5 114912.5 ;
      RECT  32317.5 114777.5 32382.5 114912.5 ;
      RECT  32127.5 115307.5 32192.5 115442.5 ;
      RECT  32507.5 115307.5 32572.5 115442.5 ;
      RECT  31965.0 115072.5 32670.0 115137.5 ;
      RECT  31965.0 115757.5 32670.0 115822.5 ;
      RECT  33022.5 115307.5 33087.5 115822.5 ;
      RECT  32832.5 114777.5 32897.5 114912.5 ;
      RECT  33022.5 114777.5 33087.5 114912.5 ;
      RECT  33022.5 114777.5 33087.5 114912.5 ;
      RECT  32832.5 114777.5 32897.5 114912.5 ;
      RECT  32832.5 115307.5 32897.5 115442.5 ;
      RECT  33022.5 115307.5 33087.5 115442.5 ;
      RECT  33022.5 115307.5 33087.5 115442.5 ;
      RECT  32832.5 115307.5 32897.5 115442.5 ;
      RECT  33022.5 115307.5 33087.5 115442.5 ;
      RECT  33212.5 115307.5 33277.5 115442.5 ;
      RECT  33212.5 115307.5 33277.5 115442.5 ;
      RECT  33022.5 115307.5 33087.5 115442.5 ;
      RECT  33002.5 115072.5 32867.5 115137.5 ;
      RECT  33022.5 115620.0 33087.5 115755.0 ;
      RECT  32832.5 114777.5 32897.5 114912.5 ;
      RECT  33022.5 114777.5 33087.5 114912.5 ;
      RECT  32832.5 115307.5 32897.5 115442.5 ;
      RECT  33212.5 115307.5 33277.5 115442.5 ;
      RECT  32670.0 115072.5 33375.0 115137.5 ;
      RECT  32670.0 115757.5 33375.0 115822.5 ;
      RECT  33727.5 115307.5 33792.5 115822.5 ;
      RECT  33537.5 114777.5 33602.5 114912.5 ;
      RECT  33727.5 114777.5 33792.5 114912.5 ;
      RECT  33727.5 114777.5 33792.5 114912.5 ;
      RECT  33537.5 114777.5 33602.5 114912.5 ;
      RECT  33537.5 115307.5 33602.5 115442.5 ;
      RECT  33727.5 115307.5 33792.5 115442.5 ;
      RECT  33727.5 115307.5 33792.5 115442.5 ;
      RECT  33537.5 115307.5 33602.5 115442.5 ;
      RECT  33727.5 115307.5 33792.5 115442.5 ;
      RECT  33917.5 115307.5 33982.5 115442.5 ;
      RECT  33917.5 115307.5 33982.5 115442.5 ;
      RECT  33727.5 115307.5 33792.5 115442.5 ;
      RECT  33707.5 115072.5 33572.5 115137.5 ;
      RECT  33727.5 115620.0 33792.5 115755.0 ;
      RECT  33537.5 114777.5 33602.5 114912.5 ;
      RECT  33727.5 114777.5 33792.5 114912.5 ;
      RECT  33537.5 115307.5 33602.5 115442.5 ;
      RECT  33917.5 115307.5 33982.5 115442.5 ;
      RECT  33375.0 115072.5 34080.0 115137.5 ;
      RECT  33375.0 115757.5 34080.0 115822.5 ;
      RECT  34432.5 115307.5 34497.5 115822.5 ;
      RECT  34242.5 114777.5 34307.5 114912.5 ;
      RECT  34432.5 114777.5 34497.5 114912.5 ;
      RECT  34432.5 114777.5 34497.5 114912.5 ;
      RECT  34242.5 114777.5 34307.5 114912.5 ;
      RECT  34242.5 115307.5 34307.5 115442.5 ;
      RECT  34432.5 115307.5 34497.5 115442.5 ;
      RECT  34432.5 115307.5 34497.5 115442.5 ;
      RECT  34242.5 115307.5 34307.5 115442.5 ;
      RECT  34432.5 115307.5 34497.5 115442.5 ;
      RECT  34622.5 115307.5 34687.5 115442.5 ;
      RECT  34622.5 115307.5 34687.5 115442.5 ;
      RECT  34432.5 115307.5 34497.5 115442.5 ;
      RECT  34412.5 115072.5 34277.5 115137.5 ;
      RECT  34432.5 115620.0 34497.5 115755.0 ;
      RECT  34242.5 114777.5 34307.5 114912.5 ;
      RECT  34432.5 114777.5 34497.5 114912.5 ;
      RECT  34242.5 115307.5 34307.5 115442.5 ;
      RECT  34622.5 115307.5 34687.5 115442.5 ;
      RECT  34080.0 115072.5 34785.0 115137.5 ;
      RECT  34080.0 115757.5 34785.0 115822.5 ;
      RECT  35137.5 115307.5 35202.5 115822.5 ;
      RECT  34947.5 114777.5 35012.5 114912.5 ;
      RECT  35137.5 114777.5 35202.5 114912.5 ;
      RECT  35137.5 114777.5 35202.5 114912.5 ;
      RECT  34947.5 114777.5 35012.5 114912.5 ;
      RECT  34947.5 115307.5 35012.5 115442.5 ;
      RECT  35137.5 115307.5 35202.5 115442.5 ;
      RECT  35137.5 115307.5 35202.5 115442.5 ;
      RECT  34947.5 115307.5 35012.5 115442.5 ;
      RECT  35137.5 115307.5 35202.5 115442.5 ;
      RECT  35327.5 115307.5 35392.5 115442.5 ;
      RECT  35327.5 115307.5 35392.5 115442.5 ;
      RECT  35137.5 115307.5 35202.5 115442.5 ;
      RECT  35117.5 115072.5 34982.5 115137.5 ;
      RECT  35137.5 115620.0 35202.5 115755.0 ;
      RECT  34947.5 114777.5 35012.5 114912.5 ;
      RECT  35137.5 114777.5 35202.5 114912.5 ;
      RECT  34947.5 115307.5 35012.5 115442.5 ;
      RECT  35327.5 115307.5 35392.5 115442.5 ;
      RECT  34785.0 115072.5 35490.0 115137.5 ;
      RECT  34785.0 115757.5 35490.0 115822.5 ;
      RECT  35842.5 115307.5 35907.5 115822.5 ;
      RECT  35652.5 114777.5 35717.5 114912.5 ;
      RECT  35842.5 114777.5 35907.5 114912.5 ;
      RECT  35842.5 114777.5 35907.5 114912.5 ;
      RECT  35652.5 114777.5 35717.5 114912.5 ;
      RECT  35652.5 115307.5 35717.5 115442.5 ;
      RECT  35842.5 115307.5 35907.5 115442.5 ;
      RECT  35842.5 115307.5 35907.5 115442.5 ;
      RECT  35652.5 115307.5 35717.5 115442.5 ;
      RECT  35842.5 115307.5 35907.5 115442.5 ;
      RECT  36032.5 115307.5 36097.5 115442.5 ;
      RECT  36032.5 115307.5 36097.5 115442.5 ;
      RECT  35842.5 115307.5 35907.5 115442.5 ;
      RECT  35822.5 115072.5 35687.5 115137.5 ;
      RECT  35842.5 115620.0 35907.5 115755.0 ;
      RECT  35652.5 114777.5 35717.5 114912.5 ;
      RECT  35842.5 114777.5 35907.5 114912.5 ;
      RECT  35652.5 115307.5 35717.5 115442.5 ;
      RECT  36032.5 115307.5 36097.5 115442.5 ;
      RECT  35490.0 115072.5 36195.0 115137.5 ;
      RECT  35490.0 115757.5 36195.0 115822.5 ;
      RECT  36547.5 115307.5 36612.5 115822.5 ;
      RECT  36357.5 114777.5 36422.5 114912.5 ;
      RECT  36547.5 114777.5 36612.5 114912.5 ;
      RECT  36547.5 114777.5 36612.5 114912.5 ;
      RECT  36357.5 114777.5 36422.5 114912.5 ;
      RECT  36357.5 115307.5 36422.5 115442.5 ;
      RECT  36547.5 115307.5 36612.5 115442.5 ;
      RECT  36547.5 115307.5 36612.5 115442.5 ;
      RECT  36357.5 115307.5 36422.5 115442.5 ;
      RECT  36547.5 115307.5 36612.5 115442.5 ;
      RECT  36737.5 115307.5 36802.5 115442.5 ;
      RECT  36737.5 115307.5 36802.5 115442.5 ;
      RECT  36547.5 115307.5 36612.5 115442.5 ;
      RECT  36527.5 115072.5 36392.5 115137.5 ;
      RECT  36547.5 115620.0 36612.5 115755.0 ;
      RECT  36357.5 114777.5 36422.5 114912.5 ;
      RECT  36547.5 114777.5 36612.5 114912.5 ;
      RECT  36357.5 115307.5 36422.5 115442.5 ;
      RECT  36737.5 115307.5 36802.5 115442.5 ;
      RECT  36195.0 115072.5 36900.0 115137.5 ;
      RECT  36195.0 115757.5 36900.0 115822.5 ;
      RECT  37252.5 115307.5 37317.5 115822.5 ;
      RECT  37062.5 114777.5 37127.5 114912.5 ;
      RECT  37252.5 114777.5 37317.5 114912.5 ;
      RECT  37252.5 114777.5 37317.5 114912.5 ;
      RECT  37062.5 114777.5 37127.5 114912.5 ;
      RECT  37062.5 115307.5 37127.5 115442.5 ;
      RECT  37252.5 115307.5 37317.5 115442.5 ;
      RECT  37252.5 115307.5 37317.5 115442.5 ;
      RECT  37062.5 115307.5 37127.5 115442.5 ;
      RECT  37252.5 115307.5 37317.5 115442.5 ;
      RECT  37442.5 115307.5 37507.5 115442.5 ;
      RECT  37442.5 115307.5 37507.5 115442.5 ;
      RECT  37252.5 115307.5 37317.5 115442.5 ;
      RECT  37232.5 115072.5 37097.5 115137.5 ;
      RECT  37252.5 115620.0 37317.5 115755.0 ;
      RECT  37062.5 114777.5 37127.5 114912.5 ;
      RECT  37252.5 114777.5 37317.5 114912.5 ;
      RECT  37062.5 115307.5 37127.5 115442.5 ;
      RECT  37442.5 115307.5 37507.5 115442.5 ;
      RECT  36900.0 115072.5 37605.0 115137.5 ;
      RECT  36900.0 115757.5 37605.0 115822.5 ;
      RECT  37957.5 115307.5 38022.5 115822.5 ;
      RECT  37767.5 114777.5 37832.5 114912.5 ;
      RECT  37957.5 114777.5 38022.5 114912.5 ;
      RECT  37957.5 114777.5 38022.5 114912.5 ;
      RECT  37767.5 114777.5 37832.5 114912.5 ;
      RECT  37767.5 115307.5 37832.5 115442.5 ;
      RECT  37957.5 115307.5 38022.5 115442.5 ;
      RECT  37957.5 115307.5 38022.5 115442.5 ;
      RECT  37767.5 115307.5 37832.5 115442.5 ;
      RECT  37957.5 115307.5 38022.5 115442.5 ;
      RECT  38147.5 115307.5 38212.5 115442.5 ;
      RECT  38147.5 115307.5 38212.5 115442.5 ;
      RECT  37957.5 115307.5 38022.5 115442.5 ;
      RECT  37937.5 115072.5 37802.5 115137.5 ;
      RECT  37957.5 115620.0 38022.5 115755.0 ;
      RECT  37767.5 114777.5 37832.5 114912.5 ;
      RECT  37957.5 114777.5 38022.5 114912.5 ;
      RECT  37767.5 115307.5 37832.5 115442.5 ;
      RECT  38147.5 115307.5 38212.5 115442.5 ;
      RECT  37605.0 115072.5 38310.0 115137.5 ;
      RECT  37605.0 115757.5 38310.0 115822.5 ;
      RECT  38662.5 115307.5 38727.5 115822.5 ;
      RECT  38472.5 114777.5 38537.5 114912.5 ;
      RECT  38662.5 114777.5 38727.5 114912.5 ;
      RECT  38662.5 114777.5 38727.5 114912.5 ;
      RECT  38472.5 114777.5 38537.5 114912.5 ;
      RECT  38472.5 115307.5 38537.5 115442.5 ;
      RECT  38662.5 115307.5 38727.5 115442.5 ;
      RECT  38662.5 115307.5 38727.5 115442.5 ;
      RECT  38472.5 115307.5 38537.5 115442.5 ;
      RECT  38662.5 115307.5 38727.5 115442.5 ;
      RECT  38852.5 115307.5 38917.5 115442.5 ;
      RECT  38852.5 115307.5 38917.5 115442.5 ;
      RECT  38662.5 115307.5 38727.5 115442.5 ;
      RECT  38642.5 115072.5 38507.5 115137.5 ;
      RECT  38662.5 115620.0 38727.5 115755.0 ;
      RECT  38472.5 114777.5 38537.5 114912.5 ;
      RECT  38662.5 114777.5 38727.5 114912.5 ;
      RECT  38472.5 115307.5 38537.5 115442.5 ;
      RECT  38852.5 115307.5 38917.5 115442.5 ;
      RECT  38310.0 115072.5 39015.0 115137.5 ;
      RECT  38310.0 115757.5 39015.0 115822.5 ;
      RECT  39367.5 115307.5 39432.5 115822.5 ;
      RECT  39177.5 114777.5 39242.5 114912.5 ;
      RECT  39367.5 114777.5 39432.5 114912.5 ;
      RECT  39367.5 114777.5 39432.5 114912.5 ;
      RECT  39177.5 114777.5 39242.5 114912.5 ;
      RECT  39177.5 115307.5 39242.5 115442.5 ;
      RECT  39367.5 115307.5 39432.5 115442.5 ;
      RECT  39367.5 115307.5 39432.5 115442.5 ;
      RECT  39177.5 115307.5 39242.5 115442.5 ;
      RECT  39367.5 115307.5 39432.5 115442.5 ;
      RECT  39557.5 115307.5 39622.5 115442.5 ;
      RECT  39557.5 115307.5 39622.5 115442.5 ;
      RECT  39367.5 115307.5 39432.5 115442.5 ;
      RECT  39347.5 115072.5 39212.5 115137.5 ;
      RECT  39367.5 115620.0 39432.5 115755.0 ;
      RECT  39177.5 114777.5 39242.5 114912.5 ;
      RECT  39367.5 114777.5 39432.5 114912.5 ;
      RECT  39177.5 115307.5 39242.5 115442.5 ;
      RECT  39557.5 115307.5 39622.5 115442.5 ;
      RECT  39015.0 115072.5 39720.0 115137.5 ;
      RECT  39015.0 115757.5 39720.0 115822.5 ;
      RECT  40072.5 115307.5 40137.5 115822.5 ;
      RECT  39882.5 114777.5 39947.5 114912.5 ;
      RECT  40072.5 114777.5 40137.5 114912.5 ;
      RECT  40072.5 114777.5 40137.5 114912.5 ;
      RECT  39882.5 114777.5 39947.5 114912.5 ;
      RECT  39882.5 115307.5 39947.5 115442.5 ;
      RECT  40072.5 115307.5 40137.5 115442.5 ;
      RECT  40072.5 115307.5 40137.5 115442.5 ;
      RECT  39882.5 115307.5 39947.5 115442.5 ;
      RECT  40072.5 115307.5 40137.5 115442.5 ;
      RECT  40262.5 115307.5 40327.5 115442.5 ;
      RECT  40262.5 115307.5 40327.5 115442.5 ;
      RECT  40072.5 115307.5 40137.5 115442.5 ;
      RECT  40052.5 115072.5 39917.5 115137.5 ;
      RECT  40072.5 115620.0 40137.5 115755.0 ;
      RECT  39882.5 114777.5 39947.5 114912.5 ;
      RECT  40072.5 114777.5 40137.5 114912.5 ;
      RECT  39882.5 115307.5 39947.5 115442.5 ;
      RECT  40262.5 115307.5 40327.5 115442.5 ;
      RECT  39720.0 115072.5 40425.0 115137.5 ;
      RECT  39720.0 115757.5 40425.0 115822.5 ;
      RECT  40777.5 115307.5 40842.5 115822.5 ;
      RECT  40587.5 114777.5 40652.5 114912.5 ;
      RECT  40777.5 114777.5 40842.5 114912.5 ;
      RECT  40777.5 114777.5 40842.5 114912.5 ;
      RECT  40587.5 114777.5 40652.5 114912.5 ;
      RECT  40587.5 115307.5 40652.5 115442.5 ;
      RECT  40777.5 115307.5 40842.5 115442.5 ;
      RECT  40777.5 115307.5 40842.5 115442.5 ;
      RECT  40587.5 115307.5 40652.5 115442.5 ;
      RECT  40777.5 115307.5 40842.5 115442.5 ;
      RECT  40967.5 115307.5 41032.5 115442.5 ;
      RECT  40967.5 115307.5 41032.5 115442.5 ;
      RECT  40777.5 115307.5 40842.5 115442.5 ;
      RECT  40757.5 115072.5 40622.5 115137.5 ;
      RECT  40777.5 115620.0 40842.5 115755.0 ;
      RECT  40587.5 114777.5 40652.5 114912.5 ;
      RECT  40777.5 114777.5 40842.5 114912.5 ;
      RECT  40587.5 115307.5 40652.5 115442.5 ;
      RECT  40967.5 115307.5 41032.5 115442.5 ;
      RECT  40425.0 115072.5 41130.0 115137.5 ;
      RECT  40425.0 115757.5 41130.0 115822.5 ;
      RECT  41482.5 115307.5 41547.5 115822.5 ;
      RECT  41292.5 114777.5 41357.5 114912.5 ;
      RECT  41482.5 114777.5 41547.5 114912.5 ;
      RECT  41482.5 114777.5 41547.5 114912.5 ;
      RECT  41292.5 114777.5 41357.5 114912.5 ;
      RECT  41292.5 115307.5 41357.5 115442.5 ;
      RECT  41482.5 115307.5 41547.5 115442.5 ;
      RECT  41482.5 115307.5 41547.5 115442.5 ;
      RECT  41292.5 115307.5 41357.5 115442.5 ;
      RECT  41482.5 115307.5 41547.5 115442.5 ;
      RECT  41672.5 115307.5 41737.5 115442.5 ;
      RECT  41672.5 115307.5 41737.5 115442.5 ;
      RECT  41482.5 115307.5 41547.5 115442.5 ;
      RECT  41462.5 115072.5 41327.5 115137.5 ;
      RECT  41482.5 115620.0 41547.5 115755.0 ;
      RECT  41292.5 114777.5 41357.5 114912.5 ;
      RECT  41482.5 114777.5 41547.5 114912.5 ;
      RECT  41292.5 115307.5 41357.5 115442.5 ;
      RECT  41672.5 115307.5 41737.5 115442.5 ;
      RECT  41130.0 115072.5 41835.0 115137.5 ;
      RECT  41130.0 115757.5 41835.0 115822.5 ;
      RECT  42187.5 115307.5 42252.5 115822.5 ;
      RECT  41997.5 114777.5 42062.5 114912.5 ;
      RECT  42187.5 114777.5 42252.5 114912.5 ;
      RECT  42187.5 114777.5 42252.5 114912.5 ;
      RECT  41997.5 114777.5 42062.5 114912.5 ;
      RECT  41997.5 115307.5 42062.5 115442.5 ;
      RECT  42187.5 115307.5 42252.5 115442.5 ;
      RECT  42187.5 115307.5 42252.5 115442.5 ;
      RECT  41997.5 115307.5 42062.5 115442.5 ;
      RECT  42187.5 115307.5 42252.5 115442.5 ;
      RECT  42377.5 115307.5 42442.5 115442.5 ;
      RECT  42377.5 115307.5 42442.5 115442.5 ;
      RECT  42187.5 115307.5 42252.5 115442.5 ;
      RECT  42167.5 115072.5 42032.5 115137.5 ;
      RECT  42187.5 115620.0 42252.5 115755.0 ;
      RECT  41997.5 114777.5 42062.5 114912.5 ;
      RECT  42187.5 114777.5 42252.5 114912.5 ;
      RECT  41997.5 115307.5 42062.5 115442.5 ;
      RECT  42377.5 115307.5 42442.5 115442.5 ;
      RECT  41835.0 115072.5 42540.0 115137.5 ;
      RECT  41835.0 115757.5 42540.0 115822.5 ;
      RECT  42892.5 115307.5 42957.5 115822.5 ;
      RECT  42702.5 114777.5 42767.5 114912.5 ;
      RECT  42892.5 114777.5 42957.5 114912.5 ;
      RECT  42892.5 114777.5 42957.5 114912.5 ;
      RECT  42702.5 114777.5 42767.5 114912.5 ;
      RECT  42702.5 115307.5 42767.5 115442.5 ;
      RECT  42892.5 115307.5 42957.5 115442.5 ;
      RECT  42892.5 115307.5 42957.5 115442.5 ;
      RECT  42702.5 115307.5 42767.5 115442.5 ;
      RECT  42892.5 115307.5 42957.5 115442.5 ;
      RECT  43082.5 115307.5 43147.5 115442.5 ;
      RECT  43082.5 115307.5 43147.5 115442.5 ;
      RECT  42892.5 115307.5 42957.5 115442.5 ;
      RECT  42872.5 115072.5 42737.5 115137.5 ;
      RECT  42892.5 115620.0 42957.5 115755.0 ;
      RECT  42702.5 114777.5 42767.5 114912.5 ;
      RECT  42892.5 114777.5 42957.5 114912.5 ;
      RECT  42702.5 115307.5 42767.5 115442.5 ;
      RECT  43082.5 115307.5 43147.5 115442.5 ;
      RECT  42540.0 115072.5 43245.0 115137.5 ;
      RECT  42540.0 115757.5 43245.0 115822.5 ;
      RECT  43597.5 115307.5 43662.5 115822.5 ;
      RECT  43407.5 114777.5 43472.5 114912.5 ;
      RECT  43597.5 114777.5 43662.5 114912.5 ;
      RECT  43597.5 114777.5 43662.5 114912.5 ;
      RECT  43407.5 114777.5 43472.5 114912.5 ;
      RECT  43407.5 115307.5 43472.5 115442.5 ;
      RECT  43597.5 115307.5 43662.5 115442.5 ;
      RECT  43597.5 115307.5 43662.5 115442.5 ;
      RECT  43407.5 115307.5 43472.5 115442.5 ;
      RECT  43597.5 115307.5 43662.5 115442.5 ;
      RECT  43787.5 115307.5 43852.5 115442.5 ;
      RECT  43787.5 115307.5 43852.5 115442.5 ;
      RECT  43597.5 115307.5 43662.5 115442.5 ;
      RECT  43577.5 115072.5 43442.5 115137.5 ;
      RECT  43597.5 115620.0 43662.5 115755.0 ;
      RECT  43407.5 114777.5 43472.5 114912.5 ;
      RECT  43597.5 114777.5 43662.5 114912.5 ;
      RECT  43407.5 115307.5 43472.5 115442.5 ;
      RECT  43787.5 115307.5 43852.5 115442.5 ;
      RECT  43245.0 115072.5 43950.0 115137.5 ;
      RECT  43245.0 115757.5 43950.0 115822.5 ;
      RECT  44302.5 115307.5 44367.5 115822.5 ;
      RECT  44112.5 114777.5 44177.5 114912.5 ;
      RECT  44302.5 114777.5 44367.5 114912.5 ;
      RECT  44302.5 114777.5 44367.5 114912.5 ;
      RECT  44112.5 114777.5 44177.5 114912.5 ;
      RECT  44112.5 115307.5 44177.5 115442.5 ;
      RECT  44302.5 115307.5 44367.5 115442.5 ;
      RECT  44302.5 115307.5 44367.5 115442.5 ;
      RECT  44112.5 115307.5 44177.5 115442.5 ;
      RECT  44302.5 115307.5 44367.5 115442.5 ;
      RECT  44492.5 115307.5 44557.5 115442.5 ;
      RECT  44492.5 115307.5 44557.5 115442.5 ;
      RECT  44302.5 115307.5 44367.5 115442.5 ;
      RECT  44282.5 115072.5 44147.5 115137.5 ;
      RECT  44302.5 115620.0 44367.5 115755.0 ;
      RECT  44112.5 114777.5 44177.5 114912.5 ;
      RECT  44302.5 114777.5 44367.5 114912.5 ;
      RECT  44112.5 115307.5 44177.5 115442.5 ;
      RECT  44492.5 115307.5 44557.5 115442.5 ;
      RECT  43950.0 115072.5 44655.0 115137.5 ;
      RECT  43950.0 115757.5 44655.0 115822.5 ;
      RECT  45007.5 115307.5 45072.5 115822.5 ;
      RECT  44817.5 114777.5 44882.5 114912.5 ;
      RECT  45007.5 114777.5 45072.5 114912.5 ;
      RECT  45007.5 114777.5 45072.5 114912.5 ;
      RECT  44817.5 114777.5 44882.5 114912.5 ;
      RECT  44817.5 115307.5 44882.5 115442.5 ;
      RECT  45007.5 115307.5 45072.5 115442.5 ;
      RECT  45007.5 115307.5 45072.5 115442.5 ;
      RECT  44817.5 115307.5 44882.5 115442.5 ;
      RECT  45007.5 115307.5 45072.5 115442.5 ;
      RECT  45197.5 115307.5 45262.5 115442.5 ;
      RECT  45197.5 115307.5 45262.5 115442.5 ;
      RECT  45007.5 115307.5 45072.5 115442.5 ;
      RECT  44987.5 115072.5 44852.5 115137.5 ;
      RECT  45007.5 115620.0 45072.5 115755.0 ;
      RECT  44817.5 114777.5 44882.5 114912.5 ;
      RECT  45007.5 114777.5 45072.5 114912.5 ;
      RECT  44817.5 115307.5 44882.5 115442.5 ;
      RECT  45197.5 115307.5 45262.5 115442.5 ;
      RECT  44655.0 115072.5 45360.0 115137.5 ;
      RECT  44655.0 115757.5 45360.0 115822.5 ;
      RECT  45712.5 115307.5 45777.5 115822.5 ;
      RECT  45522.5 114777.5 45587.5 114912.5 ;
      RECT  45712.5 114777.5 45777.5 114912.5 ;
      RECT  45712.5 114777.5 45777.5 114912.5 ;
      RECT  45522.5 114777.5 45587.5 114912.5 ;
      RECT  45522.5 115307.5 45587.5 115442.5 ;
      RECT  45712.5 115307.5 45777.5 115442.5 ;
      RECT  45712.5 115307.5 45777.5 115442.5 ;
      RECT  45522.5 115307.5 45587.5 115442.5 ;
      RECT  45712.5 115307.5 45777.5 115442.5 ;
      RECT  45902.5 115307.5 45967.5 115442.5 ;
      RECT  45902.5 115307.5 45967.5 115442.5 ;
      RECT  45712.5 115307.5 45777.5 115442.5 ;
      RECT  45692.5 115072.5 45557.5 115137.5 ;
      RECT  45712.5 115620.0 45777.5 115755.0 ;
      RECT  45522.5 114777.5 45587.5 114912.5 ;
      RECT  45712.5 114777.5 45777.5 114912.5 ;
      RECT  45522.5 115307.5 45587.5 115442.5 ;
      RECT  45902.5 115307.5 45967.5 115442.5 ;
      RECT  45360.0 115072.5 46065.0 115137.5 ;
      RECT  45360.0 115757.5 46065.0 115822.5 ;
      RECT  46417.5 115307.5 46482.5 115822.5 ;
      RECT  46227.5 114777.5 46292.5 114912.5 ;
      RECT  46417.5 114777.5 46482.5 114912.5 ;
      RECT  46417.5 114777.5 46482.5 114912.5 ;
      RECT  46227.5 114777.5 46292.5 114912.5 ;
      RECT  46227.5 115307.5 46292.5 115442.5 ;
      RECT  46417.5 115307.5 46482.5 115442.5 ;
      RECT  46417.5 115307.5 46482.5 115442.5 ;
      RECT  46227.5 115307.5 46292.5 115442.5 ;
      RECT  46417.5 115307.5 46482.5 115442.5 ;
      RECT  46607.5 115307.5 46672.5 115442.5 ;
      RECT  46607.5 115307.5 46672.5 115442.5 ;
      RECT  46417.5 115307.5 46482.5 115442.5 ;
      RECT  46397.5 115072.5 46262.5 115137.5 ;
      RECT  46417.5 115620.0 46482.5 115755.0 ;
      RECT  46227.5 114777.5 46292.5 114912.5 ;
      RECT  46417.5 114777.5 46482.5 114912.5 ;
      RECT  46227.5 115307.5 46292.5 115442.5 ;
      RECT  46607.5 115307.5 46672.5 115442.5 ;
      RECT  46065.0 115072.5 46770.0 115137.5 ;
      RECT  46065.0 115757.5 46770.0 115822.5 ;
      RECT  47122.5 115307.5 47187.5 115822.5 ;
      RECT  46932.5 114777.5 46997.5 114912.5 ;
      RECT  47122.5 114777.5 47187.5 114912.5 ;
      RECT  47122.5 114777.5 47187.5 114912.5 ;
      RECT  46932.5 114777.5 46997.5 114912.5 ;
      RECT  46932.5 115307.5 46997.5 115442.5 ;
      RECT  47122.5 115307.5 47187.5 115442.5 ;
      RECT  47122.5 115307.5 47187.5 115442.5 ;
      RECT  46932.5 115307.5 46997.5 115442.5 ;
      RECT  47122.5 115307.5 47187.5 115442.5 ;
      RECT  47312.5 115307.5 47377.5 115442.5 ;
      RECT  47312.5 115307.5 47377.5 115442.5 ;
      RECT  47122.5 115307.5 47187.5 115442.5 ;
      RECT  47102.5 115072.5 46967.5 115137.5 ;
      RECT  47122.5 115620.0 47187.5 115755.0 ;
      RECT  46932.5 114777.5 46997.5 114912.5 ;
      RECT  47122.5 114777.5 47187.5 114912.5 ;
      RECT  46932.5 115307.5 46997.5 115442.5 ;
      RECT  47312.5 115307.5 47377.5 115442.5 ;
      RECT  46770.0 115072.5 47475.0 115137.5 ;
      RECT  46770.0 115757.5 47475.0 115822.5 ;
      RECT  47827.5 115307.5 47892.5 115822.5 ;
      RECT  47637.5 114777.5 47702.5 114912.5 ;
      RECT  47827.5 114777.5 47892.5 114912.5 ;
      RECT  47827.5 114777.5 47892.5 114912.5 ;
      RECT  47637.5 114777.5 47702.5 114912.5 ;
      RECT  47637.5 115307.5 47702.5 115442.5 ;
      RECT  47827.5 115307.5 47892.5 115442.5 ;
      RECT  47827.5 115307.5 47892.5 115442.5 ;
      RECT  47637.5 115307.5 47702.5 115442.5 ;
      RECT  47827.5 115307.5 47892.5 115442.5 ;
      RECT  48017.5 115307.5 48082.5 115442.5 ;
      RECT  48017.5 115307.5 48082.5 115442.5 ;
      RECT  47827.5 115307.5 47892.5 115442.5 ;
      RECT  47807.5 115072.5 47672.5 115137.5 ;
      RECT  47827.5 115620.0 47892.5 115755.0 ;
      RECT  47637.5 114777.5 47702.5 114912.5 ;
      RECT  47827.5 114777.5 47892.5 114912.5 ;
      RECT  47637.5 115307.5 47702.5 115442.5 ;
      RECT  48017.5 115307.5 48082.5 115442.5 ;
      RECT  47475.0 115072.5 48180.0 115137.5 ;
      RECT  47475.0 115757.5 48180.0 115822.5 ;
      RECT  48532.5 115307.5 48597.5 115822.5 ;
      RECT  48342.5 114777.5 48407.5 114912.5 ;
      RECT  48532.5 114777.5 48597.5 114912.5 ;
      RECT  48532.5 114777.5 48597.5 114912.5 ;
      RECT  48342.5 114777.5 48407.5 114912.5 ;
      RECT  48342.5 115307.5 48407.5 115442.5 ;
      RECT  48532.5 115307.5 48597.5 115442.5 ;
      RECT  48532.5 115307.5 48597.5 115442.5 ;
      RECT  48342.5 115307.5 48407.5 115442.5 ;
      RECT  48532.5 115307.5 48597.5 115442.5 ;
      RECT  48722.5 115307.5 48787.5 115442.5 ;
      RECT  48722.5 115307.5 48787.5 115442.5 ;
      RECT  48532.5 115307.5 48597.5 115442.5 ;
      RECT  48512.5 115072.5 48377.5 115137.5 ;
      RECT  48532.5 115620.0 48597.5 115755.0 ;
      RECT  48342.5 114777.5 48407.5 114912.5 ;
      RECT  48532.5 114777.5 48597.5 114912.5 ;
      RECT  48342.5 115307.5 48407.5 115442.5 ;
      RECT  48722.5 115307.5 48787.5 115442.5 ;
      RECT  48180.0 115072.5 48885.0 115137.5 ;
      RECT  48180.0 115757.5 48885.0 115822.5 ;
      RECT  49237.5 115307.5 49302.5 115822.5 ;
      RECT  49047.5 114777.5 49112.5 114912.5 ;
      RECT  49237.5 114777.5 49302.5 114912.5 ;
      RECT  49237.5 114777.5 49302.5 114912.5 ;
      RECT  49047.5 114777.5 49112.5 114912.5 ;
      RECT  49047.5 115307.5 49112.5 115442.5 ;
      RECT  49237.5 115307.5 49302.5 115442.5 ;
      RECT  49237.5 115307.5 49302.5 115442.5 ;
      RECT  49047.5 115307.5 49112.5 115442.5 ;
      RECT  49237.5 115307.5 49302.5 115442.5 ;
      RECT  49427.5 115307.5 49492.5 115442.5 ;
      RECT  49427.5 115307.5 49492.5 115442.5 ;
      RECT  49237.5 115307.5 49302.5 115442.5 ;
      RECT  49217.5 115072.5 49082.5 115137.5 ;
      RECT  49237.5 115620.0 49302.5 115755.0 ;
      RECT  49047.5 114777.5 49112.5 114912.5 ;
      RECT  49237.5 114777.5 49302.5 114912.5 ;
      RECT  49047.5 115307.5 49112.5 115442.5 ;
      RECT  49427.5 115307.5 49492.5 115442.5 ;
      RECT  48885.0 115072.5 49590.0 115137.5 ;
      RECT  48885.0 115757.5 49590.0 115822.5 ;
      RECT  49942.5 115307.5 50007.5 115822.5 ;
      RECT  49752.5 114777.5 49817.5 114912.5 ;
      RECT  49942.5 114777.5 50007.5 114912.5 ;
      RECT  49942.5 114777.5 50007.5 114912.5 ;
      RECT  49752.5 114777.5 49817.5 114912.5 ;
      RECT  49752.5 115307.5 49817.5 115442.5 ;
      RECT  49942.5 115307.5 50007.5 115442.5 ;
      RECT  49942.5 115307.5 50007.5 115442.5 ;
      RECT  49752.5 115307.5 49817.5 115442.5 ;
      RECT  49942.5 115307.5 50007.5 115442.5 ;
      RECT  50132.5 115307.5 50197.5 115442.5 ;
      RECT  50132.5 115307.5 50197.5 115442.5 ;
      RECT  49942.5 115307.5 50007.5 115442.5 ;
      RECT  49922.5 115072.5 49787.5 115137.5 ;
      RECT  49942.5 115620.0 50007.5 115755.0 ;
      RECT  49752.5 114777.5 49817.5 114912.5 ;
      RECT  49942.5 114777.5 50007.5 114912.5 ;
      RECT  49752.5 115307.5 49817.5 115442.5 ;
      RECT  50132.5 115307.5 50197.5 115442.5 ;
      RECT  49590.0 115072.5 50295.0 115137.5 ;
      RECT  49590.0 115757.5 50295.0 115822.5 ;
      RECT  50647.5 115307.5 50712.5 115822.5 ;
      RECT  50457.5 114777.5 50522.5 114912.5 ;
      RECT  50647.5 114777.5 50712.5 114912.5 ;
      RECT  50647.5 114777.5 50712.5 114912.5 ;
      RECT  50457.5 114777.5 50522.5 114912.5 ;
      RECT  50457.5 115307.5 50522.5 115442.5 ;
      RECT  50647.5 115307.5 50712.5 115442.5 ;
      RECT  50647.5 115307.5 50712.5 115442.5 ;
      RECT  50457.5 115307.5 50522.5 115442.5 ;
      RECT  50647.5 115307.5 50712.5 115442.5 ;
      RECT  50837.5 115307.5 50902.5 115442.5 ;
      RECT  50837.5 115307.5 50902.5 115442.5 ;
      RECT  50647.5 115307.5 50712.5 115442.5 ;
      RECT  50627.5 115072.5 50492.5 115137.5 ;
      RECT  50647.5 115620.0 50712.5 115755.0 ;
      RECT  50457.5 114777.5 50522.5 114912.5 ;
      RECT  50647.5 114777.5 50712.5 114912.5 ;
      RECT  50457.5 115307.5 50522.5 115442.5 ;
      RECT  50837.5 115307.5 50902.5 115442.5 ;
      RECT  50295.0 115072.5 51000.0 115137.5 ;
      RECT  50295.0 115757.5 51000.0 115822.5 ;
      RECT  51352.5 115307.5 51417.5 115822.5 ;
      RECT  51162.5 114777.5 51227.5 114912.5 ;
      RECT  51352.5 114777.5 51417.5 114912.5 ;
      RECT  51352.5 114777.5 51417.5 114912.5 ;
      RECT  51162.5 114777.5 51227.5 114912.5 ;
      RECT  51162.5 115307.5 51227.5 115442.5 ;
      RECT  51352.5 115307.5 51417.5 115442.5 ;
      RECT  51352.5 115307.5 51417.5 115442.5 ;
      RECT  51162.5 115307.5 51227.5 115442.5 ;
      RECT  51352.5 115307.5 51417.5 115442.5 ;
      RECT  51542.5 115307.5 51607.5 115442.5 ;
      RECT  51542.5 115307.5 51607.5 115442.5 ;
      RECT  51352.5 115307.5 51417.5 115442.5 ;
      RECT  51332.5 115072.5 51197.5 115137.5 ;
      RECT  51352.5 115620.0 51417.5 115755.0 ;
      RECT  51162.5 114777.5 51227.5 114912.5 ;
      RECT  51352.5 114777.5 51417.5 114912.5 ;
      RECT  51162.5 115307.5 51227.5 115442.5 ;
      RECT  51542.5 115307.5 51607.5 115442.5 ;
      RECT  51000.0 115072.5 51705.0 115137.5 ;
      RECT  51000.0 115757.5 51705.0 115822.5 ;
      RECT  52057.5 115307.5 52122.5 115822.5 ;
      RECT  51867.5 114777.5 51932.5 114912.5 ;
      RECT  52057.5 114777.5 52122.5 114912.5 ;
      RECT  52057.5 114777.5 52122.5 114912.5 ;
      RECT  51867.5 114777.5 51932.5 114912.5 ;
      RECT  51867.5 115307.5 51932.5 115442.5 ;
      RECT  52057.5 115307.5 52122.5 115442.5 ;
      RECT  52057.5 115307.5 52122.5 115442.5 ;
      RECT  51867.5 115307.5 51932.5 115442.5 ;
      RECT  52057.5 115307.5 52122.5 115442.5 ;
      RECT  52247.5 115307.5 52312.5 115442.5 ;
      RECT  52247.5 115307.5 52312.5 115442.5 ;
      RECT  52057.5 115307.5 52122.5 115442.5 ;
      RECT  52037.5 115072.5 51902.5 115137.5 ;
      RECT  52057.5 115620.0 52122.5 115755.0 ;
      RECT  51867.5 114777.5 51932.5 114912.5 ;
      RECT  52057.5 114777.5 52122.5 114912.5 ;
      RECT  51867.5 115307.5 51932.5 115442.5 ;
      RECT  52247.5 115307.5 52312.5 115442.5 ;
      RECT  51705.0 115072.5 52410.0 115137.5 ;
      RECT  51705.0 115757.5 52410.0 115822.5 ;
      RECT  52762.5 115307.5 52827.5 115822.5 ;
      RECT  52572.5 114777.5 52637.5 114912.5 ;
      RECT  52762.5 114777.5 52827.5 114912.5 ;
      RECT  52762.5 114777.5 52827.5 114912.5 ;
      RECT  52572.5 114777.5 52637.5 114912.5 ;
      RECT  52572.5 115307.5 52637.5 115442.5 ;
      RECT  52762.5 115307.5 52827.5 115442.5 ;
      RECT  52762.5 115307.5 52827.5 115442.5 ;
      RECT  52572.5 115307.5 52637.5 115442.5 ;
      RECT  52762.5 115307.5 52827.5 115442.5 ;
      RECT  52952.5 115307.5 53017.5 115442.5 ;
      RECT  52952.5 115307.5 53017.5 115442.5 ;
      RECT  52762.5 115307.5 52827.5 115442.5 ;
      RECT  52742.5 115072.5 52607.5 115137.5 ;
      RECT  52762.5 115620.0 52827.5 115755.0 ;
      RECT  52572.5 114777.5 52637.5 114912.5 ;
      RECT  52762.5 114777.5 52827.5 114912.5 ;
      RECT  52572.5 115307.5 52637.5 115442.5 ;
      RECT  52952.5 115307.5 53017.5 115442.5 ;
      RECT  52410.0 115072.5 53115.0 115137.5 ;
      RECT  52410.0 115757.5 53115.0 115822.5 ;
      RECT  53467.5 115307.5 53532.5 115822.5 ;
      RECT  53277.5 114777.5 53342.5 114912.5 ;
      RECT  53467.5 114777.5 53532.5 114912.5 ;
      RECT  53467.5 114777.5 53532.5 114912.5 ;
      RECT  53277.5 114777.5 53342.5 114912.5 ;
      RECT  53277.5 115307.5 53342.5 115442.5 ;
      RECT  53467.5 115307.5 53532.5 115442.5 ;
      RECT  53467.5 115307.5 53532.5 115442.5 ;
      RECT  53277.5 115307.5 53342.5 115442.5 ;
      RECT  53467.5 115307.5 53532.5 115442.5 ;
      RECT  53657.5 115307.5 53722.5 115442.5 ;
      RECT  53657.5 115307.5 53722.5 115442.5 ;
      RECT  53467.5 115307.5 53532.5 115442.5 ;
      RECT  53447.5 115072.5 53312.5 115137.5 ;
      RECT  53467.5 115620.0 53532.5 115755.0 ;
      RECT  53277.5 114777.5 53342.5 114912.5 ;
      RECT  53467.5 114777.5 53532.5 114912.5 ;
      RECT  53277.5 115307.5 53342.5 115442.5 ;
      RECT  53657.5 115307.5 53722.5 115442.5 ;
      RECT  53115.0 115072.5 53820.0 115137.5 ;
      RECT  53115.0 115757.5 53820.0 115822.5 ;
      RECT  54172.5 115307.5 54237.5 115822.5 ;
      RECT  53982.5 114777.5 54047.5 114912.5 ;
      RECT  54172.5 114777.5 54237.5 114912.5 ;
      RECT  54172.5 114777.5 54237.5 114912.5 ;
      RECT  53982.5 114777.5 54047.5 114912.5 ;
      RECT  53982.5 115307.5 54047.5 115442.5 ;
      RECT  54172.5 115307.5 54237.5 115442.5 ;
      RECT  54172.5 115307.5 54237.5 115442.5 ;
      RECT  53982.5 115307.5 54047.5 115442.5 ;
      RECT  54172.5 115307.5 54237.5 115442.5 ;
      RECT  54362.5 115307.5 54427.5 115442.5 ;
      RECT  54362.5 115307.5 54427.5 115442.5 ;
      RECT  54172.5 115307.5 54237.5 115442.5 ;
      RECT  54152.5 115072.5 54017.5 115137.5 ;
      RECT  54172.5 115620.0 54237.5 115755.0 ;
      RECT  53982.5 114777.5 54047.5 114912.5 ;
      RECT  54172.5 114777.5 54237.5 114912.5 ;
      RECT  53982.5 115307.5 54047.5 115442.5 ;
      RECT  54362.5 115307.5 54427.5 115442.5 ;
      RECT  53820.0 115072.5 54525.0 115137.5 ;
      RECT  53820.0 115757.5 54525.0 115822.5 ;
      RECT  54877.5 115307.5 54942.5 115822.5 ;
      RECT  54687.5 114777.5 54752.5 114912.5 ;
      RECT  54877.5 114777.5 54942.5 114912.5 ;
      RECT  54877.5 114777.5 54942.5 114912.5 ;
      RECT  54687.5 114777.5 54752.5 114912.5 ;
      RECT  54687.5 115307.5 54752.5 115442.5 ;
      RECT  54877.5 115307.5 54942.5 115442.5 ;
      RECT  54877.5 115307.5 54942.5 115442.5 ;
      RECT  54687.5 115307.5 54752.5 115442.5 ;
      RECT  54877.5 115307.5 54942.5 115442.5 ;
      RECT  55067.5 115307.5 55132.5 115442.5 ;
      RECT  55067.5 115307.5 55132.5 115442.5 ;
      RECT  54877.5 115307.5 54942.5 115442.5 ;
      RECT  54857.5 115072.5 54722.5 115137.5 ;
      RECT  54877.5 115620.0 54942.5 115755.0 ;
      RECT  54687.5 114777.5 54752.5 114912.5 ;
      RECT  54877.5 114777.5 54942.5 114912.5 ;
      RECT  54687.5 115307.5 54752.5 115442.5 ;
      RECT  55067.5 115307.5 55132.5 115442.5 ;
      RECT  54525.0 115072.5 55230.0 115137.5 ;
      RECT  54525.0 115757.5 55230.0 115822.5 ;
      RECT  55582.5 115307.5 55647.5 115822.5 ;
      RECT  55392.5 114777.5 55457.5 114912.5 ;
      RECT  55582.5 114777.5 55647.5 114912.5 ;
      RECT  55582.5 114777.5 55647.5 114912.5 ;
      RECT  55392.5 114777.5 55457.5 114912.5 ;
      RECT  55392.5 115307.5 55457.5 115442.5 ;
      RECT  55582.5 115307.5 55647.5 115442.5 ;
      RECT  55582.5 115307.5 55647.5 115442.5 ;
      RECT  55392.5 115307.5 55457.5 115442.5 ;
      RECT  55582.5 115307.5 55647.5 115442.5 ;
      RECT  55772.5 115307.5 55837.5 115442.5 ;
      RECT  55772.5 115307.5 55837.5 115442.5 ;
      RECT  55582.5 115307.5 55647.5 115442.5 ;
      RECT  55562.5 115072.5 55427.5 115137.5 ;
      RECT  55582.5 115620.0 55647.5 115755.0 ;
      RECT  55392.5 114777.5 55457.5 114912.5 ;
      RECT  55582.5 114777.5 55647.5 114912.5 ;
      RECT  55392.5 115307.5 55457.5 115442.5 ;
      RECT  55772.5 115307.5 55837.5 115442.5 ;
      RECT  55230.0 115072.5 55935.0 115137.5 ;
      RECT  55230.0 115757.5 55935.0 115822.5 ;
      RECT  56287.5 115307.5 56352.5 115822.5 ;
      RECT  56097.5 114777.5 56162.5 114912.5 ;
      RECT  56287.5 114777.5 56352.5 114912.5 ;
      RECT  56287.5 114777.5 56352.5 114912.5 ;
      RECT  56097.5 114777.5 56162.5 114912.5 ;
      RECT  56097.5 115307.5 56162.5 115442.5 ;
      RECT  56287.5 115307.5 56352.5 115442.5 ;
      RECT  56287.5 115307.5 56352.5 115442.5 ;
      RECT  56097.5 115307.5 56162.5 115442.5 ;
      RECT  56287.5 115307.5 56352.5 115442.5 ;
      RECT  56477.5 115307.5 56542.5 115442.5 ;
      RECT  56477.5 115307.5 56542.5 115442.5 ;
      RECT  56287.5 115307.5 56352.5 115442.5 ;
      RECT  56267.5 115072.5 56132.5 115137.5 ;
      RECT  56287.5 115620.0 56352.5 115755.0 ;
      RECT  56097.5 114777.5 56162.5 114912.5 ;
      RECT  56287.5 114777.5 56352.5 114912.5 ;
      RECT  56097.5 115307.5 56162.5 115442.5 ;
      RECT  56477.5 115307.5 56542.5 115442.5 ;
      RECT  55935.0 115072.5 56640.0 115137.5 ;
      RECT  55935.0 115757.5 56640.0 115822.5 ;
      RECT  56992.5 115307.5 57057.5 115822.5 ;
      RECT  56802.5 114777.5 56867.5 114912.5 ;
      RECT  56992.5 114777.5 57057.5 114912.5 ;
      RECT  56992.5 114777.5 57057.5 114912.5 ;
      RECT  56802.5 114777.5 56867.5 114912.5 ;
      RECT  56802.5 115307.5 56867.5 115442.5 ;
      RECT  56992.5 115307.5 57057.5 115442.5 ;
      RECT  56992.5 115307.5 57057.5 115442.5 ;
      RECT  56802.5 115307.5 56867.5 115442.5 ;
      RECT  56992.5 115307.5 57057.5 115442.5 ;
      RECT  57182.5 115307.5 57247.5 115442.5 ;
      RECT  57182.5 115307.5 57247.5 115442.5 ;
      RECT  56992.5 115307.5 57057.5 115442.5 ;
      RECT  56972.5 115072.5 56837.5 115137.5 ;
      RECT  56992.5 115620.0 57057.5 115755.0 ;
      RECT  56802.5 114777.5 56867.5 114912.5 ;
      RECT  56992.5 114777.5 57057.5 114912.5 ;
      RECT  56802.5 115307.5 56867.5 115442.5 ;
      RECT  57182.5 115307.5 57247.5 115442.5 ;
      RECT  56640.0 115072.5 57345.0 115137.5 ;
      RECT  56640.0 115757.5 57345.0 115822.5 ;
      RECT  57697.5 115307.5 57762.5 115822.5 ;
      RECT  57507.5 114777.5 57572.5 114912.5 ;
      RECT  57697.5 114777.5 57762.5 114912.5 ;
      RECT  57697.5 114777.5 57762.5 114912.5 ;
      RECT  57507.5 114777.5 57572.5 114912.5 ;
      RECT  57507.5 115307.5 57572.5 115442.5 ;
      RECT  57697.5 115307.5 57762.5 115442.5 ;
      RECT  57697.5 115307.5 57762.5 115442.5 ;
      RECT  57507.5 115307.5 57572.5 115442.5 ;
      RECT  57697.5 115307.5 57762.5 115442.5 ;
      RECT  57887.5 115307.5 57952.5 115442.5 ;
      RECT  57887.5 115307.5 57952.5 115442.5 ;
      RECT  57697.5 115307.5 57762.5 115442.5 ;
      RECT  57677.5 115072.5 57542.5 115137.5 ;
      RECT  57697.5 115620.0 57762.5 115755.0 ;
      RECT  57507.5 114777.5 57572.5 114912.5 ;
      RECT  57697.5 114777.5 57762.5 114912.5 ;
      RECT  57507.5 115307.5 57572.5 115442.5 ;
      RECT  57887.5 115307.5 57952.5 115442.5 ;
      RECT  57345.0 115072.5 58050.0 115137.5 ;
      RECT  57345.0 115757.5 58050.0 115822.5 ;
      RECT  58402.5 115307.5 58467.5 115822.5 ;
      RECT  58212.5 114777.5 58277.5 114912.5 ;
      RECT  58402.5 114777.5 58467.5 114912.5 ;
      RECT  58402.5 114777.5 58467.5 114912.5 ;
      RECT  58212.5 114777.5 58277.5 114912.5 ;
      RECT  58212.5 115307.5 58277.5 115442.5 ;
      RECT  58402.5 115307.5 58467.5 115442.5 ;
      RECT  58402.5 115307.5 58467.5 115442.5 ;
      RECT  58212.5 115307.5 58277.5 115442.5 ;
      RECT  58402.5 115307.5 58467.5 115442.5 ;
      RECT  58592.5 115307.5 58657.5 115442.5 ;
      RECT  58592.5 115307.5 58657.5 115442.5 ;
      RECT  58402.5 115307.5 58467.5 115442.5 ;
      RECT  58382.5 115072.5 58247.5 115137.5 ;
      RECT  58402.5 115620.0 58467.5 115755.0 ;
      RECT  58212.5 114777.5 58277.5 114912.5 ;
      RECT  58402.5 114777.5 58467.5 114912.5 ;
      RECT  58212.5 115307.5 58277.5 115442.5 ;
      RECT  58592.5 115307.5 58657.5 115442.5 ;
      RECT  58050.0 115072.5 58755.0 115137.5 ;
      RECT  58050.0 115757.5 58755.0 115822.5 ;
      RECT  59107.5 115307.5 59172.5 115822.5 ;
      RECT  58917.5 114777.5 58982.5 114912.5 ;
      RECT  59107.5 114777.5 59172.5 114912.5 ;
      RECT  59107.5 114777.5 59172.5 114912.5 ;
      RECT  58917.5 114777.5 58982.5 114912.5 ;
      RECT  58917.5 115307.5 58982.5 115442.5 ;
      RECT  59107.5 115307.5 59172.5 115442.5 ;
      RECT  59107.5 115307.5 59172.5 115442.5 ;
      RECT  58917.5 115307.5 58982.5 115442.5 ;
      RECT  59107.5 115307.5 59172.5 115442.5 ;
      RECT  59297.5 115307.5 59362.5 115442.5 ;
      RECT  59297.5 115307.5 59362.5 115442.5 ;
      RECT  59107.5 115307.5 59172.5 115442.5 ;
      RECT  59087.5 115072.5 58952.5 115137.5 ;
      RECT  59107.5 115620.0 59172.5 115755.0 ;
      RECT  58917.5 114777.5 58982.5 114912.5 ;
      RECT  59107.5 114777.5 59172.5 114912.5 ;
      RECT  58917.5 115307.5 58982.5 115442.5 ;
      RECT  59297.5 115307.5 59362.5 115442.5 ;
      RECT  58755.0 115072.5 59460.0 115137.5 ;
      RECT  58755.0 115757.5 59460.0 115822.5 ;
      RECT  59812.5 115307.5 59877.5 115822.5 ;
      RECT  59622.5 114777.5 59687.5 114912.5 ;
      RECT  59812.5 114777.5 59877.5 114912.5 ;
      RECT  59812.5 114777.5 59877.5 114912.5 ;
      RECT  59622.5 114777.5 59687.5 114912.5 ;
      RECT  59622.5 115307.5 59687.5 115442.5 ;
      RECT  59812.5 115307.5 59877.5 115442.5 ;
      RECT  59812.5 115307.5 59877.5 115442.5 ;
      RECT  59622.5 115307.5 59687.5 115442.5 ;
      RECT  59812.5 115307.5 59877.5 115442.5 ;
      RECT  60002.5 115307.5 60067.5 115442.5 ;
      RECT  60002.5 115307.5 60067.5 115442.5 ;
      RECT  59812.5 115307.5 59877.5 115442.5 ;
      RECT  59792.5 115072.5 59657.5 115137.5 ;
      RECT  59812.5 115620.0 59877.5 115755.0 ;
      RECT  59622.5 114777.5 59687.5 114912.5 ;
      RECT  59812.5 114777.5 59877.5 114912.5 ;
      RECT  59622.5 115307.5 59687.5 115442.5 ;
      RECT  60002.5 115307.5 60067.5 115442.5 ;
      RECT  59460.0 115072.5 60165.0 115137.5 ;
      RECT  59460.0 115757.5 60165.0 115822.5 ;
      RECT  60517.5 115307.5 60582.5 115822.5 ;
      RECT  60327.5 114777.5 60392.5 114912.5 ;
      RECT  60517.5 114777.5 60582.5 114912.5 ;
      RECT  60517.5 114777.5 60582.5 114912.5 ;
      RECT  60327.5 114777.5 60392.5 114912.5 ;
      RECT  60327.5 115307.5 60392.5 115442.5 ;
      RECT  60517.5 115307.5 60582.5 115442.5 ;
      RECT  60517.5 115307.5 60582.5 115442.5 ;
      RECT  60327.5 115307.5 60392.5 115442.5 ;
      RECT  60517.5 115307.5 60582.5 115442.5 ;
      RECT  60707.5 115307.5 60772.5 115442.5 ;
      RECT  60707.5 115307.5 60772.5 115442.5 ;
      RECT  60517.5 115307.5 60582.5 115442.5 ;
      RECT  60497.5 115072.5 60362.5 115137.5 ;
      RECT  60517.5 115620.0 60582.5 115755.0 ;
      RECT  60327.5 114777.5 60392.5 114912.5 ;
      RECT  60517.5 114777.5 60582.5 114912.5 ;
      RECT  60327.5 115307.5 60392.5 115442.5 ;
      RECT  60707.5 115307.5 60772.5 115442.5 ;
      RECT  60165.0 115072.5 60870.0 115137.5 ;
      RECT  60165.0 115757.5 60870.0 115822.5 ;
      RECT  61222.5 115307.5 61287.5 115822.5 ;
      RECT  61032.5 114777.5 61097.5 114912.5 ;
      RECT  61222.5 114777.5 61287.5 114912.5 ;
      RECT  61222.5 114777.5 61287.5 114912.5 ;
      RECT  61032.5 114777.5 61097.5 114912.5 ;
      RECT  61032.5 115307.5 61097.5 115442.5 ;
      RECT  61222.5 115307.5 61287.5 115442.5 ;
      RECT  61222.5 115307.5 61287.5 115442.5 ;
      RECT  61032.5 115307.5 61097.5 115442.5 ;
      RECT  61222.5 115307.5 61287.5 115442.5 ;
      RECT  61412.5 115307.5 61477.5 115442.5 ;
      RECT  61412.5 115307.5 61477.5 115442.5 ;
      RECT  61222.5 115307.5 61287.5 115442.5 ;
      RECT  61202.5 115072.5 61067.5 115137.5 ;
      RECT  61222.5 115620.0 61287.5 115755.0 ;
      RECT  61032.5 114777.5 61097.5 114912.5 ;
      RECT  61222.5 114777.5 61287.5 114912.5 ;
      RECT  61032.5 115307.5 61097.5 115442.5 ;
      RECT  61412.5 115307.5 61477.5 115442.5 ;
      RECT  60870.0 115072.5 61575.0 115137.5 ;
      RECT  60870.0 115757.5 61575.0 115822.5 ;
      RECT  61927.5 115307.5 61992.5 115822.5 ;
      RECT  61737.5 114777.5 61802.5 114912.5 ;
      RECT  61927.5 114777.5 61992.5 114912.5 ;
      RECT  61927.5 114777.5 61992.5 114912.5 ;
      RECT  61737.5 114777.5 61802.5 114912.5 ;
      RECT  61737.5 115307.5 61802.5 115442.5 ;
      RECT  61927.5 115307.5 61992.5 115442.5 ;
      RECT  61927.5 115307.5 61992.5 115442.5 ;
      RECT  61737.5 115307.5 61802.5 115442.5 ;
      RECT  61927.5 115307.5 61992.5 115442.5 ;
      RECT  62117.5 115307.5 62182.5 115442.5 ;
      RECT  62117.5 115307.5 62182.5 115442.5 ;
      RECT  61927.5 115307.5 61992.5 115442.5 ;
      RECT  61907.5 115072.5 61772.5 115137.5 ;
      RECT  61927.5 115620.0 61992.5 115755.0 ;
      RECT  61737.5 114777.5 61802.5 114912.5 ;
      RECT  61927.5 114777.5 61992.5 114912.5 ;
      RECT  61737.5 115307.5 61802.5 115442.5 ;
      RECT  62117.5 115307.5 62182.5 115442.5 ;
      RECT  61575.0 115072.5 62280.0 115137.5 ;
      RECT  61575.0 115757.5 62280.0 115822.5 ;
      RECT  62632.5 115307.5 62697.5 115822.5 ;
      RECT  62442.5 114777.5 62507.5 114912.5 ;
      RECT  62632.5 114777.5 62697.5 114912.5 ;
      RECT  62632.5 114777.5 62697.5 114912.5 ;
      RECT  62442.5 114777.5 62507.5 114912.5 ;
      RECT  62442.5 115307.5 62507.5 115442.5 ;
      RECT  62632.5 115307.5 62697.5 115442.5 ;
      RECT  62632.5 115307.5 62697.5 115442.5 ;
      RECT  62442.5 115307.5 62507.5 115442.5 ;
      RECT  62632.5 115307.5 62697.5 115442.5 ;
      RECT  62822.5 115307.5 62887.5 115442.5 ;
      RECT  62822.5 115307.5 62887.5 115442.5 ;
      RECT  62632.5 115307.5 62697.5 115442.5 ;
      RECT  62612.5 115072.5 62477.5 115137.5 ;
      RECT  62632.5 115620.0 62697.5 115755.0 ;
      RECT  62442.5 114777.5 62507.5 114912.5 ;
      RECT  62632.5 114777.5 62697.5 114912.5 ;
      RECT  62442.5 115307.5 62507.5 115442.5 ;
      RECT  62822.5 115307.5 62887.5 115442.5 ;
      RECT  62280.0 115072.5 62985.0 115137.5 ;
      RECT  62280.0 115757.5 62985.0 115822.5 ;
      RECT  63337.5 115307.5 63402.5 115822.5 ;
      RECT  63147.5 114777.5 63212.5 114912.5 ;
      RECT  63337.5 114777.5 63402.5 114912.5 ;
      RECT  63337.5 114777.5 63402.5 114912.5 ;
      RECT  63147.5 114777.5 63212.5 114912.5 ;
      RECT  63147.5 115307.5 63212.5 115442.5 ;
      RECT  63337.5 115307.5 63402.5 115442.5 ;
      RECT  63337.5 115307.5 63402.5 115442.5 ;
      RECT  63147.5 115307.5 63212.5 115442.5 ;
      RECT  63337.5 115307.5 63402.5 115442.5 ;
      RECT  63527.5 115307.5 63592.5 115442.5 ;
      RECT  63527.5 115307.5 63592.5 115442.5 ;
      RECT  63337.5 115307.5 63402.5 115442.5 ;
      RECT  63317.5 115072.5 63182.5 115137.5 ;
      RECT  63337.5 115620.0 63402.5 115755.0 ;
      RECT  63147.5 114777.5 63212.5 114912.5 ;
      RECT  63337.5 114777.5 63402.5 114912.5 ;
      RECT  63147.5 115307.5 63212.5 115442.5 ;
      RECT  63527.5 115307.5 63592.5 115442.5 ;
      RECT  62985.0 115072.5 63690.0 115137.5 ;
      RECT  62985.0 115757.5 63690.0 115822.5 ;
      RECT  64042.5 115307.5 64107.5 115822.5 ;
      RECT  63852.5 114777.5 63917.5 114912.5 ;
      RECT  64042.5 114777.5 64107.5 114912.5 ;
      RECT  64042.5 114777.5 64107.5 114912.5 ;
      RECT  63852.5 114777.5 63917.5 114912.5 ;
      RECT  63852.5 115307.5 63917.5 115442.5 ;
      RECT  64042.5 115307.5 64107.5 115442.5 ;
      RECT  64042.5 115307.5 64107.5 115442.5 ;
      RECT  63852.5 115307.5 63917.5 115442.5 ;
      RECT  64042.5 115307.5 64107.5 115442.5 ;
      RECT  64232.5 115307.5 64297.5 115442.5 ;
      RECT  64232.5 115307.5 64297.5 115442.5 ;
      RECT  64042.5 115307.5 64107.5 115442.5 ;
      RECT  64022.5 115072.5 63887.5 115137.5 ;
      RECT  64042.5 115620.0 64107.5 115755.0 ;
      RECT  63852.5 114777.5 63917.5 114912.5 ;
      RECT  64042.5 114777.5 64107.5 114912.5 ;
      RECT  63852.5 115307.5 63917.5 115442.5 ;
      RECT  64232.5 115307.5 64297.5 115442.5 ;
      RECT  63690.0 115072.5 64395.0 115137.5 ;
      RECT  63690.0 115757.5 64395.0 115822.5 ;
      RECT  64747.5 115307.5 64812.5 115822.5 ;
      RECT  64557.5 114777.5 64622.5 114912.5 ;
      RECT  64747.5 114777.5 64812.5 114912.5 ;
      RECT  64747.5 114777.5 64812.5 114912.5 ;
      RECT  64557.5 114777.5 64622.5 114912.5 ;
      RECT  64557.5 115307.5 64622.5 115442.5 ;
      RECT  64747.5 115307.5 64812.5 115442.5 ;
      RECT  64747.5 115307.5 64812.5 115442.5 ;
      RECT  64557.5 115307.5 64622.5 115442.5 ;
      RECT  64747.5 115307.5 64812.5 115442.5 ;
      RECT  64937.5 115307.5 65002.5 115442.5 ;
      RECT  64937.5 115307.5 65002.5 115442.5 ;
      RECT  64747.5 115307.5 64812.5 115442.5 ;
      RECT  64727.5 115072.5 64592.5 115137.5 ;
      RECT  64747.5 115620.0 64812.5 115755.0 ;
      RECT  64557.5 114777.5 64622.5 114912.5 ;
      RECT  64747.5 114777.5 64812.5 114912.5 ;
      RECT  64557.5 115307.5 64622.5 115442.5 ;
      RECT  64937.5 115307.5 65002.5 115442.5 ;
      RECT  64395.0 115072.5 65100.0 115137.5 ;
      RECT  64395.0 115757.5 65100.0 115822.5 ;
      RECT  65452.5 115307.5 65517.5 115822.5 ;
      RECT  65262.5 114777.5 65327.5 114912.5 ;
      RECT  65452.5 114777.5 65517.5 114912.5 ;
      RECT  65452.5 114777.5 65517.5 114912.5 ;
      RECT  65262.5 114777.5 65327.5 114912.5 ;
      RECT  65262.5 115307.5 65327.5 115442.5 ;
      RECT  65452.5 115307.5 65517.5 115442.5 ;
      RECT  65452.5 115307.5 65517.5 115442.5 ;
      RECT  65262.5 115307.5 65327.5 115442.5 ;
      RECT  65452.5 115307.5 65517.5 115442.5 ;
      RECT  65642.5 115307.5 65707.5 115442.5 ;
      RECT  65642.5 115307.5 65707.5 115442.5 ;
      RECT  65452.5 115307.5 65517.5 115442.5 ;
      RECT  65432.5 115072.5 65297.5 115137.5 ;
      RECT  65452.5 115620.0 65517.5 115755.0 ;
      RECT  65262.5 114777.5 65327.5 114912.5 ;
      RECT  65452.5 114777.5 65517.5 114912.5 ;
      RECT  65262.5 115307.5 65327.5 115442.5 ;
      RECT  65642.5 115307.5 65707.5 115442.5 ;
      RECT  65100.0 115072.5 65805.0 115137.5 ;
      RECT  65100.0 115757.5 65805.0 115822.5 ;
      RECT  66157.5 115307.5 66222.5 115822.5 ;
      RECT  65967.5 114777.5 66032.5 114912.5 ;
      RECT  66157.5 114777.5 66222.5 114912.5 ;
      RECT  66157.5 114777.5 66222.5 114912.5 ;
      RECT  65967.5 114777.5 66032.5 114912.5 ;
      RECT  65967.5 115307.5 66032.5 115442.5 ;
      RECT  66157.5 115307.5 66222.5 115442.5 ;
      RECT  66157.5 115307.5 66222.5 115442.5 ;
      RECT  65967.5 115307.5 66032.5 115442.5 ;
      RECT  66157.5 115307.5 66222.5 115442.5 ;
      RECT  66347.5 115307.5 66412.5 115442.5 ;
      RECT  66347.5 115307.5 66412.5 115442.5 ;
      RECT  66157.5 115307.5 66222.5 115442.5 ;
      RECT  66137.5 115072.5 66002.5 115137.5 ;
      RECT  66157.5 115620.0 66222.5 115755.0 ;
      RECT  65967.5 114777.5 66032.5 114912.5 ;
      RECT  66157.5 114777.5 66222.5 114912.5 ;
      RECT  65967.5 115307.5 66032.5 115442.5 ;
      RECT  66347.5 115307.5 66412.5 115442.5 ;
      RECT  65805.0 115072.5 66510.0 115137.5 ;
      RECT  65805.0 115757.5 66510.0 115822.5 ;
      RECT  66862.5 115307.5 66927.5 115822.5 ;
      RECT  66672.5 114777.5 66737.5 114912.5 ;
      RECT  66862.5 114777.5 66927.5 114912.5 ;
      RECT  66862.5 114777.5 66927.5 114912.5 ;
      RECT  66672.5 114777.5 66737.5 114912.5 ;
      RECT  66672.5 115307.5 66737.5 115442.5 ;
      RECT  66862.5 115307.5 66927.5 115442.5 ;
      RECT  66862.5 115307.5 66927.5 115442.5 ;
      RECT  66672.5 115307.5 66737.5 115442.5 ;
      RECT  66862.5 115307.5 66927.5 115442.5 ;
      RECT  67052.5 115307.5 67117.5 115442.5 ;
      RECT  67052.5 115307.5 67117.5 115442.5 ;
      RECT  66862.5 115307.5 66927.5 115442.5 ;
      RECT  66842.5 115072.5 66707.5 115137.5 ;
      RECT  66862.5 115620.0 66927.5 115755.0 ;
      RECT  66672.5 114777.5 66737.5 114912.5 ;
      RECT  66862.5 114777.5 66927.5 114912.5 ;
      RECT  66672.5 115307.5 66737.5 115442.5 ;
      RECT  67052.5 115307.5 67117.5 115442.5 ;
      RECT  66510.0 115072.5 67215.0 115137.5 ;
      RECT  66510.0 115757.5 67215.0 115822.5 ;
      RECT  67567.5 115307.5 67632.5 115822.5 ;
      RECT  67377.5 114777.5 67442.5 114912.5 ;
      RECT  67567.5 114777.5 67632.5 114912.5 ;
      RECT  67567.5 114777.5 67632.5 114912.5 ;
      RECT  67377.5 114777.5 67442.5 114912.5 ;
      RECT  67377.5 115307.5 67442.5 115442.5 ;
      RECT  67567.5 115307.5 67632.5 115442.5 ;
      RECT  67567.5 115307.5 67632.5 115442.5 ;
      RECT  67377.5 115307.5 67442.5 115442.5 ;
      RECT  67567.5 115307.5 67632.5 115442.5 ;
      RECT  67757.5 115307.5 67822.5 115442.5 ;
      RECT  67757.5 115307.5 67822.5 115442.5 ;
      RECT  67567.5 115307.5 67632.5 115442.5 ;
      RECT  67547.5 115072.5 67412.5 115137.5 ;
      RECT  67567.5 115620.0 67632.5 115755.0 ;
      RECT  67377.5 114777.5 67442.5 114912.5 ;
      RECT  67567.5 114777.5 67632.5 114912.5 ;
      RECT  67377.5 115307.5 67442.5 115442.5 ;
      RECT  67757.5 115307.5 67822.5 115442.5 ;
      RECT  67215.0 115072.5 67920.0 115137.5 ;
      RECT  67215.0 115757.5 67920.0 115822.5 ;
      RECT  68272.5 115307.5 68337.5 115822.5 ;
      RECT  68082.5 114777.5 68147.5 114912.5 ;
      RECT  68272.5 114777.5 68337.5 114912.5 ;
      RECT  68272.5 114777.5 68337.5 114912.5 ;
      RECT  68082.5 114777.5 68147.5 114912.5 ;
      RECT  68082.5 115307.5 68147.5 115442.5 ;
      RECT  68272.5 115307.5 68337.5 115442.5 ;
      RECT  68272.5 115307.5 68337.5 115442.5 ;
      RECT  68082.5 115307.5 68147.5 115442.5 ;
      RECT  68272.5 115307.5 68337.5 115442.5 ;
      RECT  68462.5 115307.5 68527.5 115442.5 ;
      RECT  68462.5 115307.5 68527.5 115442.5 ;
      RECT  68272.5 115307.5 68337.5 115442.5 ;
      RECT  68252.5 115072.5 68117.5 115137.5 ;
      RECT  68272.5 115620.0 68337.5 115755.0 ;
      RECT  68082.5 114777.5 68147.5 114912.5 ;
      RECT  68272.5 114777.5 68337.5 114912.5 ;
      RECT  68082.5 115307.5 68147.5 115442.5 ;
      RECT  68462.5 115307.5 68527.5 115442.5 ;
      RECT  67920.0 115072.5 68625.0 115137.5 ;
      RECT  67920.0 115757.5 68625.0 115822.5 ;
      RECT  68977.5 115307.5 69042.5 115822.5 ;
      RECT  68787.5 114777.5 68852.5 114912.5 ;
      RECT  68977.5 114777.5 69042.5 114912.5 ;
      RECT  68977.5 114777.5 69042.5 114912.5 ;
      RECT  68787.5 114777.5 68852.5 114912.5 ;
      RECT  68787.5 115307.5 68852.5 115442.5 ;
      RECT  68977.5 115307.5 69042.5 115442.5 ;
      RECT  68977.5 115307.5 69042.5 115442.5 ;
      RECT  68787.5 115307.5 68852.5 115442.5 ;
      RECT  68977.5 115307.5 69042.5 115442.5 ;
      RECT  69167.5 115307.5 69232.5 115442.5 ;
      RECT  69167.5 115307.5 69232.5 115442.5 ;
      RECT  68977.5 115307.5 69042.5 115442.5 ;
      RECT  68957.5 115072.5 68822.5 115137.5 ;
      RECT  68977.5 115620.0 69042.5 115755.0 ;
      RECT  68787.5 114777.5 68852.5 114912.5 ;
      RECT  68977.5 114777.5 69042.5 114912.5 ;
      RECT  68787.5 115307.5 68852.5 115442.5 ;
      RECT  69167.5 115307.5 69232.5 115442.5 ;
      RECT  68625.0 115072.5 69330.0 115137.5 ;
      RECT  68625.0 115757.5 69330.0 115822.5 ;
      RECT  69682.5 115307.5 69747.5 115822.5 ;
      RECT  69492.5 114777.5 69557.5 114912.5 ;
      RECT  69682.5 114777.5 69747.5 114912.5 ;
      RECT  69682.5 114777.5 69747.5 114912.5 ;
      RECT  69492.5 114777.5 69557.5 114912.5 ;
      RECT  69492.5 115307.5 69557.5 115442.5 ;
      RECT  69682.5 115307.5 69747.5 115442.5 ;
      RECT  69682.5 115307.5 69747.5 115442.5 ;
      RECT  69492.5 115307.5 69557.5 115442.5 ;
      RECT  69682.5 115307.5 69747.5 115442.5 ;
      RECT  69872.5 115307.5 69937.5 115442.5 ;
      RECT  69872.5 115307.5 69937.5 115442.5 ;
      RECT  69682.5 115307.5 69747.5 115442.5 ;
      RECT  69662.5 115072.5 69527.5 115137.5 ;
      RECT  69682.5 115620.0 69747.5 115755.0 ;
      RECT  69492.5 114777.5 69557.5 114912.5 ;
      RECT  69682.5 114777.5 69747.5 114912.5 ;
      RECT  69492.5 115307.5 69557.5 115442.5 ;
      RECT  69872.5 115307.5 69937.5 115442.5 ;
      RECT  69330.0 115072.5 70035.0 115137.5 ;
      RECT  69330.0 115757.5 70035.0 115822.5 ;
      RECT  70387.5 115307.5 70452.5 115822.5 ;
      RECT  70197.5 114777.5 70262.5 114912.5 ;
      RECT  70387.5 114777.5 70452.5 114912.5 ;
      RECT  70387.5 114777.5 70452.5 114912.5 ;
      RECT  70197.5 114777.5 70262.5 114912.5 ;
      RECT  70197.5 115307.5 70262.5 115442.5 ;
      RECT  70387.5 115307.5 70452.5 115442.5 ;
      RECT  70387.5 115307.5 70452.5 115442.5 ;
      RECT  70197.5 115307.5 70262.5 115442.5 ;
      RECT  70387.5 115307.5 70452.5 115442.5 ;
      RECT  70577.5 115307.5 70642.5 115442.5 ;
      RECT  70577.5 115307.5 70642.5 115442.5 ;
      RECT  70387.5 115307.5 70452.5 115442.5 ;
      RECT  70367.5 115072.5 70232.5 115137.5 ;
      RECT  70387.5 115620.0 70452.5 115755.0 ;
      RECT  70197.5 114777.5 70262.5 114912.5 ;
      RECT  70387.5 114777.5 70452.5 114912.5 ;
      RECT  70197.5 115307.5 70262.5 115442.5 ;
      RECT  70577.5 115307.5 70642.5 115442.5 ;
      RECT  70035.0 115072.5 70740.0 115137.5 ;
      RECT  70035.0 115757.5 70740.0 115822.5 ;
      RECT  71092.5 115307.5 71157.5 115822.5 ;
      RECT  70902.5 114777.5 70967.5 114912.5 ;
      RECT  71092.5 114777.5 71157.5 114912.5 ;
      RECT  71092.5 114777.5 71157.5 114912.5 ;
      RECT  70902.5 114777.5 70967.5 114912.5 ;
      RECT  70902.5 115307.5 70967.5 115442.5 ;
      RECT  71092.5 115307.5 71157.5 115442.5 ;
      RECT  71092.5 115307.5 71157.5 115442.5 ;
      RECT  70902.5 115307.5 70967.5 115442.5 ;
      RECT  71092.5 115307.5 71157.5 115442.5 ;
      RECT  71282.5 115307.5 71347.5 115442.5 ;
      RECT  71282.5 115307.5 71347.5 115442.5 ;
      RECT  71092.5 115307.5 71157.5 115442.5 ;
      RECT  71072.5 115072.5 70937.5 115137.5 ;
      RECT  71092.5 115620.0 71157.5 115755.0 ;
      RECT  70902.5 114777.5 70967.5 114912.5 ;
      RECT  71092.5 114777.5 71157.5 114912.5 ;
      RECT  70902.5 115307.5 70967.5 115442.5 ;
      RECT  71282.5 115307.5 71347.5 115442.5 ;
      RECT  70740.0 115072.5 71445.0 115137.5 ;
      RECT  70740.0 115757.5 71445.0 115822.5 ;
      RECT  71797.5 115307.5 71862.5 115822.5 ;
      RECT  71607.5 114777.5 71672.5 114912.5 ;
      RECT  71797.5 114777.5 71862.5 114912.5 ;
      RECT  71797.5 114777.5 71862.5 114912.5 ;
      RECT  71607.5 114777.5 71672.5 114912.5 ;
      RECT  71607.5 115307.5 71672.5 115442.5 ;
      RECT  71797.5 115307.5 71862.5 115442.5 ;
      RECT  71797.5 115307.5 71862.5 115442.5 ;
      RECT  71607.5 115307.5 71672.5 115442.5 ;
      RECT  71797.5 115307.5 71862.5 115442.5 ;
      RECT  71987.5 115307.5 72052.5 115442.5 ;
      RECT  71987.5 115307.5 72052.5 115442.5 ;
      RECT  71797.5 115307.5 71862.5 115442.5 ;
      RECT  71777.5 115072.5 71642.5 115137.5 ;
      RECT  71797.5 115620.0 71862.5 115755.0 ;
      RECT  71607.5 114777.5 71672.5 114912.5 ;
      RECT  71797.5 114777.5 71862.5 114912.5 ;
      RECT  71607.5 115307.5 71672.5 115442.5 ;
      RECT  71987.5 115307.5 72052.5 115442.5 ;
      RECT  71445.0 115072.5 72150.0 115137.5 ;
      RECT  71445.0 115757.5 72150.0 115822.5 ;
      RECT  72502.5 115307.5 72567.5 115822.5 ;
      RECT  72312.5 114777.5 72377.5 114912.5 ;
      RECT  72502.5 114777.5 72567.5 114912.5 ;
      RECT  72502.5 114777.5 72567.5 114912.5 ;
      RECT  72312.5 114777.5 72377.5 114912.5 ;
      RECT  72312.5 115307.5 72377.5 115442.5 ;
      RECT  72502.5 115307.5 72567.5 115442.5 ;
      RECT  72502.5 115307.5 72567.5 115442.5 ;
      RECT  72312.5 115307.5 72377.5 115442.5 ;
      RECT  72502.5 115307.5 72567.5 115442.5 ;
      RECT  72692.5 115307.5 72757.5 115442.5 ;
      RECT  72692.5 115307.5 72757.5 115442.5 ;
      RECT  72502.5 115307.5 72567.5 115442.5 ;
      RECT  72482.5 115072.5 72347.5 115137.5 ;
      RECT  72502.5 115620.0 72567.5 115755.0 ;
      RECT  72312.5 114777.5 72377.5 114912.5 ;
      RECT  72502.5 114777.5 72567.5 114912.5 ;
      RECT  72312.5 115307.5 72377.5 115442.5 ;
      RECT  72692.5 115307.5 72757.5 115442.5 ;
      RECT  72150.0 115072.5 72855.0 115137.5 ;
      RECT  72150.0 115757.5 72855.0 115822.5 ;
      RECT  73207.5 115307.5 73272.5 115822.5 ;
      RECT  73017.5 114777.5 73082.5 114912.5 ;
      RECT  73207.5 114777.5 73272.5 114912.5 ;
      RECT  73207.5 114777.5 73272.5 114912.5 ;
      RECT  73017.5 114777.5 73082.5 114912.5 ;
      RECT  73017.5 115307.5 73082.5 115442.5 ;
      RECT  73207.5 115307.5 73272.5 115442.5 ;
      RECT  73207.5 115307.5 73272.5 115442.5 ;
      RECT  73017.5 115307.5 73082.5 115442.5 ;
      RECT  73207.5 115307.5 73272.5 115442.5 ;
      RECT  73397.5 115307.5 73462.5 115442.5 ;
      RECT  73397.5 115307.5 73462.5 115442.5 ;
      RECT  73207.5 115307.5 73272.5 115442.5 ;
      RECT  73187.5 115072.5 73052.5 115137.5 ;
      RECT  73207.5 115620.0 73272.5 115755.0 ;
      RECT  73017.5 114777.5 73082.5 114912.5 ;
      RECT  73207.5 114777.5 73272.5 114912.5 ;
      RECT  73017.5 115307.5 73082.5 115442.5 ;
      RECT  73397.5 115307.5 73462.5 115442.5 ;
      RECT  72855.0 115072.5 73560.0 115137.5 ;
      RECT  72855.0 115757.5 73560.0 115822.5 ;
      RECT  73912.5 115307.5 73977.5 115822.5 ;
      RECT  73722.5 114777.5 73787.5 114912.5 ;
      RECT  73912.5 114777.5 73977.5 114912.5 ;
      RECT  73912.5 114777.5 73977.5 114912.5 ;
      RECT  73722.5 114777.5 73787.5 114912.5 ;
      RECT  73722.5 115307.5 73787.5 115442.5 ;
      RECT  73912.5 115307.5 73977.5 115442.5 ;
      RECT  73912.5 115307.5 73977.5 115442.5 ;
      RECT  73722.5 115307.5 73787.5 115442.5 ;
      RECT  73912.5 115307.5 73977.5 115442.5 ;
      RECT  74102.5 115307.5 74167.5 115442.5 ;
      RECT  74102.5 115307.5 74167.5 115442.5 ;
      RECT  73912.5 115307.5 73977.5 115442.5 ;
      RECT  73892.5 115072.5 73757.5 115137.5 ;
      RECT  73912.5 115620.0 73977.5 115755.0 ;
      RECT  73722.5 114777.5 73787.5 114912.5 ;
      RECT  73912.5 114777.5 73977.5 114912.5 ;
      RECT  73722.5 115307.5 73787.5 115442.5 ;
      RECT  74102.5 115307.5 74167.5 115442.5 ;
      RECT  73560.0 115072.5 74265.0 115137.5 ;
      RECT  73560.0 115757.5 74265.0 115822.5 ;
      RECT  74617.5 115307.5 74682.5 115822.5 ;
      RECT  74427.5 114777.5 74492.5 114912.5 ;
      RECT  74617.5 114777.5 74682.5 114912.5 ;
      RECT  74617.5 114777.5 74682.5 114912.5 ;
      RECT  74427.5 114777.5 74492.5 114912.5 ;
      RECT  74427.5 115307.5 74492.5 115442.5 ;
      RECT  74617.5 115307.5 74682.5 115442.5 ;
      RECT  74617.5 115307.5 74682.5 115442.5 ;
      RECT  74427.5 115307.5 74492.5 115442.5 ;
      RECT  74617.5 115307.5 74682.5 115442.5 ;
      RECT  74807.5 115307.5 74872.5 115442.5 ;
      RECT  74807.5 115307.5 74872.5 115442.5 ;
      RECT  74617.5 115307.5 74682.5 115442.5 ;
      RECT  74597.5 115072.5 74462.5 115137.5 ;
      RECT  74617.5 115620.0 74682.5 115755.0 ;
      RECT  74427.5 114777.5 74492.5 114912.5 ;
      RECT  74617.5 114777.5 74682.5 114912.5 ;
      RECT  74427.5 115307.5 74492.5 115442.5 ;
      RECT  74807.5 115307.5 74872.5 115442.5 ;
      RECT  74265.0 115072.5 74970.0 115137.5 ;
      RECT  74265.0 115757.5 74970.0 115822.5 ;
      RECT  75322.5 115307.5 75387.5 115822.5 ;
      RECT  75132.5 114777.5 75197.5 114912.5 ;
      RECT  75322.5 114777.5 75387.5 114912.5 ;
      RECT  75322.5 114777.5 75387.5 114912.5 ;
      RECT  75132.5 114777.5 75197.5 114912.5 ;
      RECT  75132.5 115307.5 75197.5 115442.5 ;
      RECT  75322.5 115307.5 75387.5 115442.5 ;
      RECT  75322.5 115307.5 75387.5 115442.5 ;
      RECT  75132.5 115307.5 75197.5 115442.5 ;
      RECT  75322.5 115307.5 75387.5 115442.5 ;
      RECT  75512.5 115307.5 75577.5 115442.5 ;
      RECT  75512.5 115307.5 75577.5 115442.5 ;
      RECT  75322.5 115307.5 75387.5 115442.5 ;
      RECT  75302.5 115072.5 75167.5 115137.5 ;
      RECT  75322.5 115620.0 75387.5 115755.0 ;
      RECT  75132.5 114777.5 75197.5 114912.5 ;
      RECT  75322.5 114777.5 75387.5 114912.5 ;
      RECT  75132.5 115307.5 75197.5 115442.5 ;
      RECT  75512.5 115307.5 75577.5 115442.5 ;
      RECT  74970.0 115072.5 75675.0 115137.5 ;
      RECT  74970.0 115757.5 75675.0 115822.5 ;
      RECT  76027.5 115307.5 76092.5 115822.5 ;
      RECT  75837.5 114777.5 75902.5 114912.5 ;
      RECT  76027.5 114777.5 76092.5 114912.5 ;
      RECT  76027.5 114777.5 76092.5 114912.5 ;
      RECT  75837.5 114777.5 75902.5 114912.5 ;
      RECT  75837.5 115307.5 75902.5 115442.5 ;
      RECT  76027.5 115307.5 76092.5 115442.5 ;
      RECT  76027.5 115307.5 76092.5 115442.5 ;
      RECT  75837.5 115307.5 75902.5 115442.5 ;
      RECT  76027.5 115307.5 76092.5 115442.5 ;
      RECT  76217.5 115307.5 76282.5 115442.5 ;
      RECT  76217.5 115307.5 76282.5 115442.5 ;
      RECT  76027.5 115307.5 76092.5 115442.5 ;
      RECT  76007.5 115072.5 75872.5 115137.5 ;
      RECT  76027.5 115620.0 76092.5 115755.0 ;
      RECT  75837.5 114777.5 75902.5 114912.5 ;
      RECT  76027.5 114777.5 76092.5 114912.5 ;
      RECT  75837.5 115307.5 75902.5 115442.5 ;
      RECT  76217.5 115307.5 76282.5 115442.5 ;
      RECT  75675.0 115072.5 76380.0 115137.5 ;
      RECT  75675.0 115757.5 76380.0 115822.5 ;
      RECT  76732.5 115307.5 76797.5 115822.5 ;
      RECT  76542.5 114777.5 76607.5 114912.5 ;
      RECT  76732.5 114777.5 76797.5 114912.5 ;
      RECT  76732.5 114777.5 76797.5 114912.5 ;
      RECT  76542.5 114777.5 76607.5 114912.5 ;
      RECT  76542.5 115307.5 76607.5 115442.5 ;
      RECT  76732.5 115307.5 76797.5 115442.5 ;
      RECT  76732.5 115307.5 76797.5 115442.5 ;
      RECT  76542.5 115307.5 76607.5 115442.5 ;
      RECT  76732.5 115307.5 76797.5 115442.5 ;
      RECT  76922.5 115307.5 76987.5 115442.5 ;
      RECT  76922.5 115307.5 76987.5 115442.5 ;
      RECT  76732.5 115307.5 76797.5 115442.5 ;
      RECT  76712.5 115072.5 76577.5 115137.5 ;
      RECT  76732.5 115620.0 76797.5 115755.0 ;
      RECT  76542.5 114777.5 76607.5 114912.5 ;
      RECT  76732.5 114777.5 76797.5 114912.5 ;
      RECT  76542.5 115307.5 76607.5 115442.5 ;
      RECT  76922.5 115307.5 76987.5 115442.5 ;
      RECT  76380.0 115072.5 77085.0 115137.5 ;
      RECT  76380.0 115757.5 77085.0 115822.5 ;
      RECT  77437.5 115307.5 77502.5 115822.5 ;
      RECT  77247.5 114777.5 77312.5 114912.5 ;
      RECT  77437.5 114777.5 77502.5 114912.5 ;
      RECT  77437.5 114777.5 77502.5 114912.5 ;
      RECT  77247.5 114777.5 77312.5 114912.5 ;
      RECT  77247.5 115307.5 77312.5 115442.5 ;
      RECT  77437.5 115307.5 77502.5 115442.5 ;
      RECT  77437.5 115307.5 77502.5 115442.5 ;
      RECT  77247.5 115307.5 77312.5 115442.5 ;
      RECT  77437.5 115307.5 77502.5 115442.5 ;
      RECT  77627.5 115307.5 77692.5 115442.5 ;
      RECT  77627.5 115307.5 77692.5 115442.5 ;
      RECT  77437.5 115307.5 77502.5 115442.5 ;
      RECT  77417.5 115072.5 77282.5 115137.5 ;
      RECT  77437.5 115620.0 77502.5 115755.0 ;
      RECT  77247.5 114777.5 77312.5 114912.5 ;
      RECT  77437.5 114777.5 77502.5 114912.5 ;
      RECT  77247.5 115307.5 77312.5 115442.5 ;
      RECT  77627.5 115307.5 77692.5 115442.5 ;
      RECT  77085.0 115072.5 77790.0 115137.5 ;
      RECT  77085.0 115757.5 77790.0 115822.5 ;
      RECT  78142.5 115307.5 78207.5 115822.5 ;
      RECT  77952.5 114777.5 78017.5 114912.5 ;
      RECT  78142.5 114777.5 78207.5 114912.5 ;
      RECT  78142.5 114777.5 78207.5 114912.5 ;
      RECT  77952.5 114777.5 78017.5 114912.5 ;
      RECT  77952.5 115307.5 78017.5 115442.5 ;
      RECT  78142.5 115307.5 78207.5 115442.5 ;
      RECT  78142.5 115307.5 78207.5 115442.5 ;
      RECT  77952.5 115307.5 78017.5 115442.5 ;
      RECT  78142.5 115307.5 78207.5 115442.5 ;
      RECT  78332.5 115307.5 78397.5 115442.5 ;
      RECT  78332.5 115307.5 78397.5 115442.5 ;
      RECT  78142.5 115307.5 78207.5 115442.5 ;
      RECT  78122.5 115072.5 77987.5 115137.5 ;
      RECT  78142.5 115620.0 78207.5 115755.0 ;
      RECT  77952.5 114777.5 78017.5 114912.5 ;
      RECT  78142.5 114777.5 78207.5 114912.5 ;
      RECT  77952.5 115307.5 78017.5 115442.5 ;
      RECT  78332.5 115307.5 78397.5 115442.5 ;
      RECT  77790.0 115072.5 78495.0 115137.5 ;
      RECT  77790.0 115757.5 78495.0 115822.5 ;
      RECT  78847.5 115307.5 78912.5 115822.5 ;
      RECT  78657.5 114777.5 78722.5 114912.5 ;
      RECT  78847.5 114777.5 78912.5 114912.5 ;
      RECT  78847.5 114777.5 78912.5 114912.5 ;
      RECT  78657.5 114777.5 78722.5 114912.5 ;
      RECT  78657.5 115307.5 78722.5 115442.5 ;
      RECT  78847.5 115307.5 78912.5 115442.5 ;
      RECT  78847.5 115307.5 78912.5 115442.5 ;
      RECT  78657.5 115307.5 78722.5 115442.5 ;
      RECT  78847.5 115307.5 78912.5 115442.5 ;
      RECT  79037.5 115307.5 79102.5 115442.5 ;
      RECT  79037.5 115307.5 79102.5 115442.5 ;
      RECT  78847.5 115307.5 78912.5 115442.5 ;
      RECT  78827.5 115072.5 78692.5 115137.5 ;
      RECT  78847.5 115620.0 78912.5 115755.0 ;
      RECT  78657.5 114777.5 78722.5 114912.5 ;
      RECT  78847.5 114777.5 78912.5 114912.5 ;
      RECT  78657.5 115307.5 78722.5 115442.5 ;
      RECT  79037.5 115307.5 79102.5 115442.5 ;
      RECT  78495.0 115072.5 79200.0 115137.5 ;
      RECT  78495.0 115757.5 79200.0 115822.5 ;
      RECT  79552.5 115307.5 79617.5 115822.5 ;
      RECT  79362.5 114777.5 79427.5 114912.5 ;
      RECT  79552.5 114777.5 79617.5 114912.5 ;
      RECT  79552.5 114777.5 79617.5 114912.5 ;
      RECT  79362.5 114777.5 79427.5 114912.5 ;
      RECT  79362.5 115307.5 79427.5 115442.5 ;
      RECT  79552.5 115307.5 79617.5 115442.5 ;
      RECT  79552.5 115307.5 79617.5 115442.5 ;
      RECT  79362.5 115307.5 79427.5 115442.5 ;
      RECT  79552.5 115307.5 79617.5 115442.5 ;
      RECT  79742.5 115307.5 79807.5 115442.5 ;
      RECT  79742.5 115307.5 79807.5 115442.5 ;
      RECT  79552.5 115307.5 79617.5 115442.5 ;
      RECT  79532.5 115072.5 79397.5 115137.5 ;
      RECT  79552.5 115620.0 79617.5 115755.0 ;
      RECT  79362.5 114777.5 79427.5 114912.5 ;
      RECT  79552.5 114777.5 79617.5 114912.5 ;
      RECT  79362.5 115307.5 79427.5 115442.5 ;
      RECT  79742.5 115307.5 79807.5 115442.5 ;
      RECT  79200.0 115072.5 79905.0 115137.5 ;
      RECT  79200.0 115757.5 79905.0 115822.5 ;
      RECT  80257.5 115307.5 80322.5 115822.5 ;
      RECT  80067.5 114777.5 80132.5 114912.5 ;
      RECT  80257.5 114777.5 80322.5 114912.5 ;
      RECT  80257.5 114777.5 80322.5 114912.5 ;
      RECT  80067.5 114777.5 80132.5 114912.5 ;
      RECT  80067.5 115307.5 80132.5 115442.5 ;
      RECT  80257.5 115307.5 80322.5 115442.5 ;
      RECT  80257.5 115307.5 80322.5 115442.5 ;
      RECT  80067.5 115307.5 80132.5 115442.5 ;
      RECT  80257.5 115307.5 80322.5 115442.5 ;
      RECT  80447.5 115307.5 80512.5 115442.5 ;
      RECT  80447.5 115307.5 80512.5 115442.5 ;
      RECT  80257.5 115307.5 80322.5 115442.5 ;
      RECT  80237.5 115072.5 80102.5 115137.5 ;
      RECT  80257.5 115620.0 80322.5 115755.0 ;
      RECT  80067.5 114777.5 80132.5 114912.5 ;
      RECT  80257.5 114777.5 80322.5 114912.5 ;
      RECT  80067.5 115307.5 80132.5 115442.5 ;
      RECT  80447.5 115307.5 80512.5 115442.5 ;
      RECT  79905.0 115072.5 80610.0 115137.5 ;
      RECT  79905.0 115757.5 80610.0 115822.5 ;
      RECT  80962.5 115307.5 81027.5 115822.5 ;
      RECT  80772.5 114777.5 80837.5 114912.5 ;
      RECT  80962.5 114777.5 81027.5 114912.5 ;
      RECT  80962.5 114777.5 81027.5 114912.5 ;
      RECT  80772.5 114777.5 80837.5 114912.5 ;
      RECT  80772.5 115307.5 80837.5 115442.5 ;
      RECT  80962.5 115307.5 81027.5 115442.5 ;
      RECT  80962.5 115307.5 81027.5 115442.5 ;
      RECT  80772.5 115307.5 80837.5 115442.5 ;
      RECT  80962.5 115307.5 81027.5 115442.5 ;
      RECT  81152.5 115307.5 81217.5 115442.5 ;
      RECT  81152.5 115307.5 81217.5 115442.5 ;
      RECT  80962.5 115307.5 81027.5 115442.5 ;
      RECT  80942.5 115072.5 80807.5 115137.5 ;
      RECT  80962.5 115620.0 81027.5 115755.0 ;
      RECT  80772.5 114777.5 80837.5 114912.5 ;
      RECT  80962.5 114777.5 81027.5 114912.5 ;
      RECT  80772.5 115307.5 80837.5 115442.5 ;
      RECT  81152.5 115307.5 81217.5 115442.5 ;
      RECT  80610.0 115072.5 81315.0 115137.5 ;
      RECT  80610.0 115757.5 81315.0 115822.5 ;
      RECT  81667.5 115307.5 81732.5 115822.5 ;
      RECT  81477.5 114777.5 81542.5 114912.5 ;
      RECT  81667.5 114777.5 81732.5 114912.5 ;
      RECT  81667.5 114777.5 81732.5 114912.5 ;
      RECT  81477.5 114777.5 81542.5 114912.5 ;
      RECT  81477.5 115307.5 81542.5 115442.5 ;
      RECT  81667.5 115307.5 81732.5 115442.5 ;
      RECT  81667.5 115307.5 81732.5 115442.5 ;
      RECT  81477.5 115307.5 81542.5 115442.5 ;
      RECT  81667.5 115307.5 81732.5 115442.5 ;
      RECT  81857.5 115307.5 81922.5 115442.5 ;
      RECT  81857.5 115307.5 81922.5 115442.5 ;
      RECT  81667.5 115307.5 81732.5 115442.5 ;
      RECT  81647.5 115072.5 81512.5 115137.5 ;
      RECT  81667.5 115620.0 81732.5 115755.0 ;
      RECT  81477.5 114777.5 81542.5 114912.5 ;
      RECT  81667.5 114777.5 81732.5 114912.5 ;
      RECT  81477.5 115307.5 81542.5 115442.5 ;
      RECT  81857.5 115307.5 81922.5 115442.5 ;
      RECT  81315.0 115072.5 82020.0 115137.5 ;
      RECT  81315.0 115757.5 82020.0 115822.5 ;
      RECT  82372.5 115307.5 82437.5 115822.5 ;
      RECT  82182.5 114777.5 82247.5 114912.5 ;
      RECT  82372.5 114777.5 82437.5 114912.5 ;
      RECT  82372.5 114777.5 82437.5 114912.5 ;
      RECT  82182.5 114777.5 82247.5 114912.5 ;
      RECT  82182.5 115307.5 82247.5 115442.5 ;
      RECT  82372.5 115307.5 82437.5 115442.5 ;
      RECT  82372.5 115307.5 82437.5 115442.5 ;
      RECT  82182.5 115307.5 82247.5 115442.5 ;
      RECT  82372.5 115307.5 82437.5 115442.5 ;
      RECT  82562.5 115307.5 82627.5 115442.5 ;
      RECT  82562.5 115307.5 82627.5 115442.5 ;
      RECT  82372.5 115307.5 82437.5 115442.5 ;
      RECT  82352.5 115072.5 82217.5 115137.5 ;
      RECT  82372.5 115620.0 82437.5 115755.0 ;
      RECT  82182.5 114777.5 82247.5 114912.5 ;
      RECT  82372.5 114777.5 82437.5 114912.5 ;
      RECT  82182.5 115307.5 82247.5 115442.5 ;
      RECT  82562.5 115307.5 82627.5 115442.5 ;
      RECT  82020.0 115072.5 82725.0 115137.5 ;
      RECT  82020.0 115757.5 82725.0 115822.5 ;
      RECT  83077.5 115307.5 83142.5 115822.5 ;
      RECT  82887.5 114777.5 82952.5 114912.5 ;
      RECT  83077.5 114777.5 83142.5 114912.5 ;
      RECT  83077.5 114777.5 83142.5 114912.5 ;
      RECT  82887.5 114777.5 82952.5 114912.5 ;
      RECT  82887.5 115307.5 82952.5 115442.5 ;
      RECT  83077.5 115307.5 83142.5 115442.5 ;
      RECT  83077.5 115307.5 83142.5 115442.5 ;
      RECT  82887.5 115307.5 82952.5 115442.5 ;
      RECT  83077.5 115307.5 83142.5 115442.5 ;
      RECT  83267.5 115307.5 83332.5 115442.5 ;
      RECT  83267.5 115307.5 83332.5 115442.5 ;
      RECT  83077.5 115307.5 83142.5 115442.5 ;
      RECT  83057.5 115072.5 82922.5 115137.5 ;
      RECT  83077.5 115620.0 83142.5 115755.0 ;
      RECT  82887.5 114777.5 82952.5 114912.5 ;
      RECT  83077.5 114777.5 83142.5 114912.5 ;
      RECT  82887.5 115307.5 82952.5 115442.5 ;
      RECT  83267.5 115307.5 83332.5 115442.5 ;
      RECT  82725.0 115072.5 83430.0 115137.5 ;
      RECT  82725.0 115757.5 83430.0 115822.5 ;
      RECT  83782.5 115307.5 83847.5 115822.5 ;
      RECT  83592.5 114777.5 83657.5 114912.5 ;
      RECT  83782.5 114777.5 83847.5 114912.5 ;
      RECT  83782.5 114777.5 83847.5 114912.5 ;
      RECT  83592.5 114777.5 83657.5 114912.5 ;
      RECT  83592.5 115307.5 83657.5 115442.5 ;
      RECT  83782.5 115307.5 83847.5 115442.5 ;
      RECT  83782.5 115307.5 83847.5 115442.5 ;
      RECT  83592.5 115307.5 83657.5 115442.5 ;
      RECT  83782.5 115307.5 83847.5 115442.5 ;
      RECT  83972.5 115307.5 84037.5 115442.5 ;
      RECT  83972.5 115307.5 84037.5 115442.5 ;
      RECT  83782.5 115307.5 83847.5 115442.5 ;
      RECT  83762.5 115072.5 83627.5 115137.5 ;
      RECT  83782.5 115620.0 83847.5 115755.0 ;
      RECT  83592.5 114777.5 83657.5 114912.5 ;
      RECT  83782.5 114777.5 83847.5 114912.5 ;
      RECT  83592.5 115307.5 83657.5 115442.5 ;
      RECT  83972.5 115307.5 84037.5 115442.5 ;
      RECT  83430.0 115072.5 84135.0 115137.5 ;
      RECT  83430.0 115757.5 84135.0 115822.5 ;
      RECT  84487.5 115307.5 84552.5 115822.5 ;
      RECT  84297.5 114777.5 84362.5 114912.5 ;
      RECT  84487.5 114777.5 84552.5 114912.5 ;
      RECT  84487.5 114777.5 84552.5 114912.5 ;
      RECT  84297.5 114777.5 84362.5 114912.5 ;
      RECT  84297.5 115307.5 84362.5 115442.5 ;
      RECT  84487.5 115307.5 84552.5 115442.5 ;
      RECT  84487.5 115307.5 84552.5 115442.5 ;
      RECT  84297.5 115307.5 84362.5 115442.5 ;
      RECT  84487.5 115307.5 84552.5 115442.5 ;
      RECT  84677.5 115307.5 84742.5 115442.5 ;
      RECT  84677.5 115307.5 84742.5 115442.5 ;
      RECT  84487.5 115307.5 84552.5 115442.5 ;
      RECT  84467.5 115072.5 84332.5 115137.5 ;
      RECT  84487.5 115620.0 84552.5 115755.0 ;
      RECT  84297.5 114777.5 84362.5 114912.5 ;
      RECT  84487.5 114777.5 84552.5 114912.5 ;
      RECT  84297.5 115307.5 84362.5 115442.5 ;
      RECT  84677.5 115307.5 84742.5 115442.5 ;
      RECT  84135.0 115072.5 84840.0 115137.5 ;
      RECT  84135.0 115757.5 84840.0 115822.5 ;
      RECT  85192.5 115307.5 85257.5 115822.5 ;
      RECT  85002.5 114777.5 85067.5 114912.5 ;
      RECT  85192.5 114777.5 85257.5 114912.5 ;
      RECT  85192.5 114777.5 85257.5 114912.5 ;
      RECT  85002.5 114777.5 85067.5 114912.5 ;
      RECT  85002.5 115307.5 85067.5 115442.5 ;
      RECT  85192.5 115307.5 85257.5 115442.5 ;
      RECT  85192.5 115307.5 85257.5 115442.5 ;
      RECT  85002.5 115307.5 85067.5 115442.5 ;
      RECT  85192.5 115307.5 85257.5 115442.5 ;
      RECT  85382.5 115307.5 85447.5 115442.5 ;
      RECT  85382.5 115307.5 85447.5 115442.5 ;
      RECT  85192.5 115307.5 85257.5 115442.5 ;
      RECT  85172.5 115072.5 85037.5 115137.5 ;
      RECT  85192.5 115620.0 85257.5 115755.0 ;
      RECT  85002.5 114777.5 85067.5 114912.5 ;
      RECT  85192.5 114777.5 85257.5 114912.5 ;
      RECT  85002.5 115307.5 85067.5 115442.5 ;
      RECT  85382.5 115307.5 85447.5 115442.5 ;
      RECT  84840.0 115072.5 85545.0 115137.5 ;
      RECT  84840.0 115757.5 85545.0 115822.5 ;
      RECT  85897.5 115307.5 85962.5 115822.5 ;
      RECT  85707.5 114777.5 85772.5 114912.5 ;
      RECT  85897.5 114777.5 85962.5 114912.5 ;
      RECT  85897.5 114777.5 85962.5 114912.5 ;
      RECT  85707.5 114777.5 85772.5 114912.5 ;
      RECT  85707.5 115307.5 85772.5 115442.5 ;
      RECT  85897.5 115307.5 85962.5 115442.5 ;
      RECT  85897.5 115307.5 85962.5 115442.5 ;
      RECT  85707.5 115307.5 85772.5 115442.5 ;
      RECT  85897.5 115307.5 85962.5 115442.5 ;
      RECT  86087.5 115307.5 86152.5 115442.5 ;
      RECT  86087.5 115307.5 86152.5 115442.5 ;
      RECT  85897.5 115307.5 85962.5 115442.5 ;
      RECT  85877.5 115072.5 85742.5 115137.5 ;
      RECT  85897.5 115620.0 85962.5 115755.0 ;
      RECT  85707.5 114777.5 85772.5 114912.5 ;
      RECT  85897.5 114777.5 85962.5 114912.5 ;
      RECT  85707.5 115307.5 85772.5 115442.5 ;
      RECT  86087.5 115307.5 86152.5 115442.5 ;
      RECT  85545.0 115072.5 86250.0 115137.5 ;
      RECT  85545.0 115757.5 86250.0 115822.5 ;
      RECT  86602.5 115307.5 86667.5 115822.5 ;
      RECT  86412.5 114777.5 86477.5 114912.5 ;
      RECT  86602.5 114777.5 86667.5 114912.5 ;
      RECT  86602.5 114777.5 86667.5 114912.5 ;
      RECT  86412.5 114777.5 86477.5 114912.5 ;
      RECT  86412.5 115307.5 86477.5 115442.5 ;
      RECT  86602.5 115307.5 86667.5 115442.5 ;
      RECT  86602.5 115307.5 86667.5 115442.5 ;
      RECT  86412.5 115307.5 86477.5 115442.5 ;
      RECT  86602.5 115307.5 86667.5 115442.5 ;
      RECT  86792.5 115307.5 86857.5 115442.5 ;
      RECT  86792.5 115307.5 86857.5 115442.5 ;
      RECT  86602.5 115307.5 86667.5 115442.5 ;
      RECT  86582.5 115072.5 86447.5 115137.5 ;
      RECT  86602.5 115620.0 86667.5 115755.0 ;
      RECT  86412.5 114777.5 86477.5 114912.5 ;
      RECT  86602.5 114777.5 86667.5 114912.5 ;
      RECT  86412.5 115307.5 86477.5 115442.5 ;
      RECT  86792.5 115307.5 86857.5 115442.5 ;
      RECT  86250.0 115072.5 86955.0 115137.5 ;
      RECT  86250.0 115757.5 86955.0 115822.5 ;
      RECT  87307.5 115307.5 87372.5 115822.5 ;
      RECT  87117.5 114777.5 87182.5 114912.5 ;
      RECT  87307.5 114777.5 87372.5 114912.5 ;
      RECT  87307.5 114777.5 87372.5 114912.5 ;
      RECT  87117.5 114777.5 87182.5 114912.5 ;
      RECT  87117.5 115307.5 87182.5 115442.5 ;
      RECT  87307.5 115307.5 87372.5 115442.5 ;
      RECT  87307.5 115307.5 87372.5 115442.5 ;
      RECT  87117.5 115307.5 87182.5 115442.5 ;
      RECT  87307.5 115307.5 87372.5 115442.5 ;
      RECT  87497.5 115307.5 87562.5 115442.5 ;
      RECT  87497.5 115307.5 87562.5 115442.5 ;
      RECT  87307.5 115307.5 87372.5 115442.5 ;
      RECT  87287.5 115072.5 87152.5 115137.5 ;
      RECT  87307.5 115620.0 87372.5 115755.0 ;
      RECT  87117.5 114777.5 87182.5 114912.5 ;
      RECT  87307.5 114777.5 87372.5 114912.5 ;
      RECT  87117.5 115307.5 87182.5 115442.5 ;
      RECT  87497.5 115307.5 87562.5 115442.5 ;
      RECT  86955.0 115072.5 87660.0 115137.5 ;
      RECT  86955.0 115757.5 87660.0 115822.5 ;
      RECT  88012.5 115307.5 88077.5 115822.5 ;
      RECT  87822.5 114777.5 87887.5 114912.5 ;
      RECT  88012.5 114777.5 88077.5 114912.5 ;
      RECT  88012.5 114777.5 88077.5 114912.5 ;
      RECT  87822.5 114777.5 87887.5 114912.5 ;
      RECT  87822.5 115307.5 87887.5 115442.5 ;
      RECT  88012.5 115307.5 88077.5 115442.5 ;
      RECT  88012.5 115307.5 88077.5 115442.5 ;
      RECT  87822.5 115307.5 87887.5 115442.5 ;
      RECT  88012.5 115307.5 88077.5 115442.5 ;
      RECT  88202.5 115307.5 88267.5 115442.5 ;
      RECT  88202.5 115307.5 88267.5 115442.5 ;
      RECT  88012.5 115307.5 88077.5 115442.5 ;
      RECT  87992.5 115072.5 87857.5 115137.5 ;
      RECT  88012.5 115620.0 88077.5 115755.0 ;
      RECT  87822.5 114777.5 87887.5 114912.5 ;
      RECT  88012.5 114777.5 88077.5 114912.5 ;
      RECT  87822.5 115307.5 87887.5 115442.5 ;
      RECT  88202.5 115307.5 88267.5 115442.5 ;
      RECT  87660.0 115072.5 88365.0 115137.5 ;
      RECT  87660.0 115757.5 88365.0 115822.5 ;
      RECT  88717.5 115307.5 88782.5 115822.5 ;
      RECT  88527.5 114777.5 88592.5 114912.5 ;
      RECT  88717.5 114777.5 88782.5 114912.5 ;
      RECT  88717.5 114777.5 88782.5 114912.5 ;
      RECT  88527.5 114777.5 88592.5 114912.5 ;
      RECT  88527.5 115307.5 88592.5 115442.5 ;
      RECT  88717.5 115307.5 88782.5 115442.5 ;
      RECT  88717.5 115307.5 88782.5 115442.5 ;
      RECT  88527.5 115307.5 88592.5 115442.5 ;
      RECT  88717.5 115307.5 88782.5 115442.5 ;
      RECT  88907.5 115307.5 88972.5 115442.5 ;
      RECT  88907.5 115307.5 88972.5 115442.5 ;
      RECT  88717.5 115307.5 88782.5 115442.5 ;
      RECT  88697.5 115072.5 88562.5 115137.5 ;
      RECT  88717.5 115620.0 88782.5 115755.0 ;
      RECT  88527.5 114777.5 88592.5 114912.5 ;
      RECT  88717.5 114777.5 88782.5 114912.5 ;
      RECT  88527.5 115307.5 88592.5 115442.5 ;
      RECT  88907.5 115307.5 88972.5 115442.5 ;
      RECT  88365.0 115072.5 89070.0 115137.5 ;
      RECT  88365.0 115757.5 89070.0 115822.5 ;
      RECT  89422.5 115307.5 89487.5 115822.5 ;
      RECT  89232.5 114777.5 89297.5 114912.5 ;
      RECT  89422.5 114777.5 89487.5 114912.5 ;
      RECT  89422.5 114777.5 89487.5 114912.5 ;
      RECT  89232.5 114777.5 89297.5 114912.5 ;
      RECT  89232.5 115307.5 89297.5 115442.5 ;
      RECT  89422.5 115307.5 89487.5 115442.5 ;
      RECT  89422.5 115307.5 89487.5 115442.5 ;
      RECT  89232.5 115307.5 89297.5 115442.5 ;
      RECT  89422.5 115307.5 89487.5 115442.5 ;
      RECT  89612.5 115307.5 89677.5 115442.5 ;
      RECT  89612.5 115307.5 89677.5 115442.5 ;
      RECT  89422.5 115307.5 89487.5 115442.5 ;
      RECT  89402.5 115072.5 89267.5 115137.5 ;
      RECT  89422.5 115620.0 89487.5 115755.0 ;
      RECT  89232.5 114777.5 89297.5 114912.5 ;
      RECT  89422.5 114777.5 89487.5 114912.5 ;
      RECT  89232.5 115307.5 89297.5 115442.5 ;
      RECT  89612.5 115307.5 89677.5 115442.5 ;
      RECT  89070.0 115072.5 89775.0 115137.5 ;
      RECT  89070.0 115757.5 89775.0 115822.5 ;
      RECT  90127.5 115307.5 90192.5 115822.5 ;
      RECT  89937.5 114777.5 90002.5 114912.5 ;
      RECT  90127.5 114777.5 90192.5 114912.5 ;
      RECT  90127.5 114777.5 90192.5 114912.5 ;
      RECT  89937.5 114777.5 90002.5 114912.5 ;
      RECT  89937.5 115307.5 90002.5 115442.5 ;
      RECT  90127.5 115307.5 90192.5 115442.5 ;
      RECT  90127.5 115307.5 90192.5 115442.5 ;
      RECT  89937.5 115307.5 90002.5 115442.5 ;
      RECT  90127.5 115307.5 90192.5 115442.5 ;
      RECT  90317.5 115307.5 90382.5 115442.5 ;
      RECT  90317.5 115307.5 90382.5 115442.5 ;
      RECT  90127.5 115307.5 90192.5 115442.5 ;
      RECT  90107.5 115072.5 89972.5 115137.5 ;
      RECT  90127.5 115620.0 90192.5 115755.0 ;
      RECT  89937.5 114777.5 90002.5 114912.5 ;
      RECT  90127.5 114777.5 90192.5 114912.5 ;
      RECT  89937.5 115307.5 90002.5 115442.5 ;
      RECT  90317.5 115307.5 90382.5 115442.5 ;
      RECT  89775.0 115072.5 90480.0 115137.5 ;
      RECT  89775.0 115757.5 90480.0 115822.5 ;
      RECT  90832.5 115307.5 90897.5 115822.5 ;
      RECT  90642.5 114777.5 90707.5 114912.5 ;
      RECT  90832.5 114777.5 90897.5 114912.5 ;
      RECT  90832.5 114777.5 90897.5 114912.5 ;
      RECT  90642.5 114777.5 90707.5 114912.5 ;
      RECT  90642.5 115307.5 90707.5 115442.5 ;
      RECT  90832.5 115307.5 90897.5 115442.5 ;
      RECT  90832.5 115307.5 90897.5 115442.5 ;
      RECT  90642.5 115307.5 90707.5 115442.5 ;
      RECT  90832.5 115307.5 90897.5 115442.5 ;
      RECT  91022.5 115307.5 91087.5 115442.5 ;
      RECT  91022.5 115307.5 91087.5 115442.5 ;
      RECT  90832.5 115307.5 90897.5 115442.5 ;
      RECT  90812.5 115072.5 90677.5 115137.5 ;
      RECT  90832.5 115620.0 90897.5 115755.0 ;
      RECT  90642.5 114777.5 90707.5 114912.5 ;
      RECT  90832.5 114777.5 90897.5 114912.5 ;
      RECT  90642.5 115307.5 90707.5 115442.5 ;
      RECT  91022.5 115307.5 91087.5 115442.5 ;
      RECT  90480.0 115072.5 91185.0 115137.5 ;
      RECT  90480.0 115757.5 91185.0 115822.5 ;
      RECT  91537.5 115307.5 91602.5 115822.5 ;
      RECT  91347.5 114777.5 91412.5 114912.5 ;
      RECT  91537.5 114777.5 91602.5 114912.5 ;
      RECT  91537.5 114777.5 91602.5 114912.5 ;
      RECT  91347.5 114777.5 91412.5 114912.5 ;
      RECT  91347.5 115307.5 91412.5 115442.5 ;
      RECT  91537.5 115307.5 91602.5 115442.5 ;
      RECT  91537.5 115307.5 91602.5 115442.5 ;
      RECT  91347.5 115307.5 91412.5 115442.5 ;
      RECT  91537.5 115307.5 91602.5 115442.5 ;
      RECT  91727.5 115307.5 91792.5 115442.5 ;
      RECT  91727.5 115307.5 91792.5 115442.5 ;
      RECT  91537.5 115307.5 91602.5 115442.5 ;
      RECT  91517.5 115072.5 91382.5 115137.5 ;
      RECT  91537.5 115620.0 91602.5 115755.0 ;
      RECT  91347.5 114777.5 91412.5 114912.5 ;
      RECT  91537.5 114777.5 91602.5 114912.5 ;
      RECT  91347.5 115307.5 91412.5 115442.5 ;
      RECT  91727.5 115307.5 91792.5 115442.5 ;
      RECT  91185.0 115072.5 91890.0 115137.5 ;
      RECT  91185.0 115757.5 91890.0 115822.5 ;
      RECT  92242.5 115307.5 92307.5 115822.5 ;
      RECT  92052.5 114777.5 92117.5 114912.5 ;
      RECT  92242.5 114777.5 92307.5 114912.5 ;
      RECT  92242.5 114777.5 92307.5 114912.5 ;
      RECT  92052.5 114777.5 92117.5 114912.5 ;
      RECT  92052.5 115307.5 92117.5 115442.5 ;
      RECT  92242.5 115307.5 92307.5 115442.5 ;
      RECT  92242.5 115307.5 92307.5 115442.5 ;
      RECT  92052.5 115307.5 92117.5 115442.5 ;
      RECT  92242.5 115307.5 92307.5 115442.5 ;
      RECT  92432.5 115307.5 92497.5 115442.5 ;
      RECT  92432.5 115307.5 92497.5 115442.5 ;
      RECT  92242.5 115307.5 92307.5 115442.5 ;
      RECT  92222.5 115072.5 92087.5 115137.5 ;
      RECT  92242.5 115620.0 92307.5 115755.0 ;
      RECT  92052.5 114777.5 92117.5 114912.5 ;
      RECT  92242.5 114777.5 92307.5 114912.5 ;
      RECT  92052.5 115307.5 92117.5 115442.5 ;
      RECT  92432.5 115307.5 92497.5 115442.5 ;
      RECT  91890.0 115072.5 92595.0 115137.5 ;
      RECT  91890.0 115757.5 92595.0 115822.5 ;
      RECT  92947.5 115307.5 93012.5 115822.5 ;
      RECT  92757.5 114777.5 92822.5 114912.5 ;
      RECT  92947.5 114777.5 93012.5 114912.5 ;
      RECT  92947.5 114777.5 93012.5 114912.5 ;
      RECT  92757.5 114777.5 92822.5 114912.5 ;
      RECT  92757.5 115307.5 92822.5 115442.5 ;
      RECT  92947.5 115307.5 93012.5 115442.5 ;
      RECT  92947.5 115307.5 93012.5 115442.5 ;
      RECT  92757.5 115307.5 92822.5 115442.5 ;
      RECT  92947.5 115307.5 93012.5 115442.5 ;
      RECT  93137.5 115307.5 93202.5 115442.5 ;
      RECT  93137.5 115307.5 93202.5 115442.5 ;
      RECT  92947.5 115307.5 93012.5 115442.5 ;
      RECT  92927.5 115072.5 92792.5 115137.5 ;
      RECT  92947.5 115620.0 93012.5 115755.0 ;
      RECT  92757.5 114777.5 92822.5 114912.5 ;
      RECT  92947.5 114777.5 93012.5 114912.5 ;
      RECT  92757.5 115307.5 92822.5 115442.5 ;
      RECT  93137.5 115307.5 93202.5 115442.5 ;
      RECT  92595.0 115072.5 93300.0 115137.5 ;
      RECT  92595.0 115757.5 93300.0 115822.5 ;
      RECT  93652.5 115307.5 93717.5 115822.5 ;
      RECT  93462.5 114777.5 93527.5 114912.5 ;
      RECT  93652.5 114777.5 93717.5 114912.5 ;
      RECT  93652.5 114777.5 93717.5 114912.5 ;
      RECT  93462.5 114777.5 93527.5 114912.5 ;
      RECT  93462.5 115307.5 93527.5 115442.5 ;
      RECT  93652.5 115307.5 93717.5 115442.5 ;
      RECT  93652.5 115307.5 93717.5 115442.5 ;
      RECT  93462.5 115307.5 93527.5 115442.5 ;
      RECT  93652.5 115307.5 93717.5 115442.5 ;
      RECT  93842.5 115307.5 93907.5 115442.5 ;
      RECT  93842.5 115307.5 93907.5 115442.5 ;
      RECT  93652.5 115307.5 93717.5 115442.5 ;
      RECT  93632.5 115072.5 93497.5 115137.5 ;
      RECT  93652.5 115620.0 93717.5 115755.0 ;
      RECT  93462.5 114777.5 93527.5 114912.5 ;
      RECT  93652.5 114777.5 93717.5 114912.5 ;
      RECT  93462.5 115307.5 93527.5 115442.5 ;
      RECT  93842.5 115307.5 93907.5 115442.5 ;
      RECT  93300.0 115072.5 94005.0 115137.5 ;
      RECT  93300.0 115757.5 94005.0 115822.5 ;
      RECT  94357.5 115307.5 94422.5 115822.5 ;
      RECT  94167.5 114777.5 94232.5 114912.5 ;
      RECT  94357.5 114777.5 94422.5 114912.5 ;
      RECT  94357.5 114777.5 94422.5 114912.5 ;
      RECT  94167.5 114777.5 94232.5 114912.5 ;
      RECT  94167.5 115307.5 94232.5 115442.5 ;
      RECT  94357.5 115307.5 94422.5 115442.5 ;
      RECT  94357.5 115307.5 94422.5 115442.5 ;
      RECT  94167.5 115307.5 94232.5 115442.5 ;
      RECT  94357.5 115307.5 94422.5 115442.5 ;
      RECT  94547.5 115307.5 94612.5 115442.5 ;
      RECT  94547.5 115307.5 94612.5 115442.5 ;
      RECT  94357.5 115307.5 94422.5 115442.5 ;
      RECT  94337.5 115072.5 94202.5 115137.5 ;
      RECT  94357.5 115620.0 94422.5 115755.0 ;
      RECT  94167.5 114777.5 94232.5 114912.5 ;
      RECT  94357.5 114777.5 94422.5 114912.5 ;
      RECT  94167.5 115307.5 94232.5 115442.5 ;
      RECT  94547.5 115307.5 94612.5 115442.5 ;
      RECT  94005.0 115072.5 94710.0 115137.5 ;
      RECT  94005.0 115757.5 94710.0 115822.5 ;
      RECT  95062.5 115307.5 95127.5 115822.5 ;
      RECT  94872.5 114777.5 94937.5 114912.5 ;
      RECT  95062.5 114777.5 95127.5 114912.5 ;
      RECT  95062.5 114777.5 95127.5 114912.5 ;
      RECT  94872.5 114777.5 94937.5 114912.5 ;
      RECT  94872.5 115307.5 94937.5 115442.5 ;
      RECT  95062.5 115307.5 95127.5 115442.5 ;
      RECT  95062.5 115307.5 95127.5 115442.5 ;
      RECT  94872.5 115307.5 94937.5 115442.5 ;
      RECT  95062.5 115307.5 95127.5 115442.5 ;
      RECT  95252.5 115307.5 95317.5 115442.5 ;
      RECT  95252.5 115307.5 95317.5 115442.5 ;
      RECT  95062.5 115307.5 95127.5 115442.5 ;
      RECT  95042.5 115072.5 94907.5 115137.5 ;
      RECT  95062.5 115620.0 95127.5 115755.0 ;
      RECT  94872.5 114777.5 94937.5 114912.5 ;
      RECT  95062.5 114777.5 95127.5 114912.5 ;
      RECT  94872.5 115307.5 94937.5 115442.5 ;
      RECT  95252.5 115307.5 95317.5 115442.5 ;
      RECT  94710.0 115072.5 95415.0 115137.5 ;
      RECT  94710.0 115757.5 95415.0 115822.5 ;
      RECT  95767.5 115307.5 95832.5 115822.5 ;
      RECT  95577.5 114777.5 95642.5 114912.5 ;
      RECT  95767.5 114777.5 95832.5 114912.5 ;
      RECT  95767.5 114777.5 95832.5 114912.5 ;
      RECT  95577.5 114777.5 95642.5 114912.5 ;
      RECT  95577.5 115307.5 95642.5 115442.5 ;
      RECT  95767.5 115307.5 95832.5 115442.5 ;
      RECT  95767.5 115307.5 95832.5 115442.5 ;
      RECT  95577.5 115307.5 95642.5 115442.5 ;
      RECT  95767.5 115307.5 95832.5 115442.5 ;
      RECT  95957.5 115307.5 96022.5 115442.5 ;
      RECT  95957.5 115307.5 96022.5 115442.5 ;
      RECT  95767.5 115307.5 95832.5 115442.5 ;
      RECT  95747.5 115072.5 95612.5 115137.5 ;
      RECT  95767.5 115620.0 95832.5 115755.0 ;
      RECT  95577.5 114777.5 95642.5 114912.5 ;
      RECT  95767.5 114777.5 95832.5 114912.5 ;
      RECT  95577.5 115307.5 95642.5 115442.5 ;
      RECT  95957.5 115307.5 96022.5 115442.5 ;
      RECT  95415.0 115072.5 96120.0 115137.5 ;
      RECT  95415.0 115757.5 96120.0 115822.5 ;
      RECT  96472.5 115307.5 96537.5 115822.5 ;
      RECT  96282.5 114777.5 96347.5 114912.5 ;
      RECT  96472.5 114777.5 96537.5 114912.5 ;
      RECT  96472.5 114777.5 96537.5 114912.5 ;
      RECT  96282.5 114777.5 96347.5 114912.5 ;
      RECT  96282.5 115307.5 96347.5 115442.5 ;
      RECT  96472.5 115307.5 96537.5 115442.5 ;
      RECT  96472.5 115307.5 96537.5 115442.5 ;
      RECT  96282.5 115307.5 96347.5 115442.5 ;
      RECT  96472.5 115307.5 96537.5 115442.5 ;
      RECT  96662.5 115307.5 96727.5 115442.5 ;
      RECT  96662.5 115307.5 96727.5 115442.5 ;
      RECT  96472.5 115307.5 96537.5 115442.5 ;
      RECT  96452.5 115072.5 96317.5 115137.5 ;
      RECT  96472.5 115620.0 96537.5 115755.0 ;
      RECT  96282.5 114777.5 96347.5 114912.5 ;
      RECT  96472.5 114777.5 96537.5 114912.5 ;
      RECT  96282.5 115307.5 96347.5 115442.5 ;
      RECT  96662.5 115307.5 96727.5 115442.5 ;
      RECT  96120.0 115072.5 96825.0 115137.5 ;
      RECT  96120.0 115757.5 96825.0 115822.5 ;
      RECT  97177.5 115307.5 97242.5 115822.5 ;
      RECT  96987.5 114777.5 97052.5 114912.5 ;
      RECT  97177.5 114777.5 97242.5 114912.5 ;
      RECT  97177.5 114777.5 97242.5 114912.5 ;
      RECT  96987.5 114777.5 97052.5 114912.5 ;
      RECT  96987.5 115307.5 97052.5 115442.5 ;
      RECT  97177.5 115307.5 97242.5 115442.5 ;
      RECT  97177.5 115307.5 97242.5 115442.5 ;
      RECT  96987.5 115307.5 97052.5 115442.5 ;
      RECT  97177.5 115307.5 97242.5 115442.5 ;
      RECT  97367.5 115307.5 97432.5 115442.5 ;
      RECT  97367.5 115307.5 97432.5 115442.5 ;
      RECT  97177.5 115307.5 97242.5 115442.5 ;
      RECT  97157.5 115072.5 97022.5 115137.5 ;
      RECT  97177.5 115620.0 97242.5 115755.0 ;
      RECT  96987.5 114777.5 97052.5 114912.5 ;
      RECT  97177.5 114777.5 97242.5 114912.5 ;
      RECT  96987.5 115307.5 97052.5 115442.5 ;
      RECT  97367.5 115307.5 97432.5 115442.5 ;
      RECT  96825.0 115072.5 97530.0 115137.5 ;
      RECT  96825.0 115757.5 97530.0 115822.5 ;
      RECT  97882.5 115307.5 97947.5 115822.5 ;
      RECT  97692.5 114777.5 97757.5 114912.5 ;
      RECT  97882.5 114777.5 97947.5 114912.5 ;
      RECT  97882.5 114777.5 97947.5 114912.5 ;
      RECT  97692.5 114777.5 97757.5 114912.5 ;
      RECT  97692.5 115307.5 97757.5 115442.5 ;
      RECT  97882.5 115307.5 97947.5 115442.5 ;
      RECT  97882.5 115307.5 97947.5 115442.5 ;
      RECT  97692.5 115307.5 97757.5 115442.5 ;
      RECT  97882.5 115307.5 97947.5 115442.5 ;
      RECT  98072.5 115307.5 98137.5 115442.5 ;
      RECT  98072.5 115307.5 98137.5 115442.5 ;
      RECT  97882.5 115307.5 97947.5 115442.5 ;
      RECT  97862.5 115072.5 97727.5 115137.5 ;
      RECT  97882.5 115620.0 97947.5 115755.0 ;
      RECT  97692.5 114777.5 97757.5 114912.5 ;
      RECT  97882.5 114777.5 97947.5 114912.5 ;
      RECT  97692.5 115307.5 97757.5 115442.5 ;
      RECT  98072.5 115307.5 98137.5 115442.5 ;
      RECT  97530.0 115072.5 98235.0 115137.5 ;
      RECT  97530.0 115757.5 98235.0 115822.5 ;
      RECT  98587.5 115307.5 98652.5 115822.5 ;
      RECT  98397.5 114777.5 98462.5 114912.5 ;
      RECT  98587.5 114777.5 98652.5 114912.5 ;
      RECT  98587.5 114777.5 98652.5 114912.5 ;
      RECT  98397.5 114777.5 98462.5 114912.5 ;
      RECT  98397.5 115307.5 98462.5 115442.5 ;
      RECT  98587.5 115307.5 98652.5 115442.5 ;
      RECT  98587.5 115307.5 98652.5 115442.5 ;
      RECT  98397.5 115307.5 98462.5 115442.5 ;
      RECT  98587.5 115307.5 98652.5 115442.5 ;
      RECT  98777.5 115307.5 98842.5 115442.5 ;
      RECT  98777.5 115307.5 98842.5 115442.5 ;
      RECT  98587.5 115307.5 98652.5 115442.5 ;
      RECT  98567.5 115072.5 98432.5 115137.5 ;
      RECT  98587.5 115620.0 98652.5 115755.0 ;
      RECT  98397.5 114777.5 98462.5 114912.5 ;
      RECT  98587.5 114777.5 98652.5 114912.5 ;
      RECT  98397.5 115307.5 98462.5 115442.5 ;
      RECT  98777.5 115307.5 98842.5 115442.5 ;
      RECT  98235.0 115072.5 98940.0 115137.5 ;
      RECT  98235.0 115757.5 98940.0 115822.5 ;
      RECT  99292.5 115307.5 99357.5 115822.5 ;
      RECT  99102.5 114777.5 99167.5 114912.5 ;
      RECT  99292.5 114777.5 99357.5 114912.5 ;
      RECT  99292.5 114777.5 99357.5 114912.5 ;
      RECT  99102.5 114777.5 99167.5 114912.5 ;
      RECT  99102.5 115307.5 99167.5 115442.5 ;
      RECT  99292.5 115307.5 99357.5 115442.5 ;
      RECT  99292.5 115307.5 99357.5 115442.5 ;
      RECT  99102.5 115307.5 99167.5 115442.5 ;
      RECT  99292.5 115307.5 99357.5 115442.5 ;
      RECT  99482.5 115307.5 99547.5 115442.5 ;
      RECT  99482.5 115307.5 99547.5 115442.5 ;
      RECT  99292.5 115307.5 99357.5 115442.5 ;
      RECT  99272.5 115072.5 99137.5 115137.5 ;
      RECT  99292.5 115620.0 99357.5 115755.0 ;
      RECT  99102.5 114777.5 99167.5 114912.5 ;
      RECT  99292.5 114777.5 99357.5 114912.5 ;
      RECT  99102.5 115307.5 99167.5 115442.5 ;
      RECT  99482.5 115307.5 99547.5 115442.5 ;
      RECT  98940.0 115072.5 99645.0 115137.5 ;
      RECT  98940.0 115757.5 99645.0 115822.5 ;
      RECT  99997.5 115307.5 100062.5 115822.5 ;
      RECT  99807.5 114777.5 99872.5 114912.5 ;
      RECT  99997.5 114777.5 100062.5 114912.5 ;
      RECT  99997.5 114777.5 100062.5 114912.5 ;
      RECT  99807.5 114777.5 99872.5 114912.5 ;
      RECT  99807.5 115307.5 99872.5 115442.5 ;
      RECT  99997.5 115307.5 100062.5 115442.5 ;
      RECT  99997.5 115307.5 100062.5 115442.5 ;
      RECT  99807.5 115307.5 99872.5 115442.5 ;
      RECT  99997.5 115307.5 100062.5 115442.5 ;
      RECT  100187.5 115307.5 100252.5 115442.5 ;
      RECT  100187.5 115307.5 100252.5 115442.5 ;
      RECT  99997.5 115307.5 100062.5 115442.5 ;
      RECT  99977.5 115072.5 99842.5 115137.5 ;
      RECT  99997.5 115620.0 100062.5 115755.0 ;
      RECT  99807.5 114777.5 99872.5 114912.5 ;
      RECT  99997.5 114777.5 100062.5 114912.5 ;
      RECT  99807.5 115307.5 99872.5 115442.5 ;
      RECT  100187.5 115307.5 100252.5 115442.5 ;
      RECT  99645.0 115072.5 100350.0 115137.5 ;
      RECT  99645.0 115757.5 100350.0 115822.5 ;
      RECT  100702.5 115307.5 100767.5 115822.5 ;
      RECT  100512.5 114777.5 100577.5 114912.5 ;
      RECT  100702.5 114777.5 100767.5 114912.5 ;
      RECT  100702.5 114777.5 100767.5 114912.5 ;
      RECT  100512.5 114777.5 100577.5 114912.5 ;
      RECT  100512.5 115307.5 100577.5 115442.5 ;
      RECT  100702.5 115307.5 100767.5 115442.5 ;
      RECT  100702.5 115307.5 100767.5 115442.5 ;
      RECT  100512.5 115307.5 100577.5 115442.5 ;
      RECT  100702.5 115307.5 100767.5 115442.5 ;
      RECT  100892.5 115307.5 100957.5 115442.5 ;
      RECT  100892.5 115307.5 100957.5 115442.5 ;
      RECT  100702.5 115307.5 100767.5 115442.5 ;
      RECT  100682.5 115072.5 100547.5 115137.5 ;
      RECT  100702.5 115620.0 100767.5 115755.0 ;
      RECT  100512.5 114777.5 100577.5 114912.5 ;
      RECT  100702.5 114777.5 100767.5 114912.5 ;
      RECT  100512.5 115307.5 100577.5 115442.5 ;
      RECT  100892.5 115307.5 100957.5 115442.5 ;
      RECT  100350.0 115072.5 101055.0 115137.5 ;
      RECT  100350.0 115757.5 101055.0 115822.5 ;
      RECT  101407.5 115307.5 101472.5 115822.5 ;
      RECT  101217.5 114777.5 101282.5 114912.5 ;
      RECT  101407.5 114777.5 101472.5 114912.5 ;
      RECT  101407.5 114777.5 101472.5 114912.5 ;
      RECT  101217.5 114777.5 101282.5 114912.5 ;
      RECT  101217.5 115307.5 101282.5 115442.5 ;
      RECT  101407.5 115307.5 101472.5 115442.5 ;
      RECT  101407.5 115307.5 101472.5 115442.5 ;
      RECT  101217.5 115307.5 101282.5 115442.5 ;
      RECT  101407.5 115307.5 101472.5 115442.5 ;
      RECT  101597.5 115307.5 101662.5 115442.5 ;
      RECT  101597.5 115307.5 101662.5 115442.5 ;
      RECT  101407.5 115307.5 101472.5 115442.5 ;
      RECT  101387.5 115072.5 101252.5 115137.5 ;
      RECT  101407.5 115620.0 101472.5 115755.0 ;
      RECT  101217.5 114777.5 101282.5 114912.5 ;
      RECT  101407.5 114777.5 101472.5 114912.5 ;
      RECT  101217.5 115307.5 101282.5 115442.5 ;
      RECT  101597.5 115307.5 101662.5 115442.5 ;
      RECT  101055.0 115072.5 101760.0 115137.5 ;
      RECT  101055.0 115757.5 101760.0 115822.5 ;
      RECT  102112.5 115307.5 102177.5 115822.5 ;
      RECT  101922.5 114777.5 101987.5 114912.5 ;
      RECT  102112.5 114777.5 102177.5 114912.5 ;
      RECT  102112.5 114777.5 102177.5 114912.5 ;
      RECT  101922.5 114777.5 101987.5 114912.5 ;
      RECT  101922.5 115307.5 101987.5 115442.5 ;
      RECT  102112.5 115307.5 102177.5 115442.5 ;
      RECT  102112.5 115307.5 102177.5 115442.5 ;
      RECT  101922.5 115307.5 101987.5 115442.5 ;
      RECT  102112.5 115307.5 102177.5 115442.5 ;
      RECT  102302.5 115307.5 102367.5 115442.5 ;
      RECT  102302.5 115307.5 102367.5 115442.5 ;
      RECT  102112.5 115307.5 102177.5 115442.5 ;
      RECT  102092.5 115072.5 101957.5 115137.5 ;
      RECT  102112.5 115620.0 102177.5 115755.0 ;
      RECT  101922.5 114777.5 101987.5 114912.5 ;
      RECT  102112.5 114777.5 102177.5 114912.5 ;
      RECT  101922.5 115307.5 101987.5 115442.5 ;
      RECT  102302.5 115307.5 102367.5 115442.5 ;
      RECT  101760.0 115072.5 102465.0 115137.5 ;
      RECT  101760.0 115757.5 102465.0 115822.5 ;
      RECT  102817.5 115307.5 102882.5 115822.5 ;
      RECT  102627.5 114777.5 102692.5 114912.5 ;
      RECT  102817.5 114777.5 102882.5 114912.5 ;
      RECT  102817.5 114777.5 102882.5 114912.5 ;
      RECT  102627.5 114777.5 102692.5 114912.5 ;
      RECT  102627.5 115307.5 102692.5 115442.5 ;
      RECT  102817.5 115307.5 102882.5 115442.5 ;
      RECT  102817.5 115307.5 102882.5 115442.5 ;
      RECT  102627.5 115307.5 102692.5 115442.5 ;
      RECT  102817.5 115307.5 102882.5 115442.5 ;
      RECT  103007.5 115307.5 103072.5 115442.5 ;
      RECT  103007.5 115307.5 103072.5 115442.5 ;
      RECT  102817.5 115307.5 102882.5 115442.5 ;
      RECT  102797.5 115072.5 102662.5 115137.5 ;
      RECT  102817.5 115620.0 102882.5 115755.0 ;
      RECT  102627.5 114777.5 102692.5 114912.5 ;
      RECT  102817.5 114777.5 102882.5 114912.5 ;
      RECT  102627.5 115307.5 102692.5 115442.5 ;
      RECT  103007.5 115307.5 103072.5 115442.5 ;
      RECT  102465.0 115072.5 103170.0 115137.5 ;
      RECT  102465.0 115757.5 103170.0 115822.5 ;
      RECT  103522.5 115307.5 103587.5 115822.5 ;
      RECT  103332.5 114777.5 103397.5 114912.5 ;
      RECT  103522.5 114777.5 103587.5 114912.5 ;
      RECT  103522.5 114777.5 103587.5 114912.5 ;
      RECT  103332.5 114777.5 103397.5 114912.5 ;
      RECT  103332.5 115307.5 103397.5 115442.5 ;
      RECT  103522.5 115307.5 103587.5 115442.5 ;
      RECT  103522.5 115307.5 103587.5 115442.5 ;
      RECT  103332.5 115307.5 103397.5 115442.5 ;
      RECT  103522.5 115307.5 103587.5 115442.5 ;
      RECT  103712.5 115307.5 103777.5 115442.5 ;
      RECT  103712.5 115307.5 103777.5 115442.5 ;
      RECT  103522.5 115307.5 103587.5 115442.5 ;
      RECT  103502.5 115072.5 103367.5 115137.5 ;
      RECT  103522.5 115620.0 103587.5 115755.0 ;
      RECT  103332.5 114777.5 103397.5 114912.5 ;
      RECT  103522.5 114777.5 103587.5 114912.5 ;
      RECT  103332.5 115307.5 103397.5 115442.5 ;
      RECT  103712.5 115307.5 103777.5 115442.5 ;
      RECT  103170.0 115072.5 103875.0 115137.5 ;
      RECT  103170.0 115757.5 103875.0 115822.5 ;
      RECT  104227.5 115307.5 104292.5 115822.5 ;
      RECT  104037.5 114777.5 104102.5 114912.5 ;
      RECT  104227.5 114777.5 104292.5 114912.5 ;
      RECT  104227.5 114777.5 104292.5 114912.5 ;
      RECT  104037.5 114777.5 104102.5 114912.5 ;
      RECT  104037.5 115307.5 104102.5 115442.5 ;
      RECT  104227.5 115307.5 104292.5 115442.5 ;
      RECT  104227.5 115307.5 104292.5 115442.5 ;
      RECT  104037.5 115307.5 104102.5 115442.5 ;
      RECT  104227.5 115307.5 104292.5 115442.5 ;
      RECT  104417.5 115307.5 104482.5 115442.5 ;
      RECT  104417.5 115307.5 104482.5 115442.5 ;
      RECT  104227.5 115307.5 104292.5 115442.5 ;
      RECT  104207.5 115072.5 104072.5 115137.5 ;
      RECT  104227.5 115620.0 104292.5 115755.0 ;
      RECT  104037.5 114777.5 104102.5 114912.5 ;
      RECT  104227.5 114777.5 104292.5 114912.5 ;
      RECT  104037.5 115307.5 104102.5 115442.5 ;
      RECT  104417.5 115307.5 104482.5 115442.5 ;
      RECT  103875.0 115072.5 104580.0 115137.5 ;
      RECT  103875.0 115757.5 104580.0 115822.5 ;
      RECT  104932.5 115307.5 104997.5 115822.5 ;
      RECT  104742.5 114777.5 104807.5 114912.5 ;
      RECT  104932.5 114777.5 104997.5 114912.5 ;
      RECT  104932.5 114777.5 104997.5 114912.5 ;
      RECT  104742.5 114777.5 104807.5 114912.5 ;
      RECT  104742.5 115307.5 104807.5 115442.5 ;
      RECT  104932.5 115307.5 104997.5 115442.5 ;
      RECT  104932.5 115307.5 104997.5 115442.5 ;
      RECT  104742.5 115307.5 104807.5 115442.5 ;
      RECT  104932.5 115307.5 104997.5 115442.5 ;
      RECT  105122.5 115307.5 105187.5 115442.5 ;
      RECT  105122.5 115307.5 105187.5 115442.5 ;
      RECT  104932.5 115307.5 104997.5 115442.5 ;
      RECT  104912.5 115072.5 104777.5 115137.5 ;
      RECT  104932.5 115620.0 104997.5 115755.0 ;
      RECT  104742.5 114777.5 104807.5 114912.5 ;
      RECT  104932.5 114777.5 104997.5 114912.5 ;
      RECT  104742.5 115307.5 104807.5 115442.5 ;
      RECT  105122.5 115307.5 105187.5 115442.5 ;
      RECT  104580.0 115072.5 105285.0 115137.5 ;
      RECT  104580.0 115757.5 105285.0 115822.5 ;
      RECT  105637.5 115307.5 105702.5 115822.5 ;
      RECT  105447.5 114777.5 105512.5 114912.5 ;
      RECT  105637.5 114777.5 105702.5 114912.5 ;
      RECT  105637.5 114777.5 105702.5 114912.5 ;
      RECT  105447.5 114777.5 105512.5 114912.5 ;
      RECT  105447.5 115307.5 105512.5 115442.5 ;
      RECT  105637.5 115307.5 105702.5 115442.5 ;
      RECT  105637.5 115307.5 105702.5 115442.5 ;
      RECT  105447.5 115307.5 105512.5 115442.5 ;
      RECT  105637.5 115307.5 105702.5 115442.5 ;
      RECT  105827.5 115307.5 105892.5 115442.5 ;
      RECT  105827.5 115307.5 105892.5 115442.5 ;
      RECT  105637.5 115307.5 105702.5 115442.5 ;
      RECT  105617.5 115072.5 105482.5 115137.5 ;
      RECT  105637.5 115620.0 105702.5 115755.0 ;
      RECT  105447.5 114777.5 105512.5 114912.5 ;
      RECT  105637.5 114777.5 105702.5 114912.5 ;
      RECT  105447.5 115307.5 105512.5 115442.5 ;
      RECT  105827.5 115307.5 105892.5 115442.5 ;
      RECT  105285.0 115072.5 105990.0 115137.5 ;
      RECT  105285.0 115757.5 105990.0 115822.5 ;
      RECT  15750.0 115072.5 105990.0 115137.5 ;
      RECT  15750.0 115757.5 105990.0 115822.5 ;
      RECT  15900.0 25450.0 18085.0 25520.0 ;
      RECT  16235.0 25310.0 18420.0 25380.0 ;
      RECT  18720.0 25450.0 20905.0 25520.0 ;
      RECT  19055.0 25310.0 21240.0 25380.0 ;
      RECT  21540.0 25450.0 23725.0 25520.0 ;
      RECT  21875.0 25310.0 24060.0 25380.0 ;
      RECT  24360.0 25450.0 26545.0 25520.0 ;
      RECT  24695.0 25310.0 26880.0 25380.0 ;
      RECT  27180.0 25450.0 29365.0 25520.0 ;
      RECT  27515.0 25310.0 29700.0 25380.0 ;
      RECT  30000.0 25450.0 32185.0 25520.0 ;
      RECT  30335.0 25310.0 32520.0 25380.0 ;
      RECT  32820.0 25450.0 35005.0 25520.0 ;
      RECT  33155.0 25310.0 35340.0 25380.0 ;
      RECT  35640.0 25450.0 37825.0 25520.0 ;
      RECT  35975.0 25310.0 38160.0 25380.0 ;
      RECT  38460.0 25450.0 40645.0 25520.0 ;
      RECT  38795.0 25310.0 40980.0 25380.0 ;
      RECT  41280.0 25450.0 43465.0 25520.0 ;
      RECT  41615.0 25310.0 43800.0 25380.0 ;
      RECT  44100.0 25450.0 46285.0 25520.0 ;
      RECT  44435.0 25310.0 46620.0 25380.0 ;
      RECT  46920.0 25450.0 49105.0 25520.0 ;
      RECT  47255.0 25310.0 49440.0 25380.0 ;
      RECT  49740.0 25450.0 51925.0 25520.0 ;
      RECT  50075.0 25310.0 52260.0 25380.0 ;
      RECT  52560.0 25450.0 54745.0 25520.0 ;
      RECT  52895.0 25310.0 55080.0 25380.0 ;
      RECT  55380.0 25450.0 57565.0 25520.0 ;
      RECT  55715.0 25310.0 57900.0 25380.0 ;
      RECT  58200.0 25450.0 60385.0 25520.0 ;
      RECT  58535.0 25310.0 60720.0 25380.0 ;
      RECT  61020.0 25450.0 63205.0 25520.0 ;
      RECT  61355.0 25310.0 63540.0 25380.0 ;
      RECT  63840.0 25450.0 66025.0 25520.0 ;
      RECT  64175.0 25310.0 66360.0 25380.0 ;
      RECT  66660.0 25450.0 68845.0 25520.0 ;
      RECT  66995.0 25310.0 69180.0 25380.0 ;
      RECT  69480.0 25450.0 71665.0 25520.0 ;
      RECT  69815.0 25310.0 72000.0 25380.0 ;
      RECT  72300.0 25450.0 74485.0 25520.0 ;
      RECT  72635.0 25310.0 74820.0 25380.0 ;
      RECT  75120.0 25450.0 77305.0 25520.0 ;
      RECT  75455.0 25310.0 77640.0 25380.0 ;
      RECT  77940.0 25450.0 80125.0 25520.0 ;
      RECT  78275.0 25310.0 80460.0 25380.0 ;
      RECT  80760.0 25450.0 82945.0 25520.0 ;
      RECT  81095.0 25310.0 83280.0 25380.0 ;
      RECT  83580.0 25450.0 85765.0 25520.0 ;
      RECT  83915.0 25310.0 86100.0 25380.0 ;
      RECT  86400.0 25450.0 88585.0 25520.0 ;
      RECT  86735.0 25310.0 88920.0 25380.0 ;
      RECT  89220.0 25450.0 91405.0 25520.0 ;
      RECT  89555.0 25310.0 91740.0 25380.0 ;
      RECT  92040.0 25450.0 94225.0 25520.0 ;
      RECT  92375.0 25310.0 94560.0 25380.0 ;
      RECT  94860.0 25450.0 97045.0 25520.0 ;
      RECT  95195.0 25310.0 97380.0 25380.0 ;
      RECT  97680.0 25450.0 99865.0 25520.0 ;
      RECT  98015.0 25310.0 100200.0 25380.0 ;
      RECT  100500.0 25450.0 102685.0 25520.0 ;
      RECT  100835.0 25310.0 103020.0 25380.0 ;
      RECT  103320.0 25450.0 105505.0 25520.0 ;
      RECT  103655.0 25310.0 105840.0 25380.0 ;
      RECT  16165.0 27807.5 16230.0 27872.5 ;
      RECT  15900.0 27807.5 16197.5 27872.5 ;
      RECT  16165.0 27425.0 16230.0 27840.0 ;
      RECT  15975.0 26257.5 16040.0 26322.5 ;
      RECT  16007.5 26257.5 16270.0 26322.5 ;
      RECT  15975.0 26290.0 16040.0 26565.0 ;
      RECT  15975.0 26497.5 16040.0 26632.5 ;
      RECT  16165.0 26497.5 16230.0 26632.5 ;
      RECT  16165.0 26497.5 16230.0 26632.5 ;
      RECT  15975.0 26497.5 16040.0 26632.5 ;
      RECT  15975.0 27357.5 16040.0 27492.5 ;
      RECT  16165.0 27357.5 16230.0 27492.5 ;
      RECT  16165.0 27357.5 16230.0 27492.5 ;
      RECT  15975.0 27357.5 16040.0 27492.5 ;
      RECT  15902.5 27772.5 15967.5 27907.5 ;
      RECT  16237.5 26222.5 16302.5 26357.5 ;
      RECT  15975.0 27357.5 16040.0 27492.5 ;
      RECT  16165.0 26497.5 16230.0 26632.5 ;
      RECT  16422.5 26397.5 16487.5 26532.5 ;
      RECT  16422.5 26397.5 16487.5 26532.5 ;
      RECT  16870.0 27807.5 16935.0 27872.5 ;
      RECT  16605.0 27807.5 16902.5 27872.5 ;
      RECT  16870.0 27425.0 16935.0 27840.0 ;
      RECT  16680.0 26257.5 16745.0 26322.5 ;
      RECT  16712.5 26257.5 16975.0 26322.5 ;
      RECT  16680.0 26290.0 16745.0 26565.0 ;
      RECT  16680.0 26497.5 16745.0 26632.5 ;
      RECT  16870.0 26497.5 16935.0 26632.5 ;
      RECT  16870.0 26497.5 16935.0 26632.5 ;
      RECT  16680.0 26497.5 16745.0 26632.5 ;
      RECT  16680.0 27357.5 16745.0 27492.5 ;
      RECT  16870.0 27357.5 16935.0 27492.5 ;
      RECT  16870.0 27357.5 16935.0 27492.5 ;
      RECT  16680.0 27357.5 16745.0 27492.5 ;
      RECT  16607.5 27772.5 16672.5 27907.5 ;
      RECT  16942.5 26222.5 17007.5 26357.5 ;
      RECT  16680.0 27357.5 16745.0 27492.5 ;
      RECT  16870.0 26497.5 16935.0 26632.5 ;
      RECT  17127.5 26397.5 17192.5 26532.5 ;
      RECT  17127.5 26397.5 17192.5 26532.5 ;
      RECT  17575.0 27807.5 17640.0 27872.5 ;
      RECT  17310.0 27807.5 17607.5 27872.5 ;
      RECT  17575.0 27425.0 17640.0 27840.0 ;
      RECT  17385.0 26257.5 17450.0 26322.5 ;
      RECT  17417.5 26257.5 17680.0 26322.5 ;
      RECT  17385.0 26290.0 17450.0 26565.0 ;
      RECT  17385.0 26497.5 17450.0 26632.5 ;
      RECT  17575.0 26497.5 17640.0 26632.5 ;
      RECT  17575.0 26497.5 17640.0 26632.5 ;
      RECT  17385.0 26497.5 17450.0 26632.5 ;
      RECT  17385.0 27357.5 17450.0 27492.5 ;
      RECT  17575.0 27357.5 17640.0 27492.5 ;
      RECT  17575.0 27357.5 17640.0 27492.5 ;
      RECT  17385.0 27357.5 17450.0 27492.5 ;
      RECT  17312.5 27772.5 17377.5 27907.5 ;
      RECT  17647.5 26222.5 17712.5 26357.5 ;
      RECT  17385.0 27357.5 17450.0 27492.5 ;
      RECT  17575.0 26497.5 17640.0 26632.5 ;
      RECT  17832.5 26397.5 17897.5 26532.5 ;
      RECT  17832.5 26397.5 17897.5 26532.5 ;
      RECT  18280.0 27807.5 18345.0 27872.5 ;
      RECT  18015.0 27807.5 18312.5 27872.5 ;
      RECT  18280.0 27425.0 18345.0 27840.0 ;
      RECT  18090.0 26257.5 18155.0 26322.5 ;
      RECT  18122.5 26257.5 18385.0 26322.5 ;
      RECT  18090.0 26290.0 18155.0 26565.0 ;
      RECT  18090.0 26497.5 18155.0 26632.5 ;
      RECT  18280.0 26497.5 18345.0 26632.5 ;
      RECT  18280.0 26497.5 18345.0 26632.5 ;
      RECT  18090.0 26497.5 18155.0 26632.5 ;
      RECT  18090.0 27357.5 18155.0 27492.5 ;
      RECT  18280.0 27357.5 18345.0 27492.5 ;
      RECT  18280.0 27357.5 18345.0 27492.5 ;
      RECT  18090.0 27357.5 18155.0 27492.5 ;
      RECT  18017.5 27772.5 18082.5 27907.5 ;
      RECT  18352.5 26222.5 18417.5 26357.5 ;
      RECT  18090.0 27357.5 18155.0 27492.5 ;
      RECT  18280.0 26497.5 18345.0 26632.5 ;
      RECT  18537.5 26397.5 18602.5 26532.5 ;
      RECT  18537.5 26397.5 18602.5 26532.5 ;
      RECT  18985.0 27807.5 19050.0 27872.5 ;
      RECT  18720.0 27807.5 19017.5 27872.5 ;
      RECT  18985.0 27425.0 19050.0 27840.0 ;
      RECT  18795.0 26257.5 18860.0 26322.5 ;
      RECT  18827.5 26257.5 19090.0 26322.5 ;
      RECT  18795.0 26290.0 18860.0 26565.0 ;
      RECT  18795.0 26497.5 18860.0 26632.5 ;
      RECT  18985.0 26497.5 19050.0 26632.5 ;
      RECT  18985.0 26497.5 19050.0 26632.5 ;
      RECT  18795.0 26497.5 18860.0 26632.5 ;
      RECT  18795.0 27357.5 18860.0 27492.5 ;
      RECT  18985.0 27357.5 19050.0 27492.5 ;
      RECT  18985.0 27357.5 19050.0 27492.5 ;
      RECT  18795.0 27357.5 18860.0 27492.5 ;
      RECT  18722.5 27772.5 18787.5 27907.5 ;
      RECT  19057.5 26222.5 19122.5 26357.5 ;
      RECT  18795.0 27357.5 18860.0 27492.5 ;
      RECT  18985.0 26497.5 19050.0 26632.5 ;
      RECT  19242.5 26397.5 19307.5 26532.5 ;
      RECT  19242.5 26397.5 19307.5 26532.5 ;
      RECT  19690.0 27807.5 19755.0 27872.5 ;
      RECT  19425.0 27807.5 19722.5 27872.5 ;
      RECT  19690.0 27425.0 19755.0 27840.0 ;
      RECT  19500.0 26257.5 19565.0 26322.5 ;
      RECT  19532.5 26257.5 19795.0 26322.5 ;
      RECT  19500.0 26290.0 19565.0 26565.0 ;
      RECT  19500.0 26497.5 19565.0 26632.5 ;
      RECT  19690.0 26497.5 19755.0 26632.5 ;
      RECT  19690.0 26497.5 19755.0 26632.5 ;
      RECT  19500.0 26497.5 19565.0 26632.5 ;
      RECT  19500.0 27357.5 19565.0 27492.5 ;
      RECT  19690.0 27357.5 19755.0 27492.5 ;
      RECT  19690.0 27357.5 19755.0 27492.5 ;
      RECT  19500.0 27357.5 19565.0 27492.5 ;
      RECT  19427.5 27772.5 19492.5 27907.5 ;
      RECT  19762.5 26222.5 19827.5 26357.5 ;
      RECT  19500.0 27357.5 19565.0 27492.5 ;
      RECT  19690.0 26497.5 19755.0 26632.5 ;
      RECT  19947.5 26397.5 20012.5 26532.5 ;
      RECT  19947.5 26397.5 20012.5 26532.5 ;
      RECT  20395.0 27807.5 20460.0 27872.5 ;
      RECT  20130.0 27807.5 20427.5 27872.5 ;
      RECT  20395.0 27425.0 20460.0 27840.0 ;
      RECT  20205.0 26257.5 20270.0 26322.5 ;
      RECT  20237.5 26257.5 20500.0 26322.5 ;
      RECT  20205.0 26290.0 20270.0 26565.0 ;
      RECT  20205.0 26497.5 20270.0 26632.5 ;
      RECT  20395.0 26497.5 20460.0 26632.5 ;
      RECT  20395.0 26497.5 20460.0 26632.5 ;
      RECT  20205.0 26497.5 20270.0 26632.5 ;
      RECT  20205.0 27357.5 20270.0 27492.5 ;
      RECT  20395.0 27357.5 20460.0 27492.5 ;
      RECT  20395.0 27357.5 20460.0 27492.5 ;
      RECT  20205.0 27357.5 20270.0 27492.5 ;
      RECT  20132.5 27772.5 20197.5 27907.5 ;
      RECT  20467.5 26222.5 20532.5 26357.5 ;
      RECT  20205.0 27357.5 20270.0 27492.5 ;
      RECT  20395.0 26497.5 20460.0 26632.5 ;
      RECT  20652.5 26397.5 20717.5 26532.5 ;
      RECT  20652.5 26397.5 20717.5 26532.5 ;
      RECT  21100.0 27807.5 21165.0 27872.5 ;
      RECT  20835.0 27807.5 21132.5 27872.5 ;
      RECT  21100.0 27425.0 21165.0 27840.0 ;
      RECT  20910.0 26257.5 20975.0 26322.5 ;
      RECT  20942.5 26257.5 21205.0 26322.5 ;
      RECT  20910.0 26290.0 20975.0 26565.0 ;
      RECT  20910.0 26497.5 20975.0 26632.5 ;
      RECT  21100.0 26497.5 21165.0 26632.5 ;
      RECT  21100.0 26497.5 21165.0 26632.5 ;
      RECT  20910.0 26497.5 20975.0 26632.5 ;
      RECT  20910.0 27357.5 20975.0 27492.5 ;
      RECT  21100.0 27357.5 21165.0 27492.5 ;
      RECT  21100.0 27357.5 21165.0 27492.5 ;
      RECT  20910.0 27357.5 20975.0 27492.5 ;
      RECT  20837.5 27772.5 20902.5 27907.5 ;
      RECT  21172.5 26222.5 21237.5 26357.5 ;
      RECT  20910.0 27357.5 20975.0 27492.5 ;
      RECT  21100.0 26497.5 21165.0 26632.5 ;
      RECT  21357.5 26397.5 21422.5 26532.5 ;
      RECT  21357.5 26397.5 21422.5 26532.5 ;
      RECT  21805.0 27807.5 21870.0 27872.5 ;
      RECT  21540.0 27807.5 21837.5 27872.5 ;
      RECT  21805.0 27425.0 21870.0 27840.0 ;
      RECT  21615.0 26257.5 21680.0 26322.5 ;
      RECT  21647.5 26257.5 21910.0 26322.5 ;
      RECT  21615.0 26290.0 21680.0 26565.0 ;
      RECT  21615.0 26497.5 21680.0 26632.5 ;
      RECT  21805.0 26497.5 21870.0 26632.5 ;
      RECT  21805.0 26497.5 21870.0 26632.5 ;
      RECT  21615.0 26497.5 21680.0 26632.5 ;
      RECT  21615.0 27357.5 21680.0 27492.5 ;
      RECT  21805.0 27357.5 21870.0 27492.5 ;
      RECT  21805.0 27357.5 21870.0 27492.5 ;
      RECT  21615.0 27357.5 21680.0 27492.5 ;
      RECT  21542.5 27772.5 21607.5 27907.5 ;
      RECT  21877.5 26222.5 21942.5 26357.5 ;
      RECT  21615.0 27357.5 21680.0 27492.5 ;
      RECT  21805.0 26497.5 21870.0 26632.5 ;
      RECT  22062.5 26397.5 22127.5 26532.5 ;
      RECT  22062.5 26397.5 22127.5 26532.5 ;
      RECT  22510.0 27807.5 22575.0 27872.5 ;
      RECT  22245.0 27807.5 22542.5 27872.5 ;
      RECT  22510.0 27425.0 22575.0 27840.0 ;
      RECT  22320.0 26257.5 22385.0 26322.5 ;
      RECT  22352.5 26257.5 22615.0 26322.5 ;
      RECT  22320.0 26290.0 22385.0 26565.0 ;
      RECT  22320.0 26497.5 22385.0 26632.5 ;
      RECT  22510.0 26497.5 22575.0 26632.5 ;
      RECT  22510.0 26497.5 22575.0 26632.5 ;
      RECT  22320.0 26497.5 22385.0 26632.5 ;
      RECT  22320.0 27357.5 22385.0 27492.5 ;
      RECT  22510.0 27357.5 22575.0 27492.5 ;
      RECT  22510.0 27357.5 22575.0 27492.5 ;
      RECT  22320.0 27357.5 22385.0 27492.5 ;
      RECT  22247.5 27772.5 22312.5 27907.5 ;
      RECT  22582.5 26222.5 22647.5 26357.5 ;
      RECT  22320.0 27357.5 22385.0 27492.5 ;
      RECT  22510.0 26497.5 22575.0 26632.5 ;
      RECT  22767.5 26397.5 22832.5 26532.5 ;
      RECT  22767.5 26397.5 22832.5 26532.5 ;
      RECT  23215.0 27807.5 23280.0 27872.5 ;
      RECT  22950.0 27807.5 23247.5 27872.5 ;
      RECT  23215.0 27425.0 23280.0 27840.0 ;
      RECT  23025.0 26257.5 23090.0 26322.5 ;
      RECT  23057.5 26257.5 23320.0 26322.5 ;
      RECT  23025.0 26290.0 23090.0 26565.0 ;
      RECT  23025.0 26497.5 23090.0 26632.5 ;
      RECT  23215.0 26497.5 23280.0 26632.5 ;
      RECT  23215.0 26497.5 23280.0 26632.5 ;
      RECT  23025.0 26497.5 23090.0 26632.5 ;
      RECT  23025.0 27357.5 23090.0 27492.5 ;
      RECT  23215.0 27357.5 23280.0 27492.5 ;
      RECT  23215.0 27357.5 23280.0 27492.5 ;
      RECT  23025.0 27357.5 23090.0 27492.5 ;
      RECT  22952.5 27772.5 23017.5 27907.5 ;
      RECT  23287.5 26222.5 23352.5 26357.5 ;
      RECT  23025.0 27357.5 23090.0 27492.5 ;
      RECT  23215.0 26497.5 23280.0 26632.5 ;
      RECT  23472.5 26397.5 23537.5 26532.5 ;
      RECT  23472.5 26397.5 23537.5 26532.5 ;
      RECT  23920.0 27807.5 23985.0 27872.5 ;
      RECT  23655.0 27807.5 23952.5 27872.5 ;
      RECT  23920.0 27425.0 23985.0 27840.0 ;
      RECT  23730.0 26257.5 23795.0 26322.5 ;
      RECT  23762.5 26257.5 24025.0 26322.5 ;
      RECT  23730.0 26290.0 23795.0 26565.0 ;
      RECT  23730.0 26497.5 23795.0 26632.5 ;
      RECT  23920.0 26497.5 23985.0 26632.5 ;
      RECT  23920.0 26497.5 23985.0 26632.5 ;
      RECT  23730.0 26497.5 23795.0 26632.5 ;
      RECT  23730.0 27357.5 23795.0 27492.5 ;
      RECT  23920.0 27357.5 23985.0 27492.5 ;
      RECT  23920.0 27357.5 23985.0 27492.5 ;
      RECT  23730.0 27357.5 23795.0 27492.5 ;
      RECT  23657.5 27772.5 23722.5 27907.5 ;
      RECT  23992.5 26222.5 24057.5 26357.5 ;
      RECT  23730.0 27357.5 23795.0 27492.5 ;
      RECT  23920.0 26497.5 23985.0 26632.5 ;
      RECT  24177.5 26397.5 24242.5 26532.5 ;
      RECT  24177.5 26397.5 24242.5 26532.5 ;
      RECT  24625.0 27807.5 24690.0 27872.5 ;
      RECT  24360.0 27807.5 24657.5 27872.5 ;
      RECT  24625.0 27425.0 24690.0 27840.0 ;
      RECT  24435.0 26257.5 24500.0 26322.5 ;
      RECT  24467.5 26257.5 24730.0 26322.5 ;
      RECT  24435.0 26290.0 24500.0 26565.0 ;
      RECT  24435.0 26497.5 24500.0 26632.5 ;
      RECT  24625.0 26497.5 24690.0 26632.5 ;
      RECT  24625.0 26497.5 24690.0 26632.5 ;
      RECT  24435.0 26497.5 24500.0 26632.5 ;
      RECT  24435.0 27357.5 24500.0 27492.5 ;
      RECT  24625.0 27357.5 24690.0 27492.5 ;
      RECT  24625.0 27357.5 24690.0 27492.5 ;
      RECT  24435.0 27357.5 24500.0 27492.5 ;
      RECT  24362.5 27772.5 24427.5 27907.5 ;
      RECT  24697.5 26222.5 24762.5 26357.5 ;
      RECT  24435.0 27357.5 24500.0 27492.5 ;
      RECT  24625.0 26497.5 24690.0 26632.5 ;
      RECT  24882.5 26397.5 24947.5 26532.5 ;
      RECT  24882.5 26397.5 24947.5 26532.5 ;
      RECT  25330.0 27807.5 25395.0 27872.5 ;
      RECT  25065.0 27807.5 25362.5 27872.5 ;
      RECT  25330.0 27425.0 25395.0 27840.0 ;
      RECT  25140.0 26257.5 25205.0 26322.5 ;
      RECT  25172.5 26257.5 25435.0 26322.5 ;
      RECT  25140.0 26290.0 25205.0 26565.0 ;
      RECT  25140.0 26497.5 25205.0 26632.5 ;
      RECT  25330.0 26497.5 25395.0 26632.5 ;
      RECT  25330.0 26497.5 25395.0 26632.5 ;
      RECT  25140.0 26497.5 25205.0 26632.5 ;
      RECT  25140.0 27357.5 25205.0 27492.5 ;
      RECT  25330.0 27357.5 25395.0 27492.5 ;
      RECT  25330.0 27357.5 25395.0 27492.5 ;
      RECT  25140.0 27357.5 25205.0 27492.5 ;
      RECT  25067.5 27772.5 25132.5 27907.5 ;
      RECT  25402.5 26222.5 25467.5 26357.5 ;
      RECT  25140.0 27357.5 25205.0 27492.5 ;
      RECT  25330.0 26497.5 25395.0 26632.5 ;
      RECT  25587.5 26397.5 25652.5 26532.5 ;
      RECT  25587.5 26397.5 25652.5 26532.5 ;
      RECT  26035.0 27807.5 26100.0 27872.5 ;
      RECT  25770.0 27807.5 26067.5 27872.5 ;
      RECT  26035.0 27425.0 26100.0 27840.0 ;
      RECT  25845.0 26257.5 25910.0 26322.5 ;
      RECT  25877.5 26257.5 26140.0 26322.5 ;
      RECT  25845.0 26290.0 25910.0 26565.0 ;
      RECT  25845.0 26497.5 25910.0 26632.5 ;
      RECT  26035.0 26497.5 26100.0 26632.5 ;
      RECT  26035.0 26497.5 26100.0 26632.5 ;
      RECT  25845.0 26497.5 25910.0 26632.5 ;
      RECT  25845.0 27357.5 25910.0 27492.5 ;
      RECT  26035.0 27357.5 26100.0 27492.5 ;
      RECT  26035.0 27357.5 26100.0 27492.5 ;
      RECT  25845.0 27357.5 25910.0 27492.5 ;
      RECT  25772.5 27772.5 25837.5 27907.5 ;
      RECT  26107.5 26222.5 26172.5 26357.5 ;
      RECT  25845.0 27357.5 25910.0 27492.5 ;
      RECT  26035.0 26497.5 26100.0 26632.5 ;
      RECT  26292.5 26397.5 26357.5 26532.5 ;
      RECT  26292.5 26397.5 26357.5 26532.5 ;
      RECT  26740.0 27807.5 26805.0 27872.5 ;
      RECT  26475.0 27807.5 26772.5 27872.5 ;
      RECT  26740.0 27425.0 26805.0 27840.0 ;
      RECT  26550.0 26257.5 26615.0 26322.5 ;
      RECT  26582.5 26257.5 26845.0 26322.5 ;
      RECT  26550.0 26290.0 26615.0 26565.0 ;
      RECT  26550.0 26497.5 26615.0 26632.5 ;
      RECT  26740.0 26497.5 26805.0 26632.5 ;
      RECT  26740.0 26497.5 26805.0 26632.5 ;
      RECT  26550.0 26497.5 26615.0 26632.5 ;
      RECT  26550.0 27357.5 26615.0 27492.5 ;
      RECT  26740.0 27357.5 26805.0 27492.5 ;
      RECT  26740.0 27357.5 26805.0 27492.5 ;
      RECT  26550.0 27357.5 26615.0 27492.5 ;
      RECT  26477.5 27772.5 26542.5 27907.5 ;
      RECT  26812.5 26222.5 26877.5 26357.5 ;
      RECT  26550.0 27357.5 26615.0 27492.5 ;
      RECT  26740.0 26497.5 26805.0 26632.5 ;
      RECT  26997.5 26397.5 27062.5 26532.5 ;
      RECT  26997.5 26397.5 27062.5 26532.5 ;
      RECT  27445.0 27807.5 27510.0 27872.5 ;
      RECT  27180.0 27807.5 27477.5 27872.5 ;
      RECT  27445.0 27425.0 27510.0 27840.0 ;
      RECT  27255.0 26257.5 27320.0 26322.5 ;
      RECT  27287.5 26257.5 27550.0 26322.5 ;
      RECT  27255.0 26290.0 27320.0 26565.0 ;
      RECT  27255.0 26497.5 27320.0 26632.5 ;
      RECT  27445.0 26497.5 27510.0 26632.5 ;
      RECT  27445.0 26497.5 27510.0 26632.5 ;
      RECT  27255.0 26497.5 27320.0 26632.5 ;
      RECT  27255.0 27357.5 27320.0 27492.5 ;
      RECT  27445.0 27357.5 27510.0 27492.5 ;
      RECT  27445.0 27357.5 27510.0 27492.5 ;
      RECT  27255.0 27357.5 27320.0 27492.5 ;
      RECT  27182.5 27772.5 27247.5 27907.5 ;
      RECT  27517.5 26222.5 27582.5 26357.5 ;
      RECT  27255.0 27357.5 27320.0 27492.5 ;
      RECT  27445.0 26497.5 27510.0 26632.5 ;
      RECT  27702.5 26397.5 27767.5 26532.5 ;
      RECT  27702.5 26397.5 27767.5 26532.5 ;
      RECT  28150.0 27807.5 28215.0 27872.5 ;
      RECT  27885.0 27807.5 28182.5 27872.5 ;
      RECT  28150.0 27425.0 28215.0 27840.0 ;
      RECT  27960.0 26257.5 28025.0 26322.5 ;
      RECT  27992.5 26257.5 28255.0 26322.5 ;
      RECT  27960.0 26290.0 28025.0 26565.0 ;
      RECT  27960.0 26497.5 28025.0 26632.5 ;
      RECT  28150.0 26497.5 28215.0 26632.5 ;
      RECT  28150.0 26497.5 28215.0 26632.5 ;
      RECT  27960.0 26497.5 28025.0 26632.5 ;
      RECT  27960.0 27357.5 28025.0 27492.5 ;
      RECT  28150.0 27357.5 28215.0 27492.5 ;
      RECT  28150.0 27357.5 28215.0 27492.5 ;
      RECT  27960.0 27357.5 28025.0 27492.5 ;
      RECT  27887.5 27772.5 27952.5 27907.5 ;
      RECT  28222.5 26222.5 28287.5 26357.5 ;
      RECT  27960.0 27357.5 28025.0 27492.5 ;
      RECT  28150.0 26497.5 28215.0 26632.5 ;
      RECT  28407.5 26397.5 28472.5 26532.5 ;
      RECT  28407.5 26397.5 28472.5 26532.5 ;
      RECT  28855.0 27807.5 28920.0 27872.5 ;
      RECT  28590.0 27807.5 28887.5 27872.5 ;
      RECT  28855.0 27425.0 28920.0 27840.0 ;
      RECT  28665.0 26257.5 28730.0 26322.5 ;
      RECT  28697.5 26257.5 28960.0 26322.5 ;
      RECT  28665.0 26290.0 28730.0 26565.0 ;
      RECT  28665.0 26497.5 28730.0 26632.5 ;
      RECT  28855.0 26497.5 28920.0 26632.5 ;
      RECT  28855.0 26497.5 28920.0 26632.5 ;
      RECT  28665.0 26497.5 28730.0 26632.5 ;
      RECT  28665.0 27357.5 28730.0 27492.5 ;
      RECT  28855.0 27357.5 28920.0 27492.5 ;
      RECT  28855.0 27357.5 28920.0 27492.5 ;
      RECT  28665.0 27357.5 28730.0 27492.5 ;
      RECT  28592.5 27772.5 28657.5 27907.5 ;
      RECT  28927.5 26222.5 28992.5 26357.5 ;
      RECT  28665.0 27357.5 28730.0 27492.5 ;
      RECT  28855.0 26497.5 28920.0 26632.5 ;
      RECT  29112.5 26397.5 29177.5 26532.5 ;
      RECT  29112.5 26397.5 29177.5 26532.5 ;
      RECT  29560.0 27807.5 29625.0 27872.5 ;
      RECT  29295.0 27807.5 29592.5 27872.5 ;
      RECT  29560.0 27425.0 29625.0 27840.0 ;
      RECT  29370.0 26257.5 29435.0 26322.5 ;
      RECT  29402.5 26257.5 29665.0 26322.5 ;
      RECT  29370.0 26290.0 29435.0 26565.0 ;
      RECT  29370.0 26497.5 29435.0 26632.5 ;
      RECT  29560.0 26497.5 29625.0 26632.5 ;
      RECT  29560.0 26497.5 29625.0 26632.5 ;
      RECT  29370.0 26497.5 29435.0 26632.5 ;
      RECT  29370.0 27357.5 29435.0 27492.5 ;
      RECT  29560.0 27357.5 29625.0 27492.5 ;
      RECT  29560.0 27357.5 29625.0 27492.5 ;
      RECT  29370.0 27357.5 29435.0 27492.5 ;
      RECT  29297.5 27772.5 29362.5 27907.5 ;
      RECT  29632.5 26222.5 29697.5 26357.5 ;
      RECT  29370.0 27357.5 29435.0 27492.5 ;
      RECT  29560.0 26497.5 29625.0 26632.5 ;
      RECT  29817.5 26397.5 29882.5 26532.5 ;
      RECT  29817.5 26397.5 29882.5 26532.5 ;
      RECT  30265.0 27807.5 30330.0 27872.5 ;
      RECT  30000.0 27807.5 30297.5 27872.5 ;
      RECT  30265.0 27425.0 30330.0 27840.0 ;
      RECT  30075.0 26257.5 30140.0 26322.5 ;
      RECT  30107.5 26257.5 30370.0 26322.5 ;
      RECT  30075.0 26290.0 30140.0 26565.0 ;
      RECT  30075.0 26497.5 30140.0 26632.5 ;
      RECT  30265.0 26497.5 30330.0 26632.5 ;
      RECT  30265.0 26497.5 30330.0 26632.5 ;
      RECT  30075.0 26497.5 30140.0 26632.5 ;
      RECT  30075.0 27357.5 30140.0 27492.5 ;
      RECT  30265.0 27357.5 30330.0 27492.5 ;
      RECT  30265.0 27357.5 30330.0 27492.5 ;
      RECT  30075.0 27357.5 30140.0 27492.5 ;
      RECT  30002.5 27772.5 30067.5 27907.5 ;
      RECT  30337.5 26222.5 30402.5 26357.5 ;
      RECT  30075.0 27357.5 30140.0 27492.5 ;
      RECT  30265.0 26497.5 30330.0 26632.5 ;
      RECT  30522.5 26397.5 30587.5 26532.5 ;
      RECT  30522.5 26397.5 30587.5 26532.5 ;
      RECT  30970.0 27807.5 31035.0 27872.5 ;
      RECT  30705.0 27807.5 31002.5 27872.5 ;
      RECT  30970.0 27425.0 31035.0 27840.0 ;
      RECT  30780.0 26257.5 30845.0 26322.5 ;
      RECT  30812.5 26257.5 31075.0 26322.5 ;
      RECT  30780.0 26290.0 30845.0 26565.0 ;
      RECT  30780.0 26497.5 30845.0 26632.5 ;
      RECT  30970.0 26497.5 31035.0 26632.5 ;
      RECT  30970.0 26497.5 31035.0 26632.5 ;
      RECT  30780.0 26497.5 30845.0 26632.5 ;
      RECT  30780.0 27357.5 30845.0 27492.5 ;
      RECT  30970.0 27357.5 31035.0 27492.5 ;
      RECT  30970.0 27357.5 31035.0 27492.5 ;
      RECT  30780.0 27357.5 30845.0 27492.5 ;
      RECT  30707.5 27772.5 30772.5 27907.5 ;
      RECT  31042.5 26222.5 31107.5 26357.5 ;
      RECT  30780.0 27357.5 30845.0 27492.5 ;
      RECT  30970.0 26497.5 31035.0 26632.5 ;
      RECT  31227.5 26397.5 31292.5 26532.5 ;
      RECT  31227.5 26397.5 31292.5 26532.5 ;
      RECT  31675.0 27807.5 31740.0 27872.5 ;
      RECT  31410.0 27807.5 31707.5 27872.5 ;
      RECT  31675.0 27425.0 31740.0 27840.0 ;
      RECT  31485.0 26257.5 31550.0 26322.5 ;
      RECT  31517.5 26257.5 31780.0 26322.5 ;
      RECT  31485.0 26290.0 31550.0 26565.0 ;
      RECT  31485.0 26497.5 31550.0 26632.5 ;
      RECT  31675.0 26497.5 31740.0 26632.5 ;
      RECT  31675.0 26497.5 31740.0 26632.5 ;
      RECT  31485.0 26497.5 31550.0 26632.5 ;
      RECT  31485.0 27357.5 31550.0 27492.5 ;
      RECT  31675.0 27357.5 31740.0 27492.5 ;
      RECT  31675.0 27357.5 31740.0 27492.5 ;
      RECT  31485.0 27357.5 31550.0 27492.5 ;
      RECT  31412.5 27772.5 31477.5 27907.5 ;
      RECT  31747.5 26222.5 31812.5 26357.5 ;
      RECT  31485.0 27357.5 31550.0 27492.5 ;
      RECT  31675.0 26497.5 31740.0 26632.5 ;
      RECT  31932.5 26397.5 31997.5 26532.5 ;
      RECT  31932.5 26397.5 31997.5 26532.5 ;
      RECT  32380.0 27807.5 32445.0 27872.5 ;
      RECT  32115.0 27807.5 32412.5 27872.5 ;
      RECT  32380.0 27425.0 32445.0 27840.0 ;
      RECT  32190.0 26257.5 32255.0 26322.5 ;
      RECT  32222.5 26257.5 32485.0 26322.5 ;
      RECT  32190.0 26290.0 32255.0 26565.0 ;
      RECT  32190.0 26497.5 32255.0 26632.5 ;
      RECT  32380.0 26497.5 32445.0 26632.5 ;
      RECT  32380.0 26497.5 32445.0 26632.5 ;
      RECT  32190.0 26497.5 32255.0 26632.5 ;
      RECT  32190.0 27357.5 32255.0 27492.5 ;
      RECT  32380.0 27357.5 32445.0 27492.5 ;
      RECT  32380.0 27357.5 32445.0 27492.5 ;
      RECT  32190.0 27357.5 32255.0 27492.5 ;
      RECT  32117.5 27772.5 32182.5 27907.5 ;
      RECT  32452.5 26222.5 32517.5 26357.5 ;
      RECT  32190.0 27357.5 32255.0 27492.5 ;
      RECT  32380.0 26497.5 32445.0 26632.5 ;
      RECT  32637.5 26397.5 32702.5 26532.5 ;
      RECT  32637.5 26397.5 32702.5 26532.5 ;
      RECT  33085.0 27807.5 33150.0 27872.5 ;
      RECT  32820.0 27807.5 33117.5 27872.5 ;
      RECT  33085.0 27425.0 33150.0 27840.0 ;
      RECT  32895.0 26257.5 32960.0 26322.5 ;
      RECT  32927.5 26257.5 33190.0 26322.5 ;
      RECT  32895.0 26290.0 32960.0 26565.0 ;
      RECT  32895.0 26497.5 32960.0 26632.5 ;
      RECT  33085.0 26497.5 33150.0 26632.5 ;
      RECT  33085.0 26497.5 33150.0 26632.5 ;
      RECT  32895.0 26497.5 32960.0 26632.5 ;
      RECT  32895.0 27357.5 32960.0 27492.5 ;
      RECT  33085.0 27357.5 33150.0 27492.5 ;
      RECT  33085.0 27357.5 33150.0 27492.5 ;
      RECT  32895.0 27357.5 32960.0 27492.5 ;
      RECT  32822.5 27772.5 32887.5 27907.5 ;
      RECT  33157.5 26222.5 33222.5 26357.5 ;
      RECT  32895.0 27357.5 32960.0 27492.5 ;
      RECT  33085.0 26497.5 33150.0 26632.5 ;
      RECT  33342.5 26397.5 33407.5 26532.5 ;
      RECT  33342.5 26397.5 33407.5 26532.5 ;
      RECT  33790.0 27807.5 33855.0 27872.5 ;
      RECT  33525.0 27807.5 33822.5 27872.5 ;
      RECT  33790.0 27425.0 33855.0 27840.0 ;
      RECT  33600.0 26257.5 33665.0 26322.5 ;
      RECT  33632.5 26257.5 33895.0 26322.5 ;
      RECT  33600.0 26290.0 33665.0 26565.0 ;
      RECT  33600.0 26497.5 33665.0 26632.5 ;
      RECT  33790.0 26497.5 33855.0 26632.5 ;
      RECT  33790.0 26497.5 33855.0 26632.5 ;
      RECT  33600.0 26497.5 33665.0 26632.5 ;
      RECT  33600.0 27357.5 33665.0 27492.5 ;
      RECT  33790.0 27357.5 33855.0 27492.5 ;
      RECT  33790.0 27357.5 33855.0 27492.5 ;
      RECT  33600.0 27357.5 33665.0 27492.5 ;
      RECT  33527.5 27772.5 33592.5 27907.5 ;
      RECT  33862.5 26222.5 33927.5 26357.5 ;
      RECT  33600.0 27357.5 33665.0 27492.5 ;
      RECT  33790.0 26497.5 33855.0 26632.5 ;
      RECT  34047.5 26397.5 34112.5 26532.5 ;
      RECT  34047.5 26397.5 34112.5 26532.5 ;
      RECT  34495.0 27807.5 34560.0 27872.5 ;
      RECT  34230.0 27807.5 34527.5 27872.5 ;
      RECT  34495.0 27425.0 34560.0 27840.0 ;
      RECT  34305.0 26257.5 34370.0 26322.5 ;
      RECT  34337.5 26257.5 34600.0 26322.5 ;
      RECT  34305.0 26290.0 34370.0 26565.0 ;
      RECT  34305.0 26497.5 34370.0 26632.5 ;
      RECT  34495.0 26497.5 34560.0 26632.5 ;
      RECT  34495.0 26497.5 34560.0 26632.5 ;
      RECT  34305.0 26497.5 34370.0 26632.5 ;
      RECT  34305.0 27357.5 34370.0 27492.5 ;
      RECT  34495.0 27357.5 34560.0 27492.5 ;
      RECT  34495.0 27357.5 34560.0 27492.5 ;
      RECT  34305.0 27357.5 34370.0 27492.5 ;
      RECT  34232.5 27772.5 34297.5 27907.5 ;
      RECT  34567.5 26222.5 34632.5 26357.5 ;
      RECT  34305.0 27357.5 34370.0 27492.5 ;
      RECT  34495.0 26497.5 34560.0 26632.5 ;
      RECT  34752.5 26397.5 34817.5 26532.5 ;
      RECT  34752.5 26397.5 34817.5 26532.5 ;
      RECT  35200.0 27807.5 35265.0 27872.5 ;
      RECT  34935.0 27807.5 35232.5 27872.5 ;
      RECT  35200.0 27425.0 35265.0 27840.0 ;
      RECT  35010.0 26257.5 35075.0 26322.5 ;
      RECT  35042.5 26257.5 35305.0 26322.5 ;
      RECT  35010.0 26290.0 35075.0 26565.0 ;
      RECT  35010.0 26497.5 35075.0 26632.5 ;
      RECT  35200.0 26497.5 35265.0 26632.5 ;
      RECT  35200.0 26497.5 35265.0 26632.5 ;
      RECT  35010.0 26497.5 35075.0 26632.5 ;
      RECT  35010.0 27357.5 35075.0 27492.5 ;
      RECT  35200.0 27357.5 35265.0 27492.5 ;
      RECT  35200.0 27357.5 35265.0 27492.5 ;
      RECT  35010.0 27357.5 35075.0 27492.5 ;
      RECT  34937.5 27772.5 35002.5 27907.5 ;
      RECT  35272.5 26222.5 35337.5 26357.5 ;
      RECT  35010.0 27357.5 35075.0 27492.5 ;
      RECT  35200.0 26497.5 35265.0 26632.5 ;
      RECT  35457.5 26397.5 35522.5 26532.5 ;
      RECT  35457.5 26397.5 35522.5 26532.5 ;
      RECT  35905.0 27807.5 35970.0 27872.5 ;
      RECT  35640.0 27807.5 35937.5 27872.5 ;
      RECT  35905.0 27425.0 35970.0 27840.0 ;
      RECT  35715.0 26257.5 35780.0 26322.5 ;
      RECT  35747.5 26257.5 36010.0 26322.5 ;
      RECT  35715.0 26290.0 35780.0 26565.0 ;
      RECT  35715.0 26497.5 35780.0 26632.5 ;
      RECT  35905.0 26497.5 35970.0 26632.5 ;
      RECT  35905.0 26497.5 35970.0 26632.5 ;
      RECT  35715.0 26497.5 35780.0 26632.5 ;
      RECT  35715.0 27357.5 35780.0 27492.5 ;
      RECT  35905.0 27357.5 35970.0 27492.5 ;
      RECT  35905.0 27357.5 35970.0 27492.5 ;
      RECT  35715.0 27357.5 35780.0 27492.5 ;
      RECT  35642.5 27772.5 35707.5 27907.5 ;
      RECT  35977.5 26222.5 36042.5 26357.5 ;
      RECT  35715.0 27357.5 35780.0 27492.5 ;
      RECT  35905.0 26497.5 35970.0 26632.5 ;
      RECT  36162.5 26397.5 36227.5 26532.5 ;
      RECT  36162.5 26397.5 36227.5 26532.5 ;
      RECT  36610.0 27807.5 36675.0 27872.5 ;
      RECT  36345.0 27807.5 36642.5 27872.5 ;
      RECT  36610.0 27425.0 36675.0 27840.0 ;
      RECT  36420.0 26257.5 36485.0 26322.5 ;
      RECT  36452.5 26257.5 36715.0 26322.5 ;
      RECT  36420.0 26290.0 36485.0 26565.0 ;
      RECT  36420.0 26497.5 36485.0 26632.5 ;
      RECT  36610.0 26497.5 36675.0 26632.5 ;
      RECT  36610.0 26497.5 36675.0 26632.5 ;
      RECT  36420.0 26497.5 36485.0 26632.5 ;
      RECT  36420.0 27357.5 36485.0 27492.5 ;
      RECT  36610.0 27357.5 36675.0 27492.5 ;
      RECT  36610.0 27357.5 36675.0 27492.5 ;
      RECT  36420.0 27357.5 36485.0 27492.5 ;
      RECT  36347.5 27772.5 36412.5 27907.5 ;
      RECT  36682.5 26222.5 36747.5 26357.5 ;
      RECT  36420.0 27357.5 36485.0 27492.5 ;
      RECT  36610.0 26497.5 36675.0 26632.5 ;
      RECT  36867.5 26397.5 36932.5 26532.5 ;
      RECT  36867.5 26397.5 36932.5 26532.5 ;
      RECT  37315.0 27807.5 37380.0 27872.5 ;
      RECT  37050.0 27807.5 37347.5 27872.5 ;
      RECT  37315.0 27425.0 37380.0 27840.0 ;
      RECT  37125.0 26257.5 37190.0 26322.5 ;
      RECT  37157.5 26257.5 37420.0 26322.5 ;
      RECT  37125.0 26290.0 37190.0 26565.0 ;
      RECT  37125.0 26497.5 37190.0 26632.5 ;
      RECT  37315.0 26497.5 37380.0 26632.5 ;
      RECT  37315.0 26497.5 37380.0 26632.5 ;
      RECT  37125.0 26497.5 37190.0 26632.5 ;
      RECT  37125.0 27357.5 37190.0 27492.5 ;
      RECT  37315.0 27357.5 37380.0 27492.5 ;
      RECT  37315.0 27357.5 37380.0 27492.5 ;
      RECT  37125.0 27357.5 37190.0 27492.5 ;
      RECT  37052.5 27772.5 37117.5 27907.5 ;
      RECT  37387.5 26222.5 37452.5 26357.5 ;
      RECT  37125.0 27357.5 37190.0 27492.5 ;
      RECT  37315.0 26497.5 37380.0 26632.5 ;
      RECT  37572.5 26397.5 37637.5 26532.5 ;
      RECT  37572.5 26397.5 37637.5 26532.5 ;
      RECT  38020.0 27807.5 38085.0 27872.5 ;
      RECT  37755.0 27807.5 38052.5 27872.5 ;
      RECT  38020.0 27425.0 38085.0 27840.0 ;
      RECT  37830.0 26257.5 37895.0 26322.5 ;
      RECT  37862.5 26257.5 38125.0 26322.5 ;
      RECT  37830.0 26290.0 37895.0 26565.0 ;
      RECT  37830.0 26497.5 37895.0 26632.5 ;
      RECT  38020.0 26497.5 38085.0 26632.5 ;
      RECT  38020.0 26497.5 38085.0 26632.5 ;
      RECT  37830.0 26497.5 37895.0 26632.5 ;
      RECT  37830.0 27357.5 37895.0 27492.5 ;
      RECT  38020.0 27357.5 38085.0 27492.5 ;
      RECT  38020.0 27357.5 38085.0 27492.5 ;
      RECT  37830.0 27357.5 37895.0 27492.5 ;
      RECT  37757.5 27772.5 37822.5 27907.5 ;
      RECT  38092.5 26222.5 38157.5 26357.5 ;
      RECT  37830.0 27357.5 37895.0 27492.5 ;
      RECT  38020.0 26497.5 38085.0 26632.5 ;
      RECT  38277.5 26397.5 38342.5 26532.5 ;
      RECT  38277.5 26397.5 38342.5 26532.5 ;
      RECT  38725.0 27807.5 38790.0 27872.5 ;
      RECT  38460.0 27807.5 38757.5 27872.5 ;
      RECT  38725.0 27425.0 38790.0 27840.0 ;
      RECT  38535.0 26257.5 38600.0 26322.5 ;
      RECT  38567.5 26257.5 38830.0 26322.5 ;
      RECT  38535.0 26290.0 38600.0 26565.0 ;
      RECT  38535.0 26497.5 38600.0 26632.5 ;
      RECT  38725.0 26497.5 38790.0 26632.5 ;
      RECT  38725.0 26497.5 38790.0 26632.5 ;
      RECT  38535.0 26497.5 38600.0 26632.5 ;
      RECT  38535.0 27357.5 38600.0 27492.5 ;
      RECT  38725.0 27357.5 38790.0 27492.5 ;
      RECT  38725.0 27357.5 38790.0 27492.5 ;
      RECT  38535.0 27357.5 38600.0 27492.5 ;
      RECT  38462.5 27772.5 38527.5 27907.5 ;
      RECT  38797.5 26222.5 38862.5 26357.5 ;
      RECT  38535.0 27357.5 38600.0 27492.5 ;
      RECT  38725.0 26497.5 38790.0 26632.5 ;
      RECT  38982.5 26397.5 39047.5 26532.5 ;
      RECT  38982.5 26397.5 39047.5 26532.5 ;
      RECT  39430.0 27807.5 39495.0 27872.5 ;
      RECT  39165.0 27807.5 39462.5 27872.5 ;
      RECT  39430.0 27425.0 39495.0 27840.0 ;
      RECT  39240.0 26257.5 39305.0 26322.5 ;
      RECT  39272.5 26257.5 39535.0 26322.5 ;
      RECT  39240.0 26290.0 39305.0 26565.0 ;
      RECT  39240.0 26497.5 39305.0 26632.5 ;
      RECT  39430.0 26497.5 39495.0 26632.5 ;
      RECT  39430.0 26497.5 39495.0 26632.5 ;
      RECT  39240.0 26497.5 39305.0 26632.5 ;
      RECT  39240.0 27357.5 39305.0 27492.5 ;
      RECT  39430.0 27357.5 39495.0 27492.5 ;
      RECT  39430.0 27357.5 39495.0 27492.5 ;
      RECT  39240.0 27357.5 39305.0 27492.5 ;
      RECT  39167.5 27772.5 39232.5 27907.5 ;
      RECT  39502.5 26222.5 39567.5 26357.5 ;
      RECT  39240.0 27357.5 39305.0 27492.5 ;
      RECT  39430.0 26497.5 39495.0 26632.5 ;
      RECT  39687.5 26397.5 39752.5 26532.5 ;
      RECT  39687.5 26397.5 39752.5 26532.5 ;
      RECT  40135.0 27807.5 40200.0 27872.5 ;
      RECT  39870.0 27807.5 40167.5 27872.5 ;
      RECT  40135.0 27425.0 40200.0 27840.0 ;
      RECT  39945.0 26257.5 40010.0 26322.5 ;
      RECT  39977.5 26257.5 40240.0 26322.5 ;
      RECT  39945.0 26290.0 40010.0 26565.0 ;
      RECT  39945.0 26497.5 40010.0 26632.5 ;
      RECT  40135.0 26497.5 40200.0 26632.5 ;
      RECT  40135.0 26497.5 40200.0 26632.5 ;
      RECT  39945.0 26497.5 40010.0 26632.5 ;
      RECT  39945.0 27357.5 40010.0 27492.5 ;
      RECT  40135.0 27357.5 40200.0 27492.5 ;
      RECT  40135.0 27357.5 40200.0 27492.5 ;
      RECT  39945.0 27357.5 40010.0 27492.5 ;
      RECT  39872.5 27772.5 39937.5 27907.5 ;
      RECT  40207.5 26222.5 40272.5 26357.5 ;
      RECT  39945.0 27357.5 40010.0 27492.5 ;
      RECT  40135.0 26497.5 40200.0 26632.5 ;
      RECT  40392.5 26397.5 40457.5 26532.5 ;
      RECT  40392.5 26397.5 40457.5 26532.5 ;
      RECT  40840.0 27807.5 40905.0 27872.5 ;
      RECT  40575.0 27807.5 40872.5 27872.5 ;
      RECT  40840.0 27425.0 40905.0 27840.0 ;
      RECT  40650.0 26257.5 40715.0 26322.5 ;
      RECT  40682.5 26257.5 40945.0 26322.5 ;
      RECT  40650.0 26290.0 40715.0 26565.0 ;
      RECT  40650.0 26497.5 40715.0 26632.5 ;
      RECT  40840.0 26497.5 40905.0 26632.5 ;
      RECT  40840.0 26497.5 40905.0 26632.5 ;
      RECT  40650.0 26497.5 40715.0 26632.5 ;
      RECT  40650.0 27357.5 40715.0 27492.5 ;
      RECT  40840.0 27357.5 40905.0 27492.5 ;
      RECT  40840.0 27357.5 40905.0 27492.5 ;
      RECT  40650.0 27357.5 40715.0 27492.5 ;
      RECT  40577.5 27772.5 40642.5 27907.5 ;
      RECT  40912.5 26222.5 40977.5 26357.5 ;
      RECT  40650.0 27357.5 40715.0 27492.5 ;
      RECT  40840.0 26497.5 40905.0 26632.5 ;
      RECT  41097.5 26397.5 41162.5 26532.5 ;
      RECT  41097.5 26397.5 41162.5 26532.5 ;
      RECT  41545.0 27807.5 41610.0 27872.5 ;
      RECT  41280.0 27807.5 41577.5 27872.5 ;
      RECT  41545.0 27425.0 41610.0 27840.0 ;
      RECT  41355.0 26257.5 41420.0 26322.5 ;
      RECT  41387.5 26257.5 41650.0 26322.5 ;
      RECT  41355.0 26290.0 41420.0 26565.0 ;
      RECT  41355.0 26497.5 41420.0 26632.5 ;
      RECT  41545.0 26497.5 41610.0 26632.5 ;
      RECT  41545.0 26497.5 41610.0 26632.5 ;
      RECT  41355.0 26497.5 41420.0 26632.5 ;
      RECT  41355.0 27357.5 41420.0 27492.5 ;
      RECT  41545.0 27357.5 41610.0 27492.5 ;
      RECT  41545.0 27357.5 41610.0 27492.5 ;
      RECT  41355.0 27357.5 41420.0 27492.5 ;
      RECT  41282.5 27772.5 41347.5 27907.5 ;
      RECT  41617.5 26222.5 41682.5 26357.5 ;
      RECT  41355.0 27357.5 41420.0 27492.5 ;
      RECT  41545.0 26497.5 41610.0 26632.5 ;
      RECT  41802.5 26397.5 41867.5 26532.5 ;
      RECT  41802.5 26397.5 41867.5 26532.5 ;
      RECT  42250.0 27807.5 42315.0 27872.5 ;
      RECT  41985.0 27807.5 42282.5 27872.5 ;
      RECT  42250.0 27425.0 42315.0 27840.0 ;
      RECT  42060.0 26257.5 42125.0 26322.5 ;
      RECT  42092.5 26257.5 42355.0 26322.5 ;
      RECT  42060.0 26290.0 42125.0 26565.0 ;
      RECT  42060.0 26497.5 42125.0 26632.5 ;
      RECT  42250.0 26497.5 42315.0 26632.5 ;
      RECT  42250.0 26497.5 42315.0 26632.5 ;
      RECT  42060.0 26497.5 42125.0 26632.5 ;
      RECT  42060.0 27357.5 42125.0 27492.5 ;
      RECT  42250.0 27357.5 42315.0 27492.5 ;
      RECT  42250.0 27357.5 42315.0 27492.5 ;
      RECT  42060.0 27357.5 42125.0 27492.5 ;
      RECT  41987.5 27772.5 42052.5 27907.5 ;
      RECT  42322.5 26222.5 42387.5 26357.5 ;
      RECT  42060.0 27357.5 42125.0 27492.5 ;
      RECT  42250.0 26497.5 42315.0 26632.5 ;
      RECT  42507.5 26397.5 42572.5 26532.5 ;
      RECT  42507.5 26397.5 42572.5 26532.5 ;
      RECT  42955.0 27807.5 43020.0 27872.5 ;
      RECT  42690.0 27807.5 42987.5 27872.5 ;
      RECT  42955.0 27425.0 43020.0 27840.0 ;
      RECT  42765.0 26257.5 42830.0 26322.5 ;
      RECT  42797.5 26257.5 43060.0 26322.5 ;
      RECT  42765.0 26290.0 42830.0 26565.0 ;
      RECT  42765.0 26497.5 42830.0 26632.5 ;
      RECT  42955.0 26497.5 43020.0 26632.5 ;
      RECT  42955.0 26497.5 43020.0 26632.5 ;
      RECT  42765.0 26497.5 42830.0 26632.5 ;
      RECT  42765.0 27357.5 42830.0 27492.5 ;
      RECT  42955.0 27357.5 43020.0 27492.5 ;
      RECT  42955.0 27357.5 43020.0 27492.5 ;
      RECT  42765.0 27357.5 42830.0 27492.5 ;
      RECT  42692.5 27772.5 42757.5 27907.5 ;
      RECT  43027.5 26222.5 43092.5 26357.5 ;
      RECT  42765.0 27357.5 42830.0 27492.5 ;
      RECT  42955.0 26497.5 43020.0 26632.5 ;
      RECT  43212.5 26397.5 43277.5 26532.5 ;
      RECT  43212.5 26397.5 43277.5 26532.5 ;
      RECT  43660.0 27807.5 43725.0 27872.5 ;
      RECT  43395.0 27807.5 43692.5 27872.5 ;
      RECT  43660.0 27425.0 43725.0 27840.0 ;
      RECT  43470.0 26257.5 43535.0 26322.5 ;
      RECT  43502.5 26257.5 43765.0 26322.5 ;
      RECT  43470.0 26290.0 43535.0 26565.0 ;
      RECT  43470.0 26497.5 43535.0 26632.5 ;
      RECT  43660.0 26497.5 43725.0 26632.5 ;
      RECT  43660.0 26497.5 43725.0 26632.5 ;
      RECT  43470.0 26497.5 43535.0 26632.5 ;
      RECT  43470.0 27357.5 43535.0 27492.5 ;
      RECT  43660.0 27357.5 43725.0 27492.5 ;
      RECT  43660.0 27357.5 43725.0 27492.5 ;
      RECT  43470.0 27357.5 43535.0 27492.5 ;
      RECT  43397.5 27772.5 43462.5 27907.5 ;
      RECT  43732.5 26222.5 43797.5 26357.5 ;
      RECT  43470.0 27357.5 43535.0 27492.5 ;
      RECT  43660.0 26497.5 43725.0 26632.5 ;
      RECT  43917.5 26397.5 43982.5 26532.5 ;
      RECT  43917.5 26397.5 43982.5 26532.5 ;
      RECT  44365.0 27807.5 44430.0 27872.5 ;
      RECT  44100.0 27807.5 44397.5 27872.5 ;
      RECT  44365.0 27425.0 44430.0 27840.0 ;
      RECT  44175.0 26257.5 44240.0 26322.5 ;
      RECT  44207.5 26257.5 44470.0 26322.5 ;
      RECT  44175.0 26290.0 44240.0 26565.0 ;
      RECT  44175.0 26497.5 44240.0 26632.5 ;
      RECT  44365.0 26497.5 44430.0 26632.5 ;
      RECT  44365.0 26497.5 44430.0 26632.5 ;
      RECT  44175.0 26497.5 44240.0 26632.5 ;
      RECT  44175.0 27357.5 44240.0 27492.5 ;
      RECT  44365.0 27357.5 44430.0 27492.5 ;
      RECT  44365.0 27357.5 44430.0 27492.5 ;
      RECT  44175.0 27357.5 44240.0 27492.5 ;
      RECT  44102.5 27772.5 44167.5 27907.5 ;
      RECT  44437.5 26222.5 44502.5 26357.5 ;
      RECT  44175.0 27357.5 44240.0 27492.5 ;
      RECT  44365.0 26497.5 44430.0 26632.5 ;
      RECT  44622.5 26397.5 44687.5 26532.5 ;
      RECT  44622.5 26397.5 44687.5 26532.5 ;
      RECT  45070.0 27807.5 45135.0 27872.5 ;
      RECT  44805.0 27807.5 45102.5 27872.5 ;
      RECT  45070.0 27425.0 45135.0 27840.0 ;
      RECT  44880.0 26257.5 44945.0 26322.5 ;
      RECT  44912.5 26257.5 45175.0 26322.5 ;
      RECT  44880.0 26290.0 44945.0 26565.0 ;
      RECT  44880.0 26497.5 44945.0 26632.5 ;
      RECT  45070.0 26497.5 45135.0 26632.5 ;
      RECT  45070.0 26497.5 45135.0 26632.5 ;
      RECT  44880.0 26497.5 44945.0 26632.5 ;
      RECT  44880.0 27357.5 44945.0 27492.5 ;
      RECT  45070.0 27357.5 45135.0 27492.5 ;
      RECT  45070.0 27357.5 45135.0 27492.5 ;
      RECT  44880.0 27357.5 44945.0 27492.5 ;
      RECT  44807.5 27772.5 44872.5 27907.5 ;
      RECT  45142.5 26222.5 45207.5 26357.5 ;
      RECT  44880.0 27357.5 44945.0 27492.5 ;
      RECT  45070.0 26497.5 45135.0 26632.5 ;
      RECT  45327.5 26397.5 45392.5 26532.5 ;
      RECT  45327.5 26397.5 45392.5 26532.5 ;
      RECT  45775.0 27807.5 45840.0 27872.5 ;
      RECT  45510.0 27807.5 45807.5 27872.5 ;
      RECT  45775.0 27425.0 45840.0 27840.0 ;
      RECT  45585.0 26257.5 45650.0 26322.5 ;
      RECT  45617.5 26257.5 45880.0 26322.5 ;
      RECT  45585.0 26290.0 45650.0 26565.0 ;
      RECT  45585.0 26497.5 45650.0 26632.5 ;
      RECT  45775.0 26497.5 45840.0 26632.5 ;
      RECT  45775.0 26497.5 45840.0 26632.5 ;
      RECT  45585.0 26497.5 45650.0 26632.5 ;
      RECT  45585.0 27357.5 45650.0 27492.5 ;
      RECT  45775.0 27357.5 45840.0 27492.5 ;
      RECT  45775.0 27357.5 45840.0 27492.5 ;
      RECT  45585.0 27357.5 45650.0 27492.5 ;
      RECT  45512.5 27772.5 45577.5 27907.5 ;
      RECT  45847.5 26222.5 45912.5 26357.5 ;
      RECT  45585.0 27357.5 45650.0 27492.5 ;
      RECT  45775.0 26497.5 45840.0 26632.5 ;
      RECT  46032.5 26397.5 46097.5 26532.5 ;
      RECT  46032.5 26397.5 46097.5 26532.5 ;
      RECT  46480.0 27807.5 46545.0 27872.5 ;
      RECT  46215.0 27807.5 46512.5 27872.5 ;
      RECT  46480.0 27425.0 46545.0 27840.0 ;
      RECT  46290.0 26257.5 46355.0 26322.5 ;
      RECT  46322.5 26257.5 46585.0 26322.5 ;
      RECT  46290.0 26290.0 46355.0 26565.0 ;
      RECT  46290.0 26497.5 46355.0 26632.5 ;
      RECT  46480.0 26497.5 46545.0 26632.5 ;
      RECT  46480.0 26497.5 46545.0 26632.5 ;
      RECT  46290.0 26497.5 46355.0 26632.5 ;
      RECT  46290.0 27357.5 46355.0 27492.5 ;
      RECT  46480.0 27357.5 46545.0 27492.5 ;
      RECT  46480.0 27357.5 46545.0 27492.5 ;
      RECT  46290.0 27357.5 46355.0 27492.5 ;
      RECT  46217.5 27772.5 46282.5 27907.5 ;
      RECT  46552.5 26222.5 46617.5 26357.5 ;
      RECT  46290.0 27357.5 46355.0 27492.5 ;
      RECT  46480.0 26497.5 46545.0 26632.5 ;
      RECT  46737.5 26397.5 46802.5 26532.5 ;
      RECT  46737.5 26397.5 46802.5 26532.5 ;
      RECT  47185.0 27807.5 47250.0 27872.5 ;
      RECT  46920.0 27807.5 47217.5 27872.5 ;
      RECT  47185.0 27425.0 47250.0 27840.0 ;
      RECT  46995.0 26257.5 47060.0 26322.5 ;
      RECT  47027.5 26257.5 47290.0 26322.5 ;
      RECT  46995.0 26290.0 47060.0 26565.0 ;
      RECT  46995.0 26497.5 47060.0 26632.5 ;
      RECT  47185.0 26497.5 47250.0 26632.5 ;
      RECT  47185.0 26497.5 47250.0 26632.5 ;
      RECT  46995.0 26497.5 47060.0 26632.5 ;
      RECT  46995.0 27357.5 47060.0 27492.5 ;
      RECT  47185.0 27357.5 47250.0 27492.5 ;
      RECT  47185.0 27357.5 47250.0 27492.5 ;
      RECT  46995.0 27357.5 47060.0 27492.5 ;
      RECT  46922.5 27772.5 46987.5 27907.5 ;
      RECT  47257.5 26222.5 47322.5 26357.5 ;
      RECT  46995.0 27357.5 47060.0 27492.5 ;
      RECT  47185.0 26497.5 47250.0 26632.5 ;
      RECT  47442.5 26397.5 47507.5 26532.5 ;
      RECT  47442.5 26397.5 47507.5 26532.5 ;
      RECT  47890.0 27807.5 47955.0 27872.5 ;
      RECT  47625.0 27807.5 47922.5 27872.5 ;
      RECT  47890.0 27425.0 47955.0 27840.0 ;
      RECT  47700.0 26257.5 47765.0 26322.5 ;
      RECT  47732.5 26257.5 47995.0 26322.5 ;
      RECT  47700.0 26290.0 47765.0 26565.0 ;
      RECT  47700.0 26497.5 47765.0 26632.5 ;
      RECT  47890.0 26497.5 47955.0 26632.5 ;
      RECT  47890.0 26497.5 47955.0 26632.5 ;
      RECT  47700.0 26497.5 47765.0 26632.5 ;
      RECT  47700.0 27357.5 47765.0 27492.5 ;
      RECT  47890.0 27357.5 47955.0 27492.5 ;
      RECT  47890.0 27357.5 47955.0 27492.5 ;
      RECT  47700.0 27357.5 47765.0 27492.5 ;
      RECT  47627.5 27772.5 47692.5 27907.5 ;
      RECT  47962.5 26222.5 48027.5 26357.5 ;
      RECT  47700.0 27357.5 47765.0 27492.5 ;
      RECT  47890.0 26497.5 47955.0 26632.5 ;
      RECT  48147.5 26397.5 48212.5 26532.5 ;
      RECT  48147.5 26397.5 48212.5 26532.5 ;
      RECT  48595.0 27807.5 48660.0 27872.5 ;
      RECT  48330.0 27807.5 48627.5 27872.5 ;
      RECT  48595.0 27425.0 48660.0 27840.0 ;
      RECT  48405.0 26257.5 48470.0 26322.5 ;
      RECT  48437.5 26257.5 48700.0 26322.5 ;
      RECT  48405.0 26290.0 48470.0 26565.0 ;
      RECT  48405.0 26497.5 48470.0 26632.5 ;
      RECT  48595.0 26497.5 48660.0 26632.5 ;
      RECT  48595.0 26497.5 48660.0 26632.5 ;
      RECT  48405.0 26497.5 48470.0 26632.5 ;
      RECT  48405.0 27357.5 48470.0 27492.5 ;
      RECT  48595.0 27357.5 48660.0 27492.5 ;
      RECT  48595.0 27357.5 48660.0 27492.5 ;
      RECT  48405.0 27357.5 48470.0 27492.5 ;
      RECT  48332.5 27772.5 48397.5 27907.5 ;
      RECT  48667.5 26222.5 48732.5 26357.5 ;
      RECT  48405.0 27357.5 48470.0 27492.5 ;
      RECT  48595.0 26497.5 48660.0 26632.5 ;
      RECT  48852.5 26397.5 48917.5 26532.5 ;
      RECT  48852.5 26397.5 48917.5 26532.5 ;
      RECT  49300.0 27807.5 49365.0 27872.5 ;
      RECT  49035.0 27807.5 49332.5 27872.5 ;
      RECT  49300.0 27425.0 49365.0 27840.0 ;
      RECT  49110.0 26257.5 49175.0 26322.5 ;
      RECT  49142.5 26257.5 49405.0 26322.5 ;
      RECT  49110.0 26290.0 49175.0 26565.0 ;
      RECT  49110.0 26497.5 49175.0 26632.5 ;
      RECT  49300.0 26497.5 49365.0 26632.5 ;
      RECT  49300.0 26497.5 49365.0 26632.5 ;
      RECT  49110.0 26497.5 49175.0 26632.5 ;
      RECT  49110.0 27357.5 49175.0 27492.5 ;
      RECT  49300.0 27357.5 49365.0 27492.5 ;
      RECT  49300.0 27357.5 49365.0 27492.5 ;
      RECT  49110.0 27357.5 49175.0 27492.5 ;
      RECT  49037.5 27772.5 49102.5 27907.5 ;
      RECT  49372.5 26222.5 49437.5 26357.5 ;
      RECT  49110.0 27357.5 49175.0 27492.5 ;
      RECT  49300.0 26497.5 49365.0 26632.5 ;
      RECT  49557.5 26397.5 49622.5 26532.5 ;
      RECT  49557.5 26397.5 49622.5 26532.5 ;
      RECT  50005.0 27807.5 50070.0 27872.5 ;
      RECT  49740.0 27807.5 50037.5 27872.5 ;
      RECT  50005.0 27425.0 50070.0 27840.0 ;
      RECT  49815.0 26257.5 49880.0 26322.5 ;
      RECT  49847.5 26257.5 50110.0 26322.5 ;
      RECT  49815.0 26290.0 49880.0 26565.0 ;
      RECT  49815.0 26497.5 49880.0 26632.5 ;
      RECT  50005.0 26497.5 50070.0 26632.5 ;
      RECT  50005.0 26497.5 50070.0 26632.5 ;
      RECT  49815.0 26497.5 49880.0 26632.5 ;
      RECT  49815.0 27357.5 49880.0 27492.5 ;
      RECT  50005.0 27357.5 50070.0 27492.5 ;
      RECT  50005.0 27357.5 50070.0 27492.5 ;
      RECT  49815.0 27357.5 49880.0 27492.5 ;
      RECT  49742.5 27772.5 49807.5 27907.5 ;
      RECT  50077.5 26222.5 50142.5 26357.5 ;
      RECT  49815.0 27357.5 49880.0 27492.5 ;
      RECT  50005.0 26497.5 50070.0 26632.5 ;
      RECT  50262.5 26397.5 50327.5 26532.5 ;
      RECT  50262.5 26397.5 50327.5 26532.5 ;
      RECT  50710.0 27807.5 50775.0 27872.5 ;
      RECT  50445.0 27807.5 50742.5 27872.5 ;
      RECT  50710.0 27425.0 50775.0 27840.0 ;
      RECT  50520.0 26257.5 50585.0 26322.5 ;
      RECT  50552.5 26257.5 50815.0 26322.5 ;
      RECT  50520.0 26290.0 50585.0 26565.0 ;
      RECT  50520.0 26497.5 50585.0 26632.5 ;
      RECT  50710.0 26497.5 50775.0 26632.5 ;
      RECT  50710.0 26497.5 50775.0 26632.5 ;
      RECT  50520.0 26497.5 50585.0 26632.5 ;
      RECT  50520.0 27357.5 50585.0 27492.5 ;
      RECT  50710.0 27357.5 50775.0 27492.5 ;
      RECT  50710.0 27357.5 50775.0 27492.5 ;
      RECT  50520.0 27357.5 50585.0 27492.5 ;
      RECT  50447.5 27772.5 50512.5 27907.5 ;
      RECT  50782.5 26222.5 50847.5 26357.5 ;
      RECT  50520.0 27357.5 50585.0 27492.5 ;
      RECT  50710.0 26497.5 50775.0 26632.5 ;
      RECT  50967.5 26397.5 51032.5 26532.5 ;
      RECT  50967.5 26397.5 51032.5 26532.5 ;
      RECT  51415.0 27807.5 51480.0 27872.5 ;
      RECT  51150.0 27807.5 51447.5 27872.5 ;
      RECT  51415.0 27425.0 51480.0 27840.0 ;
      RECT  51225.0 26257.5 51290.0 26322.5 ;
      RECT  51257.5 26257.5 51520.0 26322.5 ;
      RECT  51225.0 26290.0 51290.0 26565.0 ;
      RECT  51225.0 26497.5 51290.0 26632.5 ;
      RECT  51415.0 26497.5 51480.0 26632.5 ;
      RECT  51415.0 26497.5 51480.0 26632.5 ;
      RECT  51225.0 26497.5 51290.0 26632.5 ;
      RECT  51225.0 27357.5 51290.0 27492.5 ;
      RECT  51415.0 27357.5 51480.0 27492.5 ;
      RECT  51415.0 27357.5 51480.0 27492.5 ;
      RECT  51225.0 27357.5 51290.0 27492.5 ;
      RECT  51152.5 27772.5 51217.5 27907.5 ;
      RECT  51487.5 26222.5 51552.5 26357.5 ;
      RECT  51225.0 27357.5 51290.0 27492.5 ;
      RECT  51415.0 26497.5 51480.0 26632.5 ;
      RECT  51672.5 26397.5 51737.5 26532.5 ;
      RECT  51672.5 26397.5 51737.5 26532.5 ;
      RECT  52120.0 27807.5 52185.0 27872.5 ;
      RECT  51855.0 27807.5 52152.5 27872.5 ;
      RECT  52120.0 27425.0 52185.0 27840.0 ;
      RECT  51930.0 26257.5 51995.0 26322.5 ;
      RECT  51962.5 26257.5 52225.0 26322.5 ;
      RECT  51930.0 26290.0 51995.0 26565.0 ;
      RECT  51930.0 26497.5 51995.0 26632.5 ;
      RECT  52120.0 26497.5 52185.0 26632.5 ;
      RECT  52120.0 26497.5 52185.0 26632.5 ;
      RECT  51930.0 26497.5 51995.0 26632.5 ;
      RECT  51930.0 27357.5 51995.0 27492.5 ;
      RECT  52120.0 27357.5 52185.0 27492.5 ;
      RECT  52120.0 27357.5 52185.0 27492.5 ;
      RECT  51930.0 27357.5 51995.0 27492.5 ;
      RECT  51857.5 27772.5 51922.5 27907.5 ;
      RECT  52192.5 26222.5 52257.5 26357.5 ;
      RECT  51930.0 27357.5 51995.0 27492.5 ;
      RECT  52120.0 26497.5 52185.0 26632.5 ;
      RECT  52377.5 26397.5 52442.5 26532.5 ;
      RECT  52377.5 26397.5 52442.5 26532.5 ;
      RECT  52825.0 27807.5 52890.0 27872.5 ;
      RECT  52560.0 27807.5 52857.5 27872.5 ;
      RECT  52825.0 27425.0 52890.0 27840.0 ;
      RECT  52635.0 26257.5 52700.0 26322.5 ;
      RECT  52667.5 26257.5 52930.0 26322.5 ;
      RECT  52635.0 26290.0 52700.0 26565.0 ;
      RECT  52635.0 26497.5 52700.0 26632.5 ;
      RECT  52825.0 26497.5 52890.0 26632.5 ;
      RECT  52825.0 26497.5 52890.0 26632.5 ;
      RECT  52635.0 26497.5 52700.0 26632.5 ;
      RECT  52635.0 27357.5 52700.0 27492.5 ;
      RECT  52825.0 27357.5 52890.0 27492.5 ;
      RECT  52825.0 27357.5 52890.0 27492.5 ;
      RECT  52635.0 27357.5 52700.0 27492.5 ;
      RECT  52562.5 27772.5 52627.5 27907.5 ;
      RECT  52897.5 26222.5 52962.5 26357.5 ;
      RECT  52635.0 27357.5 52700.0 27492.5 ;
      RECT  52825.0 26497.5 52890.0 26632.5 ;
      RECT  53082.5 26397.5 53147.5 26532.5 ;
      RECT  53082.5 26397.5 53147.5 26532.5 ;
      RECT  53530.0 27807.5 53595.0 27872.5 ;
      RECT  53265.0 27807.5 53562.5 27872.5 ;
      RECT  53530.0 27425.0 53595.0 27840.0 ;
      RECT  53340.0 26257.5 53405.0 26322.5 ;
      RECT  53372.5 26257.5 53635.0 26322.5 ;
      RECT  53340.0 26290.0 53405.0 26565.0 ;
      RECT  53340.0 26497.5 53405.0 26632.5 ;
      RECT  53530.0 26497.5 53595.0 26632.5 ;
      RECT  53530.0 26497.5 53595.0 26632.5 ;
      RECT  53340.0 26497.5 53405.0 26632.5 ;
      RECT  53340.0 27357.5 53405.0 27492.5 ;
      RECT  53530.0 27357.5 53595.0 27492.5 ;
      RECT  53530.0 27357.5 53595.0 27492.5 ;
      RECT  53340.0 27357.5 53405.0 27492.5 ;
      RECT  53267.5 27772.5 53332.5 27907.5 ;
      RECT  53602.5 26222.5 53667.5 26357.5 ;
      RECT  53340.0 27357.5 53405.0 27492.5 ;
      RECT  53530.0 26497.5 53595.0 26632.5 ;
      RECT  53787.5 26397.5 53852.5 26532.5 ;
      RECT  53787.5 26397.5 53852.5 26532.5 ;
      RECT  54235.0 27807.5 54300.0 27872.5 ;
      RECT  53970.0 27807.5 54267.5 27872.5 ;
      RECT  54235.0 27425.0 54300.0 27840.0 ;
      RECT  54045.0 26257.5 54110.0 26322.5 ;
      RECT  54077.5 26257.5 54340.0 26322.5 ;
      RECT  54045.0 26290.0 54110.0 26565.0 ;
      RECT  54045.0 26497.5 54110.0 26632.5 ;
      RECT  54235.0 26497.5 54300.0 26632.5 ;
      RECT  54235.0 26497.5 54300.0 26632.5 ;
      RECT  54045.0 26497.5 54110.0 26632.5 ;
      RECT  54045.0 27357.5 54110.0 27492.5 ;
      RECT  54235.0 27357.5 54300.0 27492.5 ;
      RECT  54235.0 27357.5 54300.0 27492.5 ;
      RECT  54045.0 27357.5 54110.0 27492.5 ;
      RECT  53972.5 27772.5 54037.5 27907.5 ;
      RECT  54307.5 26222.5 54372.5 26357.5 ;
      RECT  54045.0 27357.5 54110.0 27492.5 ;
      RECT  54235.0 26497.5 54300.0 26632.5 ;
      RECT  54492.5 26397.5 54557.5 26532.5 ;
      RECT  54492.5 26397.5 54557.5 26532.5 ;
      RECT  54940.0 27807.5 55005.0 27872.5 ;
      RECT  54675.0 27807.5 54972.5 27872.5 ;
      RECT  54940.0 27425.0 55005.0 27840.0 ;
      RECT  54750.0 26257.5 54815.0 26322.5 ;
      RECT  54782.5 26257.5 55045.0 26322.5 ;
      RECT  54750.0 26290.0 54815.0 26565.0 ;
      RECT  54750.0 26497.5 54815.0 26632.5 ;
      RECT  54940.0 26497.5 55005.0 26632.5 ;
      RECT  54940.0 26497.5 55005.0 26632.5 ;
      RECT  54750.0 26497.5 54815.0 26632.5 ;
      RECT  54750.0 27357.5 54815.0 27492.5 ;
      RECT  54940.0 27357.5 55005.0 27492.5 ;
      RECT  54940.0 27357.5 55005.0 27492.5 ;
      RECT  54750.0 27357.5 54815.0 27492.5 ;
      RECT  54677.5 27772.5 54742.5 27907.5 ;
      RECT  55012.5 26222.5 55077.5 26357.5 ;
      RECT  54750.0 27357.5 54815.0 27492.5 ;
      RECT  54940.0 26497.5 55005.0 26632.5 ;
      RECT  55197.5 26397.5 55262.5 26532.5 ;
      RECT  55197.5 26397.5 55262.5 26532.5 ;
      RECT  55645.0 27807.5 55710.0 27872.5 ;
      RECT  55380.0 27807.5 55677.5 27872.5 ;
      RECT  55645.0 27425.0 55710.0 27840.0 ;
      RECT  55455.0 26257.5 55520.0 26322.5 ;
      RECT  55487.5 26257.5 55750.0 26322.5 ;
      RECT  55455.0 26290.0 55520.0 26565.0 ;
      RECT  55455.0 26497.5 55520.0 26632.5 ;
      RECT  55645.0 26497.5 55710.0 26632.5 ;
      RECT  55645.0 26497.5 55710.0 26632.5 ;
      RECT  55455.0 26497.5 55520.0 26632.5 ;
      RECT  55455.0 27357.5 55520.0 27492.5 ;
      RECT  55645.0 27357.5 55710.0 27492.5 ;
      RECT  55645.0 27357.5 55710.0 27492.5 ;
      RECT  55455.0 27357.5 55520.0 27492.5 ;
      RECT  55382.5 27772.5 55447.5 27907.5 ;
      RECT  55717.5 26222.5 55782.5 26357.5 ;
      RECT  55455.0 27357.5 55520.0 27492.5 ;
      RECT  55645.0 26497.5 55710.0 26632.5 ;
      RECT  55902.5 26397.5 55967.5 26532.5 ;
      RECT  55902.5 26397.5 55967.5 26532.5 ;
      RECT  56350.0 27807.5 56415.0 27872.5 ;
      RECT  56085.0 27807.5 56382.5 27872.5 ;
      RECT  56350.0 27425.0 56415.0 27840.0 ;
      RECT  56160.0 26257.5 56225.0 26322.5 ;
      RECT  56192.5 26257.5 56455.0 26322.5 ;
      RECT  56160.0 26290.0 56225.0 26565.0 ;
      RECT  56160.0 26497.5 56225.0 26632.5 ;
      RECT  56350.0 26497.5 56415.0 26632.5 ;
      RECT  56350.0 26497.5 56415.0 26632.5 ;
      RECT  56160.0 26497.5 56225.0 26632.5 ;
      RECT  56160.0 27357.5 56225.0 27492.5 ;
      RECT  56350.0 27357.5 56415.0 27492.5 ;
      RECT  56350.0 27357.5 56415.0 27492.5 ;
      RECT  56160.0 27357.5 56225.0 27492.5 ;
      RECT  56087.5 27772.5 56152.5 27907.5 ;
      RECT  56422.5 26222.5 56487.5 26357.5 ;
      RECT  56160.0 27357.5 56225.0 27492.5 ;
      RECT  56350.0 26497.5 56415.0 26632.5 ;
      RECT  56607.5 26397.5 56672.5 26532.5 ;
      RECT  56607.5 26397.5 56672.5 26532.5 ;
      RECT  57055.0 27807.5 57120.0 27872.5 ;
      RECT  56790.0 27807.5 57087.5 27872.5 ;
      RECT  57055.0 27425.0 57120.0 27840.0 ;
      RECT  56865.0 26257.5 56930.0 26322.5 ;
      RECT  56897.5 26257.5 57160.0 26322.5 ;
      RECT  56865.0 26290.0 56930.0 26565.0 ;
      RECT  56865.0 26497.5 56930.0 26632.5 ;
      RECT  57055.0 26497.5 57120.0 26632.5 ;
      RECT  57055.0 26497.5 57120.0 26632.5 ;
      RECT  56865.0 26497.5 56930.0 26632.5 ;
      RECT  56865.0 27357.5 56930.0 27492.5 ;
      RECT  57055.0 27357.5 57120.0 27492.5 ;
      RECT  57055.0 27357.5 57120.0 27492.5 ;
      RECT  56865.0 27357.5 56930.0 27492.5 ;
      RECT  56792.5 27772.5 56857.5 27907.5 ;
      RECT  57127.5 26222.5 57192.5 26357.5 ;
      RECT  56865.0 27357.5 56930.0 27492.5 ;
      RECT  57055.0 26497.5 57120.0 26632.5 ;
      RECT  57312.5 26397.5 57377.5 26532.5 ;
      RECT  57312.5 26397.5 57377.5 26532.5 ;
      RECT  57760.0 27807.5 57825.0 27872.5 ;
      RECT  57495.0 27807.5 57792.5 27872.5 ;
      RECT  57760.0 27425.0 57825.0 27840.0 ;
      RECT  57570.0 26257.5 57635.0 26322.5 ;
      RECT  57602.5 26257.5 57865.0 26322.5 ;
      RECT  57570.0 26290.0 57635.0 26565.0 ;
      RECT  57570.0 26497.5 57635.0 26632.5 ;
      RECT  57760.0 26497.5 57825.0 26632.5 ;
      RECT  57760.0 26497.5 57825.0 26632.5 ;
      RECT  57570.0 26497.5 57635.0 26632.5 ;
      RECT  57570.0 27357.5 57635.0 27492.5 ;
      RECT  57760.0 27357.5 57825.0 27492.5 ;
      RECT  57760.0 27357.5 57825.0 27492.5 ;
      RECT  57570.0 27357.5 57635.0 27492.5 ;
      RECT  57497.5 27772.5 57562.5 27907.5 ;
      RECT  57832.5 26222.5 57897.5 26357.5 ;
      RECT  57570.0 27357.5 57635.0 27492.5 ;
      RECT  57760.0 26497.5 57825.0 26632.5 ;
      RECT  58017.5 26397.5 58082.5 26532.5 ;
      RECT  58017.5 26397.5 58082.5 26532.5 ;
      RECT  58465.0 27807.5 58530.0 27872.5 ;
      RECT  58200.0 27807.5 58497.5 27872.5 ;
      RECT  58465.0 27425.0 58530.0 27840.0 ;
      RECT  58275.0 26257.5 58340.0 26322.5 ;
      RECT  58307.5 26257.5 58570.0 26322.5 ;
      RECT  58275.0 26290.0 58340.0 26565.0 ;
      RECT  58275.0 26497.5 58340.0 26632.5 ;
      RECT  58465.0 26497.5 58530.0 26632.5 ;
      RECT  58465.0 26497.5 58530.0 26632.5 ;
      RECT  58275.0 26497.5 58340.0 26632.5 ;
      RECT  58275.0 27357.5 58340.0 27492.5 ;
      RECT  58465.0 27357.5 58530.0 27492.5 ;
      RECT  58465.0 27357.5 58530.0 27492.5 ;
      RECT  58275.0 27357.5 58340.0 27492.5 ;
      RECT  58202.5 27772.5 58267.5 27907.5 ;
      RECT  58537.5 26222.5 58602.5 26357.5 ;
      RECT  58275.0 27357.5 58340.0 27492.5 ;
      RECT  58465.0 26497.5 58530.0 26632.5 ;
      RECT  58722.5 26397.5 58787.5 26532.5 ;
      RECT  58722.5 26397.5 58787.5 26532.5 ;
      RECT  59170.0 27807.5 59235.0 27872.5 ;
      RECT  58905.0 27807.5 59202.5 27872.5 ;
      RECT  59170.0 27425.0 59235.0 27840.0 ;
      RECT  58980.0 26257.5 59045.0 26322.5 ;
      RECT  59012.5 26257.5 59275.0 26322.5 ;
      RECT  58980.0 26290.0 59045.0 26565.0 ;
      RECT  58980.0 26497.5 59045.0 26632.5 ;
      RECT  59170.0 26497.5 59235.0 26632.5 ;
      RECT  59170.0 26497.5 59235.0 26632.5 ;
      RECT  58980.0 26497.5 59045.0 26632.5 ;
      RECT  58980.0 27357.5 59045.0 27492.5 ;
      RECT  59170.0 27357.5 59235.0 27492.5 ;
      RECT  59170.0 27357.5 59235.0 27492.5 ;
      RECT  58980.0 27357.5 59045.0 27492.5 ;
      RECT  58907.5 27772.5 58972.5 27907.5 ;
      RECT  59242.5 26222.5 59307.5 26357.5 ;
      RECT  58980.0 27357.5 59045.0 27492.5 ;
      RECT  59170.0 26497.5 59235.0 26632.5 ;
      RECT  59427.5 26397.5 59492.5 26532.5 ;
      RECT  59427.5 26397.5 59492.5 26532.5 ;
      RECT  59875.0 27807.5 59940.0 27872.5 ;
      RECT  59610.0 27807.5 59907.5 27872.5 ;
      RECT  59875.0 27425.0 59940.0 27840.0 ;
      RECT  59685.0 26257.5 59750.0 26322.5 ;
      RECT  59717.5 26257.5 59980.0 26322.5 ;
      RECT  59685.0 26290.0 59750.0 26565.0 ;
      RECT  59685.0 26497.5 59750.0 26632.5 ;
      RECT  59875.0 26497.5 59940.0 26632.5 ;
      RECT  59875.0 26497.5 59940.0 26632.5 ;
      RECT  59685.0 26497.5 59750.0 26632.5 ;
      RECT  59685.0 27357.5 59750.0 27492.5 ;
      RECT  59875.0 27357.5 59940.0 27492.5 ;
      RECT  59875.0 27357.5 59940.0 27492.5 ;
      RECT  59685.0 27357.5 59750.0 27492.5 ;
      RECT  59612.5 27772.5 59677.5 27907.5 ;
      RECT  59947.5 26222.5 60012.5 26357.5 ;
      RECT  59685.0 27357.5 59750.0 27492.5 ;
      RECT  59875.0 26497.5 59940.0 26632.5 ;
      RECT  60132.5 26397.5 60197.5 26532.5 ;
      RECT  60132.5 26397.5 60197.5 26532.5 ;
      RECT  60580.0 27807.5 60645.0 27872.5 ;
      RECT  60315.0 27807.5 60612.5 27872.5 ;
      RECT  60580.0 27425.0 60645.0 27840.0 ;
      RECT  60390.0 26257.5 60455.0 26322.5 ;
      RECT  60422.5 26257.5 60685.0 26322.5 ;
      RECT  60390.0 26290.0 60455.0 26565.0 ;
      RECT  60390.0 26497.5 60455.0 26632.5 ;
      RECT  60580.0 26497.5 60645.0 26632.5 ;
      RECT  60580.0 26497.5 60645.0 26632.5 ;
      RECT  60390.0 26497.5 60455.0 26632.5 ;
      RECT  60390.0 27357.5 60455.0 27492.5 ;
      RECT  60580.0 27357.5 60645.0 27492.5 ;
      RECT  60580.0 27357.5 60645.0 27492.5 ;
      RECT  60390.0 27357.5 60455.0 27492.5 ;
      RECT  60317.5 27772.5 60382.5 27907.5 ;
      RECT  60652.5 26222.5 60717.5 26357.5 ;
      RECT  60390.0 27357.5 60455.0 27492.5 ;
      RECT  60580.0 26497.5 60645.0 26632.5 ;
      RECT  60837.5 26397.5 60902.5 26532.5 ;
      RECT  60837.5 26397.5 60902.5 26532.5 ;
      RECT  61285.0 27807.5 61350.0 27872.5 ;
      RECT  61020.0 27807.5 61317.5 27872.5 ;
      RECT  61285.0 27425.0 61350.0 27840.0 ;
      RECT  61095.0 26257.5 61160.0 26322.5 ;
      RECT  61127.5 26257.5 61390.0 26322.5 ;
      RECT  61095.0 26290.0 61160.0 26565.0 ;
      RECT  61095.0 26497.5 61160.0 26632.5 ;
      RECT  61285.0 26497.5 61350.0 26632.5 ;
      RECT  61285.0 26497.5 61350.0 26632.5 ;
      RECT  61095.0 26497.5 61160.0 26632.5 ;
      RECT  61095.0 27357.5 61160.0 27492.5 ;
      RECT  61285.0 27357.5 61350.0 27492.5 ;
      RECT  61285.0 27357.5 61350.0 27492.5 ;
      RECT  61095.0 27357.5 61160.0 27492.5 ;
      RECT  61022.5 27772.5 61087.5 27907.5 ;
      RECT  61357.5 26222.5 61422.5 26357.5 ;
      RECT  61095.0 27357.5 61160.0 27492.5 ;
      RECT  61285.0 26497.5 61350.0 26632.5 ;
      RECT  61542.5 26397.5 61607.5 26532.5 ;
      RECT  61542.5 26397.5 61607.5 26532.5 ;
      RECT  61990.0 27807.5 62055.0 27872.5 ;
      RECT  61725.0 27807.5 62022.5 27872.5 ;
      RECT  61990.0 27425.0 62055.0 27840.0 ;
      RECT  61800.0 26257.5 61865.0 26322.5 ;
      RECT  61832.5 26257.5 62095.0 26322.5 ;
      RECT  61800.0 26290.0 61865.0 26565.0 ;
      RECT  61800.0 26497.5 61865.0 26632.5 ;
      RECT  61990.0 26497.5 62055.0 26632.5 ;
      RECT  61990.0 26497.5 62055.0 26632.5 ;
      RECT  61800.0 26497.5 61865.0 26632.5 ;
      RECT  61800.0 27357.5 61865.0 27492.5 ;
      RECT  61990.0 27357.5 62055.0 27492.5 ;
      RECT  61990.0 27357.5 62055.0 27492.5 ;
      RECT  61800.0 27357.5 61865.0 27492.5 ;
      RECT  61727.5 27772.5 61792.5 27907.5 ;
      RECT  62062.5 26222.5 62127.5 26357.5 ;
      RECT  61800.0 27357.5 61865.0 27492.5 ;
      RECT  61990.0 26497.5 62055.0 26632.5 ;
      RECT  62247.5 26397.5 62312.5 26532.5 ;
      RECT  62247.5 26397.5 62312.5 26532.5 ;
      RECT  62695.0 27807.5 62760.0 27872.5 ;
      RECT  62430.0 27807.5 62727.5 27872.5 ;
      RECT  62695.0 27425.0 62760.0 27840.0 ;
      RECT  62505.0 26257.5 62570.0 26322.5 ;
      RECT  62537.5 26257.5 62800.0 26322.5 ;
      RECT  62505.0 26290.0 62570.0 26565.0 ;
      RECT  62505.0 26497.5 62570.0 26632.5 ;
      RECT  62695.0 26497.5 62760.0 26632.5 ;
      RECT  62695.0 26497.5 62760.0 26632.5 ;
      RECT  62505.0 26497.5 62570.0 26632.5 ;
      RECT  62505.0 27357.5 62570.0 27492.5 ;
      RECT  62695.0 27357.5 62760.0 27492.5 ;
      RECT  62695.0 27357.5 62760.0 27492.5 ;
      RECT  62505.0 27357.5 62570.0 27492.5 ;
      RECT  62432.5 27772.5 62497.5 27907.5 ;
      RECT  62767.5 26222.5 62832.5 26357.5 ;
      RECT  62505.0 27357.5 62570.0 27492.5 ;
      RECT  62695.0 26497.5 62760.0 26632.5 ;
      RECT  62952.5 26397.5 63017.5 26532.5 ;
      RECT  62952.5 26397.5 63017.5 26532.5 ;
      RECT  63400.0 27807.5 63465.0 27872.5 ;
      RECT  63135.0 27807.5 63432.5 27872.5 ;
      RECT  63400.0 27425.0 63465.0 27840.0 ;
      RECT  63210.0 26257.5 63275.0 26322.5 ;
      RECT  63242.5 26257.5 63505.0 26322.5 ;
      RECT  63210.0 26290.0 63275.0 26565.0 ;
      RECT  63210.0 26497.5 63275.0 26632.5 ;
      RECT  63400.0 26497.5 63465.0 26632.5 ;
      RECT  63400.0 26497.5 63465.0 26632.5 ;
      RECT  63210.0 26497.5 63275.0 26632.5 ;
      RECT  63210.0 27357.5 63275.0 27492.5 ;
      RECT  63400.0 27357.5 63465.0 27492.5 ;
      RECT  63400.0 27357.5 63465.0 27492.5 ;
      RECT  63210.0 27357.5 63275.0 27492.5 ;
      RECT  63137.5 27772.5 63202.5 27907.5 ;
      RECT  63472.5 26222.5 63537.5 26357.5 ;
      RECT  63210.0 27357.5 63275.0 27492.5 ;
      RECT  63400.0 26497.5 63465.0 26632.5 ;
      RECT  63657.5 26397.5 63722.5 26532.5 ;
      RECT  63657.5 26397.5 63722.5 26532.5 ;
      RECT  64105.0 27807.5 64170.0 27872.5 ;
      RECT  63840.0 27807.5 64137.5 27872.5 ;
      RECT  64105.0 27425.0 64170.0 27840.0 ;
      RECT  63915.0 26257.5 63980.0 26322.5 ;
      RECT  63947.5 26257.5 64210.0 26322.5 ;
      RECT  63915.0 26290.0 63980.0 26565.0 ;
      RECT  63915.0 26497.5 63980.0 26632.5 ;
      RECT  64105.0 26497.5 64170.0 26632.5 ;
      RECT  64105.0 26497.5 64170.0 26632.5 ;
      RECT  63915.0 26497.5 63980.0 26632.5 ;
      RECT  63915.0 27357.5 63980.0 27492.5 ;
      RECT  64105.0 27357.5 64170.0 27492.5 ;
      RECT  64105.0 27357.5 64170.0 27492.5 ;
      RECT  63915.0 27357.5 63980.0 27492.5 ;
      RECT  63842.5 27772.5 63907.5 27907.5 ;
      RECT  64177.5 26222.5 64242.5 26357.5 ;
      RECT  63915.0 27357.5 63980.0 27492.5 ;
      RECT  64105.0 26497.5 64170.0 26632.5 ;
      RECT  64362.5 26397.5 64427.5 26532.5 ;
      RECT  64362.5 26397.5 64427.5 26532.5 ;
      RECT  64810.0 27807.5 64875.0 27872.5 ;
      RECT  64545.0 27807.5 64842.5 27872.5 ;
      RECT  64810.0 27425.0 64875.0 27840.0 ;
      RECT  64620.0 26257.5 64685.0 26322.5 ;
      RECT  64652.5 26257.5 64915.0 26322.5 ;
      RECT  64620.0 26290.0 64685.0 26565.0 ;
      RECT  64620.0 26497.5 64685.0 26632.5 ;
      RECT  64810.0 26497.5 64875.0 26632.5 ;
      RECT  64810.0 26497.5 64875.0 26632.5 ;
      RECT  64620.0 26497.5 64685.0 26632.5 ;
      RECT  64620.0 27357.5 64685.0 27492.5 ;
      RECT  64810.0 27357.5 64875.0 27492.5 ;
      RECT  64810.0 27357.5 64875.0 27492.5 ;
      RECT  64620.0 27357.5 64685.0 27492.5 ;
      RECT  64547.5 27772.5 64612.5 27907.5 ;
      RECT  64882.5 26222.5 64947.5 26357.5 ;
      RECT  64620.0 27357.5 64685.0 27492.5 ;
      RECT  64810.0 26497.5 64875.0 26632.5 ;
      RECT  65067.5 26397.5 65132.5 26532.5 ;
      RECT  65067.5 26397.5 65132.5 26532.5 ;
      RECT  65515.0 27807.5 65580.0 27872.5 ;
      RECT  65250.0 27807.5 65547.5 27872.5 ;
      RECT  65515.0 27425.0 65580.0 27840.0 ;
      RECT  65325.0 26257.5 65390.0 26322.5 ;
      RECT  65357.5 26257.5 65620.0 26322.5 ;
      RECT  65325.0 26290.0 65390.0 26565.0 ;
      RECT  65325.0 26497.5 65390.0 26632.5 ;
      RECT  65515.0 26497.5 65580.0 26632.5 ;
      RECT  65515.0 26497.5 65580.0 26632.5 ;
      RECT  65325.0 26497.5 65390.0 26632.5 ;
      RECT  65325.0 27357.5 65390.0 27492.5 ;
      RECT  65515.0 27357.5 65580.0 27492.5 ;
      RECT  65515.0 27357.5 65580.0 27492.5 ;
      RECT  65325.0 27357.5 65390.0 27492.5 ;
      RECT  65252.5 27772.5 65317.5 27907.5 ;
      RECT  65587.5 26222.5 65652.5 26357.5 ;
      RECT  65325.0 27357.5 65390.0 27492.5 ;
      RECT  65515.0 26497.5 65580.0 26632.5 ;
      RECT  65772.5 26397.5 65837.5 26532.5 ;
      RECT  65772.5 26397.5 65837.5 26532.5 ;
      RECT  66220.0 27807.5 66285.0 27872.5 ;
      RECT  65955.0 27807.5 66252.5 27872.5 ;
      RECT  66220.0 27425.0 66285.0 27840.0 ;
      RECT  66030.0 26257.5 66095.0 26322.5 ;
      RECT  66062.5 26257.5 66325.0 26322.5 ;
      RECT  66030.0 26290.0 66095.0 26565.0 ;
      RECT  66030.0 26497.5 66095.0 26632.5 ;
      RECT  66220.0 26497.5 66285.0 26632.5 ;
      RECT  66220.0 26497.5 66285.0 26632.5 ;
      RECT  66030.0 26497.5 66095.0 26632.5 ;
      RECT  66030.0 27357.5 66095.0 27492.5 ;
      RECT  66220.0 27357.5 66285.0 27492.5 ;
      RECT  66220.0 27357.5 66285.0 27492.5 ;
      RECT  66030.0 27357.5 66095.0 27492.5 ;
      RECT  65957.5 27772.5 66022.5 27907.5 ;
      RECT  66292.5 26222.5 66357.5 26357.5 ;
      RECT  66030.0 27357.5 66095.0 27492.5 ;
      RECT  66220.0 26497.5 66285.0 26632.5 ;
      RECT  66477.5 26397.5 66542.5 26532.5 ;
      RECT  66477.5 26397.5 66542.5 26532.5 ;
      RECT  66925.0 27807.5 66990.0 27872.5 ;
      RECT  66660.0 27807.5 66957.5 27872.5 ;
      RECT  66925.0 27425.0 66990.0 27840.0 ;
      RECT  66735.0 26257.5 66800.0 26322.5 ;
      RECT  66767.5 26257.5 67030.0 26322.5 ;
      RECT  66735.0 26290.0 66800.0 26565.0 ;
      RECT  66735.0 26497.5 66800.0 26632.5 ;
      RECT  66925.0 26497.5 66990.0 26632.5 ;
      RECT  66925.0 26497.5 66990.0 26632.5 ;
      RECT  66735.0 26497.5 66800.0 26632.5 ;
      RECT  66735.0 27357.5 66800.0 27492.5 ;
      RECT  66925.0 27357.5 66990.0 27492.5 ;
      RECT  66925.0 27357.5 66990.0 27492.5 ;
      RECT  66735.0 27357.5 66800.0 27492.5 ;
      RECT  66662.5 27772.5 66727.5 27907.5 ;
      RECT  66997.5 26222.5 67062.5 26357.5 ;
      RECT  66735.0 27357.5 66800.0 27492.5 ;
      RECT  66925.0 26497.5 66990.0 26632.5 ;
      RECT  67182.5 26397.5 67247.5 26532.5 ;
      RECT  67182.5 26397.5 67247.5 26532.5 ;
      RECT  67630.0 27807.5 67695.0 27872.5 ;
      RECT  67365.0 27807.5 67662.5 27872.5 ;
      RECT  67630.0 27425.0 67695.0 27840.0 ;
      RECT  67440.0 26257.5 67505.0 26322.5 ;
      RECT  67472.5 26257.5 67735.0 26322.5 ;
      RECT  67440.0 26290.0 67505.0 26565.0 ;
      RECT  67440.0 26497.5 67505.0 26632.5 ;
      RECT  67630.0 26497.5 67695.0 26632.5 ;
      RECT  67630.0 26497.5 67695.0 26632.5 ;
      RECT  67440.0 26497.5 67505.0 26632.5 ;
      RECT  67440.0 27357.5 67505.0 27492.5 ;
      RECT  67630.0 27357.5 67695.0 27492.5 ;
      RECT  67630.0 27357.5 67695.0 27492.5 ;
      RECT  67440.0 27357.5 67505.0 27492.5 ;
      RECT  67367.5 27772.5 67432.5 27907.5 ;
      RECT  67702.5 26222.5 67767.5 26357.5 ;
      RECT  67440.0 27357.5 67505.0 27492.5 ;
      RECT  67630.0 26497.5 67695.0 26632.5 ;
      RECT  67887.5 26397.5 67952.5 26532.5 ;
      RECT  67887.5 26397.5 67952.5 26532.5 ;
      RECT  68335.0 27807.5 68400.0 27872.5 ;
      RECT  68070.0 27807.5 68367.5 27872.5 ;
      RECT  68335.0 27425.0 68400.0 27840.0 ;
      RECT  68145.0 26257.5 68210.0 26322.5 ;
      RECT  68177.5 26257.5 68440.0 26322.5 ;
      RECT  68145.0 26290.0 68210.0 26565.0 ;
      RECT  68145.0 26497.5 68210.0 26632.5 ;
      RECT  68335.0 26497.5 68400.0 26632.5 ;
      RECT  68335.0 26497.5 68400.0 26632.5 ;
      RECT  68145.0 26497.5 68210.0 26632.5 ;
      RECT  68145.0 27357.5 68210.0 27492.5 ;
      RECT  68335.0 27357.5 68400.0 27492.5 ;
      RECT  68335.0 27357.5 68400.0 27492.5 ;
      RECT  68145.0 27357.5 68210.0 27492.5 ;
      RECT  68072.5 27772.5 68137.5 27907.5 ;
      RECT  68407.5 26222.5 68472.5 26357.5 ;
      RECT  68145.0 27357.5 68210.0 27492.5 ;
      RECT  68335.0 26497.5 68400.0 26632.5 ;
      RECT  68592.5 26397.5 68657.5 26532.5 ;
      RECT  68592.5 26397.5 68657.5 26532.5 ;
      RECT  69040.0 27807.5 69105.0 27872.5 ;
      RECT  68775.0 27807.5 69072.5 27872.5 ;
      RECT  69040.0 27425.0 69105.0 27840.0 ;
      RECT  68850.0 26257.5 68915.0 26322.5 ;
      RECT  68882.5 26257.5 69145.0 26322.5 ;
      RECT  68850.0 26290.0 68915.0 26565.0 ;
      RECT  68850.0 26497.5 68915.0 26632.5 ;
      RECT  69040.0 26497.5 69105.0 26632.5 ;
      RECT  69040.0 26497.5 69105.0 26632.5 ;
      RECT  68850.0 26497.5 68915.0 26632.5 ;
      RECT  68850.0 27357.5 68915.0 27492.5 ;
      RECT  69040.0 27357.5 69105.0 27492.5 ;
      RECT  69040.0 27357.5 69105.0 27492.5 ;
      RECT  68850.0 27357.5 68915.0 27492.5 ;
      RECT  68777.5 27772.5 68842.5 27907.5 ;
      RECT  69112.5 26222.5 69177.5 26357.5 ;
      RECT  68850.0 27357.5 68915.0 27492.5 ;
      RECT  69040.0 26497.5 69105.0 26632.5 ;
      RECT  69297.5 26397.5 69362.5 26532.5 ;
      RECT  69297.5 26397.5 69362.5 26532.5 ;
      RECT  69745.0 27807.5 69810.0 27872.5 ;
      RECT  69480.0 27807.5 69777.5 27872.5 ;
      RECT  69745.0 27425.0 69810.0 27840.0 ;
      RECT  69555.0 26257.5 69620.0 26322.5 ;
      RECT  69587.5 26257.5 69850.0 26322.5 ;
      RECT  69555.0 26290.0 69620.0 26565.0 ;
      RECT  69555.0 26497.5 69620.0 26632.5 ;
      RECT  69745.0 26497.5 69810.0 26632.5 ;
      RECT  69745.0 26497.5 69810.0 26632.5 ;
      RECT  69555.0 26497.5 69620.0 26632.5 ;
      RECT  69555.0 27357.5 69620.0 27492.5 ;
      RECT  69745.0 27357.5 69810.0 27492.5 ;
      RECT  69745.0 27357.5 69810.0 27492.5 ;
      RECT  69555.0 27357.5 69620.0 27492.5 ;
      RECT  69482.5 27772.5 69547.5 27907.5 ;
      RECT  69817.5 26222.5 69882.5 26357.5 ;
      RECT  69555.0 27357.5 69620.0 27492.5 ;
      RECT  69745.0 26497.5 69810.0 26632.5 ;
      RECT  70002.5 26397.5 70067.5 26532.5 ;
      RECT  70002.5 26397.5 70067.5 26532.5 ;
      RECT  70450.0 27807.5 70515.0 27872.5 ;
      RECT  70185.0 27807.5 70482.5 27872.5 ;
      RECT  70450.0 27425.0 70515.0 27840.0 ;
      RECT  70260.0 26257.5 70325.0 26322.5 ;
      RECT  70292.5 26257.5 70555.0 26322.5 ;
      RECT  70260.0 26290.0 70325.0 26565.0 ;
      RECT  70260.0 26497.5 70325.0 26632.5 ;
      RECT  70450.0 26497.5 70515.0 26632.5 ;
      RECT  70450.0 26497.5 70515.0 26632.5 ;
      RECT  70260.0 26497.5 70325.0 26632.5 ;
      RECT  70260.0 27357.5 70325.0 27492.5 ;
      RECT  70450.0 27357.5 70515.0 27492.5 ;
      RECT  70450.0 27357.5 70515.0 27492.5 ;
      RECT  70260.0 27357.5 70325.0 27492.5 ;
      RECT  70187.5 27772.5 70252.5 27907.5 ;
      RECT  70522.5 26222.5 70587.5 26357.5 ;
      RECT  70260.0 27357.5 70325.0 27492.5 ;
      RECT  70450.0 26497.5 70515.0 26632.5 ;
      RECT  70707.5 26397.5 70772.5 26532.5 ;
      RECT  70707.5 26397.5 70772.5 26532.5 ;
      RECT  71155.0 27807.5 71220.0 27872.5 ;
      RECT  70890.0 27807.5 71187.5 27872.5 ;
      RECT  71155.0 27425.0 71220.0 27840.0 ;
      RECT  70965.0 26257.5 71030.0 26322.5 ;
      RECT  70997.5 26257.5 71260.0 26322.5 ;
      RECT  70965.0 26290.0 71030.0 26565.0 ;
      RECT  70965.0 26497.5 71030.0 26632.5 ;
      RECT  71155.0 26497.5 71220.0 26632.5 ;
      RECT  71155.0 26497.5 71220.0 26632.5 ;
      RECT  70965.0 26497.5 71030.0 26632.5 ;
      RECT  70965.0 27357.5 71030.0 27492.5 ;
      RECT  71155.0 27357.5 71220.0 27492.5 ;
      RECT  71155.0 27357.5 71220.0 27492.5 ;
      RECT  70965.0 27357.5 71030.0 27492.5 ;
      RECT  70892.5 27772.5 70957.5 27907.5 ;
      RECT  71227.5 26222.5 71292.5 26357.5 ;
      RECT  70965.0 27357.5 71030.0 27492.5 ;
      RECT  71155.0 26497.5 71220.0 26632.5 ;
      RECT  71412.5 26397.5 71477.5 26532.5 ;
      RECT  71412.5 26397.5 71477.5 26532.5 ;
      RECT  71860.0 27807.5 71925.0 27872.5 ;
      RECT  71595.0 27807.5 71892.5 27872.5 ;
      RECT  71860.0 27425.0 71925.0 27840.0 ;
      RECT  71670.0 26257.5 71735.0 26322.5 ;
      RECT  71702.5 26257.5 71965.0 26322.5 ;
      RECT  71670.0 26290.0 71735.0 26565.0 ;
      RECT  71670.0 26497.5 71735.0 26632.5 ;
      RECT  71860.0 26497.5 71925.0 26632.5 ;
      RECT  71860.0 26497.5 71925.0 26632.5 ;
      RECT  71670.0 26497.5 71735.0 26632.5 ;
      RECT  71670.0 27357.5 71735.0 27492.5 ;
      RECT  71860.0 27357.5 71925.0 27492.5 ;
      RECT  71860.0 27357.5 71925.0 27492.5 ;
      RECT  71670.0 27357.5 71735.0 27492.5 ;
      RECT  71597.5 27772.5 71662.5 27907.5 ;
      RECT  71932.5 26222.5 71997.5 26357.5 ;
      RECT  71670.0 27357.5 71735.0 27492.5 ;
      RECT  71860.0 26497.5 71925.0 26632.5 ;
      RECT  72117.5 26397.5 72182.5 26532.5 ;
      RECT  72117.5 26397.5 72182.5 26532.5 ;
      RECT  72565.0 27807.5 72630.0 27872.5 ;
      RECT  72300.0 27807.5 72597.5 27872.5 ;
      RECT  72565.0 27425.0 72630.0 27840.0 ;
      RECT  72375.0 26257.5 72440.0 26322.5 ;
      RECT  72407.5 26257.5 72670.0 26322.5 ;
      RECT  72375.0 26290.0 72440.0 26565.0 ;
      RECT  72375.0 26497.5 72440.0 26632.5 ;
      RECT  72565.0 26497.5 72630.0 26632.5 ;
      RECT  72565.0 26497.5 72630.0 26632.5 ;
      RECT  72375.0 26497.5 72440.0 26632.5 ;
      RECT  72375.0 27357.5 72440.0 27492.5 ;
      RECT  72565.0 27357.5 72630.0 27492.5 ;
      RECT  72565.0 27357.5 72630.0 27492.5 ;
      RECT  72375.0 27357.5 72440.0 27492.5 ;
      RECT  72302.5 27772.5 72367.5 27907.5 ;
      RECT  72637.5 26222.5 72702.5 26357.5 ;
      RECT  72375.0 27357.5 72440.0 27492.5 ;
      RECT  72565.0 26497.5 72630.0 26632.5 ;
      RECT  72822.5 26397.5 72887.5 26532.5 ;
      RECT  72822.5 26397.5 72887.5 26532.5 ;
      RECT  73270.0 27807.5 73335.0 27872.5 ;
      RECT  73005.0 27807.5 73302.5 27872.5 ;
      RECT  73270.0 27425.0 73335.0 27840.0 ;
      RECT  73080.0 26257.5 73145.0 26322.5 ;
      RECT  73112.5 26257.5 73375.0 26322.5 ;
      RECT  73080.0 26290.0 73145.0 26565.0 ;
      RECT  73080.0 26497.5 73145.0 26632.5 ;
      RECT  73270.0 26497.5 73335.0 26632.5 ;
      RECT  73270.0 26497.5 73335.0 26632.5 ;
      RECT  73080.0 26497.5 73145.0 26632.5 ;
      RECT  73080.0 27357.5 73145.0 27492.5 ;
      RECT  73270.0 27357.5 73335.0 27492.5 ;
      RECT  73270.0 27357.5 73335.0 27492.5 ;
      RECT  73080.0 27357.5 73145.0 27492.5 ;
      RECT  73007.5 27772.5 73072.5 27907.5 ;
      RECT  73342.5 26222.5 73407.5 26357.5 ;
      RECT  73080.0 27357.5 73145.0 27492.5 ;
      RECT  73270.0 26497.5 73335.0 26632.5 ;
      RECT  73527.5 26397.5 73592.5 26532.5 ;
      RECT  73527.5 26397.5 73592.5 26532.5 ;
      RECT  73975.0 27807.5 74040.0 27872.5 ;
      RECT  73710.0 27807.5 74007.5 27872.5 ;
      RECT  73975.0 27425.0 74040.0 27840.0 ;
      RECT  73785.0 26257.5 73850.0 26322.5 ;
      RECT  73817.5 26257.5 74080.0 26322.5 ;
      RECT  73785.0 26290.0 73850.0 26565.0 ;
      RECT  73785.0 26497.5 73850.0 26632.5 ;
      RECT  73975.0 26497.5 74040.0 26632.5 ;
      RECT  73975.0 26497.5 74040.0 26632.5 ;
      RECT  73785.0 26497.5 73850.0 26632.5 ;
      RECT  73785.0 27357.5 73850.0 27492.5 ;
      RECT  73975.0 27357.5 74040.0 27492.5 ;
      RECT  73975.0 27357.5 74040.0 27492.5 ;
      RECT  73785.0 27357.5 73850.0 27492.5 ;
      RECT  73712.5 27772.5 73777.5 27907.5 ;
      RECT  74047.5 26222.5 74112.5 26357.5 ;
      RECT  73785.0 27357.5 73850.0 27492.5 ;
      RECT  73975.0 26497.5 74040.0 26632.5 ;
      RECT  74232.5 26397.5 74297.5 26532.5 ;
      RECT  74232.5 26397.5 74297.5 26532.5 ;
      RECT  74680.0 27807.5 74745.0 27872.5 ;
      RECT  74415.0 27807.5 74712.5 27872.5 ;
      RECT  74680.0 27425.0 74745.0 27840.0 ;
      RECT  74490.0 26257.5 74555.0 26322.5 ;
      RECT  74522.5 26257.5 74785.0 26322.5 ;
      RECT  74490.0 26290.0 74555.0 26565.0 ;
      RECT  74490.0 26497.5 74555.0 26632.5 ;
      RECT  74680.0 26497.5 74745.0 26632.5 ;
      RECT  74680.0 26497.5 74745.0 26632.5 ;
      RECT  74490.0 26497.5 74555.0 26632.5 ;
      RECT  74490.0 27357.5 74555.0 27492.5 ;
      RECT  74680.0 27357.5 74745.0 27492.5 ;
      RECT  74680.0 27357.5 74745.0 27492.5 ;
      RECT  74490.0 27357.5 74555.0 27492.5 ;
      RECT  74417.5 27772.5 74482.5 27907.5 ;
      RECT  74752.5 26222.5 74817.5 26357.5 ;
      RECT  74490.0 27357.5 74555.0 27492.5 ;
      RECT  74680.0 26497.5 74745.0 26632.5 ;
      RECT  74937.5 26397.5 75002.5 26532.5 ;
      RECT  74937.5 26397.5 75002.5 26532.5 ;
      RECT  75385.0 27807.5 75450.0 27872.5 ;
      RECT  75120.0 27807.5 75417.5 27872.5 ;
      RECT  75385.0 27425.0 75450.0 27840.0 ;
      RECT  75195.0 26257.5 75260.0 26322.5 ;
      RECT  75227.5 26257.5 75490.0 26322.5 ;
      RECT  75195.0 26290.0 75260.0 26565.0 ;
      RECT  75195.0 26497.5 75260.0 26632.5 ;
      RECT  75385.0 26497.5 75450.0 26632.5 ;
      RECT  75385.0 26497.5 75450.0 26632.5 ;
      RECT  75195.0 26497.5 75260.0 26632.5 ;
      RECT  75195.0 27357.5 75260.0 27492.5 ;
      RECT  75385.0 27357.5 75450.0 27492.5 ;
      RECT  75385.0 27357.5 75450.0 27492.5 ;
      RECT  75195.0 27357.5 75260.0 27492.5 ;
      RECT  75122.5 27772.5 75187.5 27907.5 ;
      RECT  75457.5 26222.5 75522.5 26357.5 ;
      RECT  75195.0 27357.5 75260.0 27492.5 ;
      RECT  75385.0 26497.5 75450.0 26632.5 ;
      RECT  75642.5 26397.5 75707.5 26532.5 ;
      RECT  75642.5 26397.5 75707.5 26532.5 ;
      RECT  76090.0 27807.5 76155.0 27872.5 ;
      RECT  75825.0 27807.5 76122.5 27872.5 ;
      RECT  76090.0 27425.0 76155.0 27840.0 ;
      RECT  75900.0 26257.5 75965.0 26322.5 ;
      RECT  75932.5 26257.5 76195.0 26322.5 ;
      RECT  75900.0 26290.0 75965.0 26565.0 ;
      RECT  75900.0 26497.5 75965.0 26632.5 ;
      RECT  76090.0 26497.5 76155.0 26632.5 ;
      RECT  76090.0 26497.5 76155.0 26632.5 ;
      RECT  75900.0 26497.5 75965.0 26632.5 ;
      RECT  75900.0 27357.5 75965.0 27492.5 ;
      RECT  76090.0 27357.5 76155.0 27492.5 ;
      RECT  76090.0 27357.5 76155.0 27492.5 ;
      RECT  75900.0 27357.5 75965.0 27492.5 ;
      RECT  75827.5 27772.5 75892.5 27907.5 ;
      RECT  76162.5 26222.5 76227.5 26357.5 ;
      RECT  75900.0 27357.5 75965.0 27492.5 ;
      RECT  76090.0 26497.5 76155.0 26632.5 ;
      RECT  76347.5 26397.5 76412.5 26532.5 ;
      RECT  76347.5 26397.5 76412.5 26532.5 ;
      RECT  76795.0 27807.5 76860.0 27872.5 ;
      RECT  76530.0 27807.5 76827.5 27872.5 ;
      RECT  76795.0 27425.0 76860.0 27840.0 ;
      RECT  76605.0 26257.5 76670.0 26322.5 ;
      RECT  76637.5 26257.5 76900.0 26322.5 ;
      RECT  76605.0 26290.0 76670.0 26565.0 ;
      RECT  76605.0 26497.5 76670.0 26632.5 ;
      RECT  76795.0 26497.5 76860.0 26632.5 ;
      RECT  76795.0 26497.5 76860.0 26632.5 ;
      RECT  76605.0 26497.5 76670.0 26632.5 ;
      RECT  76605.0 27357.5 76670.0 27492.5 ;
      RECT  76795.0 27357.5 76860.0 27492.5 ;
      RECT  76795.0 27357.5 76860.0 27492.5 ;
      RECT  76605.0 27357.5 76670.0 27492.5 ;
      RECT  76532.5 27772.5 76597.5 27907.5 ;
      RECT  76867.5 26222.5 76932.5 26357.5 ;
      RECT  76605.0 27357.5 76670.0 27492.5 ;
      RECT  76795.0 26497.5 76860.0 26632.5 ;
      RECT  77052.5 26397.5 77117.5 26532.5 ;
      RECT  77052.5 26397.5 77117.5 26532.5 ;
      RECT  77500.0 27807.5 77565.0 27872.5 ;
      RECT  77235.0 27807.5 77532.5 27872.5 ;
      RECT  77500.0 27425.0 77565.0 27840.0 ;
      RECT  77310.0 26257.5 77375.0 26322.5 ;
      RECT  77342.5 26257.5 77605.0 26322.5 ;
      RECT  77310.0 26290.0 77375.0 26565.0 ;
      RECT  77310.0 26497.5 77375.0 26632.5 ;
      RECT  77500.0 26497.5 77565.0 26632.5 ;
      RECT  77500.0 26497.5 77565.0 26632.5 ;
      RECT  77310.0 26497.5 77375.0 26632.5 ;
      RECT  77310.0 27357.5 77375.0 27492.5 ;
      RECT  77500.0 27357.5 77565.0 27492.5 ;
      RECT  77500.0 27357.5 77565.0 27492.5 ;
      RECT  77310.0 27357.5 77375.0 27492.5 ;
      RECT  77237.5 27772.5 77302.5 27907.5 ;
      RECT  77572.5 26222.5 77637.5 26357.5 ;
      RECT  77310.0 27357.5 77375.0 27492.5 ;
      RECT  77500.0 26497.5 77565.0 26632.5 ;
      RECT  77757.5 26397.5 77822.5 26532.5 ;
      RECT  77757.5 26397.5 77822.5 26532.5 ;
      RECT  78205.0 27807.5 78270.0 27872.5 ;
      RECT  77940.0 27807.5 78237.5 27872.5 ;
      RECT  78205.0 27425.0 78270.0 27840.0 ;
      RECT  78015.0 26257.5 78080.0 26322.5 ;
      RECT  78047.5 26257.5 78310.0 26322.5 ;
      RECT  78015.0 26290.0 78080.0 26565.0 ;
      RECT  78015.0 26497.5 78080.0 26632.5 ;
      RECT  78205.0 26497.5 78270.0 26632.5 ;
      RECT  78205.0 26497.5 78270.0 26632.5 ;
      RECT  78015.0 26497.5 78080.0 26632.5 ;
      RECT  78015.0 27357.5 78080.0 27492.5 ;
      RECT  78205.0 27357.5 78270.0 27492.5 ;
      RECT  78205.0 27357.5 78270.0 27492.5 ;
      RECT  78015.0 27357.5 78080.0 27492.5 ;
      RECT  77942.5 27772.5 78007.5 27907.5 ;
      RECT  78277.5 26222.5 78342.5 26357.5 ;
      RECT  78015.0 27357.5 78080.0 27492.5 ;
      RECT  78205.0 26497.5 78270.0 26632.5 ;
      RECT  78462.5 26397.5 78527.5 26532.5 ;
      RECT  78462.5 26397.5 78527.5 26532.5 ;
      RECT  78910.0 27807.5 78975.0 27872.5 ;
      RECT  78645.0 27807.5 78942.5 27872.5 ;
      RECT  78910.0 27425.0 78975.0 27840.0 ;
      RECT  78720.0 26257.5 78785.0 26322.5 ;
      RECT  78752.5 26257.5 79015.0 26322.5 ;
      RECT  78720.0 26290.0 78785.0 26565.0 ;
      RECT  78720.0 26497.5 78785.0 26632.5 ;
      RECT  78910.0 26497.5 78975.0 26632.5 ;
      RECT  78910.0 26497.5 78975.0 26632.5 ;
      RECT  78720.0 26497.5 78785.0 26632.5 ;
      RECT  78720.0 27357.5 78785.0 27492.5 ;
      RECT  78910.0 27357.5 78975.0 27492.5 ;
      RECT  78910.0 27357.5 78975.0 27492.5 ;
      RECT  78720.0 27357.5 78785.0 27492.5 ;
      RECT  78647.5 27772.5 78712.5 27907.5 ;
      RECT  78982.5 26222.5 79047.5 26357.5 ;
      RECT  78720.0 27357.5 78785.0 27492.5 ;
      RECT  78910.0 26497.5 78975.0 26632.5 ;
      RECT  79167.5 26397.5 79232.5 26532.5 ;
      RECT  79167.5 26397.5 79232.5 26532.5 ;
      RECT  79615.0 27807.5 79680.0 27872.5 ;
      RECT  79350.0 27807.5 79647.5 27872.5 ;
      RECT  79615.0 27425.0 79680.0 27840.0 ;
      RECT  79425.0 26257.5 79490.0 26322.5 ;
      RECT  79457.5 26257.5 79720.0 26322.5 ;
      RECT  79425.0 26290.0 79490.0 26565.0 ;
      RECT  79425.0 26497.5 79490.0 26632.5 ;
      RECT  79615.0 26497.5 79680.0 26632.5 ;
      RECT  79615.0 26497.5 79680.0 26632.5 ;
      RECT  79425.0 26497.5 79490.0 26632.5 ;
      RECT  79425.0 27357.5 79490.0 27492.5 ;
      RECT  79615.0 27357.5 79680.0 27492.5 ;
      RECT  79615.0 27357.5 79680.0 27492.5 ;
      RECT  79425.0 27357.5 79490.0 27492.5 ;
      RECT  79352.5 27772.5 79417.5 27907.5 ;
      RECT  79687.5 26222.5 79752.5 26357.5 ;
      RECT  79425.0 27357.5 79490.0 27492.5 ;
      RECT  79615.0 26497.5 79680.0 26632.5 ;
      RECT  79872.5 26397.5 79937.5 26532.5 ;
      RECT  79872.5 26397.5 79937.5 26532.5 ;
      RECT  80320.0 27807.5 80385.0 27872.5 ;
      RECT  80055.0 27807.5 80352.5 27872.5 ;
      RECT  80320.0 27425.0 80385.0 27840.0 ;
      RECT  80130.0 26257.5 80195.0 26322.5 ;
      RECT  80162.5 26257.5 80425.0 26322.5 ;
      RECT  80130.0 26290.0 80195.0 26565.0 ;
      RECT  80130.0 26497.5 80195.0 26632.5 ;
      RECT  80320.0 26497.5 80385.0 26632.5 ;
      RECT  80320.0 26497.5 80385.0 26632.5 ;
      RECT  80130.0 26497.5 80195.0 26632.5 ;
      RECT  80130.0 27357.5 80195.0 27492.5 ;
      RECT  80320.0 27357.5 80385.0 27492.5 ;
      RECT  80320.0 27357.5 80385.0 27492.5 ;
      RECT  80130.0 27357.5 80195.0 27492.5 ;
      RECT  80057.5 27772.5 80122.5 27907.5 ;
      RECT  80392.5 26222.5 80457.5 26357.5 ;
      RECT  80130.0 27357.5 80195.0 27492.5 ;
      RECT  80320.0 26497.5 80385.0 26632.5 ;
      RECT  80577.5 26397.5 80642.5 26532.5 ;
      RECT  80577.5 26397.5 80642.5 26532.5 ;
      RECT  81025.0 27807.5 81090.0 27872.5 ;
      RECT  80760.0 27807.5 81057.5 27872.5 ;
      RECT  81025.0 27425.0 81090.0 27840.0 ;
      RECT  80835.0 26257.5 80900.0 26322.5 ;
      RECT  80867.5 26257.5 81130.0 26322.5 ;
      RECT  80835.0 26290.0 80900.0 26565.0 ;
      RECT  80835.0 26497.5 80900.0 26632.5 ;
      RECT  81025.0 26497.5 81090.0 26632.5 ;
      RECT  81025.0 26497.5 81090.0 26632.5 ;
      RECT  80835.0 26497.5 80900.0 26632.5 ;
      RECT  80835.0 27357.5 80900.0 27492.5 ;
      RECT  81025.0 27357.5 81090.0 27492.5 ;
      RECT  81025.0 27357.5 81090.0 27492.5 ;
      RECT  80835.0 27357.5 80900.0 27492.5 ;
      RECT  80762.5 27772.5 80827.5 27907.5 ;
      RECT  81097.5 26222.5 81162.5 26357.5 ;
      RECT  80835.0 27357.5 80900.0 27492.5 ;
      RECT  81025.0 26497.5 81090.0 26632.5 ;
      RECT  81282.5 26397.5 81347.5 26532.5 ;
      RECT  81282.5 26397.5 81347.5 26532.5 ;
      RECT  81730.0 27807.5 81795.0 27872.5 ;
      RECT  81465.0 27807.5 81762.5 27872.5 ;
      RECT  81730.0 27425.0 81795.0 27840.0 ;
      RECT  81540.0 26257.5 81605.0 26322.5 ;
      RECT  81572.5 26257.5 81835.0 26322.5 ;
      RECT  81540.0 26290.0 81605.0 26565.0 ;
      RECT  81540.0 26497.5 81605.0 26632.5 ;
      RECT  81730.0 26497.5 81795.0 26632.5 ;
      RECT  81730.0 26497.5 81795.0 26632.5 ;
      RECT  81540.0 26497.5 81605.0 26632.5 ;
      RECT  81540.0 27357.5 81605.0 27492.5 ;
      RECT  81730.0 27357.5 81795.0 27492.5 ;
      RECT  81730.0 27357.5 81795.0 27492.5 ;
      RECT  81540.0 27357.5 81605.0 27492.5 ;
      RECT  81467.5 27772.5 81532.5 27907.5 ;
      RECT  81802.5 26222.5 81867.5 26357.5 ;
      RECT  81540.0 27357.5 81605.0 27492.5 ;
      RECT  81730.0 26497.5 81795.0 26632.5 ;
      RECT  81987.5 26397.5 82052.5 26532.5 ;
      RECT  81987.5 26397.5 82052.5 26532.5 ;
      RECT  82435.0 27807.5 82500.0 27872.5 ;
      RECT  82170.0 27807.5 82467.5 27872.5 ;
      RECT  82435.0 27425.0 82500.0 27840.0 ;
      RECT  82245.0 26257.5 82310.0 26322.5 ;
      RECT  82277.5 26257.5 82540.0 26322.5 ;
      RECT  82245.0 26290.0 82310.0 26565.0 ;
      RECT  82245.0 26497.5 82310.0 26632.5 ;
      RECT  82435.0 26497.5 82500.0 26632.5 ;
      RECT  82435.0 26497.5 82500.0 26632.5 ;
      RECT  82245.0 26497.5 82310.0 26632.5 ;
      RECT  82245.0 27357.5 82310.0 27492.5 ;
      RECT  82435.0 27357.5 82500.0 27492.5 ;
      RECT  82435.0 27357.5 82500.0 27492.5 ;
      RECT  82245.0 27357.5 82310.0 27492.5 ;
      RECT  82172.5 27772.5 82237.5 27907.5 ;
      RECT  82507.5 26222.5 82572.5 26357.5 ;
      RECT  82245.0 27357.5 82310.0 27492.5 ;
      RECT  82435.0 26497.5 82500.0 26632.5 ;
      RECT  82692.5 26397.5 82757.5 26532.5 ;
      RECT  82692.5 26397.5 82757.5 26532.5 ;
      RECT  83140.0 27807.5 83205.0 27872.5 ;
      RECT  82875.0 27807.5 83172.5 27872.5 ;
      RECT  83140.0 27425.0 83205.0 27840.0 ;
      RECT  82950.0 26257.5 83015.0 26322.5 ;
      RECT  82982.5 26257.5 83245.0 26322.5 ;
      RECT  82950.0 26290.0 83015.0 26565.0 ;
      RECT  82950.0 26497.5 83015.0 26632.5 ;
      RECT  83140.0 26497.5 83205.0 26632.5 ;
      RECT  83140.0 26497.5 83205.0 26632.5 ;
      RECT  82950.0 26497.5 83015.0 26632.5 ;
      RECT  82950.0 27357.5 83015.0 27492.5 ;
      RECT  83140.0 27357.5 83205.0 27492.5 ;
      RECT  83140.0 27357.5 83205.0 27492.5 ;
      RECT  82950.0 27357.5 83015.0 27492.5 ;
      RECT  82877.5 27772.5 82942.5 27907.5 ;
      RECT  83212.5 26222.5 83277.5 26357.5 ;
      RECT  82950.0 27357.5 83015.0 27492.5 ;
      RECT  83140.0 26497.5 83205.0 26632.5 ;
      RECT  83397.5 26397.5 83462.5 26532.5 ;
      RECT  83397.5 26397.5 83462.5 26532.5 ;
      RECT  83845.0 27807.5 83910.0 27872.5 ;
      RECT  83580.0 27807.5 83877.5 27872.5 ;
      RECT  83845.0 27425.0 83910.0 27840.0 ;
      RECT  83655.0 26257.5 83720.0 26322.5 ;
      RECT  83687.5 26257.5 83950.0 26322.5 ;
      RECT  83655.0 26290.0 83720.0 26565.0 ;
      RECT  83655.0 26497.5 83720.0 26632.5 ;
      RECT  83845.0 26497.5 83910.0 26632.5 ;
      RECT  83845.0 26497.5 83910.0 26632.5 ;
      RECT  83655.0 26497.5 83720.0 26632.5 ;
      RECT  83655.0 27357.5 83720.0 27492.5 ;
      RECT  83845.0 27357.5 83910.0 27492.5 ;
      RECT  83845.0 27357.5 83910.0 27492.5 ;
      RECT  83655.0 27357.5 83720.0 27492.5 ;
      RECT  83582.5 27772.5 83647.5 27907.5 ;
      RECT  83917.5 26222.5 83982.5 26357.5 ;
      RECT  83655.0 27357.5 83720.0 27492.5 ;
      RECT  83845.0 26497.5 83910.0 26632.5 ;
      RECT  84102.5 26397.5 84167.5 26532.5 ;
      RECT  84102.5 26397.5 84167.5 26532.5 ;
      RECT  84550.0 27807.5 84615.0 27872.5 ;
      RECT  84285.0 27807.5 84582.5 27872.5 ;
      RECT  84550.0 27425.0 84615.0 27840.0 ;
      RECT  84360.0 26257.5 84425.0 26322.5 ;
      RECT  84392.5 26257.5 84655.0 26322.5 ;
      RECT  84360.0 26290.0 84425.0 26565.0 ;
      RECT  84360.0 26497.5 84425.0 26632.5 ;
      RECT  84550.0 26497.5 84615.0 26632.5 ;
      RECT  84550.0 26497.5 84615.0 26632.5 ;
      RECT  84360.0 26497.5 84425.0 26632.5 ;
      RECT  84360.0 27357.5 84425.0 27492.5 ;
      RECT  84550.0 27357.5 84615.0 27492.5 ;
      RECT  84550.0 27357.5 84615.0 27492.5 ;
      RECT  84360.0 27357.5 84425.0 27492.5 ;
      RECT  84287.5 27772.5 84352.5 27907.5 ;
      RECT  84622.5 26222.5 84687.5 26357.5 ;
      RECT  84360.0 27357.5 84425.0 27492.5 ;
      RECT  84550.0 26497.5 84615.0 26632.5 ;
      RECT  84807.5 26397.5 84872.5 26532.5 ;
      RECT  84807.5 26397.5 84872.5 26532.5 ;
      RECT  85255.0 27807.5 85320.0 27872.5 ;
      RECT  84990.0 27807.5 85287.5 27872.5 ;
      RECT  85255.0 27425.0 85320.0 27840.0 ;
      RECT  85065.0 26257.5 85130.0 26322.5 ;
      RECT  85097.5 26257.5 85360.0 26322.5 ;
      RECT  85065.0 26290.0 85130.0 26565.0 ;
      RECT  85065.0 26497.5 85130.0 26632.5 ;
      RECT  85255.0 26497.5 85320.0 26632.5 ;
      RECT  85255.0 26497.5 85320.0 26632.5 ;
      RECT  85065.0 26497.5 85130.0 26632.5 ;
      RECT  85065.0 27357.5 85130.0 27492.5 ;
      RECT  85255.0 27357.5 85320.0 27492.5 ;
      RECT  85255.0 27357.5 85320.0 27492.5 ;
      RECT  85065.0 27357.5 85130.0 27492.5 ;
      RECT  84992.5 27772.5 85057.5 27907.5 ;
      RECT  85327.5 26222.5 85392.5 26357.5 ;
      RECT  85065.0 27357.5 85130.0 27492.5 ;
      RECT  85255.0 26497.5 85320.0 26632.5 ;
      RECT  85512.5 26397.5 85577.5 26532.5 ;
      RECT  85512.5 26397.5 85577.5 26532.5 ;
      RECT  85960.0 27807.5 86025.0 27872.5 ;
      RECT  85695.0 27807.5 85992.5 27872.5 ;
      RECT  85960.0 27425.0 86025.0 27840.0 ;
      RECT  85770.0 26257.5 85835.0 26322.5 ;
      RECT  85802.5 26257.5 86065.0 26322.5 ;
      RECT  85770.0 26290.0 85835.0 26565.0 ;
      RECT  85770.0 26497.5 85835.0 26632.5 ;
      RECT  85960.0 26497.5 86025.0 26632.5 ;
      RECT  85960.0 26497.5 86025.0 26632.5 ;
      RECT  85770.0 26497.5 85835.0 26632.5 ;
      RECT  85770.0 27357.5 85835.0 27492.5 ;
      RECT  85960.0 27357.5 86025.0 27492.5 ;
      RECT  85960.0 27357.5 86025.0 27492.5 ;
      RECT  85770.0 27357.5 85835.0 27492.5 ;
      RECT  85697.5 27772.5 85762.5 27907.5 ;
      RECT  86032.5 26222.5 86097.5 26357.5 ;
      RECT  85770.0 27357.5 85835.0 27492.5 ;
      RECT  85960.0 26497.5 86025.0 26632.5 ;
      RECT  86217.5 26397.5 86282.5 26532.5 ;
      RECT  86217.5 26397.5 86282.5 26532.5 ;
      RECT  86665.0 27807.5 86730.0 27872.5 ;
      RECT  86400.0 27807.5 86697.5 27872.5 ;
      RECT  86665.0 27425.0 86730.0 27840.0 ;
      RECT  86475.0 26257.5 86540.0 26322.5 ;
      RECT  86507.5 26257.5 86770.0 26322.5 ;
      RECT  86475.0 26290.0 86540.0 26565.0 ;
      RECT  86475.0 26497.5 86540.0 26632.5 ;
      RECT  86665.0 26497.5 86730.0 26632.5 ;
      RECT  86665.0 26497.5 86730.0 26632.5 ;
      RECT  86475.0 26497.5 86540.0 26632.5 ;
      RECT  86475.0 27357.5 86540.0 27492.5 ;
      RECT  86665.0 27357.5 86730.0 27492.5 ;
      RECT  86665.0 27357.5 86730.0 27492.5 ;
      RECT  86475.0 27357.5 86540.0 27492.5 ;
      RECT  86402.5 27772.5 86467.5 27907.5 ;
      RECT  86737.5 26222.5 86802.5 26357.5 ;
      RECT  86475.0 27357.5 86540.0 27492.5 ;
      RECT  86665.0 26497.5 86730.0 26632.5 ;
      RECT  86922.5 26397.5 86987.5 26532.5 ;
      RECT  86922.5 26397.5 86987.5 26532.5 ;
      RECT  87370.0 27807.5 87435.0 27872.5 ;
      RECT  87105.0 27807.5 87402.5 27872.5 ;
      RECT  87370.0 27425.0 87435.0 27840.0 ;
      RECT  87180.0 26257.5 87245.0 26322.5 ;
      RECT  87212.5 26257.5 87475.0 26322.5 ;
      RECT  87180.0 26290.0 87245.0 26565.0 ;
      RECT  87180.0 26497.5 87245.0 26632.5 ;
      RECT  87370.0 26497.5 87435.0 26632.5 ;
      RECT  87370.0 26497.5 87435.0 26632.5 ;
      RECT  87180.0 26497.5 87245.0 26632.5 ;
      RECT  87180.0 27357.5 87245.0 27492.5 ;
      RECT  87370.0 27357.5 87435.0 27492.5 ;
      RECT  87370.0 27357.5 87435.0 27492.5 ;
      RECT  87180.0 27357.5 87245.0 27492.5 ;
      RECT  87107.5 27772.5 87172.5 27907.5 ;
      RECT  87442.5 26222.5 87507.5 26357.5 ;
      RECT  87180.0 27357.5 87245.0 27492.5 ;
      RECT  87370.0 26497.5 87435.0 26632.5 ;
      RECT  87627.5 26397.5 87692.5 26532.5 ;
      RECT  87627.5 26397.5 87692.5 26532.5 ;
      RECT  88075.0 27807.5 88140.0 27872.5 ;
      RECT  87810.0 27807.5 88107.5 27872.5 ;
      RECT  88075.0 27425.0 88140.0 27840.0 ;
      RECT  87885.0 26257.5 87950.0 26322.5 ;
      RECT  87917.5 26257.5 88180.0 26322.5 ;
      RECT  87885.0 26290.0 87950.0 26565.0 ;
      RECT  87885.0 26497.5 87950.0 26632.5 ;
      RECT  88075.0 26497.5 88140.0 26632.5 ;
      RECT  88075.0 26497.5 88140.0 26632.5 ;
      RECT  87885.0 26497.5 87950.0 26632.5 ;
      RECT  87885.0 27357.5 87950.0 27492.5 ;
      RECT  88075.0 27357.5 88140.0 27492.5 ;
      RECT  88075.0 27357.5 88140.0 27492.5 ;
      RECT  87885.0 27357.5 87950.0 27492.5 ;
      RECT  87812.5 27772.5 87877.5 27907.5 ;
      RECT  88147.5 26222.5 88212.5 26357.5 ;
      RECT  87885.0 27357.5 87950.0 27492.5 ;
      RECT  88075.0 26497.5 88140.0 26632.5 ;
      RECT  88332.5 26397.5 88397.5 26532.5 ;
      RECT  88332.5 26397.5 88397.5 26532.5 ;
      RECT  88780.0 27807.5 88845.0 27872.5 ;
      RECT  88515.0 27807.5 88812.5 27872.5 ;
      RECT  88780.0 27425.0 88845.0 27840.0 ;
      RECT  88590.0 26257.5 88655.0 26322.5 ;
      RECT  88622.5 26257.5 88885.0 26322.5 ;
      RECT  88590.0 26290.0 88655.0 26565.0 ;
      RECT  88590.0 26497.5 88655.0 26632.5 ;
      RECT  88780.0 26497.5 88845.0 26632.5 ;
      RECT  88780.0 26497.5 88845.0 26632.5 ;
      RECT  88590.0 26497.5 88655.0 26632.5 ;
      RECT  88590.0 27357.5 88655.0 27492.5 ;
      RECT  88780.0 27357.5 88845.0 27492.5 ;
      RECT  88780.0 27357.5 88845.0 27492.5 ;
      RECT  88590.0 27357.5 88655.0 27492.5 ;
      RECT  88517.5 27772.5 88582.5 27907.5 ;
      RECT  88852.5 26222.5 88917.5 26357.5 ;
      RECT  88590.0 27357.5 88655.0 27492.5 ;
      RECT  88780.0 26497.5 88845.0 26632.5 ;
      RECT  89037.5 26397.5 89102.5 26532.5 ;
      RECT  89037.5 26397.5 89102.5 26532.5 ;
      RECT  89485.0 27807.5 89550.0 27872.5 ;
      RECT  89220.0 27807.5 89517.5 27872.5 ;
      RECT  89485.0 27425.0 89550.0 27840.0 ;
      RECT  89295.0 26257.5 89360.0 26322.5 ;
      RECT  89327.5 26257.5 89590.0 26322.5 ;
      RECT  89295.0 26290.0 89360.0 26565.0 ;
      RECT  89295.0 26497.5 89360.0 26632.5 ;
      RECT  89485.0 26497.5 89550.0 26632.5 ;
      RECT  89485.0 26497.5 89550.0 26632.5 ;
      RECT  89295.0 26497.5 89360.0 26632.5 ;
      RECT  89295.0 27357.5 89360.0 27492.5 ;
      RECT  89485.0 27357.5 89550.0 27492.5 ;
      RECT  89485.0 27357.5 89550.0 27492.5 ;
      RECT  89295.0 27357.5 89360.0 27492.5 ;
      RECT  89222.5 27772.5 89287.5 27907.5 ;
      RECT  89557.5 26222.5 89622.5 26357.5 ;
      RECT  89295.0 27357.5 89360.0 27492.5 ;
      RECT  89485.0 26497.5 89550.0 26632.5 ;
      RECT  89742.5 26397.5 89807.5 26532.5 ;
      RECT  89742.5 26397.5 89807.5 26532.5 ;
      RECT  90190.0 27807.5 90255.0 27872.5 ;
      RECT  89925.0 27807.5 90222.5 27872.5 ;
      RECT  90190.0 27425.0 90255.0 27840.0 ;
      RECT  90000.0 26257.5 90065.0 26322.5 ;
      RECT  90032.5 26257.5 90295.0 26322.5 ;
      RECT  90000.0 26290.0 90065.0 26565.0 ;
      RECT  90000.0 26497.5 90065.0 26632.5 ;
      RECT  90190.0 26497.5 90255.0 26632.5 ;
      RECT  90190.0 26497.5 90255.0 26632.5 ;
      RECT  90000.0 26497.5 90065.0 26632.5 ;
      RECT  90000.0 27357.5 90065.0 27492.5 ;
      RECT  90190.0 27357.5 90255.0 27492.5 ;
      RECT  90190.0 27357.5 90255.0 27492.5 ;
      RECT  90000.0 27357.5 90065.0 27492.5 ;
      RECT  89927.5 27772.5 89992.5 27907.5 ;
      RECT  90262.5 26222.5 90327.5 26357.5 ;
      RECT  90000.0 27357.5 90065.0 27492.5 ;
      RECT  90190.0 26497.5 90255.0 26632.5 ;
      RECT  90447.5 26397.5 90512.5 26532.5 ;
      RECT  90447.5 26397.5 90512.5 26532.5 ;
      RECT  90895.0 27807.5 90960.0 27872.5 ;
      RECT  90630.0 27807.5 90927.5 27872.5 ;
      RECT  90895.0 27425.0 90960.0 27840.0 ;
      RECT  90705.0 26257.5 90770.0 26322.5 ;
      RECT  90737.5 26257.5 91000.0 26322.5 ;
      RECT  90705.0 26290.0 90770.0 26565.0 ;
      RECT  90705.0 26497.5 90770.0 26632.5 ;
      RECT  90895.0 26497.5 90960.0 26632.5 ;
      RECT  90895.0 26497.5 90960.0 26632.5 ;
      RECT  90705.0 26497.5 90770.0 26632.5 ;
      RECT  90705.0 27357.5 90770.0 27492.5 ;
      RECT  90895.0 27357.5 90960.0 27492.5 ;
      RECT  90895.0 27357.5 90960.0 27492.5 ;
      RECT  90705.0 27357.5 90770.0 27492.5 ;
      RECT  90632.5 27772.5 90697.5 27907.5 ;
      RECT  90967.5 26222.5 91032.5 26357.5 ;
      RECT  90705.0 27357.5 90770.0 27492.5 ;
      RECT  90895.0 26497.5 90960.0 26632.5 ;
      RECT  91152.5 26397.5 91217.5 26532.5 ;
      RECT  91152.5 26397.5 91217.5 26532.5 ;
      RECT  91600.0 27807.5 91665.0 27872.5 ;
      RECT  91335.0 27807.5 91632.5 27872.5 ;
      RECT  91600.0 27425.0 91665.0 27840.0 ;
      RECT  91410.0 26257.5 91475.0 26322.5 ;
      RECT  91442.5 26257.5 91705.0 26322.5 ;
      RECT  91410.0 26290.0 91475.0 26565.0 ;
      RECT  91410.0 26497.5 91475.0 26632.5 ;
      RECT  91600.0 26497.5 91665.0 26632.5 ;
      RECT  91600.0 26497.5 91665.0 26632.5 ;
      RECT  91410.0 26497.5 91475.0 26632.5 ;
      RECT  91410.0 27357.5 91475.0 27492.5 ;
      RECT  91600.0 27357.5 91665.0 27492.5 ;
      RECT  91600.0 27357.5 91665.0 27492.5 ;
      RECT  91410.0 27357.5 91475.0 27492.5 ;
      RECT  91337.5 27772.5 91402.5 27907.5 ;
      RECT  91672.5 26222.5 91737.5 26357.5 ;
      RECT  91410.0 27357.5 91475.0 27492.5 ;
      RECT  91600.0 26497.5 91665.0 26632.5 ;
      RECT  91857.5 26397.5 91922.5 26532.5 ;
      RECT  91857.5 26397.5 91922.5 26532.5 ;
      RECT  92305.0 27807.5 92370.0 27872.5 ;
      RECT  92040.0 27807.5 92337.5 27872.5 ;
      RECT  92305.0 27425.0 92370.0 27840.0 ;
      RECT  92115.0 26257.5 92180.0 26322.5 ;
      RECT  92147.5 26257.5 92410.0 26322.5 ;
      RECT  92115.0 26290.0 92180.0 26565.0 ;
      RECT  92115.0 26497.5 92180.0 26632.5 ;
      RECT  92305.0 26497.5 92370.0 26632.5 ;
      RECT  92305.0 26497.5 92370.0 26632.5 ;
      RECT  92115.0 26497.5 92180.0 26632.5 ;
      RECT  92115.0 27357.5 92180.0 27492.5 ;
      RECT  92305.0 27357.5 92370.0 27492.5 ;
      RECT  92305.0 27357.5 92370.0 27492.5 ;
      RECT  92115.0 27357.5 92180.0 27492.5 ;
      RECT  92042.5 27772.5 92107.5 27907.5 ;
      RECT  92377.5 26222.5 92442.5 26357.5 ;
      RECT  92115.0 27357.5 92180.0 27492.5 ;
      RECT  92305.0 26497.5 92370.0 26632.5 ;
      RECT  92562.5 26397.5 92627.5 26532.5 ;
      RECT  92562.5 26397.5 92627.5 26532.5 ;
      RECT  93010.0 27807.5 93075.0 27872.5 ;
      RECT  92745.0 27807.5 93042.5 27872.5 ;
      RECT  93010.0 27425.0 93075.0 27840.0 ;
      RECT  92820.0 26257.5 92885.0 26322.5 ;
      RECT  92852.5 26257.5 93115.0 26322.5 ;
      RECT  92820.0 26290.0 92885.0 26565.0 ;
      RECT  92820.0 26497.5 92885.0 26632.5 ;
      RECT  93010.0 26497.5 93075.0 26632.5 ;
      RECT  93010.0 26497.5 93075.0 26632.5 ;
      RECT  92820.0 26497.5 92885.0 26632.5 ;
      RECT  92820.0 27357.5 92885.0 27492.5 ;
      RECT  93010.0 27357.5 93075.0 27492.5 ;
      RECT  93010.0 27357.5 93075.0 27492.5 ;
      RECT  92820.0 27357.5 92885.0 27492.5 ;
      RECT  92747.5 27772.5 92812.5 27907.5 ;
      RECT  93082.5 26222.5 93147.5 26357.5 ;
      RECT  92820.0 27357.5 92885.0 27492.5 ;
      RECT  93010.0 26497.5 93075.0 26632.5 ;
      RECT  93267.5 26397.5 93332.5 26532.5 ;
      RECT  93267.5 26397.5 93332.5 26532.5 ;
      RECT  93715.0 27807.5 93780.0 27872.5 ;
      RECT  93450.0 27807.5 93747.5 27872.5 ;
      RECT  93715.0 27425.0 93780.0 27840.0 ;
      RECT  93525.0 26257.5 93590.0 26322.5 ;
      RECT  93557.5 26257.5 93820.0 26322.5 ;
      RECT  93525.0 26290.0 93590.0 26565.0 ;
      RECT  93525.0 26497.5 93590.0 26632.5 ;
      RECT  93715.0 26497.5 93780.0 26632.5 ;
      RECT  93715.0 26497.5 93780.0 26632.5 ;
      RECT  93525.0 26497.5 93590.0 26632.5 ;
      RECT  93525.0 27357.5 93590.0 27492.5 ;
      RECT  93715.0 27357.5 93780.0 27492.5 ;
      RECT  93715.0 27357.5 93780.0 27492.5 ;
      RECT  93525.0 27357.5 93590.0 27492.5 ;
      RECT  93452.5 27772.5 93517.5 27907.5 ;
      RECT  93787.5 26222.5 93852.5 26357.5 ;
      RECT  93525.0 27357.5 93590.0 27492.5 ;
      RECT  93715.0 26497.5 93780.0 26632.5 ;
      RECT  93972.5 26397.5 94037.5 26532.5 ;
      RECT  93972.5 26397.5 94037.5 26532.5 ;
      RECT  94420.0 27807.5 94485.0 27872.5 ;
      RECT  94155.0 27807.5 94452.5 27872.5 ;
      RECT  94420.0 27425.0 94485.0 27840.0 ;
      RECT  94230.0 26257.5 94295.0 26322.5 ;
      RECT  94262.5 26257.5 94525.0 26322.5 ;
      RECT  94230.0 26290.0 94295.0 26565.0 ;
      RECT  94230.0 26497.5 94295.0 26632.5 ;
      RECT  94420.0 26497.5 94485.0 26632.5 ;
      RECT  94420.0 26497.5 94485.0 26632.5 ;
      RECT  94230.0 26497.5 94295.0 26632.5 ;
      RECT  94230.0 27357.5 94295.0 27492.5 ;
      RECT  94420.0 27357.5 94485.0 27492.5 ;
      RECT  94420.0 27357.5 94485.0 27492.5 ;
      RECT  94230.0 27357.5 94295.0 27492.5 ;
      RECT  94157.5 27772.5 94222.5 27907.5 ;
      RECT  94492.5 26222.5 94557.5 26357.5 ;
      RECT  94230.0 27357.5 94295.0 27492.5 ;
      RECT  94420.0 26497.5 94485.0 26632.5 ;
      RECT  94677.5 26397.5 94742.5 26532.5 ;
      RECT  94677.5 26397.5 94742.5 26532.5 ;
      RECT  95125.0 27807.5 95190.0 27872.5 ;
      RECT  94860.0 27807.5 95157.5 27872.5 ;
      RECT  95125.0 27425.0 95190.0 27840.0 ;
      RECT  94935.0 26257.5 95000.0 26322.5 ;
      RECT  94967.5 26257.5 95230.0 26322.5 ;
      RECT  94935.0 26290.0 95000.0 26565.0 ;
      RECT  94935.0 26497.5 95000.0 26632.5 ;
      RECT  95125.0 26497.5 95190.0 26632.5 ;
      RECT  95125.0 26497.5 95190.0 26632.5 ;
      RECT  94935.0 26497.5 95000.0 26632.5 ;
      RECT  94935.0 27357.5 95000.0 27492.5 ;
      RECT  95125.0 27357.5 95190.0 27492.5 ;
      RECT  95125.0 27357.5 95190.0 27492.5 ;
      RECT  94935.0 27357.5 95000.0 27492.5 ;
      RECT  94862.5 27772.5 94927.5 27907.5 ;
      RECT  95197.5 26222.5 95262.5 26357.5 ;
      RECT  94935.0 27357.5 95000.0 27492.5 ;
      RECT  95125.0 26497.5 95190.0 26632.5 ;
      RECT  95382.5 26397.5 95447.5 26532.5 ;
      RECT  95382.5 26397.5 95447.5 26532.5 ;
      RECT  95830.0 27807.5 95895.0 27872.5 ;
      RECT  95565.0 27807.5 95862.5 27872.5 ;
      RECT  95830.0 27425.0 95895.0 27840.0 ;
      RECT  95640.0 26257.5 95705.0 26322.5 ;
      RECT  95672.5 26257.5 95935.0 26322.5 ;
      RECT  95640.0 26290.0 95705.0 26565.0 ;
      RECT  95640.0 26497.5 95705.0 26632.5 ;
      RECT  95830.0 26497.5 95895.0 26632.5 ;
      RECT  95830.0 26497.5 95895.0 26632.5 ;
      RECT  95640.0 26497.5 95705.0 26632.5 ;
      RECT  95640.0 27357.5 95705.0 27492.5 ;
      RECT  95830.0 27357.5 95895.0 27492.5 ;
      RECT  95830.0 27357.5 95895.0 27492.5 ;
      RECT  95640.0 27357.5 95705.0 27492.5 ;
      RECT  95567.5 27772.5 95632.5 27907.5 ;
      RECT  95902.5 26222.5 95967.5 26357.5 ;
      RECT  95640.0 27357.5 95705.0 27492.5 ;
      RECT  95830.0 26497.5 95895.0 26632.5 ;
      RECT  96087.5 26397.5 96152.5 26532.5 ;
      RECT  96087.5 26397.5 96152.5 26532.5 ;
      RECT  96535.0 27807.5 96600.0 27872.5 ;
      RECT  96270.0 27807.5 96567.5 27872.5 ;
      RECT  96535.0 27425.0 96600.0 27840.0 ;
      RECT  96345.0 26257.5 96410.0 26322.5 ;
      RECT  96377.5 26257.5 96640.0 26322.5 ;
      RECT  96345.0 26290.0 96410.0 26565.0 ;
      RECT  96345.0 26497.5 96410.0 26632.5 ;
      RECT  96535.0 26497.5 96600.0 26632.5 ;
      RECT  96535.0 26497.5 96600.0 26632.5 ;
      RECT  96345.0 26497.5 96410.0 26632.5 ;
      RECT  96345.0 27357.5 96410.0 27492.5 ;
      RECT  96535.0 27357.5 96600.0 27492.5 ;
      RECT  96535.0 27357.5 96600.0 27492.5 ;
      RECT  96345.0 27357.5 96410.0 27492.5 ;
      RECT  96272.5 27772.5 96337.5 27907.5 ;
      RECT  96607.5 26222.5 96672.5 26357.5 ;
      RECT  96345.0 27357.5 96410.0 27492.5 ;
      RECT  96535.0 26497.5 96600.0 26632.5 ;
      RECT  96792.5 26397.5 96857.5 26532.5 ;
      RECT  96792.5 26397.5 96857.5 26532.5 ;
      RECT  97240.0 27807.5 97305.0 27872.5 ;
      RECT  96975.0 27807.5 97272.5 27872.5 ;
      RECT  97240.0 27425.0 97305.0 27840.0 ;
      RECT  97050.0 26257.5 97115.0 26322.5 ;
      RECT  97082.5 26257.5 97345.0 26322.5 ;
      RECT  97050.0 26290.0 97115.0 26565.0 ;
      RECT  97050.0 26497.5 97115.0 26632.5 ;
      RECT  97240.0 26497.5 97305.0 26632.5 ;
      RECT  97240.0 26497.5 97305.0 26632.5 ;
      RECT  97050.0 26497.5 97115.0 26632.5 ;
      RECT  97050.0 27357.5 97115.0 27492.5 ;
      RECT  97240.0 27357.5 97305.0 27492.5 ;
      RECT  97240.0 27357.5 97305.0 27492.5 ;
      RECT  97050.0 27357.5 97115.0 27492.5 ;
      RECT  96977.5 27772.5 97042.5 27907.5 ;
      RECT  97312.5 26222.5 97377.5 26357.5 ;
      RECT  97050.0 27357.5 97115.0 27492.5 ;
      RECT  97240.0 26497.5 97305.0 26632.5 ;
      RECT  97497.5 26397.5 97562.5 26532.5 ;
      RECT  97497.5 26397.5 97562.5 26532.5 ;
      RECT  97945.0 27807.5 98010.0 27872.5 ;
      RECT  97680.0 27807.5 97977.5 27872.5 ;
      RECT  97945.0 27425.0 98010.0 27840.0 ;
      RECT  97755.0 26257.5 97820.0 26322.5 ;
      RECT  97787.5 26257.5 98050.0 26322.5 ;
      RECT  97755.0 26290.0 97820.0 26565.0 ;
      RECT  97755.0 26497.5 97820.0 26632.5 ;
      RECT  97945.0 26497.5 98010.0 26632.5 ;
      RECT  97945.0 26497.5 98010.0 26632.5 ;
      RECT  97755.0 26497.5 97820.0 26632.5 ;
      RECT  97755.0 27357.5 97820.0 27492.5 ;
      RECT  97945.0 27357.5 98010.0 27492.5 ;
      RECT  97945.0 27357.5 98010.0 27492.5 ;
      RECT  97755.0 27357.5 97820.0 27492.5 ;
      RECT  97682.5 27772.5 97747.5 27907.5 ;
      RECT  98017.5 26222.5 98082.5 26357.5 ;
      RECT  97755.0 27357.5 97820.0 27492.5 ;
      RECT  97945.0 26497.5 98010.0 26632.5 ;
      RECT  98202.5 26397.5 98267.5 26532.5 ;
      RECT  98202.5 26397.5 98267.5 26532.5 ;
      RECT  98650.0 27807.5 98715.0 27872.5 ;
      RECT  98385.0 27807.5 98682.5 27872.5 ;
      RECT  98650.0 27425.0 98715.0 27840.0 ;
      RECT  98460.0 26257.5 98525.0 26322.5 ;
      RECT  98492.5 26257.5 98755.0 26322.5 ;
      RECT  98460.0 26290.0 98525.0 26565.0 ;
      RECT  98460.0 26497.5 98525.0 26632.5 ;
      RECT  98650.0 26497.5 98715.0 26632.5 ;
      RECT  98650.0 26497.5 98715.0 26632.5 ;
      RECT  98460.0 26497.5 98525.0 26632.5 ;
      RECT  98460.0 27357.5 98525.0 27492.5 ;
      RECT  98650.0 27357.5 98715.0 27492.5 ;
      RECT  98650.0 27357.5 98715.0 27492.5 ;
      RECT  98460.0 27357.5 98525.0 27492.5 ;
      RECT  98387.5 27772.5 98452.5 27907.5 ;
      RECT  98722.5 26222.5 98787.5 26357.5 ;
      RECT  98460.0 27357.5 98525.0 27492.5 ;
      RECT  98650.0 26497.5 98715.0 26632.5 ;
      RECT  98907.5 26397.5 98972.5 26532.5 ;
      RECT  98907.5 26397.5 98972.5 26532.5 ;
      RECT  99355.0 27807.5 99420.0 27872.5 ;
      RECT  99090.0 27807.5 99387.5 27872.5 ;
      RECT  99355.0 27425.0 99420.0 27840.0 ;
      RECT  99165.0 26257.5 99230.0 26322.5 ;
      RECT  99197.5 26257.5 99460.0 26322.5 ;
      RECT  99165.0 26290.0 99230.0 26565.0 ;
      RECT  99165.0 26497.5 99230.0 26632.5 ;
      RECT  99355.0 26497.5 99420.0 26632.5 ;
      RECT  99355.0 26497.5 99420.0 26632.5 ;
      RECT  99165.0 26497.5 99230.0 26632.5 ;
      RECT  99165.0 27357.5 99230.0 27492.5 ;
      RECT  99355.0 27357.5 99420.0 27492.5 ;
      RECT  99355.0 27357.5 99420.0 27492.5 ;
      RECT  99165.0 27357.5 99230.0 27492.5 ;
      RECT  99092.5 27772.5 99157.5 27907.5 ;
      RECT  99427.5 26222.5 99492.5 26357.5 ;
      RECT  99165.0 27357.5 99230.0 27492.5 ;
      RECT  99355.0 26497.5 99420.0 26632.5 ;
      RECT  99612.5 26397.5 99677.5 26532.5 ;
      RECT  99612.5 26397.5 99677.5 26532.5 ;
      RECT  100060.0 27807.5 100125.0 27872.5 ;
      RECT  99795.0 27807.5 100092.5 27872.5 ;
      RECT  100060.0 27425.0 100125.0 27840.0 ;
      RECT  99870.0 26257.5 99935.0 26322.5 ;
      RECT  99902.5 26257.5 100165.0 26322.5 ;
      RECT  99870.0 26290.0 99935.0 26565.0 ;
      RECT  99870.0 26497.5 99935.0 26632.5 ;
      RECT  100060.0 26497.5 100125.0 26632.5 ;
      RECT  100060.0 26497.5 100125.0 26632.5 ;
      RECT  99870.0 26497.5 99935.0 26632.5 ;
      RECT  99870.0 27357.5 99935.0 27492.5 ;
      RECT  100060.0 27357.5 100125.0 27492.5 ;
      RECT  100060.0 27357.5 100125.0 27492.5 ;
      RECT  99870.0 27357.5 99935.0 27492.5 ;
      RECT  99797.5 27772.5 99862.5 27907.5 ;
      RECT  100132.5 26222.5 100197.5 26357.5 ;
      RECT  99870.0 27357.5 99935.0 27492.5 ;
      RECT  100060.0 26497.5 100125.0 26632.5 ;
      RECT  100317.5 26397.5 100382.5 26532.5 ;
      RECT  100317.5 26397.5 100382.5 26532.5 ;
      RECT  100765.0 27807.5 100830.0 27872.5 ;
      RECT  100500.0 27807.5 100797.5 27872.5 ;
      RECT  100765.0 27425.0 100830.0 27840.0 ;
      RECT  100575.0 26257.5 100640.0 26322.5 ;
      RECT  100607.5 26257.5 100870.0 26322.5 ;
      RECT  100575.0 26290.0 100640.0 26565.0 ;
      RECT  100575.0 26497.5 100640.0 26632.5 ;
      RECT  100765.0 26497.5 100830.0 26632.5 ;
      RECT  100765.0 26497.5 100830.0 26632.5 ;
      RECT  100575.0 26497.5 100640.0 26632.5 ;
      RECT  100575.0 27357.5 100640.0 27492.5 ;
      RECT  100765.0 27357.5 100830.0 27492.5 ;
      RECT  100765.0 27357.5 100830.0 27492.5 ;
      RECT  100575.0 27357.5 100640.0 27492.5 ;
      RECT  100502.5 27772.5 100567.5 27907.5 ;
      RECT  100837.5 26222.5 100902.5 26357.5 ;
      RECT  100575.0 27357.5 100640.0 27492.5 ;
      RECT  100765.0 26497.5 100830.0 26632.5 ;
      RECT  101022.5 26397.5 101087.5 26532.5 ;
      RECT  101022.5 26397.5 101087.5 26532.5 ;
      RECT  101470.0 27807.5 101535.0 27872.5 ;
      RECT  101205.0 27807.5 101502.5 27872.5 ;
      RECT  101470.0 27425.0 101535.0 27840.0 ;
      RECT  101280.0 26257.5 101345.0 26322.5 ;
      RECT  101312.5 26257.5 101575.0 26322.5 ;
      RECT  101280.0 26290.0 101345.0 26565.0 ;
      RECT  101280.0 26497.5 101345.0 26632.5 ;
      RECT  101470.0 26497.5 101535.0 26632.5 ;
      RECT  101470.0 26497.5 101535.0 26632.5 ;
      RECT  101280.0 26497.5 101345.0 26632.5 ;
      RECT  101280.0 27357.5 101345.0 27492.5 ;
      RECT  101470.0 27357.5 101535.0 27492.5 ;
      RECT  101470.0 27357.5 101535.0 27492.5 ;
      RECT  101280.0 27357.5 101345.0 27492.5 ;
      RECT  101207.5 27772.5 101272.5 27907.5 ;
      RECT  101542.5 26222.5 101607.5 26357.5 ;
      RECT  101280.0 27357.5 101345.0 27492.5 ;
      RECT  101470.0 26497.5 101535.0 26632.5 ;
      RECT  101727.5 26397.5 101792.5 26532.5 ;
      RECT  101727.5 26397.5 101792.5 26532.5 ;
      RECT  102175.0 27807.5 102240.0 27872.5 ;
      RECT  101910.0 27807.5 102207.5 27872.5 ;
      RECT  102175.0 27425.0 102240.0 27840.0 ;
      RECT  101985.0 26257.5 102050.0 26322.5 ;
      RECT  102017.5 26257.5 102280.0 26322.5 ;
      RECT  101985.0 26290.0 102050.0 26565.0 ;
      RECT  101985.0 26497.5 102050.0 26632.5 ;
      RECT  102175.0 26497.5 102240.0 26632.5 ;
      RECT  102175.0 26497.5 102240.0 26632.5 ;
      RECT  101985.0 26497.5 102050.0 26632.5 ;
      RECT  101985.0 27357.5 102050.0 27492.5 ;
      RECT  102175.0 27357.5 102240.0 27492.5 ;
      RECT  102175.0 27357.5 102240.0 27492.5 ;
      RECT  101985.0 27357.5 102050.0 27492.5 ;
      RECT  101912.5 27772.5 101977.5 27907.5 ;
      RECT  102247.5 26222.5 102312.5 26357.5 ;
      RECT  101985.0 27357.5 102050.0 27492.5 ;
      RECT  102175.0 26497.5 102240.0 26632.5 ;
      RECT  102432.5 26397.5 102497.5 26532.5 ;
      RECT  102432.5 26397.5 102497.5 26532.5 ;
      RECT  102880.0 27807.5 102945.0 27872.5 ;
      RECT  102615.0 27807.5 102912.5 27872.5 ;
      RECT  102880.0 27425.0 102945.0 27840.0 ;
      RECT  102690.0 26257.5 102755.0 26322.5 ;
      RECT  102722.5 26257.5 102985.0 26322.5 ;
      RECT  102690.0 26290.0 102755.0 26565.0 ;
      RECT  102690.0 26497.5 102755.0 26632.5 ;
      RECT  102880.0 26497.5 102945.0 26632.5 ;
      RECT  102880.0 26497.5 102945.0 26632.5 ;
      RECT  102690.0 26497.5 102755.0 26632.5 ;
      RECT  102690.0 27357.5 102755.0 27492.5 ;
      RECT  102880.0 27357.5 102945.0 27492.5 ;
      RECT  102880.0 27357.5 102945.0 27492.5 ;
      RECT  102690.0 27357.5 102755.0 27492.5 ;
      RECT  102617.5 27772.5 102682.5 27907.5 ;
      RECT  102952.5 26222.5 103017.5 26357.5 ;
      RECT  102690.0 27357.5 102755.0 27492.5 ;
      RECT  102880.0 26497.5 102945.0 26632.5 ;
      RECT  103137.5 26397.5 103202.5 26532.5 ;
      RECT  103137.5 26397.5 103202.5 26532.5 ;
      RECT  103585.0 27807.5 103650.0 27872.5 ;
      RECT  103320.0 27807.5 103617.5 27872.5 ;
      RECT  103585.0 27425.0 103650.0 27840.0 ;
      RECT  103395.0 26257.5 103460.0 26322.5 ;
      RECT  103427.5 26257.5 103690.0 26322.5 ;
      RECT  103395.0 26290.0 103460.0 26565.0 ;
      RECT  103395.0 26497.5 103460.0 26632.5 ;
      RECT  103585.0 26497.5 103650.0 26632.5 ;
      RECT  103585.0 26497.5 103650.0 26632.5 ;
      RECT  103395.0 26497.5 103460.0 26632.5 ;
      RECT  103395.0 27357.5 103460.0 27492.5 ;
      RECT  103585.0 27357.5 103650.0 27492.5 ;
      RECT  103585.0 27357.5 103650.0 27492.5 ;
      RECT  103395.0 27357.5 103460.0 27492.5 ;
      RECT  103322.5 27772.5 103387.5 27907.5 ;
      RECT  103657.5 26222.5 103722.5 26357.5 ;
      RECT  103395.0 27357.5 103460.0 27492.5 ;
      RECT  103585.0 26497.5 103650.0 26632.5 ;
      RECT  103842.5 26397.5 103907.5 26532.5 ;
      RECT  103842.5 26397.5 103907.5 26532.5 ;
      RECT  104290.0 27807.5 104355.0 27872.5 ;
      RECT  104025.0 27807.5 104322.5 27872.5 ;
      RECT  104290.0 27425.0 104355.0 27840.0 ;
      RECT  104100.0 26257.5 104165.0 26322.5 ;
      RECT  104132.5 26257.5 104395.0 26322.5 ;
      RECT  104100.0 26290.0 104165.0 26565.0 ;
      RECT  104100.0 26497.5 104165.0 26632.5 ;
      RECT  104290.0 26497.5 104355.0 26632.5 ;
      RECT  104290.0 26497.5 104355.0 26632.5 ;
      RECT  104100.0 26497.5 104165.0 26632.5 ;
      RECT  104100.0 27357.5 104165.0 27492.5 ;
      RECT  104290.0 27357.5 104355.0 27492.5 ;
      RECT  104290.0 27357.5 104355.0 27492.5 ;
      RECT  104100.0 27357.5 104165.0 27492.5 ;
      RECT  104027.5 27772.5 104092.5 27907.5 ;
      RECT  104362.5 26222.5 104427.5 26357.5 ;
      RECT  104100.0 27357.5 104165.0 27492.5 ;
      RECT  104290.0 26497.5 104355.0 26632.5 ;
      RECT  104547.5 26397.5 104612.5 26532.5 ;
      RECT  104547.5 26397.5 104612.5 26532.5 ;
      RECT  104995.0 27807.5 105060.0 27872.5 ;
      RECT  104730.0 27807.5 105027.5 27872.5 ;
      RECT  104995.0 27425.0 105060.0 27840.0 ;
      RECT  104805.0 26257.5 104870.0 26322.5 ;
      RECT  104837.5 26257.5 105100.0 26322.5 ;
      RECT  104805.0 26290.0 104870.0 26565.0 ;
      RECT  104805.0 26497.5 104870.0 26632.5 ;
      RECT  104995.0 26497.5 105060.0 26632.5 ;
      RECT  104995.0 26497.5 105060.0 26632.5 ;
      RECT  104805.0 26497.5 104870.0 26632.5 ;
      RECT  104805.0 27357.5 104870.0 27492.5 ;
      RECT  104995.0 27357.5 105060.0 27492.5 ;
      RECT  104995.0 27357.5 105060.0 27492.5 ;
      RECT  104805.0 27357.5 104870.0 27492.5 ;
      RECT  104732.5 27772.5 104797.5 27907.5 ;
      RECT  105067.5 26222.5 105132.5 26357.5 ;
      RECT  104805.0 27357.5 104870.0 27492.5 ;
      RECT  104995.0 26497.5 105060.0 26632.5 ;
      RECT  105252.5 26397.5 105317.5 26532.5 ;
      RECT  105252.5 26397.5 105317.5 26532.5 ;
      RECT  105700.0 27807.5 105765.0 27872.5 ;
      RECT  105435.0 27807.5 105732.5 27872.5 ;
      RECT  105700.0 27425.0 105765.0 27840.0 ;
      RECT  105510.0 26257.5 105575.0 26322.5 ;
      RECT  105542.5 26257.5 105805.0 26322.5 ;
      RECT  105510.0 26290.0 105575.0 26565.0 ;
      RECT  105510.0 26497.5 105575.0 26632.5 ;
      RECT  105700.0 26497.5 105765.0 26632.5 ;
      RECT  105700.0 26497.5 105765.0 26632.5 ;
      RECT  105510.0 26497.5 105575.0 26632.5 ;
      RECT  105510.0 27357.5 105575.0 27492.5 ;
      RECT  105700.0 27357.5 105765.0 27492.5 ;
      RECT  105700.0 27357.5 105765.0 27492.5 ;
      RECT  105510.0 27357.5 105575.0 27492.5 ;
      RECT  105437.5 27772.5 105502.5 27907.5 ;
      RECT  105772.5 26222.5 105837.5 26357.5 ;
      RECT  105510.0 27357.5 105575.0 27492.5 ;
      RECT  105700.0 26497.5 105765.0 26632.5 ;
      RECT  105957.5 26397.5 106022.5 26532.5 ;
      RECT  105957.5 26397.5 106022.5 26532.5 ;
      RECT  16170.0 26012.5 16035.0 26077.5 ;
      RECT  16875.0 25872.5 16740.0 25937.5 ;
      RECT  17580.0 25732.5 17445.0 25797.5 ;
      RECT  18285.0 25592.5 18150.0 25657.5 ;
      RECT  18990.0 26012.5 18855.0 26077.5 ;
      RECT  19695.0 25872.5 19560.0 25937.5 ;
      RECT  20400.0 25732.5 20265.0 25797.5 ;
      RECT  21105.0 25592.5 20970.0 25657.5 ;
      RECT  21810.0 26012.5 21675.0 26077.5 ;
      RECT  22515.0 25872.5 22380.0 25937.5 ;
      RECT  23220.0 25732.5 23085.0 25797.5 ;
      RECT  23925.0 25592.5 23790.0 25657.5 ;
      RECT  24630.0 26012.5 24495.0 26077.5 ;
      RECT  25335.0 25872.5 25200.0 25937.5 ;
      RECT  26040.0 25732.5 25905.0 25797.5 ;
      RECT  26745.0 25592.5 26610.0 25657.5 ;
      RECT  27450.0 26012.5 27315.0 26077.5 ;
      RECT  28155.0 25872.5 28020.0 25937.5 ;
      RECT  28860.0 25732.5 28725.0 25797.5 ;
      RECT  29565.0 25592.5 29430.0 25657.5 ;
      RECT  30270.0 26012.5 30135.0 26077.5 ;
      RECT  30975.0 25872.5 30840.0 25937.5 ;
      RECT  31680.0 25732.5 31545.0 25797.5 ;
      RECT  32385.0 25592.5 32250.0 25657.5 ;
      RECT  33090.0 26012.5 32955.0 26077.5 ;
      RECT  33795.0 25872.5 33660.0 25937.5 ;
      RECT  34500.0 25732.5 34365.0 25797.5 ;
      RECT  35205.0 25592.5 35070.0 25657.5 ;
      RECT  35910.0 26012.5 35775.0 26077.5 ;
      RECT  36615.0 25872.5 36480.0 25937.5 ;
      RECT  37320.0 25732.5 37185.0 25797.5 ;
      RECT  38025.0 25592.5 37890.0 25657.5 ;
      RECT  38730.0 26012.5 38595.0 26077.5 ;
      RECT  39435.0 25872.5 39300.0 25937.5 ;
      RECT  40140.0 25732.5 40005.0 25797.5 ;
      RECT  40845.0 25592.5 40710.0 25657.5 ;
      RECT  41550.0 26012.5 41415.0 26077.5 ;
      RECT  42255.0 25872.5 42120.0 25937.5 ;
      RECT  42960.0 25732.5 42825.0 25797.5 ;
      RECT  43665.0 25592.5 43530.0 25657.5 ;
      RECT  44370.0 26012.5 44235.0 26077.5 ;
      RECT  45075.0 25872.5 44940.0 25937.5 ;
      RECT  45780.0 25732.5 45645.0 25797.5 ;
      RECT  46485.0 25592.5 46350.0 25657.5 ;
      RECT  47190.0 26012.5 47055.0 26077.5 ;
      RECT  47895.0 25872.5 47760.0 25937.5 ;
      RECT  48600.0 25732.5 48465.0 25797.5 ;
      RECT  49305.0 25592.5 49170.0 25657.5 ;
      RECT  50010.0 26012.5 49875.0 26077.5 ;
      RECT  50715.0 25872.5 50580.0 25937.5 ;
      RECT  51420.0 25732.5 51285.0 25797.5 ;
      RECT  52125.0 25592.5 51990.0 25657.5 ;
      RECT  52830.0 26012.5 52695.0 26077.5 ;
      RECT  53535.0 25872.5 53400.0 25937.5 ;
      RECT  54240.0 25732.5 54105.0 25797.5 ;
      RECT  54945.0 25592.5 54810.0 25657.5 ;
      RECT  55650.0 26012.5 55515.0 26077.5 ;
      RECT  56355.0 25872.5 56220.0 25937.5 ;
      RECT  57060.0 25732.5 56925.0 25797.5 ;
      RECT  57765.0 25592.5 57630.0 25657.5 ;
      RECT  58470.0 26012.5 58335.0 26077.5 ;
      RECT  59175.0 25872.5 59040.0 25937.5 ;
      RECT  59880.0 25732.5 59745.0 25797.5 ;
      RECT  60585.0 25592.5 60450.0 25657.5 ;
      RECT  61290.0 26012.5 61155.0 26077.5 ;
      RECT  61995.0 25872.5 61860.0 25937.5 ;
      RECT  62700.0 25732.5 62565.0 25797.5 ;
      RECT  63405.0 25592.5 63270.0 25657.5 ;
      RECT  64110.0 26012.5 63975.0 26077.5 ;
      RECT  64815.0 25872.5 64680.0 25937.5 ;
      RECT  65520.0 25732.5 65385.0 25797.5 ;
      RECT  66225.0 25592.5 66090.0 25657.5 ;
      RECT  66930.0 26012.5 66795.0 26077.5 ;
      RECT  67635.0 25872.5 67500.0 25937.5 ;
      RECT  68340.0 25732.5 68205.0 25797.5 ;
      RECT  69045.0 25592.5 68910.0 25657.5 ;
      RECT  69750.0 26012.5 69615.0 26077.5 ;
      RECT  70455.0 25872.5 70320.0 25937.5 ;
      RECT  71160.0 25732.5 71025.0 25797.5 ;
      RECT  71865.0 25592.5 71730.0 25657.5 ;
      RECT  72570.0 26012.5 72435.0 26077.5 ;
      RECT  73275.0 25872.5 73140.0 25937.5 ;
      RECT  73980.0 25732.5 73845.0 25797.5 ;
      RECT  74685.0 25592.5 74550.0 25657.5 ;
      RECT  75390.0 26012.5 75255.0 26077.5 ;
      RECT  76095.0 25872.5 75960.0 25937.5 ;
      RECT  76800.0 25732.5 76665.0 25797.5 ;
      RECT  77505.0 25592.5 77370.0 25657.5 ;
      RECT  78210.0 26012.5 78075.0 26077.5 ;
      RECT  78915.0 25872.5 78780.0 25937.5 ;
      RECT  79620.0 25732.5 79485.0 25797.5 ;
      RECT  80325.0 25592.5 80190.0 25657.5 ;
      RECT  81030.0 26012.5 80895.0 26077.5 ;
      RECT  81735.0 25872.5 81600.0 25937.5 ;
      RECT  82440.0 25732.5 82305.0 25797.5 ;
      RECT  83145.0 25592.5 83010.0 25657.5 ;
      RECT  83850.0 26012.5 83715.0 26077.5 ;
      RECT  84555.0 25872.5 84420.0 25937.5 ;
      RECT  85260.0 25732.5 85125.0 25797.5 ;
      RECT  85965.0 25592.5 85830.0 25657.5 ;
      RECT  86670.0 26012.5 86535.0 26077.5 ;
      RECT  87375.0 25872.5 87240.0 25937.5 ;
      RECT  88080.0 25732.5 87945.0 25797.5 ;
      RECT  88785.0 25592.5 88650.0 25657.5 ;
      RECT  89490.0 26012.5 89355.0 26077.5 ;
      RECT  90195.0 25872.5 90060.0 25937.5 ;
      RECT  90900.0 25732.5 90765.0 25797.5 ;
      RECT  91605.0 25592.5 91470.0 25657.5 ;
      RECT  92310.0 26012.5 92175.0 26077.5 ;
      RECT  93015.0 25872.5 92880.0 25937.5 ;
      RECT  93720.0 25732.5 93585.0 25797.5 ;
      RECT  94425.0 25592.5 94290.0 25657.5 ;
      RECT  95130.0 26012.5 94995.0 26077.5 ;
      RECT  95835.0 25872.5 95700.0 25937.5 ;
      RECT  96540.0 25732.5 96405.0 25797.5 ;
      RECT  97245.0 25592.5 97110.0 25657.5 ;
      RECT  97950.0 26012.5 97815.0 26077.5 ;
      RECT  98655.0 25872.5 98520.0 25937.5 ;
      RECT  99360.0 25732.5 99225.0 25797.5 ;
      RECT  100065.0 25592.5 99930.0 25657.5 ;
      RECT  100770.0 26012.5 100635.0 26077.5 ;
      RECT  101475.0 25872.5 101340.0 25937.5 ;
      RECT  102180.0 25732.5 102045.0 25797.5 ;
      RECT  102885.0 25592.5 102750.0 25657.5 ;
      RECT  103590.0 26012.5 103455.0 26077.5 ;
      RECT  104295.0 25872.5 104160.0 25937.5 ;
      RECT  105000.0 25732.5 104865.0 25797.5 ;
      RECT  105705.0 25592.5 105570.0 25657.5 ;
      RECT  16035.0 25452.5 15900.0 25517.5 ;
      RECT  16235.0 25312.5 16100.0 25377.5 ;
      RECT  16740.0 25452.5 16605.0 25517.5 ;
      RECT  16940.0 25312.5 16805.0 25377.5 ;
      RECT  17445.0 25452.5 17310.0 25517.5 ;
      RECT  17645.0 25312.5 17510.0 25377.5 ;
      RECT  18150.0 25452.5 18015.0 25517.5 ;
      RECT  18350.0 25312.5 18215.0 25377.5 ;
      RECT  18855.0 25452.5 18720.0 25517.5 ;
      RECT  19055.0 25312.5 18920.0 25377.5 ;
      RECT  19560.0 25452.5 19425.0 25517.5 ;
      RECT  19760.0 25312.5 19625.0 25377.5 ;
      RECT  20265.0 25452.5 20130.0 25517.5 ;
      RECT  20465.0 25312.5 20330.0 25377.5 ;
      RECT  20970.0 25452.5 20835.0 25517.5 ;
      RECT  21170.0 25312.5 21035.0 25377.5 ;
      RECT  21675.0 25452.5 21540.0 25517.5 ;
      RECT  21875.0 25312.5 21740.0 25377.5 ;
      RECT  22380.0 25452.5 22245.0 25517.5 ;
      RECT  22580.0 25312.5 22445.0 25377.5 ;
      RECT  23085.0 25452.5 22950.0 25517.5 ;
      RECT  23285.0 25312.5 23150.0 25377.5 ;
      RECT  23790.0 25452.5 23655.0 25517.5 ;
      RECT  23990.0 25312.5 23855.0 25377.5 ;
      RECT  24495.0 25452.5 24360.0 25517.5 ;
      RECT  24695.0 25312.5 24560.0 25377.5 ;
      RECT  25200.0 25452.5 25065.0 25517.5 ;
      RECT  25400.0 25312.5 25265.0 25377.5 ;
      RECT  25905.0 25452.5 25770.0 25517.5 ;
      RECT  26105.0 25312.5 25970.0 25377.5 ;
      RECT  26610.0 25452.5 26475.0 25517.5 ;
      RECT  26810.0 25312.5 26675.0 25377.5 ;
      RECT  27315.0 25452.5 27180.0 25517.5 ;
      RECT  27515.0 25312.5 27380.0 25377.5 ;
      RECT  28020.0 25452.5 27885.0 25517.5 ;
      RECT  28220.0 25312.5 28085.0 25377.5 ;
      RECT  28725.0 25452.5 28590.0 25517.5 ;
      RECT  28925.0 25312.5 28790.0 25377.5 ;
      RECT  29430.0 25452.5 29295.0 25517.5 ;
      RECT  29630.0 25312.5 29495.0 25377.5 ;
      RECT  30135.0 25452.5 30000.0 25517.5 ;
      RECT  30335.0 25312.5 30200.0 25377.5 ;
      RECT  30840.0 25452.5 30705.0 25517.5 ;
      RECT  31040.0 25312.5 30905.0 25377.5 ;
      RECT  31545.0 25452.5 31410.0 25517.5 ;
      RECT  31745.0 25312.5 31610.0 25377.5 ;
      RECT  32250.0 25452.5 32115.0 25517.5 ;
      RECT  32450.0 25312.5 32315.0 25377.5 ;
      RECT  32955.0 25452.5 32820.0 25517.5 ;
      RECT  33155.0 25312.5 33020.0 25377.5 ;
      RECT  33660.0 25452.5 33525.0 25517.5 ;
      RECT  33860.0 25312.5 33725.0 25377.5 ;
      RECT  34365.0 25452.5 34230.0 25517.5 ;
      RECT  34565.0 25312.5 34430.0 25377.5 ;
      RECT  35070.0 25452.5 34935.0 25517.5 ;
      RECT  35270.0 25312.5 35135.0 25377.5 ;
      RECT  35775.0 25452.5 35640.0 25517.5 ;
      RECT  35975.0 25312.5 35840.0 25377.5 ;
      RECT  36480.0 25452.5 36345.0 25517.5 ;
      RECT  36680.0 25312.5 36545.0 25377.5 ;
      RECT  37185.0 25452.5 37050.0 25517.5 ;
      RECT  37385.0 25312.5 37250.0 25377.5 ;
      RECT  37890.0 25452.5 37755.0 25517.5 ;
      RECT  38090.0 25312.5 37955.0 25377.5 ;
      RECT  38595.0 25452.5 38460.0 25517.5 ;
      RECT  38795.0 25312.5 38660.0 25377.5 ;
      RECT  39300.0 25452.5 39165.0 25517.5 ;
      RECT  39500.0 25312.5 39365.0 25377.5 ;
      RECT  40005.0 25452.5 39870.0 25517.5 ;
      RECT  40205.0 25312.5 40070.0 25377.5 ;
      RECT  40710.0 25452.5 40575.0 25517.5 ;
      RECT  40910.0 25312.5 40775.0 25377.5 ;
      RECT  41415.0 25452.5 41280.0 25517.5 ;
      RECT  41615.0 25312.5 41480.0 25377.5 ;
      RECT  42120.0 25452.5 41985.0 25517.5 ;
      RECT  42320.0 25312.5 42185.0 25377.5 ;
      RECT  42825.0 25452.5 42690.0 25517.5 ;
      RECT  43025.0 25312.5 42890.0 25377.5 ;
      RECT  43530.0 25452.5 43395.0 25517.5 ;
      RECT  43730.0 25312.5 43595.0 25377.5 ;
      RECT  44235.0 25452.5 44100.0 25517.5 ;
      RECT  44435.0 25312.5 44300.0 25377.5 ;
      RECT  44940.0 25452.5 44805.0 25517.5 ;
      RECT  45140.0 25312.5 45005.0 25377.5 ;
      RECT  45645.0 25452.5 45510.0 25517.5 ;
      RECT  45845.0 25312.5 45710.0 25377.5 ;
      RECT  46350.0 25452.5 46215.0 25517.5 ;
      RECT  46550.0 25312.5 46415.0 25377.5 ;
      RECT  47055.0 25452.5 46920.0 25517.5 ;
      RECT  47255.0 25312.5 47120.0 25377.5 ;
      RECT  47760.0 25452.5 47625.0 25517.5 ;
      RECT  47960.0 25312.5 47825.0 25377.5 ;
      RECT  48465.0 25452.5 48330.0 25517.5 ;
      RECT  48665.0 25312.5 48530.0 25377.5 ;
      RECT  49170.0 25452.5 49035.0 25517.5 ;
      RECT  49370.0 25312.5 49235.0 25377.5 ;
      RECT  49875.0 25452.5 49740.0 25517.5 ;
      RECT  50075.0 25312.5 49940.0 25377.5 ;
      RECT  50580.0 25452.5 50445.0 25517.5 ;
      RECT  50780.0 25312.5 50645.0 25377.5 ;
      RECT  51285.0 25452.5 51150.0 25517.5 ;
      RECT  51485.0 25312.5 51350.0 25377.5 ;
      RECT  51990.0 25452.5 51855.0 25517.5 ;
      RECT  52190.0 25312.5 52055.0 25377.5 ;
      RECT  52695.0 25452.5 52560.0 25517.5 ;
      RECT  52895.0 25312.5 52760.0 25377.5 ;
      RECT  53400.0 25452.5 53265.0 25517.5 ;
      RECT  53600.0 25312.5 53465.0 25377.5 ;
      RECT  54105.0 25452.5 53970.0 25517.5 ;
      RECT  54305.0 25312.5 54170.0 25377.5 ;
      RECT  54810.0 25452.5 54675.0 25517.5 ;
      RECT  55010.0 25312.5 54875.0 25377.5 ;
      RECT  55515.0 25452.5 55380.0 25517.5 ;
      RECT  55715.0 25312.5 55580.0 25377.5 ;
      RECT  56220.0 25452.5 56085.0 25517.5 ;
      RECT  56420.0 25312.5 56285.0 25377.5 ;
      RECT  56925.0 25452.5 56790.0 25517.5 ;
      RECT  57125.0 25312.5 56990.0 25377.5 ;
      RECT  57630.0 25452.5 57495.0 25517.5 ;
      RECT  57830.0 25312.5 57695.0 25377.5 ;
      RECT  58335.0 25452.5 58200.0 25517.5 ;
      RECT  58535.0 25312.5 58400.0 25377.5 ;
      RECT  59040.0 25452.5 58905.0 25517.5 ;
      RECT  59240.0 25312.5 59105.0 25377.5 ;
      RECT  59745.0 25452.5 59610.0 25517.5 ;
      RECT  59945.0 25312.5 59810.0 25377.5 ;
      RECT  60450.0 25452.5 60315.0 25517.5 ;
      RECT  60650.0 25312.5 60515.0 25377.5 ;
      RECT  61155.0 25452.5 61020.0 25517.5 ;
      RECT  61355.0 25312.5 61220.0 25377.5 ;
      RECT  61860.0 25452.5 61725.0 25517.5 ;
      RECT  62060.0 25312.5 61925.0 25377.5 ;
      RECT  62565.0 25452.5 62430.0 25517.5 ;
      RECT  62765.0 25312.5 62630.0 25377.5 ;
      RECT  63270.0 25452.5 63135.0 25517.5 ;
      RECT  63470.0 25312.5 63335.0 25377.5 ;
      RECT  63975.0 25452.5 63840.0 25517.5 ;
      RECT  64175.0 25312.5 64040.0 25377.5 ;
      RECT  64680.0 25452.5 64545.0 25517.5 ;
      RECT  64880.0 25312.5 64745.0 25377.5 ;
      RECT  65385.0 25452.5 65250.0 25517.5 ;
      RECT  65585.0 25312.5 65450.0 25377.5 ;
      RECT  66090.0 25452.5 65955.0 25517.5 ;
      RECT  66290.0 25312.5 66155.0 25377.5 ;
      RECT  66795.0 25452.5 66660.0 25517.5 ;
      RECT  66995.0 25312.5 66860.0 25377.5 ;
      RECT  67500.0 25452.5 67365.0 25517.5 ;
      RECT  67700.0 25312.5 67565.0 25377.5 ;
      RECT  68205.0 25452.5 68070.0 25517.5 ;
      RECT  68405.0 25312.5 68270.0 25377.5 ;
      RECT  68910.0 25452.5 68775.0 25517.5 ;
      RECT  69110.0 25312.5 68975.0 25377.5 ;
      RECT  69615.0 25452.5 69480.0 25517.5 ;
      RECT  69815.0 25312.5 69680.0 25377.5 ;
      RECT  70320.0 25452.5 70185.0 25517.5 ;
      RECT  70520.0 25312.5 70385.0 25377.5 ;
      RECT  71025.0 25452.5 70890.0 25517.5 ;
      RECT  71225.0 25312.5 71090.0 25377.5 ;
      RECT  71730.0 25452.5 71595.0 25517.5 ;
      RECT  71930.0 25312.5 71795.0 25377.5 ;
      RECT  72435.0 25452.5 72300.0 25517.5 ;
      RECT  72635.0 25312.5 72500.0 25377.5 ;
      RECT  73140.0 25452.5 73005.0 25517.5 ;
      RECT  73340.0 25312.5 73205.0 25377.5 ;
      RECT  73845.0 25452.5 73710.0 25517.5 ;
      RECT  74045.0 25312.5 73910.0 25377.5 ;
      RECT  74550.0 25452.5 74415.0 25517.5 ;
      RECT  74750.0 25312.5 74615.0 25377.5 ;
      RECT  75255.0 25452.5 75120.0 25517.5 ;
      RECT  75455.0 25312.5 75320.0 25377.5 ;
      RECT  75960.0 25452.5 75825.0 25517.5 ;
      RECT  76160.0 25312.5 76025.0 25377.5 ;
      RECT  76665.0 25452.5 76530.0 25517.5 ;
      RECT  76865.0 25312.5 76730.0 25377.5 ;
      RECT  77370.0 25452.5 77235.0 25517.5 ;
      RECT  77570.0 25312.5 77435.0 25377.5 ;
      RECT  78075.0 25452.5 77940.0 25517.5 ;
      RECT  78275.0 25312.5 78140.0 25377.5 ;
      RECT  78780.0 25452.5 78645.0 25517.5 ;
      RECT  78980.0 25312.5 78845.0 25377.5 ;
      RECT  79485.0 25452.5 79350.0 25517.5 ;
      RECT  79685.0 25312.5 79550.0 25377.5 ;
      RECT  80190.0 25452.5 80055.0 25517.5 ;
      RECT  80390.0 25312.5 80255.0 25377.5 ;
      RECT  80895.0 25452.5 80760.0 25517.5 ;
      RECT  81095.0 25312.5 80960.0 25377.5 ;
      RECT  81600.0 25452.5 81465.0 25517.5 ;
      RECT  81800.0 25312.5 81665.0 25377.5 ;
      RECT  82305.0 25452.5 82170.0 25517.5 ;
      RECT  82505.0 25312.5 82370.0 25377.5 ;
      RECT  83010.0 25452.5 82875.0 25517.5 ;
      RECT  83210.0 25312.5 83075.0 25377.5 ;
      RECT  83715.0 25452.5 83580.0 25517.5 ;
      RECT  83915.0 25312.5 83780.0 25377.5 ;
      RECT  84420.0 25452.5 84285.0 25517.5 ;
      RECT  84620.0 25312.5 84485.0 25377.5 ;
      RECT  85125.0 25452.5 84990.0 25517.5 ;
      RECT  85325.0 25312.5 85190.0 25377.5 ;
      RECT  85830.0 25452.5 85695.0 25517.5 ;
      RECT  86030.0 25312.5 85895.0 25377.5 ;
      RECT  86535.0 25452.5 86400.0 25517.5 ;
      RECT  86735.0 25312.5 86600.0 25377.5 ;
      RECT  87240.0 25452.5 87105.0 25517.5 ;
      RECT  87440.0 25312.5 87305.0 25377.5 ;
      RECT  87945.0 25452.5 87810.0 25517.5 ;
      RECT  88145.0 25312.5 88010.0 25377.5 ;
      RECT  88650.0 25452.5 88515.0 25517.5 ;
      RECT  88850.0 25312.5 88715.0 25377.5 ;
      RECT  89355.0 25452.5 89220.0 25517.5 ;
      RECT  89555.0 25312.5 89420.0 25377.5 ;
      RECT  90060.0 25452.5 89925.0 25517.5 ;
      RECT  90260.0 25312.5 90125.0 25377.5 ;
      RECT  90765.0 25452.5 90630.0 25517.5 ;
      RECT  90965.0 25312.5 90830.0 25377.5 ;
      RECT  91470.0 25452.5 91335.0 25517.5 ;
      RECT  91670.0 25312.5 91535.0 25377.5 ;
      RECT  92175.0 25452.5 92040.0 25517.5 ;
      RECT  92375.0 25312.5 92240.0 25377.5 ;
      RECT  92880.0 25452.5 92745.0 25517.5 ;
      RECT  93080.0 25312.5 92945.0 25377.5 ;
      RECT  93585.0 25452.5 93450.0 25517.5 ;
      RECT  93785.0 25312.5 93650.0 25377.5 ;
      RECT  94290.0 25452.5 94155.0 25517.5 ;
      RECT  94490.0 25312.5 94355.0 25377.5 ;
      RECT  94995.0 25452.5 94860.0 25517.5 ;
      RECT  95195.0 25312.5 95060.0 25377.5 ;
      RECT  95700.0 25452.5 95565.0 25517.5 ;
      RECT  95900.0 25312.5 95765.0 25377.5 ;
      RECT  96405.0 25452.5 96270.0 25517.5 ;
      RECT  96605.0 25312.5 96470.0 25377.5 ;
      RECT  97110.0 25452.5 96975.0 25517.5 ;
      RECT  97310.0 25312.5 97175.0 25377.5 ;
      RECT  97815.0 25452.5 97680.0 25517.5 ;
      RECT  98015.0 25312.5 97880.0 25377.5 ;
      RECT  98520.0 25452.5 98385.0 25517.5 ;
      RECT  98720.0 25312.5 98585.0 25377.5 ;
      RECT  99225.0 25452.5 99090.0 25517.5 ;
      RECT  99425.0 25312.5 99290.0 25377.5 ;
      RECT  99930.0 25452.5 99795.0 25517.5 ;
      RECT  100130.0 25312.5 99995.0 25377.5 ;
      RECT  100635.0 25452.5 100500.0 25517.5 ;
      RECT  100835.0 25312.5 100700.0 25377.5 ;
      RECT  101340.0 25452.5 101205.0 25517.5 ;
      RECT  101540.0 25312.5 101405.0 25377.5 ;
      RECT  102045.0 25452.5 101910.0 25517.5 ;
      RECT  102245.0 25312.5 102110.0 25377.5 ;
      RECT  102750.0 25452.5 102615.0 25517.5 ;
      RECT  102950.0 25312.5 102815.0 25377.5 ;
      RECT  103455.0 25452.5 103320.0 25517.5 ;
      RECT  103655.0 25312.5 103520.0 25377.5 ;
      RECT  104160.0 25452.5 104025.0 25517.5 ;
      RECT  104360.0 25312.5 104225.0 25377.5 ;
      RECT  104865.0 25452.5 104730.0 25517.5 ;
      RECT  105065.0 25312.5 104930.0 25377.5 ;
      RECT  105570.0 25452.5 105435.0 25517.5 ;
      RECT  105770.0 25312.5 105635.0 25377.5 ;
      RECT  15750.0 26010.0 105990.0 26080.0 ;
      RECT  15750.0 25870.0 105990.0 25940.0 ;
      RECT  15750.0 25730.0 105990.0 25800.0 ;
      RECT  15750.0 25590.0 105990.0 25660.0 ;
      RECT  7862.5 630.0 7927.5 695.0 ;
      RECT  7862.5 1152.5 7927.5 1217.5 ;
      RECT  7625.0 630.0 7895.0 695.0 ;
      RECT  7862.5 662.5 7927.5 1185.0 ;
      RECT  7895.0 1152.5 8140.0 1217.5 ;
      RECT  6755.0 630.0 7395.0 695.0 ;
      RECT  7862.5 2065.0 7927.5 2130.0 ;
      RECT  7862.5 2497.5 7927.5 2562.5 ;
      RECT  7625.0 2065.0 7895.0 2130.0 ;
      RECT  7862.5 2097.5 7927.5 2530.0 ;
      RECT  7895.0 2497.5 8415.0 2562.5 ;
      RECT  7030.0 2065.0 7395.0 2130.0 ;
      RECT  6755.0 2827.5 8690.0 2892.5 ;
      RECT  7030.0 4172.5 8965.0 4237.5 ;
      RECT  8140.0 642.5 9265.0 707.5 ;
      RECT  8415.0 427.5 9522.5 492.5 ;
      RECT  8690.0 2052.5 9265.0 2117.5 ;
      RECT  8415.0 2267.5 9522.5 2332.5 ;
      RECT  8140.0 3332.5 9265.0 3397.5 ;
      RECT  8965.0 3117.5 9522.5 3182.5 ;
      RECT  8690.0 4742.5 9265.0 4807.5 ;
      RECT  8965.0 4957.5 9522.5 5022.5 ;
      RECT  9970.0 642.5 10035.0 707.5 ;
      RECT  9970.0 630.0 10035.0 695.0 ;
      RECT  9752.5 642.5 10002.5 707.5 ;
      RECT  9970.0 662.5 10035.0 675.0 ;
      RECT  10002.5 630.0 10250.0 695.0 ;
      RECT  9970.0 2052.5 10035.0 2117.5 ;
      RECT  9970.0 2065.0 10035.0 2130.0 ;
      RECT  9752.5 2052.5 10002.5 2117.5 ;
      RECT  9970.0 2085.0 10035.0 2097.5 ;
      RECT  10002.5 2065.0 10250.0 2130.0 ;
      RECT  9970.0 3332.5 10035.0 3397.5 ;
      RECT  9970.0 3320.0 10035.0 3385.0 ;
      RECT  9752.5 3332.5 10002.5 3397.5 ;
      RECT  9970.0 3352.5 10035.0 3365.0 ;
      RECT  10002.5 3320.0 10250.0 3385.0 ;
      RECT  9970.0 4742.5 10035.0 4807.5 ;
      RECT  9970.0 4755.0 10035.0 4820.0 ;
      RECT  9752.5 4742.5 10002.5 4807.5 ;
      RECT  9970.0 4775.0 10035.0 4787.5 ;
      RECT  10002.5 4755.0 10250.0 4820.0 ;
      RECT  7697.5 1195.0 7762.5 1380.0 ;
      RECT  7697.5 35.0 7762.5 220.0 ;
      RECT  7337.5 152.5 7402.5 2.5 ;
      RECT  7337.5 1037.5 7402.5 1412.5 ;
      RECT  7527.5 152.5 7592.5 1037.5 ;
      RECT  7337.5 1037.5 7402.5 1172.5 ;
      RECT  7527.5 1037.5 7592.5 1172.5 ;
      RECT  7527.5 1037.5 7592.5 1172.5 ;
      RECT  7337.5 1037.5 7402.5 1172.5 ;
      RECT  7337.5 152.5 7402.5 287.5 ;
      RECT  7527.5 152.5 7592.5 287.5 ;
      RECT  7527.5 152.5 7592.5 287.5 ;
      RECT  7337.5 152.5 7402.5 287.5 ;
      RECT  7697.5 1127.5 7762.5 1262.5 ;
      RECT  7697.5 152.5 7762.5 287.5 ;
      RECT  7395.0 595.0 7460.0 730.0 ;
      RECT  7395.0 595.0 7460.0 730.0 ;
      RECT  7560.0 630.0 7625.0 695.0 ;
      RECT  7270.0 1347.5 7830.0 1412.5 ;
      RECT  7270.0 2.5 7830.0 67.5 ;
      RECT  7697.5 1565.0 7762.5 1380.0 ;
      RECT  7697.5 2725.0 7762.5 2540.0 ;
      RECT  7337.5 2607.5 7402.5 2757.5 ;
      RECT  7337.5 1722.5 7402.5 1347.5 ;
      RECT  7527.5 2607.5 7592.5 1722.5 ;
      RECT  7337.5 1722.5 7402.5 1587.5 ;
      RECT  7527.5 1722.5 7592.5 1587.5 ;
      RECT  7527.5 1722.5 7592.5 1587.5 ;
      RECT  7337.5 1722.5 7402.5 1587.5 ;
      RECT  7337.5 2607.5 7402.5 2472.5 ;
      RECT  7527.5 2607.5 7592.5 2472.5 ;
      RECT  7527.5 2607.5 7592.5 2472.5 ;
      RECT  7337.5 2607.5 7402.5 2472.5 ;
      RECT  7697.5 1632.5 7762.5 1497.5 ;
      RECT  7697.5 2607.5 7762.5 2472.5 ;
      RECT  7395.0 2165.0 7460.0 2030.0 ;
      RECT  7395.0 2165.0 7460.0 2030.0 ;
      RECT  7560.0 2130.0 7625.0 2065.0 ;
      RECT  7270.0 1412.5 7830.0 1347.5 ;
      RECT  7270.0 2757.5 7830.0 2692.5 ;
      RECT  10552.5 1195.0 10617.5 1380.0 ;
      RECT  10552.5 35.0 10617.5 220.0 ;
      RECT  10192.5 152.5 10257.5 2.5 ;
      RECT  10192.5 1037.5 10257.5 1412.5 ;
      RECT  10382.5 152.5 10447.5 1037.5 ;
      RECT  10192.5 1037.5 10257.5 1172.5 ;
      RECT  10382.5 1037.5 10447.5 1172.5 ;
      RECT  10382.5 1037.5 10447.5 1172.5 ;
      RECT  10192.5 1037.5 10257.5 1172.5 ;
      RECT  10192.5 152.5 10257.5 287.5 ;
      RECT  10382.5 152.5 10447.5 287.5 ;
      RECT  10382.5 152.5 10447.5 287.5 ;
      RECT  10192.5 152.5 10257.5 287.5 ;
      RECT  10552.5 1127.5 10617.5 1262.5 ;
      RECT  10552.5 152.5 10617.5 287.5 ;
      RECT  10250.0 595.0 10315.0 730.0 ;
      RECT  10250.0 595.0 10315.0 730.0 ;
      RECT  10415.0 630.0 10480.0 695.0 ;
      RECT  10125.0 1347.5 10685.0 1412.5 ;
      RECT  10125.0 2.5 10685.0 67.5 ;
      RECT  10552.5 1565.0 10617.5 1380.0 ;
      RECT  10552.5 2725.0 10617.5 2540.0 ;
      RECT  10192.5 2607.5 10257.5 2757.5 ;
      RECT  10192.5 1722.5 10257.5 1347.5 ;
      RECT  10382.5 2607.5 10447.5 1722.5 ;
      RECT  10192.5 1722.5 10257.5 1587.5 ;
      RECT  10382.5 1722.5 10447.5 1587.5 ;
      RECT  10382.5 1722.5 10447.5 1587.5 ;
      RECT  10192.5 1722.5 10257.5 1587.5 ;
      RECT  10192.5 2607.5 10257.5 2472.5 ;
      RECT  10382.5 2607.5 10447.5 2472.5 ;
      RECT  10382.5 2607.5 10447.5 2472.5 ;
      RECT  10192.5 2607.5 10257.5 2472.5 ;
      RECT  10552.5 1632.5 10617.5 1497.5 ;
      RECT  10552.5 2607.5 10617.5 2472.5 ;
      RECT  10250.0 2165.0 10315.0 2030.0 ;
      RECT  10250.0 2165.0 10315.0 2030.0 ;
      RECT  10415.0 2130.0 10480.0 2065.0 ;
      RECT  10125.0 1412.5 10685.0 1347.5 ;
      RECT  10125.0 2757.5 10685.0 2692.5 ;
      RECT  10552.5 3885.0 10617.5 4070.0 ;
      RECT  10552.5 2725.0 10617.5 2910.0 ;
      RECT  10192.5 2842.5 10257.5 2692.5 ;
      RECT  10192.5 3727.5 10257.5 4102.5 ;
      RECT  10382.5 2842.5 10447.5 3727.5 ;
      RECT  10192.5 3727.5 10257.5 3862.5 ;
      RECT  10382.5 3727.5 10447.5 3862.5 ;
      RECT  10382.5 3727.5 10447.5 3862.5 ;
      RECT  10192.5 3727.5 10257.5 3862.5 ;
      RECT  10192.5 2842.5 10257.5 2977.5 ;
      RECT  10382.5 2842.5 10447.5 2977.5 ;
      RECT  10382.5 2842.5 10447.5 2977.5 ;
      RECT  10192.5 2842.5 10257.5 2977.5 ;
      RECT  10552.5 3817.5 10617.5 3952.5 ;
      RECT  10552.5 2842.5 10617.5 2977.5 ;
      RECT  10250.0 3285.0 10315.0 3420.0 ;
      RECT  10250.0 3285.0 10315.0 3420.0 ;
      RECT  10415.0 3320.0 10480.0 3385.0 ;
      RECT  10125.0 4037.5 10685.0 4102.5 ;
      RECT  10125.0 2692.5 10685.0 2757.5 ;
      RECT  10552.5 4255.0 10617.5 4070.0 ;
      RECT  10552.5 5415.0 10617.5 5230.0 ;
      RECT  10192.5 5297.5 10257.5 5447.5 ;
      RECT  10192.5 4412.5 10257.5 4037.5 ;
      RECT  10382.5 5297.5 10447.5 4412.5 ;
      RECT  10192.5 4412.5 10257.5 4277.5 ;
      RECT  10382.5 4412.5 10447.5 4277.5 ;
      RECT  10382.5 4412.5 10447.5 4277.5 ;
      RECT  10192.5 4412.5 10257.5 4277.5 ;
      RECT  10192.5 5297.5 10257.5 5162.5 ;
      RECT  10382.5 5297.5 10447.5 5162.5 ;
      RECT  10382.5 5297.5 10447.5 5162.5 ;
      RECT  10192.5 5297.5 10257.5 5162.5 ;
      RECT  10552.5 4322.5 10617.5 4187.5 ;
      RECT  10552.5 5297.5 10617.5 5162.5 ;
      RECT  10250.0 4855.0 10315.0 4720.0 ;
      RECT  10250.0 4855.0 10315.0 4720.0 ;
      RECT  10415.0 4820.0 10480.0 4755.0 ;
      RECT  10125.0 4102.5 10685.0 4037.5 ;
      RECT  10125.0 5447.5 10685.0 5382.5 ;
      RECT  9272.5 197.5 9337.5 2.5 ;
      RECT  9272.5 1037.5 9337.5 1412.5 ;
      RECT  9652.5 1037.5 9717.5 1412.5 ;
      RECT  9822.5 1195.0 9887.5 1380.0 ;
      RECT  9822.5 35.0 9887.5 220.0 ;
      RECT  9272.5 1037.5 9337.5 1172.5 ;
      RECT  9462.5 1037.5 9527.5 1172.5 ;
      RECT  9462.5 1037.5 9527.5 1172.5 ;
      RECT  9272.5 1037.5 9337.5 1172.5 ;
      RECT  9462.5 1037.5 9527.5 1172.5 ;
      RECT  9652.5 1037.5 9717.5 1172.5 ;
      RECT  9652.5 1037.5 9717.5 1172.5 ;
      RECT  9462.5 1037.5 9527.5 1172.5 ;
      RECT  9272.5 197.5 9337.5 332.5 ;
      RECT  9462.5 197.5 9527.5 332.5 ;
      RECT  9462.5 197.5 9527.5 332.5 ;
      RECT  9272.5 197.5 9337.5 332.5 ;
      RECT  9462.5 197.5 9527.5 332.5 ;
      RECT  9652.5 197.5 9717.5 332.5 ;
      RECT  9652.5 197.5 9717.5 332.5 ;
      RECT  9462.5 197.5 9527.5 332.5 ;
      RECT  9822.5 1127.5 9887.5 1262.5 ;
      RECT  9822.5 152.5 9887.5 287.5 ;
      RECT  9657.5 427.5 9522.5 492.5 ;
      RECT  9400.0 642.5 9265.0 707.5 ;
      RECT  9462.5 1037.5 9527.5 1172.5 ;
      RECT  9652.5 197.5 9717.5 332.5 ;
      RECT  9752.5 642.5 9617.5 707.5 ;
      RECT  9265.0 642.5 9400.0 707.5 ;
      RECT  9522.5 427.5 9657.5 492.5 ;
      RECT  9617.5 642.5 9752.5 707.5 ;
      RECT  9205.0 1347.5 10125.0 1412.5 ;
      RECT  9205.0 2.5 10125.0 67.5 ;
      RECT  9272.5 2562.5 9337.5 2757.5 ;
      RECT  9272.5 1722.5 9337.5 1347.5 ;
      RECT  9652.5 1722.5 9717.5 1347.5 ;
      RECT  9822.5 1565.0 9887.5 1380.0 ;
      RECT  9822.5 2725.0 9887.5 2540.0 ;
      RECT  9272.5 1722.5 9337.5 1587.5 ;
      RECT  9462.5 1722.5 9527.5 1587.5 ;
      RECT  9462.5 1722.5 9527.5 1587.5 ;
      RECT  9272.5 1722.5 9337.5 1587.5 ;
      RECT  9462.5 1722.5 9527.5 1587.5 ;
      RECT  9652.5 1722.5 9717.5 1587.5 ;
      RECT  9652.5 1722.5 9717.5 1587.5 ;
      RECT  9462.5 1722.5 9527.5 1587.5 ;
      RECT  9272.5 2562.5 9337.5 2427.5 ;
      RECT  9462.5 2562.5 9527.5 2427.5 ;
      RECT  9462.5 2562.5 9527.5 2427.5 ;
      RECT  9272.5 2562.5 9337.5 2427.5 ;
      RECT  9462.5 2562.5 9527.5 2427.5 ;
      RECT  9652.5 2562.5 9717.5 2427.5 ;
      RECT  9652.5 2562.5 9717.5 2427.5 ;
      RECT  9462.5 2562.5 9527.5 2427.5 ;
      RECT  9822.5 1632.5 9887.5 1497.5 ;
      RECT  9822.5 2607.5 9887.5 2472.5 ;
      RECT  9657.5 2332.5 9522.5 2267.5 ;
      RECT  9400.0 2117.5 9265.0 2052.5 ;
      RECT  9462.5 1722.5 9527.5 1587.5 ;
      RECT  9652.5 2562.5 9717.5 2427.5 ;
      RECT  9752.5 2117.5 9617.5 2052.5 ;
      RECT  9265.0 2117.5 9400.0 2052.5 ;
      RECT  9522.5 2332.5 9657.5 2267.5 ;
      RECT  9617.5 2117.5 9752.5 2052.5 ;
      RECT  9205.0 1412.5 10125.0 1347.5 ;
      RECT  9205.0 2757.5 10125.0 2692.5 ;
      RECT  9272.5 2887.5 9337.5 2692.5 ;
      RECT  9272.5 3727.5 9337.5 4102.5 ;
      RECT  9652.5 3727.5 9717.5 4102.5 ;
      RECT  9822.5 3885.0 9887.5 4070.0 ;
      RECT  9822.5 2725.0 9887.5 2910.0 ;
      RECT  9272.5 3727.5 9337.5 3862.5 ;
      RECT  9462.5 3727.5 9527.5 3862.5 ;
      RECT  9462.5 3727.5 9527.5 3862.5 ;
      RECT  9272.5 3727.5 9337.5 3862.5 ;
      RECT  9462.5 3727.5 9527.5 3862.5 ;
      RECT  9652.5 3727.5 9717.5 3862.5 ;
      RECT  9652.5 3727.5 9717.5 3862.5 ;
      RECT  9462.5 3727.5 9527.5 3862.5 ;
      RECT  9272.5 2887.5 9337.5 3022.5 ;
      RECT  9462.5 2887.5 9527.5 3022.5 ;
      RECT  9462.5 2887.5 9527.5 3022.5 ;
      RECT  9272.5 2887.5 9337.5 3022.5 ;
      RECT  9462.5 2887.5 9527.5 3022.5 ;
      RECT  9652.5 2887.5 9717.5 3022.5 ;
      RECT  9652.5 2887.5 9717.5 3022.5 ;
      RECT  9462.5 2887.5 9527.5 3022.5 ;
      RECT  9822.5 3817.5 9887.5 3952.5 ;
      RECT  9822.5 2842.5 9887.5 2977.5 ;
      RECT  9657.5 3117.5 9522.5 3182.5 ;
      RECT  9400.0 3332.5 9265.0 3397.5 ;
      RECT  9462.5 3727.5 9527.5 3862.5 ;
      RECT  9652.5 2887.5 9717.5 3022.5 ;
      RECT  9752.5 3332.5 9617.5 3397.5 ;
      RECT  9265.0 3332.5 9400.0 3397.5 ;
      RECT  9522.5 3117.5 9657.5 3182.5 ;
      RECT  9617.5 3332.5 9752.5 3397.5 ;
      RECT  9205.0 4037.5 10125.0 4102.5 ;
      RECT  9205.0 2692.5 10125.0 2757.5 ;
      RECT  9272.5 5252.5 9337.5 5447.5 ;
      RECT  9272.5 4412.5 9337.5 4037.5 ;
      RECT  9652.5 4412.5 9717.5 4037.5 ;
      RECT  9822.5 4255.0 9887.5 4070.0 ;
      RECT  9822.5 5415.0 9887.5 5230.0 ;
      RECT  9272.5 4412.5 9337.5 4277.5 ;
      RECT  9462.5 4412.5 9527.5 4277.5 ;
      RECT  9462.5 4412.5 9527.5 4277.5 ;
      RECT  9272.5 4412.5 9337.5 4277.5 ;
      RECT  9462.5 4412.5 9527.5 4277.5 ;
      RECT  9652.5 4412.5 9717.5 4277.5 ;
      RECT  9652.5 4412.5 9717.5 4277.5 ;
      RECT  9462.5 4412.5 9527.5 4277.5 ;
      RECT  9272.5 5252.5 9337.5 5117.5 ;
      RECT  9462.5 5252.5 9527.5 5117.5 ;
      RECT  9462.5 5252.5 9527.5 5117.5 ;
      RECT  9272.5 5252.5 9337.5 5117.5 ;
      RECT  9462.5 5252.5 9527.5 5117.5 ;
      RECT  9652.5 5252.5 9717.5 5117.5 ;
      RECT  9652.5 5252.5 9717.5 5117.5 ;
      RECT  9462.5 5252.5 9527.5 5117.5 ;
      RECT  9822.5 4322.5 9887.5 4187.5 ;
      RECT  9822.5 5297.5 9887.5 5162.5 ;
      RECT  9657.5 5022.5 9522.5 4957.5 ;
      RECT  9400.0 4807.5 9265.0 4742.5 ;
      RECT  9462.5 4412.5 9527.5 4277.5 ;
      RECT  9652.5 5252.5 9717.5 5117.5 ;
      RECT  9752.5 4807.5 9617.5 4742.5 ;
      RECT  9265.0 4807.5 9400.0 4742.5 ;
      RECT  9522.5 5022.5 9657.5 4957.5 ;
      RECT  9617.5 4807.5 9752.5 4742.5 ;
      RECT  9205.0 4102.5 10125.0 4037.5 ;
      RECT  9205.0 5447.5 10125.0 5382.5 ;
      RECT  8207.5 1152.5 8072.5 1217.5 ;
      RECT  6822.5 630.0 6687.5 695.0 ;
      RECT  8482.5 2497.5 8347.5 2562.5 ;
      RECT  7097.5 2065.0 6962.5 2130.0 ;
      RECT  6822.5 2827.5 6687.5 2892.5 ;
      RECT  8757.5 2827.5 8622.5 2892.5 ;
      RECT  7097.5 4172.5 6962.5 4237.5 ;
      RECT  9032.5 4172.5 8897.5 4237.5 ;
      RECT  8207.5 642.5 8072.5 707.5 ;
      RECT  8482.5 427.5 8347.5 492.5 ;
      RECT  8757.5 2052.5 8622.5 2117.5 ;
      RECT  8482.5 2267.5 8347.5 2332.5 ;
      RECT  8207.5 3332.5 8072.5 3397.5 ;
      RECT  9032.5 3117.5 8897.5 3182.5 ;
      RECT  8757.5 4742.5 8622.5 4807.5 ;
      RECT  9032.5 4957.5 8897.5 5022.5 ;
      RECT  10480.0 630.0 10685.0 695.0 ;
      RECT  10480.0 2065.0 10685.0 2130.0 ;
      RECT  10480.0 3320.0 10685.0 3385.0 ;
      RECT  10480.0 4755.0 10685.0 4820.0 ;
      RECT  6720.0 1347.5 10685.0 1412.5 ;
      RECT  6720.0 4037.5 10685.0 4102.5 ;
      RECT  6720.0 2.5 10685.0 67.5 ;
      RECT  6720.0 2692.5 10685.0 2757.5 ;
      RECT  6720.0 5382.5 10685.0 5447.5 ;
      RECT  15750.0 20285.0 16455.0 25170.0 ;
      RECT  18570.0 20285.0 19275.0 25170.0 ;
      RECT  21390.0 20285.0 22095.0 25170.0 ;
      RECT  24210.0 20285.0 24915.0 25170.0 ;
      RECT  27030.0 20285.0 27735.0 25170.0 ;
      RECT  29850.0 20285.0 30555.0 25170.0 ;
      RECT  32670.0 20285.0 33375.0 25170.0 ;
      RECT  35490.0 20285.0 36195.0 25170.0 ;
      RECT  38310.0 20285.0 39015.0 25170.0 ;
      RECT  41130.0 20285.0 41835.0 25170.0 ;
      RECT  43950.0 20285.0 44655.0 25170.0 ;
      RECT  46770.0 20285.0 47475.0 25170.0 ;
      RECT  49590.0 20285.0 50295.0 25170.0 ;
      RECT  52410.0 20285.0 53115.0 25170.0 ;
      RECT  55230.0 20285.0 55935.0 25170.0 ;
      RECT  58050.0 20285.0 58755.0 25170.0 ;
      RECT  60870.0 20285.0 61575.0 25170.0 ;
      RECT  63690.0 20285.0 64395.0 25170.0 ;
      RECT  66510.0 20285.0 67215.0 25170.0 ;
      RECT  69330.0 20285.0 70035.0 25170.0 ;
      RECT  72150.0 20285.0 72855.0 25170.0 ;
      RECT  74970.0 20285.0 75675.0 25170.0 ;
      RECT  77790.0 20285.0 78495.0 25170.0 ;
      RECT  80610.0 20285.0 81315.0 25170.0 ;
      RECT  83430.0 20285.0 84135.0 25170.0 ;
      RECT  86250.0 20285.0 86955.0 25170.0 ;
      RECT  89070.0 20285.0 89775.0 25170.0 ;
      RECT  91890.0 20285.0 92595.0 25170.0 ;
      RECT  94710.0 20285.0 95415.0 25170.0 ;
      RECT  97530.0 20285.0 98235.0 25170.0 ;
      RECT  100350.0 20285.0 101055.0 25170.0 ;
      RECT  103170.0 20285.0 103875.0 25170.0 ;
      RECT  15750.0 20402.5 105990.0 20467.5 ;
      RECT  15750.0 24975.0 105990.0 25040.0 ;
      RECT  15750.0 20532.5 105990.0 20597.5 ;
      RECT  15750.0 16110.0 16455.0 20285.0 ;
      RECT  18570.0 16110.0 19275.0 20285.0 ;
      RECT  21390.0 16110.0 22095.0 20285.0 ;
      RECT  24210.0 16110.0 24915.0 20285.0 ;
      RECT  27030.0 16110.0 27735.0 20285.0 ;
      RECT  29850.0 16110.0 30555.0 20285.0 ;
      RECT  32670.0 16110.0 33375.0 20285.0 ;
      RECT  35490.0 16110.0 36195.0 20285.0 ;
      RECT  38310.0 16110.0 39015.0 20285.0 ;
      RECT  41130.0 16110.0 41835.0 20285.0 ;
      RECT  43950.0 16110.0 44655.0 20285.0 ;
      RECT  46770.0 16110.0 47475.0 20285.0 ;
      RECT  49590.0 16110.0 50295.0 20285.0 ;
      RECT  52410.0 16110.0 53115.0 20285.0 ;
      RECT  55230.0 16110.0 55935.0 20285.0 ;
      RECT  58050.0 16110.0 58755.0 20285.0 ;
      RECT  60870.0 16110.0 61575.0 20285.0 ;
      RECT  63690.0 16110.0 64395.0 20285.0 ;
      RECT  66510.0 16110.0 67215.0 20285.0 ;
      RECT  69330.0 16110.0 70035.0 20285.0 ;
      RECT  72150.0 16110.0 72855.0 20285.0 ;
      RECT  74970.0 16110.0 75675.0 20285.0 ;
      RECT  77790.0 16110.0 78495.0 20285.0 ;
      RECT  80610.0 16110.0 81315.0 20285.0 ;
      RECT  83430.0 16110.0 84135.0 20285.0 ;
      RECT  86250.0 16110.0 86955.0 20285.0 ;
      RECT  89070.0 16110.0 89775.0 20285.0 ;
      RECT  91890.0 16110.0 92595.0 20285.0 ;
      RECT  94710.0 16110.0 95415.0 20285.0 ;
      RECT  97530.0 16110.0 98235.0 20285.0 ;
      RECT  100350.0 16110.0 101055.0 20285.0 ;
      RECT  103170.0 16110.0 103875.0 20285.0 ;
      RECT  15750.0 16377.5 105990.0 16442.5 ;
      RECT  15750.0 16507.5 105990.0 16572.5 ;
      RECT  15750.0 17310.0 105990.0 17375.0 ;
      RECT  15750.0 9670.0 16455.0 16110.0 ;
      RECT  18570.0 9670.0 19275.0 16110.0 ;
      RECT  21390.0 9670.0 22095.0 16110.0 ;
      RECT  24210.0 9670.0 24915.0 16110.0 ;
      RECT  27030.0 9670.0 27735.0 16110.0 ;
      RECT  29850.0 9670.0 30555.0 16110.0 ;
      RECT  32670.0 9670.0 33375.0 16110.0 ;
      RECT  35490.0 9670.0 36195.0 16110.0 ;
      RECT  38310.0 9670.0 39015.0 16110.0 ;
      RECT  41130.0 9670.0 41835.0 16110.0 ;
      RECT  43950.0 9670.0 44655.0 16110.0 ;
      RECT  46770.0 9670.0 47475.0 16110.0 ;
      RECT  49590.0 9670.0 50295.0 16110.0 ;
      RECT  52410.0 9670.0 53115.0 16110.0 ;
      RECT  55230.0 9670.0 55935.0 16110.0 ;
      RECT  58050.0 9670.0 58755.0 16110.0 ;
      RECT  60870.0 9670.0 61575.0 16110.0 ;
      RECT  63690.0 9670.0 64395.0 16110.0 ;
      RECT  66510.0 9670.0 67215.0 16110.0 ;
      RECT  69330.0 9670.0 70035.0 16110.0 ;
      RECT  72150.0 9670.0 72855.0 16110.0 ;
      RECT  74970.0 9670.0 75675.0 16110.0 ;
      RECT  77790.0 9670.0 78495.0 16110.0 ;
      RECT  80610.0 9670.0 81315.0 16110.0 ;
      RECT  83430.0 9670.0 84135.0 16110.0 ;
      RECT  86250.0 9670.0 86955.0 16110.0 ;
      RECT  89070.0 9670.0 89775.0 16110.0 ;
      RECT  91890.0 9670.0 92595.0 16110.0 ;
      RECT  94710.0 9670.0 95415.0 16110.0 ;
      RECT  97530.0 9670.0 98235.0 16110.0 ;
      RECT  100350.0 9670.0 101055.0 16110.0 ;
      RECT  103170.0 9670.0 103875.0 16110.0 ;
      RECT  15750.0 9875.0 105990.0 9940.0 ;
      RECT  15750.0 12880.0 105990.0 12945.0 ;
      RECT  15750.0 15840.0 105990.0 15905.0 ;
      RECT  15750.0 10890.0 105990.0 10955.0 ;
      RECT  15750.0 13850.0 105990.0 13915.0 ;
      RECT  15750.0 10035.0 105990.0 10100.0 ;
      RECT  15750.0 9670.0 16455.0 6695.0 ;
      RECT  18570.0 9670.0 19275.0 6695.0 ;
      RECT  21390.0 9670.0 22095.0 6695.0 ;
      RECT  24210.0 9670.0 24915.0 6695.0 ;
      RECT  27030.0 9670.0 27735.0 6695.0 ;
      RECT  29850.0 9670.0 30555.0 6695.0 ;
      RECT  32670.0 9670.0 33375.0 6695.0 ;
      RECT  35490.0 9670.0 36195.0 6695.0 ;
      RECT  38310.0 9670.0 39015.0 6695.0 ;
      RECT  41130.0 9670.0 41835.0 6695.0 ;
      RECT  43950.0 9670.0 44655.0 6695.0 ;
      RECT  46770.0 9670.0 47475.0 6695.0 ;
      RECT  49590.0 9670.0 50295.0 6695.0 ;
      RECT  52410.0 9670.0 53115.0 6695.0 ;
      RECT  55230.0 9670.0 55935.0 6695.0 ;
      RECT  58050.0 9670.0 58755.0 6695.0 ;
      RECT  60870.0 9670.0 61575.0 6695.0 ;
      RECT  63690.0 9670.0 64395.0 6695.0 ;
      RECT  66510.0 9670.0 67215.0 6695.0 ;
      RECT  69330.0 9670.0 70035.0 6695.0 ;
      RECT  72150.0 9670.0 72855.0 6695.0 ;
      RECT  74970.0 9670.0 75675.0 6695.0 ;
      RECT  77790.0 9670.0 78495.0 6695.0 ;
      RECT  80610.0 9670.0 81315.0 6695.0 ;
      RECT  83430.0 9670.0 84135.0 6695.0 ;
      RECT  86250.0 9670.0 86955.0 6695.0 ;
      RECT  89070.0 9670.0 89775.0 6695.0 ;
      RECT  91890.0 9670.0 92595.0 6695.0 ;
      RECT  94710.0 9670.0 95415.0 6695.0 ;
      RECT  97530.0 9670.0 98235.0 6695.0 ;
      RECT  100350.0 9670.0 101055.0 6695.0 ;
      RECT  103170.0 9670.0 103875.0 6695.0 ;
      RECT  15750.0 9302.5 103875.0 9237.5 ;
      RECT  15750.0 7755.0 103875.0 7690.0 ;
      RECT  15750.0 7885.0 103875.0 7820.0 ;
      RECT  15750.0 9172.5 103875.0 9107.5 ;
      RECT  8017.5 28670.0 8082.5 28735.0 ;
      RECT  8017.5 28610.0 8082.5 28675.0 ;
      RECT  7832.5 28670.0 8050.0 28735.0 ;
      RECT  8017.5 28642.5 8082.5 28702.5 ;
      RECT  8050.0 28610.0 8265.0 28675.0 ;
      RECT  8017.5 29985.0 8082.5 30050.0 ;
      RECT  8017.5 30045.0 8082.5 30110.0 ;
      RECT  7832.5 29985.0 8050.0 30050.0 ;
      RECT  8017.5 30017.5 8082.5 30077.5 ;
      RECT  8050.0 30045.0 8265.0 30110.0 ;
      RECT  8017.5 31360.0 8082.5 31425.0 ;
      RECT  8017.5 31300.0 8082.5 31365.0 ;
      RECT  7832.5 31360.0 8050.0 31425.0 ;
      RECT  8017.5 31332.5 8082.5 31392.5 ;
      RECT  8050.0 31300.0 8265.0 31365.0 ;
      RECT  8017.5 32675.0 8082.5 32740.0 ;
      RECT  8017.5 32735.0 8082.5 32800.0 ;
      RECT  7832.5 32675.0 8050.0 32740.0 ;
      RECT  8017.5 32707.5 8082.5 32767.5 ;
      RECT  8050.0 32735.0 8265.0 32800.0 ;
      RECT  8017.5 34050.0 8082.5 34115.0 ;
      RECT  8017.5 33990.0 8082.5 34055.0 ;
      RECT  7832.5 34050.0 8050.0 34115.0 ;
      RECT  8017.5 34022.5 8082.5 34082.5 ;
      RECT  8050.0 33990.0 8265.0 34055.0 ;
      RECT  8017.5 35365.0 8082.5 35430.0 ;
      RECT  8017.5 35425.0 8082.5 35490.0 ;
      RECT  7832.5 35365.0 8050.0 35430.0 ;
      RECT  8017.5 35397.5 8082.5 35457.5 ;
      RECT  8050.0 35425.0 8265.0 35490.0 ;
      RECT  8017.5 36740.0 8082.5 36805.0 ;
      RECT  8017.5 36680.0 8082.5 36745.0 ;
      RECT  7832.5 36740.0 8050.0 36805.0 ;
      RECT  8017.5 36712.5 8082.5 36772.5 ;
      RECT  8050.0 36680.0 8265.0 36745.0 ;
      RECT  8017.5 38055.0 8082.5 38120.0 ;
      RECT  8017.5 38115.0 8082.5 38180.0 ;
      RECT  7832.5 38055.0 8050.0 38120.0 ;
      RECT  8017.5 38087.5 8082.5 38147.5 ;
      RECT  8050.0 38115.0 8265.0 38180.0 ;
      RECT  8017.5 39430.0 8082.5 39495.0 ;
      RECT  8017.5 39370.0 8082.5 39435.0 ;
      RECT  7832.5 39430.0 8050.0 39495.0 ;
      RECT  8017.5 39402.5 8082.5 39462.5 ;
      RECT  8050.0 39370.0 8265.0 39435.0 ;
      RECT  8017.5 40745.0 8082.5 40810.0 ;
      RECT  8017.5 40805.0 8082.5 40870.0 ;
      RECT  7832.5 40745.0 8050.0 40810.0 ;
      RECT  8017.5 40777.5 8082.5 40837.5 ;
      RECT  8050.0 40805.0 8265.0 40870.0 ;
      RECT  8017.5 42120.0 8082.5 42185.0 ;
      RECT  8017.5 42060.0 8082.5 42125.0 ;
      RECT  7832.5 42120.0 8050.0 42185.0 ;
      RECT  8017.5 42092.5 8082.5 42152.5 ;
      RECT  8050.0 42060.0 8265.0 42125.0 ;
      RECT  8017.5 43435.0 8082.5 43500.0 ;
      RECT  8017.5 43495.0 8082.5 43560.0 ;
      RECT  7832.5 43435.0 8050.0 43500.0 ;
      RECT  8017.5 43467.5 8082.5 43527.5 ;
      RECT  8050.0 43495.0 8265.0 43560.0 ;
      RECT  8017.5 44810.0 8082.5 44875.0 ;
      RECT  8017.5 44750.0 8082.5 44815.0 ;
      RECT  7832.5 44810.0 8050.0 44875.0 ;
      RECT  8017.5 44782.5 8082.5 44842.5 ;
      RECT  8050.0 44750.0 8265.0 44815.0 ;
      RECT  8017.5 46125.0 8082.5 46190.0 ;
      RECT  8017.5 46185.0 8082.5 46250.0 ;
      RECT  7832.5 46125.0 8050.0 46190.0 ;
      RECT  8017.5 46157.5 8082.5 46217.5 ;
      RECT  8050.0 46185.0 8265.0 46250.0 ;
      RECT  8017.5 47500.0 8082.5 47565.0 ;
      RECT  8017.5 47440.0 8082.5 47505.0 ;
      RECT  7832.5 47500.0 8050.0 47565.0 ;
      RECT  8017.5 47472.5 8082.5 47532.5 ;
      RECT  8050.0 47440.0 8265.0 47505.0 ;
      RECT  8017.5 48815.0 8082.5 48880.0 ;
      RECT  8017.5 48875.0 8082.5 48940.0 ;
      RECT  7832.5 48815.0 8050.0 48880.0 ;
      RECT  8017.5 48847.5 8082.5 48907.5 ;
      RECT  8050.0 48875.0 8265.0 48940.0 ;
      RECT  8017.5 50190.0 8082.5 50255.0 ;
      RECT  8017.5 50130.0 8082.5 50195.0 ;
      RECT  7832.5 50190.0 8050.0 50255.0 ;
      RECT  8017.5 50162.5 8082.5 50222.5 ;
      RECT  8050.0 50130.0 8265.0 50195.0 ;
      RECT  8017.5 51505.0 8082.5 51570.0 ;
      RECT  8017.5 51565.0 8082.5 51630.0 ;
      RECT  7832.5 51505.0 8050.0 51570.0 ;
      RECT  8017.5 51537.5 8082.5 51597.5 ;
      RECT  8050.0 51565.0 8265.0 51630.0 ;
      RECT  8017.5 52880.0 8082.5 52945.0 ;
      RECT  8017.5 52820.0 8082.5 52885.0 ;
      RECT  7832.5 52880.0 8050.0 52945.0 ;
      RECT  8017.5 52852.5 8082.5 52912.5 ;
      RECT  8050.0 52820.0 8265.0 52885.0 ;
      RECT  8017.5 54195.0 8082.5 54260.0 ;
      RECT  8017.5 54255.0 8082.5 54320.0 ;
      RECT  7832.5 54195.0 8050.0 54260.0 ;
      RECT  8017.5 54227.5 8082.5 54287.5 ;
      RECT  8050.0 54255.0 8265.0 54320.0 ;
      RECT  8017.5 55570.0 8082.5 55635.0 ;
      RECT  8017.5 55510.0 8082.5 55575.0 ;
      RECT  7832.5 55570.0 8050.0 55635.0 ;
      RECT  8017.5 55542.5 8082.5 55602.5 ;
      RECT  8050.0 55510.0 8265.0 55575.0 ;
      RECT  8017.5 56885.0 8082.5 56950.0 ;
      RECT  8017.5 56945.0 8082.5 57010.0 ;
      RECT  7832.5 56885.0 8050.0 56950.0 ;
      RECT  8017.5 56917.5 8082.5 56977.5 ;
      RECT  8050.0 56945.0 8265.0 57010.0 ;
      RECT  8017.5 58260.0 8082.5 58325.0 ;
      RECT  8017.5 58200.0 8082.5 58265.0 ;
      RECT  7832.5 58260.0 8050.0 58325.0 ;
      RECT  8017.5 58232.5 8082.5 58292.5 ;
      RECT  8050.0 58200.0 8265.0 58265.0 ;
      RECT  8017.5 59575.0 8082.5 59640.0 ;
      RECT  8017.5 59635.0 8082.5 59700.0 ;
      RECT  7832.5 59575.0 8050.0 59640.0 ;
      RECT  8017.5 59607.5 8082.5 59667.5 ;
      RECT  8050.0 59635.0 8265.0 59700.0 ;
      RECT  8017.5 60950.0 8082.5 61015.0 ;
      RECT  8017.5 60890.0 8082.5 60955.0 ;
      RECT  7832.5 60950.0 8050.0 61015.0 ;
      RECT  8017.5 60922.5 8082.5 60982.5 ;
      RECT  8050.0 60890.0 8265.0 60955.0 ;
      RECT  8017.5 62265.0 8082.5 62330.0 ;
      RECT  8017.5 62325.0 8082.5 62390.0 ;
      RECT  7832.5 62265.0 8050.0 62330.0 ;
      RECT  8017.5 62297.5 8082.5 62357.5 ;
      RECT  8050.0 62325.0 8265.0 62390.0 ;
      RECT  8017.5 63640.0 8082.5 63705.0 ;
      RECT  8017.5 63580.0 8082.5 63645.0 ;
      RECT  7832.5 63640.0 8050.0 63705.0 ;
      RECT  8017.5 63612.5 8082.5 63672.5 ;
      RECT  8050.0 63580.0 8265.0 63645.0 ;
      RECT  8017.5 64955.0 8082.5 65020.0 ;
      RECT  8017.5 65015.0 8082.5 65080.0 ;
      RECT  7832.5 64955.0 8050.0 65020.0 ;
      RECT  8017.5 64987.5 8082.5 65047.5 ;
      RECT  8050.0 65015.0 8265.0 65080.0 ;
      RECT  8017.5 66330.0 8082.5 66395.0 ;
      RECT  8017.5 66270.0 8082.5 66335.0 ;
      RECT  7832.5 66330.0 8050.0 66395.0 ;
      RECT  8017.5 66302.5 8082.5 66362.5 ;
      RECT  8050.0 66270.0 8265.0 66335.0 ;
      RECT  8017.5 67645.0 8082.5 67710.0 ;
      RECT  8017.5 67705.0 8082.5 67770.0 ;
      RECT  7832.5 67645.0 8050.0 67710.0 ;
      RECT  8017.5 67677.5 8082.5 67737.5 ;
      RECT  8050.0 67705.0 8265.0 67770.0 ;
      RECT  8017.5 69020.0 8082.5 69085.0 ;
      RECT  8017.5 68960.0 8082.5 69025.0 ;
      RECT  7832.5 69020.0 8050.0 69085.0 ;
      RECT  8017.5 68992.5 8082.5 69052.5 ;
      RECT  8050.0 68960.0 8265.0 69025.0 ;
      RECT  8017.5 70335.0 8082.5 70400.0 ;
      RECT  8017.5 70395.0 8082.5 70460.0 ;
      RECT  7832.5 70335.0 8050.0 70400.0 ;
      RECT  8017.5 70367.5 8082.5 70427.5 ;
      RECT  8050.0 70395.0 8265.0 70460.0 ;
      RECT  8017.5 71710.0 8082.5 71775.0 ;
      RECT  8017.5 71650.0 8082.5 71715.0 ;
      RECT  7832.5 71710.0 8050.0 71775.0 ;
      RECT  8017.5 71682.5 8082.5 71742.5 ;
      RECT  8050.0 71650.0 8265.0 71715.0 ;
      RECT  8017.5 73025.0 8082.5 73090.0 ;
      RECT  8017.5 73085.0 8082.5 73150.0 ;
      RECT  7832.5 73025.0 8050.0 73090.0 ;
      RECT  8017.5 73057.5 8082.5 73117.5 ;
      RECT  8050.0 73085.0 8265.0 73150.0 ;
      RECT  8017.5 74400.0 8082.5 74465.0 ;
      RECT  8017.5 74340.0 8082.5 74405.0 ;
      RECT  7832.5 74400.0 8050.0 74465.0 ;
      RECT  8017.5 74372.5 8082.5 74432.5 ;
      RECT  8050.0 74340.0 8265.0 74405.0 ;
      RECT  8017.5 75715.0 8082.5 75780.0 ;
      RECT  8017.5 75775.0 8082.5 75840.0 ;
      RECT  7832.5 75715.0 8050.0 75780.0 ;
      RECT  8017.5 75747.5 8082.5 75807.5 ;
      RECT  8050.0 75775.0 8265.0 75840.0 ;
      RECT  8017.5 77090.0 8082.5 77155.0 ;
      RECT  8017.5 77030.0 8082.5 77095.0 ;
      RECT  7832.5 77090.0 8050.0 77155.0 ;
      RECT  8017.5 77062.5 8082.5 77122.5 ;
      RECT  8050.0 77030.0 8265.0 77095.0 ;
      RECT  8017.5 78405.0 8082.5 78470.0 ;
      RECT  8017.5 78465.0 8082.5 78530.0 ;
      RECT  7832.5 78405.0 8050.0 78470.0 ;
      RECT  8017.5 78437.5 8082.5 78497.5 ;
      RECT  8050.0 78465.0 8265.0 78530.0 ;
      RECT  8017.5 79780.0 8082.5 79845.0 ;
      RECT  8017.5 79720.0 8082.5 79785.0 ;
      RECT  7832.5 79780.0 8050.0 79845.0 ;
      RECT  8017.5 79752.5 8082.5 79812.5 ;
      RECT  8050.0 79720.0 8265.0 79785.0 ;
      RECT  8017.5 81095.0 8082.5 81160.0 ;
      RECT  8017.5 81155.0 8082.5 81220.0 ;
      RECT  7832.5 81095.0 8050.0 81160.0 ;
      RECT  8017.5 81127.5 8082.5 81187.5 ;
      RECT  8050.0 81155.0 8265.0 81220.0 ;
      RECT  8017.5 82470.0 8082.5 82535.0 ;
      RECT  8017.5 82410.0 8082.5 82475.0 ;
      RECT  7832.5 82470.0 8050.0 82535.0 ;
      RECT  8017.5 82442.5 8082.5 82502.5 ;
      RECT  8050.0 82410.0 8265.0 82475.0 ;
      RECT  8017.5 83785.0 8082.5 83850.0 ;
      RECT  8017.5 83845.0 8082.5 83910.0 ;
      RECT  7832.5 83785.0 8050.0 83850.0 ;
      RECT  8017.5 83817.5 8082.5 83877.5 ;
      RECT  8050.0 83845.0 8265.0 83910.0 ;
      RECT  8017.5 85160.0 8082.5 85225.0 ;
      RECT  8017.5 85100.0 8082.5 85165.0 ;
      RECT  7832.5 85160.0 8050.0 85225.0 ;
      RECT  8017.5 85132.5 8082.5 85192.5 ;
      RECT  8050.0 85100.0 8265.0 85165.0 ;
      RECT  8017.5 86475.0 8082.5 86540.0 ;
      RECT  8017.5 86535.0 8082.5 86600.0 ;
      RECT  7832.5 86475.0 8050.0 86540.0 ;
      RECT  8017.5 86507.5 8082.5 86567.5 ;
      RECT  8050.0 86535.0 8265.0 86600.0 ;
      RECT  8017.5 87850.0 8082.5 87915.0 ;
      RECT  8017.5 87790.0 8082.5 87855.0 ;
      RECT  7832.5 87850.0 8050.0 87915.0 ;
      RECT  8017.5 87822.5 8082.5 87882.5 ;
      RECT  8050.0 87790.0 8265.0 87855.0 ;
      RECT  8017.5 89165.0 8082.5 89230.0 ;
      RECT  8017.5 89225.0 8082.5 89290.0 ;
      RECT  7832.5 89165.0 8050.0 89230.0 ;
      RECT  8017.5 89197.5 8082.5 89257.5 ;
      RECT  8050.0 89225.0 8265.0 89290.0 ;
      RECT  8017.5 90540.0 8082.5 90605.0 ;
      RECT  8017.5 90480.0 8082.5 90545.0 ;
      RECT  7832.5 90540.0 8050.0 90605.0 ;
      RECT  8017.5 90512.5 8082.5 90572.5 ;
      RECT  8050.0 90480.0 8265.0 90545.0 ;
      RECT  8017.5 91855.0 8082.5 91920.0 ;
      RECT  8017.5 91915.0 8082.5 91980.0 ;
      RECT  7832.5 91855.0 8050.0 91920.0 ;
      RECT  8017.5 91887.5 8082.5 91947.5 ;
      RECT  8050.0 91915.0 8265.0 91980.0 ;
      RECT  8017.5 93230.0 8082.5 93295.0 ;
      RECT  8017.5 93170.0 8082.5 93235.0 ;
      RECT  7832.5 93230.0 8050.0 93295.0 ;
      RECT  8017.5 93202.5 8082.5 93262.5 ;
      RECT  8050.0 93170.0 8265.0 93235.0 ;
      RECT  8017.5 94545.0 8082.5 94610.0 ;
      RECT  8017.5 94605.0 8082.5 94670.0 ;
      RECT  7832.5 94545.0 8050.0 94610.0 ;
      RECT  8017.5 94577.5 8082.5 94637.5 ;
      RECT  8050.0 94605.0 8265.0 94670.0 ;
      RECT  8017.5 95920.0 8082.5 95985.0 ;
      RECT  8017.5 95860.0 8082.5 95925.0 ;
      RECT  7832.5 95920.0 8050.0 95985.0 ;
      RECT  8017.5 95892.5 8082.5 95952.5 ;
      RECT  8050.0 95860.0 8265.0 95925.0 ;
      RECT  8017.5 97235.0 8082.5 97300.0 ;
      RECT  8017.5 97295.0 8082.5 97360.0 ;
      RECT  7832.5 97235.0 8050.0 97300.0 ;
      RECT  8017.5 97267.5 8082.5 97327.5 ;
      RECT  8050.0 97295.0 8265.0 97360.0 ;
      RECT  8017.5 98610.0 8082.5 98675.0 ;
      RECT  8017.5 98550.0 8082.5 98615.0 ;
      RECT  7832.5 98610.0 8050.0 98675.0 ;
      RECT  8017.5 98582.5 8082.5 98642.5 ;
      RECT  8050.0 98550.0 8265.0 98615.0 ;
      RECT  8017.5 99925.0 8082.5 99990.0 ;
      RECT  8017.5 99985.0 8082.5 100050.0 ;
      RECT  7832.5 99925.0 8050.0 99990.0 ;
      RECT  8017.5 99957.5 8082.5 100017.5 ;
      RECT  8050.0 99985.0 8265.0 100050.0 ;
      RECT  8017.5 101300.0 8082.5 101365.0 ;
      RECT  8017.5 101240.0 8082.5 101305.0 ;
      RECT  7832.5 101300.0 8050.0 101365.0 ;
      RECT  8017.5 101272.5 8082.5 101332.5 ;
      RECT  8050.0 101240.0 8265.0 101305.0 ;
      RECT  8017.5 102615.0 8082.5 102680.0 ;
      RECT  8017.5 102675.0 8082.5 102740.0 ;
      RECT  7832.5 102615.0 8050.0 102680.0 ;
      RECT  8017.5 102647.5 8082.5 102707.5 ;
      RECT  8050.0 102675.0 8265.0 102740.0 ;
      RECT  8017.5 103990.0 8082.5 104055.0 ;
      RECT  8017.5 103930.0 8082.5 103995.0 ;
      RECT  7832.5 103990.0 8050.0 104055.0 ;
      RECT  8017.5 103962.5 8082.5 104022.5 ;
      RECT  8050.0 103930.0 8265.0 103995.0 ;
      RECT  8017.5 105305.0 8082.5 105370.0 ;
      RECT  8017.5 105365.0 8082.5 105430.0 ;
      RECT  7832.5 105305.0 8050.0 105370.0 ;
      RECT  8017.5 105337.5 8082.5 105397.5 ;
      RECT  8050.0 105365.0 8265.0 105430.0 ;
      RECT  8017.5 106680.0 8082.5 106745.0 ;
      RECT  8017.5 106620.0 8082.5 106685.0 ;
      RECT  7832.5 106680.0 8050.0 106745.0 ;
      RECT  8017.5 106652.5 8082.5 106712.5 ;
      RECT  8050.0 106620.0 8265.0 106685.0 ;
      RECT  8017.5 107995.0 8082.5 108060.0 ;
      RECT  8017.5 108055.0 8082.5 108120.0 ;
      RECT  7832.5 107995.0 8050.0 108060.0 ;
      RECT  8017.5 108027.5 8082.5 108087.5 ;
      RECT  8050.0 108055.0 8265.0 108120.0 ;
      RECT  8017.5 109370.0 8082.5 109435.0 ;
      RECT  8017.5 109310.0 8082.5 109375.0 ;
      RECT  7832.5 109370.0 8050.0 109435.0 ;
      RECT  8017.5 109342.5 8082.5 109402.5 ;
      RECT  8050.0 109310.0 8265.0 109375.0 ;
      RECT  8017.5 110685.0 8082.5 110750.0 ;
      RECT  8017.5 110745.0 8082.5 110810.0 ;
      RECT  7832.5 110685.0 8050.0 110750.0 ;
      RECT  8017.5 110717.5 8082.5 110777.5 ;
      RECT  8050.0 110745.0 8265.0 110810.0 ;
      RECT  8017.5 112060.0 8082.5 112125.0 ;
      RECT  8017.5 112000.0 8082.5 112065.0 ;
      RECT  7832.5 112060.0 8050.0 112125.0 ;
      RECT  8017.5 112032.5 8082.5 112092.5 ;
      RECT  8050.0 112000.0 8265.0 112065.0 ;
      RECT  8017.5 113375.0 8082.5 113440.0 ;
      RECT  8017.5 113435.0 8082.5 113500.0 ;
      RECT  7832.5 113375.0 8050.0 113440.0 ;
      RECT  8017.5 113407.5 8082.5 113467.5 ;
      RECT  8050.0 113435.0 8265.0 113500.0 ;
      RECT  5065.0 12470.0 7130.0 12535.0 ;
      RECT  5240.0 13905.0 7130.0 13970.0 ;
      RECT  5415.0 15160.0 7130.0 15225.0 ;
      RECT  5590.0 16595.0 7130.0 16660.0 ;
      RECT  5765.0 17850.0 7130.0 17915.0 ;
      RECT  5940.0 19285.0 7130.0 19350.0 ;
      RECT  6115.0 20540.0 7130.0 20605.0 ;
      RECT  6290.0 21975.0 7130.0 22040.0 ;
      RECT  6465.0 23230.0 7130.0 23295.0 ;
      RECT  6640.0 24665.0 7130.0 24730.0 ;
      RECT  6815.0 25920.0 7130.0 25985.0 ;
      RECT  6990.0 27355.0 7130.0 27420.0 ;
      RECT  5065.0 28670.0 7257.5 28735.0 ;
      RECT  5765.0 28530.0 7447.5 28595.0 ;
      RECT  6465.0 28390.0 7637.5 28455.0 ;
      RECT  5065.0 29985.0 7257.5 30050.0 ;
      RECT  5765.0 30125.0 7447.5 30190.0 ;
      RECT  6640.0 30265.0 7637.5 30330.0 ;
      RECT  5065.0 31360.0 7257.5 31425.0 ;
      RECT  5765.0 31220.0 7447.5 31285.0 ;
      RECT  6815.0 31080.0 7637.5 31145.0 ;
      RECT  5065.0 32675.0 7257.5 32740.0 ;
      RECT  5765.0 32815.0 7447.5 32880.0 ;
      RECT  6990.0 32955.0 7637.5 33020.0 ;
      RECT  5065.0 34050.0 7257.5 34115.0 ;
      RECT  5940.0 33910.0 7447.5 33975.0 ;
      RECT  6465.0 33770.0 7637.5 33835.0 ;
      RECT  5065.0 35365.0 7257.5 35430.0 ;
      RECT  5940.0 35505.0 7447.5 35570.0 ;
      RECT  6640.0 35645.0 7637.5 35710.0 ;
      RECT  5065.0 36740.0 7257.5 36805.0 ;
      RECT  5940.0 36600.0 7447.5 36665.0 ;
      RECT  6815.0 36460.0 7637.5 36525.0 ;
      RECT  5065.0 38055.0 7257.5 38120.0 ;
      RECT  5940.0 38195.0 7447.5 38260.0 ;
      RECT  6990.0 38335.0 7637.5 38400.0 ;
      RECT  5065.0 39430.0 7257.5 39495.0 ;
      RECT  6115.0 39290.0 7447.5 39355.0 ;
      RECT  6465.0 39150.0 7637.5 39215.0 ;
      RECT  5065.0 40745.0 7257.5 40810.0 ;
      RECT  6115.0 40885.0 7447.5 40950.0 ;
      RECT  6640.0 41025.0 7637.5 41090.0 ;
      RECT  5065.0 42120.0 7257.5 42185.0 ;
      RECT  6115.0 41980.0 7447.5 42045.0 ;
      RECT  6815.0 41840.0 7637.5 41905.0 ;
      RECT  5065.0 43435.0 7257.5 43500.0 ;
      RECT  6115.0 43575.0 7447.5 43640.0 ;
      RECT  6990.0 43715.0 7637.5 43780.0 ;
      RECT  5065.0 44810.0 7257.5 44875.0 ;
      RECT  6290.0 44670.0 7447.5 44735.0 ;
      RECT  6465.0 44530.0 7637.5 44595.0 ;
      RECT  5065.0 46125.0 7257.5 46190.0 ;
      RECT  6290.0 46265.0 7447.5 46330.0 ;
      RECT  6640.0 46405.0 7637.5 46470.0 ;
      RECT  5065.0 47500.0 7257.5 47565.0 ;
      RECT  6290.0 47360.0 7447.5 47425.0 ;
      RECT  6815.0 47220.0 7637.5 47285.0 ;
      RECT  5065.0 48815.0 7257.5 48880.0 ;
      RECT  6290.0 48955.0 7447.5 49020.0 ;
      RECT  6990.0 49095.0 7637.5 49160.0 ;
      RECT  5240.0 50190.0 7257.5 50255.0 ;
      RECT  5765.0 50050.0 7447.5 50115.0 ;
      RECT  6465.0 49910.0 7637.5 49975.0 ;
      RECT  5240.0 51505.0 7257.5 51570.0 ;
      RECT  5765.0 51645.0 7447.5 51710.0 ;
      RECT  6640.0 51785.0 7637.5 51850.0 ;
      RECT  5240.0 52880.0 7257.5 52945.0 ;
      RECT  5765.0 52740.0 7447.5 52805.0 ;
      RECT  6815.0 52600.0 7637.5 52665.0 ;
      RECT  5240.0 54195.0 7257.5 54260.0 ;
      RECT  5765.0 54335.0 7447.5 54400.0 ;
      RECT  6990.0 54475.0 7637.5 54540.0 ;
      RECT  5240.0 55570.0 7257.5 55635.0 ;
      RECT  5940.0 55430.0 7447.5 55495.0 ;
      RECT  6465.0 55290.0 7637.5 55355.0 ;
      RECT  5240.0 56885.0 7257.5 56950.0 ;
      RECT  5940.0 57025.0 7447.5 57090.0 ;
      RECT  6640.0 57165.0 7637.5 57230.0 ;
      RECT  5240.0 58260.0 7257.5 58325.0 ;
      RECT  5940.0 58120.0 7447.5 58185.0 ;
      RECT  6815.0 57980.0 7637.5 58045.0 ;
      RECT  5240.0 59575.0 7257.5 59640.0 ;
      RECT  5940.0 59715.0 7447.5 59780.0 ;
      RECT  6990.0 59855.0 7637.5 59920.0 ;
      RECT  5240.0 60950.0 7257.5 61015.0 ;
      RECT  6115.0 60810.0 7447.5 60875.0 ;
      RECT  6465.0 60670.0 7637.5 60735.0 ;
      RECT  5240.0 62265.0 7257.5 62330.0 ;
      RECT  6115.0 62405.0 7447.5 62470.0 ;
      RECT  6640.0 62545.0 7637.5 62610.0 ;
      RECT  5240.0 63640.0 7257.5 63705.0 ;
      RECT  6115.0 63500.0 7447.5 63565.0 ;
      RECT  6815.0 63360.0 7637.5 63425.0 ;
      RECT  5240.0 64955.0 7257.5 65020.0 ;
      RECT  6115.0 65095.0 7447.5 65160.0 ;
      RECT  6990.0 65235.0 7637.5 65300.0 ;
      RECT  5240.0 66330.0 7257.5 66395.0 ;
      RECT  6290.0 66190.0 7447.5 66255.0 ;
      RECT  6465.0 66050.0 7637.5 66115.0 ;
      RECT  5240.0 67645.0 7257.5 67710.0 ;
      RECT  6290.0 67785.0 7447.5 67850.0 ;
      RECT  6640.0 67925.0 7637.5 67990.0 ;
      RECT  5240.0 69020.0 7257.5 69085.0 ;
      RECT  6290.0 68880.0 7447.5 68945.0 ;
      RECT  6815.0 68740.0 7637.5 68805.0 ;
      RECT  5240.0 70335.0 7257.5 70400.0 ;
      RECT  6290.0 70475.0 7447.5 70540.0 ;
      RECT  6990.0 70615.0 7637.5 70680.0 ;
      RECT  5415.0 71710.0 7257.5 71775.0 ;
      RECT  5765.0 71570.0 7447.5 71635.0 ;
      RECT  6465.0 71430.0 7637.5 71495.0 ;
      RECT  5415.0 73025.0 7257.5 73090.0 ;
      RECT  5765.0 73165.0 7447.5 73230.0 ;
      RECT  6640.0 73305.0 7637.5 73370.0 ;
      RECT  5415.0 74400.0 7257.5 74465.0 ;
      RECT  5765.0 74260.0 7447.5 74325.0 ;
      RECT  6815.0 74120.0 7637.5 74185.0 ;
      RECT  5415.0 75715.0 7257.5 75780.0 ;
      RECT  5765.0 75855.0 7447.5 75920.0 ;
      RECT  6990.0 75995.0 7637.5 76060.0 ;
      RECT  5415.0 77090.0 7257.5 77155.0 ;
      RECT  5940.0 76950.0 7447.5 77015.0 ;
      RECT  6465.0 76810.0 7637.5 76875.0 ;
      RECT  5415.0 78405.0 7257.5 78470.0 ;
      RECT  5940.0 78545.0 7447.5 78610.0 ;
      RECT  6640.0 78685.0 7637.5 78750.0 ;
      RECT  5415.0 79780.0 7257.5 79845.0 ;
      RECT  5940.0 79640.0 7447.5 79705.0 ;
      RECT  6815.0 79500.0 7637.5 79565.0 ;
      RECT  5415.0 81095.0 7257.5 81160.0 ;
      RECT  5940.0 81235.0 7447.5 81300.0 ;
      RECT  6990.0 81375.0 7637.5 81440.0 ;
      RECT  5415.0 82470.0 7257.5 82535.0 ;
      RECT  6115.0 82330.0 7447.5 82395.0 ;
      RECT  6465.0 82190.0 7637.5 82255.0 ;
      RECT  5415.0 83785.0 7257.5 83850.0 ;
      RECT  6115.0 83925.0 7447.5 83990.0 ;
      RECT  6640.0 84065.0 7637.5 84130.0 ;
      RECT  5415.0 85160.0 7257.5 85225.0 ;
      RECT  6115.0 85020.0 7447.5 85085.0 ;
      RECT  6815.0 84880.0 7637.5 84945.0 ;
      RECT  5415.0 86475.0 7257.5 86540.0 ;
      RECT  6115.0 86615.0 7447.5 86680.0 ;
      RECT  6990.0 86755.0 7637.5 86820.0 ;
      RECT  5415.0 87850.0 7257.5 87915.0 ;
      RECT  6290.0 87710.0 7447.5 87775.0 ;
      RECT  6465.0 87570.0 7637.5 87635.0 ;
      RECT  5415.0 89165.0 7257.5 89230.0 ;
      RECT  6290.0 89305.0 7447.5 89370.0 ;
      RECT  6640.0 89445.0 7637.5 89510.0 ;
      RECT  5415.0 90540.0 7257.5 90605.0 ;
      RECT  6290.0 90400.0 7447.5 90465.0 ;
      RECT  6815.0 90260.0 7637.5 90325.0 ;
      RECT  5415.0 91855.0 7257.5 91920.0 ;
      RECT  6290.0 91995.0 7447.5 92060.0 ;
      RECT  6990.0 92135.0 7637.5 92200.0 ;
      RECT  5590.0 93230.0 7257.5 93295.0 ;
      RECT  5765.0 93090.0 7447.5 93155.0 ;
      RECT  6465.0 92950.0 7637.5 93015.0 ;
      RECT  5590.0 94545.0 7257.5 94610.0 ;
      RECT  5765.0 94685.0 7447.5 94750.0 ;
      RECT  6640.0 94825.0 7637.5 94890.0 ;
      RECT  5590.0 95920.0 7257.5 95985.0 ;
      RECT  5765.0 95780.0 7447.5 95845.0 ;
      RECT  6815.0 95640.0 7637.5 95705.0 ;
      RECT  5590.0 97235.0 7257.5 97300.0 ;
      RECT  5765.0 97375.0 7447.5 97440.0 ;
      RECT  6990.0 97515.0 7637.5 97580.0 ;
      RECT  5590.0 98610.0 7257.5 98675.0 ;
      RECT  5940.0 98470.0 7447.5 98535.0 ;
      RECT  6465.0 98330.0 7637.5 98395.0 ;
      RECT  5590.0 99925.0 7257.5 99990.0 ;
      RECT  5940.0 100065.0 7447.5 100130.0 ;
      RECT  6640.0 100205.0 7637.5 100270.0 ;
      RECT  5590.0 101300.0 7257.5 101365.0 ;
      RECT  5940.0 101160.0 7447.5 101225.0 ;
      RECT  6815.0 101020.0 7637.5 101085.0 ;
      RECT  5590.0 102615.0 7257.5 102680.0 ;
      RECT  5940.0 102755.0 7447.5 102820.0 ;
      RECT  6990.0 102895.0 7637.5 102960.0 ;
      RECT  5590.0 103990.0 7257.5 104055.0 ;
      RECT  6115.0 103850.0 7447.5 103915.0 ;
      RECT  6465.0 103710.0 7637.5 103775.0 ;
      RECT  5590.0 105305.0 7257.5 105370.0 ;
      RECT  6115.0 105445.0 7447.5 105510.0 ;
      RECT  6640.0 105585.0 7637.5 105650.0 ;
      RECT  5590.0 106680.0 7257.5 106745.0 ;
      RECT  6115.0 106540.0 7447.5 106605.0 ;
      RECT  6815.0 106400.0 7637.5 106465.0 ;
      RECT  5590.0 107995.0 7257.5 108060.0 ;
      RECT  6115.0 108135.0 7447.5 108200.0 ;
      RECT  6990.0 108275.0 7637.5 108340.0 ;
      RECT  5590.0 109370.0 7257.5 109435.0 ;
      RECT  6290.0 109230.0 7447.5 109295.0 ;
      RECT  6465.0 109090.0 7637.5 109155.0 ;
      RECT  5590.0 110685.0 7257.5 110750.0 ;
      RECT  6290.0 110825.0 7447.5 110890.0 ;
      RECT  6640.0 110965.0 7637.5 111030.0 ;
      RECT  5590.0 112060.0 7257.5 112125.0 ;
      RECT  6290.0 111920.0 7447.5 111985.0 ;
      RECT  6815.0 111780.0 7637.5 111845.0 ;
      RECT  5590.0 113375.0 7257.5 113440.0 ;
      RECT  6290.0 113515.0 7447.5 113580.0 ;
      RECT  6990.0 113655.0 7637.5 113720.0 ;
      RECT  9952.5 12470.0 9887.5 12535.0 ;
      RECT  9952.5 12992.5 9887.5 13057.5 ;
      RECT  10190.0 12470.0 9920.0 12535.0 ;
      RECT  9952.5 12502.5 9887.5 13025.0 ;
      RECT  9920.0 12992.5 9675.0 13057.5 ;
      RECT  11060.0 12470.0 10420.0 12535.0 ;
      RECT  9952.5 13905.0 9887.5 13970.0 ;
      RECT  9952.5 14337.5 9887.5 14402.5 ;
      RECT  10190.0 13905.0 9920.0 13970.0 ;
      RECT  9952.5 13937.5 9887.5 14370.0 ;
      RECT  9920.0 14337.5 9400.0 14402.5 ;
      RECT  10785.0 13905.0 10420.0 13970.0 ;
      RECT  11060.0 14667.5 9125.0 14732.5 ;
      RECT  10785.0 16012.5 8850.0 16077.5 ;
      RECT  9675.0 12482.5 8550.0 12547.5 ;
      RECT  9400.0 12267.5 8292.5 12332.5 ;
      RECT  9125.0 13892.5 8550.0 13957.5 ;
      RECT  9400.0 14107.5 8292.5 14172.5 ;
      RECT  9675.0 15172.5 8550.0 15237.5 ;
      RECT  8850.0 14957.5 8292.5 15022.5 ;
      RECT  9125.0 16582.5 8550.0 16647.5 ;
      RECT  8850.0 16797.5 8292.5 16862.5 ;
      RECT  7845.0 12482.5 7780.0 12547.5 ;
      RECT  7845.0 12470.0 7780.0 12535.0 ;
      RECT  8062.5 12482.5 7812.5 12547.5 ;
      RECT  7845.0 12502.5 7780.0 12515.0 ;
      RECT  7812.5 12470.0 7565.0 12535.0 ;
      RECT  7845.0 13892.5 7780.0 13957.5 ;
      RECT  7845.0 13905.0 7780.0 13970.0 ;
      RECT  8062.5 13892.5 7812.5 13957.5 ;
      RECT  7845.0 13925.0 7780.0 13937.5 ;
      RECT  7812.5 13905.0 7565.0 13970.0 ;
      RECT  7845.0 15172.5 7780.0 15237.5 ;
      RECT  7845.0 15160.0 7780.0 15225.0 ;
      RECT  8062.5 15172.5 7812.5 15237.5 ;
      RECT  7845.0 15192.5 7780.0 15205.0 ;
      RECT  7812.5 15160.0 7565.0 15225.0 ;
      RECT  7845.0 16582.5 7780.0 16647.5 ;
      RECT  7845.0 16595.0 7780.0 16660.0 ;
      RECT  8062.5 16582.5 7812.5 16647.5 ;
      RECT  7845.0 16615.0 7780.0 16627.5 ;
      RECT  7812.5 16595.0 7565.0 16660.0 ;
      RECT  10117.5 13035.0 10052.5 13220.0 ;
      RECT  10117.5 11875.0 10052.5 12060.0 ;
      RECT  10477.5 11992.5 10412.5 11842.5 ;
      RECT  10477.5 12877.5 10412.5 13252.5 ;
      RECT  10287.5 11992.5 10222.5 12877.5 ;
      RECT  10477.5 12877.5 10412.5 13012.5 ;
      RECT  10287.5 12877.5 10222.5 13012.5 ;
      RECT  10287.5 12877.5 10222.5 13012.5 ;
      RECT  10477.5 12877.5 10412.5 13012.5 ;
      RECT  10477.5 11992.5 10412.5 12127.5 ;
      RECT  10287.5 11992.5 10222.5 12127.5 ;
      RECT  10287.5 11992.5 10222.5 12127.5 ;
      RECT  10477.5 11992.5 10412.5 12127.5 ;
      RECT  10117.5 12967.5 10052.5 13102.5 ;
      RECT  10117.5 11992.5 10052.5 12127.5 ;
      RECT  10420.0 12435.0 10355.0 12570.0 ;
      RECT  10420.0 12435.0 10355.0 12570.0 ;
      RECT  10255.0 12470.0 10190.0 12535.0 ;
      RECT  10545.0 13187.5 9985.0 13252.5 ;
      RECT  10545.0 11842.5 9985.0 11907.5 ;
      RECT  10117.5 13405.0 10052.5 13220.0 ;
      RECT  10117.5 14565.0 10052.5 14380.0 ;
      RECT  10477.5 14447.5 10412.5 14597.5 ;
      RECT  10477.5 13562.5 10412.5 13187.5 ;
      RECT  10287.5 14447.5 10222.5 13562.5 ;
      RECT  10477.5 13562.5 10412.5 13427.5 ;
      RECT  10287.5 13562.5 10222.5 13427.5 ;
      RECT  10287.5 13562.5 10222.5 13427.5 ;
      RECT  10477.5 13562.5 10412.5 13427.5 ;
      RECT  10477.5 14447.5 10412.5 14312.5 ;
      RECT  10287.5 14447.5 10222.5 14312.5 ;
      RECT  10287.5 14447.5 10222.5 14312.5 ;
      RECT  10477.5 14447.5 10412.5 14312.5 ;
      RECT  10117.5 13472.5 10052.5 13337.5 ;
      RECT  10117.5 14447.5 10052.5 14312.5 ;
      RECT  10420.0 14005.0 10355.0 13870.0 ;
      RECT  10420.0 14005.0 10355.0 13870.0 ;
      RECT  10255.0 13970.0 10190.0 13905.0 ;
      RECT  10545.0 13252.5 9985.0 13187.5 ;
      RECT  10545.0 14597.5 9985.0 14532.5 ;
      RECT  7262.5 13035.0 7197.5 13220.0 ;
      RECT  7262.5 11875.0 7197.5 12060.0 ;
      RECT  7622.5 11992.5 7557.5 11842.5 ;
      RECT  7622.5 12877.5 7557.5 13252.5 ;
      RECT  7432.5 11992.5 7367.5 12877.5 ;
      RECT  7622.5 12877.5 7557.5 13012.5 ;
      RECT  7432.5 12877.5 7367.5 13012.5 ;
      RECT  7432.5 12877.5 7367.5 13012.5 ;
      RECT  7622.5 12877.5 7557.5 13012.5 ;
      RECT  7622.5 11992.5 7557.5 12127.5 ;
      RECT  7432.5 11992.5 7367.5 12127.5 ;
      RECT  7432.5 11992.5 7367.5 12127.5 ;
      RECT  7622.5 11992.5 7557.5 12127.5 ;
      RECT  7262.5 12967.5 7197.5 13102.5 ;
      RECT  7262.5 11992.5 7197.5 12127.5 ;
      RECT  7565.0 12435.0 7500.0 12570.0 ;
      RECT  7565.0 12435.0 7500.0 12570.0 ;
      RECT  7400.0 12470.0 7335.0 12535.0 ;
      RECT  7690.0 13187.5 7130.0 13252.5 ;
      RECT  7690.0 11842.5 7130.0 11907.5 ;
      RECT  7262.5 13405.0 7197.5 13220.0 ;
      RECT  7262.5 14565.0 7197.5 14380.0 ;
      RECT  7622.5 14447.5 7557.5 14597.5 ;
      RECT  7622.5 13562.5 7557.5 13187.5 ;
      RECT  7432.5 14447.5 7367.5 13562.5 ;
      RECT  7622.5 13562.5 7557.5 13427.5 ;
      RECT  7432.5 13562.5 7367.5 13427.5 ;
      RECT  7432.5 13562.5 7367.5 13427.5 ;
      RECT  7622.5 13562.5 7557.5 13427.5 ;
      RECT  7622.5 14447.5 7557.5 14312.5 ;
      RECT  7432.5 14447.5 7367.5 14312.5 ;
      RECT  7432.5 14447.5 7367.5 14312.5 ;
      RECT  7622.5 14447.5 7557.5 14312.5 ;
      RECT  7262.5 13472.5 7197.5 13337.5 ;
      RECT  7262.5 14447.5 7197.5 14312.5 ;
      RECT  7565.0 14005.0 7500.0 13870.0 ;
      RECT  7565.0 14005.0 7500.0 13870.0 ;
      RECT  7400.0 13970.0 7335.0 13905.0 ;
      RECT  7690.0 13252.5 7130.0 13187.5 ;
      RECT  7690.0 14597.5 7130.0 14532.5 ;
      RECT  7262.5 15725.0 7197.5 15910.0 ;
      RECT  7262.5 14565.0 7197.5 14750.0 ;
      RECT  7622.5 14682.5 7557.5 14532.5 ;
      RECT  7622.5 15567.5 7557.5 15942.5 ;
      RECT  7432.5 14682.5 7367.5 15567.5 ;
      RECT  7622.5 15567.5 7557.5 15702.5 ;
      RECT  7432.5 15567.5 7367.5 15702.5 ;
      RECT  7432.5 15567.5 7367.5 15702.5 ;
      RECT  7622.5 15567.5 7557.5 15702.5 ;
      RECT  7622.5 14682.5 7557.5 14817.5 ;
      RECT  7432.5 14682.5 7367.5 14817.5 ;
      RECT  7432.5 14682.5 7367.5 14817.5 ;
      RECT  7622.5 14682.5 7557.5 14817.5 ;
      RECT  7262.5 15657.5 7197.5 15792.5 ;
      RECT  7262.5 14682.5 7197.5 14817.5 ;
      RECT  7565.0 15125.0 7500.0 15260.0 ;
      RECT  7565.0 15125.0 7500.0 15260.0 ;
      RECT  7400.0 15160.0 7335.0 15225.0 ;
      RECT  7690.0 15877.5 7130.0 15942.5 ;
      RECT  7690.0 14532.5 7130.0 14597.5 ;
      RECT  7262.5 16095.0 7197.5 15910.0 ;
      RECT  7262.5 17255.0 7197.5 17070.0 ;
      RECT  7622.5 17137.5 7557.5 17287.5 ;
      RECT  7622.5 16252.5 7557.5 15877.5 ;
      RECT  7432.5 17137.5 7367.5 16252.5 ;
      RECT  7622.5 16252.5 7557.5 16117.5 ;
      RECT  7432.5 16252.5 7367.5 16117.5 ;
      RECT  7432.5 16252.5 7367.5 16117.5 ;
      RECT  7622.5 16252.5 7557.5 16117.5 ;
      RECT  7622.5 17137.5 7557.5 17002.5 ;
      RECT  7432.5 17137.5 7367.5 17002.5 ;
      RECT  7432.5 17137.5 7367.5 17002.5 ;
      RECT  7622.5 17137.5 7557.5 17002.5 ;
      RECT  7262.5 16162.5 7197.5 16027.5 ;
      RECT  7262.5 17137.5 7197.5 17002.5 ;
      RECT  7565.0 16695.0 7500.0 16560.0 ;
      RECT  7565.0 16695.0 7500.0 16560.0 ;
      RECT  7400.0 16660.0 7335.0 16595.0 ;
      RECT  7690.0 15942.5 7130.0 15877.5 ;
      RECT  7690.0 17287.5 7130.0 17222.5 ;
      RECT  8542.5 12037.5 8477.5 11842.5 ;
      RECT  8542.5 12877.5 8477.5 13252.5 ;
      RECT  8162.5 12877.5 8097.5 13252.5 ;
      RECT  7992.5 13035.0 7927.5 13220.0 ;
      RECT  7992.5 11875.0 7927.5 12060.0 ;
      RECT  8542.5 12877.5 8477.5 13012.5 ;
      RECT  8352.5 12877.5 8287.5 13012.5 ;
      RECT  8352.5 12877.5 8287.5 13012.5 ;
      RECT  8542.5 12877.5 8477.5 13012.5 ;
      RECT  8352.5 12877.5 8287.5 13012.5 ;
      RECT  8162.5 12877.5 8097.5 13012.5 ;
      RECT  8162.5 12877.5 8097.5 13012.5 ;
      RECT  8352.5 12877.5 8287.5 13012.5 ;
      RECT  8542.5 12037.5 8477.5 12172.5 ;
      RECT  8352.5 12037.5 8287.5 12172.5 ;
      RECT  8352.5 12037.5 8287.5 12172.5 ;
      RECT  8542.5 12037.5 8477.5 12172.5 ;
      RECT  8352.5 12037.5 8287.5 12172.5 ;
      RECT  8162.5 12037.5 8097.5 12172.5 ;
      RECT  8162.5 12037.5 8097.5 12172.5 ;
      RECT  8352.5 12037.5 8287.5 12172.5 ;
      RECT  7992.5 12967.5 7927.5 13102.5 ;
      RECT  7992.5 11992.5 7927.5 12127.5 ;
      RECT  8157.5 12267.5 8292.5 12332.5 ;
      RECT  8415.0 12482.5 8550.0 12547.5 ;
      RECT  8352.5 12877.5 8287.5 13012.5 ;
      RECT  8162.5 12037.5 8097.5 12172.5 ;
      RECT  8062.5 12482.5 8197.5 12547.5 ;
      RECT  8550.0 12482.5 8415.0 12547.5 ;
      RECT  8292.5 12267.5 8157.5 12332.5 ;
      RECT  8197.5 12482.5 8062.5 12547.5 ;
      RECT  8610.0 13187.5 7690.0 13252.5 ;
      RECT  8610.0 11842.5 7690.0 11907.5 ;
      RECT  8542.5 14402.5 8477.5 14597.5 ;
      RECT  8542.5 13562.5 8477.5 13187.5 ;
      RECT  8162.5 13562.5 8097.5 13187.5 ;
      RECT  7992.5 13405.0 7927.5 13220.0 ;
      RECT  7992.5 14565.0 7927.5 14380.0 ;
      RECT  8542.5 13562.5 8477.5 13427.5 ;
      RECT  8352.5 13562.5 8287.5 13427.5 ;
      RECT  8352.5 13562.5 8287.5 13427.5 ;
      RECT  8542.5 13562.5 8477.5 13427.5 ;
      RECT  8352.5 13562.5 8287.5 13427.5 ;
      RECT  8162.5 13562.5 8097.5 13427.5 ;
      RECT  8162.5 13562.5 8097.5 13427.5 ;
      RECT  8352.5 13562.5 8287.5 13427.5 ;
      RECT  8542.5 14402.5 8477.5 14267.5 ;
      RECT  8352.5 14402.5 8287.5 14267.5 ;
      RECT  8352.5 14402.5 8287.5 14267.5 ;
      RECT  8542.5 14402.5 8477.5 14267.5 ;
      RECT  8352.5 14402.5 8287.5 14267.5 ;
      RECT  8162.5 14402.5 8097.5 14267.5 ;
      RECT  8162.5 14402.5 8097.5 14267.5 ;
      RECT  8352.5 14402.5 8287.5 14267.5 ;
      RECT  7992.5 13472.5 7927.5 13337.5 ;
      RECT  7992.5 14447.5 7927.5 14312.5 ;
      RECT  8157.5 14172.5 8292.5 14107.5 ;
      RECT  8415.0 13957.5 8550.0 13892.5 ;
      RECT  8352.5 13562.5 8287.5 13427.5 ;
      RECT  8162.5 14402.5 8097.5 14267.5 ;
      RECT  8062.5 13957.5 8197.5 13892.5 ;
      RECT  8550.0 13957.5 8415.0 13892.5 ;
      RECT  8292.5 14172.5 8157.5 14107.5 ;
      RECT  8197.5 13957.5 8062.5 13892.5 ;
      RECT  8610.0 13252.5 7690.0 13187.5 ;
      RECT  8610.0 14597.5 7690.0 14532.5 ;
      RECT  8542.5 14727.5 8477.5 14532.5 ;
      RECT  8542.5 15567.5 8477.5 15942.5 ;
      RECT  8162.5 15567.5 8097.5 15942.5 ;
      RECT  7992.5 15725.0 7927.5 15910.0 ;
      RECT  7992.5 14565.0 7927.5 14750.0 ;
      RECT  8542.5 15567.5 8477.5 15702.5 ;
      RECT  8352.5 15567.5 8287.5 15702.5 ;
      RECT  8352.5 15567.5 8287.5 15702.5 ;
      RECT  8542.5 15567.5 8477.5 15702.5 ;
      RECT  8352.5 15567.5 8287.5 15702.5 ;
      RECT  8162.5 15567.5 8097.5 15702.5 ;
      RECT  8162.5 15567.5 8097.5 15702.5 ;
      RECT  8352.5 15567.5 8287.5 15702.5 ;
      RECT  8542.5 14727.5 8477.5 14862.5 ;
      RECT  8352.5 14727.5 8287.5 14862.5 ;
      RECT  8352.5 14727.5 8287.5 14862.5 ;
      RECT  8542.5 14727.5 8477.5 14862.5 ;
      RECT  8352.5 14727.5 8287.5 14862.5 ;
      RECT  8162.5 14727.5 8097.5 14862.5 ;
      RECT  8162.5 14727.5 8097.5 14862.5 ;
      RECT  8352.5 14727.5 8287.5 14862.5 ;
      RECT  7992.5 15657.5 7927.5 15792.5 ;
      RECT  7992.5 14682.5 7927.5 14817.5 ;
      RECT  8157.5 14957.5 8292.5 15022.5 ;
      RECT  8415.0 15172.5 8550.0 15237.5 ;
      RECT  8352.5 15567.5 8287.5 15702.5 ;
      RECT  8162.5 14727.5 8097.5 14862.5 ;
      RECT  8062.5 15172.5 8197.5 15237.5 ;
      RECT  8550.0 15172.5 8415.0 15237.5 ;
      RECT  8292.5 14957.5 8157.5 15022.5 ;
      RECT  8197.5 15172.5 8062.5 15237.5 ;
      RECT  8610.0 15877.5 7690.0 15942.5 ;
      RECT  8610.0 14532.5 7690.0 14597.5 ;
      RECT  8542.5 17092.5 8477.5 17287.5 ;
      RECT  8542.5 16252.5 8477.5 15877.5 ;
      RECT  8162.5 16252.5 8097.5 15877.5 ;
      RECT  7992.5 16095.0 7927.5 15910.0 ;
      RECT  7992.5 17255.0 7927.5 17070.0 ;
      RECT  8542.5 16252.5 8477.5 16117.5 ;
      RECT  8352.5 16252.5 8287.5 16117.5 ;
      RECT  8352.5 16252.5 8287.5 16117.5 ;
      RECT  8542.5 16252.5 8477.5 16117.5 ;
      RECT  8352.5 16252.5 8287.5 16117.5 ;
      RECT  8162.5 16252.5 8097.5 16117.5 ;
      RECT  8162.5 16252.5 8097.5 16117.5 ;
      RECT  8352.5 16252.5 8287.5 16117.5 ;
      RECT  8542.5 17092.5 8477.5 16957.5 ;
      RECT  8352.5 17092.5 8287.5 16957.5 ;
      RECT  8352.5 17092.5 8287.5 16957.5 ;
      RECT  8542.5 17092.5 8477.5 16957.5 ;
      RECT  8352.5 17092.5 8287.5 16957.5 ;
      RECT  8162.5 17092.5 8097.5 16957.5 ;
      RECT  8162.5 17092.5 8097.5 16957.5 ;
      RECT  8352.5 17092.5 8287.5 16957.5 ;
      RECT  7992.5 16162.5 7927.5 16027.5 ;
      RECT  7992.5 17137.5 7927.5 17002.5 ;
      RECT  8157.5 16862.5 8292.5 16797.5 ;
      RECT  8415.0 16647.5 8550.0 16582.5 ;
      RECT  8352.5 16252.5 8287.5 16117.5 ;
      RECT  8162.5 17092.5 8097.5 16957.5 ;
      RECT  8062.5 16647.5 8197.5 16582.5 ;
      RECT  8550.0 16647.5 8415.0 16582.5 ;
      RECT  8292.5 16862.5 8157.5 16797.5 ;
      RECT  8197.5 16647.5 8062.5 16582.5 ;
      RECT  8610.0 15942.5 7690.0 15877.5 ;
      RECT  8610.0 17287.5 7690.0 17222.5 ;
      RECT  9607.5 12992.5 9742.5 13057.5 ;
      RECT  10992.5 12470.0 11127.5 12535.0 ;
      RECT  9332.5 14337.5 9467.5 14402.5 ;
      RECT  10717.5 13905.0 10852.5 13970.0 ;
      RECT  10992.5 14667.5 11127.5 14732.5 ;
      RECT  9057.5 14667.5 9192.5 14732.5 ;
      RECT  10717.5 16012.5 10852.5 16077.5 ;
      RECT  8782.5 16012.5 8917.5 16077.5 ;
      RECT  9607.5 12482.5 9742.5 12547.5 ;
      RECT  9332.5 12267.5 9467.5 12332.5 ;
      RECT  9057.5 13892.5 9192.5 13957.5 ;
      RECT  9332.5 14107.5 9467.5 14172.5 ;
      RECT  9607.5 15172.5 9742.5 15237.5 ;
      RECT  8782.5 14957.5 8917.5 15022.5 ;
      RECT  9057.5 16582.5 9192.5 16647.5 ;
      RECT  8782.5 16797.5 8917.5 16862.5 ;
      RECT  7335.0 12470.0 7130.0 12535.0 ;
      RECT  7335.0 13905.0 7130.0 13970.0 ;
      RECT  7335.0 15160.0 7130.0 15225.0 ;
      RECT  7335.0 16595.0 7130.0 16660.0 ;
      RECT  11095.0 13187.5 7130.0 13252.5 ;
      RECT  11095.0 15877.5 7130.0 15942.5 ;
      RECT  11095.0 11842.5 7130.0 11907.5 ;
      RECT  11095.0 14532.5 7130.0 14597.5 ;
      RECT  11095.0 17222.5 7130.0 17287.5 ;
      RECT  9952.5 17850.0 9887.5 17915.0 ;
      RECT  9952.5 18372.5 9887.5 18437.5 ;
      RECT  10190.0 17850.0 9920.0 17915.0 ;
      RECT  9952.5 17882.5 9887.5 18405.0 ;
      RECT  9920.0 18372.5 9675.0 18437.5 ;
      RECT  11060.0 17850.0 10420.0 17915.0 ;
      RECT  9952.5 19285.0 9887.5 19350.0 ;
      RECT  9952.5 19717.5 9887.5 19782.5 ;
      RECT  10190.0 19285.0 9920.0 19350.0 ;
      RECT  9952.5 19317.5 9887.5 19750.0 ;
      RECT  9920.0 19717.5 9400.0 19782.5 ;
      RECT  10785.0 19285.0 10420.0 19350.0 ;
      RECT  11060.0 20047.5 9125.0 20112.5 ;
      RECT  10785.0 21392.5 8850.0 21457.5 ;
      RECT  9675.0 17862.5 8550.0 17927.5 ;
      RECT  9400.0 17647.5 8292.5 17712.5 ;
      RECT  9125.0 19272.5 8550.0 19337.5 ;
      RECT  9400.0 19487.5 8292.5 19552.5 ;
      RECT  9675.0 20552.5 8550.0 20617.5 ;
      RECT  8850.0 20337.5 8292.5 20402.5 ;
      RECT  9125.0 21962.5 8550.0 22027.5 ;
      RECT  8850.0 22177.5 8292.5 22242.5 ;
      RECT  7845.0 17862.5 7780.0 17927.5 ;
      RECT  7845.0 17850.0 7780.0 17915.0 ;
      RECT  8062.5 17862.5 7812.5 17927.5 ;
      RECT  7845.0 17882.5 7780.0 17895.0 ;
      RECT  7812.5 17850.0 7565.0 17915.0 ;
      RECT  7845.0 19272.5 7780.0 19337.5 ;
      RECT  7845.0 19285.0 7780.0 19350.0 ;
      RECT  8062.5 19272.5 7812.5 19337.5 ;
      RECT  7845.0 19305.0 7780.0 19317.5 ;
      RECT  7812.5 19285.0 7565.0 19350.0 ;
      RECT  7845.0 20552.5 7780.0 20617.5 ;
      RECT  7845.0 20540.0 7780.0 20605.0 ;
      RECT  8062.5 20552.5 7812.5 20617.5 ;
      RECT  7845.0 20572.5 7780.0 20585.0 ;
      RECT  7812.5 20540.0 7565.0 20605.0 ;
      RECT  7845.0 21962.5 7780.0 22027.5 ;
      RECT  7845.0 21975.0 7780.0 22040.0 ;
      RECT  8062.5 21962.5 7812.5 22027.5 ;
      RECT  7845.0 21995.0 7780.0 22007.5 ;
      RECT  7812.5 21975.0 7565.0 22040.0 ;
      RECT  10117.5 18415.0 10052.5 18600.0 ;
      RECT  10117.5 17255.0 10052.5 17440.0 ;
      RECT  10477.5 17372.5 10412.5 17222.5 ;
      RECT  10477.5 18257.5 10412.5 18632.5 ;
      RECT  10287.5 17372.5 10222.5 18257.5 ;
      RECT  10477.5 18257.5 10412.5 18392.5 ;
      RECT  10287.5 18257.5 10222.5 18392.5 ;
      RECT  10287.5 18257.5 10222.5 18392.5 ;
      RECT  10477.5 18257.5 10412.5 18392.5 ;
      RECT  10477.5 17372.5 10412.5 17507.5 ;
      RECT  10287.5 17372.5 10222.5 17507.5 ;
      RECT  10287.5 17372.5 10222.5 17507.5 ;
      RECT  10477.5 17372.5 10412.5 17507.5 ;
      RECT  10117.5 18347.5 10052.5 18482.5 ;
      RECT  10117.5 17372.5 10052.5 17507.5 ;
      RECT  10420.0 17815.0 10355.0 17950.0 ;
      RECT  10420.0 17815.0 10355.0 17950.0 ;
      RECT  10255.0 17850.0 10190.0 17915.0 ;
      RECT  10545.0 18567.5 9985.0 18632.5 ;
      RECT  10545.0 17222.5 9985.0 17287.5 ;
      RECT  10117.5 18785.0 10052.5 18600.0 ;
      RECT  10117.5 19945.0 10052.5 19760.0 ;
      RECT  10477.5 19827.5 10412.5 19977.5 ;
      RECT  10477.5 18942.5 10412.5 18567.5 ;
      RECT  10287.5 19827.5 10222.5 18942.5 ;
      RECT  10477.5 18942.5 10412.5 18807.5 ;
      RECT  10287.5 18942.5 10222.5 18807.5 ;
      RECT  10287.5 18942.5 10222.5 18807.5 ;
      RECT  10477.5 18942.5 10412.5 18807.5 ;
      RECT  10477.5 19827.5 10412.5 19692.5 ;
      RECT  10287.5 19827.5 10222.5 19692.5 ;
      RECT  10287.5 19827.5 10222.5 19692.5 ;
      RECT  10477.5 19827.5 10412.5 19692.5 ;
      RECT  10117.5 18852.5 10052.5 18717.5 ;
      RECT  10117.5 19827.5 10052.5 19692.5 ;
      RECT  10420.0 19385.0 10355.0 19250.0 ;
      RECT  10420.0 19385.0 10355.0 19250.0 ;
      RECT  10255.0 19350.0 10190.0 19285.0 ;
      RECT  10545.0 18632.5 9985.0 18567.5 ;
      RECT  10545.0 19977.5 9985.0 19912.5 ;
      RECT  7262.5 18415.0 7197.5 18600.0 ;
      RECT  7262.5 17255.0 7197.5 17440.0 ;
      RECT  7622.5 17372.5 7557.5 17222.5 ;
      RECT  7622.5 18257.5 7557.5 18632.5 ;
      RECT  7432.5 17372.5 7367.5 18257.5 ;
      RECT  7622.5 18257.5 7557.5 18392.5 ;
      RECT  7432.5 18257.5 7367.5 18392.5 ;
      RECT  7432.5 18257.5 7367.5 18392.5 ;
      RECT  7622.5 18257.5 7557.5 18392.5 ;
      RECT  7622.5 17372.5 7557.5 17507.5 ;
      RECT  7432.5 17372.5 7367.5 17507.5 ;
      RECT  7432.5 17372.5 7367.5 17507.5 ;
      RECT  7622.5 17372.5 7557.5 17507.5 ;
      RECT  7262.5 18347.5 7197.5 18482.5 ;
      RECT  7262.5 17372.5 7197.5 17507.5 ;
      RECT  7565.0 17815.0 7500.0 17950.0 ;
      RECT  7565.0 17815.0 7500.0 17950.0 ;
      RECT  7400.0 17850.0 7335.0 17915.0 ;
      RECT  7690.0 18567.5 7130.0 18632.5 ;
      RECT  7690.0 17222.5 7130.0 17287.5 ;
      RECT  7262.5 18785.0 7197.5 18600.0 ;
      RECT  7262.5 19945.0 7197.5 19760.0 ;
      RECT  7622.5 19827.5 7557.5 19977.5 ;
      RECT  7622.5 18942.5 7557.5 18567.5 ;
      RECT  7432.5 19827.5 7367.5 18942.5 ;
      RECT  7622.5 18942.5 7557.5 18807.5 ;
      RECT  7432.5 18942.5 7367.5 18807.5 ;
      RECT  7432.5 18942.5 7367.5 18807.5 ;
      RECT  7622.5 18942.5 7557.5 18807.5 ;
      RECT  7622.5 19827.5 7557.5 19692.5 ;
      RECT  7432.5 19827.5 7367.5 19692.5 ;
      RECT  7432.5 19827.5 7367.5 19692.5 ;
      RECT  7622.5 19827.5 7557.5 19692.5 ;
      RECT  7262.5 18852.5 7197.5 18717.5 ;
      RECT  7262.5 19827.5 7197.5 19692.5 ;
      RECT  7565.0 19385.0 7500.0 19250.0 ;
      RECT  7565.0 19385.0 7500.0 19250.0 ;
      RECT  7400.0 19350.0 7335.0 19285.0 ;
      RECT  7690.0 18632.5 7130.0 18567.5 ;
      RECT  7690.0 19977.5 7130.0 19912.5 ;
      RECT  7262.5 21105.0 7197.5 21290.0 ;
      RECT  7262.5 19945.0 7197.5 20130.0 ;
      RECT  7622.5 20062.5 7557.5 19912.5 ;
      RECT  7622.5 20947.5 7557.5 21322.5 ;
      RECT  7432.5 20062.5 7367.5 20947.5 ;
      RECT  7622.5 20947.5 7557.5 21082.5 ;
      RECT  7432.5 20947.5 7367.5 21082.5 ;
      RECT  7432.5 20947.5 7367.5 21082.5 ;
      RECT  7622.5 20947.5 7557.5 21082.5 ;
      RECT  7622.5 20062.5 7557.5 20197.5 ;
      RECT  7432.5 20062.5 7367.5 20197.5 ;
      RECT  7432.5 20062.5 7367.5 20197.5 ;
      RECT  7622.5 20062.5 7557.5 20197.5 ;
      RECT  7262.5 21037.5 7197.5 21172.5 ;
      RECT  7262.5 20062.5 7197.5 20197.5 ;
      RECT  7565.0 20505.0 7500.0 20640.0 ;
      RECT  7565.0 20505.0 7500.0 20640.0 ;
      RECT  7400.0 20540.0 7335.0 20605.0 ;
      RECT  7690.0 21257.5 7130.0 21322.5 ;
      RECT  7690.0 19912.5 7130.0 19977.5 ;
      RECT  7262.5 21475.0 7197.5 21290.0 ;
      RECT  7262.5 22635.0 7197.5 22450.0 ;
      RECT  7622.5 22517.5 7557.5 22667.5 ;
      RECT  7622.5 21632.5 7557.5 21257.5 ;
      RECT  7432.5 22517.5 7367.5 21632.5 ;
      RECT  7622.5 21632.5 7557.5 21497.5 ;
      RECT  7432.5 21632.5 7367.5 21497.5 ;
      RECT  7432.5 21632.5 7367.5 21497.5 ;
      RECT  7622.5 21632.5 7557.5 21497.5 ;
      RECT  7622.5 22517.5 7557.5 22382.5 ;
      RECT  7432.5 22517.5 7367.5 22382.5 ;
      RECT  7432.5 22517.5 7367.5 22382.5 ;
      RECT  7622.5 22517.5 7557.5 22382.5 ;
      RECT  7262.5 21542.5 7197.5 21407.5 ;
      RECT  7262.5 22517.5 7197.5 22382.5 ;
      RECT  7565.0 22075.0 7500.0 21940.0 ;
      RECT  7565.0 22075.0 7500.0 21940.0 ;
      RECT  7400.0 22040.0 7335.0 21975.0 ;
      RECT  7690.0 21322.5 7130.0 21257.5 ;
      RECT  7690.0 22667.5 7130.0 22602.5 ;
      RECT  8542.5 17417.5 8477.5 17222.5 ;
      RECT  8542.5 18257.5 8477.5 18632.5 ;
      RECT  8162.5 18257.5 8097.5 18632.5 ;
      RECT  7992.5 18415.0 7927.5 18600.0 ;
      RECT  7992.5 17255.0 7927.5 17440.0 ;
      RECT  8542.5 18257.5 8477.5 18392.5 ;
      RECT  8352.5 18257.5 8287.5 18392.5 ;
      RECT  8352.5 18257.5 8287.5 18392.5 ;
      RECT  8542.5 18257.5 8477.5 18392.5 ;
      RECT  8352.5 18257.5 8287.5 18392.5 ;
      RECT  8162.5 18257.5 8097.5 18392.5 ;
      RECT  8162.5 18257.5 8097.5 18392.5 ;
      RECT  8352.5 18257.5 8287.5 18392.5 ;
      RECT  8542.5 17417.5 8477.5 17552.5 ;
      RECT  8352.5 17417.5 8287.5 17552.5 ;
      RECT  8352.5 17417.5 8287.5 17552.5 ;
      RECT  8542.5 17417.5 8477.5 17552.5 ;
      RECT  8352.5 17417.5 8287.5 17552.5 ;
      RECT  8162.5 17417.5 8097.5 17552.5 ;
      RECT  8162.5 17417.5 8097.5 17552.5 ;
      RECT  8352.5 17417.5 8287.5 17552.5 ;
      RECT  7992.5 18347.5 7927.5 18482.5 ;
      RECT  7992.5 17372.5 7927.5 17507.5 ;
      RECT  8157.5 17647.5 8292.5 17712.5 ;
      RECT  8415.0 17862.5 8550.0 17927.5 ;
      RECT  8352.5 18257.5 8287.5 18392.5 ;
      RECT  8162.5 17417.5 8097.5 17552.5 ;
      RECT  8062.5 17862.5 8197.5 17927.5 ;
      RECT  8550.0 17862.5 8415.0 17927.5 ;
      RECT  8292.5 17647.5 8157.5 17712.5 ;
      RECT  8197.5 17862.5 8062.5 17927.5 ;
      RECT  8610.0 18567.5 7690.0 18632.5 ;
      RECT  8610.0 17222.5 7690.0 17287.5 ;
      RECT  8542.5 19782.5 8477.5 19977.5 ;
      RECT  8542.5 18942.5 8477.5 18567.5 ;
      RECT  8162.5 18942.5 8097.5 18567.5 ;
      RECT  7992.5 18785.0 7927.5 18600.0 ;
      RECT  7992.5 19945.0 7927.5 19760.0 ;
      RECT  8542.5 18942.5 8477.5 18807.5 ;
      RECT  8352.5 18942.5 8287.5 18807.5 ;
      RECT  8352.5 18942.5 8287.5 18807.5 ;
      RECT  8542.5 18942.5 8477.5 18807.5 ;
      RECT  8352.5 18942.5 8287.5 18807.5 ;
      RECT  8162.5 18942.5 8097.5 18807.5 ;
      RECT  8162.5 18942.5 8097.5 18807.5 ;
      RECT  8352.5 18942.5 8287.5 18807.5 ;
      RECT  8542.5 19782.5 8477.5 19647.5 ;
      RECT  8352.5 19782.5 8287.5 19647.5 ;
      RECT  8352.5 19782.5 8287.5 19647.5 ;
      RECT  8542.5 19782.5 8477.5 19647.5 ;
      RECT  8352.5 19782.5 8287.5 19647.5 ;
      RECT  8162.5 19782.5 8097.5 19647.5 ;
      RECT  8162.5 19782.5 8097.5 19647.5 ;
      RECT  8352.5 19782.5 8287.5 19647.5 ;
      RECT  7992.5 18852.5 7927.5 18717.5 ;
      RECT  7992.5 19827.5 7927.5 19692.5 ;
      RECT  8157.5 19552.5 8292.5 19487.5 ;
      RECT  8415.0 19337.5 8550.0 19272.5 ;
      RECT  8352.5 18942.5 8287.5 18807.5 ;
      RECT  8162.5 19782.5 8097.5 19647.5 ;
      RECT  8062.5 19337.5 8197.5 19272.5 ;
      RECT  8550.0 19337.5 8415.0 19272.5 ;
      RECT  8292.5 19552.5 8157.5 19487.5 ;
      RECT  8197.5 19337.5 8062.5 19272.5 ;
      RECT  8610.0 18632.5 7690.0 18567.5 ;
      RECT  8610.0 19977.5 7690.0 19912.5 ;
      RECT  8542.5 20107.5 8477.5 19912.5 ;
      RECT  8542.5 20947.5 8477.5 21322.5 ;
      RECT  8162.5 20947.5 8097.5 21322.5 ;
      RECT  7992.5 21105.0 7927.5 21290.0 ;
      RECT  7992.5 19945.0 7927.5 20130.0 ;
      RECT  8542.5 20947.5 8477.5 21082.5 ;
      RECT  8352.5 20947.5 8287.5 21082.5 ;
      RECT  8352.5 20947.5 8287.5 21082.5 ;
      RECT  8542.5 20947.5 8477.5 21082.5 ;
      RECT  8352.5 20947.5 8287.5 21082.5 ;
      RECT  8162.5 20947.5 8097.5 21082.5 ;
      RECT  8162.5 20947.5 8097.5 21082.5 ;
      RECT  8352.5 20947.5 8287.5 21082.5 ;
      RECT  8542.5 20107.5 8477.5 20242.5 ;
      RECT  8352.5 20107.5 8287.5 20242.5 ;
      RECT  8352.5 20107.5 8287.5 20242.5 ;
      RECT  8542.5 20107.5 8477.5 20242.5 ;
      RECT  8352.5 20107.5 8287.5 20242.5 ;
      RECT  8162.5 20107.5 8097.5 20242.5 ;
      RECT  8162.5 20107.5 8097.5 20242.5 ;
      RECT  8352.5 20107.5 8287.5 20242.5 ;
      RECT  7992.5 21037.5 7927.5 21172.5 ;
      RECT  7992.5 20062.5 7927.5 20197.5 ;
      RECT  8157.5 20337.5 8292.5 20402.5 ;
      RECT  8415.0 20552.5 8550.0 20617.5 ;
      RECT  8352.5 20947.5 8287.5 21082.5 ;
      RECT  8162.5 20107.5 8097.5 20242.5 ;
      RECT  8062.5 20552.5 8197.5 20617.5 ;
      RECT  8550.0 20552.5 8415.0 20617.5 ;
      RECT  8292.5 20337.5 8157.5 20402.5 ;
      RECT  8197.5 20552.5 8062.5 20617.5 ;
      RECT  8610.0 21257.5 7690.0 21322.5 ;
      RECT  8610.0 19912.5 7690.0 19977.5 ;
      RECT  8542.5 22472.5 8477.5 22667.5 ;
      RECT  8542.5 21632.5 8477.5 21257.5 ;
      RECT  8162.5 21632.5 8097.5 21257.5 ;
      RECT  7992.5 21475.0 7927.5 21290.0 ;
      RECT  7992.5 22635.0 7927.5 22450.0 ;
      RECT  8542.5 21632.5 8477.5 21497.5 ;
      RECT  8352.5 21632.5 8287.5 21497.5 ;
      RECT  8352.5 21632.5 8287.5 21497.5 ;
      RECT  8542.5 21632.5 8477.5 21497.5 ;
      RECT  8352.5 21632.5 8287.5 21497.5 ;
      RECT  8162.5 21632.5 8097.5 21497.5 ;
      RECT  8162.5 21632.5 8097.5 21497.5 ;
      RECT  8352.5 21632.5 8287.5 21497.5 ;
      RECT  8542.5 22472.5 8477.5 22337.5 ;
      RECT  8352.5 22472.5 8287.5 22337.5 ;
      RECT  8352.5 22472.5 8287.5 22337.5 ;
      RECT  8542.5 22472.5 8477.5 22337.5 ;
      RECT  8352.5 22472.5 8287.5 22337.5 ;
      RECT  8162.5 22472.5 8097.5 22337.5 ;
      RECT  8162.5 22472.5 8097.5 22337.5 ;
      RECT  8352.5 22472.5 8287.5 22337.5 ;
      RECT  7992.5 21542.5 7927.5 21407.5 ;
      RECT  7992.5 22517.5 7927.5 22382.5 ;
      RECT  8157.5 22242.5 8292.5 22177.5 ;
      RECT  8415.0 22027.5 8550.0 21962.5 ;
      RECT  8352.5 21632.5 8287.5 21497.5 ;
      RECT  8162.5 22472.5 8097.5 22337.5 ;
      RECT  8062.5 22027.5 8197.5 21962.5 ;
      RECT  8550.0 22027.5 8415.0 21962.5 ;
      RECT  8292.5 22242.5 8157.5 22177.5 ;
      RECT  8197.5 22027.5 8062.5 21962.5 ;
      RECT  8610.0 21322.5 7690.0 21257.5 ;
      RECT  8610.0 22667.5 7690.0 22602.5 ;
      RECT  9607.5 18372.5 9742.5 18437.5 ;
      RECT  10992.5 17850.0 11127.5 17915.0 ;
      RECT  9332.5 19717.5 9467.5 19782.5 ;
      RECT  10717.5 19285.0 10852.5 19350.0 ;
      RECT  10992.5 20047.5 11127.5 20112.5 ;
      RECT  9057.5 20047.5 9192.5 20112.5 ;
      RECT  10717.5 21392.5 10852.5 21457.5 ;
      RECT  8782.5 21392.5 8917.5 21457.5 ;
      RECT  9607.5 17862.5 9742.5 17927.5 ;
      RECT  9332.5 17647.5 9467.5 17712.5 ;
      RECT  9057.5 19272.5 9192.5 19337.5 ;
      RECT  9332.5 19487.5 9467.5 19552.5 ;
      RECT  9607.5 20552.5 9742.5 20617.5 ;
      RECT  8782.5 20337.5 8917.5 20402.5 ;
      RECT  9057.5 21962.5 9192.5 22027.5 ;
      RECT  8782.5 22177.5 8917.5 22242.5 ;
      RECT  7335.0 17850.0 7130.0 17915.0 ;
      RECT  7335.0 19285.0 7130.0 19350.0 ;
      RECT  7335.0 20540.0 7130.0 20605.0 ;
      RECT  7335.0 21975.0 7130.0 22040.0 ;
      RECT  11095.0 18567.5 7130.0 18632.5 ;
      RECT  11095.0 21257.5 7130.0 21322.5 ;
      RECT  11095.0 17222.5 7130.0 17287.5 ;
      RECT  11095.0 19912.5 7130.0 19977.5 ;
      RECT  11095.0 22602.5 7130.0 22667.5 ;
      RECT  9952.5 23230.0 9887.5 23295.0 ;
      RECT  9952.5 23752.5 9887.5 23817.5 ;
      RECT  10190.0 23230.0 9920.0 23295.0 ;
      RECT  9952.5 23262.5 9887.5 23785.0 ;
      RECT  9920.0 23752.5 9675.0 23817.5 ;
      RECT  11060.0 23230.0 10420.0 23295.0 ;
      RECT  9952.5 24665.0 9887.5 24730.0 ;
      RECT  9952.5 25097.5 9887.5 25162.5 ;
      RECT  10190.0 24665.0 9920.0 24730.0 ;
      RECT  9952.5 24697.5 9887.5 25130.0 ;
      RECT  9920.0 25097.5 9400.0 25162.5 ;
      RECT  10785.0 24665.0 10420.0 24730.0 ;
      RECT  11060.0 25427.5 9125.0 25492.5 ;
      RECT  10785.0 26772.5 8850.0 26837.5 ;
      RECT  9675.0 23242.5 8550.0 23307.5 ;
      RECT  9400.0 23027.5 8292.5 23092.5 ;
      RECT  9125.0 24652.5 8550.0 24717.5 ;
      RECT  9400.0 24867.5 8292.5 24932.5 ;
      RECT  9675.0 25932.5 8550.0 25997.5 ;
      RECT  8850.0 25717.5 8292.5 25782.5 ;
      RECT  9125.0 27342.5 8550.0 27407.5 ;
      RECT  8850.0 27557.5 8292.5 27622.5 ;
      RECT  7845.0 23242.5 7780.0 23307.5 ;
      RECT  7845.0 23230.0 7780.0 23295.0 ;
      RECT  8062.5 23242.5 7812.5 23307.5 ;
      RECT  7845.0 23262.5 7780.0 23275.0 ;
      RECT  7812.5 23230.0 7565.0 23295.0 ;
      RECT  7845.0 24652.5 7780.0 24717.5 ;
      RECT  7845.0 24665.0 7780.0 24730.0 ;
      RECT  8062.5 24652.5 7812.5 24717.5 ;
      RECT  7845.0 24685.0 7780.0 24697.5 ;
      RECT  7812.5 24665.0 7565.0 24730.0 ;
      RECT  7845.0 25932.5 7780.0 25997.5 ;
      RECT  7845.0 25920.0 7780.0 25985.0 ;
      RECT  8062.5 25932.5 7812.5 25997.5 ;
      RECT  7845.0 25952.5 7780.0 25965.0 ;
      RECT  7812.5 25920.0 7565.0 25985.0 ;
      RECT  7845.0 27342.5 7780.0 27407.5 ;
      RECT  7845.0 27355.0 7780.0 27420.0 ;
      RECT  8062.5 27342.5 7812.5 27407.5 ;
      RECT  7845.0 27375.0 7780.0 27387.5 ;
      RECT  7812.5 27355.0 7565.0 27420.0 ;
      RECT  10117.5 23795.0 10052.5 23980.0 ;
      RECT  10117.5 22635.0 10052.5 22820.0 ;
      RECT  10477.5 22752.5 10412.5 22602.5 ;
      RECT  10477.5 23637.5 10412.5 24012.5 ;
      RECT  10287.5 22752.5 10222.5 23637.5 ;
      RECT  10477.5 23637.5 10412.5 23772.5 ;
      RECT  10287.5 23637.5 10222.5 23772.5 ;
      RECT  10287.5 23637.5 10222.5 23772.5 ;
      RECT  10477.5 23637.5 10412.5 23772.5 ;
      RECT  10477.5 22752.5 10412.5 22887.5 ;
      RECT  10287.5 22752.5 10222.5 22887.5 ;
      RECT  10287.5 22752.5 10222.5 22887.5 ;
      RECT  10477.5 22752.5 10412.5 22887.5 ;
      RECT  10117.5 23727.5 10052.5 23862.5 ;
      RECT  10117.5 22752.5 10052.5 22887.5 ;
      RECT  10420.0 23195.0 10355.0 23330.0 ;
      RECT  10420.0 23195.0 10355.0 23330.0 ;
      RECT  10255.0 23230.0 10190.0 23295.0 ;
      RECT  10545.0 23947.5 9985.0 24012.5 ;
      RECT  10545.0 22602.5 9985.0 22667.5 ;
      RECT  10117.5 24165.0 10052.5 23980.0 ;
      RECT  10117.5 25325.0 10052.5 25140.0 ;
      RECT  10477.5 25207.5 10412.5 25357.5 ;
      RECT  10477.5 24322.5 10412.5 23947.5 ;
      RECT  10287.5 25207.5 10222.5 24322.5 ;
      RECT  10477.5 24322.5 10412.5 24187.5 ;
      RECT  10287.5 24322.5 10222.5 24187.5 ;
      RECT  10287.5 24322.5 10222.5 24187.5 ;
      RECT  10477.5 24322.5 10412.5 24187.5 ;
      RECT  10477.5 25207.5 10412.5 25072.5 ;
      RECT  10287.5 25207.5 10222.5 25072.5 ;
      RECT  10287.5 25207.5 10222.5 25072.5 ;
      RECT  10477.5 25207.5 10412.5 25072.5 ;
      RECT  10117.5 24232.5 10052.5 24097.5 ;
      RECT  10117.5 25207.5 10052.5 25072.5 ;
      RECT  10420.0 24765.0 10355.0 24630.0 ;
      RECT  10420.0 24765.0 10355.0 24630.0 ;
      RECT  10255.0 24730.0 10190.0 24665.0 ;
      RECT  10545.0 24012.5 9985.0 23947.5 ;
      RECT  10545.0 25357.5 9985.0 25292.5 ;
      RECT  7262.5 23795.0 7197.5 23980.0 ;
      RECT  7262.5 22635.0 7197.5 22820.0 ;
      RECT  7622.5 22752.5 7557.5 22602.5 ;
      RECT  7622.5 23637.5 7557.5 24012.5 ;
      RECT  7432.5 22752.5 7367.5 23637.5 ;
      RECT  7622.5 23637.5 7557.5 23772.5 ;
      RECT  7432.5 23637.5 7367.5 23772.5 ;
      RECT  7432.5 23637.5 7367.5 23772.5 ;
      RECT  7622.5 23637.5 7557.5 23772.5 ;
      RECT  7622.5 22752.5 7557.5 22887.5 ;
      RECT  7432.5 22752.5 7367.5 22887.5 ;
      RECT  7432.5 22752.5 7367.5 22887.5 ;
      RECT  7622.5 22752.5 7557.5 22887.5 ;
      RECT  7262.5 23727.5 7197.5 23862.5 ;
      RECT  7262.5 22752.5 7197.5 22887.5 ;
      RECT  7565.0 23195.0 7500.0 23330.0 ;
      RECT  7565.0 23195.0 7500.0 23330.0 ;
      RECT  7400.0 23230.0 7335.0 23295.0 ;
      RECT  7690.0 23947.5 7130.0 24012.5 ;
      RECT  7690.0 22602.5 7130.0 22667.5 ;
      RECT  7262.5 24165.0 7197.5 23980.0 ;
      RECT  7262.5 25325.0 7197.5 25140.0 ;
      RECT  7622.5 25207.5 7557.5 25357.5 ;
      RECT  7622.5 24322.5 7557.5 23947.5 ;
      RECT  7432.5 25207.5 7367.5 24322.5 ;
      RECT  7622.5 24322.5 7557.5 24187.5 ;
      RECT  7432.5 24322.5 7367.5 24187.5 ;
      RECT  7432.5 24322.5 7367.5 24187.5 ;
      RECT  7622.5 24322.5 7557.5 24187.5 ;
      RECT  7622.5 25207.5 7557.5 25072.5 ;
      RECT  7432.5 25207.5 7367.5 25072.5 ;
      RECT  7432.5 25207.5 7367.5 25072.5 ;
      RECT  7622.5 25207.5 7557.5 25072.5 ;
      RECT  7262.5 24232.5 7197.5 24097.5 ;
      RECT  7262.5 25207.5 7197.5 25072.5 ;
      RECT  7565.0 24765.0 7500.0 24630.0 ;
      RECT  7565.0 24765.0 7500.0 24630.0 ;
      RECT  7400.0 24730.0 7335.0 24665.0 ;
      RECT  7690.0 24012.5 7130.0 23947.5 ;
      RECT  7690.0 25357.5 7130.0 25292.5 ;
      RECT  7262.5 26485.0 7197.5 26670.0 ;
      RECT  7262.5 25325.0 7197.5 25510.0 ;
      RECT  7622.5 25442.5 7557.5 25292.5 ;
      RECT  7622.5 26327.5 7557.5 26702.5 ;
      RECT  7432.5 25442.5 7367.5 26327.5 ;
      RECT  7622.5 26327.5 7557.5 26462.5 ;
      RECT  7432.5 26327.5 7367.5 26462.5 ;
      RECT  7432.5 26327.5 7367.5 26462.5 ;
      RECT  7622.5 26327.5 7557.5 26462.5 ;
      RECT  7622.5 25442.5 7557.5 25577.5 ;
      RECT  7432.5 25442.5 7367.5 25577.5 ;
      RECT  7432.5 25442.5 7367.5 25577.5 ;
      RECT  7622.5 25442.5 7557.5 25577.5 ;
      RECT  7262.5 26417.5 7197.5 26552.5 ;
      RECT  7262.5 25442.5 7197.5 25577.5 ;
      RECT  7565.0 25885.0 7500.0 26020.0 ;
      RECT  7565.0 25885.0 7500.0 26020.0 ;
      RECT  7400.0 25920.0 7335.0 25985.0 ;
      RECT  7690.0 26637.5 7130.0 26702.5 ;
      RECT  7690.0 25292.5 7130.0 25357.5 ;
      RECT  7262.5 26855.0 7197.5 26670.0 ;
      RECT  7262.5 28015.0 7197.5 27830.0 ;
      RECT  7622.5 27897.5 7557.5 28047.5 ;
      RECT  7622.5 27012.5 7557.5 26637.5 ;
      RECT  7432.5 27897.5 7367.5 27012.5 ;
      RECT  7622.5 27012.5 7557.5 26877.5 ;
      RECT  7432.5 27012.5 7367.5 26877.5 ;
      RECT  7432.5 27012.5 7367.5 26877.5 ;
      RECT  7622.5 27012.5 7557.5 26877.5 ;
      RECT  7622.5 27897.5 7557.5 27762.5 ;
      RECT  7432.5 27897.5 7367.5 27762.5 ;
      RECT  7432.5 27897.5 7367.5 27762.5 ;
      RECT  7622.5 27897.5 7557.5 27762.5 ;
      RECT  7262.5 26922.5 7197.5 26787.5 ;
      RECT  7262.5 27897.5 7197.5 27762.5 ;
      RECT  7565.0 27455.0 7500.0 27320.0 ;
      RECT  7565.0 27455.0 7500.0 27320.0 ;
      RECT  7400.0 27420.0 7335.0 27355.0 ;
      RECT  7690.0 26702.5 7130.0 26637.5 ;
      RECT  7690.0 28047.5 7130.0 27982.5 ;
      RECT  8542.5 22797.5 8477.5 22602.5 ;
      RECT  8542.5 23637.5 8477.5 24012.5 ;
      RECT  8162.5 23637.5 8097.5 24012.5 ;
      RECT  7992.5 23795.0 7927.5 23980.0 ;
      RECT  7992.5 22635.0 7927.5 22820.0 ;
      RECT  8542.5 23637.5 8477.5 23772.5 ;
      RECT  8352.5 23637.5 8287.5 23772.5 ;
      RECT  8352.5 23637.5 8287.5 23772.5 ;
      RECT  8542.5 23637.5 8477.5 23772.5 ;
      RECT  8352.5 23637.5 8287.5 23772.5 ;
      RECT  8162.5 23637.5 8097.5 23772.5 ;
      RECT  8162.5 23637.5 8097.5 23772.5 ;
      RECT  8352.5 23637.5 8287.5 23772.5 ;
      RECT  8542.5 22797.5 8477.5 22932.5 ;
      RECT  8352.5 22797.5 8287.5 22932.5 ;
      RECT  8352.5 22797.5 8287.5 22932.5 ;
      RECT  8542.5 22797.5 8477.5 22932.5 ;
      RECT  8352.5 22797.5 8287.5 22932.5 ;
      RECT  8162.5 22797.5 8097.5 22932.5 ;
      RECT  8162.5 22797.5 8097.5 22932.5 ;
      RECT  8352.5 22797.5 8287.5 22932.5 ;
      RECT  7992.5 23727.5 7927.5 23862.5 ;
      RECT  7992.5 22752.5 7927.5 22887.5 ;
      RECT  8157.5 23027.5 8292.5 23092.5 ;
      RECT  8415.0 23242.5 8550.0 23307.5 ;
      RECT  8352.5 23637.5 8287.5 23772.5 ;
      RECT  8162.5 22797.5 8097.5 22932.5 ;
      RECT  8062.5 23242.5 8197.5 23307.5 ;
      RECT  8550.0 23242.5 8415.0 23307.5 ;
      RECT  8292.5 23027.5 8157.5 23092.5 ;
      RECT  8197.5 23242.5 8062.5 23307.5 ;
      RECT  8610.0 23947.5 7690.0 24012.5 ;
      RECT  8610.0 22602.5 7690.0 22667.5 ;
      RECT  8542.5 25162.5 8477.5 25357.5 ;
      RECT  8542.5 24322.5 8477.5 23947.5 ;
      RECT  8162.5 24322.5 8097.5 23947.5 ;
      RECT  7992.5 24165.0 7927.5 23980.0 ;
      RECT  7992.5 25325.0 7927.5 25140.0 ;
      RECT  8542.5 24322.5 8477.5 24187.5 ;
      RECT  8352.5 24322.5 8287.5 24187.5 ;
      RECT  8352.5 24322.5 8287.5 24187.5 ;
      RECT  8542.5 24322.5 8477.5 24187.5 ;
      RECT  8352.5 24322.5 8287.5 24187.5 ;
      RECT  8162.5 24322.5 8097.5 24187.5 ;
      RECT  8162.5 24322.5 8097.5 24187.5 ;
      RECT  8352.5 24322.5 8287.5 24187.5 ;
      RECT  8542.5 25162.5 8477.5 25027.5 ;
      RECT  8352.5 25162.5 8287.5 25027.5 ;
      RECT  8352.5 25162.5 8287.5 25027.5 ;
      RECT  8542.5 25162.5 8477.5 25027.5 ;
      RECT  8352.5 25162.5 8287.5 25027.5 ;
      RECT  8162.5 25162.5 8097.5 25027.5 ;
      RECT  8162.5 25162.5 8097.5 25027.5 ;
      RECT  8352.5 25162.5 8287.5 25027.5 ;
      RECT  7992.5 24232.5 7927.5 24097.5 ;
      RECT  7992.5 25207.5 7927.5 25072.5 ;
      RECT  8157.5 24932.5 8292.5 24867.5 ;
      RECT  8415.0 24717.5 8550.0 24652.5 ;
      RECT  8352.5 24322.5 8287.5 24187.5 ;
      RECT  8162.5 25162.5 8097.5 25027.5 ;
      RECT  8062.5 24717.5 8197.5 24652.5 ;
      RECT  8550.0 24717.5 8415.0 24652.5 ;
      RECT  8292.5 24932.5 8157.5 24867.5 ;
      RECT  8197.5 24717.5 8062.5 24652.5 ;
      RECT  8610.0 24012.5 7690.0 23947.5 ;
      RECT  8610.0 25357.5 7690.0 25292.5 ;
      RECT  8542.5 25487.5 8477.5 25292.5 ;
      RECT  8542.5 26327.5 8477.5 26702.5 ;
      RECT  8162.5 26327.5 8097.5 26702.5 ;
      RECT  7992.5 26485.0 7927.5 26670.0 ;
      RECT  7992.5 25325.0 7927.5 25510.0 ;
      RECT  8542.5 26327.5 8477.5 26462.5 ;
      RECT  8352.5 26327.5 8287.5 26462.5 ;
      RECT  8352.5 26327.5 8287.5 26462.5 ;
      RECT  8542.5 26327.5 8477.5 26462.5 ;
      RECT  8352.5 26327.5 8287.5 26462.5 ;
      RECT  8162.5 26327.5 8097.5 26462.5 ;
      RECT  8162.5 26327.5 8097.5 26462.5 ;
      RECT  8352.5 26327.5 8287.5 26462.5 ;
      RECT  8542.5 25487.5 8477.5 25622.5 ;
      RECT  8352.5 25487.5 8287.5 25622.5 ;
      RECT  8352.5 25487.5 8287.5 25622.5 ;
      RECT  8542.5 25487.5 8477.5 25622.5 ;
      RECT  8352.5 25487.5 8287.5 25622.5 ;
      RECT  8162.5 25487.5 8097.5 25622.5 ;
      RECT  8162.5 25487.5 8097.5 25622.5 ;
      RECT  8352.5 25487.5 8287.5 25622.5 ;
      RECT  7992.5 26417.5 7927.5 26552.5 ;
      RECT  7992.5 25442.5 7927.5 25577.5 ;
      RECT  8157.5 25717.5 8292.5 25782.5 ;
      RECT  8415.0 25932.5 8550.0 25997.5 ;
      RECT  8352.5 26327.5 8287.5 26462.5 ;
      RECT  8162.5 25487.5 8097.5 25622.5 ;
      RECT  8062.5 25932.5 8197.5 25997.5 ;
      RECT  8550.0 25932.5 8415.0 25997.5 ;
      RECT  8292.5 25717.5 8157.5 25782.5 ;
      RECT  8197.5 25932.5 8062.5 25997.5 ;
      RECT  8610.0 26637.5 7690.0 26702.5 ;
      RECT  8610.0 25292.5 7690.0 25357.5 ;
      RECT  8542.5 27852.5 8477.5 28047.5 ;
      RECT  8542.5 27012.5 8477.5 26637.5 ;
      RECT  8162.5 27012.5 8097.5 26637.5 ;
      RECT  7992.5 26855.0 7927.5 26670.0 ;
      RECT  7992.5 28015.0 7927.5 27830.0 ;
      RECT  8542.5 27012.5 8477.5 26877.5 ;
      RECT  8352.5 27012.5 8287.5 26877.5 ;
      RECT  8352.5 27012.5 8287.5 26877.5 ;
      RECT  8542.5 27012.5 8477.5 26877.5 ;
      RECT  8352.5 27012.5 8287.5 26877.5 ;
      RECT  8162.5 27012.5 8097.5 26877.5 ;
      RECT  8162.5 27012.5 8097.5 26877.5 ;
      RECT  8352.5 27012.5 8287.5 26877.5 ;
      RECT  8542.5 27852.5 8477.5 27717.5 ;
      RECT  8352.5 27852.5 8287.5 27717.5 ;
      RECT  8352.5 27852.5 8287.5 27717.5 ;
      RECT  8542.5 27852.5 8477.5 27717.5 ;
      RECT  8352.5 27852.5 8287.5 27717.5 ;
      RECT  8162.5 27852.5 8097.5 27717.5 ;
      RECT  8162.5 27852.5 8097.5 27717.5 ;
      RECT  8352.5 27852.5 8287.5 27717.5 ;
      RECT  7992.5 26922.5 7927.5 26787.5 ;
      RECT  7992.5 27897.5 7927.5 27762.5 ;
      RECT  8157.5 27622.5 8292.5 27557.5 ;
      RECT  8415.0 27407.5 8550.0 27342.5 ;
      RECT  8352.5 27012.5 8287.5 26877.5 ;
      RECT  8162.5 27852.5 8097.5 27717.5 ;
      RECT  8062.5 27407.5 8197.5 27342.5 ;
      RECT  8550.0 27407.5 8415.0 27342.5 ;
      RECT  8292.5 27622.5 8157.5 27557.5 ;
      RECT  8197.5 27407.5 8062.5 27342.5 ;
      RECT  8610.0 26702.5 7690.0 26637.5 ;
      RECT  8610.0 28047.5 7690.0 27982.5 ;
      RECT  9607.5 23752.5 9742.5 23817.5 ;
      RECT  10992.5 23230.0 11127.5 23295.0 ;
      RECT  9332.5 25097.5 9467.5 25162.5 ;
      RECT  10717.5 24665.0 10852.5 24730.0 ;
      RECT  10992.5 25427.5 11127.5 25492.5 ;
      RECT  9057.5 25427.5 9192.5 25492.5 ;
      RECT  10717.5 26772.5 10852.5 26837.5 ;
      RECT  8782.5 26772.5 8917.5 26837.5 ;
      RECT  9607.5 23242.5 9742.5 23307.5 ;
      RECT  9332.5 23027.5 9467.5 23092.5 ;
      RECT  9057.5 24652.5 9192.5 24717.5 ;
      RECT  9332.5 24867.5 9467.5 24932.5 ;
      RECT  9607.5 25932.5 9742.5 25997.5 ;
      RECT  8782.5 25717.5 8917.5 25782.5 ;
      RECT  9057.5 27342.5 9192.5 27407.5 ;
      RECT  8782.5 27557.5 8917.5 27622.5 ;
      RECT  7335.0 23230.0 7130.0 23295.0 ;
      RECT  7335.0 24665.0 7130.0 24730.0 ;
      RECT  7335.0 25920.0 7130.0 25985.0 ;
      RECT  7335.0 27355.0 7130.0 27420.0 ;
      RECT  11095.0 23947.5 7130.0 24012.5 ;
      RECT  11095.0 26637.5 7130.0 26702.5 ;
      RECT  11095.0 22602.5 7130.0 22667.5 ;
      RECT  11095.0 25292.5 7130.0 25357.5 ;
      RECT  11095.0 27982.5 7130.0 28047.5 ;
      RECT  7197.5 28177.5 7262.5 27982.5 ;
      RECT  7197.5 29017.5 7262.5 29392.5 ;
      RECT  7577.5 29017.5 7642.5 29392.5 ;
      RECT  7937.5 29175.0 8002.5 29360.0 ;
      RECT  7937.5 28015.0 8002.5 28200.0 ;
      RECT  7197.5 29017.5 7262.5 29152.5 ;
      RECT  7387.5 29017.5 7452.5 29152.5 ;
      RECT  7387.5 29017.5 7452.5 29152.5 ;
      RECT  7197.5 29017.5 7262.5 29152.5 ;
      RECT  7387.5 29017.5 7452.5 29152.5 ;
      RECT  7577.5 29017.5 7642.5 29152.5 ;
      RECT  7577.5 29017.5 7642.5 29152.5 ;
      RECT  7387.5 29017.5 7452.5 29152.5 ;
      RECT  7577.5 29017.5 7642.5 29152.5 ;
      RECT  7767.5 29017.5 7832.5 29152.5 ;
      RECT  7767.5 29017.5 7832.5 29152.5 ;
      RECT  7577.5 29017.5 7642.5 29152.5 ;
      RECT  7197.5 28177.5 7262.5 28312.5 ;
      RECT  7387.5 28177.5 7452.5 28312.5 ;
      RECT  7387.5 28177.5 7452.5 28312.5 ;
      RECT  7197.5 28177.5 7262.5 28312.5 ;
      RECT  7387.5 28177.5 7452.5 28312.5 ;
      RECT  7577.5 28177.5 7642.5 28312.5 ;
      RECT  7577.5 28177.5 7642.5 28312.5 ;
      RECT  7387.5 28177.5 7452.5 28312.5 ;
      RECT  7577.5 28177.5 7642.5 28312.5 ;
      RECT  7767.5 28177.5 7832.5 28312.5 ;
      RECT  7767.5 28177.5 7832.5 28312.5 ;
      RECT  7577.5 28177.5 7642.5 28312.5 ;
      RECT  7937.5 29107.5 8002.5 29242.5 ;
      RECT  7937.5 28132.5 8002.5 28267.5 ;
      RECT  7772.5 28390.0 7637.5 28455.0 ;
      RECT  7582.5 28530.0 7447.5 28595.0 ;
      RECT  7392.5 28670.0 7257.5 28735.0 ;
      RECT  7387.5 29017.5 7452.5 29152.5 ;
      RECT  7767.5 29017.5 7832.5 29152.5 ;
      RECT  7767.5 28177.5 7832.5 28312.5 ;
      RECT  7767.5 28635.0 7832.5 28770.0 ;
      RECT  7257.5 28670.0 7392.5 28735.0 ;
      RECT  7447.5 28530.0 7582.5 28595.0 ;
      RECT  7637.5 28390.0 7772.5 28455.0 ;
      RECT  7767.5 28635.0 7832.5 28770.0 ;
      RECT  7130.0 29327.5 8140.0 29392.5 ;
      RECT  7130.0 27982.5 8140.0 28047.5 ;
      RECT  7197.5 30542.5 7262.5 30737.5 ;
      RECT  7197.5 29702.5 7262.5 29327.5 ;
      RECT  7577.5 29702.5 7642.5 29327.5 ;
      RECT  7937.5 29545.0 8002.5 29360.0 ;
      RECT  7937.5 30705.0 8002.5 30520.0 ;
      RECT  7197.5 29702.5 7262.5 29567.5 ;
      RECT  7387.5 29702.5 7452.5 29567.5 ;
      RECT  7387.5 29702.5 7452.5 29567.5 ;
      RECT  7197.5 29702.5 7262.5 29567.5 ;
      RECT  7387.5 29702.5 7452.5 29567.5 ;
      RECT  7577.5 29702.5 7642.5 29567.5 ;
      RECT  7577.5 29702.5 7642.5 29567.5 ;
      RECT  7387.5 29702.5 7452.5 29567.5 ;
      RECT  7577.5 29702.5 7642.5 29567.5 ;
      RECT  7767.5 29702.5 7832.5 29567.5 ;
      RECT  7767.5 29702.5 7832.5 29567.5 ;
      RECT  7577.5 29702.5 7642.5 29567.5 ;
      RECT  7197.5 30542.5 7262.5 30407.5 ;
      RECT  7387.5 30542.5 7452.5 30407.5 ;
      RECT  7387.5 30542.5 7452.5 30407.5 ;
      RECT  7197.5 30542.5 7262.5 30407.5 ;
      RECT  7387.5 30542.5 7452.5 30407.5 ;
      RECT  7577.5 30542.5 7642.5 30407.5 ;
      RECT  7577.5 30542.5 7642.5 30407.5 ;
      RECT  7387.5 30542.5 7452.5 30407.5 ;
      RECT  7577.5 30542.5 7642.5 30407.5 ;
      RECT  7767.5 30542.5 7832.5 30407.5 ;
      RECT  7767.5 30542.5 7832.5 30407.5 ;
      RECT  7577.5 30542.5 7642.5 30407.5 ;
      RECT  7937.5 29612.5 8002.5 29477.5 ;
      RECT  7937.5 30587.5 8002.5 30452.5 ;
      RECT  7772.5 30330.0 7637.5 30265.0 ;
      RECT  7582.5 30190.0 7447.5 30125.0 ;
      RECT  7392.5 30050.0 7257.5 29985.0 ;
      RECT  7387.5 29702.5 7452.5 29567.5 ;
      RECT  7767.5 29702.5 7832.5 29567.5 ;
      RECT  7767.5 30542.5 7832.5 30407.5 ;
      RECT  7767.5 30085.0 7832.5 29950.0 ;
      RECT  7257.5 30050.0 7392.5 29985.0 ;
      RECT  7447.5 30190.0 7582.5 30125.0 ;
      RECT  7637.5 30330.0 7772.5 30265.0 ;
      RECT  7767.5 30085.0 7832.5 29950.0 ;
      RECT  7130.0 29392.5 8140.0 29327.5 ;
      RECT  7130.0 30737.5 8140.0 30672.5 ;
      RECT  7197.5 30867.5 7262.5 30672.5 ;
      RECT  7197.5 31707.5 7262.5 32082.5 ;
      RECT  7577.5 31707.5 7642.5 32082.5 ;
      RECT  7937.5 31865.0 8002.5 32050.0 ;
      RECT  7937.5 30705.0 8002.5 30890.0 ;
      RECT  7197.5 31707.5 7262.5 31842.5 ;
      RECT  7387.5 31707.5 7452.5 31842.5 ;
      RECT  7387.5 31707.5 7452.5 31842.5 ;
      RECT  7197.5 31707.5 7262.5 31842.5 ;
      RECT  7387.5 31707.5 7452.5 31842.5 ;
      RECT  7577.5 31707.5 7642.5 31842.5 ;
      RECT  7577.5 31707.5 7642.5 31842.5 ;
      RECT  7387.5 31707.5 7452.5 31842.5 ;
      RECT  7577.5 31707.5 7642.5 31842.5 ;
      RECT  7767.5 31707.5 7832.5 31842.5 ;
      RECT  7767.5 31707.5 7832.5 31842.5 ;
      RECT  7577.5 31707.5 7642.5 31842.5 ;
      RECT  7197.5 30867.5 7262.5 31002.5 ;
      RECT  7387.5 30867.5 7452.5 31002.5 ;
      RECT  7387.5 30867.5 7452.5 31002.5 ;
      RECT  7197.5 30867.5 7262.5 31002.5 ;
      RECT  7387.5 30867.5 7452.5 31002.5 ;
      RECT  7577.5 30867.5 7642.5 31002.5 ;
      RECT  7577.5 30867.5 7642.5 31002.5 ;
      RECT  7387.5 30867.5 7452.5 31002.5 ;
      RECT  7577.5 30867.5 7642.5 31002.5 ;
      RECT  7767.5 30867.5 7832.5 31002.5 ;
      RECT  7767.5 30867.5 7832.5 31002.5 ;
      RECT  7577.5 30867.5 7642.5 31002.5 ;
      RECT  7937.5 31797.5 8002.5 31932.5 ;
      RECT  7937.5 30822.5 8002.5 30957.5 ;
      RECT  7772.5 31080.0 7637.5 31145.0 ;
      RECT  7582.5 31220.0 7447.5 31285.0 ;
      RECT  7392.5 31360.0 7257.5 31425.0 ;
      RECT  7387.5 31707.5 7452.5 31842.5 ;
      RECT  7767.5 31707.5 7832.5 31842.5 ;
      RECT  7767.5 30867.5 7832.5 31002.5 ;
      RECT  7767.5 31325.0 7832.5 31460.0 ;
      RECT  7257.5 31360.0 7392.5 31425.0 ;
      RECT  7447.5 31220.0 7582.5 31285.0 ;
      RECT  7637.5 31080.0 7772.5 31145.0 ;
      RECT  7767.5 31325.0 7832.5 31460.0 ;
      RECT  7130.0 32017.5 8140.0 32082.5 ;
      RECT  7130.0 30672.5 8140.0 30737.5 ;
      RECT  7197.5 33232.5 7262.5 33427.5 ;
      RECT  7197.5 32392.5 7262.5 32017.5 ;
      RECT  7577.5 32392.5 7642.5 32017.5 ;
      RECT  7937.5 32235.0 8002.5 32050.0 ;
      RECT  7937.5 33395.0 8002.5 33210.0 ;
      RECT  7197.5 32392.5 7262.5 32257.5 ;
      RECT  7387.5 32392.5 7452.5 32257.5 ;
      RECT  7387.5 32392.5 7452.5 32257.5 ;
      RECT  7197.5 32392.5 7262.5 32257.5 ;
      RECT  7387.5 32392.5 7452.5 32257.5 ;
      RECT  7577.5 32392.5 7642.5 32257.5 ;
      RECT  7577.5 32392.5 7642.5 32257.5 ;
      RECT  7387.5 32392.5 7452.5 32257.5 ;
      RECT  7577.5 32392.5 7642.5 32257.5 ;
      RECT  7767.5 32392.5 7832.5 32257.5 ;
      RECT  7767.5 32392.5 7832.5 32257.5 ;
      RECT  7577.5 32392.5 7642.5 32257.5 ;
      RECT  7197.5 33232.5 7262.5 33097.5 ;
      RECT  7387.5 33232.5 7452.5 33097.5 ;
      RECT  7387.5 33232.5 7452.5 33097.5 ;
      RECT  7197.5 33232.5 7262.5 33097.5 ;
      RECT  7387.5 33232.5 7452.5 33097.5 ;
      RECT  7577.5 33232.5 7642.5 33097.5 ;
      RECT  7577.5 33232.5 7642.5 33097.5 ;
      RECT  7387.5 33232.5 7452.5 33097.5 ;
      RECT  7577.5 33232.5 7642.5 33097.5 ;
      RECT  7767.5 33232.5 7832.5 33097.5 ;
      RECT  7767.5 33232.5 7832.5 33097.5 ;
      RECT  7577.5 33232.5 7642.5 33097.5 ;
      RECT  7937.5 32302.5 8002.5 32167.5 ;
      RECT  7937.5 33277.5 8002.5 33142.5 ;
      RECT  7772.5 33020.0 7637.5 32955.0 ;
      RECT  7582.5 32880.0 7447.5 32815.0 ;
      RECT  7392.5 32740.0 7257.5 32675.0 ;
      RECT  7387.5 32392.5 7452.5 32257.5 ;
      RECT  7767.5 32392.5 7832.5 32257.5 ;
      RECT  7767.5 33232.5 7832.5 33097.5 ;
      RECT  7767.5 32775.0 7832.5 32640.0 ;
      RECT  7257.5 32740.0 7392.5 32675.0 ;
      RECT  7447.5 32880.0 7582.5 32815.0 ;
      RECT  7637.5 33020.0 7772.5 32955.0 ;
      RECT  7767.5 32775.0 7832.5 32640.0 ;
      RECT  7130.0 32082.5 8140.0 32017.5 ;
      RECT  7130.0 33427.5 8140.0 33362.5 ;
      RECT  7197.5 33557.5 7262.5 33362.5 ;
      RECT  7197.5 34397.5 7262.5 34772.5 ;
      RECT  7577.5 34397.5 7642.5 34772.5 ;
      RECT  7937.5 34555.0 8002.5 34740.0 ;
      RECT  7937.5 33395.0 8002.5 33580.0 ;
      RECT  7197.5 34397.5 7262.5 34532.5 ;
      RECT  7387.5 34397.5 7452.5 34532.5 ;
      RECT  7387.5 34397.5 7452.5 34532.5 ;
      RECT  7197.5 34397.5 7262.5 34532.5 ;
      RECT  7387.5 34397.5 7452.5 34532.5 ;
      RECT  7577.5 34397.5 7642.5 34532.5 ;
      RECT  7577.5 34397.5 7642.5 34532.5 ;
      RECT  7387.5 34397.5 7452.5 34532.5 ;
      RECT  7577.5 34397.5 7642.5 34532.5 ;
      RECT  7767.5 34397.5 7832.5 34532.5 ;
      RECT  7767.5 34397.5 7832.5 34532.5 ;
      RECT  7577.5 34397.5 7642.5 34532.5 ;
      RECT  7197.5 33557.5 7262.5 33692.5 ;
      RECT  7387.5 33557.5 7452.5 33692.5 ;
      RECT  7387.5 33557.5 7452.5 33692.5 ;
      RECT  7197.5 33557.5 7262.5 33692.5 ;
      RECT  7387.5 33557.5 7452.5 33692.5 ;
      RECT  7577.5 33557.5 7642.5 33692.5 ;
      RECT  7577.5 33557.5 7642.5 33692.5 ;
      RECT  7387.5 33557.5 7452.5 33692.5 ;
      RECT  7577.5 33557.5 7642.5 33692.5 ;
      RECT  7767.5 33557.5 7832.5 33692.5 ;
      RECT  7767.5 33557.5 7832.5 33692.5 ;
      RECT  7577.5 33557.5 7642.5 33692.5 ;
      RECT  7937.5 34487.5 8002.5 34622.5 ;
      RECT  7937.5 33512.5 8002.5 33647.5 ;
      RECT  7772.5 33770.0 7637.5 33835.0 ;
      RECT  7582.5 33910.0 7447.5 33975.0 ;
      RECT  7392.5 34050.0 7257.5 34115.0 ;
      RECT  7387.5 34397.5 7452.5 34532.5 ;
      RECT  7767.5 34397.5 7832.5 34532.5 ;
      RECT  7767.5 33557.5 7832.5 33692.5 ;
      RECT  7767.5 34015.0 7832.5 34150.0 ;
      RECT  7257.5 34050.0 7392.5 34115.0 ;
      RECT  7447.5 33910.0 7582.5 33975.0 ;
      RECT  7637.5 33770.0 7772.5 33835.0 ;
      RECT  7767.5 34015.0 7832.5 34150.0 ;
      RECT  7130.0 34707.5 8140.0 34772.5 ;
      RECT  7130.0 33362.5 8140.0 33427.5 ;
      RECT  7197.5 35922.5 7262.5 36117.5 ;
      RECT  7197.5 35082.5 7262.5 34707.5 ;
      RECT  7577.5 35082.5 7642.5 34707.5 ;
      RECT  7937.5 34925.0 8002.5 34740.0 ;
      RECT  7937.5 36085.0 8002.5 35900.0 ;
      RECT  7197.5 35082.5 7262.5 34947.5 ;
      RECT  7387.5 35082.5 7452.5 34947.5 ;
      RECT  7387.5 35082.5 7452.5 34947.5 ;
      RECT  7197.5 35082.5 7262.5 34947.5 ;
      RECT  7387.5 35082.5 7452.5 34947.5 ;
      RECT  7577.5 35082.5 7642.5 34947.5 ;
      RECT  7577.5 35082.5 7642.5 34947.5 ;
      RECT  7387.5 35082.5 7452.5 34947.5 ;
      RECT  7577.5 35082.5 7642.5 34947.5 ;
      RECT  7767.5 35082.5 7832.5 34947.5 ;
      RECT  7767.5 35082.5 7832.5 34947.5 ;
      RECT  7577.5 35082.5 7642.5 34947.5 ;
      RECT  7197.5 35922.5 7262.5 35787.5 ;
      RECT  7387.5 35922.5 7452.5 35787.5 ;
      RECT  7387.5 35922.5 7452.5 35787.5 ;
      RECT  7197.5 35922.5 7262.5 35787.5 ;
      RECT  7387.5 35922.5 7452.5 35787.5 ;
      RECT  7577.5 35922.5 7642.5 35787.5 ;
      RECT  7577.5 35922.5 7642.5 35787.5 ;
      RECT  7387.5 35922.5 7452.5 35787.5 ;
      RECT  7577.5 35922.5 7642.5 35787.5 ;
      RECT  7767.5 35922.5 7832.5 35787.5 ;
      RECT  7767.5 35922.5 7832.5 35787.5 ;
      RECT  7577.5 35922.5 7642.5 35787.5 ;
      RECT  7937.5 34992.5 8002.5 34857.5 ;
      RECT  7937.5 35967.5 8002.5 35832.5 ;
      RECT  7772.5 35710.0 7637.5 35645.0 ;
      RECT  7582.5 35570.0 7447.5 35505.0 ;
      RECT  7392.5 35430.0 7257.5 35365.0 ;
      RECT  7387.5 35082.5 7452.5 34947.5 ;
      RECT  7767.5 35082.5 7832.5 34947.5 ;
      RECT  7767.5 35922.5 7832.5 35787.5 ;
      RECT  7767.5 35465.0 7832.5 35330.0 ;
      RECT  7257.5 35430.0 7392.5 35365.0 ;
      RECT  7447.5 35570.0 7582.5 35505.0 ;
      RECT  7637.5 35710.0 7772.5 35645.0 ;
      RECT  7767.5 35465.0 7832.5 35330.0 ;
      RECT  7130.0 34772.5 8140.0 34707.5 ;
      RECT  7130.0 36117.5 8140.0 36052.5 ;
      RECT  7197.5 36247.5 7262.5 36052.5 ;
      RECT  7197.5 37087.5 7262.5 37462.5 ;
      RECT  7577.5 37087.5 7642.5 37462.5 ;
      RECT  7937.5 37245.0 8002.5 37430.0 ;
      RECT  7937.5 36085.0 8002.5 36270.0 ;
      RECT  7197.5 37087.5 7262.5 37222.5 ;
      RECT  7387.5 37087.5 7452.5 37222.5 ;
      RECT  7387.5 37087.5 7452.5 37222.5 ;
      RECT  7197.5 37087.5 7262.5 37222.5 ;
      RECT  7387.5 37087.5 7452.5 37222.5 ;
      RECT  7577.5 37087.5 7642.5 37222.5 ;
      RECT  7577.5 37087.5 7642.5 37222.5 ;
      RECT  7387.5 37087.5 7452.5 37222.5 ;
      RECT  7577.5 37087.5 7642.5 37222.5 ;
      RECT  7767.5 37087.5 7832.5 37222.5 ;
      RECT  7767.5 37087.5 7832.5 37222.5 ;
      RECT  7577.5 37087.5 7642.5 37222.5 ;
      RECT  7197.5 36247.5 7262.5 36382.5 ;
      RECT  7387.5 36247.5 7452.5 36382.5 ;
      RECT  7387.5 36247.5 7452.5 36382.5 ;
      RECT  7197.5 36247.5 7262.5 36382.5 ;
      RECT  7387.5 36247.5 7452.5 36382.5 ;
      RECT  7577.5 36247.5 7642.5 36382.5 ;
      RECT  7577.5 36247.5 7642.5 36382.5 ;
      RECT  7387.5 36247.5 7452.5 36382.5 ;
      RECT  7577.5 36247.5 7642.5 36382.5 ;
      RECT  7767.5 36247.5 7832.5 36382.5 ;
      RECT  7767.5 36247.5 7832.5 36382.5 ;
      RECT  7577.5 36247.5 7642.5 36382.5 ;
      RECT  7937.5 37177.5 8002.5 37312.5 ;
      RECT  7937.5 36202.5 8002.5 36337.5 ;
      RECT  7772.5 36460.0 7637.5 36525.0 ;
      RECT  7582.5 36600.0 7447.5 36665.0 ;
      RECT  7392.5 36740.0 7257.5 36805.0 ;
      RECT  7387.5 37087.5 7452.5 37222.5 ;
      RECT  7767.5 37087.5 7832.5 37222.5 ;
      RECT  7767.5 36247.5 7832.5 36382.5 ;
      RECT  7767.5 36705.0 7832.5 36840.0 ;
      RECT  7257.5 36740.0 7392.5 36805.0 ;
      RECT  7447.5 36600.0 7582.5 36665.0 ;
      RECT  7637.5 36460.0 7772.5 36525.0 ;
      RECT  7767.5 36705.0 7832.5 36840.0 ;
      RECT  7130.0 37397.5 8140.0 37462.5 ;
      RECT  7130.0 36052.5 8140.0 36117.5 ;
      RECT  7197.5 38612.5 7262.5 38807.5 ;
      RECT  7197.5 37772.5 7262.5 37397.5 ;
      RECT  7577.5 37772.5 7642.5 37397.5 ;
      RECT  7937.5 37615.0 8002.5 37430.0 ;
      RECT  7937.5 38775.0 8002.5 38590.0 ;
      RECT  7197.5 37772.5 7262.5 37637.5 ;
      RECT  7387.5 37772.5 7452.5 37637.5 ;
      RECT  7387.5 37772.5 7452.5 37637.5 ;
      RECT  7197.5 37772.5 7262.5 37637.5 ;
      RECT  7387.5 37772.5 7452.5 37637.5 ;
      RECT  7577.5 37772.5 7642.5 37637.5 ;
      RECT  7577.5 37772.5 7642.5 37637.5 ;
      RECT  7387.5 37772.5 7452.5 37637.5 ;
      RECT  7577.5 37772.5 7642.5 37637.5 ;
      RECT  7767.5 37772.5 7832.5 37637.5 ;
      RECT  7767.5 37772.5 7832.5 37637.5 ;
      RECT  7577.5 37772.5 7642.5 37637.5 ;
      RECT  7197.5 38612.5 7262.5 38477.5 ;
      RECT  7387.5 38612.5 7452.5 38477.5 ;
      RECT  7387.5 38612.5 7452.5 38477.5 ;
      RECT  7197.5 38612.5 7262.5 38477.5 ;
      RECT  7387.5 38612.5 7452.5 38477.5 ;
      RECT  7577.5 38612.5 7642.5 38477.5 ;
      RECT  7577.5 38612.5 7642.5 38477.5 ;
      RECT  7387.5 38612.5 7452.5 38477.5 ;
      RECT  7577.5 38612.5 7642.5 38477.5 ;
      RECT  7767.5 38612.5 7832.5 38477.5 ;
      RECT  7767.5 38612.5 7832.5 38477.5 ;
      RECT  7577.5 38612.5 7642.5 38477.5 ;
      RECT  7937.5 37682.5 8002.5 37547.5 ;
      RECT  7937.5 38657.5 8002.5 38522.5 ;
      RECT  7772.5 38400.0 7637.5 38335.0 ;
      RECT  7582.5 38260.0 7447.5 38195.0 ;
      RECT  7392.5 38120.0 7257.5 38055.0 ;
      RECT  7387.5 37772.5 7452.5 37637.5 ;
      RECT  7767.5 37772.5 7832.5 37637.5 ;
      RECT  7767.5 38612.5 7832.5 38477.5 ;
      RECT  7767.5 38155.0 7832.5 38020.0 ;
      RECT  7257.5 38120.0 7392.5 38055.0 ;
      RECT  7447.5 38260.0 7582.5 38195.0 ;
      RECT  7637.5 38400.0 7772.5 38335.0 ;
      RECT  7767.5 38155.0 7832.5 38020.0 ;
      RECT  7130.0 37462.5 8140.0 37397.5 ;
      RECT  7130.0 38807.5 8140.0 38742.5 ;
      RECT  7197.5 38937.5 7262.5 38742.5 ;
      RECT  7197.5 39777.5 7262.5 40152.5 ;
      RECT  7577.5 39777.5 7642.5 40152.5 ;
      RECT  7937.5 39935.0 8002.5 40120.0 ;
      RECT  7937.5 38775.0 8002.5 38960.0 ;
      RECT  7197.5 39777.5 7262.5 39912.5 ;
      RECT  7387.5 39777.5 7452.5 39912.5 ;
      RECT  7387.5 39777.5 7452.5 39912.5 ;
      RECT  7197.5 39777.5 7262.5 39912.5 ;
      RECT  7387.5 39777.5 7452.5 39912.5 ;
      RECT  7577.5 39777.5 7642.5 39912.5 ;
      RECT  7577.5 39777.5 7642.5 39912.5 ;
      RECT  7387.5 39777.5 7452.5 39912.5 ;
      RECT  7577.5 39777.5 7642.5 39912.5 ;
      RECT  7767.5 39777.5 7832.5 39912.5 ;
      RECT  7767.5 39777.5 7832.5 39912.5 ;
      RECT  7577.5 39777.5 7642.5 39912.5 ;
      RECT  7197.5 38937.5 7262.5 39072.5 ;
      RECT  7387.5 38937.5 7452.5 39072.5 ;
      RECT  7387.5 38937.5 7452.5 39072.5 ;
      RECT  7197.5 38937.5 7262.5 39072.5 ;
      RECT  7387.5 38937.5 7452.5 39072.5 ;
      RECT  7577.5 38937.5 7642.5 39072.5 ;
      RECT  7577.5 38937.5 7642.5 39072.5 ;
      RECT  7387.5 38937.5 7452.5 39072.5 ;
      RECT  7577.5 38937.5 7642.5 39072.5 ;
      RECT  7767.5 38937.5 7832.5 39072.5 ;
      RECT  7767.5 38937.5 7832.5 39072.5 ;
      RECT  7577.5 38937.5 7642.5 39072.5 ;
      RECT  7937.5 39867.5 8002.5 40002.5 ;
      RECT  7937.5 38892.5 8002.5 39027.5 ;
      RECT  7772.5 39150.0 7637.5 39215.0 ;
      RECT  7582.5 39290.0 7447.5 39355.0 ;
      RECT  7392.5 39430.0 7257.5 39495.0 ;
      RECT  7387.5 39777.5 7452.5 39912.5 ;
      RECT  7767.5 39777.5 7832.5 39912.5 ;
      RECT  7767.5 38937.5 7832.5 39072.5 ;
      RECT  7767.5 39395.0 7832.5 39530.0 ;
      RECT  7257.5 39430.0 7392.5 39495.0 ;
      RECT  7447.5 39290.0 7582.5 39355.0 ;
      RECT  7637.5 39150.0 7772.5 39215.0 ;
      RECT  7767.5 39395.0 7832.5 39530.0 ;
      RECT  7130.0 40087.5 8140.0 40152.5 ;
      RECT  7130.0 38742.5 8140.0 38807.5 ;
      RECT  7197.5 41302.5 7262.5 41497.5 ;
      RECT  7197.5 40462.5 7262.5 40087.5 ;
      RECT  7577.5 40462.5 7642.5 40087.5 ;
      RECT  7937.5 40305.0 8002.5 40120.0 ;
      RECT  7937.5 41465.0 8002.5 41280.0 ;
      RECT  7197.5 40462.5 7262.5 40327.5 ;
      RECT  7387.5 40462.5 7452.5 40327.5 ;
      RECT  7387.5 40462.5 7452.5 40327.5 ;
      RECT  7197.5 40462.5 7262.5 40327.5 ;
      RECT  7387.5 40462.5 7452.5 40327.5 ;
      RECT  7577.5 40462.5 7642.5 40327.5 ;
      RECT  7577.5 40462.5 7642.5 40327.5 ;
      RECT  7387.5 40462.5 7452.5 40327.5 ;
      RECT  7577.5 40462.5 7642.5 40327.5 ;
      RECT  7767.5 40462.5 7832.5 40327.5 ;
      RECT  7767.5 40462.5 7832.5 40327.5 ;
      RECT  7577.5 40462.5 7642.5 40327.5 ;
      RECT  7197.5 41302.5 7262.5 41167.5 ;
      RECT  7387.5 41302.5 7452.5 41167.5 ;
      RECT  7387.5 41302.5 7452.5 41167.5 ;
      RECT  7197.5 41302.5 7262.5 41167.5 ;
      RECT  7387.5 41302.5 7452.5 41167.5 ;
      RECT  7577.5 41302.5 7642.5 41167.5 ;
      RECT  7577.5 41302.5 7642.5 41167.5 ;
      RECT  7387.5 41302.5 7452.5 41167.5 ;
      RECT  7577.5 41302.5 7642.5 41167.5 ;
      RECT  7767.5 41302.5 7832.5 41167.5 ;
      RECT  7767.5 41302.5 7832.5 41167.5 ;
      RECT  7577.5 41302.5 7642.5 41167.5 ;
      RECT  7937.5 40372.5 8002.5 40237.5 ;
      RECT  7937.5 41347.5 8002.5 41212.5 ;
      RECT  7772.5 41090.0 7637.5 41025.0 ;
      RECT  7582.5 40950.0 7447.5 40885.0 ;
      RECT  7392.5 40810.0 7257.5 40745.0 ;
      RECT  7387.5 40462.5 7452.5 40327.5 ;
      RECT  7767.5 40462.5 7832.5 40327.5 ;
      RECT  7767.5 41302.5 7832.5 41167.5 ;
      RECT  7767.5 40845.0 7832.5 40710.0 ;
      RECT  7257.5 40810.0 7392.5 40745.0 ;
      RECT  7447.5 40950.0 7582.5 40885.0 ;
      RECT  7637.5 41090.0 7772.5 41025.0 ;
      RECT  7767.5 40845.0 7832.5 40710.0 ;
      RECT  7130.0 40152.5 8140.0 40087.5 ;
      RECT  7130.0 41497.5 8140.0 41432.5 ;
      RECT  7197.5 41627.5 7262.5 41432.5 ;
      RECT  7197.5 42467.5 7262.5 42842.5 ;
      RECT  7577.5 42467.5 7642.5 42842.5 ;
      RECT  7937.5 42625.0 8002.5 42810.0 ;
      RECT  7937.5 41465.0 8002.5 41650.0 ;
      RECT  7197.5 42467.5 7262.5 42602.5 ;
      RECT  7387.5 42467.5 7452.5 42602.5 ;
      RECT  7387.5 42467.5 7452.5 42602.5 ;
      RECT  7197.5 42467.5 7262.5 42602.5 ;
      RECT  7387.5 42467.5 7452.5 42602.5 ;
      RECT  7577.5 42467.5 7642.5 42602.5 ;
      RECT  7577.5 42467.5 7642.5 42602.5 ;
      RECT  7387.5 42467.5 7452.5 42602.5 ;
      RECT  7577.5 42467.5 7642.5 42602.5 ;
      RECT  7767.5 42467.5 7832.5 42602.5 ;
      RECT  7767.5 42467.5 7832.5 42602.5 ;
      RECT  7577.5 42467.5 7642.5 42602.5 ;
      RECT  7197.5 41627.5 7262.5 41762.5 ;
      RECT  7387.5 41627.5 7452.5 41762.5 ;
      RECT  7387.5 41627.5 7452.5 41762.5 ;
      RECT  7197.5 41627.5 7262.5 41762.5 ;
      RECT  7387.5 41627.5 7452.5 41762.5 ;
      RECT  7577.5 41627.5 7642.5 41762.5 ;
      RECT  7577.5 41627.5 7642.5 41762.5 ;
      RECT  7387.5 41627.5 7452.5 41762.5 ;
      RECT  7577.5 41627.5 7642.5 41762.5 ;
      RECT  7767.5 41627.5 7832.5 41762.5 ;
      RECT  7767.5 41627.5 7832.5 41762.5 ;
      RECT  7577.5 41627.5 7642.5 41762.5 ;
      RECT  7937.5 42557.5 8002.5 42692.5 ;
      RECT  7937.5 41582.5 8002.5 41717.5 ;
      RECT  7772.5 41840.0 7637.5 41905.0 ;
      RECT  7582.5 41980.0 7447.5 42045.0 ;
      RECT  7392.5 42120.0 7257.5 42185.0 ;
      RECT  7387.5 42467.5 7452.5 42602.5 ;
      RECT  7767.5 42467.5 7832.5 42602.5 ;
      RECT  7767.5 41627.5 7832.5 41762.5 ;
      RECT  7767.5 42085.0 7832.5 42220.0 ;
      RECT  7257.5 42120.0 7392.5 42185.0 ;
      RECT  7447.5 41980.0 7582.5 42045.0 ;
      RECT  7637.5 41840.0 7772.5 41905.0 ;
      RECT  7767.5 42085.0 7832.5 42220.0 ;
      RECT  7130.0 42777.5 8140.0 42842.5 ;
      RECT  7130.0 41432.5 8140.0 41497.5 ;
      RECT  7197.5 43992.5 7262.5 44187.5 ;
      RECT  7197.5 43152.5 7262.5 42777.5 ;
      RECT  7577.5 43152.5 7642.5 42777.5 ;
      RECT  7937.5 42995.0 8002.5 42810.0 ;
      RECT  7937.5 44155.0 8002.5 43970.0 ;
      RECT  7197.5 43152.5 7262.5 43017.5 ;
      RECT  7387.5 43152.5 7452.5 43017.5 ;
      RECT  7387.5 43152.5 7452.5 43017.5 ;
      RECT  7197.5 43152.5 7262.5 43017.5 ;
      RECT  7387.5 43152.5 7452.5 43017.5 ;
      RECT  7577.5 43152.5 7642.5 43017.5 ;
      RECT  7577.5 43152.5 7642.5 43017.5 ;
      RECT  7387.5 43152.5 7452.5 43017.5 ;
      RECT  7577.5 43152.5 7642.5 43017.5 ;
      RECT  7767.5 43152.5 7832.5 43017.5 ;
      RECT  7767.5 43152.5 7832.5 43017.5 ;
      RECT  7577.5 43152.5 7642.5 43017.5 ;
      RECT  7197.5 43992.5 7262.5 43857.5 ;
      RECT  7387.5 43992.5 7452.5 43857.5 ;
      RECT  7387.5 43992.5 7452.5 43857.5 ;
      RECT  7197.5 43992.5 7262.5 43857.5 ;
      RECT  7387.5 43992.5 7452.5 43857.5 ;
      RECT  7577.5 43992.5 7642.5 43857.5 ;
      RECT  7577.5 43992.5 7642.5 43857.5 ;
      RECT  7387.5 43992.5 7452.5 43857.5 ;
      RECT  7577.5 43992.5 7642.5 43857.5 ;
      RECT  7767.5 43992.5 7832.5 43857.5 ;
      RECT  7767.5 43992.5 7832.5 43857.5 ;
      RECT  7577.5 43992.5 7642.5 43857.5 ;
      RECT  7937.5 43062.5 8002.5 42927.5 ;
      RECT  7937.5 44037.5 8002.5 43902.5 ;
      RECT  7772.5 43780.0 7637.5 43715.0 ;
      RECT  7582.5 43640.0 7447.5 43575.0 ;
      RECT  7392.5 43500.0 7257.5 43435.0 ;
      RECT  7387.5 43152.5 7452.5 43017.5 ;
      RECT  7767.5 43152.5 7832.5 43017.5 ;
      RECT  7767.5 43992.5 7832.5 43857.5 ;
      RECT  7767.5 43535.0 7832.5 43400.0 ;
      RECT  7257.5 43500.0 7392.5 43435.0 ;
      RECT  7447.5 43640.0 7582.5 43575.0 ;
      RECT  7637.5 43780.0 7772.5 43715.0 ;
      RECT  7767.5 43535.0 7832.5 43400.0 ;
      RECT  7130.0 42842.5 8140.0 42777.5 ;
      RECT  7130.0 44187.5 8140.0 44122.5 ;
      RECT  7197.5 44317.5 7262.5 44122.5 ;
      RECT  7197.5 45157.5 7262.5 45532.5 ;
      RECT  7577.5 45157.5 7642.5 45532.5 ;
      RECT  7937.5 45315.0 8002.5 45500.0 ;
      RECT  7937.5 44155.0 8002.5 44340.0 ;
      RECT  7197.5 45157.5 7262.5 45292.5 ;
      RECT  7387.5 45157.5 7452.5 45292.5 ;
      RECT  7387.5 45157.5 7452.5 45292.5 ;
      RECT  7197.5 45157.5 7262.5 45292.5 ;
      RECT  7387.5 45157.5 7452.5 45292.5 ;
      RECT  7577.5 45157.5 7642.5 45292.5 ;
      RECT  7577.5 45157.5 7642.5 45292.5 ;
      RECT  7387.5 45157.5 7452.5 45292.5 ;
      RECT  7577.5 45157.5 7642.5 45292.5 ;
      RECT  7767.5 45157.5 7832.5 45292.5 ;
      RECT  7767.5 45157.5 7832.5 45292.5 ;
      RECT  7577.5 45157.5 7642.5 45292.5 ;
      RECT  7197.5 44317.5 7262.5 44452.5 ;
      RECT  7387.5 44317.5 7452.5 44452.5 ;
      RECT  7387.5 44317.5 7452.5 44452.5 ;
      RECT  7197.5 44317.5 7262.5 44452.5 ;
      RECT  7387.5 44317.5 7452.5 44452.5 ;
      RECT  7577.5 44317.5 7642.5 44452.5 ;
      RECT  7577.5 44317.5 7642.5 44452.5 ;
      RECT  7387.5 44317.5 7452.5 44452.5 ;
      RECT  7577.5 44317.5 7642.5 44452.5 ;
      RECT  7767.5 44317.5 7832.5 44452.5 ;
      RECT  7767.5 44317.5 7832.5 44452.5 ;
      RECT  7577.5 44317.5 7642.5 44452.5 ;
      RECT  7937.5 45247.5 8002.5 45382.5 ;
      RECT  7937.5 44272.5 8002.5 44407.5 ;
      RECT  7772.5 44530.0 7637.5 44595.0 ;
      RECT  7582.5 44670.0 7447.5 44735.0 ;
      RECT  7392.5 44810.0 7257.5 44875.0 ;
      RECT  7387.5 45157.5 7452.5 45292.5 ;
      RECT  7767.5 45157.5 7832.5 45292.5 ;
      RECT  7767.5 44317.5 7832.5 44452.5 ;
      RECT  7767.5 44775.0 7832.5 44910.0 ;
      RECT  7257.5 44810.0 7392.5 44875.0 ;
      RECT  7447.5 44670.0 7582.5 44735.0 ;
      RECT  7637.5 44530.0 7772.5 44595.0 ;
      RECT  7767.5 44775.0 7832.5 44910.0 ;
      RECT  7130.0 45467.5 8140.0 45532.5 ;
      RECT  7130.0 44122.5 8140.0 44187.5 ;
      RECT  7197.5 46682.5 7262.5 46877.5 ;
      RECT  7197.5 45842.5 7262.5 45467.5 ;
      RECT  7577.5 45842.5 7642.5 45467.5 ;
      RECT  7937.5 45685.0 8002.5 45500.0 ;
      RECT  7937.5 46845.0 8002.5 46660.0 ;
      RECT  7197.5 45842.5 7262.5 45707.5 ;
      RECT  7387.5 45842.5 7452.5 45707.5 ;
      RECT  7387.5 45842.5 7452.5 45707.5 ;
      RECT  7197.5 45842.5 7262.5 45707.5 ;
      RECT  7387.5 45842.5 7452.5 45707.5 ;
      RECT  7577.5 45842.5 7642.5 45707.5 ;
      RECT  7577.5 45842.5 7642.5 45707.5 ;
      RECT  7387.5 45842.5 7452.5 45707.5 ;
      RECT  7577.5 45842.5 7642.5 45707.5 ;
      RECT  7767.5 45842.5 7832.5 45707.5 ;
      RECT  7767.5 45842.5 7832.5 45707.5 ;
      RECT  7577.5 45842.5 7642.5 45707.5 ;
      RECT  7197.5 46682.5 7262.5 46547.5 ;
      RECT  7387.5 46682.5 7452.5 46547.5 ;
      RECT  7387.5 46682.5 7452.5 46547.5 ;
      RECT  7197.5 46682.5 7262.5 46547.5 ;
      RECT  7387.5 46682.5 7452.5 46547.5 ;
      RECT  7577.5 46682.5 7642.5 46547.5 ;
      RECT  7577.5 46682.5 7642.5 46547.5 ;
      RECT  7387.5 46682.5 7452.5 46547.5 ;
      RECT  7577.5 46682.5 7642.5 46547.5 ;
      RECT  7767.5 46682.5 7832.5 46547.5 ;
      RECT  7767.5 46682.5 7832.5 46547.5 ;
      RECT  7577.5 46682.5 7642.5 46547.5 ;
      RECT  7937.5 45752.5 8002.5 45617.5 ;
      RECT  7937.5 46727.5 8002.5 46592.5 ;
      RECT  7772.5 46470.0 7637.5 46405.0 ;
      RECT  7582.5 46330.0 7447.5 46265.0 ;
      RECT  7392.5 46190.0 7257.5 46125.0 ;
      RECT  7387.5 45842.5 7452.5 45707.5 ;
      RECT  7767.5 45842.5 7832.5 45707.5 ;
      RECT  7767.5 46682.5 7832.5 46547.5 ;
      RECT  7767.5 46225.0 7832.5 46090.0 ;
      RECT  7257.5 46190.0 7392.5 46125.0 ;
      RECT  7447.5 46330.0 7582.5 46265.0 ;
      RECT  7637.5 46470.0 7772.5 46405.0 ;
      RECT  7767.5 46225.0 7832.5 46090.0 ;
      RECT  7130.0 45532.5 8140.0 45467.5 ;
      RECT  7130.0 46877.5 8140.0 46812.5 ;
      RECT  7197.5 47007.5 7262.5 46812.5 ;
      RECT  7197.5 47847.5 7262.5 48222.5 ;
      RECT  7577.5 47847.5 7642.5 48222.5 ;
      RECT  7937.5 48005.0 8002.5 48190.0 ;
      RECT  7937.5 46845.0 8002.5 47030.0 ;
      RECT  7197.5 47847.5 7262.5 47982.5 ;
      RECT  7387.5 47847.5 7452.5 47982.5 ;
      RECT  7387.5 47847.5 7452.5 47982.5 ;
      RECT  7197.5 47847.5 7262.5 47982.5 ;
      RECT  7387.5 47847.5 7452.5 47982.5 ;
      RECT  7577.5 47847.5 7642.5 47982.5 ;
      RECT  7577.5 47847.5 7642.5 47982.5 ;
      RECT  7387.5 47847.5 7452.5 47982.5 ;
      RECT  7577.5 47847.5 7642.5 47982.5 ;
      RECT  7767.5 47847.5 7832.5 47982.5 ;
      RECT  7767.5 47847.5 7832.5 47982.5 ;
      RECT  7577.5 47847.5 7642.5 47982.5 ;
      RECT  7197.5 47007.5 7262.5 47142.5 ;
      RECT  7387.5 47007.5 7452.5 47142.5 ;
      RECT  7387.5 47007.5 7452.5 47142.5 ;
      RECT  7197.5 47007.5 7262.5 47142.5 ;
      RECT  7387.5 47007.5 7452.5 47142.5 ;
      RECT  7577.5 47007.5 7642.5 47142.5 ;
      RECT  7577.5 47007.5 7642.5 47142.5 ;
      RECT  7387.5 47007.5 7452.5 47142.5 ;
      RECT  7577.5 47007.5 7642.5 47142.5 ;
      RECT  7767.5 47007.5 7832.5 47142.5 ;
      RECT  7767.5 47007.5 7832.5 47142.5 ;
      RECT  7577.5 47007.5 7642.5 47142.5 ;
      RECT  7937.5 47937.5 8002.5 48072.5 ;
      RECT  7937.5 46962.5 8002.5 47097.5 ;
      RECT  7772.5 47220.0 7637.5 47285.0 ;
      RECT  7582.5 47360.0 7447.5 47425.0 ;
      RECT  7392.5 47500.0 7257.5 47565.0 ;
      RECT  7387.5 47847.5 7452.5 47982.5 ;
      RECT  7767.5 47847.5 7832.5 47982.5 ;
      RECT  7767.5 47007.5 7832.5 47142.5 ;
      RECT  7767.5 47465.0 7832.5 47600.0 ;
      RECT  7257.5 47500.0 7392.5 47565.0 ;
      RECT  7447.5 47360.0 7582.5 47425.0 ;
      RECT  7637.5 47220.0 7772.5 47285.0 ;
      RECT  7767.5 47465.0 7832.5 47600.0 ;
      RECT  7130.0 48157.5 8140.0 48222.5 ;
      RECT  7130.0 46812.5 8140.0 46877.5 ;
      RECT  7197.5 49372.5 7262.5 49567.5 ;
      RECT  7197.5 48532.5 7262.5 48157.5 ;
      RECT  7577.5 48532.5 7642.5 48157.5 ;
      RECT  7937.5 48375.0 8002.5 48190.0 ;
      RECT  7937.5 49535.0 8002.5 49350.0 ;
      RECT  7197.5 48532.5 7262.5 48397.5 ;
      RECT  7387.5 48532.5 7452.5 48397.5 ;
      RECT  7387.5 48532.5 7452.5 48397.5 ;
      RECT  7197.5 48532.5 7262.5 48397.5 ;
      RECT  7387.5 48532.5 7452.5 48397.5 ;
      RECT  7577.5 48532.5 7642.5 48397.5 ;
      RECT  7577.5 48532.5 7642.5 48397.5 ;
      RECT  7387.5 48532.5 7452.5 48397.5 ;
      RECT  7577.5 48532.5 7642.5 48397.5 ;
      RECT  7767.5 48532.5 7832.5 48397.5 ;
      RECT  7767.5 48532.5 7832.5 48397.5 ;
      RECT  7577.5 48532.5 7642.5 48397.5 ;
      RECT  7197.5 49372.5 7262.5 49237.5 ;
      RECT  7387.5 49372.5 7452.5 49237.5 ;
      RECT  7387.5 49372.5 7452.5 49237.5 ;
      RECT  7197.5 49372.5 7262.5 49237.5 ;
      RECT  7387.5 49372.5 7452.5 49237.5 ;
      RECT  7577.5 49372.5 7642.5 49237.5 ;
      RECT  7577.5 49372.5 7642.5 49237.5 ;
      RECT  7387.5 49372.5 7452.5 49237.5 ;
      RECT  7577.5 49372.5 7642.5 49237.5 ;
      RECT  7767.5 49372.5 7832.5 49237.5 ;
      RECT  7767.5 49372.5 7832.5 49237.5 ;
      RECT  7577.5 49372.5 7642.5 49237.5 ;
      RECT  7937.5 48442.5 8002.5 48307.5 ;
      RECT  7937.5 49417.5 8002.5 49282.5 ;
      RECT  7772.5 49160.0 7637.5 49095.0 ;
      RECT  7582.5 49020.0 7447.5 48955.0 ;
      RECT  7392.5 48880.0 7257.5 48815.0 ;
      RECT  7387.5 48532.5 7452.5 48397.5 ;
      RECT  7767.5 48532.5 7832.5 48397.5 ;
      RECT  7767.5 49372.5 7832.5 49237.5 ;
      RECT  7767.5 48915.0 7832.5 48780.0 ;
      RECT  7257.5 48880.0 7392.5 48815.0 ;
      RECT  7447.5 49020.0 7582.5 48955.0 ;
      RECT  7637.5 49160.0 7772.5 49095.0 ;
      RECT  7767.5 48915.0 7832.5 48780.0 ;
      RECT  7130.0 48222.5 8140.0 48157.5 ;
      RECT  7130.0 49567.5 8140.0 49502.5 ;
      RECT  7197.5 49697.5 7262.5 49502.5 ;
      RECT  7197.5 50537.5 7262.5 50912.5 ;
      RECT  7577.5 50537.5 7642.5 50912.5 ;
      RECT  7937.5 50695.0 8002.5 50880.0 ;
      RECT  7937.5 49535.0 8002.5 49720.0 ;
      RECT  7197.5 50537.5 7262.5 50672.5 ;
      RECT  7387.5 50537.5 7452.5 50672.5 ;
      RECT  7387.5 50537.5 7452.5 50672.5 ;
      RECT  7197.5 50537.5 7262.5 50672.5 ;
      RECT  7387.5 50537.5 7452.5 50672.5 ;
      RECT  7577.5 50537.5 7642.5 50672.5 ;
      RECT  7577.5 50537.5 7642.5 50672.5 ;
      RECT  7387.5 50537.5 7452.5 50672.5 ;
      RECT  7577.5 50537.5 7642.5 50672.5 ;
      RECT  7767.5 50537.5 7832.5 50672.5 ;
      RECT  7767.5 50537.5 7832.5 50672.5 ;
      RECT  7577.5 50537.5 7642.5 50672.5 ;
      RECT  7197.5 49697.5 7262.5 49832.5 ;
      RECT  7387.5 49697.5 7452.5 49832.5 ;
      RECT  7387.5 49697.5 7452.5 49832.5 ;
      RECT  7197.5 49697.5 7262.5 49832.5 ;
      RECT  7387.5 49697.5 7452.5 49832.5 ;
      RECT  7577.5 49697.5 7642.5 49832.5 ;
      RECT  7577.5 49697.5 7642.5 49832.5 ;
      RECT  7387.5 49697.5 7452.5 49832.5 ;
      RECT  7577.5 49697.5 7642.5 49832.5 ;
      RECT  7767.5 49697.5 7832.5 49832.5 ;
      RECT  7767.5 49697.5 7832.5 49832.5 ;
      RECT  7577.5 49697.5 7642.5 49832.5 ;
      RECT  7937.5 50627.5 8002.5 50762.5 ;
      RECT  7937.5 49652.5 8002.5 49787.5 ;
      RECT  7772.5 49910.0 7637.5 49975.0 ;
      RECT  7582.5 50050.0 7447.5 50115.0 ;
      RECT  7392.5 50190.0 7257.5 50255.0 ;
      RECT  7387.5 50537.5 7452.5 50672.5 ;
      RECT  7767.5 50537.5 7832.5 50672.5 ;
      RECT  7767.5 49697.5 7832.5 49832.5 ;
      RECT  7767.5 50155.0 7832.5 50290.0 ;
      RECT  7257.5 50190.0 7392.5 50255.0 ;
      RECT  7447.5 50050.0 7582.5 50115.0 ;
      RECT  7637.5 49910.0 7772.5 49975.0 ;
      RECT  7767.5 50155.0 7832.5 50290.0 ;
      RECT  7130.0 50847.5 8140.0 50912.5 ;
      RECT  7130.0 49502.5 8140.0 49567.5 ;
      RECT  7197.5 52062.5 7262.5 52257.5 ;
      RECT  7197.5 51222.5 7262.5 50847.5 ;
      RECT  7577.5 51222.5 7642.5 50847.5 ;
      RECT  7937.5 51065.0 8002.5 50880.0 ;
      RECT  7937.5 52225.0 8002.5 52040.0 ;
      RECT  7197.5 51222.5 7262.5 51087.5 ;
      RECT  7387.5 51222.5 7452.5 51087.5 ;
      RECT  7387.5 51222.5 7452.5 51087.5 ;
      RECT  7197.5 51222.5 7262.5 51087.5 ;
      RECT  7387.5 51222.5 7452.5 51087.5 ;
      RECT  7577.5 51222.5 7642.5 51087.5 ;
      RECT  7577.5 51222.5 7642.5 51087.5 ;
      RECT  7387.5 51222.5 7452.5 51087.5 ;
      RECT  7577.5 51222.5 7642.5 51087.5 ;
      RECT  7767.5 51222.5 7832.5 51087.5 ;
      RECT  7767.5 51222.5 7832.5 51087.5 ;
      RECT  7577.5 51222.5 7642.5 51087.5 ;
      RECT  7197.5 52062.5 7262.5 51927.5 ;
      RECT  7387.5 52062.5 7452.5 51927.5 ;
      RECT  7387.5 52062.5 7452.5 51927.5 ;
      RECT  7197.5 52062.5 7262.5 51927.5 ;
      RECT  7387.5 52062.5 7452.5 51927.5 ;
      RECT  7577.5 52062.5 7642.5 51927.5 ;
      RECT  7577.5 52062.5 7642.5 51927.5 ;
      RECT  7387.5 52062.5 7452.5 51927.5 ;
      RECT  7577.5 52062.5 7642.5 51927.5 ;
      RECT  7767.5 52062.5 7832.5 51927.5 ;
      RECT  7767.5 52062.5 7832.5 51927.5 ;
      RECT  7577.5 52062.5 7642.5 51927.5 ;
      RECT  7937.5 51132.5 8002.5 50997.5 ;
      RECT  7937.5 52107.5 8002.5 51972.5 ;
      RECT  7772.5 51850.0 7637.5 51785.0 ;
      RECT  7582.5 51710.0 7447.5 51645.0 ;
      RECT  7392.5 51570.0 7257.5 51505.0 ;
      RECT  7387.5 51222.5 7452.5 51087.5 ;
      RECT  7767.5 51222.5 7832.5 51087.5 ;
      RECT  7767.5 52062.5 7832.5 51927.5 ;
      RECT  7767.5 51605.0 7832.5 51470.0 ;
      RECT  7257.5 51570.0 7392.5 51505.0 ;
      RECT  7447.5 51710.0 7582.5 51645.0 ;
      RECT  7637.5 51850.0 7772.5 51785.0 ;
      RECT  7767.5 51605.0 7832.5 51470.0 ;
      RECT  7130.0 50912.5 8140.0 50847.5 ;
      RECT  7130.0 52257.5 8140.0 52192.5 ;
      RECT  7197.5 52387.5 7262.5 52192.5 ;
      RECT  7197.5 53227.5 7262.5 53602.5 ;
      RECT  7577.5 53227.5 7642.5 53602.5 ;
      RECT  7937.5 53385.0 8002.5 53570.0 ;
      RECT  7937.5 52225.0 8002.5 52410.0 ;
      RECT  7197.5 53227.5 7262.5 53362.5 ;
      RECT  7387.5 53227.5 7452.5 53362.5 ;
      RECT  7387.5 53227.5 7452.5 53362.5 ;
      RECT  7197.5 53227.5 7262.5 53362.5 ;
      RECT  7387.5 53227.5 7452.5 53362.5 ;
      RECT  7577.5 53227.5 7642.5 53362.5 ;
      RECT  7577.5 53227.5 7642.5 53362.5 ;
      RECT  7387.5 53227.5 7452.5 53362.5 ;
      RECT  7577.5 53227.5 7642.5 53362.5 ;
      RECT  7767.5 53227.5 7832.5 53362.5 ;
      RECT  7767.5 53227.5 7832.5 53362.5 ;
      RECT  7577.5 53227.5 7642.5 53362.5 ;
      RECT  7197.5 52387.5 7262.5 52522.5 ;
      RECT  7387.5 52387.5 7452.5 52522.5 ;
      RECT  7387.5 52387.5 7452.5 52522.5 ;
      RECT  7197.5 52387.5 7262.5 52522.5 ;
      RECT  7387.5 52387.5 7452.5 52522.5 ;
      RECT  7577.5 52387.5 7642.5 52522.5 ;
      RECT  7577.5 52387.5 7642.5 52522.5 ;
      RECT  7387.5 52387.5 7452.5 52522.5 ;
      RECT  7577.5 52387.5 7642.5 52522.5 ;
      RECT  7767.5 52387.5 7832.5 52522.5 ;
      RECT  7767.5 52387.5 7832.5 52522.5 ;
      RECT  7577.5 52387.5 7642.5 52522.5 ;
      RECT  7937.5 53317.5 8002.5 53452.5 ;
      RECT  7937.5 52342.5 8002.5 52477.5 ;
      RECT  7772.5 52600.0 7637.5 52665.0 ;
      RECT  7582.5 52740.0 7447.5 52805.0 ;
      RECT  7392.5 52880.0 7257.5 52945.0 ;
      RECT  7387.5 53227.5 7452.5 53362.5 ;
      RECT  7767.5 53227.5 7832.5 53362.5 ;
      RECT  7767.5 52387.5 7832.5 52522.5 ;
      RECT  7767.5 52845.0 7832.5 52980.0 ;
      RECT  7257.5 52880.0 7392.5 52945.0 ;
      RECT  7447.5 52740.0 7582.5 52805.0 ;
      RECT  7637.5 52600.0 7772.5 52665.0 ;
      RECT  7767.5 52845.0 7832.5 52980.0 ;
      RECT  7130.0 53537.5 8140.0 53602.5 ;
      RECT  7130.0 52192.5 8140.0 52257.5 ;
      RECT  7197.5 54752.5 7262.5 54947.5 ;
      RECT  7197.5 53912.5 7262.5 53537.5 ;
      RECT  7577.5 53912.5 7642.5 53537.5 ;
      RECT  7937.5 53755.0 8002.5 53570.0 ;
      RECT  7937.5 54915.0 8002.5 54730.0 ;
      RECT  7197.5 53912.5 7262.5 53777.5 ;
      RECT  7387.5 53912.5 7452.5 53777.5 ;
      RECT  7387.5 53912.5 7452.5 53777.5 ;
      RECT  7197.5 53912.5 7262.5 53777.5 ;
      RECT  7387.5 53912.5 7452.5 53777.5 ;
      RECT  7577.5 53912.5 7642.5 53777.5 ;
      RECT  7577.5 53912.5 7642.5 53777.5 ;
      RECT  7387.5 53912.5 7452.5 53777.5 ;
      RECT  7577.5 53912.5 7642.5 53777.5 ;
      RECT  7767.5 53912.5 7832.5 53777.5 ;
      RECT  7767.5 53912.5 7832.5 53777.5 ;
      RECT  7577.5 53912.5 7642.5 53777.5 ;
      RECT  7197.5 54752.5 7262.5 54617.5 ;
      RECT  7387.5 54752.5 7452.5 54617.5 ;
      RECT  7387.5 54752.5 7452.5 54617.5 ;
      RECT  7197.5 54752.5 7262.5 54617.5 ;
      RECT  7387.5 54752.5 7452.5 54617.5 ;
      RECT  7577.5 54752.5 7642.5 54617.5 ;
      RECT  7577.5 54752.5 7642.5 54617.5 ;
      RECT  7387.5 54752.5 7452.5 54617.5 ;
      RECT  7577.5 54752.5 7642.5 54617.5 ;
      RECT  7767.5 54752.5 7832.5 54617.5 ;
      RECT  7767.5 54752.5 7832.5 54617.5 ;
      RECT  7577.5 54752.5 7642.5 54617.5 ;
      RECT  7937.5 53822.5 8002.5 53687.5 ;
      RECT  7937.5 54797.5 8002.5 54662.5 ;
      RECT  7772.5 54540.0 7637.5 54475.0 ;
      RECT  7582.5 54400.0 7447.5 54335.0 ;
      RECT  7392.5 54260.0 7257.5 54195.0 ;
      RECT  7387.5 53912.5 7452.5 53777.5 ;
      RECT  7767.5 53912.5 7832.5 53777.5 ;
      RECT  7767.5 54752.5 7832.5 54617.5 ;
      RECT  7767.5 54295.0 7832.5 54160.0 ;
      RECT  7257.5 54260.0 7392.5 54195.0 ;
      RECT  7447.5 54400.0 7582.5 54335.0 ;
      RECT  7637.5 54540.0 7772.5 54475.0 ;
      RECT  7767.5 54295.0 7832.5 54160.0 ;
      RECT  7130.0 53602.5 8140.0 53537.5 ;
      RECT  7130.0 54947.5 8140.0 54882.5 ;
      RECT  7197.5 55077.5 7262.5 54882.5 ;
      RECT  7197.5 55917.5 7262.5 56292.5 ;
      RECT  7577.5 55917.5 7642.5 56292.5 ;
      RECT  7937.5 56075.0 8002.5 56260.0 ;
      RECT  7937.5 54915.0 8002.5 55100.0 ;
      RECT  7197.5 55917.5 7262.5 56052.5 ;
      RECT  7387.5 55917.5 7452.5 56052.5 ;
      RECT  7387.5 55917.5 7452.5 56052.5 ;
      RECT  7197.5 55917.5 7262.5 56052.5 ;
      RECT  7387.5 55917.5 7452.5 56052.5 ;
      RECT  7577.5 55917.5 7642.5 56052.5 ;
      RECT  7577.5 55917.5 7642.5 56052.5 ;
      RECT  7387.5 55917.5 7452.5 56052.5 ;
      RECT  7577.5 55917.5 7642.5 56052.5 ;
      RECT  7767.5 55917.5 7832.5 56052.5 ;
      RECT  7767.5 55917.5 7832.5 56052.5 ;
      RECT  7577.5 55917.5 7642.5 56052.5 ;
      RECT  7197.5 55077.5 7262.5 55212.5 ;
      RECT  7387.5 55077.5 7452.5 55212.5 ;
      RECT  7387.5 55077.5 7452.5 55212.5 ;
      RECT  7197.5 55077.5 7262.5 55212.5 ;
      RECT  7387.5 55077.5 7452.5 55212.5 ;
      RECT  7577.5 55077.5 7642.5 55212.5 ;
      RECT  7577.5 55077.5 7642.5 55212.5 ;
      RECT  7387.5 55077.5 7452.5 55212.5 ;
      RECT  7577.5 55077.5 7642.5 55212.5 ;
      RECT  7767.5 55077.5 7832.5 55212.5 ;
      RECT  7767.5 55077.5 7832.5 55212.5 ;
      RECT  7577.5 55077.5 7642.5 55212.5 ;
      RECT  7937.5 56007.5 8002.5 56142.5 ;
      RECT  7937.5 55032.5 8002.5 55167.5 ;
      RECT  7772.5 55290.0 7637.5 55355.0 ;
      RECT  7582.5 55430.0 7447.5 55495.0 ;
      RECT  7392.5 55570.0 7257.5 55635.0 ;
      RECT  7387.5 55917.5 7452.5 56052.5 ;
      RECT  7767.5 55917.5 7832.5 56052.5 ;
      RECT  7767.5 55077.5 7832.5 55212.5 ;
      RECT  7767.5 55535.0 7832.5 55670.0 ;
      RECT  7257.5 55570.0 7392.5 55635.0 ;
      RECT  7447.5 55430.0 7582.5 55495.0 ;
      RECT  7637.5 55290.0 7772.5 55355.0 ;
      RECT  7767.5 55535.0 7832.5 55670.0 ;
      RECT  7130.0 56227.5 8140.0 56292.5 ;
      RECT  7130.0 54882.5 8140.0 54947.5 ;
      RECT  7197.5 57442.5 7262.5 57637.5 ;
      RECT  7197.5 56602.5 7262.5 56227.5 ;
      RECT  7577.5 56602.5 7642.5 56227.5 ;
      RECT  7937.5 56445.0 8002.5 56260.0 ;
      RECT  7937.5 57605.0 8002.5 57420.0 ;
      RECT  7197.5 56602.5 7262.5 56467.5 ;
      RECT  7387.5 56602.5 7452.5 56467.5 ;
      RECT  7387.5 56602.5 7452.5 56467.5 ;
      RECT  7197.5 56602.5 7262.5 56467.5 ;
      RECT  7387.5 56602.5 7452.5 56467.5 ;
      RECT  7577.5 56602.5 7642.5 56467.5 ;
      RECT  7577.5 56602.5 7642.5 56467.5 ;
      RECT  7387.5 56602.5 7452.5 56467.5 ;
      RECT  7577.5 56602.5 7642.5 56467.5 ;
      RECT  7767.5 56602.5 7832.5 56467.5 ;
      RECT  7767.5 56602.5 7832.5 56467.5 ;
      RECT  7577.5 56602.5 7642.5 56467.5 ;
      RECT  7197.5 57442.5 7262.5 57307.5 ;
      RECT  7387.5 57442.5 7452.5 57307.5 ;
      RECT  7387.5 57442.5 7452.5 57307.5 ;
      RECT  7197.5 57442.5 7262.5 57307.5 ;
      RECT  7387.5 57442.5 7452.5 57307.5 ;
      RECT  7577.5 57442.5 7642.5 57307.5 ;
      RECT  7577.5 57442.5 7642.5 57307.5 ;
      RECT  7387.5 57442.5 7452.5 57307.5 ;
      RECT  7577.5 57442.5 7642.5 57307.5 ;
      RECT  7767.5 57442.5 7832.5 57307.5 ;
      RECT  7767.5 57442.5 7832.5 57307.5 ;
      RECT  7577.5 57442.5 7642.5 57307.5 ;
      RECT  7937.5 56512.5 8002.5 56377.5 ;
      RECT  7937.5 57487.5 8002.5 57352.5 ;
      RECT  7772.5 57230.0 7637.5 57165.0 ;
      RECT  7582.5 57090.0 7447.5 57025.0 ;
      RECT  7392.5 56950.0 7257.5 56885.0 ;
      RECT  7387.5 56602.5 7452.5 56467.5 ;
      RECT  7767.5 56602.5 7832.5 56467.5 ;
      RECT  7767.5 57442.5 7832.5 57307.5 ;
      RECT  7767.5 56985.0 7832.5 56850.0 ;
      RECT  7257.5 56950.0 7392.5 56885.0 ;
      RECT  7447.5 57090.0 7582.5 57025.0 ;
      RECT  7637.5 57230.0 7772.5 57165.0 ;
      RECT  7767.5 56985.0 7832.5 56850.0 ;
      RECT  7130.0 56292.5 8140.0 56227.5 ;
      RECT  7130.0 57637.5 8140.0 57572.5 ;
      RECT  7197.5 57767.5 7262.5 57572.5 ;
      RECT  7197.5 58607.5 7262.5 58982.5 ;
      RECT  7577.5 58607.5 7642.5 58982.5 ;
      RECT  7937.5 58765.0 8002.5 58950.0 ;
      RECT  7937.5 57605.0 8002.5 57790.0 ;
      RECT  7197.5 58607.5 7262.5 58742.5 ;
      RECT  7387.5 58607.5 7452.5 58742.5 ;
      RECT  7387.5 58607.5 7452.5 58742.5 ;
      RECT  7197.5 58607.5 7262.5 58742.5 ;
      RECT  7387.5 58607.5 7452.5 58742.5 ;
      RECT  7577.5 58607.5 7642.5 58742.5 ;
      RECT  7577.5 58607.5 7642.5 58742.5 ;
      RECT  7387.5 58607.5 7452.5 58742.5 ;
      RECT  7577.5 58607.5 7642.5 58742.5 ;
      RECT  7767.5 58607.5 7832.5 58742.5 ;
      RECT  7767.5 58607.5 7832.5 58742.5 ;
      RECT  7577.5 58607.5 7642.5 58742.5 ;
      RECT  7197.5 57767.5 7262.5 57902.5 ;
      RECT  7387.5 57767.5 7452.5 57902.5 ;
      RECT  7387.5 57767.5 7452.5 57902.5 ;
      RECT  7197.5 57767.5 7262.5 57902.5 ;
      RECT  7387.5 57767.5 7452.5 57902.5 ;
      RECT  7577.5 57767.5 7642.5 57902.5 ;
      RECT  7577.5 57767.5 7642.5 57902.5 ;
      RECT  7387.5 57767.5 7452.5 57902.5 ;
      RECT  7577.5 57767.5 7642.5 57902.5 ;
      RECT  7767.5 57767.5 7832.5 57902.5 ;
      RECT  7767.5 57767.5 7832.5 57902.5 ;
      RECT  7577.5 57767.5 7642.5 57902.5 ;
      RECT  7937.5 58697.5 8002.5 58832.5 ;
      RECT  7937.5 57722.5 8002.5 57857.5 ;
      RECT  7772.5 57980.0 7637.5 58045.0 ;
      RECT  7582.5 58120.0 7447.5 58185.0 ;
      RECT  7392.5 58260.0 7257.5 58325.0 ;
      RECT  7387.5 58607.5 7452.5 58742.5 ;
      RECT  7767.5 58607.5 7832.5 58742.5 ;
      RECT  7767.5 57767.5 7832.5 57902.5 ;
      RECT  7767.5 58225.0 7832.5 58360.0 ;
      RECT  7257.5 58260.0 7392.5 58325.0 ;
      RECT  7447.5 58120.0 7582.5 58185.0 ;
      RECT  7637.5 57980.0 7772.5 58045.0 ;
      RECT  7767.5 58225.0 7832.5 58360.0 ;
      RECT  7130.0 58917.5 8140.0 58982.5 ;
      RECT  7130.0 57572.5 8140.0 57637.5 ;
      RECT  7197.5 60132.5 7262.5 60327.5 ;
      RECT  7197.5 59292.5 7262.5 58917.5 ;
      RECT  7577.5 59292.5 7642.5 58917.5 ;
      RECT  7937.5 59135.0 8002.5 58950.0 ;
      RECT  7937.5 60295.0 8002.5 60110.0 ;
      RECT  7197.5 59292.5 7262.5 59157.5 ;
      RECT  7387.5 59292.5 7452.5 59157.5 ;
      RECT  7387.5 59292.5 7452.5 59157.5 ;
      RECT  7197.5 59292.5 7262.5 59157.5 ;
      RECT  7387.5 59292.5 7452.5 59157.5 ;
      RECT  7577.5 59292.5 7642.5 59157.5 ;
      RECT  7577.5 59292.5 7642.5 59157.5 ;
      RECT  7387.5 59292.5 7452.5 59157.5 ;
      RECT  7577.5 59292.5 7642.5 59157.5 ;
      RECT  7767.5 59292.5 7832.5 59157.5 ;
      RECT  7767.5 59292.5 7832.5 59157.5 ;
      RECT  7577.5 59292.5 7642.5 59157.5 ;
      RECT  7197.5 60132.5 7262.5 59997.5 ;
      RECT  7387.5 60132.5 7452.5 59997.5 ;
      RECT  7387.5 60132.5 7452.5 59997.5 ;
      RECT  7197.5 60132.5 7262.5 59997.5 ;
      RECT  7387.5 60132.5 7452.5 59997.5 ;
      RECT  7577.5 60132.5 7642.5 59997.5 ;
      RECT  7577.5 60132.5 7642.5 59997.5 ;
      RECT  7387.5 60132.5 7452.5 59997.5 ;
      RECT  7577.5 60132.5 7642.5 59997.5 ;
      RECT  7767.5 60132.5 7832.5 59997.5 ;
      RECT  7767.5 60132.5 7832.5 59997.5 ;
      RECT  7577.5 60132.5 7642.5 59997.5 ;
      RECT  7937.5 59202.5 8002.5 59067.5 ;
      RECT  7937.5 60177.5 8002.5 60042.5 ;
      RECT  7772.5 59920.0 7637.5 59855.0 ;
      RECT  7582.5 59780.0 7447.5 59715.0 ;
      RECT  7392.5 59640.0 7257.5 59575.0 ;
      RECT  7387.5 59292.5 7452.5 59157.5 ;
      RECT  7767.5 59292.5 7832.5 59157.5 ;
      RECT  7767.5 60132.5 7832.5 59997.5 ;
      RECT  7767.5 59675.0 7832.5 59540.0 ;
      RECT  7257.5 59640.0 7392.5 59575.0 ;
      RECT  7447.5 59780.0 7582.5 59715.0 ;
      RECT  7637.5 59920.0 7772.5 59855.0 ;
      RECT  7767.5 59675.0 7832.5 59540.0 ;
      RECT  7130.0 58982.5 8140.0 58917.5 ;
      RECT  7130.0 60327.5 8140.0 60262.5 ;
      RECT  7197.5 60457.5 7262.5 60262.5 ;
      RECT  7197.5 61297.5 7262.5 61672.5 ;
      RECT  7577.5 61297.5 7642.5 61672.5 ;
      RECT  7937.5 61455.0 8002.5 61640.0 ;
      RECT  7937.5 60295.0 8002.5 60480.0 ;
      RECT  7197.5 61297.5 7262.5 61432.5 ;
      RECT  7387.5 61297.5 7452.5 61432.5 ;
      RECT  7387.5 61297.5 7452.5 61432.5 ;
      RECT  7197.5 61297.5 7262.5 61432.5 ;
      RECT  7387.5 61297.5 7452.5 61432.5 ;
      RECT  7577.5 61297.5 7642.5 61432.5 ;
      RECT  7577.5 61297.5 7642.5 61432.5 ;
      RECT  7387.5 61297.5 7452.5 61432.5 ;
      RECT  7577.5 61297.5 7642.5 61432.5 ;
      RECT  7767.5 61297.5 7832.5 61432.5 ;
      RECT  7767.5 61297.5 7832.5 61432.5 ;
      RECT  7577.5 61297.5 7642.5 61432.5 ;
      RECT  7197.5 60457.5 7262.5 60592.5 ;
      RECT  7387.5 60457.5 7452.5 60592.5 ;
      RECT  7387.5 60457.5 7452.5 60592.5 ;
      RECT  7197.5 60457.5 7262.5 60592.5 ;
      RECT  7387.5 60457.5 7452.5 60592.5 ;
      RECT  7577.5 60457.5 7642.5 60592.5 ;
      RECT  7577.5 60457.5 7642.5 60592.5 ;
      RECT  7387.5 60457.5 7452.5 60592.5 ;
      RECT  7577.5 60457.5 7642.5 60592.5 ;
      RECT  7767.5 60457.5 7832.5 60592.5 ;
      RECT  7767.5 60457.5 7832.5 60592.5 ;
      RECT  7577.5 60457.5 7642.5 60592.5 ;
      RECT  7937.5 61387.5 8002.5 61522.5 ;
      RECT  7937.5 60412.5 8002.5 60547.5 ;
      RECT  7772.5 60670.0 7637.5 60735.0 ;
      RECT  7582.5 60810.0 7447.5 60875.0 ;
      RECT  7392.5 60950.0 7257.5 61015.0 ;
      RECT  7387.5 61297.5 7452.5 61432.5 ;
      RECT  7767.5 61297.5 7832.5 61432.5 ;
      RECT  7767.5 60457.5 7832.5 60592.5 ;
      RECT  7767.5 60915.0 7832.5 61050.0 ;
      RECT  7257.5 60950.0 7392.5 61015.0 ;
      RECT  7447.5 60810.0 7582.5 60875.0 ;
      RECT  7637.5 60670.0 7772.5 60735.0 ;
      RECT  7767.5 60915.0 7832.5 61050.0 ;
      RECT  7130.0 61607.5 8140.0 61672.5 ;
      RECT  7130.0 60262.5 8140.0 60327.5 ;
      RECT  7197.5 62822.5 7262.5 63017.5 ;
      RECT  7197.5 61982.5 7262.5 61607.5 ;
      RECT  7577.5 61982.5 7642.5 61607.5 ;
      RECT  7937.5 61825.0 8002.5 61640.0 ;
      RECT  7937.5 62985.0 8002.5 62800.0 ;
      RECT  7197.5 61982.5 7262.5 61847.5 ;
      RECT  7387.5 61982.5 7452.5 61847.5 ;
      RECT  7387.5 61982.5 7452.5 61847.5 ;
      RECT  7197.5 61982.5 7262.5 61847.5 ;
      RECT  7387.5 61982.5 7452.5 61847.5 ;
      RECT  7577.5 61982.5 7642.5 61847.5 ;
      RECT  7577.5 61982.5 7642.5 61847.5 ;
      RECT  7387.5 61982.5 7452.5 61847.5 ;
      RECT  7577.5 61982.5 7642.5 61847.5 ;
      RECT  7767.5 61982.5 7832.5 61847.5 ;
      RECT  7767.5 61982.5 7832.5 61847.5 ;
      RECT  7577.5 61982.5 7642.5 61847.5 ;
      RECT  7197.5 62822.5 7262.5 62687.5 ;
      RECT  7387.5 62822.5 7452.5 62687.5 ;
      RECT  7387.5 62822.5 7452.5 62687.5 ;
      RECT  7197.5 62822.5 7262.5 62687.5 ;
      RECT  7387.5 62822.5 7452.5 62687.5 ;
      RECT  7577.5 62822.5 7642.5 62687.5 ;
      RECT  7577.5 62822.5 7642.5 62687.5 ;
      RECT  7387.5 62822.5 7452.5 62687.5 ;
      RECT  7577.5 62822.5 7642.5 62687.5 ;
      RECT  7767.5 62822.5 7832.5 62687.5 ;
      RECT  7767.5 62822.5 7832.5 62687.5 ;
      RECT  7577.5 62822.5 7642.5 62687.5 ;
      RECT  7937.5 61892.5 8002.5 61757.5 ;
      RECT  7937.5 62867.5 8002.5 62732.5 ;
      RECT  7772.5 62610.0 7637.5 62545.0 ;
      RECT  7582.5 62470.0 7447.5 62405.0 ;
      RECT  7392.5 62330.0 7257.5 62265.0 ;
      RECT  7387.5 61982.5 7452.5 61847.5 ;
      RECT  7767.5 61982.5 7832.5 61847.5 ;
      RECT  7767.5 62822.5 7832.5 62687.5 ;
      RECT  7767.5 62365.0 7832.5 62230.0 ;
      RECT  7257.5 62330.0 7392.5 62265.0 ;
      RECT  7447.5 62470.0 7582.5 62405.0 ;
      RECT  7637.5 62610.0 7772.5 62545.0 ;
      RECT  7767.5 62365.0 7832.5 62230.0 ;
      RECT  7130.0 61672.5 8140.0 61607.5 ;
      RECT  7130.0 63017.5 8140.0 62952.5 ;
      RECT  7197.5 63147.5 7262.5 62952.5 ;
      RECT  7197.5 63987.5 7262.5 64362.5 ;
      RECT  7577.5 63987.5 7642.5 64362.5 ;
      RECT  7937.5 64145.0 8002.5 64330.0 ;
      RECT  7937.5 62985.0 8002.5 63170.0 ;
      RECT  7197.5 63987.5 7262.5 64122.5 ;
      RECT  7387.5 63987.5 7452.5 64122.5 ;
      RECT  7387.5 63987.5 7452.5 64122.5 ;
      RECT  7197.5 63987.5 7262.5 64122.5 ;
      RECT  7387.5 63987.5 7452.5 64122.5 ;
      RECT  7577.5 63987.5 7642.5 64122.5 ;
      RECT  7577.5 63987.5 7642.5 64122.5 ;
      RECT  7387.5 63987.5 7452.5 64122.5 ;
      RECT  7577.5 63987.5 7642.5 64122.5 ;
      RECT  7767.5 63987.5 7832.5 64122.5 ;
      RECT  7767.5 63987.5 7832.5 64122.5 ;
      RECT  7577.5 63987.5 7642.5 64122.5 ;
      RECT  7197.5 63147.5 7262.5 63282.5 ;
      RECT  7387.5 63147.5 7452.5 63282.5 ;
      RECT  7387.5 63147.5 7452.5 63282.5 ;
      RECT  7197.5 63147.5 7262.5 63282.5 ;
      RECT  7387.5 63147.5 7452.5 63282.5 ;
      RECT  7577.5 63147.5 7642.5 63282.5 ;
      RECT  7577.5 63147.5 7642.5 63282.5 ;
      RECT  7387.5 63147.5 7452.5 63282.5 ;
      RECT  7577.5 63147.5 7642.5 63282.5 ;
      RECT  7767.5 63147.5 7832.5 63282.5 ;
      RECT  7767.5 63147.5 7832.5 63282.5 ;
      RECT  7577.5 63147.5 7642.5 63282.5 ;
      RECT  7937.5 64077.5 8002.5 64212.5 ;
      RECT  7937.5 63102.5 8002.5 63237.5 ;
      RECT  7772.5 63360.0 7637.5 63425.0 ;
      RECT  7582.5 63500.0 7447.5 63565.0 ;
      RECT  7392.5 63640.0 7257.5 63705.0 ;
      RECT  7387.5 63987.5 7452.5 64122.5 ;
      RECT  7767.5 63987.5 7832.5 64122.5 ;
      RECT  7767.5 63147.5 7832.5 63282.5 ;
      RECT  7767.5 63605.0 7832.5 63740.0 ;
      RECT  7257.5 63640.0 7392.5 63705.0 ;
      RECT  7447.5 63500.0 7582.5 63565.0 ;
      RECT  7637.5 63360.0 7772.5 63425.0 ;
      RECT  7767.5 63605.0 7832.5 63740.0 ;
      RECT  7130.0 64297.5 8140.0 64362.5 ;
      RECT  7130.0 62952.5 8140.0 63017.5 ;
      RECT  7197.5 65512.5 7262.5 65707.5 ;
      RECT  7197.5 64672.5 7262.5 64297.5 ;
      RECT  7577.5 64672.5 7642.5 64297.5 ;
      RECT  7937.5 64515.0 8002.5 64330.0 ;
      RECT  7937.5 65675.0 8002.5 65490.0 ;
      RECT  7197.5 64672.5 7262.5 64537.5 ;
      RECT  7387.5 64672.5 7452.5 64537.5 ;
      RECT  7387.5 64672.5 7452.5 64537.5 ;
      RECT  7197.5 64672.5 7262.5 64537.5 ;
      RECT  7387.5 64672.5 7452.5 64537.5 ;
      RECT  7577.5 64672.5 7642.5 64537.5 ;
      RECT  7577.5 64672.5 7642.5 64537.5 ;
      RECT  7387.5 64672.5 7452.5 64537.5 ;
      RECT  7577.5 64672.5 7642.5 64537.5 ;
      RECT  7767.5 64672.5 7832.5 64537.5 ;
      RECT  7767.5 64672.5 7832.5 64537.5 ;
      RECT  7577.5 64672.5 7642.5 64537.5 ;
      RECT  7197.5 65512.5 7262.5 65377.5 ;
      RECT  7387.5 65512.5 7452.5 65377.5 ;
      RECT  7387.5 65512.5 7452.5 65377.5 ;
      RECT  7197.5 65512.5 7262.5 65377.5 ;
      RECT  7387.5 65512.5 7452.5 65377.5 ;
      RECT  7577.5 65512.5 7642.5 65377.5 ;
      RECT  7577.5 65512.5 7642.5 65377.5 ;
      RECT  7387.5 65512.5 7452.5 65377.5 ;
      RECT  7577.5 65512.5 7642.5 65377.5 ;
      RECT  7767.5 65512.5 7832.5 65377.5 ;
      RECT  7767.5 65512.5 7832.5 65377.5 ;
      RECT  7577.5 65512.5 7642.5 65377.5 ;
      RECT  7937.5 64582.5 8002.5 64447.5 ;
      RECT  7937.5 65557.5 8002.5 65422.5 ;
      RECT  7772.5 65300.0 7637.5 65235.0 ;
      RECT  7582.5 65160.0 7447.5 65095.0 ;
      RECT  7392.5 65020.0 7257.5 64955.0 ;
      RECT  7387.5 64672.5 7452.5 64537.5 ;
      RECT  7767.5 64672.5 7832.5 64537.5 ;
      RECT  7767.5 65512.5 7832.5 65377.5 ;
      RECT  7767.5 65055.0 7832.5 64920.0 ;
      RECT  7257.5 65020.0 7392.5 64955.0 ;
      RECT  7447.5 65160.0 7582.5 65095.0 ;
      RECT  7637.5 65300.0 7772.5 65235.0 ;
      RECT  7767.5 65055.0 7832.5 64920.0 ;
      RECT  7130.0 64362.5 8140.0 64297.5 ;
      RECT  7130.0 65707.5 8140.0 65642.5 ;
      RECT  7197.5 65837.5 7262.5 65642.5 ;
      RECT  7197.5 66677.5 7262.5 67052.5 ;
      RECT  7577.5 66677.5 7642.5 67052.5 ;
      RECT  7937.5 66835.0 8002.5 67020.0 ;
      RECT  7937.5 65675.0 8002.5 65860.0 ;
      RECT  7197.5 66677.5 7262.5 66812.5 ;
      RECT  7387.5 66677.5 7452.5 66812.5 ;
      RECT  7387.5 66677.5 7452.5 66812.5 ;
      RECT  7197.5 66677.5 7262.5 66812.5 ;
      RECT  7387.5 66677.5 7452.5 66812.5 ;
      RECT  7577.5 66677.5 7642.5 66812.5 ;
      RECT  7577.5 66677.5 7642.5 66812.5 ;
      RECT  7387.5 66677.5 7452.5 66812.5 ;
      RECT  7577.5 66677.5 7642.5 66812.5 ;
      RECT  7767.5 66677.5 7832.5 66812.5 ;
      RECT  7767.5 66677.5 7832.5 66812.5 ;
      RECT  7577.5 66677.5 7642.5 66812.5 ;
      RECT  7197.5 65837.5 7262.5 65972.5 ;
      RECT  7387.5 65837.5 7452.5 65972.5 ;
      RECT  7387.5 65837.5 7452.5 65972.5 ;
      RECT  7197.5 65837.5 7262.5 65972.5 ;
      RECT  7387.5 65837.5 7452.5 65972.5 ;
      RECT  7577.5 65837.5 7642.5 65972.5 ;
      RECT  7577.5 65837.5 7642.5 65972.5 ;
      RECT  7387.5 65837.5 7452.5 65972.5 ;
      RECT  7577.5 65837.5 7642.5 65972.5 ;
      RECT  7767.5 65837.5 7832.5 65972.5 ;
      RECT  7767.5 65837.5 7832.5 65972.5 ;
      RECT  7577.5 65837.5 7642.5 65972.5 ;
      RECT  7937.5 66767.5 8002.5 66902.5 ;
      RECT  7937.5 65792.5 8002.5 65927.5 ;
      RECT  7772.5 66050.0 7637.5 66115.0 ;
      RECT  7582.5 66190.0 7447.5 66255.0 ;
      RECT  7392.5 66330.0 7257.5 66395.0 ;
      RECT  7387.5 66677.5 7452.5 66812.5 ;
      RECT  7767.5 66677.5 7832.5 66812.5 ;
      RECT  7767.5 65837.5 7832.5 65972.5 ;
      RECT  7767.5 66295.0 7832.5 66430.0 ;
      RECT  7257.5 66330.0 7392.5 66395.0 ;
      RECT  7447.5 66190.0 7582.5 66255.0 ;
      RECT  7637.5 66050.0 7772.5 66115.0 ;
      RECT  7767.5 66295.0 7832.5 66430.0 ;
      RECT  7130.0 66987.5 8140.0 67052.5 ;
      RECT  7130.0 65642.5 8140.0 65707.5 ;
      RECT  7197.5 68202.5 7262.5 68397.5 ;
      RECT  7197.5 67362.5 7262.5 66987.5 ;
      RECT  7577.5 67362.5 7642.5 66987.5 ;
      RECT  7937.5 67205.0 8002.5 67020.0 ;
      RECT  7937.5 68365.0 8002.5 68180.0 ;
      RECT  7197.5 67362.5 7262.5 67227.5 ;
      RECT  7387.5 67362.5 7452.5 67227.5 ;
      RECT  7387.5 67362.5 7452.5 67227.5 ;
      RECT  7197.5 67362.5 7262.5 67227.5 ;
      RECT  7387.5 67362.5 7452.5 67227.5 ;
      RECT  7577.5 67362.5 7642.5 67227.5 ;
      RECT  7577.5 67362.5 7642.5 67227.5 ;
      RECT  7387.5 67362.5 7452.5 67227.5 ;
      RECT  7577.5 67362.5 7642.5 67227.5 ;
      RECT  7767.5 67362.5 7832.5 67227.5 ;
      RECT  7767.5 67362.5 7832.5 67227.5 ;
      RECT  7577.5 67362.5 7642.5 67227.5 ;
      RECT  7197.5 68202.5 7262.5 68067.5 ;
      RECT  7387.5 68202.5 7452.5 68067.5 ;
      RECT  7387.5 68202.5 7452.5 68067.5 ;
      RECT  7197.5 68202.5 7262.5 68067.5 ;
      RECT  7387.5 68202.5 7452.5 68067.5 ;
      RECT  7577.5 68202.5 7642.5 68067.5 ;
      RECT  7577.5 68202.5 7642.5 68067.5 ;
      RECT  7387.5 68202.5 7452.5 68067.5 ;
      RECT  7577.5 68202.5 7642.5 68067.5 ;
      RECT  7767.5 68202.5 7832.5 68067.5 ;
      RECT  7767.5 68202.5 7832.5 68067.5 ;
      RECT  7577.5 68202.5 7642.5 68067.5 ;
      RECT  7937.5 67272.5 8002.5 67137.5 ;
      RECT  7937.5 68247.5 8002.5 68112.5 ;
      RECT  7772.5 67990.0 7637.5 67925.0 ;
      RECT  7582.5 67850.0 7447.5 67785.0 ;
      RECT  7392.5 67710.0 7257.5 67645.0 ;
      RECT  7387.5 67362.5 7452.5 67227.5 ;
      RECT  7767.5 67362.5 7832.5 67227.5 ;
      RECT  7767.5 68202.5 7832.5 68067.5 ;
      RECT  7767.5 67745.0 7832.5 67610.0 ;
      RECT  7257.5 67710.0 7392.5 67645.0 ;
      RECT  7447.5 67850.0 7582.5 67785.0 ;
      RECT  7637.5 67990.0 7772.5 67925.0 ;
      RECT  7767.5 67745.0 7832.5 67610.0 ;
      RECT  7130.0 67052.5 8140.0 66987.5 ;
      RECT  7130.0 68397.5 8140.0 68332.5 ;
      RECT  7197.5 68527.5 7262.5 68332.5 ;
      RECT  7197.5 69367.5 7262.5 69742.5 ;
      RECT  7577.5 69367.5 7642.5 69742.5 ;
      RECT  7937.5 69525.0 8002.5 69710.0 ;
      RECT  7937.5 68365.0 8002.5 68550.0 ;
      RECT  7197.5 69367.5 7262.5 69502.5 ;
      RECT  7387.5 69367.5 7452.5 69502.5 ;
      RECT  7387.5 69367.5 7452.5 69502.5 ;
      RECT  7197.5 69367.5 7262.5 69502.5 ;
      RECT  7387.5 69367.5 7452.5 69502.5 ;
      RECT  7577.5 69367.5 7642.5 69502.5 ;
      RECT  7577.5 69367.5 7642.5 69502.5 ;
      RECT  7387.5 69367.5 7452.5 69502.5 ;
      RECT  7577.5 69367.5 7642.5 69502.5 ;
      RECT  7767.5 69367.5 7832.5 69502.5 ;
      RECT  7767.5 69367.5 7832.5 69502.5 ;
      RECT  7577.5 69367.5 7642.5 69502.5 ;
      RECT  7197.5 68527.5 7262.5 68662.5 ;
      RECT  7387.5 68527.5 7452.5 68662.5 ;
      RECT  7387.5 68527.5 7452.5 68662.5 ;
      RECT  7197.5 68527.5 7262.5 68662.5 ;
      RECT  7387.5 68527.5 7452.5 68662.5 ;
      RECT  7577.5 68527.5 7642.5 68662.5 ;
      RECT  7577.5 68527.5 7642.5 68662.5 ;
      RECT  7387.5 68527.5 7452.5 68662.5 ;
      RECT  7577.5 68527.5 7642.5 68662.5 ;
      RECT  7767.5 68527.5 7832.5 68662.5 ;
      RECT  7767.5 68527.5 7832.5 68662.5 ;
      RECT  7577.5 68527.5 7642.5 68662.5 ;
      RECT  7937.5 69457.5 8002.5 69592.5 ;
      RECT  7937.5 68482.5 8002.5 68617.5 ;
      RECT  7772.5 68740.0 7637.5 68805.0 ;
      RECT  7582.5 68880.0 7447.5 68945.0 ;
      RECT  7392.5 69020.0 7257.5 69085.0 ;
      RECT  7387.5 69367.5 7452.5 69502.5 ;
      RECT  7767.5 69367.5 7832.5 69502.5 ;
      RECT  7767.5 68527.5 7832.5 68662.5 ;
      RECT  7767.5 68985.0 7832.5 69120.0 ;
      RECT  7257.5 69020.0 7392.5 69085.0 ;
      RECT  7447.5 68880.0 7582.5 68945.0 ;
      RECT  7637.5 68740.0 7772.5 68805.0 ;
      RECT  7767.5 68985.0 7832.5 69120.0 ;
      RECT  7130.0 69677.5 8140.0 69742.5 ;
      RECT  7130.0 68332.5 8140.0 68397.5 ;
      RECT  7197.5 70892.5 7262.5 71087.5 ;
      RECT  7197.5 70052.5 7262.5 69677.5 ;
      RECT  7577.5 70052.5 7642.5 69677.5 ;
      RECT  7937.5 69895.0 8002.5 69710.0 ;
      RECT  7937.5 71055.0 8002.5 70870.0 ;
      RECT  7197.5 70052.5 7262.5 69917.5 ;
      RECT  7387.5 70052.5 7452.5 69917.5 ;
      RECT  7387.5 70052.5 7452.5 69917.5 ;
      RECT  7197.5 70052.5 7262.5 69917.5 ;
      RECT  7387.5 70052.5 7452.5 69917.5 ;
      RECT  7577.5 70052.5 7642.5 69917.5 ;
      RECT  7577.5 70052.5 7642.5 69917.5 ;
      RECT  7387.5 70052.5 7452.5 69917.5 ;
      RECT  7577.5 70052.5 7642.5 69917.5 ;
      RECT  7767.5 70052.5 7832.5 69917.5 ;
      RECT  7767.5 70052.5 7832.5 69917.5 ;
      RECT  7577.5 70052.5 7642.5 69917.5 ;
      RECT  7197.5 70892.5 7262.5 70757.5 ;
      RECT  7387.5 70892.5 7452.5 70757.5 ;
      RECT  7387.5 70892.5 7452.5 70757.5 ;
      RECT  7197.5 70892.5 7262.5 70757.5 ;
      RECT  7387.5 70892.5 7452.5 70757.5 ;
      RECT  7577.5 70892.5 7642.5 70757.5 ;
      RECT  7577.5 70892.5 7642.5 70757.5 ;
      RECT  7387.5 70892.5 7452.5 70757.5 ;
      RECT  7577.5 70892.5 7642.5 70757.5 ;
      RECT  7767.5 70892.5 7832.5 70757.5 ;
      RECT  7767.5 70892.5 7832.5 70757.5 ;
      RECT  7577.5 70892.5 7642.5 70757.5 ;
      RECT  7937.5 69962.5 8002.5 69827.5 ;
      RECT  7937.5 70937.5 8002.5 70802.5 ;
      RECT  7772.5 70680.0 7637.5 70615.0 ;
      RECT  7582.5 70540.0 7447.5 70475.0 ;
      RECT  7392.5 70400.0 7257.5 70335.0 ;
      RECT  7387.5 70052.5 7452.5 69917.5 ;
      RECT  7767.5 70052.5 7832.5 69917.5 ;
      RECT  7767.5 70892.5 7832.5 70757.5 ;
      RECT  7767.5 70435.0 7832.5 70300.0 ;
      RECT  7257.5 70400.0 7392.5 70335.0 ;
      RECT  7447.5 70540.0 7582.5 70475.0 ;
      RECT  7637.5 70680.0 7772.5 70615.0 ;
      RECT  7767.5 70435.0 7832.5 70300.0 ;
      RECT  7130.0 69742.5 8140.0 69677.5 ;
      RECT  7130.0 71087.5 8140.0 71022.5 ;
      RECT  7197.5 71217.5 7262.5 71022.5 ;
      RECT  7197.5 72057.5 7262.5 72432.5 ;
      RECT  7577.5 72057.5 7642.5 72432.5 ;
      RECT  7937.5 72215.0 8002.5 72400.0 ;
      RECT  7937.5 71055.0 8002.5 71240.0 ;
      RECT  7197.5 72057.5 7262.5 72192.5 ;
      RECT  7387.5 72057.5 7452.5 72192.5 ;
      RECT  7387.5 72057.5 7452.5 72192.5 ;
      RECT  7197.5 72057.5 7262.5 72192.5 ;
      RECT  7387.5 72057.5 7452.5 72192.5 ;
      RECT  7577.5 72057.5 7642.5 72192.5 ;
      RECT  7577.5 72057.5 7642.5 72192.5 ;
      RECT  7387.5 72057.5 7452.5 72192.5 ;
      RECT  7577.5 72057.5 7642.5 72192.5 ;
      RECT  7767.5 72057.5 7832.5 72192.5 ;
      RECT  7767.5 72057.5 7832.5 72192.5 ;
      RECT  7577.5 72057.5 7642.5 72192.5 ;
      RECT  7197.5 71217.5 7262.5 71352.5 ;
      RECT  7387.5 71217.5 7452.5 71352.5 ;
      RECT  7387.5 71217.5 7452.5 71352.5 ;
      RECT  7197.5 71217.5 7262.5 71352.5 ;
      RECT  7387.5 71217.5 7452.5 71352.5 ;
      RECT  7577.5 71217.5 7642.5 71352.5 ;
      RECT  7577.5 71217.5 7642.5 71352.5 ;
      RECT  7387.5 71217.5 7452.5 71352.5 ;
      RECT  7577.5 71217.5 7642.5 71352.5 ;
      RECT  7767.5 71217.5 7832.5 71352.5 ;
      RECT  7767.5 71217.5 7832.5 71352.5 ;
      RECT  7577.5 71217.5 7642.5 71352.5 ;
      RECT  7937.5 72147.5 8002.5 72282.5 ;
      RECT  7937.5 71172.5 8002.5 71307.5 ;
      RECT  7772.5 71430.0 7637.5 71495.0 ;
      RECT  7582.5 71570.0 7447.5 71635.0 ;
      RECT  7392.5 71710.0 7257.5 71775.0 ;
      RECT  7387.5 72057.5 7452.5 72192.5 ;
      RECT  7767.5 72057.5 7832.5 72192.5 ;
      RECT  7767.5 71217.5 7832.5 71352.5 ;
      RECT  7767.5 71675.0 7832.5 71810.0 ;
      RECT  7257.5 71710.0 7392.5 71775.0 ;
      RECT  7447.5 71570.0 7582.5 71635.0 ;
      RECT  7637.5 71430.0 7772.5 71495.0 ;
      RECT  7767.5 71675.0 7832.5 71810.0 ;
      RECT  7130.0 72367.5 8140.0 72432.5 ;
      RECT  7130.0 71022.5 8140.0 71087.5 ;
      RECT  7197.5 73582.5 7262.5 73777.5 ;
      RECT  7197.5 72742.5 7262.5 72367.5 ;
      RECT  7577.5 72742.5 7642.5 72367.5 ;
      RECT  7937.5 72585.0 8002.5 72400.0 ;
      RECT  7937.5 73745.0 8002.5 73560.0 ;
      RECT  7197.5 72742.5 7262.5 72607.5 ;
      RECT  7387.5 72742.5 7452.5 72607.5 ;
      RECT  7387.5 72742.5 7452.5 72607.5 ;
      RECT  7197.5 72742.5 7262.5 72607.5 ;
      RECT  7387.5 72742.5 7452.5 72607.5 ;
      RECT  7577.5 72742.5 7642.5 72607.5 ;
      RECT  7577.5 72742.5 7642.5 72607.5 ;
      RECT  7387.5 72742.5 7452.5 72607.5 ;
      RECT  7577.5 72742.5 7642.5 72607.5 ;
      RECT  7767.5 72742.5 7832.5 72607.5 ;
      RECT  7767.5 72742.5 7832.5 72607.5 ;
      RECT  7577.5 72742.5 7642.5 72607.5 ;
      RECT  7197.5 73582.5 7262.5 73447.5 ;
      RECT  7387.5 73582.5 7452.5 73447.5 ;
      RECT  7387.5 73582.5 7452.5 73447.5 ;
      RECT  7197.5 73582.5 7262.5 73447.5 ;
      RECT  7387.5 73582.5 7452.5 73447.5 ;
      RECT  7577.5 73582.5 7642.5 73447.5 ;
      RECT  7577.5 73582.5 7642.5 73447.5 ;
      RECT  7387.5 73582.5 7452.5 73447.5 ;
      RECT  7577.5 73582.5 7642.5 73447.5 ;
      RECT  7767.5 73582.5 7832.5 73447.5 ;
      RECT  7767.5 73582.5 7832.5 73447.5 ;
      RECT  7577.5 73582.5 7642.5 73447.5 ;
      RECT  7937.5 72652.5 8002.5 72517.5 ;
      RECT  7937.5 73627.5 8002.5 73492.5 ;
      RECT  7772.5 73370.0 7637.5 73305.0 ;
      RECT  7582.5 73230.0 7447.5 73165.0 ;
      RECT  7392.5 73090.0 7257.5 73025.0 ;
      RECT  7387.5 72742.5 7452.5 72607.5 ;
      RECT  7767.5 72742.5 7832.5 72607.5 ;
      RECT  7767.5 73582.5 7832.5 73447.5 ;
      RECT  7767.5 73125.0 7832.5 72990.0 ;
      RECT  7257.5 73090.0 7392.5 73025.0 ;
      RECT  7447.5 73230.0 7582.5 73165.0 ;
      RECT  7637.5 73370.0 7772.5 73305.0 ;
      RECT  7767.5 73125.0 7832.5 72990.0 ;
      RECT  7130.0 72432.5 8140.0 72367.5 ;
      RECT  7130.0 73777.5 8140.0 73712.5 ;
      RECT  7197.5 73907.5 7262.5 73712.5 ;
      RECT  7197.5 74747.5 7262.5 75122.5 ;
      RECT  7577.5 74747.5 7642.5 75122.5 ;
      RECT  7937.5 74905.0 8002.5 75090.0 ;
      RECT  7937.5 73745.0 8002.5 73930.0 ;
      RECT  7197.5 74747.5 7262.5 74882.5 ;
      RECT  7387.5 74747.5 7452.5 74882.5 ;
      RECT  7387.5 74747.5 7452.5 74882.5 ;
      RECT  7197.5 74747.5 7262.5 74882.5 ;
      RECT  7387.5 74747.5 7452.5 74882.5 ;
      RECT  7577.5 74747.5 7642.5 74882.5 ;
      RECT  7577.5 74747.5 7642.5 74882.5 ;
      RECT  7387.5 74747.5 7452.5 74882.5 ;
      RECT  7577.5 74747.5 7642.5 74882.5 ;
      RECT  7767.5 74747.5 7832.5 74882.5 ;
      RECT  7767.5 74747.5 7832.5 74882.5 ;
      RECT  7577.5 74747.5 7642.5 74882.5 ;
      RECT  7197.5 73907.5 7262.5 74042.5 ;
      RECT  7387.5 73907.5 7452.5 74042.5 ;
      RECT  7387.5 73907.5 7452.5 74042.5 ;
      RECT  7197.5 73907.5 7262.5 74042.5 ;
      RECT  7387.5 73907.5 7452.5 74042.5 ;
      RECT  7577.5 73907.5 7642.5 74042.5 ;
      RECT  7577.5 73907.5 7642.5 74042.5 ;
      RECT  7387.5 73907.5 7452.5 74042.5 ;
      RECT  7577.5 73907.5 7642.5 74042.5 ;
      RECT  7767.5 73907.5 7832.5 74042.5 ;
      RECT  7767.5 73907.5 7832.5 74042.5 ;
      RECT  7577.5 73907.5 7642.5 74042.5 ;
      RECT  7937.5 74837.5 8002.5 74972.5 ;
      RECT  7937.5 73862.5 8002.5 73997.5 ;
      RECT  7772.5 74120.0 7637.5 74185.0 ;
      RECT  7582.5 74260.0 7447.5 74325.0 ;
      RECT  7392.5 74400.0 7257.5 74465.0 ;
      RECT  7387.5 74747.5 7452.5 74882.5 ;
      RECT  7767.5 74747.5 7832.5 74882.5 ;
      RECT  7767.5 73907.5 7832.5 74042.5 ;
      RECT  7767.5 74365.0 7832.5 74500.0 ;
      RECT  7257.5 74400.0 7392.5 74465.0 ;
      RECT  7447.5 74260.0 7582.5 74325.0 ;
      RECT  7637.5 74120.0 7772.5 74185.0 ;
      RECT  7767.5 74365.0 7832.5 74500.0 ;
      RECT  7130.0 75057.5 8140.0 75122.5 ;
      RECT  7130.0 73712.5 8140.0 73777.5 ;
      RECT  7197.5 76272.5 7262.5 76467.5 ;
      RECT  7197.5 75432.5 7262.5 75057.5 ;
      RECT  7577.5 75432.5 7642.5 75057.5 ;
      RECT  7937.5 75275.0 8002.5 75090.0 ;
      RECT  7937.5 76435.0 8002.5 76250.0 ;
      RECT  7197.5 75432.5 7262.5 75297.5 ;
      RECT  7387.5 75432.5 7452.5 75297.5 ;
      RECT  7387.5 75432.5 7452.5 75297.5 ;
      RECT  7197.5 75432.5 7262.5 75297.5 ;
      RECT  7387.5 75432.5 7452.5 75297.5 ;
      RECT  7577.5 75432.5 7642.5 75297.5 ;
      RECT  7577.5 75432.5 7642.5 75297.5 ;
      RECT  7387.5 75432.5 7452.5 75297.5 ;
      RECT  7577.5 75432.5 7642.5 75297.5 ;
      RECT  7767.5 75432.5 7832.5 75297.5 ;
      RECT  7767.5 75432.5 7832.5 75297.5 ;
      RECT  7577.5 75432.5 7642.5 75297.5 ;
      RECT  7197.5 76272.5 7262.5 76137.5 ;
      RECT  7387.5 76272.5 7452.5 76137.5 ;
      RECT  7387.5 76272.5 7452.5 76137.5 ;
      RECT  7197.5 76272.5 7262.5 76137.5 ;
      RECT  7387.5 76272.5 7452.5 76137.5 ;
      RECT  7577.5 76272.5 7642.5 76137.5 ;
      RECT  7577.5 76272.5 7642.5 76137.5 ;
      RECT  7387.5 76272.5 7452.5 76137.5 ;
      RECT  7577.5 76272.5 7642.5 76137.5 ;
      RECT  7767.5 76272.5 7832.5 76137.5 ;
      RECT  7767.5 76272.5 7832.5 76137.5 ;
      RECT  7577.5 76272.5 7642.5 76137.5 ;
      RECT  7937.5 75342.5 8002.5 75207.5 ;
      RECT  7937.5 76317.5 8002.5 76182.5 ;
      RECT  7772.5 76060.0 7637.5 75995.0 ;
      RECT  7582.5 75920.0 7447.5 75855.0 ;
      RECT  7392.5 75780.0 7257.5 75715.0 ;
      RECT  7387.5 75432.5 7452.5 75297.5 ;
      RECT  7767.5 75432.5 7832.5 75297.5 ;
      RECT  7767.5 76272.5 7832.5 76137.5 ;
      RECT  7767.5 75815.0 7832.5 75680.0 ;
      RECT  7257.5 75780.0 7392.5 75715.0 ;
      RECT  7447.5 75920.0 7582.5 75855.0 ;
      RECT  7637.5 76060.0 7772.5 75995.0 ;
      RECT  7767.5 75815.0 7832.5 75680.0 ;
      RECT  7130.0 75122.5 8140.0 75057.5 ;
      RECT  7130.0 76467.5 8140.0 76402.5 ;
      RECT  7197.5 76597.5 7262.5 76402.5 ;
      RECT  7197.5 77437.5 7262.5 77812.5 ;
      RECT  7577.5 77437.5 7642.5 77812.5 ;
      RECT  7937.5 77595.0 8002.5 77780.0 ;
      RECT  7937.5 76435.0 8002.5 76620.0 ;
      RECT  7197.5 77437.5 7262.5 77572.5 ;
      RECT  7387.5 77437.5 7452.5 77572.5 ;
      RECT  7387.5 77437.5 7452.5 77572.5 ;
      RECT  7197.5 77437.5 7262.5 77572.5 ;
      RECT  7387.5 77437.5 7452.5 77572.5 ;
      RECT  7577.5 77437.5 7642.5 77572.5 ;
      RECT  7577.5 77437.5 7642.5 77572.5 ;
      RECT  7387.5 77437.5 7452.5 77572.5 ;
      RECT  7577.5 77437.5 7642.5 77572.5 ;
      RECT  7767.5 77437.5 7832.5 77572.5 ;
      RECT  7767.5 77437.5 7832.5 77572.5 ;
      RECT  7577.5 77437.5 7642.5 77572.5 ;
      RECT  7197.5 76597.5 7262.5 76732.5 ;
      RECT  7387.5 76597.5 7452.5 76732.5 ;
      RECT  7387.5 76597.5 7452.5 76732.5 ;
      RECT  7197.5 76597.5 7262.5 76732.5 ;
      RECT  7387.5 76597.5 7452.5 76732.5 ;
      RECT  7577.5 76597.5 7642.5 76732.5 ;
      RECT  7577.5 76597.5 7642.5 76732.5 ;
      RECT  7387.5 76597.5 7452.5 76732.5 ;
      RECT  7577.5 76597.5 7642.5 76732.5 ;
      RECT  7767.5 76597.5 7832.5 76732.5 ;
      RECT  7767.5 76597.5 7832.5 76732.5 ;
      RECT  7577.5 76597.5 7642.5 76732.5 ;
      RECT  7937.5 77527.5 8002.5 77662.5 ;
      RECT  7937.5 76552.5 8002.5 76687.5 ;
      RECT  7772.5 76810.0 7637.5 76875.0 ;
      RECT  7582.5 76950.0 7447.5 77015.0 ;
      RECT  7392.5 77090.0 7257.5 77155.0 ;
      RECT  7387.5 77437.5 7452.5 77572.5 ;
      RECT  7767.5 77437.5 7832.5 77572.5 ;
      RECT  7767.5 76597.5 7832.5 76732.5 ;
      RECT  7767.5 77055.0 7832.5 77190.0 ;
      RECT  7257.5 77090.0 7392.5 77155.0 ;
      RECT  7447.5 76950.0 7582.5 77015.0 ;
      RECT  7637.5 76810.0 7772.5 76875.0 ;
      RECT  7767.5 77055.0 7832.5 77190.0 ;
      RECT  7130.0 77747.5 8140.0 77812.5 ;
      RECT  7130.0 76402.5 8140.0 76467.5 ;
      RECT  7197.5 78962.5 7262.5 79157.5 ;
      RECT  7197.5 78122.5 7262.5 77747.5 ;
      RECT  7577.5 78122.5 7642.5 77747.5 ;
      RECT  7937.5 77965.0 8002.5 77780.0 ;
      RECT  7937.5 79125.0 8002.5 78940.0 ;
      RECT  7197.5 78122.5 7262.5 77987.5 ;
      RECT  7387.5 78122.5 7452.5 77987.5 ;
      RECT  7387.5 78122.5 7452.5 77987.5 ;
      RECT  7197.5 78122.5 7262.5 77987.5 ;
      RECT  7387.5 78122.5 7452.5 77987.5 ;
      RECT  7577.5 78122.5 7642.5 77987.5 ;
      RECT  7577.5 78122.5 7642.5 77987.5 ;
      RECT  7387.5 78122.5 7452.5 77987.5 ;
      RECT  7577.5 78122.5 7642.5 77987.5 ;
      RECT  7767.5 78122.5 7832.5 77987.5 ;
      RECT  7767.5 78122.5 7832.5 77987.5 ;
      RECT  7577.5 78122.5 7642.5 77987.5 ;
      RECT  7197.5 78962.5 7262.5 78827.5 ;
      RECT  7387.5 78962.5 7452.5 78827.5 ;
      RECT  7387.5 78962.5 7452.5 78827.5 ;
      RECT  7197.5 78962.5 7262.5 78827.5 ;
      RECT  7387.5 78962.5 7452.5 78827.5 ;
      RECT  7577.5 78962.5 7642.5 78827.5 ;
      RECT  7577.5 78962.5 7642.5 78827.5 ;
      RECT  7387.5 78962.5 7452.5 78827.5 ;
      RECT  7577.5 78962.5 7642.5 78827.5 ;
      RECT  7767.5 78962.5 7832.5 78827.5 ;
      RECT  7767.5 78962.5 7832.5 78827.5 ;
      RECT  7577.5 78962.5 7642.5 78827.5 ;
      RECT  7937.5 78032.5 8002.5 77897.5 ;
      RECT  7937.5 79007.5 8002.5 78872.5 ;
      RECT  7772.5 78750.0 7637.5 78685.0 ;
      RECT  7582.5 78610.0 7447.5 78545.0 ;
      RECT  7392.5 78470.0 7257.5 78405.0 ;
      RECT  7387.5 78122.5 7452.5 77987.5 ;
      RECT  7767.5 78122.5 7832.5 77987.5 ;
      RECT  7767.5 78962.5 7832.5 78827.5 ;
      RECT  7767.5 78505.0 7832.5 78370.0 ;
      RECT  7257.5 78470.0 7392.5 78405.0 ;
      RECT  7447.5 78610.0 7582.5 78545.0 ;
      RECT  7637.5 78750.0 7772.5 78685.0 ;
      RECT  7767.5 78505.0 7832.5 78370.0 ;
      RECT  7130.0 77812.5 8140.0 77747.5 ;
      RECT  7130.0 79157.5 8140.0 79092.5 ;
      RECT  7197.5 79287.5 7262.5 79092.5 ;
      RECT  7197.5 80127.5 7262.5 80502.5 ;
      RECT  7577.5 80127.5 7642.5 80502.5 ;
      RECT  7937.5 80285.0 8002.5 80470.0 ;
      RECT  7937.5 79125.0 8002.5 79310.0 ;
      RECT  7197.5 80127.5 7262.5 80262.5 ;
      RECT  7387.5 80127.5 7452.5 80262.5 ;
      RECT  7387.5 80127.5 7452.5 80262.5 ;
      RECT  7197.5 80127.5 7262.5 80262.5 ;
      RECT  7387.5 80127.5 7452.5 80262.5 ;
      RECT  7577.5 80127.5 7642.5 80262.5 ;
      RECT  7577.5 80127.5 7642.5 80262.5 ;
      RECT  7387.5 80127.5 7452.5 80262.5 ;
      RECT  7577.5 80127.5 7642.5 80262.5 ;
      RECT  7767.5 80127.5 7832.5 80262.5 ;
      RECT  7767.5 80127.5 7832.5 80262.5 ;
      RECT  7577.5 80127.5 7642.5 80262.5 ;
      RECT  7197.5 79287.5 7262.5 79422.5 ;
      RECT  7387.5 79287.5 7452.5 79422.5 ;
      RECT  7387.5 79287.5 7452.5 79422.5 ;
      RECT  7197.5 79287.5 7262.5 79422.5 ;
      RECT  7387.5 79287.5 7452.5 79422.5 ;
      RECT  7577.5 79287.5 7642.5 79422.5 ;
      RECT  7577.5 79287.5 7642.5 79422.5 ;
      RECT  7387.5 79287.5 7452.5 79422.5 ;
      RECT  7577.5 79287.5 7642.5 79422.5 ;
      RECT  7767.5 79287.5 7832.5 79422.5 ;
      RECT  7767.5 79287.5 7832.5 79422.5 ;
      RECT  7577.5 79287.5 7642.5 79422.5 ;
      RECT  7937.5 80217.5 8002.5 80352.5 ;
      RECT  7937.5 79242.5 8002.5 79377.5 ;
      RECT  7772.5 79500.0 7637.5 79565.0 ;
      RECT  7582.5 79640.0 7447.5 79705.0 ;
      RECT  7392.5 79780.0 7257.5 79845.0 ;
      RECT  7387.5 80127.5 7452.5 80262.5 ;
      RECT  7767.5 80127.5 7832.5 80262.5 ;
      RECT  7767.5 79287.5 7832.5 79422.5 ;
      RECT  7767.5 79745.0 7832.5 79880.0 ;
      RECT  7257.5 79780.0 7392.5 79845.0 ;
      RECT  7447.5 79640.0 7582.5 79705.0 ;
      RECT  7637.5 79500.0 7772.5 79565.0 ;
      RECT  7767.5 79745.0 7832.5 79880.0 ;
      RECT  7130.0 80437.5 8140.0 80502.5 ;
      RECT  7130.0 79092.5 8140.0 79157.5 ;
      RECT  7197.5 81652.5 7262.5 81847.5 ;
      RECT  7197.5 80812.5 7262.5 80437.5 ;
      RECT  7577.5 80812.5 7642.5 80437.5 ;
      RECT  7937.5 80655.0 8002.5 80470.0 ;
      RECT  7937.5 81815.0 8002.5 81630.0 ;
      RECT  7197.5 80812.5 7262.5 80677.5 ;
      RECT  7387.5 80812.5 7452.5 80677.5 ;
      RECT  7387.5 80812.5 7452.5 80677.5 ;
      RECT  7197.5 80812.5 7262.5 80677.5 ;
      RECT  7387.5 80812.5 7452.5 80677.5 ;
      RECT  7577.5 80812.5 7642.5 80677.5 ;
      RECT  7577.5 80812.5 7642.5 80677.5 ;
      RECT  7387.5 80812.5 7452.5 80677.5 ;
      RECT  7577.5 80812.5 7642.5 80677.5 ;
      RECT  7767.5 80812.5 7832.5 80677.5 ;
      RECT  7767.5 80812.5 7832.5 80677.5 ;
      RECT  7577.5 80812.5 7642.5 80677.5 ;
      RECT  7197.5 81652.5 7262.5 81517.5 ;
      RECT  7387.5 81652.5 7452.5 81517.5 ;
      RECT  7387.5 81652.5 7452.5 81517.5 ;
      RECT  7197.5 81652.5 7262.5 81517.5 ;
      RECT  7387.5 81652.5 7452.5 81517.5 ;
      RECT  7577.5 81652.5 7642.5 81517.5 ;
      RECT  7577.5 81652.5 7642.5 81517.5 ;
      RECT  7387.5 81652.5 7452.5 81517.5 ;
      RECT  7577.5 81652.5 7642.5 81517.5 ;
      RECT  7767.5 81652.5 7832.5 81517.5 ;
      RECT  7767.5 81652.5 7832.5 81517.5 ;
      RECT  7577.5 81652.5 7642.5 81517.5 ;
      RECT  7937.5 80722.5 8002.5 80587.5 ;
      RECT  7937.5 81697.5 8002.5 81562.5 ;
      RECT  7772.5 81440.0 7637.5 81375.0 ;
      RECT  7582.5 81300.0 7447.5 81235.0 ;
      RECT  7392.5 81160.0 7257.5 81095.0 ;
      RECT  7387.5 80812.5 7452.5 80677.5 ;
      RECT  7767.5 80812.5 7832.5 80677.5 ;
      RECT  7767.5 81652.5 7832.5 81517.5 ;
      RECT  7767.5 81195.0 7832.5 81060.0 ;
      RECT  7257.5 81160.0 7392.5 81095.0 ;
      RECT  7447.5 81300.0 7582.5 81235.0 ;
      RECT  7637.5 81440.0 7772.5 81375.0 ;
      RECT  7767.5 81195.0 7832.5 81060.0 ;
      RECT  7130.0 80502.5 8140.0 80437.5 ;
      RECT  7130.0 81847.5 8140.0 81782.5 ;
      RECT  7197.5 81977.5 7262.5 81782.5 ;
      RECT  7197.5 82817.5 7262.5 83192.5 ;
      RECT  7577.5 82817.5 7642.5 83192.5 ;
      RECT  7937.5 82975.0 8002.5 83160.0 ;
      RECT  7937.5 81815.0 8002.5 82000.0 ;
      RECT  7197.5 82817.5 7262.5 82952.5 ;
      RECT  7387.5 82817.5 7452.5 82952.5 ;
      RECT  7387.5 82817.5 7452.5 82952.5 ;
      RECT  7197.5 82817.5 7262.5 82952.5 ;
      RECT  7387.5 82817.5 7452.5 82952.5 ;
      RECT  7577.5 82817.5 7642.5 82952.5 ;
      RECT  7577.5 82817.5 7642.5 82952.5 ;
      RECT  7387.5 82817.5 7452.5 82952.5 ;
      RECT  7577.5 82817.5 7642.5 82952.5 ;
      RECT  7767.5 82817.5 7832.5 82952.5 ;
      RECT  7767.5 82817.5 7832.5 82952.5 ;
      RECT  7577.5 82817.5 7642.5 82952.5 ;
      RECT  7197.5 81977.5 7262.5 82112.5 ;
      RECT  7387.5 81977.5 7452.5 82112.5 ;
      RECT  7387.5 81977.5 7452.5 82112.5 ;
      RECT  7197.5 81977.5 7262.5 82112.5 ;
      RECT  7387.5 81977.5 7452.5 82112.5 ;
      RECT  7577.5 81977.5 7642.5 82112.5 ;
      RECT  7577.5 81977.5 7642.5 82112.5 ;
      RECT  7387.5 81977.5 7452.5 82112.5 ;
      RECT  7577.5 81977.5 7642.5 82112.5 ;
      RECT  7767.5 81977.5 7832.5 82112.5 ;
      RECT  7767.5 81977.5 7832.5 82112.5 ;
      RECT  7577.5 81977.5 7642.5 82112.5 ;
      RECT  7937.5 82907.5 8002.5 83042.5 ;
      RECT  7937.5 81932.5 8002.5 82067.5 ;
      RECT  7772.5 82190.0 7637.5 82255.0 ;
      RECT  7582.5 82330.0 7447.5 82395.0 ;
      RECT  7392.5 82470.0 7257.5 82535.0 ;
      RECT  7387.5 82817.5 7452.5 82952.5 ;
      RECT  7767.5 82817.5 7832.5 82952.5 ;
      RECT  7767.5 81977.5 7832.5 82112.5 ;
      RECT  7767.5 82435.0 7832.5 82570.0 ;
      RECT  7257.5 82470.0 7392.5 82535.0 ;
      RECT  7447.5 82330.0 7582.5 82395.0 ;
      RECT  7637.5 82190.0 7772.5 82255.0 ;
      RECT  7767.5 82435.0 7832.5 82570.0 ;
      RECT  7130.0 83127.5 8140.0 83192.5 ;
      RECT  7130.0 81782.5 8140.0 81847.5 ;
      RECT  7197.5 84342.5 7262.5 84537.5 ;
      RECT  7197.5 83502.5 7262.5 83127.5 ;
      RECT  7577.5 83502.5 7642.5 83127.5 ;
      RECT  7937.5 83345.0 8002.5 83160.0 ;
      RECT  7937.5 84505.0 8002.5 84320.0 ;
      RECT  7197.5 83502.5 7262.5 83367.5 ;
      RECT  7387.5 83502.5 7452.5 83367.5 ;
      RECT  7387.5 83502.5 7452.5 83367.5 ;
      RECT  7197.5 83502.5 7262.5 83367.5 ;
      RECT  7387.5 83502.5 7452.5 83367.5 ;
      RECT  7577.5 83502.5 7642.5 83367.5 ;
      RECT  7577.5 83502.5 7642.5 83367.5 ;
      RECT  7387.5 83502.5 7452.5 83367.5 ;
      RECT  7577.5 83502.5 7642.5 83367.5 ;
      RECT  7767.5 83502.5 7832.5 83367.5 ;
      RECT  7767.5 83502.5 7832.5 83367.5 ;
      RECT  7577.5 83502.5 7642.5 83367.5 ;
      RECT  7197.5 84342.5 7262.5 84207.5 ;
      RECT  7387.5 84342.5 7452.5 84207.5 ;
      RECT  7387.5 84342.5 7452.5 84207.5 ;
      RECT  7197.5 84342.5 7262.5 84207.5 ;
      RECT  7387.5 84342.5 7452.5 84207.5 ;
      RECT  7577.5 84342.5 7642.5 84207.5 ;
      RECT  7577.5 84342.5 7642.5 84207.5 ;
      RECT  7387.5 84342.5 7452.5 84207.5 ;
      RECT  7577.5 84342.5 7642.5 84207.5 ;
      RECT  7767.5 84342.5 7832.5 84207.5 ;
      RECT  7767.5 84342.5 7832.5 84207.5 ;
      RECT  7577.5 84342.5 7642.5 84207.5 ;
      RECT  7937.5 83412.5 8002.5 83277.5 ;
      RECT  7937.5 84387.5 8002.5 84252.5 ;
      RECT  7772.5 84130.0 7637.5 84065.0 ;
      RECT  7582.5 83990.0 7447.5 83925.0 ;
      RECT  7392.5 83850.0 7257.5 83785.0 ;
      RECT  7387.5 83502.5 7452.5 83367.5 ;
      RECT  7767.5 83502.5 7832.5 83367.5 ;
      RECT  7767.5 84342.5 7832.5 84207.5 ;
      RECT  7767.5 83885.0 7832.5 83750.0 ;
      RECT  7257.5 83850.0 7392.5 83785.0 ;
      RECT  7447.5 83990.0 7582.5 83925.0 ;
      RECT  7637.5 84130.0 7772.5 84065.0 ;
      RECT  7767.5 83885.0 7832.5 83750.0 ;
      RECT  7130.0 83192.5 8140.0 83127.5 ;
      RECT  7130.0 84537.5 8140.0 84472.5 ;
      RECT  7197.5 84667.5 7262.5 84472.5 ;
      RECT  7197.5 85507.5 7262.5 85882.5 ;
      RECT  7577.5 85507.5 7642.5 85882.5 ;
      RECT  7937.5 85665.0 8002.5 85850.0 ;
      RECT  7937.5 84505.0 8002.5 84690.0 ;
      RECT  7197.5 85507.5 7262.5 85642.5 ;
      RECT  7387.5 85507.5 7452.5 85642.5 ;
      RECT  7387.5 85507.5 7452.5 85642.5 ;
      RECT  7197.5 85507.5 7262.5 85642.5 ;
      RECT  7387.5 85507.5 7452.5 85642.5 ;
      RECT  7577.5 85507.5 7642.5 85642.5 ;
      RECT  7577.5 85507.5 7642.5 85642.5 ;
      RECT  7387.5 85507.5 7452.5 85642.5 ;
      RECT  7577.5 85507.5 7642.5 85642.5 ;
      RECT  7767.5 85507.5 7832.5 85642.5 ;
      RECT  7767.5 85507.5 7832.5 85642.5 ;
      RECT  7577.5 85507.5 7642.5 85642.5 ;
      RECT  7197.5 84667.5 7262.5 84802.5 ;
      RECT  7387.5 84667.5 7452.5 84802.5 ;
      RECT  7387.5 84667.5 7452.5 84802.5 ;
      RECT  7197.5 84667.5 7262.5 84802.5 ;
      RECT  7387.5 84667.5 7452.5 84802.5 ;
      RECT  7577.5 84667.5 7642.5 84802.5 ;
      RECT  7577.5 84667.5 7642.5 84802.5 ;
      RECT  7387.5 84667.5 7452.5 84802.5 ;
      RECT  7577.5 84667.5 7642.5 84802.5 ;
      RECT  7767.5 84667.5 7832.5 84802.5 ;
      RECT  7767.5 84667.5 7832.5 84802.5 ;
      RECT  7577.5 84667.5 7642.5 84802.5 ;
      RECT  7937.5 85597.5 8002.5 85732.5 ;
      RECT  7937.5 84622.5 8002.5 84757.5 ;
      RECT  7772.5 84880.0 7637.5 84945.0 ;
      RECT  7582.5 85020.0 7447.5 85085.0 ;
      RECT  7392.5 85160.0 7257.5 85225.0 ;
      RECT  7387.5 85507.5 7452.5 85642.5 ;
      RECT  7767.5 85507.5 7832.5 85642.5 ;
      RECT  7767.5 84667.5 7832.5 84802.5 ;
      RECT  7767.5 85125.0 7832.5 85260.0 ;
      RECT  7257.5 85160.0 7392.5 85225.0 ;
      RECT  7447.5 85020.0 7582.5 85085.0 ;
      RECT  7637.5 84880.0 7772.5 84945.0 ;
      RECT  7767.5 85125.0 7832.5 85260.0 ;
      RECT  7130.0 85817.5 8140.0 85882.5 ;
      RECT  7130.0 84472.5 8140.0 84537.5 ;
      RECT  7197.5 87032.5 7262.5 87227.5 ;
      RECT  7197.5 86192.5 7262.5 85817.5 ;
      RECT  7577.5 86192.5 7642.5 85817.5 ;
      RECT  7937.5 86035.0 8002.5 85850.0 ;
      RECT  7937.5 87195.0 8002.5 87010.0 ;
      RECT  7197.5 86192.5 7262.5 86057.5 ;
      RECT  7387.5 86192.5 7452.5 86057.5 ;
      RECT  7387.5 86192.5 7452.5 86057.5 ;
      RECT  7197.5 86192.5 7262.5 86057.5 ;
      RECT  7387.5 86192.5 7452.5 86057.5 ;
      RECT  7577.5 86192.5 7642.5 86057.5 ;
      RECT  7577.5 86192.5 7642.5 86057.5 ;
      RECT  7387.5 86192.5 7452.5 86057.5 ;
      RECT  7577.5 86192.5 7642.5 86057.5 ;
      RECT  7767.5 86192.5 7832.5 86057.5 ;
      RECT  7767.5 86192.5 7832.5 86057.5 ;
      RECT  7577.5 86192.5 7642.5 86057.5 ;
      RECT  7197.5 87032.5 7262.5 86897.5 ;
      RECT  7387.5 87032.5 7452.5 86897.5 ;
      RECT  7387.5 87032.5 7452.5 86897.5 ;
      RECT  7197.5 87032.5 7262.5 86897.5 ;
      RECT  7387.5 87032.5 7452.5 86897.5 ;
      RECT  7577.5 87032.5 7642.5 86897.5 ;
      RECT  7577.5 87032.5 7642.5 86897.5 ;
      RECT  7387.5 87032.5 7452.5 86897.5 ;
      RECT  7577.5 87032.5 7642.5 86897.5 ;
      RECT  7767.5 87032.5 7832.5 86897.5 ;
      RECT  7767.5 87032.5 7832.5 86897.5 ;
      RECT  7577.5 87032.5 7642.5 86897.5 ;
      RECT  7937.5 86102.5 8002.5 85967.5 ;
      RECT  7937.5 87077.5 8002.5 86942.5 ;
      RECT  7772.5 86820.0 7637.5 86755.0 ;
      RECT  7582.5 86680.0 7447.5 86615.0 ;
      RECT  7392.5 86540.0 7257.5 86475.0 ;
      RECT  7387.5 86192.5 7452.5 86057.5 ;
      RECT  7767.5 86192.5 7832.5 86057.5 ;
      RECT  7767.5 87032.5 7832.5 86897.5 ;
      RECT  7767.5 86575.0 7832.5 86440.0 ;
      RECT  7257.5 86540.0 7392.5 86475.0 ;
      RECT  7447.5 86680.0 7582.5 86615.0 ;
      RECT  7637.5 86820.0 7772.5 86755.0 ;
      RECT  7767.5 86575.0 7832.5 86440.0 ;
      RECT  7130.0 85882.5 8140.0 85817.5 ;
      RECT  7130.0 87227.5 8140.0 87162.5 ;
      RECT  7197.5 87357.5 7262.5 87162.5 ;
      RECT  7197.5 88197.5 7262.5 88572.5 ;
      RECT  7577.5 88197.5 7642.5 88572.5 ;
      RECT  7937.5 88355.0 8002.5 88540.0 ;
      RECT  7937.5 87195.0 8002.5 87380.0 ;
      RECT  7197.5 88197.5 7262.5 88332.5 ;
      RECT  7387.5 88197.5 7452.5 88332.5 ;
      RECT  7387.5 88197.5 7452.5 88332.5 ;
      RECT  7197.5 88197.5 7262.5 88332.5 ;
      RECT  7387.5 88197.5 7452.5 88332.5 ;
      RECT  7577.5 88197.5 7642.5 88332.5 ;
      RECT  7577.5 88197.5 7642.5 88332.5 ;
      RECT  7387.5 88197.5 7452.5 88332.5 ;
      RECT  7577.5 88197.5 7642.5 88332.5 ;
      RECT  7767.5 88197.5 7832.5 88332.5 ;
      RECT  7767.5 88197.5 7832.5 88332.5 ;
      RECT  7577.5 88197.5 7642.5 88332.5 ;
      RECT  7197.5 87357.5 7262.5 87492.5 ;
      RECT  7387.5 87357.5 7452.5 87492.5 ;
      RECT  7387.5 87357.5 7452.5 87492.5 ;
      RECT  7197.5 87357.5 7262.5 87492.5 ;
      RECT  7387.5 87357.5 7452.5 87492.5 ;
      RECT  7577.5 87357.5 7642.5 87492.5 ;
      RECT  7577.5 87357.5 7642.5 87492.5 ;
      RECT  7387.5 87357.5 7452.5 87492.5 ;
      RECT  7577.5 87357.5 7642.5 87492.5 ;
      RECT  7767.5 87357.5 7832.5 87492.5 ;
      RECT  7767.5 87357.5 7832.5 87492.5 ;
      RECT  7577.5 87357.5 7642.5 87492.5 ;
      RECT  7937.5 88287.5 8002.5 88422.5 ;
      RECT  7937.5 87312.5 8002.5 87447.5 ;
      RECT  7772.5 87570.0 7637.5 87635.0 ;
      RECT  7582.5 87710.0 7447.5 87775.0 ;
      RECT  7392.5 87850.0 7257.5 87915.0 ;
      RECT  7387.5 88197.5 7452.5 88332.5 ;
      RECT  7767.5 88197.5 7832.5 88332.5 ;
      RECT  7767.5 87357.5 7832.5 87492.5 ;
      RECT  7767.5 87815.0 7832.5 87950.0 ;
      RECT  7257.5 87850.0 7392.5 87915.0 ;
      RECT  7447.5 87710.0 7582.5 87775.0 ;
      RECT  7637.5 87570.0 7772.5 87635.0 ;
      RECT  7767.5 87815.0 7832.5 87950.0 ;
      RECT  7130.0 88507.5 8140.0 88572.5 ;
      RECT  7130.0 87162.5 8140.0 87227.5 ;
      RECT  7197.5 89722.5 7262.5 89917.5 ;
      RECT  7197.5 88882.5 7262.5 88507.5 ;
      RECT  7577.5 88882.5 7642.5 88507.5 ;
      RECT  7937.5 88725.0 8002.5 88540.0 ;
      RECT  7937.5 89885.0 8002.5 89700.0 ;
      RECT  7197.5 88882.5 7262.5 88747.5 ;
      RECT  7387.5 88882.5 7452.5 88747.5 ;
      RECT  7387.5 88882.5 7452.5 88747.5 ;
      RECT  7197.5 88882.5 7262.5 88747.5 ;
      RECT  7387.5 88882.5 7452.5 88747.5 ;
      RECT  7577.5 88882.5 7642.5 88747.5 ;
      RECT  7577.5 88882.5 7642.5 88747.5 ;
      RECT  7387.5 88882.5 7452.5 88747.5 ;
      RECT  7577.5 88882.5 7642.5 88747.5 ;
      RECT  7767.5 88882.5 7832.5 88747.5 ;
      RECT  7767.5 88882.5 7832.5 88747.5 ;
      RECT  7577.5 88882.5 7642.5 88747.5 ;
      RECT  7197.5 89722.5 7262.5 89587.5 ;
      RECT  7387.5 89722.5 7452.5 89587.5 ;
      RECT  7387.5 89722.5 7452.5 89587.5 ;
      RECT  7197.5 89722.5 7262.5 89587.5 ;
      RECT  7387.5 89722.5 7452.5 89587.5 ;
      RECT  7577.5 89722.5 7642.5 89587.5 ;
      RECT  7577.5 89722.5 7642.5 89587.5 ;
      RECT  7387.5 89722.5 7452.5 89587.5 ;
      RECT  7577.5 89722.5 7642.5 89587.5 ;
      RECT  7767.5 89722.5 7832.5 89587.5 ;
      RECT  7767.5 89722.5 7832.5 89587.5 ;
      RECT  7577.5 89722.5 7642.5 89587.5 ;
      RECT  7937.5 88792.5 8002.5 88657.5 ;
      RECT  7937.5 89767.5 8002.5 89632.5 ;
      RECT  7772.5 89510.0 7637.5 89445.0 ;
      RECT  7582.5 89370.0 7447.5 89305.0 ;
      RECT  7392.5 89230.0 7257.5 89165.0 ;
      RECT  7387.5 88882.5 7452.5 88747.5 ;
      RECT  7767.5 88882.5 7832.5 88747.5 ;
      RECT  7767.5 89722.5 7832.5 89587.5 ;
      RECT  7767.5 89265.0 7832.5 89130.0 ;
      RECT  7257.5 89230.0 7392.5 89165.0 ;
      RECT  7447.5 89370.0 7582.5 89305.0 ;
      RECT  7637.5 89510.0 7772.5 89445.0 ;
      RECT  7767.5 89265.0 7832.5 89130.0 ;
      RECT  7130.0 88572.5 8140.0 88507.5 ;
      RECT  7130.0 89917.5 8140.0 89852.5 ;
      RECT  7197.5 90047.5 7262.5 89852.5 ;
      RECT  7197.5 90887.5 7262.5 91262.5 ;
      RECT  7577.5 90887.5 7642.5 91262.5 ;
      RECT  7937.5 91045.0 8002.5 91230.0 ;
      RECT  7937.5 89885.0 8002.5 90070.0 ;
      RECT  7197.5 90887.5 7262.5 91022.5 ;
      RECT  7387.5 90887.5 7452.5 91022.5 ;
      RECT  7387.5 90887.5 7452.5 91022.5 ;
      RECT  7197.5 90887.5 7262.5 91022.5 ;
      RECT  7387.5 90887.5 7452.5 91022.5 ;
      RECT  7577.5 90887.5 7642.5 91022.5 ;
      RECT  7577.5 90887.5 7642.5 91022.5 ;
      RECT  7387.5 90887.5 7452.5 91022.5 ;
      RECT  7577.5 90887.5 7642.5 91022.5 ;
      RECT  7767.5 90887.5 7832.5 91022.5 ;
      RECT  7767.5 90887.5 7832.5 91022.5 ;
      RECT  7577.5 90887.5 7642.5 91022.5 ;
      RECT  7197.5 90047.5 7262.5 90182.5 ;
      RECT  7387.5 90047.5 7452.5 90182.5 ;
      RECT  7387.5 90047.5 7452.5 90182.5 ;
      RECT  7197.5 90047.5 7262.5 90182.5 ;
      RECT  7387.5 90047.5 7452.5 90182.5 ;
      RECT  7577.5 90047.5 7642.5 90182.5 ;
      RECT  7577.5 90047.5 7642.5 90182.5 ;
      RECT  7387.5 90047.5 7452.5 90182.5 ;
      RECT  7577.5 90047.5 7642.5 90182.5 ;
      RECT  7767.5 90047.5 7832.5 90182.5 ;
      RECT  7767.5 90047.5 7832.5 90182.5 ;
      RECT  7577.5 90047.5 7642.5 90182.5 ;
      RECT  7937.5 90977.5 8002.5 91112.5 ;
      RECT  7937.5 90002.5 8002.5 90137.5 ;
      RECT  7772.5 90260.0 7637.5 90325.0 ;
      RECT  7582.5 90400.0 7447.5 90465.0 ;
      RECT  7392.5 90540.0 7257.5 90605.0 ;
      RECT  7387.5 90887.5 7452.5 91022.5 ;
      RECT  7767.5 90887.5 7832.5 91022.5 ;
      RECT  7767.5 90047.5 7832.5 90182.5 ;
      RECT  7767.5 90505.0 7832.5 90640.0 ;
      RECT  7257.5 90540.0 7392.5 90605.0 ;
      RECT  7447.5 90400.0 7582.5 90465.0 ;
      RECT  7637.5 90260.0 7772.5 90325.0 ;
      RECT  7767.5 90505.0 7832.5 90640.0 ;
      RECT  7130.0 91197.5 8140.0 91262.5 ;
      RECT  7130.0 89852.5 8140.0 89917.5 ;
      RECT  7197.5 92412.5 7262.5 92607.5 ;
      RECT  7197.5 91572.5 7262.5 91197.5 ;
      RECT  7577.5 91572.5 7642.5 91197.5 ;
      RECT  7937.5 91415.0 8002.5 91230.0 ;
      RECT  7937.5 92575.0 8002.5 92390.0 ;
      RECT  7197.5 91572.5 7262.5 91437.5 ;
      RECT  7387.5 91572.5 7452.5 91437.5 ;
      RECT  7387.5 91572.5 7452.5 91437.5 ;
      RECT  7197.5 91572.5 7262.5 91437.5 ;
      RECT  7387.5 91572.5 7452.5 91437.5 ;
      RECT  7577.5 91572.5 7642.5 91437.5 ;
      RECT  7577.5 91572.5 7642.5 91437.5 ;
      RECT  7387.5 91572.5 7452.5 91437.5 ;
      RECT  7577.5 91572.5 7642.5 91437.5 ;
      RECT  7767.5 91572.5 7832.5 91437.5 ;
      RECT  7767.5 91572.5 7832.5 91437.5 ;
      RECT  7577.5 91572.5 7642.5 91437.5 ;
      RECT  7197.5 92412.5 7262.5 92277.5 ;
      RECT  7387.5 92412.5 7452.5 92277.5 ;
      RECT  7387.5 92412.5 7452.5 92277.5 ;
      RECT  7197.5 92412.5 7262.5 92277.5 ;
      RECT  7387.5 92412.5 7452.5 92277.5 ;
      RECT  7577.5 92412.5 7642.5 92277.5 ;
      RECT  7577.5 92412.5 7642.5 92277.5 ;
      RECT  7387.5 92412.5 7452.5 92277.5 ;
      RECT  7577.5 92412.5 7642.5 92277.5 ;
      RECT  7767.5 92412.5 7832.5 92277.5 ;
      RECT  7767.5 92412.5 7832.5 92277.5 ;
      RECT  7577.5 92412.5 7642.5 92277.5 ;
      RECT  7937.5 91482.5 8002.5 91347.5 ;
      RECT  7937.5 92457.5 8002.5 92322.5 ;
      RECT  7772.5 92200.0 7637.5 92135.0 ;
      RECT  7582.5 92060.0 7447.5 91995.0 ;
      RECT  7392.5 91920.0 7257.5 91855.0 ;
      RECT  7387.5 91572.5 7452.5 91437.5 ;
      RECT  7767.5 91572.5 7832.5 91437.5 ;
      RECT  7767.5 92412.5 7832.5 92277.5 ;
      RECT  7767.5 91955.0 7832.5 91820.0 ;
      RECT  7257.5 91920.0 7392.5 91855.0 ;
      RECT  7447.5 92060.0 7582.5 91995.0 ;
      RECT  7637.5 92200.0 7772.5 92135.0 ;
      RECT  7767.5 91955.0 7832.5 91820.0 ;
      RECT  7130.0 91262.5 8140.0 91197.5 ;
      RECT  7130.0 92607.5 8140.0 92542.5 ;
      RECT  7197.5 92737.5 7262.5 92542.5 ;
      RECT  7197.5 93577.5 7262.5 93952.5 ;
      RECT  7577.5 93577.5 7642.5 93952.5 ;
      RECT  7937.5 93735.0 8002.5 93920.0 ;
      RECT  7937.5 92575.0 8002.5 92760.0 ;
      RECT  7197.5 93577.5 7262.5 93712.5 ;
      RECT  7387.5 93577.5 7452.5 93712.5 ;
      RECT  7387.5 93577.5 7452.5 93712.5 ;
      RECT  7197.5 93577.5 7262.5 93712.5 ;
      RECT  7387.5 93577.5 7452.5 93712.5 ;
      RECT  7577.5 93577.5 7642.5 93712.5 ;
      RECT  7577.5 93577.5 7642.5 93712.5 ;
      RECT  7387.5 93577.5 7452.5 93712.5 ;
      RECT  7577.5 93577.5 7642.5 93712.5 ;
      RECT  7767.5 93577.5 7832.5 93712.5 ;
      RECT  7767.5 93577.5 7832.5 93712.5 ;
      RECT  7577.5 93577.5 7642.5 93712.5 ;
      RECT  7197.5 92737.5 7262.5 92872.5 ;
      RECT  7387.5 92737.5 7452.5 92872.5 ;
      RECT  7387.5 92737.5 7452.5 92872.5 ;
      RECT  7197.5 92737.5 7262.5 92872.5 ;
      RECT  7387.5 92737.5 7452.5 92872.5 ;
      RECT  7577.5 92737.5 7642.5 92872.5 ;
      RECT  7577.5 92737.5 7642.5 92872.5 ;
      RECT  7387.5 92737.5 7452.5 92872.5 ;
      RECT  7577.5 92737.5 7642.5 92872.5 ;
      RECT  7767.5 92737.5 7832.5 92872.5 ;
      RECT  7767.5 92737.5 7832.5 92872.5 ;
      RECT  7577.5 92737.5 7642.5 92872.5 ;
      RECT  7937.5 93667.5 8002.5 93802.5 ;
      RECT  7937.5 92692.5 8002.5 92827.5 ;
      RECT  7772.5 92950.0 7637.5 93015.0 ;
      RECT  7582.5 93090.0 7447.5 93155.0 ;
      RECT  7392.5 93230.0 7257.5 93295.0 ;
      RECT  7387.5 93577.5 7452.5 93712.5 ;
      RECT  7767.5 93577.5 7832.5 93712.5 ;
      RECT  7767.5 92737.5 7832.5 92872.5 ;
      RECT  7767.5 93195.0 7832.5 93330.0 ;
      RECT  7257.5 93230.0 7392.5 93295.0 ;
      RECT  7447.5 93090.0 7582.5 93155.0 ;
      RECT  7637.5 92950.0 7772.5 93015.0 ;
      RECT  7767.5 93195.0 7832.5 93330.0 ;
      RECT  7130.0 93887.5 8140.0 93952.5 ;
      RECT  7130.0 92542.5 8140.0 92607.5 ;
      RECT  7197.5 95102.5 7262.5 95297.5 ;
      RECT  7197.5 94262.5 7262.5 93887.5 ;
      RECT  7577.5 94262.5 7642.5 93887.5 ;
      RECT  7937.5 94105.0 8002.5 93920.0 ;
      RECT  7937.5 95265.0 8002.5 95080.0 ;
      RECT  7197.5 94262.5 7262.5 94127.5 ;
      RECT  7387.5 94262.5 7452.5 94127.5 ;
      RECT  7387.5 94262.5 7452.5 94127.5 ;
      RECT  7197.5 94262.5 7262.5 94127.5 ;
      RECT  7387.5 94262.5 7452.5 94127.5 ;
      RECT  7577.5 94262.5 7642.5 94127.5 ;
      RECT  7577.5 94262.5 7642.5 94127.5 ;
      RECT  7387.5 94262.5 7452.5 94127.5 ;
      RECT  7577.5 94262.5 7642.5 94127.5 ;
      RECT  7767.5 94262.5 7832.5 94127.5 ;
      RECT  7767.5 94262.5 7832.5 94127.5 ;
      RECT  7577.5 94262.5 7642.5 94127.5 ;
      RECT  7197.5 95102.5 7262.5 94967.5 ;
      RECT  7387.5 95102.5 7452.5 94967.5 ;
      RECT  7387.5 95102.5 7452.5 94967.5 ;
      RECT  7197.5 95102.5 7262.5 94967.5 ;
      RECT  7387.5 95102.5 7452.5 94967.5 ;
      RECT  7577.5 95102.5 7642.5 94967.5 ;
      RECT  7577.5 95102.5 7642.5 94967.5 ;
      RECT  7387.5 95102.5 7452.5 94967.5 ;
      RECT  7577.5 95102.5 7642.5 94967.5 ;
      RECT  7767.5 95102.5 7832.5 94967.5 ;
      RECT  7767.5 95102.5 7832.5 94967.5 ;
      RECT  7577.5 95102.5 7642.5 94967.5 ;
      RECT  7937.5 94172.5 8002.5 94037.5 ;
      RECT  7937.5 95147.5 8002.5 95012.5 ;
      RECT  7772.5 94890.0 7637.5 94825.0 ;
      RECT  7582.5 94750.0 7447.5 94685.0 ;
      RECT  7392.5 94610.0 7257.5 94545.0 ;
      RECT  7387.5 94262.5 7452.5 94127.5 ;
      RECT  7767.5 94262.5 7832.5 94127.5 ;
      RECT  7767.5 95102.5 7832.5 94967.5 ;
      RECT  7767.5 94645.0 7832.5 94510.0 ;
      RECT  7257.5 94610.0 7392.5 94545.0 ;
      RECT  7447.5 94750.0 7582.5 94685.0 ;
      RECT  7637.5 94890.0 7772.5 94825.0 ;
      RECT  7767.5 94645.0 7832.5 94510.0 ;
      RECT  7130.0 93952.5 8140.0 93887.5 ;
      RECT  7130.0 95297.5 8140.0 95232.5 ;
      RECT  7197.5 95427.5 7262.5 95232.5 ;
      RECT  7197.5 96267.5 7262.5 96642.5 ;
      RECT  7577.5 96267.5 7642.5 96642.5 ;
      RECT  7937.5 96425.0 8002.5 96610.0 ;
      RECT  7937.5 95265.0 8002.5 95450.0 ;
      RECT  7197.5 96267.5 7262.5 96402.5 ;
      RECT  7387.5 96267.5 7452.5 96402.5 ;
      RECT  7387.5 96267.5 7452.5 96402.5 ;
      RECT  7197.5 96267.5 7262.5 96402.5 ;
      RECT  7387.5 96267.5 7452.5 96402.5 ;
      RECT  7577.5 96267.5 7642.5 96402.5 ;
      RECT  7577.5 96267.5 7642.5 96402.5 ;
      RECT  7387.5 96267.5 7452.5 96402.5 ;
      RECT  7577.5 96267.5 7642.5 96402.5 ;
      RECT  7767.5 96267.5 7832.5 96402.5 ;
      RECT  7767.5 96267.5 7832.5 96402.5 ;
      RECT  7577.5 96267.5 7642.5 96402.5 ;
      RECT  7197.5 95427.5 7262.5 95562.5 ;
      RECT  7387.5 95427.5 7452.5 95562.5 ;
      RECT  7387.5 95427.5 7452.5 95562.5 ;
      RECT  7197.5 95427.5 7262.5 95562.5 ;
      RECT  7387.5 95427.5 7452.5 95562.5 ;
      RECT  7577.5 95427.5 7642.5 95562.5 ;
      RECT  7577.5 95427.5 7642.5 95562.5 ;
      RECT  7387.5 95427.5 7452.5 95562.5 ;
      RECT  7577.5 95427.5 7642.5 95562.5 ;
      RECT  7767.5 95427.5 7832.5 95562.5 ;
      RECT  7767.5 95427.5 7832.5 95562.5 ;
      RECT  7577.5 95427.5 7642.5 95562.5 ;
      RECT  7937.5 96357.5 8002.5 96492.5 ;
      RECT  7937.5 95382.5 8002.5 95517.5 ;
      RECT  7772.5 95640.0 7637.5 95705.0 ;
      RECT  7582.5 95780.0 7447.5 95845.0 ;
      RECT  7392.5 95920.0 7257.5 95985.0 ;
      RECT  7387.5 96267.5 7452.5 96402.5 ;
      RECT  7767.5 96267.5 7832.5 96402.5 ;
      RECT  7767.5 95427.5 7832.5 95562.5 ;
      RECT  7767.5 95885.0 7832.5 96020.0 ;
      RECT  7257.5 95920.0 7392.5 95985.0 ;
      RECT  7447.5 95780.0 7582.5 95845.0 ;
      RECT  7637.5 95640.0 7772.5 95705.0 ;
      RECT  7767.5 95885.0 7832.5 96020.0 ;
      RECT  7130.0 96577.5 8140.0 96642.5 ;
      RECT  7130.0 95232.5 8140.0 95297.5 ;
      RECT  7197.5 97792.5 7262.5 97987.5 ;
      RECT  7197.5 96952.5 7262.5 96577.5 ;
      RECT  7577.5 96952.5 7642.5 96577.5 ;
      RECT  7937.5 96795.0 8002.5 96610.0 ;
      RECT  7937.5 97955.0 8002.5 97770.0 ;
      RECT  7197.5 96952.5 7262.5 96817.5 ;
      RECT  7387.5 96952.5 7452.5 96817.5 ;
      RECT  7387.5 96952.5 7452.5 96817.5 ;
      RECT  7197.5 96952.5 7262.5 96817.5 ;
      RECT  7387.5 96952.5 7452.5 96817.5 ;
      RECT  7577.5 96952.5 7642.5 96817.5 ;
      RECT  7577.5 96952.5 7642.5 96817.5 ;
      RECT  7387.5 96952.5 7452.5 96817.5 ;
      RECT  7577.5 96952.5 7642.5 96817.5 ;
      RECT  7767.5 96952.5 7832.5 96817.5 ;
      RECT  7767.5 96952.5 7832.5 96817.5 ;
      RECT  7577.5 96952.5 7642.5 96817.5 ;
      RECT  7197.5 97792.5 7262.5 97657.5 ;
      RECT  7387.5 97792.5 7452.5 97657.5 ;
      RECT  7387.5 97792.5 7452.5 97657.5 ;
      RECT  7197.5 97792.5 7262.5 97657.5 ;
      RECT  7387.5 97792.5 7452.5 97657.5 ;
      RECT  7577.5 97792.5 7642.5 97657.5 ;
      RECT  7577.5 97792.5 7642.5 97657.5 ;
      RECT  7387.5 97792.5 7452.5 97657.5 ;
      RECT  7577.5 97792.5 7642.5 97657.5 ;
      RECT  7767.5 97792.5 7832.5 97657.5 ;
      RECT  7767.5 97792.5 7832.5 97657.5 ;
      RECT  7577.5 97792.5 7642.5 97657.5 ;
      RECT  7937.5 96862.5 8002.5 96727.5 ;
      RECT  7937.5 97837.5 8002.5 97702.5 ;
      RECT  7772.5 97580.0 7637.5 97515.0 ;
      RECT  7582.5 97440.0 7447.5 97375.0 ;
      RECT  7392.5 97300.0 7257.5 97235.0 ;
      RECT  7387.5 96952.5 7452.5 96817.5 ;
      RECT  7767.5 96952.5 7832.5 96817.5 ;
      RECT  7767.5 97792.5 7832.5 97657.5 ;
      RECT  7767.5 97335.0 7832.5 97200.0 ;
      RECT  7257.5 97300.0 7392.5 97235.0 ;
      RECT  7447.5 97440.0 7582.5 97375.0 ;
      RECT  7637.5 97580.0 7772.5 97515.0 ;
      RECT  7767.5 97335.0 7832.5 97200.0 ;
      RECT  7130.0 96642.5 8140.0 96577.5 ;
      RECT  7130.0 97987.5 8140.0 97922.5 ;
      RECT  7197.5 98117.5 7262.5 97922.5 ;
      RECT  7197.5 98957.5 7262.5 99332.5 ;
      RECT  7577.5 98957.5 7642.5 99332.5 ;
      RECT  7937.5 99115.0 8002.5 99300.0 ;
      RECT  7937.5 97955.0 8002.5 98140.0 ;
      RECT  7197.5 98957.5 7262.5 99092.5 ;
      RECT  7387.5 98957.5 7452.5 99092.5 ;
      RECT  7387.5 98957.5 7452.5 99092.5 ;
      RECT  7197.5 98957.5 7262.5 99092.5 ;
      RECT  7387.5 98957.5 7452.5 99092.5 ;
      RECT  7577.5 98957.5 7642.5 99092.5 ;
      RECT  7577.5 98957.5 7642.5 99092.5 ;
      RECT  7387.5 98957.5 7452.5 99092.5 ;
      RECT  7577.5 98957.5 7642.5 99092.5 ;
      RECT  7767.5 98957.5 7832.5 99092.5 ;
      RECT  7767.5 98957.5 7832.5 99092.5 ;
      RECT  7577.5 98957.5 7642.5 99092.5 ;
      RECT  7197.5 98117.5 7262.5 98252.5 ;
      RECT  7387.5 98117.5 7452.5 98252.5 ;
      RECT  7387.5 98117.5 7452.5 98252.5 ;
      RECT  7197.5 98117.5 7262.5 98252.5 ;
      RECT  7387.5 98117.5 7452.5 98252.5 ;
      RECT  7577.5 98117.5 7642.5 98252.5 ;
      RECT  7577.5 98117.5 7642.5 98252.5 ;
      RECT  7387.5 98117.5 7452.5 98252.5 ;
      RECT  7577.5 98117.5 7642.5 98252.5 ;
      RECT  7767.5 98117.5 7832.5 98252.5 ;
      RECT  7767.5 98117.5 7832.5 98252.5 ;
      RECT  7577.5 98117.5 7642.5 98252.5 ;
      RECT  7937.5 99047.5 8002.5 99182.5 ;
      RECT  7937.5 98072.5 8002.5 98207.5 ;
      RECT  7772.5 98330.0 7637.5 98395.0 ;
      RECT  7582.5 98470.0 7447.5 98535.0 ;
      RECT  7392.5 98610.0 7257.5 98675.0 ;
      RECT  7387.5 98957.5 7452.5 99092.5 ;
      RECT  7767.5 98957.5 7832.5 99092.5 ;
      RECT  7767.5 98117.5 7832.5 98252.5 ;
      RECT  7767.5 98575.0 7832.5 98710.0 ;
      RECT  7257.5 98610.0 7392.5 98675.0 ;
      RECT  7447.5 98470.0 7582.5 98535.0 ;
      RECT  7637.5 98330.0 7772.5 98395.0 ;
      RECT  7767.5 98575.0 7832.5 98710.0 ;
      RECT  7130.0 99267.5 8140.0 99332.5 ;
      RECT  7130.0 97922.5 8140.0 97987.5 ;
      RECT  7197.5 100482.5 7262.5 100677.5 ;
      RECT  7197.5 99642.5 7262.5 99267.5 ;
      RECT  7577.5 99642.5 7642.5 99267.5 ;
      RECT  7937.5 99485.0 8002.5 99300.0 ;
      RECT  7937.5 100645.0 8002.5 100460.0 ;
      RECT  7197.5 99642.5 7262.5 99507.5 ;
      RECT  7387.5 99642.5 7452.5 99507.5 ;
      RECT  7387.5 99642.5 7452.5 99507.5 ;
      RECT  7197.5 99642.5 7262.5 99507.5 ;
      RECT  7387.5 99642.5 7452.5 99507.5 ;
      RECT  7577.5 99642.5 7642.5 99507.5 ;
      RECT  7577.5 99642.5 7642.5 99507.5 ;
      RECT  7387.5 99642.5 7452.5 99507.5 ;
      RECT  7577.5 99642.5 7642.5 99507.5 ;
      RECT  7767.5 99642.5 7832.5 99507.5 ;
      RECT  7767.5 99642.5 7832.5 99507.5 ;
      RECT  7577.5 99642.5 7642.5 99507.5 ;
      RECT  7197.5 100482.5 7262.5 100347.5 ;
      RECT  7387.5 100482.5 7452.5 100347.5 ;
      RECT  7387.5 100482.5 7452.5 100347.5 ;
      RECT  7197.5 100482.5 7262.5 100347.5 ;
      RECT  7387.5 100482.5 7452.5 100347.5 ;
      RECT  7577.5 100482.5 7642.5 100347.5 ;
      RECT  7577.5 100482.5 7642.5 100347.5 ;
      RECT  7387.5 100482.5 7452.5 100347.5 ;
      RECT  7577.5 100482.5 7642.5 100347.5 ;
      RECT  7767.5 100482.5 7832.5 100347.5 ;
      RECT  7767.5 100482.5 7832.5 100347.5 ;
      RECT  7577.5 100482.5 7642.5 100347.5 ;
      RECT  7937.5 99552.5 8002.5 99417.5 ;
      RECT  7937.5 100527.5 8002.5 100392.5 ;
      RECT  7772.5 100270.0 7637.5 100205.0 ;
      RECT  7582.5 100130.0 7447.5 100065.0 ;
      RECT  7392.5 99990.0 7257.5 99925.0 ;
      RECT  7387.5 99642.5 7452.5 99507.5 ;
      RECT  7767.5 99642.5 7832.5 99507.5 ;
      RECT  7767.5 100482.5 7832.5 100347.5 ;
      RECT  7767.5 100025.0 7832.5 99890.0 ;
      RECT  7257.5 99990.0 7392.5 99925.0 ;
      RECT  7447.5 100130.0 7582.5 100065.0 ;
      RECT  7637.5 100270.0 7772.5 100205.0 ;
      RECT  7767.5 100025.0 7832.5 99890.0 ;
      RECT  7130.0 99332.5 8140.0 99267.5 ;
      RECT  7130.0 100677.5 8140.0 100612.5 ;
      RECT  7197.5 100807.5 7262.5 100612.5 ;
      RECT  7197.5 101647.5 7262.5 102022.5 ;
      RECT  7577.5 101647.5 7642.5 102022.5 ;
      RECT  7937.5 101805.0 8002.5 101990.0 ;
      RECT  7937.5 100645.0 8002.5 100830.0 ;
      RECT  7197.5 101647.5 7262.5 101782.5 ;
      RECT  7387.5 101647.5 7452.5 101782.5 ;
      RECT  7387.5 101647.5 7452.5 101782.5 ;
      RECT  7197.5 101647.5 7262.5 101782.5 ;
      RECT  7387.5 101647.5 7452.5 101782.5 ;
      RECT  7577.5 101647.5 7642.5 101782.5 ;
      RECT  7577.5 101647.5 7642.5 101782.5 ;
      RECT  7387.5 101647.5 7452.5 101782.5 ;
      RECT  7577.5 101647.5 7642.5 101782.5 ;
      RECT  7767.5 101647.5 7832.5 101782.5 ;
      RECT  7767.5 101647.5 7832.5 101782.5 ;
      RECT  7577.5 101647.5 7642.5 101782.5 ;
      RECT  7197.5 100807.5 7262.5 100942.5 ;
      RECT  7387.5 100807.5 7452.5 100942.5 ;
      RECT  7387.5 100807.5 7452.5 100942.5 ;
      RECT  7197.5 100807.5 7262.5 100942.5 ;
      RECT  7387.5 100807.5 7452.5 100942.5 ;
      RECT  7577.5 100807.5 7642.5 100942.5 ;
      RECT  7577.5 100807.5 7642.5 100942.5 ;
      RECT  7387.5 100807.5 7452.5 100942.5 ;
      RECT  7577.5 100807.5 7642.5 100942.5 ;
      RECT  7767.5 100807.5 7832.5 100942.5 ;
      RECT  7767.5 100807.5 7832.5 100942.5 ;
      RECT  7577.5 100807.5 7642.5 100942.5 ;
      RECT  7937.5 101737.5 8002.5 101872.5 ;
      RECT  7937.5 100762.5 8002.5 100897.5 ;
      RECT  7772.5 101020.0 7637.5 101085.0 ;
      RECT  7582.5 101160.0 7447.5 101225.0 ;
      RECT  7392.5 101300.0 7257.5 101365.0 ;
      RECT  7387.5 101647.5 7452.5 101782.5 ;
      RECT  7767.5 101647.5 7832.5 101782.5 ;
      RECT  7767.5 100807.5 7832.5 100942.5 ;
      RECT  7767.5 101265.0 7832.5 101400.0 ;
      RECT  7257.5 101300.0 7392.5 101365.0 ;
      RECT  7447.5 101160.0 7582.5 101225.0 ;
      RECT  7637.5 101020.0 7772.5 101085.0 ;
      RECT  7767.5 101265.0 7832.5 101400.0 ;
      RECT  7130.0 101957.5 8140.0 102022.5 ;
      RECT  7130.0 100612.5 8140.0 100677.5 ;
      RECT  7197.5 103172.5 7262.5 103367.5 ;
      RECT  7197.5 102332.5 7262.5 101957.5 ;
      RECT  7577.5 102332.5 7642.5 101957.5 ;
      RECT  7937.5 102175.0 8002.5 101990.0 ;
      RECT  7937.5 103335.0 8002.5 103150.0 ;
      RECT  7197.5 102332.5 7262.5 102197.5 ;
      RECT  7387.5 102332.5 7452.5 102197.5 ;
      RECT  7387.5 102332.5 7452.5 102197.5 ;
      RECT  7197.5 102332.5 7262.5 102197.5 ;
      RECT  7387.5 102332.5 7452.5 102197.5 ;
      RECT  7577.5 102332.5 7642.5 102197.5 ;
      RECT  7577.5 102332.5 7642.5 102197.5 ;
      RECT  7387.5 102332.5 7452.5 102197.5 ;
      RECT  7577.5 102332.5 7642.5 102197.5 ;
      RECT  7767.5 102332.5 7832.5 102197.5 ;
      RECT  7767.5 102332.5 7832.5 102197.5 ;
      RECT  7577.5 102332.5 7642.5 102197.5 ;
      RECT  7197.5 103172.5 7262.5 103037.5 ;
      RECT  7387.5 103172.5 7452.5 103037.5 ;
      RECT  7387.5 103172.5 7452.5 103037.5 ;
      RECT  7197.5 103172.5 7262.5 103037.5 ;
      RECT  7387.5 103172.5 7452.5 103037.5 ;
      RECT  7577.5 103172.5 7642.5 103037.5 ;
      RECT  7577.5 103172.5 7642.5 103037.5 ;
      RECT  7387.5 103172.5 7452.5 103037.5 ;
      RECT  7577.5 103172.5 7642.5 103037.5 ;
      RECT  7767.5 103172.5 7832.5 103037.5 ;
      RECT  7767.5 103172.5 7832.5 103037.5 ;
      RECT  7577.5 103172.5 7642.5 103037.5 ;
      RECT  7937.5 102242.5 8002.5 102107.5 ;
      RECT  7937.5 103217.5 8002.5 103082.5 ;
      RECT  7772.5 102960.0 7637.5 102895.0 ;
      RECT  7582.5 102820.0 7447.5 102755.0 ;
      RECT  7392.5 102680.0 7257.5 102615.0 ;
      RECT  7387.5 102332.5 7452.5 102197.5 ;
      RECT  7767.5 102332.5 7832.5 102197.5 ;
      RECT  7767.5 103172.5 7832.5 103037.5 ;
      RECT  7767.5 102715.0 7832.5 102580.0 ;
      RECT  7257.5 102680.0 7392.5 102615.0 ;
      RECT  7447.5 102820.0 7582.5 102755.0 ;
      RECT  7637.5 102960.0 7772.5 102895.0 ;
      RECT  7767.5 102715.0 7832.5 102580.0 ;
      RECT  7130.0 102022.5 8140.0 101957.5 ;
      RECT  7130.0 103367.5 8140.0 103302.5 ;
      RECT  7197.5 103497.5 7262.5 103302.5 ;
      RECT  7197.5 104337.5 7262.5 104712.5 ;
      RECT  7577.5 104337.5 7642.5 104712.5 ;
      RECT  7937.5 104495.0 8002.5 104680.0 ;
      RECT  7937.5 103335.0 8002.5 103520.0 ;
      RECT  7197.5 104337.5 7262.5 104472.5 ;
      RECT  7387.5 104337.5 7452.5 104472.5 ;
      RECT  7387.5 104337.5 7452.5 104472.5 ;
      RECT  7197.5 104337.5 7262.5 104472.5 ;
      RECT  7387.5 104337.5 7452.5 104472.5 ;
      RECT  7577.5 104337.5 7642.5 104472.5 ;
      RECT  7577.5 104337.5 7642.5 104472.5 ;
      RECT  7387.5 104337.5 7452.5 104472.5 ;
      RECT  7577.5 104337.5 7642.5 104472.5 ;
      RECT  7767.5 104337.5 7832.5 104472.5 ;
      RECT  7767.5 104337.5 7832.5 104472.5 ;
      RECT  7577.5 104337.5 7642.5 104472.5 ;
      RECT  7197.5 103497.5 7262.5 103632.5 ;
      RECT  7387.5 103497.5 7452.5 103632.5 ;
      RECT  7387.5 103497.5 7452.5 103632.5 ;
      RECT  7197.5 103497.5 7262.5 103632.5 ;
      RECT  7387.5 103497.5 7452.5 103632.5 ;
      RECT  7577.5 103497.5 7642.5 103632.5 ;
      RECT  7577.5 103497.5 7642.5 103632.5 ;
      RECT  7387.5 103497.5 7452.5 103632.5 ;
      RECT  7577.5 103497.5 7642.5 103632.5 ;
      RECT  7767.5 103497.5 7832.5 103632.5 ;
      RECT  7767.5 103497.5 7832.5 103632.5 ;
      RECT  7577.5 103497.5 7642.5 103632.5 ;
      RECT  7937.5 104427.5 8002.5 104562.5 ;
      RECT  7937.5 103452.5 8002.5 103587.5 ;
      RECT  7772.5 103710.0 7637.5 103775.0 ;
      RECT  7582.5 103850.0 7447.5 103915.0 ;
      RECT  7392.5 103990.0 7257.5 104055.0 ;
      RECT  7387.5 104337.5 7452.5 104472.5 ;
      RECT  7767.5 104337.5 7832.5 104472.5 ;
      RECT  7767.5 103497.5 7832.5 103632.5 ;
      RECT  7767.5 103955.0 7832.5 104090.0 ;
      RECT  7257.5 103990.0 7392.5 104055.0 ;
      RECT  7447.5 103850.0 7582.5 103915.0 ;
      RECT  7637.5 103710.0 7772.5 103775.0 ;
      RECT  7767.5 103955.0 7832.5 104090.0 ;
      RECT  7130.0 104647.5 8140.0 104712.5 ;
      RECT  7130.0 103302.5 8140.0 103367.5 ;
      RECT  7197.5 105862.5 7262.5 106057.5 ;
      RECT  7197.5 105022.5 7262.5 104647.5 ;
      RECT  7577.5 105022.5 7642.5 104647.5 ;
      RECT  7937.5 104865.0 8002.5 104680.0 ;
      RECT  7937.5 106025.0 8002.5 105840.0 ;
      RECT  7197.5 105022.5 7262.5 104887.5 ;
      RECT  7387.5 105022.5 7452.5 104887.5 ;
      RECT  7387.5 105022.5 7452.5 104887.5 ;
      RECT  7197.5 105022.5 7262.5 104887.5 ;
      RECT  7387.5 105022.5 7452.5 104887.5 ;
      RECT  7577.5 105022.5 7642.5 104887.5 ;
      RECT  7577.5 105022.5 7642.5 104887.5 ;
      RECT  7387.5 105022.5 7452.5 104887.5 ;
      RECT  7577.5 105022.5 7642.5 104887.5 ;
      RECT  7767.5 105022.5 7832.5 104887.5 ;
      RECT  7767.5 105022.5 7832.5 104887.5 ;
      RECT  7577.5 105022.5 7642.5 104887.5 ;
      RECT  7197.5 105862.5 7262.5 105727.5 ;
      RECT  7387.5 105862.5 7452.5 105727.5 ;
      RECT  7387.5 105862.5 7452.5 105727.5 ;
      RECT  7197.5 105862.5 7262.5 105727.5 ;
      RECT  7387.5 105862.5 7452.5 105727.5 ;
      RECT  7577.5 105862.5 7642.5 105727.5 ;
      RECT  7577.5 105862.5 7642.5 105727.5 ;
      RECT  7387.5 105862.5 7452.5 105727.5 ;
      RECT  7577.5 105862.5 7642.5 105727.5 ;
      RECT  7767.5 105862.5 7832.5 105727.5 ;
      RECT  7767.5 105862.5 7832.5 105727.5 ;
      RECT  7577.5 105862.5 7642.5 105727.5 ;
      RECT  7937.5 104932.5 8002.5 104797.5 ;
      RECT  7937.5 105907.5 8002.5 105772.5 ;
      RECT  7772.5 105650.0 7637.5 105585.0 ;
      RECT  7582.5 105510.0 7447.5 105445.0 ;
      RECT  7392.5 105370.0 7257.5 105305.0 ;
      RECT  7387.5 105022.5 7452.5 104887.5 ;
      RECT  7767.5 105022.5 7832.5 104887.5 ;
      RECT  7767.5 105862.5 7832.5 105727.5 ;
      RECT  7767.5 105405.0 7832.5 105270.0 ;
      RECT  7257.5 105370.0 7392.5 105305.0 ;
      RECT  7447.5 105510.0 7582.5 105445.0 ;
      RECT  7637.5 105650.0 7772.5 105585.0 ;
      RECT  7767.5 105405.0 7832.5 105270.0 ;
      RECT  7130.0 104712.5 8140.0 104647.5 ;
      RECT  7130.0 106057.5 8140.0 105992.5 ;
      RECT  7197.5 106187.5 7262.5 105992.5 ;
      RECT  7197.5 107027.5 7262.5 107402.5 ;
      RECT  7577.5 107027.5 7642.5 107402.5 ;
      RECT  7937.5 107185.0 8002.5 107370.0 ;
      RECT  7937.5 106025.0 8002.5 106210.0 ;
      RECT  7197.5 107027.5 7262.5 107162.5 ;
      RECT  7387.5 107027.5 7452.5 107162.5 ;
      RECT  7387.5 107027.5 7452.5 107162.5 ;
      RECT  7197.5 107027.5 7262.5 107162.5 ;
      RECT  7387.5 107027.5 7452.5 107162.5 ;
      RECT  7577.5 107027.5 7642.5 107162.5 ;
      RECT  7577.5 107027.5 7642.5 107162.5 ;
      RECT  7387.5 107027.5 7452.5 107162.5 ;
      RECT  7577.5 107027.5 7642.5 107162.5 ;
      RECT  7767.5 107027.5 7832.5 107162.5 ;
      RECT  7767.5 107027.5 7832.5 107162.5 ;
      RECT  7577.5 107027.5 7642.5 107162.5 ;
      RECT  7197.5 106187.5 7262.5 106322.5 ;
      RECT  7387.5 106187.5 7452.5 106322.5 ;
      RECT  7387.5 106187.5 7452.5 106322.5 ;
      RECT  7197.5 106187.5 7262.5 106322.5 ;
      RECT  7387.5 106187.5 7452.5 106322.5 ;
      RECT  7577.5 106187.5 7642.5 106322.5 ;
      RECT  7577.5 106187.5 7642.5 106322.5 ;
      RECT  7387.5 106187.5 7452.5 106322.5 ;
      RECT  7577.5 106187.5 7642.5 106322.5 ;
      RECT  7767.5 106187.5 7832.5 106322.5 ;
      RECT  7767.5 106187.5 7832.5 106322.5 ;
      RECT  7577.5 106187.5 7642.5 106322.5 ;
      RECT  7937.5 107117.5 8002.5 107252.5 ;
      RECT  7937.5 106142.5 8002.5 106277.5 ;
      RECT  7772.5 106400.0 7637.5 106465.0 ;
      RECT  7582.5 106540.0 7447.5 106605.0 ;
      RECT  7392.5 106680.0 7257.5 106745.0 ;
      RECT  7387.5 107027.5 7452.5 107162.5 ;
      RECT  7767.5 107027.5 7832.5 107162.5 ;
      RECT  7767.5 106187.5 7832.5 106322.5 ;
      RECT  7767.5 106645.0 7832.5 106780.0 ;
      RECT  7257.5 106680.0 7392.5 106745.0 ;
      RECT  7447.5 106540.0 7582.5 106605.0 ;
      RECT  7637.5 106400.0 7772.5 106465.0 ;
      RECT  7767.5 106645.0 7832.5 106780.0 ;
      RECT  7130.0 107337.5 8140.0 107402.5 ;
      RECT  7130.0 105992.5 8140.0 106057.5 ;
      RECT  7197.5 108552.5 7262.5 108747.5 ;
      RECT  7197.5 107712.5 7262.5 107337.5 ;
      RECT  7577.5 107712.5 7642.5 107337.5 ;
      RECT  7937.5 107555.0 8002.5 107370.0 ;
      RECT  7937.5 108715.0 8002.5 108530.0 ;
      RECT  7197.5 107712.5 7262.5 107577.5 ;
      RECT  7387.5 107712.5 7452.5 107577.5 ;
      RECT  7387.5 107712.5 7452.5 107577.5 ;
      RECT  7197.5 107712.5 7262.5 107577.5 ;
      RECT  7387.5 107712.5 7452.5 107577.5 ;
      RECT  7577.5 107712.5 7642.5 107577.5 ;
      RECT  7577.5 107712.5 7642.5 107577.5 ;
      RECT  7387.5 107712.5 7452.5 107577.5 ;
      RECT  7577.5 107712.5 7642.5 107577.5 ;
      RECT  7767.5 107712.5 7832.5 107577.5 ;
      RECT  7767.5 107712.5 7832.5 107577.5 ;
      RECT  7577.5 107712.5 7642.5 107577.5 ;
      RECT  7197.5 108552.5 7262.5 108417.5 ;
      RECT  7387.5 108552.5 7452.5 108417.5 ;
      RECT  7387.5 108552.5 7452.5 108417.5 ;
      RECT  7197.5 108552.5 7262.5 108417.5 ;
      RECT  7387.5 108552.5 7452.5 108417.5 ;
      RECT  7577.5 108552.5 7642.5 108417.5 ;
      RECT  7577.5 108552.5 7642.5 108417.5 ;
      RECT  7387.5 108552.5 7452.5 108417.5 ;
      RECT  7577.5 108552.5 7642.5 108417.5 ;
      RECT  7767.5 108552.5 7832.5 108417.5 ;
      RECT  7767.5 108552.5 7832.5 108417.5 ;
      RECT  7577.5 108552.5 7642.5 108417.5 ;
      RECT  7937.5 107622.5 8002.5 107487.5 ;
      RECT  7937.5 108597.5 8002.5 108462.5 ;
      RECT  7772.5 108340.0 7637.5 108275.0 ;
      RECT  7582.5 108200.0 7447.5 108135.0 ;
      RECT  7392.5 108060.0 7257.5 107995.0 ;
      RECT  7387.5 107712.5 7452.5 107577.5 ;
      RECT  7767.5 107712.5 7832.5 107577.5 ;
      RECT  7767.5 108552.5 7832.5 108417.5 ;
      RECT  7767.5 108095.0 7832.5 107960.0 ;
      RECT  7257.5 108060.0 7392.5 107995.0 ;
      RECT  7447.5 108200.0 7582.5 108135.0 ;
      RECT  7637.5 108340.0 7772.5 108275.0 ;
      RECT  7767.5 108095.0 7832.5 107960.0 ;
      RECT  7130.0 107402.5 8140.0 107337.5 ;
      RECT  7130.0 108747.5 8140.0 108682.5 ;
      RECT  7197.5 108877.5 7262.5 108682.5 ;
      RECT  7197.5 109717.5 7262.5 110092.5 ;
      RECT  7577.5 109717.5 7642.5 110092.5 ;
      RECT  7937.5 109875.0 8002.5 110060.0 ;
      RECT  7937.5 108715.0 8002.5 108900.0 ;
      RECT  7197.5 109717.5 7262.5 109852.5 ;
      RECT  7387.5 109717.5 7452.5 109852.5 ;
      RECT  7387.5 109717.5 7452.5 109852.5 ;
      RECT  7197.5 109717.5 7262.5 109852.5 ;
      RECT  7387.5 109717.5 7452.5 109852.5 ;
      RECT  7577.5 109717.5 7642.5 109852.5 ;
      RECT  7577.5 109717.5 7642.5 109852.5 ;
      RECT  7387.5 109717.5 7452.5 109852.5 ;
      RECT  7577.5 109717.5 7642.5 109852.5 ;
      RECT  7767.5 109717.5 7832.5 109852.5 ;
      RECT  7767.5 109717.5 7832.5 109852.5 ;
      RECT  7577.5 109717.5 7642.5 109852.5 ;
      RECT  7197.5 108877.5 7262.5 109012.5 ;
      RECT  7387.5 108877.5 7452.5 109012.5 ;
      RECT  7387.5 108877.5 7452.5 109012.5 ;
      RECT  7197.5 108877.5 7262.5 109012.5 ;
      RECT  7387.5 108877.5 7452.5 109012.5 ;
      RECT  7577.5 108877.5 7642.5 109012.5 ;
      RECT  7577.5 108877.5 7642.5 109012.5 ;
      RECT  7387.5 108877.5 7452.5 109012.5 ;
      RECT  7577.5 108877.5 7642.5 109012.5 ;
      RECT  7767.5 108877.5 7832.5 109012.5 ;
      RECT  7767.5 108877.5 7832.5 109012.5 ;
      RECT  7577.5 108877.5 7642.5 109012.5 ;
      RECT  7937.5 109807.5 8002.5 109942.5 ;
      RECT  7937.5 108832.5 8002.5 108967.5 ;
      RECT  7772.5 109090.0 7637.5 109155.0 ;
      RECT  7582.5 109230.0 7447.5 109295.0 ;
      RECT  7392.5 109370.0 7257.5 109435.0 ;
      RECT  7387.5 109717.5 7452.5 109852.5 ;
      RECT  7767.5 109717.5 7832.5 109852.5 ;
      RECT  7767.5 108877.5 7832.5 109012.5 ;
      RECT  7767.5 109335.0 7832.5 109470.0 ;
      RECT  7257.5 109370.0 7392.5 109435.0 ;
      RECT  7447.5 109230.0 7582.5 109295.0 ;
      RECT  7637.5 109090.0 7772.5 109155.0 ;
      RECT  7767.5 109335.0 7832.5 109470.0 ;
      RECT  7130.0 110027.5 8140.0 110092.5 ;
      RECT  7130.0 108682.5 8140.0 108747.5 ;
      RECT  7197.5 111242.5 7262.5 111437.5 ;
      RECT  7197.5 110402.5 7262.5 110027.5 ;
      RECT  7577.5 110402.5 7642.5 110027.5 ;
      RECT  7937.5 110245.0 8002.5 110060.0 ;
      RECT  7937.5 111405.0 8002.5 111220.0 ;
      RECT  7197.5 110402.5 7262.5 110267.5 ;
      RECT  7387.5 110402.5 7452.5 110267.5 ;
      RECT  7387.5 110402.5 7452.5 110267.5 ;
      RECT  7197.5 110402.5 7262.5 110267.5 ;
      RECT  7387.5 110402.5 7452.5 110267.5 ;
      RECT  7577.5 110402.5 7642.5 110267.5 ;
      RECT  7577.5 110402.5 7642.5 110267.5 ;
      RECT  7387.5 110402.5 7452.5 110267.5 ;
      RECT  7577.5 110402.5 7642.5 110267.5 ;
      RECT  7767.5 110402.5 7832.5 110267.5 ;
      RECT  7767.5 110402.5 7832.5 110267.5 ;
      RECT  7577.5 110402.5 7642.5 110267.5 ;
      RECT  7197.5 111242.5 7262.5 111107.5 ;
      RECT  7387.5 111242.5 7452.5 111107.5 ;
      RECT  7387.5 111242.5 7452.5 111107.5 ;
      RECT  7197.5 111242.5 7262.5 111107.5 ;
      RECT  7387.5 111242.5 7452.5 111107.5 ;
      RECT  7577.5 111242.5 7642.5 111107.5 ;
      RECT  7577.5 111242.5 7642.5 111107.5 ;
      RECT  7387.5 111242.5 7452.5 111107.5 ;
      RECT  7577.5 111242.5 7642.5 111107.5 ;
      RECT  7767.5 111242.5 7832.5 111107.5 ;
      RECT  7767.5 111242.5 7832.5 111107.5 ;
      RECT  7577.5 111242.5 7642.5 111107.5 ;
      RECT  7937.5 110312.5 8002.5 110177.5 ;
      RECT  7937.5 111287.5 8002.5 111152.5 ;
      RECT  7772.5 111030.0 7637.5 110965.0 ;
      RECT  7582.5 110890.0 7447.5 110825.0 ;
      RECT  7392.5 110750.0 7257.5 110685.0 ;
      RECT  7387.5 110402.5 7452.5 110267.5 ;
      RECT  7767.5 110402.5 7832.5 110267.5 ;
      RECT  7767.5 111242.5 7832.5 111107.5 ;
      RECT  7767.5 110785.0 7832.5 110650.0 ;
      RECT  7257.5 110750.0 7392.5 110685.0 ;
      RECT  7447.5 110890.0 7582.5 110825.0 ;
      RECT  7637.5 111030.0 7772.5 110965.0 ;
      RECT  7767.5 110785.0 7832.5 110650.0 ;
      RECT  7130.0 110092.5 8140.0 110027.5 ;
      RECT  7130.0 111437.5 8140.0 111372.5 ;
      RECT  7197.5 111567.5 7262.5 111372.5 ;
      RECT  7197.5 112407.5 7262.5 112782.5 ;
      RECT  7577.5 112407.5 7642.5 112782.5 ;
      RECT  7937.5 112565.0 8002.5 112750.0 ;
      RECT  7937.5 111405.0 8002.5 111590.0 ;
      RECT  7197.5 112407.5 7262.5 112542.5 ;
      RECT  7387.5 112407.5 7452.5 112542.5 ;
      RECT  7387.5 112407.5 7452.5 112542.5 ;
      RECT  7197.5 112407.5 7262.5 112542.5 ;
      RECT  7387.5 112407.5 7452.5 112542.5 ;
      RECT  7577.5 112407.5 7642.5 112542.5 ;
      RECT  7577.5 112407.5 7642.5 112542.5 ;
      RECT  7387.5 112407.5 7452.5 112542.5 ;
      RECT  7577.5 112407.5 7642.5 112542.5 ;
      RECT  7767.5 112407.5 7832.5 112542.5 ;
      RECT  7767.5 112407.5 7832.5 112542.5 ;
      RECT  7577.5 112407.5 7642.5 112542.5 ;
      RECT  7197.5 111567.5 7262.5 111702.5 ;
      RECT  7387.5 111567.5 7452.5 111702.5 ;
      RECT  7387.5 111567.5 7452.5 111702.5 ;
      RECT  7197.5 111567.5 7262.5 111702.5 ;
      RECT  7387.5 111567.5 7452.5 111702.5 ;
      RECT  7577.5 111567.5 7642.5 111702.5 ;
      RECT  7577.5 111567.5 7642.5 111702.5 ;
      RECT  7387.5 111567.5 7452.5 111702.5 ;
      RECT  7577.5 111567.5 7642.5 111702.5 ;
      RECT  7767.5 111567.5 7832.5 111702.5 ;
      RECT  7767.5 111567.5 7832.5 111702.5 ;
      RECT  7577.5 111567.5 7642.5 111702.5 ;
      RECT  7937.5 112497.5 8002.5 112632.5 ;
      RECT  7937.5 111522.5 8002.5 111657.5 ;
      RECT  7772.5 111780.0 7637.5 111845.0 ;
      RECT  7582.5 111920.0 7447.5 111985.0 ;
      RECT  7392.5 112060.0 7257.5 112125.0 ;
      RECT  7387.5 112407.5 7452.5 112542.5 ;
      RECT  7767.5 112407.5 7832.5 112542.5 ;
      RECT  7767.5 111567.5 7832.5 111702.5 ;
      RECT  7767.5 112025.0 7832.5 112160.0 ;
      RECT  7257.5 112060.0 7392.5 112125.0 ;
      RECT  7447.5 111920.0 7582.5 111985.0 ;
      RECT  7637.5 111780.0 7772.5 111845.0 ;
      RECT  7767.5 112025.0 7832.5 112160.0 ;
      RECT  7130.0 112717.5 8140.0 112782.5 ;
      RECT  7130.0 111372.5 8140.0 111437.5 ;
      RECT  7197.5 113932.5 7262.5 114127.5 ;
      RECT  7197.5 113092.5 7262.5 112717.5 ;
      RECT  7577.5 113092.5 7642.5 112717.5 ;
      RECT  7937.5 112935.0 8002.5 112750.0 ;
      RECT  7937.5 114095.0 8002.5 113910.0 ;
      RECT  7197.5 113092.5 7262.5 112957.5 ;
      RECT  7387.5 113092.5 7452.5 112957.5 ;
      RECT  7387.5 113092.5 7452.5 112957.5 ;
      RECT  7197.5 113092.5 7262.5 112957.5 ;
      RECT  7387.5 113092.5 7452.5 112957.5 ;
      RECT  7577.5 113092.5 7642.5 112957.5 ;
      RECT  7577.5 113092.5 7642.5 112957.5 ;
      RECT  7387.5 113092.5 7452.5 112957.5 ;
      RECT  7577.5 113092.5 7642.5 112957.5 ;
      RECT  7767.5 113092.5 7832.5 112957.5 ;
      RECT  7767.5 113092.5 7832.5 112957.5 ;
      RECT  7577.5 113092.5 7642.5 112957.5 ;
      RECT  7197.5 113932.5 7262.5 113797.5 ;
      RECT  7387.5 113932.5 7452.5 113797.5 ;
      RECT  7387.5 113932.5 7452.5 113797.5 ;
      RECT  7197.5 113932.5 7262.5 113797.5 ;
      RECT  7387.5 113932.5 7452.5 113797.5 ;
      RECT  7577.5 113932.5 7642.5 113797.5 ;
      RECT  7577.5 113932.5 7642.5 113797.5 ;
      RECT  7387.5 113932.5 7452.5 113797.5 ;
      RECT  7577.5 113932.5 7642.5 113797.5 ;
      RECT  7767.5 113932.5 7832.5 113797.5 ;
      RECT  7767.5 113932.5 7832.5 113797.5 ;
      RECT  7577.5 113932.5 7642.5 113797.5 ;
      RECT  7937.5 113002.5 8002.5 112867.5 ;
      RECT  7937.5 113977.5 8002.5 113842.5 ;
      RECT  7772.5 113720.0 7637.5 113655.0 ;
      RECT  7582.5 113580.0 7447.5 113515.0 ;
      RECT  7392.5 113440.0 7257.5 113375.0 ;
      RECT  7387.5 113092.5 7452.5 112957.5 ;
      RECT  7767.5 113092.5 7832.5 112957.5 ;
      RECT  7767.5 113932.5 7832.5 113797.5 ;
      RECT  7767.5 113475.0 7832.5 113340.0 ;
      RECT  7257.5 113440.0 7392.5 113375.0 ;
      RECT  7447.5 113580.0 7582.5 113515.0 ;
      RECT  7637.5 113720.0 7772.5 113655.0 ;
      RECT  7767.5 113475.0 7832.5 113340.0 ;
      RECT  7130.0 112782.5 8140.0 112717.5 ;
      RECT  7130.0 114127.5 8140.0 114062.5 ;
      RECT  8567.5 29175.0 8632.5 29360.0 ;
      RECT  8567.5 28015.0 8632.5 28200.0 ;
      RECT  8207.5 28132.5 8272.5 27982.5 ;
      RECT  8207.5 29017.5 8272.5 29392.5 ;
      RECT  8397.5 28132.5 8462.5 29017.5 ;
      RECT  8207.5 29017.5 8272.5 29152.5 ;
      RECT  8397.5 29017.5 8462.5 29152.5 ;
      RECT  8397.5 29017.5 8462.5 29152.5 ;
      RECT  8207.5 29017.5 8272.5 29152.5 ;
      RECT  8207.5 28132.5 8272.5 28267.5 ;
      RECT  8397.5 28132.5 8462.5 28267.5 ;
      RECT  8397.5 28132.5 8462.5 28267.5 ;
      RECT  8207.5 28132.5 8272.5 28267.5 ;
      RECT  8567.5 29107.5 8632.5 29242.5 ;
      RECT  8567.5 28132.5 8632.5 28267.5 ;
      RECT  8265.0 28575.0 8330.0 28710.0 ;
      RECT  8265.0 28575.0 8330.0 28710.0 ;
      RECT  8430.0 28610.0 8495.0 28675.0 ;
      RECT  8140.0 29327.5 8700.0 29392.5 ;
      RECT  8140.0 27982.5 8700.0 28047.5 ;
      RECT  8567.5 29545.0 8632.5 29360.0 ;
      RECT  8567.5 30705.0 8632.5 30520.0 ;
      RECT  8207.5 30587.5 8272.5 30737.5 ;
      RECT  8207.5 29702.5 8272.5 29327.5 ;
      RECT  8397.5 30587.5 8462.5 29702.5 ;
      RECT  8207.5 29702.5 8272.5 29567.5 ;
      RECT  8397.5 29702.5 8462.5 29567.5 ;
      RECT  8397.5 29702.5 8462.5 29567.5 ;
      RECT  8207.5 29702.5 8272.5 29567.5 ;
      RECT  8207.5 30587.5 8272.5 30452.5 ;
      RECT  8397.5 30587.5 8462.5 30452.5 ;
      RECT  8397.5 30587.5 8462.5 30452.5 ;
      RECT  8207.5 30587.5 8272.5 30452.5 ;
      RECT  8567.5 29612.5 8632.5 29477.5 ;
      RECT  8567.5 30587.5 8632.5 30452.5 ;
      RECT  8265.0 30145.0 8330.0 30010.0 ;
      RECT  8265.0 30145.0 8330.0 30010.0 ;
      RECT  8430.0 30110.0 8495.0 30045.0 ;
      RECT  8140.0 29392.5 8700.0 29327.5 ;
      RECT  8140.0 30737.5 8700.0 30672.5 ;
      RECT  8567.5 31865.0 8632.5 32050.0 ;
      RECT  8567.5 30705.0 8632.5 30890.0 ;
      RECT  8207.5 30822.5 8272.5 30672.5 ;
      RECT  8207.5 31707.5 8272.5 32082.5 ;
      RECT  8397.5 30822.5 8462.5 31707.5 ;
      RECT  8207.5 31707.5 8272.5 31842.5 ;
      RECT  8397.5 31707.5 8462.5 31842.5 ;
      RECT  8397.5 31707.5 8462.5 31842.5 ;
      RECT  8207.5 31707.5 8272.5 31842.5 ;
      RECT  8207.5 30822.5 8272.5 30957.5 ;
      RECT  8397.5 30822.5 8462.5 30957.5 ;
      RECT  8397.5 30822.5 8462.5 30957.5 ;
      RECT  8207.5 30822.5 8272.5 30957.5 ;
      RECT  8567.5 31797.5 8632.5 31932.5 ;
      RECT  8567.5 30822.5 8632.5 30957.5 ;
      RECT  8265.0 31265.0 8330.0 31400.0 ;
      RECT  8265.0 31265.0 8330.0 31400.0 ;
      RECT  8430.0 31300.0 8495.0 31365.0 ;
      RECT  8140.0 32017.5 8700.0 32082.5 ;
      RECT  8140.0 30672.5 8700.0 30737.5 ;
      RECT  8567.5 32235.0 8632.5 32050.0 ;
      RECT  8567.5 33395.0 8632.5 33210.0 ;
      RECT  8207.5 33277.5 8272.5 33427.5 ;
      RECT  8207.5 32392.5 8272.5 32017.5 ;
      RECT  8397.5 33277.5 8462.5 32392.5 ;
      RECT  8207.5 32392.5 8272.5 32257.5 ;
      RECT  8397.5 32392.5 8462.5 32257.5 ;
      RECT  8397.5 32392.5 8462.5 32257.5 ;
      RECT  8207.5 32392.5 8272.5 32257.5 ;
      RECT  8207.5 33277.5 8272.5 33142.5 ;
      RECT  8397.5 33277.5 8462.5 33142.5 ;
      RECT  8397.5 33277.5 8462.5 33142.5 ;
      RECT  8207.5 33277.5 8272.5 33142.5 ;
      RECT  8567.5 32302.5 8632.5 32167.5 ;
      RECT  8567.5 33277.5 8632.5 33142.5 ;
      RECT  8265.0 32835.0 8330.0 32700.0 ;
      RECT  8265.0 32835.0 8330.0 32700.0 ;
      RECT  8430.0 32800.0 8495.0 32735.0 ;
      RECT  8140.0 32082.5 8700.0 32017.5 ;
      RECT  8140.0 33427.5 8700.0 33362.5 ;
      RECT  8567.5 34555.0 8632.5 34740.0 ;
      RECT  8567.5 33395.0 8632.5 33580.0 ;
      RECT  8207.5 33512.5 8272.5 33362.5 ;
      RECT  8207.5 34397.5 8272.5 34772.5 ;
      RECT  8397.5 33512.5 8462.5 34397.5 ;
      RECT  8207.5 34397.5 8272.5 34532.5 ;
      RECT  8397.5 34397.5 8462.5 34532.5 ;
      RECT  8397.5 34397.5 8462.5 34532.5 ;
      RECT  8207.5 34397.5 8272.5 34532.5 ;
      RECT  8207.5 33512.5 8272.5 33647.5 ;
      RECT  8397.5 33512.5 8462.5 33647.5 ;
      RECT  8397.5 33512.5 8462.5 33647.5 ;
      RECT  8207.5 33512.5 8272.5 33647.5 ;
      RECT  8567.5 34487.5 8632.5 34622.5 ;
      RECT  8567.5 33512.5 8632.5 33647.5 ;
      RECT  8265.0 33955.0 8330.0 34090.0 ;
      RECT  8265.0 33955.0 8330.0 34090.0 ;
      RECT  8430.0 33990.0 8495.0 34055.0 ;
      RECT  8140.0 34707.5 8700.0 34772.5 ;
      RECT  8140.0 33362.5 8700.0 33427.5 ;
      RECT  8567.5 34925.0 8632.5 34740.0 ;
      RECT  8567.5 36085.0 8632.5 35900.0 ;
      RECT  8207.5 35967.5 8272.5 36117.5 ;
      RECT  8207.5 35082.5 8272.5 34707.5 ;
      RECT  8397.5 35967.5 8462.5 35082.5 ;
      RECT  8207.5 35082.5 8272.5 34947.5 ;
      RECT  8397.5 35082.5 8462.5 34947.5 ;
      RECT  8397.5 35082.5 8462.5 34947.5 ;
      RECT  8207.5 35082.5 8272.5 34947.5 ;
      RECT  8207.5 35967.5 8272.5 35832.5 ;
      RECT  8397.5 35967.5 8462.5 35832.5 ;
      RECT  8397.5 35967.5 8462.5 35832.5 ;
      RECT  8207.5 35967.5 8272.5 35832.5 ;
      RECT  8567.5 34992.5 8632.5 34857.5 ;
      RECT  8567.5 35967.5 8632.5 35832.5 ;
      RECT  8265.0 35525.0 8330.0 35390.0 ;
      RECT  8265.0 35525.0 8330.0 35390.0 ;
      RECT  8430.0 35490.0 8495.0 35425.0 ;
      RECT  8140.0 34772.5 8700.0 34707.5 ;
      RECT  8140.0 36117.5 8700.0 36052.5 ;
      RECT  8567.5 37245.0 8632.5 37430.0 ;
      RECT  8567.5 36085.0 8632.5 36270.0 ;
      RECT  8207.5 36202.5 8272.5 36052.5 ;
      RECT  8207.5 37087.5 8272.5 37462.5 ;
      RECT  8397.5 36202.5 8462.5 37087.5 ;
      RECT  8207.5 37087.5 8272.5 37222.5 ;
      RECT  8397.5 37087.5 8462.5 37222.5 ;
      RECT  8397.5 37087.5 8462.5 37222.5 ;
      RECT  8207.5 37087.5 8272.5 37222.5 ;
      RECT  8207.5 36202.5 8272.5 36337.5 ;
      RECT  8397.5 36202.5 8462.5 36337.5 ;
      RECT  8397.5 36202.5 8462.5 36337.5 ;
      RECT  8207.5 36202.5 8272.5 36337.5 ;
      RECT  8567.5 37177.5 8632.5 37312.5 ;
      RECT  8567.5 36202.5 8632.5 36337.5 ;
      RECT  8265.0 36645.0 8330.0 36780.0 ;
      RECT  8265.0 36645.0 8330.0 36780.0 ;
      RECT  8430.0 36680.0 8495.0 36745.0 ;
      RECT  8140.0 37397.5 8700.0 37462.5 ;
      RECT  8140.0 36052.5 8700.0 36117.5 ;
      RECT  8567.5 37615.0 8632.5 37430.0 ;
      RECT  8567.5 38775.0 8632.5 38590.0 ;
      RECT  8207.5 38657.5 8272.5 38807.5 ;
      RECT  8207.5 37772.5 8272.5 37397.5 ;
      RECT  8397.5 38657.5 8462.5 37772.5 ;
      RECT  8207.5 37772.5 8272.5 37637.5 ;
      RECT  8397.5 37772.5 8462.5 37637.5 ;
      RECT  8397.5 37772.5 8462.5 37637.5 ;
      RECT  8207.5 37772.5 8272.5 37637.5 ;
      RECT  8207.5 38657.5 8272.5 38522.5 ;
      RECT  8397.5 38657.5 8462.5 38522.5 ;
      RECT  8397.5 38657.5 8462.5 38522.5 ;
      RECT  8207.5 38657.5 8272.5 38522.5 ;
      RECT  8567.5 37682.5 8632.5 37547.5 ;
      RECT  8567.5 38657.5 8632.5 38522.5 ;
      RECT  8265.0 38215.0 8330.0 38080.0 ;
      RECT  8265.0 38215.0 8330.0 38080.0 ;
      RECT  8430.0 38180.0 8495.0 38115.0 ;
      RECT  8140.0 37462.5 8700.0 37397.5 ;
      RECT  8140.0 38807.5 8700.0 38742.5 ;
      RECT  8567.5 39935.0 8632.5 40120.0 ;
      RECT  8567.5 38775.0 8632.5 38960.0 ;
      RECT  8207.5 38892.5 8272.5 38742.5 ;
      RECT  8207.5 39777.5 8272.5 40152.5 ;
      RECT  8397.5 38892.5 8462.5 39777.5 ;
      RECT  8207.5 39777.5 8272.5 39912.5 ;
      RECT  8397.5 39777.5 8462.5 39912.5 ;
      RECT  8397.5 39777.5 8462.5 39912.5 ;
      RECT  8207.5 39777.5 8272.5 39912.5 ;
      RECT  8207.5 38892.5 8272.5 39027.5 ;
      RECT  8397.5 38892.5 8462.5 39027.5 ;
      RECT  8397.5 38892.5 8462.5 39027.5 ;
      RECT  8207.5 38892.5 8272.5 39027.5 ;
      RECT  8567.5 39867.5 8632.5 40002.5 ;
      RECT  8567.5 38892.5 8632.5 39027.5 ;
      RECT  8265.0 39335.0 8330.0 39470.0 ;
      RECT  8265.0 39335.0 8330.0 39470.0 ;
      RECT  8430.0 39370.0 8495.0 39435.0 ;
      RECT  8140.0 40087.5 8700.0 40152.5 ;
      RECT  8140.0 38742.5 8700.0 38807.5 ;
      RECT  8567.5 40305.0 8632.5 40120.0 ;
      RECT  8567.5 41465.0 8632.5 41280.0 ;
      RECT  8207.5 41347.5 8272.5 41497.5 ;
      RECT  8207.5 40462.5 8272.5 40087.5 ;
      RECT  8397.5 41347.5 8462.5 40462.5 ;
      RECT  8207.5 40462.5 8272.5 40327.5 ;
      RECT  8397.5 40462.5 8462.5 40327.5 ;
      RECT  8397.5 40462.5 8462.5 40327.5 ;
      RECT  8207.5 40462.5 8272.5 40327.5 ;
      RECT  8207.5 41347.5 8272.5 41212.5 ;
      RECT  8397.5 41347.5 8462.5 41212.5 ;
      RECT  8397.5 41347.5 8462.5 41212.5 ;
      RECT  8207.5 41347.5 8272.5 41212.5 ;
      RECT  8567.5 40372.5 8632.5 40237.5 ;
      RECT  8567.5 41347.5 8632.5 41212.5 ;
      RECT  8265.0 40905.0 8330.0 40770.0 ;
      RECT  8265.0 40905.0 8330.0 40770.0 ;
      RECT  8430.0 40870.0 8495.0 40805.0 ;
      RECT  8140.0 40152.5 8700.0 40087.5 ;
      RECT  8140.0 41497.5 8700.0 41432.5 ;
      RECT  8567.5 42625.0 8632.5 42810.0 ;
      RECT  8567.5 41465.0 8632.5 41650.0 ;
      RECT  8207.5 41582.5 8272.5 41432.5 ;
      RECT  8207.5 42467.5 8272.5 42842.5 ;
      RECT  8397.5 41582.5 8462.5 42467.5 ;
      RECT  8207.5 42467.5 8272.5 42602.5 ;
      RECT  8397.5 42467.5 8462.5 42602.5 ;
      RECT  8397.5 42467.5 8462.5 42602.5 ;
      RECT  8207.5 42467.5 8272.5 42602.5 ;
      RECT  8207.5 41582.5 8272.5 41717.5 ;
      RECT  8397.5 41582.5 8462.5 41717.5 ;
      RECT  8397.5 41582.5 8462.5 41717.5 ;
      RECT  8207.5 41582.5 8272.5 41717.5 ;
      RECT  8567.5 42557.5 8632.5 42692.5 ;
      RECT  8567.5 41582.5 8632.5 41717.5 ;
      RECT  8265.0 42025.0 8330.0 42160.0 ;
      RECT  8265.0 42025.0 8330.0 42160.0 ;
      RECT  8430.0 42060.0 8495.0 42125.0 ;
      RECT  8140.0 42777.5 8700.0 42842.5 ;
      RECT  8140.0 41432.5 8700.0 41497.5 ;
      RECT  8567.5 42995.0 8632.5 42810.0 ;
      RECT  8567.5 44155.0 8632.5 43970.0 ;
      RECT  8207.5 44037.5 8272.5 44187.5 ;
      RECT  8207.5 43152.5 8272.5 42777.5 ;
      RECT  8397.5 44037.5 8462.5 43152.5 ;
      RECT  8207.5 43152.5 8272.5 43017.5 ;
      RECT  8397.5 43152.5 8462.5 43017.5 ;
      RECT  8397.5 43152.5 8462.5 43017.5 ;
      RECT  8207.5 43152.5 8272.5 43017.5 ;
      RECT  8207.5 44037.5 8272.5 43902.5 ;
      RECT  8397.5 44037.5 8462.5 43902.5 ;
      RECT  8397.5 44037.5 8462.5 43902.5 ;
      RECT  8207.5 44037.5 8272.5 43902.5 ;
      RECT  8567.5 43062.5 8632.5 42927.5 ;
      RECT  8567.5 44037.5 8632.5 43902.5 ;
      RECT  8265.0 43595.0 8330.0 43460.0 ;
      RECT  8265.0 43595.0 8330.0 43460.0 ;
      RECT  8430.0 43560.0 8495.0 43495.0 ;
      RECT  8140.0 42842.5 8700.0 42777.5 ;
      RECT  8140.0 44187.5 8700.0 44122.5 ;
      RECT  8567.5 45315.0 8632.5 45500.0 ;
      RECT  8567.5 44155.0 8632.5 44340.0 ;
      RECT  8207.5 44272.5 8272.5 44122.5 ;
      RECT  8207.5 45157.5 8272.5 45532.5 ;
      RECT  8397.5 44272.5 8462.5 45157.5 ;
      RECT  8207.5 45157.5 8272.5 45292.5 ;
      RECT  8397.5 45157.5 8462.5 45292.5 ;
      RECT  8397.5 45157.5 8462.5 45292.5 ;
      RECT  8207.5 45157.5 8272.5 45292.5 ;
      RECT  8207.5 44272.5 8272.5 44407.5 ;
      RECT  8397.5 44272.5 8462.5 44407.5 ;
      RECT  8397.5 44272.5 8462.5 44407.5 ;
      RECT  8207.5 44272.5 8272.5 44407.5 ;
      RECT  8567.5 45247.5 8632.5 45382.5 ;
      RECT  8567.5 44272.5 8632.5 44407.5 ;
      RECT  8265.0 44715.0 8330.0 44850.0 ;
      RECT  8265.0 44715.0 8330.0 44850.0 ;
      RECT  8430.0 44750.0 8495.0 44815.0 ;
      RECT  8140.0 45467.5 8700.0 45532.5 ;
      RECT  8140.0 44122.5 8700.0 44187.5 ;
      RECT  8567.5 45685.0 8632.5 45500.0 ;
      RECT  8567.5 46845.0 8632.5 46660.0 ;
      RECT  8207.5 46727.5 8272.5 46877.5 ;
      RECT  8207.5 45842.5 8272.5 45467.5 ;
      RECT  8397.5 46727.5 8462.5 45842.5 ;
      RECT  8207.5 45842.5 8272.5 45707.5 ;
      RECT  8397.5 45842.5 8462.5 45707.5 ;
      RECT  8397.5 45842.5 8462.5 45707.5 ;
      RECT  8207.5 45842.5 8272.5 45707.5 ;
      RECT  8207.5 46727.5 8272.5 46592.5 ;
      RECT  8397.5 46727.5 8462.5 46592.5 ;
      RECT  8397.5 46727.5 8462.5 46592.5 ;
      RECT  8207.5 46727.5 8272.5 46592.5 ;
      RECT  8567.5 45752.5 8632.5 45617.5 ;
      RECT  8567.5 46727.5 8632.5 46592.5 ;
      RECT  8265.0 46285.0 8330.0 46150.0 ;
      RECT  8265.0 46285.0 8330.0 46150.0 ;
      RECT  8430.0 46250.0 8495.0 46185.0 ;
      RECT  8140.0 45532.5 8700.0 45467.5 ;
      RECT  8140.0 46877.5 8700.0 46812.5 ;
      RECT  8567.5 48005.0 8632.5 48190.0 ;
      RECT  8567.5 46845.0 8632.5 47030.0 ;
      RECT  8207.5 46962.5 8272.5 46812.5 ;
      RECT  8207.5 47847.5 8272.5 48222.5 ;
      RECT  8397.5 46962.5 8462.5 47847.5 ;
      RECT  8207.5 47847.5 8272.5 47982.5 ;
      RECT  8397.5 47847.5 8462.5 47982.5 ;
      RECT  8397.5 47847.5 8462.5 47982.5 ;
      RECT  8207.5 47847.5 8272.5 47982.5 ;
      RECT  8207.5 46962.5 8272.5 47097.5 ;
      RECT  8397.5 46962.5 8462.5 47097.5 ;
      RECT  8397.5 46962.5 8462.5 47097.5 ;
      RECT  8207.5 46962.5 8272.5 47097.5 ;
      RECT  8567.5 47937.5 8632.5 48072.5 ;
      RECT  8567.5 46962.5 8632.5 47097.5 ;
      RECT  8265.0 47405.0 8330.0 47540.0 ;
      RECT  8265.0 47405.0 8330.0 47540.0 ;
      RECT  8430.0 47440.0 8495.0 47505.0 ;
      RECT  8140.0 48157.5 8700.0 48222.5 ;
      RECT  8140.0 46812.5 8700.0 46877.5 ;
      RECT  8567.5 48375.0 8632.5 48190.0 ;
      RECT  8567.5 49535.0 8632.5 49350.0 ;
      RECT  8207.5 49417.5 8272.5 49567.5 ;
      RECT  8207.5 48532.5 8272.5 48157.5 ;
      RECT  8397.5 49417.5 8462.5 48532.5 ;
      RECT  8207.5 48532.5 8272.5 48397.5 ;
      RECT  8397.5 48532.5 8462.5 48397.5 ;
      RECT  8397.5 48532.5 8462.5 48397.5 ;
      RECT  8207.5 48532.5 8272.5 48397.5 ;
      RECT  8207.5 49417.5 8272.5 49282.5 ;
      RECT  8397.5 49417.5 8462.5 49282.5 ;
      RECT  8397.5 49417.5 8462.5 49282.5 ;
      RECT  8207.5 49417.5 8272.5 49282.5 ;
      RECT  8567.5 48442.5 8632.5 48307.5 ;
      RECT  8567.5 49417.5 8632.5 49282.5 ;
      RECT  8265.0 48975.0 8330.0 48840.0 ;
      RECT  8265.0 48975.0 8330.0 48840.0 ;
      RECT  8430.0 48940.0 8495.0 48875.0 ;
      RECT  8140.0 48222.5 8700.0 48157.5 ;
      RECT  8140.0 49567.5 8700.0 49502.5 ;
      RECT  8567.5 50695.0 8632.5 50880.0 ;
      RECT  8567.5 49535.0 8632.5 49720.0 ;
      RECT  8207.5 49652.5 8272.5 49502.5 ;
      RECT  8207.5 50537.5 8272.5 50912.5 ;
      RECT  8397.5 49652.5 8462.5 50537.5 ;
      RECT  8207.5 50537.5 8272.5 50672.5 ;
      RECT  8397.5 50537.5 8462.5 50672.5 ;
      RECT  8397.5 50537.5 8462.5 50672.5 ;
      RECT  8207.5 50537.5 8272.5 50672.5 ;
      RECT  8207.5 49652.5 8272.5 49787.5 ;
      RECT  8397.5 49652.5 8462.5 49787.5 ;
      RECT  8397.5 49652.5 8462.5 49787.5 ;
      RECT  8207.5 49652.5 8272.5 49787.5 ;
      RECT  8567.5 50627.5 8632.5 50762.5 ;
      RECT  8567.5 49652.5 8632.5 49787.5 ;
      RECT  8265.0 50095.0 8330.0 50230.0 ;
      RECT  8265.0 50095.0 8330.0 50230.0 ;
      RECT  8430.0 50130.0 8495.0 50195.0 ;
      RECT  8140.0 50847.5 8700.0 50912.5 ;
      RECT  8140.0 49502.5 8700.0 49567.5 ;
      RECT  8567.5 51065.0 8632.5 50880.0 ;
      RECT  8567.5 52225.0 8632.5 52040.0 ;
      RECT  8207.5 52107.5 8272.5 52257.5 ;
      RECT  8207.5 51222.5 8272.5 50847.5 ;
      RECT  8397.5 52107.5 8462.5 51222.5 ;
      RECT  8207.5 51222.5 8272.5 51087.5 ;
      RECT  8397.5 51222.5 8462.5 51087.5 ;
      RECT  8397.5 51222.5 8462.5 51087.5 ;
      RECT  8207.5 51222.5 8272.5 51087.5 ;
      RECT  8207.5 52107.5 8272.5 51972.5 ;
      RECT  8397.5 52107.5 8462.5 51972.5 ;
      RECT  8397.5 52107.5 8462.5 51972.5 ;
      RECT  8207.5 52107.5 8272.5 51972.5 ;
      RECT  8567.5 51132.5 8632.5 50997.5 ;
      RECT  8567.5 52107.5 8632.5 51972.5 ;
      RECT  8265.0 51665.0 8330.0 51530.0 ;
      RECT  8265.0 51665.0 8330.0 51530.0 ;
      RECT  8430.0 51630.0 8495.0 51565.0 ;
      RECT  8140.0 50912.5 8700.0 50847.5 ;
      RECT  8140.0 52257.5 8700.0 52192.5 ;
      RECT  8567.5 53385.0 8632.5 53570.0 ;
      RECT  8567.5 52225.0 8632.5 52410.0 ;
      RECT  8207.5 52342.5 8272.5 52192.5 ;
      RECT  8207.5 53227.5 8272.5 53602.5 ;
      RECT  8397.5 52342.5 8462.5 53227.5 ;
      RECT  8207.5 53227.5 8272.5 53362.5 ;
      RECT  8397.5 53227.5 8462.5 53362.5 ;
      RECT  8397.5 53227.5 8462.5 53362.5 ;
      RECT  8207.5 53227.5 8272.5 53362.5 ;
      RECT  8207.5 52342.5 8272.5 52477.5 ;
      RECT  8397.5 52342.5 8462.5 52477.5 ;
      RECT  8397.5 52342.5 8462.5 52477.5 ;
      RECT  8207.5 52342.5 8272.5 52477.5 ;
      RECT  8567.5 53317.5 8632.5 53452.5 ;
      RECT  8567.5 52342.5 8632.5 52477.5 ;
      RECT  8265.0 52785.0 8330.0 52920.0 ;
      RECT  8265.0 52785.0 8330.0 52920.0 ;
      RECT  8430.0 52820.0 8495.0 52885.0 ;
      RECT  8140.0 53537.5 8700.0 53602.5 ;
      RECT  8140.0 52192.5 8700.0 52257.5 ;
      RECT  8567.5 53755.0 8632.5 53570.0 ;
      RECT  8567.5 54915.0 8632.5 54730.0 ;
      RECT  8207.5 54797.5 8272.5 54947.5 ;
      RECT  8207.5 53912.5 8272.5 53537.5 ;
      RECT  8397.5 54797.5 8462.5 53912.5 ;
      RECT  8207.5 53912.5 8272.5 53777.5 ;
      RECT  8397.5 53912.5 8462.5 53777.5 ;
      RECT  8397.5 53912.5 8462.5 53777.5 ;
      RECT  8207.5 53912.5 8272.5 53777.5 ;
      RECT  8207.5 54797.5 8272.5 54662.5 ;
      RECT  8397.5 54797.5 8462.5 54662.5 ;
      RECT  8397.5 54797.5 8462.5 54662.5 ;
      RECT  8207.5 54797.5 8272.5 54662.5 ;
      RECT  8567.5 53822.5 8632.5 53687.5 ;
      RECT  8567.5 54797.5 8632.5 54662.5 ;
      RECT  8265.0 54355.0 8330.0 54220.0 ;
      RECT  8265.0 54355.0 8330.0 54220.0 ;
      RECT  8430.0 54320.0 8495.0 54255.0 ;
      RECT  8140.0 53602.5 8700.0 53537.5 ;
      RECT  8140.0 54947.5 8700.0 54882.5 ;
      RECT  8567.5 56075.0 8632.5 56260.0 ;
      RECT  8567.5 54915.0 8632.5 55100.0 ;
      RECT  8207.5 55032.5 8272.5 54882.5 ;
      RECT  8207.5 55917.5 8272.5 56292.5 ;
      RECT  8397.5 55032.5 8462.5 55917.5 ;
      RECT  8207.5 55917.5 8272.5 56052.5 ;
      RECT  8397.5 55917.5 8462.5 56052.5 ;
      RECT  8397.5 55917.5 8462.5 56052.5 ;
      RECT  8207.5 55917.5 8272.5 56052.5 ;
      RECT  8207.5 55032.5 8272.5 55167.5 ;
      RECT  8397.5 55032.5 8462.5 55167.5 ;
      RECT  8397.5 55032.5 8462.5 55167.5 ;
      RECT  8207.5 55032.5 8272.5 55167.5 ;
      RECT  8567.5 56007.5 8632.5 56142.5 ;
      RECT  8567.5 55032.5 8632.5 55167.5 ;
      RECT  8265.0 55475.0 8330.0 55610.0 ;
      RECT  8265.0 55475.0 8330.0 55610.0 ;
      RECT  8430.0 55510.0 8495.0 55575.0 ;
      RECT  8140.0 56227.5 8700.0 56292.5 ;
      RECT  8140.0 54882.5 8700.0 54947.5 ;
      RECT  8567.5 56445.0 8632.5 56260.0 ;
      RECT  8567.5 57605.0 8632.5 57420.0 ;
      RECT  8207.5 57487.5 8272.5 57637.5 ;
      RECT  8207.5 56602.5 8272.5 56227.5 ;
      RECT  8397.5 57487.5 8462.5 56602.5 ;
      RECT  8207.5 56602.5 8272.5 56467.5 ;
      RECT  8397.5 56602.5 8462.5 56467.5 ;
      RECT  8397.5 56602.5 8462.5 56467.5 ;
      RECT  8207.5 56602.5 8272.5 56467.5 ;
      RECT  8207.5 57487.5 8272.5 57352.5 ;
      RECT  8397.5 57487.5 8462.5 57352.5 ;
      RECT  8397.5 57487.5 8462.5 57352.5 ;
      RECT  8207.5 57487.5 8272.5 57352.5 ;
      RECT  8567.5 56512.5 8632.5 56377.5 ;
      RECT  8567.5 57487.5 8632.5 57352.5 ;
      RECT  8265.0 57045.0 8330.0 56910.0 ;
      RECT  8265.0 57045.0 8330.0 56910.0 ;
      RECT  8430.0 57010.0 8495.0 56945.0 ;
      RECT  8140.0 56292.5 8700.0 56227.5 ;
      RECT  8140.0 57637.5 8700.0 57572.5 ;
      RECT  8567.5 58765.0 8632.5 58950.0 ;
      RECT  8567.5 57605.0 8632.5 57790.0 ;
      RECT  8207.5 57722.5 8272.5 57572.5 ;
      RECT  8207.5 58607.5 8272.5 58982.5 ;
      RECT  8397.5 57722.5 8462.5 58607.5 ;
      RECT  8207.5 58607.5 8272.5 58742.5 ;
      RECT  8397.5 58607.5 8462.5 58742.5 ;
      RECT  8397.5 58607.5 8462.5 58742.5 ;
      RECT  8207.5 58607.5 8272.5 58742.5 ;
      RECT  8207.5 57722.5 8272.5 57857.5 ;
      RECT  8397.5 57722.5 8462.5 57857.5 ;
      RECT  8397.5 57722.5 8462.5 57857.5 ;
      RECT  8207.5 57722.5 8272.5 57857.5 ;
      RECT  8567.5 58697.5 8632.5 58832.5 ;
      RECT  8567.5 57722.5 8632.5 57857.5 ;
      RECT  8265.0 58165.0 8330.0 58300.0 ;
      RECT  8265.0 58165.0 8330.0 58300.0 ;
      RECT  8430.0 58200.0 8495.0 58265.0 ;
      RECT  8140.0 58917.5 8700.0 58982.5 ;
      RECT  8140.0 57572.5 8700.0 57637.5 ;
      RECT  8567.5 59135.0 8632.5 58950.0 ;
      RECT  8567.5 60295.0 8632.5 60110.0 ;
      RECT  8207.5 60177.5 8272.5 60327.5 ;
      RECT  8207.5 59292.5 8272.5 58917.5 ;
      RECT  8397.5 60177.5 8462.5 59292.5 ;
      RECT  8207.5 59292.5 8272.5 59157.5 ;
      RECT  8397.5 59292.5 8462.5 59157.5 ;
      RECT  8397.5 59292.5 8462.5 59157.5 ;
      RECT  8207.5 59292.5 8272.5 59157.5 ;
      RECT  8207.5 60177.5 8272.5 60042.5 ;
      RECT  8397.5 60177.5 8462.5 60042.5 ;
      RECT  8397.5 60177.5 8462.5 60042.5 ;
      RECT  8207.5 60177.5 8272.5 60042.5 ;
      RECT  8567.5 59202.5 8632.5 59067.5 ;
      RECT  8567.5 60177.5 8632.5 60042.5 ;
      RECT  8265.0 59735.0 8330.0 59600.0 ;
      RECT  8265.0 59735.0 8330.0 59600.0 ;
      RECT  8430.0 59700.0 8495.0 59635.0 ;
      RECT  8140.0 58982.5 8700.0 58917.5 ;
      RECT  8140.0 60327.5 8700.0 60262.5 ;
      RECT  8567.5 61455.0 8632.5 61640.0 ;
      RECT  8567.5 60295.0 8632.5 60480.0 ;
      RECT  8207.5 60412.5 8272.5 60262.5 ;
      RECT  8207.5 61297.5 8272.5 61672.5 ;
      RECT  8397.5 60412.5 8462.5 61297.5 ;
      RECT  8207.5 61297.5 8272.5 61432.5 ;
      RECT  8397.5 61297.5 8462.5 61432.5 ;
      RECT  8397.5 61297.5 8462.5 61432.5 ;
      RECT  8207.5 61297.5 8272.5 61432.5 ;
      RECT  8207.5 60412.5 8272.5 60547.5 ;
      RECT  8397.5 60412.5 8462.5 60547.5 ;
      RECT  8397.5 60412.5 8462.5 60547.5 ;
      RECT  8207.5 60412.5 8272.5 60547.5 ;
      RECT  8567.5 61387.5 8632.5 61522.5 ;
      RECT  8567.5 60412.5 8632.5 60547.5 ;
      RECT  8265.0 60855.0 8330.0 60990.0 ;
      RECT  8265.0 60855.0 8330.0 60990.0 ;
      RECT  8430.0 60890.0 8495.0 60955.0 ;
      RECT  8140.0 61607.5 8700.0 61672.5 ;
      RECT  8140.0 60262.5 8700.0 60327.5 ;
      RECT  8567.5 61825.0 8632.5 61640.0 ;
      RECT  8567.5 62985.0 8632.5 62800.0 ;
      RECT  8207.5 62867.5 8272.5 63017.5 ;
      RECT  8207.5 61982.5 8272.5 61607.5 ;
      RECT  8397.5 62867.5 8462.5 61982.5 ;
      RECT  8207.5 61982.5 8272.5 61847.5 ;
      RECT  8397.5 61982.5 8462.5 61847.5 ;
      RECT  8397.5 61982.5 8462.5 61847.5 ;
      RECT  8207.5 61982.5 8272.5 61847.5 ;
      RECT  8207.5 62867.5 8272.5 62732.5 ;
      RECT  8397.5 62867.5 8462.5 62732.5 ;
      RECT  8397.5 62867.5 8462.5 62732.5 ;
      RECT  8207.5 62867.5 8272.5 62732.5 ;
      RECT  8567.5 61892.5 8632.5 61757.5 ;
      RECT  8567.5 62867.5 8632.5 62732.5 ;
      RECT  8265.0 62425.0 8330.0 62290.0 ;
      RECT  8265.0 62425.0 8330.0 62290.0 ;
      RECT  8430.0 62390.0 8495.0 62325.0 ;
      RECT  8140.0 61672.5 8700.0 61607.5 ;
      RECT  8140.0 63017.5 8700.0 62952.5 ;
      RECT  8567.5 64145.0 8632.5 64330.0 ;
      RECT  8567.5 62985.0 8632.5 63170.0 ;
      RECT  8207.5 63102.5 8272.5 62952.5 ;
      RECT  8207.5 63987.5 8272.5 64362.5 ;
      RECT  8397.5 63102.5 8462.5 63987.5 ;
      RECT  8207.5 63987.5 8272.5 64122.5 ;
      RECT  8397.5 63987.5 8462.5 64122.5 ;
      RECT  8397.5 63987.5 8462.5 64122.5 ;
      RECT  8207.5 63987.5 8272.5 64122.5 ;
      RECT  8207.5 63102.5 8272.5 63237.5 ;
      RECT  8397.5 63102.5 8462.5 63237.5 ;
      RECT  8397.5 63102.5 8462.5 63237.5 ;
      RECT  8207.5 63102.5 8272.5 63237.5 ;
      RECT  8567.5 64077.5 8632.5 64212.5 ;
      RECT  8567.5 63102.5 8632.5 63237.5 ;
      RECT  8265.0 63545.0 8330.0 63680.0 ;
      RECT  8265.0 63545.0 8330.0 63680.0 ;
      RECT  8430.0 63580.0 8495.0 63645.0 ;
      RECT  8140.0 64297.5 8700.0 64362.5 ;
      RECT  8140.0 62952.5 8700.0 63017.5 ;
      RECT  8567.5 64515.0 8632.5 64330.0 ;
      RECT  8567.5 65675.0 8632.5 65490.0 ;
      RECT  8207.5 65557.5 8272.5 65707.5 ;
      RECT  8207.5 64672.5 8272.5 64297.5 ;
      RECT  8397.5 65557.5 8462.5 64672.5 ;
      RECT  8207.5 64672.5 8272.5 64537.5 ;
      RECT  8397.5 64672.5 8462.5 64537.5 ;
      RECT  8397.5 64672.5 8462.5 64537.5 ;
      RECT  8207.5 64672.5 8272.5 64537.5 ;
      RECT  8207.5 65557.5 8272.5 65422.5 ;
      RECT  8397.5 65557.5 8462.5 65422.5 ;
      RECT  8397.5 65557.5 8462.5 65422.5 ;
      RECT  8207.5 65557.5 8272.5 65422.5 ;
      RECT  8567.5 64582.5 8632.5 64447.5 ;
      RECT  8567.5 65557.5 8632.5 65422.5 ;
      RECT  8265.0 65115.0 8330.0 64980.0 ;
      RECT  8265.0 65115.0 8330.0 64980.0 ;
      RECT  8430.0 65080.0 8495.0 65015.0 ;
      RECT  8140.0 64362.5 8700.0 64297.5 ;
      RECT  8140.0 65707.5 8700.0 65642.5 ;
      RECT  8567.5 66835.0 8632.5 67020.0 ;
      RECT  8567.5 65675.0 8632.5 65860.0 ;
      RECT  8207.5 65792.5 8272.5 65642.5 ;
      RECT  8207.5 66677.5 8272.5 67052.5 ;
      RECT  8397.5 65792.5 8462.5 66677.5 ;
      RECT  8207.5 66677.5 8272.5 66812.5 ;
      RECT  8397.5 66677.5 8462.5 66812.5 ;
      RECT  8397.5 66677.5 8462.5 66812.5 ;
      RECT  8207.5 66677.5 8272.5 66812.5 ;
      RECT  8207.5 65792.5 8272.5 65927.5 ;
      RECT  8397.5 65792.5 8462.5 65927.5 ;
      RECT  8397.5 65792.5 8462.5 65927.5 ;
      RECT  8207.5 65792.5 8272.5 65927.5 ;
      RECT  8567.5 66767.5 8632.5 66902.5 ;
      RECT  8567.5 65792.5 8632.5 65927.5 ;
      RECT  8265.0 66235.0 8330.0 66370.0 ;
      RECT  8265.0 66235.0 8330.0 66370.0 ;
      RECT  8430.0 66270.0 8495.0 66335.0 ;
      RECT  8140.0 66987.5 8700.0 67052.5 ;
      RECT  8140.0 65642.5 8700.0 65707.5 ;
      RECT  8567.5 67205.0 8632.5 67020.0 ;
      RECT  8567.5 68365.0 8632.5 68180.0 ;
      RECT  8207.5 68247.5 8272.5 68397.5 ;
      RECT  8207.5 67362.5 8272.5 66987.5 ;
      RECT  8397.5 68247.5 8462.5 67362.5 ;
      RECT  8207.5 67362.5 8272.5 67227.5 ;
      RECT  8397.5 67362.5 8462.5 67227.5 ;
      RECT  8397.5 67362.5 8462.5 67227.5 ;
      RECT  8207.5 67362.5 8272.5 67227.5 ;
      RECT  8207.5 68247.5 8272.5 68112.5 ;
      RECT  8397.5 68247.5 8462.5 68112.5 ;
      RECT  8397.5 68247.5 8462.5 68112.5 ;
      RECT  8207.5 68247.5 8272.5 68112.5 ;
      RECT  8567.5 67272.5 8632.5 67137.5 ;
      RECT  8567.5 68247.5 8632.5 68112.5 ;
      RECT  8265.0 67805.0 8330.0 67670.0 ;
      RECT  8265.0 67805.0 8330.0 67670.0 ;
      RECT  8430.0 67770.0 8495.0 67705.0 ;
      RECT  8140.0 67052.5 8700.0 66987.5 ;
      RECT  8140.0 68397.5 8700.0 68332.5 ;
      RECT  8567.5 69525.0 8632.5 69710.0 ;
      RECT  8567.5 68365.0 8632.5 68550.0 ;
      RECT  8207.5 68482.5 8272.5 68332.5 ;
      RECT  8207.5 69367.5 8272.5 69742.5 ;
      RECT  8397.5 68482.5 8462.5 69367.5 ;
      RECT  8207.5 69367.5 8272.5 69502.5 ;
      RECT  8397.5 69367.5 8462.5 69502.5 ;
      RECT  8397.5 69367.5 8462.5 69502.5 ;
      RECT  8207.5 69367.5 8272.5 69502.5 ;
      RECT  8207.5 68482.5 8272.5 68617.5 ;
      RECT  8397.5 68482.5 8462.5 68617.5 ;
      RECT  8397.5 68482.5 8462.5 68617.5 ;
      RECT  8207.5 68482.5 8272.5 68617.5 ;
      RECT  8567.5 69457.5 8632.5 69592.5 ;
      RECT  8567.5 68482.5 8632.5 68617.5 ;
      RECT  8265.0 68925.0 8330.0 69060.0 ;
      RECT  8265.0 68925.0 8330.0 69060.0 ;
      RECT  8430.0 68960.0 8495.0 69025.0 ;
      RECT  8140.0 69677.5 8700.0 69742.5 ;
      RECT  8140.0 68332.5 8700.0 68397.5 ;
      RECT  8567.5 69895.0 8632.5 69710.0 ;
      RECT  8567.5 71055.0 8632.5 70870.0 ;
      RECT  8207.5 70937.5 8272.5 71087.5 ;
      RECT  8207.5 70052.5 8272.5 69677.5 ;
      RECT  8397.5 70937.5 8462.5 70052.5 ;
      RECT  8207.5 70052.5 8272.5 69917.5 ;
      RECT  8397.5 70052.5 8462.5 69917.5 ;
      RECT  8397.5 70052.5 8462.5 69917.5 ;
      RECT  8207.5 70052.5 8272.5 69917.5 ;
      RECT  8207.5 70937.5 8272.5 70802.5 ;
      RECT  8397.5 70937.5 8462.5 70802.5 ;
      RECT  8397.5 70937.5 8462.5 70802.5 ;
      RECT  8207.5 70937.5 8272.5 70802.5 ;
      RECT  8567.5 69962.5 8632.5 69827.5 ;
      RECT  8567.5 70937.5 8632.5 70802.5 ;
      RECT  8265.0 70495.0 8330.0 70360.0 ;
      RECT  8265.0 70495.0 8330.0 70360.0 ;
      RECT  8430.0 70460.0 8495.0 70395.0 ;
      RECT  8140.0 69742.5 8700.0 69677.5 ;
      RECT  8140.0 71087.5 8700.0 71022.5 ;
      RECT  8567.5 72215.0 8632.5 72400.0 ;
      RECT  8567.5 71055.0 8632.5 71240.0 ;
      RECT  8207.5 71172.5 8272.5 71022.5 ;
      RECT  8207.5 72057.5 8272.5 72432.5 ;
      RECT  8397.5 71172.5 8462.5 72057.5 ;
      RECT  8207.5 72057.5 8272.5 72192.5 ;
      RECT  8397.5 72057.5 8462.5 72192.5 ;
      RECT  8397.5 72057.5 8462.5 72192.5 ;
      RECT  8207.5 72057.5 8272.5 72192.5 ;
      RECT  8207.5 71172.5 8272.5 71307.5 ;
      RECT  8397.5 71172.5 8462.5 71307.5 ;
      RECT  8397.5 71172.5 8462.5 71307.5 ;
      RECT  8207.5 71172.5 8272.5 71307.5 ;
      RECT  8567.5 72147.5 8632.5 72282.5 ;
      RECT  8567.5 71172.5 8632.5 71307.5 ;
      RECT  8265.0 71615.0 8330.0 71750.0 ;
      RECT  8265.0 71615.0 8330.0 71750.0 ;
      RECT  8430.0 71650.0 8495.0 71715.0 ;
      RECT  8140.0 72367.5 8700.0 72432.5 ;
      RECT  8140.0 71022.5 8700.0 71087.5 ;
      RECT  8567.5 72585.0 8632.5 72400.0 ;
      RECT  8567.5 73745.0 8632.5 73560.0 ;
      RECT  8207.5 73627.5 8272.5 73777.5 ;
      RECT  8207.5 72742.5 8272.5 72367.5 ;
      RECT  8397.5 73627.5 8462.5 72742.5 ;
      RECT  8207.5 72742.5 8272.5 72607.5 ;
      RECT  8397.5 72742.5 8462.5 72607.5 ;
      RECT  8397.5 72742.5 8462.5 72607.5 ;
      RECT  8207.5 72742.5 8272.5 72607.5 ;
      RECT  8207.5 73627.5 8272.5 73492.5 ;
      RECT  8397.5 73627.5 8462.5 73492.5 ;
      RECT  8397.5 73627.5 8462.5 73492.5 ;
      RECT  8207.5 73627.5 8272.5 73492.5 ;
      RECT  8567.5 72652.5 8632.5 72517.5 ;
      RECT  8567.5 73627.5 8632.5 73492.5 ;
      RECT  8265.0 73185.0 8330.0 73050.0 ;
      RECT  8265.0 73185.0 8330.0 73050.0 ;
      RECT  8430.0 73150.0 8495.0 73085.0 ;
      RECT  8140.0 72432.5 8700.0 72367.5 ;
      RECT  8140.0 73777.5 8700.0 73712.5 ;
      RECT  8567.5 74905.0 8632.5 75090.0 ;
      RECT  8567.5 73745.0 8632.5 73930.0 ;
      RECT  8207.5 73862.5 8272.5 73712.5 ;
      RECT  8207.5 74747.5 8272.5 75122.5 ;
      RECT  8397.5 73862.5 8462.5 74747.5 ;
      RECT  8207.5 74747.5 8272.5 74882.5 ;
      RECT  8397.5 74747.5 8462.5 74882.5 ;
      RECT  8397.5 74747.5 8462.5 74882.5 ;
      RECT  8207.5 74747.5 8272.5 74882.5 ;
      RECT  8207.5 73862.5 8272.5 73997.5 ;
      RECT  8397.5 73862.5 8462.5 73997.5 ;
      RECT  8397.5 73862.5 8462.5 73997.5 ;
      RECT  8207.5 73862.5 8272.5 73997.5 ;
      RECT  8567.5 74837.5 8632.5 74972.5 ;
      RECT  8567.5 73862.5 8632.5 73997.5 ;
      RECT  8265.0 74305.0 8330.0 74440.0 ;
      RECT  8265.0 74305.0 8330.0 74440.0 ;
      RECT  8430.0 74340.0 8495.0 74405.0 ;
      RECT  8140.0 75057.5 8700.0 75122.5 ;
      RECT  8140.0 73712.5 8700.0 73777.5 ;
      RECT  8567.5 75275.0 8632.5 75090.0 ;
      RECT  8567.5 76435.0 8632.5 76250.0 ;
      RECT  8207.5 76317.5 8272.5 76467.5 ;
      RECT  8207.5 75432.5 8272.5 75057.5 ;
      RECT  8397.5 76317.5 8462.5 75432.5 ;
      RECT  8207.5 75432.5 8272.5 75297.5 ;
      RECT  8397.5 75432.5 8462.5 75297.5 ;
      RECT  8397.5 75432.5 8462.5 75297.5 ;
      RECT  8207.5 75432.5 8272.5 75297.5 ;
      RECT  8207.5 76317.5 8272.5 76182.5 ;
      RECT  8397.5 76317.5 8462.5 76182.5 ;
      RECT  8397.5 76317.5 8462.5 76182.5 ;
      RECT  8207.5 76317.5 8272.5 76182.5 ;
      RECT  8567.5 75342.5 8632.5 75207.5 ;
      RECT  8567.5 76317.5 8632.5 76182.5 ;
      RECT  8265.0 75875.0 8330.0 75740.0 ;
      RECT  8265.0 75875.0 8330.0 75740.0 ;
      RECT  8430.0 75840.0 8495.0 75775.0 ;
      RECT  8140.0 75122.5 8700.0 75057.5 ;
      RECT  8140.0 76467.5 8700.0 76402.5 ;
      RECT  8567.5 77595.0 8632.5 77780.0 ;
      RECT  8567.5 76435.0 8632.5 76620.0 ;
      RECT  8207.5 76552.5 8272.5 76402.5 ;
      RECT  8207.5 77437.5 8272.5 77812.5 ;
      RECT  8397.5 76552.5 8462.5 77437.5 ;
      RECT  8207.5 77437.5 8272.5 77572.5 ;
      RECT  8397.5 77437.5 8462.5 77572.5 ;
      RECT  8397.5 77437.5 8462.5 77572.5 ;
      RECT  8207.5 77437.5 8272.5 77572.5 ;
      RECT  8207.5 76552.5 8272.5 76687.5 ;
      RECT  8397.5 76552.5 8462.5 76687.5 ;
      RECT  8397.5 76552.5 8462.5 76687.5 ;
      RECT  8207.5 76552.5 8272.5 76687.5 ;
      RECT  8567.5 77527.5 8632.5 77662.5 ;
      RECT  8567.5 76552.5 8632.5 76687.5 ;
      RECT  8265.0 76995.0 8330.0 77130.0 ;
      RECT  8265.0 76995.0 8330.0 77130.0 ;
      RECT  8430.0 77030.0 8495.0 77095.0 ;
      RECT  8140.0 77747.5 8700.0 77812.5 ;
      RECT  8140.0 76402.5 8700.0 76467.5 ;
      RECT  8567.5 77965.0 8632.5 77780.0 ;
      RECT  8567.5 79125.0 8632.5 78940.0 ;
      RECT  8207.5 79007.5 8272.5 79157.5 ;
      RECT  8207.5 78122.5 8272.5 77747.5 ;
      RECT  8397.5 79007.5 8462.5 78122.5 ;
      RECT  8207.5 78122.5 8272.5 77987.5 ;
      RECT  8397.5 78122.5 8462.5 77987.5 ;
      RECT  8397.5 78122.5 8462.5 77987.5 ;
      RECT  8207.5 78122.5 8272.5 77987.5 ;
      RECT  8207.5 79007.5 8272.5 78872.5 ;
      RECT  8397.5 79007.5 8462.5 78872.5 ;
      RECT  8397.5 79007.5 8462.5 78872.5 ;
      RECT  8207.5 79007.5 8272.5 78872.5 ;
      RECT  8567.5 78032.5 8632.5 77897.5 ;
      RECT  8567.5 79007.5 8632.5 78872.5 ;
      RECT  8265.0 78565.0 8330.0 78430.0 ;
      RECT  8265.0 78565.0 8330.0 78430.0 ;
      RECT  8430.0 78530.0 8495.0 78465.0 ;
      RECT  8140.0 77812.5 8700.0 77747.5 ;
      RECT  8140.0 79157.5 8700.0 79092.5 ;
      RECT  8567.5 80285.0 8632.5 80470.0 ;
      RECT  8567.5 79125.0 8632.5 79310.0 ;
      RECT  8207.5 79242.5 8272.5 79092.5 ;
      RECT  8207.5 80127.5 8272.5 80502.5 ;
      RECT  8397.5 79242.5 8462.5 80127.5 ;
      RECT  8207.5 80127.5 8272.5 80262.5 ;
      RECT  8397.5 80127.5 8462.5 80262.5 ;
      RECT  8397.5 80127.5 8462.5 80262.5 ;
      RECT  8207.5 80127.5 8272.5 80262.5 ;
      RECT  8207.5 79242.5 8272.5 79377.5 ;
      RECT  8397.5 79242.5 8462.5 79377.5 ;
      RECT  8397.5 79242.5 8462.5 79377.5 ;
      RECT  8207.5 79242.5 8272.5 79377.5 ;
      RECT  8567.5 80217.5 8632.5 80352.5 ;
      RECT  8567.5 79242.5 8632.5 79377.5 ;
      RECT  8265.0 79685.0 8330.0 79820.0 ;
      RECT  8265.0 79685.0 8330.0 79820.0 ;
      RECT  8430.0 79720.0 8495.0 79785.0 ;
      RECT  8140.0 80437.5 8700.0 80502.5 ;
      RECT  8140.0 79092.5 8700.0 79157.5 ;
      RECT  8567.5 80655.0 8632.5 80470.0 ;
      RECT  8567.5 81815.0 8632.5 81630.0 ;
      RECT  8207.5 81697.5 8272.5 81847.5 ;
      RECT  8207.5 80812.5 8272.5 80437.5 ;
      RECT  8397.5 81697.5 8462.5 80812.5 ;
      RECT  8207.5 80812.5 8272.5 80677.5 ;
      RECT  8397.5 80812.5 8462.5 80677.5 ;
      RECT  8397.5 80812.5 8462.5 80677.5 ;
      RECT  8207.5 80812.5 8272.5 80677.5 ;
      RECT  8207.5 81697.5 8272.5 81562.5 ;
      RECT  8397.5 81697.5 8462.5 81562.5 ;
      RECT  8397.5 81697.5 8462.5 81562.5 ;
      RECT  8207.5 81697.5 8272.5 81562.5 ;
      RECT  8567.5 80722.5 8632.5 80587.5 ;
      RECT  8567.5 81697.5 8632.5 81562.5 ;
      RECT  8265.0 81255.0 8330.0 81120.0 ;
      RECT  8265.0 81255.0 8330.0 81120.0 ;
      RECT  8430.0 81220.0 8495.0 81155.0 ;
      RECT  8140.0 80502.5 8700.0 80437.5 ;
      RECT  8140.0 81847.5 8700.0 81782.5 ;
      RECT  8567.5 82975.0 8632.5 83160.0 ;
      RECT  8567.5 81815.0 8632.5 82000.0 ;
      RECT  8207.5 81932.5 8272.5 81782.5 ;
      RECT  8207.5 82817.5 8272.5 83192.5 ;
      RECT  8397.5 81932.5 8462.5 82817.5 ;
      RECT  8207.5 82817.5 8272.5 82952.5 ;
      RECT  8397.5 82817.5 8462.5 82952.5 ;
      RECT  8397.5 82817.5 8462.5 82952.5 ;
      RECT  8207.5 82817.5 8272.5 82952.5 ;
      RECT  8207.5 81932.5 8272.5 82067.5 ;
      RECT  8397.5 81932.5 8462.5 82067.5 ;
      RECT  8397.5 81932.5 8462.5 82067.5 ;
      RECT  8207.5 81932.5 8272.5 82067.5 ;
      RECT  8567.5 82907.5 8632.5 83042.5 ;
      RECT  8567.5 81932.5 8632.5 82067.5 ;
      RECT  8265.0 82375.0 8330.0 82510.0 ;
      RECT  8265.0 82375.0 8330.0 82510.0 ;
      RECT  8430.0 82410.0 8495.0 82475.0 ;
      RECT  8140.0 83127.5 8700.0 83192.5 ;
      RECT  8140.0 81782.5 8700.0 81847.5 ;
      RECT  8567.5 83345.0 8632.5 83160.0 ;
      RECT  8567.5 84505.0 8632.5 84320.0 ;
      RECT  8207.5 84387.5 8272.5 84537.5 ;
      RECT  8207.5 83502.5 8272.5 83127.5 ;
      RECT  8397.5 84387.5 8462.5 83502.5 ;
      RECT  8207.5 83502.5 8272.5 83367.5 ;
      RECT  8397.5 83502.5 8462.5 83367.5 ;
      RECT  8397.5 83502.5 8462.5 83367.5 ;
      RECT  8207.5 83502.5 8272.5 83367.5 ;
      RECT  8207.5 84387.5 8272.5 84252.5 ;
      RECT  8397.5 84387.5 8462.5 84252.5 ;
      RECT  8397.5 84387.5 8462.5 84252.5 ;
      RECT  8207.5 84387.5 8272.5 84252.5 ;
      RECT  8567.5 83412.5 8632.5 83277.5 ;
      RECT  8567.5 84387.5 8632.5 84252.5 ;
      RECT  8265.0 83945.0 8330.0 83810.0 ;
      RECT  8265.0 83945.0 8330.0 83810.0 ;
      RECT  8430.0 83910.0 8495.0 83845.0 ;
      RECT  8140.0 83192.5 8700.0 83127.5 ;
      RECT  8140.0 84537.5 8700.0 84472.5 ;
      RECT  8567.5 85665.0 8632.5 85850.0 ;
      RECT  8567.5 84505.0 8632.5 84690.0 ;
      RECT  8207.5 84622.5 8272.5 84472.5 ;
      RECT  8207.5 85507.5 8272.5 85882.5 ;
      RECT  8397.5 84622.5 8462.5 85507.5 ;
      RECT  8207.5 85507.5 8272.5 85642.5 ;
      RECT  8397.5 85507.5 8462.5 85642.5 ;
      RECT  8397.5 85507.5 8462.5 85642.5 ;
      RECT  8207.5 85507.5 8272.5 85642.5 ;
      RECT  8207.5 84622.5 8272.5 84757.5 ;
      RECT  8397.5 84622.5 8462.5 84757.5 ;
      RECT  8397.5 84622.5 8462.5 84757.5 ;
      RECT  8207.5 84622.5 8272.5 84757.5 ;
      RECT  8567.5 85597.5 8632.5 85732.5 ;
      RECT  8567.5 84622.5 8632.5 84757.5 ;
      RECT  8265.0 85065.0 8330.0 85200.0 ;
      RECT  8265.0 85065.0 8330.0 85200.0 ;
      RECT  8430.0 85100.0 8495.0 85165.0 ;
      RECT  8140.0 85817.5 8700.0 85882.5 ;
      RECT  8140.0 84472.5 8700.0 84537.5 ;
      RECT  8567.5 86035.0 8632.5 85850.0 ;
      RECT  8567.5 87195.0 8632.5 87010.0 ;
      RECT  8207.5 87077.5 8272.5 87227.5 ;
      RECT  8207.5 86192.5 8272.5 85817.5 ;
      RECT  8397.5 87077.5 8462.5 86192.5 ;
      RECT  8207.5 86192.5 8272.5 86057.5 ;
      RECT  8397.5 86192.5 8462.5 86057.5 ;
      RECT  8397.5 86192.5 8462.5 86057.5 ;
      RECT  8207.5 86192.5 8272.5 86057.5 ;
      RECT  8207.5 87077.5 8272.5 86942.5 ;
      RECT  8397.5 87077.5 8462.5 86942.5 ;
      RECT  8397.5 87077.5 8462.5 86942.5 ;
      RECT  8207.5 87077.5 8272.5 86942.5 ;
      RECT  8567.5 86102.5 8632.5 85967.5 ;
      RECT  8567.5 87077.5 8632.5 86942.5 ;
      RECT  8265.0 86635.0 8330.0 86500.0 ;
      RECT  8265.0 86635.0 8330.0 86500.0 ;
      RECT  8430.0 86600.0 8495.0 86535.0 ;
      RECT  8140.0 85882.5 8700.0 85817.5 ;
      RECT  8140.0 87227.5 8700.0 87162.5 ;
      RECT  8567.5 88355.0 8632.5 88540.0 ;
      RECT  8567.5 87195.0 8632.5 87380.0 ;
      RECT  8207.5 87312.5 8272.5 87162.5 ;
      RECT  8207.5 88197.5 8272.5 88572.5 ;
      RECT  8397.5 87312.5 8462.5 88197.5 ;
      RECT  8207.5 88197.5 8272.5 88332.5 ;
      RECT  8397.5 88197.5 8462.5 88332.5 ;
      RECT  8397.5 88197.5 8462.5 88332.5 ;
      RECT  8207.5 88197.5 8272.5 88332.5 ;
      RECT  8207.5 87312.5 8272.5 87447.5 ;
      RECT  8397.5 87312.5 8462.5 87447.5 ;
      RECT  8397.5 87312.5 8462.5 87447.5 ;
      RECT  8207.5 87312.5 8272.5 87447.5 ;
      RECT  8567.5 88287.5 8632.5 88422.5 ;
      RECT  8567.5 87312.5 8632.5 87447.5 ;
      RECT  8265.0 87755.0 8330.0 87890.0 ;
      RECT  8265.0 87755.0 8330.0 87890.0 ;
      RECT  8430.0 87790.0 8495.0 87855.0 ;
      RECT  8140.0 88507.5 8700.0 88572.5 ;
      RECT  8140.0 87162.5 8700.0 87227.5 ;
      RECT  8567.5 88725.0 8632.5 88540.0 ;
      RECT  8567.5 89885.0 8632.5 89700.0 ;
      RECT  8207.5 89767.5 8272.5 89917.5 ;
      RECT  8207.5 88882.5 8272.5 88507.5 ;
      RECT  8397.5 89767.5 8462.5 88882.5 ;
      RECT  8207.5 88882.5 8272.5 88747.5 ;
      RECT  8397.5 88882.5 8462.5 88747.5 ;
      RECT  8397.5 88882.5 8462.5 88747.5 ;
      RECT  8207.5 88882.5 8272.5 88747.5 ;
      RECT  8207.5 89767.5 8272.5 89632.5 ;
      RECT  8397.5 89767.5 8462.5 89632.5 ;
      RECT  8397.5 89767.5 8462.5 89632.5 ;
      RECT  8207.5 89767.5 8272.5 89632.5 ;
      RECT  8567.5 88792.5 8632.5 88657.5 ;
      RECT  8567.5 89767.5 8632.5 89632.5 ;
      RECT  8265.0 89325.0 8330.0 89190.0 ;
      RECT  8265.0 89325.0 8330.0 89190.0 ;
      RECT  8430.0 89290.0 8495.0 89225.0 ;
      RECT  8140.0 88572.5 8700.0 88507.5 ;
      RECT  8140.0 89917.5 8700.0 89852.5 ;
      RECT  8567.5 91045.0 8632.5 91230.0 ;
      RECT  8567.5 89885.0 8632.5 90070.0 ;
      RECT  8207.5 90002.5 8272.5 89852.5 ;
      RECT  8207.5 90887.5 8272.5 91262.5 ;
      RECT  8397.5 90002.5 8462.5 90887.5 ;
      RECT  8207.5 90887.5 8272.5 91022.5 ;
      RECT  8397.5 90887.5 8462.5 91022.5 ;
      RECT  8397.5 90887.5 8462.5 91022.5 ;
      RECT  8207.5 90887.5 8272.5 91022.5 ;
      RECT  8207.5 90002.5 8272.5 90137.5 ;
      RECT  8397.5 90002.5 8462.5 90137.5 ;
      RECT  8397.5 90002.5 8462.5 90137.5 ;
      RECT  8207.5 90002.5 8272.5 90137.5 ;
      RECT  8567.5 90977.5 8632.5 91112.5 ;
      RECT  8567.5 90002.5 8632.5 90137.5 ;
      RECT  8265.0 90445.0 8330.0 90580.0 ;
      RECT  8265.0 90445.0 8330.0 90580.0 ;
      RECT  8430.0 90480.0 8495.0 90545.0 ;
      RECT  8140.0 91197.5 8700.0 91262.5 ;
      RECT  8140.0 89852.5 8700.0 89917.5 ;
      RECT  8567.5 91415.0 8632.5 91230.0 ;
      RECT  8567.5 92575.0 8632.5 92390.0 ;
      RECT  8207.5 92457.5 8272.5 92607.5 ;
      RECT  8207.5 91572.5 8272.5 91197.5 ;
      RECT  8397.5 92457.5 8462.5 91572.5 ;
      RECT  8207.5 91572.5 8272.5 91437.5 ;
      RECT  8397.5 91572.5 8462.5 91437.5 ;
      RECT  8397.5 91572.5 8462.5 91437.5 ;
      RECT  8207.5 91572.5 8272.5 91437.5 ;
      RECT  8207.5 92457.5 8272.5 92322.5 ;
      RECT  8397.5 92457.5 8462.5 92322.5 ;
      RECT  8397.5 92457.5 8462.5 92322.5 ;
      RECT  8207.5 92457.5 8272.5 92322.5 ;
      RECT  8567.5 91482.5 8632.5 91347.5 ;
      RECT  8567.5 92457.5 8632.5 92322.5 ;
      RECT  8265.0 92015.0 8330.0 91880.0 ;
      RECT  8265.0 92015.0 8330.0 91880.0 ;
      RECT  8430.0 91980.0 8495.0 91915.0 ;
      RECT  8140.0 91262.5 8700.0 91197.5 ;
      RECT  8140.0 92607.5 8700.0 92542.5 ;
      RECT  8567.5 93735.0 8632.5 93920.0 ;
      RECT  8567.5 92575.0 8632.5 92760.0 ;
      RECT  8207.5 92692.5 8272.5 92542.5 ;
      RECT  8207.5 93577.5 8272.5 93952.5 ;
      RECT  8397.5 92692.5 8462.5 93577.5 ;
      RECT  8207.5 93577.5 8272.5 93712.5 ;
      RECT  8397.5 93577.5 8462.5 93712.5 ;
      RECT  8397.5 93577.5 8462.5 93712.5 ;
      RECT  8207.5 93577.5 8272.5 93712.5 ;
      RECT  8207.5 92692.5 8272.5 92827.5 ;
      RECT  8397.5 92692.5 8462.5 92827.5 ;
      RECT  8397.5 92692.5 8462.5 92827.5 ;
      RECT  8207.5 92692.5 8272.5 92827.5 ;
      RECT  8567.5 93667.5 8632.5 93802.5 ;
      RECT  8567.5 92692.5 8632.5 92827.5 ;
      RECT  8265.0 93135.0 8330.0 93270.0 ;
      RECT  8265.0 93135.0 8330.0 93270.0 ;
      RECT  8430.0 93170.0 8495.0 93235.0 ;
      RECT  8140.0 93887.5 8700.0 93952.5 ;
      RECT  8140.0 92542.5 8700.0 92607.5 ;
      RECT  8567.5 94105.0 8632.5 93920.0 ;
      RECT  8567.5 95265.0 8632.5 95080.0 ;
      RECT  8207.5 95147.5 8272.5 95297.5 ;
      RECT  8207.5 94262.5 8272.5 93887.5 ;
      RECT  8397.5 95147.5 8462.5 94262.5 ;
      RECT  8207.5 94262.5 8272.5 94127.5 ;
      RECT  8397.5 94262.5 8462.5 94127.5 ;
      RECT  8397.5 94262.5 8462.5 94127.5 ;
      RECT  8207.5 94262.5 8272.5 94127.5 ;
      RECT  8207.5 95147.5 8272.5 95012.5 ;
      RECT  8397.5 95147.5 8462.5 95012.5 ;
      RECT  8397.5 95147.5 8462.5 95012.5 ;
      RECT  8207.5 95147.5 8272.5 95012.5 ;
      RECT  8567.5 94172.5 8632.5 94037.5 ;
      RECT  8567.5 95147.5 8632.5 95012.5 ;
      RECT  8265.0 94705.0 8330.0 94570.0 ;
      RECT  8265.0 94705.0 8330.0 94570.0 ;
      RECT  8430.0 94670.0 8495.0 94605.0 ;
      RECT  8140.0 93952.5 8700.0 93887.5 ;
      RECT  8140.0 95297.5 8700.0 95232.5 ;
      RECT  8567.5 96425.0 8632.5 96610.0 ;
      RECT  8567.5 95265.0 8632.5 95450.0 ;
      RECT  8207.5 95382.5 8272.5 95232.5 ;
      RECT  8207.5 96267.5 8272.5 96642.5 ;
      RECT  8397.5 95382.5 8462.5 96267.5 ;
      RECT  8207.5 96267.5 8272.5 96402.5 ;
      RECT  8397.5 96267.5 8462.5 96402.5 ;
      RECT  8397.5 96267.5 8462.5 96402.5 ;
      RECT  8207.5 96267.5 8272.5 96402.5 ;
      RECT  8207.5 95382.5 8272.5 95517.5 ;
      RECT  8397.5 95382.5 8462.5 95517.5 ;
      RECT  8397.5 95382.5 8462.5 95517.5 ;
      RECT  8207.5 95382.5 8272.5 95517.5 ;
      RECT  8567.5 96357.5 8632.5 96492.5 ;
      RECT  8567.5 95382.5 8632.5 95517.5 ;
      RECT  8265.0 95825.0 8330.0 95960.0 ;
      RECT  8265.0 95825.0 8330.0 95960.0 ;
      RECT  8430.0 95860.0 8495.0 95925.0 ;
      RECT  8140.0 96577.5 8700.0 96642.5 ;
      RECT  8140.0 95232.5 8700.0 95297.5 ;
      RECT  8567.5 96795.0 8632.5 96610.0 ;
      RECT  8567.5 97955.0 8632.5 97770.0 ;
      RECT  8207.5 97837.5 8272.5 97987.5 ;
      RECT  8207.5 96952.5 8272.5 96577.5 ;
      RECT  8397.5 97837.5 8462.5 96952.5 ;
      RECT  8207.5 96952.5 8272.5 96817.5 ;
      RECT  8397.5 96952.5 8462.5 96817.5 ;
      RECT  8397.5 96952.5 8462.5 96817.5 ;
      RECT  8207.5 96952.5 8272.5 96817.5 ;
      RECT  8207.5 97837.5 8272.5 97702.5 ;
      RECT  8397.5 97837.5 8462.5 97702.5 ;
      RECT  8397.5 97837.5 8462.5 97702.5 ;
      RECT  8207.5 97837.5 8272.5 97702.5 ;
      RECT  8567.5 96862.5 8632.5 96727.5 ;
      RECT  8567.5 97837.5 8632.5 97702.5 ;
      RECT  8265.0 97395.0 8330.0 97260.0 ;
      RECT  8265.0 97395.0 8330.0 97260.0 ;
      RECT  8430.0 97360.0 8495.0 97295.0 ;
      RECT  8140.0 96642.5 8700.0 96577.5 ;
      RECT  8140.0 97987.5 8700.0 97922.5 ;
      RECT  8567.5 99115.0 8632.5 99300.0 ;
      RECT  8567.5 97955.0 8632.5 98140.0 ;
      RECT  8207.5 98072.5 8272.5 97922.5 ;
      RECT  8207.5 98957.5 8272.5 99332.5 ;
      RECT  8397.5 98072.5 8462.5 98957.5 ;
      RECT  8207.5 98957.5 8272.5 99092.5 ;
      RECT  8397.5 98957.5 8462.5 99092.5 ;
      RECT  8397.5 98957.5 8462.5 99092.5 ;
      RECT  8207.5 98957.5 8272.5 99092.5 ;
      RECT  8207.5 98072.5 8272.5 98207.5 ;
      RECT  8397.5 98072.5 8462.5 98207.5 ;
      RECT  8397.5 98072.5 8462.5 98207.5 ;
      RECT  8207.5 98072.5 8272.5 98207.5 ;
      RECT  8567.5 99047.5 8632.5 99182.5 ;
      RECT  8567.5 98072.5 8632.5 98207.5 ;
      RECT  8265.0 98515.0 8330.0 98650.0 ;
      RECT  8265.0 98515.0 8330.0 98650.0 ;
      RECT  8430.0 98550.0 8495.0 98615.0 ;
      RECT  8140.0 99267.5 8700.0 99332.5 ;
      RECT  8140.0 97922.5 8700.0 97987.5 ;
      RECT  8567.5 99485.0 8632.5 99300.0 ;
      RECT  8567.5 100645.0 8632.5 100460.0 ;
      RECT  8207.5 100527.5 8272.5 100677.5 ;
      RECT  8207.5 99642.5 8272.5 99267.5 ;
      RECT  8397.5 100527.5 8462.5 99642.5 ;
      RECT  8207.5 99642.5 8272.5 99507.5 ;
      RECT  8397.5 99642.5 8462.5 99507.5 ;
      RECT  8397.5 99642.5 8462.5 99507.5 ;
      RECT  8207.5 99642.5 8272.5 99507.5 ;
      RECT  8207.5 100527.5 8272.5 100392.5 ;
      RECT  8397.5 100527.5 8462.5 100392.5 ;
      RECT  8397.5 100527.5 8462.5 100392.5 ;
      RECT  8207.5 100527.5 8272.5 100392.5 ;
      RECT  8567.5 99552.5 8632.5 99417.5 ;
      RECT  8567.5 100527.5 8632.5 100392.5 ;
      RECT  8265.0 100085.0 8330.0 99950.0 ;
      RECT  8265.0 100085.0 8330.0 99950.0 ;
      RECT  8430.0 100050.0 8495.0 99985.0 ;
      RECT  8140.0 99332.5 8700.0 99267.5 ;
      RECT  8140.0 100677.5 8700.0 100612.5 ;
      RECT  8567.5 101805.0 8632.5 101990.0 ;
      RECT  8567.5 100645.0 8632.5 100830.0 ;
      RECT  8207.5 100762.5 8272.5 100612.5 ;
      RECT  8207.5 101647.5 8272.5 102022.5 ;
      RECT  8397.5 100762.5 8462.5 101647.5 ;
      RECT  8207.5 101647.5 8272.5 101782.5 ;
      RECT  8397.5 101647.5 8462.5 101782.5 ;
      RECT  8397.5 101647.5 8462.5 101782.5 ;
      RECT  8207.5 101647.5 8272.5 101782.5 ;
      RECT  8207.5 100762.5 8272.5 100897.5 ;
      RECT  8397.5 100762.5 8462.5 100897.5 ;
      RECT  8397.5 100762.5 8462.5 100897.5 ;
      RECT  8207.5 100762.5 8272.5 100897.5 ;
      RECT  8567.5 101737.5 8632.5 101872.5 ;
      RECT  8567.5 100762.5 8632.5 100897.5 ;
      RECT  8265.0 101205.0 8330.0 101340.0 ;
      RECT  8265.0 101205.0 8330.0 101340.0 ;
      RECT  8430.0 101240.0 8495.0 101305.0 ;
      RECT  8140.0 101957.5 8700.0 102022.5 ;
      RECT  8140.0 100612.5 8700.0 100677.5 ;
      RECT  8567.5 102175.0 8632.5 101990.0 ;
      RECT  8567.5 103335.0 8632.5 103150.0 ;
      RECT  8207.5 103217.5 8272.5 103367.5 ;
      RECT  8207.5 102332.5 8272.5 101957.5 ;
      RECT  8397.5 103217.5 8462.5 102332.5 ;
      RECT  8207.5 102332.5 8272.5 102197.5 ;
      RECT  8397.5 102332.5 8462.5 102197.5 ;
      RECT  8397.5 102332.5 8462.5 102197.5 ;
      RECT  8207.5 102332.5 8272.5 102197.5 ;
      RECT  8207.5 103217.5 8272.5 103082.5 ;
      RECT  8397.5 103217.5 8462.5 103082.5 ;
      RECT  8397.5 103217.5 8462.5 103082.5 ;
      RECT  8207.5 103217.5 8272.5 103082.5 ;
      RECT  8567.5 102242.5 8632.5 102107.5 ;
      RECT  8567.5 103217.5 8632.5 103082.5 ;
      RECT  8265.0 102775.0 8330.0 102640.0 ;
      RECT  8265.0 102775.0 8330.0 102640.0 ;
      RECT  8430.0 102740.0 8495.0 102675.0 ;
      RECT  8140.0 102022.5 8700.0 101957.5 ;
      RECT  8140.0 103367.5 8700.0 103302.5 ;
      RECT  8567.5 104495.0 8632.5 104680.0 ;
      RECT  8567.5 103335.0 8632.5 103520.0 ;
      RECT  8207.5 103452.5 8272.5 103302.5 ;
      RECT  8207.5 104337.5 8272.5 104712.5 ;
      RECT  8397.5 103452.5 8462.5 104337.5 ;
      RECT  8207.5 104337.5 8272.5 104472.5 ;
      RECT  8397.5 104337.5 8462.5 104472.5 ;
      RECT  8397.5 104337.5 8462.5 104472.5 ;
      RECT  8207.5 104337.5 8272.5 104472.5 ;
      RECT  8207.5 103452.5 8272.5 103587.5 ;
      RECT  8397.5 103452.5 8462.5 103587.5 ;
      RECT  8397.5 103452.5 8462.5 103587.5 ;
      RECT  8207.5 103452.5 8272.5 103587.5 ;
      RECT  8567.5 104427.5 8632.5 104562.5 ;
      RECT  8567.5 103452.5 8632.5 103587.5 ;
      RECT  8265.0 103895.0 8330.0 104030.0 ;
      RECT  8265.0 103895.0 8330.0 104030.0 ;
      RECT  8430.0 103930.0 8495.0 103995.0 ;
      RECT  8140.0 104647.5 8700.0 104712.5 ;
      RECT  8140.0 103302.5 8700.0 103367.5 ;
      RECT  8567.5 104865.0 8632.5 104680.0 ;
      RECT  8567.5 106025.0 8632.5 105840.0 ;
      RECT  8207.5 105907.5 8272.5 106057.5 ;
      RECT  8207.5 105022.5 8272.5 104647.5 ;
      RECT  8397.5 105907.5 8462.5 105022.5 ;
      RECT  8207.5 105022.5 8272.5 104887.5 ;
      RECT  8397.5 105022.5 8462.5 104887.5 ;
      RECT  8397.5 105022.5 8462.5 104887.5 ;
      RECT  8207.5 105022.5 8272.5 104887.5 ;
      RECT  8207.5 105907.5 8272.5 105772.5 ;
      RECT  8397.5 105907.5 8462.5 105772.5 ;
      RECT  8397.5 105907.5 8462.5 105772.5 ;
      RECT  8207.5 105907.5 8272.5 105772.5 ;
      RECT  8567.5 104932.5 8632.5 104797.5 ;
      RECT  8567.5 105907.5 8632.5 105772.5 ;
      RECT  8265.0 105465.0 8330.0 105330.0 ;
      RECT  8265.0 105465.0 8330.0 105330.0 ;
      RECT  8430.0 105430.0 8495.0 105365.0 ;
      RECT  8140.0 104712.5 8700.0 104647.5 ;
      RECT  8140.0 106057.5 8700.0 105992.5 ;
      RECT  8567.5 107185.0 8632.5 107370.0 ;
      RECT  8567.5 106025.0 8632.5 106210.0 ;
      RECT  8207.5 106142.5 8272.5 105992.5 ;
      RECT  8207.5 107027.5 8272.5 107402.5 ;
      RECT  8397.5 106142.5 8462.5 107027.5 ;
      RECT  8207.5 107027.5 8272.5 107162.5 ;
      RECT  8397.5 107027.5 8462.5 107162.5 ;
      RECT  8397.5 107027.5 8462.5 107162.5 ;
      RECT  8207.5 107027.5 8272.5 107162.5 ;
      RECT  8207.5 106142.5 8272.5 106277.5 ;
      RECT  8397.5 106142.5 8462.5 106277.5 ;
      RECT  8397.5 106142.5 8462.5 106277.5 ;
      RECT  8207.5 106142.5 8272.5 106277.5 ;
      RECT  8567.5 107117.5 8632.5 107252.5 ;
      RECT  8567.5 106142.5 8632.5 106277.5 ;
      RECT  8265.0 106585.0 8330.0 106720.0 ;
      RECT  8265.0 106585.0 8330.0 106720.0 ;
      RECT  8430.0 106620.0 8495.0 106685.0 ;
      RECT  8140.0 107337.5 8700.0 107402.5 ;
      RECT  8140.0 105992.5 8700.0 106057.5 ;
      RECT  8567.5 107555.0 8632.5 107370.0 ;
      RECT  8567.5 108715.0 8632.5 108530.0 ;
      RECT  8207.5 108597.5 8272.5 108747.5 ;
      RECT  8207.5 107712.5 8272.5 107337.5 ;
      RECT  8397.5 108597.5 8462.5 107712.5 ;
      RECT  8207.5 107712.5 8272.5 107577.5 ;
      RECT  8397.5 107712.5 8462.5 107577.5 ;
      RECT  8397.5 107712.5 8462.5 107577.5 ;
      RECT  8207.5 107712.5 8272.5 107577.5 ;
      RECT  8207.5 108597.5 8272.5 108462.5 ;
      RECT  8397.5 108597.5 8462.5 108462.5 ;
      RECT  8397.5 108597.5 8462.5 108462.5 ;
      RECT  8207.5 108597.5 8272.5 108462.5 ;
      RECT  8567.5 107622.5 8632.5 107487.5 ;
      RECT  8567.5 108597.5 8632.5 108462.5 ;
      RECT  8265.0 108155.0 8330.0 108020.0 ;
      RECT  8265.0 108155.0 8330.0 108020.0 ;
      RECT  8430.0 108120.0 8495.0 108055.0 ;
      RECT  8140.0 107402.5 8700.0 107337.5 ;
      RECT  8140.0 108747.5 8700.0 108682.5 ;
      RECT  8567.5 109875.0 8632.5 110060.0 ;
      RECT  8567.5 108715.0 8632.5 108900.0 ;
      RECT  8207.5 108832.5 8272.5 108682.5 ;
      RECT  8207.5 109717.5 8272.5 110092.5 ;
      RECT  8397.5 108832.5 8462.5 109717.5 ;
      RECT  8207.5 109717.5 8272.5 109852.5 ;
      RECT  8397.5 109717.5 8462.5 109852.5 ;
      RECT  8397.5 109717.5 8462.5 109852.5 ;
      RECT  8207.5 109717.5 8272.5 109852.5 ;
      RECT  8207.5 108832.5 8272.5 108967.5 ;
      RECT  8397.5 108832.5 8462.5 108967.5 ;
      RECT  8397.5 108832.5 8462.5 108967.5 ;
      RECT  8207.5 108832.5 8272.5 108967.5 ;
      RECT  8567.5 109807.5 8632.5 109942.5 ;
      RECT  8567.5 108832.5 8632.5 108967.5 ;
      RECT  8265.0 109275.0 8330.0 109410.0 ;
      RECT  8265.0 109275.0 8330.0 109410.0 ;
      RECT  8430.0 109310.0 8495.0 109375.0 ;
      RECT  8140.0 110027.5 8700.0 110092.5 ;
      RECT  8140.0 108682.5 8700.0 108747.5 ;
      RECT  8567.5 110245.0 8632.5 110060.0 ;
      RECT  8567.5 111405.0 8632.5 111220.0 ;
      RECT  8207.5 111287.5 8272.5 111437.5 ;
      RECT  8207.5 110402.5 8272.5 110027.5 ;
      RECT  8397.5 111287.5 8462.5 110402.5 ;
      RECT  8207.5 110402.5 8272.5 110267.5 ;
      RECT  8397.5 110402.5 8462.5 110267.5 ;
      RECT  8397.5 110402.5 8462.5 110267.5 ;
      RECT  8207.5 110402.5 8272.5 110267.5 ;
      RECT  8207.5 111287.5 8272.5 111152.5 ;
      RECT  8397.5 111287.5 8462.5 111152.5 ;
      RECT  8397.5 111287.5 8462.5 111152.5 ;
      RECT  8207.5 111287.5 8272.5 111152.5 ;
      RECT  8567.5 110312.5 8632.5 110177.5 ;
      RECT  8567.5 111287.5 8632.5 111152.5 ;
      RECT  8265.0 110845.0 8330.0 110710.0 ;
      RECT  8265.0 110845.0 8330.0 110710.0 ;
      RECT  8430.0 110810.0 8495.0 110745.0 ;
      RECT  8140.0 110092.5 8700.0 110027.5 ;
      RECT  8140.0 111437.5 8700.0 111372.5 ;
      RECT  8567.5 112565.0 8632.5 112750.0 ;
      RECT  8567.5 111405.0 8632.5 111590.0 ;
      RECT  8207.5 111522.5 8272.5 111372.5 ;
      RECT  8207.5 112407.5 8272.5 112782.5 ;
      RECT  8397.5 111522.5 8462.5 112407.5 ;
      RECT  8207.5 112407.5 8272.5 112542.5 ;
      RECT  8397.5 112407.5 8462.5 112542.5 ;
      RECT  8397.5 112407.5 8462.5 112542.5 ;
      RECT  8207.5 112407.5 8272.5 112542.5 ;
      RECT  8207.5 111522.5 8272.5 111657.5 ;
      RECT  8397.5 111522.5 8462.5 111657.5 ;
      RECT  8397.5 111522.5 8462.5 111657.5 ;
      RECT  8207.5 111522.5 8272.5 111657.5 ;
      RECT  8567.5 112497.5 8632.5 112632.5 ;
      RECT  8567.5 111522.5 8632.5 111657.5 ;
      RECT  8265.0 111965.0 8330.0 112100.0 ;
      RECT  8265.0 111965.0 8330.0 112100.0 ;
      RECT  8430.0 112000.0 8495.0 112065.0 ;
      RECT  8140.0 112717.5 8700.0 112782.5 ;
      RECT  8140.0 111372.5 8700.0 111437.5 ;
      RECT  8567.5 112935.0 8632.5 112750.0 ;
      RECT  8567.5 114095.0 8632.5 113910.0 ;
      RECT  8207.5 113977.5 8272.5 114127.5 ;
      RECT  8207.5 113092.5 8272.5 112717.5 ;
      RECT  8397.5 113977.5 8462.5 113092.5 ;
      RECT  8207.5 113092.5 8272.5 112957.5 ;
      RECT  8397.5 113092.5 8462.5 112957.5 ;
      RECT  8397.5 113092.5 8462.5 112957.5 ;
      RECT  8207.5 113092.5 8272.5 112957.5 ;
      RECT  8207.5 113977.5 8272.5 113842.5 ;
      RECT  8397.5 113977.5 8462.5 113842.5 ;
      RECT  8397.5 113977.5 8462.5 113842.5 ;
      RECT  8207.5 113977.5 8272.5 113842.5 ;
      RECT  8567.5 113002.5 8632.5 112867.5 ;
      RECT  8567.5 113977.5 8632.5 113842.5 ;
      RECT  8265.0 113535.0 8330.0 113400.0 ;
      RECT  8265.0 113535.0 8330.0 113400.0 ;
      RECT  8430.0 113500.0 8495.0 113435.0 ;
      RECT  8140.0 112782.5 8700.0 112717.5 ;
      RECT  8140.0 114127.5 8700.0 114062.5 ;
      RECT  5132.5 12470.0 4997.5 12535.0 ;
      RECT  5307.5 13905.0 5172.5 13970.0 ;
      RECT  5482.5 15160.0 5347.5 15225.0 ;
      RECT  5657.5 16595.0 5522.5 16660.0 ;
      RECT  5832.5 17850.0 5697.5 17915.0 ;
      RECT  6007.5 19285.0 5872.5 19350.0 ;
      RECT  6182.5 20540.0 6047.5 20605.0 ;
      RECT  6357.5 21975.0 6222.5 22040.0 ;
      RECT  6532.5 23230.0 6397.5 23295.0 ;
      RECT  6707.5 24665.0 6572.5 24730.0 ;
      RECT  6882.5 25920.0 6747.5 25985.0 ;
      RECT  7057.5 27355.0 6922.5 27420.0 ;
      RECT  5132.5 28670.0 4997.5 28735.0 ;
      RECT  5832.5 28530.0 5697.5 28595.0 ;
      RECT  6532.5 28390.0 6397.5 28455.0 ;
      RECT  5132.5 29985.0 4997.5 30050.0 ;
      RECT  5832.5 30125.0 5697.5 30190.0 ;
      RECT  6707.5 30265.0 6572.5 30330.0 ;
      RECT  5132.5 31360.0 4997.5 31425.0 ;
      RECT  5832.5 31220.0 5697.5 31285.0 ;
      RECT  6882.5 31080.0 6747.5 31145.0 ;
      RECT  5132.5 32675.0 4997.5 32740.0 ;
      RECT  5832.5 32815.0 5697.5 32880.0 ;
      RECT  7057.5 32955.0 6922.5 33020.0 ;
      RECT  5132.5 34050.0 4997.5 34115.0 ;
      RECT  6007.5 33910.0 5872.5 33975.0 ;
      RECT  6532.5 33770.0 6397.5 33835.0 ;
      RECT  5132.5 35365.0 4997.5 35430.0 ;
      RECT  6007.5 35505.0 5872.5 35570.0 ;
      RECT  6707.5 35645.0 6572.5 35710.0 ;
      RECT  5132.5 36740.0 4997.5 36805.0 ;
      RECT  6007.5 36600.0 5872.5 36665.0 ;
      RECT  6882.5 36460.0 6747.5 36525.0 ;
      RECT  5132.5 38055.0 4997.5 38120.0 ;
      RECT  6007.5 38195.0 5872.5 38260.0 ;
      RECT  7057.5 38335.0 6922.5 38400.0 ;
      RECT  5132.5 39430.0 4997.5 39495.0 ;
      RECT  6182.5 39290.0 6047.5 39355.0 ;
      RECT  6532.5 39150.0 6397.5 39215.0 ;
      RECT  5132.5 40745.0 4997.5 40810.0 ;
      RECT  6182.5 40885.0 6047.5 40950.0 ;
      RECT  6707.5 41025.0 6572.5 41090.0 ;
      RECT  5132.5 42120.0 4997.5 42185.0 ;
      RECT  6182.5 41980.0 6047.5 42045.0 ;
      RECT  6882.5 41840.0 6747.5 41905.0 ;
      RECT  5132.5 43435.0 4997.5 43500.0 ;
      RECT  6182.5 43575.0 6047.5 43640.0 ;
      RECT  7057.5 43715.0 6922.5 43780.0 ;
      RECT  5132.5 44810.0 4997.5 44875.0 ;
      RECT  6357.5 44670.0 6222.5 44735.0 ;
      RECT  6532.5 44530.0 6397.5 44595.0 ;
      RECT  5132.5 46125.0 4997.5 46190.0 ;
      RECT  6357.5 46265.0 6222.5 46330.0 ;
      RECT  6707.5 46405.0 6572.5 46470.0 ;
      RECT  5132.5 47500.0 4997.5 47565.0 ;
      RECT  6357.5 47360.0 6222.5 47425.0 ;
      RECT  6882.5 47220.0 6747.5 47285.0 ;
      RECT  5132.5 48815.0 4997.5 48880.0 ;
      RECT  6357.5 48955.0 6222.5 49020.0 ;
      RECT  7057.5 49095.0 6922.5 49160.0 ;
      RECT  5307.5 50190.0 5172.5 50255.0 ;
      RECT  5832.5 50050.0 5697.5 50115.0 ;
      RECT  6532.5 49910.0 6397.5 49975.0 ;
      RECT  5307.5 51505.0 5172.5 51570.0 ;
      RECT  5832.5 51645.0 5697.5 51710.0 ;
      RECT  6707.5 51785.0 6572.5 51850.0 ;
      RECT  5307.5 52880.0 5172.5 52945.0 ;
      RECT  5832.5 52740.0 5697.5 52805.0 ;
      RECT  6882.5 52600.0 6747.5 52665.0 ;
      RECT  5307.5 54195.0 5172.5 54260.0 ;
      RECT  5832.5 54335.0 5697.5 54400.0 ;
      RECT  7057.5 54475.0 6922.5 54540.0 ;
      RECT  5307.5 55570.0 5172.5 55635.0 ;
      RECT  6007.5 55430.0 5872.5 55495.0 ;
      RECT  6532.5 55290.0 6397.5 55355.0 ;
      RECT  5307.5 56885.0 5172.5 56950.0 ;
      RECT  6007.5 57025.0 5872.5 57090.0 ;
      RECT  6707.5 57165.0 6572.5 57230.0 ;
      RECT  5307.5 58260.0 5172.5 58325.0 ;
      RECT  6007.5 58120.0 5872.5 58185.0 ;
      RECT  6882.5 57980.0 6747.5 58045.0 ;
      RECT  5307.5 59575.0 5172.5 59640.0 ;
      RECT  6007.5 59715.0 5872.5 59780.0 ;
      RECT  7057.5 59855.0 6922.5 59920.0 ;
      RECT  5307.5 60950.0 5172.5 61015.0 ;
      RECT  6182.5 60810.0 6047.5 60875.0 ;
      RECT  6532.5 60670.0 6397.5 60735.0 ;
      RECT  5307.5 62265.0 5172.5 62330.0 ;
      RECT  6182.5 62405.0 6047.5 62470.0 ;
      RECT  6707.5 62545.0 6572.5 62610.0 ;
      RECT  5307.5 63640.0 5172.5 63705.0 ;
      RECT  6182.5 63500.0 6047.5 63565.0 ;
      RECT  6882.5 63360.0 6747.5 63425.0 ;
      RECT  5307.5 64955.0 5172.5 65020.0 ;
      RECT  6182.5 65095.0 6047.5 65160.0 ;
      RECT  7057.5 65235.0 6922.5 65300.0 ;
      RECT  5307.5 66330.0 5172.5 66395.0 ;
      RECT  6357.5 66190.0 6222.5 66255.0 ;
      RECT  6532.5 66050.0 6397.5 66115.0 ;
      RECT  5307.5 67645.0 5172.5 67710.0 ;
      RECT  6357.5 67785.0 6222.5 67850.0 ;
      RECT  6707.5 67925.0 6572.5 67990.0 ;
      RECT  5307.5 69020.0 5172.5 69085.0 ;
      RECT  6357.5 68880.0 6222.5 68945.0 ;
      RECT  6882.5 68740.0 6747.5 68805.0 ;
      RECT  5307.5 70335.0 5172.5 70400.0 ;
      RECT  6357.5 70475.0 6222.5 70540.0 ;
      RECT  7057.5 70615.0 6922.5 70680.0 ;
      RECT  5482.5 71710.0 5347.5 71775.0 ;
      RECT  5832.5 71570.0 5697.5 71635.0 ;
      RECT  6532.5 71430.0 6397.5 71495.0 ;
      RECT  5482.5 73025.0 5347.5 73090.0 ;
      RECT  5832.5 73165.0 5697.5 73230.0 ;
      RECT  6707.5 73305.0 6572.5 73370.0 ;
      RECT  5482.5 74400.0 5347.5 74465.0 ;
      RECT  5832.5 74260.0 5697.5 74325.0 ;
      RECT  6882.5 74120.0 6747.5 74185.0 ;
      RECT  5482.5 75715.0 5347.5 75780.0 ;
      RECT  5832.5 75855.0 5697.5 75920.0 ;
      RECT  7057.5 75995.0 6922.5 76060.0 ;
      RECT  5482.5 77090.0 5347.5 77155.0 ;
      RECT  6007.5 76950.0 5872.5 77015.0 ;
      RECT  6532.5 76810.0 6397.5 76875.0 ;
      RECT  5482.5 78405.0 5347.5 78470.0 ;
      RECT  6007.5 78545.0 5872.5 78610.0 ;
      RECT  6707.5 78685.0 6572.5 78750.0 ;
      RECT  5482.5 79780.0 5347.5 79845.0 ;
      RECT  6007.5 79640.0 5872.5 79705.0 ;
      RECT  6882.5 79500.0 6747.5 79565.0 ;
      RECT  5482.5 81095.0 5347.5 81160.0 ;
      RECT  6007.5 81235.0 5872.5 81300.0 ;
      RECT  7057.5 81375.0 6922.5 81440.0 ;
      RECT  5482.5 82470.0 5347.5 82535.0 ;
      RECT  6182.5 82330.0 6047.5 82395.0 ;
      RECT  6532.5 82190.0 6397.5 82255.0 ;
      RECT  5482.5 83785.0 5347.5 83850.0 ;
      RECT  6182.5 83925.0 6047.5 83990.0 ;
      RECT  6707.5 84065.0 6572.5 84130.0 ;
      RECT  5482.5 85160.0 5347.5 85225.0 ;
      RECT  6182.5 85020.0 6047.5 85085.0 ;
      RECT  6882.5 84880.0 6747.5 84945.0 ;
      RECT  5482.5 86475.0 5347.5 86540.0 ;
      RECT  6182.5 86615.0 6047.5 86680.0 ;
      RECT  7057.5 86755.0 6922.5 86820.0 ;
      RECT  5482.5 87850.0 5347.5 87915.0 ;
      RECT  6357.5 87710.0 6222.5 87775.0 ;
      RECT  6532.5 87570.0 6397.5 87635.0 ;
      RECT  5482.5 89165.0 5347.5 89230.0 ;
      RECT  6357.5 89305.0 6222.5 89370.0 ;
      RECT  6707.5 89445.0 6572.5 89510.0 ;
      RECT  5482.5 90540.0 5347.5 90605.0 ;
      RECT  6357.5 90400.0 6222.5 90465.0 ;
      RECT  6882.5 90260.0 6747.5 90325.0 ;
      RECT  5482.5 91855.0 5347.5 91920.0 ;
      RECT  6357.5 91995.0 6222.5 92060.0 ;
      RECT  7057.5 92135.0 6922.5 92200.0 ;
      RECT  5657.5 93230.0 5522.5 93295.0 ;
      RECT  5832.5 93090.0 5697.5 93155.0 ;
      RECT  6532.5 92950.0 6397.5 93015.0 ;
      RECT  5657.5 94545.0 5522.5 94610.0 ;
      RECT  5832.5 94685.0 5697.5 94750.0 ;
      RECT  6707.5 94825.0 6572.5 94890.0 ;
      RECT  5657.5 95920.0 5522.5 95985.0 ;
      RECT  5832.5 95780.0 5697.5 95845.0 ;
      RECT  6882.5 95640.0 6747.5 95705.0 ;
      RECT  5657.5 97235.0 5522.5 97300.0 ;
      RECT  5832.5 97375.0 5697.5 97440.0 ;
      RECT  7057.5 97515.0 6922.5 97580.0 ;
      RECT  5657.5 98610.0 5522.5 98675.0 ;
      RECT  6007.5 98470.0 5872.5 98535.0 ;
      RECT  6532.5 98330.0 6397.5 98395.0 ;
      RECT  5657.5 99925.0 5522.5 99990.0 ;
      RECT  6007.5 100065.0 5872.5 100130.0 ;
      RECT  6707.5 100205.0 6572.5 100270.0 ;
      RECT  5657.5 101300.0 5522.5 101365.0 ;
      RECT  6007.5 101160.0 5872.5 101225.0 ;
      RECT  6882.5 101020.0 6747.5 101085.0 ;
      RECT  5657.5 102615.0 5522.5 102680.0 ;
      RECT  6007.5 102755.0 5872.5 102820.0 ;
      RECT  7057.5 102895.0 6922.5 102960.0 ;
      RECT  5657.5 103990.0 5522.5 104055.0 ;
      RECT  6182.5 103850.0 6047.5 103915.0 ;
      RECT  6532.5 103710.0 6397.5 103775.0 ;
      RECT  5657.5 105305.0 5522.5 105370.0 ;
      RECT  6182.5 105445.0 6047.5 105510.0 ;
      RECT  6707.5 105585.0 6572.5 105650.0 ;
      RECT  5657.5 106680.0 5522.5 106745.0 ;
      RECT  6182.5 106540.0 6047.5 106605.0 ;
      RECT  6882.5 106400.0 6747.5 106465.0 ;
      RECT  5657.5 107995.0 5522.5 108060.0 ;
      RECT  6182.5 108135.0 6047.5 108200.0 ;
      RECT  7057.5 108275.0 6922.5 108340.0 ;
      RECT  5657.5 109370.0 5522.5 109435.0 ;
      RECT  6357.5 109230.0 6222.5 109295.0 ;
      RECT  6532.5 109090.0 6397.5 109155.0 ;
      RECT  5657.5 110685.0 5522.5 110750.0 ;
      RECT  6357.5 110825.0 6222.5 110890.0 ;
      RECT  6707.5 110965.0 6572.5 111030.0 ;
      RECT  5657.5 112060.0 5522.5 112125.0 ;
      RECT  6357.5 111920.0 6222.5 111985.0 ;
      RECT  6882.5 111780.0 6747.5 111845.0 ;
      RECT  5657.5 113375.0 5522.5 113440.0 ;
      RECT  6357.5 113515.0 6222.5 113580.0 ;
      RECT  7057.5 113655.0 6922.5 113720.0 ;
      RECT  8430.0 28610.0 8495.0 28675.0 ;
      RECT  8430.0 30045.0 8495.0 30110.0 ;
      RECT  8430.0 31300.0 8495.0 31365.0 ;
      RECT  8430.0 32735.0 8495.0 32800.0 ;
      RECT  8430.0 33990.0 8495.0 34055.0 ;
      RECT  8430.0 35425.0 8495.0 35490.0 ;
      RECT  8430.0 36680.0 8495.0 36745.0 ;
      RECT  8430.0 38115.0 8495.0 38180.0 ;
      RECT  8430.0 39370.0 8495.0 39435.0 ;
      RECT  8430.0 40805.0 8495.0 40870.0 ;
      RECT  8430.0 42060.0 8495.0 42125.0 ;
      RECT  8430.0 43495.0 8495.0 43560.0 ;
      RECT  8430.0 44750.0 8495.0 44815.0 ;
      RECT  8430.0 46185.0 8495.0 46250.0 ;
      RECT  8430.0 47440.0 8495.0 47505.0 ;
      RECT  8430.0 48875.0 8495.0 48940.0 ;
      RECT  8430.0 50130.0 8495.0 50195.0 ;
      RECT  8430.0 51565.0 8495.0 51630.0 ;
      RECT  8430.0 52820.0 8495.0 52885.0 ;
      RECT  8430.0 54255.0 8495.0 54320.0 ;
      RECT  8430.0 55510.0 8495.0 55575.0 ;
      RECT  8430.0 56945.0 8495.0 57010.0 ;
      RECT  8430.0 58200.0 8495.0 58265.0 ;
      RECT  8430.0 59635.0 8495.0 59700.0 ;
      RECT  8430.0 60890.0 8495.0 60955.0 ;
      RECT  8430.0 62325.0 8495.0 62390.0 ;
      RECT  8430.0 63580.0 8495.0 63645.0 ;
      RECT  8430.0 65015.0 8495.0 65080.0 ;
      RECT  8430.0 66270.0 8495.0 66335.0 ;
      RECT  8430.0 67705.0 8495.0 67770.0 ;
      RECT  8430.0 68960.0 8495.0 69025.0 ;
      RECT  8430.0 70395.0 8495.0 70460.0 ;
      RECT  8430.0 71650.0 8495.0 71715.0 ;
      RECT  8430.0 73085.0 8495.0 73150.0 ;
      RECT  8430.0 74340.0 8495.0 74405.0 ;
      RECT  8430.0 75775.0 8495.0 75840.0 ;
      RECT  8430.0 77030.0 8495.0 77095.0 ;
      RECT  8430.0 78465.0 8495.0 78530.0 ;
      RECT  8430.0 79720.0 8495.0 79785.0 ;
      RECT  8430.0 81155.0 8495.0 81220.0 ;
      RECT  8430.0 82410.0 8495.0 82475.0 ;
      RECT  8430.0 83845.0 8495.0 83910.0 ;
      RECT  8430.0 85100.0 8495.0 85165.0 ;
      RECT  8430.0 86535.0 8495.0 86600.0 ;
      RECT  8430.0 87790.0 8495.0 87855.0 ;
      RECT  8430.0 89225.0 8495.0 89290.0 ;
      RECT  8430.0 90480.0 8495.0 90545.0 ;
      RECT  8430.0 91915.0 8495.0 91980.0 ;
      RECT  8430.0 93170.0 8495.0 93235.0 ;
      RECT  8430.0 94605.0 8495.0 94670.0 ;
      RECT  8430.0 95860.0 8495.0 95925.0 ;
      RECT  8430.0 97295.0 8495.0 97360.0 ;
      RECT  8430.0 98550.0 8495.0 98615.0 ;
      RECT  8430.0 99985.0 8495.0 100050.0 ;
      RECT  8430.0 101240.0 8495.0 101305.0 ;
      RECT  8430.0 102675.0 8495.0 102740.0 ;
      RECT  8430.0 103930.0 8495.0 103995.0 ;
      RECT  8430.0 105365.0 8495.0 105430.0 ;
      RECT  8430.0 106620.0 8495.0 106685.0 ;
      RECT  8430.0 108055.0 8495.0 108120.0 ;
      RECT  8430.0 109310.0 8495.0 109375.0 ;
      RECT  8430.0 110745.0 8495.0 110810.0 ;
      RECT  8430.0 112000.0 8495.0 112065.0 ;
      RECT  8430.0 113435.0 8495.0 113500.0 ;
      RECT  5030.0 13187.5 11095.0 13252.5 ;
      RECT  5030.0 15877.5 11095.0 15942.5 ;
      RECT  5030.0 18567.5 11095.0 18632.5 ;
      RECT  5030.0 21257.5 11095.0 21322.5 ;
      RECT  5030.0 23947.5 11095.0 24012.5 ;
      RECT  5030.0 26637.5 11095.0 26702.5 ;
      RECT  5030.0 29327.5 11095.0 29392.5 ;
      RECT  5030.0 32017.5 11095.0 32082.5 ;
      RECT  5030.0 34707.5 11095.0 34772.5 ;
      RECT  5030.0 37397.5 11095.0 37462.5 ;
      RECT  5030.0 40087.5 11095.0 40152.5 ;
      RECT  5030.0 42777.5 11095.0 42842.5 ;
      RECT  5030.0 45467.5 11095.0 45532.5 ;
      RECT  5030.0 48157.5 11095.0 48222.5 ;
      RECT  5030.0 50847.5 11095.0 50912.5 ;
      RECT  5030.0 53537.5 11095.0 53602.5 ;
      RECT  5030.0 56227.5 11095.0 56292.5 ;
      RECT  5030.0 58917.5 11095.0 58982.5 ;
      RECT  5030.0 61607.5 11095.0 61672.5 ;
      RECT  5030.0 64297.5 11095.0 64362.5 ;
      RECT  5030.0 66987.5 11095.0 67052.5 ;
      RECT  5030.0 69677.5 11095.0 69742.5 ;
      RECT  5030.0 72367.5 11095.0 72432.5 ;
      RECT  5030.0 75057.5 11095.0 75122.5 ;
      RECT  5030.0 77747.5 11095.0 77812.5 ;
      RECT  5030.0 80437.5 11095.0 80502.5 ;
      RECT  5030.0 83127.5 11095.0 83192.5 ;
      RECT  5030.0 85817.5 11095.0 85882.5 ;
      RECT  5030.0 88507.5 11095.0 88572.5 ;
      RECT  5030.0 91197.5 11095.0 91262.5 ;
      RECT  5030.0 93887.5 11095.0 93952.5 ;
      RECT  5030.0 96577.5 11095.0 96642.5 ;
      RECT  5030.0 99267.5 11095.0 99332.5 ;
      RECT  5030.0 101957.5 11095.0 102022.5 ;
      RECT  5030.0 104647.5 11095.0 104712.5 ;
      RECT  5030.0 107337.5 11095.0 107402.5 ;
      RECT  5030.0 110027.5 11095.0 110092.5 ;
      RECT  5030.0 112717.5 11095.0 112782.5 ;
      RECT  5030.0 11842.5 11095.0 11907.5 ;
      RECT  5030.0 14532.5 11095.0 14597.5 ;
      RECT  5030.0 17222.5 11095.0 17287.5 ;
      RECT  5030.0 19912.5 11095.0 19977.5 ;
      RECT  5030.0 22602.5 11095.0 22667.5 ;
      RECT  5030.0 25292.5 11095.0 25357.5 ;
      RECT  5030.0 27982.5 11095.0 28047.5 ;
      RECT  5030.0 30672.5 11095.0 30737.5 ;
      RECT  5030.0 33362.5 11095.0 33427.5 ;
      RECT  5030.0 36052.5 11095.0 36117.5 ;
      RECT  5030.0 38742.5 11095.0 38807.5 ;
      RECT  5030.0 41432.5 11095.0 41497.5 ;
      RECT  5030.0 44122.5 11095.0 44187.5 ;
      RECT  5030.0 46812.5 11095.0 46877.5 ;
      RECT  5030.0 49502.5 11095.0 49567.5 ;
      RECT  5030.0 52192.5 11095.0 52257.5 ;
      RECT  5030.0 54882.5 11095.0 54947.5 ;
      RECT  5030.0 57572.5 11095.0 57637.5 ;
      RECT  5030.0 60262.5 11095.0 60327.5 ;
      RECT  5030.0 62952.5 11095.0 63017.5 ;
      RECT  5030.0 65642.5 11095.0 65707.5 ;
      RECT  5030.0 68332.5 11095.0 68397.5 ;
      RECT  5030.0 71022.5 11095.0 71087.5 ;
      RECT  5030.0 73712.5 11095.0 73777.5 ;
      RECT  5030.0 76402.5 11095.0 76467.5 ;
      RECT  5030.0 79092.5 11095.0 79157.5 ;
      RECT  5030.0 81782.5 11095.0 81847.5 ;
      RECT  5030.0 84472.5 11095.0 84537.5 ;
      RECT  5030.0 87162.5 11095.0 87227.5 ;
      RECT  5030.0 89852.5 11095.0 89917.5 ;
      RECT  5030.0 92542.5 11095.0 92607.5 ;
      RECT  5030.0 95232.5 11095.0 95297.5 ;
      RECT  5030.0 97922.5 11095.0 97987.5 ;
      RECT  5030.0 100612.5 11095.0 100677.5 ;
      RECT  5030.0 103302.5 11095.0 103367.5 ;
      RECT  5030.0 105992.5 11095.0 106057.5 ;
      RECT  5030.0 108682.5 11095.0 108747.5 ;
      RECT  5030.0 111372.5 11095.0 111437.5 ;
      RECT  5030.0 114062.5 11095.0 114127.5 ;
      RECT  8930.0 28610.0 9280.0 28675.0 ;
      RECT  9445.0 28622.5 9510.0 28687.5 ;
      RECT  9445.0 28610.0 9510.0 28675.0 ;
      RECT  9445.0 28655.0 9510.0 28675.0 ;
      RECT  9477.5 28622.5 9775.0 28687.5 ;
      RECT  9775.0 28622.5 9910.0 28687.5 ;
      RECT  10480.0 28622.5 10545.0 28687.5 ;
      RECT  10480.0 28610.0 10545.0 28675.0 ;
      RECT  10262.5 28622.5 10512.5 28687.5 ;
      RECT  10480.0 28642.5 10545.0 28655.0 ;
      RECT  10512.5 28610.0 10760.0 28675.0 ;
      RECT  8930.0 30045.0 9280.0 30110.0 ;
      RECT  9445.0 30032.5 9510.0 30097.5 ;
      RECT  9445.0 30045.0 9510.0 30110.0 ;
      RECT  9445.0 30065.0 9510.0 30110.0 ;
      RECT  9477.5 30032.5 9775.0 30097.5 ;
      RECT  9775.0 30032.5 9910.0 30097.5 ;
      RECT  10480.0 30032.5 10545.0 30097.5 ;
      RECT  10480.0 30045.0 10545.0 30110.0 ;
      RECT  10262.5 30032.5 10512.5 30097.5 ;
      RECT  10480.0 30065.0 10545.0 30077.5 ;
      RECT  10512.5 30045.0 10760.0 30110.0 ;
      RECT  8930.0 31300.0 9280.0 31365.0 ;
      RECT  9445.0 31312.5 9510.0 31377.5 ;
      RECT  9445.0 31300.0 9510.0 31365.0 ;
      RECT  9445.0 31345.0 9510.0 31365.0 ;
      RECT  9477.5 31312.5 9775.0 31377.5 ;
      RECT  9775.0 31312.5 9910.0 31377.5 ;
      RECT  10480.0 31312.5 10545.0 31377.5 ;
      RECT  10480.0 31300.0 10545.0 31365.0 ;
      RECT  10262.5 31312.5 10512.5 31377.5 ;
      RECT  10480.0 31332.5 10545.0 31345.0 ;
      RECT  10512.5 31300.0 10760.0 31365.0 ;
      RECT  8930.0 32735.0 9280.0 32800.0 ;
      RECT  9445.0 32722.5 9510.0 32787.5 ;
      RECT  9445.0 32735.0 9510.0 32800.0 ;
      RECT  9445.0 32755.0 9510.0 32800.0 ;
      RECT  9477.5 32722.5 9775.0 32787.5 ;
      RECT  9775.0 32722.5 9910.0 32787.5 ;
      RECT  10480.0 32722.5 10545.0 32787.5 ;
      RECT  10480.0 32735.0 10545.0 32800.0 ;
      RECT  10262.5 32722.5 10512.5 32787.5 ;
      RECT  10480.0 32755.0 10545.0 32767.5 ;
      RECT  10512.5 32735.0 10760.0 32800.0 ;
      RECT  8930.0 33990.0 9280.0 34055.0 ;
      RECT  9445.0 34002.5 9510.0 34067.5 ;
      RECT  9445.0 33990.0 9510.0 34055.0 ;
      RECT  9445.0 34035.0 9510.0 34055.0 ;
      RECT  9477.5 34002.5 9775.0 34067.5 ;
      RECT  9775.0 34002.5 9910.0 34067.5 ;
      RECT  10480.0 34002.5 10545.0 34067.5 ;
      RECT  10480.0 33990.0 10545.0 34055.0 ;
      RECT  10262.5 34002.5 10512.5 34067.5 ;
      RECT  10480.0 34022.5 10545.0 34035.0 ;
      RECT  10512.5 33990.0 10760.0 34055.0 ;
      RECT  8930.0 35425.0 9280.0 35490.0 ;
      RECT  9445.0 35412.5 9510.0 35477.5 ;
      RECT  9445.0 35425.0 9510.0 35490.0 ;
      RECT  9445.0 35445.0 9510.0 35490.0 ;
      RECT  9477.5 35412.5 9775.0 35477.5 ;
      RECT  9775.0 35412.5 9910.0 35477.5 ;
      RECT  10480.0 35412.5 10545.0 35477.5 ;
      RECT  10480.0 35425.0 10545.0 35490.0 ;
      RECT  10262.5 35412.5 10512.5 35477.5 ;
      RECT  10480.0 35445.0 10545.0 35457.5 ;
      RECT  10512.5 35425.0 10760.0 35490.0 ;
      RECT  8930.0 36680.0 9280.0 36745.0 ;
      RECT  9445.0 36692.5 9510.0 36757.5 ;
      RECT  9445.0 36680.0 9510.0 36745.0 ;
      RECT  9445.0 36725.0 9510.0 36745.0 ;
      RECT  9477.5 36692.5 9775.0 36757.5 ;
      RECT  9775.0 36692.5 9910.0 36757.5 ;
      RECT  10480.0 36692.5 10545.0 36757.5 ;
      RECT  10480.0 36680.0 10545.0 36745.0 ;
      RECT  10262.5 36692.5 10512.5 36757.5 ;
      RECT  10480.0 36712.5 10545.0 36725.0 ;
      RECT  10512.5 36680.0 10760.0 36745.0 ;
      RECT  8930.0 38115.0 9280.0 38180.0 ;
      RECT  9445.0 38102.5 9510.0 38167.5 ;
      RECT  9445.0 38115.0 9510.0 38180.0 ;
      RECT  9445.0 38135.0 9510.0 38180.0 ;
      RECT  9477.5 38102.5 9775.0 38167.5 ;
      RECT  9775.0 38102.5 9910.0 38167.5 ;
      RECT  10480.0 38102.5 10545.0 38167.5 ;
      RECT  10480.0 38115.0 10545.0 38180.0 ;
      RECT  10262.5 38102.5 10512.5 38167.5 ;
      RECT  10480.0 38135.0 10545.0 38147.5 ;
      RECT  10512.5 38115.0 10760.0 38180.0 ;
      RECT  8930.0 39370.0 9280.0 39435.0 ;
      RECT  9445.0 39382.5 9510.0 39447.5 ;
      RECT  9445.0 39370.0 9510.0 39435.0 ;
      RECT  9445.0 39415.0 9510.0 39435.0 ;
      RECT  9477.5 39382.5 9775.0 39447.5 ;
      RECT  9775.0 39382.5 9910.0 39447.5 ;
      RECT  10480.0 39382.5 10545.0 39447.5 ;
      RECT  10480.0 39370.0 10545.0 39435.0 ;
      RECT  10262.5 39382.5 10512.5 39447.5 ;
      RECT  10480.0 39402.5 10545.0 39415.0 ;
      RECT  10512.5 39370.0 10760.0 39435.0 ;
      RECT  8930.0 40805.0 9280.0 40870.0 ;
      RECT  9445.0 40792.5 9510.0 40857.5 ;
      RECT  9445.0 40805.0 9510.0 40870.0 ;
      RECT  9445.0 40825.0 9510.0 40870.0 ;
      RECT  9477.5 40792.5 9775.0 40857.5 ;
      RECT  9775.0 40792.5 9910.0 40857.5 ;
      RECT  10480.0 40792.5 10545.0 40857.5 ;
      RECT  10480.0 40805.0 10545.0 40870.0 ;
      RECT  10262.5 40792.5 10512.5 40857.5 ;
      RECT  10480.0 40825.0 10545.0 40837.5 ;
      RECT  10512.5 40805.0 10760.0 40870.0 ;
      RECT  8930.0 42060.0 9280.0 42125.0 ;
      RECT  9445.0 42072.5 9510.0 42137.5 ;
      RECT  9445.0 42060.0 9510.0 42125.0 ;
      RECT  9445.0 42105.0 9510.0 42125.0 ;
      RECT  9477.5 42072.5 9775.0 42137.5 ;
      RECT  9775.0 42072.5 9910.0 42137.5 ;
      RECT  10480.0 42072.5 10545.0 42137.5 ;
      RECT  10480.0 42060.0 10545.0 42125.0 ;
      RECT  10262.5 42072.5 10512.5 42137.5 ;
      RECT  10480.0 42092.5 10545.0 42105.0 ;
      RECT  10512.5 42060.0 10760.0 42125.0 ;
      RECT  8930.0 43495.0 9280.0 43560.0 ;
      RECT  9445.0 43482.5 9510.0 43547.5 ;
      RECT  9445.0 43495.0 9510.0 43560.0 ;
      RECT  9445.0 43515.0 9510.0 43560.0 ;
      RECT  9477.5 43482.5 9775.0 43547.5 ;
      RECT  9775.0 43482.5 9910.0 43547.5 ;
      RECT  10480.0 43482.5 10545.0 43547.5 ;
      RECT  10480.0 43495.0 10545.0 43560.0 ;
      RECT  10262.5 43482.5 10512.5 43547.5 ;
      RECT  10480.0 43515.0 10545.0 43527.5 ;
      RECT  10512.5 43495.0 10760.0 43560.0 ;
      RECT  8930.0 44750.0 9280.0 44815.0 ;
      RECT  9445.0 44762.5 9510.0 44827.5 ;
      RECT  9445.0 44750.0 9510.0 44815.0 ;
      RECT  9445.0 44795.0 9510.0 44815.0 ;
      RECT  9477.5 44762.5 9775.0 44827.5 ;
      RECT  9775.0 44762.5 9910.0 44827.5 ;
      RECT  10480.0 44762.5 10545.0 44827.5 ;
      RECT  10480.0 44750.0 10545.0 44815.0 ;
      RECT  10262.5 44762.5 10512.5 44827.5 ;
      RECT  10480.0 44782.5 10545.0 44795.0 ;
      RECT  10512.5 44750.0 10760.0 44815.0 ;
      RECT  8930.0 46185.0 9280.0 46250.0 ;
      RECT  9445.0 46172.5 9510.0 46237.5 ;
      RECT  9445.0 46185.0 9510.0 46250.0 ;
      RECT  9445.0 46205.0 9510.0 46250.0 ;
      RECT  9477.5 46172.5 9775.0 46237.5 ;
      RECT  9775.0 46172.5 9910.0 46237.5 ;
      RECT  10480.0 46172.5 10545.0 46237.5 ;
      RECT  10480.0 46185.0 10545.0 46250.0 ;
      RECT  10262.5 46172.5 10512.5 46237.5 ;
      RECT  10480.0 46205.0 10545.0 46217.5 ;
      RECT  10512.5 46185.0 10760.0 46250.0 ;
      RECT  8930.0 47440.0 9280.0 47505.0 ;
      RECT  9445.0 47452.5 9510.0 47517.5 ;
      RECT  9445.0 47440.0 9510.0 47505.0 ;
      RECT  9445.0 47485.0 9510.0 47505.0 ;
      RECT  9477.5 47452.5 9775.0 47517.5 ;
      RECT  9775.0 47452.5 9910.0 47517.5 ;
      RECT  10480.0 47452.5 10545.0 47517.5 ;
      RECT  10480.0 47440.0 10545.0 47505.0 ;
      RECT  10262.5 47452.5 10512.5 47517.5 ;
      RECT  10480.0 47472.5 10545.0 47485.0 ;
      RECT  10512.5 47440.0 10760.0 47505.0 ;
      RECT  8930.0 48875.0 9280.0 48940.0 ;
      RECT  9445.0 48862.5 9510.0 48927.5 ;
      RECT  9445.0 48875.0 9510.0 48940.0 ;
      RECT  9445.0 48895.0 9510.0 48940.0 ;
      RECT  9477.5 48862.5 9775.0 48927.5 ;
      RECT  9775.0 48862.5 9910.0 48927.5 ;
      RECT  10480.0 48862.5 10545.0 48927.5 ;
      RECT  10480.0 48875.0 10545.0 48940.0 ;
      RECT  10262.5 48862.5 10512.5 48927.5 ;
      RECT  10480.0 48895.0 10545.0 48907.5 ;
      RECT  10512.5 48875.0 10760.0 48940.0 ;
      RECT  8930.0 50130.0 9280.0 50195.0 ;
      RECT  9445.0 50142.5 9510.0 50207.5 ;
      RECT  9445.0 50130.0 9510.0 50195.0 ;
      RECT  9445.0 50175.0 9510.0 50195.0 ;
      RECT  9477.5 50142.5 9775.0 50207.5 ;
      RECT  9775.0 50142.5 9910.0 50207.5 ;
      RECT  10480.0 50142.5 10545.0 50207.5 ;
      RECT  10480.0 50130.0 10545.0 50195.0 ;
      RECT  10262.5 50142.5 10512.5 50207.5 ;
      RECT  10480.0 50162.5 10545.0 50175.0 ;
      RECT  10512.5 50130.0 10760.0 50195.0 ;
      RECT  8930.0 51565.0 9280.0 51630.0 ;
      RECT  9445.0 51552.5 9510.0 51617.5 ;
      RECT  9445.0 51565.0 9510.0 51630.0 ;
      RECT  9445.0 51585.0 9510.0 51630.0 ;
      RECT  9477.5 51552.5 9775.0 51617.5 ;
      RECT  9775.0 51552.5 9910.0 51617.5 ;
      RECT  10480.0 51552.5 10545.0 51617.5 ;
      RECT  10480.0 51565.0 10545.0 51630.0 ;
      RECT  10262.5 51552.5 10512.5 51617.5 ;
      RECT  10480.0 51585.0 10545.0 51597.5 ;
      RECT  10512.5 51565.0 10760.0 51630.0 ;
      RECT  8930.0 52820.0 9280.0 52885.0 ;
      RECT  9445.0 52832.5 9510.0 52897.5 ;
      RECT  9445.0 52820.0 9510.0 52885.0 ;
      RECT  9445.0 52865.0 9510.0 52885.0 ;
      RECT  9477.5 52832.5 9775.0 52897.5 ;
      RECT  9775.0 52832.5 9910.0 52897.5 ;
      RECT  10480.0 52832.5 10545.0 52897.5 ;
      RECT  10480.0 52820.0 10545.0 52885.0 ;
      RECT  10262.5 52832.5 10512.5 52897.5 ;
      RECT  10480.0 52852.5 10545.0 52865.0 ;
      RECT  10512.5 52820.0 10760.0 52885.0 ;
      RECT  8930.0 54255.0 9280.0 54320.0 ;
      RECT  9445.0 54242.5 9510.0 54307.5 ;
      RECT  9445.0 54255.0 9510.0 54320.0 ;
      RECT  9445.0 54275.0 9510.0 54320.0 ;
      RECT  9477.5 54242.5 9775.0 54307.5 ;
      RECT  9775.0 54242.5 9910.0 54307.5 ;
      RECT  10480.0 54242.5 10545.0 54307.5 ;
      RECT  10480.0 54255.0 10545.0 54320.0 ;
      RECT  10262.5 54242.5 10512.5 54307.5 ;
      RECT  10480.0 54275.0 10545.0 54287.5 ;
      RECT  10512.5 54255.0 10760.0 54320.0 ;
      RECT  8930.0 55510.0 9280.0 55575.0 ;
      RECT  9445.0 55522.5 9510.0 55587.5 ;
      RECT  9445.0 55510.0 9510.0 55575.0 ;
      RECT  9445.0 55555.0 9510.0 55575.0 ;
      RECT  9477.5 55522.5 9775.0 55587.5 ;
      RECT  9775.0 55522.5 9910.0 55587.5 ;
      RECT  10480.0 55522.5 10545.0 55587.5 ;
      RECT  10480.0 55510.0 10545.0 55575.0 ;
      RECT  10262.5 55522.5 10512.5 55587.5 ;
      RECT  10480.0 55542.5 10545.0 55555.0 ;
      RECT  10512.5 55510.0 10760.0 55575.0 ;
      RECT  8930.0 56945.0 9280.0 57010.0 ;
      RECT  9445.0 56932.5 9510.0 56997.5 ;
      RECT  9445.0 56945.0 9510.0 57010.0 ;
      RECT  9445.0 56965.0 9510.0 57010.0 ;
      RECT  9477.5 56932.5 9775.0 56997.5 ;
      RECT  9775.0 56932.5 9910.0 56997.5 ;
      RECT  10480.0 56932.5 10545.0 56997.5 ;
      RECT  10480.0 56945.0 10545.0 57010.0 ;
      RECT  10262.5 56932.5 10512.5 56997.5 ;
      RECT  10480.0 56965.0 10545.0 56977.5 ;
      RECT  10512.5 56945.0 10760.0 57010.0 ;
      RECT  8930.0 58200.0 9280.0 58265.0 ;
      RECT  9445.0 58212.5 9510.0 58277.5 ;
      RECT  9445.0 58200.0 9510.0 58265.0 ;
      RECT  9445.0 58245.0 9510.0 58265.0 ;
      RECT  9477.5 58212.5 9775.0 58277.5 ;
      RECT  9775.0 58212.5 9910.0 58277.5 ;
      RECT  10480.0 58212.5 10545.0 58277.5 ;
      RECT  10480.0 58200.0 10545.0 58265.0 ;
      RECT  10262.5 58212.5 10512.5 58277.5 ;
      RECT  10480.0 58232.5 10545.0 58245.0 ;
      RECT  10512.5 58200.0 10760.0 58265.0 ;
      RECT  8930.0 59635.0 9280.0 59700.0 ;
      RECT  9445.0 59622.5 9510.0 59687.5 ;
      RECT  9445.0 59635.0 9510.0 59700.0 ;
      RECT  9445.0 59655.0 9510.0 59700.0 ;
      RECT  9477.5 59622.5 9775.0 59687.5 ;
      RECT  9775.0 59622.5 9910.0 59687.5 ;
      RECT  10480.0 59622.5 10545.0 59687.5 ;
      RECT  10480.0 59635.0 10545.0 59700.0 ;
      RECT  10262.5 59622.5 10512.5 59687.5 ;
      RECT  10480.0 59655.0 10545.0 59667.5 ;
      RECT  10512.5 59635.0 10760.0 59700.0 ;
      RECT  8930.0 60890.0 9280.0 60955.0 ;
      RECT  9445.0 60902.5 9510.0 60967.5 ;
      RECT  9445.0 60890.0 9510.0 60955.0 ;
      RECT  9445.0 60935.0 9510.0 60955.0 ;
      RECT  9477.5 60902.5 9775.0 60967.5 ;
      RECT  9775.0 60902.5 9910.0 60967.5 ;
      RECT  10480.0 60902.5 10545.0 60967.5 ;
      RECT  10480.0 60890.0 10545.0 60955.0 ;
      RECT  10262.5 60902.5 10512.5 60967.5 ;
      RECT  10480.0 60922.5 10545.0 60935.0 ;
      RECT  10512.5 60890.0 10760.0 60955.0 ;
      RECT  8930.0 62325.0 9280.0 62390.0 ;
      RECT  9445.0 62312.5 9510.0 62377.5 ;
      RECT  9445.0 62325.0 9510.0 62390.0 ;
      RECT  9445.0 62345.0 9510.0 62390.0 ;
      RECT  9477.5 62312.5 9775.0 62377.5 ;
      RECT  9775.0 62312.5 9910.0 62377.5 ;
      RECT  10480.0 62312.5 10545.0 62377.5 ;
      RECT  10480.0 62325.0 10545.0 62390.0 ;
      RECT  10262.5 62312.5 10512.5 62377.5 ;
      RECT  10480.0 62345.0 10545.0 62357.5 ;
      RECT  10512.5 62325.0 10760.0 62390.0 ;
      RECT  8930.0 63580.0 9280.0 63645.0 ;
      RECT  9445.0 63592.5 9510.0 63657.5 ;
      RECT  9445.0 63580.0 9510.0 63645.0 ;
      RECT  9445.0 63625.0 9510.0 63645.0 ;
      RECT  9477.5 63592.5 9775.0 63657.5 ;
      RECT  9775.0 63592.5 9910.0 63657.5 ;
      RECT  10480.0 63592.5 10545.0 63657.5 ;
      RECT  10480.0 63580.0 10545.0 63645.0 ;
      RECT  10262.5 63592.5 10512.5 63657.5 ;
      RECT  10480.0 63612.5 10545.0 63625.0 ;
      RECT  10512.5 63580.0 10760.0 63645.0 ;
      RECT  8930.0 65015.0 9280.0 65080.0 ;
      RECT  9445.0 65002.5 9510.0 65067.5 ;
      RECT  9445.0 65015.0 9510.0 65080.0 ;
      RECT  9445.0 65035.0 9510.0 65080.0 ;
      RECT  9477.5 65002.5 9775.0 65067.5 ;
      RECT  9775.0 65002.5 9910.0 65067.5 ;
      RECT  10480.0 65002.5 10545.0 65067.5 ;
      RECT  10480.0 65015.0 10545.0 65080.0 ;
      RECT  10262.5 65002.5 10512.5 65067.5 ;
      RECT  10480.0 65035.0 10545.0 65047.5 ;
      RECT  10512.5 65015.0 10760.0 65080.0 ;
      RECT  8930.0 66270.0 9280.0 66335.0 ;
      RECT  9445.0 66282.5 9510.0 66347.5 ;
      RECT  9445.0 66270.0 9510.0 66335.0 ;
      RECT  9445.0 66315.0 9510.0 66335.0 ;
      RECT  9477.5 66282.5 9775.0 66347.5 ;
      RECT  9775.0 66282.5 9910.0 66347.5 ;
      RECT  10480.0 66282.5 10545.0 66347.5 ;
      RECT  10480.0 66270.0 10545.0 66335.0 ;
      RECT  10262.5 66282.5 10512.5 66347.5 ;
      RECT  10480.0 66302.5 10545.0 66315.0 ;
      RECT  10512.5 66270.0 10760.0 66335.0 ;
      RECT  8930.0 67705.0 9280.0 67770.0 ;
      RECT  9445.0 67692.5 9510.0 67757.5 ;
      RECT  9445.0 67705.0 9510.0 67770.0 ;
      RECT  9445.0 67725.0 9510.0 67770.0 ;
      RECT  9477.5 67692.5 9775.0 67757.5 ;
      RECT  9775.0 67692.5 9910.0 67757.5 ;
      RECT  10480.0 67692.5 10545.0 67757.5 ;
      RECT  10480.0 67705.0 10545.0 67770.0 ;
      RECT  10262.5 67692.5 10512.5 67757.5 ;
      RECT  10480.0 67725.0 10545.0 67737.5 ;
      RECT  10512.5 67705.0 10760.0 67770.0 ;
      RECT  8930.0 68960.0 9280.0 69025.0 ;
      RECT  9445.0 68972.5 9510.0 69037.5 ;
      RECT  9445.0 68960.0 9510.0 69025.0 ;
      RECT  9445.0 69005.0 9510.0 69025.0 ;
      RECT  9477.5 68972.5 9775.0 69037.5 ;
      RECT  9775.0 68972.5 9910.0 69037.5 ;
      RECT  10480.0 68972.5 10545.0 69037.5 ;
      RECT  10480.0 68960.0 10545.0 69025.0 ;
      RECT  10262.5 68972.5 10512.5 69037.5 ;
      RECT  10480.0 68992.5 10545.0 69005.0 ;
      RECT  10512.5 68960.0 10760.0 69025.0 ;
      RECT  8930.0 70395.0 9280.0 70460.0 ;
      RECT  9445.0 70382.5 9510.0 70447.5 ;
      RECT  9445.0 70395.0 9510.0 70460.0 ;
      RECT  9445.0 70415.0 9510.0 70460.0 ;
      RECT  9477.5 70382.5 9775.0 70447.5 ;
      RECT  9775.0 70382.5 9910.0 70447.5 ;
      RECT  10480.0 70382.5 10545.0 70447.5 ;
      RECT  10480.0 70395.0 10545.0 70460.0 ;
      RECT  10262.5 70382.5 10512.5 70447.5 ;
      RECT  10480.0 70415.0 10545.0 70427.5 ;
      RECT  10512.5 70395.0 10760.0 70460.0 ;
      RECT  8930.0 71650.0 9280.0 71715.0 ;
      RECT  9445.0 71662.5 9510.0 71727.5 ;
      RECT  9445.0 71650.0 9510.0 71715.0 ;
      RECT  9445.0 71695.0 9510.0 71715.0 ;
      RECT  9477.5 71662.5 9775.0 71727.5 ;
      RECT  9775.0 71662.5 9910.0 71727.5 ;
      RECT  10480.0 71662.5 10545.0 71727.5 ;
      RECT  10480.0 71650.0 10545.0 71715.0 ;
      RECT  10262.5 71662.5 10512.5 71727.5 ;
      RECT  10480.0 71682.5 10545.0 71695.0 ;
      RECT  10512.5 71650.0 10760.0 71715.0 ;
      RECT  8930.0 73085.0 9280.0 73150.0 ;
      RECT  9445.0 73072.5 9510.0 73137.5 ;
      RECT  9445.0 73085.0 9510.0 73150.0 ;
      RECT  9445.0 73105.0 9510.0 73150.0 ;
      RECT  9477.5 73072.5 9775.0 73137.5 ;
      RECT  9775.0 73072.5 9910.0 73137.5 ;
      RECT  10480.0 73072.5 10545.0 73137.5 ;
      RECT  10480.0 73085.0 10545.0 73150.0 ;
      RECT  10262.5 73072.5 10512.5 73137.5 ;
      RECT  10480.0 73105.0 10545.0 73117.5 ;
      RECT  10512.5 73085.0 10760.0 73150.0 ;
      RECT  8930.0 74340.0 9280.0 74405.0 ;
      RECT  9445.0 74352.5 9510.0 74417.5 ;
      RECT  9445.0 74340.0 9510.0 74405.0 ;
      RECT  9445.0 74385.0 9510.0 74405.0 ;
      RECT  9477.5 74352.5 9775.0 74417.5 ;
      RECT  9775.0 74352.5 9910.0 74417.5 ;
      RECT  10480.0 74352.5 10545.0 74417.5 ;
      RECT  10480.0 74340.0 10545.0 74405.0 ;
      RECT  10262.5 74352.5 10512.5 74417.5 ;
      RECT  10480.0 74372.5 10545.0 74385.0 ;
      RECT  10512.5 74340.0 10760.0 74405.0 ;
      RECT  8930.0 75775.0 9280.0 75840.0 ;
      RECT  9445.0 75762.5 9510.0 75827.5 ;
      RECT  9445.0 75775.0 9510.0 75840.0 ;
      RECT  9445.0 75795.0 9510.0 75840.0 ;
      RECT  9477.5 75762.5 9775.0 75827.5 ;
      RECT  9775.0 75762.5 9910.0 75827.5 ;
      RECT  10480.0 75762.5 10545.0 75827.5 ;
      RECT  10480.0 75775.0 10545.0 75840.0 ;
      RECT  10262.5 75762.5 10512.5 75827.5 ;
      RECT  10480.0 75795.0 10545.0 75807.5 ;
      RECT  10512.5 75775.0 10760.0 75840.0 ;
      RECT  8930.0 77030.0 9280.0 77095.0 ;
      RECT  9445.0 77042.5 9510.0 77107.5 ;
      RECT  9445.0 77030.0 9510.0 77095.0 ;
      RECT  9445.0 77075.0 9510.0 77095.0 ;
      RECT  9477.5 77042.5 9775.0 77107.5 ;
      RECT  9775.0 77042.5 9910.0 77107.5 ;
      RECT  10480.0 77042.5 10545.0 77107.5 ;
      RECT  10480.0 77030.0 10545.0 77095.0 ;
      RECT  10262.5 77042.5 10512.5 77107.5 ;
      RECT  10480.0 77062.5 10545.0 77075.0 ;
      RECT  10512.5 77030.0 10760.0 77095.0 ;
      RECT  8930.0 78465.0 9280.0 78530.0 ;
      RECT  9445.0 78452.5 9510.0 78517.5 ;
      RECT  9445.0 78465.0 9510.0 78530.0 ;
      RECT  9445.0 78485.0 9510.0 78530.0 ;
      RECT  9477.5 78452.5 9775.0 78517.5 ;
      RECT  9775.0 78452.5 9910.0 78517.5 ;
      RECT  10480.0 78452.5 10545.0 78517.5 ;
      RECT  10480.0 78465.0 10545.0 78530.0 ;
      RECT  10262.5 78452.5 10512.5 78517.5 ;
      RECT  10480.0 78485.0 10545.0 78497.5 ;
      RECT  10512.5 78465.0 10760.0 78530.0 ;
      RECT  8930.0 79720.0 9280.0 79785.0 ;
      RECT  9445.0 79732.5 9510.0 79797.5 ;
      RECT  9445.0 79720.0 9510.0 79785.0 ;
      RECT  9445.0 79765.0 9510.0 79785.0 ;
      RECT  9477.5 79732.5 9775.0 79797.5 ;
      RECT  9775.0 79732.5 9910.0 79797.5 ;
      RECT  10480.0 79732.5 10545.0 79797.5 ;
      RECT  10480.0 79720.0 10545.0 79785.0 ;
      RECT  10262.5 79732.5 10512.5 79797.5 ;
      RECT  10480.0 79752.5 10545.0 79765.0 ;
      RECT  10512.5 79720.0 10760.0 79785.0 ;
      RECT  8930.0 81155.0 9280.0 81220.0 ;
      RECT  9445.0 81142.5 9510.0 81207.5 ;
      RECT  9445.0 81155.0 9510.0 81220.0 ;
      RECT  9445.0 81175.0 9510.0 81220.0 ;
      RECT  9477.5 81142.5 9775.0 81207.5 ;
      RECT  9775.0 81142.5 9910.0 81207.5 ;
      RECT  10480.0 81142.5 10545.0 81207.5 ;
      RECT  10480.0 81155.0 10545.0 81220.0 ;
      RECT  10262.5 81142.5 10512.5 81207.5 ;
      RECT  10480.0 81175.0 10545.0 81187.5 ;
      RECT  10512.5 81155.0 10760.0 81220.0 ;
      RECT  8930.0 82410.0 9280.0 82475.0 ;
      RECT  9445.0 82422.5 9510.0 82487.5 ;
      RECT  9445.0 82410.0 9510.0 82475.0 ;
      RECT  9445.0 82455.0 9510.0 82475.0 ;
      RECT  9477.5 82422.5 9775.0 82487.5 ;
      RECT  9775.0 82422.5 9910.0 82487.5 ;
      RECT  10480.0 82422.5 10545.0 82487.5 ;
      RECT  10480.0 82410.0 10545.0 82475.0 ;
      RECT  10262.5 82422.5 10512.5 82487.5 ;
      RECT  10480.0 82442.5 10545.0 82455.0 ;
      RECT  10512.5 82410.0 10760.0 82475.0 ;
      RECT  8930.0 83845.0 9280.0 83910.0 ;
      RECT  9445.0 83832.5 9510.0 83897.5 ;
      RECT  9445.0 83845.0 9510.0 83910.0 ;
      RECT  9445.0 83865.0 9510.0 83910.0 ;
      RECT  9477.5 83832.5 9775.0 83897.5 ;
      RECT  9775.0 83832.5 9910.0 83897.5 ;
      RECT  10480.0 83832.5 10545.0 83897.5 ;
      RECT  10480.0 83845.0 10545.0 83910.0 ;
      RECT  10262.5 83832.5 10512.5 83897.5 ;
      RECT  10480.0 83865.0 10545.0 83877.5 ;
      RECT  10512.5 83845.0 10760.0 83910.0 ;
      RECT  8930.0 85100.0 9280.0 85165.0 ;
      RECT  9445.0 85112.5 9510.0 85177.5 ;
      RECT  9445.0 85100.0 9510.0 85165.0 ;
      RECT  9445.0 85145.0 9510.0 85165.0 ;
      RECT  9477.5 85112.5 9775.0 85177.5 ;
      RECT  9775.0 85112.5 9910.0 85177.5 ;
      RECT  10480.0 85112.5 10545.0 85177.5 ;
      RECT  10480.0 85100.0 10545.0 85165.0 ;
      RECT  10262.5 85112.5 10512.5 85177.5 ;
      RECT  10480.0 85132.5 10545.0 85145.0 ;
      RECT  10512.5 85100.0 10760.0 85165.0 ;
      RECT  8930.0 86535.0 9280.0 86600.0 ;
      RECT  9445.0 86522.5 9510.0 86587.5 ;
      RECT  9445.0 86535.0 9510.0 86600.0 ;
      RECT  9445.0 86555.0 9510.0 86600.0 ;
      RECT  9477.5 86522.5 9775.0 86587.5 ;
      RECT  9775.0 86522.5 9910.0 86587.5 ;
      RECT  10480.0 86522.5 10545.0 86587.5 ;
      RECT  10480.0 86535.0 10545.0 86600.0 ;
      RECT  10262.5 86522.5 10512.5 86587.5 ;
      RECT  10480.0 86555.0 10545.0 86567.5 ;
      RECT  10512.5 86535.0 10760.0 86600.0 ;
      RECT  8930.0 87790.0 9280.0 87855.0 ;
      RECT  9445.0 87802.5 9510.0 87867.5 ;
      RECT  9445.0 87790.0 9510.0 87855.0 ;
      RECT  9445.0 87835.0 9510.0 87855.0 ;
      RECT  9477.5 87802.5 9775.0 87867.5 ;
      RECT  9775.0 87802.5 9910.0 87867.5 ;
      RECT  10480.0 87802.5 10545.0 87867.5 ;
      RECT  10480.0 87790.0 10545.0 87855.0 ;
      RECT  10262.5 87802.5 10512.5 87867.5 ;
      RECT  10480.0 87822.5 10545.0 87835.0 ;
      RECT  10512.5 87790.0 10760.0 87855.0 ;
      RECT  8930.0 89225.0 9280.0 89290.0 ;
      RECT  9445.0 89212.5 9510.0 89277.5 ;
      RECT  9445.0 89225.0 9510.0 89290.0 ;
      RECT  9445.0 89245.0 9510.0 89290.0 ;
      RECT  9477.5 89212.5 9775.0 89277.5 ;
      RECT  9775.0 89212.5 9910.0 89277.5 ;
      RECT  10480.0 89212.5 10545.0 89277.5 ;
      RECT  10480.0 89225.0 10545.0 89290.0 ;
      RECT  10262.5 89212.5 10512.5 89277.5 ;
      RECT  10480.0 89245.0 10545.0 89257.5 ;
      RECT  10512.5 89225.0 10760.0 89290.0 ;
      RECT  8930.0 90480.0 9280.0 90545.0 ;
      RECT  9445.0 90492.5 9510.0 90557.5 ;
      RECT  9445.0 90480.0 9510.0 90545.0 ;
      RECT  9445.0 90525.0 9510.0 90545.0 ;
      RECT  9477.5 90492.5 9775.0 90557.5 ;
      RECT  9775.0 90492.5 9910.0 90557.5 ;
      RECT  10480.0 90492.5 10545.0 90557.5 ;
      RECT  10480.0 90480.0 10545.0 90545.0 ;
      RECT  10262.5 90492.5 10512.5 90557.5 ;
      RECT  10480.0 90512.5 10545.0 90525.0 ;
      RECT  10512.5 90480.0 10760.0 90545.0 ;
      RECT  8930.0 91915.0 9280.0 91980.0 ;
      RECT  9445.0 91902.5 9510.0 91967.5 ;
      RECT  9445.0 91915.0 9510.0 91980.0 ;
      RECT  9445.0 91935.0 9510.0 91980.0 ;
      RECT  9477.5 91902.5 9775.0 91967.5 ;
      RECT  9775.0 91902.5 9910.0 91967.5 ;
      RECT  10480.0 91902.5 10545.0 91967.5 ;
      RECT  10480.0 91915.0 10545.0 91980.0 ;
      RECT  10262.5 91902.5 10512.5 91967.5 ;
      RECT  10480.0 91935.0 10545.0 91947.5 ;
      RECT  10512.5 91915.0 10760.0 91980.0 ;
      RECT  8930.0 93170.0 9280.0 93235.0 ;
      RECT  9445.0 93182.5 9510.0 93247.5 ;
      RECT  9445.0 93170.0 9510.0 93235.0 ;
      RECT  9445.0 93215.0 9510.0 93235.0 ;
      RECT  9477.5 93182.5 9775.0 93247.5 ;
      RECT  9775.0 93182.5 9910.0 93247.5 ;
      RECT  10480.0 93182.5 10545.0 93247.5 ;
      RECT  10480.0 93170.0 10545.0 93235.0 ;
      RECT  10262.5 93182.5 10512.5 93247.5 ;
      RECT  10480.0 93202.5 10545.0 93215.0 ;
      RECT  10512.5 93170.0 10760.0 93235.0 ;
      RECT  8930.0 94605.0 9280.0 94670.0 ;
      RECT  9445.0 94592.5 9510.0 94657.5 ;
      RECT  9445.0 94605.0 9510.0 94670.0 ;
      RECT  9445.0 94625.0 9510.0 94670.0 ;
      RECT  9477.5 94592.5 9775.0 94657.5 ;
      RECT  9775.0 94592.5 9910.0 94657.5 ;
      RECT  10480.0 94592.5 10545.0 94657.5 ;
      RECT  10480.0 94605.0 10545.0 94670.0 ;
      RECT  10262.5 94592.5 10512.5 94657.5 ;
      RECT  10480.0 94625.0 10545.0 94637.5 ;
      RECT  10512.5 94605.0 10760.0 94670.0 ;
      RECT  8930.0 95860.0 9280.0 95925.0 ;
      RECT  9445.0 95872.5 9510.0 95937.5 ;
      RECT  9445.0 95860.0 9510.0 95925.0 ;
      RECT  9445.0 95905.0 9510.0 95925.0 ;
      RECT  9477.5 95872.5 9775.0 95937.5 ;
      RECT  9775.0 95872.5 9910.0 95937.5 ;
      RECT  10480.0 95872.5 10545.0 95937.5 ;
      RECT  10480.0 95860.0 10545.0 95925.0 ;
      RECT  10262.5 95872.5 10512.5 95937.5 ;
      RECT  10480.0 95892.5 10545.0 95905.0 ;
      RECT  10512.5 95860.0 10760.0 95925.0 ;
      RECT  8930.0 97295.0 9280.0 97360.0 ;
      RECT  9445.0 97282.5 9510.0 97347.5 ;
      RECT  9445.0 97295.0 9510.0 97360.0 ;
      RECT  9445.0 97315.0 9510.0 97360.0 ;
      RECT  9477.5 97282.5 9775.0 97347.5 ;
      RECT  9775.0 97282.5 9910.0 97347.5 ;
      RECT  10480.0 97282.5 10545.0 97347.5 ;
      RECT  10480.0 97295.0 10545.0 97360.0 ;
      RECT  10262.5 97282.5 10512.5 97347.5 ;
      RECT  10480.0 97315.0 10545.0 97327.5 ;
      RECT  10512.5 97295.0 10760.0 97360.0 ;
      RECT  8930.0 98550.0 9280.0 98615.0 ;
      RECT  9445.0 98562.5 9510.0 98627.5 ;
      RECT  9445.0 98550.0 9510.0 98615.0 ;
      RECT  9445.0 98595.0 9510.0 98615.0 ;
      RECT  9477.5 98562.5 9775.0 98627.5 ;
      RECT  9775.0 98562.5 9910.0 98627.5 ;
      RECT  10480.0 98562.5 10545.0 98627.5 ;
      RECT  10480.0 98550.0 10545.0 98615.0 ;
      RECT  10262.5 98562.5 10512.5 98627.5 ;
      RECT  10480.0 98582.5 10545.0 98595.0 ;
      RECT  10512.5 98550.0 10760.0 98615.0 ;
      RECT  8930.0 99985.0 9280.0 100050.0 ;
      RECT  9445.0 99972.5 9510.0 100037.5 ;
      RECT  9445.0 99985.0 9510.0 100050.0 ;
      RECT  9445.0 100005.0 9510.0 100050.0 ;
      RECT  9477.5 99972.5 9775.0 100037.5 ;
      RECT  9775.0 99972.5 9910.0 100037.5 ;
      RECT  10480.0 99972.5 10545.0 100037.5 ;
      RECT  10480.0 99985.0 10545.0 100050.0 ;
      RECT  10262.5 99972.5 10512.5 100037.5 ;
      RECT  10480.0 100005.0 10545.0 100017.5 ;
      RECT  10512.5 99985.0 10760.0 100050.0 ;
      RECT  8930.0 101240.0 9280.0 101305.0 ;
      RECT  9445.0 101252.5 9510.0 101317.5 ;
      RECT  9445.0 101240.0 9510.0 101305.0 ;
      RECT  9445.0 101285.0 9510.0 101305.0 ;
      RECT  9477.5 101252.5 9775.0 101317.5 ;
      RECT  9775.0 101252.5 9910.0 101317.5 ;
      RECT  10480.0 101252.5 10545.0 101317.5 ;
      RECT  10480.0 101240.0 10545.0 101305.0 ;
      RECT  10262.5 101252.5 10512.5 101317.5 ;
      RECT  10480.0 101272.5 10545.0 101285.0 ;
      RECT  10512.5 101240.0 10760.0 101305.0 ;
      RECT  8930.0 102675.0 9280.0 102740.0 ;
      RECT  9445.0 102662.5 9510.0 102727.5 ;
      RECT  9445.0 102675.0 9510.0 102740.0 ;
      RECT  9445.0 102695.0 9510.0 102740.0 ;
      RECT  9477.5 102662.5 9775.0 102727.5 ;
      RECT  9775.0 102662.5 9910.0 102727.5 ;
      RECT  10480.0 102662.5 10545.0 102727.5 ;
      RECT  10480.0 102675.0 10545.0 102740.0 ;
      RECT  10262.5 102662.5 10512.5 102727.5 ;
      RECT  10480.0 102695.0 10545.0 102707.5 ;
      RECT  10512.5 102675.0 10760.0 102740.0 ;
      RECT  8930.0 103930.0 9280.0 103995.0 ;
      RECT  9445.0 103942.5 9510.0 104007.5 ;
      RECT  9445.0 103930.0 9510.0 103995.0 ;
      RECT  9445.0 103975.0 9510.0 103995.0 ;
      RECT  9477.5 103942.5 9775.0 104007.5 ;
      RECT  9775.0 103942.5 9910.0 104007.5 ;
      RECT  10480.0 103942.5 10545.0 104007.5 ;
      RECT  10480.0 103930.0 10545.0 103995.0 ;
      RECT  10262.5 103942.5 10512.5 104007.5 ;
      RECT  10480.0 103962.5 10545.0 103975.0 ;
      RECT  10512.5 103930.0 10760.0 103995.0 ;
      RECT  8930.0 105365.0 9280.0 105430.0 ;
      RECT  9445.0 105352.5 9510.0 105417.5 ;
      RECT  9445.0 105365.0 9510.0 105430.0 ;
      RECT  9445.0 105385.0 9510.0 105430.0 ;
      RECT  9477.5 105352.5 9775.0 105417.5 ;
      RECT  9775.0 105352.5 9910.0 105417.5 ;
      RECT  10480.0 105352.5 10545.0 105417.5 ;
      RECT  10480.0 105365.0 10545.0 105430.0 ;
      RECT  10262.5 105352.5 10512.5 105417.5 ;
      RECT  10480.0 105385.0 10545.0 105397.5 ;
      RECT  10512.5 105365.0 10760.0 105430.0 ;
      RECT  8930.0 106620.0 9280.0 106685.0 ;
      RECT  9445.0 106632.5 9510.0 106697.5 ;
      RECT  9445.0 106620.0 9510.0 106685.0 ;
      RECT  9445.0 106665.0 9510.0 106685.0 ;
      RECT  9477.5 106632.5 9775.0 106697.5 ;
      RECT  9775.0 106632.5 9910.0 106697.5 ;
      RECT  10480.0 106632.5 10545.0 106697.5 ;
      RECT  10480.0 106620.0 10545.0 106685.0 ;
      RECT  10262.5 106632.5 10512.5 106697.5 ;
      RECT  10480.0 106652.5 10545.0 106665.0 ;
      RECT  10512.5 106620.0 10760.0 106685.0 ;
      RECT  8930.0 108055.0 9280.0 108120.0 ;
      RECT  9445.0 108042.5 9510.0 108107.5 ;
      RECT  9445.0 108055.0 9510.0 108120.0 ;
      RECT  9445.0 108075.0 9510.0 108120.0 ;
      RECT  9477.5 108042.5 9775.0 108107.5 ;
      RECT  9775.0 108042.5 9910.0 108107.5 ;
      RECT  10480.0 108042.5 10545.0 108107.5 ;
      RECT  10480.0 108055.0 10545.0 108120.0 ;
      RECT  10262.5 108042.5 10512.5 108107.5 ;
      RECT  10480.0 108075.0 10545.0 108087.5 ;
      RECT  10512.5 108055.0 10760.0 108120.0 ;
      RECT  8930.0 109310.0 9280.0 109375.0 ;
      RECT  9445.0 109322.5 9510.0 109387.5 ;
      RECT  9445.0 109310.0 9510.0 109375.0 ;
      RECT  9445.0 109355.0 9510.0 109375.0 ;
      RECT  9477.5 109322.5 9775.0 109387.5 ;
      RECT  9775.0 109322.5 9910.0 109387.5 ;
      RECT  10480.0 109322.5 10545.0 109387.5 ;
      RECT  10480.0 109310.0 10545.0 109375.0 ;
      RECT  10262.5 109322.5 10512.5 109387.5 ;
      RECT  10480.0 109342.5 10545.0 109355.0 ;
      RECT  10512.5 109310.0 10760.0 109375.0 ;
      RECT  8930.0 110745.0 9280.0 110810.0 ;
      RECT  9445.0 110732.5 9510.0 110797.5 ;
      RECT  9445.0 110745.0 9510.0 110810.0 ;
      RECT  9445.0 110765.0 9510.0 110810.0 ;
      RECT  9477.5 110732.5 9775.0 110797.5 ;
      RECT  9775.0 110732.5 9910.0 110797.5 ;
      RECT  10480.0 110732.5 10545.0 110797.5 ;
      RECT  10480.0 110745.0 10545.0 110810.0 ;
      RECT  10262.5 110732.5 10512.5 110797.5 ;
      RECT  10480.0 110765.0 10545.0 110777.5 ;
      RECT  10512.5 110745.0 10760.0 110810.0 ;
      RECT  8930.0 112000.0 9280.0 112065.0 ;
      RECT  9445.0 112012.5 9510.0 112077.5 ;
      RECT  9445.0 112000.0 9510.0 112065.0 ;
      RECT  9445.0 112045.0 9510.0 112065.0 ;
      RECT  9477.5 112012.5 9775.0 112077.5 ;
      RECT  9775.0 112012.5 9910.0 112077.5 ;
      RECT  10480.0 112012.5 10545.0 112077.5 ;
      RECT  10480.0 112000.0 10545.0 112065.0 ;
      RECT  10262.5 112012.5 10512.5 112077.5 ;
      RECT  10480.0 112032.5 10545.0 112045.0 ;
      RECT  10512.5 112000.0 10760.0 112065.0 ;
      RECT  8930.0 113435.0 9280.0 113500.0 ;
      RECT  9445.0 113422.5 9510.0 113487.5 ;
      RECT  9445.0 113435.0 9510.0 113500.0 ;
      RECT  9445.0 113455.0 9510.0 113500.0 ;
      RECT  9477.5 113422.5 9775.0 113487.5 ;
      RECT  9775.0 113422.5 9910.0 113487.5 ;
      RECT  10480.0 113422.5 10545.0 113487.5 ;
      RECT  10480.0 113435.0 10545.0 113500.0 ;
      RECT  10262.5 113422.5 10512.5 113487.5 ;
      RECT  10480.0 113455.0 10545.0 113467.5 ;
      RECT  10512.5 113435.0 10760.0 113500.0 ;
      RECT  9582.5 29175.0 9647.5 29360.0 ;
      RECT  9582.5 28015.0 9647.5 28200.0 ;
      RECT  9222.5 28132.5 9287.5 27982.5 ;
      RECT  9222.5 29017.5 9287.5 29392.5 ;
      RECT  9412.5 28132.5 9477.5 29017.5 ;
      RECT  9222.5 29017.5 9287.5 29152.5 ;
      RECT  9412.5 29017.5 9477.5 29152.5 ;
      RECT  9412.5 29017.5 9477.5 29152.5 ;
      RECT  9222.5 29017.5 9287.5 29152.5 ;
      RECT  9222.5 28132.5 9287.5 28267.5 ;
      RECT  9412.5 28132.5 9477.5 28267.5 ;
      RECT  9412.5 28132.5 9477.5 28267.5 ;
      RECT  9222.5 28132.5 9287.5 28267.5 ;
      RECT  9582.5 29107.5 9647.5 29242.5 ;
      RECT  9582.5 28132.5 9647.5 28267.5 ;
      RECT  9280.0 28575.0 9345.0 28710.0 ;
      RECT  9280.0 28575.0 9345.0 28710.0 ;
      RECT  9445.0 28610.0 9510.0 28675.0 ;
      RECT  9155.0 29327.5 9715.0 29392.5 ;
      RECT  9155.0 27982.5 9715.0 28047.5 ;
      RECT  9782.5 28177.5 9847.5 27982.5 ;
      RECT  9782.5 29017.5 9847.5 29392.5 ;
      RECT  10162.5 29017.5 10227.5 29392.5 ;
      RECT  10332.5 29175.0 10397.5 29360.0 ;
      RECT  10332.5 28015.0 10397.5 28200.0 ;
      RECT  9782.5 29017.5 9847.5 29152.5 ;
      RECT  9972.5 29017.5 10037.5 29152.5 ;
      RECT  9972.5 29017.5 10037.5 29152.5 ;
      RECT  9782.5 29017.5 9847.5 29152.5 ;
      RECT  9972.5 29017.5 10037.5 29152.5 ;
      RECT  10162.5 29017.5 10227.5 29152.5 ;
      RECT  10162.5 29017.5 10227.5 29152.5 ;
      RECT  9972.5 29017.5 10037.5 29152.5 ;
      RECT  9782.5 28177.5 9847.5 28312.5 ;
      RECT  9972.5 28177.5 10037.5 28312.5 ;
      RECT  9972.5 28177.5 10037.5 28312.5 ;
      RECT  9782.5 28177.5 9847.5 28312.5 ;
      RECT  9972.5 28177.5 10037.5 28312.5 ;
      RECT  10162.5 28177.5 10227.5 28312.5 ;
      RECT  10162.5 28177.5 10227.5 28312.5 ;
      RECT  9972.5 28177.5 10037.5 28312.5 ;
      RECT  10332.5 29107.5 10397.5 29242.5 ;
      RECT  10332.5 28132.5 10397.5 28267.5 ;
      RECT  10167.5 28407.5 10032.5 28472.5 ;
      RECT  9910.0 28622.5 9775.0 28687.5 ;
      RECT  9972.5 29017.5 10037.5 29152.5 ;
      RECT  10162.5 28177.5 10227.5 28312.5 ;
      RECT  10262.5 28622.5 10127.5 28687.5 ;
      RECT  9775.0 28622.5 9910.0 28687.5 ;
      RECT  10032.5 28407.5 10167.5 28472.5 ;
      RECT  10127.5 28622.5 10262.5 28687.5 ;
      RECT  9715.0 29327.5 10635.0 29392.5 ;
      RECT  9715.0 27982.5 10635.0 28047.5 ;
      RECT  11062.5 29175.0 11127.5 29360.0 ;
      RECT  11062.5 28015.0 11127.5 28200.0 ;
      RECT  10702.5 28132.5 10767.5 27982.5 ;
      RECT  10702.5 29017.5 10767.5 29392.5 ;
      RECT  10892.5 28132.5 10957.5 29017.5 ;
      RECT  10702.5 29017.5 10767.5 29152.5 ;
      RECT  10892.5 29017.5 10957.5 29152.5 ;
      RECT  10892.5 29017.5 10957.5 29152.5 ;
      RECT  10702.5 29017.5 10767.5 29152.5 ;
      RECT  10702.5 28132.5 10767.5 28267.5 ;
      RECT  10892.5 28132.5 10957.5 28267.5 ;
      RECT  10892.5 28132.5 10957.5 28267.5 ;
      RECT  10702.5 28132.5 10767.5 28267.5 ;
      RECT  11062.5 29107.5 11127.5 29242.5 ;
      RECT  11062.5 28132.5 11127.5 28267.5 ;
      RECT  10760.0 28575.0 10825.0 28710.0 ;
      RECT  10760.0 28575.0 10825.0 28710.0 ;
      RECT  10925.0 28610.0 10990.0 28675.0 ;
      RECT  10635.0 29327.5 11195.0 29392.5 ;
      RECT  10635.0 27982.5 11195.0 28047.5 ;
      RECT  8897.5 28575.0 8962.5 28710.0 ;
      RECT  9037.5 28302.5 9102.5 28437.5 ;
      RECT  10032.5 28407.5 9897.5 28472.5 ;
      RECT  9582.5 29545.0 9647.5 29360.0 ;
      RECT  9582.5 30705.0 9647.5 30520.0 ;
      RECT  9222.5 30587.5 9287.5 30737.5 ;
      RECT  9222.5 29702.5 9287.5 29327.5 ;
      RECT  9412.5 30587.5 9477.5 29702.5 ;
      RECT  9222.5 29702.5 9287.5 29567.5 ;
      RECT  9412.5 29702.5 9477.5 29567.5 ;
      RECT  9412.5 29702.5 9477.5 29567.5 ;
      RECT  9222.5 29702.5 9287.5 29567.5 ;
      RECT  9222.5 30587.5 9287.5 30452.5 ;
      RECT  9412.5 30587.5 9477.5 30452.5 ;
      RECT  9412.5 30587.5 9477.5 30452.5 ;
      RECT  9222.5 30587.5 9287.5 30452.5 ;
      RECT  9582.5 29612.5 9647.5 29477.5 ;
      RECT  9582.5 30587.5 9647.5 30452.5 ;
      RECT  9280.0 30145.0 9345.0 30010.0 ;
      RECT  9280.0 30145.0 9345.0 30010.0 ;
      RECT  9445.0 30110.0 9510.0 30045.0 ;
      RECT  9155.0 29392.5 9715.0 29327.5 ;
      RECT  9155.0 30737.5 9715.0 30672.5 ;
      RECT  9782.5 30542.5 9847.5 30737.5 ;
      RECT  9782.5 29702.5 9847.5 29327.5 ;
      RECT  10162.5 29702.5 10227.5 29327.5 ;
      RECT  10332.5 29545.0 10397.5 29360.0 ;
      RECT  10332.5 30705.0 10397.5 30520.0 ;
      RECT  9782.5 29702.5 9847.5 29567.5 ;
      RECT  9972.5 29702.5 10037.5 29567.5 ;
      RECT  9972.5 29702.5 10037.5 29567.5 ;
      RECT  9782.5 29702.5 9847.5 29567.5 ;
      RECT  9972.5 29702.5 10037.5 29567.5 ;
      RECT  10162.5 29702.5 10227.5 29567.5 ;
      RECT  10162.5 29702.5 10227.5 29567.5 ;
      RECT  9972.5 29702.5 10037.5 29567.5 ;
      RECT  9782.5 30542.5 9847.5 30407.5 ;
      RECT  9972.5 30542.5 10037.5 30407.5 ;
      RECT  9972.5 30542.5 10037.5 30407.5 ;
      RECT  9782.5 30542.5 9847.5 30407.5 ;
      RECT  9972.5 30542.5 10037.5 30407.5 ;
      RECT  10162.5 30542.5 10227.5 30407.5 ;
      RECT  10162.5 30542.5 10227.5 30407.5 ;
      RECT  9972.5 30542.5 10037.5 30407.5 ;
      RECT  10332.5 29612.5 10397.5 29477.5 ;
      RECT  10332.5 30587.5 10397.5 30452.5 ;
      RECT  10167.5 30312.5 10032.5 30247.5 ;
      RECT  9910.0 30097.5 9775.0 30032.5 ;
      RECT  9972.5 29702.5 10037.5 29567.5 ;
      RECT  10162.5 30542.5 10227.5 30407.5 ;
      RECT  10262.5 30097.5 10127.5 30032.5 ;
      RECT  9775.0 30097.5 9910.0 30032.5 ;
      RECT  10032.5 30312.5 10167.5 30247.5 ;
      RECT  10127.5 30097.5 10262.5 30032.5 ;
      RECT  9715.0 29392.5 10635.0 29327.5 ;
      RECT  9715.0 30737.5 10635.0 30672.5 ;
      RECT  11062.5 29545.0 11127.5 29360.0 ;
      RECT  11062.5 30705.0 11127.5 30520.0 ;
      RECT  10702.5 30587.5 10767.5 30737.5 ;
      RECT  10702.5 29702.5 10767.5 29327.5 ;
      RECT  10892.5 30587.5 10957.5 29702.5 ;
      RECT  10702.5 29702.5 10767.5 29567.5 ;
      RECT  10892.5 29702.5 10957.5 29567.5 ;
      RECT  10892.5 29702.5 10957.5 29567.5 ;
      RECT  10702.5 29702.5 10767.5 29567.5 ;
      RECT  10702.5 30587.5 10767.5 30452.5 ;
      RECT  10892.5 30587.5 10957.5 30452.5 ;
      RECT  10892.5 30587.5 10957.5 30452.5 ;
      RECT  10702.5 30587.5 10767.5 30452.5 ;
      RECT  11062.5 29612.5 11127.5 29477.5 ;
      RECT  11062.5 30587.5 11127.5 30452.5 ;
      RECT  10760.0 30145.0 10825.0 30010.0 ;
      RECT  10760.0 30145.0 10825.0 30010.0 ;
      RECT  10925.0 30110.0 10990.0 30045.0 ;
      RECT  10635.0 29392.5 11195.0 29327.5 ;
      RECT  10635.0 30737.5 11195.0 30672.5 ;
      RECT  8897.5 30010.0 8962.5 30145.0 ;
      RECT  9037.5 30282.5 9102.5 30417.5 ;
      RECT  10032.5 30247.5 9897.5 30312.5 ;
      RECT  9582.5 31865.0 9647.5 32050.0 ;
      RECT  9582.5 30705.0 9647.5 30890.0 ;
      RECT  9222.5 30822.5 9287.5 30672.5 ;
      RECT  9222.5 31707.5 9287.5 32082.5 ;
      RECT  9412.5 30822.5 9477.5 31707.5 ;
      RECT  9222.5 31707.5 9287.5 31842.5 ;
      RECT  9412.5 31707.5 9477.5 31842.5 ;
      RECT  9412.5 31707.5 9477.5 31842.5 ;
      RECT  9222.5 31707.5 9287.5 31842.5 ;
      RECT  9222.5 30822.5 9287.5 30957.5 ;
      RECT  9412.5 30822.5 9477.5 30957.5 ;
      RECT  9412.5 30822.5 9477.5 30957.5 ;
      RECT  9222.5 30822.5 9287.5 30957.5 ;
      RECT  9582.5 31797.5 9647.5 31932.5 ;
      RECT  9582.5 30822.5 9647.5 30957.5 ;
      RECT  9280.0 31265.0 9345.0 31400.0 ;
      RECT  9280.0 31265.0 9345.0 31400.0 ;
      RECT  9445.0 31300.0 9510.0 31365.0 ;
      RECT  9155.0 32017.5 9715.0 32082.5 ;
      RECT  9155.0 30672.5 9715.0 30737.5 ;
      RECT  9782.5 30867.5 9847.5 30672.5 ;
      RECT  9782.5 31707.5 9847.5 32082.5 ;
      RECT  10162.5 31707.5 10227.5 32082.5 ;
      RECT  10332.5 31865.0 10397.5 32050.0 ;
      RECT  10332.5 30705.0 10397.5 30890.0 ;
      RECT  9782.5 31707.5 9847.5 31842.5 ;
      RECT  9972.5 31707.5 10037.5 31842.5 ;
      RECT  9972.5 31707.5 10037.5 31842.5 ;
      RECT  9782.5 31707.5 9847.5 31842.5 ;
      RECT  9972.5 31707.5 10037.5 31842.5 ;
      RECT  10162.5 31707.5 10227.5 31842.5 ;
      RECT  10162.5 31707.5 10227.5 31842.5 ;
      RECT  9972.5 31707.5 10037.5 31842.5 ;
      RECT  9782.5 30867.5 9847.5 31002.5 ;
      RECT  9972.5 30867.5 10037.5 31002.5 ;
      RECT  9972.5 30867.5 10037.5 31002.5 ;
      RECT  9782.5 30867.5 9847.5 31002.5 ;
      RECT  9972.5 30867.5 10037.5 31002.5 ;
      RECT  10162.5 30867.5 10227.5 31002.5 ;
      RECT  10162.5 30867.5 10227.5 31002.5 ;
      RECT  9972.5 30867.5 10037.5 31002.5 ;
      RECT  10332.5 31797.5 10397.5 31932.5 ;
      RECT  10332.5 30822.5 10397.5 30957.5 ;
      RECT  10167.5 31097.5 10032.5 31162.5 ;
      RECT  9910.0 31312.5 9775.0 31377.5 ;
      RECT  9972.5 31707.5 10037.5 31842.5 ;
      RECT  10162.5 30867.5 10227.5 31002.5 ;
      RECT  10262.5 31312.5 10127.5 31377.5 ;
      RECT  9775.0 31312.5 9910.0 31377.5 ;
      RECT  10032.5 31097.5 10167.5 31162.5 ;
      RECT  10127.5 31312.5 10262.5 31377.5 ;
      RECT  9715.0 32017.5 10635.0 32082.5 ;
      RECT  9715.0 30672.5 10635.0 30737.5 ;
      RECT  11062.5 31865.0 11127.5 32050.0 ;
      RECT  11062.5 30705.0 11127.5 30890.0 ;
      RECT  10702.5 30822.5 10767.5 30672.5 ;
      RECT  10702.5 31707.5 10767.5 32082.5 ;
      RECT  10892.5 30822.5 10957.5 31707.5 ;
      RECT  10702.5 31707.5 10767.5 31842.5 ;
      RECT  10892.5 31707.5 10957.5 31842.5 ;
      RECT  10892.5 31707.5 10957.5 31842.5 ;
      RECT  10702.5 31707.5 10767.5 31842.5 ;
      RECT  10702.5 30822.5 10767.5 30957.5 ;
      RECT  10892.5 30822.5 10957.5 30957.5 ;
      RECT  10892.5 30822.5 10957.5 30957.5 ;
      RECT  10702.5 30822.5 10767.5 30957.5 ;
      RECT  11062.5 31797.5 11127.5 31932.5 ;
      RECT  11062.5 30822.5 11127.5 30957.5 ;
      RECT  10760.0 31265.0 10825.0 31400.0 ;
      RECT  10760.0 31265.0 10825.0 31400.0 ;
      RECT  10925.0 31300.0 10990.0 31365.0 ;
      RECT  10635.0 32017.5 11195.0 32082.5 ;
      RECT  10635.0 30672.5 11195.0 30737.5 ;
      RECT  8897.5 31265.0 8962.5 31400.0 ;
      RECT  9037.5 30992.5 9102.5 31127.5 ;
      RECT  10032.5 31097.5 9897.5 31162.5 ;
      RECT  9582.5 32235.0 9647.5 32050.0 ;
      RECT  9582.5 33395.0 9647.5 33210.0 ;
      RECT  9222.5 33277.5 9287.5 33427.5 ;
      RECT  9222.5 32392.5 9287.5 32017.5 ;
      RECT  9412.5 33277.5 9477.5 32392.5 ;
      RECT  9222.5 32392.5 9287.5 32257.5 ;
      RECT  9412.5 32392.5 9477.5 32257.5 ;
      RECT  9412.5 32392.5 9477.5 32257.5 ;
      RECT  9222.5 32392.5 9287.5 32257.5 ;
      RECT  9222.5 33277.5 9287.5 33142.5 ;
      RECT  9412.5 33277.5 9477.5 33142.5 ;
      RECT  9412.5 33277.5 9477.5 33142.5 ;
      RECT  9222.5 33277.5 9287.5 33142.5 ;
      RECT  9582.5 32302.5 9647.5 32167.5 ;
      RECT  9582.5 33277.5 9647.5 33142.5 ;
      RECT  9280.0 32835.0 9345.0 32700.0 ;
      RECT  9280.0 32835.0 9345.0 32700.0 ;
      RECT  9445.0 32800.0 9510.0 32735.0 ;
      RECT  9155.0 32082.5 9715.0 32017.5 ;
      RECT  9155.0 33427.5 9715.0 33362.5 ;
      RECT  9782.5 33232.5 9847.5 33427.5 ;
      RECT  9782.5 32392.5 9847.5 32017.5 ;
      RECT  10162.5 32392.5 10227.5 32017.5 ;
      RECT  10332.5 32235.0 10397.5 32050.0 ;
      RECT  10332.5 33395.0 10397.5 33210.0 ;
      RECT  9782.5 32392.5 9847.5 32257.5 ;
      RECT  9972.5 32392.5 10037.5 32257.5 ;
      RECT  9972.5 32392.5 10037.5 32257.5 ;
      RECT  9782.5 32392.5 9847.5 32257.5 ;
      RECT  9972.5 32392.5 10037.5 32257.5 ;
      RECT  10162.5 32392.5 10227.5 32257.5 ;
      RECT  10162.5 32392.5 10227.5 32257.5 ;
      RECT  9972.5 32392.5 10037.5 32257.5 ;
      RECT  9782.5 33232.5 9847.5 33097.5 ;
      RECT  9972.5 33232.5 10037.5 33097.5 ;
      RECT  9972.5 33232.5 10037.5 33097.5 ;
      RECT  9782.5 33232.5 9847.5 33097.5 ;
      RECT  9972.5 33232.5 10037.5 33097.5 ;
      RECT  10162.5 33232.5 10227.5 33097.5 ;
      RECT  10162.5 33232.5 10227.5 33097.5 ;
      RECT  9972.5 33232.5 10037.5 33097.5 ;
      RECT  10332.5 32302.5 10397.5 32167.5 ;
      RECT  10332.5 33277.5 10397.5 33142.5 ;
      RECT  10167.5 33002.5 10032.5 32937.5 ;
      RECT  9910.0 32787.5 9775.0 32722.5 ;
      RECT  9972.5 32392.5 10037.5 32257.5 ;
      RECT  10162.5 33232.5 10227.5 33097.5 ;
      RECT  10262.5 32787.5 10127.5 32722.5 ;
      RECT  9775.0 32787.5 9910.0 32722.5 ;
      RECT  10032.5 33002.5 10167.5 32937.5 ;
      RECT  10127.5 32787.5 10262.5 32722.5 ;
      RECT  9715.0 32082.5 10635.0 32017.5 ;
      RECT  9715.0 33427.5 10635.0 33362.5 ;
      RECT  11062.5 32235.0 11127.5 32050.0 ;
      RECT  11062.5 33395.0 11127.5 33210.0 ;
      RECT  10702.5 33277.5 10767.5 33427.5 ;
      RECT  10702.5 32392.5 10767.5 32017.5 ;
      RECT  10892.5 33277.5 10957.5 32392.5 ;
      RECT  10702.5 32392.5 10767.5 32257.5 ;
      RECT  10892.5 32392.5 10957.5 32257.5 ;
      RECT  10892.5 32392.5 10957.5 32257.5 ;
      RECT  10702.5 32392.5 10767.5 32257.5 ;
      RECT  10702.5 33277.5 10767.5 33142.5 ;
      RECT  10892.5 33277.5 10957.5 33142.5 ;
      RECT  10892.5 33277.5 10957.5 33142.5 ;
      RECT  10702.5 33277.5 10767.5 33142.5 ;
      RECT  11062.5 32302.5 11127.5 32167.5 ;
      RECT  11062.5 33277.5 11127.5 33142.5 ;
      RECT  10760.0 32835.0 10825.0 32700.0 ;
      RECT  10760.0 32835.0 10825.0 32700.0 ;
      RECT  10925.0 32800.0 10990.0 32735.0 ;
      RECT  10635.0 32082.5 11195.0 32017.5 ;
      RECT  10635.0 33427.5 11195.0 33362.5 ;
      RECT  8897.5 32700.0 8962.5 32835.0 ;
      RECT  9037.5 32972.5 9102.5 33107.5 ;
      RECT  10032.5 32937.5 9897.5 33002.5 ;
      RECT  9582.5 34555.0 9647.5 34740.0 ;
      RECT  9582.5 33395.0 9647.5 33580.0 ;
      RECT  9222.5 33512.5 9287.5 33362.5 ;
      RECT  9222.5 34397.5 9287.5 34772.5 ;
      RECT  9412.5 33512.5 9477.5 34397.5 ;
      RECT  9222.5 34397.5 9287.5 34532.5 ;
      RECT  9412.5 34397.5 9477.5 34532.5 ;
      RECT  9412.5 34397.5 9477.5 34532.5 ;
      RECT  9222.5 34397.5 9287.5 34532.5 ;
      RECT  9222.5 33512.5 9287.5 33647.5 ;
      RECT  9412.5 33512.5 9477.5 33647.5 ;
      RECT  9412.5 33512.5 9477.5 33647.5 ;
      RECT  9222.5 33512.5 9287.5 33647.5 ;
      RECT  9582.5 34487.5 9647.5 34622.5 ;
      RECT  9582.5 33512.5 9647.5 33647.5 ;
      RECT  9280.0 33955.0 9345.0 34090.0 ;
      RECT  9280.0 33955.0 9345.0 34090.0 ;
      RECT  9445.0 33990.0 9510.0 34055.0 ;
      RECT  9155.0 34707.5 9715.0 34772.5 ;
      RECT  9155.0 33362.5 9715.0 33427.5 ;
      RECT  9782.5 33557.5 9847.5 33362.5 ;
      RECT  9782.5 34397.5 9847.5 34772.5 ;
      RECT  10162.5 34397.5 10227.5 34772.5 ;
      RECT  10332.5 34555.0 10397.5 34740.0 ;
      RECT  10332.5 33395.0 10397.5 33580.0 ;
      RECT  9782.5 34397.5 9847.5 34532.5 ;
      RECT  9972.5 34397.5 10037.5 34532.5 ;
      RECT  9972.5 34397.5 10037.5 34532.5 ;
      RECT  9782.5 34397.5 9847.5 34532.5 ;
      RECT  9972.5 34397.5 10037.5 34532.5 ;
      RECT  10162.5 34397.5 10227.5 34532.5 ;
      RECT  10162.5 34397.5 10227.5 34532.5 ;
      RECT  9972.5 34397.5 10037.5 34532.5 ;
      RECT  9782.5 33557.5 9847.5 33692.5 ;
      RECT  9972.5 33557.5 10037.5 33692.5 ;
      RECT  9972.5 33557.5 10037.5 33692.5 ;
      RECT  9782.5 33557.5 9847.5 33692.5 ;
      RECT  9972.5 33557.5 10037.5 33692.5 ;
      RECT  10162.5 33557.5 10227.5 33692.5 ;
      RECT  10162.5 33557.5 10227.5 33692.5 ;
      RECT  9972.5 33557.5 10037.5 33692.5 ;
      RECT  10332.5 34487.5 10397.5 34622.5 ;
      RECT  10332.5 33512.5 10397.5 33647.5 ;
      RECT  10167.5 33787.5 10032.5 33852.5 ;
      RECT  9910.0 34002.5 9775.0 34067.5 ;
      RECT  9972.5 34397.5 10037.5 34532.5 ;
      RECT  10162.5 33557.5 10227.5 33692.5 ;
      RECT  10262.5 34002.5 10127.5 34067.5 ;
      RECT  9775.0 34002.5 9910.0 34067.5 ;
      RECT  10032.5 33787.5 10167.5 33852.5 ;
      RECT  10127.5 34002.5 10262.5 34067.5 ;
      RECT  9715.0 34707.5 10635.0 34772.5 ;
      RECT  9715.0 33362.5 10635.0 33427.5 ;
      RECT  11062.5 34555.0 11127.5 34740.0 ;
      RECT  11062.5 33395.0 11127.5 33580.0 ;
      RECT  10702.5 33512.5 10767.5 33362.5 ;
      RECT  10702.5 34397.5 10767.5 34772.5 ;
      RECT  10892.5 33512.5 10957.5 34397.5 ;
      RECT  10702.5 34397.5 10767.5 34532.5 ;
      RECT  10892.5 34397.5 10957.5 34532.5 ;
      RECT  10892.5 34397.5 10957.5 34532.5 ;
      RECT  10702.5 34397.5 10767.5 34532.5 ;
      RECT  10702.5 33512.5 10767.5 33647.5 ;
      RECT  10892.5 33512.5 10957.5 33647.5 ;
      RECT  10892.5 33512.5 10957.5 33647.5 ;
      RECT  10702.5 33512.5 10767.5 33647.5 ;
      RECT  11062.5 34487.5 11127.5 34622.5 ;
      RECT  11062.5 33512.5 11127.5 33647.5 ;
      RECT  10760.0 33955.0 10825.0 34090.0 ;
      RECT  10760.0 33955.0 10825.0 34090.0 ;
      RECT  10925.0 33990.0 10990.0 34055.0 ;
      RECT  10635.0 34707.5 11195.0 34772.5 ;
      RECT  10635.0 33362.5 11195.0 33427.5 ;
      RECT  8897.5 33955.0 8962.5 34090.0 ;
      RECT  9037.5 33682.5 9102.5 33817.5 ;
      RECT  10032.5 33787.5 9897.5 33852.5 ;
      RECT  9582.5 34925.0 9647.5 34740.0 ;
      RECT  9582.5 36085.0 9647.5 35900.0 ;
      RECT  9222.5 35967.5 9287.5 36117.5 ;
      RECT  9222.5 35082.5 9287.5 34707.5 ;
      RECT  9412.5 35967.5 9477.5 35082.5 ;
      RECT  9222.5 35082.5 9287.5 34947.5 ;
      RECT  9412.5 35082.5 9477.5 34947.5 ;
      RECT  9412.5 35082.5 9477.5 34947.5 ;
      RECT  9222.5 35082.5 9287.5 34947.5 ;
      RECT  9222.5 35967.5 9287.5 35832.5 ;
      RECT  9412.5 35967.5 9477.5 35832.5 ;
      RECT  9412.5 35967.5 9477.5 35832.5 ;
      RECT  9222.5 35967.5 9287.5 35832.5 ;
      RECT  9582.5 34992.5 9647.5 34857.5 ;
      RECT  9582.5 35967.5 9647.5 35832.5 ;
      RECT  9280.0 35525.0 9345.0 35390.0 ;
      RECT  9280.0 35525.0 9345.0 35390.0 ;
      RECT  9445.0 35490.0 9510.0 35425.0 ;
      RECT  9155.0 34772.5 9715.0 34707.5 ;
      RECT  9155.0 36117.5 9715.0 36052.5 ;
      RECT  9782.5 35922.5 9847.5 36117.5 ;
      RECT  9782.5 35082.5 9847.5 34707.5 ;
      RECT  10162.5 35082.5 10227.5 34707.5 ;
      RECT  10332.5 34925.0 10397.5 34740.0 ;
      RECT  10332.5 36085.0 10397.5 35900.0 ;
      RECT  9782.5 35082.5 9847.5 34947.5 ;
      RECT  9972.5 35082.5 10037.5 34947.5 ;
      RECT  9972.5 35082.5 10037.5 34947.5 ;
      RECT  9782.5 35082.5 9847.5 34947.5 ;
      RECT  9972.5 35082.5 10037.5 34947.5 ;
      RECT  10162.5 35082.5 10227.5 34947.5 ;
      RECT  10162.5 35082.5 10227.5 34947.5 ;
      RECT  9972.5 35082.5 10037.5 34947.5 ;
      RECT  9782.5 35922.5 9847.5 35787.5 ;
      RECT  9972.5 35922.5 10037.5 35787.5 ;
      RECT  9972.5 35922.5 10037.5 35787.5 ;
      RECT  9782.5 35922.5 9847.5 35787.5 ;
      RECT  9972.5 35922.5 10037.5 35787.5 ;
      RECT  10162.5 35922.5 10227.5 35787.5 ;
      RECT  10162.5 35922.5 10227.5 35787.5 ;
      RECT  9972.5 35922.5 10037.5 35787.5 ;
      RECT  10332.5 34992.5 10397.5 34857.5 ;
      RECT  10332.5 35967.5 10397.5 35832.5 ;
      RECT  10167.5 35692.5 10032.5 35627.5 ;
      RECT  9910.0 35477.5 9775.0 35412.5 ;
      RECT  9972.5 35082.5 10037.5 34947.5 ;
      RECT  10162.5 35922.5 10227.5 35787.5 ;
      RECT  10262.5 35477.5 10127.5 35412.5 ;
      RECT  9775.0 35477.5 9910.0 35412.5 ;
      RECT  10032.5 35692.5 10167.5 35627.5 ;
      RECT  10127.5 35477.5 10262.5 35412.5 ;
      RECT  9715.0 34772.5 10635.0 34707.5 ;
      RECT  9715.0 36117.5 10635.0 36052.5 ;
      RECT  11062.5 34925.0 11127.5 34740.0 ;
      RECT  11062.5 36085.0 11127.5 35900.0 ;
      RECT  10702.5 35967.5 10767.5 36117.5 ;
      RECT  10702.5 35082.5 10767.5 34707.5 ;
      RECT  10892.5 35967.5 10957.5 35082.5 ;
      RECT  10702.5 35082.5 10767.5 34947.5 ;
      RECT  10892.5 35082.5 10957.5 34947.5 ;
      RECT  10892.5 35082.5 10957.5 34947.5 ;
      RECT  10702.5 35082.5 10767.5 34947.5 ;
      RECT  10702.5 35967.5 10767.5 35832.5 ;
      RECT  10892.5 35967.5 10957.5 35832.5 ;
      RECT  10892.5 35967.5 10957.5 35832.5 ;
      RECT  10702.5 35967.5 10767.5 35832.5 ;
      RECT  11062.5 34992.5 11127.5 34857.5 ;
      RECT  11062.5 35967.5 11127.5 35832.5 ;
      RECT  10760.0 35525.0 10825.0 35390.0 ;
      RECT  10760.0 35525.0 10825.0 35390.0 ;
      RECT  10925.0 35490.0 10990.0 35425.0 ;
      RECT  10635.0 34772.5 11195.0 34707.5 ;
      RECT  10635.0 36117.5 11195.0 36052.5 ;
      RECT  8897.5 35390.0 8962.5 35525.0 ;
      RECT  9037.5 35662.5 9102.5 35797.5 ;
      RECT  10032.5 35627.5 9897.5 35692.5 ;
      RECT  9582.5 37245.0 9647.5 37430.0 ;
      RECT  9582.5 36085.0 9647.5 36270.0 ;
      RECT  9222.5 36202.5 9287.5 36052.5 ;
      RECT  9222.5 37087.5 9287.5 37462.5 ;
      RECT  9412.5 36202.5 9477.5 37087.5 ;
      RECT  9222.5 37087.5 9287.5 37222.5 ;
      RECT  9412.5 37087.5 9477.5 37222.5 ;
      RECT  9412.5 37087.5 9477.5 37222.5 ;
      RECT  9222.5 37087.5 9287.5 37222.5 ;
      RECT  9222.5 36202.5 9287.5 36337.5 ;
      RECT  9412.5 36202.5 9477.5 36337.5 ;
      RECT  9412.5 36202.5 9477.5 36337.5 ;
      RECT  9222.5 36202.5 9287.5 36337.5 ;
      RECT  9582.5 37177.5 9647.5 37312.5 ;
      RECT  9582.5 36202.5 9647.5 36337.5 ;
      RECT  9280.0 36645.0 9345.0 36780.0 ;
      RECT  9280.0 36645.0 9345.0 36780.0 ;
      RECT  9445.0 36680.0 9510.0 36745.0 ;
      RECT  9155.0 37397.5 9715.0 37462.5 ;
      RECT  9155.0 36052.5 9715.0 36117.5 ;
      RECT  9782.5 36247.5 9847.5 36052.5 ;
      RECT  9782.5 37087.5 9847.5 37462.5 ;
      RECT  10162.5 37087.5 10227.5 37462.5 ;
      RECT  10332.5 37245.0 10397.5 37430.0 ;
      RECT  10332.5 36085.0 10397.5 36270.0 ;
      RECT  9782.5 37087.5 9847.5 37222.5 ;
      RECT  9972.5 37087.5 10037.5 37222.5 ;
      RECT  9972.5 37087.5 10037.5 37222.5 ;
      RECT  9782.5 37087.5 9847.5 37222.5 ;
      RECT  9972.5 37087.5 10037.5 37222.5 ;
      RECT  10162.5 37087.5 10227.5 37222.5 ;
      RECT  10162.5 37087.5 10227.5 37222.5 ;
      RECT  9972.5 37087.5 10037.5 37222.5 ;
      RECT  9782.5 36247.5 9847.5 36382.5 ;
      RECT  9972.5 36247.5 10037.5 36382.5 ;
      RECT  9972.5 36247.5 10037.5 36382.5 ;
      RECT  9782.5 36247.5 9847.5 36382.5 ;
      RECT  9972.5 36247.5 10037.5 36382.5 ;
      RECT  10162.5 36247.5 10227.5 36382.5 ;
      RECT  10162.5 36247.5 10227.5 36382.5 ;
      RECT  9972.5 36247.5 10037.5 36382.5 ;
      RECT  10332.5 37177.5 10397.5 37312.5 ;
      RECT  10332.5 36202.5 10397.5 36337.5 ;
      RECT  10167.5 36477.5 10032.5 36542.5 ;
      RECT  9910.0 36692.5 9775.0 36757.5 ;
      RECT  9972.5 37087.5 10037.5 37222.5 ;
      RECT  10162.5 36247.5 10227.5 36382.5 ;
      RECT  10262.5 36692.5 10127.5 36757.5 ;
      RECT  9775.0 36692.5 9910.0 36757.5 ;
      RECT  10032.5 36477.5 10167.5 36542.5 ;
      RECT  10127.5 36692.5 10262.5 36757.5 ;
      RECT  9715.0 37397.5 10635.0 37462.5 ;
      RECT  9715.0 36052.5 10635.0 36117.5 ;
      RECT  11062.5 37245.0 11127.5 37430.0 ;
      RECT  11062.5 36085.0 11127.5 36270.0 ;
      RECT  10702.5 36202.5 10767.5 36052.5 ;
      RECT  10702.5 37087.5 10767.5 37462.5 ;
      RECT  10892.5 36202.5 10957.5 37087.5 ;
      RECT  10702.5 37087.5 10767.5 37222.5 ;
      RECT  10892.5 37087.5 10957.5 37222.5 ;
      RECT  10892.5 37087.5 10957.5 37222.5 ;
      RECT  10702.5 37087.5 10767.5 37222.5 ;
      RECT  10702.5 36202.5 10767.5 36337.5 ;
      RECT  10892.5 36202.5 10957.5 36337.5 ;
      RECT  10892.5 36202.5 10957.5 36337.5 ;
      RECT  10702.5 36202.5 10767.5 36337.5 ;
      RECT  11062.5 37177.5 11127.5 37312.5 ;
      RECT  11062.5 36202.5 11127.5 36337.5 ;
      RECT  10760.0 36645.0 10825.0 36780.0 ;
      RECT  10760.0 36645.0 10825.0 36780.0 ;
      RECT  10925.0 36680.0 10990.0 36745.0 ;
      RECT  10635.0 37397.5 11195.0 37462.5 ;
      RECT  10635.0 36052.5 11195.0 36117.5 ;
      RECT  8897.5 36645.0 8962.5 36780.0 ;
      RECT  9037.5 36372.5 9102.5 36507.5 ;
      RECT  10032.5 36477.5 9897.5 36542.5 ;
      RECT  9582.5 37615.0 9647.5 37430.0 ;
      RECT  9582.5 38775.0 9647.5 38590.0 ;
      RECT  9222.5 38657.5 9287.5 38807.5 ;
      RECT  9222.5 37772.5 9287.5 37397.5 ;
      RECT  9412.5 38657.5 9477.5 37772.5 ;
      RECT  9222.5 37772.5 9287.5 37637.5 ;
      RECT  9412.5 37772.5 9477.5 37637.5 ;
      RECT  9412.5 37772.5 9477.5 37637.5 ;
      RECT  9222.5 37772.5 9287.5 37637.5 ;
      RECT  9222.5 38657.5 9287.5 38522.5 ;
      RECT  9412.5 38657.5 9477.5 38522.5 ;
      RECT  9412.5 38657.5 9477.5 38522.5 ;
      RECT  9222.5 38657.5 9287.5 38522.5 ;
      RECT  9582.5 37682.5 9647.5 37547.5 ;
      RECT  9582.5 38657.5 9647.5 38522.5 ;
      RECT  9280.0 38215.0 9345.0 38080.0 ;
      RECT  9280.0 38215.0 9345.0 38080.0 ;
      RECT  9445.0 38180.0 9510.0 38115.0 ;
      RECT  9155.0 37462.5 9715.0 37397.5 ;
      RECT  9155.0 38807.5 9715.0 38742.5 ;
      RECT  9782.5 38612.5 9847.5 38807.5 ;
      RECT  9782.5 37772.5 9847.5 37397.5 ;
      RECT  10162.5 37772.5 10227.5 37397.5 ;
      RECT  10332.5 37615.0 10397.5 37430.0 ;
      RECT  10332.5 38775.0 10397.5 38590.0 ;
      RECT  9782.5 37772.5 9847.5 37637.5 ;
      RECT  9972.5 37772.5 10037.5 37637.5 ;
      RECT  9972.5 37772.5 10037.5 37637.5 ;
      RECT  9782.5 37772.5 9847.5 37637.5 ;
      RECT  9972.5 37772.5 10037.5 37637.5 ;
      RECT  10162.5 37772.5 10227.5 37637.5 ;
      RECT  10162.5 37772.5 10227.5 37637.5 ;
      RECT  9972.5 37772.5 10037.5 37637.5 ;
      RECT  9782.5 38612.5 9847.5 38477.5 ;
      RECT  9972.5 38612.5 10037.5 38477.5 ;
      RECT  9972.5 38612.5 10037.5 38477.5 ;
      RECT  9782.5 38612.5 9847.5 38477.5 ;
      RECT  9972.5 38612.5 10037.5 38477.5 ;
      RECT  10162.5 38612.5 10227.5 38477.5 ;
      RECT  10162.5 38612.5 10227.5 38477.5 ;
      RECT  9972.5 38612.5 10037.5 38477.5 ;
      RECT  10332.5 37682.5 10397.5 37547.5 ;
      RECT  10332.5 38657.5 10397.5 38522.5 ;
      RECT  10167.5 38382.5 10032.5 38317.5 ;
      RECT  9910.0 38167.5 9775.0 38102.5 ;
      RECT  9972.5 37772.5 10037.5 37637.5 ;
      RECT  10162.5 38612.5 10227.5 38477.5 ;
      RECT  10262.5 38167.5 10127.5 38102.5 ;
      RECT  9775.0 38167.5 9910.0 38102.5 ;
      RECT  10032.5 38382.5 10167.5 38317.5 ;
      RECT  10127.5 38167.5 10262.5 38102.5 ;
      RECT  9715.0 37462.5 10635.0 37397.5 ;
      RECT  9715.0 38807.5 10635.0 38742.5 ;
      RECT  11062.5 37615.0 11127.5 37430.0 ;
      RECT  11062.5 38775.0 11127.5 38590.0 ;
      RECT  10702.5 38657.5 10767.5 38807.5 ;
      RECT  10702.5 37772.5 10767.5 37397.5 ;
      RECT  10892.5 38657.5 10957.5 37772.5 ;
      RECT  10702.5 37772.5 10767.5 37637.5 ;
      RECT  10892.5 37772.5 10957.5 37637.5 ;
      RECT  10892.5 37772.5 10957.5 37637.5 ;
      RECT  10702.5 37772.5 10767.5 37637.5 ;
      RECT  10702.5 38657.5 10767.5 38522.5 ;
      RECT  10892.5 38657.5 10957.5 38522.5 ;
      RECT  10892.5 38657.5 10957.5 38522.5 ;
      RECT  10702.5 38657.5 10767.5 38522.5 ;
      RECT  11062.5 37682.5 11127.5 37547.5 ;
      RECT  11062.5 38657.5 11127.5 38522.5 ;
      RECT  10760.0 38215.0 10825.0 38080.0 ;
      RECT  10760.0 38215.0 10825.0 38080.0 ;
      RECT  10925.0 38180.0 10990.0 38115.0 ;
      RECT  10635.0 37462.5 11195.0 37397.5 ;
      RECT  10635.0 38807.5 11195.0 38742.5 ;
      RECT  8897.5 38080.0 8962.5 38215.0 ;
      RECT  9037.5 38352.5 9102.5 38487.5 ;
      RECT  10032.5 38317.5 9897.5 38382.5 ;
      RECT  9582.5 39935.0 9647.5 40120.0 ;
      RECT  9582.5 38775.0 9647.5 38960.0 ;
      RECT  9222.5 38892.5 9287.5 38742.5 ;
      RECT  9222.5 39777.5 9287.5 40152.5 ;
      RECT  9412.5 38892.5 9477.5 39777.5 ;
      RECT  9222.5 39777.5 9287.5 39912.5 ;
      RECT  9412.5 39777.5 9477.5 39912.5 ;
      RECT  9412.5 39777.5 9477.5 39912.5 ;
      RECT  9222.5 39777.5 9287.5 39912.5 ;
      RECT  9222.5 38892.5 9287.5 39027.5 ;
      RECT  9412.5 38892.5 9477.5 39027.5 ;
      RECT  9412.5 38892.5 9477.5 39027.5 ;
      RECT  9222.5 38892.5 9287.5 39027.5 ;
      RECT  9582.5 39867.5 9647.5 40002.5 ;
      RECT  9582.5 38892.5 9647.5 39027.5 ;
      RECT  9280.0 39335.0 9345.0 39470.0 ;
      RECT  9280.0 39335.0 9345.0 39470.0 ;
      RECT  9445.0 39370.0 9510.0 39435.0 ;
      RECT  9155.0 40087.5 9715.0 40152.5 ;
      RECT  9155.0 38742.5 9715.0 38807.5 ;
      RECT  9782.5 38937.5 9847.5 38742.5 ;
      RECT  9782.5 39777.5 9847.5 40152.5 ;
      RECT  10162.5 39777.5 10227.5 40152.5 ;
      RECT  10332.5 39935.0 10397.5 40120.0 ;
      RECT  10332.5 38775.0 10397.5 38960.0 ;
      RECT  9782.5 39777.5 9847.5 39912.5 ;
      RECT  9972.5 39777.5 10037.5 39912.5 ;
      RECT  9972.5 39777.5 10037.5 39912.5 ;
      RECT  9782.5 39777.5 9847.5 39912.5 ;
      RECT  9972.5 39777.5 10037.5 39912.5 ;
      RECT  10162.5 39777.5 10227.5 39912.5 ;
      RECT  10162.5 39777.5 10227.5 39912.5 ;
      RECT  9972.5 39777.5 10037.5 39912.5 ;
      RECT  9782.5 38937.5 9847.5 39072.5 ;
      RECT  9972.5 38937.5 10037.5 39072.5 ;
      RECT  9972.5 38937.5 10037.5 39072.5 ;
      RECT  9782.5 38937.5 9847.5 39072.5 ;
      RECT  9972.5 38937.5 10037.5 39072.5 ;
      RECT  10162.5 38937.5 10227.5 39072.5 ;
      RECT  10162.5 38937.5 10227.5 39072.5 ;
      RECT  9972.5 38937.5 10037.5 39072.5 ;
      RECT  10332.5 39867.5 10397.5 40002.5 ;
      RECT  10332.5 38892.5 10397.5 39027.5 ;
      RECT  10167.5 39167.5 10032.5 39232.5 ;
      RECT  9910.0 39382.5 9775.0 39447.5 ;
      RECT  9972.5 39777.5 10037.5 39912.5 ;
      RECT  10162.5 38937.5 10227.5 39072.5 ;
      RECT  10262.5 39382.5 10127.5 39447.5 ;
      RECT  9775.0 39382.5 9910.0 39447.5 ;
      RECT  10032.5 39167.5 10167.5 39232.5 ;
      RECT  10127.5 39382.5 10262.5 39447.5 ;
      RECT  9715.0 40087.5 10635.0 40152.5 ;
      RECT  9715.0 38742.5 10635.0 38807.5 ;
      RECT  11062.5 39935.0 11127.5 40120.0 ;
      RECT  11062.5 38775.0 11127.5 38960.0 ;
      RECT  10702.5 38892.5 10767.5 38742.5 ;
      RECT  10702.5 39777.5 10767.5 40152.5 ;
      RECT  10892.5 38892.5 10957.5 39777.5 ;
      RECT  10702.5 39777.5 10767.5 39912.5 ;
      RECT  10892.5 39777.5 10957.5 39912.5 ;
      RECT  10892.5 39777.5 10957.5 39912.5 ;
      RECT  10702.5 39777.5 10767.5 39912.5 ;
      RECT  10702.5 38892.5 10767.5 39027.5 ;
      RECT  10892.5 38892.5 10957.5 39027.5 ;
      RECT  10892.5 38892.5 10957.5 39027.5 ;
      RECT  10702.5 38892.5 10767.5 39027.5 ;
      RECT  11062.5 39867.5 11127.5 40002.5 ;
      RECT  11062.5 38892.5 11127.5 39027.5 ;
      RECT  10760.0 39335.0 10825.0 39470.0 ;
      RECT  10760.0 39335.0 10825.0 39470.0 ;
      RECT  10925.0 39370.0 10990.0 39435.0 ;
      RECT  10635.0 40087.5 11195.0 40152.5 ;
      RECT  10635.0 38742.5 11195.0 38807.5 ;
      RECT  8897.5 39335.0 8962.5 39470.0 ;
      RECT  9037.5 39062.5 9102.5 39197.5 ;
      RECT  10032.5 39167.5 9897.5 39232.5 ;
      RECT  9582.5 40305.0 9647.5 40120.0 ;
      RECT  9582.5 41465.0 9647.5 41280.0 ;
      RECT  9222.5 41347.5 9287.5 41497.5 ;
      RECT  9222.5 40462.5 9287.5 40087.5 ;
      RECT  9412.5 41347.5 9477.5 40462.5 ;
      RECT  9222.5 40462.5 9287.5 40327.5 ;
      RECT  9412.5 40462.5 9477.5 40327.5 ;
      RECT  9412.5 40462.5 9477.5 40327.5 ;
      RECT  9222.5 40462.5 9287.5 40327.5 ;
      RECT  9222.5 41347.5 9287.5 41212.5 ;
      RECT  9412.5 41347.5 9477.5 41212.5 ;
      RECT  9412.5 41347.5 9477.5 41212.5 ;
      RECT  9222.5 41347.5 9287.5 41212.5 ;
      RECT  9582.5 40372.5 9647.5 40237.5 ;
      RECT  9582.5 41347.5 9647.5 41212.5 ;
      RECT  9280.0 40905.0 9345.0 40770.0 ;
      RECT  9280.0 40905.0 9345.0 40770.0 ;
      RECT  9445.0 40870.0 9510.0 40805.0 ;
      RECT  9155.0 40152.5 9715.0 40087.5 ;
      RECT  9155.0 41497.5 9715.0 41432.5 ;
      RECT  9782.5 41302.5 9847.5 41497.5 ;
      RECT  9782.5 40462.5 9847.5 40087.5 ;
      RECT  10162.5 40462.5 10227.5 40087.5 ;
      RECT  10332.5 40305.0 10397.5 40120.0 ;
      RECT  10332.5 41465.0 10397.5 41280.0 ;
      RECT  9782.5 40462.5 9847.5 40327.5 ;
      RECT  9972.5 40462.5 10037.5 40327.5 ;
      RECT  9972.5 40462.5 10037.5 40327.5 ;
      RECT  9782.5 40462.5 9847.5 40327.5 ;
      RECT  9972.5 40462.5 10037.5 40327.5 ;
      RECT  10162.5 40462.5 10227.5 40327.5 ;
      RECT  10162.5 40462.5 10227.5 40327.5 ;
      RECT  9972.5 40462.5 10037.5 40327.5 ;
      RECT  9782.5 41302.5 9847.5 41167.5 ;
      RECT  9972.5 41302.5 10037.5 41167.5 ;
      RECT  9972.5 41302.5 10037.5 41167.5 ;
      RECT  9782.5 41302.5 9847.5 41167.5 ;
      RECT  9972.5 41302.5 10037.5 41167.5 ;
      RECT  10162.5 41302.5 10227.5 41167.5 ;
      RECT  10162.5 41302.5 10227.5 41167.5 ;
      RECT  9972.5 41302.5 10037.5 41167.5 ;
      RECT  10332.5 40372.5 10397.5 40237.5 ;
      RECT  10332.5 41347.5 10397.5 41212.5 ;
      RECT  10167.5 41072.5 10032.5 41007.5 ;
      RECT  9910.0 40857.5 9775.0 40792.5 ;
      RECT  9972.5 40462.5 10037.5 40327.5 ;
      RECT  10162.5 41302.5 10227.5 41167.5 ;
      RECT  10262.5 40857.5 10127.5 40792.5 ;
      RECT  9775.0 40857.5 9910.0 40792.5 ;
      RECT  10032.5 41072.5 10167.5 41007.5 ;
      RECT  10127.5 40857.5 10262.5 40792.5 ;
      RECT  9715.0 40152.5 10635.0 40087.5 ;
      RECT  9715.0 41497.5 10635.0 41432.5 ;
      RECT  11062.5 40305.0 11127.5 40120.0 ;
      RECT  11062.5 41465.0 11127.5 41280.0 ;
      RECT  10702.5 41347.5 10767.5 41497.5 ;
      RECT  10702.5 40462.5 10767.5 40087.5 ;
      RECT  10892.5 41347.5 10957.5 40462.5 ;
      RECT  10702.5 40462.5 10767.5 40327.5 ;
      RECT  10892.5 40462.5 10957.5 40327.5 ;
      RECT  10892.5 40462.5 10957.5 40327.5 ;
      RECT  10702.5 40462.5 10767.5 40327.5 ;
      RECT  10702.5 41347.5 10767.5 41212.5 ;
      RECT  10892.5 41347.5 10957.5 41212.5 ;
      RECT  10892.5 41347.5 10957.5 41212.5 ;
      RECT  10702.5 41347.5 10767.5 41212.5 ;
      RECT  11062.5 40372.5 11127.5 40237.5 ;
      RECT  11062.5 41347.5 11127.5 41212.5 ;
      RECT  10760.0 40905.0 10825.0 40770.0 ;
      RECT  10760.0 40905.0 10825.0 40770.0 ;
      RECT  10925.0 40870.0 10990.0 40805.0 ;
      RECT  10635.0 40152.5 11195.0 40087.5 ;
      RECT  10635.0 41497.5 11195.0 41432.5 ;
      RECT  8897.5 40770.0 8962.5 40905.0 ;
      RECT  9037.5 41042.5 9102.5 41177.5 ;
      RECT  10032.5 41007.5 9897.5 41072.5 ;
      RECT  9582.5 42625.0 9647.5 42810.0 ;
      RECT  9582.5 41465.0 9647.5 41650.0 ;
      RECT  9222.5 41582.5 9287.5 41432.5 ;
      RECT  9222.5 42467.5 9287.5 42842.5 ;
      RECT  9412.5 41582.5 9477.5 42467.5 ;
      RECT  9222.5 42467.5 9287.5 42602.5 ;
      RECT  9412.5 42467.5 9477.5 42602.5 ;
      RECT  9412.5 42467.5 9477.5 42602.5 ;
      RECT  9222.5 42467.5 9287.5 42602.5 ;
      RECT  9222.5 41582.5 9287.5 41717.5 ;
      RECT  9412.5 41582.5 9477.5 41717.5 ;
      RECT  9412.5 41582.5 9477.5 41717.5 ;
      RECT  9222.5 41582.5 9287.5 41717.5 ;
      RECT  9582.5 42557.5 9647.5 42692.5 ;
      RECT  9582.5 41582.5 9647.5 41717.5 ;
      RECT  9280.0 42025.0 9345.0 42160.0 ;
      RECT  9280.0 42025.0 9345.0 42160.0 ;
      RECT  9445.0 42060.0 9510.0 42125.0 ;
      RECT  9155.0 42777.5 9715.0 42842.5 ;
      RECT  9155.0 41432.5 9715.0 41497.5 ;
      RECT  9782.5 41627.5 9847.5 41432.5 ;
      RECT  9782.5 42467.5 9847.5 42842.5 ;
      RECT  10162.5 42467.5 10227.5 42842.5 ;
      RECT  10332.5 42625.0 10397.5 42810.0 ;
      RECT  10332.5 41465.0 10397.5 41650.0 ;
      RECT  9782.5 42467.5 9847.5 42602.5 ;
      RECT  9972.5 42467.5 10037.5 42602.5 ;
      RECT  9972.5 42467.5 10037.5 42602.5 ;
      RECT  9782.5 42467.5 9847.5 42602.5 ;
      RECT  9972.5 42467.5 10037.5 42602.5 ;
      RECT  10162.5 42467.5 10227.5 42602.5 ;
      RECT  10162.5 42467.5 10227.5 42602.5 ;
      RECT  9972.5 42467.5 10037.5 42602.5 ;
      RECT  9782.5 41627.5 9847.5 41762.5 ;
      RECT  9972.5 41627.5 10037.5 41762.5 ;
      RECT  9972.5 41627.5 10037.5 41762.5 ;
      RECT  9782.5 41627.5 9847.5 41762.5 ;
      RECT  9972.5 41627.5 10037.5 41762.5 ;
      RECT  10162.5 41627.5 10227.5 41762.5 ;
      RECT  10162.5 41627.5 10227.5 41762.5 ;
      RECT  9972.5 41627.5 10037.5 41762.5 ;
      RECT  10332.5 42557.5 10397.5 42692.5 ;
      RECT  10332.5 41582.5 10397.5 41717.5 ;
      RECT  10167.5 41857.5 10032.5 41922.5 ;
      RECT  9910.0 42072.5 9775.0 42137.5 ;
      RECT  9972.5 42467.5 10037.5 42602.5 ;
      RECT  10162.5 41627.5 10227.5 41762.5 ;
      RECT  10262.5 42072.5 10127.5 42137.5 ;
      RECT  9775.0 42072.5 9910.0 42137.5 ;
      RECT  10032.5 41857.5 10167.5 41922.5 ;
      RECT  10127.5 42072.5 10262.5 42137.5 ;
      RECT  9715.0 42777.5 10635.0 42842.5 ;
      RECT  9715.0 41432.5 10635.0 41497.5 ;
      RECT  11062.5 42625.0 11127.5 42810.0 ;
      RECT  11062.5 41465.0 11127.5 41650.0 ;
      RECT  10702.5 41582.5 10767.5 41432.5 ;
      RECT  10702.5 42467.5 10767.5 42842.5 ;
      RECT  10892.5 41582.5 10957.5 42467.5 ;
      RECT  10702.5 42467.5 10767.5 42602.5 ;
      RECT  10892.5 42467.5 10957.5 42602.5 ;
      RECT  10892.5 42467.5 10957.5 42602.5 ;
      RECT  10702.5 42467.5 10767.5 42602.5 ;
      RECT  10702.5 41582.5 10767.5 41717.5 ;
      RECT  10892.5 41582.5 10957.5 41717.5 ;
      RECT  10892.5 41582.5 10957.5 41717.5 ;
      RECT  10702.5 41582.5 10767.5 41717.5 ;
      RECT  11062.5 42557.5 11127.5 42692.5 ;
      RECT  11062.5 41582.5 11127.5 41717.5 ;
      RECT  10760.0 42025.0 10825.0 42160.0 ;
      RECT  10760.0 42025.0 10825.0 42160.0 ;
      RECT  10925.0 42060.0 10990.0 42125.0 ;
      RECT  10635.0 42777.5 11195.0 42842.5 ;
      RECT  10635.0 41432.5 11195.0 41497.5 ;
      RECT  8897.5 42025.0 8962.5 42160.0 ;
      RECT  9037.5 41752.5 9102.5 41887.5 ;
      RECT  10032.5 41857.5 9897.5 41922.5 ;
      RECT  9582.5 42995.0 9647.5 42810.0 ;
      RECT  9582.5 44155.0 9647.5 43970.0 ;
      RECT  9222.5 44037.5 9287.5 44187.5 ;
      RECT  9222.5 43152.5 9287.5 42777.5 ;
      RECT  9412.5 44037.5 9477.5 43152.5 ;
      RECT  9222.5 43152.5 9287.5 43017.5 ;
      RECT  9412.5 43152.5 9477.5 43017.5 ;
      RECT  9412.5 43152.5 9477.5 43017.5 ;
      RECT  9222.5 43152.5 9287.5 43017.5 ;
      RECT  9222.5 44037.5 9287.5 43902.5 ;
      RECT  9412.5 44037.5 9477.5 43902.5 ;
      RECT  9412.5 44037.5 9477.5 43902.5 ;
      RECT  9222.5 44037.5 9287.5 43902.5 ;
      RECT  9582.5 43062.5 9647.5 42927.5 ;
      RECT  9582.5 44037.5 9647.5 43902.5 ;
      RECT  9280.0 43595.0 9345.0 43460.0 ;
      RECT  9280.0 43595.0 9345.0 43460.0 ;
      RECT  9445.0 43560.0 9510.0 43495.0 ;
      RECT  9155.0 42842.5 9715.0 42777.5 ;
      RECT  9155.0 44187.5 9715.0 44122.5 ;
      RECT  9782.5 43992.5 9847.5 44187.5 ;
      RECT  9782.5 43152.5 9847.5 42777.5 ;
      RECT  10162.5 43152.5 10227.5 42777.5 ;
      RECT  10332.5 42995.0 10397.5 42810.0 ;
      RECT  10332.5 44155.0 10397.5 43970.0 ;
      RECT  9782.5 43152.5 9847.5 43017.5 ;
      RECT  9972.5 43152.5 10037.5 43017.5 ;
      RECT  9972.5 43152.5 10037.5 43017.5 ;
      RECT  9782.5 43152.5 9847.5 43017.5 ;
      RECT  9972.5 43152.5 10037.5 43017.5 ;
      RECT  10162.5 43152.5 10227.5 43017.5 ;
      RECT  10162.5 43152.5 10227.5 43017.5 ;
      RECT  9972.5 43152.5 10037.5 43017.5 ;
      RECT  9782.5 43992.5 9847.5 43857.5 ;
      RECT  9972.5 43992.5 10037.5 43857.5 ;
      RECT  9972.5 43992.5 10037.5 43857.5 ;
      RECT  9782.5 43992.5 9847.5 43857.5 ;
      RECT  9972.5 43992.5 10037.5 43857.5 ;
      RECT  10162.5 43992.5 10227.5 43857.5 ;
      RECT  10162.5 43992.5 10227.5 43857.5 ;
      RECT  9972.5 43992.5 10037.5 43857.5 ;
      RECT  10332.5 43062.5 10397.5 42927.5 ;
      RECT  10332.5 44037.5 10397.5 43902.5 ;
      RECT  10167.5 43762.5 10032.5 43697.5 ;
      RECT  9910.0 43547.5 9775.0 43482.5 ;
      RECT  9972.5 43152.5 10037.5 43017.5 ;
      RECT  10162.5 43992.5 10227.5 43857.5 ;
      RECT  10262.5 43547.5 10127.5 43482.5 ;
      RECT  9775.0 43547.5 9910.0 43482.5 ;
      RECT  10032.5 43762.5 10167.5 43697.5 ;
      RECT  10127.5 43547.5 10262.5 43482.5 ;
      RECT  9715.0 42842.5 10635.0 42777.5 ;
      RECT  9715.0 44187.5 10635.0 44122.5 ;
      RECT  11062.5 42995.0 11127.5 42810.0 ;
      RECT  11062.5 44155.0 11127.5 43970.0 ;
      RECT  10702.5 44037.5 10767.5 44187.5 ;
      RECT  10702.5 43152.5 10767.5 42777.5 ;
      RECT  10892.5 44037.5 10957.5 43152.5 ;
      RECT  10702.5 43152.5 10767.5 43017.5 ;
      RECT  10892.5 43152.5 10957.5 43017.5 ;
      RECT  10892.5 43152.5 10957.5 43017.5 ;
      RECT  10702.5 43152.5 10767.5 43017.5 ;
      RECT  10702.5 44037.5 10767.5 43902.5 ;
      RECT  10892.5 44037.5 10957.5 43902.5 ;
      RECT  10892.5 44037.5 10957.5 43902.5 ;
      RECT  10702.5 44037.5 10767.5 43902.5 ;
      RECT  11062.5 43062.5 11127.5 42927.5 ;
      RECT  11062.5 44037.5 11127.5 43902.5 ;
      RECT  10760.0 43595.0 10825.0 43460.0 ;
      RECT  10760.0 43595.0 10825.0 43460.0 ;
      RECT  10925.0 43560.0 10990.0 43495.0 ;
      RECT  10635.0 42842.5 11195.0 42777.5 ;
      RECT  10635.0 44187.5 11195.0 44122.5 ;
      RECT  8897.5 43460.0 8962.5 43595.0 ;
      RECT  9037.5 43732.5 9102.5 43867.5 ;
      RECT  10032.5 43697.5 9897.5 43762.5 ;
      RECT  9582.5 45315.0 9647.5 45500.0 ;
      RECT  9582.5 44155.0 9647.5 44340.0 ;
      RECT  9222.5 44272.5 9287.5 44122.5 ;
      RECT  9222.5 45157.5 9287.5 45532.5 ;
      RECT  9412.5 44272.5 9477.5 45157.5 ;
      RECT  9222.5 45157.5 9287.5 45292.5 ;
      RECT  9412.5 45157.5 9477.5 45292.5 ;
      RECT  9412.5 45157.5 9477.5 45292.5 ;
      RECT  9222.5 45157.5 9287.5 45292.5 ;
      RECT  9222.5 44272.5 9287.5 44407.5 ;
      RECT  9412.5 44272.5 9477.5 44407.5 ;
      RECT  9412.5 44272.5 9477.5 44407.5 ;
      RECT  9222.5 44272.5 9287.5 44407.5 ;
      RECT  9582.5 45247.5 9647.5 45382.5 ;
      RECT  9582.5 44272.5 9647.5 44407.5 ;
      RECT  9280.0 44715.0 9345.0 44850.0 ;
      RECT  9280.0 44715.0 9345.0 44850.0 ;
      RECT  9445.0 44750.0 9510.0 44815.0 ;
      RECT  9155.0 45467.5 9715.0 45532.5 ;
      RECT  9155.0 44122.5 9715.0 44187.5 ;
      RECT  9782.5 44317.5 9847.5 44122.5 ;
      RECT  9782.5 45157.5 9847.5 45532.5 ;
      RECT  10162.5 45157.5 10227.5 45532.5 ;
      RECT  10332.5 45315.0 10397.5 45500.0 ;
      RECT  10332.5 44155.0 10397.5 44340.0 ;
      RECT  9782.5 45157.5 9847.5 45292.5 ;
      RECT  9972.5 45157.5 10037.5 45292.5 ;
      RECT  9972.5 45157.5 10037.5 45292.5 ;
      RECT  9782.5 45157.5 9847.5 45292.5 ;
      RECT  9972.5 45157.5 10037.5 45292.5 ;
      RECT  10162.5 45157.5 10227.5 45292.5 ;
      RECT  10162.5 45157.5 10227.5 45292.5 ;
      RECT  9972.5 45157.5 10037.5 45292.5 ;
      RECT  9782.5 44317.5 9847.5 44452.5 ;
      RECT  9972.5 44317.5 10037.5 44452.5 ;
      RECT  9972.5 44317.5 10037.5 44452.5 ;
      RECT  9782.5 44317.5 9847.5 44452.5 ;
      RECT  9972.5 44317.5 10037.5 44452.5 ;
      RECT  10162.5 44317.5 10227.5 44452.5 ;
      RECT  10162.5 44317.5 10227.5 44452.5 ;
      RECT  9972.5 44317.5 10037.5 44452.5 ;
      RECT  10332.5 45247.5 10397.5 45382.5 ;
      RECT  10332.5 44272.5 10397.5 44407.5 ;
      RECT  10167.5 44547.5 10032.5 44612.5 ;
      RECT  9910.0 44762.5 9775.0 44827.5 ;
      RECT  9972.5 45157.5 10037.5 45292.5 ;
      RECT  10162.5 44317.5 10227.5 44452.5 ;
      RECT  10262.5 44762.5 10127.5 44827.5 ;
      RECT  9775.0 44762.5 9910.0 44827.5 ;
      RECT  10032.5 44547.5 10167.5 44612.5 ;
      RECT  10127.5 44762.5 10262.5 44827.5 ;
      RECT  9715.0 45467.5 10635.0 45532.5 ;
      RECT  9715.0 44122.5 10635.0 44187.5 ;
      RECT  11062.5 45315.0 11127.5 45500.0 ;
      RECT  11062.5 44155.0 11127.5 44340.0 ;
      RECT  10702.5 44272.5 10767.5 44122.5 ;
      RECT  10702.5 45157.5 10767.5 45532.5 ;
      RECT  10892.5 44272.5 10957.5 45157.5 ;
      RECT  10702.5 45157.5 10767.5 45292.5 ;
      RECT  10892.5 45157.5 10957.5 45292.5 ;
      RECT  10892.5 45157.5 10957.5 45292.5 ;
      RECT  10702.5 45157.5 10767.5 45292.5 ;
      RECT  10702.5 44272.5 10767.5 44407.5 ;
      RECT  10892.5 44272.5 10957.5 44407.5 ;
      RECT  10892.5 44272.5 10957.5 44407.5 ;
      RECT  10702.5 44272.5 10767.5 44407.5 ;
      RECT  11062.5 45247.5 11127.5 45382.5 ;
      RECT  11062.5 44272.5 11127.5 44407.5 ;
      RECT  10760.0 44715.0 10825.0 44850.0 ;
      RECT  10760.0 44715.0 10825.0 44850.0 ;
      RECT  10925.0 44750.0 10990.0 44815.0 ;
      RECT  10635.0 45467.5 11195.0 45532.5 ;
      RECT  10635.0 44122.5 11195.0 44187.5 ;
      RECT  8897.5 44715.0 8962.5 44850.0 ;
      RECT  9037.5 44442.5 9102.5 44577.5 ;
      RECT  10032.5 44547.5 9897.5 44612.5 ;
      RECT  9582.5 45685.0 9647.5 45500.0 ;
      RECT  9582.5 46845.0 9647.5 46660.0 ;
      RECT  9222.5 46727.5 9287.5 46877.5 ;
      RECT  9222.5 45842.5 9287.5 45467.5 ;
      RECT  9412.5 46727.5 9477.5 45842.5 ;
      RECT  9222.5 45842.5 9287.5 45707.5 ;
      RECT  9412.5 45842.5 9477.5 45707.5 ;
      RECT  9412.5 45842.5 9477.5 45707.5 ;
      RECT  9222.5 45842.5 9287.5 45707.5 ;
      RECT  9222.5 46727.5 9287.5 46592.5 ;
      RECT  9412.5 46727.5 9477.5 46592.5 ;
      RECT  9412.5 46727.5 9477.5 46592.5 ;
      RECT  9222.5 46727.5 9287.5 46592.5 ;
      RECT  9582.5 45752.5 9647.5 45617.5 ;
      RECT  9582.5 46727.5 9647.5 46592.5 ;
      RECT  9280.0 46285.0 9345.0 46150.0 ;
      RECT  9280.0 46285.0 9345.0 46150.0 ;
      RECT  9445.0 46250.0 9510.0 46185.0 ;
      RECT  9155.0 45532.5 9715.0 45467.5 ;
      RECT  9155.0 46877.5 9715.0 46812.5 ;
      RECT  9782.5 46682.5 9847.5 46877.5 ;
      RECT  9782.5 45842.5 9847.5 45467.5 ;
      RECT  10162.5 45842.5 10227.5 45467.5 ;
      RECT  10332.5 45685.0 10397.5 45500.0 ;
      RECT  10332.5 46845.0 10397.5 46660.0 ;
      RECT  9782.5 45842.5 9847.5 45707.5 ;
      RECT  9972.5 45842.5 10037.5 45707.5 ;
      RECT  9972.5 45842.5 10037.5 45707.5 ;
      RECT  9782.5 45842.5 9847.5 45707.5 ;
      RECT  9972.5 45842.5 10037.5 45707.5 ;
      RECT  10162.5 45842.5 10227.5 45707.5 ;
      RECT  10162.5 45842.5 10227.5 45707.5 ;
      RECT  9972.5 45842.5 10037.5 45707.5 ;
      RECT  9782.5 46682.5 9847.5 46547.5 ;
      RECT  9972.5 46682.5 10037.5 46547.5 ;
      RECT  9972.5 46682.5 10037.5 46547.5 ;
      RECT  9782.5 46682.5 9847.5 46547.5 ;
      RECT  9972.5 46682.5 10037.5 46547.5 ;
      RECT  10162.5 46682.5 10227.5 46547.5 ;
      RECT  10162.5 46682.5 10227.5 46547.5 ;
      RECT  9972.5 46682.5 10037.5 46547.5 ;
      RECT  10332.5 45752.5 10397.5 45617.5 ;
      RECT  10332.5 46727.5 10397.5 46592.5 ;
      RECT  10167.5 46452.5 10032.5 46387.5 ;
      RECT  9910.0 46237.5 9775.0 46172.5 ;
      RECT  9972.5 45842.5 10037.5 45707.5 ;
      RECT  10162.5 46682.5 10227.5 46547.5 ;
      RECT  10262.5 46237.5 10127.5 46172.5 ;
      RECT  9775.0 46237.5 9910.0 46172.5 ;
      RECT  10032.5 46452.5 10167.5 46387.5 ;
      RECT  10127.5 46237.5 10262.5 46172.5 ;
      RECT  9715.0 45532.5 10635.0 45467.5 ;
      RECT  9715.0 46877.5 10635.0 46812.5 ;
      RECT  11062.5 45685.0 11127.5 45500.0 ;
      RECT  11062.5 46845.0 11127.5 46660.0 ;
      RECT  10702.5 46727.5 10767.5 46877.5 ;
      RECT  10702.5 45842.5 10767.5 45467.5 ;
      RECT  10892.5 46727.5 10957.5 45842.5 ;
      RECT  10702.5 45842.5 10767.5 45707.5 ;
      RECT  10892.5 45842.5 10957.5 45707.5 ;
      RECT  10892.5 45842.5 10957.5 45707.5 ;
      RECT  10702.5 45842.5 10767.5 45707.5 ;
      RECT  10702.5 46727.5 10767.5 46592.5 ;
      RECT  10892.5 46727.5 10957.5 46592.5 ;
      RECT  10892.5 46727.5 10957.5 46592.5 ;
      RECT  10702.5 46727.5 10767.5 46592.5 ;
      RECT  11062.5 45752.5 11127.5 45617.5 ;
      RECT  11062.5 46727.5 11127.5 46592.5 ;
      RECT  10760.0 46285.0 10825.0 46150.0 ;
      RECT  10760.0 46285.0 10825.0 46150.0 ;
      RECT  10925.0 46250.0 10990.0 46185.0 ;
      RECT  10635.0 45532.5 11195.0 45467.5 ;
      RECT  10635.0 46877.5 11195.0 46812.5 ;
      RECT  8897.5 46150.0 8962.5 46285.0 ;
      RECT  9037.5 46422.5 9102.5 46557.5 ;
      RECT  10032.5 46387.5 9897.5 46452.5 ;
      RECT  9582.5 48005.0 9647.5 48190.0 ;
      RECT  9582.5 46845.0 9647.5 47030.0 ;
      RECT  9222.5 46962.5 9287.5 46812.5 ;
      RECT  9222.5 47847.5 9287.5 48222.5 ;
      RECT  9412.5 46962.5 9477.5 47847.5 ;
      RECT  9222.5 47847.5 9287.5 47982.5 ;
      RECT  9412.5 47847.5 9477.5 47982.5 ;
      RECT  9412.5 47847.5 9477.5 47982.5 ;
      RECT  9222.5 47847.5 9287.5 47982.5 ;
      RECT  9222.5 46962.5 9287.5 47097.5 ;
      RECT  9412.5 46962.5 9477.5 47097.5 ;
      RECT  9412.5 46962.5 9477.5 47097.5 ;
      RECT  9222.5 46962.5 9287.5 47097.5 ;
      RECT  9582.5 47937.5 9647.5 48072.5 ;
      RECT  9582.5 46962.5 9647.5 47097.5 ;
      RECT  9280.0 47405.0 9345.0 47540.0 ;
      RECT  9280.0 47405.0 9345.0 47540.0 ;
      RECT  9445.0 47440.0 9510.0 47505.0 ;
      RECT  9155.0 48157.5 9715.0 48222.5 ;
      RECT  9155.0 46812.5 9715.0 46877.5 ;
      RECT  9782.5 47007.5 9847.5 46812.5 ;
      RECT  9782.5 47847.5 9847.5 48222.5 ;
      RECT  10162.5 47847.5 10227.5 48222.5 ;
      RECT  10332.5 48005.0 10397.5 48190.0 ;
      RECT  10332.5 46845.0 10397.5 47030.0 ;
      RECT  9782.5 47847.5 9847.5 47982.5 ;
      RECT  9972.5 47847.5 10037.5 47982.5 ;
      RECT  9972.5 47847.5 10037.5 47982.5 ;
      RECT  9782.5 47847.5 9847.5 47982.5 ;
      RECT  9972.5 47847.5 10037.5 47982.5 ;
      RECT  10162.5 47847.5 10227.5 47982.5 ;
      RECT  10162.5 47847.5 10227.5 47982.5 ;
      RECT  9972.5 47847.5 10037.5 47982.5 ;
      RECT  9782.5 47007.5 9847.5 47142.5 ;
      RECT  9972.5 47007.5 10037.5 47142.5 ;
      RECT  9972.5 47007.5 10037.5 47142.5 ;
      RECT  9782.5 47007.5 9847.5 47142.5 ;
      RECT  9972.5 47007.5 10037.5 47142.5 ;
      RECT  10162.5 47007.5 10227.5 47142.5 ;
      RECT  10162.5 47007.5 10227.5 47142.5 ;
      RECT  9972.5 47007.5 10037.5 47142.5 ;
      RECT  10332.5 47937.5 10397.5 48072.5 ;
      RECT  10332.5 46962.5 10397.5 47097.5 ;
      RECT  10167.5 47237.5 10032.5 47302.5 ;
      RECT  9910.0 47452.5 9775.0 47517.5 ;
      RECT  9972.5 47847.5 10037.5 47982.5 ;
      RECT  10162.5 47007.5 10227.5 47142.5 ;
      RECT  10262.5 47452.5 10127.5 47517.5 ;
      RECT  9775.0 47452.5 9910.0 47517.5 ;
      RECT  10032.5 47237.5 10167.5 47302.5 ;
      RECT  10127.5 47452.5 10262.5 47517.5 ;
      RECT  9715.0 48157.5 10635.0 48222.5 ;
      RECT  9715.0 46812.5 10635.0 46877.5 ;
      RECT  11062.5 48005.0 11127.5 48190.0 ;
      RECT  11062.5 46845.0 11127.5 47030.0 ;
      RECT  10702.5 46962.5 10767.5 46812.5 ;
      RECT  10702.5 47847.5 10767.5 48222.5 ;
      RECT  10892.5 46962.5 10957.5 47847.5 ;
      RECT  10702.5 47847.5 10767.5 47982.5 ;
      RECT  10892.5 47847.5 10957.5 47982.5 ;
      RECT  10892.5 47847.5 10957.5 47982.5 ;
      RECT  10702.5 47847.5 10767.5 47982.5 ;
      RECT  10702.5 46962.5 10767.5 47097.5 ;
      RECT  10892.5 46962.5 10957.5 47097.5 ;
      RECT  10892.5 46962.5 10957.5 47097.5 ;
      RECT  10702.5 46962.5 10767.5 47097.5 ;
      RECT  11062.5 47937.5 11127.5 48072.5 ;
      RECT  11062.5 46962.5 11127.5 47097.5 ;
      RECT  10760.0 47405.0 10825.0 47540.0 ;
      RECT  10760.0 47405.0 10825.0 47540.0 ;
      RECT  10925.0 47440.0 10990.0 47505.0 ;
      RECT  10635.0 48157.5 11195.0 48222.5 ;
      RECT  10635.0 46812.5 11195.0 46877.5 ;
      RECT  8897.5 47405.0 8962.5 47540.0 ;
      RECT  9037.5 47132.5 9102.5 47267.5 ;
      RECT  10032.5 47237.5 9897.5 47302.5 ;
      RECT  9582.5 48375.0 9647.5 48190.0 ;
      RECT  9582.5 49535.0 9647.5 49350.0 ;
      RECT  9222.5 49417.5 9287.5 49567.5 ;
      RECT  9222.5 48532.5 9287.5 48157.5 ;
      RECT  9412.5 49417.5 9477.5 48532.5 ;
      RECT  9222.5 48532.5 9287.5 48397.5 ;
      RECT  9412.5 48532.5 9477.5 48397.5 ;
      RECT  9412.5 48532.5 9477.5 48397.5 ;
      RECT  9222.5 48532.5 9287.5 48397.5 ;
      RECT  9222.5 49417.5 9287.5 49282.5 ;
      RECT  9412.5 49417.5 9477.5 49282.5 ;
      RECT  9412.5 49417.5 9477.5 49282.5 ;
      RECT  9222.5 49417.5 9287.5 49282.5 ;
      RECT  9582.5 48442.5 9647.5 48307.5 ;
      RECT  9582.5 49417.5 9647.5 49282.5 ;
      RECT  9280.0 48975.0 9345.0 48840.0 ;
      RECT  9280.0 48975.0 9345.0 48840.0 ;
      RECT  9445.0 48940.0 9510.0 48875.0 ;
      RECT  9155.0 48222.5 9715.0 48157.5 ;
      RECT  9155.0 49567.5 9715.0 49502.5 ;
      RECT  9782.5 49372.5 9847.5 49567.5 ;
      RECT  9782.5 48532.5 9847.5 48157.5 ;
      RECT  10162.5 48532.5 10227.5 48157.5 ;
      RECT  10332.5 48375.0 10397.5 48190.0 ;
      RECT  10332.5 49535.0 10397.5 49350.0 ;
      RECT  9782.5 48532.5 9847.5 48397.5 ;
      RECT  9972.5 48532.5 10037.5 48397.5 ;
      RECT  9972.5 48532.5 10037.5 48397.5 ;
      RECT  9782.5 48532.5 9847.5 48397.5 ;
      RECT  9972.5 48532.5 10037.5 48397.5 ;
      RECT  10162.5 48532.5 10227.5 48397.5 ;
      RECT  10162.5 48532.5 10227.5 48397.5 ;
      RECT  9972.5 48532.5 10037.5 48397.5 ;
      RECT  9782.5 49372.5 9847.5 49237.5 ;
      RECT  9972.5 49372.5 10037.5 49237.5 ;
      RECT  9972.5 49372.5 10037.5 49237.5 ;
      RECT  9782.5 49372.5 9847.5 49237.5 ;
      RECT  9972.5 49372.5 10037.5 49237.5 ;
      RECT  10162.5 49372.5 10227.5 49237.5 ;
      RECT  10162.5 49372.5 10227.5 49237.5 ;
      RECT  9972.5 49372.5 10037.5 49237.5 ;
      RECT  10332.5 48442.5 10397.5 48307.5 ;
      RECT  10332.5 49417.5 10397.5 49282.5 ;
      RECT  10167.5 49142.5 10032.5 49077.5 ;
      RECT  9910.0 48927.5 9775.0 48862.5 ;
      RECT  9972.5 48532.5 10037.5 48397.5 ;
      RECT  10162.5 49372.5 10227.5 49237.5 ;
      RECT  10262.5 48927.5 10127.5 48862.5 ;
      RECT  9775.0 48927.5 9910.0 48862.5 ;
      RECT  10032.5 49142.5 10167.5 49077.5 ;
      RECT  10127.5 48927.5 10262.5 48862.5 ;
      RECT  9715.0 48222.5 10635.0 48157.5 ;
      RECT  9715.0 49567.5 10635.0 49502.5 ;
      RECT  11062.5 48375.0 11127.5 48190.0 ;
      RECT  11062.5 49535.0 11127.5 49350.0 ;
      RECT  10702.5 49417.5 10767.5 49567.5 ;
      RECT  10702.5 48532.5 10767.5 48157.5 ;
      RECT  10892.5 49417.5 10957.5 48532.5 ;
      RECT  10702.5 48532.5 10767.5 48397.5 ;
      RECT  10892.5 48532.5 10957.5 48397.5 ;
      RECT  10892.5 48532.5 10957.5 48397.5 ;
      RECT  10702.5 48532.5 10767.5 48397.5 ;
      RECT  10702.5 49417.5 10767.5 49282.5 ;
      RECT  10892.5 49417.5 10957.5 49282.5 ;
      RECT  10892.5 49417.5 10957.5 49282.5 ;
      RECT  10702.5 49417.5 10767.5 49282.5 ;
      RECT  11062.5 48442.5 11127.5 48307.5 ;
      RECT  11062.5 49417.5 11127.5 49282.5 ;
      RECT  10760.0 48975.0 10825.0 48840.0 ;
      RECT  10760.0 48975.0 10825.0 48840.0 ;
      RECT  10925.0 48940.0 10990.0 48875.0 ;
      RECT  10635.0 48222.5 11195.0 48157.5 ;
      RECT  10635.0 49567.5 11195.0 49502.5 ;
      RECT  8897.5 48840.0 8962.5 48975.0 ;
      RECT  9037.5 49112.5 9102.5 49247.5 ;
      RECT  10032.5 49077.5 9897.5 49142.5 ;
      RECT  9582.5 50695.0 9647.5 50880.0 ;
      RECT  9582.5 49535.0 9647.5 49720.0 ;
      RECT  9222.5 49652.5 9287.5 49502.5 ;
      RECT  9222.5 50537.5 9287.5 50912.5 ;
      RECT  9412.5 49652.5 9477.5 50537.5 ;
      RECT  9222.5 50537.5 9287.5 50672.5 ;
      RECT  9412.5 50537.5 9477.5 50672.5 ;
      RECT  9412.5 50537.5 9477.5 50672.5 ;
      RECT  9222.5 50537.5 9287.5 50672.5 ;
      RECT  9222.5 49652.5 9287.5 49787.5 ;
      RECT  9412.5 49652.5 9477.5 49787.5 ;
      RECT  9412.5 49652.5 9477.5 49787.5 ;
      RECT  9222.5 49652.5 9287.5 49787.5 ;
      RECT  9582.5 50627.5 9647.5 50762.5 ;
      RECT  9582.5 49652.5 9647.5 49787.5 ;
      RECT  9280.0 50095.0 9345.0 50230.0 ;
      RECT  9280.0 50095.0 9345.0 50230.0 ;
      RECT  9445.0 50130.0 9510.0 50195.0 ;
      RECT  9155.0 50847.5 9715.0 50912.5 ;
      RECT  9155.0 49502.5 9715.0 49567.5 ;
      RECT  9782.5 49697.5 9847.5 49502.5 ;
      RECT  9782.5 50537.5 9847.5 50912.5 ;
      RECT  10162.5 50537.5 10227.5 50912.5 ;
      RECT  10332.5 50695.0 10397.5 50880.0 ;
      RECT  10332.5 49535.0 10397.5 49720.0 ;
      RECT  9782.5 50537.5 9847.5 50672.5 ;
      RECT  9972.5 50537.5 10037.5 50672.5 ;
      RECT  9972.5 50537.5 10037.5 50672.5 ;
      RECT  9782.5 50537.5 9847.5 50672.5 ;
      RECT  9972.5 50537.5 10037.5 50672.5 ;
      RECT  10162.5 50537.5 10227.5 50672.5 ;
      RECT  10162.5 50537.5 10227.5 50672.5 ;
      RECT  9972.5 50537.5 10037.5 50672.5 ;
      RECT  9782.5 49697.5 9847.5 49832.5 ;
      RECT  9972.5 49697.5 10037.5 49832.5 ;
      RECT  9972.5 49697.5 10037.5 49832.5 ;
      RECT  9782.5 49697.5 9847.5 49832.5 ;
      RECT  9972.5 49697.5 10037.5 49832.5 ;
      RECT  10162.5 49697.5 10227.5 49832.5 ;
      RECT  10162.5 49697.5 10227.5 49832.5 ;
      RECT  9972.5 49697.5 10037.5 49832.5 ;
      RECT  10332.5 50627.5 10397.5 50762.5 ;
      RECT  10332.5 49652.5 10397.5 49787.5 ;
      RECT  10167.5 49927.5 10032.5 49992.5 ;
      RECT  9910.0 50142.5 9775.0 50207.5 ;
      RECT  9972.5 50537.5 10037.5 50672.5 ;
      RECT  10162.5 49697.5 10227.5 49832.5 ;
      RECT  10262.5 50142.5 10127.5 50207.5 ;
      RECT  9775.0 50142.5 9910.0 50207.5 ;
      RECT  10032.5 49927.5 10167.5 49992.5 ;
      RECT  10127.5 50142.5 10262.5 50207.5 ;
      RECT  9715.0 50847.5 10635.0 50912.5 ;
      RECT  9715.0 49502.5 10635.0 49567.5 ;
      RECT  11062.5 50695.0 11127.5 50880.0 ;
      RECT  11062.5 49535.0 11127.5 49720.0 ;
      RECT  10702.5 49652.5 10767.5 49502.5 ;
      RECT  10702.5 50537.5 10767.5 50912.5 ;
      RECT  10892.5 49652.5 10957.5 50537.5 ;
      RECT  10702.5 50537.5 10767.5 50672.5 ;
      RECT  10892.5 50537.5 10957.5 50672.5 ;
      RECT  10892.5 50537.5 10957.5 50672.5 ;
      RECT  10702.5 50537.5 10767.5 50672.5 ;
      RECT  10702.5 49652.5 10767.5 49787.5 ;
      RECT  10892.5 49652.5 10957.5 49787.5 ;
      RECT  10892.5 49652.5 10957.5 49787.5 ;
      RECT  10702.5 49652.5 10767.5 49787.5 ;
      RECT  11062.5 50627.5 11127.5 50762.5 ;
      RECT  11062.5 49652.5 11127.5 49787.5 ;
      RECT  10760.0 50095.0 10825.0 50230.0 ;
      RECT  10760.0 50095.0 10825.0 50230.0 ;
      RECT  10925.0 50130.0 10990.0 50195.0 ;
      RECT  10635.0 50847.5 11195.0 50912.5 ;
      RECT  10635.0 49502.5 11195.0 49567.5 ;
      RECT  8897.5 50095.0 8962.5 50230.0 ;
      RECT  9037.5 49822.5 9102.5 49957.5 ;
      RECT  10032.5 49927.5 9897.5 49992.5 ;
      RECT  9582.5 51065.0 9647.5 50880.0 ;
      RECT  9582.5 52225.0 9647.5 52040.0 ;
      RECT  9222.5 52107.5 9287.5 52257.5 ;
      RECT  9222.5 51222.5 9287.5 50847.5 ;
      RECT  9412.5 52107.5 9477.5 51222.5 ;
      RECT  9222.5 51222.5 9287.5 51087.5 ;
      RECT  9412.5 51222.5 9477.5 51087.5 ;
      RECT  9412.5 51222.5 9477.5 51087.5 ;
      RECT  9222.5 51222.5 9287.5 51087.5 ;
      RECT  9222.5 52107.5 9287.5 51972.5 ;
      RECT  9412.5 52107.5 9477.5 51972.5 ;
      RECT  9412.5 52107.5 9477.5 51972.5 ;
      RECT  9222.5 52107.5 9287.5 51972.5 ;
      RECT  9582.5 51132.5 9647.5 50997.5 ;
      RECT  9582.5 52107.5 9647.5 51972.5 ;
      RECT  9280.0 51665.0 9345.0 51530.0 ;
      RECT  9280.0 51665.0 9345.0 51530.0 ;
      RECT  9445.0 51630.0 9510.0 51565.0 ;
      RECT  9155.0 50912.5 9715.0 50847.5 ;
      RECT  9155.0 52257.5 9715.0 52192.5 ;
      RECT  9782.5 52062.5 9847.5 52257.5 ;
      RECT  9782.5 51222.5 9847.5 50847.5 ;
      RECT  10162.5 51222.5 10227.5 50847.5 ;
      RECT  10332.5 51065.0 10397.5 50880.0 ;
      RECT  10332.5 52225.0 10397.5 52040.0 ;
      RECT  9782.5 51222.5 9847.5 51087.5 ;
      RECT  9972.5 51222.5 10037.5 51087.5 ;
      RECT  9972.5 51222.5 10037.5 51087.5 ;
      RECT  9782.5 51222.5 9847.5 51087.5 ;
      RECT  9972.5 51222.5 10037.5 51087.5 ;
      RECT  10162.5 51222.5 10227.5 51087.5 ;
      RECT  10162.5 51222.5 10227.5 51087.5 ;
      RECT  9972.5 51222.5 10037.5 51087.5 ;
      RECT  9782.5 52062.5 9847.5 51927.5 ;
      RECT  9972.5 52062.5 10037.5 51927.5 ;
      RECT  9972.5 52062.5 10037.5 51927.5 ;
      RECT  9782.5 52062.5 9847.5 51927.5 ;
      RECT  9972.5 52062.5 10037.5 51927.5 ;
      RECT  10162.5 52062.5 10227.5 51927.5 ;
      RECT  10162.5 52062.5 10227.5 51927.5 ;
      RECT  9972.5 52062.5 10037.5 51927.5 ;
      RECT  10332.5 51132.5 10397.5 50997.5 ;
      RECT  10332.5 52107.5 10397.5 51972.5 ;
      RECT  10167.5 51832.5 10032.5 51767.5 ;
      RECT  9910.0 51617.5 9775.0 51552.5 ;
      RECT  9972.5 51222.5 10037.5 51087.5 ;
      RECT  10162.5 52062.5 10227.5 51927.5 ;
      RECT  10262.5 51617.5 10127.5 51552.5 ;
      RECT  9775.0 51617.5 9910.0 51552.5 ;
      RECT  10032.5 51832.5 10167.5 51767.5 ;
      RECT  10127.5 51617.5 10262.5 51552.5 ;
      RECT  9715.0 50912.5 10635.0 50847.5 ;
      RECT  9715.0 52257.5 10635.0 52192.5 ;
      RECT  11062.5 51065.0 11127.5 50880.0 ;
      RECT  11062.5 52225.0 11127.5 52040.0 ;
      RECT  10702.5 52107.5 10767.5 52257.5 ;
      RECT  10702.5 51222.5 10767.5 50847.5 ;
      RECT  10892.5 52107.5 10957.5 51222.5 ;
      RECT  10702.5 51222.5 10767.5 51087.5 ;
      RECT  10892.5 51222.5 10957.5 51087.5 ;
      RECT  10892.5 51222.5 10957.5 51087.5 ;
      RECT  10702.5 51222.5 10767.5 51087.5 ;
      RECT  10702.5 52107.5 10767.5 51972.5 ;
      RECT  10892.5 52107.5 10957.5 51972.5 ;
      RECT  10892.5 52107.5 10957.5 51972.5 ;
      RECT  10702.5 52107.5 10767.5 51972.5 ;
      RECT  11062.5 51132.5 11127.5 50997.5 ;
      RECT  11062.5 52107.5 11127.5 51972.5 ;
      RECT  10760.0 51665.0 10825.0 51530.0 ;
      RECT  10760.0 51665.0 10825.0 51530.0 ;
      RECT  10925.0 51630.0 10990.0 51565.0 ;
      RECT  10635.0 50912.5 11195.0 50847.5 ;
      RECT  10635.0 52257.5 11195.0 52192.5 ;
      RECT  8897.5 51530.0 8962.5 51665.0 ;
      RECT  9037.5 51802.5 9102.5 51937.5 ;
      RECT  10032.5 51767.5 9897.5 51832.5 ;
      RECT  9582.5 53385.0 9647.5 53570.0 ;
      RECT  9582.5 52225.0 9647.5 52410.0 ;
      RECT  9222.5 52342.5 9287.5 52192.5 ;
      RECT  9222.5 53227.5 9287.5 53602.5 ;
      RECT  9412.5 52342.5 9477.5 53227.5 ;
      RECT  9222.5 53227.5 9287.5 53362.5 ;
      RECT  9412.5 53227.5 9477.5 53362.5 ;
      RECT  9412.5 53227.5 9477.5 53362.5 ;
      RECT  9222.5 53227.5 9287.5 53362.5 ;
      RECT  9222.5 52342.5 9287.5 52477.5 ;
      RECT  9412.5 52342.5 9477.5 52477.5 ;
      RECT  9412.5 52342.5 9477.5 52477.5 ;
      RECT  9222.5 52342.5 9287.5 52477.5 ;
      RECT  9582.5 53317.5 9647.5 53452.5 ;
      RECT  9582.5 52342.5 9647.5 52477.5 ;
      RECT  9280.0 52785.0 9345.0 52920.0 ;
      RECT  9280.0 52785.0 9345.0 52920.0 ;
      RECT  9445.0 52820.0 9510.0 52885.0 ;
      RECT  9155.0 53537.5 9715.0 53602.5 ;
      RECT  9155.0 52192.5 9715.0 52257.5 ;
      RECT  9782.5 52387.5 9847.5 52192.5 ;
      RECT  9782.5 53227.5 9847.5 53602.5 ;
      RECT  10162.5 53227.5 10227.5 53602.5 ;
      RECT  10332.5 53385.0 10397.5 53570.0 ;
      RECT  10332.5 52225.0 10397.5 52410.0 ;
      RECT  9782.5 53227.5 9847.5 53362.5 ;
      RECT  9972.5 53227.5 10037.5 53362.5 ;
      RECT  9972.5 53227.5 10037.5 53362.5 ;
      RECT  9782.5 53227.5 9847.5 53362.5 ;
      RECT  9972.5 53227.5 10037.5 53362.5 ;
      RECT  10162.5 53227.5 10227.5 53362.5 ;
      RECT  10162.5 53227.5 10227.5 53362.5 ;
      RECT  9972.5 53227.5 10037.5 53362.5 ;
      RECT  9782.5 52387.5 9847.5 52522.5 ;
      RECT  9972.5 52387.5 10037.5 52522.5 ;
      RECT  9972.5 52387.5 10037.5 52522.5 ;
      RECT  9782.5 52387.5 9847.5 52522.5 ;
      RECT  9972.5 52387.5 10037.5 52522.5 ;
      RECT  10162.5 52387.5 10227.5 52522.5 ;
      RECT  10162.5 52387.5 10227.5 52522.5 ;
      RECT  9972.5 52387.5 10037.5 52522.5 ;
      RECT  10332.5 53317.5 10397.5 53452.5 ;
      RECT  10332.5 52342.5 10397.5 52477.5 ;
      RECT  10167.5 52617.5 10032.5 52682.5 ;
      RECT  9910.0 52832.5 9775.0 52897.5 ;
      RECT  9972.5 53227.5 10037.5 53362.5 ;
      RECT  10162.5 52387.5 10227.5 52522.5 ;
      RECT  10262.5 52832.5 10127.5 52897.5 ;
      RECT  9775.0 52832.5 9910.0 52897.5 ;
      RECT  10032.5 52617.5 10167.5 52682.5 ;
      RECT  10127.5 52832.5 10262.5 52897.5 ;
      RECT  9715.0 53537.5 10635.0 53602.5 ;
      RECT  9715.0 52192.5 10635.0 52257.5 ;
      RECT  11062.5 53385.0 11127.5 53570.0 ;
      RECT  11062.5 52225.0 11127.5 52410.0 ;
      RECT  10702.5 52342.5 10767.5 52192.5 ;
      RECT  10702.5 53227.5 10767.5 53602.5 ;
      RECT  10892.5 52342.5 10957.5 53227.5 ;
      RECT  10702.5 53227.5 10767.5 53362.5 ;
      RECT  10892.5 53227.5 10957.5 53362.5 ;
      RECT  10892.5 53227.5 10957.5 53362.5 ;
      RECT  10702.5 53227.5 10767.5 53362.5 ;
      RECT  10702.5 52342.5 10767.5 52477.5 ;
      RECT  10892.5 52342.5 10957.5 52477.5 ;
      RECT  10892.5 52342.5 10957.5 52477.5 ;
      RECT  10702.5 52342.5 10767.5 52477.5 ;
      RECT  11062.5 53317.5 11127.5 53452.5 ;
      RECT  11062.5 52342.5 11127.5 52477.5 ;
      RECT  10760.0 52785.0 10825.0 52920.0 ;
      RECT  10760.0 52785.0 10825.0 52920.0 ;
      RECT  10925.0 52820.0 10990.0 52885.0 ;
      RECT  10635.0 53537.5 11195.0 53602.5 ;
      RECT  10635.0 52192.5 11195.0 52257.5 ;
      RECT  8897.5 52785.0 8962.5 52920.0 ;
      RECT  9037.5 52512.5 9102.5 52647.5 ;
      RECT  10032.5 52617.5 9897.5 52682.5 ;
      RECT  9582.5 53755.0 9647.5 53570.0 ;
      RECT  9582.5 54915.0 9647.5 54730.0 ;
      RECT  9222.5 54797.5 9287.5 54947.5 ;
      RECT  9222.5 53912.5 9287.5 53537.5 ;
      RECT  9412.5 54797.5 9477.5 53912.5 ;
      RECT  9222.5 53912.5 9287.5 53777.5 ;
      RECT  9412.5 53912.5 9477.5 53777.5 ;
      RECT  9412.5 53912.5 9477.5 53777.5 ;
      RECT  9222.5 53912.5 9287.5 53777.5 ;
      RECT  9222.5 54797.5 9287.5 54662.5 ;
      RECT  9412.5 54797.5 9477.5 54662.5 ;
      RECT  9412.5 54797.5 9477.5 54662.5 ;
      RECT  9222.5 54797.5 9287.5 54662.5 ;
      RECT  9582.5 53822.5 9647.5 53687.5 ;
      RECT  9582.5 54797.5 9647.5 54662.5 ;
      RECT  9280.0 54355.0 9345.0 54220.0 ;
      RECT  9280.0 54355.0 9345.0 54220.0 ;
      RECT  9445.0 54320.0 9510.0 54255.0 ;
      RECT  9155.0 53602.5 9715.0 53537.5 ;
      RECT  9155.0 54947.5 9715.0 54882.5 ;
      RECT  9782.5 54752.5 9847.5 54947.5 ;
      RECT  9782.5 53912.5 9847.5 53537.5 ;
      RECT  10162.5 53912.5 10227.5 53537.5 ;
      RECT  10332.5 53755.0 10397.5 53570.0 ;
      RECT  10332.5 54915.0 10397.5 54730.0 ;
      RECT  9782.5 53912.5 9847.5 53777.5 ;
      RECT  9972.5 53912.5 10037.5 53777.5 ;
      RECT  9972.5 53912.5 10037.5 53777.5 ;
      RECT  9782.5 53912.5 9847.5 53777.5 ;
      RECT  9972.5 53912.5 10037.5 53777.5 ;
      RECT  10162.5 53912.5 10227.5 53777.5 ;
      RECT  10162.5 53912.5 10227.5 53777.5 ;
      RECT  9972.5 53912.5 10037.5 53777.5 ;
      RECT  9782.5 54752.5 9847.5 54617.5 ;
      RECT  9972.5 54752.5 10037.5 54617.5 ;
      RECT  9972.5 54752.5 10037.5 54617.5 ;
      RECT  9782.5 54752.5 9847.5 54617.5 ;
      RECT  9972.5 54752.5 10037.5 54617.5 ;
      RECT  10162.5 54752.5 10227.5 54617.5 ;
      RECT  10162.5 54752.5 10227.5 54617.5 ;
      RECT  9972.5 54752.5 10037.5 54617.5 ;
      RECT  10332.5 53822.5 10397.5 53687.5 ;
      RECT  10332.5 54797.5 10397.5 54662.5 ;
      RECT  10167.5 54522.5 10032.5 54457.5 ;
      RECT  9910.0 54307.5 9775.0 54242.5 ;
      RECT  9972.5 53912.5 10037.5 53777.5 ;
      RECT  10162.5 54752.5 10227.5 54617.5 ;
      RECT  10262.5 54307.5 10127.5 54242.5 ;
      RECT  9775.0 54307.5 9910.0 54242.5 ;
      RECT  10032.5 54522.5 10167.5 54457.5 ;
      RECT  10127.5 54307.5 10262.5 54242.5 ;
      RECT  9715.0 53602.5 10635.0 53537.5 ;
      RECT  9715.0 54947.5 10635.0 54882.5 ;
      RECT  11062.5 53755.0 11127.5 53570.0 ;
      RECT  11062.5 54915.0 11127.5 54730.0 ;
      RECT  10702.5 54797.5 10767.5 54947.5 ;
      RECT  10702.5 53912.5 10767.5 53537.5 ;
      RECT  10892.5 54797.5 10957.5 53912.5 ;
      RECT  10702.5 53912.5 10767.5 53777.5 ;
      RECT  10892.5 53912.5 10957.5 53777.5 ;
      RECT  10892.5 53912.5 10957.5 53777.5 ;
      RECT  10702.5 53912.5 10767.5 53777.5 ;
      RECT  10702.5 54797.5 10767.5 54662.5 ;
      RECT  10892.5 54797.5 10957.5 54662.5 ;
      RECT  10892.5 54797.5 10957.5 54662.5 ;
      RECT  10702.5 54797.5 10767.5 54662.5 ;
      RECT  11062.5 53822.5 11127.5 53687.5 ;
      RECT  11062.5 54797.5 11127.5 54662.5 ;
      RECT  10760.0 54355.0 10825.0 54220.0 ;
      RECT  10760.0 54355.0 10825.0 54220.0 ;
      RECT  10925.0 54320.0 10990.0 54255.0 ;
      RECT  10635.0 53602.5 11195.0 53537.5 ;
      RECT  10635.0 54947.5 11195.0 54882.5 ;
      RECT  8897.5 54220.0 8962.5 54355.0 ;
      RECT  9037.5 54492.5 9102.5 54627.5 ;
      RECT  10032.5 54457.5 9897.5 54522.5 ;
      RECT  9582.5 56075.0 9647.5 56260.0 ;
      RECT  9582.5 54915.0 9647.5 55100.0 ;
      RECT  9222.5 55032.5 9287.5 54882.5 ;
      RECT  9222.5 55917.5 9287.5 56292.5 ;
      RECT  9412.5 55032.5 9477.5 55917.5 ;
      RECT  9222.5 55917.5 9287.5 56052.5 ;
      RECT  9412.5 55917.5 9477.5 56052.5 ;
      RECT  9412.5 55917.5 9477.5 56052.5 ;
      RECT  9222.5 55917.5 9287.5 56052.5 ;
      RECT  9222.5 55032.5 9287.5 55167.5 ;
      RECT  9412.5 55032.5 9477.5 55167.5 ;
      RECT  9412.5 55032.5 9477.5 55167.5 ;
      RECT  9222.5 55032.5 9287.5 55167.5 ;
      RECT  9582.5 56007.5 9647.5 56142.5 ;
      RECT  9582.5 55032.5 9647.5 55167.5 ;
      RECT  9280.0 55475.0 9345.0 55610.0 ;
      RECT  9280.0 55475.0 9345.0 55610.0 ;
      RECT  9445.0 55510.0 9510.0 55575.0 ;
      RECT  9155.0 56227.5 9715.0 56292.5 ;
      RECT  9155.0 54882.5 9715.0 54947.5 ;
      RECT  9782.5 55077.5 9847.5 54882.5 ;
      RECT  9782.5 55917.5 9847.5 56292.5 ;
      RECT  10162.5 55917.5 10227.5 56292.5 ;
      RECT  10332.5 56075.0 10397.5 56260.0 ;
      RECT  10332.5 54915.0 10397.5 55100.0 ;
      RECT  9782.5 55917.5 9847.5 56052.5 ;
      RECT  9972.5 55917.5 10037.5 56052.5 ;
      RECT  9972.5 55917.5 10037.5 56052.5 ;
      RECT  9782.5 55917.5 9847.5 56052.5 ;
      RECT  9972.5 55917.5 10037.5 56052.5 ;
      RECT  10162.5 55917.5 10227.5 56052.5 ;
      RECT  10162.5 55917.5 10227.5 56052.5 ;
      RECT  9972.5 55917.5 10037.5 56052.5 ;
      RECT  9782.5 55077.5 9847.5 55212.5 ;
      RECT  9972.5 55077.5 10037.5 55212.5 ;
      RECT  9972.5 55077.5 10037.5 55212.5 ;
      RECT  9782.5 55077.5 9847.5 55212.5 ;
      RECT  9972.5 55077.5 10037.5 55212.5 ;
      RECT  10162.5 55077.5 10227.5 55212.5 ;
      RECT  10162.5 55077.5 10227.5 55212.5 ;
      RECT  9972.5 55077.5 10037.5 55212.5 ;
      RECT  10332.5 56007.5 10397.5 56142.5 ;
      RECT  10332.5 55032.5 10397.5 55167.5 ;
      RECT  10167.5 55307.5 10032.5 55372.5 ;
      RECT  9910.0 55522.5 9775.0 55587.5 ;
      RECT  9972.5 55917.5 10037.5 56052.5 ;
      RECT  10162.5 55077.5 10227.5 55212.5 ;
      RECT  10262.5 55522.5 10127.5 55587.5 ;
      RECT  9775.0 55522.5 9910.0 55587.5 ;
      RECT  10032.5 55307.5 10167.5 55372.5 ;
      RECT  10127.5 55522.5 10262.5 55587.5 ;
      RECT  9715.0 56227.5 10635.0 56292.5 ;
      RECT  9715.0 54882.5 10635.0 54947.5 ;
      RECT  11062.5 56075.0 11127.5 56260.0 ;
      RECT  11062.5 54915.0 11127.5 55100.0 ;
      RECT  10702.5 55032.5 10767.5 54882.5 ;
      RECT  10702.5 55917.5 10767.5 56292.5 ;
      RECT  10892.5 55032.5 10957.5 55917.5 ;
      RECT  10702.5 55917.5 10767.5 56052.5 ;
      RECT  10892.5 55917.5 10957.5 56052.5 ;
      RECT  10892.5 55917.5 10957.5 56052.5 ;
      RECT  10702.5 55917.5 10767.5 56052.5 ;
      RECT  10702.5 55032.5 10767.5 55167.5 ;
      RECT  10892.5 55032.5 10957.5 55167.5 ;
      RECT  10892.5 55032.5 10957.5 55167.5 ;
      RECT  10702.5 55032.5 10767.5 55167.5 ;
      RECT  11062.5 56007.5 11127.5 56142.5 ;
      RECT  11062.5 55032.5 11127.5 55167.5 ;
      RECT  10760.0 55475.0 10825.0 55610.0 ;
      RECT  10760.0 55475.0 10825.0 55610.0 ;
      RECT  10925.0 55510.0 10990.0 55575.0 ;
      RECT  10635.0 56227.5 11195.0 56292.5 ;
      RECT  10635.0 54882.5 11195.0 54947.5 ;
      RECT  8897.5 55475.0 8962.5 55610.0 ;
      RECT  9037.5 55202.5 9102.5 55337.5 ;
      RECT  10032.5 55307.5 9897.5 55372.5 ;
      RECT  9582.5 56445.0 9647.5 56260.0 ;
      RECT  9582.5 57605.0 9647.5 57420.0 ;
      RECT  9222.5 57487.5 9287.5 57637.5 ;
      RECT  9222.5 56602.5 9287.5 56227.5 ;
      RECT  9412.5 57487.5 9477.5 56602.5 ;
      RECT  9222.5 56602.5 9287.5 56467.5 ;
      RECT  9412.5 56602.5 9477.5 56467.5 ;
      RECT  9412.5 56602.5 9477.5 56467.5 ;
      RECT  9222.5 56602.5 9287.5 56467.5 ;
      RECT  9222.5 57487.5 9287.5 57352.5 ;
      RECT  9412.5 57487.5 9477.5 57352.5 ;
      RECT  9412.5 57487.5 9477.5 57352.5 ;
      RECT  9222.5 57487.5 9287.5 57352.5 ;
      RECT  9582.5 56512.5 9647.5 56377.5 ;
      RECT  9582.5 57487.5 9647.5 57352.5 ;
      RECT  9280.0 57045.0 9345.0 56910.0 ;
      RECT  9280.0 57045.0 9345.0 56910.0 ;
      RECT  9445.0 57010.0 9510.0 56945.0 ;
      RECT  9155.0 56292.5 9715.0 56227.5 ;
      RECT  9155.0 57637.5 9715.0 57572.5 ;
      RECT  9782.5 57442.5 9847.5 57637.5 ;
      RECT  9782.5 56602.5 9847.5 56227.5 ;
      RECT  10162.5 56602.5 10227.5 56227.5 ;
      RECT  10332.5 56445.0 10397.5 56260.0 ;
      RECT  10332.5 57605.0 10397.5 57420.0 ;
      RECT  9782.5 56602.5 9847.5 56467.5 ;
      RECT  9972.5 56602.5 10037.5 56467.5 ;
      RECT  9972.5 56602.5 10037.5 56467.5 ;
      RECT  9782.5 56602.5 9847.5 56467.5 ;
      RECT  9972.5 56602.5 10037.5 56467.5 ;
      RECT  10162.5 56602.5 10227.5 56467.5 ;
      RECT  10162.5 56602.5 10227.5 56467.5 ;
      RECT  9972.5 56602.5 10037.5 56467.5 ;
      RECT  9782.5 57442.5 9847.5 57307.5 ;
      RECT  9972.5 57442.5 10037.5 57307.5 ;
      RECT  9972.5 57442.5 10037.5 57307.5 ;
      RECT  9782.5 57442.5 9847.5 57307.5 ;
      RECT  9972.5 57442.5 10037.5 57307.5 ;
      RECT  10162.5 57442.5 10227.5 57307.5 ;
      RECT  10162.5 57442.5 10227.5 57307.5 ;
      RECT  9972.5 57442.5 10037.5 57307.5 ;
      RECT  10332.5 56512.5 10397.5 56377.5 ;
      RECT  10332.5 57487.5 10397.5 57352.5 ;
      RECT  10167.5 57212.5 10032.5 57147.5 ;
      RECT  9910.0 56997.5 9775.0 56932.5 ;
      RECT  9972.5 56602.5 10037.5 56467.5 ;
      RECT  10162.5 57442.5 10227.5 57307.5 ;
      RECT  10262.5 56997.5 10127.5 56932.5 ;
      RECT  9775.0 56997.5 9910.0 56932.5 ;
      RECT  10032.5 57212.5 10167.5 57147.5 ;
      RECT  10127.5 56997.5 10262.5 56932.5 ;
      RECT  9715.0 56292.5 10635.0 56227.5 ;
      RECT  9715.0 57637.5 10635.0 57572.5 ;
      RECT  11062.5 56445.0 11127.5 56260.0 ;
      RECT  11062.5 57605.0 11127.5 57420.0 ;
      RECT  10702.5 57487.5 10767.5 57637.5 ;
      RECT  10702.5 56602.5 10767.5 56227.5 ;
      RECT  10892.5 57487.5 10957.5 56602.5 ;
      RECT  10702.5 56602.5 10767.5 56467.5 ;
      RECT  10892.5 56602.5 10957.5 56467.5 ;
      RECT  10892.5 56602.5 10957.5 56467.5 ;
      RECT  10702.5 56602.5 10767.5 56467.5 ;
      RECT  10702.5 57487.5 10767.5 57352.5 ;
      RECT  10892.5 57487.5 10957.5 57352.5 ;
      RECT  10892.5 57487.5 10957.5 57352.5 ;
      RECT  10702.5 57487.5 10767.5 57352.5 ;
      RECT  11062.5 56512.5 11127.5 56377.5 ;
      RECT  11062.5 57487.5 11127.5 57352.5 ;
      RECT  10760.0 57045.0 10825.0 56910.0 ;
      RECT  10760.0 57045.0 10825.0 56910.0 ;
      RECT  10925.0 57010.0 10990.0 56945.0 ;
      RECT  10635.0 56292.5 11195.0 56227.5 ;
      RECT  10635.0 57637.5 11195.0 57572.5 ;
      RECT  8897.5 56910.0 8962.5 57045.0 ;
      RECT  9037.5 57182.5 9102.5 57317.5 ;
      RECT  10032.5 57147.5 9897.5 57212.5 ;
      RECT  9582.5 58765.0 9647.5 58950.0 ;
      RECT  9582.5 57605.0 9647.5 57790.0 ;
      RECT  9222.5 57722.5 9287.5 57572.5 ;
      RECT  9222.5 58607.5 9287.5 58982.5 ;
      RECT  9412.5 57722.5 9477.5 58607.5 ;
      RECT  9222.5 58607.5 9287.5 58742.5 ;
      RECT  9412.5 58607.5 9477.5 58742.5 ;
      RECT  9412.5 58607.5 9477.5 58742.5 ;
      RECT  9222.5 58607.5 9287.5 58742.5 ;
      RECT  9222.5 57722.5 9287.5 57857.5 ;
      RECT  9412.5 57722.5 9477.5 57857.5 ;
      RECT  9412.5 57722.5 9477.5 57857.5 ;
      RECT  9222.5 57722.5 9287.5 57857.5 ;
      RECT  9582.5 58697.5 9647.5 58832.5 ;
      RECT  9582.5 57722.5 9647.5 57857.5 ;
      RECT  9280.0 58165.0 9345.0 58300.0 ;
      RECT  9280.0 58165.0 9345.0 58300.0 ;
      RECT  9445.0 58200.0 9510.0 58265.0 ;
      RECT  9155.0 58917.5 9715.0 58982.5 ;
      RECT  9155.0 57572.5 9715.0 57637.5 ;
      RECT  9782.5 57767.5 9847.5 57572.5 ;
      RECT  9782.5 58607.5 9847.5 58982.5 ;
      RECT  10162.5 58607.5 10227.5 58982.5 ;
      RECT  10332.5 58765.0 10397.5 58950.0 ;
      RECT  10332.5 57605.0 10397.5 57790.0 ;
      RECT  9782.5 58607.5 9847.5 58742.5 ;
      RECT  9972.5 58607.5 10037.5 58742.5 ;
      RECT  9972.5 58607.5 10037.5 58742.5 ;
      RECT  9782.5 58607.5 9847.5 58742.5 ;
      RECT  9972.5 58607.5 10037.5 58742.5 ;
      RECT  10162.5 58607.5 10227.5 58742.5 ;
      RECT  10162.5 58607.5 10227.5 58742.5 ;
      RECT  9972.5 58607.5 10037.5 58742.5 ;
      RECT  9782.5 57767.5 9847.5 57902.5 ;
      RECT  9972.5 57767.5 10037.5 57902.5 ;
      RECT  9972.5 57767.5 10037.5 57902.5 ;
      RECT  9782.5 57767.5 9847.5 57902.5 ;
      RECT  9972.5 57767.5 10037.5 57902.5 ;
      RECT  10162.5 57767.5 10227.5 57902.5 ;
      RECT  10162.5 57767.5 10227.5 57902.5 ;
      RECT  9972.5 57767.5 10037.5 57902.5 ;
      RECT  10332.5 58697.5 10397.5 58832.5 ;
      RECT  10332.5 57722.5 10397.5 57857.5 ;
      RECT  10167.5 57997.5 10032.5 58062.5 ;
      RECT  9910.0 58212.5 9775.0 58277.5 ;
      RECT  9972.5 58607.5 10037.5 58742.5 ;
      RECT  10162.5 57767.5 10227.5 57902.5 ;
      RECT  10262.5 58212.5 10127.5 58277.5 ;
      RECT  9775.0 58212.5 9910.0 58277.5 ;
      RECT  10032.5 57997.5 10167.5 58062.5 ;
      RECT  10127.5 58212.5 10262.5 58277.5 ;
      RECT  9715.0 58917.5 10635.0 58982.5 ;
      RECT  9715.0 57572.5 10635.0 57637.5 ;
      RECT  11062.5 58765.0 11127.5 58950.0 ;
      RECT  11062.5 57605.0 11127.5 57790.0 ;
      RECT  10702.5 57722.5 10767.5 57572.5 ;
      RECT  10702.5 58607.5 10767.5 58982.5 ;
      RECT  10892.5 57722.5 10957.5 58607.5 ;
      RECT  10702.5 58607.5 10767.5 58742.5 ;
      RECT  10892.5 58607.5 10957.5 58742.5 ;
      RECT  10892.5 58607.5 10957.5 58742.5 ;
      RECT  10702.5 58607.5 10767.5 58742.5 ;
      RECT  10702.5 57722.5 10767.5 57857.5 ;
      RECT  10892.5 57722.5 10957.5 57857.5 ;
      RECT  10892.5 57722.5 10957.5 57857.5 ;
      RECT  10702.5 57722.5 10767.5 57857.5 ;
      RECT  11062.5 58697.5 11127.5 58832.5 ;
      RECT  11062.5 57722.5 11127.5 57857.5 ;
      RECT  10760.0 58165.0 10825.0 58300.0 ;
      RECT  10760.0 58165.0 10825.0 58300.0 ;
      RECT  10925.0 58200.0 10990.0 58265.0 ;
      RECT  10635.0 58917.5 11195.0 58982.5 ;
      RECT  10635.0 57572.5 11195.0 57637.5 ;
      RECT  8897.5 58165.0 8962.5 58300.0 ;
      RECT  9037.5 57892.5 9102.5 58027.5 ;
      RECT  10032.5 57997.5 9897.5 58062.5 ;
      RECT  9582.5 59135.0 9647.5 58950.0 ;
      RECT  9582.5 60295.0 9647.5 60110.0 ;
      RECT  9222.5 60177.5 9287.5 60327.5 ;
      RECT  9222.5 59292.5 9287.5 58917.5 ;
      RECT  9412.5 60177.5 9477.5 59292.5 ;
      RECT  9222.5 59292.5 9287.5 59157.5 ;
      RECT  9412.5 59292.5 9477.5 59157.5 ;
      RECT  9412.5 59292.5 9477.5 59157.5 ;
      RECT  9222.5 59292.5 9287.5 59157.5 ;
      RECT  9222.5 60177.5 9287.5 60042.5 ;
      RECT  9412.5 60177.5 9477.5 60042.5 ;
      RECT  9412.5 60177.5 9477.5 60042.5 ;
      RECT  9222.5 60177.5 9287.5 60042.5 ;
      RECT  9582.5 59202.5 9647.5 59067.5 ;
      RECT  9582.5 60177.5 9647.5 60042.5 ;
      RECT  9280.0 59735.0 9345.0 59600.0 ;
      RECT  9280.0 59735.0 9345.0 59600.0 ;
      RECT  9445.0 59700.0 9510.0 59635.0 ;
      RECT  9155.0 58982.5 9715.0 58917.5 ;
      RECT  9155.0 60327.5 9715.0 60262.5 ;
      RECT  9782.5 60132.5 9847.5 60327.5 ;
      RECT  9782.5 59292.5 9847.5 58917.5 ;
      RECT  10162.5 59292.5 10227.5 58917.5 ;
      RECT  10332.5 59135.0 10397.5 58950.0 ;
      RECT  10332.5 60295.0 10397.5 60110.0 ;
      RECT  9782.5 59292.5 9847.5 59157.5 ;
      RECT  9972.5 59292.5 10037.5 59157.5 ;
      RECT  9972.5 59292.5 10037.5 59157.5 ;
      RECT  9782.5 59292.5 9847.5 59157.5 ;
      RECT  9972.5 59292.5 10037.5 59157.5 ;
      RECT  10162.5 59292.5 10227.5 59157.5 ;
      RECT  10162.5 59292.5 10227.5 59157.5 ;
      RECT  9972.5 59292.5 10037.5 59157.5 ;
      RECT  9782.5 60132.5 9847.5 59997.5 ;
      RECT  9972.5 60132.5 10037.5 59997.5 ;
      RECT  9972.5 60132.5 10037.5 59997.5 ;
      RECT  9782.5 60132.5 9847.5 59997.5 ;
      RECT  9972.5 60132.5 10037.5 59997.5 ;
      RECT  10162.5 60132.5 10227.5 59997.5 ;
      RECT  10162.5 60132.5 10227.5 59997.5 ;
      RECT  9972.5 60132.5 10037.5 59997.5 ;
      RECT  10332.5 59202.5 10397.5 59067.5 ;
      RECT  10332.5 60177.5 10397.5 60042.5 ;
      RECT  10167.5 59902.5 10032.5 59837.5 ;
      RECT  9910.0 59687.5 9775.0 59622.5 ;
      RECT  9972.5 59292.5 10037.5 59157.5 ;
      RECT  10162.5 60132.5 10227.5 59997.5 ;
      RECT  10262.5 59687.5 10127.5 59622.5 ;
      RECT  9775.0 59687.5 9910.0 59622.5 ;
      RECT  10032.5 59902.5 10167.5 59837.5 ;
      RECT  10127.5 59687.5 10262.5 59622.5 ;
      RECT  9715.0 58982.5 10635.0 58917.5 ;
      RECT  9715.0 60327.5 10635.0 60262.5 ;
      RECT  11062.5 59135.0 11127.5 58950.0 ;
      RECT  11062.5 60295.0 11127.5 60110.0 ;
      RECT  10702.5 60177.5 10767.5 60327.5 ;
      RECT  10702.5 59292.5 10767.5 58917.5 ;
      RECT  10892.5 60177.5 10957.5 59292.5 ;
      RECT  10702.5 59292.5 10767.5 59157.5 ;
      RECT  10892.5 59292.5 10957.5 59157.5 ;
      RECT  10892.5 59292.5 10957.5 59157.5 ;
      RECT  10702.5 59292.5 10767.5 59157.5 ;
      RECT  10702.5 60177.5 10767.5 60042.5 ;
      RECT  10892.5 60177.5 10957.5 60042.5 ;
      RECT  10892.5 60177.5 10957.5 60042.5 ;
      RECT  10702.5 60177.5 10767.5 60042.5 ;
      RECT  11062.5 59202.5 11127.5 59067.5 ;
      RECT  11062.5 60177.5 11127.5 60042.5 ;
      RECT  10760.0 59735.0 10825.0 59600.0 ;
      RECT  10760.0 59735.0 10825.0 59600.0 ;
      RECT  10925.0 59700.0 10990.0 59635.0 ;
      RECT  10635.0 58982.5 11195.0 58917.5 ;
      RECT  10635.0 60327.5 11195.0 60262.5 ;
      RECT  8897.5 59600.0 8962.5 59735.0 ;
      RECT  9037.5 59872.5 9102.5 60007.5 ;
      RECT  10032.5 59837.5 9897.5 59902.5 ;
      RECT  9582.5 61455.0 9647.5 61640.0 ;
      RECT  9582.5 60295.0 9647.5 60480.0 ;
      RECT  9222.5 60412.5 9287.5 60262.5 ;
      RECT  9222.5 61297.5 9287.5 61672.5 ;
      RECT  9412.5 60412.5 9477.5 61297.5 ;
      RECT  9222.5 61297.5 9287.5 61432.5 ;
      RECT  9412.5 61297.5 9477.5 61432.5 ;
      RECT  9412.5 61297.5 9477.5 61432.5 ;
      RECT  9222.5 61297.5 9287.5 61432.5 ;
      RECT  9222.5 60412.5 9287.5 60547.5 ;
      RECT  9412.5 60412.5 9477.5 60547.5 ;
      RECT  9412.5 60412.5 9477.5 60547.5 ;
      RECT  9222.5 60412.5 9287.5 60547.5 ;
      RECT  9582.5 61387.5 9647.5 61522.5 ;
      RECT  9582.5 60412.5 9647.5 60547.5 ;
      RECT  9280.0 60855.0 9345.0 60990.0 ;
      RECT  9280.0 60855.0 9345.0 60990.0 ;
      RECT  9445.0 60890.0 9510.0 60955.0 ;
      RECT  9155.0 61607.5 9715.0 61672.5 ;
      RECT  9155.0 60262.5 9715.0 60327.5 ;
      RECT  9782.5 60457.5 9847.5 60262.5 ;
      RECT  9782.5 61297.5 9847.5 61672.5 ;
      RECT  10162.5 61297.5 10227.5 61672.5 ;
      RECT  10332.5 61455.0 10397.5 61640.0 ;
      RECT  10332.5 60295.0 10397.5 60480.0 ;
      RECT  9782.5 61297.5 9847.5 61432.5 ;
      RECT  9972.5 61297.5 10037.5 61432.5 ;
      RECT  9972.5 61297.5 10037.5 61432.5 ;
      RECT  9782.5 61297.5 9847.5 61432.5 ;
      RECT  9972.5 61297.5 10037.5 61432.5 ;
      RECT  10162.5 61297.5 10227.5 61432.5 ;
      RECT  10162.5 61297.5 10227.5 61432.5 ;
      RECT  9972.5 61297.5 10037.5 61432.5 ;
      RECT  9782.5 60457.5 9847.5 60592.5 ;
      RECT  9972.5 60457.5 10037.5 60592.5 ;
      RECT  9972.5 60457.5 10037.5 60592.5 ;
      RECT  9782.5 60457.5 9847.5 60592.5 ;
      RECT  9972.5 60457.5 10037.5 60592.5 ;
      RECT  10162.5 60457.5 10227.5 60592.5 ;
      RECT  10162.5 60457.5 10227.5 60592.5 ;
      RECT  9972.5 60457.5 10037.5 60592.5 ;
      RECT  10332.5 61387.5 10397.5 61522.5 ;
      RECT  10332.5 60412.5 10397.5 60547.5 ;
      RECT  10167.5 60687.5 10032.5 60752.5 ;
      RECT  9910.0 60902.5 9775.0 60967.5 ;
      RECT  9972.5 61297.5 10037.5 61432.5 ;
      RECT  10162.5 60457.5 10227.5 60592.5 ;
      RECT  10262.5 60902.5 10127.5 60967.5 ;
      RECT  9775.0 60902.5 9910.0 60967.5 ;
      RECT  10032.5 60687.5 10167.5 60752.5 ;
      RECT  10127.5 60902.5 10262.5 60967.5 ;
      RECT  9715.0 61607.5 10635.0 61672.5 ;
      RECT  9715.0 60262.5 10635.0 60327.5 ;
      RECT  11062.5 61455.0 11127.5 61640.0 ;
      RECT  11062.5 60295.0 11127.5 60480.0 ;
      RECT  10702.5 60412.5 10767.5 60262.5 ;
      RECT  10702.5 61297.5 10767.5 61672.5 ;
      RECT  10892.5 60412.5 10957.5 61297.5 ;
      RECT  10702.5 61297.5 10767.5 61432.5 ;
      RECT  10892.5 61297.5 10957.5 61432.5 ;
      RECT  10892.5 61297.5 10957.5 61432.5 ;
      RECT  10702.5 61297.5 10767.5 61432.5 ;
      RECT  10702.5 60412.5 10767.5 60547.5 ;
      RECT  10892.5 60412.5 10957.5 60547.5 ;
      RECT  10892.5 60412.5 10957.5 60547.5 ;
      RECT  10702.5 60412.5 10767.5 60547.5 ;
      RECT  11062.5 61387.5 11127.5 61522.5 ;
      RECT  11062.5 60412.5 11127.5 60547.5 ;
      RECT  10760.0 60855.0 10825.0 60990.0 ;
      RECT  10760.0 60855.0 10825.0 60990.0 ;
      RECT  10925.0 60890.0 10990.0 60955.0 ;
      RECT  10635.0 61607.5 11195.0 61672.5 ;
      RECT  10635.0 60262.5 11195.0 60327.5 ;
      RECT  8897.5 60855.0 8962.5 60990.0 ;
      RECT  9037.5 60582.5 9102.5 60717.5 ;
      RECT  10032.5 60687.5 9897.5 60752.5 ;
      RECT  9582.5 61825.0 9647.5 61640.0 ;
      RECT  9582.5 62985.0 9647.5 62800.0 ;
      RECT  9222.5 62867.5 9287.5 63017.5 ;
      RECT  9222.5 61982.5 9287.5 61607.5 ;
      RECT  9412.5 62867.5 9477.5 61982.5 ;
      RECT  9222.5 61982.5 9287.5 61847.5 ;
      RECT  9412.5 61982.5 9477.5 61847.5 ;
      RECT  9412.5 61982.5 9477.5 61847.5 ;
      RECT  9222.5 61982.5 9287.5 61847.5 ;
      RECT  9222.5 62867.5 9287.5 62732.5 ;
      RECT  9412.5 62867.5 9477.5 62732.5 ;
      RECT  9412.5 62867.5 9477.5 62732.5 ;
      RECT  9222.5 62867.5 9287.5 62732.5 ;
      RECT  9582.5 61892.5 9647.5 61757.5 ;
      RECT  9582.5 62867.5 9647.5 62732.5 ;
      RECT  9280.0 62425.0 9345.0 62290.0 ;
      RECT  9280.0 62425.0 9345.0 62290.0 ;
      RECT  9445.0 62390.0 9510.0 62325.0 ;
      RECT  9155.0 61672.5 9715.0 61607.5 ;
      RECT  9155.0 63017.5 9715.0 62952.5 ;
      RECT  9782.5 62822.5 9847.5 63017.5 ;
      RECT  9782.5 61982.5 9847.5 61607.5 ;
      RECT  10162.5 61982.5 10227.5 61607.5 ;
      RECT  10332.5 61825.0 10397.5 61640.0 ;
      RECT  10332.5 62985.0 10397.5 62800.0 ;
      RECT  9782.5 61982.5 9847.5 61847.5 ;
      RECT  9972.5 61982.5 10037.5 61847.5 ;
      RECT  9972.5 61982.5 10037.5 61847.5 ;
      RECT  9782.5 61982.5 9847.5 61847.5 ;
      RECT  9972.5 61982.5 10037.5 61847.5 ;
      RECT  10162.5 61982.5 10227.5 61847.5 ;
      RECT  10162.5 61982.5 10227.5 61847.5 ;
      RECT  9972.5 61982.5 10037.5 61847.5 ;
      RECT  9782.5 62822.5 9847.5 62687.5 ;
      RECT  9972.5 62822.5 10037.5 62687.5 ;
      RECT  9972.5 62822.5 10037.5 62687.5 ;
      RECT  9782.5 62822.5 9847.5 62687.5 ;
      RECT  9972.5 62822.5 10037.5 62687.5 ;
      RECT  10162.5 62822.5 10227.5 62687.5 ;
      RECT  10162.5 62822.5 10227.5 62687.5 ;
      RECT  9972.5 62822.5 10037.5 62687.5 ;
      RECT  10332.5 61892.5 10397.5 61757.5 ;
      RECT  10332.5 62867.5 10397.5 62732.5 ;
      RECT  10167.5 62592.5 10032.5 62527.5 ;
      RECT  9910.0 62377.5 9775.0 62312.5 ;
      RECT  9972.5 61982.5 10037.5 61847.5 ;
      RECT  10162.5 62822.5 10227.5 62687.5 ;
      RECT  10262.5 62377.5 10127.5 62312.5 ;
      RECT  9775.0 62377.5 9910.0 62312.5 ;
      RECT  10032.5 62592.5 10167.5 62527.5 ;
      RECT  10127.5 62377.5 10262.5 62312.5 ;
      RECT  9715.0 61672.5 10635.0 61607.5 ;
      RECT  9715.0 63017.5 10635.0 62952.5 ;
      RECT  11062.5 61825.0 11127.5 61640.0 ;
      RECT  11062.5 62985.0 11127.5 62800.0 ;
      RECT  10702.5 62867.5 10767.5 63017.5 ;
      RECT  10702.5 61982.5 10767.5 61607.5 ;
      RECT  10892.5 62867.5 10957.5 61982.5 ;
      RECT  10702.5 61982.5 10767.5 61847.5 ;
      RECT  10892.5 61982.5 10957.5 61847.5 ;
      RECT  10892.5 61982.5 10957.5 61847.5 ;
      RECT  10702.5 61982.5 10767.5 61847.5 ;
      RECT  10702.5 62867.5 10767.5 62732.5 ;
      RECT  10892.5 62867.5 10957.5 62732.5 ;
      RECT  10892.5 62867.5 10957.5 62732.5 ;
      RECT  10702.5 62867.5 10767.5 62732.5 ;
      RECT  11062.5 61892.5 11127.5 61757.5 ;
      RECT  11062.5 62867.5 11127.5 62732.5 ;
      RECT  10760.0 62425.0 10825.0 62290.0 ;
      RECT  10760.0 62425.0 10825.0 62290.0 ;
      RECT  10925.0 62390.0 10990.0 62325.0 ;
      RECT  10635.0 61672.5 11195.0 61607.5 ;
      RECT  10635.0 63017.5 11195.0 62952.5 ;
      RECT  8897.5 62290.0 8962.5 62425.0 ;
      RECT  9037.5 62562.5 9102.5 62697.5 ;
      RECT  10032.5 62527.5 9897.5 62592.5 ;
      RECT  9582.5 64145.0 9647.5 64330.0 ;
      RECT  9582.5 62985.0 9647.5 63170.0 ;
      RECT  9222.5 63102.5 9287.5 62952.5 ;
      RECT  9222.5 63987.5 9287.5 64362.5 ;
      RECT  9412.5 63102.5 9477.5 63987.5 ;
      RECT  9222.5 63987.5 9287.5 64122.5 ;
      RECT  9412.5 63987.5 9477.5 64122.5 ;
      RECT  9412.5 63987.5 9477.5 64122.5 ;
      RECT  9222.5 63987.5 9287.5 64122.5 ;
      RECT  9222.5 63102.5 9287.5 63237.5 ;
      RECT  9412.5 63102.5 9477.5 63237.5 ;
      RECT  9412.5 63102.5 9477.5 63237.5 ;
      RECT  9222.5 63102.5 9287.5 63237.5 ;
      RECT  9582.5 64077.5 9647.5 64212.5 ;
      RECT  9582.5 63102.5 9647.5 63237.5 ;
      RECT  9280.0 63545.0 9345.0 63680.0 ;
      RECT  9280.0 63545.0 9345.0 63680.0 ;
      RECT  9445.0 63580.0 9510.0 63645.0 ;
      RECT  9155.0 64297.5 9715.0 64362.5 ;
      RECT  9155.0 62952.5 9715.0 63017.5 ;
      RECT  9782.5 63147.5 9847.5 62952.5 ;
      RECT  9782.5 63987.5 9847.5 64362.5 ;
      RECT  10162.5 63987.5 10227.5 64362.5 ;
      RECT  10332.5 64145.0 10397.5 64330.0 ;
      RECT  10332.5 62985.0 10397.5 63170.0 ;
      RECT  9782.5 63987.5 9847.5 64122.5 ;
      RECT  9972.5 63987.5 10037.5 64122.5 ;
      RECT  9972.5 63987.5 10037.5 64122.5 ;
      RECT  9782.5 63987.5 9847.5 64122.5 ;
      RECT  9972.5 63987.5 10037.5 64122.5 ;
      RECT  10162.5 63987.5 10227.5 64122.5 ;
      RECT  10162.5 63987.5 10227.5 64122.5 ;
      RECT  9972.5 63987.5 10037.5 64122.5 ;
      RECT  9782.5 63147.5 9847.5 63282.5 ;
      RECT  9972.5 63147.5 10037.5 63282.5 ;
      RECT  9972.5 63147.5 10037.5 63282.5 ;
      RECT  9782.5 63147.5 9847.5 63282.5 ;
      RECT  9972.5 63147.5 10037.5 63282.5 ;
      RECT  10162.5 63147.5 10227.5 63282.5 ;
      RECT  10162.5 63147.5 10227.5 63282.5 ;
      RECT  9972.5 63147.5 10037.5 63282.5 ;
      RECT  10332.5 64077.5 10397.5 64212.5 ;
      RECT  10332.5 63102.5 10397.5 63237.5 ;
      RECT  10167.5 63377.5 10032.5 63442.5 ;
      RECT  9910.0 63592.5 9775.0 63657.5 ;
      RECT  9972.5 63987.5 10037.5 64122.5 ;
      RECT  10162.5 63147.5 10227.5 63282.5 ;
      RECT  10262.5 63592.5 10127.5 63657.5 ;
      RECT  9775.0 63592.5 9910.0 63657.5 ;
      RECT  10032.5 63377.5 10167.5 63442.5 ;
      RECT  10127.5 63592.5 10262.5 63657.5 ;
      RECT  9715.0 64297.5 10635.0 64362.5 ;
      RECT  9715.0 62952.5 10635.0 63017.5 ;
      RECT  11062.5 64145.0 11127.5 64330.0 ;
      RECT  11062.5 62985.0 11127.5 63170.0 ;
      RECT  10702.5 63102.5 10767.5 62952.5 ;
      RECT  10702.5 63987.5 10767.5 64362.5 ;
      RECT  10892.5 63102.5 10957.5 63987.5 ;
      RECT  10702.5 63987.5 10767.5 64122.5 ;
      RECT  10892.5 63987.5 10957.5 64122.5 ;
      RECT  10892.5 63987.5 10957.5 64122.5 ;
      RECT  10702.5 63987.5 10767.5 64122.5 ;
      RECT  10702.5 63102.5 10767.5 63237.5 ;
      RECT  10892.5 63102.5 10957.5 63237.5 ;
      RECT  10892.5 63102.5 10957.5 63237.5 ;
      RECT  10702.5 63102.5 10767.5 63237.5 ;
      RECT  11062.5 64077.5 11127.5 64212.5 ;
      RECT  11062.5 63102.5 11127.5 63237.5 ;
      RECT  10760.0 63545.0 10825.0 63680.0 ;
      RECT  10760.0 63545.0 10825.0 63680.0 ;
      RECT  10925.0 63580.0 10990.0 63645.0 ;
      RECT  10635.0 64297.5 11195.0 64362.5 ;
      RECT  10635.0 62952.5 11195.0 63017.5 ;
      RECT  8897.5 63545.0 8962.5 63680.0 ;
      RECT  9037.5 63272.5 9102.5 63407.5 ;
      RECT  10032.5 63377.5 9897.5 63442.5 ;
      RECT  9582.5 64515.0 9647.5 64330.0 ;
      RECT  9582.5 65675.0 9647.5 65490.0 ;
      RECT  9222.5 65557.5 9287.5 65707.5 ;
      RECT  9222.5 64672.5 9287.5 64297.5 ;
      RECT  9412.5 65557.5 9477.5 64672.5 ;
      RECT  9222.5 64672.5 9287.5 64537.5 ;
      RECT  9412.5 64672.5 9477.5 64537.5 ;
      RECT  9412.5 64672.5 9477.5 64537.5 ;
      RECT  9222.5 64672.5 9287.5 64537.5 ;
      RECT  9222.5 65557.5 9287.5 65422.5 ;
      RECT  9412.5 65557.5 9477.5 65422.5 ;
      RECT  9412.5 65557.5 9477.5 65422.5 ;
      RECT  9222.5 65557.5 9287.5 65422.5 ;
      RECT  9582.5 64582.5 9647.5 64447.5 ;
      RECT  9582.5 65557.5 9647.5 65422.5 ;
      RECT  9280.0 65115.0 9345.0 64980.0 ;
      RECT  9280.0 65115.0 9345.0 64980.0 ;
      RECT  9445.0 65080.0 9510.0 65015.0 ;
      RECT  9155.0 64362.5 9715.0 64297.5 ;
      RECT  9155.0 65707.5 9715.0 65642.5 ;
      RECT  9782.5 65512.5 9847.5 65707.5 ;
      RECT  9782.5 64672.5 9847.5 64297.5 ;
      RECT  10162.5 64672.5 10227.5 64297.5 ;
      RECT  10332.5 64515.0 10397.5 64330.0 ;
      RECT  10332.5 65675.0 10397.5 65490.0 ;
      RECT  9782.5 64672.5 9847.5 64537.5 ;
      RECT  9972.5 64672.5 10037.5 64537.5 ;
      RECT  9972.5 64672.5 10037.5 64537.5 ;
      RECT  9782.5 64672.5 9847.5 64537.5 ;
      RECT  9972.5 64672.5 10037.5 64537.5 ;
      RECT  10162.5 64672.5 10227.5 64537.5 ;
      RECT  10162.5 64672.5 10227.5 64537.5 ;
      RECT  9972.5 64672.5 10037.5 64537.5 ;
      RECT  9782.5 65512.5 9847.5 65377.5 ;
      RECT  9972.5 65512.5 10037.5 65377.5 ;
      RECT  9972.5 65512.5 10037.5 65377.5 ;
      RECT  9782.5 65512.5 9847.5 65377.5 ;
      RECT  9972.5 65512.5 10037.5 65377.5 ;
      RECT  10162.5 65512.5 10227.5 65377.5 ;
      RECT  10162.5 65512.5 10227.5 65377.5 ;
      RECT  9972.5 65512.5 10037.5 65377.5 ;
      RECT  10332.5 64582.5 10397.5 64447.5 ;
      RECT  10332.5 65557.5 10397.5 65422.5 ;
      RECT  10167.5 65282.5 10032.5 65217.5 ;
      RECT  9910.0 65067.5 9775.0 65002.5 ;
      RECT  9972.5 64672.5 10037.5 64537.5 ;
      RECT  10162.5 65512.5 10227.5 65377.5 ;
      RECT  10262.5 65067.5 10127.5 65002.5 ;
      RECT  9775.0 65067.5 9910.0 65002.5 ;
      RECT  10032.5 65282.5 10167.5 65217.5 ;
      RECT  10127.5 65067.5 10262.5 65002.5 ;
      RECT  9715.0 64362.5 10635.0 64297.5 ;
      RECT  9715.0 65707.5 10635.0 65642.5 ;
      RECT  11062.5 64515.0 11127.5 64330.0 ;
      RECT  11062.5 65675.0 11127.5 65490.0 ;
      RECT  10702.5 65557.5 10767.5 65707.5 ;
      RECT  10702.5 64672.5 10767.5 64297.5 ;
      RECT  10892.5 65557.5 10957.5 64672.5 ;
      RECT  10702.5 64672.5 10767.5 64537.5 ;
      RECT  10892.5 64672.5 10957.5 64537.5 ;
      RECT  10892.5 64672.5 10957.5 64537.5 ;
      RECT  10702.5 64672.5 10767.5 64537.5 ;
      RECT  10702.5 65557.5 10767.5 65422.5 ;
      RECT  10892.5 65557.5 10957.5 65422.5 ;
      RECT  10892.5 65557.5 10957.5 65422.5 ;
      RECT  10702.5 65557.5 10767.5 65422.5 ;
      RECT  11062.5 64582.5 11127.5 64447.5 ;
      RECT  11062.5 65557.5 11127.5 65422.5 ;
      RECT  10760.0 65115.0 10825.0 64980.0 ;
      RECT  10760.0 65115.0 10825.0 64980.0 ;
      RECT  10925.0 65080.0 10990.0 65015.0 ;
      RECT  10635.0 64362.5 11195.0 64297.5 ;
      RECT  10635.0 65707.5 11195.0 65642.5 ;
      RECT  8897.5 64980.0 8962.5 65115.0 ;
      RECT  9037.5 65252.5 9102.5 65387.5 ;
      RECT  10032.5 65217.5 9897.5 65282.5 ;
      RECT  9582.5 66835.0 9647.5 67020.0 ;
      RECT  9582.5 65675.0 9647.5 65860.0 ;
      RECT  9222.5 65792.5 9287.5 65642.5 ;
      RECT  9222.5 66677.5 9287.5 67052.5 ;
      RECT  9412.5 65792.5 9477.5 66677.5 ;
      RECT  9222.5 66677.5 9287.5 66812.5 ;
      RECT  9412.5 66677.5 9477.5 66812.5 ;
      RECT  9412.5 66677.5 9477.5 66812.5 ;
      RECT  9222.5 66677.5 9287.5 66812.5 ;
      RECT  9222.5 65792.5 9287.5 65927.5 ;
      RECT  9412.5 65792.5 9477.5 65927.5 ;
      RECT  9412.5 65792.5 9477.5 65927.5 ;
      RECT  9222.5 65792.5 9287.5 65927.5 ;
      RECT  9582.5 66767.5 9647.5 66902.5 ;
      RECT  9582.5 65792.5 9647.5 65927.5 ;
      RECT  9280.0 66235.0 9345.0 66370.0 ;
      RECT  9280.0 66235.0 9345.0 66370.0 ;
      RECT  9445.0 66270.0 9510.0 66335.0 ;
      RECT  9155.0 66987.5 9715.0 67052.5 ;
      RECT  9155.0 65642.5 9715.0 65707.5 ;
      RECT  9782.5 65837.5 9847.5 65642.5 ;
      RECT  9782.5 66677.5 9847.5 67052.5 ;
      RECT  10162.5 66677.5 10227.5 67052.5 ;
      RECT  10332.5 66835.0 10397.5 67020.0 ;
      RECT  10332.5 65675.0 10397.5 65860.0 ;
      RECT  9782.5 66677.5 9847.5 66812.5 ;
      RECT  9972.5 66677.5 10037.5 66812.5 ;
      RECT  9972.5 66677.5 10037.5 66812.5 ;
      RECT  9782.5 66677.5 9847.5 66812.5 ;
      RECT  9972.5 66677.5 10037.5 66812.5 ;
      RECT  10162.5 66677.5 10227.5 66812.5 ;
      RECT  10162.5 66677.5 10227.5 66812.5 ;
      RECT  9972.5 66677.5 10037.5 66812.5 ;
      RECT  9782.5 65837.5 9847.5 65972.5 ;
      RECT  9972.5 65837.5 10037.5 65972.5 ;
      RECT  9972.5 65837.5 10037.5 65972.5 ;
      RECT  9782.5 65837.5 9847.5 65972.5 ;
      RECT  9972.5 65837.5 10037.5 65972.5 ;
      RECT  10162.5 65837.5 10227.5 65972.5 ;
      RECT  10162.5 65837.5 10227.5 65972.5 ;
      RECT  9972.5 65837.5 10037.5 65972.5 ;
      RECT  10332.5 66767.5 10397.5 66902.5 ;
      RECT  10332.5 65792.5 10397.5 65927.5 ;
      RECT  10167.5 66067.5 10032.5 66132.5 ;
      RECT  9910.0 66282.5 9775.0 66347.5 ;
      RECT  9972.5 66677.5 10037.5 66812.5 ;
      RECT  10162.5 65837.5 10227.5 65972.5 ;
      RECT  10262.5 66282.5 10127.5 66347.5 ;
      RECT  9775.0 66282.5 9910.0 66347.5 ;
      RECT  10032.5 66067.5 10167.5 66132.5 ;
      RECT  10127.5 66282.5 10262.5 66347.5 ;
      RECT  9715.0 66987.5 10635.0 67052.5 ;
      RECT  9715.0 65642.5 10635.0 65707.5 ;
      RECT  11062.5 66835.0 11127.5 67020.0 ;
      RECT  11062.5 65675.0 11127.5 65860.0 ;
      RECT  10702.5 65792.5 10767.5 65642.5 ;
      RECT  10702.5 66677.5 10767.5 67052.5 ;
      RECT  10892.5 65792.5 10957.5 66677.5 ;
      RECT  10702.5 66677.5 10767.5 66812.5 ;
      RECT  10892.5 66677.5 10957.5 66812.5 ;
      RECT  10892.5 66677.5 10957.5 66812.5 ;
      RECT  10702.5 66677.5 10767.5 66812.5 ;
      RECT  10702.5 65792.5 10767.5 65927.5 ;
      RECT  10892.5 65792.5 10957.5 65927.5 ;
      RECT  10892.5 65792.5 10957.5 65927.5 ;
      RECT  10702.5 65792.5 10767.5 65927.5 ;
      RECT  11062.5 66767.5 11127.5 66902.5 ;
      RECT  11062.5 65792.5 11127.5 65927.5 ;
      RECT  10760.0 66235.0 10825.0 66370.0 ;
      RECT  10760.0 66235.0 10825.0 66370.0 ;
      RECT  10925.0 66270.0 10990.0 66335.0 ;
      RECT  10635.0 66987.5 11195.0 67052.5 ;
      RECT  10635.0 65642.5 11195.0 65707.5 ;
      RECT  8897.5 66235.0 8962.5 66370.0 ;
      RECT  9037.5 65962.5 9102.5 66097.5 ;
      RECT  10032.5 66067.5 9897.5 66132.5 ;
      RECT  9582.5 67205.0 9647.5 67020.0 ;
      RECT  9582.5 68365.0 9647.5 68180.0 ;
      RECT  9222.5 68247.5 9287.5 68397.5 ;
      RECT  9222.5 67362.5 9287.5 66987.5 ;
      RECT  9412.5 68247.5 9477.5 67362.5 ;
      RECT  9222.5 67362.5 9287.5 67227.5 ;
      RECT  9412.5 67362.5 9477.5 67227.5 ;
      RECT  9412.5 67362.5 9477.5 67227.5 ;
      RECT  9222.5 67362.5 9287.5 67227.5 ;
      RECT  9222.5 68247.5 9287.5 68112.5 ;
      RECT  9412.5 68247.5 9477.5 68112.5 ;
      RECT  9412.5 68247.5 9477.5 68112.5 ;
      RECT  9222.5 68247.5 9287.5 68112.5 ;
      RECT  9582.5 67272.5 9647.5 67137.5 ;
      RECT  9582.5 68247.5 9647.5 68112.5 ;
      RECT  9280.0 67805.0 9345.0 67670.0 ;
      RECT  9280.0 67805.0 9345.0 67670.0 ;
      RECT  9445.0 67770.0 9510.0 67705.0 ;
      RECT  9155.0 67052.5 9715.0 66987.5 ;
      RECT  9155.0 68397.5 9715.0 68332.5 ;
      RECT  9782.5 68202.5 9847.5 68397.5 ;
      RECT  9782.5 67362.5 9847.5 66987.5 ;
      RECT  10162.5 67362.5 10227.5 66987.5 ;
      RECT  10332.5 67205.0 10397.5 67020.0 ;
      RECT  10332.5 68365.0 10397.5 68180.0 ;
      RECT  9782.5 67362.5 9847.5 67227.5 ;
      RECT  9972.5 67362.5 10037.5 67227.5 ;
      RECT  9972.5 67362.5 10037.5 67227.5 ;
      RECT  9782.5 67362.5 9847.5 67227.5 ;
      RECT  9972.5 67362.5 10037.5 67227.5 ;
      RECT  10162.5 67362.5 10227.5 67227.5 ;
      RECT  10162.5 67362.5 10227.5 67227.5 ;
      RECT  9972.5 67362.5 10037.5 67227.5 ;
      RECT  9782.5 68202.5 9847.5 68067.5 ;
      RECT  9972.5 68202.5 10037.5 68067.5 ;
      RECT  9972.5 68202.5 10037.5 68067.5 ;
      RECT  9782.5 68202.5 9847.5 68067.5 ;
      RECT  9972.5 68202.5 10037.5 68067.5 ;
      RECT  10162.5 68202.5 10227.5 68067.5 ;
      RECT  10162.5 68202.5 10227.5 68067.5 ;
      RECT  9972.5 68202.5 10037.5 68067.5 ;
      RECT  10332.5 67272.5 10397.5 67137.5 ;
      RECT  10332.5 68247.5 10397.5 68112.5 ;
      RECT  10167.5 67972.5 10032.5 67907.5 ;
      RECT  9910.0 67757.5 9775.0 67692.5 ;
      RECT  9972.5 67362.5 10037.5 67227.5 ;
      RECT  10162.5 68202.5 10227.5 68067.5 ;
      RECT  10262.5 67757.5 10127.5 67692.5 ;
      RECT  9775.0 67757.5 9910.0 67692.5 ;
      RECT  10032.5 67972.5 10167.5 67907.5 ;
      RECT  10127.5 67757.5 10262.5 67692.5 ;
      RECT  9715.0 67052.5 10635.0 66987.5 ;
      RECT  9715.0 68397.5 10635.0 68332.5 ;
      RECT  11062.5 67205.0 11127.5 67020.0 ;
      RECT  11062.5 68365.0 11127.5 68180.0 ;
      RECT  10702.5 68247.5 10767.5 68397.5 ;
      RECT  10702.5 67362.5 10767.5 66987.5 ;
      RECT  10892.5 68247.5 10957.5 67362.5 ;
      RECT  10702.5 67362.5 10767.5 67227.5 ;
      RECT  10892.5 67362.5 10957.5 67227.5 ;
      RECT  10892.5 67362.5 10957.5 67227.5 ;
      RECT  10702.5 67362.5 10767.5 67227.5 ;
      RECT  10702.5 68247.5 10767.5 68112.5 ;
      RECT  10892.5 68247.5 10957.5 68112.5 ;
      RECT  10892.5 68247.5 10957.5 68112.5 ;
      RECT  10702.5 68247.5 10767.5 68112.5 ;
      RECT  11062.5 67272.5 11127.5 67137.5 ;
      RECT  11062.5 68247.5 11127.5 68112.5 ;
      RECT  10760.0 67805.0 10825.0 67670.0 ;
      RECT  10760.0 67805.0 10825.0 67670.0 ;
      RECT  10925.0 67770.0 10990.0 67705.0 ;
      RECT  10635.0 67052.5 11195.0 66987.5 ;
      RECT  10635.0 68397.5 11195.0 68332.5 ;
      RECT  8897.5 67670.0 8962.5 67805.0 ;
      RECT  9037.5 67942.5 9102.5 68077.5 ;
      RECT  10032.5 67907.5 9897.5 67972.5 ;
      RECT  9582.5 69525.0 9647.5 69710.0 ;
      RECT  9582.5 68365.0 9647.5 68550.0 ;
      RECT  9222.5 68482.5 9287.5 68332.5 ;
      RECT  9222.5 69367.5 9287.5 69742.5 ;
      RECT  9412.5 68482.5 9477.5 69367.5 ;
      RECT  9222.5 69367.5 9287.5 69502.5 ;
      RECT  9412.5 69367.5 9477.5 69502.5 ;
      RECT  9412.5 69367.5 9477.5 69502.5 ;
      RECT  9222.5 69367.5 9287.5 69502.5 ;
      RECT  9222.5 68482.5 9287.5 68617.5 ;
      RECT  9412.5 68482.5 9477.5 68617.5 ;
      RECT  9412.5 68482.5 9477.5 68617.5 ;
      RECT  9222.5 68482.5 9287.5 68617.5 ;
      RECT  9582.5 69457.5 9647.5 69592.5 ;
      RECT  9582.5 68482.5 9647.5 68617.5 ;
      RECT  9280.0 68925.0 9345.0 69060.0 ;
      RECT  9280.0 68925.0 9345.0 69060.0 ;
      RECT  9445.0 68960.0 9510.0 69025.0 ;
      RECT  9155.0 69677.5 9715.0 69742.5 ;
      RECT  9155.0 68332.5 9715.0 68397.5 ;
      RECT  9782.5 68527.5 9847.5 68332.5 ;
      RECT  9782.5 69367.5 9847.5 69742.5 ;
      RECT  10162.5 69367.5 10227.5 69742.5 ;
      RECT  10332.5 69525.0 10397.5 69710.0 ;
      RECT  10332.5 68365.0 10397.5 68550.0 ;
      RECT  9782.5 69367.5 9847.5 69502.5 ;
      RECT  9972.5 69367.5 10037.5 69502.5 ;
      RECT  9972.5 69367.5 10037.5 69502.5 ;
      RECT  9782.5 69367.5 9847.5 69502.5 ;
      RECT  9972.5 69367.5 10037.5 69502.5 ;
      RECT  10162.5 69367.5 10227.5 69502.5 ;
      RECT  10162.5 69367.5 10227.5 69502.5 ;
      RECT  9972.5 69367.5 10037.5 69502.5 ;
      RECT  9782.5 68527.5 9847.5 68662.5 ;
      RECT  9972.5 68527.5 10037.5 68662.5 ;
      RECT  9972.5 68527.5 10037.5 68662.5 ;
      RECT  9782.5 68527.5 9847.5 68662.5 ;
      RECT  9972.5 68527.5 10037.5 68662.5 ;
      RECT  10162.5 68527.5 10227.5 68662.5 ;
      RECT  10162.5 68527.5 10227.5 68662.5 ;
      RECT  9972.5 68527.5 10037.5 68662.5 ;
      RECT  10332.5 69457.5 10397.5 69592.5 ;
      RECT  10332.5 68482.5 10397.5 68617.5 ;
      RECT  10167.5 68757.5 10032.5 68822.5 ;
      RECT  9910.0 68972.5 9775.0 69037.5 ;
      RECT  9972.5 69367.5 10037.5 69502.5 ;
      RECT  10162.5 68527.5 10227.5 68662.5 ;
      RECT  10262.5 68972.5 10127.5 69037.5 ;
      RECT  9775.0 68972.5 9910.0 69037.5 ;
      RECT  10032.5 68757.5 10167.5 68822.5 ;
      RECT  10127.5 68972.5 10262.5 69037.5 ;
      RECT  9715.0 69677.5 10635.0 69742.5 ;
      RECT  9715.0 68332.5 10635.0 68397.5 ;
      RECT  11062.5 69525.0 11127.5 69710.0 ;
      RECT  11062.5 68365.0 11127.5 68550.0 ;
      RECT  10702.5 68482.5 10767.5 68332.5 ;
      RECT  10702.5 69367.5 10767.5 69742.5 ;
      RECT  10892.5 68482.5 10957.5 69367.5 ;
      RECT  10702.5 69367.5 10767.5 69502.5 ;
      RECT  10892.5 69367.5 10957.5 69502.5 ;
      RECT  10892.5 69367.5 10957.5 69502.5 ;
      RECT  10702.5 69367.5 10767.5 69502.5 ;
      RECT  10702.5 68482.5 10767.5 68617.5 ;
      RECT  10892.5 68482.5 10957.5 68617.5 ;
      RECT  10892.5 68482.5 10957.5 68617.5 ;
      RECT  10702.5 68482.5 10767.5 68617.5 ;
      RECT  11062.5 69457.5 11127.5 69592.5 ;
      RECT  11062.5 68482.5 11127.5 68617.5 ;
      RECT  10760.0 68925.0 10825.0 69060.0 ;
      RECT  10760.0 68925.0 10825.0 69060.0 ;
      RECT  10925.0 68960.0 10990.0 69025.0 ;
      RECT  10635.0 69677.5 11195.0 69742.5 ;
      RECT  10635.0 68332.5 11195.0 68397.5 ;
      RECT  8897.5 68925.0 8962.5 69060.0 ;
      RECT  9037.5 68652.5 9102.5 68787.5 ;
      RECT  10032.5 68757.5 9897.5 68822.5 ;
      RECT  9582.5 69895.0 9647.5 69710.0 ;
      RECT  9582.5 71055.0 9647.5 70870.0 ;
      RECT  9222.5 70937.5 9287.5 71087.5 ;
      RECT  9222.5 70052.5 9287.5 69677.5 ;
      RECT  9412.5 70937.5 9477.5 70052.5 ;
      RECT  9222.5 70052.5 9287.5 69917.5 ;
      RECT  9412.5 70052.5 9477.5 69917.5 ;
      RECT  9412.5 70052.5 9477.5 69917.5 ;
      RECT  9222.5 70052.5 9287.5 69917.5 ;
      RECT  9222.5 70937.5 9287.5 70802.5 ;
      RECT  9412.5 70937.5 9477.5 70802.5 ;
      RECT  9412.5 70937.5 9477.5 70802.5 ;
      RECT  9222.5 70937.5 9287.5 70802.5 ;
      RECT  9582.5 69962.5 9647.5 69827.5 ;
      RECT  9582.5 70937.5 9647.5 70802.5 ;
      RECT  9280.0 70495.0 9345.0 70360.0 ;
      RECT  9280.0 70495.0 9345.0 70360.0 ;
      RECT  9445.0 70460.0 9510.0 70395.0 ;
      RECT  9155.0 69742.5 9715.0 69677.5 ;
      RECT  9155.0 71087.5 9715.0 71022.5 ;
      RECT  9782.5 70892.5 9847.5 71087.5 ;
      RECT  9782.5 70052.5 9847.5 69677.5 ;
      RECT  10162.5 70052.5 10227.5 69677.5 ;
      RECT  10332.5 69895.0 10397.5 69710.0 ;
      RECT  10332.5 71055.0 10397.5 70870.0 ;
      RECT  9782.5 70052.5 9847.5 69917.5 ;
      RECT  9972.5 70052.5 10037.5 69917.5 ;
      RECT  9972.5 70052.5 10037.5 69917.5 ;
      RECT  9782.5 70052.5 9847.5 69917.5 ;
      RECT  9972.5 70052.5 10037.5 69917.5 ;
      RECT  10162.5 70052.5 10227.5 69917.5 ;
      RECT  10162.5 70052.5 10227.5 69917.5 ;
      RECT  9972.5 70052.5 10037.5 69917.5 ;
      RECT  9782.5 70892.5 9847.5 70757.5 ;
      RECT  9972.5 70892.5 10037.5 70757.5 ;
      RECT  9972.5 70892.5 10037.5 70757.5 ;
      RECT  9782.5 70892.5 9847.5 70757.5 ;
      RECT  9972.5 70892.5 10037.5 70757.5 ;
      RECT  10162.5 70892.5 10227.5 70757.5 ;
      RECT  10162.5 70892.5 10227.5 70757.5 ;
      RECT  9972.5 70892.5 10037.5 70757.5 ;
      RECT  10332.5 69962.5 10397.5 69827.5 ;
      RECT  10332.5 70937.5 10397.5 70802.5 ;
      RECT  10167.5 70662.5 10032.5 70597.5 ;
      RECT  9910.0 70447.5 9775.0 70382.5 ;
      RECT  9972.5 70052.5 10037.5 69917.5 ;
      RECT  10162.5 70892.5 10227.5 70757.5 ;
      RECT  10262.5 70447.5 10127.5 70382.5 ;
      RECT  9775.0 70447.5 9910.0 70382.5 ;
      RECT  10032.5 70662.5 10167.5 70597.5 ;
      RECT  10127.5 70447.5 10262.5 70382.5 ;
      RECT  9715.0 69742.5 10635.0 69677.5 ;
      RECT  9715.0 71087.5 10635.0 71022.5 ;
      RECT  11062.5 69895.0 11127.5 69710.0 ;
      RECT  11062.5 71055.0 11127.5 70870.0 ;
      RECT  10702.5 70937.5 10767.5 71087.5 ;
      RECT  10702.5 70052.5 10767.5 69677.5 ;
      RECT  10892.5 70937.5 10957.5 70052.5 ;
      RECT  10702.5 70052.5 10767.5 69917.5 ;
      RECT  10892.5 70052.5 10957.5 69917.5 ;
      RECT  10892.5 70052.5 10957.5 69917.5 ;
      RECT  10702.5 70052.5 10767.5 69917.5 ;
      RECT  10702.5 70937.5 10767.5 70802.5 ;
      RECT  10892.5 70937.5 10957.5 70802.5 ;
      RECT  10892.5 70937.5 10957.5 70802.5 ;
      RECT  10702.5 70937.5 10767.5 70802.5 ;
      RECT  11062.5 69962.5 11127.5 69827.5 ;
      RECT  11062.5 70937.5 11127.5 70802.5 ;
      RECT  10760.0 70495.0 10825.0 70360.0 ;
      RECT  10760.0 70495.0 10825.0 70360.0 ;
      RECT  10925.0 70460.0 10990.0 70395.0 ;
      RECT  10635.0 69742.5 11195.0 69677.5 ;
      RECT  10635.0 71087.5 11195.0 71022.5 ;
      RECT  8897.5 70360.0 8962.5 70495.0 ;
      RECT  9037.5 70632.5 9102.5 70767.5 ;
      RECT  10032.5 70597.5 9897.5 70662.5 ;
      RECT  9582.5 72215.0 9647.5 72400.0 ;
      RECT  9582.5 71055.0 9647.5 71240.0 ;
      RECT  9222.5 71172.5 9287.5 71022.5 ;
      RECT  9222.5 72057.5 9287.5 72432.5 ;
      RECT  9412.5 71172.5 9477.5 72057.5 ;
      RECT  9222.5 72057.5 9287.5 72192.5 ;
      RECT  9412.5 72057.5 9477.5 72192.5 ;
      RECT  9412.5 72057.5 9477.5 72192.5 ;
      RECT  9222.5 72057.5 9287.5 72192.5 ;
      RECT  9222.5 71172.5 9287.5 71307.5 ;
      RECT  9412.5 71172.5 9477.5 71307.5 ;
      RECT  9412.5 71172.5 9477.5 71307.5 ;
      RECT  9222.5 71172.5 9287.5 71307.5 ;
      RECT  9582.5 72147.5 9647.5 72282.5 ;
      RECT  9582.5 71172.5 9647.5 71307.5 ;
      RECT  9280.0 71615.0 9345.0 71750.0 ;
      RECT  9280.0 71615.0 9345.0 71750.0 ;
      RECT  9445.0 71650.0 9510.0 71715.0 ;
      RECT  9155.0 72367.5 9715.0 72432.5 ;
      RECT  9155.0 71022.5 9715.0 71087.5 ;
      RECT  9782.5 71217.5 9847.5 71022.5 ;
      RECT  9782.5 72057.5 9847.5 72432.5 ;
      RECT  10162.5 72057.5 10227.5 72432.5 ;
      RECT  10332.5 72215.0 10397.5 72400.0 ;
      RECT  10332.5 71055.0 10397.5 71240.0 ;
      RECT  9782.5 72057.5 9847.5 72192.5 ;
      RECT  9972.5 72057.5 10037.5 72192.5 ;
      RECT  9972.5 72057.5 10037.5 72192.5 ;
      RECT  9782.5 72057.5 9847.5 72192.5 ;
      RECT  9972.5 72057.5 10037.5 72192.5 ;
      RECT  10162.5 72057.5 10227.5 72192.5 ;
      RECT  10162.5 72057.5 10227.5 72192.5 ;
      RECT  9972.5 72057.5 10037.5 72192.5 ;
      RECT  9782.5 71217.5 9847.5 71352.5 ;
      RECT  9972.5 71217.5 10037.5 71352.5 ;
      RECT  9972.5 71217.5 10037.5 71352.5 ;
      RECT  9782.5 71217.5 9847.5 71352.5 ;
      RECT  9972.5 71217.5 10037.5 71352.5 ;
      RECT  10162.5 71217.5 10227.5 71352.5 ;
      RECT  10162.5 71217.5 10227.5 71352.5 ;
      RECT  9972.5 71217.5 10037.5 71352.5 ;
      RECT  10332.5 72147.5 10397.5 72282.5 ;
      RECT  10332.5 71172.5 10397.5 71307.5 ;
      RECT  10167.5 71447.5 10032.5 71512.5 ;
      RECT  9910.0 71662.5 9775.0 71727.5 ;
      RECT  9972.5 72057.5 10037.5 72192.5 ;
      RECT  10162.5 71217.5 10227.5 71352.5 ;
      RECT  10262.5 71662.5 10127.5 71727.5 ;
      RECT  9775.0 71662.5 9910.0 71727.5 ;
      RECT  10032.5 71447.5 10167.5 71512.5 ;
      RECT  10127.5 71662.5 10262.5 71727.5 ;
      RECT  9715.0 72367.5 10635.0 72432.5 ;
      RECT  9715.0 71022.5 10635.0 71087.5 ;
      RECT  11062.5 72215.0 11127.5 72400.0 ;
      RECT  11062.5 71055.0 11127.5 71240.0 ;
      RECT  10702.5 71172.5 10767.5 71022.5 ;
      RECT  10702.5 72057.5 10767.5 72432.5 ;
      RECT  10892.5 71172.5 10957.5 72057.5 ;
      RECT  10702.5 72057.5 10767.5 72192.5 ;
      RECT  10892.5 72057.5 10957.5 72192.5 ;
      RECT  10892.5 72057.5 10957.5 72192.5 ;
      RECT  10702.5 72057.5 10767.5 72192.5 ;
      RECT  10702.5 71172.5 10767.5 71307.5 ;
      RECT  10892.5 71172.5 10957.5 71307.5 ;
      RECT  10892.5 71172.5 10957.5 71307.5 ;
      RECT  10702.5 71172.5 10767.5 71307.5 ;
      RECT  11062.5 72147.5 11127.5 72282.5 ;
      RECT  11062.5 71172.5 11127.5 71307.5 ;
      RECT  10760.0 71615.0 10825.0 71750.0 ;
      RECT  10760.0 71615.0 10825.0 71750.0 ;
      RECT  10925.0 71650.0 10990.0 71715.0 ;
      RECT  10635.0 72367.5 11195.0 72432.5 ;
      RECT  10635.0 71022.5 11195.0 71087.5 ;
      RECT  8897.5 71615.0 8962.5 71750.0 ;
      RECT  9037.5 71342.5 9102.5 71477.5 ;
      RECT  10032.5 71447.5 9897.5 71512.5 ;
      RECT  9582.5 72585.0 9647.5 72400.0 ;
      RECT  9582.5 73745.0 9647.5 73560.0 ;
      RECT  9222.5 73627.5 9287.5 73777.5 ;
      RECT  9222.5 72742.5 9287.5 72367.5 ;
      RECT  9412.5 73627.5 9477.5 72742.5 ;
      RECT  9222.5 72742.5 9287.5 72607.5 ;
      RECT  9412.5 72742.5 9477.5 72607.5 ;
      RECT  9412.5 72742.5 9477.5 72607.5 ;
      RECT  9222.5 72742.5 9287.5 72607.5 ;
      RECT  9222.5 73627.5 9287.5 73492.5 ;
      RECT  9412.5 73627.5 9477.5 73492.5 ;
      RECT  9412.5 73627.5 9477.5 73492.5 ;
      RECT  9222.5 73627.5 9287.5 73492.5 ;
      RECT  9582.5 72652.5 9647.5 72517.5 ;
      RECT  9582.5 73627.5 9647.5 73492.5 ;
      RECT  9280.0 73185.0 9345.0 73050.0 ;
      RECT  9280.0 73185.0 9345.0 73050.0 ;
      RECT  9445.0 73150.0 9510.0 73085.0 ;
      RECT  9155.0 72432.5 9715.0 72367.5 ;
      RECT  9155.0 73777.5 9715.0 73712.5 ;
      RECT  9782.5 73582.5 9847.5 73777.5 ;
      RECT  9782.5 72742.5 9847.5 72367.5 ;
      RECT  10162.5 72742.5 10227.5 72367.5 ;
      RECT  10332.5 72585.0 10397.5 72400.0 ;
      RECT  10332.5 73745.0 10397.5 73560.0 ;
      RECT  9782.5 72742.5 9847.5 72607.5 ;
      RECT  9972.5 72742.5 10037.5 72607.5 ;
      RECT  9972.5 72742.5 10037.5 72607.5 ;
      RECT  9782.5 72742.5 9847.5 72607.5 ;
      RECT  9972.5 72742.5 10037.5 72607.5 ;
      RECT  10162.5 72742.5 10227.5 72607.5 ;
      RECT  10162.5 72742.5 10227.5 72607.5 ;
      RECT  9972.5 72742.5 10037.5 72607.5 ;
      RECT  9782.5 73582.5 9847.5 73447.5 ;
      RECT  9972.5 73582.5 10037.5 73447.5 ;
      RECT  9972.5 73582.5 10037.5 73447.5 ;
      RECT  9782.5 73582.5 9847.5 73447.5 ;
      RECT  9972.5 73582.5 10037.5 73447.5 ;
      RECT  10162.5 73582.5 10227.5 73447.5 ;
      RECT  10162.5 73582.5 10227.5 73447.5 ;
      RECT  9972.5 73582.5 10037.5 73447.5 ;
      RECT  10332.5 72652.5 10397.5 72517.5 ;
      RECT  10332.5 73627.5 10397.5 73492.5 ;
      RECT  10167.5 73352.5 10032.5 73287.5 ;
      RECT  9910.0 73137.5 9775.0 73072.5 ;
      RECT  9972.5 72742.5 10037.5 72607.5 ;
      RECT  10162.5 73582.5 10227.5 73447.5 ;
      RECT  10262.5 73137.5 10127.5 73072.5 ;
      RECT  9775.0 73137.5 9910.0 73072.5 ;
      RECT  10032.5 73352.5 10167.5 73287.5 ;
      RECT  10127.5 73137.5 10262.5 73072.5 ;
      RECT  9715.0 72432.5 10635.0 72367.5 ;
      RECT  9715.0 73777.5 10635.0 73712.5 ;
      RECT  11062.5 72585.0 11127.5 72400.0 ;
      RECT  11062.5 73745.0 11127.5 73560.0 ;
      RECT  10702.5 73627.5 10767.5 73777.5 ;
      RECT  10702.5 72742.5 10767.5 72367.5 ;
      RECT  10892.5 73627.5 10957.5 72742.5 ;
      RECT  10702.5 72742.5 10767.5 72607.5 ;
      RECT  10892.5 72742.5 10957.5 72607.5 ;
      RECT  10892.5 72742.5 10957.5 72607.5 ;
      RECT  10702.5 72742.5 10767.5 72607.5 ;
      RECT  10702.5 73627.5 10767.5 73492.5 ;
      RECT  10892.5 73627.5 10957.5 73492.5 ;
      RECT  10892.5 73627.5 10957.5 73492.5 ;
      RECT  10702.5 73627.5 10767.5 73492.5 ;
      RECT  11062.5 72652.5 11127.5 72517.5 ;
      RECT  11062.5 73627.5 11127.5 73492.5 ;
      RECT  10760.0 73185.0 10825.0 73050.0 ;
      RECT  10760.0 73185.0 10825.0 73050.0 ;
      RECT  10925.0 73150.0 10990.0 73085.0 ;
      RECT  10635.0 72432.5 11195.0 72367.5 ;
      RECT  10635.0 73777.5 11195.0 73712.5 ;
      RECT  8897.5 73050.0 8962.5 73185.0 ;
      RECT  9037.5 73322.5 9102.5 73457.5 ;
      RECT  10032.5 73287.5 9897.5 73352.5 ;
      RECT  9582.5 74905.0 9647.5 75090.0 ;
      RECT  9582.5 73745.0 9647.5 73930.0 ;
      RECT  9222.5 73862.5 9287.5 73712.5 ;
      RECT  9222.5 74747.5 9287.5 75122.5 ;
      RECT  9412.5 73862.5 9477.5 74747.5 ;
      RECT  9222.5 74747.5 9287.5 74882.5 ;
      RECT  9412.5 74747.5 9477.5 74882.5 ;
      RECT  9412.5 74747.5 9477.5 74882.5 ;
      RECT  9222.5 74747.5 9287.5 74882.5 ;
      RECT  9222.5 73862.5 9287.5 73997.5 ;
      RECT  9412.5 73862.5 9477.5 73997.5 ;
      RECT  9412.5 73862.5 9477.5 73997.5 ;
      RECT  9222.5 73862.5 9287.5 73997.5 ;
      RECT  9582.5 74837.5 9647.5 74972.5 ;
      RECT  9582.5 73862.5 9647.5 73997.5 ;
      RECT  9280.0 74305.0 9345.0 74440.0 ;
      RECT  9280.0 74305.0 9345.0 74440.0 ;
      RECT  9445.0 74340.0 9510.0 74405.0 ;
      RECT  9155.0 75057.5 9715.0 75122.5 ;
      RECT  9155.0 73712.5 9715.0 73777.5 ;
      RECT  9782.5 73907.5 9847.5 73712.5 ;
      RECT  9782.5 74747.5 9847.5 75122.5 ;
      RECT  10162.5 74747.5 10227.5 75122.5 ;
      RECT  10332.5 74905.0 10397.5 75090.0 ;
      RECT  10332.5 73745.0 10397.5 73930.0 ;
      RECT  9782.5 74747.5 9847.5 74882.5 ;
      RECT  9972.5 74747.5 10037.5 74882.5 ;
      RECT  9972.5 74747.5 10037.5 74882.5 ;
      RECT  9782.5 74747.5 9847.5 74882.5 ;
      RECT  9972.5 74747.5 10037.5 74882.5 ;
      RECT  10162.5 74747.5 10227.5 74882.5 ;
      RECT  10162.5 74747.5 10227.5 74882.5 ;
      RECT  9972.5 74747.5 10037.5 74882.5 ;
      RECT  9782.5 73907.5 9847.5 74042.5 ;
      RECT  9972.5 73907.5 10037.5 74042.5 ;
      RECT  9972.5 73907.5 10037.5 74042.5 ;
      RECT  9782.5 73907.5 9847.5 74042.5 ;
      RECT  9972.5 73907.5 10037.5 74042.5 ;
      RECT  10162.5 73907.5 10227.5 74042.5 ;
      RECT  10162.5 73907.5 10227.5 74042.5 ;
      RECT  9972.5 73907.5 10037.5 74042.5 ;
      RECT  10332.5 74837.5 10397.5 74972.5 ;
      RECT  10332.5 73862.5 10397.5 73997.5 ;
      RECT  10167.5 74137.5 10032.5 74202.5 ;
      RECT  9910.0 74352.5 9775.0 74417.5 ;
      RECT  9972.5 74747.5 10037.5 74882.5 ;
      RECT  10162.5 73907.5 10227.5 74042.5 ;
      RECT  10262.5 74352.5 10127.5 74417.5 ;
      RECT  9775.0 74352.5 9910.0 74417.5 ;
      RECT  10032.5 74137.5 10167.5 74202.5 ;
      RECT  10127.5 74352.5 10262.5 74417.5 ;
      RECT  9715.0 75057.5 10635.0 75122.5 ;
      RECT  9715.0 73712.5 10635.0 73777.5 ;
      RECT  11062.5 74905.0 11127.5 75090.0 ;
      RECT  11062.5 73745.0 11127.5 73930.0 ;
      RECT  10702.5 73862.5 10767.5 73712.5 ;
      RECT  10702.5 74747.5 10767.5 75122.5 ;
      RECT  10892.5 73862.5 10957.5 74747.5 ;
      RECT  10702.5 74747.5 10767.5 74882.5 ;
      RECT  10892.5 74747.5 10957.5 74882.5 ;
      RECT  10892.5 74747.5 10957.5 74882.5 ;
      RECT  10702.5 74747.5 10767.5 74882.5 ;
      RECT  10702.5 73862.5 10767.5 73997.5 ;
      RECT  10892.5 73862.5 10957.5 73997.5 ;
      RECT  10892.5 73862.5 10957.5 73997.5 ;
      RECT  10702.5 73862.5 10767.5 73997.5 ;
      RECT  11062.5 74837.5 11127.5 74972.5 ;
      RECT  11062.5 73862.5 11127.5 73997.5 ;
      RECT  10760.0 74305.0 10825.0 74440.0 ;
      RECT  10760.0 74305.0 10825.0 74440.0 ;
      RECT  10925.0 74340.0 10990.0 74405.0 ;
      RECT  10635.0 75057.5 11195.0 75122.5 ;
      RECT  10635.0 73712.5 11195.0 73777.5 ;
      RECT  8897.5 74305.0 8962.5 74440.0 ;
      RECT  9037.5 74032.5 9102.5 74167.5 ;
      RECT  10032.5 74137.5 9897.5 74202.5 ;
      RECT  9582.5 75275.0 9647.5 75090.0 ;
      RECT  9582.5 76435.0 9647.5 76250.0 ;
      RECT  9222.5 76317.5 9287.5 76467.5 ;
      RECT  9222.5 75432.5 9287.5 75057.5 ;
      RECT  9412.5 76317.5 9477.5 75432.5 ;
      RECT  9222.5 75432.5 9287.5 75297.5 ;
      RECT  9412.5 75432.5 9477.5 75297.5 ;
      RECT  9412.5 75432.5 9477.5 75297.5 ;
      RECT  9222.5 75432.5 9287.5 75297.5 ;
      RECT  9222.5 76317.5 9287.5 76182.5 ;
      RECT  9412.5 76317.5 9477.5 76182.5 ;
      RECT  9412.5 76317.5 9477.5 76182.5 ;
      RECT  9222.5 76317.5 9287.5 76182.5 ;
      RECT  9582.5 75342.5 9647.5 75207.5 ;
      RECT  9582.5 76317.5 9647.5 76182.5 ;
      RECT  9280.0 75875.0 9345.0 75740.0 ;
      RECT  9280.0 75875.0 9345.0 75740.0 ;
      RECT  9445.0 75840.0 9510.0 75775.0 ;
      RECT  9155.0 75122.5 9715.0 75057.5 ;
      RECT  9155.0 76467.5 9715.0 76402.5 ;
      RECT  9782.5 76272.5 9847.5 76467.5 ;
      RECT  9782.5 75432.5 9847.5 75057.5 ;
      RECT  10162.5 75432.5 10227.5 75057.5 ;
      RECT  10332.5 75275.0 10397.5 75090.0 ;
      RECT  10332.5 76435.0 10397.5 76250.0 ;
      RECT  9782.5 75432.5 9847.5 75297.5 ;
      RECT  9972.5 75432.5 10037.5 75297.5 ;
      RECT  9972.5 75432.5 10037.5 75297.5 ;
      RECT  9782.5 75432.5 9847.5 75297.5 ;
      RECT  9972.5 75432.5 10037.5 75297.5 ;
      RECT  10162.5 75432.5 10227.5 75297.5 ;
      RECT  10162.5 75432.5 10227.5 75297.5 ;
      RECT  9972.5 75432.5 10037.5 75297.5 ;
      RECT  9782.5 76272.5 9847.5 76137.5 ;
      RECT  9972.5 76272.5 10037.5 76137.5 ;
      RECT  9972.5 76272.5 10037.5 76137.5 ;
      RECT  9782.5 76272.5 9847.5 76137.5 ;
      RECT  9972.5 76272.5 10037.5 76137.5 ;
      RECT  10162.5 76272.5 10227.5 76137.5 ;
      RECT  10162.5 76272.5 10227.5 76137.5 ;
      RECT  9972.5 76272.5 10037.5 76137.5 ;
      RECT  10332.5 75342.5 10397.5 75207.5 ;
      RECT  10332.5 76317.5 10397.5 76182.5 ;
      RECT  10167.5 76042.5 10032.5 75977.5 ;
      RECT  9910.0 75827.5 9775.0 75762.5 ;
      RECT  9972.5 75432.5 10037.5 75297.5 ;
      RECT  10162.5 76272.5 10227.5 76137.5 ;
      RECT  10262.5 75827.5 10127.5 75762.5 ;
      RECT  9775.0 75827.5 9910.0 75762.5 ;
      RECT  10032.5 76042.5 10167.5 75977.5 ;
      RECT  10127.5 75827.5 10262.5 75762.5 ;
      RECT  9715.0 75122.5 10635.0 75057.5 ;
      RECT  9715.0 76467.5 10635.0 76402.5 ;
      RECT  11062.5 75275.0 11127.5 75090.0 ;
      RECT  11062.5 76435.0 11127.5 76250.0 ;
      RECT  10702.5 76317.5 10767.5 76467.5 ;
      RECT  10702.5 75432.5 10767.5 75057.5 ;
      RECT  10892.5 76317.5 10957.5 75432.5 ;
      RECT  10702.5 75432.5 10767.5 75297.5 ;
      RECT  10892.5 75432.5 10957.5 75297.5 ;
      RECT  10892.5 75432.5 10957.5 75297.5 ;
      RECT  10702.5 75432.5 10767.5 75297.5 ;
      RECT  10702.5 76317.5 10767.5 76182.5 ;
      RECT  10892.5 76317.5 10957.5 76182.5 ;
      RECT  10892.5 76317.5 10957.5 76182.5 ;
      RECT  10702.5 76317.5 10767.5 76182.5 ;
      RECT  11062.5 75342.5 11127.5 75207.5 ;
      RECT  11062.5 76317.5 11127.5 76182.5 ;
      RECT  10760.0 75875.0 10825.0 75740.0 ;
      RECT  10760.0 75875.0 10825.0 75740.0 ;
      RECT  10925.0 75840.0 10990.0 75775.0 ;
      RECT  10635.0 75122.5 11195.0 75057.5 ;
      RECT  10635.0 76467.5 11195.0 76402.5 ;
      RECT  8897.5 75740.0 8962.5 75875.0 ;
      RECT  9037.5 76012.5 9102.5 76147.5 ;
      RECT  10032.5 75977.5 9897.5 76042.5 ;
      RECT  9582.5 77595.0 9647.5 77780.0 ;
      RECT  9582.5 76435.0 9647.5 76620.0 ;
      RECT  9222.5 76552.5 9287.5 76402.5 ;
      RECT  9222.5 77437.5 9287.5 77812.5 ;
      RECT  9412.5 76552.5 9477.5 77437.5 ;
      RECT  9222.5 77437.5 9287.5 77572.5 ;
      RECT  9412.5 77437.5 9477.5 77572.5 ;
      RECT  9412.5 77437.5 9477.5 77572.5 ;
      RECT  9222.5 77437.5 9287.5 77572.5 ;
      RECT  9222.5 76552.5 9287.5 76687.5 ;
      RECT  9412.5 76552.5 9477.5 76687.5 ;
      RECT  9412.5 76552.5 9477.5 76687.5 ;
      RECT  9222.5 76552.5 9287.5 76687.5 ;
      RECT  9582.5 77527.5 9647.5 77662.5 ;
      RECT  9582.5 76552.5 9647.5 76687.5 ;
      RECT  9280.0 76995.0 9345.0 77130.0 ;
      RECT  9280.0 76995.0 9345.0 77130.0 ;
      RECT  9445.0 77030.0 9510.0 77095.0 ;
      RECT  9155.0 77747.5 9715.0 77812.5 ;
      RECT  9155.0 76402.5 9715.0 76467.5 ;
      RECT  9782.5 76597.5 9847.5 76402.5 ;
      RECT  9782.5 77437.5 9847.5 77812.5 ;
      RECT  10162.5 77437.5 10227.5 77812.5 ;
      RECT  10332.5 77595.0 10397.5 77780.0 ;
      RECT  10332.5 76435.0 10397.5 76620.0 ;
      RECT  9782.5 77437.5 9847.5 77572.5 ;
      RECT  9972.5 77437.5 10037.5 77572.5 ;
      RECT  9972.5 77437.5 10037.5 77572.5 ;
      RECT  9782.5 77437.5 9847.5 77572.5 ;
      RECT  9972.5 77437.5 10037.5 77572.5 ;
      RECT  10162.5 77437.5 10227.5 77572.5 ;
      RECT  10162.5 77437.5 10227.5 77572.5 ;
      RECT  9972.5 77437.5 10037.5 77572.5 ;
      RECT  9782.5 76597.5 9847.5 76732.5 ;
      RECT  9972.5 76597.5 10037.5 76732.5 ;
      RECT  9972.5 76597.5 10037.5 76732.5 ;
      RECT  9782.5 76597.5 9847.5 76732.5 ;
      RECT  9972.5 76597.5 10037.5 76732.5 ;
      RECT  10162.5 76597.5 10227.5 76732.5 ;
      RECT  10162.5 76597.5 10227.5 76732.5 ;
      RECT  9972.5 76597.5 10037.5 76732.5 ;
      RECT  10332.5 77527.5 10397.5 77662.5 ;
      RECT  10332.5 76552.5 10397.5 76687.5 ;
      RECT  10167.5 76827.5 10032.5 76892.5 ;
      RECT  9910.0 77042.5 9775.0 77107.5 ;
      RECT  9972.5 77437.5 10037.5 77572.5 ;
      RECT  10162.5 76597.5 10227.5 76732.5 ;
      RECT  10262.5 77042.5 10127.5 77107.5 ;
      RECT  9775.0 77042.5 9910.0 77107.5 ;
      RECT  10032.5 76827.5 10167.5 76892.5 ;
      RECT  10127.5 77042.5 10262.5 77107.5 ;
      RECT  9715.0 77747.5 10635.0 77812.5 ;
      RECT  9715.0 76402.5 10635.0 76467.5 ;
      RECT  11062.5 77595.0 11127.5 77780.0 ;
      RECT  11062.5 76435.0 11127.5 76620.0 ;
      RECT  10702.5 76552.5 10767.5 76402.5 ;
      RECT  10702.5 77437.5 10767.5 77812.5 ;
      RECT  10892.5 76552.5 10957.5 77437.5 ;
      RECT  10702.5 77437.5 10767.5 77572.5 ;
      RECT  10892.5 77437.5 10957.5 77572.5 ;
      RECT  10892.5 77437.5 10957.5 77572.5 ;
      RECT  10702.5 77437.5 10767.5 77572.5 ;
      RECT  10702.5 76552.5 10767.5 76687.5 ;
      RECT  10892.5 76552.5 10957.5 76687.5 ;
      RECT  10892.5 76552.5 10957.5 76687.5 ;
      RECT  10702.5 76552.5 10767.5 76687.5 ;
      RECT  11062.5 77527.5 11127.5 77662.5 ;
      RECT  11062.5 76552.5 11127.5 76687.5 ;
      RECT  10760.0 76995.0 10825.0 77130.0 ;
      RECT  10760.0 76995.0 10825.0 77130.0 ;
      RECT  10925.0 77030.0 10990.0 77095.0 ;
      RECT  10635.0 77747.5 11195.0 77812.5 ;
      RECT  10635.0 76402.5 11195.0 76467.5 ;
      RECT  8897.5 76995.0 8962.5 77130.0 ;
      RECT  9037.5 76722.5 9102.5 76857.5 ;
      RECT  10032.5 76827.5 9897.5 76892.5 ;
      RECT  9582.5 77965.0 9647.5 77780.0 ;
      RECT  9582.5 79125.0 9647.5 78940.0 ;
      RECT  9222.5 79007.5 9287.5 79157.5 ;
      RECT  9222.5 78122.5 9287.5 77747.5 ;
      RECT  9412.5 79007.5 9477.5 78122.5 ;
      RECT  9222.5 78122.5 9287.5 77987.5 ;
      RECT  9412.5 78122.5 9477.5 77987.5 ;
      RECT  9412.5 78122.5 9477.5 77987.5 ;
      RECT  9222.5 78122.5 9287.5 77987.5 ;
      RECT  9222.5 79007.5 9287.5 78872.5 ;
      RECT  9412.5 79007.5 9477.5 78872.5 ;
      RECT  9412.5 79007.5 9477.5 78872.5 ;
      RECT  9222.5 79007.5 9287.5 78872.5 ;
      RECT  9582.5 78032.5 9647.5 77897.5 ;
      RECT  9582.5 79007.5 9647.5 78872.5 ;
      RECT  9280.0 78565.0 9345.0 78430.0 ;
      RECT  9280.0 78565.0 9345.0 78430.0 ;
      RECT  9445.0 78530.0 9510.0 78465.0 ;
      RECT  9155.0 77812.5 9715.0 77747.5 ;
      RECT  9155.0 79157.5 9715.0 79092.5 ;
      RECT  9782.5 78962.5 9847.5 79157.5 ;
      RECT  9782.5 78122.5 9847.5 77747.5 ;
      RECT  10162.5 78122.5 10227.5 77747.5 ;
      RECT  10332.5 77965.0 10397.5 77780.0 ;
      RECT  10332.5 79125.0 10397.5 78940.0 ;
      RECT  9782.5 78122.5 9847.5 77987.5 ;
      RECT  9972.5 78122.5 10037.5 77987.5 ;
      RECT  9972.5 78122.5 10037.5 77987.5 ;
      RECT  9782.5 78122.5 9847.5 77987.5 ;
      RECT  9972.5 78122.5 10037.5 77987.5 ;
      RECT  10162.5 78122.5 10227.5 77987.5 ;
      RECT  10162.5 78122.5 10227.5 77987.5 ;
      RECT  9972.5 78122.5 10037.5 77987.5 ;
      RECT  9782.5 78962.5 9847.5 78827.5 ;
      RECT  9972.5 78962.5 10037.5 78827.5 ;
      RECT  9972.5 78962.5 10037.5 78827.5 ;
      RECT  9782.5 78962.5 9847.5 78827.5 ;
      RECT  9972.5 78962.5 10037.5 78827.5 ;
      RECT  10162.5 78962.5 10227.5 78827.5 ;
      RECT  10162.5 78962.5 10227.5 78827.5 ;
      RECT  9972.5 78962.5 10037.5 78827.5 ;
      RECT  10332.5 78032.5 10397.5 77897.5 ;
      RECT  10332.5 79007.5 10397.5 78872.5 ;
      RECT  10167.5 78732.5 10032.5 78667.5 ;
      RECT  9910.0 78517.5 9775.0 78452.5 ;
      RECT  9972.5 78122.5 10037.5 77987.5 ;
      RECT  10162.5 78962.5 10227.5 78827.5 ;
      RECT  10262.5 78517.5 10127.5 78452.5 ;
      RECT  9775.0 78517.5 9910.0 78452.5 ;
      RECT  10032.5 78732.5 10167.5 78667.5 ;
      RECT  10127.5 78517.5 10262.5 78452.5 ;
      RECT  9715.0 77812.5 10635.0 77747.5 ;
      RECT  9715.0 79157.5 10635.0 79092.5 ;
      RECT  11062.5 77965.0 11127.5 77780.0 ;
      RECT  11062.5 79125.0 11127.5 78940.0 ;
      RECT  10702.5 79007.5 10767.5 79157.5 ;
      RECT  10702.5 78122.5 10767.5 77747.5 ;
      RECT  10892.5 79007.5 10957.5 78122.5 ;
      RECT  10702.5 78122.5 10767.5 77987.5 ;
      RECT  10892.5 78122.5 10957.5 77987.5 ;
      RECT  10892.5 78122.5 10957.5 77987.5 ;
      RECT  10702.5 78122.5 10767.5 77987.5 ;
      RECT  10702.5 79007.5 10767.5 78872.5 ;
      RECT  10892.5 79007.5 10957.5 78872.5 ;
      RECT  10892.5 79007.5 10957.5 78872.5 ;
      RECT  10702.5 79007.5 10767.5 78872.5 ;
      RECT  11062.5 78032.5 11127.5 77897.5 ;
      RECT  11062.5 79007.5 11127.5 78872.5 ;
      RECT  10760.0 78565.0 10825.0 78430.0 ;
      RECT  10760.0 78565.0 10825.0 78430.0 ;
      RECT  10925.0 78530.0 10990.0 78465.0 ;
      RECT  10635.0 77812.5 11195.0 77747.5 ;
      RECT  10635.0 79157.5 11195.0 79092.5 ;
      RECT  8897.5 78430.0 8962.5 78565.0 ;
      RECT  9037.5 78702.5 9102.5 78837.5 ;
      RECT  10032.5 78667.5 9897.5 78732.5 ;
      RECT  9582.5 80285.0 9647.5 80470.0 ;
      RECT  9582.5 79125.0 9647.5 79310.0 ;
      RECT  9222.5 79242.5 9287.5 79092.5 ;
      RECT  9222.5 80127.5 9287.5 80502.5 ;
      RECT  9412.5 79242.5 9477.5 80127.5 ;
      RECT  9222.5 80127.5 9287.5 80262.5 ;
      RECT  9412.5 80127.5 9477.5 80262.5 ;
      RECT  9412.5 80127.5 9477.5 80262.5 ;
      RECT  9222.5 80127.5 9287.5 80262.5 ;
      RECT  9222.5 79242.5 9287.5 79377.5 ;
      RECT  9412.5 79242.5 9477.5 79377.5 ;
      RECT  9412.5 79242.5 9477.5 79377.5 ;
      RECT  9222.5 79242.5 9287.5 79377.5 ;
      RECT  9582.5 80217.5 9647.5 80352.5 ;
      RECT  9582.5 79242.5 9647.5 79377.5 ;
      RECT  9280.0 79685.0 9345.0 79820.0 ;
      RECT  9280.0 79685.0 9345.0 79820.0 ;
      RECT  9445.0 79720.0 9510.0 79785.0 ;
      RECT  9155.0 80437.5 9715.0 80502.5 ;
      RECT  9155.0 79092.5 9715.0 79157.5 ;
      RECT  9782.5 79287.5 9847.5 79092.5 ;
      RECT  9782.5 80127.5 9847.5 80502.5 ;
      RECT  10162.5 80127.5 10227.5 80502.5 ;
      RECT  10332.5 80285.0 10397.5 80470.0 ;
      RECT  10332.5 79125.0 10397.5 79310.0 ;
      RECT  9782.5 80127.5 9847.5 80262.5 ;
      RECT  9972.5 80127.5 10037.5 80262.5 ;
      RECT  9972.5 80127.5 10037.5 80262.5 ;
      RECT  9782.5 80127.5 9847.5 80262.5 ;
      RECT  9972.5 80127.5 10037.5 80262.5 ;
      RECT  10162.5 80127.5 10227.5 80262.5 ;
      RECT  10162.5 80127.5 10227.5 80262.5 ;
      RECT  9972.5 80127.5 10037.5 80262.5 ;
      RECT  9782.5 79287.5 9847.5 79422.5 ;
      RECT  9972.5 79287.5 10037.5 79422.5 ;
      RECT  9972.5 79287.5 10037.5 79422.5 ;
      RECT  9782.5 79287.5 9847.5 79422.5 ;
      RECT  9972.5 79287.5 10037.5 79422.5 ;
      RECT  10162.5 79287.5 10227.5 79422.5 ;
      RECT  10162.5 79287.5 10227.5 79422.5 ;
      RECT  9972.5 79287.5 10037.5 79422.5 ;
      RECT  10332.5 80217.5 10397.5 80352.5 ;
      RECT  10332.5 79242.5 10397.5 79377.5 ;
      RECT  10167.5 79517.5 10032.5 79582.5 ;
      RECT  9910.0 79732.5 9775.0 79797.5 ;
      RECT  9972.5 80127.5 10037.5 80262.5 ;
      RECT  10162.5 79287.5 10227.5 79422.5 ;
      RECT  10262.5 79732.5 10127.5 79797.5 ;
      RECT  9775.0 79732.5 9910.0 79797.5 ;
      RECT  10032.5 79517.5 10167.5 79582.5 ;
      RECT  10127.5 79732.5 10262.5 79797.5 ;
      RECT  9715.0 80437.5 10635.0 80502.5 ;
      RECT  9715.0 79092.5 10635.0 79157.5 ;
      RECT  11062.5 80285.0 11127.5 80470.0 ;
      RECT  11062.5 79125.0 11127.5 79310.0 ;
      RECT  10702.5 79242.5 10767.5 79092.5 ;
      RECT  10702.5 80127.5 10767.5 80502.5 ;
      RECT  10892.5 79242.5 10957.5 80127.5 ;
      RECT  10702.5 80127.5 10767.5 80262.5 ;
      RECT  10892.5 80127.5 10957.5 80262.5 ;
      RECT  10892.5 80127.5 10957.5 80262.5 ;
      RECT  10702.5 80127.5 10767.5 80262.5 ;
      RECT  10702.5 79242.5 10767.5 79377.5 ;
      RECT  10892.5 79242.5 10957.5 79377.5 ;
      RECT  10892.5 79242.5 10957.5 79377.5 ;
      RECT  10702.5 79242.5 10767.5 79377.5 ;
      RECT  11062.5 80217.5 11127.5 80352.5 ;
      RECT  11062.5 79242.5 11127.5 79377.5 ;
      RECT  10760.0 79685.0 10825.0 79820.0 ;
      RECT  10760.0 79685.0 10825.0 79820.0 ;
      RECT  10925.0 79720.0 10990.0 79785.0 ;
      RECT  10635.0 80437.5 11195.0 80502.5 ;
      RECT  10635.0 79092.5 11195.0 79157.5 ;
      RECT  8897.5 79685.0 8962.5 79820.0 ;
      RECT  9037.5 79412.5 9102.5 79547.5 ;
      RECT  10032.5 79517.5 9897.5 79582.5 ;
      RECT  9582.5 80655.0 9647.5 80470.0 ;
      RECT  9582.5 81815.0 9647.5 81630.0 ;
      RECT  9222.5 81697.5 9287.5 81847.5 ;
      RECT  9222.5 80812.5 9287.5 80437.5 ;
      RECT  9412.5 81697.5 9477.5 80812.5 ;
      RECT  9222.5 80812.5 9287.5 80677.5 ;
      RECT  9412.5 80812.5 9477.5 80677.5 ;
      RECT  9412.5 80812.5 9477.5 80677.5 ;
      RECT  9222.5 80812.5 9287.5 80677.5 ;
      RECT  9222.5 81697.5 9287.5 81562.5 ;
      RECT  9412.5 81697.5 9477.5 81562.5 ;
      RECT  9412.5 81697.5 9477.5 81562.5 ;
      RECT  9222.5 81697.5 9287.5 81562.5 ;
      RECT  9582.5 80722.5 9647.5 80587.5 ;
      RECT  9582.5 81697.5 9647.5 81562.5 ;
      RECT  9280.0 81255.0 9345.0 81120.0 ;
      RECT  9280.0 81255.0 9345.0 81120.0 ;
      RECT  9445.0 81220.0 9510.0 81155.0 ;
      RECT  9155.0 80502.5 9715.0 80437.5 ;
      RECT  9155.0 81847.5 9715.0 81782.5 ;
      RECT  9782.5 81652.5 9847.5 81847.5 ;
      RECT  9782.5 80812.5 9847.5 80437.5 ;
      RECT  10162.5 80812.5 10227.5 80437.5 ;
      RECT  10332.5 80655.0 10397.5 80470.0 ;
      RECT  10332.5 81815.0 10397.5 81630.0 ;
      RECT  9782.5 80812.5 9847.5 80677.5 ;
      RECT  9972.5 80812.5 10037.5 80677.5 ;
      RECT  9972.5 80812.5 10037.5 80677.5 ;
      RECT  9782.5 80812.5 9847.5 80677.5 ;
      RECT  9972.5 80812.5 10037.5 80677.5 ;
      RECT  10162.5 80812.5 10227.5 80677.5 ;
      RECT  10162.5 80812.5 10227.5 80677.5 ;
      RECT  9972.5 80812.5 10037.5 80677.5 ;
      RECT  9782.5 81652.5 9847.5 81517.5 ;
      RECT  9972.5 81652.5 10037.5 81517.5 ;
      RECT  9972.5 81652.5 10037.5 81517.5 ;
      RECT  9782.5 81652.5 9847.5 81517.5 ;
      RECT  9972.5 81652.5 10037.5 81517.5 ;
      RECT  10162.5 81652.5 10227.5 81517.5 ;
      RECT  10162.5 81652.5 10227.5 81517.5 ;
      RECT  9972.5 81652.5 10037.5 81517.5 ;
      RECT  10332.5 80722.5 10397.5 80587.5 ;
      RECT  10332.5 81697.5 10397.5 81562.5 ;
      RECT  10167.5 81422.5 10032.5 81357.5 ;
      RECT  9910.0 81207.5 9775.0 81142.5 ;
      RECT  9972.5 80812.5 10037.5 80677.5 ;
      RECT  10162.5 81652.5 10227.5 81517.5 ;
      RECT  10262.5 81207.5 10127.5 81142.5 ;
      RECT  9775.0 81207.5 9910.0 81142.5 ;
      RECT  10032.5 81422.5 10167.5 81357.5 ;
      RECT  10127.5 81207.5 10262.5 81142.5 ;
      RECT  9715.0 80502.5 10635.0 80437.5 ;
      RECT  9715.0 81847.5 10635.0 81782.5 ;
      RECT  11062.5 80655.0 11127.5 80470.0 ;
      RECT  11062.5 81815.0 11127.5 81630.0 ;
      RECT  10702.5 81697.5 10767.5 81847.5 ;
      RECT  10702.5 80812.5 10767.5 80437.5 ;
      RECT  10892.5 81697.5 10957.5 80812.5 ;
      RECT  10702.5 80812.5 10767.5 80677.5 ;
      RECT  10892.5 80812.5 10957.5 80677.5 ;
      RECT  10892.5 80812.5 10957.5 80677.5 ;
      RECT  10702.5 80812.5 10767.5 80677.5 ;
      RECT  10702.5 81697.5 10767.5 81562.5 ;
      RECT  10892.5 81697.5 10957.5 81562.5 ;
      RECT  10892.5 81697.5 10957.5 81562.5 ;
      RECT  10702.5 81697.5 10767.5 81562.5 ;
      RECT  11062.5 80722.5 11127.5 80587.5 ;
      RECT  11062.5 81697.5 11127.5 81562.5 ;
      RECT  10760.0 81255.0 10825.0 81120.0 ;
      RECT  10760.0 81255.0 10825.0 81120.0 ;
      RECT  10925.0 81220.0 10990.0 81155.0 ;
      RECT  10635.0 80502.5 11195.0 80437.5 ;
      RECT  10635.0 81847.5 11195.0 81782.5 ;
      RECT  8897.5 81120.0 8962.5 81255.0 ;
      RECT  9037.5 81392.5 9102.5 81527.5 ;
      RECT  10032.5 81357.5 9897.5 81422.5 ;
      RECT  9582.5 82975.0 9647.5 83160.0 ;
      RECT  9582.5 81815.0 9647.5 82000.0 ;
      RECT  9222.5 81932.5 9287.5 81782.5 ;
      RECT  9222.5 82817.5 9287.5 83192.5 ;
      RECT  9412.5 81932.5 9477.5 82817.5 ;
      RECT  9222.5 82817.5 9287.5 82952.5 ;
      RECT  9412.5 82817.5 9477.5 82952.5 ;
      RECT  9412.5 82817.5 9477.5 82952.5 ;
      RECT  9222.5 82817.5 9287.5 82952.5 ;
      RECT  9222.5 81932.5 9287.5 82067.5 ;
      RECT  9412.5 81932.5 9477.5 82067.5 ;
      RECT  9412.5 81932.5 9477.5 82067.5 ;
      RECT  9222.5 81932.5 9287.5 82067.5 ;
      RECT  9582.5 82907.5 9647.5 83042.5 ;
      RECT  9582.5 81932.5 9647.5 82067.5 ;
      RECT  9280.0 82375.0 9345.0 82510.0 ;
      RECT  9280.0 82375.0 9345.0 82510.0 ;
      RECT  9445.0 82410.0 9510.0 82475.0 ;
      RECT  9155.0 83127.5 9715.0 83192.5 ;
      RECT  9155.0 81782.5 9715.0 81847.5 ;
      RECT  9782.5 81977.5 9847.5 81782.5 ;
      RECT  9782.5 82817.5 9847.5 83192.5 ;
      RECT  10162.5 82817.5 10227.5 83192.5 ;
      RECT  10332.5 82975.0 10397.5 83160.0 ;
      RECT  10332.5 81815.0 10397.5 82000.0 ;
      RECT  9782.5 82817.5 9847.5 82952.5 ;
      RECT  9972.5 82817.5 10037.5 82952.5 ;
      RECT  9972.5 82817.5 10037.5 82952.5 ;
      RECT  9782.5 82817.5 9847.5 82952.5 ;
      RECT  9972.5 82817.5 10037.5 82952.5 ;
      RECT  10162.5 82817.5 10227.5 82952.5 ;
      RECT  10162.5 82817.5 10227.5 82952.5 ;
      RECT  9972.5 82817.5 10037.5 82952.5 ;
      RECT  9782.5 81977.5 9847.5 82112.5 ;
      RECT  9972.5 81977.5 10037.5 82112.5 ;
      RECT  9972.5 81977.5 10037.5 82112.5 ;
      RECT  9782.5 81977.5 9847.5 82112.5 ;
      RECT  9972.5 81977.5 10037.5 82112.5 ;
      RECT  10162.5 81977.5 10227.5 82112.5 ;
      RECT  10162.5 81977.5 10227.5 82112.5 ;
      RECT  9972.5 81977.5 10037.5 82112.5 ;
      RECT  10332.5 82907.5 10397.5 83042.5 ;
      RECT  10332.5 81932.5 10397.5 82067.5 ;
      RECT  10167.5 82207.5 10032.5 82272.5 ;
      RECT  9910.0 82422.5 9775.0 82487.5 ;
      RECT  9972.5 82817.5 10037.5 82952.5 ;
      RECT  10162.5 81977.5 10227.5 82112.5 ;
      RECT  10262.5 82422.5 10127.5 82487.5 ;
      RECT  9775.0 82422.5 9910.0 82487.5 ;
      RECT  10032.5 82207.5 10167.5 82272.5 ;
      RECT  10127.5 82422.5 10262.5 82487.5 ;
      RECT  9715.0 83127.5 10635.0 83192.5 ;
      RECT  9715.0 81782.5 10635.0 81847.5 ;
      RECT  11062.5 82975.0 11127.5 83160.0 ;
      RECT  11062.5 81815.0 11127.5 82000.0 ;
      RECT  10702.5 81932.5 10767.5 81782.5 ;
      RECT  10702.5 82817.5 10767.5 83192.5 ;
      RECT  10892.5 81932.5 10957.5 82817.5 ;
      RECT  10702.5 82817.5 10767.5 82952.5 ;
      RECT  10892.5 82817.5 10957.5 82952.5 ;
      RECT  10892.5 82817.5 10957.5 82952.5 ;
      RECT  10702.5 82817.5 10767.5 82952.5 ;
      RECT  10702.5 81932.5 10767.5 82067.5 ;
      RECT  10892.5 81932.5 10957.5 82067.5 ;
      RECT  10892.5 81932.5 10957.5 82067.5 ;
      RECT  10702.5 81932.5 10767.5 82067.5 ;
      RECT  11062.5 82907.5 11127.5 83042.5 ;
      RECT  11062.5 81932.5 11127.5 82067.5 ;
      RECT  10760.0 82375.0 10825.0 82510.0 ;
      RECT  10760.0 82375.0 10825.0 82510.0 ;
      RECT  10925.0 82410.0 10990.0 82475.0 ;
      RECT  10635.0 83127.5 11195.0 83192.5 ;
      RECT  10635.0 81782.5 11195.0 81847.5 ;
      RECT  8897.5 82375.0 8962.5 82510.0 ;
      RECT  9037.5 82102.5 9102.5 82237.5 ;
      RECT  10032.5 82207.5 9897.5 82272.5 ;
      RECT  9582.5 83345.0 9647.5 83160.0 ;
      RECT  9582.5 84505.0 9647.5 84320.0 ;
      RECT  9222.5 84387.5 9287.5 84537.5 ;
      RECT  9222.5 83502.5 9287.5 83127.5 ;
      RECT  9412.5 84387.5 9477.5 83502.5 ;
      RECT  9222.5 83502.5 9287.5 83367.5 ;
      RECT  9412.5 83502.5 9477.5 83367.5 ;
      RECT  9412.5 83502.5 9477.5 83367.5 ;
      RECT  9222.5 83502.5 9287.5 83367.5 ;
      RECT  9222.5 84387.5 9287.5 84252.5 ;
      RECT  9412.5 84387.5 9477.5 84252.5 ;
      RECT  9412.5 84387.5 9477.5 84252.5 ;
      RECT  9222.5 84387.5 9287.5 84252.5 ;
      RECT  9582.5 83412.5 9647.5 83277.5 ;
      RECT  9582.5 84387.5 9647.5 84252.5 ;
      RECT  9280.0 83945.0 9345.0 83810.0 ;
      RECT  9280.0 83945.0 9345.0 83810.0 ;
      RECT  9445.0 83910.0 9510.0 83845.0 ;
      RECT  9155.0 83192.5 9715.0 83127.5 ;
      RECT  9155.0 84537.5 9715.0 84472.5 ;
      RECT  9782.5 84342.5 9847.5 84537.5 ;
      RECT  9782.5 83502.5 9847.5 83127.5 ;
      RECT  10162.5 83502.5 10227.5 83127.5 ;
      RECT  10332.5 83345.0 10397.5 83160.0 ;
      RECT  10332.5 84505.0 10397.5 84320.0 ;
      RECT  9782.5 83502.5 9847.5 83367.5 ;
      RECT  9972.5 83502.5 10037.5 83367.5 ;
      RECT  9972.5 83502.5 10037.5 83367.5 ;
      RECT  9782.5 83502.5 9847.5 83367.5 ;
      RECT  9972.5 83502.5 10037.5 83367.5 ;
      RECT  10162.5 83502.5 10227.5 83367.5 ;
      RECT  10162.5 83502.5 10227.5 83367.5 ;
      RECT  9972.5 83502.5 10037.5 83367.5 ;
      RECT  9782.5 84342.5 9847.5 84207.5 ;
      RECT  9972.5 84342.5 10037.5 84207.5 ;
      RECT  9972.5 84342.5 10037.5 84207.5 ;
      RECT  9782.5 84342.5 9847.5 84207.5 ;
      RECT  9972.5 84342.5 10037.5 84207.5 ;
      RECT  10162.5 84342.5 10227.5 84207.5 ;
      RECT  10162.5 84342.5 10227.5 84207.5 ;
      RECT  9972.5 84342.5 10037.5 84207.5 ;
      RECT  10332.5 83412.5 10397.5 83277.5 ;
      RECT  10332.5 84387.5 10397.5 84252.5 ;
      RECT  10167.5 84112.5 10032.5 84047.5 ;
      RECT  9910.0 83897.5 9775.0 83832.5 ;
      RECT  9972.5 83502.5 10037.5 83367.5 ;
      RECT  10162.5 84342.5 10227.5 84207.5 ;
      RECT  10262.5 83897.5 10127.5 83832.5 ;
      RECT  9775.0 83897.5 9910.0 83832.5 ;
      RECT  10032.5 84112.5 10167.5 84047.5 ;
      RECT  10127.5 83897.5 10262.5 83832.5 ;
      RECT  9715.0 83192.5 10635.0 83127.5 ;
      RECT  9715.0 84537.5 10635.0 84472.5 ;
      RECT  11062.5 83345.0 11127.5 83160.0 ;
      RECT  11062.5 84505.0 11127.5 84320.0 ;
      RECT  10702.5 84387.5 10767.5 84537.5 ;
      RECT  10702.5 83502.5 10767.5 83127.5 ;
      RECT  10892.5 84387.5 10957.5 83502.5 ;
      RECT  10702.5 83502.5 10767.5 83367.5 ;
      RECT  10892.5 83502.5 10957.5 83367.5 ;
      RECT  10892.5 83502.5 10957.5 83367.5 ;
      RECT  10702.5 83502.5 10767.5 83367.5 ;
      RECT  10702.5 84387.5 10767.5 84252.5 ;
      RECT  10892.5 84387.5 10957.5 84252.5 ;
      RECT  10892.5 84387.5 10957.5 84252.5 ;
      RECT  10702.5 84387.5 10767.5 84252.5 ;
      RECT  11062.5 83412.5 11127.5 83277.5 ;
      RECT  11062.5 84387.5 11127.5 84252.5 ;
      RECT  10760.0 83945.0 10825.0 83810.0 ;
      RECT  10760.0 83945.0 10825.0 83810.0 ;
      RECT  10925.0 83910.0 10990.0 83845.0 ;
      RECT  10635.0 83192.5 11195.0 83127.5 ;
      RECT  10635.0 84537.5 11195.0 84472.5 ;
      RECT  8897.5 83810.0 8962.5 83945.0 ;
      RECT  9037.5 84082.5 9102.5 84217.5 ;
      RECT  10032.5 84047.5 9897.5 84112.5 ;
      RECT  9582.5 85665.0 9647.5 85850.0 ;
      RECT  9582.5 84505.0 9647.5 84690.0 ;
      RECT  9222.5 84622.5 9287.5 84472.5 ;
      RECT  9222.5 85507.5 9287.5 85882.5 ;
      RECT  9412.5 84622.5 9477.5 85507.5 ;
      RECT  9222.5 85507.5 9287.5 85642.5 ;
      RECT  9412.5 85507.5 9477.5 85642.5 ;
      RECT  9412.5 85507.5 9477.5 85642.5 ;
      RECT  9222.5 85507.5 9287.5 85642.5 ;
      RECT  9222.5 84622.5 9287.5 84757.5 ;
      RECT  9412.5 84622.5 9477.5 84757.5 ;
      RECT  9412.5 84622.5 9477.5 84757.5 ;
      RECT  9222.5 84622.5 9287.5 84757.5 ;
      RECT  9582.5 85597.5 9647.5 85732.5 ;
      RECT  9582.5 84622.5 9647.5 84757.5 ;
      RECT  9280.0 85065.0 9345.0 85200.0 ;
      RECT  9280.0 85065.0 9345.0 85200.0 ;
      RECT  9445.0 85100.0 9510.0 85165.0 ;
      RECT  9155.0 85817.5 9715.0 85882.5 ;
      RECT  9155.0 84472.5 9715.0 84537.5 ;
      RECT  9782.5 84667.5 9847.5 84472.5 ;
      RECT  9782.5 85507.5 9847.5 85882.5 ;
      RECT  10162.5 85507.5 10227.5 85882.5 ;
      RECT  10332.5 85665.0 10397.5 85850.0 ;
      RECT  10332.5 84505.0 10397.5 84690.0 ;
      RECT  9782.5 85507.5 9847.5 85642.5 ;
      RECT  9972.5 85507.5 10037.5 85642.5 ;
      RECT  9972.5 85507.5 10037.5 85642.5 ;
      RECT  9782.5 85507.5 9847.5 85642.5 ;
      RECT  9972.5 85507.5 10037.5 85642.5 ;
      RECT  10162.5 85507.5 10227.5 85642.5 ;
      RECT  10162.5 85507.5 10227.5 85642.5 ;
      RECT  9972.5 85507.5 10037.5 85642.5 ;
      RECT  9782.5 84667.5 9847.5 84802.5 ;
      RECT  9972.5 84667.5 10037.5 84802.5 ;
      RECT  9972.5 84667.5 10037.5 84802.5 ;
      RECT  9782.5 84667.5 9847.5 84802.5 ;
      RECT  9972.5 84667.5 10037.5 84802.5 ;
      RECT  10162.5 84667.5 10227.5 84802.5 ;
      RECT  10162.5 84667.5 10227.5 84802.5 ;
      RECT  9972.5 84667.5 10037.5 84802.5 ;
      RECT  10332.5 85597.5 10397.5 85732.5 ;
      RECT  10332.5 84622.5 10397.5 84757.5 ;
      RECT  10167.5 84897.5 10032.5 84962.5 ;
      RECT  9910.0 85112.5 9775.0 85177.5 ;
      RECT  9972.5 85507.5 10037.5 85642.5 ;
      RECT  10162.5 84667.5 10227.5 84802.5 ;
      RECT  10262.5 85112.5 10127.5 85177.5 ;
      RECT  9775.0 85112.5 9910.0 85177.5 ;
      RECT  10032.5 84897.5 10167.5 84962.5 ;
      RECT  10127.5 85112.5 10262.5 85177.5 ;
      RECT  9715.0 85817.5 10635.0 85882.5 ;
      RECT  9715.0 84472.5 10635.0 84537.5 ;
      RECT  11062.5 85665.0 11127.5 85850.0 ;
      RECT  11062.5 84505.0 11127.5 84690.0 ;
      RECT  10702.5 84622.5 10767.5 84472.5 ;
      RECT  10702.5 85507.5 10767.5 85882.5 ;
      RECT  10892.5 84622.5 10957.5 85507.5 ;
      RECT  10702.5 85507.5 10767.5 85642.5 ;
      RECT  10892.5 85507.5 10957.5 85642.5 ;
      RECT  10892.5 85507.5 10957.5 85642.5 ;
      RECT  10702.5 85507.5 10767.5 85642.5 ;
      RECT  10702.5 84622.5 10767.5 84757.5 ;
      RECT  10892.5 84622.5 10957.5 84757.5 ;
      RECT  10892.5 84622.5 10957.5 84757.5 ;
      RECT  10702.5 84622.5 10767.5 84757.5 ;
      RECT  11062.5 85597.5 11127.5 85732.5 ;
      RECT  11062.5 84622.5 11127.5 84757.5 ;
      RECT  10760.0 85065.0 10825.0 85200.0 ;
      RECT  10760.0 85065.0 10825.0 85200.0 ;
      RECT  10925.0 85100.0 10990.0 85165.0 ;
      RECT  10635.0 85817.5 11195.0 85882.5 ;
      RECT  10635.0 84472.5 11195.0 84537.5 ;
      RECT  8897.5 85065.0 8962.5 85200.0 ;
      RECT  9037.5 84792.5 9102.5 84927.5 ;
      RECT  10032.5 84897.5 9897.5 84962.5 ;
      RECT  9582.5 86035.0 9647.5 85850.0 ;
      RECT  9582.5 87195.0 9647.5 87010.0 ;
      RECT  9222.5 87077.5 9287.5 87227.5 ;
      RECT  9222.5 86192.5 9287.5 85817.5 ;
      RECT  9412.5 87077.5 9477.5 86192.5 ;
      RECT  9222.5 86192.5 9287.5 86057.5 ;
      RECT  9412.5 86192.5 9477.5 86057.5 ;
      RECT  9412.5 86192.5 9477.5 86057.5 ;
      RECT  9222.5 86192.5 9287.5 86057.5 ;
      RECT  9222.5 87077.5 9287.5 86942.5 ;
      RECT  9412.5 87077.5 9477.5 86942.5 ;
      RECT  9412.5 87077.5 9477.5 86942.5 ;
      RECT  9222.5 87077.5 9287.5 86942.5 ;
      RECT  9582.5 86102.5 9647.5 85967.5 ;
      RECT  9582.5 87077.5 9647.5 86942.5 ;
      RECT  9280.0 86635.0 9345.0 86500.0 ;
      RECT  9280.0 86635.0 9345.0 86500.0 ;
      RECT  9445.0 86600.0 9510.0 86535.0 ;
      RECT  9155.0 85882.5 9715.0 85817.5 ;
      RECT  9155.0 87227.5 9715.0 87162.5 ;
      RECT  9782.5 87032.5 9847.5 87227.5 ;
      RECT  9782.5 86192.5 9847.5 85817.5 ;
      RECT  10162.5 86192.5 10227.5 85817.5 ;
      RECT  10332.5 86035.0 10397.5 85850.0 ;
      RECT  10332.5 87195.0 10397.5 87010.0 ;
      RECT  9782.5 86192.5 9847.5 86057.5 ;
      RECT  9972.5 86192.5 10037.5 86057.5 ;
      RECT  9972.5 86192.5 10037.5 86057.5 ;
      RECT  9782.5 86192.5 9847.5 86057.5 ;
      RECT  9972.5 86192.5 10037.5 86057.5 ;
      RECT  10162.5 86192.5 10227.5 86057.5 ;
      RECT  10162.5 86192.5 10227.5 86057.5 ;
      RECT  9972.5 86192.5 10037.5 86057.5 ;
      RECT  9782.5 87032.5 9847.5 86897.5 ;
      RECT  9972.5 87032.5 10037.5 86897.5 ;
      RECT  9972.5 87032.5 10037.5 86897.5 ;
      RECT  9782.5 87032.5 9847.5 86897.5 ;
      RECT  9972.5 87032.5 10037.5 86897.5 ;
      RECT  10162.5 87032.5 10227.5 86897.5 ;
      RECT  10162.5 87032.5 10227.5 86897.5 ;
      RECT  9972.5 87032.5 10037.5 86897.5 ;
      RECT  10332.5 86102.5 10397.5 85967.5 ;
      RECT  10332.5 87077.5 10397.5 86942.5 ;
      RECT  10167.5 86802.5 10032.5 86737.5 ;
      RECT  9910.0 86587.5 9775.0 86522.5 ;
      RECT  9972.5 86192.5 10037.5 86057.5 ;
      RECT  10162.5 87032.5 10227.5 86897.5 ;
      RECT  10262.5 86587.5 10127.5 86522.5 ;
      RECT  9775.0 86587.5 9910.0 86522.5 ;
      RECT  10032.5 86802.5 10167.5 86737.5 ;
      RECT  10127.5 86587.5 10262.5 86522.5 ;
      RECT  9715.0 85882.5 10635.0 85817.5 ;
      RECT  9715.0 87227.5 10635.0 87162.5 ;
      RECT  11062.5 86035.0 11127.5 85850.0 ;
      RECT  11062.5 87195.0 11127.5 87010.0 ;
      RECT  10702.5 87077.5 10767.5 87227.5 ;
      RECT  10702.5 86192.5 10767.5 85817.5 ;
      RECT  10892.5 87077.5 10957.5 86192.5 ;
      RECT  10702.5 86192.5 10767.5 86057.5 ;
      RECT  10892.5 86192.5 10957.5 86057.5 ;
      RECT  10892.5 86192.5 10957.5 86057.5 ;
      RECT  10702.5 86192.5 10767.5 86057.5 ;
      RECT  10702.5 87077.5 10767.5 86942.5 ;
      RECT  10892.5 87077.5 10957.5 86942.5 ;
      RECT  10892.5 87077.5 10957.5 86942.5 ;
      RECT  10702.5 87077.5 10767.5 86942.5 ;
      RECT  11062.5 86102.5 11127.5 85967.5 ;
      RECT  11062.5 87077.5 11127.5 86942.5 ;
      RECT  10760.0 86635.0 10825.0 86500.0 ;
      RECT  10760.0 86635.0 10825.0 86500.0 ;
      RECT  10925.0 86600.0 10990.0 86535.0 ;
      RECT  10635.0 85882.5 11195.0 85817.5 ;
      RECT  10635.0 87227.5 11195.0 87162.5 ;
      RECT  8897.5 86500.0 8962.5 86635.0 ;
      RECT  9037.5 86772.5 9102.5 86907.5 ;
      RECT  10032.5 86737.5 9897.5 86802.5 ;
      RECT  9582.5 88355.0 9647.5 88540.0 ;
      RECT  9582.5 87195.0 9647.5 87380.0 ;
      RECT  9222.5 87312.5 9287.5 87162.5 ;
      RECT  9222.5 88197.5 9287.5 88572.5 ;
      RECT  9412.5 87312.5 9477.5 88197.5 ;
      RECT  9222.5 88197.5 9287.5 88332.5 ;
      RECT  9412.5 88197.5 9477.5 88332.5 ;
      RECT  9412.5 88197.5 9477.5 88332.5 ;
      RECT  9222.5 88197.5 9287.5 88332.5 ;
      RECT  9222.5 87312.5 9287.5 87447.5 ;
      RECT  9412.5 87312.5 9477.5 87447.5 ;
      RECT  9412.5 87312.5 9477.5 87447.5 ;
      RECT  9222.5 87312.5 9287.5 87447.5 ;
      RECT  9582.5 88287.5 9647.5 88422.5 ;
      RECT  9582.5 87312.5 9647.5 87447.5 ;
      RECT  9280.0 87755.0 9345.0 87890.0 ;
      RECT  9280.0 87755.0 9345.0 87890.0 ;
      RECT  9445.0 87790.0 9510.0 87855.0 ;
      RECT  9155.0 88507.5 9715.0 88572.5 ;
      RECT  9155.0 87162.5 9715.0 87227.5 ;
      RECT  9782.5 87357.5 9847.5 87162.5 ;
      RECT  9782.5 88197.5 9847.5 88572.5 ;
      RECT  10162.5 88197.5 10227.5 88572.5 ;
      RECT  10332.5 88355.0 10397.5 88540.0 ;
      RECT  10332.5 87195.0 10397.5 87380.0 ;
      RECT  9782.5 88197.5 9847.5 88332.5 ;
      RECT  9972.5 88197.5 10037.5 88332.5 ;
      RECT  9972.5 88197.5 10037.5 88332.5 ;
      RECT  9782.5 88197.5 9847.5 88332.5 ;
      RECT  9972.5 88197.5 10037.5 88332.5 ;
      RECT  10162.5 88197.5 10227.5 88332.5 ;
      RECT  10162.5 88197.5 10227.5 88332.5 ;
      RECT  9972.5 88197.5 10037.5 88332.5 ;
      RECT  9782.5 87357.5 9847.5 87492.5 ;
      RECT  9972.5 87357.5 10037.5 87492.5 ;
      RECT  9972.5 87357.5 10037.5 87492.5 ;
      RECT  9782.5 87357.5 9847.5 87492.5 ;
      RECT  9972.5 87357.5 10037.5 87492.5 ;
      RECT  10162.5 87357.5 10227.5 87492.5 ;
      RECT  10162.5 87357.5 10227.5 87492.5 ;
      RECT  9972.5 87357.5 10037.5 87492.5 ;
      RECT  10332.5 88287.5 10397.5 88422.5 ;
      RECT  10332.5 87312.5 10397.5 87447.5 ;
      RECT  10167.5 87587.5 10032.5 87652.5 ;
      RECT  9910.0 87802.5 9775.0 87867.5 ;
      RECT  9972.5 88197.5 10037.5 88332.5 ;
      RECT  10162.5 87357.5 10227.5 87492.5 ;
      RECT  10262.5 87802.5 10127.5 87867.5 ;
      RECT  9775.0 87802.5 9910.0 87867.5 ;
      RECT  10032.5 87587.5 10167.5 87652.5 ;
      RECT  10127.5 87802.5 10262.5 87867.5 ;
      RECT  9715.0 88507.5 10635.0 88572.5 ;
      RECT  9715.0 87162.5 10635.0 87227.5 ;
      RECT  11062.5 88355.0 11127.5 88540.0 ;
      RECT  11062.5 87195.0 11127.5 87380.0 ;
      RECT  10702.5 87312.5 10767.5 87162.5 ;
      RECT  10702.5 88197.5 10767.5 88572.5 ;
      RECT  10892.5 87312.5 10957.5 88197.5 ;
      RECT  10702.5 88197.5 10767.5 88332.5 ;
      RECT  10892.5 88197.5 10957.5 88332.5 ;
      RECT  10892.5 88197.5 10957.5 88332.5 ;
      RECT  10702.5 88197.5 10767.5 88332.5 ;
      RECT  10702.5 87312.5 10767.5 87447.5 ;
      RECT  10892.5 87312.5 10957.5 87447.5 ;
      RECT  10892.5 87312.5 10957.5 87447.5 ;
      RECT  10702.5 87312.5 10767.5 87447.5 ;
      RECT  11062.5 88287.5 11127.5 88422.5 ;
      RECT  11062.5 87312.5 11127.5 87447.5 ;
      RECT  10760.0 87755.0 10825.0 87890.0 ;
      RECT  10760.0 87755.0 10825.0 87890.0 ;
      RECT  10925.0 87790.0 10990.0 87855.0 ;
      RECT  10635.0 88507.5 11195.0 88572.5 ;
      RECT  10635.0 87162.5 11195.0 87227.5 ;
      RECT  8897.5 87755.0 8962.5 87890.0 ;
      RECT  9037.5 87482.5 9102.5 87617.5 ;
      RECT  10032.5 87587.5 9897.5 87652.5 ;
      RECT  9582.5 88725.0 9647.5 88540.0 ;
      RECT  9582.5 89885.0 9647.5 89700.0 ;
      RECT  9222.5 89767.5 9287.5 89917.5 ;
      RECT  9222.5 88882.5 9287.5 88507.5 ;
      RECT  9412.5 89767.5 9477.5 88882.5 ;
      RECT  9222.5 88882.5 9287.5 88747.5 ;
      RECT  9412.5 88882.5 9477.5 88747.5 ;
      RECT  9412.5 88882.5 9477.5 88747.5 ;
      RECT  9222.5 88882.5 9287.5 88747.5 ;
      RECT  9222.5 89767.5 9287.5 89632.5 ;
      RECT  9412.5 89767.5 9477.5 89632.5 ;
      RECT  9412.5 89767.5 9477.5 89632.5 ;
      RECT  9222.5 89767.5 9287.5 89632.5 ;
      RECT  9582.5 88792.5 9647.5 88657.5 ;
      RECT  9582.5 89767.5 9647.5 89632.5 ;
      RECT  9280.0 89325.0 9345.0 89190.0 ;
      RECT  9280.0 89325.0 9345.0 89190.0 ;
      RECT  9445.0 89290.0 9510.0 89225.0 ;
      RECT  9155.0 88572.5 9715.0 88507.5 ;
      RECT  9155.0 89917.5 9715.0 89852.5 ;
      RECT  9782.5 89722.5 9847.5 89917.5 ;
      RECT  9782.5 88882.5 9847.5 88507.5 ;
      RECT  10162.5 88882.5 10227.5 88507.5 ;
      RECT  10332.5 88725.0 10397.5 88540.0 ;
      RECT  10332.5 89885.0 10397.5 89700.0 ;
      RECT  9782.5 88882.5 9847.5 88747.5 ;
      RECT  9972.5 88882.5 10037.5 88747.5 ;
      RECT  9972.5 88882.5 10037.5 88747.5 ;
      RECT  9782.5 88882.5 9847.5 88747.5 ;
      RECT  9972.5 88882.5 10037.5 88747.5 ;
      RECT  10162.5 88882.5 10227.5 88747.5 ;
      RECT  10162.5 88882.5 10227.5 88747.5 ;
      RECT  9972.5 88882.5 10037.5 88747.5 ;
      RECT  9782.5 89722.5 9847.5 89587.5 ;
      RECT  9972.5 89722.5 10037.5 89587.5 ;
      RECT  9972.5 89722.5 10037.5 89587.5 ;
      RECT  9782.5 89722.5 9847.5 89587.5 ;
      RECT  9972.5 89722.5 10037.5 89587.5 ;
      RECT  10162.5 89722.5 10227.5 89587.5 ;
      RECT  10162.5 89722.5 10227.5 89587.5 ;
      RECT  9972.5 89722.5 10037.5 89587.5 ;
      RECT  10332.5 88792.5 10397.5 88657.5 ;
      RECT  10332.5 89767.5 10397.5 89632.5 ;
      RECT  10167.5 89492.5 10032.5 89427.5 ;
      RECT  9910.0 89277.5 9775.0 89212.5 ;
      RECT  9972.5 88882.5 10037.5 88747.5 ;
      RECT  10162.5 89722.5 10227.5 89587.5 ;
      RECT  10262.5 89277.5 10127.5 89212.5 ;
      RECT  9775.0 89277.5 9910.0 89212.5 ;
      RECT  10032.5 89492.5 10167.5 89427.5 ;
      RECT  10127.5 89277.5 10262.5 89212.5 ;
      RECT  9715.0 88572.5 10635.0 88507.5 ;
      RECT  9715.0 89917.5 10635.0 89852.5 ;
      RECT  11062.5 88725.0 11127.5 88540.0 ;
      RECT  11062.5 89885.0 11127.5 89700.0 ;
      RECT  10702.5 89767.5 10767.5 89917.5 ;
      RECT  10702.5 88882.5 10767.5 88507.5 ;
      RECT  10892.5 89767.5 10957.5 88882.5 ;
      RECT  10702.5 88882.5 10767.5 88747.5 ;
      RECT  10892.5 88882.5 10957.5 88747.5 ;
      RECT  10892.5 88882.5 10957.5 88747.5 ;
      RECT  10702.5 88882.5 10767.5 88747.5 ;
      RECT  10702.5 89767.5 10767.5 89632.5 ;
      RECT  10892.5 89767.5 10957.5 89632.5 ;
      RECT  10892.5 89767.5 10957.5 89632.5 ;
      RECT  10702.5 89767.5 10767.5 89632.5 ;
      RECT  11062.5 88792.5 11127.5 88657.5 ;
      RECT  11062.5 89767.5 11127.5 89632.5 ;
      RECT  10760.0 89325.0 10825.0 89190.0 ;
      RECT  10760.0 89325.0 10825.0 89190.0 ;
      RECT  10925.0 89290.0 10990.0 89225.0 ;
      RECT  10635.0 88572.5 11195.0 88507.5 ;
      RECT  10635.0 89917.5 11195.0 89852.5 ;
      RECT  8897.5 89190.0 8962.5 89325.0 ;
      RECT  9037.5 89462.5 9102.5 89597.5 ;
      RECT  10032.5 89427.5 9897.5 89492.5 ;
      RECT  9582.5 91045.0 9647.5 91230.0 ;
      RECT  9582.5 89885.0 9647.5 90070.0 ;
      RECT  9222.5 90002.5 9287.5 89852.5 ;
      RECT  9222.5 90887.5 9287.5 91262.5 ;
      RECT  9412.5 90002.5 9477.5 90887.5 ;
      RECT  9222.5 90887.5 9287.5 91022.5 ;
      RECT  9412.5 90887.5 9477.5 91022.5 ;
      RECT  9412.5 90887.5 9477.5 91022.5 ;
      RECT  9222.5 90887.5 9287.5 91022.5 ;
      RECT  9222.5 90002.5 9287.5 90137.5 ;
      RECT  9412.5 90002.5 9477.5 90137.5 ;
      RECT  9412.5 90002.5 9477.5 90137.5 ;
      RECT  9222.5 90002.5 9287.5 90137.5 ;
      RECT  9582.5 90977.5 9647.5 91112.5 ;
      RECT  9582.5 90002.5 9647.5 90137.5 ;
      RECT  9280.0 90445.0 9345.0 90580.0 ;
      RECT  9280.0 90445.0 9345.0 90580.0 ;
      RECT  9445.0 90480.0 9510.0 90545.0 ;
      RECT  9155.0 91197.5 9715.0 91262.5 ;
      RECT  9155.0 89852.5 9715.0 89917.5 ;
      RECT  9782.5 90047.5 9847.5 89852.5 ;
      RECT  9782.5 90887.5 9847.5 91262.5 ;
      RECT  10162.5 90887.5 10227.5 91262.5 ;
      RECT  10332.5 91045.0 10397.5 91230.0 ;
      RECT  10332.5 89885.0 10397.5 90070.0 ;
      RECT  9782.5 90887.5 9847.5 91022.5 ;
      RECT  9972.5 90887.5 10037.5 91022.5 ;
      RECT  9972.5 90887.5 10037.5 91022.5 ;
      RECT  9782.5 90887.5 9847.5 91022.5 ;
      RECT  9972.5 90887.5 10037.5 91022.5 ;
      RECT  10162.5 90887.5 10227.5 91022.5 ;
      RECT  10162.5 90887.5 10227.5 91022.5 ;
      RECT  9972.5 90887.5 10037.5 91022.5 ;
      RECT  9782.5 90047.5 9847.5 90182.5 ;
      RECT  9972.5 90047.5 10037.5 90182.5 ;
      RECT  9972.5 90047.5 10037.5 90182.5 ;
      RECT  9782.5 90047.5 9847.5 90182.5 ;
      RECT  9972.5 90047.5 10037.5 90182.5 ;
      RECT  10162.5 90047.5 10227.5 90182.5 ;
      RECT  10162.5 90047.5 10227.5 90182.5 ;
      RECT  9972.5 90047.5 10037.5 90182.5 ;
      RECT  10332.5 90977.5 10397.5 91112.5 ;
      RECT  10332.5 90002.5 10397.5 90137.5 ;
      RECT  10167.5 90277.5 10032.5 90342.5 ;
      RECT  9910.0 90492.5 9775.0 90557.5 ;
      RECT  9972.5 90887.5 10037.5 91022.5 ;
      RECT  10162.5 90047.5 10227.5 90182.5 ;
      RECT  10262.5 90492.5 10127.5 90557.5 ;
      RECT  9775.0 90492.5 9910.0 90557.5 ;
      RECT  10032.5 90277.5 10167.5 90342.5 ;
      RECT  10127.5 90492.5 10262.5 90557.5 ;
      RECT  9715.0 91197.5 10635.0 91262.5 ;
      RECT  9715.0 89852.5 10635.0 89917.5 ;
      RECT  11062.5 91045.0 11127.5 91230.0 ;
      RECT  11062.5 89885.0 11127.5 90070.0 ;
      RECT  10702.5 90002.5 10767.5 89852.5 ;
      RECT  10702.5 90887.5 10767.5 91262.5 ;
      RECT  10892.5 90002.5 10957.5 90887.5 ;
      RECT  10702.5 90887.5 10767.5 91022.5 ;
      RECT  10892.5 90887.5 10957.5 91022.5 ;
      RECT  10892.5 90887.5 10957.5 91022.5 ;
      RECT  10702.5 90887.5 10767.5 91022.5 ;
      RECT  10702.5 90002.5 10767.5 90137.5 ;
      RECT  10892.5 90002.5 10957.5 90137.5 ;
      RECT  10892.5 90002.5 10957.5 90137.5 ;
      RECT  10702.5 90002.5 10767.5 90137.5 ;
      RECT  11062.5 90977.5 11127.5 91112.5 ;
      RECT  11062.5 90002.5 11127.5 90137.5 ;
      RECT  10760.0 90445.0 10825.0 90580.0 ;
      RECT  10760.0 90445.0 10825.0 90580.0 ;
      RECT  10925.0 90480.0 10990.0 90545.0 ;
      RECT  10635.0 91197.5 11195.0 91262.5 ;
      RECT  10635.0 89852.5 11195.0 89917.5 ;
      RECT  8897.5 90445.0 8962.5 90580.0 ;
      RECT  9037.5 90172.5 9102.5 90307.5 ;
      RECT  10032.5 90277.5 9897.5 90342.5 ;
      RECT  9582.5 91415.0 9647.5 91230.0 ;
      RECT  9582.5 92575.0 9647.5 92390.0 ;
      RECT  9222.5 92457.5 9287.5 92607.5 ;
      RECT  9222.5 91572.5 9287.5 91197.5 ;
      RECT  9412.5 92457.5 9477.5 91572.5 ;
      RECT  9222.5 91572.5 9287.5 91437.5 ;
      RECT  9412.5 91572.5 9477.5 91437.5 ;
      RECT  9412.5 91572.5 9477.5 91437.5 ;
      RECT  9222.5 91572.5 9287.5 91437.5 ;
      RECT  9222.5 92457.5 9287.5 92322.5 ;
      RECT  9412.5 92457.5 9477.5 92322.5 ;
      RECT  9412.5 92457.5 9477.5 92322.5 ;
      RECT  9222.5 92457.5 9287.5 92322.5 ;
      RECT  9582.5 91482.5 9647.5 91347.5 ;
      RECT  9582.5 92457.5 9647.5 92322.5 ;
      RECT  9280.0 92015.0 9345.0 91880.0 ;
      RECT  9280.0 92015.0 9345.0 91880.0 ;
      RECT  9445.0 91980.0 9510.0 91915.0 ;
      RECT  9155.0 91262.5 9715.0 91197.5 ;
      RECT  9155.0 92607.5 9715.0 92542.5 ;
      RECT  9782.5 92412.5 9847.5 92607.5 ;
      RECT  9782.5 91572.5 9847.5 91197.5 ;
      RECT  10162.5 91572.5 10227.5 91197.5 ;
      RECT  10332.5 91415.0 10397.5 91230.0 ;
      RECT  10332.5 92575.0 10397.5 92390.0 ;
      RECT  9782.5 91572.5 9847.5 91437.5 ;
      RECT  9972.5 91572.5 10037.5 91437.5 ;
      RECT  9972.5 91572.5 10037.5 91437.5 ;
      RECT  9782.5 91572.5 9847.5 91437.5 ;
      RECT  9972.5 91572.5 10037.5 91437.5 ;
      RECT  10162.5 91572.5 10227.5 91437.5 ;
      RECT  10162.5 91572.5 10227.5 91437.5 ;
      RECT  9972.5 91572.5 10037.5 91437.5 ;
      RECT  9782.5 92412.5 9847.5 92277.5 ;
      RECT  9972.5 92412.5 10037.5 92277.5 ;
      RECT  9972.5 92412.5 10037.5 92277.5 ;
      RECT  9782.5 92412.5 9847.5 92277.5 ;
      RECT  9972.5 92412.5 10037.5 92277.5 ;
      RECT  10162.5 92412.5 10227.5 92277.5 ;
      RECT  10162.5 92412.5 10227.5 92277.5 ;
      RECT  9972.5 92412.5 10037.5 92277.5 ;
      RECT  10332.5 91482.5 10397.5 91347.5 ;
      RECT  10332.5 92457.5 10397.5 92322.5 ;
      RECT  10167.5 92182.5 10032.5 92117.5 ;
      RECT  9910.0 91967.5 9775.0 91902.5 ;
      RECT  9972.5 91572.5 10037.5 91437.5 ;
      RECT  10162.5 92412.5 10227.5 92277.5 ;
      RECT  10262.5 91967.5 10127.5 91902.5 ;
      RECT  9775.0 91967.5 9910.0 91902.5 ;
      RECT  10032.5 92182.5 10167.5 92117.5 ;
      RECT  10127.5 91967.5 10262.5 91902.5 ;
      RECT  9715.0 91262.5 10635.0 91197.5 ;
      RECT  9715.0 92607.5 10635.0 92542.5 ;
      RECT  11062.5 91415.0 11127.5 91230.0 ;
      RECT  11062.5 92575.0 11127.5 92390.0 ;
      RECT  10702.5 92457.5 10767.5 92607.5 ;
      RECT  10702.5 91572.5 10767.5 91197.5 ;
      RECT  10892.5 92457.5 10957.5 91572.5 ;
      RECT  10702.5 91572.5 10767.5 91437.5 ;
      RECT  10892.5 91572.5 10957.5 91437.5 ;
      RECT  10892.5 91572.5 10957.5 91437.5 ;
      RECT  10702.5 91572.5 10767.5 91437.5 ;
      RECT  10702.5 92457.5 10767.5 92322.5 ;
      RECT  10892.5 92457.5 10957.5 92322.5 ;
      RECT  10892.5 92457.5 10957.5 92322.5 ;
      RECT  10702.5 92457.5 10767.5 92322.5 ;
      RECT  11062.5 91482.5 11127.5 91347.5 ;
      RECT  11062.5 92457.5 11127.5 92322.5 ;
      RECT  10760.0 92015.0 10825.0 91880.0 ;
      RECT  10760.0 92015.0 10825.0 91880.0 ;
      RECT  10925.0 91980.0 10990.0 91915.0 ;
      RECT  10635.0 91262.5 11195.0 91197.5 ;
      RECT  10635.0 92607.5 11195.0 92542.5 ;
      RECT  8897.5 91880.0 8962.5 92015.0 ;
      RECT  9037.5 92152.5 9102.5 92287.5 ;
      RECT  10032.5 92117.5 9897.5 92182.5 ;
      RECT  9582.5 93735.0 9647.5 93920.0 ;
      RECT  9582.5 92575.0 9647.5 92760.0 ;
      RECT  9222.5 92692.5 9287.5 92542.5 ;
      RECT  9222.5 93577.5 9287.5 93952.5 ;
      RECT  9412.5 92692.5 9477.5 93577.5 ;
      RECT  9222.5 93577.5 9287.5 93712.5 ;
      RECT  9412.5 93577.5 9477.5 93712.5 ;
      RECT  9412.5 93577.5 9477.5 93712.5 ;
      RECT  9222.5 93577.5 9287.5 93712.5 ;
      RECT  9222.5 92692.5 9287.5 92827.5 ;
      RECT  9412.5 92692.5 9477.5 92827.5 ;
      RECT  9412.5 92692.5 9477.5 92827.5 ;
      RECT  9222.5 92692.5 9287.5 92827.5 ;
      RECT  9582.5 93667.5 9647.5 93802.5 ;
      RECT  9582.5 92692.5 9647.5 92827.5 ;
      RECT  9280.0 93135.0 9345.0 93270.0 ;
      RECT  9280.0 93135.0 9345.0 93270.0 ;
      RECT  9445.0 93170.0 9510.0 93235.0 ;
      RECT  9155.0 93887.5 9715.0 93952.5 ;
      RECT  9155.0 92542.5 9715.0 92607.5 ;
      RECT  9782.5 92737.5 9847.5 92542.5 ;
      RECT  9782.5 93577.5 9847.5 93952.5 ;
      RECT  10162.5 93577.5 10227.5 93952.5 ;
      RECT  10332.5 93735.0 10397.5 93920.0 ;
      RECT  10332.5 92575.0 10397.5 92760.0 ;
      RECT  9782.5 93577.5 9847.5 93712.5 ;
      RECT  9972.5 93577.5 10037.5 93712.5 ;
      RECT  9972.5 93577.5 10037.5 93712.5 ;
      RECT  9782.5 93577.5 9847.5 93712.5 ;
      RECT  9972.5 93577.5 10037.5 93712.5 ;
      RECT  10162.5 93577.5 10227.5 93712.5 ;
      RECT  10162.5 93577.5 10227.5 93712.5 ;
      RECT  9972.5 93577.5 10037.5 93712.5 ;
      RECT  9782.5 92737.5 9847.5 92872.5 ;
      RECT  9972.5 92737.5 10037.5 92872.5 ;
      RECT  9972.5 92737.5 10037.5 92872.5 ;
      RECT  9782.5 92737.5 9847.5 92872.5 ;
      RECT  9972.5 92737.5 10037.5 92872.5 ;
      RECT  10162.5 92737.5 10227.5 92872.5 ;
      RECT  10162.5 92737.5 10227.5 92872.5 ;
      RECT  9972.5 92737.5 10037.5 92872.5 ;
      RECT  10332.5 93667.5 10397.5 93802.5 ;
      RECT  10332.5 92692.5 10397.5 92827.5 ;
      RECT  10167.5 92967.5 10032.5 93032.5 ;
      RECT  9910.0 93182.5 9775.0 93247.5 ;
      RECT  9972.5 93577.5 10037.5 93712.5 ;
      RECT  10162.5 92737.5 10227.5 92872.5 ;
      RECT  10262.5 93182.5 10127.5 93247.5 ;
      RECT  9775.0 93182.5 9910.0 93247.5 ;
      RECT  10032.5 92967.5 10167.5 93032.5 ;
      RECT  10127.5 93182.5 10262.5 93247.5 ;
      RECT  9715.0 93887.5 10635.0 93952.5 ;
      RECT  9715.0 92542.5 10635.0 92607.5 ;
      RECT  11062.5 93735.0 11127.5 93920.0 ;
      RECT  11062.5 92575.0 11127.5 92760.0 ;
      RECT  10702.5 92692.5 10767.5 92542.5 ;
      RECT  10702.5 93577.5 10767.5 93952.5 ;
      RECT  10892.5 92692.5 10957.5 93577.5 ;
      RECT  10702.5 93577.5 10767.5 93712.5 ;
      RECT  10892.5 93577.5 10957.5 93712.5 ;
      RECT  10892.5 93577.5 10957.5 93712.5 ;
      RECT  10702.5 93577.5 10767.5 93712.5 ;
      RECT  10702.5 92692.5 10767.5 92827.5 ;
      RECT  10892.5 92692.5 10957.5 92827.5 ;
      RECT  10892.5 92692.5 10957.5 92827.5 ;
      RECT  10702.5 92692.5 10767.5 92827.5 ;
      RECT  11062.5 93667.5 11127.5 93802.5 ;
      RECT  11062.5 92692.5 11127.5 92827.5 ;
      RECT  10760.0 93135.0 10825.0 93270.0 ;
      RECT  10760.0 93135.0 10825.0 93270.0 ;
      RECT  10925.0 93170.0 10990.0 93235.0 ;
      RECT  10635.0 93887.5 11195.0 93952.5 ;
      RECT  10635.0 92542.5 11195.0 92607.5 ;
      RECT  8897.5 93135.0 8962.5 93270.0 ;
      RECT  9037.5 92862.5 9102.5 92997.5 ;
      RECT  10032.5 92967.5 9897.5 93032.5 ;
      RECT  9582.5 94105.0 9647.5 93920.0 ;
      RECT  9582.5 95265.0 9647.5 95080.0 ;
      RECT  9222.5 95147.5 9287.5 95297.5 ;
      RECT  9222.5 94262.5 9287.5 93887.5 ;
      RECT  9412.5 95147.5 9477.5 94262.5 ;
      RECT  9222.5 94262.5 9287.5 94127.5 ;
      RECT  9412.5 94262.5 9477.5 94127.5 ;
      RECT  9412.5 94262.5 9477.5 94127.5 ;
      RECT  9222.5 94262.5 9287.5 94127.5 ;
      RECT  9222.5 95147.5 9287.5 95012.5 ;
      RECT  9412.5 95147.5 9477.5 95012.5 ;
      RECT  9412.5 95147.5 9477.5 95012.5 ;
      RECT  9222.5 95147.5 9287.5 95012.5 ;
      RECT  9582.5 94172.5 9647.5 94037.5 ;
      RECT  9582.5 95147.5 9647.5 95012.5 ;
      RECT  9280.0 94705.0 9345.0 94570.0 ;
      RECT  9280.0 94705.0 9345.0 94570.0 ;
      RECT  9445.0 94670.0 9510.0 94605.0 ;
      RECT  9155.0 93952.5 9715.0 93887.5 ;
      RECT  9155.0 95297.5 9715.0 95232.5 ;
      RECT  9782.5 95102.5 9847.5 95297.5 ;
      RECT  9782.5 94262.5 9847.5 93887.5 ;
      RECT  10162.5 94262.5 10227.5 93887.5 ;
      RECT  10332.5 94105.0 10397.5 93920.0 ;
      RECT  10332.5 95265.0 10397.5 95080.0 ;
      RECT  9782.5 94262.5 9847.5 94127.5 ;
      RECT  9972.5 94262.5 10037.5 94127.5 ;
      RECT  9972.5 94262.5 10037.5 94127.5 ;
      RECT  9782.5 94262.5 9847.5 94127.5 ;
      RECT  9972.5 94262.5 10037.5 94127.5 ;
      RECT  10162.5 94262.5 10227.5 94127.5 ;
      RECT  10162.5 94262.5 10227.5 94127.5 ;
      RECT  9972.5 94262.5 10037.5 94127.5 ;
      RECT  9782.5 95102.5 9847.5 94967.5 ;
      RECT  9972.5 95102.5 10037.5 94967.5 ;
      RECT  9972.5 95102.5 10037.5 94967.5 ;
      RECT  9782.5 95102.5 9847.5 94967.5 ;
      RECT  9972.5 95102.5 10037.5 94967.5 ;
      RECT  10162.5 95102.5 10227.5 94967.5 ;
      RECT  10162.5 95102.5 10227.5 94967.5 ;
      RECT  9972.5 95102.5 10037.5 94967.5 ;
      RECT  10332.5 94172.5 10397.5 94037.5 ;
      RECT  10332.5 95147.5 10397.5 95012.5 ;
      RECT  10167.5 94872.5 10032.5 94807.5 ;
      RECT  9910.0 94657.5 9775.0 94592.5 ;
      RECT  9972.5 94262.5 10037.5 94127.5 ;
      RECT  10162.5 95102.5 10227.5 94967.5 ;
      RECT  10262.5 94657.5 10127.5 94592.5 ;
      RECT  9775.0 94657.5 9910.0 94592.5 ;
      RECT  10032.5 94872.5 10167.5 94807.5 ;
      RECT  10127.5 94657.5 10262.5 94592.5 ;
      RECT  9715.0 93952.5 10635.0 93887.5 ;
      RECT  9715.0 95297.5 10635.0 95232.5 ;
      RECT  11062.5 94105.0 11127.5 93920.0 ;
      RECT  11062.5 95265.0 11127.5 95080.0 ;
      RECT  10702.5 95147.5 10767.5 95297.5 ;
      RECT  10702.5 94262.5 10767.5 93887.5 ;
      RECT  10892.5 95147.5 10957.5 94262.5 ;
      RECT  10702.5 94262.5 10767.5 94127.5 ;
      RECT  10892.5 94262.5 10957.5 94127.5 ;
      RECT  10892.5 94262.5 10957.5 94127.5 ;
      RECT  10702.5 94262.5 10767.5 94127.5 ;
      RECT  10702.5 95147.5 10767.5 95012.5 ;
      RECT  10892.5 95147.5 10957.5 95012.5 ;
      RECT  10892.5 95147.5 10957.5 95012.5 ;
      RECT  10702.5 95147.5 10767.5 95012.5 ;
      RECT  11062.5 94172.5 11127.5 94037.5 ;
      RECT  11062.5 95147.5 11127.5 95012.5 ;
      RECT  10760.0 94705.0 10825.0 94570.0 ;
      RECT  10760.0 94705.0 10825.0 94570.0 ;
      RECT  10925.0 94670.0 10990.0 94605.0 ;
      RECT  10635.0 93952.5 11195.0 93887.5 ;
      RECT  10635.0 95297.5 11195.0 95232.5 ;
      RECT  8897.5 94570.0 8962.5 94705.0 ;
      RECT  9037.5 94842.5 9102.5 94977.5 ;
      RECT  10032.5 94807.5 9897.5 94872.5 ;
      RECT  9582.5 96425.0 9647.5 96610.0 ;
      RECT  9582.5 95265.0 9647.5 95450.0 ;
      RECT  9222.5 95382.5 9287.5 95232.5 ;
      RECT  9222.5 96267.5 9287.5 96642.5 ;
      RECT  9412.5 95382.5 9477.5 96267.5 ;
      RECT  9222.5 96267.5 9287.5 96402.5 ;
      RECT  9412.5 96267.5 9477.5 96402.5 ;
      RECT  9412.5 96267.5 9477.5 96402.5 ;
      RECT  9222.5 96267.5 9287.5 96402.5 ;
      RECT  9222.5 95382.5 9287.5 95517.5 ;
      RECT  9412.5 95382.5 9477.5 95517.5 ;
      RECT  9412.5 95382.5 9477.5 95517.5 ;
      RECT  9222.5 95382.5 9287.5 95517.5 ;
      RECT  9582.5 96357.5 9647.5 96492.5 ;
      RECT  9582.5 95382.5 9647.5 95517.5 ;
      RECT  9280.0 95825.0 9345.0 95960.0 ;
      RECT  9280.0 95825.0 9345.0 95960.0 ;
      RECT  9445.0 95860.0 9510.0 95925.0 ;
      RECT  9155.0 96577.5 9715.0 96642.5 ;
      RECT  9155.0 95232.5 9715.0 95297.5 ;
      RECT  9782.5 95427.5 9847.5 95232.5 ;
      RECT  9782.5 96267.5 9847.5 96642.5 ;
      RECT  10162.5 96267.5 10227.5 96642.5 ;
      RECT  10332.5 96425.0 10397.5 96610.0 ;
      RECT  10332.5 95265.0 10397.5 95450.0 ;
      RECT  9782.5 96267.5 9847.5 96402.5 ;
      RECT  9972.5 96267.5 10037.5 96402.5 ;
      RECT  9972.5 96267.5 10037.5 96402.5 ;
      RECT  9782.5 96267.5 9847.5 96402.5 ;
      RECT  9972.5 96267.5 10037.5 96402.5 ;
      RECT  10162.5 96267.5 10227.5 96402.5 ;
      RECT  10162.5 96267.5 10227.5 96402.5 ;
      RECT  9972.5 96267.5 10037.5 96402.5 ;
      RECT  9782.5 95427.5 9847.5 95562.5 ;
      RECT  9972.5 95427.5 10037.5 95562.5 ;
      RECT  9972.5 95427.5 10037.5 95562.5 ;
      RECT  9782.5 95427.5 9847.5 95562.5 ;
      RECT  9972.5 95427.5 10037.5 95562.5 ;
      RECT  10162.5 95427.5 10227.5 95562.5 ;
      RECT  10162.5 95427.5 10227.5 95562.5 ;
      RECT  9972.5 95427.5 10037.5 95562.5 ;
      RECT  10332.5 96357.5 10397.5 96492.5 ;
      RECT  10332.5 95382.5 10397.5 95517.5 ;
      RECT  10167.5 95657.5 10032.5 95722.5 ;
      RECT  9910.0 95872.5 9775.0 95937.5 ;
      RECT  9972.5 96267.5 10037.5 96402.5 ;
      RECT  10162.5 95427.5 10227.5 95562.5 ;
      RECT  10262.5 95872.5 10127.5 95937.5 ;
      RECT  9775.0 95872.5 9910.0 95937.5 ;
      RECT  10032.5 95657.5 10167.5 95722.5 ;
      RECT  10127.5 95872.5 10262.5 95937.5 ;
      RECT  9715.0 96577.5 10635.0 96642.5 ;
      RECT  9715.0 95232.5 10635.0 95297.5 ;
      RECT  11062.5 96425.0 11127.5 96610.0 ;
      RECT  11062.5 95265.0 11127.5 95450.0 ;
      RECT  10702.5 95382.5 10767.5 95232.5 ;
      RECT  10702.5 96267.5 10767.5 96642.5 ;
      RECT  10892.5 95382.5 10957.5 96267.5 ;
      RECT  10702.5 96267.5 10767.5 96402.5 ;
      RECT  10892.5 96267.5 10957.5 96402.5 ;
      RECT  10892.5 96267.5 10957.5 96402.5 ;
      RECT  10702.5 96267.5 10767.5 96402.5 ;
      RECT  10702.5 95382.5 10767.5 95517.5 ;
      RECT  10892.5 95382.5 10957.5 95517.5 ;
      RECT  10892.5 95382.5 10957.5 95517.5 ;
      RECT  10702.5 95382.5 10767.5 95517.5 ;
      RECT  11062.5 96357.5 11127.5 96492.5 ;
      RECT  11062.5 95382.5 11127.5 95517.5 ;
      RECT  10760.0 95825.0 10825.0 95960.0 ;
      RECT  10760.0 95825.0 10825.0 95960.0 ;
      RECT  10925.0 95860.0 10990.0 95925.0 ;
      RECT  10635.0 96577.5 11195.0 96642.5 ;
      RECT  10635.0 95232.5 11195.0 95297.5 ;
      RECT  8897.5 95825.0 8962.5 95960.0 ;
      RECT  9037.5 95552.5 9102.5 95687.5 ;
      RECT  10032.5 95657.5 9897.5 95722.5 ;
      RECT  9582.5 96795.0 9647.5 96610.0 ;
      RECT  9582.5 97955.0 9647.5 97770.0 ;
      RECT  9222.5 97837.5 9287.5 97987.5 ;
      RECT  9222.5 96952.5 9287.5 96577.5 ;
      RECT  9412.5 97837.5 9477.5 96952.5 ;
      RECT  9222.5 96952.5 9287.5 96817.5 ;
      RECT  9412.5 96952.5 9477.5 96817.5 ;
      RECT  9412.5 96952.5 9477.5 96817.5 ;
      RECT  9222.5 96952.5 9287.5 96817.5 ;
      RECT  9222.5 97837.5 9287.5 97702.5 ;
      RECT  9412.5 97837.5 9477.5 97702.5 ;
      RECT  9412.5 97837.5 9477.5 97702.5 ;
      RECT  9222.5 97837.5 9287.5 97702.5 ;
      RECT  9582.5 96862.5 9647.5 96727.5 ;
      RECT  9582.5 97837.5 9647.5 97702.5 ;
      RECT  9280.0 97395.0 9345.0 97260.0 ;
      RECT  9280.0 97395.0 9345.0 97260.0 ;
      RECT  9445.0 97360.0 9510.0 97295.0 ;
      RECT  9155.0 96642.5 9715.0 96577.5 ;
      RECT  9155.0 97987.5 9715.0 97922.5 ;
      RECT  9782.5 97792.5 9847.5 97987.5 ;
      RECT  9782.5 96952.5 9847.5 96577.5 ;
      RECT  10162.5 96952.5 10227.5 96577.5 ;
      RECT  10332.5 96795.0 10397.5 96610.0 ;
      RECT  10332.5 97955.0 10397.5 97770.0 ;
      RECT  9782.5 96952.5 9847.5 96817.5 ;
      RECT  9972.5 96952.5 10037.5 96817.5 ;
      RECT  9972.5 96952.5 10037.5 96817.5 ;
      RECT  9782.5 96952.5 9847.5 96817.5 ;
      RECT  9972.5 96952.5 10037.5 96817.5 ;
      RECT  10162.5 96952.5 10227.5 96817.5 ;
      RECT  10162.5 96952.5 10227.5 96817.5 ;
      RECT  9972.5 96952.5 10037.5 96817.5 ;
      RECT  9782.5 97792.5 9847.5 97657.5 ;
      RECT  9972.5 97792.5 10037.5 97657.5 ;
      RECT  9972.5 97792.5 10037.5 97657.5 ;
      RECT  9782.5 97792.5 9847.5 97657.5 ;
      RECT  9972.5 97792.5 10037.5 97657.5 ;
      RECT  10162.5 97792.5 10227.5 97657.5 ;
      RECT  10162.5 97792.5 10227.5 97657.5 ;
      RECT  9972.5 97792.5 10037.5 97657.5 ;
      RECT  10332.5 96862.5 10397.5 96727.5 ;
      RECT  10332.5 97837.5 10397.5 97702.5 ;
      RECT  10167.5 97562.5 10032.5 97497.5 ;
      RECT  9910.0 97347.5 9775.0 97282.5 ;
      RECT  9972.5 96952.5 10037.5 96817.5 ;
      RECT  10162.5 97792.5 10227.5 97657.5 ;
      RECT  10262.5 97347.5 10127.5 97282.5 ;
      RECT  9775.0 97347.5 9910.0 97282.5 ;
      RECT  10032.5 97562.5 10167.5 97497.5 ;
      RECT  10127.5 97347.5 10262.5 97282.5 ;
      RECT  9715.0 96642.5 10635.0 96577.5 ;
      RECT  9715.0 97987.5 10635.0 97922.5 ;
      RECT  11062.5 96795.0 11127.5 96610.0 ;
      RECT  11062.5 97955.0 11127.5 97770.0 ;
      RECT  10702.5 97837.5 10767.5 97987.5 ;
      RECT  10702.5 96952.5 10767.5 96577.5 ;
      RECT  10892.5 97837.5 10957.5 96952.5 ;
      RECT  10702.5 96952.5 10767.5 96817.5 ;
      RECT  10892.5 96952.5 10957.5 96817.5 ;
      RECT  10892.5 96952.5 10957.5 96817.5 ;
      RECT  10702.5 96952.5 10767.5 96817.5 ;
      RECT  10702.5 97837.5 10767.5 97702.5 ;
      RECT  10892.5 97837.5 10957.5 97702.5 ;
      RECT  10892.5 97837.5 10957.5 97702.5 ;
      RECT  10702.5 97837.5 10767.5 97702.5 ;
      RECT  11062.5 96862.5 11127.5 96727.5 ;
      RECT  11062.5 97837.5 11127.5 97702.5 ;
      RECT  10760.0 97395.0 10825.0 97260.0 ;
      RECT  10760.0 97395.0 10825.0 97260.0 ;
      RECT  10925.0 97360.0 10990.0 97295.0 ;
      RECT  10635.0 96642.5 11195.0 96577.5 ;
      RECT  10635.0 97987.5 11195.0 97922.5 ;
      RECT  8897.5 97260.0 8962.5 97395.0 ;
      RECT  9037.5 97532.5 9102.5 97667.5 ;
      RECT  10032.5 97497.5 9897.5 97562.5 ;
      RECT  9582.5 99115.0 9647.5 99300.0 ;
      RECT  9582.5 97955.0 9647.5 98140.0 ;
      RECT  9222.5 98072.5 9287.5 97922.5 ;
      RECT  9222.5 98957.5 9287.5 99332.5 ;
      RECT  9412.5 98072.5 9477.5 98957.5 ;
      RECT  9222.5 98957.5 9287.5 99092.5 ;
      RECT  9412.5 98957.5 9477.5 99092.5 ;
      RECT  9412.5 98957.5 9477.5 99092.5 ;
      RECT  9222.5 98957.5 9287.5 99092.5 ;
      RECT  9222.5 98072.5 9287.5 98207.5 ;
      RECT  9412.5 98072.5 9477.5 98207.5 ;
      RECT  9412.5 98072.5 9477.5 98207.5 ;
      RECT  9222.5 98072.5 9287.5 98207.5 ;
      RECT  9582.5 99047.5 9647.5 99182.5 ;
      RECT  9582.5 98072.5 9647.5 98207.5 ;
      RECT  9280.0 98515.0 9345.0 98650.0 ;
      RECT  9280.0 98515.0 9345.0 98650.0 ;
      RECT  9445.0 98550.0 9510.0 98615.0 ;
      RECT  9155.0 99267.5 9715.0 99332.5 ;
      RECT  9155.0 97922.5 9715.0 97987.5 ;
      RECT  9782.5 98117.5 9847.5 97922.5 ;
      RECT  9782.5 98957.5 9847.5 99332.5 ;
      RECT  10162.5 98957.5 10227.5 99332.5 ;
      RECT  10332.5 99115.0 10397.5 99300.0 ;
      RECT  10332.5 97955.0 10397.5 98140.0 ;
      RECT  9782.5 98957.5 9847.5 99092.5 ;
      RECT  9972.5 98957.5 10037.5 99092.5 ;
      RECT  9972.5 98957.5 10037.5 99092.5 ;
      RECT  9782.5 98957.5 9847.5 99092.5 ;
      RECT  9972.5 98957.5 10037.5 99092.5 ;
      RECT  10162.5 98957.5 10227.5 99092.5 ;
      RECT  10162.5 98957.5 10227.5 99092.5 ;
      RECT  9972.5 98957.5 10037.5 99092.5 ;
      RECT  9782.5 98117.5 9847.5 98252.5 ;
      RECT  9972.5 98117.5 10037.5 98252.5 ;
      RECT  9972.5 98117.5 10037.5 98252.5 ;
      RECT  9782.5 98117.5 9847.5 98252.5 ;
      RECT  9972.5 98117.5 10037.5 98252.5 ;
      RECT  10162.5 98117.5 10227.5 98252.5 ;
      RECT  10162.5 98117.5 10227.5 98252.5 ;
      RECT  9972.5 98117.5 10037.5 98252.5 ;
      RECT  10332.5 99047.5 10397.5 99182.5 ;
      RECT  10332.5 98072.5 10397.5 98207.5 ;
      RECT  10167.5 98347.5 10032.5 98412.5 ;
      RECT  9910.0 98562.5 9775.0 98627.5 ;
      RECT  9972.5 98957.5 10037.5 99092.5 ;
      RECT  10162.5 98117.5 10227.5 98252.5 ;
      RECT  10262.5 98562.5 10127.5 98627.5 ;
      RECT  9775.0 98562.5 9910.0 98627.5 ;
      RECT  10032.5 98347.5 10167.5 98412.5 ;
      RECT  10127.5 98562.5 10262.5 98627.5 ;
      RECT  9715.0 99267.5 10635.0 99332.5 ;
      RECT  9715.0 97922.5 10635.0 97987.5 ;
      RECT  11062.5 99115.0 11127.5 99300.0 ;
      RECT  11062.5 97955.0 11127.5 98140.0 ;
      RECT  10702.5 98072.5 10767.5 97922.5 ;
      RECT  10702.5 98957.5 10767.5 99332.5 ;
      RECT  10892.5 98072.5 10957.5 98957.5 ;
      RECT  10702.5 98957.5 10767.5 99092.5 ;
      RECT  10892.5 98957.5 10957.5 99092.5 ;
      RECT  10892.5 98957.5 10957.5 99092.5 ;
      RECT  10702.5 98957.5 10767.5 99092.5 ;
      RECT  10702.5 98072.5 10767.5 98207.5 ;
      RECT  10892.5 98072.5 10957.5 98207.5 ;
      RECT  10892.5 98072.5 10957.5 98207.5 ;
      RECT  10702.5 98072.5 10767.5 98207.5 ;
      RECT  11062.5 99047.5 11127.5 99182.5 ;
      RECT  11062.5 98072.5 11127.5 98207.5 ;
      RECT  10760.0 98515.0 10825.0 98650.0 ;
      RECT  10760.0 98515.0 10825.0 98650.0 ;
      RECT  10925.0 98550.0 10990.0 98615.0 ;
      RECT  10635.0 99267.5 11195.0 99332.5 ;
      RECT  10635.0 97922.5 11195.0 97987.5 ;
      RECT  8897.5 98515.0 8962.5 98650.0 ;
      RECT  9037.5 98242.5 9102.5 98377.5 ;
      RECT  10032.5 98347.5 9897.5 98412.5 ;
      RECT  9582.5 99485.0 9647.5 99300.0 ;
      RECT  9582.5 100645.0 9647.5 100460.0 ;
      RECT  9222.5 100527.5 9287.5 100677.5 ;
      RECT  9222.5 99642.5 9287.5 99267.5 ;
      RECT  9412.5 100527.5 9477.5 99642.5 ;
      RECT  9222.5 99642.5 9287.5 99507.5 ;
      RECT  9412.5 99642.5 9477.5 99507.5 ;
      RECT  9412.5 99642.5 9477.5 99507.5 ;
      RECT  9222.5 99642.5 9287.5 99507.5 ;
      RECT  9222.5 100527.5 9287.5 100392.5 ;
      RECT  9412.5 100527.5 9477.5 100392.5 ;
      RECT  9412.5 100527.5 9477.5 100392.5 ;
      RECT  9222.5 100527.5 9287.5 100392.5 ;
      RECT  9582.5 99552.5 9647.5 99417.5 ;
      RECT  9582.5 100527.5 9647.5 100392.5 ;
      RECT  9280.0 100085.0 9345.0 99950.0 ;
      RECT  9280.0 100085.0 9345.0 99950.0 ;
      RECT  9445.0 100050.0 9510.0 99985.0 ;
      RECT  9155.0 99332.5 9715.0 99267.5 ;
      RECT  9155.0 100677.5 9715.0 100612.5 ;
      RECT  9782.5 100482.5 9847.5 100677.5 ;
      RECT  9782.5 99642.5 9847.5 99267.5 ;
      RECT  10162.5 99642.5 10227.5 99267.5 ;
      RECT  10332.5 99485.0 10397.5 99300.0 ;
      RECT  10332.5 100645.0 10397.5 100460.0 ;
      RECT  9782.5 99642.5 9847.5 99507.5 ;
      RECT  9972.5 99642.5 10037.5 99507.5 ;
      RECT  9972.5 99642.5 10037.5 99507.5 ;
      RECT  9782.5 99642.5 9847.5 99507.5 ;
      RECT  9972.5 99642.5 10037.5 99507.5 ;
      RECT  10162.5 99642.5 10227.5 99507.5 ;
      RECT  10162.5 99642.5 10227.5 99507.5 ;
      RECT  9972.5 99642.5 10037.5 99507.5 ;
      RECT  9782.5 100482.5 9847.5 100347.5 ;
      RECT  9972.5 100482.5 10037.5 100347.5 ;
      RECT  9972.5 100482.5 10037.5 100347.5 ;
      RECT  9782.5 100482.5 9847.5 100347.5 ;
      RECT  9972.5 100482.5 10037.5 100347.5 ;
      RECT  10162.5 100482.5 10227.5 100347.5 ;
      RECT  10162.5 100482.5 10227.5 100347.5 ;
      RECT  9972.5 100482.5 10037.5 100347.5 ;
      RECT  10332.5 99552.5 10397.5 99417.5 ;
      RECT  10332.5 100527.5 10397.5 100392.5 ;
      RECT  10167.5 100252.5 10032.5 100187.5 ;
      RECT  9910.0 100037.5 9775.0 99972.5 ;
      RECT  9972.5 99642.5 10037.5 99507.5 ;
      RECT  10162.5 100482.5 10227.5 100347.5 ;
      RECT  10262.5 100037.5 10127.5 99972.5 ;
      RECT  9775.0 100037.5 9910.0 99972.5 ;
      RECT  10032.5 100252.5 10167.5 100187.5 ;
      RECT  10127.5 100037.5 10262.5 99972.5 ;
      RECT  9715.0 99332.5 10635.0 99267.5 ;
      RECT  9715.0 100677.5 10635.0 100612.5 ;
      RECT  11062.5 99485.0 11127.5 99300.0 ;
      RECT  11062.5 100645.0 11127.5 100460.0 ;
      RECT  10702.5 100527.5 10767.5 100677.5 ;
      RECT  10702.5 99642.5 10767.5 99267.5 ;
      RECT  10892.5 100527.5 10957.5 99642.5 ;
      RECT  10702.5 99642.5 10767.5 99507.5 ;
      RECT  10892.5 99642.5 10957.5 99507.5 ;
      RECT  10892.5 99642.5 10957.5 99507.5 ;
      RECT  10702.5 99642.5 10767.5 99507.5 ;
      RECT  10702.5 100527.5 10767.5 100392.5 ;
      RECT  10892.5 100527.5 10957.5 100392.5 ;
      RECT  10892.5 100527.5 10957.5 100392.5 ;
      RECT  10702.5 100527.5 10767.5 100392.5 ;
      RECT  11062.5 99552.5 11127.5 99417.5 ;
      RECT  11062.5 100527.5 11127.5 100392.5 ;
      RECT  10760.0 100085.0 10825.0 99950.0 ;
      RECT  10760.0 100085.0 10825.0 99950.0 ;
      RECT  10925.0 100050.0 10990.0 99985.0 ;
      RECT  10635.0 99332.5 11195.0 99267.5 ;
      RECT  10635.0 100677.5 11195.0 100612.5 ;
      RECT  8897.5 99950.0 8962.5 100085.0 ;
      RECT  9037.5 100222.5 9102.5 100357.5 ;
      RECT  10032.5 100187.5 9897.5 100252.5 ;
      RECT  9582.5 101805.0 9647.5 101990.0 ;
      RECT  9582.5 100645.0 9647.5 100830.0 ;
      RECT  9222.5 100762.5 9287.5 100612.5 ;
      RECT  9222.5 101647.5 9287.5 102022.5 ;
      RECT  9412.5 100762.5 9477.5 101647.5 ;
      RECT  9222.5 101647.5 9287.5 101782.5 ;
      RECT  9412.5 101647.5 9477.5 101782.5 ;
      RECT  9412.5 101647.5 9477.5 101782.5 ;
      RECT  9222.5 101647.5 9287.5 101782.5 ;
      RECT  9222.5 100762.5 9287.5 100897.5 ;
      RECT  9412.5 100762.5 9477.5 100897.5 ;
      RECT  9412.5 100762.5 9477.5 100897.5 ;
      RECT  9222.5 100762.5 9287.5 100897.5 ;
      RECT  9582.5 101737.5 9647.5 101872.5 ;
      RECT  9582.5 100762.5 9647.5 100897.5 ;
      RECT  9280.0 101205.0 9345.0 101340.0 ;
      RECT  9280.0 101205.0 9345.0 101340.0 ;
      RECT  9445.0 101240.0 9510.0 101305.0 ;
      RECT  9155.0 101957.5 9715.0 102022.5 ;
      RECT  9155.0 100612.5 9715.0 100677.5 ;
      RECT  9782.5 100807.5 9847.5 100612.5 ;
      RECT  9782.5 101647.5 9847.5 102022.5 ;
      RECT  10162.5 101647.5 10227.5 102022.5 ;
      RECT  10332.5 101805.0 10397.5 101990.0 ;
      RECT  10332.5 100645.0 10397.5 100830.0 ;
      RECT  9782.5 101647.5 9847.5 101782.5 ;
      RECT  9972.5 101647.5 10037.5 101782.5 ;
      RECT  9972.5 101647.5 10037.5 101782.5 ;
      RECT  9782.5 101647.5 9847.5 101782.5 ;
      RECT  9972.5 101647.5 10037.5 101782.5 ;
      RECT  10162.5 101647.5 10227.5 101782.5 ;
      RECT  10162.5 101647.5 10227.5 101782.5 ;
      RECT  9972.5 101647.5 10037.5 101782.5 ;
      RECT  9782.5 100807.5 9847.5 100942.5 ;
      RECT  9972.5 100807.5 10037.5 100942.5 ;
      RECT  9972.5 100807.5 10037.5 100942.5 ;
      RECT  9782.5 100807.5 9847.5 100942.5 ;
      RECT  9972.5 100807.5 10037.5 100942.5 ;
      RECT  10162.5 100807.5 10227.5 100942.5 ;
      RECT  10162.5 100807.5 10227.5 100942.5 ;
      RECT  9972.5 100807.5 10037.5 100942.5 ;
      RECT  10332.5 101737.5 10397.5 101872.5 ;
      RECT  10332.5 100762.5 10397.5 100897.5 ;
      RECT  10167.5 101037.5 10032.5 101102.5 ;
      RECT  9910.0 101252.5 9775.0 101317.5 ;
      RECT  9972.5 101647.5 10037.5 101782.5 ;
      RECT  10162.5 100807.5 10227.5 100942.5 ;
      RECT  10262.5 101252.5 10127.5 101317.5 ;
      RECT  9775.0 101252.5 9910.0 101317.5 ;
      RECT  10032.5 101037.5 10167.5 101102.5 ;
      RECT  10127.5 101252.5 10262.5 101317.5 ;
      RECT  9715.0 101957.5 10635.0 102022.5 ;
      RECT  9715.0 100612.5 10635.0 100677.5 ;
      RECT  11062.5 101805.0 11127.5 101990.0 ;
      RECT  11062.5 100645.0 11127.5 100830.0 ;
      RECT  10702.5 100762.5 10767.5 100612.5 ;
      RECT  10702.5 101647.5 10767.5 102022.5 ;
      RECT  10892.5 100762.5 10957.5 101647.5 ;
      RECT  10702.5 101647.5 10767.5 101782.5 ;
      RECT  10892.5 101647.5 10957.5 101782.5 ;
      RECT  10892.5 101647.5 10957.5 101782.5 ;
      RECT  10702.5 101647.5 10767.5 101782.5 ;
      RECT  10702.5 100762.5 10767.5 100897.5 ;
      RECT  10892.5 100762.5 10957.5 100897.5 ;
      RECT  10892.5 100762.5 10957.5 100897.5 ;
      RECT  10702.5 100762.5 10767.5 100897.5 ;
      RECT  11062.5 101737.5 11127.5 101872.5 ;
      RECT  11062.5 100762.5 11127.5 100897.5 ;
      RECT  10760.0 101205.0 10825.0 101340.0 ;
      RECT  10760.0 101205.0 10825.0 101340.0 ;
      RECT  10925.0 101240.0 10990.0 101305.0 ;
      RECT  10635.0 101957.5 11195.0 102022.5 ;
      RECT  10635.0 100612.5 11195.0 100677.5 ;
      RECT  8897.5 101205.0 8962.5 101340.0 ;
      RECT  9037.5 100932.5 9102.5 101067.5 ;
      RECT  10032.5 101037.5 9897.5 101102.5 ;
      RECT  9582.5 102175.0 9647.5 101990.0 ;
      RECT  9582.5 103335.0 9647.5 103150.0 ;
      RECT  9222.5 103217.5 9287.5 103367.5 ;
      RECT  9222.5 102332.5 9287.5 101957.5 ;
      RECT  9412.5 103217.5 9477.5 102332.5 ;
      RECT  9222.5 102332.5 9287.5 102197.5 ;
      RECT  9412.5 102332.5 9477.5 102197.5 ;
      RECT  9412.5 102332.5 9477.5 102197.5 ;
      RECT  9222.5 102332.5 9287.5 102197.5 ;
      RECT  9222.5 103217.5 9287.5 103082.5 ;
      RECT  9412.5 103217.5 9477.5 103082.5 ;
      RECT  9412.5 103217.5 9477.5 103082.5 ;
      RECT  9222.5 103217.5 9287.5 103082.5 ;
      RECT  9582.5 102242.5 9647.5 102107.5 ;
      RECT  9582.5 103217.5 9647.5 103082.5 ;
      RECT  9280.0 102775.0 9345.0 102640.0 ;
      RECT  9280.0 102775.0 9345.0 102640.0 ;
      RECT  9445.0 102740.0 9510.0 102675.0 ;
      RECT  9155.0 102022.5 9715.0 101957.5 ;
      RECT  9155.0 103367.5 9715.0 103302.5 ;
      RECT  9782.5 103172.5 9847.5 103367.5 ;
      RECT  9782.5 102332.5 9847.5 101957.5 ;
      RECT  10162.5 102332.5 10227.5 101957.5 ;
      RECT  10332.5 102175.0 10397.5 101990.0 ;
      RECT  10332.5 103335.0 10397.5 103150.0 ;
      RECT  9782.5 102332.5 9847.5 102197.5 ;
      RECT  9972.5 102332.5 10037.5 102197.5 ;
      RECT  9972.5 102332.5 10037.5 102197.5 ;
      RECT  9782.5 102332.5 9847.5 102197.5 ;
      RECT  9972.5 102332.5 10037.5 102197.5 ;
      RECT  10162.5 102332.5 10227.5 102197.5 ;
      RECT  10162.5 102332.5 10227.5 102197.5 ;
      RECT  9972.5 102332.5 10037.5 102197.5 ;
      RECT  9782.5 103172.5 9847.5 103037.5 ;
      RECT  9972.5 103172.5 10037.5 103037.5 ;
      RECT  9972.5 103172.5 10037.5 103037.5 ;
      RECT  9782.5 103172.5 9847.5 103037.5 ;
      RECT  9972.5 103172.5 10037.5 103037.5 ;
      RECT  10162.5 103172.5 10227.5 103037.5 ;
      RECT  10162.5 103172.5 10227.5 103037.5 ;
      RECT  9972.5 103172.5 10037.5 103037.5 ;
      RECT  10332.5 102242.5 10397.5 102107.5 ;
      RECT  10332.5 103217.5 10397.5 103082.5 ;
      RECT  10167.5 102942.5 10032.5 102877.5 ;
      RECT  9910.0 102727.5 9775.0 102662.5 ;
      RECT  9972.5 102332.5 10037.5 102197.5 ;
      RECT  10162.5 103172.5 10227.5 103037.5 ;
      RECT  10262.5 102727.5 10127.5 102662.5 ;
      RECT  9775.0 102727.5 9910.0 102662.5 ;
      RECT  10032.5 102942.5 10167.5 102877.5 ;
      RECT  10127.5 102727.5 10262.5 102662.5 ;
      RECT  9715.0 102022.5 10635.0 101957.5 ;
      RECT  9715.0 103367.5 10635.0 103302.5 ;
      RECT  11062.5 102175.0 11127.5 101990.0 ;
      RECT  11062.5 103335.0 11127.5 103150.0 ;
      RECT  10702.5 103217.5 10767.5 103367.5 ;
      RECT  10702.5 102332.5 10767.5 101957.5 ;
      RECT  10892.5 103217.5 10957.5 102332.5 ;
      RECT  10702.5 102332.5 10767.5 102197.5 ;
      RECT  10892.5 102332.5 10957.5 102197.5 ;
      RECT  10892.5 102332.5 10957.5 102197.5 ;
      RECT  10702.5 102332.5 10767.5 102197.5 ;
      RECT  10702.5 103217.5 10767.5 103082.5 ;
      RECT  10892.5 103217.5 10957.5 103082.5 ;
      RECT  10892.5 103217.5 10957.5 103082.5 ;
      RECT  10702.5 103217.5 10767.5 103082.5 ;
      RECT  11062.5 102242.5 11127.5 102107.5 ;
      RECT  11062.5 103217.5 11127.5 103082.5 ;
      RECT  10760.0 102775.0 10825.0 102640.0 ;
      RECT  10760.0 102775.0 10825.0 102640.0 ;
      RECT  10925.0 102740.0 10990.0 102675.0 ;
      RECT  10635.0 102022.5 11195.0 101957.5 ;
      RECT  10635.0 103367.5 11195.0 103302.5 ;
      RECT  8897.5 102640.0 8962.5 102775.0 ;
      RECT  9037.5 102912.5 9102.5 103047.5 ;
      RECT  10032.5 102877.5 9897.5 102942.5 ;
      RECT  9582.5 104495.0 9647.5 104680.0 ;
      RECT  9582.5 103335.0 9647.5 103520.0 ;
      RECT  9222.5 103452.5 9287.5 103302.5 ;
      RECT  9222.5 104337.5 9287.5 104712.5 ;
      RECT  9412.5 103452.5 9477.5 104337.5 ;
      RECT  9222.5 104337.5 9287.5 104472.5 ;
      RECT  9412.5 104337.5 9477.5 104472.5 ;
      RECT  9412.5 104337.5 9477.5 104472.5 ;
      RECT  9222.5 104337.5 9287.5 104472.5 ;
      RECT  9222.5 103452.5 9287.5 103587.5 ;
      RECT  9412.5 103452.5 9477.5 103587.5 ;
      RECT  9412.5 103452.5 9477.5 103587.5 ;
      RECT  9222.5 103452.5 9287.5 103587.5 ;
      RECT  9582.5 104427.5 9647.5 104562.5 ;
      RECT  9582.5 103452.5 9647.5 103587.5 ;
      RECT  9280.0 103895.0 9345.0 104030.0 ;
      RECT  9280.0 103895.0 9345.0 104030.0 ;
      RECT  9445.0 103930.0 9510.0 103995.0 ;
      RECT  9155.0 104647.5 9715.0 104712.5 ;
      RECT  9155.0 103302.5 9715.0 103367.5 ;
      RECT  9782.5 103497.5 9847.5 103302.5 ;
      RECT  9782.5 104337.5 9847.5 104712.5 ;
      RECT  10162.5 104337.5 10227.5 104712.5 ;
      RECT  10332.5 104495.0 10397.5 104680.0 ;
      RECT  10332.5 103335.0 10397.5 103520.0 ;
      RECT  9782.5 104337.5 9847.5 104472.5 ;
      RECT  9972.5 104337.5 10037.5 104472.5 ;
      RECT  9972.5 104337.5 10037.5 104472.5 ;
      RECT  9782.5 104337.5 9847.5 104472.5 ;
      RECT  9972.5 104337.5 10037.5 104472.5 ;
      RECT  10162.5 104337.5 10227.5 104472.5 ;
      RECT  10162.5 104337.5 10227.5 104472.5 ;
      RECT  9972.5 104337.5 10037.5 104472.5 ;
      RECT  9782.5 103497.5 9847.5 103632.5 ;
      RECT  9972.5 103497.5 10037.5 103632.5 ;
      RECT  9972.5 103497.5 10037.5 103632.5 ;
      RECT  9782.5 103497.5 9847.5 103632.5 ;
      RECT  9972.5 103497.5 10037.5 103632.5 ;
      RECT  10162.5 103497.5 10227.5 103632.5 ;
      RECT  10162.5 103497.5 10227.5 103632.5 ;
      RECT  9972.5 103497.5 10037.5 103632.5 ;
      RECT  10332.5 104427.5 10397.5 104562.5 ;
      RECT  10332.5 103452.5 10397.5 103587.5 ;
      RECT  10167.5 103727.5 10032.5 103792.5 ;
      RECT  9910.0 103942.5 9775.0 104007.5 ;
      RECT  9972.5 104337.5 10037.5 104472.5 ;
      RECT  10162.5 103497.5 10227.5 103632.5 ;
      RECT  10262.5 103942.5 10127.5 104007.5 ;
      RECT  9775.0 103942.5 9910.0 104007.5 ;
      RECT  10032.5 103727.5 10167.5 103792.5 ;
      RECT  10127.5 103942.5 10262.5 104007.5 ;
      RECT  9715.0 104647.5 10635.0 104712.5 ;
      RECT  9715.0 103302.5 10635.0 103367.5 ;
      RECT  11062.5 104495.0 11127.5 104680.0 ;
      RECT  11062.5 103335.0 11127.5 103520.0 ;
      RECT  10702.5 103452.5 10767.5 103302.5 ;
      RECT  10702.5 104337.5 10767.5 104712.5 ;
      RECT  10892.5 103452.5 10957.5 104337.5 ;
      RECT  10702.5 104337.5 10767.5 104472.5 ;
      RECT  10892.5 104337.5 10957.5 104472.5 ;
      RECT  10892.5 104337.5 10957.5 104472.5 ;
      RECT  10702.5 104337.5 10767.5 104472.5 ;
      RECT  10702.5 103452.5 10767.5 103587.5 ;
      RECT  10892.5 103452.5 10957.5 103587.5 ;
      RECT  10892.5 103452.5 10957.5 103587.5 ;
      RECT  10702.5 103452.5 10767.5 103587.5 ;
      RECT  11062.5 104427.5 11127.5 104562.5 ;
      RECT  11062.5 103452.5 11127.5 103587.5 ;
      RECT  10760.0 103895.0 10825.0 104030.0 ;
      RECT  10760.0 103895.0 10825.0 104030.0 ;
      RECT  10925.0 103930.0 10990.0 103995.0 ;
      RECT  10635.0 104647.5 11195.0 104712.5 ;
      RECT  10635.0 103302.5 11195.0 103367.5 ;
      RECT  8897.5 103895.0 8962.5 104030.0 ;
      RECT  9037.5 103622.5 9102.5 103757.5 ;
      RECT  10032.5 103727.5 9897.5 103792.5 ;
      RECT  9582.5 104865.0 9647.5 104680.0 ;
      RECT  9582.5 106025.0 9647.5 105840.0 ;
      RECT  9222.5 105907.5 9287.5 106057.5 ;
      RECT  9222.5 105022.5 9287.5 104647.5 ;
      RECT  9412.5 105907.5 9477.5 105022.5 ;
      RECT  9222.5 105022.5 9287.5 104887.5 ;
      RECT  9412.5 105022.5 9477.5 104887.5 ;
      RECT  9412.5 105022.5 9477.5 104887.5 ;
      RECT  9222.5 105022.5 9287.5 104887.5 ;
      RECT  9222.5 105907.5 9287.5 105772.5 ;
      RECT  9412.5 105907.5 9477.5 105772.5 ;
      RECT  9412.5 105907.5 9477.5 105772.5 ;
      RECT  9222.5 105907.5 9287.5 105772.5 ;
      RECT  9582.5 104932.5 9647.5 104797.5 ;
      RECT  9582.5 105907.5 9647.5 105772.5 ;
      RECT  9280.0 105465.0 9345.0 105330.0 ;
      RECT  9280.0 105465.0 9345.0 105330.0 ;
      RECT  9445.0 105430.0 9510.0 105365.0 ;
      RECT  9155.0 104712.5 9715.0 104647.5 ;
      RECT  9155.0 106057.5 9715.0 105992.5 ;
      RECT  9782.5 105862.5 9847.5 106057.5 ;
      RECT  9782.5 105022.5 9847.5 104647.5 ;
      RECT  10162.5 105022.5 10227.5 104647.5 ;
      RECT  10332.5 104865.0 10397.5 104680.0 ;
      RECT  10332.5 106025.0 10397.5 105840.0 ;
      RECT  9782.5 105022.5 9847.5 104887.5 ;
      RECT  9972.5 105022.5 10037.5 104887.5 ;
      RECT  9972.5 105022.5 10037.5 104887.5 ;
      RECT  9782.5 105022.5 9847.5 104887.5 ;
      RECT  9972.5 105022.5 10037.5 104887.5 ;
      RECT  10162.5 105022.5 10227.5 104887.5 ;
      RECT  10162.5 105022.5 10227.5 104887.5 ;
      RECT  9972.5 105022.5 10037.5 104887.5 ;
      RECT  9782.5 105862.5 9847.5 105727.5 ;
      RECT  9972.5 105862.5 10037.5 105727.5 ;
      RECT  9972.5 105862.5 10037.5 105727.5 ;
      RECT  9782.5 105862.5 9847.5 105727.5 ;
      RECT  9972.5 105862.5 10037.5 105727.5 ;
      RECT  10162.5 105862.5 10227.5 105727.5 ;
      RECT  10162.5 105862.5 10227.5 105727.5 ;
      RECT  9972.5 105862.5 10037.5 105727.5 ;
      RECT  10332.5 104932.5 10397.5 104797.5 ;
      RECT  10332.5 105907.5 10397.5 105772.5 ;
      RECT  10167.5 105632.5 10032.5 105567.5 ;
      RECT  9910.0 105417.5 9775.0 105352.5 ;
      RECT  9972.5 105022.5 10037.5 104887.5 ;
      RECT  10162.5 105862.5 10227.5 105727.5 ;
      RECT  10262.5 105417.5 10127.5 105352.5 ;
      RECT  9775.0 105417.5 9910.0 105352.5 ;
      RECT  10032.5 105632.5 10167.5 105567.5 ;
      RECT  10127.5 105417.5 10262.5 105352.5 ;
      RECT  9715.0 104712.5 10635.0 104647.5 ;
      RECT  9715.0 106057.5 10635.0 105992.5 ;
      RECT  11062.5 104865.0 11127.5 104680.0 ;
      RECT  11062.5 106025.0 11127.5 105840.0 ;
      RECT  10702.5 105907.5 10767.5 106057.5 ;
      RECT  10702.5 105022.5 10767.5 104647.5 ;
      RECT  10892.5 105907.5 10957.5 105022.5 ;
      RECT  10702.5 105022.5 10767.5 104887.5 ;
      RECT  10892.5 105022.5 10957.5 104887.5 ;
      RECT  10892.5 105022.5 10957.5 104887.5 ;
      RECT  10702.5 105022.5 10767.5 104887.5 ;
      RECT  10702.5 105907.5 10767.5 105772.5 ;
      RECT  10892.5 105907.5 10957.5 105772.5 ;
      RECT  10892.5 105907.5 10957.5 105772.5 ;
      RECT  10702.5 105907.5 10767.5 105772.5 ;
      RECT  11062.5 104932.5 11127.5 104797.5 ;
      RECT  11062.5 105907.5 11127.5 105772.5 ;
      RECT  10760.0 105465.0 10825.0 105330.0 ;
      RECT  10760.0 105465.0 10825.0 105330.0 ;
      RECT  10925.0 105430.0 10990.0 105365.0 ;
      RECT  10635.0 104712.5 11195.0 104647.5 ;
      RECT  10635.0 106057.5 11195.0 105992.5 ;
      RECT  8897.5 105330.0 8962.5 105465.0 ;
      RECT  9037.5 105602.5 9102.5 105737.5 ;
      RECT  10032.5 105567.5 9897.5 105632.5 ;
      RECT  9582.5 107185.0 9647.5 107370.0 ;
      RECT  9582.5 106025.0 9647.5 106210.0 ;
      RECT  9222.5 106142.5 9287.5 105992.5 ;
      RECT  9222.5 107027.5 9287.5 107402.5 ;
      RECT  9412.5 106142.5 9477.5 107027.5 ;
      RECT  9222.5 107027.5 9287.5 107162.5 ;
      RECT  9412.5 107027.5 9477.5 107162.5 ;
      RECT  9412.5 107027.5 9477.5 107162.5 ;
      RECT  9222.5 107027.5 9287.5 107162.5 ;
      RECT  9222.5 106142.5 9287.5 106277.5 ;
      RECT  9412.5 106142.5 9477.5 106277.5 ;
      RECT  9412.5 106142.5 9477.5 106277.5 ;
      RECT  9222.5 106142.5 9287.5 106277.5 ;
      RECT  9582.5 107117.5 9647.5 107252.5 ;
      RECT  9582.5 106142.5 9647.5 106277.5 ;
      RECT  9280.0 106585.0 9345.0 106720.0 ;
      RECT  9280.0 106585.0 9345.0 106720.0 ;
      RECT  9445.0 106620.0 9510.0 106685.0 ;
      RECT  9155.0 107337.5 9715.0 107402.5 ;
      RECT  9155.0 105992.5 9715.0 106057.5 ;
      RECT  9782.5 106187.5 9847.5 105992.5 ;
      RECT  9782.5 107027.5 9847.5 107402.5 ;
      RECT  10162.5 107027.5 10227.5 107402.5 ;
      RECT  10332.5 107185.0 10397.5 107370.0 ;
      RECT  10332.5 106025.0 10397.5 106210.0 ;
      RECT  9782.5 107027.5 9847.5 107162.5 ;
      RECT  9972.5 107027.5 10037.5 107162.5 ;
      RECT  9972.5 107027.5 10037.5 107162.5 ;
      RECT  9782.5 107027.5 9847.5 107162.5 ;
      RECT  9972.5 107027.5 10037.5 107162.5 ;
      RECT  10162.5 107027.5 10227.5 107162.5 ;
      RECT  10162.5 107027.5 10227.5 107162.5 ;
      RECT  9972.5 107027.5 10037.5 107162.5 ;
      RECT  9782.5 106187.5 9847.5 106322.5 ;
      RECT  9972.5 106187.5 10037.5 106322.5 ;
      RECT  9972.5 106187.5 10037.5 106322.5 ;
      RECT  9782.5 106187.5 9847.5 106322.5 ;
      RECT  9972.5 106187.5 10037.5 106322.5 ;
      RECT  10162.5 106187.5 10227.5 106322.5 ;
      RECT  10162.5 106187.5 10227.5 106322.5 ;
      RECT  9972.5 106187.5 10037.5 106322.5 ;
      RECT  10332.5 107117.5 10397.5 107252.5 ;
      RECT  10332.5 106142.5 10397.5 106277.5 ;
      RECT  10167.5 106417.5 10032.5 106482.5 ;
      RECT  9910.0 106632.5 9775.0 106697.5 ;
      RECT  9972.5 107027.5 10037.5 107162.5 ;
      RECT  10162.5 106187.5 10227.5 106322.5 ;
      RECT  10262.5 106632.5 10127.5 106697.5 ;
      RECT  9775.0 106632.5 9910.0 106697.5 ;
      RECT  10032.5 106417.5 10167.5 106482.5 ;
      RECT  10127.5 106632.5 10262.5 106697.5 ;
      RECT  9715.0 107337.5 10635.0 107402.5 ;
      RECT  9715.0 105992.5 10635.0 106057.5 ;
      RECT  11062.5 107185.0 11127.5 107370.0 ;
      RECT  11062.5 106025.0 11127.5 106210.0 ;
      RECT  10702.5 106142.5 10767.5 105992.5 ;
      RECT  10702.5 107027.5 10767.5 107402.5 ;
      RECT  10892.5 106142.5 10957.5 107027.5 ;
      RECT  10702.5 107027.5 10767.5 107162.5 ;
      RECT  10892.5 107027.5 10957.5 107162.5 ;
      RECT  10892.5 107027.5 10957.5 107162.5 ;
      RECT  10702.5 107027.5 10767.5 107162.5 ;
      RECT  10702.5 106142.5 10767.5 106277.5 ;
      RECT  10892.5 106142.5 10957.5 106277.5 ;
      RECT  10892.5 106142.5 10957.5 106277.5 ;
      RECT  10702.5 106142.5 10767.5 106277.5 ;
      RECT  11062.5 107117.5 11127.5 107252.5 ;
      RECT  11062.5 106142.5 11127.5 106277.5 ;
      RECT  10760.0 106585.0 10825.0 106720.0 ;
      RECT  10760.0 106585.0 10825.0 106720.0 ;
      RECT  10925.0 106620.0 10990.0 106685.0 ;
      RECT  10635.0 107337.5 11195.0 107402.5 ;
      RECT  10635.0 105992.5 11195.0 106057.5 ;
      RECT  8897.5 106585.0 8962.5 106720.0 ;
      RECT  9037.5 106312.5 9102.5 106447.5 ;
      RECT  10032.5 106417.5 9897.5 106482.5 ;
      RECT  9582.5 107555.0 9647.5 107370.0 ;
      RECT  9582.5 108715.0 9647.5 108530.0 ;
      RECT  9222.5 108597.5 9287.5 108747.5 ;
      RECT  9222.5 107712.5 9287.5 107337.5 ;
      RECT  9412.5 108597.5 9477.5 107712.5 ;
      RECT  9222.5 107712.5 9287.5 107577.5 ;
      RECT  9412.5 107712.5 9477.5 107577.5 ;
      RECT  9412.5 107712.5 9477.5 107577.5 ;
      RECT  9222.5 107712.5 9287.5 107577.5 ;
      RECT  9222.5 108597.5 9287.5 108462.5 ;
      RECT  9412.5 108597.5 9477.5 108462.5 ;
      RECT  9412.5 108597.5 9477.5 108462.5 ;
      RECT  9222.5 108597.5 9287.5 108462.5 ;
      RECT  9582.5 107622.5 9647.5 107487.5 ;
      RECT  9582.5 108597.5 9647.5 108462.5 ;
      RECT  9280.0 108155.0 9345.0 108020.0 ;
      RECT  9280.0 108155.0 9345.0 108020.0 ;
      RECT  9445.0 108120.0 9510.0 108055.0 ;
      RECT  9155.0 107402.5 9715.0 107337.5 ;
      RECT  9155.0 108747.5 9715.0 108682.5 ;
      RECT  9782.5 108552.5 9847.5 108747.5 ;
      RECT  9782.5 107712.5 9847.5 107337.5 ;
      RECT  10162.5 107712.5 10227.5 107337.5 ;
      RECT  10332.5 107555.0 10397.5 107370.0 ;
      RECT  10332.5 108715.0 10397.5 108530.0 ;
      RECT  9782.5 107712.5 9847.5 107577.5 ;
      RECT  9972.5 107712.5 10037.5 107577.5 ;
      RECT  9972.5 107712.5 10037.5 107577.5 ;
      RECT  9782.5 107712.5 9847.5 107577.5 ;
      RECT  9972.5 107712.5 10037.5 107577.5 ;
      RECT  10162.5 107712.5 10227.5 107577.5 ;
      RECT  10162.5 107712.5 10227.5 107577.5 ;
      RECT  9972.5 107712.5 10037.5 107577.5 ;
      RECT  9782.5 108552.5 9847.5 108417.5 ;
      RECT  9972.5 108552.5 10037.5 108417.5 ;
      RECT  9972.5 108552.5 10037.5 108417.5 ;
      RECT  9782.5 108552.5 9847.5 108417.5 ;
      RECT  9972.5 108552.5 10037.5 108417.5 ;
      RECT  10162.5 108552.5 10227.5 108417.5 ;
      RECT  10162.5 108552.5 10227.5 108417.5 ;
      RECT  9972.5 108552.5 10037.5 108417.5 ;
      RECT  10332.5 107622.5 10397.5 107487.5 ;
      RECT  10332.5 108597.5 10397.5 108462.5 ;
      RECT  10167.5 108322.5 10032.5 108257.5 ;
      RECT  9910.0 108107.5 9775.0 108042.5 ;
      RECT  9972.5 107712.5 10037.5 107577.5 ;
      RECT  10162.5 108552.5 10227.5 108417.5 ;
      RECT  10262.5 108107.5 10127.5 108042.5 ;
      RECT  9775.0 108107.5 9910.0 108042.5 ;
      RECT  10032.5 108322.5 10167.5 108257.5 ;
      RECT  10127.5 108107.5 10262.5 108042.5 ;
      RECT  9715.0 107402.5 10635.0 107337.5 ;
      RECT  9715.0 108747.5 10635.0 108682.5 ;
      RECT  11062.5 107555.0 11127.5 107370.0 ;
      RECT  11062.5 108715.0 11127.5 108530.0 ;
      RECT  10702.5 108597.5 10767.5 108747.5 ;
      RECT  10702.5 107712.5 10767.5 107337.5 ;
      RECT  10892.5 108597.5 10957.5 107712.5 ;
      RECT  10702.5 107712.5 10767.5 107577.5 ;
      RECT  10892.5 107712.5 10957.5 107577.5 ;
      RECT  10892.5 107712.5 10957.5 107577.5 ;
      RECT  10702.5 107712.5 10767.5 107577.5 ;
      RECT  10702.5 108597.5 10767.5 108462.5 ;
      RECT  10892.5 108597.5 10957.5 108462.5 ;
      RECT  10892.5 108597.5 10957.5 108462.5 ;
      RECT  10702.5 108597.5 10767.5 108462.5 ;
      RECT  11062.5 107622.5 11127.5 107487.5 ;
      RECT  11062.5 108597.5 11127.5 108462.5 ;
      RECT  10760.0 108155.0 10825.0 108020.0 ;
      RECT  10760.0 108155.0 10825.0 108020.0 ;
      RECT  10925.0 108120.0 10990.0 108055.0 ;
      RECT  10635.0 107402.5 11195.0 107337.5 ;
      RECT  10635.0 108747.5 11195.0 108682.5 ;
      RECT  8897.5 108020.0 8962.5 108155.0 ;
      RECT  9037.5 108292.5 9102.5 108427.5 ;
      RECT  10032.5 108257.5 9897.5 108322.5 ;
      RECT  9582.5 109875.0 9647.5 110060.0 ;
      RECT  9582.5 108715.0 9647.5 108900.0 ;
      RECT  9222.5 108832.5 9287.5 108682.5 ;
      RECT  9222.5 109717.5 9287.5 110092.5 ;
      RECT  9412.5 108832.5 9477.5 109717.5 ;
      RECT  9222.5 109717.5 9287.5 109852.5 ;
      RECT  9412.5 109717.5 9477.5 109852.5 ;
      RECT  9412.5 109717.5 9477.5 109852.5 ;
      RECT  9222.5 109717.5 9287.5 109852.5 ;
      RECT  9222.5 108832.5 9287.5 108967.5 ;
      RECT  9412.5 108832.5 9477.5 108967.5 ;
      RECT  9412.5 108832.5 9477.5 108967.5 ;
      RECT  9222.5 108832.5 9287.5 108967.5 ;
      RECT  9582.5 109807.5 9647.5 109942.5 ;
      RECT  9582.5 108832.5 9647.5 108967.5 ;
      RECT  9280.0 109275.0 9345.0 109410.0 ;
      RECT  9280.0 109275.0 9345.0 109410.0 ;
      RECT  9445.0 109310.0 9510.0 109375.0 ;
      RECT  9155.0 110027.5 9715.0 110092.5 ;
      RECT  9155.0 108682.5 9715.0 108747.5 ;
      RECT  9782.5 108877.5 9847.5 108682.5 ;
      RECT  9782.5 109717.5 9847.5 110092.5 ;
      RECT  10162.5 109717.5 10227.5 110092.5 ;
      RECT  10332.5 109875.0 10397.5 110060.0 ;
      RECT  10332.5 108715.0 10397.5 108900.0 ;
      RECT  9782.5 109717.5 9847.5 109852.5 ;
      RECT  9972.5 109717.5 10037.5 109852.5 ;
      RECT  9972.5 109717.5 10037.5 109852.5 ;
      RECT  9782.5 109717.5 9847.5 109852.5 ;
      RECT  9972.5 109717.5 10037.5 109852.5 ;
      RECT  10162.5 109717.5 10227.5 109852.5 ;
      RECT  10162.5 109717.5 10227.5 109852.5 ;
      RECT  9972.5 109717.5 10037.5 109852.5 ;
      RECT  9782.5 108877.5 9847.5 109012.5 ;
      RECT  9972.5 108877.5 10037.5 109012.5 ;
      RECT  9972.5 108877.5 10037.5 109012.5 ;
      RECT  9782.5 108877.5 9847.5 109012.5 ;
      RECT  9972.5 108877.5 10037.5 109012.5 ;
      RECT  10162.5 108877.5 10227.5 109012.5 ;
      RECT  10162.5 108877.5 10227.5 109012.5 ;
      RECT  9972.5 108877.5 10037.5 109012.5 ;
      RECT  10332.5 109807.5 10397.5 109942.5 ;
      RECT  10332.5 108832.5 10397.5 108967.5 ;
      RECT  10167.5 109107.5 10032.5 109172.5 ;
      RECT  9910.0 109322.5 9775.0 109387.5 ;
      RECT  9972.5 109717.5 10037.5 109852.5 ;
      RECT  10162.5 108877.5 10227.5 109012.5 ;
      RECT  10262.5 109322.5 10127.5 109387.5 ;
      RECT  9775.0 109322.5 9910.0 109387.5 ;
      RECT  10032.5 109107.5 10167.5 109172.5 ;
      RECT  10127.5 109322.5 10262.5 109387.5 ;
      RECT  9715.0 110027.5 10635.0 110092.5 ;
      RECT  9715.0 108682.5 10635.0 108747.5 ;
      RECT  11062.5 109875.0 11127.5 110060.0 ;
      RECT  11062.5 108715.0 11127.5 108900.0 ;
      RECT  10702.5 108832.5 10767.5 108682.5 ;
      RECT  10702.5 109717.5 10767.5 110092.5 ;
      RECT  10892.5 108832.5 10957.5 109717.5 ;
      RECT  10702.5 109717.5 10767.5 109852.5 ;
      RECT  10892.5 109717.5 10957.5 109852.5 ;
      RECT  10892.5 109717.5 10957.5 109852.5 ;
      RECT  10702.5 109717.5 10767.5 109852.5 ;
      RECT  10702.5 108832.5 10767.5 108967.5 ;
      RECT  10892.5 108832.5 10957.5 108967.5 ;
      RECT  10892.5 108832.5 10957.5 108967.5 ;
      RECT  10702.5 108832.5 10767.5 108967.5 ;
      RECT  11062.5 109807.5 11127.5 109942.5 ;
      RECT  11062.5 108832.5 11127.5 108967.5 ;
      RECT  10760.0 109275.0 10825.0 109410.0 ;
      RECT  10760.0 109275.0 10825.0 109410.0 ;
      RECT  10925.0 109310.0 10990.0 109375.0 ;
      RECT  10635.0 110027.5 11195.0 110092.5 ;
      RECT  10635.0 108682.5 11195.0 108747.5 ;
      RECT  8897.5 109275.0 8962.5 109410.0 ;
      RECT  9037.5 109002.5 9102.5 109137.5 ;
      RECT  10032.5 109107.5 9897.5 109172.5 ;
      RECT  9582.5 110245.0 9647.5 110060.0 ;
      RECT  9582.5 111405.0 9647.5 111220.0 ;
      RECT  9222.5 111287.5 9287.5 111437.5 ;
      RECT  9222.5 110402.5 9287.5 110027.5 ;
      RECT  9412.5 111287.5 9477.5 110402.5 ;
      RECT  9222.5 110402.5 9287.5 110267.5 ;
      RECT  9412.5 110402.5 9477.5 110267.5 ;
      RECT  9412.5 110402.5 9477.5 110267.5 ;
      RECT  9222.5 110402.5 9287.5 110267.5 ;
      RECT  9222.5 111287.5 9287.5 111152.5 ;
      RECT  9412.5 111287.5 9477.5 111152.5 ;
      RECT  9412.5 111287.5 9477.5 111152.5 ;
      RECT  9222.5 111287.5 9287.5 111152.5 ;
      RECT  9582.5 110312.5 9647.5 110177.5 ;
      RECT  9582.5 111287.5 9647.5 111152.5 ;
      RECT  9280.0 110845.0 9345.0 110710.0 ;
      RECT  9280.0 110845.0 9345.0 110710.0 ;
      RECT  9445.0 110810.0 9510.0 110745.0 ;
      RECT  9155.0 110092.5 9715.0 110027.5 ;
      RECT  9155.0 111437.5 9715.0 111372.5 ;
      RECT  9782.5 111242.5 9847.5 111437.5 ;
      RECT  9782.5 110402.5 9847.5 110027.5 ;
      RECT  10162.5 110402.5 10227.5 110027.5 ;
      RECT  10332.5 110245.0 10397.5 110060.0 ;
      RECT  10332.5 111405.0 10397.5 111220.0 ;
      RECT  9782.5 110402.5 9847.5 110267.5 ;
      RECT  9972.5 110402.5 10037.5 110267.5 ;
      RECT  9972.5 110402.5 10037.5 110267.5 ;
      RECT  9782.5 110402.5 9847.5 110267.5 ;
      RECT  9972.5 110402.5 10037.5 110267.5 ;
      RECT  10162.5 110402.5 10227.5 110267.5 ;
      RECT  10162.5 110402.5 10227.5 110267.5 ;
      RECT  9972.5 110402.5 10037.5 110267.5 ;
      RECT  9782.5 111242.5 9847.5 111107.5 ;
      RECT  9972.5 111242.5 10037.5 111107.5 ;
      RECT  9972.5 111242.5 10037.5 111107.5 ;
      RECT  9782.5 111242.5 9847.5 111107.5 ;
      RECT  9972.5 111242.5 10037.5 111107.5 ;
      RECT  10162.5 111242.5 10227.5 111107.5 ;
      RECT  10162.5 111242.5 10227.5 111107.5 ;
      RECT  9972.5 111242.5 10037.5 111107.5 ;
      RECT  10332.5 110312.5 10397.5 110177.5 ;
      RECT  10332.5 111287.5 10397.5 111152.5 ;
      RECT  10167.5 111012.5 10032.5 110947.5 ;
      RECT  9910.0 110797.5 9775.0 110732.5 ;
      RECT  9972.5 110402.5 10037.5 110267.5 ;
      RECT  10162.5 111242.5 10227.5 111107.5 ;
      RECT  10262.5 110797.5 10127.5 110732.5 ;
      RECT  9775.0 110797.5 9910.0 110732.5 ;
      RECT  10032.5 111012.5 10167.5 110947.5 ;
      RECT  10127.5 110797.5 10262.5 110732.5 ;
      RECT  9715.0 110092.5 10635.0 110027.5 ;
      RECT  9715.0 111437.5 10635.0 111372.5 ;
      RECT  11062.5 110245.0 11127.5 110060.0 ;
      RECT  11062.5 111405.0 11127.5 111220.0 ;
      RECT  10702.5 111287.5 10767.5 111437.5 ;
      RECT  10702.5 110402.5 10767.5 110027.5 ;
      RECT  10892.5 111287.5 10957.5 110402.5 ;
      RECT  10702.5 110402.5 10767.5 110267.5 ;
      RECT  10892.5 110402.5 10957.5 110267.5 ;
      RECT  10892.5 110402.5 10957.5 110267.5 ;
      RECT  10702.5 110402.5 10767.5 110267.5 ;
      RECT  10702.5 111287.5 10767.5 111152.5 ;
      RECT  10892.5 111287.5 10957.5 111152.5 ;
      RECT  10892.5 111287.5 10957.5 111152.5 ;
      RECT  10702.5 111287.5 10767.5 111152.5 ;
      RECT  11062.5 110312.5 11127.5 110177.5 ;
      RECT  11062.5 111287.5 11127.5 111152.5 ;
      RECT  10760.0 110845.0 10825.0 110710.0 ;
      RECT  10760.0 110845.0 10825.0 110710.0 ;
      RECT  10925.0 110810.0 10990.0 110745.0 ;
      RECT  10635.0 110092.5 11195.0 110027.5 ;
      RECT  10635.0 111437.5 11195.0 111372.5 ;
      RECT  8897.5 110710.0 8962.5 110845.0 ;
      RECT  9037.5 110982.5 9102.5 111117.5 ;
      RECT  10032.5 110947.5 9897.5 111012.5 ;
      RECT  9582.5 112565.0 9647.5 112750.0 ;
      RECT  9582.5 111405.0 9647.5 111590.0 ;
      RECT  9222.5 111522.5 9287.5 111372.5 ;
      RECT  9222.5 112407.5 9287.5 112782.5 ;
      RECT  9412.5 111522.5 9477.5 112407.5 ;
      RECT  9222.5 112407.5 9287.5 112542.5 ;
      RECT  9412.5 112407.5 9477.5 112542.5 ;
      RECT  9412.5 112407.5 9477.5 112542.5 ;
      RECT  9222.5 112407.5 9287.5 112542.5 ;
      RECT  9222.5 111522.5 9287.5 111657.5 ;
      RECT  9412.5 111522.5 9477.5 111657.5 ;
      RECT  9412.5 111522.5 9477.5 111657.5 ;
      RECT  9222.5 111522.5 9287.5 111657.5 ;
      RECT  9582.5 112497.5 9647.5 112632.5 ;
      RECT  9582.5 111522.5 9647.5 111657.5 ;
      RECT  9280.0 111965.0 9345.0 112100.0 ;
      RECT  9280.0 111965.0 9345.0 112100.0 ;
      RECT  9445.0 112000.0 9510.0 112065.0 ;
      RECT  9155.0 112717.5 9715.0 112782.5 ;
      RECT  9155.0 111372.5 9715.0 111437.5 ;
      RECT  9782.5 111567.5 9847.5 111372.5 ;
      RECT  9782.5 112407.5 9847.5 112782.5 ;
      RECT  10162.5 112407.5 10227.5 112782.5 ;
      RECT  10332.5 112565.0 10397.5 112750.0 ;
      RECT  10332.5 111405.0 10397.5 111590.0 ;
      RECT  9782.5 112407.5 9847.5 112542.5 ;
      RECT  9972.5 112407.5 10037.5 112542.5 ;
      RECT  9972.5 112407.5 10037.5 112542.5 ;
      RECT  9782.5 112407.5 9847.5 112542.5 ;
      RECT  9972.5 112407.5 10037.5 112542.5 ;
      RECT  10162.5 112407.5 10227.5 112542.5 ;
      RECT  10162.5 112407.5 10227.5 112542.5 ;
      RECT  9972.5 112407.5 10037.5 112542.5 ;
      RECT  9782.5 111567.5 9847.5 111702.5 ;
      RECT  9972.5 111567.5 10037.5 111702.5 ;
      RECT  9972.5 111567.5 10037.5 111702.5 ;
      RECT  9782.5 111567.5 9847.5 111702.5 ;
      RECT  9972.5 111567.5 10037.5 111702.5 ;
      RECT  10162.5 111567.5 10227.5 111702.5 ;
      RECT  10162.5 111567.5 10227.5 111702.5 ;
      RECT  9972.5 111567.5 10037.5 111702.5 ;
      RECT  10332.5 112497.5 10397.5 112632.5 ;
      RECT  10332.5 111522.5 10397.5 111657.5 ;
      RECT  10167.5 111797.5 10032.5 111862.5 ;
      RECT  9910.0 112012.5 9775.0 112077.5 ;
      RECT  9972.5 112407.5 10037.5 112542.5 ;
      RECT  10162.5 111567.5 10227.5 111702.5 ;
      RECT  10262.5 112012.5 10127.5 112077.5 ;
      RECT  9775.0 112012.5 9910.0 112077.5 ;
      RECT  10032.5 111797.5 10167.5 111862.5 ;
      RECT  10127.5 112012.5 10262.5 112077.5 ;
      RECT  9715.0 112717.5 10635.0 112782.5 ;
      RECT  9715.0 111372.5 10635.0 111437.5 ;
      RECT  11062.5 112565.0 11127.5 112750.0 ;
      RECT  11062.5 111405.0 11127.5 111590.0 ;
      RECT  10702.5 111522.5 10767.5 111372.5 ;
      RECT  10702.5 112407.5 10767.5 112782.5 ;
      RECT  10892.5 111522.5 10957.5 112407.5 ;
      RECT  10702.5 112407.5 10767.5 112542.5 ;
      RECT  10892.5 112407.5 10957.5 112542.5 ;
      RECT  10892.5 112407.5 10957.5 112542.5 ;
      RECT  10702.5 112407.5 10767.5 112542.5 ;
      RECT  10702.5 111522.5 10767.5 111657.5 ;
      RECT  10892.5 111522.5 10957.5 111657.5 ;
      RECT  10892.5 111522.5 10957.5 111657.5 ;
      RECT  10702.5 111522.5 10767.5 111657.5 ;
      RECT  11062.5 112497.5 11127.5 112632.5 ;
      RECT  11062.5 111522.5 11127.5 111657.5 ;
      RECT  10760.0 111965.0 10825.0 112100.0 ;
      RECT  10760.0 111965.0 10825.0 112100.0 ;
      RECT  10925.0 112000.0 10990.0 112065.0 ;
      RECT  10635.0 112717.5 11195.0 112782.5 ;
      RECT  10635.0 111372.5 11195.0 111437.5 ;
      RECT  8897.5 111965.0 8962.5 112100.0 ;
      RECT  9037.5 111692.5 9102.5 111827.5 ;
      RECT  10032.5 111797.5 9897.5 111862.5 ;
      RECT  9582.5 112935.0 9647.5 112750.0 ;
      RECT  9582.5 114095.0 9647.5 113910.0 ;
      RECT  9222.5 113977.5 9287.5 114127.5 ;
      RECT  9222.5 113092.5 9287.5 112717.5 ;
      RECT  9412.5 113977.5 9477.5 113092.5 ;
      RECT  9222.5 113092.5 9287.5 112957.5 ;
      RECT  9412.5 113092.5 9477.5 112957.5 ;
      RECT  9412.5 113092.5 9477.5 112957.5 ;
      RECT  9222.5 113092.5 9287.5 112957.5 ;
      RECT  9222.5 113977.5 9287.5 113842.5 ;
      RECT  9412.5 113977.5 9477.5 113842.5 ;
      RECT  9412.5 113977.5 9477.5 113842.5 ;
      RECT  9222.5 113977.5 9287.5 113842.5 ;
      RECT  9582.5 113002.5 9647.5 112867.5 ;
      RECT  9582.5 113977.5 9647.5 113842.5 ;
      RECT  9280.0 113535.0 9345.0 113400.0 ;
      RECT  9280.0 113535.0 9345.0 113400.0 ;
      RECT  9445.0 113500.0 9510.0 113435.0 ;
      RECT  9155.0 112782.5 9715.0 112717.5 ;
      RECT  9155.0 114127.5 9715.0 114062.5 ;
      RECT  9782.5 113932.5 9847.5 114127.5 ;
      RECT  9782.5 113092.5 9847.5 112717.5 ;
      RECT  10162.5 113092.5 10227.5 112717.5 ;
      RECT  10332.5 112935.0 10397.5 112750.0 ;
      RECT  10332.5 114095.0 10397.5 113910.0 ;
      RECT  9782.5 113092.5 9847.5 112957.5 ;
      RECT  9972.5 113092.5 10037.5 112957.5 ;
      RECT  9972.5 113092.5 10037.5 112957.5 ;
      RECT  9782.5 113092.5 9847.5 112957.5 ;
      RECT  9972.5 113092.5 10037.5 112957.5 ;
      RECT  10162.5 113092.5 10227.5 112957.5 ;
      RECT  10162.5 113092.5 10227.5 112957.5 ;
      RECT  9972.5 113092.5 10037.5 112957.5 ;
      RECT  9782.5 113932.5 9847.5 113797.5 ;
      RECT  9972.5 113932.5 10037.5 113797.5 ;
      RECT  9972.5 113932.5 10037.5 113797.5 ;
      RECT  9782.5 113932.5 9847.5 113797.5 ;
      RECT  9972.5 113932.5 10037.5 113797.5 ;
      RECT  10162.5 113932.5 10227.5 113797.5 ;
      RECT  10162.5 113932.5 10227.5 113797.5 ;
      RECT  9972.5 113932.5 10037.5 113797.5 ;
      RECT  10332.5 113002.5 10397.5 112867.5 ;
      RECT  10332.5 113977.5 10397.5 113842.5 ;
      RECT  10167.5 113702.5 10032.5 113637.5 ;
      RECT  9910.0 113487.5 9775.0 113422.5 ;
      RECT  9972.5 113092.5 10037.5 112957.5 ;
      RECT  10162.5 113932.5 10227.5 113797.5 ;
      RECT  10262.5 113487.5 10127.5 113422.5 ;
      RECT  9775.0 113487.5 9910.0 113422.5 ;
      RECT  10032.5 113702.5 10167.5 113637.5 ;
      RECT  10127.5 113487.5 10262.5 113422.5 ;
      RECT  9715.0 112782.5 10635.0 112717.5 ;
      RECT  9715.0 114127.5 10635.0 114062.5 ;
      RECT  11062.5 112935.0 11127.5 112750.0 ;
      RECT  11062.5 114095.0 11127.5 113910.0 ;
      RECT  10702.5 113977.5 10767.5 114127.5 ;
      RECT  10702.5 113092.5 10767.5 112717.5 ;
      RECT  10892.5 113977.5 10957.5 113092.5 ;
      RECT  10702.5 113092.5 10767.5 112957.5 ;
      RECT  10892.5 113092.5 10957.5 112957.5 ;
      RECT  10892.5 113092.5 10957.5 112957.5 ;
      RECT  10702.5 113092.5 10767.5 112957.5 ;
      RECT  10702.5 113977.5 10767.5 113842.5 ;
      RECT  10892.5 113977.5 10957.5 113842.5 ;
      RECT  10892.5 113977.5 10957.5 113842.5 ;
      RECT  10702.5 113977.5 10767.5 113842.5 ;
      RECT  11062.5 113002.5 11127.5 112867.5 ;
      RECT  11062.5 113977.5 11127.5 113842.5 ;
      RECT  10760.0 113535.0 10825.0 113400.0 ;
      RECT  10760.0 113535.0 10825.0 113400.0 ;
      RECT  10925.0 113500.0 10990.0 113435.0 ;
      RECT  10635.0 112782.5 11195.0 112717.5 ;
      RECT  10635.0 114127.5 11195.0 114062.5 ;
      RECT  8897.5 113400.0 8962.5 113535.0 ;
      RECT  9037.5 113672.5 9102.5 113807.5 ;
      RECT  10032.5 113637.5 9897.5 113702.5 ;
      RECT  8700.0 28337.5 9070.0 28402.5 ;
      RECT  8700.0 30317.5 9070.0 30382.5 ;
      RECT  8700.0 31027.5 9070.0 31092.5 ;
      RECT  8700.0 33007.5 9070.0 33072.5 ;
      RECT  8700.0 33717.5 9070.0 33782.5 ;
      RECT  8700.0 35697.5 9070.0 35762.5 ;
      RECT  8700.0 36407.5 9070.0 36472.5 ;
      RECT  8700.0 38387.5 9070.0 38452.5 ;
      RECT  8700.0 39097.5 9070.0 39162.5 ;
      RECT  8700.0 41077.5 9070.0 41142.5 ;
      RECT  8700.0 41787.5 9070.0 41852.5 ;
      RECT  8700.0 43767.5 9070.0 43832.5 ;
      RECT  8700.0 44477.5 9070.0 44542.5 ;
      RECT  8700.0 46457.5 9070.0 46522.5 ;
      RECT  8700.0 47167.5 9070.0 47232.5 ;
      RECT  8700.0 49147.5 9070.0 49212.5 ;
      RECT  8700.0 49857.5 9070.0 49922.5 ;
      RECT  8700.0 51837.5 9070.0 51902.5 ;
      RECT  8700.0 52547.5 9070.0 52612.5 ;
      RECT  8700.0 54527.5 9070.0 54592.5 ;
      RECT  8700.0 55237.5 9070.0 55302.5 ;
      RECT  8700.0 57217.5 9070.0 57282.5 ;
      RECT  8700.0 57927.5 9070.0 57992.5 ;
      RECT  8700.0 59907.5 9070.0 59972.5 ;
      RECT  8700.0 60617.5 9070.0 60682.5 ;
      RECT  8700.0 62597.5 9070.0 62662.5 ;
      RECT  8700.0 63307.5 9070.0 63372.5 ;
      RECT  8700.0 65287.5 9070.0 65352.5 ;
      RECT  8700.0 65997.5 9070.0 66062.5 ;
      RECT  8700.0 67977.5 9070.0 68042.5 ;
      RECT  8700.0 68687.5 9070.0 68752.5 ;
      RECT  8700.0 70667.5 9070.0 70732.5 ;
      RECT  8700.0 71377.5 9070.0 71442.5 ;
      RECT  8700.0 73357.5 9070.0 73422.5 ;
      RECT  8700.0 74067.5 9070.0 74132.5 ;
      RECT  8700.0 76047.5 9070.0 76112.5 ;
      RECT  8700.0 76757.5 9070.0 76822.5 ;
      RECT  8700.0 78737.5 9070.0 78802.5 ;
      RECT  8700.0 79447.5 9070.0 79512.5 ;
      RECT  8700.0 81427.5 9070.0 81492.5 ;
      RECT  8700.0 82137.5 9070.0 82202.5 ;
      RECT  8700.0 84117.5 9070.0 84182.5 ;
      RECT  8700.0 84827.5 9070.0 84892.5 ;
      RECT  8700.0 86807.5 9070.0 86872.5 ;
      RECT  8700.0 87517.5 9070.0 87582.5 ;
      RECT  8700.0 89497.5 9070.0 89562.5 ;
      RECT  8700.0 90207.5 9070.0 90272.5 ;
      RECT  8700.0 92187.5 9070.0 92252.5 ;
      RECT  8700.0 92897.5 9070.0 92962.5 ;
      RECT  8700.0 94877.5 9070.0 94942.5 ;
      RECT  8700.0 95587.5 9070.0 95652.5 ;
      RECT  8700.0 97567.5 9070.0 97632.5 ;
      RECT  8700.0 98277.5 9070.0 98342.5 ;
      RECT  8700.0 100257.5 9070.0 100322.5 ;
      RECT  8700.0 100967.5 9070.0 101032.5 ;
      RECT  8700.0 102947.5 9070.0 103012.5 ;
      RECT  8700.0 103657.5 9070.0 103722.5 ;
      RECT  8700.0 105637.5 9070.0 105702.5 ;
      RECT  8700.0 106347.5 9070.0 106412.5 ;
      RECT  8700.0 108327.5 9070.0 108392.5 ;
      RECT  8700.0 109037.5 9070.0 109102.5 ;
      RECT  8700.0 111017.5 9070.0 111082.5 ;
      RECT  8700.0 111727.5 9070.0 111792.5 ;
      RECT  8700.0 113707.5 9070.0 113772.5 ;
      RECT  10925.0 28610.0 10990.0 28675.0 ;
      RECT  10925.0 30045.0 10990.0 30110.0 ;
      RECT  10925.0 31300.0 10990.0 31365.0 ;
      RECT  10925.0 32735.0 10990.0 32800.0 ;
      RECT  10925.0 33990.0 10990.0 34055.0 ;
      RECT  10925.0 35425.0 10990.0 35490.0 ;
      RECT  10925.0 36680.0 10990.0 36745.0 ;
      RECT  10925.0 38115.0 10990.0 38180.0 ;
      RECT  10925.0 39370.0 10990.0 39435.0 ;
      RECT  10925.0 40805.0 10990.0 40870.0 ;
      RECT  10925.0 42060.0 10990.0 42125.0 ;
      RECT  10925.0 43495.0 10990.0 43560.0 ;
      RECT  10925.0 44750.0 10990.0 44815.0 ;
      RECT  10925.0 46185.0 10990.0 46250.0 ;
      RECT  10925.0 47440.0 10990.0 47505.0 ;
      RECT  10925.0 48875.0 10990.0 48940.0 ;
      RECT  10925.0 50130.0 10990.0 50195.0 ;
      RECT  10925.0 51565.0 10990.0 51630.0 ;
      RECT  10925.0 52820.0 10990.0 52885.0 ;
      RECT  10925.0 54255.0 10990.0 54320.0 ;
      RECT  10925.0 55510.0 10990.0 55575.0 ;
      RECT  10925.0 56945.0 10990.0 57010.0 ;
      RECT  10925.0 58200.0 10990.0 58265.0 ;
      RECT  10925.0 59635.0 10990.0 59700.0 ;
      RECT  10925.0 60890.0 10990.0 60955.0 ;
      RECT  10925.0 62325.0 10990.0 62390.0 ;
      RECT  10925.0 63580.0 10990.0 63645.0 ;
      RECT  10925.0 65015.0 10990.0 65080.0 ;
      RECT  10925.0 66270.0 10990.0 66335.0 ;
      RECT  10925.0 67705.0 10990.0 67770.0 ;
      RECT  10925.0 68960.0 10990.0 69025.0 ;
      RECT  10925.0 70395.0 10990.0 70460.0 ;
      RECT  10925.0 71650.0 10990.0 71715.0 ;
      RECT  10925.0 73085.0 10990.0 73150.0 ;
      RECT  10925.0 74340.0 10990.0 74405.0 ;
      RECT  10925.0 75775.0 10990.0 75840.0 ;
      RECT  10925.0 77030.0 10990.0 77095.0 ;
      RECT  10925.0 78465.0 10990.0 78530.0 ;
      RECT  10925.0 79720.0 10990.0 79785.0 ;
      RECT  10925.0 81155.0 10990.0 81220.0 ;
      RECT  10925.0 82410.0 10990.0 82475.0 ;
      RECT  10925.0 83845.0 10990.0 83910.0 ;
      RECT  10925.0 85100.0 10990.0 85165.0 ;
      RECT  10925.0 86535.0 10990.0 86600.0 ;
      RECT  10925.0 87790.0 10990.0 87855.0 ;
      RECT  10925.0 89225.0 10990.0 89290.0 ;
      RECT  10925.0 90480.0 10990.0 90545.0 ;
      RECT  10925.0 91915.0 10990.0 91980.0 ;
      RECT  10925.0 93170.0 10990.0 93235.0 ;
      RECT  10925.0 94605.0 10990.0 94670.0 ;
      RECT  10925.0 95860.0 10990.0 95925.0 ;
      RECT  10925.0 97295.0 10990.0 97360.0 ;
      RECT  10925.0 98550.0 10990.0 98615.0 ;
      RECT  10925.0 99985.0 10990.0 100050.0 ;
      RECT  10925.0 101240.0 10990.0 101305.0 ;
      RECT  10925.0 102675.0 10990.0 102740.0 ;
      RECT  10925.0 103930.0 10990.0 103995.0 ;
      RECT  10925.0 105365.0 10990.0 105430.0 ;
      RECT  10925.0 106620.0 10990.0 106685.0 ;
      RECT  10925.0 108055.0 10990.0 108120.0 ;
      RECT  10925.0 109310.0 10990.0 109375.0 ;
      RECT  10925.0 110745.0 10990.0 110810.0 ;
      RECT  10925.0 112000.0 10990.0 112065.0 ;
      RECT  10925.0 113435.0 10990.0 113500.0 ;
      RECT  8700.0 29327.5 9155.0 29392.5 ;
      RECT  8700.0 32017.5 9155.0 32082.5 ;
      RECT  8700.0 34707.5 9155.0 34772.5 ;
      RECT  8700.0 37397.5 9155.0 37462.5 ;
      RECT  8700.0 40087.5 9155.0 40152.5 ;
      RECT  8700.0 42777.5 9155.0 42842.5 ;
      RECT  8700.0 45467.5 9155.0 45532.5 ;
      RECT  8700.0 48157.5 9155.0 48222.5 ;
      RECT  8700.0 50847.5 9155.0 50912.5 ;
      RECT  8700.0 53537.5 9155.0 53602.5 ;
      RECT  8700.0 56227.5 9155.0 56292.5 ;
      RECT  8700.0 58917.5 9155.0 58982.5 ;
      RECT  8700.0 61607.5 9155.0 61672.5 ;
      RECT  8700.0 64297.5 9155.0 64362.5 ;
      RECT  8700.0 66987.5 9155.0 67052.5 ;
      RECT  8700.0 69677.5 9155.0 69742.5 ;
      RECT  8700.0 72367.5 9155.0 72432.5 ;
      RECT  8700.0 75057.5 9155.0 75122.5 ;
      RECT  8700.0 77747.5 9155.0 77812.5 ;
      RECT  8700.0 80437.5 9155.0 80502.5 ;
      RECT  8700.0 83127.5 9155.0 83192.5 ;
      RECT  8700.0 85817.5 9155.0 85882.5 ;
      RECT  8700.0 88507.5 9155.0 88572.5 ;
      RECT  8700.0 91197.5 9155.0 91262.5 ;
      RECT  8700.0 93887.5 9155.0 93952.5 ;
      RECT  8700.0 96577.5 9155.0 96642.5 ;
      RECT  8700.0 99267.5 9155.0 99332.5 ;
      RECT  8700.0 101957.5 9155.0 102022.5 ;
      RECT  8700.0 104647.5 9155.0 104712.5 ;
      RECT  8700.0 107337.5 9155.0 107402.5 ;
      RECT  8700.0 110027.5 9155.0 110092.5 ;
      RECT  8700.0 112717.5 9155.0 112782.5 ;
      RECT  8700.0 27982.5 9155.0 28047.5 ;
      RECT  8700.0 30672.5 9155.0 30737.5 ;
      RECT  8700.0 33362.5 9155.0 33427.5 ;
      RECT  8700.0 36052.5 9155.0 36117.5 ;
      RECT  8700.0 38742.5 9155.0 38807.5 ;
      RECT  8700.0 41432.5 9155.0 41497.5 ;
      RECT  8700.0 44122.5 9155.0 44187.5 ;
      RECT  8700.0 46812.5 9155.0 46877.5 ;
      RECT  8700.0 49502.5 9155.0 49567.5 ;
      RECT  8700.0 52192.5 9155.0 52257.5 ;
      RECT  8700.0 54882.5 9155.0 54947.5 ;
      RECT  8700.0 57572.5 9155.0 57637.5 ;
      RECT  8700.0 60262.5 9155.0 60327.5 ;
      RECT  8700.0 62952.5 9155.0 63017.5 ;
      RECT  8700.0 65642.5 9155.0 65707.5 ;
      RECT  8700.0 68332.5 9155.0 68397.5 ;
      RECT  8700.0 71022.5 9155.0 71087.5 ;
      RECT  8700.0 73712.5 9155.0 73777.5 ;
      RECT  8700.0 76402.5 9155.0 76467.5 ;
      RECT  8700.0 79092.5 9155.0 79157.5 ;
      RECT  8700.0 81782.5 9155.0 81847.5 ;
      RECT  8700.0 84472.5 9155.0 84537.5 ;
      RECT  8700.0 87162.5 9155.0 87227.5 ;
      RECT  8700.0 89852.5 9155.0 89917.5 ;
      RECT  8700.0 92542.5 9155.0 92607.5 ;
      RECT  8700.0 95232.5 9155.0 95297.5 ;
      RECT  8700.0 97922.5 9155.0 97987.5 ;
      RECT  8700.0 100612.5 9155.0 100677.5 ;
      RECT  8700.0 103302.5 9155.0 103367.5 ;
      RECT  8700.0 105992.5 9155.0 106057.5 ;
      RECT  8700.0 108682.5 9155.0 108747.5 ;
      RECT  8700.0 111372.5 9155.0 111437.5 ;
      RECT  8700.0 114062.5 9155.0 114127.5 ;
      RECT  4655.0 11465.0 11095.0 10760.0 ;
      RECT  4655.0 10055.0 11095.0 10760.0 ;
      RECT  4655.0 10055.0 11095.0 9350.0 ;
      RECT  4655.0 8645.0 11095.0 9350.0 ;
      RECT  4655.0 8645.0 11095.0 7940.0 ;
      RECT  4655.0 7235.0 11095.0 7940.0 ;
      RECT  4655.0 7235.0 11095.0 6530.0 ;
      RECT  4655.0 5825.0 11095.0 6530.0 ;
      RECT  4860.0 11465.0 4925.0 5825.0 ;
      RECT  7865.0 11465.0 7930.0 5825.0 ;
      RECT  10825.0 11465.0 10890.0 5825.0 ;
      RECT  5875.0 11465.0 5940.0 5825.0 ;
      RECT  8835.0 11465.0 8900.0 5825.0 ;
      RECT  5020.0 11465.0 5085.0 5825.0 ;
      RECT  13657.5 28047.5 13792.5 27982.5 ;
      RECT  13657.5 30737.5 13792.5 30672.5 ;
      RECT  13657.5 33427.5 13792.5 33362.5 ;
      RECT  13657.5 36117.5 13792.5 36052.5 ;
      RECT  13657.5 38807.5 13792.5 38742.5 ;
      RECT  13657.5 41497.5 13792.5 41432.5 ;
      RECT  13657.5 44187.5 13792.5 44122.5 ;
      RECT  13657.5 46877.5 13792.5 46812.5 ;
      RECT  13657.5 49567.5 13792.5 49502.5 ;
      RECT  13657.5 52257.5 13792.5 52192.5 ;
      RECT  13657.5 54947.5 13792.5 54882.5 ;
      RECT  13657.5 57637.5 13792.5 57572.5 ;
      RECT  13657.5 60327.5 13792.5 60262.5 ;
      RECT  13657.5 63017.5 13792.5 62952.5 ;
      RECT  13657.5 65707.5 13792.5 65642.5 ;
      RECT  13657.5 68397.5 13792.5 68332.5 ;
      RECT  13657.5 71087.5 13792.5 71022.5 ;
      RECT  13657.5 73777.5 13792.5 73712.5 ;
      RECT  13657.5 76467.5 13792.5 76402.5 ;
      RECT  13657.5 79157.5 13792.5 79092.5 ;
      RECT  13657.5 81847.5 13792.5 81782.5 ;
      RECT  13657.5 84537.5 13792.5 84472.5 ;
      RECT  13657.5 87227.5 13792.5 87162.5 ;
      RECT  13657.5 89917.5 13792.5 89852.5 ;
      RECT  13657.5 92607.5 13792.5 92542.5 ;
      RECT  13657.5 95297.5 13792.5 95232.5 ;
      RECT  13657.5 97987.5 13792.5 97922.5 ;
      RECT  13657.5 100677.5 13792.5 100612.5 ;
      RECT  13657.5 103367.5 13792.5 103302.5 ;
      RECT  13657.5 106057.5 13792.5 105992.5 ;
      RECT  13657.5 108747.5 13792.5 108682.5 ;
      RECT  13657.5 111437.5 13792.5 111372.5 ;
      RECT  13657.5 114127.5 13792.5 114062.5 ;
      RECT  11095.0 12047.5 10960.0 12112.5 ;
      RECT  11505.0 12047.5 11370.0 12112.5 ;
      RECT  10820.0 13392.5 10685.0 13457.5 ;
      RECT  11710.0 13392.5 11575.0 13457.5 ;
      RECT  11095.0 17427.5 10960.0 17492.5 ;
      RECT  11915.0 17427.5 11780.0 17492.5 ;
      RECT  10820.0 18772.5 10685.0 18837.5 ;
      RECT  12120.0 18772.5 11985.0 18837.5 ;
      RECT  11095.0 22807.5 10960.0 22872.5 ;
      RECT  12325.0 22807.5 12190.0 22872.5 ;
      RECT  10820.0 24152.5 10685.0 24217.5 ;
      RECT  12530.0 24152.5 12395.0 24217.5 ;
      RECT  11300.0 11842.5 11165.0 11907.5 ;
      RECT  11300.0 14532.5 11165.0 14597.5 ;
      RECT  11300.0 17222.5 11165.0 17287.5 ;
      RECT  11300.0 19912.5 11165.0 19977.5 ;
      RECT  11300.0 22602.5 11165.0 22667.5 ;
      RECT  11300.0 25292.5 11165.0 25357.5 ;
      RECT  12735.0 26012.5 12600.0 26077.5 ;
      RECT  12940.0 25872.5 12805.0 25937.5 ;
      RECT  13145.0 25732.5 13010.0 25797.5 ;
      RECT  13350.0 25592.5 13215.0 25657.5 ;
      RECT  12735.0 630.0 12600.0 695.0 ;
      RECT  12940.0 2065.0 12805.0 2130.0 ;
      RECT  13145.0 3320.0 13010.0 3385.0 ;
      RECT  13350.0 4755.0 13215.0 4820.0 ;
      RECT  13657.5 67.5 13792.5 2.5 ;
      RECT  13657.5 2757.5 13792.5 2692.5 ;
      RECT  13657.5 5447.5 13792.5 5382.5 ;
      RECT  11162.5 11080.0 11027.5 11145.0 ;
      RECT  11505.0 11080.0 11370.0 11145.0 ;
      RECT  11162.5 10375.0 11027.5 10440.0 ;
      RECT  11710.0 10375.0 11575.0 10440.0 ;
      RECT  11162.5 9670.0 11027.5 9735.0 ;
      RECT  11915.0 9670.0 11780.0 9735.0 ;
      RECT  11162.5 8965.0 11027.5 9030.0 ;
      RECT  12120.0 8965.0 11985.0 9030.0 ;
      RECT  11162.5 8260.0 11027.5 8325.0 ;
      RECT  12325.0 8260.0 12190.0 8325.0 ;
      RECT  11162.5 7555.0 11027.5 7620.0 ;
      RECT  12530.0 7555.0 12395.0 7620.0 ;
      RECT  11230.0 11432.5 11095.0 11497.5 ;
      RECT  13792.5 11432.5 13657.5 11497.5 ;
      RECT  11230.0 10727.5 11095.0 10792.5 ;
      RECT  13792.5 10727.5 13657.5 10792.5 ;
      RECT  11230.0 10022.5 11095.0 10087.5 ;
      RECT  13792.5 10022.5 13657.5 10087.5 ;
      RECT  11230.0 9317.5 11095.0 9382.5 ;
      RECT  13792.5 9317.5 13657.5 9382.5 ;
      RECT  11230.0 8612.5 11095.0 8677.5 ;
      RECT  13792.5 8612.5 13657.5 8677.5 ;
      RECT  11230.0 7907.5 11095.0 7972.5 ;
      RECT  13792.5 7907.5 13657.5 7972.5 ;
      RECT  11230.0 7202.5 11095.0 7267.5 ;
      RECT  13792.5 7202.5 13657.5 7267.5 ;
      RECT  11230.0 6497.5 11095.0 6562.5 ;
      RECT  13792.5 6497.5 13657.5 6562.5 ;
      RECT  11230.0 5792.5 11095.0 5857.5 ;
      RECT  13792.5 5792.5 13657.5 5857.5 ;
      RECT  14930.0 9875.0 14795.0 9940.0 ;
      RECT  14520.0 7690.0 14385.0 7755.0 ;
      RECT  14725.0 9237.5 14590.0 9302.5 ;
      RECT  14930.0 115072.5 14795.0 115137.5 ;
      RECT  15135.0 16377.5 15000.0 16442.5 ;
      RECT  15340.0 20402.5 15205.0 20467.5 ;
      RECT  14315.0 11637.5 14180.0 11702.5 ;
      RECT  8997.5 114267.5 8862.5 114332.5 ;
      RECT  14315.0 114267.5 14180.0 114332.5 ;
      RECT  14007.5 9107.5 13872.5 9172.5 ;
      RECT  14007.5 20532.5 13872.5 20597.5 ;
      RECT  14007.5 10035.0 13872.5 10100.0 ;
      RECT  14007.5 17310.0 13872.5 17375.0 ;
      RECT  106185.0 35.0 106535.0 115822.5 ;
      RECT  4175.0 35.0 4525.0 115822.5 ;
      RECT  3455.0 28445.0 3390.0 28510.0 ;
      RECT  3422.5 28445.0 3407.5 28510.0 ;
      RECT  3455.0 28477.5 3390.0 29062.5 ;
      RECT  3455.0 29607.5 3390.0 30002.5 ;
      RECT  3455.0 30927.5 3390.0 31512.5 ;
      RECT  2657.5 31365.0 2280.0 31430.0 ;
      RECT  2657.5 34325.0 2280.0 34390.0 ;
      RECT  2657.5 29375.0 2280.0 29440.0 ;
      RECT  2657.5 32335.0 2280.0 32400.0 ;
      RECT  3440.0 28445.0 3375.0 28510.0 ;
      RECT  3455.0 29575.0 3390.0 29640.0 ;
      RECT  2005.0 40260.0 1940.0 41025.0 ;
      RECT  3455.0 33610.0 3390.0 35040.0 ;
      RECT  2485.0 28360.0 2280.0 28425.0 ;
      RECT  1962.5 35040.0 1897.5 36977.5 ;
      RECT  1747.5 35450.0 1682.5 37235.0 ;
      RECT  3380.0 36475.0 3315.0 37045.0 ;
      RECT  3520.0 36270.0 3455.0 37235.0 ;
      RECT  3660.0 35655.0 3595.0 37425.0 ;
      RECT  3380.0 37985.0 3315.0 38050.0 ;
      RECT  3380.0 37520.0 3315.0 38017.5 ;
      RECT  3407.5 37985.0 3347.5 38050.0 ;
      RECT  3475.0 38150.0 3410.0 38215.0 ;
      RECT  3442.5 38150.0 3407.5 38215.0 ;
      RECT  3475.0 38182.5 3410.0 41722.5 ;
      RECT  690.0 36475.0 625.0 37605.0 ;
      RECT  830.0 35655.0 765.0 37795.0 ;
      RECT  970.0 35860.0 905.0 37985.0 ;
      RECT  690.0 38545.0 625.0 38610.0 ;
      RECT  690.0 38080.0 625.0 38577.5 ;
      RECT  717.5 38545.0 657.5 38610.0 ;
      RECT  750.0 38742.5 685.0 39137.5 ;
      RECT  750.0 39302.5 685.0 39697.5 ;
      RECT  2005.0 40227.5 1940.0 40292.5 ;
      RECT  1972.5 40227.5 1940.0 40292.5 ;
      RECT  2005.0 40135.0 1940.0 40260.0 ;
      RECT  2005.0 39542.5 1940.0 39937.5 ;
      RECT  1962.5 37400.0 1897.5 37770.0 ;
      RECT  2017.5 38475.0 1952.5 38915.0 ;
      RECT  750.0 39862.5 685.0 40100.0 ;
      RECT  2005.0 39140.0 1940.0 39377.5 ;
      RECT  4067.5 28155.0 4002.5 40260.0 ;
      RECT  4067.5 35245.0 4002.5 36850.0 ;
      RECT  2722.5 28155.0 2657.5 40260.0 ;
      RECT  2722.5 36065.0 2657.5 36850.0 ;
      RECT  1377.5 36850.0 1312.5 40260.0 ;
      RECT  1377.5 35245.0 1312.5 36850.0 ;
      RECT  32.5 36850.0 -32.5 40260.0 ;
      RECT  32.5 36065.0 -32.5 36850.0 ;
      RECT  32.5 40227.5 -32.5 40292.5 ;
      RECT  32.5 40055.0 -32.5 40260.0 ;
      RECT  8.881784197e-13 40227.5 -45.0 40292.5 ;
      RECT  165.0 28155.0 870.0 34595.0 ;
      RECT  1575.0 28155.0 870.0 34595.0 ;
      RECT  1575.0 28155.0 2280.0 34595.0 ;
      RECT  165.0 28360.0 2280.0 28425.0 ;
      RECT  165.0 31365.0 2280.0 31430.0 ;
      RECT  165.0 34325.0 2280.0 34390.0 ;
      RECT  165.0 29375.0 2280.0 29440.0 ;
      RECT  165.0 32335.0 2280.0 32400.0 ;
      RECT  165.0 28520.0 2280.0 28585.0 ;
      RECT  2875.0 28772.5 2690.0 28837.5 ;
      RECT  4035.0 28772.5 3850.0 28837.5 ;
      RECT  2832.5 28222.5 2657.5 28667.5 ;
      RECT  3917.5 28412.5 3032.5 28477.5 ;
      RECT  2965.0 28222.5 2800.0 28287.5 ;
      RECT  2965.0 28602.5 2800.0 28667.5 ;
      RECT  3032.5 28222.5 2897.5 28287.5 ;
      RECT  3032.5 28602.5 2897.5 28667.5 ;
      RECT  3032.5 28412.5 2897.5 28477.5 ;
      RECT  3032.5 28412.5 2897.5 28477.5 ;
      RECT  2832.5 28222.5 2767.5 28667.5 ;
      RECT  4015.0 28222.5 3850.0 28287.5 ;
      RECT  4015.0 28602.5 3850.0 28667.5 ;
      RECT  3917.5 28222.5 3782.5 28287.5 ;
      RECT  3917.5 28602.5 3782.5 28667.5 ;
      RECT  3917.5 28412.5 3782.5 28477.5 ;
      RECT  3917.5 28412.5 3782.5 28477.5 ;
      RECT  4047.5 28222.5 3982.5 28667.5 ;
      RECT  2942.5 28772.5 2807.5 28837.5 ;
      RECT  3917.5 28772.5 3782.5 28837.5 ;
      RECT  3475.0 28280.0 3340.0 28345.0 ;
      RECT  3475.0 28280.0 3340.0 28345.0 ;
      RECT  3440.0 28445.0 3375.0 28510.0 ;
      RECT  2722.5 28155.0 2657.5 28905.0 ;
      RECT  4067.5 28155.0 4002.5 28905.0 ;
      RECT  2875.0 29712.5 2690.0 29777.5 ;
      RECT  4035.0 29712.5 3850.0 29777.5 ;
      RECT  2877.5 28972.5 2657.5 29417.5 ;
      RECT  3702.5 29542.5 3207.5 29607.5 ;
      RECT  3010.0 28972.5 2845.0 29037.5 ;
      RECT  3010.0 29352.5 2845.0 29417.5 ;
      RECT  3175.0 29162.5 3010.0 29227.5 ;
      RECT  3175.0 29542.5 3010.0 29607.5 ;
      RECT  3077.5 28972.5 2942.5 29037.5 ;
      RECT  3077.5 29352.5 2942.5 29417.5 ;
      RECT  3077.5 29162.5 2942.5 29227.5 ;
      RECT  3077.5 29542.5 2942.5 29607.5 ;
      RECT  3207.5 29162.5 3142.5 29607.5 ;
      RECT  2877.5 28972.5 2812.5 29417.5 ;
      RECT  4000.0 28972.5 3835.0 29037.5 ;
      RECT  4000.0 29352.5 3835.0 29417.5 ;
      RECT  3835.0 29162.5 3670.0 29227.5 ;
      RECT  3835.0 29542.5 3670.0 29607.5 ;
      RECT  3902.5 28972.5 3767.5 29037.5 ;
      RECT  3902.5 29352.5 3767.5 29417.5 ;
      RECT  3902.5 29162.5 3767.5 29227.5 ;
      RECT  3902.5 29542.5 3767.5 29607.5 ;
      RECT  3702.5 29162.5 3637.5 29607.5 ;
      RECT  4032.5 28972.5 3967.5 29417.5 ;
      RECT  2942.5 29712.5 2807.5 29777.5 ;
      RECT  3917.5 29712.5 3782.5 29777.5 ;
      RECT  3490.0 29030.0 3355.0 29095.0 ;
      RECT  3490.0 29030.0 3355.0 29095.0 ;
      RECT  3455.0 29575.0 3390.0 29640.0 ;
      RECT  2722.5 28905.0 2657.5 29845.0 ;
      RECT  4067.5 28905.0 4002.5 29845.0 ;
      RECT  2875.0 31222.5 2690.0 31287.5 ;
      RECT  4035.0 31222.5 3850.0 31287.5 ;
      RECT  2877.5 29912.5 2657.5 31117.5 ;
      RECT  3702.5 30862.5 3207.5 30927.5 ;
      RECT  3010.0 29912.5 2845.0 29977.5 ;
      RECT  3010.0 30292.5 2845.0 30357.5 ;
      RECT  3010.0 30672.5 2845.0 30737.5 ;
      RECT  3010.0 31052.5 2845.0 31117.5 ;
      RECT  3175.0 30102.5 3010.0 30167.5 ;
      RECT  3175.0 30482.5 3010.0 30547.5 ;
      RECT  3175.0 30862.5 3010.0 30927.5 ;
      RECT  3077.5 29912.5 2942.5 29977.5 ;
      RECT  3077.5 30292.5 2942.5 30357.5 ;
      RECT  3077.5 30672.5 2942.5 30737.5 ;
      RECT  3077.5 31052.5 2942.5 31117.5 ;
      RECT  3077.5 30102.5 2942.5 30167.5 ;
      RECT  3077.5 30482.5 2942.5 30547.5 ;
      RECT  3077.5 30862.5 2942.5 30927.5 ;
      RECT  3207.5 30102.5 3142.5 30927.5 ;
      RECT  2877.5 29912.5 2812.5 31117.5 ;
      RECT  4000.0 29912.5 3835.0 29977.5 ;
      RECT  4000.0 30292.5 3835.0 30357.5 ;
      RECT  4000.0 30672.5 3835.0 30737.5 ;
      RECT  4000.0 31052.5 3835.0 31117.5 ;
      RECT  3835.0 30102.5 3670.0 30167.5 ;
      RECT  3835.0 30482.5 3670.0 30547.5 ;
      RECT  3835.0 30862.5 3670.0 30927.5 ;
      RECT  3902.5 29912.5 3767.5 29977.5 ;
      RECT  3902.5 30292.5 3767.5 30357.5 ;
      RECT  3902.5 30672.5 3767.5 30737.5 ;
      RECT  3902.5 31052.5 3767.5 31117.5 ;
      RECT  3902.5 30102.5 3767.5 30167.5 ;
      RECT  3902.5 30482.5 3767.5 30547.5 ;
      RECT  3902.5 30862.5 3767.5 30927.5 ;
      RECT  3702.5 30102.5 3637.5 30927.5 ;
      RECT  4032.5 29912.5 3967.5 31117.5 ;
      RECT  2942.5 31222.5 2807.5 31287.5 ;
      RECT  3917.5 31222.5 3782.5 31287.5 ;
      RECT  3490.0 29970.0 3355.0 30035.0 ;
      RECT  3490.0 29970.0 3355.0 30035.0 ;
      RECT  3455.0 30895.0 3390.0 30960.0 ;
      RECT  2722.5 29845.0 2657.5 31355.0 ;
      RECT  4067.5 29845.0 4002.5 31355.0 ;
      RECT  2875.0 33872.5 2690.0 33937.5 ;
      RECT  4035.0 33872.5 3850.0 33937.5 ;
      RECT  2877.5 31422.5 2657.5 33767.5 ;
      RECT  3702.5 33512.5 3207.5 33577.5 ;
      RECT  3010.0 31422.5 2845.0 31487.5 ;
      RECT  3010.0 31802.5 2845.0 31867.5 ;
      RECT  3010.0 32182.5 2845.0 32247.5 ;
      RECT  3010.0 32562.5 2845.0 32627.5 ;
      RECT  3010.0 32942.5 2845.0 33007.5 ;
      RECT  3010.0 33322.5 2845.0 33387.5 ;
      RECT  3010.0 33702.5 2845.0 33767.5 ;
      RECT  3175.0 31612.5 3010.0 31677.5 ;
      RECT  3175.0 31992.5 3010.0 32057.5 ;
      RECT  3175.0 32372.5 3010.0 32437.5 ;
      RECT  3175.0 32752.5 3010.0 32817.5 ;
      RECT  3175.0 33132.5 3010.0 33197.5 ;
      RECT  3175.0 33512.5 3010.0 33577.5 ;
      RECT  3077.5 31422.5 2942.5 31487.5 ;
      RECT  3077.5 31802.5 2942.5 31867.5 ;
      RECT  3077.5 32182.5 2942.5 32247.5 ;
      RECT  3077.5 32562.5 2942.5 32627.5 ;
      RECT  3077.5 32942.5 2942.5 33007.5 ;
      RECT  3077.5 33322.5 2942.5 33387.5 ;
      RECT  3077.5 33702.5 2942.5 33767.5 ;
      RECT  3077.5 31612.5 2942.5 31677.5 ;
      RECT  3077.5 31992.5 2942.5 32057.5 ;
      RECT  3077.5 32372.5 2942.5 32437.5 ;
      RECT  3077.5 32752.5 2942.5 32817.5 ;
      RECT  3077.5 33132.5 2942.5 33197.5 ;
      RECT  3077.5 33512.5 2942.5 33577.5 ;
      RECT  3207.5 31612.5 3142.5 33577.5 ;
      RECT  2877.5 31422.5 2812.5 33767.5 ;
      RECT  4000.0 31422.5 3835.0 31487.5 ;
      RECT  4000.0 31802.5 3835.0 31867.5 ;
      RECT  4000.0 32182.5 3835.0 32247.5 ;
      RECT  4000.0 32562.5 3835.0 32627.5 ;
      RECT  4000.0 32942.5 3835.0 33007.5 ;
      RECT  4000.0 33322.5 3835.0 33387.5 ;
      RECT  4000.0 33702.5 3835.0 33767.5 ;
      RECT  3835.0 31612.5 3670.0 31677.5 ;
      RECT  3835.0 31992.5 3670.0 32057.5 ;
      RECT  3835.0 32372.5 3670.0 32437.5 ;
      RECT  3835.0 32752.5 3670.0 32817.5 ;
      RECT  3835.0 33132.5 3670.0 33197.5 ;
      RECT  3835.0 33512.5 3670.0 33577.5 ;
      RECT  3902.5 31422.5 3767.5 31487.5 ;
      RECT  3902.5 31802.5 3767.5 31867.5 ;
      RECT  3902.5 32182.5 3767.5 32247.5 ;
      RECT  3902.5 32562.5 3767.5 32627.5 ;
      RECT  3902.5 32942.5 3767.5 33007.5 ;
      RECT  3902.5 33322.5 3767.5 33387.5 ;
      RECT  3902.5 33702.5 3767.5 33767.5 ;
      RECT  3902.5 31612.5 3767.5 31677.5 ;
      RECT  3902.5 31992.5 3767.5 32057.5 ;
      RECT  3902.5 32372.5 3767.5 32437.5 ;
      RECT  3902.5 32752.5 3767.5 32817.5 ;
      RECT  3902.5 33132.5 3767.5 33197.5 ;
      RECT  3902.5 33512.5 3767.5 33577.5 ;
      RECT  3702.5 31612.5 3637.5 33577.5 ;
      RECT  4032.5 31422.5 3967.5 33767.5 ;
      RECT  2942.5 33872.5 2807.5 33937.5 ;
      RECT  3917.5 33872.5 3782.5 33937.5 ;
      RECT  3490.0 31480.0 3355.0 31545.0 ;
      RECT  3490.0 31480.0 3355.0 31545.0 ;
      RECT  3455.0 33545.0 3390.0 33610.0 ;
      RECT  2722.5 31355.0 2657.5 34005.0 ;
      RECT  4067.5 31355.0 4002.5 34005.0 ;
      RECT  3872.5 36917.5 4067.5 36982.5 ;
      RECT  3032.5 36917.5 2657.5 36982.5 ;
      RECT  3032.5 37297.5 2657.5 37362.5 ;
      RECT  2875.0 37657.5 2690.0 37722.5 ;
      RECT  4035.0 37657.5 3850.0 37722.5 ;
      RECT  3032.5 36917.5 2897.5 36982.5 ;
      RECT  3032.5 37107.5 2897.5 37172.5 ;
      RECT  3032.5 37107.5 2897.5 37172.5 ;
      RECT  3032.5 36917.5 2897.5 36982.5 ;
      RECT  3032.5 37107.5 2897.5 37172.5 ;
      RECT  3032.5 37297.5 2897.5 37362.5 ;
      RECT  3032.5 37297.5 2897.5 37362.5 ;
      RECT  3032.5 37107.5 2897.5 37172.5 ;
      RECT  3032.5 37297.5 2897.5 37362.5 ;
      RECT  3032.5 37487.5 2897.5 37552.5 ;
      RECT  3032.5 37487.5 2897.5 37552.5 ;
      RECT  3032.5 37297.5 2897.5 37362.5 ;
      RECT  3872.5 36917.5 3737.5 36982.5 ;
      RECT  3872.5 37107.5 3737.5 37172.5 ;
      RECT  3872.5 37107.5 3737.5 37172.5 ;
      RECT  3872.5 36917.5 3737.5 36982.5 ;
      RECT  3872.5 37107.5 3737.5 37172.5 ;
      RECT  3872.5 37297.5 3737.5 37362.5 ;
      RECT  3872.5 37297.5 3737.5 37362.5 ;
      RECT  3872.5 37107.5 3737.5 37172.5 ;
      RECT  3872.5 37297.5 3737.5 37362.5 ;
      RECT  3872.5 37487.5 3737.5 37552.5 ;
      RECT  3872.5 37487.5 3737.5 37552.5 ;
      RECT  3872.5 37297.5 3737.5 37362.5 ;
      RECT  2942.5 37657.5 2807.5 37722.5 ;
      RECT  3917.5 37657.5 3782.5 37722.5 ;
      RECT  3660.0 37492.5 3595.0 37357.5 ;
      RECT  3520.0 37302.5 3455.0 37167.5 ;
      RECT  3380.0 37112.5 3315.0 36977.5 ;
      RECT  3032.5 37107.5 2897.5 37172.5 ;
      RECT  3032.5 37487.5 2897.5 37552.5 ;
      RECT  3872.5 37487.5 3737.5 37552.5 ;
      RECT  3415.0 37487.5 3280.0 37552.5 ;
      RECT  3380.0 36977.5 3315.0 37112.5 ;
      RECT  3520.0 37167.5 3455.0 37302.5 ;
      RECT  3660.0 37357.5 3595.0 37492.5 ;
      RECT  3415.0 37487.5 3280.0 37552.5 ;
      RECT  2722.5 36850.0 2657.5 37860.0 ;
      RECT  4067.5 36850.0 4002.5 37860.0 ;
      RECT  2875.0 38287.5 2690.0 38352.5 ;
      RECT  4035.0 38287.5 3850.0 38352.5 ;
      RECT  3917.5 37927.5 4067.5 37992.5 ;
      RECT  3032.5 37927.5 2657.5 37992.5 ;
      RECT  3917.5 38117.5 3032.5 38182.5 ;
      RECT  3032.5 37927.5 2897.5 37992.5 ;
      RECT  3032.5 38117.5 2897.5 38182.5 ;
      RECT  3032.5 38117.5 2897.5 38182.5 ;
      RECT  3032.5 37927.5 2897.5 37992.5 ;
      RECT  3917.5 37927.5 3782.5 37992.5 ;
      RECT  3917.5 38117.5 3782.5 38182.5 ;
      RECT  3917.5 38117.5 3782.5 38182.5 ;
      RECT  3917.5 37927.5 3782.5 37992.5 ;
      RECT  2942.5 38287.5 2807.5 38352.5 ;
      RECT  3917.5 38287.5 3782.5 38352.5 ;
      RECT  3475.0 37985.0 3340.0 38050.0 ;
      RECT  3475.0 37985.0 3340.0 38050.0 ;
      RECT  3440.0 38150.0 3375.0 38215.0 ;
      RECT  2722.5 37860.0 2657.5 38420.0 ;
      RECT  4067.5 37860.0 4002.5 38420.0 ;
      RECT  1462.5 36917.5 1312.5 36982.5 ;
      RECT  1462.5 37297.5 1312.5 37362.5 ;
      RECT  2280.0 36917.5 2722.5 36982.5 ;
      RECT  2505.0 37467.5 2690.0 37532.5 ;
      RECT  1345.0 37467.5 1530.0 37532.5 ;
      RECT  2280.0 36917.5 2415.0 36982.5 ;
      RECT  2280.0 37107.5 2415.0 37172.5 ;
      RECT  2280.0 37107.5 2415.0 37172.5 ;
      RECT  2280.0 36917.5 2415.0 36982.5 ;
      RECT  2280.0 37107.5 2415.0 37172.5 ;
      RECT  2280.0 37297.5 2415.0 37362.5 ;
      RECT  2280.0 37297.5 2415.0 37362.5 ;
      RECT  2280.0 37107.5 2415.0 37172.5 ;
      RECT  1462.5 36917.5 1597.5 36982.5 ;
      RECT  1462.5 37107.5 1597.5 37172.5 ;
      RECT  1462.5 37107.5 1597.5 37172.5 ;
      RECT  1462.5 36917.5 1597.5 36982.5 ;
      RECT  1462.5 37107.5 1597.5 37172.5 ;
      RECT  1462.5 37297.5 1597.5 37362.5 ;
      RECT  1462.5 37297.5 1597.5 37362.5 ;
      RECT  1462.5 37107.5 1597.5 37172.5 ;
      RECT  2437.5 37467.5 2572.5 37532.5 ;
      RECT  1462.5 37467.5 1597.5 37532.5 ;
      RECT  1682.5 37302.5 1747.5 37167.5 ;
      RECT  1897.5 37045.0 1962.5 36910.0 ;
      RECT  2280.0 37297.5 2415.0 37362.5 ;
      RECT  1497.5 37207.5 1562.5 37072.5 ;
      RECT  1897.5 37467.5 1962.5 37332.5 ;
      RECT  1897.5 36910.0 1962.5 37045.0 ;
      RECT  1682.5 37167.5 1747.5 37302.5 ;
      RECT  1897.5 37332.5 1962.5 37467.5 ;
      RECT  2657.5 36850.0 2722.5 37770.0 ;
      RECT  1312.5 36850.0 1377.5 37770.0 ;
      RECT  1507.5 38062.5 1312.5 38127.5 ;
      RECT  2347.5 38062.5 2722.5 38127.5 ;
      RECT  2347.5 38442.5 2722.5 38507.5 ;
      RECT  2505.0 38612.5 2690.0 38677.5 ;
      RECT  1345.0 38612.5 1530.0 38677.5 ;
      RECT  2347.5 38062.5 2482.5 38127.5 ;
      RECT  2347.5 38252.5 2482.5 38317.5 ;
      RECT  2347.5 38252.5 2482.5 38317.5 ;
      RECT  2347.5 38062.5 2482.5 38127.5 ;
      RECT  2347.5 38252.5 2482.5 38317.5 ;
      RECT  2347.5 38442.5 2482.5 38507.5 ;
      RECT  2347.5 38442.5 2482.5 38507.5 ;
      RECT  2347.5 38252.5 2482.5 38317.5 ;
      RECT  1507.5 38062.5 1642.5 38127.5 ;
      RECT  1507.5 38252.5 1642.5 38317.5 ;
      RECT  1507.5 38252.5 1642.5 38317.5 ;
      RECT  1507.5 38062.5 1642.5 38127.5 ;
      RECT  1507.5 38252.5 1642.5 38317.5 ;
      RECT  1507.5 38442.5 1642.5 38507.5 ;
      RECT  1507.5 38442.5 1642.5 38507.5 ;
      RECT  1507.5 38252.5 1642.5 38317.5 ;
      RECT  2437.5 38612.5 2572.5 38677.5 ;
      RECT  1462.5 38612.5 1597.5 38677.5 ;
      RECT  1737.5 38447.5 1802.5 38312.5 ;
      RECT  1952.5 38190.0 2017.5 38055.0 ;
      RECT  2347.5 38252.5 2482.5 38317.5 ;
      RECT  1507.5 38442.5 1642.5 38507.5 ;
      RECT  1952.5 38542.5 2017.5 38407.5 ;
      RECT  1952.5 38055.0 2017.5 38190.0 ;
      RECT  1737.5 38312.5 1802.5 38447.5 ;
      RECT  1952.5 38407.5 2017.5 38542.5 ;
      RECT  2657.5 37995.0 2722.5 38915.0 ;
      RECT  1312.5 37995.0 1377.5 38915.0 ;
      RECT  2505.0 39272.5 2690.0 39207.5 ;
      RECT  1345.0 39272.5 1530.0 39207.5 ;
      RECT  1462.5 39632.5 1312.5 39567.5 ;
      RECT  2347.5 39632.5 2722.5 39567.5 ;
      RECT  1462.5 39442.5 2347.5 39377.5 ;
      RECT  2347.5 39632.5 2482.5 39567.5 ;
      RECT  2347.5 39442.5 2482.5 39377.5 ;
      RECT  2347.5 39442.5 2482.5 39377.5 ;
      RECT  2347.5 39632.5 2482.5 39567.5 ;
      RECT  1462.5 39632.5 1597.5 39567.5 ;
      RECT  1462.5 39442.5 1597.5 39377.5 ;
      RECT  1462.5 39442.5 1597.5 39377.5 ;
      RECT  1462.5 39632.5 1597.5 39567.5 ;
      RECT  2437.5 39272.5 2572.5 39207.5 ;
      RECT  1462.5 39272.5 1597.5 39207.5 ;
      RECT  1905.0 39575.0 2040.0 39510.0 ;
      RECT  1905.0 39575.0 2040.0 39510.0 ;
      RECT  1940.0 39410.0 2005.0 39345.0 ;
      RECT  2657.5 39700.0 2722.5 39140.0 ;
      RECT  1312.5 39700.0 1377.5 39140.0 ;
      RECT  2505.0 39832.5 2690.0 39767.5 ;
      RECT  1345.0 39832.5 1530.0 39767.5 ;
      RECT  1462.5 40192.5 1312.5 40127.5 ;
      RECT  2347.5 40192.5 2722.5 40127.5 ;
      RECT  1462.5 40002.5 2347.5 39937.5 ;
      RECT  2347.5 40192.5 2482.5 40127.5 ;
      RECT  2347.5 40002.5 2482.5 39937.5 ;
      RECT  2347.5 40002.5 2482.5 39937.5 ;
      RECT  2347.5 40192.5 2482.5 40127.5 ;
      RECT  1462.5 40192.5 1597.5 40127.5 ;
      RECT  1462.5 40002.5 1597.5 39937.5 ;
      RECT  1462.5 40002.5 1597.5 39937.5 ;
      RECT  1462.5 40192.5 1597.5 40127.5 ;
      RECT  2437.5 39832.5 2572.5 39767.5 ;
      RECT  1462.5 39832.5 1597.5 39767.5 ;
      RECT  1905.0 40135.0 2040.0 40070.0 ;
      RECT  1905.0 40135.0 2040.0 40070.0 ;
      RECT  1940.0 39970.0 2005.0 39905.0 ;
      RECT  2657.5 40260.0 2722.5 39700.0 ;
      RECT  1312.5 40260.0 1377.5 39700.0 ;
      RECT  1182.5 37477.5 1377.5 37542.5 ;
      RECT  342.5 37477.5 -32.5 37542.5 ;
      RECT  342.5 37857.5 -32.5 37922.5 ;
      RECT  185.0 38217.5 8.881784197e-13 38282.5 ;
      RECT  1345.0 38217.5 1160.0 38282.5 ;
      RECT  342.5 37477.5 207.5 37542.5 ;
      RECT  342.5 37667.5 207.5 37732.5 ;
      RECT  342.5 37667.5 207.5 37732.5 ;
      RECT  342.5 37477.5 207.5 37542.5 ;
      RECT  342.5 37667.5 207.5 37732.5 ;
      RECT  342.5 37857.5 207.5 37922.5 ;
      RECT  342.5 37857.5 207.5 37922.5 ;
      RECT  342.5 37667.5 207.5 37732.5 ;
      RECT  342.5 37857.5 207.5 37922.5 ;
      RECT  342.5 38047.5 207.5 38112.5 ;
      RECT  342.5 38047.5 207.5 38112.5 ;
      RECT  342.5 37857.5 207.5 37922.5 ;
      RECT  1182.5 37477.5 1047.5 37542.5 ;
      RECT  1182.5 37667.5 1047.5 37732.5 ;
      RECT  1182.5 37667.5 1047.5 37732.5 ;
      RECT  1182.5 37477.5 1047.5 37542.5 ;
      RECT  1182.5 37667.5 1047.5 37732.5 ;
      RECT  1182.5 37857.5 1047.5 37922.5 ;
      RECT  1182.5 37857.5 1047.5 37922.5 ;
      RECT  1182.5 37667.5 1047.5 37732.5 ;
      RECT  1182.5 37857.5 1047.5 37922.5 ;
      RECT  1182.5 38047.5 1047.5 38112.5 ;
      RECT  1182.5 38047.5 1047.5 38112.5 ;
      RECT  1182.5 37857.5 1047.5 37922.5 ;
      RECT  252.5 38217.5 117.5 38282.5 ;
      RECT  1227.5 38217.5 1092.5 38282.5 ;
      RECT  970.0 38052.5 905.0 37917.5 ;
      RECT  830.0 37862.5 765.0 37727.5 ;
      RECT  690.0 37672.5 625.0 37537.5 ;
      RECT  342.5 37667.5 207.5 37732.5 ;
      RECT  342.5 38047.5 207.5 38112.5 ;
      RECT  1182.5 38047.5 1047.5 38112.5 ;
      RECT  725.0 38047.5 590.0 38112.5 ;
      RECT  690.0 37537.5 625.0 37672.5 ;
      RECT  830.0 37727.5 765.0 37862.5 ;
      RECT  970.0 37917.5 905.0 38052.5 ;
      RECT  725.0 38047.5 590.0 38112.5 ;
      RECT  32.5 37410.0 -32.5 38420.0 ;
      RECT  1377.5 37410.0 1312.5 38420.0 ;
      RECT  185.0 38847.5 8.881784197e-13 38912.5 ;
      RECT  1345.0 38847.5 1160.0 38912.5 ;
      RECT  1227.5 38487.5 1377.5 38552.5 ;
      RECT  342.5 38487.5 -32.5 38552.5 ;
      RECT  1227.5 38677.5 342.5 38742.5 ;
      RECT  342.5 38487.5 207.5 38552.5 ;
      RECT  342.5 38677.5 207.5 38742.5 ;
      RECT  342.5 38677.5 207.5 38742.5 ;
      RECT  342.5 38487.5 207.5 38552.5 ;
      RECT  1227.5 38487.5 1092.5 38552.5 ;
      RECT  1227.5 38677.5 1092.5 38742.5 ;
      RECT  1227.5 38677.5 1092.5 38742.5 ;
      RECT  1227.5 38487.5 1092.5 38552.5 ;
      RECT  252.5 38847.5 117.5 38912.5 ;
      RECT  1227.5 38847.5 1092.5 38912.5 ;
      RECT  785.0 38545.0 650.0 38610.0 ;
      RECT  785.0 38545.0 650.0 38610.0 ;
      RECT  750.0 38710.0 685.0 38775.0 ;
      RECT  32.5 38420.0 -32.5 38980.0 ;
      RECT  1377.5 38420.0 1312.5 38980.0 ;
      RECT  185.0 39407.5 8.881784197e-13 39472.5 ;
      RECT  1345.0 39407.5 1160.0 39472.5 ;
      RECT  1227.5 39047.5 1377.5 39112.5 ;
      RECT  342.5 39047.5 -32.5 39112.5 ;
      RECT  1227.5 39237.5 342.5 39302.5 ;
      RECT  342.5 39047.5 207.5 39112.5 ;
      RECT  342.5 39237.5 207.5 39302.5 ;
      RECT  342.5 39237.5 207.5 39302.5 ;
      RECT  342.5 39047.5 207.5 39112.5 ;
      RECT  1227.5 39047.5 1092.5 39112.5 ;
      RECT  1227.5 39237.5 1092.5 39302.5 ;
      RECT  1227.5 39237.5 1092.5 39302.5 ;
      RECT  1227.5 39047.5 1092.5 39112.5 ;
      RECT  252.5 39407.5 117.5 39472.5 ;
      RECT  1227.5 39407.5 1092.5 39472.5 ;
      RECT  785.0 39105.0 650.0 39170.0 ;
      RECT  785.0 39105.0 650.0 39170.0 ;
      RECT  750.0 39270.0 685.0 39335.0 ;
      RECT  32.5 38980.0 -32.5 39540.0 ;
      RECT  1377.5 38980.0 1312.5 39540.0 ;
      RECT  185.0 39967.5 8.881784197e-13 40032.5 ;
      RECT  1345.0 39967.5 1160.0 40032.5 ;
      RECT  1227.5 39607.5 1377.5 39672.5 ;
      RECT  342.5 39607.5 -32.5 39672.5 ;
      RECT  1227.5 39797.5 342.5 39862.5 ;
      RECT  342.5 39607.5 207.5 39672.5 ;
      RECT  342.5 39797.5 207.5 39862.5 ;
      RECT  342.5 39797.5 207.5 39862.5 ;
      RECT  342.5 39607.5 207.5 39672.5 ;
      RECT  1227.5 39607.5 1092.5 39672.5 ;
      RECT  1227.5 39797.5 1092.5 39862.5 ;
      RECT  1227.5 39797.5 1092.5 39862.5 ;
      RECT  1227.5 39607.5 1092.5 39672.5 ;
      RECT  252.5 39967.5 117.5 40032.5 ;
      RECT  1227.5 39967.5 1092.5 40032.5 ;
      RECT  785.0 39665.0 650.0 39730.0 ;
      RECT  785.0 39665.0 650.0 39730.0 ;
      RECT  750.0 39830.0 685.0 39895.0 ;
      RECT  32.5 39540.0 -32.5 40100.0 ;
      RECT  1377.5 39540.0 1312.5 40100.0 ;
      RECT  1377.5 47142.5 1312.5 60675.0 ;
      RECT  1312.5 42832.5 1025.0 42897.5 ;
      RECT  1312.5 45242.5 1025.0 45307.5 ;
      RECT  1312.5 45522.5 1025.0 45587.5 ;
      RECT  1312.5 47932.5 1025.0 47997.5 ;
      RECT  1312.5 48212.5 1025.0 48277.5 ;
      RECT  1312.5 50622.5 1025.0 50687.5 ;
      RECT  1312.5 50902.5 1025.0 50967.5 ;
      RECT  1312.5 53312.5 1025.0 53377.5 ;
      RECT  1312.5 53592.5 1025.0 53657.5 ;
      RECT  1312.5 56002.5 1025.0 56067.5 ;
      RECT  1312.5 56282.5 1025.0 56347.5 ;
      RECT  1312.5 58692.5 1025.0 58757.5 ;
      RECT  1312.5 58972.5 1025.0 59037.5 ;
      RECT  1377.5 40787.5 935.0 40852.5 ;
      RECT  935.0 40787.5 230.0 40852.5 ;
      RECT  20.0 44037.5 935.0 44102.5 ;
      RECT  20.0 46727.5 935.0 46792.5 ;
      RECT  20.0 49417.5 935.0 49482.5 ;
      RECT  20.0 52107.5 935.0 52172.5 ;
      RECT  20.0 54797.5 935.0 54862.5 ;
      RECT  20.0 57487.5 935.0 57552.5 ;
      RECT  20.0 60177.5 935.0 60242.5 ;
      RECT  20.0 41347.5 935.0 41412.5 ;
      RECT  2005.0 42360.0 1940.0 43060.0 ;
      RECT  2005.0 42552.5 1940.0 42617.5 ;
      RECT  2005.0 42360.0 1940.0 42585.0 ;
      RECT  1972.5 42552.5 1025.0 42617.5 ;
      RECT  2690.0 42422.5 2465.0 42487.5 ;
      RECT  2430.0 41552.5 2365.0 41617.5 ;
      RECT  2005.0 41552.5 1940.0 41617.5 ;
      RECT  2430.0 41585.0 2365.0 42232.5 ;
      RECT  2397.5 41552.5 1972.5 41617.5 ;
      RECT  2005.0 41255.0 1940.0 41585.0 ;
      RECT  1972.5 41552.5 1172.5 41617.5 ;
      RECT  1172.5 40955.0 750.0 41020.0 ;
      RECT  2040.0 41190.0 1905.0 41255.0 ;
      RECT  2005.0 43060.0 1940.0 43265.0 ;
      RECT  2505.0 40952.5 2690.0 40887.5 ;
      RECT  1345.0 40952.5 1530.0 40887.5 ;
      RECT  1462.5 41312.5 1312.5 41247.5 ;
      RECT  2347.5 41312.5 2722.5 41247.5 ;
      RECT  1462.5 41122.5 2347.5 41057.5 ;
      RECT  2347.5 41312.5 2482.5 41247.5 ;
      RECT  2347.5 41122.5 2482.5 41057.5 ;
      RECT  2347.5 41122.5 2482.5 41057.5 ;
      RECT  2347.5 41312.5 2482.5 41247.5 ;
      RECT  1462.5 41312.5 1597.5 41247.5 ;
      RECT  1462.5 41122.5 1597.5 41057.5 ;
      RECT  1462.5 41122.5 1597.5 41057.5 ;
      RECT  1462.5 41312.5 1597.5 41247.5 ;
      RECT  2437.5 40952.5 2572.5 40887.5 ;
      RECT  1462.5 40952.5 1597.5 40887.5 ;
      RECT  1905.0 41255.0 2040.0 41190.0 ;
      RECT  1905.0 41255.0 2040.0 41190.0 ;
      RECT  1940.0 41090.0 2005.0 41025.0 ;
      RECT  2657.5 41380.0 2722.5 40820.0 ;
      RECT  1312.5 41380.0 1377.5 40820.0 ;
      RECT  2330.0 42232.5 2465.0 42297.5 ;
      RECT  2330.0 42422.5 2465.0 42487.5 ;
      RECT  2330.0 42422.5 2465.0 42487.5 ;
      RECT  2330.0 42232.5 2465.0 42297.5 ;
      RECT  1312.5 47077.5 1377.5 47142.5 ;
      RECT  4002.5 47077.5 4067.5 47142.5 ;
      RECT  1312.5 46980.0 1377.5 47110.0 ;
      RECT  1345.0 47077.5 4035.0 47142.5 ;
      RECT  4002.5 46980.0 4067.5 47110.0 ;
      RECT  2875.0 43487.5 2690.0 43552.5 ;
      RECT  4035.0 43487.5 3850.0 43552.5 ;
      RECT  3917.5 43127.5 4067.5 43192.5 ;
      RECT  3032.5 43127.5 2657.5 43192.5 ;
      RECT  3917.5 43317.5 3032.5 43382.5 ;
      RECT  3032.5 43127.5 2897.5 43192.5 ;
      RECT  3032.5 43317.5 2897.5 43382.5 ;
      RECT  3032.5 43317.5 2897.5 43382.5 ;
      RECT  3032.5 43127.5 2897.5 43192.5 ;
      RECT  3917.5 43127.5 3782.5 43192.5 ;
      RECT  3917.5 43317.5 3782.5 43382.5 ;
      RECT  3917.5 43317.5 3782.5 43382.5 ;
      RECT  3917.5 43127.5 3782.5 43192.5 ;
      RECT  2942.5 43487.5 2807.5 43552.5 ;
      RECT  3917.5 43487.5 3782.5 43552.5 ;
      RECT  3475.0 43185.0 3340.0 43250.0 ;
      RECT  3475.0 43185.0 3340.0 43250.0 ;
      RECT  3440.0 43350.0 3375.0 43415.0 ;
      RECT  2722.5 43060.0 2657.5 43620.0 ;
      RECT  4067.5 43060.0 4002.5 43620.0 ;
      RECT  2875.0 44047.5 2690.0 44112.5 ;
      RECT  4035.0 44047.5 3850.0 44112.5 ;
      RECT  3917.5 43687.5 4067.5 43752.5 ;
      RECT  3032.5 43687.5 2657.5 43752.5 ;
      RECT  3917.5 43877.5 3032.5 43942.5 ;
      RECT  3032.5 43687.5 2897.5 43752.5 ;
      RECT  3032.5 43877.5 2897.5 43942.5 ;
      RECT  3032.5 43877.5 2897.5 43942.5 ;
      RECT  3032.5 43687.5 2897.5 43752.5 ;
      RECT  3917.5 43687.5 3782.5 43752.5 ;
      RECT  3917.5 43877.5 3782.5 43942.5 ;
      RECT  3917.5 43877.5 3782.5 43942.5 ;
      RECT  3917.5 43687.5 3782.5 43752.5 ;
      RECT  2942.5 44047.5 2807.5 44112.5 ;
      RECT  3917.5 44047.5 3782.5 44112.5 ;
      RECT  3475.0 43745.0 3340.0 43810.0 ;
      RECT  3475.0 43745.0 3340.0 43810.0 ;
      RECT  3440.0 43910.0 3375.0 43975.0 ;
      RECT  2722.5 43620.0 2657.5 44180.0 ;
      RECT  4067.5 43620.0 4002.5 44180.0 ;
      RECT  3340.0 43745.0 3475.0 43810.0 ;
      RECT  2875.0 44607.5 2690.0 44672.5 ;
      RECT  4035.0 44607.5 3850.0 44672.5 ;
      RECT  3917.5 44247.5 4067.5 44312.5 ;
      RECT  3032.5 44247.5 2657.5 44312.5 ;
      RECT  3917.5 44437.5 3032.5 44502.5 ;
      RECT  3032.5 44247.5 2897.5 44312.5 ;
      RECT  3032.5 44437.5 2897.5 44502.5 ;
      RECT  3032.5 44437.5 2897.5 44502.5 ;
      RECT  3032.5 44247.5 2897.5 44312.5 ;
      RECT  3917.5 44247.5 3782.5 44312.5 ;
      RECT  3917.5 44437.5 3782.5 44502.5 ;
      RECT  3917.5 44437.5 3782.5 44502.5 ;
      RECT  3917.5 44247.5 3782.5 44312.5 ;
      RECT  2942.5 44607.5 2807.5 44672.5 ;
      RECT  3917.5 44607.5 3782.5 44672.5 ;
      RECT  3475.0 44305.0 3340.0 44370.0 ;
      RECT  3475.0 44305.0 3340.0 44370.0 ;
      RECT  3440.0 44470.0 3375.0 44535.0 ;
      RECT  2722.5 44180.0 2657.5 44740.0 ;
      RECT  4067.5 44180.0 4002.5 44740.0 ;
      RECT  3340.0 44305.0 3475.0 44370.0 ;
      RECT  2875.0 45167.5 2690.0 45232.5 ;
      RECT  4035.0 45167.5 3850.0 45232.5 ;
      RECT  3917.5 44807.5 4067.5 44872.5 ;
      RECT  3032.5 44807.5 2657.5 44872.5 ;
      RECT  3917.5 44997.5 3032.5 45062.5 ;
      RECT  3032.5 44807.5 2897.5 44872.5 ;
      RECT  3032.5 44997.5 2897.5 45062.5 ;
      RECT  3032.5 44997.5 2897.5 45062.5 ;
      RECT  3032.5 44807.5 2897.5 44872.5 ;
      RECT  3917.5 44807.5 3782.5 44872.5 ;
      RECT  3917.5 44997.5 3782.5 45062.5 ;
      RECT  3917.5 44997.5 3782.5 45062.5 ;
      RECT  3917.5 44807.5 3782.5 44872.5 ;
      RECT  2942.5 45167.5 2807.5 45232.5 ;
      RECT  3917.5 45167.5 3782.5 45232.5 ;
      RECT  3475.0 44865.0 3340.0 44930.0 ;
      RECT  3475.0 44865.0 3340.0 44930.0 ;
      RECT  3440.0 45030.0 3375.0 45095.0 ;
      RECT  2722.5 44740.0 2657.5 45300.0 ;
      RECT  4067.5 44740.0 4002.5 45300.0 ;
      RECT  3340.0 44865.0 3475.0 44930.0 ;
      RECT  2875.0 45727.5 2690.0 45792.5 ;
      RECT  4035.0 45727.5 3850.0 45792.5 ;
      RECT  3917.5 45367.5 4067.5 45432.5 ;
      RECT  3032.5 45367.5 2657.5 45432.5 ;
      RECT  3917.5 45557.5 3032.5 45622.5 ;
      RECT  3032.5 45367.5 2897.5 45432.5 ;
      RECT  3032.5 45557.5 2897.5 45622.5 ;
      RECT  3032.5 45557.5 2897.5 45622.5 ;
      RECT  3032.5 45367.5 2897.5 45432.5 ;
      RECT  3917.5 45367.5 3782.5 45432.5 ;
      RECT  3917.5 45557.5 3782.5 45622.5 ;
      RECT  3917.5 45557.5 3782.5 45622.5 ;
      RECT  3917.5 45367.5 3782.5 45432.5 ;
      RECT  2942.5 45727.5 2807.5 45792.5 ;
      RECT  3917.5 45727.5 3782.5 45792.5 ;
      RECT  3475.0 45425.0 3340.0 45490.0 ;
      RECT  3475.0 45425.0 3340.0 45490.0 ;
      RECT  3440.0 45590.0 3375.0 45655.0 ;
      RECT  2722.5 45300.0 2657.5 45860.0 ;
      RECT  4067.5 45300.0 4002.5 45860.0 ;
      RECT  3340.0 45425.0 3475.0 45490.0 ;
      RECT  2875.0 46287.5 2690.0 46352.5 ;
      RECT  4035.0 46287.5 3850.0 46352.5 ;
      RECT  3917.5 45927.5 4067.5 45992.5 ;
      RECT  3032.5 45927.5 2657.5 45992.5 ;
      RECT  3917.5 46117.5 3032.5 46182.5 ;
      RECT  3032.5 45927.5 2897.5 45992.5 ;
      RECT  3032.5 46117.5 2897.5 46182.5 ;
      RECT  3032.5 46117.5 2897.5 46182.5 ;
      RECT  3032.5 45927.5 2897.5 45992.5 ;
      RECT  3917.5 45927.5 3782.5 45992.5 ;
      RECT  3917.5 46117.5 3782.5 46182.5 ;
      RECT  3917.5 46117.5 3782.5 46182.5 ;
      RECT  3917.5 45927.5 3782.5 45992.5 ;
      RECT  2942.5 46287.5 2807.5 46352.5 ;
      RECT  3917.5 46287.5 3782.5 46352.5 ;
      RECT  3475.0 45985.0 3340.0 46050.0 ;
      RECT  3475.0 45985.0 3340.0 46050.0 ;
      RECT  3440.0 46150.0 3375.0 46215.0 ;
      RECT  2722.5 45860.0 2657.5 46420.0 ;
      RECT  4067.5 45860.0 4002.5 46420.0 ;
      RECT  3340.0 45985.0 3475.0 46050.0 ;
      RECT  2875.0 46847.5 2690.0 46912.5 ;
      RECT  4035.0 46847.5 3850.0 46912.5 ;
      RECT  3917.5 46487.5 4067.5 46552.5 ;
      RECT  3032.5 46487.5 2657.5 46552.5 ;
      RECT  3917.5 46677.5 3032.5 46742.5 ;
      RECT  3032.5 46487.5 2897.5 46552.5 ;
      RECT  3032.5 46677.5 2897.5 46742.5 ;
      RECT  3032.5 46677.5 2897.5 46742.5 ;
      RECT  3032.5 46487.5 2897.5 46552.5 ;
      RECT  3917.5 46487.5 3782.5 46552.5 ;
      RECT  3917.5 46677.5 3782.5 46742.5 ;
      RECT  3917.5 46677.5 3782.5 46742.5 ;
      RECT  3917.5 46487.5 3782.5 46552.5 ;
      RECT  2942.5 46847.5 2807.5 46912.5 ;
      RECT  3917.5 46847.5 3782.5 46912.5 ;
      RECT  3475.0 46545.0 3340.0 46610.0 ;
      RECT  3475.0 46545.0 3340.0 46610.0 ;
      RECT  3440.0 46710.0 3375.0 46775.0 ;
      RECT  2722.5 46420.0 2657.5 46980.0 ;
      RECT  4067.5 46420.0 4002.5 46980.0 ;
      RECT  3340.0 46545.0 3475.0 46610.0 ;
      RECT  2505.0 45992.5 2690.0 45927.5 ;
      RECT  1345.0 45992.5 1530.0 45927.5 ;
      RECT  1462.5 46352.5 1312.5 46287.5 ;
      RECT  2347.5 46352.5 2722.5 46287.5 ;
      RECT  1462.5 46162.5 2347.5 46097.5 ;
      RECT  2347.5 46352.5 2482.5 46287.5 ;
      RECT  2347.5 46162.5 2482.5 46097.5 ;
      RECT  2347.5 46162.5 2482.5 46097.5 ;
      RECT  2347.5 46352.5 2482.5 46287.5 ;
      RECT  1462.5 46352.5 1597.5 46287.5 ;
      RECT  1462.5 46162.5 1597.5 46097.5 ;
      RECT  1462.5 46162.5 1597.5 46097.5 ;
      RECT  1462.5 46352.5 1597.5 46287.5 ;
      RECT  2437.5 45992.5 2572.5 45927.5 ;
      RECT  1462.5 45992.5 1597.5 45927.5 ;
      RECT  1905.0 46295.0 2040.0 46230.0 ;
      RECT  1905.0 46295.0 2040.0 46230.0 ;
      RECT  1940.0 46130.0 2005.0 46065.0 ;
      RECT  2657.5 46420.0 2722.5 45860.0 ;
      RECT  1312.5 46420.0 1377.5 45860.0 ;
      RECT  1905.0 46230.0 2040.0 46295.0 ;
      RECT  2505.0 45432.5 2690.0 45367.5 ;
      RECT  1345.0 45432.5 1530.0 45367.5 ;
      RECT  1462.5 45792.5 1312.5 45727.5 ;
      RECT  2347.5 45792.5 2722.5 45727.5 ;
      RECT  1462.5 45602.5 2347.5 45537.5 ;
      RECT  2347.5 45792.5 2482.5 45727.5 ;
      RECT  2347.5 45602.5 2482.5 45537.5 ;
      RECT  2347.5 45602.5 2482.5 45537.5 ;
      RECT  2347.5 45792.5 2482.5 45727.5 ;
      RECT  1462.5 45792.5 1597.5 45727.5 ;
      RECT  1462.5 45602.5 1597.5 45537.5 ;
      RECT  1462.5 45602.5 1597.5 45537.5 ;
      RECT  1462.5 45792.5 1597.5 45727.5 ;
      RECT  2437.5 45432.5 2572.5 45367.5 ;
      RECT  1462.5 45432.5 1597.5 45367.5 ;
      RECT  1905.0 45735.0 2040.0 45670.0 ;
      RECT  1905.0 45735.0 2040.0 45670.0 ;
      RECT  1940.0 45570.0 2005.0 45505.0 ;
      RECT  2657.5 45860.0 2722.5 45300.0 ;
      RECT  1312.5 45860.0 1377.5 45300.0 ;
      RECT  1905.0 45670.0 2040.0 45735.0 ;
      RECT  2505.0 44872.5 2690.0 44807.5 ;
      RECT  1345.0 44872.5 1530.0 44807.5 ;
      RECT  1462.5 45232.5 1312.5 45167.5 ;
      RECT  2347.5 45232.5 2722.5 45167.5 ;
      RECT  1462.5 45042.5 2347.5 44977.5 ;
      RECT  2347.5 45232.5 2482.5 45167.5 ;
      RECT  2347.5 45042.5 2482.5 44977.5 ;
      RECT  2347.5 45042.5 2482.5 44977.5 ;
      RECT  2347.5 45232.5 2482.5 45167.5 ;
      RECT  1462.5 45232.5 1597.5 45167.5 ;
      RECT  1462.5 45042.5 1597.5 44977.5 ;
      RECT  1462.5 45042.5 1597.5 44977.5 ;
      RECT  1462.5 45232.5 1597.5 45167.5 ;
      RECT  2437.5 44872.5 2572.5 44807.5 ;
      RECT  1462.5 44872.5 1597.5 44807.5 ;
      RECT  1905.0 45175.0 2040.0 45110.0 ;
      RECT  1905.0 45175.0 2040.0 45110.0 ;
      RECT  1940.0 45010.0 2005.0 44945.0 ;
      RECT  2657.5 45300.0 2722.5 44740.0 ;
      RECT  1312.5 45300.0 1377.5 44740.0 ;
      RECT  1905.0 45110.0 2040.0 45175.0 ;
      RECT  2505.0 44312.5 2690.0 44247.5 ;
      RECT  1345.0 44312.5 1530.0 44247.5 ;
      RECT  1462.5 44672.5 1312.5 44607.5 ;
      RECT  2347.5 44672.5 2722.5 44607.5 ;
      RECT  1462.5 44482.5 2347.5 44417.5 ;
      RECT  2347.5 44672.5 2482.5 44607.5 ;
      RECT  2347.5 44482.5 2482.5 44417.5 ;
      RECT  2347.5 44482.5 2482.5 44417.5 ;
      RECT  2347.5 44672.5 2482.5 44607.5 ;
      RECT  1462.5 44672.5 1597.5 44607.5 ;
      RECT  1462.5 44482.5 1597.5 44417.5 ;
      RECT  1462.5 44482.5 1597.5 44417.5 ;
      RECT  1462.5 44672.5 1597.5 44607.5 ;
      RECT  2437.5 44312.5 2572.5 44247.5 ;
      RECT  1462.5 44312.5 1597.5 44247.5 ;
      RECT  1905.0 44615.0 2040.0 44550.0 ;
      RECT  1905.0 44615.0 2040.0 44550.0 ;
      RECT  1940.0 44450.0 2005.0 44385.0 ;
      RECT  2657.5 44740.0 2722.5 44180.0 ;
      RECT  1312.5 44740.0 1377.5 44180.0 ;
      RECT  1905.0 44550.0 2040.0 44615.0 ;
      RECT  2505.0 43752.5 2690.0 43687.5 ;
      RECT  1345.0 43752.5 1530.0 43687.5 ;
      RECT  1462.5 44112.5 1312.5 44047.5 ;
      RECT  2347.5 44112.5 2722.5 44047.5 ;
      RECT  1462.5 43922.5 2347.5 43857.5 ;
      RECT  2347.5 44112.5 2482.5 44047.5 ;
      RECT  2347.5 43922.5 2482.5 43857.5 ;
      RECT  2347.5 43922.5 2482.5 43857.5 ;
      RECT  2347.5 44112.5 2482.5 44047.5 ;
      RECT  1462.5 44112.5 1597.5 44047.5 ;
      RECT  1462.5 43922.5 1597.5 43857.5 ;
      RECT  1462.5 43922.5 1597.5 43857.5 ;
      RECT  1462.5 44112.5 1597.5 44047.5 ;
      RECT  2437.5 43752.5 2572.5 43687.5 ;
      RECT  1462.5 43752.5 1597.5 43687.5 ;
      RECT  1905.0 44055.0 2040.0 43990.0 ;
      RECT  1905.0 44055.0 2040.0 43990.0 ;
      RECT  1940.0 43890.0 2005.0 43825.0 ;
      RECT  2657.5 44180.0 2722.5 43620.0 ;
      RECT  1312.5 44180.0 1377.5 43620.0 ;
      RECT  1905.0 43990.0 2040.0 44055.0 ;
      RECT  2505.0 43192.5 2690.0 43127.5 ;
      RECT  1345.0 43192.5 1530.0 43127.5 ;
      RECT  1462.5 43552.5 1312.5 43487.5 ;
      RECT  2347.5 43552.5 2722.5 43487.5 ;
      RECT  1462.5 43362.5 2347.5 43297.5 ;
      RECT  2347.5 43552.5 2482.5 43487.5 ;
      RECT  2347.5 43362.5 2482.5 43297.5 ;
      RECT  2347.5 43362.5 2482.5 43297.5 ;
      RECT  2347.5 43552.5 2482.5 43487.5 ;
      RECT  1462.5 43552.5 1597.5 43487.5 ;
      RECT  1462.5 43362.5 1597.5 43297.5 ;
      RECT  1462.5 43362.5 1597.5 43297.5 ;
      RECT  1462.5 43552.5 1597.5 43487.5 ;
      RECT  2437.5 43192.5 2572.5 43127.5 ;
      RECT  1462.5 43192.5 1597.5 43127.5 ;
      RECT  1905.0 43495.0 2040.0 43430.0 ;
      RECT  1905.0 43495.0 2040.0 43430.0 ;
      RECT  1940.0 43330.0 2005.0 43265.0 ;
      RECT  2657.5 43620.0 2722.5 43060.0 ;
      RECT  1312.5 43620.0 1377.5 43060.0 ;
      RECT  1905.0 43430.0 2040.0 43495.0 ;
      RECT  3340.0 43350.0 3475.0 43415.0 ;
      RECT  3340.0 45030.0 3475.0 45095.0 ;
      RECT  3340.0 46710.0 3475.0 46775.0 ;
      RECT  1905.0 44945.0 2040.0 45010.0 ;
      RECT  3340.0 43185.0 3475.0 43250.0 ;
      RECT  1940.0 43060.0 2005.0 43265.0 ;
      RECT  2657.5 43060.0 2722.5 46980.0 ;
      RECT  1312.5 43060.0 1377.5 46980.0 ;
      RECT  4002.5 43060.0 4067.5 46980.0 ;
      RECT  935.0 42725.0 225.0 41380.0 ;
      RECT  935.0 42725.0 230.0 44070.0 ;
      RECT  935.0 45415.0 230.0 44070.0 ;
      RECT  935.0 45415.0 230.0 46760.0 ;
      RECT  935.0 48105.0 230.0 46760.0 ;
      RECT  935.0 48105.0 230.0 49450.0 ;
      RECT  935.0 50795.0 230.0 49450.0 ;
      RECT  935.0 50795.0 230.0 52140.0 ;
      RECT  935.0 53485.0 230.0 52140.0 ;
      RECT  935.0 53485.0 230.0 54830.0 ;
      RECT  935.0 56175.0 230.0 54830.0 ;
      RECT  935.0 56175.0 230.0 57520.0 ;
      RECT  935.0 58865.0 230.0 57520.0 ;
      RECT  935.0 58865.0 230.0 60210.0 ;
      RECT  1025.0 42832.5 140.0 42897.5 ;
      RECT  1025.0 45242.5 140.0 45307.5 ;
      RECT  1025.0 45522.5 140.0 45587.5 ;
      RECT  1025.0 47932.5 140.0 47997.5 ;
      RECT  1025.0 48212.5 140.0 48277.5 ;
      RECT  1025.0 50622.5 140.0 50687.5 ;
      RECT  1025.0 50902.5 140.0 50967.5 ;
      RECT  1025.0 53312.5 140.0 53377.5 ;
      RECT  1025.0 53592.5 140.0 53657.5 ;
      RECT  1025.0 56002.5 140.0 56067.5 ;
      RECT  1025.0 56282.5 140.0 56347.5 ;
      RECT  1025.0 58692.5 140.0 58757.5 ;
      RECT  1025.0 58972.5 140.0 59037.5 ;
      RECT  1025.0 44037.5 140.0 44102.5 ;
      RECT  1025.0 46727.5 140.0 46792.5 ;
      RECT  1025.0 49417.5 140.0 49482.5 ;
      RECT  1025.0 52107.5 140.0 52172.5 ;
      RECT  1025.0 54797.5 140.0 54862.5 ;
      RECT  1025.0 57487.5 140.0 57552.5 ;
      RECT  1025.0 60177.5 140.0 60242.5 ;
      RECT  1025.0 42692.5 140.0 42757.5 ;
      RECT  1025.0 45382.5 140.0 45447.5 ;
      RECT  1025.0 48072.5 140.0 48137.5 ;
      RECT  1025.0 50762.5 140.0 50827.5 ;
      RECT  1025.0 53452.5 140.0 53517.5 ;
      RECT  1025.0 56142.5 140.0 56207.5 ;
      RECT  1025.0 58832.5 140.0 58897.5 ;
      RECT  1345.0 42797.5 1280.0 42932.5 ;
      RECT  1345.0 45207.5 1280.0 45342.5 ;
      RECT  1345.0 45487.5 1280.0 45622.5 ;
      RECT  1345.0 47897.5 1280.0 48032.5 ;
      RECT  1345.0 48177.5 1280.0 48312.5 ;
      RECT  1345.0 50587.5 1280.0 50722.5 ;
      RECT  1345.0 50867.5 1280.0 51002.5 ;
      RECT  1345.0 53277.5 1280.0 53412.5 ;
      RECT  1345.0 53557.5 1280.0 53692.5 ;
      RECT  1345.0 55967.5 1280.0 56102.5 ;
      RECT  1345.0 56247.5 1280.0 56382.5 ;
      RECT  1345.0 58657.5 1280.0 58792.5 ;
      RECT  1345.0 58937.5 1280.0 59072.5 ;
      RECT  1342.5 43060.0 1277.5 43195.0 ;
      RECT  1377.5 40685.0 1312.5 40820.0 ;
      RECT  867.5 40787.5 1002.5 40852.5 ;
      RECT  162.5 40787.5 297.5 40852.5 ;
      RECT  2005.0 42292.5 1940.0 42427.5 ;
      RECT  1105.0 41552.5 1240.0 41617.5 ;
      RECT  1105.0 40955.0 1240.0 41020.0 ;
      RECT  682.5 40955.0 817.5 41020.0 ;
      RECT  3475.0 40260.0 3410.0 43185.0 ;
      RECT  2005.0 40260.0 1940.0 41025.0 ;
      RECT  20.0 40260.0 -45.0 60297.5 ;
      RECT  2722.5 40260.0 2657.5 43060.0 ;
      RECT  1377.5 40260.0 1312.5 40820.0 ;
      RECT  4067.5 40260.0 4002.5 43060.0 ;
      RECT  3455.0 35107.5 3390.0 34972.5 ;
      RECT  3455.0 31027.5 3390.0 30892.5 ;
      RECT  2517.5 28460.0 2452.5 28325.0 ;
      RECT  1962.5 35107.5 1897.5 34972.5 ;
      RECT  1747.5 35517.5 1682.5 35382.5 ;
      RECT  2017.5 38055.0 1952.5 37920.0 ;
      RECT  1802.5 38312.5 1737.5 38177.5 ;
      RECT  3380.0 36542.5 3315.0 36407.5 ;
      RECT  3520.0 36337.5 3455.0 36202.5 ;
      RECT  3660.0 35722.5 3595.0 35587.5 ;
      RECT  690.0 36542.5 625.0 36407.5 ;
      RECT  830.0 35722.5 765.0 35587.5 ;
      RECT  970.0 35927.5 905.0 35792.5 ;
      RECT  1997.5 37737.5 1862.5 37802.5 ;
      RECT  2052.5 38882.5 1917.5 38947.5 ;
      RECT  785.0 40067.5 650.0 40132.5 ;
      RECT  2040.0 39107.5 1905.0 39172.5 ;
      RECT  4067.5 35312.5 4002.5 35177.5 ;
      RECT  2722.5 36132.5 2657.5 35997.5 ;
      RECT  1377.5 35312.5 1312.5 35177.5 ;
      RECT  32.5 36132.5 -32.5 35997.5 ;
      RECT  3475.0 28155.0 3340.0 28345.0 ;
      RECT  2722.5 28155.0 2657.5 28220.0 ;
      RECT  4067.5 28155.0 4002.5 28220.0 ;
      RECT  4417.5 36032.5 4282.5 36097.5 ;
   LAYER  metal2 ;
      RECT  15237.5 38935.0 15307.5 39140.0 ;
      RECT  15032.5 39895.0 15102.5 40100.0 ;
      RECT  14622.5 37565.0 14692.5 37770.0 ;
      RECT  14417.5 38710.0 14487.5 38915.0 ;
      RECT  14827.5 36270.0 14897.5 36475.0 ;
      RECT  14212.5 34835.0 14282.5 35040.0 ;
      RECT  4035.0 36030.0 4350.0 36100.0 ;
      RECT  13797.5 35040.0 13867.5 35245.0 ;
      RECT  14212.5 35.0 14282.5 115822.5 ;
      RECT  14417.5 35.0 14487.5 115822.5 ;
      RECT  14622.5 35.0 14692.5 115822.5 ;
      RECT  14827.5 35.0 14897.5 115822.5 ;
      RECT  15032.5 35.0 15102.5 115822.5 ;
      RECT  15237.5 35.0 15307.5 115822.5 ;
      RECT  11402.5 35.0 11472.5 28015.0 ;
      RECT  11607.5 35.0 11677.5 28015.0 ;
      RECT  11812.5 35.0 11882.5 28015.0 ;
      RECT  12017.5 35.0 12087.5 28015.0 ;
      RECT  12222.5 35.0 12292.5 28015.0 ;
      RECT  12427.5 35.0 12497.5 28015.0 ;
      RECT  12632.5 35.0 12702.5 28015.0 ;
      RECT  12837.5 35.0 12907.5 28015.0 ;
      RECT  13042.5 35.0 13112.5 28015.0 ;
      RECT  13247.5 35.0 13317.5 28015.0 ;
      RECT  15900.0 114250.0 15970.0 114655.0 ;
      RECT  16235.0 114250.0 16305.0 114655.0 ;
      RECT  16605.0 114250.0 16675.0 114655.0 ;
      RECT  16940.0 114250.0 17010.0 114655.0 ;
      RECT  17310.0 114250.0 17380.0 114655.0 ;
      RECT  17645.0 114250.0 17715.0 114655.0 ;
      RECT  18015.0 114250.0 18085.0 114655.0 ;
      RECT  18350.0 114250.0 18420.0 114655.0 ;
      RECT  18720.0 114250.0 18790.0 114655.0 ;
      RECT  19055.0 114250.0 19125.0 114655.0 ;
      RECT  19425.0 114250.0 19495.0 114655.0 ;
      RECT  19760.0 114250.0 19830.0 114655.0 ;
      RECT  20130.0 114250.0 20200.0 114655.0 ;
      RECT  20465.0 114250.0 20535.0 114655.0 ;
      RECT  20835.0 114250.0 20905.0 114655.0 ;
      RECT  21170.0 114250.0 21240.0 114655.0 ;
      RECT  21540.0 114250.0 21610.0 114655.0 ;
      RECT  21875.0 114250.0 21945.0 114655.0 ;
      RECT  22245.0 114250.0 22315.0 114655.0 ;
      RECT  22580.0 114250.0 22650.0 114655.0 ;
      RECT  22950.0 114250.0 23020.0 114655.0 ;
      RECT  23285.0 114250.0 23355.0 114655.0 ;
      RECT  23655.0 114250.0 23725.0 114655.0 ;
      RECT  23990.0 114250.0 24060.0 114655.0 ;
      RECT  24360.0 114250.0 24430.0 114655.0 ;
      RECT  24695.0 114250.0 24765.0 114655.0 ;
      RECT  25065.0 114250.0 25135.0 114655.0 ;
      RECT  25400.0 114250.0 25470.0 114655.0 ;
      RECT  25770.0 114250.0 25840.0 114655.0 ;
      RECT  26105.0 114250.0 26175.0 114655.0 ;
      RECT  26475.0 114250.0 26545.0 114655.0 ;
      RECT  26810.0 114250.0 26880.0 114655.0 ;
      RECT  27180.0 114250.0 27250.0 114655.0 ;
      RECT  27515.0 114250.0 27585.0 114655.0 ;
      RECT  27885.0 114250.0 27955.0 114655.0 ;
      RECT  28220.0 114250.0 28290.0 114655.0 ;
      RECT  28590.0 114250.0 28660.0 114655.0 ;
      RECT  28925.0 114250.0 28995.0 114655.0 ;
      RECT  29295.0 114250.0 29365.0 114655.0 ;
      RECT  29630.0 114250.0 29700.0 114655.0 ;
      RECT  30000.0 114250.0 30070.0 114655.0 ;
      RECT  30335.0 114250.0 30405.0 114655.0 ;
      RECT  30705.0 114250.0 30775.0 114655.0 ;
      RECT  31040.0 114250.0 31110.0 114655.0 ;
      RECT  31410.0 114250.0 31480.0 114655.0 ;
      RECT  31745.0 114250.0 31815.0 114655.0 ;
      RECT  32115.0 114250.0 32185.0 114655.0 ;
      RECT  32450.0 114250.0 32520.0 114655.0 ;
      RECT  32820.0 114250.0 32890.0 114655.0 ;
      RECT  33155.0 114250.0 33225.0 114655.0 ;
      RECT  33525.0 114250.0 33595.0 114655.0 ;
      RECT  33860.0 114250.0 33930.0 114655.0 ;
      RECT  34230.0 114250.0 34300.0 114655.0 ;
      RECT  34565.0 114250.0 34635.0 114655.0 ;
      RECT  34935.0 114250.0 35005.0 114655.0 ;
      RECT  35270.0 114250.0 35340.0 114655.0 ;
      RECT  35640.0 114250.0 35710.0 114655.0 ;
      RECT  35975.0 114250.0 36045.0 114655.0 ;
      RECT  36345.0 114250.0 36415.0 114655.0 ;
      RECT  36680.0 114250.0 36750.0 114655.0 ;
      RECT  37050.0 114250.0 37120.0 114655.0 ;
      RECT  37385.0 114250.0 37455.0 114655.0 ;
      RECT  37755.0 114250.0 37825.0 114655.0 ;
      RECT  38090.0 114250.0 38160.0 114655.0 ;
      RECT  38460.0 114250.0 38530.0 114655.0 ;
      RECT  38795.0 114250.0 38865.0 114655.0 ;
      RECT  39165.0 114250.0 39235.0 114655.0 ;
      RECT  39500.0 114250.0 39570.0 114655.0 ;
      RECT  39870.0 114250.0 39940.0 114655.0 ;
      RECT  40205.0 114250.0 40275.0 114655.0 ;
      RECT  40575.0 114250.0 40645.0 114655.0 ;
      RECT  40910.0 114250.0 40980.0 114655.0 ;
      RECT  41280.0 114250.0 41350.0 114655.0 ;
      RECT  41615.0 114250.0 41685.0 114655.0 ;
      RECT  41985.0 114250.0 42055.0 114655.0 ;
      RECT  42320.0 114250.0 42390.0 114655.0 ;
      RECT  42690.0 114250.0 42760.0 114655.0 ;
      RECT  43025.0 114250.0 43095.0 114655.0 ;
      RECT  43395.0 114250.0 43465.0 114655.0 ;
      RECT  43730.0 114250.0 43800.0 114655.0 ;
      RECT  44100.0 114250.0 44170.0 114655.0 ;
      RECT  44435.0 114250.0 44505.0 114655.0 ;
      RECT  44805.0 114250.0 44875.0 114655.0 ;
      RECT  45140.0 114250.0 45210.0 114655.0 ;
      RECT  45510.0 114250.0 45580.0 114655.0 ;
      RECT  45845.0 114250.0 45915.0 114655.0 ;
      RECT  46215.0 114250.0 46285.0 114655.0 ;
      RECT  46550.0 114250.0 46620.0 114655.0 ;
      RECT  46920.0 114250.0 46990.0 114655.0 ;
      RECT  47255.0 114250.0 47325.0 114655.0 ;
      RECT  47625.0 114250.0 47695.0 114655.0 ;
      RECT  47960.0 114250.0 48030.0 114655.0 ;
      RECT  48330.0 114250.0 48400.0 114655.0 ;
      RECT  48665.0 114250.0 48735.0 114655.0 ;
      RECT  49035.0 114250.0 49105.0 114655.0 ;
      RECT  49370.0 114250.0 49440.0 114655.0 ;
      RECT  49740.0 114250.0 49810.0 114655.0 ;
      RECT  50075.0 114250.0 50145.0 114655.0 ;
      RECT  50445.0 114250.0 50515.0 114655.0 ;
      RECT  50780.0 114250.0 50850.0 114655.0 ;
      RECT  51150.0 114250.0 51220.0 114655.0 ;
      RECT  51485.0 114250.0 51555.0 114655.0 ;
      RECT  51855.0 114250.0 51925.0 114655.0 ;
      RECT  52190.0 114250.0 52260.0 114655.0 ;
      RECT  52560.0 114250.0 52630.0 114655.0 ;
      RECT  52895.0 114250.0 52965.0 114655.0 ;
      RECT  53265.0 114250.0 53335.0 114655.0 ;
      RECT  53600.0 114250.0 53670.0 114655.0 ;
      RECT  53970.0 114250.0 54040.0 114655.0 ;
      RECT  54305.0 114250.0 54375.0 114655.0 ;
      RECT  54675.0 114250.0 54745.0 114655.0 ;
      RECT  55010.0 114250.0 55080.0 114655.0 ;
      RECT  55380.0 114250.0 55450.0 114655.0 ;
      RECT  55715.0 114250.0 55785.0 114655.0 ;
      RECT  56085.0 114250.0 56155.0 114655.0 ;
      RECT  56420.0 114250.0 56490.0 114655.0 ;
      RECT  56790.0 114250.0 56860.0 114655.0 ;
      RECT  57125.0 114250.0 57195.0 114655.0 ;
      RECT  57495.0 114250.0 57565.0 114655.0 ;
      RECT  57830.0 114250.0 57900.0 114655.0 ;
      RECT  58200.0 114250.0 58270.0 114655.0 ;
      RECT  58535.0 114250.0 58605.0 114655.0 ;
      RECT  58905.0 114250.0 58975.0 114655.0 ;
      RECT  59240.0 114250.0 59310.0 114655.0 ;
      RECT  59610.0 114250.0 59680.0 114655.0 ;
      RECT  59945.0 114250.0 60015.0 114655.0 ;
      RECT  60315.0 114250.0 60385.0 114655.0 ;
      RECT  60650.0 114250.0 60720.0 114655.0 ;
      RECT  61020.0 114250.0 61090.0 114655.0 ;
      RECT  61355.0 114250.0 61425.0 114655.0 ;
      RECT  61725.0 114250.0 61795.0 114655.0 ;
      RECT  62060.0 114250.0 62130.0 114655.0 ;
      RECT  62430.0 114250.0 62500.0 114655.0 ;
      RECT  62765.0 114250.0 62835.0 114655.0 ;
      RECT  63135.0 114250.0 63205.0 114655.0 ;
      RECT  63470.0 114250.0 63540.0 114655.0 ;
      RECT  63840.0 114250.0 63910.0 114655.0 ;
      RECT  64175.0 114250.0 64245.0 114655.0 ;
      RECT  64545.0 114250.0 64615.0 114655.0 ;
      RECT  64880.0 114250.0 64950.0 114655.0 ;
      RECT  65250.0 114250.0 65320.0 114655.0 ;
      RECT  65585.0 114250.0 65655.0 114655.0 ;
      RECT  65955.0 114250.0 66025.0 114655.0 ;
      RECT  66290.0 114250.0 66360.0 114655.0 ;
      RECT  66660.0 114250.0 66730.0 114655.0 ;
      RECT  66995.0 114250.0 67065.0 114655.0 ;
      RECT  67365.0 114250.0 67435.0 114655.0 ;
      RECT  67700.0 114250.0 67770.0 114655.0 ;
      RECT  68070.0 114250.0 68140.0 114655.0 ;
      RECT  68405.0 114250.0 68475.0 114655.0 ;
      RECT  68775.0 114250.0 68845.0 114655.0 ;
      RECT  69110.0 114250.0 69180.0 114655.0 ;
      RECT  69480.0 114250.0 69550.0 114655.0 ;
      RECT  69815.0 114250.0 69885.0 114655.0 ;
      RECT  70185.0 114250.0 70255.0 114655.0 ;
      RECT  70520.0 114250.0 70590.0 114655.0 ;
      RECT  70890.0 114250.0 70960.0 114655.0 ;
      RECT  71225.0 114250.0 71295.0 114655.0 ;
      RECT  71595.0 114250.0 71665.0 114655.0 ;
      RECT  71930.0 114250.0 72000.0 114655.0 ;
      RECT  72300.0 114250.0 72370.0 114655.0 ;
      RECT  72635.0 114250.0 72705.0 114655.0 ;
      RECT  73005.0 114250.0 73075.0 114655.0 ;
      RECT  73340.0 114250.0 73410.0 114655.0 ;
      RECT  73710.0 114250.0 73780.0 114655.0 ;
      RECT  74045.0 114250.0 74115.0 114655.0 ;
      RECT  74415.0 114250.0 74485.0 114655.0 ;
      RECT  74750.0 114250.0 74820.0 114655.0 ;
      RECT  75120.0 114250.0 75190.0 114655.0 ;
      RECT  75455.0 114250.0 75525.0 114655.0 ;
      RECT  75825.0 114250.0 75895.0 114655.0 ;
      RECT  76160.0 114250.0 76230.0 114655.0 ;
      RECT  76530.0 114250.0 76600.0 114655.0 ;
      RECT  76865.0 114250.0 76935.0 114655.0 ;
      RECT  77235.0 114250.0 77305.0 114655.0 ;
      RECT  77570.0 114250.0 77640.0 114655.0 ;
      RECT  77940.0 114250.0 78010.0 114655.0 ;
      RECT  78275.0 114250.0 78345.0 114655.0 ;
      RECT  78645.0 114250.0 78715.0 114655.0 ;
      RECT  78980.0 114250.0 79050.0 114655.0 ;
      RECT  79350.0 114250.0 79420.0 114655.0 ;
      RECT  79685.0 114250.0 79755.0 114655.0 ;
      RECT  80055.0 114250.0 80125.0 114655.0 ;
      RECT  80390.0 114250.0 80460.0 114655.0 ;
      RECT  80760.0 114250.0 80830.0 114655.0 ;
      RECT  81095.0 114250.0 81165.0 114655.0 ;
      RECT  81465.0 114250.0 81535.0 114655.0 ;
      RECT  81800.0 114250.0 81870.0 114655.0 ;
      RECT  82170.0 114250.0 82240.0 114655.0 ;
      RECT  82505.0 114250.0 82575.0 114655.0 ;
      RECT  82875.0 114250.0 82945.0 114655.0 ;
      RECT  83210.0 114250.0 83280.0 114655.0 ;
      RECT  83580.0 114250.0 83650.0 114655.0 ;
      RECT  83915.0 114250.0 83985.0 114655.0 ;
      RECT  84285.0 114250.0 84355.0 114655.0 ;
      RECT  84620.0 114250.0 84690.0 114655.0 ;
      RECT  84990.0 114250.0 85060.0 114655.0 ;
      RECT  85325.0 114250.0 85395.0 114655.0 ;
      RECT  85695.0 114250.0 85765.0 114655.0 ;
      RECT  86030.0 114250.0 86100.0 114655.0 ;
      RECT  86400.0 114250.0 86470.0 114655.0 ;
      RECT  86735.0 114250.0 86805.0 114655.0 ;
      RECT  87105.0 114250.0 87175.0 114655.0 ;
      RECT  87440.0 114250.0 87510.0 114655.0 ;
      RECT  87810.0 114250.0 87880.0 114655.0 ;
      RECT  88145.0 114250.0 88215.0 114655.0 ;
      RECT  88515.0 114250.0 88585.0 114655.0 ;
      RECT  88850.0 114250.0 88920.0 114655.0 ;
      RECT  89220.0 114250.0 89290.0 114655.0 ;
      RECT  89555.0 114250.0 89625.0 114655.0 ;
      RECT  89925.0 114250.0 89995.0 114655.0 ;
      RECT  90260.0 114250.0 90330.0 114655.0 ;
      RECT  90630.0 114250.0 90700.0 114655.0 ;
      RECT  90965.0 114250.0 91035.0 114655.0 ;
      RECT  91335.0 114250.0 91405.0 114655.0 ;
      RECT  91670.0 114250.0 91740.0 114655.0 ;
      RECT  92040.0 114250.0 92110.0 114655.0 ;
      RECT  92375.0 114250.0 92445.0 114655.0 ;
      RECT  92745.0 114250.0 92815.0 114655.0 ;
      RECT  93080.0 114250.0 93150.0 114655.0 ;
      RECT  93450.0 114250.0 93520.0 114655.0 ;
      RECT  93785.0 114250.0 93855.0 114655.0 ;
      RECT  94155.0 114250.0 94225.0 114655.0 ;
      RECT  94490.0 114250.0 94560.0 114655.0 ;
      RECT  94860.0 114250.0 94930.0 114655.0 ;
      RECT  95195.0 114250.0 95265.0 114655.0 ;
      RECT  95565.0 114250.0 95635.0 114655.0 ;
      RECT  95900.0 114250.0 95970.0 114655.0 ;
      RECT  96270.0 114250.0 96340.0 114655.0 ;
      RECT  96605.0 114250.0 96675.0 114655.0 ;
      RECT  96975.0 114250.0 97045.0 114655.0 ;
      RECT  97310.0 114250.0 97380.0 114655.0 ;
      RECT  97680.0 114250.0 97750.0 114655.0 ;
      RECT  98015.0 114250.0 98085.0 114655.0 ;
      RECT  98385.0 114250.0 98455.0 114655.0 ;
      RECT  98720.0 114250.0 98790.0 114655.0 ;
      RECT  99090.0 114250.0 99160.0 114655.0 ;
      RECT  99425.0 114250.0 99495.0 114655.0 ;
      RECT  99795.0 114250.0 99865.0 114655.0 ;
      RECT  100130.0 114250.0 100200.0 114655.0 ;
      RECT  100500.0 114250.0 100570.0 114655.0 ;
      RECT  100835.0 114250.0 100905.0 114655.0 ;
      RECT  101205.0 114250.0 101275.0 114655.0 ;
      RECT  101540.0 114250.0 101610.0 114655.0 ;
      RECT  101910.0 114250.0 101980.0 114655.0 ;
      RECT  102245.0 114250.0 102315.0 114655.0 ;
      RECT  102615.0 114250.0 102685.0 114655.0 ;
      RECT  102950.0 114250.0 103020.0 114655.0 ;
      RECT  103320.0 114250.0 103390.0 114655.0 ;
      RECT  103655.0 114250.0 103725.0 114655.0 ;
      RECT  104025.0 114250.0 104095.0 114655.0 ;
      RECT  104360.0 114250.0 104430.0 114655.0 ;
      RECT  104730.0 114250.0 104800.0 114655.0 ;
      RECT  105065.0 114250.0 105135.0 114655.0 ;
      RECT  105435.0 114250.0 105505.0 114655.0 ;
      RECT  105770.0 114250.0 105840.0 114655.0 ;
      RECT  16067.5 6520.0 16137.5 6590.0 ;
      RECT  15892.5 6520.0 16102.5 6590.0 ;
      RECT  16067.5 6555.0 16137.5 6695.0 ;
      RECT  18887.5 6520.0 18957.5 6590.0 ;
      RECT  18712.5 6520.0 18922.5 6590.0 ;
      RECT  18887.5 6555.0 18957.5 6695.0 ;
      RECT  21707.5 6520.0 21777.5 6590.0 ;
      RECT  21532.5 6520.0 21742.5 6590.0 ;
      RECT  21707.5 6555.0 21777.5 6695.0 ;
      RECT  24527.5 6520.0 24597.5 6590.0 ;
      RECT  24352.5 6520.0 24562.5 6590.0 ;
      RECT  24527.5 6555.0 24597.5 6695.0 ;
      RECT  27347.5 6520.0 27417.5 6590.0 ;
      RECT  27172.5 6520.0 27382.5 6590.0 ;
      RECT  27347.5 6555.0 27417.5 6695.0 ;
      RECT  30167.5 6520.0 30237.5 6590.0 ;
      RECT  29992.5 6520.0 30202.5 6590.0 ;
      RECT  30167.5 6555.0 30237.5 6695.0 ;
      RECT  32987.5 6520.0 33057.5 6590.0 ;
      RECT  32812.5 6520.0 33022.5 6590.0 ;
      RECT  32987.5 6555.0 33057.5 6695.0 ;
      RECT  35807.5 6520.0 35877.5 6590.0 ;
      RECT  35632.5 6520.0 35842.5 6590.0 ;
      RECT  35807.5 6555.0 35877.5 6695.0 ;
      RECT  38627.5 6520.0 38697.5 6590.0 ;
      RECT  38452.5 6520.0 38662.5 6590.0 ;
      RECT  38627.5 6555.0 38697.5 6695.0 ;
      RECT  41447.5 6520.0 41517.5 6590.0 ;
      RECT  41272.5 6520.0 41482.5 6590.0 ;
      RECT  41447.5 6555.0 41517.5 6695.0 ;
      RECT  44267.5 6520.0 44337.5 6590.0 ;
      RECT  44092.5 6520.0 44302.5 6590.0 ;
      RECT  44267.5 6555.0 44337.5 6695.0 ;
      RECT  47087.5 6520.0 47157.5 6590.0 ;
      RECT  46912.5 6520.0 47122.5 6590.0 ;
      RECT  47087.5 6555.0 47157.5 6695.0 ;
      RECT  49907.5 6520.0 49977.5 6590.0 ;
      RECT  49732.5 6520.0 49942.5 6590.0 ;
      RECT  49907.5 6555.0 49977.5 6695.0 ;
      RECT  52727.5 6520.0 52797.5 6590.0 ;
      RECT  52552.5 6520.0 52762.5 6590.0 ;
      RECT  52727.5 6555.0 52797.5 6695.0 ;
      RECT  55547.5 6520.0 55617.5 6590.0 ;
      RECT  55372.5 6520.0 55582.5 6590.0 ;
      RECT  55547.5 6555.0 55617.5 6695.0 ;
      RECT  58367.5 6520.0 58437.5 6590.0 ;
      RECT  58192.5 6520.0 58402.5 6590.0 ;
      RECT  58367.5 6555.0 58437.5 6695.0 ;
      RECT  61187.5 6520.0 61257.5 6590.0 ;
      RECT  61012.5 6520.0 61222.5 6590.0 ;
      RECT  61187.5 6555.0 61257.5 6695.0 ;
      RECT  64007.5 6520.0 64077.5 6590.0 ;
      RECT  63832.5 6520.0 64042.5 6590.0 ;
      RECT  64007.5 6555.0 64077.5 6695.0 ;
      RECT  66827.5 6520.0 66897.5 6590.0 ;
      RECT  66652.5 6520.0 66862.5 6590.0 ;
      RECT  66827.5 6555.0 66897.5 6695.0 ;
      RECT  69647.5 6520.0 69717.5 6590.0 ;
      RECT  69472.5 6520.0 69682.5 6590.0 ;
      RECT  69647.5 6555.0 69717.5 6695.0 ;
      RECT  72467.5 6520.0 72537.5 6590.0 ;
      RECT  72292.5 6520.0 72502.5 6590.0 ;
      RECT  72467.5 6555.0 72537.5 6695.0 ;
      RECT  75287.5 6520.0 75357.5 6590.0 ;
      RECT  75112.5 6520.0 75322.5 6590.0 ;
      RECT  75287.5 6555.0 75357.5 6695.0 ;
      RECT  78107.5 6520.0 78177.5 6590.0 ;
      RECT  77932.5 6520.0 78142.5 6590.0 ;
      RECT  78107.5 6555.0 78177.5 6695.0 ;
      RECT  80927.5 6520.0 80997.5 6590.0 ;
      RECT  80752.5 6520.0 80962.5 6590.0 ;
      RECT  80927.5 6555.0 80997.5 6695.0 ;
      RECT  83747.5 6520.0 83817.5 6590.0 ;
      RECT  83572.5 6520.0 83782.5 6590.0 ;
      RECT  83747.5 6555.0 83817.5 6695.0 ;
      RECT  86567.5 6520.0 86637.5 6590.0 ;
      RECT  86392.5 6520.0 86602.5 6590.0 ;
      RECT  86567.5 6555.0 86637.5 6695.0 ;
      RECT  89387.5 6520.0 89457.5 6590.0 ;
      RECT  89212.5 6520.0 89422.5 6590.0 ;
      RECT  89387.5 6555.0 89457.5 6695.0 ;
      RECT  92207.5 6520.0 92277.5 6590.0 ;
      RECT  92032.5 6520.0 92242.5 6590.0 ;
      RECT  92207.5 6555.0 92277.5 6695.0 ;
      RECT  95027.5 6520.0 95097.5 6590.0 ;
      RECT  94852.5 6520.0 95062.5 6590.0 ;
      RECT  95027.5 6555.0 95097.5 6695.0 ;
      RECT  97847.5 6520.0 97917.5 6590.0 ;
      RECT  97672.5 6520.0 97882.5 6590.0 ;
      RECT  97847.5 6555.0 97917.5 6695.0 ;
      RECT  100667.5 6520.0 100737.5 6590.0 ;
      RECT  100492.5 6520.0 100702.5 6590.0 ;
      RECT  100667.5 6555.0 100737.5 6695.0 ;
      RECT  103487.5 6520.0 103557.5 6590.0 ;
      RECT  103312.5 6520.0 103522.5 6590.0 ;
      RECT  103487.5 6555.0 103557.5 6695.0 ;
      RECT  8895.0 114095.0 8965.0 114300.0 ;
      RECT  15750.0 28015.0 16455.0 29360.0 ;
      RECT  15750.0 30705.0 16455.0 29360.0 ;
      RECT  15750.0 30705.0 16455.0 32050.0 ;
      RECT  15750.0 33395.0 16455.0 32050.0 ;
      RECT  15750.0 33395.0 16455.0 34740.0 ;
      RECT  15750.0 36085.0 16455.0 34740.0 ;
      RECT  15750.0 36085.0 16455.0 37430.0 ;
      RECT  15750.0 38775.0 16455.0 37430.0 ;
      RECT  15750.0 38775.0 16455.0 40120.0 ;
      RECT  15750.0 41465.0 16455.0 40120.0 ;
      RECT  15750.0 41465.0 16455.0 42810.0 ;
      RECT  15750.0 44155.0 16455.0 42810.0 ;
      RECT  15750.0 44155.0 16455.0 45500.0 ;
      RECT  15750.0 46845.0 16455.0 45500.0 ;
      RECT  15750.0 46845.0 16455.0 48190.0 ;
      RECT  15750.0 49535.0 16455.0 48190.0 ;
      RECT  15750.0 49535.0 16455.0 50880.0 ;
      RECT  15750.0 52225.0 16455.0 50880.0 ;
      RECT  15750.0 52225.0 16455.0 53570.0 ;
      RECT  15750.0 54915.0 16455.0 53570.0 ;
      RECT  15750.0 54915.0 16455.0 56260.0 ;
      RECT  15750.0 57605.0 16455.0 56260.0 ;
      RECT  15750.0 57605.0 16455.0 58950.0 ;
      RECT  15750.0 60295.0 16455.0 58950.0 ;
      RECT  15750.0 60295.0 16455.0 61640.0 ;
      RECT  15750.0 62985.0 16455.0 61640.0 ;
      RECT  15750.0 62985.0 16455.0 64330.0 ;
      RECT  15750.0 65675.0 16455.0 64330.0 ;
      RECT  15750.0 65675.0 16455.0 67020.0 ;
      RECT  15750.0 68365.0 16455.0 67020.0 ;
      RECT  15750.0 68365.0 16455.0 69710.0 ;
      RECT  15750.0 71055.0 16455.0 69710.0 ;
      RECT  15750.0 71055.0 16455.0 72400.0 ;
      RECT  15750.0 73745.0 16455.0 72400.0 ;
      RECT  15750.0 73745.0 16455.0 75090.0 ;
      RECT  15750.0 76435.0 16455.0 75090.0 ;
      RECT  15750.0 76435.0 16455.0 77780.0 ;
      RECT  15750.0 79125.0 16455.0 77780.0 ;
      RECT  15750.0 79125.0 16455.0 80470.0 ;
      RECT  15750.0 81815.0 16455.0 80470.0 ;
      RECT  15750.0 81815.0 16455.0 83160.0 ;
      RECT  15750.0 84505.0 16455.0 83160.0 ;
      RECT  15750.0 84505.0 16455.0 85850.0 ;
      RECT  15750.0 87195.0 16455.0 85850.0 ;
      RECT  15750.0 87195.0 16455.0 88540.0 ;
      RECT  15750.0 89885.0 16455.0 88540.0 ;
      RECT  15750.0 89885.0 16455.0 91230.0 ;
      RECT  15750.0 92575.0 16455.0 91230.0 ;
      RECT  15750.0 92575.0 16455.0 93920.0 ;
      RECT  15750.0 95265.0 16455.0 93920.0 ;
      RECT  15750.0 95265.0 16455.0 96610.0 ;
      RECT  15750.0 97955.0 16455.0 96610.0 ;
      RECT  15750.0 97955.0 16455.0 99300.0 ;
      RECT  15750.0 100645.0 16455.0 99300.0 ;
      RECT  15750.0 100645.0 16455.0 101990.0 ;
      RECT  15750.0 103335.0 16455.0 101990.0 ;
      RECT  15750.0 103335.0 16455.0 104680.0 ;
      RECT  15750.0 106025.0 16455.0 104680.0 ;
      RECT  15750.0 106025.0 16455.0 107370.0 ;
      RECT  15750.0 108715.0 16455.0 107370.0 ;
      RECT  15750.0 108715.0 16455.0 110060.0 ;
      RECT  15750.0 111405.0 16455.0 110060.0 ;
      RECT  15750.0 111405.0 16455.0 112750.0 ;
      RECT  15750.0 114095.0 16455.0 112750.0 ;
      RECT  16455.0 28015.0 17160.0 29360.0 ;
      RECT  16455.0 30705.0 17160.0 29360.0 ;
      RECT  16455.0 30705.0 17160.0 32050.0 ;
      RECT  16455.0 33395.0 17160.0 32050.0 ;
      RECT  16455.0 33395.0 17160.0 34740.0 ;
      RECT  16455.0 36085.0 17160.0 34740.0 ;
      RECT  16455.0 36085.0 17160.0 37430.0 ;
      RECT  16455.0 38775.0 17160.0 37430.0 ;
      RECT  16455.0 38775.0 17160.0 40120.0 ;
      RECT  16455.0 41465.0 17160.0 40120.0 ;
      RECT  16455.0 41465.0 17160.0 42810.0 ;
      RECT  16455.0 44155.0 17160.0 42810.0 ;
      RECT  16455.0 44155.0 17160.0 45500.0 ;
      RECT  16455.0 46845.0 17160.0 45500.0 ;
      RECT  16455.0 46845.0 17160.0 48190.0 ;
      RECT  16455.0 49535.0 17160.0 48190.0 ;
      RECT  16455.0 49535.0 17160.0 50880.0 ;
      RECT  16455.0 52225.0 17160.0 50880.0 ;
      RECT  16455.0 52225.0 17160.0 53570.0 ;
      RECT  16455.0 54915.0 17160.0 53570.0 ;
      RECT  16455.0 54915.0 17160.0 56260.0 ;
      RECT  16455.0 57605.0 17160.0 56260.0 ;
      RECT  16455.0 57605.0 17160.0 58950.0 ;
      RECT  16455.0 60295.0 17160.0 58950.0 ;
      RECT  16455.0 60295.0 17160.0 61640.0 ;
      RECT  16455.0 62985.0 17160.0 61640.0 ;
      RECT  16455.0 62985.0 17160.0 64330.0 ;
      RECT  16455.0 65675.0 17160.0 64330.0 ;
      RECT  16455.0 65675.0 17160.0 67020.0 ;
      RECT  16455.0 68365.0 17160.0 67020.0 ;
      RECT  16455.0 68365.0 17160.0 69710.0 ;
      RECT  16455.0 71055.0 17160.0 69710.0 ;
      RECT  16455.0 71055.0 17160.0 72400.0 ;
      RECT  16455.0 73745.0 17160.0 72400.0 ;
      RECT  16455.0 73745.0 17160.0 75090.0 ;
      RECT  16455.0 76435.0 17160.0 75090.0 ;
      RECT  16455.0 76435.0 17160.0 77780.0 ;
      RECT  16455.0 79125.0 17160.0 77780.0 ;
      RECT  16455.0 79125.0 17160.0 80470.0 ;
      RECT  16455.0 81815.0 17160.0 80470.0 ;
      RECT  16455.0 81815.0 17160.0 83160.0 ;
      RECT  16455.0 84505.0 17160.0 83160.0 ;
      RECT  16455.0 84505.0 17160.0 85850.0 ;
      RECT  16455.0 87195.0 17160.0 85850.0 ;
      RECT  16455.0 87195.0 17160.0 88540.0 ;
      RECT  16455.0 89885.0 17160.0 88540.0 ;
      RECT  16455.0 89885.0 17160.0 91230.0 ;
      RECT  16455.0 92575.0 17160.0 91230.0 ;
      RECT  16455.0 92575.0 17160.0 93920.0 ;
      RECT  16455.0 95265.0 17160.0 93920.0 ;
      RECT  16455.0 95265.0 17160.0 96610.0 ;
      RECT  16455.0 97955.0 17160.0 96610.0 ;
      RECT  16455.0 97955.0 17160.0 99300.0 ;
      RECT  16455.0 100645.0 17160.0 99300.0 ;
      RECT  16455.0 100645.0 17160.0 101990.0 ;
      RECT  16455.0 103335.0 17160.0 101990.0 ;
      RECT  16455.0 103335.0 17160.0 104680.0 ;
      RECT  16455.0 106025.0 17160.0 104680.0 ;
      RECT  16455.0 106025.0 17160.0 107370.0 ;
      RECT  16455.0 108715.0 17160.0 107370.0 ;
      RECT  16455.0 108715.0 17160.0 110060.0 ;
      RECT  16455.0 111405.0 17160.0 110060.0 ;
      RECT  16455.0 111405.0 17160.0 112750.0 ;
      RECT  16455.0 114095.0 17160.0 112750.0 ;
      RECT  17160.0 28015.0 17865.0 29360.0 ;
      RECT  17160.0 30705.0 17865.0 29360.0 ;
      RECT  17160.0 30705.0 17865.0 32050.0 ;
      RECT  17160.0 33395.0 17865.0 32050.0 ;
      RECT  17160.0 33395.0 17865.0 34740.0 ;
      RECT  17160.0 36085.0 17865.0 34740.0 ;
      RECT  17160.0 36085.0 17865.0 37430.0 ;
      RECT  17160.0 38775.0 17865.0 37430.0 ;
      RECT  17160.0 38775.0 17865.0 40120.0 ;
      RECT  17160.0 41465.0 17865.0 40120.0 ;
      RECT  17160.0 41465.0 17865.0 42810.0 ;
      RECT  17160.0 44155.0 17865.0 42810.0 ;
      RECT  17160.0 44155.0 17865.0 45500.0 ;
      RECT  17160.0 46845.0 17865.0 45500.0 ;
      RECT  17160.0 46845.0 17865.0 48190.0 ;
      RECT  17160.0 49535.0 17865.0 48190.0 ;
      RECT  17160.0 49535.0 17865.0 50880.0 ;
      RECT  17160.0 52225.0 17865.0 50880.0 ;
      RECT  17160.0 52225.0 17865.0 53570.0 ;
      RECT  17160.0 54915.0 17865.0 53570.0 ;
      RECT  17160.0 54915.0 17865.0 56260.0 ;
      RECT  17160.0 57605.0 17865.0 56260.0 ;
      RECT  17160.0 57605.0 17865.0 58950.0 ;
      RECT  17160.0 60295.0 17865.0 58950.0 ;
      RECT  17160.0 60295.0 17865.0 61640.0 ;
      RECT  17160.0 62985.0 17865.0 61640.0 ;
      RECT  17160.0 62985.0 17865.0 64330.0 ;
      RECT  17160.0 65675.0 17865.0 64330.0 ;
      RECT  17160.0 65675.0 17865.0 67020.0 ;
      RECT  17160.0 68365.0 17865.0 67020.0 ;
      RECT  17160.0 68365.0 17865.0 69710.0 ;
      RECT  17160.0 71055.0 17865.0 69710.0 ;
      RECT  17160.0 71055.0 17865.0 72400.0 ;
      RECT  17160.0 73745.0 17865.0 72400.0 ;
      RECT  17160.0 73745.0 17865.0 75090.0 ;
      RECT  17160.0 76435.0 17865.0 75090.0 ;
      RECT  17160.0 76435.0 17865.0 77780.0 ;
      RECT  17160.0 79125.0 17865.0 77780.0 ;
      RECT  17160.0 79125.0 17865.0 80470.0 ;
      RECT  17160.0 81815.0 17865.0 80470.0 ;
      RECT  17160.0 81815.0 17865.0 83160.0 ;
      RECT  17160.0 84505.0 17865.0 83160.0 ;
      RECT  17160.0 84505.0 17865.0 85850.0 ;
      RECT  17160.0 87195.0 17865.0 85850.0 ;
      RECT  17160.0 87195.0 17865.0 88540.0 ;
      RECT  17160.0 89885.0 17865.0 88540.0 ;
      RECT  17160.0 89885.0 17865.0 91230.0 ;
      RECT  17160.0 92575.0 17865.0 91230.0 ;
      RECT  17160.0 92575.0 17865.0 93920.0 ;
      RECT  17160.0 95265.0 17865.0 93920.0 ;
      RECT  17160.0 95265.0 17865.0 96610.0 ;
      RECT  17160.0 97955.0 17865.0 96610.0 ;
      RECT  17160.0 97955.0 17865.0 99300.0 ;
      RECT  17160.0 100645.0 17865.0 99300.0 ;
      RECT  17160.0 100645.0 17865.0 101990.0 ;
      RECT  17160.0 103335.0 17865.0 101990.0 ;
      RECT  17160.0 103335.0 17865.0 104680.0 ;
      RECT  17160.0 106025.0 17865.0 104680.0 ;
      RECT  17160.0 106025.0 17865.0 107370.0 ;
      RECT  17160.0 108715.0 17865.0 107370.0 ;
      RECT  17160.0 108715.0 17865.0 110060.0 ;
      RECT  17160.0 111405.0 17865.0 110060.0 ;
      RECT  17160.0 111405.0 17865.0 112750.0 ;
      RECT  17160.0 114095.0 17865.0 112750.0 ;
      RECT  17865.0 28015.0 18570.0 29360.0 ;
      RECT  17865.0 30705.0 18570.0 29360.0 ;
      RECT  17865.0 30705.0 18570.0 32050.0 ;
      RECT  17865.0 33395.0 18570.0 32050.0 ;
      RECT  17865.0 33395.0 18570.0 34740.0 ;
      RECT  17865.0 36085.0 18570.0 34740.0 ;
      RECT  17865.0 36085.0 18570.0 37430.0 ;
      RECT  17865.0 38775.0 18570.0 37430.0 ;
      RECT  17865.0 38775.0 18570.0 40120.0 ;
      RECT  17865.0 41465.0 18570.0 40120.0 ;
      RECT  17865.0 41465.0 18570.0 42810.0 ;
      RECT  17865.0 44155.0 18570.0 42810.0 ;
      RECT  17865.0 44155.0 18570.0 45500.0 ;
      RECT  17865.0 46845.0 18570.0 45500.0 ;
      RECT  17865.0 46845.0 18570.0 48190.0 ;
      RECT  17865.0 49535.0 18570.0 48190.0 ;
      RECT  17865.0 49535.0 18570.0 50880.0 ;
      RECT  17865.0 52225.0 18570.0 50880.0 ;
      RECT  17865.0 52225.0 18570.0 53570.0 ;
      RECT  17865.0 54915.0 18570.0 53570.0 ;
      RECT  17865.0 54915.0 18570.0 56260.0 ;
      RECT  17865.0 57605.0 18570.0 56260.0 ;
      RECT  17865.0 57605.0 18570.0 58950.0 ;
      RECT  17865.0 60295.0 18570.0 58950.0 ;
      RECT  17865.0 60295.0 18570.0 61640.0 ;
      RECT  17865.0 62985.0 18570.0 61640.0 ;
      RECT  17865.0 62985.0 18570.0 64330.0 ;
      RECT  17865.0 65675.0 18570.0 64330.0 ;
      RECT  17865.0 65675.0 18570.0 67020.0 ;
      RECT  17865.0 68365.0 18570.0 67020.0 ;
      RECT  17865.0 68365.0 18570.0 69710.0 ;
      RECT  17865.0 71055.0 18570.0 69710.0 ;
      RECT  17865.0 71055.0 18570.0 72400.0 ;
      RECT  17865.0 73745.0 18570.0 72400.0 ;
      RECT  17865.0 73745.0 18570.0 75090.0 ;
      RECT  17865.0 76435.0 18570.0 75090.0 ;
      RECT  17865.0 76435.0 18570.0 77780.0 ;
      RECT  17865.0 79125.0 18570.0 77780.0 ;
      RECT  17865.0 79125.0 18570.0 80470.0 ;
      RECT  17865.0 81815.0 18570.0 80470.0 ;
      RECT  17865.0 81815.0 18570.0 83160.0 ;
      RECT  17865.0 84505.0 18570.0 83160.0 ;
      RECT  17865.0 84505.0 18570.0 85850.0 ;
      RECT  17865.0 87195.0 18570.0 85850.0 ;
      RECT  17865.0 87195.0 18570.0 88540.0 ;
      RECT  17865.0 89885.0 18570.0 88540.0 ;
      RECT  17865.0 89885.0 18570.0 91230.0 ;
      RECT  17865.0 92575.0 18570.0 91230.0 ;
      RECT  17865.0 92575.0 18570.0 93920.0 ;
      RECT  17865.0 95265.0 18570.0 93920.0 ;
      RECT  17865.0 95265.0 18570.0 96610.0 ;
      RECT  17865.0 97955.0 18570.0 96610.0 ;
      RECT  17865.0 97955.0 18570.0 99300.0 ;
      RECT  17865.0 100645.0 18570.0 99300.0 ;
      RECT  17865.0 100645.0 18570.0 101990.0 ;
      RECT  17865.0 103335.0 18570.0 101990.0 ;
      RECT  17865.0 103335.0 18570.0 104680.0 ;
      RECT  17865.0 106025.0 18570.0 104680.0 ;
      RECT  17865.0 106025.0 18570.0 107370.0 ;
      RECT  17865.0 108715.0 18570.0 107370.0 ;
      RECT  17865.0 108715.0 18570.0 110060.0 ;
      RECT  17865.0 111405.0 18570.0 110060.0 ;
      RECT  17865.0 111405.0 18570.0 112750.0 ;
      RECT  17865.0 114095.0 18570.0 112750.0 ;
      RECT  18570.0 28015.0 19275.0 29360.0 ;
      RECT  18570.0 30705.0 19275.0 29360.0 ;
      RECT  18570.0 30705.0 19275.0 32050.0 ;
      RECT  18570.0 33395.0 19275.0 32050.0 ;
      RECT  18570.0 33395.0 19275.0 34740.0 ;
      RECT  18570.0 36085.0 19275.0 34740.0 ;
      RECT  18570.0 36085.0 19275.0 37430.0 ;
      RECT  18570.0 38775.0 19275.0 37430.0 ;
      RECT  18570.0 38775.0 19275.0 40120.0 ;
      RECT  18570.0 41465.0 19275.0 40120.0 ;
      RECT  18570.0 41465.0 19275.0 42810.0 ;
      RECT  18570.0 44155.0 19275.0 42810.0 ;
      RECT  18570.0 44155.0 19275.0 45500.0 ;
      RECT  18570.0 46845.0 19275.0 45500.0 ;
      RECT  18570.0 46845.0 19275.0 48190.0 ;
      RECT  18570.0 49535.0 19275.0 48190.0 ;
      RECT  18570.0 49535.0 19275.0 50880.0 ;
      RECT  18570.0 52225.0 19275.0 50880.0 ;
      RECT  18570.0 52225.0 19275.0 53570.0 ;
      RECT  18570.0 54915.0 19275.0 53570.0 ;
      RECT  18570.0 54915.0 19275.0 56260.0 ;
      RECT  18570.0 57605.0 19275.0 56260.0 ;
      RECT  18570.0 57605.0 19275.0 58950.0 ;
      RECT  18570.0 60295.0 19275.0 58950.0 ;
      RECT  18570.0 60295.0 19275.0 61640.0 ;
      RECT  18570.0 62985.0 19275.0 61640.0 ;
      RECT  18570.0 62985.0 19275.0 64330.0 ;
      RECT  18570.0 65675.0 19275.0 64330.0 ;
      RECT  18570.0 65675.0 19275.0 67020.0 ;
      RECT  18570.0 68365.0 19275.0 67020.0 ;
      RECT  18570.0 68365.0 19275.0 69710.0 ;
      RECT  18570.0 71055.0 19275.0 69710.0 ;
      RECT  18570.0 71055.0 19275.0 72400.0 ;
      RECT  18570.0 73745.0 19275.0 72400.0 ;
      RECT  18570.0 73745.0 19275.0 75090.0 ;
      RECT  18570.0 76435.0 19275.0 75090.0 ;
      RECT  18570.0 76435.0 19275.0 77780.0 ;
      RECT  18570.0 79125.0 19275.0 77780.0 ;
      RECT  18570.0 79125.0 19275.0 80470.0 ;
      RECT  18570.0 81815.0 19275.0 80470.0 ;
      RECT  18570.0 81815.0 19275.0 83160.0 ;
      RECT  18570.0 84505.0 19275.0 83160.0 ;
      RECT  18570.0 84505.0 19275.0 85850.0 ;
      RECT  18570.0 87195.0 19275.0 85850.0 ;
      RECT  18570.0 87195.0 19275.0 88540.0 ;
      RECT  18570.0 89885.0 19275.0 88540.0 ;
      RECT  18570.0 89885.0 19275.0 91230.0 ;
      RECT  18570.0 92575.0 19275.0 91230.0 ;
      RECT  18570.0 92575.0 19275.0 93920.0 ;
      RECT  18570.0 95265.0 19275.0 93920.0 ;
      RECT  18570.0 95265.0 19275.0 96610.0 ;
      RECT  18570.0 97955.0 19275.0 96610.0 ;
      RECT  18570.0 97955.0 19275.0 99300.0 ;
      RECT  18570.0 100645.0 19275.0 99300.0 ;
      RECT  18570.0 100645.0 19275.0 101990.0 ;
      RECT  18570.0 103335.0 19275.0 101990.0 ;
      RECT  18570.0 103335.0 19275.0 104680.0 ;
      RECT  18570.0 106025.0 19275.0 104680.0 ;
      RECT  18570.0 106025.0 19275.0 107370.0 ;
      RECT  18570.0 108715.0 19275.0 107370.0 ;
      RECT  18570.0 108715.0 19275.0 110060.0 ;
      RECT  18570.0 111405.0 19275.0 110060.0 ;
      RECT  18570.0 111405.0 19275.0 112750.0 ;
      RECT  18570.0 114095.0 19275.0 112750.0 ;
      RECT  19275.0 28015.0 19980.0 29360.0 ;
      RECT  19275.0 30705.0 19980.0 29360.0 ;
      RECT  19275.0 30705.0 19980.0 32050.0 ;
      RECT  19275.0 33395.0 19980.0 32050.0 ;
      RECT  19275.0 33395.0 19980.0 34740.0 ;
      RECT  19275.0 36085.0 19980.0 34740.0 ;
      RECT  19275.0 36085.0 19980.0 37430.0 ;
      RECT  19275.0 38775.0 19980.0 37430.0 ;
      RECT  19275.0 38775.0 19980.0 40120.0 ;
      RECT  19275.0 41465.0 19980.0 40120.0 ;
      RECT  19275.0 41465.0 19980.0 42810.0 ;
      RECT  19275.0 44155.0 19980.0 42810.0 ;
      RECT  19275.0 44155.0 19980.0 45500.0 ;
      RECT  19275.0 46845.0 19980.0 45500.0 ;
      RECT  19275.0 46845.0 19980.0 48190.0 ;
      RECT  19275.0 49535.0 19980.0 48190.0 ;
      RECT  19275.0 49535.0 19980.0 50880.0 ;
      RECT  19275.0 52225.0 19980.0 50880.0 ;
      RECT  19275.0 52225.0 19980.0 53570.0 ;
      RECT  19275.0 54915.0 19980.0 53570.0 ;
      RECT  19275.0 54915.0 19980.0 56260.0 ;
      RECT  19275.0 57605.0 19980.0 56260.0 ;
      RECT  19275.0 57605.0 19980.0 58950.0 ;
      RECT  19275.0 60295.0 19980.0 58950.0 ;
      RECT  19275.0 60295.0 19980.0 61640.0 ;
      RECT  19275.0 62985.0 19980.0 61640.0 ;
      RECT  19275.0 62985.0 19980.0 64330.0 ;
      RECT  19275.0 65675.0 19980.0 64330.0 ;
      RECT  19275.0 65675.0 19980.0 67020.0 ;
      RECT  19275.0 68365.0 19980.0 67020.0 ;
      RECT  19275.0 68365.0 19980.0 69710.0 ;
      RECT  19275.0 71055.0 19980.0 69710.0 ;
      RECT  19275.0 71055.0 19980.0 72400.0 ;
      RECT  19275.0 73745.0 19980.0 72400.0 ;
      RECT  19275.0 73745.0 19980.0 75090.0 ;
      RECT  19275.0 76435.0 19980.0 75090.0 ;
      RECT  19275.0 76435.0 19980.0 77780.0 ;
      RECT  19275.0 79125.0 19980.0 77780.0 ;
      RECT  19275.0 79125.0 19980.0 80470.0 ;
      RECT  19275.0 81815.0 19980.0 80470.0 ;
      RECT  19275.0 81815.0 19980.0 83160.0 ;
      RECT  19275.0 84505.0 19980.0 83160.0 ;
      RECT  19275.0 84505.0 19980.0 85850.0 ;
      RECT  19275.0 87195.0 19980.0 85850.0 ;
      RECT  19275.0 87195.0 19980.0 88540.0 ;
      RECT  19275.0 89885.0 19980.0 88540.0 ;
      RECT  19275.0 89885.0 19980.0 91230.0 ;
      RECT  19275.0 92575.0 19980.0 91230.0 ;
      RECT  19275.0 92575.0 19980.0 93920.0 ;
      RECT  19275.0 95265.0 19980.0 93920.0 ;
      RECT  19275.0 95265.0 19980.0 96610.0 ;
      RECT  19275.0 97955.0 19980.0 96610.0 ;
      RECT  19275.0 97955.0 19980.0 99300.0 ;
      RECT  19275.0 100645.0 19980.0 99300.0 ;
      RECT  19275.0 100645.0 19980.0 101990.0 ;
      RECT  19275.0 103335.0 19980.0 101990.0 ;
      RECT  19275.0 103335.0 19980.0 104680.0 ;
      RECT  19275.0 106025.0 19980.0 104680.0 ;
      RECT  19275.0 106025.0 19980.0 107370.0 ;
      RECT  19275.0 108715.0 19980.0 107370.0 ;
      RECT  19275.0 108715.0 19980.0 110060.0 ;
      RECT  19275.0 111405.0 19980.0 110060.0 ;
      RECT  19275.0 111405.0 19980.0 112750.0 ;
      RECT  19275.0 114095.0 19980.0 112750.0 ;
      RECT  19980.0 28015.0 20685.0 29360.0 ;
      RECT  19980.0 30705.0 20685.0 29360.0 ;
      RECT  19980.0 30705.0 20685.0 32050.0 ;
      RECT  19980.0 33395.0 20685.0 32050.0 ;
      RECT  19980.0 33395.0 20685.0 34740.0 ;
      RECT  19980.0 36085.0 20685.0 34740.0 ;
      RECT  19980.0 36085.0 20685.0 37430.0 ;
      RECT  19980.0 38775.0 20685.0 37430.0 ;
      RECT  19980.0 38775.0 20685.0 40120.0 ;
      RECT  19980.0 41465.0 20685.0 40120.0 ;
      RECT  19980.0 41465.0 20685.0 42810.0 ;
      RECT  19980.0 44155.0 20685.0 42810.0 ;
      RECT  19980.0 44155.0 20685.0 45500.0 ;
      RECT  19980.0 46845.0 20685.0 45500.0 ;
      RECT  19980.0 46845.0 20685.0 48190.0 ;
      RECT  19980.0 49535.0 20685.0 48190.0 ;
      RECT  19980.0 49535.0 20685.0 50880.0 ;
      RECT  19980.0 52225.0 20685.0 50880.0 ;
      RECT  19980.0 52225.0 20685.0 53570.0 ;
      RECT  19980.0 54915.0 20685.0 53570.0 ;
      RECT  19980.0 54915.0 20685.0 56260.0 ;
      RECT  19980.0 57605.0 20685.0 56260.0 ;
      RECT  19980.0 57605.0 20685.0 58950.0 ;
      RECT  19980.0 60295.0 20685.0 58950.0 ;
      RECT  19980.0 60295.0 20685.0 61640.0 ;
      RECT  19980.0 62985.0 20685.0 61640.0 ;
      RECT  19980.0 62985.0 20685.0 64330.0 ;
      RECT  19980.0 65675.0 20685.0 64330.0 ;
      RECT  19980.0 65675.0 20685.0 67020.0 ;
      RECT  19980.0 68365.0 20685.0 67020.0 ;
      RECT  19980.0 68365.0 20685.0 69710.0 ;
      RECT  19980.0 71055.0 20685.0 69710.0 ;
      RECT  19980.0 71055.0 20685.0 72400.0 ;
      RECT  19980.0 73745.0 20685.0 72400.0 ;
      RECT  19980.0 73745.0 20685.0 75090.0 ;
      RECT  19980.0 76435.0 20685.0 75090.0 ;
      RECT  19980.0 76435.0 20685.0 77780.0 ;
      RECT  19980.0 79125.0 20685.0 77780.0 ;
      RECT  19980.0 79125.0 20685.0 80470.0 ;
      RECT  19980.0 81815.0 20685.0 80470.0 ;
      RECT  19980.0 81815.0 20685.0 83160.0 ;
      RECT  19980.0 84505.0 20685.0 83160.0 ;
      RECT  19980.0 84505.0 20685.0 85850.0 ;
      RECT  19980.0 87195.0 20685.0 85850.0 ;
      RECT  19980.0 87195.0 20685.0 88540.0 ;
      RECT  19980.0 89885.0 20685.0 88540.0 ;
      RECT  19980.0 89885.0 20685.0 91230.0 ;
      RECT  19980.0 92575.0 20685.0 91230.0 ;
      RECT  19980.0 92575.0 20685.0 93920.0 ;
      RECT  19980.0 95265.0 20685.0 93920.0 ;
      RECT  19980.0 95265.0 20685.0 96610.0 ;
      RECT  19980.0 97955.0 20685.0 96610.0 ;
      RECT  19980.0 97955.0 20685.0 99300.0 ;
      RECT  19980.0 100645.0 20685.0 99300.0 ;
      RECT  19980.0 100645.0 20685.0 101990.0 ;
      RECT  19980.0 103335.0 20685.0 101990.0 ;
      RECT  19980.0 103335.0 20685.0 104680.0 ;
      RECT  19980.0 106025.0 20685.0 104680.0 ;
      RECT  19980.0 106025.0 20685.0 107370.0 ;
      RECT  19980.0 108715.0 20685.0 107370.0 ;
      RECT  19980.0 108715.0 20685.0 110060.0 ;
      RECT  19980.0 111405.0 20685.0 110060.0 ;
      RECT  19980.0 111405.0 20685.0 112750.0 ;
      RECT  19980.0 114095.0 20685.0 112750.0 ;
      RECT  20685.0 28015.0 21390.0 29360.0 ;
      RECT  20685.0 30705.0 21390.0 29360.0 ;
      RECT  20685.0 30705.0 21390.0 32050.0 ;
      RECT  20685.0 33395.0 21390.0 32050.0 ;
      RECT  20685.0 33395.0 21390.0 34740.0 ;
      RECT  20685.0 36085.0 21390.0 34740.0 ;
      RECT  20685.0 36085.0 21390.0 37430.0 ;
      RECT  20685.0 38775.0 21390.0 37430.0 ;
      RECT  20685.0 38775.0 21390.0 40120.0 ;
      RECT  20685.0 41465.0 21390.0 40120.0 ;
      RECT  20685.0 41465.0 21390.0 42810.0 ;
      RECT  20685.0 44155.0 21390.0 42810.0 ;
      RECT  20685.0 44155.0 21390.0 45500.0 ;
      RECT  20685.0 46845.0 21390.0 45500.0 ;
      RECT  20685.0 46845.0 21390.0 48190.0 ;
      RECT  20685.0 49535.0 21390.0 48190.0 ;
      RECT  20685.0 49535.0 21390.0 50880.0 ;
      RECT  20685.0 52225.0 21390.0 50880.0 ;
      RECT  20685.0 52225.0 21390.0 53570.0 ;
      RECT  20685.0 54915.0 21390.0 53570.0 ;
      RECT  20685.0 54915.0 21390.0 56260.0 ;
      RECT  20685.0 57605.0 21390.0 56260.0 ;
      RECT  20685.0 57605.0 21390.0 58950.0 ;
      RECT  20685.0 60295.0 21390.0 58950.0 ;
      RECT  20685.0 60295.0 21390.0 61640.0 ;
      RECT  20685.0 62985.0 21390.0 61640.0 ;
      RECT  20685.0 62985.0 21390.0 64330.0 ;
      RECT  20685.0 65675.0 21390.0 64330.0 ;
      RECT  20685.0 65675.0 21390.0 67020.0 ;
      RECT  20685.0 68365.0 21390.0 67020.0 ;
      RECT  20685.0 68365.0 21390.0 69710.0 ;
      RECT  20685.0 71055.0 21390.0 69710.0 ;
      RECT  20685.0 71055.0 21390.0 72400.0 ;
      RECT  20685.0 73745.0 21390.0 72400.0 ;
      RECT  20685.0 73745.0 21390.0 75090.0 ;
      RECT  20685.0 76435.0 21390.0 75090.0 ;
      RECT  20685.0 76435.0 21390.0 77780.0 ;
      RECT  20685.0 79125.0 21390.0 77780.0 ;
      RECT  20685.0 79125.0 21390.0 80470.0 ;
      RECT  20685.0 81815.0 21390.0 80470.0 ;
      RECT  20685.0 81815.0 21390.0 83160.0 ;
      RECT  20685.0 84505.0 21390.0 83160.0 ;
      RECT  20685.0 84505.0 21390.0 85850.0 ;
      RECT  20685.0 87195.0 21390.0 85850.0 ;
      RECT  20685.0 87195.0 21390.0 88540.0 ;
      RECT  20685.0 89885.0 21390.0 88540.0 ;
      RECT  20685.0 89885.0 21390.0 91230.0 ;
      RECT  20685.0 92575.0 21390.0 91230.0 ;
      RECT  20685.0 92575.0 21390.0 93920.0 ;
      RECT  20685.0 95265.0 21390.0 93920.0 ;
      RECT  20685.0 95265.0 21390.0 96610.0 ;
      RECT  20685.0 97955.0 21390.0 96610.0 ;
      RECT  20685.0 97955.0 21390.0 99300.0 ;
      RECT  20685.0 100645.0 21390.0 99300.0 ;
      RECT  20685.0 100645.0 21390.0 101990.0 ;
      RECT  20685.0 103335.0 21390.0 101990.0 ;
      RECT  20685.0 103335.0 21390.0 104680.0 ;
      RECT  20685.0 106025.0 21390.0 104680.0 ;
      RECT  20685.0 106025.0 21390.0 107370.0 ;
      RECT  20685.0 108715.0 21390.0 107370.0 ;
      RECT  20685.0 108715.0 21390.0 110060.0 ;
      RECT  20685.0 111405.0 21390.0 110060.0 ;
      RECT  20685.0 111405.0 21390.0 112750.0 ;
      RECT  20685.0 114095.0 21390.0 112750.0 ;
      RECT  21390.0 28015.0 22095.0 29360.0 ;
      RECT  21390.0 30705.0 22095.0 29360.0 ;
      RECT  21390.0 30705.0 22095.0 32050.0 ;
      RECT  21390.0 33395.0 22095.0 32050.0 ;
      RECT  21390.0 33395.0 22095.0 34740.0 ;
      RECT  21390.0 36085.0 22095.0 34740.0 ;
      RECT  21390.0 36085.0 22095.0 37430.0 ;
      RECT  21390.0 38775.0 22095.0 37430.0 ;
      RECT  21390.0 38775.0 22095.0 40120.0 ;
      RECT  21390.0 41465.0 22095.0 40120.0 ;
      RECT  21390.0 41465.0 22095.0 42810.0 ;
      RECT  21390.0 44155.0 22095.0 42810.0 ;
      RECT  21390.0 44155.0 22095.0 45500.0 ;
      RECT  21390.0 46845.0 22095.0 45500.0 ;
      RECT  21390.0 46845.0 22095.0 48190.0 ;
      RECT  21390.0 49535.0 22095.0 48190.0 ;
      RECT  21390.0 49535.0 22095.0 50880.0 ;
      RECT  21390.0 52225.0 22095.0 50880.0 ;
      RECT  21390.0 52225.0 22095.0 53570.0 ;
      RECT  21390.0 54915.0 22095.0 53570.0 ;
      RECT  21390.0 54915.0 22095.0 56260.0 ;
      RECT  21390.0 57605.0 22095.0 56260.0 ;
      RECT  21390.0 57605.0 22095.0 58950.0 ;
      RECT  21390.0 60295.0 22095.0 58950.0 ;
      RECT  21390.0 60295.0 22095.0 61640.0 ;
      RECT  21390.0 62985.0 22095.0 61640.0 ;
      RECT  21390.0 62985.0 22095.0 64330.0 ;
      RECT  21390.0 65675.0 22095.0 64330.0 ;
      RECT  21390.0 65675.0 22095.0 67020.0 ;
      RECT  21390.0 68365.0 22095.0 67020.0 ;
      RECT  21390.0 68365.0 22095.0 69710.0 ;
      RECT  21390.0 71055.0 22095.0 69710.0 ;
      RECT  21390.0 71055.0 22095.0 72400.0 ;
      RECT  21390.0 73745.0 22095.0 72400.0 ;
      RECT  21390.0 73745.0 22095.0 75090.0 ;
      RECT  21390.0 76435.0 22095.0 75090.0 ;
      RECT  21390.0 76435.0 22095.0 77780.0 ;
      RECT  21390.0 79125.0 22095.0 77780.0 ;
      RECT  21390.0 79125.0 22095.0 80470.0 ;
      RECT  21390.0 81815.0 22095.0 80470.0 ;
      RECT  21390.0 81815.0 22095.0 83160.0 ;
      RECT  21390.0 84505.0 22095.0 83160.0 ;
      RECT  21390.0 84505.0 22095.0 85850.0 ;
      RECT  21390.0 87195.0 22095.0 85850.0 ;
      RECT  21390.0 87195.0 22095.0 88540.0 ;
      RECT  21390.0 89885.0 22095.0 88540.0 ;
      RECT  21390.0 89885.0 22095.0 91230.0 ;
      RECT  21390.0 92575.0 22095.0 91230.0 ;
      RECT  21390.0 92575.0 22095.0 93920.0 ;
      RECT  21390.0 95265.0 22095.0 93920.0 ;
      RECT  21390.0 95265.0 22095.0 96610.0 ;
      RECT  21390.0 97955.0 22095.0 96610.0 ;
      RECT  21390.0 97955.0 22095.0 99300.0 ;
      RECT  21390.0 100645.0 22095.0 99300.0 ;
      RECT  21390.0 100645.0 22095.0 101990.0 ;
      RECT  21390.0 103335.0 22095.0 101990.0 ;
      RECT  21390.0 103335.0 22095.0 104680.0 ;
      RECT  21390.0 106025.0 22095.0 104680.0 ;
      RECT  21390.0 106025.0 22095.0 107370.0 ;
      RECT  21390.0 108715.0 22095.0 107370.0 ;
      RECT  21390.0 108715.0 22095.0 110060.0 ;
      RECT  21390.0 111405.0 22095.0 110060.0 ;
      RECT  21390.0 111405.0 22095.0 112750.0 ;
      RECT  21390.0 114095.0 22095.0 112750.0 ;
      RECT  22095.0 28015.0 22800.0 29360.0 ;
      RECT  22095.0 30705.0 22800.0 29360.0 ;
      RECT  22095.0 30705.0 22800.0 32050.0 ;
      RECT  22095.0 33395.0 22800.0 32050.0 ;
      RECT  22095.0 33395.0 22800.0 34740.0 ;
      RECT  22095.0 36085.0 22800.0 34740.0 ;
      RECT  22095.0 36085.0 22800.0 37430.0 ;
      RECT  22095.0 38775.0 22800.0 37430.0 ;
      RECT  22095.0 38775.0 22800.0 40120.0 ;
      RECT  22095.0 41465.0 22800.0 40120.0 ;
      RECT  22095.0 41465.0 22800.0 42810.0 ;
      RECT  22095.0 44155.0 22800.0 42810.0 ;
      RECT  22095.0 44155.0 22800.0 45500.0 ;
      RECT  22095.0 46845.0 22800.0 45500.0 ;
      RECT  22095.0 46845.0 22800.0 48190.0 ;
      RECT  22095.0 49535.0 22800.0 48190.0 ;
      RECT  22095.0 49535.0 22800.0 50880.0 ;
      RECT  22095.0 52225.0 22800.0 50880.0 ;
      RECT  22095.0 52225.0 22800.0 53570.0 ;
      RECT  22095.0 54915.0 22800.0 53570.0 ;
      RECT  22095.0 54915.0 22800.0 56260.0 ;
      RECT  22095.0 57605.0 22800.0 56260.0 ;
      RECT  22095.0 57605.0 22800.0 58950.0 ;
      RECT  22095.0 60295.0 22800.0 58950.0 ;
      RECT  22095.0 60295.0 22800.0 61640.0 ;
      RECT  22095.0 62985.0 22800.0 61640.0 ;
      RECT  22095.0 62985.0 22800.0 64330.0 ;
      RECT  22095.0 65675.0 22800.0 64330.0 ;
      RECT  22095.0 65675.0 22800.0 67020.0 ;
      RECT  22095.0 68365.0 22800.0 67020.0 ;
      RECT  22095.0 68365.0 22800.0 69710.0 ;
      RECT  22095.0 71055.0 22800.0 69710.0 ;
      RECT  22095.0 71055.0 22800.0 72400.0 ;
      RECT  22095.0 73745.0 22800.0 72400.0 ;
      RECT  22095.0 73745.0 22800.0 75090.0 ;
      RECT  22095.0 76435.0 22800.0 75090.0 ;
      RECT  22095.0 76435.0 22800.0 77780.0 ;
      RECT  22095.0 79125.0 22800.0 77780.0 ;
      RECT  22095.0 79125.0 22800.0 80470.0 ;
      RECT  22095.0 81815.0 22800.0 80470.0 ;
      RECT  22095.0 81815.0 22800.0 83160.0 ;
      RECT  22095.0 84505.0 22800.0 83160.0 ;
      RECT  22095.0 84505.0 22800.0 85850.0 ;
      RECT  22095.0 87195.0 22800.0 85850.0 ;
      RECT  22095.0 87195.0 22800.0 88540.0 ;
      RECT  22095.0 89885.0 22800.0 88540.0 ;
      RECT  22095.0 89885.0 22800.0 91230.0 ;
      RECT  22095.0 92575.0 22800.0 91230.0 ;
      RECT  22095.0 92575.0 22800.0 93920.0 ;
      RECT  22095.0 95265.0 22800.0 93920.0 ;
      RECT  22095.0 95265.0 22800.0 96610.0 ;
      RECT  22095.0 97955.0 22800.0 96610.0 ;
      RECT  22095.0 97955.0 22800.0 99300.0 ;
      RECT  22095.0 100645.0 22800.0 99300.0 ;
      RECT  22095.0 100645.0 22800.0 101990.0 ;
      RECT  22095.0 103335.0 22800.0 101990.0 ;
      RECT  22095.0 103335.0 22800.0 104680.0 ;
      RECT  22095.0 106025.0 22800.0 104680.0 ;
      RECT  22095.0 106025.0 22800.0 107370.0 ;
      RECT  22095.0 108715.0 22800.0 107370.0 ;
      RECT  22095.0 108715.0 22800.0 110060.0 ;
      RECT  22095.0 111405.0 22800.0 110060.0 ;
      RECT  22095.0 111405.0 22800.0 112750.0 ;
      RECT  22095.0 114095.0 22800.0 112750.0 ;
      RECT  22800.0 28015.0 23505.0 29360.0 ;
      RECT  22800.0 30705.0 23505.0 29360.0 ;
      RECT  22800.0 30705.0 23505.0 32050.0 ;
      RECT  22800.0 33395.0 23505.0 32050.0 ;
      RECT  22800.0 33395.0 23505.0 34740.0 ;
      RECT  22800.0 36085.0 23505.0 34740.0 ;
      RECT  22800.0 36085.0 23505.0 37430.0 ;
      RECT  22800.0 38775.0 23505.0 37430.0 ;
      RECT  22800.0 38775.0 23505.0 40120.0 ;
      RECT  22800.0 41465.0 23505.0 40120.0 ;
      RECT  22800.0 41465.0 23505.0 42810.0 ;
      RECT  22800.0 44155.0 23505.0 42810.0 ;
      RECT  22800.0 44155.0 23505.0 45500.0 ;
      RECT  22800.0 46845.0 23505.0 45500.0 ;
      RECT  22800.0 46845.0 23505.0 48190.0 ;
      RECT  22800.0 49535.0 23505.0 48190.0 ;
      RECT  22800.0 49535.0 23505.0 50880.0 ;
      RECT  22800.0 52225.0 23505.0 50880.0 ;
      RECT  22800.0 52225.0 23505.0 53570.0 ;
      RECT  22800.0 54915.0 23505.0 53570.0 ;
      RECT  22800.0 54915.0 23505.0 56260.0 ;
      RECT  22800.0 57605.0 23505.0 56260.0 ;
      RECT  22800.0 57605.0 23505.0 58950.0 ;
      RECT  22800.0 60295.0 23505.0 58950.0 ;
      RECT  22800.0 60295.0 23505.0 61640.0 ;
      RECT  22800.0 62985.0 23505.0 61640.0 ;
      RECT  22800.0 62985.0 23505.0 64330.0 ;
      RECT  22800.0 65675.0 23505.0 64330.0 ;
      RECT  22800.0 65675.0 23505.0 67020.0 ;
      RECT  22800.0 68365.0 23505.0 67020.0 ;
      RECT  22800.0 68365.0 23505.0 69710.0 ;
      RECT  22800.0 71055.0 23505.0 69710.0 ;
      RECT  22800.0 71055.0 23505.0 72400.0 ;
      RECT  22800.0 73745.0 23505.0 72400.0 ;
      RECT  22800.0 73745.0 23505.0 75090.0 ;
      RECT  22800.0 76435.0 23505.0 75090.0 ;
      RECT  22800.0 76435.0 23505.0 77780.0 ;
      RECT  22800.0 79125.0 23505.0 77780.0 ;
      RECT  22800.0 79125.0 23505.0 80470.0 ;
      RECT  22800.0 81815.0 23505.0 80470.0 ;
      RECT  22800.0 81815.0 23505.0 83160.0 ;
      RECT  22800.0 84505.0 23505.0 83160.0 ;
      RECT  22800.0 84505.0 23505.0 85850.0 ;
      RECT  22800.0 87195.0 23505.0 85850.0 ;
      RECT  22800.0 87195.0 23505.0 88540.0 ;
      RECT  22800.0 89885.0 23505.0 88540.0 ;
      RECT  22800.0 89885.0 23505.0 91230.0 ;
      RECT  22800.0 92575.0 23505.0 91230.0 ;
      RECT  22800.0 92575.0 23505.0 93920.0 ;
      RECT  22800.0 95265.0 23505.0 93920.0 ;
      RECT  22800.0 95265.0 23505.0 96610.0 ;
      RECT  22800.0 97955.0 23505.0 96610.0 ;
      RECT  22800.0 97955.0 23505.0 99300.0 ;
      RECT  22800.0 100645.0 23505.0 99300.0 ;
      RECT  22800.0 100645.0 23505.0 101990.0 ;
      RECT  22800.0 103335.0 23505.0 101990.0 ;
      RECT  22800.0 103335.0 23505.0 104680.0 ;
      RECT  22800.0 106025.0 23505.0 104680.0 ;
      RECT  22800.0 106025.0 23505.0 107370.0 ;
      RECT  22800.0 108715.0 23505.0 107370.0 ;
      RECT  22800.0 108715.0 23505.0 110060.0 ;
      RECT  22800.0 111405.0 23505.0 110060.0 ;
      RECT  22800.0 111405.0 23505.0 112750.0 ;
      RECT  22800.0 114095.0 23505.0 112750.0 ;
      RECT  23505.0 28015.0 24210.0 29360.0 ;
      RECT  23505.0 30705.0 24210.0 29360.0 ;
      RECT  23505.0 30705.0 24210.0 32050.0 ;
      RECT  23505.0 33395.0 24210.0 32050.0 ;
      RECT  23505.0 33395.0 24210.0 34740.0 ;
      RECT  23505.0 36085.0 24210.0 34740.0 ;
      RECT  23505.0 36085.0 24210.0 37430.0 ;
      RECT  23505.0 38775.0 24210.0 37430.0 ;
      RECT  23505.0 38775.0 24210.0 40120.0 ;
      RECT  23505.0 41465.0 24210.0 40120.0 ;
      RECT  23505.0 41465.0 24210.0 42810.0 ;
      RECT  23505.0 44155.0 24210.0 42810.0 ;
      RECT  23505.0 44155.0 24210.0 45500.0 ;
      RECT  23505.0 46845.0 24210.0 45500.0 ;
      RECT  23505.0 46845.0 24210.0 48190.0 ;
      RECT  23505.0 49535.0 24210.0 48190.0 ;
      RECT  23505.0 49535.0 24210.0 50880.0 ;
      RECT  23505.0 52225.0 24210.0 50880.0 ;
      RECT  23505.0 52225.0 24210.0 53570.0 ;
      RECT  23505.0 54915.0 24210.0 53570.0 ;
      RECT  23505.0 54915.0 24210.0 56260.0 ;
      RECT  23505.0 57605.0 24210.0 56260.0 ;
      RECT  23505.0 57605.0 24210.0 58950.0 ;
      RECT  23505.0 60295.0 24210.0 58950.0 ;
      RECT  23505.0 60295.0 24210.0 61640.0 ;
      RECT  23505.0 62985.0 24210.0 61640.0 ;
      RECT  23505.0 62985.0 24210.0 64330.0 ;
      RECT  23505.0 65675.0 24210.0 64330.0 ;
      RECT  23505.0 65675.0 24210.0 67020.0 ;
      RECT  23505.0 68365.0 24210.0 67020.0 ;
      RECT  23505.0 68365.0 24210.0 69710.0 ;
      RECT  23505.0 71055.0 24210.0 69710.0 ;
      RECT  23505.0 71055.0 24210.0 72400.0 ;
      RECT  23505.0 73745.0 24210.0 72400.0 ;
      RECT  23505.0 73745.0 24210.0 75090.0 ;
      RECT  23505.0 76435.0 24210.0 75090.0 ;
      RECT  23505.0 76435.0 24210.0 77780.0 ;
      RECT  23505.0 79125.0 24210.0 77780.0 ;
      RECT  23505.0 79125.0 24210.0 80470.0 ;
      RECT  23505.0 81815.0 24210.0 80470.0 ;
      RECT  23505.0 81815.0 24210.0 83160.0 ;
      RECT  23505.0 84505.0 24210.0 83160.0 ;
      RECT  23505.0 84505.0 24210.0 85850.0 ;
      RECT  23505.0 87195.0 24210.0 85850.0 ;
      RECT  23505.0 87195.0 24210.0 88540.0 ;
      RECT  23505.0 89885.0 24210.0 88540.0 ;
      RECT  23505.0 89885.0 24210.0 91230.0 ;
      RECT  23505.0 92575.0 24210.0 91230.0 ;
      RECT  23505.0 92575.0 24210.0 93920.0 ;
      RECT  23505.0 95265.0 24210.0 93920.0 ;
      RECT  23505.0 95265.0 24210.0 96610.0 ;
      RECT  23505.0 97955.0 24210.0 96610.0 ;
      RECT  23505.0 97955.0 24210.0 99300.0 ;
      RECT  23505.0 100645.0 24210.0 99300.0 ;
      RECT  23505.0 100645.0 24210.0 101990.0 ;
      RECT  23505.0 103335.0 24210.0 101990.0 ;
      RECT  23505.0 103335.0 24210.0 104680.0 ;
      RECT  23505.0 106025.0 24210.0 104680.0 ;
      RECT  23505.0 106025.0 24210.0 107370.0 ;
      RECT  23505.0 108715.0 24210.0 107370.0 ;
      RECT  23505.0 108715.0 24210.0 110060.0 ;
      RECT  23505.0 111405.0 24210.0 110060.0 ;
      RECT  23505.0 111405.0 24210.0 112750.0 ;
      RECT  23505.0 114095.0 24210.0 112750.0 ;
      RECT  24210.0 28015.0 24915.0 29360.0 ;
      RECT  24210.0 30705.0 24915.0 29360.0 ;
      RECT  24210.0 30705.0 24915.0 32050.0 ;
      RECT  24210.0 33395.0 24915.0 32050.0 ;
      RECT  24210.0 33395.0 24915.0 34740.0 ;
      RECT  24210.0 36085.0 24915.0 34740.0 ;
      RECT  24210.0 36085.0 24915.0 37430.0 ;
      RECT  24210.0 38775.0 24915.0 37430.0 ;
      RECT  24210.0 38775.0 24915.0 40120.0 ;
      RECT  24210.0 41465.0 24915.0 40120.0 ;
      RECT  24210.0 41465.0 24915.0 42810.0 ;
      RECT  24210.0 44155.0 24915.0 42810.0 ;
      RECT  24210.0 44155.0 24915.0 45500.0 ;
      RECT  24210.0 46845.0 24915.0 45500.0 ;
      RECT  24210.0 46845.0 24915.0 48190.0 ;
      RECT  24210.0 49535.0 24915.0 48190.0 ;
      RECT  24210.0 49535.0 24915.0 50880.0 ;
      RECT  24210.0 52225.0 24915.0 50880.0 ;
      RECT  24210.0 52225.0 24915.0 53570.0 ;
      RECT  24210.0 54915.0 24915.0 53570.0 ;
      RECT  24210.0 54915.0 24915.0 56260.0 ;
      RECT  24210.0 57605.0 24915.0 56260.0 ;
      RECT  24210.0 57605.0 24915.0 58950.0 ;
      RECT  24210.0 60295.0 24915.0 58950.0 ;
      RECT  24210.0 60295.0 24915.0 61640.0 ;
      RECT  24210.0 62985.0 24915.0 61640.0 ;
      RECT  24210.0 62985.0 24915.0 64330.0 ;
      RECT  24210.0 65675.0 24915.0 64330.0 ;
      RECT  24210.0 65675.0 24915.0 67020.0 ;
      RECT  24210.0 68365.0 24915.0 67020.0 ;
      RECT  24210.0 68365.0 24915.0 69710.0 ;
      RECT  24210.0 71055.0 24915.0 69710.0 ;
      RECT  24210.0 71055.0 24915.0 72400.0 ;
      RECT  24210.0 73745.0 24915.0 72400.0 ;
      RECT  24210.0 73745.0 24915.0 75090.0 ;
      RECT  24210.0 76435.0 24915.0 75090.0 ;
      RECT  24210.0 76435.0 24915.0 77780.0 ;
      RECT  24210.0 79125.0 24915.0 77780.0 ;
      RECT  24210.0 79125.0 24915.0 80470.0 ;
      RECT  24210.0 81815.0 24915.0 80470.0 ;
      RECT  24210.0 81815.0 24915.0 83160.0 ;
      RECT  24210.0 84505.0 24915.0 83160.0 ;
      RECT  24210.0 84505.0 24915.0 85850.0 ;
      RECT  24210.0 87195.0 24915.0 85850.0 ;
      RECT  24210.0 87195.0 24915.0 88540.0 ;
      RECT  24210.0 89885.0 24915.0 88540.0 ;
      RECT  24210.0 89885.0 24915.0 91230.0 ;
      RECT  24210.0 92575.0 24915.0 91230.0 ;
      RECT  24210.0 92575.0 24915.0 93920.0 ;
      RECT  24210.0 95265.0 24915.0 93920.0 ;
      RECT  24210.0 95265.0 24915.0 96610.0 ;
      RECT  24210.0 97955.0 24915.0 96610.0 ;
      RECT  24210.0 97955.0 24915.0 99300.0 ;
      RECT  24210.0 100645.0 24915.0 99300.0 ;
      RECT  24210.0 100645.0 24915.0 101990.0 ;
      RECT  24210.0 103335.0 24915.0 101990.0 ;
      RECT  24210.0 103335.0 24915.0 104680.0 ;
      RECT  24210.0 106025.0 24915.0 104680.0 ;
      RECT  24210.0 106025.0 24915.0 107370.0 ;
      RECT  24210.0 108715.0 24915.0 107370.0 ;
      RECT  24210.0 108715.0 24915.0 110060.0 ;
      RECT  24210.0 111405.0 24915.0 110060.0 ;
      RECT  24210.0 111405.0 24915.0 112750.0 ;
      RECT  24210.0 114095.0 24915.0 112750.0 ;
      RECT  24915.0 28015.0 25620.0 29360.0 ;
      RECT  24915.0 30705.0 25620.0 29360.0 ;
      RECT  24915.0 30705.0 25620.0 32050.0 ;
      RECT  24915.0 33395.0 25620.0 32050.0 ;
      RECT  24915.0 33395.0 25620.0 34740.0 ;
      RECT  24915.0 36085.0 25620.0 34740.0 ;
      RECT  24915.0 36085.0 25620.0 37430.0 ;
      RECT  24915.0 38775.0 25620.0 37430.0 ;
      RECT  24915.0 38775.0 25620.0 40120.0 ;
      RECT  24915.0 41465.0 25620.0 40120.0 ;
      RECT  24915.0 41465.0 25620.0 42810.0 ;
      RECT  24915.0 44155.0 25620.0 42810.0 ;
      RECT  24915.0 44155.0 25620.0 45500.0 ;
      RECT  24915.0 46845.0 25620.0 45500.0 ;
      RECT  24915.0 46845.0 25620.0 48190.0 ;
      RECT  24915.0 49535.0 25620.0 48190.0 ;
      RECT  24915.0 49535.0 25620.0 50880.0 ;
      RECT  24915.0 52225.0 25620.0 50880.0 ;
      RECT  24915.0 52225.0 25620.0 53570.0 ;
      RECT  24915.0 54915.0 25620.0 53570.0 ;
      RECT  24915.0 54915.0 25620.0 56260.0 ;
      RECT  24915.0 57605.0 25620.0 56260.0 ;
      RECT  24915.0 57605.0 25620.0 58950.0 ;
      RECT  24915.0 60295.0 25620.0 58950.0 ;
      RECT  24915.0 60295.0 25620.0 61640.0 ;
      RECT  24915.0 62985.0 25620.0 61640.0 ;
      RECT  24915.0 62985.0 25620.0 64330.0 ;
      RECT  24915.0 65675.0 25620.0 64330.0 ;
      RECT  24915.0 65675.0 25620.0 67020.0 ;
      RECT  24915.0 68365.0 25620.0 67020.0 ;
      RECT  24915.0 68365.0 25620.0 69710.0 ;
      RECT  24915.0 71055.0 25620.0 69710.0 ;
      RECT  24915.0 71055.0 25620.0 72400.0 ;
      RECT  24915.0 73745.0 25620.0 72400.0 ;
      RECT  24915.0 73745.0 25620.0 75090.0 ;
      RECT  24915.0 76435.0 25620.0 75090.0 ;
      RECT  24915.0 76435.0 25620.0 77780.0 ;
      RECT  24915.0 79125.0 25620.0 77780.0 ;
      RECT  24915.0 79125.0 25620.0 80470.0 ;
      RECT  24915.0 81815.0 25620.0 80470.0 ;
      RECT  24915.0 81815.0 25620.0 83160.0 ;
      RECT  24915.0 84505.0 25620.0 83160.0 ;
      RECT  24915.0 84505.0 25620.0 85850.0 ;
      RECT  24915.0 87195.0 25620.0 85850.0 ;
      RECT  24915.0 87195.0 25620.0 88540.0 ;
      RECT  24915.0 89885.0 25620.0 88540.0 ;
      RECT  24915.0 89885.0 25620.0 91230.0 ;
      RECT  24915.0 92575.0 25620.0 91230.0 ;
      RECT  24915.0 92575.0 25620.0 93920.0 ;
      RECT  24915.0 95265.0 25620.0 93920.0 ;
      RECT  24915.0 95265.0 25620.0 96610.0 ;
      RECT  24915.0 97955.0 25620.0 96610.0 ;
      RECT  24915.0 97955.0 25620.0 99300.0 ;
      RECT  24915.0 100645.0 25620.0 99300.0 ;
      RECT  24915.0 100645.0 25620.0 101990.0 ;
      RECT  24915.0 103335.0 25620.0 101990.0 ;
      RECT  24915.0 103335.0 25620.0 104680.0 ;
      RECT  24915.0 106025.0 25620.0 104680.0 ;
      RECT  24915.0 106025.0 25620.0 107370.0 ;
      RECT  24915.0 108715.0 25620.0 107370.0 ;
      RECT  24915.0 108715.0 25620.0 110060.0 ;
      RECT  24915.0 111405.0 25620.0 110060.0 ;
      RECT  24915.0 111405.0 25620.0 112750.0 ;
      RECT  24915.0 114095.0 25620.0 112750.0 ;
      RECT  25620.0 28015.0 26325.0 29360.0 ;
      RECT  25620.0 30705.0 26325.0 29360.0 ;
      RECT  25620.0 30705.0 26325.0 32050.0 ;
      RECT  25620.0 33395.0 26325.0 32050.0 ;
      RECT  25620.0 33395.0 26325.0 34740.0 ;
      RECT  25620.0 36085.0 26325.0 34740.0 ;
      RECT  25620.0 36085.0 26325.0 37430.0 ;
      RECT  25620.0 38775.0 26325.0 37430.0 ;
      RECT  25620.0 38775.0 26325.0 40120.0 ;
      RECT  25620.0 41465.0 26325.0 40120.0 ;
      RECT  25620.0 41465.0 26325.0 42810.0 ;
      RECT  25620.0 44155.0 26325.0 42810.0 ;
      RECT  25620.0 44155.0 26325.0 45500.0 ;
      RECT  25620.0 46845.0 26325.0 45500.0 ;
      RECT  25620.0 46845.0 26325.0 48190.0 ;
      RECT  25620.0 49535.0 26325.0 48190.0 ;
      RECT  25620.0 49535.0 26325.0 50880.0 ;
      RECT  25620.0 52225.0 26325.0 50880.0 ;
      RECT  25620.0 52225.0 26325.0 53570.0 ;
      RECT  25620.0 54915.0 26325.0 53570.0 ;
      RECT  25620.0 54915.0 26325.0 56260.0 ;
      RECT  25620.0 57605.0 26325.0 56260.0 ;
      RECT  25620.0 57605.0 26325.0 58950.0 ;
      RECT  25620.0 60295.0 26325.0 58950.0 ;
      RECT  25620.0 60295.0 26325.0 61640.0 ;
      RECT  25620.0 62985.0 26325.0 61640.0 ;
      RECT  25620.0 62985.0 26325.0 64330.0 ;
      RECT  25620.0 65675.0 26325.0 64330.0 ;
      RECT  25620.0 65675.0 26325.0 67020.0 ;
      RECT  25620.0 68365.0 26325.0 67020.0 ;
      RECT  25620.0 68365.0 26325.0 69710.0 ;
      RECT  25620.0 71055.0 26325.0 69710.0 ;
      RECT  25620.0 71055.0 26325.0 72400.0 ;
      RECT  25620.0 73745.0 26325.0 72400.0 ;
      RECT  25620.0 73745.0 26325.0 75090.0 ;
      RECT  25620.0 76435.0 26325.0 75090.0 ;
      RECT  25620.0 76435.0 26325.0 77780.0 ;
      RECT  25620.0 79125.0 26325.0 77780.0 ;
      RECT  25620.0 79125.0 26325.0 80470.0 ;
      RECT  25620.0 81815.0 26325.0 80470.0 ;
      RECT  25620.0 81815.0 26325.0 83160.0 ;
      RECT  25620.0 84505.0 26325.0 83160.0 ;
      RECT  25620.0 84505.0 26325.0 85850.0 ;
      RECT  25620.0 87195.0 26325.0 85850.0 ;
      RECT  25620.0 87195.0 26325.0 88540.0 ;
      RECT  25620.0 89885.0 26325.0 88540.0 ;
      RECT  25620.0 89885.0 26325.0 91230.0 ;
      RECT  25620.0 92575.0 26325.0 91230.0 ;
      RECT  25620.0 92575.0 26325.0 93920.0 ;
      RECT  25620.0 95265.0 26325.0 93920.0 ;
      RECT  25620.0 95265.0 26325.0 96610.0 ;
      RECT  25620.0 97955.0 26325.0 96610.0 ;
      RECT  25620.0 97955.0 26325.0 99300.0 ;
      RECT  25620.0 100645.0 26325.0 99300.0 ;
      RECT  25620.0 100645.0 26325.0 101990.0 ;
      RECT  25620.0 103335.0 26325.0 101990.0 ;
      RECT  25620.0 103335.0 26325.0 104680.0 ;
      RECT  25620.0 106025.0 26325.0 104680.0 ;
      RECT  25620.0 106025.0 26325.0 107370.0 ;
      RECT  25620.0 108715.0 26325.0 107370.0 ;
      RECT  25620.0 108715.0 26325.0 110060.0 ;
      RECT  25620.0 111405.0 26325.0 110060.0 ;
      RECT  25620.0 111405.0 26325.0 112750.0 ;
      RECT  25620.0 114095.0 26325.0 112750.0 ;
      RECT  26325.0 28015.0 27030.0 29360.0 ;
      RECT  26325.0 30705.0 27030.0 29360.0 ;
      RECT  26325.0 30705.0 27030.0 32050.0 ;
      RECT  26325.0 33395.0 27030.0 32050.0 ;
      RECT  26325.0 33395.0 27030.0 34740.0 ;
      RECT  26325.0 36085.0 27030.0 34740.0 ;
      RECT  26325.0 36085.0 27030.0 37430.0 ;
      RECT  26325.0 38775.0 27030.0 37430.0 ;
      RECT  26325.0 38775.0 27030.0 40120.0 ;
      RECT  26325.0 41465.0 27030.0 40120.0 ;
      RECT  26325.0 41465.0 27030.0 42810.0 ;
      RECT  26325.0 44155.0 27030.0 42810.0 ;
      RECT  26325.0 44155.0 27030.0 45500.0 ;
      RECT  26325.0 46845.0 27030.0 45500.0 ;
      RECT  26325.0 46845.0 27030.0 48190.0 ;
      RECT  26325.0 49535.0 27030.0 48190.0 ;
      RECT  26325.0 49535.0 27030.0 50880.0 ;
      RECT  26325.0 52225.0 27030.0 50880.0 ;
      RECT  26325.0 52225.0 27030.0 53570.0 ;
      RECT  26325.0 54915.0 27030.0 53570.0 ;
      RECT  26325.0 54915.0 27030.0 56260.0 ;
      RECT  26325.0 57605.0 27030.0 56260.0 ;
      RECT  26325.0 57605.0 27030.0 58950.0 ;
      RECT  26325.0 60295.0 27030.0 58950.0 ;
      RECT  26325.0 60295.0 27030.0 61640.0 ;
      RECT  26325.0 62985.0 27030.0 61640.0 ;
      RECT  26325.0 62985.0 27030.0 64330.0 ;
      RECT  26325.0 65675.0 27030.0 64330.0 ;
      RECT  26325.0 65675.0 27030.0 67020.0 ;
      RECT  26325.0 68365.0 27030.0 67020.0 ;
      RECT  26325.0 68365.0 27030.0 69710.0 ;
      RECT  26325.0 71055.0 27030.0 69710.0 ;
      RECT  26325.0 71055.0 27030.0 72400.0 ;
      RECT  26325.0 73745.0 27030.0 72400.0 ;
      RECT  26325.0 73745.0 27030.0 75090.0 ;
      RECT  26325.0 76435.0 27030.0 75090.0 ;
      RECT  26325.0 76435.0 27030.0 77780.0 ;
      RECT  26325.0 79125.0 27030.0 77780.0 ;
      RECT  26325.0 79125.0 27030.0 80470.0 ;
      RECT  26325.0 81815.0 27030.0 80470.0 ;
      RECT  26325.0 81815.0 27030.0 83160.0 ;
      RECT  26325.0 84505.0 27030.0 83160.0 ;
      RECT  26325.0 84505.0 27030.0 85850.0 ;
      RECT  26325.0 87195.0 27030.0 85850.0 ;
      RECT  26325.0 87195.0 27030.0 88540.0 ;
      RECT  26325.0 89885.0 27030.0 88540.0 ;
      RECT  26325.0 89885.0 27030.0 91230.0 ;
      RECT  26325.0 92575.0 27030.0 91230.0 ;
      RECT  26325.0 92575.0 27030.0 93920.0 ;
      RECT  26325.0 95265.0 27030.0 93920.0 ;
      RECT  26325.0 95265.0 27030.0 96610.0 ;
      RECT  26325.0 97955.0 27030.0 96610.0 ;
      RECT  26325.0 97955.0 27030.0 99300.0 ;
      RECT  26325.0 100645.0 27030.0 99300.0 ;
      RECT  26325.0 100645.0 27030.0 101990.0 ;
      RECT  26325.0 103335.0 27030.0 101990.0 ;
      RECT  26325.0 103335.0 27030.0 104680.0 ;
      RECT  26325.0 106025.0 27030.0 104680.0 ;
      RECT  26325.0 106025.0 27030.0 107370.0 ;
      RECT  26325.0 108715.0 27030.0 107370.0 ;
      RECT  26325.0 108715.0 27030.0 110060.0 ;
      RECT  26325.0 111405.0 27030.0 110060.0 ;
      RECT  26325.0 111405.0 27030.0 112750.0 ;
      RECT  26325.0 114095.0 27030.0 112750.0 ;
      RECT  27030.0 28015.0 27735.0 29360.0 ;
      RECT  27030.0 30705.0 27735.0 29360.0 ;
      RECT  27030.0 30705.0 27735.0 32050.0 ;
      RECT  27030.0 33395.0 27735.0 32050.0 ;
      RECT  27030.0 33395.0 27735.0 34740.0 ;
      RECT  27030.0 36085.0 27735.0 34740.0 ;
      RECT  27030.0 36085.0 27735.0 37430.0 ;
      RECT  27030.0 38775.0 27735.0 37430.0 ;
      RECT  27030.0 38775.0 27735.0 40120.0 ;
      RECT  27030.0 41465.0 27735.0 40120.0 ;
      RECT  27030.0 41465.0 27735.0 42810.0 ;
      RECT  27030.0 44155.0 27735.0 42810.0 ;
      RECT  27030.0 44155.0 27735.0 45500.0 ;
      RECT  27030.0 46845.0 27735.0 45500.0 ;
      RECT  27030.0 46845.0 27735.0 48190.0 ;
      RECT  27030.0 49535.0 27735.0 48190.0 ;
      RECT  27030.0 49535.0 27735.0 50880.0 ;
      RECT  27030.0 52225.0 27735.0 50880.0 ;
      RECT  27030.0 52225.0 27735.0 53570.0 ;
      RECT  27030.0 54915.0 27735.0 53570.0 ;
      RECT  27030.0 54915.0 27735.0 56260.0 ;
      RECT  27030.0 57605.0 27735.0 56260.0 ;
      RECT  27030.0 57605.0 27735.0 58950.0 ;
      RECT  27030.0 60295.0 27735.0 58950.0 ;
      RECT  27030.0 60295.0 27735.0 61640.0 ;
      RECT  27030.0 62985.0 27735.0 61640.0 ;
      RECT  27030.0 62985.0 27735.0 64330.0 ;
      RECT  27030.0 65675.0 27735.0 64330.0 ;
      RECT  27030.0 65675.0 27735.0 67020.0 ;
      RECT  27030.0 68365.0 27735.0 67020.0 ;
      RECT  27030.0 68365.0 27735.0 69710.0 ;
      RECT  27030.0 71055.0 27735.0 69710.0 ;
      RECT  27030.0 71055.0 27735.0 72400.0 ;
      RECT  27030.0 73745.0 27735.0 72400.0 ;
      RECT  27030.0 73745.0 27735.0 75090.0 ;
      RECT  27030.0 76435.0 27735.0 75090.0 ;
      RECT  27030.0 76435.0 27735.0 77780.0 ;
      RECT  27030.0 79125.0 27735.0 77780.0 ;
      RECT  27030.0 79125.0 27735.0 80470.0 ;
      RECT  27030.0 81815.0 27735.0 80470.0 ;
      RECT  27030.0 81815.0 27735.0 83160.0 ;
      RECT  27030.0 84505.0 27735.0 83160.0 ;
      RECT  27030.0 84505.0 27735.0 85850.0 ;
      RECT  27030.0 87195.0 27735.0 85850.0 ;
      RECT  27030.0 87195.0 27735.0 88540.0 ;
      RECT  27030.0 89885.0 27735.0 88540.0 ;
      RECT  27030.0 89885.0 27735.0 91230.0 ;
      RECT  27030.0 92575.0 27735.0 91230.0 ;
      RECT  27030.0 92575.0 27735.0 93920.0 ;
      RECT  27030.0 95265.0 27735.0 93920.0 ;
      RECT  27030.0 95265.0 27735.0 96610.0 ;
      RECT  27030.0 97955.0 27735.0 96610.0 ;
      RECT  27030.0 97955.0 27735.0 99300.0 ;
      RECT  27030.0 100645.0 27735.0 99300.0 ;
      RECT  27030.0 100645.0 27735.0 101990.0 ;
      RECT  27030.0 103335.0 27735.0 101990.0 ;
      RECT  27030.0 103335.0 27735.0 104680.0 ;
      RECT  27030.0 106025.0 27735.0 104680.0 ;
      RECT  27030.0 106025.0 27735.0 107370.0 ;
      RECT  27030.0 108715.0 27735.0 107370.0 ;
      RECT  27030.0 108715.0 27735.0 110060.0 ;
      RECT  27030.0 111405.0 27735.0 110060.0 ;
      RECT  27030.0 111405.0 27735.0 112750.0 ;
      RECT  27030.0 114095.0 27735.0 112750.0 ;
      RECT  27735.0 28015.0 28440.0 29360.0 ;
      RECT  27735.0 30705.0 28440.0 29360.0 ;
      RECT  27735.0 30705.0 28440.0 32050.0 ;
      RECT  27735.0 33395.0 28440.0 32050.0 ;
      RECT  27735.0 33395.0 28440.0 34740.0 ;
      RECT  27735.0 36085.0 28440.0 34740.0 ;
      RECT  27735.0 36085.0 28440.0 37430.0 ;
      RECT  27735.0 38775.0 28440.0 37430.0 ;
      RECT  27735.0 38775.0 28440.0 40120.0 ;
      RECT  27735.0 41465.0 28440.0 40120.0 ;
      RECT  27735.0 41465.0 28440.0 42810.0 ;
      RECT  27735.0 44155.0 28440.0 42810.0 ;
      RECT  27735.0 44155.0 28440.0 45500.0 ;
      RECT  27735.0 46845.0 28440.0 45500.0 ;
      RECT  27735.0 46845.0 28440.0 48190.0 ;
      RECT  27735.0 49535.0 28440.0 48190.0 ;
      RECT  27735.0 49535.0 28440.0 50880.0 ;
      RECT  27735.0 52225.0 28440.0 50880.0 ;
      RECT  27735.0 52225.0 28440.0 53570.0 ;
      RECT  27735.0 54915.0 28440.0 53570.0 ;
      RECT  27735.0 54915.0 28440.0 56260.0 ;
      RECT  27735.0 57605.0 28440.0 56260.0 ;
      RECT  27735.0 57605.0 28440.0 58950.0 ;
      RECT  27735.0 60295.0 28440.0 58950.0 ;
      RECT  27735.0 60295.0 28440.0 61640.0 ;
      RECT  27735.0 62985.0 28440.0 61640.0 ;
      RECT  27735.0 62985.0 28440.0 64330.0 ;
      RECT  27735.0 65675.0 28440.0 64330.0 ;
      RECT  27735.0 65675.0 28440.0 67020.0 ;
      RECT  27735.0 68365.0 28440.0 67020.0 ;
      RECT  27735.0 68365.0 28440.0 69710.0 ;
      RECT  27735.0 71055.0 28440.0 69710.0 ;
      RECT  27735.0 71055.0 28440.0 72400.0 ;
      RECT  27735.0 73745.0 28440.0 72400.0 ;
      RECT  27735.0 73745.0 28440.0 75090.0 ;
      RECT  27735.0 76435.0 28440.0 75090.0 ;
      RECT  27735.0 76435.0 28440.0 77780.0 ;
      RECT  27735.0 79125.0 28440.0 77780.0 ;
      RECT  27735.0 79125.0 28440.0 80470.0 ;
      RECT  27735.0 81815.0 28440.0 80470.0 ;
      RECT  27735.0 81815.0 28440.0 83160.0 ;
      RECT  27735.0 84505.0 28440.0 83160.0 ;
      RECT  27735.0 84505.0 28440.0 85850.0 ;
      RECT  27735.0 87195.0 28440.0 85850.0 ;
      RECT  27735.0 87195.0 28440.0 88540.0 ;
      RECT  27735.0 89885.0 28440.0 88540.0 ;
      RECT  27735.0 89885.0 28440.0 91230.0 ;
      RECT  27735.0 92575.0 28440.0 91230.0 ;
      RECT  27735.0 92575.0 28440.0 93920.0 ;
      RECT  27735.0 95265.0 28440.0 93920.0 ;
      RECT  27735.0 95265.0 28440.0 96610.0 ;
      RECT  27735.0 97955.0 28440.0 96610.0 ;
      RECT  27735.0 97955.0 28440.0 99300.0 ;
      RECT  27735.0 100645.0 28440.0 99300.0 ;
      RECT  27735.0 100645.0 28440.0 101990.0 ;
      RECT  27735.0 103335.0 28440.0 101990.0 ;
      RECT  27735.0 103335.0 28440.0 104680.0 ;
      RECT  27735.0 106025.0 28440.0 104680.0 ;
      RECT  27735.0 106025.0 28440.0 107370.0 ;
      RECT  27735.0 108715.0 28440.0 107370.0 ;
      RECT  27735.0 108715.0 28440.0 110060.0 ;
      RECT  27735.0 111405.0 28440.0 110060.0 ;
      RECT  27735.0 111405.0 28440.0 112750.0 ;
      RECT  27735.0 114095.0 28440.0 112750.0 ;
      RECT  28440.0 28015.0 29145.0 29360.0 ;
      RECT  28440.0 30705.0 29145.0 29360.0 ;
      RECT  28440.0 30705.0 29145.0 32050.0 ;
      RECT  28440.0 33395.0 29145.0 32050.0 ;
      RECT  28440.0 33395.0 29145.0 34740.0 ;
      RECT  28440.0 36085.0 29145.0 34740.0 ;
      RECT  28440.0 36085.0 29145.0 37430.0 ;
      RECT  28440.0 38775.0 29145.0 37430.0 ;
      RECT  28440.0 38775.0 29145.0 40120.0 ;
      RECT  28440.0 41465.0 29145.0 40120.0 ;
      RECT  28440.0 41465.0 29145.0 42810.0 ;
      RECT  28440.0 44155.0 29145.0 42810.0 ;
      RECT  28440.0 44155.0 29145.0 45500.0 ;
      RECT  28440.0 46845.0 29145.0 45500.0 ;
      RECT  28440.0 46845.0 29145.0 48190.0 ;
      RECT  28440.0 49535.0 29145.0 48190.0 ;
      RECT  28440.0 49535.0 29145.0 50880.0 ;
      RECT  28440.0 52225.0 29145.0 50880.0 ;
      RECT  28440.0 52225.0 29145.0 53570.0 ;
      RECT  28440.0 54915.0 29145.0 53570.0 ;
      RECT  28440.0 54915.0 29145.0 56260.0 ;
      RECT  28440.0 57605.0 29145.0 56260.0 ;
      RECT  28440.0 57605.0 29145.0 58950.0 ;
      RECT  28440.0 60295.0 29145.0 58950.0 ;
      RECT  28440.0 60295.0 29145.0 61640.0 ;
      RECT  28440.0 62985.0 29145.0 61640.0 ;
      RECT  28440.0 62985.0 29145.0 64330.0 ;
      RECT  28440.0 65675.0 29145.0 64330.0 ;
      RECT  28440.0 65675.0 29145.0 67020.0 ;
      RECT  28440.0 68365.0 29145.0 67020.0 ;
      RECT  28440.0 68365.0 29145.0 69710.0 ;
      RECT  28440.0 71055.0 29145.0 69710.0 ;
      RECT  28440.0 71055.0 29145.0 72400.0 ;
      RECT  28440.0 73745.0 29145.0 72400.0 ;
      RECT  28440.0 73745.0 29145.0 75090.0 ;
      RECT  28440.0 76435.0 29145.0 75090.0 ;
      RECT  28440.0 76435.0 29145.0 77780.0 ;
      RECT  28440.0 79125.0 29145.0 77780.0 ;
      RECT  28440.0 79125.0 29145.0 80470.0 ;
      RECT  28440.0 81815.0 29145.0 80470.0 ;
      RECT  28440.0 81815.0 29145.0 83160.0 ;
      RECT  28440.0 84505.0 29145.0 83160.0 ;
      RECT  28440.0 84505.0 29145.0 85850.0 ;
      RECT  28440.0 87195.0 29145.0 85850.0 ;
      RECT  28440.0 87195.0 29145.0 88540.0 ;
      RECT  28440.0 89885.0 29145.0 88540.0 ;
      RECT  28440.0 89885.0 29145.0 91230.0 ;
      RECT  28440.0 92575.0 29145.0 91230.0 ;
      RECT  28440.0 92575.0 29145.0 93920.0 ;
      RECT  28440.0 95265.0 29145.0 93920.0 ;
      RECT  28440.0 95265.0 29145.0 96610.0 ;
      RECT  28440.0 97955.0 29145.0 96610.0 ;
      RECT  28440.0 97955.0 29145.0 99300.0 ;
      RECT  28440.0 100645.0 29145.0 99300.0 ;
      RECT  28440.0 100645.0 29145.0 101990.0 ;
      RECT  28440.0 103335.0 29145.0 101990.0 ;
      RECT  28440.0 103335.0 29145.0 104680.0 ;
      RECT  28440.0 106025.0 29145.0 104680.0 ;
      RECT  28440.0 106025.0 29145.0 107370.0 ;
      RECT  28440.0 108715.0 29145.0 107370.0 ;
      RECT  28440.0 108715.0 29145.0 110060.0 ;
      RECT  28440.0 111405.0 29145.0 110060.0 ;
      RECT  28440.0 111405.0 29145.0 112750.0 ;
      RECT  28440.0 114095.0 29145.0 112750.0 ;
      RECT  29145.0 28015.0 29850.0 29360.0 ;
      RECT  29145.0 30705.0 29850.0 29360.0 ;
      RECT  29145.0 30705.0 29850.0 32050.0 ;
      RECT  29145.0 33395.0 29850.0 32050.0 ;
      RECT  29145.0 33395.0 29850.0 34740.0 ;
      RECT  29145.0 36085.0 29850.0 34740.0 ;
      RECT  29145.0 36085.0 29850.0 37430.0 ;
      RECT  29145.0 38775.0 29850.0 37430.0 ;
      RECT  29145.0 38775.0 29850.0 40120.0 ;
      RECT  29145.0 41465.0 29850.0 40120.0 ;
      RECT  29145.0 41465.0 29850.0 42810.0 ;
      RECT  29145.0 44155.0 29850.0 42810.0 ;
      RECT  29145.0 44155.0 29850.0 45500.0 ;
      RECT  29145.0 46845.0 29850.0 45500.0 ;
      RECT  29145.0 46845.0 29850.0 48190.0 ;
      RECT  29145.0 49535.0 29850.0 48190.0 ;
      RECT  29145.0 49535.0 29850.0 50880.0 ;
      RECT  29145.0 52225.0 29850.0 50880.0 ;
      RECT  29145.0 52225.0 29850.0 53570.0 ;
      RECT  29145.0 54915.0 29850.0 53570.0 ;
      RECT  29145.0 54915.0 29850.0 56260.0 ;
      RECT  29145.0 57605.0 29850.0 56260.0 ;
      RECT  29145.0 57605.0 29850.0 58950.0 ;
      RECT  29145.0 60295.0 29850.0 58950.0 ;
      RECT  29145.0 60295.0 29850.0 61640.0 ;
      RECT  29145.0 62985.0 29850.0 61640.0 ;
      RECT  29145.0 62985.0 29850.0 64330.0 ;
      RECT  29145.0 65675.0 29850.0 64330.0 ;
      RECT  29145.0 65675.0 29850.0 67020.0 ;
      RECT  29145.0 68365.0 29850.0 67020.0 ;
      RECT  29145.0 68365.0 29850.0 69710.0 ;
      RECT  29145.0 71055.0 29850.0 69710.0 ;
      RECT  29145.0 71055.0 29850.0 72400.0 ;
      RECT  29145.0 73745.0 29850.0 72400.0 ;
      RECT  29145.0 73745.0 29850.0 75090.0 ;
      RECT  29145.0 76435.0 29850.0 75090.0 ;
      RECT  29145.0 76435.0 29850.0 77780.0 ;
      RECT  29145.0 79125.0 29850.0 77780.0 ;
      RECT  29145.0 79125.0 29850.0 80470.0 ;
      RECT  29145.0 81815.0 29850.0 80470.0 ;
      RECT  29145.0 81815.0 29850.0 83160.0 ;
      RECT  29145.0 84505.0 29850.0 83160.0 ;
      RECT  29145.0 84505.0 29850.0 85850.0 ;
      RECT  29145.0 87195.0 29850.0 85850.0 ;
      RECT  29145.0 87195.0 29850.0 88540.0 ;
      RECT  29145.0 89885.0 29850.0 88540.0 ;
      RECT  29145.0 89885.0 29850.0 91230.0 ;
      RECT  29145.0 92575.0 29850.0 91230.0 ;
      RECT  29145.0 92575.0 29850.0 93920.0 ;
      RECT  29145.0 95265.0 29850.0 93920.0 ;
      RECT  29145.0 95265.0 29850.0 96610.0 ;
      RECT  29145.0 97955.0 29850.0 96610.0 ;
      RECT  29145.0 97955.0 29850.0 99300.0 ;
      RECT  29145.0 100645.0 29850.0 99300.0 ;
      RECT  29145.0 100645.0 29850.0 101990.0 ;
      RECT  29145.0 103335.0 29850.0 101990.0 ;
      RECT  29145.0 103335.0 29850.0 104680.0 ;
      RECT  29145.0 106025.0 29850.0 104680.0 ;
      RECT  29145.0 106025.0 29850.0 107370.0 ;
      RECT  29145.0 108715.0 29850.0 107370.0 ;
      RECT  29145.0 108715.0 29850.0 110060.0 ;
      RECT  29145.0 111405.0 29850.0 110060.0 ;
      RECT  29145.0 111405.0 29850.0 112750.0 ;
      RECT  29145.0 114095.0 29850.0 112750.0 ;
      RECT  29850.0 28015.0 30555.0 29360.0 ;
      RECT  29850.0 30705.0 30555.0 29360.0 ;
      RECT  29850.0 30705.0 30555.0 32050.0 ;
      RECT  29850.0 33395.0 30555.0 32050.0 ;
      RECT  29850.0 33395.0 30555.0 34740.0 ;
      RECT  29850.0 36085.0 30555.0 34740.0 ;
      RECT  29850.0 36085.0 30555.0 37430.0 ;
      RECT  29850.0 38775.0 30555.0 37430.0 ;
      RECT  29850.0 38775.0 30555.0 40120.0 ;
      RECT  29850.0 41465.0 30555.0 40120.0 ;
      RECT  29850.0 41465.0 30555.0 42810.0 ;
      RECT  29850.0 44155.0 30555.0 42810.0 ;
      RECT  29850.0 44155.0 30555.0 45500.0 ;
      RECT  29850.0 46845.0 30555.0 45500.0 ;
      RECT  29850.0 46845.0 30555.0 48190.0 ;
      RECT  29850.0 49535.0 30555.0 48190.0 ;
      RECT  29850.0 49535.0 30555.0 50880.0 ;
      RECT  29850.0 52225.0 30555.0 50880.0 ;
      RECT  29850.0 52225.0 30555.0 53570.0 ;
      RECT  29850.0 54915.0 30555.0 53570.0 ;
      RECT  29850.0 54915.0 30555.0 56260.0 ;
      RECT  29850.0 57605.0 30555.0 56260.0 ;
      RECT  29850.0 57605.0 30555.0 58950.0 ;
      RECT  29850.0 60295.0 30555.0 58950.0 ;
      RECT  29850.0 60295.0 30555.0 61640.0 ;
      RECT  29850.0 62985.0 30555.0 61640.0 ;
      RECT  29850.0 62985.0 30555.0 64330.0 ;
      RECT  29850.0 65675.0 30555.0 64330.0 ;
      RECT  29850.0 65675.0 30555.0 67020.0 ;
      RECT  29850.0 68365.0 30555.0 67020.0 ;
      RECT  29850.0 68365.0 30555.0 69710.0 ;
      RECT  29850.0 71055.0 30555.0 69710.0 ;
      RECT  29850.0 71055.0 30555.0 72400.0 ;
      RECT  29850.0 73745.0 30555.0 72400.0 ;
      RECT  29850.0 73745.0 30555.0 75090.0 ;
      RECT  29850.0 76435.0 30555.0 75090.0 ;
      RECT  29850.0 76435.0 30555.0 77780.0 ;
      RECT  29850.0 79125.0 30555.0 77780.0 ;
      RECT  29850.0 79125.0 30555.0 80470.0 ;
      RECT  29850.0 81815.0 30555.0 80470.0 ;
      RECT  29850.0 81815.0 30555.0 83160.0 ;
      RECT  29850.0 84505.0 30555.0 83160.0 ;
      RECT  29850.0 84505.0 30555.0 85850.0 ;
      RECT  29850.0 87195.0 30555.0 85850.0 ;
      RECT  29850.0 87195.0 30555.0 88540.0 ;
      RECT  29850.0 89885.0 30555.0 88540.0 ;
      RECT  29850.0 89885.0 30555.0 91230.0 ;
      RECT  29850.0 92575.0 30555.0 91230.0 ;
      RECT  29850.0 92575.0 30555.0 93920.0 ;
      RECT  29850.0 95265.0 30555.0 93920.0 ;
      RECT  29850.0 95265.0 30555.0 96610.0 ;
      RECT  29850.0 97955.0 30555.0 96610.0 ;
      RECT  29850.0 97955.0 30555.0 99300.0 ;
      RECT  29850.0 100645.0 30555.0 99300.0 ;
      RECT  29850.0 100645.0 30555.0 101990.0 ;
      RECT  29850.0 103335.0 30555.0 101990.0 ;
      RECT  29850.0 103335.0 30555.0 104680.0 ;
      RECT  29850.0 106025.0 30555.0 104680.0 ;
      RECT  29850.0 106025.0 30555.0 107370.0 ;
      RECT  29850.0 108715.0 30555.0 107370.0 ;
      RECT  29850.0 108715.0 30555.0 110060.0 ;
      RECT  29850.0 111405.0 30555.0 110060.0 ;
      RECT  29850.0 111405.0 30555.0 112750.0 ;
      RECT  29850.0 114095.0 30555.0 112750.0 ;
      RECT  30555.0 28015.0 31260.0 29360.0 ;
      RECT  30555.0 30705.0 31260.0 29360.0 ;
      RECT  30555.0 30705.0 31260.0 32050.0 ;
      RECT  30555.0 33395.0 31260.0 32050.0 ;
      RECT  30555.0 33395.0 31260.0 34740.0 ;
      RECT  30555.0 36085.0 31260.0 34740.0 ;
      RECT  30555.0 36085.0 31260.0 37430.0 ;
      RECT  30555.0 38775.0 31260.0 37430.0 ;
      RECT  30555.0 38775.0 31260.0 40120.0 ;
      RECT  30555.0 41465.0 31260.0 40120.0 ;
      RECT  30555.0 41465.0 31260.0 42810.0 ;
      RECT  30555.0 44155.0 31260.0 42810.0 ;
      RECT  30555.0 44155.0 31260.0 45500.0 ;
      RECT  30555.0 46845.0 31260.0 45500.0 ;
      RECT  30555.0 46845.0 31260.0 48190.0 ;
      RECT  30555.0 49535.0 31260.0 48190.0 ;
      RECT  30555.0 49535.0 31260.0 50880.0 ;
      RECT  30555.0 52225.0 31260.0 50880.0 ;
      RECT  30555.0 52225.0 31260.0 53570.0 ;
      RECT  30555.0 54915.0 31260.0 53570.0 ;
      RECT  30555.0 54915.0 31260.0 56260.0 ;
      RECT  30555.0 57605.0 31260.0 56260.0 ;
      RECT  30555.0 57605.0 31260.0 58950.0 ;
      RECT  30555.0 60295.0 31260.0 58950.0 ;
      RECT  30555.0 60295.0 31260.0 61640.0 ;
      RECT  30555.0 62985.0 31260.0 61640.0 ;
      RECT  30555.0 62985.0 31260.0 64330.0 ;
      RECT  30555.0 65675.0 31260.0 64330.0 ;
      RECT  30555.0 65675.0 31260.0 67020.0 ;
      RECT  30555.0 68365.0 31260.0 67020.0 ;
      RECT  30555.0 68365.0 31260.0 69710.0 ;
      RECT  30555.0 71055.0 31260.0 69710.0 ;
      RECT  30555.0 71055.0 31260.0 72400.0 ;
      RECT  30555.0 73745.0 31260.0 72400.0 ;
      RECT  30555.0 73745.0 31260.0 75090.0 ;
      RECT  30555.0 76435.0 31260.0 75090.0 ;
      RECT  30555.0 76435.0 31260.0 77780.0 ;
      RECT  30555.0 79125.0 31260.0 77780.0 ;
      RECT  30555.0 79125.0 31260.0 80470.0 ;
      RECT  30555.0 81815.0 31260.0 80470.0 ;
      RECT  30555.0 81815.0 31260.0 83160.0 ;
      RECT  30555.0 84505.0 31260.0 83160.0 ;
      RECT  30555.0 84505.0 31260.0 85850.0 ;
      RECT  30555.0 87195.0 31260.0 85850.0 ;
      RECT  30555.0 87195.0 31260.0 88540.0 ;
      RECT  30555.0 89885.0 31260.0 88540.0 ;
      RECT  30555.0 89885.0 31260.0 91230.0 ;
      RECT  30555.0 92575.0 31260.0 91230.0 ;
      RECT  30555.0 92575.0 31260.0 93920.0 ;
      RECT  30555.0 95265.0 31260.0 93920.0 ;
      RECT  30555.0 95265.0 31260.0 96610.0 ;
      RECT  30555.0 97955.0 31260.0 96610.0 ;
      RECT  30555.0 97955.0 31260.0 99300.0 ;
      RECT  30555.0 100645.0 31260.0 99300.0 ;
      RECT  30555.0 100645.0 31260.0 101990.0 ;
      RECT  30555.0 103335.0 31260.0 101990.0 ;
      RECT  30555.0 103335.0 31260.0 104680.0 ;
      RECT  30555.0 106025.0 31260.0 104680.0 ;
      RECT  30555.0 106025.0 31260.0 107370.0 ;
      RECT  30555.0 108715.0 31260.0 107370.0 ;
      RECT  30555.0 108715.0 31260.0 110060.0 ;
      RECT  30555.0 111405.0 31260.0 110060.0 ;
      RECT  30555.0 111405.0 31260.0 112750.0 ;
      RECT  30555.0 114095.0 31260.0 112750.0 ;
      RECT  31260.0 28015.0 31965.0 29360.0 ;
      RECT  31260.0 30705.0 31965.0 29360.0 ;
      RECT  31260.0 30705.0 31965.0 32050.0 ;
      RECT  31260.0 33395.0 31965.0 32050.0 ;
      RECT  31260.0 33395.0 31965.0 34740.0 ;
      RECT  31260.0 36085.0 31965.0 34740.0 ;
      RECT  31260.0 36085.0 31965.0 37430.0 ;
      RECT  31260.0 38775.0 31965.0 37430.0 ;
      RECT  31260.0 38775.0 31965.0 40120.0 ;
      RECT  31260.0 41465.0 31965.0 40120.0 ;
      RECT  31260.0 41465.0 31965.0 42810.0 ;
      RECT  31260.0 44155.0 31965.0 42810.0 ;
      RECT  31260.0 44155.0 31965.0 45500.0 ;
      RECT  31260.0 46845.0 31965.0 45500.0 ;
      RECT  31260.0 46845.0 31965.0 48190.0 ;
      RECT  31260.0 49535.0 31965.0 48190.0 ;
      RECT  31260.0 49535.0 31965.0 50880.0 ;
      RECT  31260.0 52225.0 31965.0 50880.0 ;
      RECT  31260.0 52225.0 31965.0 53570.0 ;
      RECT  31260.0 54915.0 31965.0 53570.0 ;
      RECT  31260.0 54915.0 31965.0 56260.0 ;
      RECT  31260.0 57605.0 31965.0 56260.0 ;
      RECT  31260.0 57605.0 31965.0 58950.0 ;
      RECT  31260.0 60295.0 31965.0 58950.0 ;
      RECT  31260.0 60295.0 31965.0 61640.0 ;
      RECT  31260.0 62985.0 31965.0 61640.0 ;
      RECT  31260.0 62985.0 31965.0 64330.0 ;
      RECT  31260.0 65675.0 31965.0 64330.0 ;
      RECT  31260.0 65675.0 31965.0 67020.0 ;
      RECT  31260.0 68365.0 31965.0 67020.0 ;
      RECT  31260.0 68365.0 31965.0 69710.0 ;
      RECT  31260.0 71055.0 31965.0 69710.0 ;
      RECT  31260.0 71055.0 31965.0 72400.0 ;
      RECT  31260.0 73745.0 31965.0 72400.0 ;
      RECT  31260.0 73745.0 31965.0 75090.0 ;
      RECT  31260.0 76435.0 31965.0 75090.0 ;
      RECT  31260.0 76435.0 31965.0 77780.0 ;
      RECT  31260.0 79125.0 31965.0 77780.0 ;
      RECT  31260.0 79125.0 31965.0 80470.0 ;
      RECT  31260.0 81815.0 31965.0 80470.0 ;
      RECT  31260.0 81815.0 31965.0 83160.0 ;
      RECT  31260.0 84505.0 31965.0 83160.0 ;
      RECT  31260.0 84505.0 31965.0 85850.0 ;
      RECT  31260.0 87195.0 31965.0 85850.0 ;
      RECT  31260.0 87195.0 31965.0 88540.0 ;
      RECT  31260.0 89885.0 31965.0 88540.0 ;
      RECT  31260.0 89885.0 31965.0 91230.0 ;
      RECT  31260.0 92575.0 31965.0 91230.0 ;
      RECT  31260.0 92575.0 31965.0 93920.0 ;
      RECT  31260.0 95265.0 31965.0 93920.0 ;
      RECT  31260.0 95265.0 31965.0 96610.0 ;
      RECT  31260.0 97955.0 31965.0 96610.0 ;
      RECT  31260.0 97955.0 31965.0 99300.0 ;
      RECT  31260.0 100645.0 31965.0 99300.0 ;
      RECT  31260.0 100645.0 31965.0 101990.0 ;
      RECT  31260.0 103335.0 31965.0 101990.0 ;
      RECT  31260.0 103335.0 31965.0 104680.0 ;
      RECT  31260.0 106025.0 31965.0 104680.0 ;
      RECT  31260.0 106025.0 31965.0 107370.0 ;
      RECT  31260.0 108715.0 31965.0 107370.0 ;
      RECT  31260.0 108715.0 31965.0 110060.0 ;
      RECT  31260.0 111405.0 31965.0 110060.0 ;
      RECT  31260.0 111405.0 31965.0 112750.0 ;
      RECT  31260.0 114095.0 31965.0 112750.0 ;
      RECT  31965.0 28015.0 32670.0 29360.0 ;
      RECT  31965.0 30705.0 32670.0 29360.0 ;
      RECT  31965.0 30705.0 32670.0 32050.0 ;
      RECT  31965.0 33395.0 32670.0 32050.0 ;
      RECT  31965.0 33395.0 32670.0 34740.0 ;
      RECT  31965.0 36085.0 32670.0 34740.0 ;
      RECT  31965.0 36085.0 32670.0 37430.0 ;
      RECT  31965.0 38775.0 32670.0 37430.0 ;
      RECT  31965.0 38775.0 32670.0 40120.0 ;
      RECT  31965.0 41465.0 32670.0 40120.0 ;
      RECT  31965.0 41465.0 32670.0 42810.0 ;
      RECT  31965.0 44155.0 32670.0 42810.0 ;
      RECT  31965.0 44155.0 32670.0 45500.0 ;
      RECT  31965.0 46845.0 32670.0 45500.0 ;
      RECT  31965.0 46845.0 32670.0 48190.0 ;
      RECT  31965.0 49535.0 32670.0 48190.0 ;
      RECT  31965.0 49535.0 32670.0 50880.0 ;
      RECT  31965.0 52225.0 32670.0 50880.0 ;
      RECT  31965.0 52225.0 32670.0 53570.0 ;
      RECT  31965.0 54915.0 32670.0 53570.0 ;
      RECT  31965.0 54915.0 32670.0 56260.0 ;
      RECT  31965.0 57605.0 32670.0 56260.0 ;
      RECT  31965.0 57605.0 32670.0 58950.0 ;
      RECT  31965.0 60295.0 32670.0 58950.0 ;
      RECT  31965.0 60295.0 32670.0 61640.0 ;
      RECT  31965.0 62985.0 32670.0 61640.0 ;
      RECT  31965.0 62985.0 32670.0 64330.0 ;
      RECT  31965.0 65675.0 32670.0 64330.0 ;
      RECT  31965.0 65675.0 32670.0 67020.0 ;
      RECT  31965.0 68365.0 32670.0 67020.0 ;
      RECT  31965.0 68365.0 32670.0 69710.0 ;
      RECT  31965.0 71055.0 32670.0 69710.0 ;
      RECT  31965.0 71055.0 32670.0 72400.0 ;
      RECT  31965.0 73745.0 32670.0 72400.0 ;
      RECT  31965.0 73745.0 32670.0 75090.0 ;
      RECT  31965.0 76435.0 32670.0 75090.0 ;
      RECT  31965.0 76435.0 32670.0 77780.0 ;
      RECT  31965.0 79125.0 32670.0 77780.0 ;
      RECT  31965.0 79125.0 32670.0 80470.0 ;
      RECT  31965.0 81815.0 32670.0 80470.0 ;
      RECT  31965.0 81815.0 32670.0 83160.0 ;
      RECT  31965.0 84505.0 32670.0 83160.0 ;
      RECT  31965.0 84505.0 32670.0 85850.0 ;
      RECT  31965.0 87195.0 32670.0 85850.0 ;
      RECT  31965.0 87195.0 32670.0 88540.0 ;
      RECT  31965.0 89885.0 32670.0 88540.0 ;
      RECT  31965.0 89885.0 32670.0 91230.0 ;
      RECT  31965.0 92575.0 32670.0 91230.0 ;
      RECT  31965.0 92575.0 32670.0 93920.0 ;
      RECT  31965.0 95265.0 32670.0 93920.0 ;
      RECT  31965.0 95265.0 32670.0 96610.0 ;
      RECT  31965.0 97955.0 32670.0 96610.0 ;
      RECT  31965.0 97955.0 32670.0 99300.0 ;
      RECT  31965.0 100645.0 32670.0 99300.0 ;
      RECT  31965.0 100645.0 32670.0 101990.0 ;
      RECT  31965.0 103335.0 32670.0 101990.0 ;
      RECT  31965.0 103335.0 32670.0 104680.0 ;
      RECT  31965.0 106025.0 32670.0 104680.0 ;
      RECT  31965.0 106025.0 32670.0 107370.0 ;
      RECT  31965.0 108715.0 32670.0 107370.0 ;
      RECT  31965.0 108715.0 32670.0 110060.0 ;
      RECT  31965.0 111405.0 32670.0 110060.0 ;
      RECT  31965.0 111405.0 32670.0 112750.0 ;
      RECT  31965.0 114095.0 32670.0 112750.0 ;
      RECT  32670.0 28015.0 33375.0 29360.0 ;
      RECT  32670.0 30705.0 33375.0 29360.0 ;
      RECT  32670.0 30705.0 33375.0 32050.0 ;
      RECT  32670.0 33395.0 33375.0 32050.0 ;
      RECT  32670.0 33395.0 33375.0 34740.0 ;
      RECT  32670.0 36085.0 33375.0 34740.0 ;
      RECT  32670.0 36085.0 33375.0 37430.0 ;
      RECT  32670.0 38775.0 33375.0 37430.0 ;
      RECT  32670.0 38775.0 33375.0 40120.0 ;
      RECT  32670.0 41465.0 33375.0 40120.0 ;
      RECT  32670.0 41465.0 33375.0 42810.0 ;
      RECT  32670.0 44155.0 33375.0 42810.0 ;
      RECT  32670.0 44155.0 33375.0 45500.0 ;
      RECT  32670.0 46845.0 33375.0 45500.0 ;
      RECT  32670.0 46845.0 33375.0 48190.0 ;
      RECT  32670.0 49535.0 33375.0 48190.0 ;
      RECT  32670.0 49535.0 33375.0 50880.0 ;
      RECT  32670.0 52225.0 33375.0 50880.0 ;
      RECT  32670.0 52225.0 33375.0 53570.0 ;
      RECT  32670.0 54915.0 33375.0 53570.0 ;
      RECT  32670.0 54915.0 33375.0 56260.0 ;
      RECT  32670.0 57605.0 33375.0 56260.0 ;
      RECT  32670.0 57605.0 33375.0 58950.0 ;
      RECT  32670.0 60295.0 33375.0 58950.0 ;
      RECT  32670.0 60295.0 33375.0 61640.0 ;
      RECT  32670.0 62985.0 33375.0 61640.0 ;
      RECT  32670.0 62985.0 33375.0 64330.0 ;
      RECT  32670.0 65675.0 33375.0 64330.0 ;
      RECT  32670.0 65675.0 33375.0 67020.0 ;
      RECT  32670.0 68365.0 33375.0 67020.0 ;
      RECT  32670.0 68365.0 33375.0 69710.0 ;
      RECT  32670.0 71055.0 33375.0 69710.0 ;
      RECT  32670.0 71055.0 33375.0 72400.0 ;
      RECT  32670.0 73745.0 33375.0 72400.0 ;
      RECT  32670.0 73745.0 33375.0 75090.0 ;
      RECT  32670.0 76435.0 33375.0 75090.0 ;
      RECT  32670.0 76435.0 33375.0 77780.0 ;
      RECT  32670.0 79125.0 33375.0 77780.0 ;
      RECT  32670.0 79125.0 33375.0 80470.0 ;
      RECT  32670.0 81815.0 33375.0 80470.0 ;
      RECT  32670.0 81815.0 33375.0 83160.0 ;
      RECT  32670.0 84505.0 33375.0 83160.0 ;
      RECT  32670.0 84505.0 33375.0 85850.0 ;
      RECT  32670.0 87195.0 33375.0 85850.0 ;
      RECT  32670.0 87195.0 33375.0 88540.0 ;
      RECT  32670.0 89885.0 33375.0 88540.0 ;
      RECT  32670.0 89885.0 33375.0 91230.0 ;
      RECT  32670.0 92575.0 33375.0 91230.0 ;
      RECT  32670.0 92575.0 33375.0 93920.0 ;
      RECT  32670.0 95265.0 33375.0 93920.0 ;
      RECT  32670.0 95265.0 33375.0 96610.0 ;
      RECT  32670.0 97955.0 33375.0 96610.0 ;
      RECT  32670.0 97955.0 33375.0 99300.0 ;
      RECT  32670.0 100645.0 33375.0 99300.0 ;
      RECT  32670.0 100645.0 33375.0 101990.0 ;
      RECT  32670.0 103335.0 33375.0 101990.0 ;
      RECT  32670.0 103335.0 33375.0 104680.0 ;
      RECT  32670.0 106025.0 33375.0 104680.0 ;
      RECT  32670.0 106025.0 33375.0 107370.0 ;
      RECT  32670.0 108715.0 33375.0 107370.0 ;
      RECT  32670.0 108715.0 33375.0 110060.0 ;
      RECT  32670.0 111405.0 33375.0 110060.0 ;
      RECT  32670.0 111405.0 33375.0 112750.0 ;
      RECT  32670.0 114095.0 33375.0 112750.0 ;
      RECT  33375.0 28015.0 34080.0 29360.0 ;
      RECT  33375.0 30705.0 34080.0 29360.0 ;
      RECT  33375.0 30705.0 34080.0 32050.0 ;
      RECT  33375.0 33395.0 34080.0 32050.0 ;
      RECT  33375.0 33395.0 34080.0 34740.0 ;
      RECT  33375.0 36085.0 34080.0 34740.0 ;
      RECT  33375.0 36085.0 34080.0 37430.0 ;
      RECT  33375.0 38775.0 34080.0 37430.0 ;
      RECT  33375.0 38775.0 34080.0 40120.0 ;
      RECT  33375.0 41465.0 34080.0 40120.0 ;
      RECT  33375.0 41465.0 34080.0 42810.0 ;
      RECT  33375.0 44155.0 34080.0 42810.0 ;
      RECT  33375.0 44155.0 34080.0 45500.0 ;
      RECT  33375.0 46845.0 34080.0 45500.0 ;
      RECT  33375.0 46845.0 34080.0 48190.0 ;
      RECT  33375.0 49535.0 34080.0 48190.0 ;
      RECT  33375.0 49535.0 34080.0 50880.0 ;
      RECT  33375.0 52225.0 34080.0 50880.0 ;
      RECT  33375.0 52225.0 34080.0 53570.0 ;
      RECT  33375.0 54915.0 34080.0 53570.0 ;
      RECT  33375.0 54915.0 34080.0 56260.0 ;
      RECT  33375.0 57605.0 34080.0 56260.0 ;
      RECT  33375.0 57605.0 34080.0 58950.0 ;
      RECT  33375.0 60295.0 34080.0 58950.0 ;
      RECT  33375.0 60295.0 34080.0 61640.0 ;
      RECT  33375.0 62985.0 34080.0 61640.0 ;
      RECT  33375.0 62985.0 34080.0 64330.0 ;
      RECT  33375.0 65675.0 34080.0 64330.0 ;
      RECT  33375.0 65675.0 34080.0 67020.0 ;
      RECT  33375.0 68365.0 34080.0 67020.0 ;
      RECT  33375.0 68365.0 34080.0 69710.0 ;
      RECT  33375.0 71055.0 34080.0 69710.0 ;
      RECT  33375.0 71055.0 34080.0 72400.0 ;
      RECT  33375.0 73745.0 34080.0 72400.0 ;
      RECT  33375.0 73745.0 34080.0 75090.0 ;
      RECT  33375.0 76435.0 34080.0 75090.0 ;
      RECT  33375.0 76435.0 34080.0 77780.0 ;
      RECT  33375.0 79125.0 34080.0 77780.0 ;
      RECT  33375.0 79125.0 34080.0 80470.0 ;
      RECT  33375.0 81815.0 34080.0 80470.0 ;
      RECT  33375.0 81815.0 34080.0 83160.0 ;
      RECT  33375.0 84505.0 34080.0 83160.0 ;
      RECT  33375.0 84505.0 34080.0 85850.0 ;
      RECT  33375.0 87195.0 34080.0 85850.0 ;
      RECT  33375.0 87195.0 34080.0 88540.0 ;
      RECT  33375.0 89885.0 34080.0 88540.0 ;
      RECT  33375.0 89885.0 34080.0 91230.0 ;
      RECT  33375.0 92575.0 34080.0 91230.0 ;
      RECT  33375.0 92575.0 34080.0 93920.0 ;
      RECT  33375.0 95265.0 34080.0 93920.0 ;
      RECT  33375.0 95265.0 34080.0 96610.0 ;
      RECT  33375.0 97955.0 34080.0 96610.0 ;
      RECT  33375.0 97955.0 34080.0 99300.0 ;
      RECT  33375.0 100645.0 34080.0 99300.0 ;
      RECT  33375.0 100645.0 34080.0 101990.0 ;
      RECT  33375.0 103335.0 34080.0 101990.0 ;
      RECT  33375.0 103335.0 34080.0 104680.0 ;
      RECT  33375.0 106025.0 34080.0 104680.0 ;
      RECT  33375.0 106025.0 34080.0 107370.0 ;
      RECT  33375.0 108715.0 34080.0 107370.0 ;
      RECT  33375.0 108715.0 34080.0 110060.0 ;
      RECT  33375.0 111405.0 34080.0 110060.0 ;
      RECT  33375.0 111405.0 34080.0 112750.0 ;
      RECT  33375.0 114095.0 34080.0 112750.0 ;
      RECT  34080.0 28015.0 34785.0 29360.0 ;
      RECT  34080.0 30705.0 34785.0 29360.0 ;
      RECT  34080.0 30705.0 34785.0 32050.0 ;
      RECT  34080.0 33395.0 34785.0 32050.0 ;
      RECT  34080.0 33395.0 34785.0 34740.0 ;
      RECT  34080.0 36085.0 34785.0 34740.0 ;
      RECT  34080.0 36085.0 34785.0 37430.0 ;
      RECT  34080.0 38775.0 34785.0 37430.0 ;
      RECT  34080.0 38775.0 34785.0 40120.0 ;
      RECT  34080.0 41465.0 34785.0 40120.0 ;
      RECT  34080.0 41465.0 34785.0 42810.0 ;
      RECT  34080.0 44155.0 34785.0 42810.0 ;
      RECT  34080.0 44155.0 34785.0 45500.0 ;
      RECT  34080.0 46845.0 34785.0 45500.0 ;
      RECT  34080.0 46845.0 34785.0 48190.0 ;
      RECT  34080.0 49535.0 34785.0 48190.0 ;
      RECT  34080.0 49535.0 34785.0 50880.0 ;
      RECT  34080.0 52225.0 34785.0 50880.0 ;
      RECT  34080.0 52225.0 34785.0 53570.0 ;
      RECT  34080.0 54915.0 34785.0 53570.0 ;
      RECT  34080.0 54915.0 34785.0 56260.0 ;
      RECT  34080.0 57605.0 34785.0 56260.0 ;
      RECT  34080.0 57605.0 34785.0 58950.0 ;
      RECT  34080.0 60295.0 34785.0 58950.0 ;
      RECT  34080.0 60295.0 34785.0 61640.0 ;
      RECT  34080.0 62985.0 34785.0 61640.0 ;
      RECT  34080.0 62985.0 34785.0 64330.0 ;
      RECT  34080.0 65675.0 34785.0 64330.0 ;
      RECT  34080.0 65675.0 34785.0 67020.0 ;
      RECT  34080.0 68365.0 34785.0 67020.0 ;
      RECT  34080.0 68365.0 34785.0 69710.0 ;
      RECT  34080.0 71055.0 34785.0 69710.0 ;
      RECT  34080.0 71055.0 34785.0 72400.0 ;
      RECT  34080.0 73745.0 34785.0 72400.0 ;
      RECT  34080.0 73745.0 34785.0 75090.0 ;
      RECT  34080.0 76435.0 34785.0 75090.0 ;
      RECT  34080.0 76435.0 34785.0 77780.0 ;
      RECT  34080.0 79125.0 34785.0 77780.0 ;
      RECT  34080.0 79125.0 34785.0 80470.0 ;
      RECT  34080.0 81815.0 34785.0 80470.0 ;
      RECT  34080.0 81815.0 34785.0 83160.0 ;
      RECT  34080.0 84505.0 34785.0 83160.0 ;
      RECT  34080.0 84505.0 34785.0 85850.0 ;
      RECT  34080.0 87195.0 34785.0 85850.0 ;
      RECT  34080.0 87195.0 34785.0 88540.0 ;
      RECT  34080.0 89885.0 34785.0 88540.0 ;
      RECT  34080.0 89885.0 34785.0 91230.0 ;
      RECT  34080.0 92575.0 34785.0 91230.0 ;
      RECT  34080.0 92575.0 34785.0 93920.0 ;
      RECT  34080.0 95265.0 34785.0 93920.0 ;
      RECT  34080.0 95265.0 34785.0 96610.0 ;
      RECT  34080.0 97955.0 34785.0 96610.0 ;
      RECT  34080.0 97955.0 34785.0 99300.0 ;
      RECT  34080.0 100645.0 34785.0 99300.0 ;
      RECT  34080.0 100645.0 34785.0 101990.0 ;
      RECT  34080.0 103335.0 34785.0 101990.0 ;
      RECT  34080.0 103335.0 34785.0 104680.0 ;
      RECT  34080.0 106025.0 34785.0 104680.0 ;
      RECT  34080.0 106025.0 34785.0 107370.0 ;
      RECT  34080.0 108715.0 34785.0 107370.0 ;
      RECT  34080.0 108715.0 34785.0 110060.0 ;
      RECT  34080.0 111405.0 34785.0 110060.0 ;
      RECT  34080.0 111405.0 34785.0 112750.0 ;
      RECT  34080.0 114095.0 34785.0 112750.0 ;
      RECT  34785.0 28015.0 35490.0 29360.0 ;
      RECT  34785.0 30705.0 35490.0 29360.0 ;
      RECT  34785.0 30705.0 35490.0 32050.0 ;
      RECT  34785.0 33395.0 35490.0 32050.0 ;
      RECT  34785.0 33395.0 35490.0 34740.0 ;
      RECT  34785.0 36085.0 35490.0 34740.0 ;
      RECT  34785.0 36085.0 35490.0 37430.0 ;
      RECT  34785.0 38775.0 35490.0 37430.0 ;
      RECT  34785.0 38775.0 35490.0 40120.0 ;
      RECT  34785.0 41465.0 35490.0 40120.0 ;
      RECT  34785.0 41465.0 35490.0 42810.0 ;
      RECT  34785.0 44155.0 35490.0 42810.0 ;
      RECT  34785.0 44155.0 35490.0 45500.0 ;
      RECT  34785.0 46845.0 35490.0 45500.0 ;
      RECT  34785.0 46845.0 35490.0 48190.0 ;
      RECT  34785.0 49535.0 35490.0 48190.0 ;
      RECT  34785.0 49535.0 35490.0 50880.0 ;
      RECT  34785.0 52225.0 35490.0 50880.0 ;
      RECT  34785.0 52225.0 35490.0 53570.0 ;
      RECT  34785.0 54915.0 35490.0 53570.0 ;
      RECT  34785.0 54915.0 35490.0 56260.0 ;
      RECT  34785.0 57605.0 35490.0 56260.0 ;
      RECT  34785.0 57605.0 35490.0 58950.0 ;
      RECT  34785.0 60295.0 35490.0 58950.0 ;
      RECT  34785.0 60295.0 35490.0 61640.0 ;
      RECT  34785.0 62985.0 35490.0 61640.0 ;
      RECT  34785.0 62985.0 35490.0 64330.0 ;
      RECT  34785.0 65675.0 35490.0 64330.0 ;
      RECT  34785.0 65675.0 35490.0 67020.0 ;
      RECT  34785.0 68365.0 35490.0 67020.0 ;
      RECT  34785.0 68365.0 35490.0 69710.0 ;
      RECT  34785.0 71055.0 35490.0 69710.0 ;
      RECT  34785.0 71055.0 35490.0 72400.0 ;
      RECT  34785.0 73745.0 35490.0 72400.0 ;
      RECT  34785.0 73745.0 35490.0 75090.0 ;
      RECT  34785.0 76435.0 35490.0 75090.0 ;
      RECT  34785.0 76435.0 35490.0 77780.0 ;
      RECT  34785.0 79125.0 35490.0 77780.0 ;
      RECT  34785.0 79125.0 35490.0 80470.0 ;
      RECT  34785.0 81815.0 35490.0 80470.0 ;
      RECT  34785.0 81815.0 35490.0 83160.0 ;
      RECT  34785.0 84505.0 35490.0 83160.0 ;
      RECT  34785.0 84505.0 35490.0 85850.0 ;
      RECT  34785.0 87195.0 35490.0 85850.0 ;
      RECT  34785.0 87195.0 35490.0 88540.0 ;
      RECT  34785.0 89885.0 35490.0 88540.0 ;
      RECT  34785.0 89885.0 35490.0 91230.0 ;
      RECT  34785.0 92575.0 35490.0 91230.0 ;
      RECT  34785.0 92575.0 35490.0 93920.0 ;
      RECT  34785.0 95265.0 35490.0 93920.0 ;
      RECT  34785.0 95265.0 35490.0 96610.0 ;
      RECT  34785.0 97955.0 35490.0 96610.0 ;
      RECT  34785.0 97955.0 35490.0 99300.0 ;
      RECT  34785.0 100645.0 35490.0 99300.0 ;
      RECT  34785.0 100645.0 35490.0 101990.0 ;
      RECT  34785.0 103335.0 35490.0 101990.0 ;
      RECT  34785.0 103335.0 35490.0 104680.0 ;
      RECT  34785.0 106025.0 35490.0 104680.0 ;
      RECT  34785.0 106025.0 35490.0 107370.0 ;
      RECT  34785.0 108715.0 35490.0 107370.0 ;
      RECT  34785.0 108715.0 35490.0 110060.0 ;
      RECT  34785.0 111405.0 35490.0 110060.0 ;
      RECT  34785.0 111405.0 35490.0 112750.0 ;
      RECT  34785.0 114095.0 35490.0 112750.0 ;
      RECT  35490.0 28015.0 36195.0 29360.0 ;
      RECT  35490.0 30705.0 36195.0 29360.0 ;
      RECT  35490.0 30705.0 36195.0 32050.0 ;
      RECT  35490.0 33395.0 36195.0 32050.0 ;
      RECT  35490.0 33395.0 36195.0 34740.0 ;
      RECT  35490.0 36085.0 36195.0 34740.0 ;
      RECT  35490.0 36085.0 36195.0 37430.0 ;
      RECT  35490.0 38775.0 36195.0 37430.0 ;
      RECT  35490.0 38775.0 36195.0 40120.0 ;
      RECT  35490.0 41465.0 36195.0 40120.0 ;
      RECT  35490.0 41465.0 36195.0 42810.0 ;
      RECT  35490.0 44155.0 36195.0 42810.0 ;
      RECT  35490.0 44155.0 36195.0 45500.0 ;
      RECT  35490.0 46845.0 36195.0 45500.0 ;
      RECT  35490.0 46845.0 36195.0 48190.0 ;
      RECT  35490.0 49535.0 36195.0 48190.0 ;
      RECT  35490.0 49535.0 36195.0 50880.0 ;
      RECT  35490.0 52225.0 36195.0 50880.0 ;
      RECT  35490.0 52225.0 36195.0 53570.0 ;
      RECT  35490.0 54915.0 36195.0 53570.0 ;
      RECT  35490.0 54915.0 36195.0 56260.0 ;
      RECT  35490.0 57605.0 36195.0 56260.0 ;
      RECT  35490.0 57605.0 36195.0 58950.0 ;
      RECT  35490.0 60295.0 36195.0 58950.0 ;
      RECT  35490.0 60295.0 36195.0 61640.0 ;
      RECT  35490.0 62985.0 36195.0 61640.0 ;
      RECT  35490.0 62985.0 36195.0 64330.0 ;
      RECT  35490.0 65675.0 36195.0 64330.0 ;
      RECT  35490.0 65675.0 36195.0 67020.0 ;
      RECT  35490.0 68365.0 36195.0 67020.0 ;
      RECT  35490.0 68365.0 36195.0 69710.0 ;
      RECT  35490.0 71055.0 36195.0 69710.0 ;
      RECT  35490.0 71055.0 36195.0 72400.0 ;
      RECT  35490.0 73745.0 36195.0 72400.0 ;
      RECT  35490.0 73745.0 36195.0 75090.0 ;
      RECT  35490.0 76435.0 36195.0 75090.0 ;
      RECT  35490.0 76435.0 36195.0 77780.0 ;
      RECT  35490.0 79125.0 36195.0 77780.0 ;
      RECT  35490.0 79125.0 36195.0 80470.0 ;
      RECT  35490.0 81815.0 36195.0 80470.0 ;
      RECT  35490.0 81815.0 36195.0 83160.0 ;
      RECT  35490.0 84505.0 36195.0 83160.0 ;
      RECT  35490.0 84505.0 36195.0 85850.0 ;
      RECT  35490.0 87195.0 36195.0 85850.0 ;
      RECT  35490.0 87195.0 36195.0 88540.0 ;
      RECT  35490.0 89885.0 36195.0 88540.0 ;
      RECT  35490.0 89885.0 36195.0 91230.0 ;
      RECT  35490.0 92575.0 36195.0 91230.0 ;
      RECT  35490.0 92575.0 36195.0 93920.0 ;
      RECT  35490.0 95265.0 36195.0 93920.0 ;
      RECT  35490.0 95265.0 36195.0 96610.0 ;
      RECT  35490.0 97955.0 36195.0 96610.0 ;
      RECT  35490.0 97955.0 36195.0 99300.0 ;
      RECT  35490.0 100645.0 36195.0 99300.0 ;
      RECT  35490.0 100645.0 36195.0 101990.0 ;
      RECT  35490.0 103335.0 36195.0 101990.0 ;
      RECT  35490.0 103335.0 36195.0 104680.0 ;
      RECT  35490.0 106025.0 36195.0 104680.0 ;
      RECT  35490.0 106025.0 36195.0 107370.0 ;
      RECT  35490.0 108715.0 36195.0 107370.0 ;
      RECT  35490.0 108715.0 36195.0 110060.0 ;
      RECT  35490.0 111405.0 36195.0 110060.0 ;
      RECT  35490.0 111405.0 36195.0 112750.0 ;
      RECT  35490.0 114095.0 36195.0 112750.0 ;
      RECT  36195.0 28015.0 36900.0 29360.0 ;
      RECT  36195.0 30705.0 36900.0 29360.0 ;
      RECT  36195.0 30705.0 36900.0 32050.0 ;
      RECT  36195.0 33395.0 36900.0 32050.0 ;
      RECT  36195.0 33395.0 36900.0 34740.0 ;
      RECT  36195.0 36085.0 36900.0 34740.0 ;
      RECT  36195.0 36085.0 36900.0 37430.0 ;
      RECT  36195.0 38775.0 36900.0 37430.0 ;
      RECT  36195.0 38775.0 36900.0 40120.0 ;
      RECT  36195.0 41465.0 36900.0 40120.0 ;
      RECT  36195.0 41465.0 36900.0 42810.0 ;
      RECT  36195.0 44155.0 36900.0 42810.0 ;
      RECT  36195.0 44155.0 36900.0 45500.0 ;
      RECT  36195.0 46845.0 36900.0 45500.0 ;
      RECT  36195.0 46845.0 36900.0 48190.0 ;
      RECT  36195.0 49535.0 36900.0 48190.0 ;
      RECT  36195.0 49535.0 36900.0 50880.0 ;
      RECT  36195.0 52225.0 36900.0 50880.0 ;
      RECT  36195.0 52225.0 36900.0 53570.0 ;
      RECT  36195.0 54915.0 36900.0 53570.0 ;
      RECT  36195.0 54915.0 36900.0 56260.0 ;
      RECT  36195.0 57605.0 36900.0 56260.0 ;
      RECT  36195.0 57605.0 36900.0 58950.0 ;
      RECT  36195.0 60295.0 36900.0 58950.0 ;
      RECT  36195.0 60295.0 36900.0 61640.0 ;
      RECT  36195.0 62985.0 36900.0 61640.0 ;
      RECT  36195.0 62985.0 36900.0 64330.0 ;
      RECT  36195.0 65675.0 36900.0 64330.0 ;
      RECT  36195.0 65675.0 36900.0 67020.0 ;
      RECT  36195.0 68365.0 36900.0 67020.0 ;
      RECT  36195.0 68365.0 36900.0 69710.0 ;
      RECT  36195.0 71055.0 36900.0 69710.0 ;
      RECT  36195.0 71055.0 36900.0 72400.0 ;
      RECT  36195.0 73745.0 36900.0 72400.0 ;
      RECT  36195.0 73745.0 36900.0 75090.0 ;
      RECT  36195.0 76435.0 36900.0 75090.0 ;
      RECT  36195.0 76435.0 36900.0 77780.0 ;
      RECT  36195.0 79125.0 36900.0 77780.0 ;
      RECT  36195.0 79125.0 36900.0 80470.0 ;
      RECT  36195.0 81815.0 36900.0 80470.0 ;
      RECT  36195.0 81815.0 36900.0 83160.0 ;
      RECT  36195.0 84505.0 36900.0 83160.0 ;
      RECT  36195.0 84505.0 36900.0 85850.0 ;
      RECT  36195.0 87195.0 36900.0 85850.0 ;
      RECT  36195.0 87195.0 36900.0 88540.0 ;
      RECT  36195.0 89885.0 36900.0 88540.0 ;
      RECT  36195.0 89885.0 36900.0 91230.0 ;
      RECT  36195.0 92575.0 36900.0 91230.0 ;
      RECT  36195.0 92575.0 36900.0 93920.0 ;
      RECT  36195.0 95265.0 36900.0 93920.0 ;
      RECT  36195.0 95265.0 36900.0 96610.0 ;
      RECT  36195.0 97955.0 36900.0 96610.0 ;
      RECT  36195.0 97955.0 36900.0 99300.0 ;
      RECT  36195.0 100645.0 36900.0 99300.0 ;
      RECT  36195.0 100645.0 36900.0 101990.0 ;
      RECT  36195.0 103335.0 36900.0 101990.0 ;
      RECT  36195.0 103335.0 36900.0 104680.0 ;
      RECT  36195.0 106025.0 36900.0 104680.0 ;
      RECT  36195.0 106025.0 36900.0 107370.0 ;
      RECT  36195.0 108715.0 36900.0 107370.0 ;
      RECT  36195.0 108715.0 36900.0 110060.0 ;
      RECT  36195.0 111405.0 36900.0 110060.0 ;
      RECT  36195.0 111405.0 36900.0 112750.0 ;
      RECT  36195.0 114095.0 36900.0 112750.0 ;
      RECT  36900.0 28015.0 37605.0 29360.0 ;
      RECT  36900.0 30705.0 37605.0 29360.0 ;
      RECT  36900.0 30705.0 37605.0 32050.0 ;
      RECT  36900.0 33395.0 37605.0 32050.0 ;
      RECT  36900.0 33395.0 37605.0 34740.0 ;
      RECT  36900.0 36085.0 37605.0 34740.0 ;
      RECT  36900.0 36085.0 37605.0 37430.0 ;
      RECT  36900.0 38775.0 37605.0 37430.0 ;
      RECT  36900.0 38775.0 37605.0 40120.0 ;
      RECT  36900.0 41465.0 37605.0 40120.0 ;
      RECT  36900.0 41465.0 37605.0 42810.0 ;
      RECT  36900.0 44155.0 37605.0 42810.0 ;
      RECT  36900.0 44155.0 37605.0 45500.0 ;
      RECT  36900.0 46845.0 37605.0 45500.0 ;
      RECT  36900.0 46845.0 37605.0 48190.0 ;
      RECT  36900.0 49535.0 37605.0 48190.0 ;
      RECT  36900.0 49535.0 37605.0 50880.0 ;
      RECT  36900.0 52225.0 37605.0 50880.0 ;
      RECT  36900.0 52225.0 37605.0 53570.0 ;
      RECT  36900.0 54915.0 37605.0 53570.0 ;
      RECT  36900.0 54915.0 37605.0 56260.0 ;
      RECT  36900.0 57605.0 37605.0 56260.0 ;
      RECT  36900.0 57605.0 37605.0 58950.0 ;
      RECT  36900.0 60295.0 37605.0 58950.0 ;
      RECT  36900.0 60295.0 37605.0 61640.0 ;
      RECT  36900.0 62985.0 37605.0 61640.0 ;
      RECT  36900.0 62985.0 37605.0 64330.0 ;
      RECT  36900.0 65675.0 37605.0 64330.0 ;
      RECT  36900.0 65675.0 37605.0 67020.0 ;
      RECT  36900.0 68365.0 37605.0 67020.0 ;
      RECT  36900.0 68365.0 37605.0 69710.0 ;
      RECT  36900.0 71055.0 37605.0 69710.0 ;
      RECT  36900.0 71055.0 37605.0 72400.0 ;
      RECT  36900.0 73745.0 37605.0 72400.0 ;
      RECT  36900.0 73745.0 37605.0 75090.0 ;
      RECT  36900.0 76435.0 37605.0 75090.0 ;
      RECT  36900.0 76435.0 37605.0 77780.0 ;
      RECT  36900.0 79125.0 37605.0 77780.0 ;
      RECT  36900.0 79125.0 37605.0 80470.0 ;
      RECT  36900.0 81815.0 37605.0 80470.0 ;
      RECT  36900.0 81815.0 37605.0 83160.0 ;
      RECT  36900.0 84505.0 37605.0 83160.0 ;
      RECT  36900.0 84505.0 37605.0 85850.0 ;
      RECT  36900.0 87195.0 37605.0 85850.0 ;
      RECT  36900.0 87195.0 37605.0 88540.0 ;
      RECT  36900.0 89885.0 37605.0 88540.0 ;
      RECT  36900.0 89885.0 37605.0 91230.0 ;
      RECT  36900.0 92575.0 37605.0 91230.0 ;
      RECT  36900.0 92575.0 37605.0 93920.0 ;
      RECT  36900.0 95265.0 37605.0 93920.0 ;
      RECT  36900.0 95265.0 37605.0 96610.0 ;
      RECT  36900.0 97955.0 37605.0 96610.0 ;
      RECT  36900.0 97955.0 37605.0 99300.0 ;
      RECT  36900.0 100645.0 37605.0 99300.0 ;
      RECT  36900.0 100645.0 37605.0 101990.0 ;
      RECT  36900.0 103335.0 37605.0 101990.0 ;
      RECT  36900.0 103335.0 37605.0 104680.0 ;
      RECT  36900.0 106025.0 37605.0 104680.0 ;
      RECT  36900.0 106025.0 37605.0 107370.0 ;
      RECT  36900.0 108715.0 37605.0 107370.0 ;
      RECT  36900.0 108715.0 37605.0 110060.0 ;
      RECT  36900.0 111405.0 37605.0 110060.0 ;
      RECT  36900.0 111405.0 37605.0 112750.0 ;
      RECT  36900.0 114095.0 37605.0 112750.0 ;
      RECT  37605.0 28015.0 38310.0 29360.0 ;
      RECT  37605.0 30705.0 38310.0 29360.0 ;
      RECT  37605.0 30705.0 38310.0 32050.0 ;
      RECT  37605.0 33395.0 38310.0 32050.0 ;
      RECT  37605.0 33395.0 38310.0 34740.0 ;
      RECT  37605.0 36085.0 38310.0 34740.0 ;
      RECT  37605.0 36085.0 38310.0 37430.0 ;
      RECT  37605.0 38775.0 38310.0 37430.0 ;
      RECT  37605.0 38775.0 38310.0 40120.0 ;
      RECT  37605.0 41465.0 38310.0 40120.0 ;
      RECT  37605.0 41465.0 38310.0 42810.0 ;
      RECT  37605.0 44155.0 38310.0 42810.0 ;
      RECT  37605.0 44155.0 38310.0 45500.0 ;
      RECT  37605.0 46845.0 38310.0 45500.0 ;
      RECT  37605.0 46845.0 38310.0 48190.0 ;
      RECT  37605.0 49535.0 38310.0 48190.0 ;
      RECT  37605.0 49535.0 38310.0 50880.0 ;
      RECT  37605.0 52225.0 38310.0 50880.0 ;
      RECT  37605.0 52225.0 38310.0 53570.0 ;
      RECT  37605.0 54915.0 38310.0 53570.0 ;
      RECT  37605.0 54915.0 38310.0 56260.0 ;
      RECT  37605.0 57605.0 38310.0 56260.0 ;
      RECT  37605.0 57605.0 38310.0 58950.0 ;
      RECT  37605.0 60295.0 38310.0 58950.0 ;
      RECT  37605.0 60295.0 38310.0 61640.0 ;
      RECT  37605.0 62985.0 38310.0 61640.0 ;
      RECT  37605.0 62985.0 38310.0 64330.0 ;
      RECT  37605.0 65675.0 38310.0 64330.0 ;
      RECT  37605.0 65675.0 38310.0 67020.0 ;
      RECT  37605.0 68365.0 38310.0 67020.0 ;
      RECT  37605.0 68365.0 38310.0 69710.0 ;
      RECT  37605.0 71055.0 38310.0 69710.0 ;
      RECT  37605.0 71055.0 38310.0 72400.0 ;
      RECT  37605.0 73745.0 38310.0 72400.0 ;
      RECT  37605.0 73745.0 38310.0 75090.0 ;
      RECT  37605.0 76435.0 38310.0 75090.0 ;
      RECT  37605.0 76435.0 38310.0 77780.0 ;
      RECT  37605.0 79125.0 38310.0 77780.0 ;
      RECT  37605.0 79125.0 38310.0 80470.0 ;
      RECT  37605.0 81815.0 38310.0 80470.0 ;
      RECT  37605.0 81815.0 38310.0 83160.0 ;
      RECT  37605.0 84505.0 38310.0 83160.0 ;
      RECT  37605.0 84505.0 38310.0 85850.0 ;
      RECT  37605.0 87195.0 38310.0 85850.0 ;
      RECT  37605.0 87195.0 38310.0 88540.0 ;
      RECT  37605.0 89885.0 38310.0 88540.0 ;
      RECT  37605.0 89885.0 38310.0 91230.0 ;
      RECT  37605.0 92575.0 38310.0 91230.0 ;
      RECT  37605.0 92575.0 38310.0 93920.0 ;
      RECT  37605.0 95265.0 38310.0 93920.0 ;
      RECT  37605.0 95265.0 38310.0 96610.0 ;
      RECT  37605.0 97955.0 38310.0 96610.0 ;
      RECT  37605.0 97955.0 38310.0 99300.0 ;
      RECT  37605.0 100645.0 38310.0 99300.0 ;
      RECT  37605.0 100645.0 38310.0 101990.0 ;
      RECT  37605.0 103335.0 38310.0 101990.0 ;
      RECT  37605.0 103335.0 38310.0 104680.0 ;
      RECT  37605.0 106025.0 38310.0 104680.0 ;
      RECT  37605.0 106025.0 38310.0 107370.0 ;
      RECT  37605.0 108715.0 38310.0 107370.0 ;
      RECT  37605.0 108715.0 38310.0 110060.0 ;
      RECT  37605.0 111405.0 38310.0 110060.0 ;
      RECT  37605.0 111405.0 38310.0 112750.0 ;
      RECT  37605.0 114095.0 38310.0 112750.0 ;
      RECT  38310.0 28015.0 39015.0 29360.0 ;
      RECT  38310.0 30705.0 39015.0 29360.0 ;
      RECT  38310.0 30705.0 39015.0 32050.0 ;
      RECT  38310.0 33395.0 39015.0 32050.0 ;
      RECT  38310.0 33395.0 39015.0 34740.0 ;
      RECT  38310.0 36085.0 39015.0 34740.0 ;
      RECT  38310.0 36085.0 39015.0 37430.0 ;
      RECT  38310.0 38775.0 39015.0 37430.0 ;
      RECT  38310.0 38775.0 39015.0 40120.0 ;
      RECT  38310.0 41465.0 39015.0 40120.0 ;
      RECT  38310.0 41465.0 39015.0 42810.0 ;
      RECT  38310.0 44155.0 39015.0 42810.0 ;
      RECT  38310.0 44155.0 39015.0 45500.0 ;
      RECT  38310.0 46845.0 39015.0 45500.0 ;
      RECT  38310.0 46845.0 39015.0 48190.0 ;
      RECT  38310.0 49535.0 39015.0 48190.0 ;
      RECT  38310.0 49535.0 39015.0 50880.0 ;
      RECT  38310.0 52225.0 39015.0 50880.0 ;
      RECT  38310.0 52225.0 39015.0 53570.0 ;
      RECT  38310.0 54915.0 39015.0 53570.0 ;
      RECT  38310.0 54915.0 39015.0 56260.0 ;
      RECT  38310.0 57605.0 39015.0 56260.0 ;
      RECT  38310.0 57605.0 39015.0 58950.0 ;
      RECT  38310.0 60295.0 39015.0 58950.0 ;
      RECT  38310.0 60295.0 39015.0 61640.0 ;
      RECT  38310.0 62985.0 39015.0 61640.0 ;
      RECT  38310.0 62985.0 39015.0 64330.0 ;
      RECT  38310.0 65675.0 39015.0 64330.0 ;
      RECT  38310.0 65675.0 39015.0 67020.0 ;
      RECT  38310.0 68365.0 39015.0 67020.0 ;
      RECT  38310.0 68365.0 39015.0 69710.0 ;
      RECT  38310.0 71055.0 39015.0 69710.0 ;
      RECT  38310.0 71055.0 39015.0 72400.0 ;
      RECT  38310.0 73745.0 39015.0 72400.0 ;
      RECT  38310.0 73745.0 39015.0 75090.0 ;
      RECT  38310.0 76435.0 39015.0 75090.0 ;
      RECT  38310.0 76435.0 39015.0 77780.0 ;
      RECT  38310.0 79125.0 39015.0 77780.0 ;
      RECT  38310.0 79125.0 39015.0 80470.0 ;
      RECT  38310.0 81815.0 39015.0 80470.0 ;
      RECT  38310.0 81815.0 39015.0 83160.0 ;
      RECT  38310.0 84505.0 39015.0 83160.0 ;
      RECT  38310.0 84505.0 39015.0 85850.0 ;
      RECT  38310.0 87195.0 39015.0 85850.0 ;
      RECT  38310.0 87195.0 39015.0 88540.0 ;
      RECT  38310.0 89885.0 39015.0 88540.0 ;
      RECT  38310.0 89885.0 39015.0 91230.0 ;
      RECT  38310.0 92575.0 39015.0 91230.0 ;
      RECT  38310.0 92575.0 39015.0 93920.0 ;
      RECT  38310.0 95265.0 39015.0 93920.0 ;
      RECT  38310.0 95265.0 39015.0 96610.0 ;
      RECT  38310.0 97955.0 39015.0 96610.0 ;
      RECT  38310.0 97955.0 39015.0 99300.0 ;
      RECT  38310.0 100645.0 39015.0 99300.0 ;
      RECT  38310.0 100645.0 39015.0 101990.0 ;
      RECT  38310.0 103335.0 39015.0 101990.0 ;
      RECT  38310.0 103335.0 39015.0 104680.0 ;
      RECT  38310.0 106025.0 39015.0 104680.0 ;
      RECT  38310.0 106025.0 39015.0 107370.0 ;
      RECT  38310.0 108715.0 39015.0 107370.0 ;
      RECT  38310.0 108715.0 39015.0 110060.0 ;
      RECT  38310.0 111405.0 39015.0 110060.0 ;
      RECT  38310.0 111405.0 39015.0 112750.0 ;
      RECT  38310.0 114095.0 39015.0 112750.0 ;
      RECT  39015.0 28015.0 39720.0 29360.0 ;
      RECT  39015.0 30705.0 39720.0 29360.0 ;
      RECT  39015.0 30705.0 39720.0 32050.0 ;
      RECT  39015.0 33395.0 39720.0 32050.0 ;
      RECT  39015.0 33395.0 39720.0 34740.0 ;
      RECT  39015.0 36085.0 39720.0 34740.0 ;
      RECT  39015.0 36085.0 39720.0 37430.0 ;
      RECT  39015.0 38775.0 39720.0 37430.0 ;
      RECT  39015.0 38775.0 39720.0 40120.0 ;
      RECT  39015.0 41465.0 39720.0 40120.0 ;
      RECT  39015.0 41465.0 39720.0 42810.0 ;
      RECT  39015.0 44155.0 39720.0 42810.0 ;
      RECT  39015.0 44155.0 39720.0 45500.0 ;
      RECT  39015.0 46845.0 39720.0 45500.0 ;
      RECT  39015.0 46845.0 39720.0 48190.0 ;
      RECT  39015.0 49535.0 39720.0 48190.0 ;
      RECT  39015.0 49535.0 39720.0 50880.0 ;
      RECT  39015.0 52225.0 39720.0 50880.0 ;
      RECT  39015.0 52225.0 39720.0 53570.0 ;
      RECT  39015.0 54915.0 39720.0 53570.0 ;
      RECT  39015.0 54915.0 39720.0 56260.0 ;
      RECT  39015.0 57605.0 39720.0 56260.0 ;
      RECT  39015.0 57605.0 39720.0 58950.0 ;
      RECT  39015.0 60295.0 39720.0 58950.0 ;
      RECT  39015.0 60295.0 39720.0 61640.0 ;
      RECT  39015.0 62985.0 39720.0 61640.0 ;
      RECT  39015.0 62985.0 39720.0 64330.0 ;
      RECT  39015.0 65675.0 39720.0 64330.0 ;
      RECT  39015.0 65675.0 39720.0 67020.0 ;
      RECT  39015.0 68365.0 39720.0 67020.0 ;
      RECT  39015.0 68365.0 39720.0 69710.0 ;
      RECT  39015.0 71055.0 39720.0 69710.0 ;
      RECT  39015.0 71055.0 39720.0 72400.0 ;
      RECT  39015.0 73745.0 39720.0 72400.0 ;
      RECT  39015.0 73745.0 39720.0 75090.0 ;
      RECT  39015.0 76435.0 39720.0 75090.0 ;
      RECT  39015.0 76435.0 39720.0 77780.0 ;
      RECT  39015.0 79125.0 39720.0 77780.0 ;
      RECT  39015.0 79125.0 39720.0 80470.0 ;
      RECT  39015.0 81815.0 39720.0 80470.0 ;
      RECT  39015.0 81815.0 39720.0 83160.0 ;
      RECT  39015.0 84505.0 39720.0 83160.0 ;
      RECT  39015.0 84505.0 39720.0 85850.0 ;
      RECT  39015.0 87195.0 39720.0 85850.0 ;
      RECT  39015.0 87195.0 39720.0 88540.0 ;
      RECT  39015.0 89885.0 39720.0 88540.0 ;
      RECT  39015.0 89885.0 39720.0 91230.0 ;
      RECT  39015.0 92575.0 39720.0 91230.0 ;
      RECT  39015.0 92575.0 39720.0 93920.0 ;
      RECT  39015.0 95265.0 39720.0 93920.0 ;
      RECT  39015.0 95265.0 39720.0 96610.0 ;
      RECT  39015.0 97955.0 39720.0 96610.0 ;
      RECT  39015.0 97955.0 39720.0 99300.0 ;
      RECT  39015.0 100645.0 39720.0 99300.0 ;
      RECT  39015.0 100645.0 39720.0 101990.0 ;
      RECT  39015.0 103335.0 39720.0 101990.0 ;
      RECT  39015.0 103335.0 39720.0 104680.0 ;
      RECT  39015.0 106025.0 39720.0 104680.0 ;
      RECT  39015.0 106025.0 39720.0 107370.0 ;
      RECT  39015.0 108715.0 39720.0 107370.0 ;
      RECT  39015.0 108715.0 39720.0 110060.0 ;
      RECT  39015.0 111405.0 39720.0 110060.0 ;
      RECT  39015.0 111405.0 39720.0 112750.0 ;
      RECT  39015.0 114095.0 39720.0 112750.0 ;
      RECT  39720.0 28015.0 40425.0 29360.0 ;
      RECT  39720.0 30705.0 40425.0 29360.0 ;
      RECT  39720.0 30705.0 40425.0 32050.0 ;
      RECT  39720.0 33395.0 40425.0 32050.0 ;
      RECT  39720.0 33395.0 40425.0 34740.0 ;
      RECT  39720.0 36085.0 40425.0 34740.0 ;
      RECT  39720.0 36085.0 40425.0 37430.0 ;
      RECT  39720.0 38775.0 40425.0 37430.0 ;
      RECT  39720.0 38775.0 40425.0 40120.0 ;
      RECT  39720.0 41465.0 40425.0 40120.0 ;
      RECT  39720.0 41465.0 40425.0 42810.0 ;
      RECT  39720.0 44155.0 40425.0 42810.0 ;
      RECT  39720.0 44155.0 40425.0 45500.0 ;
      RECT  39720.0 46845.0 40425.0 45500.0 ;
      RECT  39720.0 46845.0 40425.0 48190.0 ;
      RECT  39720.0 49535.0 40425.0 48190.0 ;
      RECT  39720.0 49535.0 40425.0 50880.0 ;
      RECT  39720.0 52225.0 40425.0 50880.0 ;
      RECT  39720.0 52225.0 40425.0 53570.0 ;
      RECT  39720.0 54915.0 40425.0 53570.0 ;
      RECT  39720.0 54915.0 40425.0 56260.0 ;
      RECT  39720.0 57605.0 40425.0 56260.0 ;
      RECT  39720.0 57605.0 40425.0 58950.0 ;
      RECT  39720.0 60295.0 40425.0 58950.0 ;
      RECT  39720.0 60295.0 40425.0 61640.0 ;
      RECT  39720.0 62985.0 40425.0 61640.0 ;
      RECT  39720.0 62985.0 40425.0 64330.0 ;
      RECT  39720.0 65675.0 40425.0 64330.0 ;
      RECT  39720.0 65675.0 40425.0 67020.0 ;
      RECT  39720.0 68365.0 40425.0 67020.0 ;
      RECT  39720.0 68365.0 40425.0 69710.0 ;
      RECT  39720.0 71055.0 40425.0 69710.0 ;
      RECT  39720.0 71055.0 40425.0 72400.0 ;
      RECT  39720.0 73745.0 40425.0 72400.0 ;
      RECT  39720.0 73745.0 40425.0 75090.0 ;
      RECT  39720.0 76435.0 40425.0 75090.0 ;
      RECT  39720.0 76435.0 40425.0 77780.0 ;
      RECT  39720.0 79125.0 40425.0 77780.0 ;
      RECT  39720.0 79125.0 40425.0 80470.0 ;
      RECT  39720.0 81815.0 40425.0 80470.0 ;
      RECT  39720.0 81815.0 40425.0 83160.0 ;
      RECT  39720.0 84505.0 40425.0 83160.0 ;
      RECT  39720.0 84505.0 40425.0 85850.0 ;
      RECT  39720.0 87195.0 40425.0 85850.0 ;
      RECT  39720.0 87195.0 40425.0 88540.0 ;
      RECT  39720.0 89885.0 40425.0 88540.0 ;
      RECT  39720.0 89885.0 40425.0 91230.0 ;
      RECT  39720.0 92575.0 40425.0 91230.0 ;
      RECT  39720.0 92575.0 40425.0 93920.0 ;
      RECT  39720.0 95265.0 40425.0 93920.0 ;
      RECT  39720.0 95265.0 40425.0 96610.0 ;
      RECT  39720.0 97955.0 40425.0 96610.0 ;
      RECT  39720.0 97955.0 40425.0 99300.0 ;
      RECT  39720.0 100645.0 40425.0 99300.0 ;
      RECT  39720.0 100645.0 40425.0 101990.0 ;
      RECT  39720.0 103335.0 40425.0 101990.0 ;
      RECT  39720.0 103335.0 40425.0 104680.0 ;
      RECT  39720.0 106025.0 40425.0 104680.0 ;
      RECT  39720.0 106025.0 40425.0 107370.0 ;
      RECT  39720.0 108715.0 40425.0 107370.0 ;
      RECT  39720.0 108715.0 40425.0 110060.0 ;
      RECT  39720.0 111405.0 40425.0 110060.0 ;
      RECT  39720.0 111405.0 40425.0 112750.0 ;
      RECT  39720.0 114095.0 40425.0 112750.0 ;
      RECT  40425.0 28015.0 41130.0 29360.0 ;
      RECT  40425.0 30705.0 41130.0 29360.0 ;
      RECT  40425.0 30705.0 41130.0 32050.0 ;
      RECT  40425.0 33395.0 41130.0 32050.0 ;
      RECT  40425.0 33395.0 41130.0 34740.0 ;
      RECT  40425.0 36085.0 41130.0 34740.0 ;
      RECT  40425.0 36085.0 41130.0 37430.0 ;
      RECT  40425.0 38775.0 41130.0 37430.0 ;
      RECT  40425.0 38775.0 41130.0 40120.0 ;
      RECT  40425.0 41465.0 41130.0 40120.0 ;
      RECT  40425.0 41465.0 41130.0 42810.0 ;
      RECT  40425.0 44155.0 41130.0 42810.0 ;
      RECT  40425.0 44155.0 41130.0 45500.0 ;
      RECT  40425.0 46845.0 41130.0 45500.0 ;
      RECT  40425.0 46845.0 41130.0 48190.0 ;
      RECT  40425.0 49535.0 41130.0 48190.0 ;
      RECT  40425.0 49535.0 41130.0 50880.0 ;
      RECT  40425.0 52225.0 41130.0 50880.0 ;
      RECT  40425.0 52225.0 41130.0 53570.0 ;
      RECT  40425.0 54915.0 41130.0 53570.0 ;
      RECT  40425.0 54915.0 41130.0 56260.0 ;
      RECT  40425.0 57605.0 41130.0 56260.0 ;
      RECT  40425.0 57605.0 41130.0 58950.0 ;
      RECT  40425.0 60295.0 41130.0 58950.0 ;
      RECT  40425.0 60295.0 41130.0 61640.0 ;
      RECT  40425.0 62985.0 41130.0 61640.0 ;
      RECT  40425.0 62985.0 41130.0 64330.0 ;
      RECT  40425.0 65675.0 41130.0 64330.0 ;
      RECT  40425.0 65675.0 41130.0 67020.0 ;
      RECT  40425.0 68365.0 41130.0 67020.0 ;
      RECT  40425.0 68365.0 41130.0 69710.0 ;
      RECT  40425.0 71055.0 41130.0 69710.0 ;
      RECT  40425.0 71055.0 41130.0 72400.0 ;
      RECT  40425.0 73745.0 41130.0 72400.0 ;
      RECT  40425.0 73745.0 41130.0 75090.0 ;
      RECT  40425.0 76435.0 41130.0 75090.0 ;
      RECT  40425.0 76435.0 41130.0 77780.0 ;
      RECT  40425.0 79125.0 41130.0 77780.0 ;
      RECT  40425.0 79125.0 41130.0 80470.0 ;
      RECT  40425.0 81815.0 41130.0 80470.0 ;
      RECT  40425.0 81815.0 41130.0 83160.0 ;
      RECT  40425.0 84505.0 41130.0 83160.0 ;
      RECT  40425.0 84505.0 41130.0 85850.0 ;
      RECT  40425.0 87195.0 41130.0 85850.0 ;
      RECT  40425.0 87195.0 41130.0 88540.0 ;
      RECT  40425.0 89885.0 41130.0 88540.0 ;
      RECT  40425.0 89885.0 41130.0 91230.0 ;
      RECT  40425.0 92575.0 41130.0 91230.0 ;
      RECT  40425.0 92575.0 41130.0 93920.0 ;
      RECT  40425.0 95265.0 41130.0 93920.0 ;
      RECT  40425.0 95265.0 41130.0 96610.0 ;
      RECT  40425.0 97955.0 41130.0 96610.0 ;
      RECT  40425.0 97955.0 41130.0 99300.0 ;
      RECT  40425.0 100645.0 41130.0 99300.0 ;
      RECT  40425.0 100645.0 41130.0 101990.0 ;
      RECT  40425.0 103335.0 41130.0 101990.0 ;
      RECT  40425.0 103335.0 41130.0 104680.0 ;
      RECT  40425.0 106025.0 41130.0 104680.0 ;
      RECT  40425.0 106025.0 41130.0 107370.0 ;
      RECT  40425.0 108715.0 41130.0 107370.0 ;
      RECT  40425.0 108715.0 41130.0 110060.0 ;
      RECT  40425.0 111405.0 41130.0 110060.0 ;
      RECT  40425.0 111405.0 41130.0 112750.0 ;
      RECT  40425.0 114095.0 41130.0 112750.0 ;
      RECT  41130.0 28015.0 41835.0 29360.0 ;
      RECT  41130.0 30705.0 41835.0 29360.0 ;
      RECT  41130.0 30705.0 41835.0 32050.0 ;
      RECT  41130.0 33395.0 41835.0 32050.0 ;
      RECT  41130.0 33395.0 41835.0 34740.0 ;
      RECT  41130.0 36085.0 41835.0 34740.0 ;
      RECT  41130.0 36085.0 41835.0 37430.0 ;
      RECT  41130.0 38775.0 41835.0 37430.0 ;
      RECT  41130.0 38775.0 41835.0 40120.0 ;
      RECT  41130.0 41465.0 41835.0 40120.0 ;
      RECT  41130.0 41465.0 41835.0 42810.0 ;
      RECT  41130.0 44155.0 41835.0 42810.0 ;
      RECT  41130.0 44155.0 41835.0 45500.0 ;
      RECT  41130.0 46845.0 41835.0 45500.0 ;
      RECT  41130.0 46845.0 41835.0 48190.0 ;
      RECT  41130.0 49535.0 41835.0 48190.0 ;
      RECT  41130.0 49535.0 41835.0 50880.0 ;
      RECT  41130.0 52225.0 41835.0 50880.0 ;
      RECT  41130.0 52225.0 41835.0 53570.0 ;
      RECT  41130.0 54915.0 41835.0 53570.0 ;
      RECT  41130.0 54915.0 41835.0 56260.0 ;
      RECT  41130.0 57605.0 41835.0 56260.0 ;
      RECT  41130.0 57605.0 41835.0 58950.0 ;
      RECT  41130.0 60295.0 41835.0 58950.0 ;
      RECT  41130.0 60295.0 41835.0 61640.0 ;
      RECT  41130.0 62985.0 41835.0 61640.0 ;
      RECT  41130.0 62985.0 41835.0 64330.0 ;
      RECT  41130.0 65675.0 41835.0 64330.0 ;
      RECT  41130.0 65675.0 41835.0 67020.0 ;
      RECT  41130.0 68365.0 41835.0 67020.0 ;
      RECT  41130.0 68365.0 41835.0 69710.0 ;
      RECT  41130.0 71055.0 41835.0 69710.0 ;
      RECT  41130.0 71055.0 41835.0 72400.0 ;
      RECT  41130.0 73745.0 41835.0 72400.0 ;
      RECT  41130.0 73745.0 41835.0 75090.0 ;
      RECT  41130.0 76435.0 41835.0 75090.0 ;
      RECT  41130.0 76435.0 41835.0 77780.0 ;
      RECT  41130.0 79125.0 41835.0 77780.0 ;
      RECT  41130.0 79125.0 41835.0 80470.0 ;
      RECT  41130.0 81815.0 41835.0 80470.0 ;
      RECT  41130.0 81815.0 41835.0 83160.0 ;
      RECT  41130.0 84505.0 41835.0 83160.0 ;
      RECT  41130.0 84505.0 41835.0 85850.0 ;
      RECT  41130.0 87195.0 41835.0 85850.0 ;
      RECT  41130.0 87195.0 41835.0 88540.0 ;
      RECT  41130.0 89885.0 41835.0 88540.0 ;
      RECT  41130.0 89885.0 41835.0 91230.0 ;
      RECT  41130.0 92575.0 41835.0 91230.0 ;
      RECT  41130.0 92575.0 41835.0 93920.0 ;
      RECT  41130.0 95265.0 41835.0 93920.0 ;
      RECT  41130.0 95265.0 41835.0 96610.0 ;
      RECT  41130.0 97955.0 41835.0 96610.0 ;
      RECT  41130.0 97955.0 41835.0 99300.0 ;
      RECT  41130.0 100645.0 41835.0 99300.0 ;
      RECT  41130.0 100645.0 41835.0 101990.0 ;
      RECT  41130.0 103335.0 41835.0 101990.0 ;
      RECT  41130.0 103335.0 41835.0 104680.0 ;
      RECT  41130.0 106025.0 41835.0 104680.0 ;
      RECT  41130.0 106025.0 41835.0 107370.0 ;
      RECT  41130.0 108715.0 41835.0 107370.0 ;
      RECT  41130.0 108715.0 41835.0 110060.0 ;
      RECT  41130.0 111405.0 41835.0 110060.0 ;
      RECT  41130.0 111405.0 41835.0 112750.0 ;
      RECT  41130.0 114095.0 41835.0 112750.0 ;
      RECT  41835.0 28015.0 42540.0 29360.0 ;
      RECT  41835.0 30705.0 42540.0 29360.0 ;
      RECT  41835.0 30705.0 42540.0 32050.0 ;
      RECT  41835.0 33395.0 42540.0 32050.0 ;
      RECT  41835.0 33395.0 42540.0 34740.0 ;
      RECT  41835.0 36085.0 42540.0 34740.0 ;
      RECT  41835.0 36085.0 42540.0 37430.0 ;
      RECT  41835.0 38775.0 42540.0 37430.0 ;
      RECT  41835.0 38775.0 42540.0 40120.0 ;
      RECT  41835.0 41465.0 42540.0 40120.0 ;
      RECT  41835.0 41465.0 42540.0 42810.0 ;
      RECT  41835.0 44155.0 42540.0 42810.0 ;
      RECT  41835.0 44155.0 42540.0 45500.0 ;
      RECT  41835.0 46845.0 42540.0 45500.0 ;
      RECT  41835.0 46845.0 42540.0 48190.0 ;
      RECT  41835.0 49535.0 42540.0 48190.0 ;
      RECT  41835.0 49535.0 42540.0 50880.0 ;
      RECT  41835.0 52225.0 42540.0 50880.0 ;
      RECT  41835.0 52225.0 42540.0 53570.0 ;
      RECT  41835.0 54915.0 42540.0 53570.0 ;
      RECT  41835.0 54915.0 42540.0 56260.0 ;
      RECT  41835.0 57605.0 42540.0 56260.0 ;
      RECT  41835.0 57605.0 42540.0 58950.0 ;
      RECT  41835.0 60295.0 42540.0 58950.0 ;
      RECT  41835.0 60295.0 42540.0 61640.0 ;
      RECT  41835.0 62985.0 42540.0 61640.0 ;
      RECT  41835.0 62985.0 42540.0 64330.0 ;
      RECT  41835.0 65675.0 42540.0 64330.0 ;
      RECT  41835.0 65675.0 42540.0 67020.0 ;
      RECT  41835.0 68365.0 42540.0 67020.0 ;
      RECT  41835.0 68365.0 42540.0 69710.0 ;
      RECT  41835.0 71055.0 42540.0 69710.0 ;
      RECT  41835.0 71055.0 42540.0 72400.0 ;
      RECT  41835.0 73745.0 42540.0 72400.0 ;
      RECT  41835.0 73745.0 42540.0 75090.0 ;
      RECT  41835.0 76435.0 42540.0 75090.0 ;
      RECT  41835.0 76435.0 42540.0 77780.0 ;
      RECT  41835.0 79125.0 42540.0 77780.0 ;
      RECT  41835.0 79125.0 42540.0 80470.0 ;
      RECT  41835.0 81815.0 42540.0 80470.0 ;
      RECT  41835.0 81815.0 42540.0 83160.0 ;
      RECT  41835.0 84505.0 42540.0 83160.0 ;
      RECT  41835.0 84505.0 42540.0 85850.0 ;
      RECT  41835.0 87195.0 42540.0 85850.0 ;
      RECT  41835.0 87195.0 42540.0 88540.0 ;
      RECT  41835.0 89885.0 42540.0 88540.0 ;
      RECT  41835.0 89885.0 42540.0 91230.0 ;
      RECT  41835.0 92575.0 42540.0 91230.0 ;
      RECT  41835.0 92575.0 42540.0 93920.0 ;
      RECT  41835.0 95265.0 42540.0 93920.0 ;
      RECT  41835.0 95265.0 42540.0 96610.0 ;
      RECT  41835.0 97955.0 42540.0 96610.0 ;
      RECT  41835.0 97955.0 42540.0 99300.0 ;
      RECT  41835.0 100645.0 42540.0 99300.0 ;
      RECT  41835.0 100645.0 42540.0 101990.0 ;
      RECT  41835.0 103335.0 42540.0 101990.0 ;
      RECT  41835.0 103335.0 42540.0 104680.0 ;
      RECT  41835.0 106025.0 42540.0 104680.0 ;
      RECT  41835.0 106025.0 42540.0 107370.0 ;
      RECT  41835.0 108715.0 42540.0 107370.0 ;
      RECT  41835.0 108715.0 42540.0 110060.0 ;
      RECT  41835.0 111405.0 42540.0 110060.0 ;
      RECT  41835.0 111405.0 42540.0 112750.0 ;
      RECT  41835.0 114095.0 42540.0 112750.0 ;
      RECT  42540.0 28015.0 43245.0 29360.0 ;
      RECT  42540.0 30705.0 43245.0 29360.0 ;
      RECT  42540.0 30705.0 43245.0 32050.0 ;
      RECT  42540.0 33395.0 43245.0 32050.0 ;
      RECT  42540.0 33395.0 43245.0 34740.0 ;
      RECT  42540.0 36085.0 43245.0 34740.0 ;
      RECT  42540.0 36085.0 43245.0 37430.0 ;
      RECT  42540.0 38775.0 43245.0 37430.0 ;
      RECT  42540.0 38775.0 43245.0 40120.0 ;
      RECT  42540.0 41465.0 43245.0 40120.0 ;
      RECT  42540.0 41465.0 43245.0 42810.0 ;
      RECT  42540.0 44155.0 43245.0 42810.0 ;
      RECT  42540.0 44155.0 43245.0 45500.0 ;
      RECT  42540.0 46845.0 43245.0 45500.0 ;
      RECT  42540.0 46845.0 43245.0 48190.0 ;
      RECT  42540.0 49535.0 43245.0 48190.0 ;
      RECT  42540.0 49535.0 43245.0 50880.0 ;
      RECT  42540.0 52225.0 43245.0 50880.0 ;
      RECT  42540.0 52225.0 43245.0 53570.0 ;
      RECT  42540.0 54915.0 43245.0 53570.0 ;
      RECT  42540.0 54915.0 43245.0 56260.0 ;
      RECT  42540.0 57605.0 43245.0 56260.0 ;
      RECT  42540.0 57605.0 43245.0 58950.0 ;
      RECT  42540.0 60295.0 43245.0 58950.0 ;
      RECT  42540.0 60295.0 43245.0 61640.0 ;
      RECT  42540.0 62985.0 43245.0 61640.0 ;
      RECT  42540.0 62985.0 43245.0 64330.0 ;
      RECT  42540.0 65675.0 43245.0 64330.0 ;
      RECT  42540.0 65675.0 43245.0 67020.0 ;
      RECT  42540.0 68365.0 43245.0 67020.0 ;
      RECT  42540.0 68365.0 43245.0 69710.0 ;
      RECT  42540.0 71055.0 43245.0 69710.0 ;
      RECT  42540.0 71055.0 43245.0 72400.0 ;
      RECT  42540.0 73745.0 43245.0 72400.0 ;
      RECT  42540.0 73745.0 43245.0 75090.0 ;
      RECT  42540.0 76435.0 43245.0 75090.0 ;
      RECT  42540.0 76435.0 43245.0 77780.0 ;
      RECT  42540.0 79125.0 43245.0 77780.0 ;
      RECT  42540.0 79125.0 43245.0 80470.0 ;
      RECT  42540.0 81815.0 43245.0 80470.0 ;
      RECT  42540.0 81815.0 43245.0 83160.0 ;
      RECT  42540.0 84505.0 43245.0 83160.0 ;
      RECT  42540.0 84505.0 43245.0 85850.0 ;
      RECT  42540.0 87195.0 43245.0 85850.0 ;
      RECT  42540.0 87195.0 43245.0 88540.0 ;
      RECT  42540.0 89885.0 43245.0 88540.0 ;
      RECT  42540.0 89885.0 43245.0 91230.0 ;
      RECT  42540.0 92575.0 43245.0 91230.0 ;
      RECT  42540.0 92575.0 43245.0 93920.0 ;
      RECT  42540.0 95265.0 43245.0 93920.0 ;
      RECT  42540.0 95265.0 43245.0 96610.0 ;
      RECT  42540.0 97955.0 43245.0 96610.0 ;
      RECT  42540.0 97955.0 43245.0 99300.0 ;
      RECT  42540.0 100645.0 43245.0 99300.0 ;
      RECT  42540.0 100645.0 43245.0 101990.0 ;
      RECT  42540.0 103335.0 43245.0 101990.0 ;
      RECT  42540.0 103335.0 43245.0 104680.0 ;
      RECT  42540.0 106025.0 43245.0 104680.0 ;
      RECT  42540.0 106025.0 43245.0 107370.0 ;
      RECT  42540.0 108715.0 43245.0 107370.0 ;
      RECT  42540.0 108715.0 43245.0 110060.0 ;
      RECT  42540.0 111405.0 43245.0 110060.0 ;
      RECT  42540.0 111405.0 43245.0 112750.0 ;
      RECT  42540.0 114095.0 43245.0 112750.0 ;
      RECT  43245.0 28015.0 43950.0 29360.0 ;
      RECT  43245.0 30705.0 43950.0 29360.0 ;
      RECT  43245.0 30705.0 43950.0 32050.0 ;
      RECT  43245.0 33395.0 43950.0 32050.0 ;
      RECT  43245.0 33395.0 43950.0 34740.0 ;
      RECT  43245.0 36085.0 43950.0 34740.0 ;
      RECT  43245.0 36085.0 43950.0 37430.0 ;
      RECT  43245.0 38775.0 43950.0 37430.0 ;
      RECT  43245.0 38775.0 43950.0 40120.0 ;
      RECT  43245.0 41465.0 43950.0 40120.0 ;
      RECT  43245.0 41465.0 43950.0 42810.0 ;
      RECT  43245.0 44155.0 43950.0 42810.0 ;
      RECT  43245.0 44155.0 43950.0 45500.0 ;
      RECT  43245.0 46845.0 43950.0 45500.0 ;
      RECT  43245.0 46845.0 43950.0 48190.0 ;
      RECT  43245.0 49535.0 43950.0 48190.0 ;
      RECT  43245.0 49535.0 43950.0 50880.0 ;
      RECT  43245.0 52225.0 43950.0 50880.0 ;
      RECT  43245.0 52225.0 43950.0 53570.0 ;
      RECT  43245.0 54915.0 43950.0 53570.0 ;
      RECT  43245.0 54915.0 43950.0 56260.0 ;
      RECT  43245.0 57605.0 43950.0 56260.0 ;
      RECT  43245.0 57605.0 43950.0 58950.0 ;
      RECT  43245.0 60295.0 43950.0 58950.0 ;
      RECT  43245.0 60295.0 43950.0 61640.0 ;
      RECT  43245.0 62985.0 43950.0 61640.0 ;
      RECT  43245.0 62985.0 43950.0 64330.0 ;
      RECT  43245.0 65675.0 43950.0 64330.0 ;
      RECT  43245.0 65675.0 43950.0 67020.0 ;
      RECT  43245.0 68365.0 43950.0 67020.0 ;
      RECT  43245.0 68365.0 43950.0 69710.0 ;
      RECT  43245.0 71055.0 43950.0 69710.0 ;
      RECT  43245.0 71055.0 43950.0 72400.0 ;
      RECT  43245.0 73745.0 43950.0 72400.0 ;
      RECT  43245.0 73745.0 43950.0 75090.0 ;
      RECT  43245.0 76435.0 43950.0 75090.0 ;
      RECT  43245.0 76435.0 43950.0 77780.0 ;
      RECT  43245.0 79125.0 43950.0 77780.0 ;
      RECT  43245.0 79125.0 43950.0 80470.0 ;
      RECT  43245.0 81815.0 43950.0 80470.0 ;
      RECT  43245.0 81815.0 43950.0 83160.0 ;
      RECT  43245.0 84505.0 43950.0 83160.0 ;
      RECT  43245.0 84505.0 43950.0 85850.0 ;
      RECT  43245.0 87195.0 43950.0 85850.0 ;
      RECT  43245.0 87195.0 43950.0 88540.0 ;
      RECT  43245.0 89885.0 43950.0 88540.0 ;
      RECT  43245.0 89885.0 43950.0 91230.0 ;
      RECT  43245.0 92575.0 43950.0 91230.0 ;
      RECT  43245.0 92575.0 43950.0 93920.0 ;
      RECT  43245.0 95265.0 43950.0 93920.0 ;
      RECT  43245.0 95265.0 43950.0 96610.0 ;
      RECT  43245.0 97955.0 43950.0 96610.0 ;
      RECT  43245.0 97955.0 43950.0 99300.0 ;
      RECT  43245.0 100645.0 43950.0 99300.0 ;
      RECT  43245.0 100645.0 43950.0 101990.0 ;
      RECT  43245.0 103335.0 43950.0 101990.0 ;
      RECT  43245.0 103335.0 43950.0 104680.0 ;
      RECT  43245.0 106025.0 43950.0 104680.0 ;
      RECT  43245.0 106025.0 43950.0 107370.0 ;
      RECT  43245.0 108715.0 43950.0 107370.0 ;
      RECT  43245.0 108715.0 43950.0 110060.0 ;
      RECT  43245.0 111405.0 43950.0 110060.0 ;
      RECT  43245.0 111405.0 43950.0 112750.0 ;
      RECT  43245.0 114095.0 43950.0 112750.0 ;
      RECT  43950.0 28015.0 44655.0 29360.0 ;
      RECT  43950.0 30705.0 44655.0 29360.0 ;
      RECT  43950.0 30705.0 44655.0 32050.0 ;
      RECT  43950.0 33395.0 44655.0 32050.0 ;
      RECT  43950.0 33395.0 44655.0 34740.0 ;
      RECT  43950.0 36085.0 44655.0 34740.0 ;
      RECT  43950.0 36085.0 44655.0 37430.0 ;
      RECT  43950.0 38775.0 44655.0 37430.0 ;
      RECT  43950.0 38775.0 44655.0 40120.0 ;
      RECT  43950.0 41465.0 44655.0 40120.0 ;
      RECT  43950.0 41465.0 44655.0 42810.0 ;
      RECT  43950.0 44155.0 44655.0 42810.0 ;
      RECT  43950.0 44155.0 44655.0 45500.0 ;
      RECT  43950.0 46845.0 44655.0 45500.0 ;
      RECT  43950.0 46845.0 44655.0 48190.0 ;
      RECT  43950.0 49535.0 44655.0 48190.0 ;
      RECT  43950.0 49535.0 44655.0 50880.0 ;
      RECT  43950.0 52225.0 44655.0 50880.0 ;
      RECT  43950.0 52225.0 44655.0 53570.0 ;
      RECT  43950.0 54915.0 44655.0 53570.0 ;
      RECT  43950.0 54915.0 44655.0 56260.0 ;
      RECT  43950.0 57605.0 44655.0 56260.0 ;
      RECT  43950.0 57605.0 44655.0 58950.0 ;
      RECT  43950.0 60295.0 44655.0 58950.0 ;
      RECT  43950.0 60295.0 44655.0 61640.0 ;
      RECT  43950.0 62985.0 44655.0 61640.0 ;
      RECT  43950.0 62985.0 44655.0 64330.0 ;
      RECT  43950.0 65675.0 44655.0 64330.0 ;
      RECT  43950.0 65675.0 44655.0 67020.0 ;
      RECT  43950.0 68365.0 44655.0 67020.0 ;
      RECT  43950.0 68365.0 44655.0 69710.0 ;
      RECT  43950.0 71055.0 44655.0 69710.0 ;
      RECT  43950.0 71055.0 44655.0 72400.0 ;
      RECT  43950.0 73745.0 44655.0 72400.0 ;
      RECT  43950.0 73745.0 44655.0 75090.0 ;
      RECT  43950.0 76435.0 44655.0 75090.0 ;
      RECT  43950.0 76435.0 44655.0 77780.0 ;
      RECT  43950.0 79125.0 44655.0 77780.0 ;
      RECT  43950.0 79125.0 44655.0 80470.0 ;
      RECT  43950.0 81815.0 44655.0 80470.0 ;
      RECT  43950.0 81815.0 44655.0 83160.0 ;
      RECT  43950.0 84505.0 44655.0 83160.0 ;
      RECT  43950.0 84505.0 44655.0 85850.0 ;
      RECT  43950.0 87195.0 44655.0 85850.0 ;
      RECT  43950.0 87195.0 44655.0 88540.0 ;
      RECT  43950.0 89885.0 44655.0 88540.0 ;
      RECT  43950.0 89885.0 44655.0 91230.0 ;
      RECT  43950.0 92575.0 44655.0 91230.0 ;
      RECT  43950.0 92575.0 44655.0 93920.0 ;
      RECT  43950.0 95265.0 44655.0 93920.0 ;
      RECT  43950.0 95265.0 44655.0 96610.0 ;
      RECT  43950.0 97955.0 44655.0 96610.0 ;
      RECT  43950.0 97955.0 44655.0 99300.0 ;
      RECT  43950.0 100645.0 44655.0 99300.0 ;
      RECT  43950.0 100645.0 44655.0 101990.0 ;
      RECT  43950.0 103335.0 44655.0 101990.0 ;
      RECT  43950.0 103335.0 44655.0 104680.0 ;
      RECT  43950.0 106025.0 44655.0 104680.0 ;
      RECT  43950.0 106025.0 44655.0 107370.0 ;
      RECT  43950.0 108715.0 44655.0 107370.0 ;
      RECT  43950.0 108715.0 44655.0 110060.0 ;
      RECT  43950.0 111405.0 44655.0 110060.0 ;
      RECT  43950.0 111405.0 44655.0 112750.0 ;
      RECT  43950.0 114095.0 44655.0 112750.0 ;
      RECT  44655.0 28015.0 45360.0 29360.0 ;
      RECT  44655.0 30705.0 45360.0 29360.0 ;
      RECT  44655.0 30705.0 45360.0 32050.0 ;
      RECT  44655.0 33395.0 45360.0 32050.0 ;
      RECT  44655.0 33395.0 45360.0 34740.0 ;
      RECT  44655.0 36085.0 45360.0 34740.0 ;
      RECT  44655.0 36085.0 45360.0 37430.0 ;
      RECT  44655.0 38775.0 45360.0 37430.0 ;
      RECT  44655.0 38775.0 45360.0 40120.0 ;
      RECT  44655.0 41465.0 45360.0 40120.0 ;
      RECT  44655.0 41465.0 45360.0 42810.0 ;
      RECT  44655.0 44155.0 45360.0 42810.0 ;
      RECT  44655.0 44155.0 45360.0 45500.0 ;
      RECT  44655.0 46845.0 45360.0 45500.0 ;
      RECT  44655.0 46845.0 45360.0 48190.0 ;
      RECT  44655.0 49535.0 45360.0 48190.0 ;
      RECT  44655.0 49535.0 45360.0 50880.0 ;
      RECT  44655.0 52225.0 45360.0 50880.0 ;
      RECT  44655.0 52225.0 45360.0 53570.0 ;
      RECT  44655.0 54915.0 45360.0 53570.0 ;
      RECT  44655.0 54915.0 45360.0 56260.0 ;
      RECT  44655.0 57605.0 45360.0 56260.0 ;
      RECT  44655.0 57605.0 45360.0 58950.0 ;
      RECT  44655.0 60295.0 45360.0 58950.0 ;
      RECT  44655.0 60295.0 45360.0 61640.0 ;
      RECT  44655.0 62985.0 45360.0 61640.0 ;
      RECT  44655.0 62985.0 45360.0 64330.0 ;
      RECT  44655.0 65675.0 45360.0 64330.0 ;
      RECT  44655.0 65675.0 45360.0 67020.0 ;
      RECT  44655.0 68365.0 45360.0 67020.0 ;
      RECT  44655.0 68365.0 45360.0 69710.0 ;
      RECT  44655.0 71055.0 45360.0 69710.0 ;
      RECT  44655.0 71055.0 45360.0 72400.0 ;
      RECT  44655.0 73745.0 45360.0 72400.0 ;
      RECT  44655.0 73745.0 45360.0 75090.0 ;
      RECT  44655.0 76435.0 45360.0 75090.0 ;
      RECT  44655.0 76435.0 45360.0 77780.0 ;
      RECT  44655.0 79125.0 45360.0 77780.0 ;
      RECT  44655.0 79125.0 45360.0 80470.0 ;
      RECT  44655.0 81815.0 45360.0 80470.0 ;
      RECT  44655.0 81815.0 45360.0 83160.0 ;
      RECT  44655.0 84505.0 45360.0 83160.0 ;
      RECT  44655.0 84505.0 45360.0 85850.0 ;
      RECT  44655.0 87195.0 45360.0 85850.0 ;
      RECT  44655.0 87195.0 45360.0 88540.0 ;
      RECT  44655.0 89885.0 45360.0 88540.0 ;
      RECT  44655.0 89885.0 45360.0 91230.0 ;
      RECT  44655.0 92575.0 45360.0 91230.0 ;
      RECT  44655.0 92575.0 45360.0 93920.0 ;
      RECT  44655.0 95265.0 45360.0 93920.0 ;
      RECT  44655.0 95265.0 45360.0 96610.0 ;
      RECT  44655.0 97955.0 45360.0 96610.0 ;
      RECT  44655.0 97955.0 45360.0 99300.0 ;
      RECT  44655.0 100645.0 45360.0 99300.0 ;
      RECT  44655.0 100645.0 45360.0 101990.0 ;
      RECT  44655.0 103335.0 45360.0 101990.0 ;
      RECT  44655.0 103335.0 45360.0 104680.0 ;
      RECT  44655.0 106025.0 45360.0 104680.0 ;
      RECT  44655.0 106025.0 45360.0 107370.0 ;
      RECT  44655.0 108715.0 45360.0 107370.0 ;
      RECT  44655.0 108715.0 45360.0 110060.0 ;
      RECT  44655.0 111405.0 45360.0 110060.0 ;
      RECT  44655.0 111405.0 45360.0 112750.0 ;
      RECT  44655.0 114095.0 45360.0 112750.0 ;
      RECT  45360.0 28015.0 46065.0 29360.0 ;
      RECT  45360.0 30705.0 46065.0 29360.0 ;
      RECT  45360.0 30705.0 46065.0 32050.0 ;
      RECT  45360.0 33395.0 46065.0 32050.0 ;
      RECT  45360.0 33395.0 46065.0 34740.0 ;
      RECT  45360.0 36085.0 46065.0 34740.0 ;
      RECT  45360.0 36085.0 46065.0 37430.0 ;
      RECT  45360.0 38775.0 46065.0 37430.0 ;
      RECT  45360.0 38775.0 46065.0 40120.0 ;
      RECT  45360.0 41465.0 46065.0 40120.0 ;
      RECT  45360.0 41465.0 46065.0 42810.0 ;
      RECT  45360.0 44155.0 46065.0 42810.0 ;
      RECT  45360.0 44155.0 46065.0 45500.0 ;
      RECT  45360.0 46845.0 46065.0 45500.0 ;
      RECT  45360.0 46845.0 46065.0 48190.0 ;
      RECT  45360.0 49535.0 46065.0 48190.0 ;
      RECT  45360.0 49535.0 46065.0 50880.0 ;
      RECT  45360.0 52225.0 46065.0 50880.0 ;
      RECT  45360.0 52225.0 46065.0 53570.0 ;
      RECT  45360.0 54915.0 46065.0 53570.0 ;
      RECT  45360.0 54915.0 46065.0 56260.0 ;
      RECT  45360.0 57605.0 46065.0 56260.0 ;
      RECT  45360.0 57605.0 46065.0 58950.0 ;
      RECT  45360.0 60295.0 46065.0 58950.0 ;
      RECT  45360.0 60295.0 46065.0 61640.0 ;
      RECT  45360.0 62985.0 46065.0 61640.0 ;
      RECT  45360.0 62985.0 46065.0 64330.0 ;
      RECT  45360.0 65675.0 46065.0 64330.0 ;
      RECT  45360.0 65675.0 46065.0 67020.0 ;
      RECT  45360.0 68365.0 46065.0 67020.0 ;
      RECT  45360.0 68365.0 46065.0 69710.0 ;
      RECT  45360.0 71055.0 46065.0 69710.0 ;
      RECT  45360.0 71055.0 46065.0 72400.0 ;
      RECT  45360.0 73745.0 46065.0 72400.0 ;
      RECT  45360.0 73745.0 46065.0 75090.0 ;
      RECT  45360.0 76435.0 46065.0 75090.0 ;
      RECT  45360.0 76435.0 46065.0 77780.0 ;
      RECT  45360.0 79125.0 46065.0 77780.0 ;
      RECT  45360.0 79125.0 46065.0 80470.0 ;
      RECT  45360.0 81815.0 46065.0 80470.0 ;
      RECT  45360.0 81815.0 46065.0 83160.0 ;
      RECT  45360.0 84505.0 46065.0 83160.0 ;
      RECT  45360.0 84505.0 46065.0 85850.0 ;
      RECT  45360.0 87195.0 46065.0 85850.0 ;
      RECT  45360.0 87195.0 46065.0 88540.0 ;
      RECT  45360.0 89885.0 46065.0 88540.0 ;
      RECT  45360.0 89885.0 46065.0 91230.0 ;
      RECT  45360.0 92575.0 46065.0 91230.0 ;
      RECT  45360.0 92575.0 46065.0 93920.0 ;
      RECT  45360.0 95265.0 46065.0 93920.0 ;
      RECT  45360.0 95265.0 46065.0 96610.0 ;
      RECT  45360.0 97955.0 46065.0 96610.0 ;
      RECT  45360.0 97955.0 46065.0 99300.0 ;
      RECT  45360.0 100645.0 46065.0 99300.0 ;
      RECT  45360.0 100645.0 46065.0 101990.0 ;
      RECT  45360.0 103335.0 46065.0 101990.0 ;
      RECT  45360.0 103335.0 46065.0 104680.0 ;
      RECT  45360.0 106025.0 46065.0 104680.0 ;
      RECT  45360.0 106025.0 46065.0 107370.0 ;
      RECT  45360.0 108715.0 46065.0 107370.0 ;
      RECT  45360.0 108715.0 46065.0 110060.0 ;
      RECT  45360.0 111405.0 46065.0 110060.0 ;
      RECT  45360.0 111405.0 46065.0 112750.0 ;
      RECT  45360.0 114095.0 46065.0 112750.0 ;
      RECT  46065.0 28015.0 46770.0 29360.0 ;
      RECT  46065.0 30705.0 46770.0 29360.0 ;
      RECT  46065.0 30705.0 46770.0 32050.0 ;
      RECT  46065.0 33395.0 46770.0 32050.0 ;
      RECT  46065.0 33395.0 46770.0 34740.0 ;
      RECT  46065.0 36085.0 46770.0 34740.0 ;
      RECT  46065.0 36085.0 46770.0 37430.0 ;
      RECT  46065.0 38775.0 46770.0 37430.0 ;
      RECT  46065.0 38775.0 46770.0 40120.0 ;
      RECT  46065.0 41465.0 46770.0 40120.0 ;
      RECT  46065.0 41465.0 46770.0 42810.0 ;
      RECT  46065.0 44155.0 46770.0 42810.0 ;
      RECT  46065.0 44155.0 46770.0 45500.0 ;
      RECT  46065.0 46845.0 46770.0 45500.0 ;
      RECT  46065.0 46845.0 46770.0 48190.0 ;
      RECT  46065.0 49535.0 46770.0 48190.0 ;
      RECT  46065.0 49535.0 46770.0 50880.0 ;
      RECT  46065.0 52225.0 46770.0 50880.0 ;
      RECT  46065.0 52225.0 46770.0 53570.0 ;
      RECT  46065.0 54915.0 46770.0 53570.0 ;
      RECT  46065.0 54915.0 46770.0 56260.0 ;
      RECT  46065.0 57605.0 46770.0 56260.0 ;
      RECT  46065.0 57605.0 46770.0 58950.0 ;
      RECT  46065.0 60295.0 46770.0 58950.0 ;
      RECT  46065.0 60295.0 46770.0 61640.0 ;
      RECT  46065.0 62985.0 46770.0 61640.0 ;
      RECT  46065.0 62985.0 46770.0 64330.0 ;
      RECT  46065.0 65675.0 46770.0 64330.0 ;
      RECT  46065.0 65675.0 46770.0 67020.0 ;
      RECT  46065.0 68365.0 46770.0 67020.0 ;
      RECT  46065.0 68365.0 46770.0 69710.0 ;
      RECT  46065.0 71055.0 46770.0 69710.0 ;
      RECT  46065.0 71055.0 46770.0 72400.0 ;
      RECT  46065.0 73745.0 46770.0 72400.0 ;
      RECT  46065.0 73745.0 46770.0 75090.0 ;
      RECT  46065.0 76435.0 46770.0 75090.0 ;
      RECT  46065.0 76435.0 46770.0 77780.0 ;
      RECT  46065.0 79125.0 46770.0 77780.0 ;
      RECT  46065.0 79125.0 46770.0 80470.0 ;
      RECT  46065.0 81815.0 46770.0 80470.0 ;
      RECT  46065.0 81815.0 46770.0 83160.0 ;
      RECT  46065.0 84505.0 46770.0 83160.0 ;
      RECT  46065.0 84505.0 46770.0 85850.0 ;
      RECT  46065.0 87195.0 46770.0 85850.0 ;
      RECT  46065.0 87195.0 46770.0 88540.0 ;
      RECT  46065.0 89885.0 46770.0 88540.0 ;
      RECT  46065.0 89885.0 46770.0 91230.0 ;
      RECT  46065.0 92575.0 46770.0 91230.0 ;
      RECT  46065.0 92575.0 46770.0 93920.0 ;
      RECT  46065.0 95265.0 46770.0 93920.0 ;
      RECT  46065.0 95265.0 46770.0 96610.0 ;
      RECT  46065.0 97955.0 46770.0 96610.0 ;
      RECT  46065.0 97955.0 46770.0 99300.0 ;
      RECT  46065.0 100645.0 46770.0 99300.0 ;
      RECT  46065.0 100645.0 46770.0 101990.0 ;
      RECT  46065.0 103335.0 46770.0 101990.0 ;
      RECT  46065.0 103335.0 46770.0 104680.0 ;
      RECT  46065.0 106025.0 46770.0 104680.0 ;
      RECT  46065.0 106025.0 46770.0 107370.0 ;
      RECT  46065.0 108715.0 46770.0 107370.0 ;
      RECT  46065.0 108715.0 46770.0 110060.0 ;
      RECT  46065.0 111405.0 46770.0 110060.0 ;
      RECT  46065.0 111405.0 46770.0 112750.0 ;
      RECT  46065.0 114095.0 46770.0 112750.0 ;
      RECT  46770.0 28015.0 47475.0 29360.0 ;
      RECT  46770.0 30705.0 47475.0 29360.0 ;
      RECT  46770.0 30705.0 47475.0 32050.0 ;
      RECT  46770.0 33395.0 47475.0 32050.0 ;
      RECT  46770.0 33395.0 47475.0 34740.0 ;
      RECT  46770.0 36085.0 47475.0 34740.0 ;
      RECT  46770.0 36085.0 47475.0 37430.0 ;
      RECT  46770.0 38775.0 47475.0 37430.0 ;
      RECT  46770.0 38775.0 47475.0 40120.0 ;
      RECT  46770.0 41465.0 47475.0 40120.0 ;
      RECT  46770.0 41465.0 47475.0 42810.0 ;
      RECT  46770.0 44155.0 47475.0 42810.0 ;
      RECT  46770.0 44155.0 47475.0 45500.0 ;
      RECT  46770.0 46845.0 47475.0 45500.0 ;
      RECT  46770.0 46845.0 47475.0 48190.0 ;
      RECT  46770.0 49535.0 47475.0 48190.0 ;
      RECT  46770.0 49535.0 47475.0 50880.0 ;
      RECT  46770.0 52225.0 47475.0 50880.0 ;
      RECT  46770.0 52225.0 47475.0 53570.0 ;
      RECT  46770.0 54915.0 47475.0 53570.0 ;
      RECT  46770.0 54915.0 47475.0 56260.0 ;
      RECT  46770.0 57605.0 47475.0 56260.0 ;
      RECT  46770.0 57605.0 47475.0 58950.0 ;
      RECT  46770.0 60295.0 47475.0 58950.0 ;
      RECT  46770.0 60295.0 47475.0 61640.0 ;
      RECT  46770.0 62985.0 47475.0 61640.0 ;
      RECT  46770.0 62985.0 47475.0 64330.0 ;
      RECT  46770.0 65675.0 47475.0 64330.0 ;
      RECT  46770.0 65675.0 47475.0 67020.0 ;
      RECT  46770.0 68365.0 47475.0 67020.0 ;
      RECT  46770.0 68365.0 47475.0 69710.0 ;
      RECT  46770.0 71055.0 47475.0 69710.0 ;
      RECT  46770.0 71055.0 47475.0 72400.0 ;
      RECT  46770.0 73745.0 47475.0 72400.0 ;
      RECT  46770.0 73745.0 47475.0 75090.0 ;
      RECT  46770.0 76435.0 47475.0 75090.0 ;
      RECT  46770.0 76435.0 47475.0 77780.0 ;
      RECT  46770.0 79125.0 47475.0 77780.0 ;
      RECT  46770.0 79125.0 47475.0 80470.0 ;
      RECT  46770.0 81815.0 47475.0 80470.0 ;
      RECT  46770.0 81815.0 47475.0 83160.0 ;
      RECT  46770.0 84505.0 47475.0 83160.0 ;
      RECT  46770.0 84505.0 47475.0 85850.0 ;
      RECT  46770.0 87195.0 47475.0 85850.0 ;
      RECT  46770.0 87195.0 47475.0 88540.0 ;
      RECT  46770.0 89885.0 47475.0 88540.0 ;
      RECT  46770.0 89885.0 47475.0 91230.0 ;
      RECT  46770.0 92575.0 47475.0 91230.0 ;
      RECT  46770.0 92575.0 47475.0 93920.0 ;
      RECT  46770.0 95265.0 47475.0 93920.0 ;
      RECT  46770.0 95265.0 47475.0 96610.0 ;
      RECT  46770.0 97955.0 47475.0 96610.0 ;
      RECT  46770.0 97955.0 47475.0 99300.0 ;
      RECT  46770.0 100645.0 47475.0 99300.0 ;
      RECT  46770.0 100645.0 47475.0 101990.0 ;
      RECT  46770.0 103335.0 47475.0 101990.0 ;
      RECT  46770.0 103335.0 47475.0 104680.0 ;
      RECT  46770.0 106025.0 47475.0 104680.0 ;
      RECT  46770.0 106025.0 47475.0 107370.0 ;
      RECT  46770.0 108715.0 47475.0 107370.0 ;
      RECT  46770.0 108715.0 47475.0 110060.0 ;
      RECT  46770.0 111405.0 47475.0 110060.0 ;
      RECT  46770.0 111405.0 47475.0 112750.0 ;
      RECT  46770.0 114095.0 47475.0 112750.0 ;
      RECT  47475.0 28015.0 48180.0 29360.0 ;
      RECT  47475.0 30705.0 48180.0 29360.0 ;
      RECT  47475.0 30705.0 48180.0 32050.0 ;
      RECT  47475.0 33395.0 48180.0 32050.0 ;
      RECT  47475.0 33395.0 48180.0 34740.0 ;
      RECT  47475.0 36085.0 48180.0 34740.0 ;
      RECT  47475.0 36085.0 48180.0 37430.0 ;
      RECT  47475.0 38775.0 48180.0 37430.0 ;
      RECT  47475.0 38775.0 48180.0 40120.0 ;
      RECT  47475.0 41465.0 48180.0 40120.0 ;
      RECT  47475.0 41465.0 48180.0 42810.0 ;
      RECT  47475.0 44155.0 48180.0 42810.0 ;
      RECT  47475.0 44155.0 48180.0 45500.0 ;
      RECT  47475.0 46845.0 48180.0 45500.0 ;
      RECT  47475.0 46845.0 48180.0 48190.0 ;
      RECT  47475.0 49535.0 48180.0 48190.0 ;
      RECT  47475.0 49535.0 48180.0 50880.0 ;
      RECT  47475.0 52225.0 48180.0 50880.0 ;
      RECT  47475.0 52225.0 48180.0 53570.0 ;
      RECT  47475.0 54915.0 48180.0 53570.0 ;
      RECT  47475.0 54915.0 48180.0 56260.0 ;
      RECT  47475.0 57605.0 48180.0 56260.0 ;
      RECT  47475.0 57605.0 48180.0 58950.0 ;
      RECT  47475.0 60295.0 48180.0 58950.0 ;
      RECT  47475.0 60295.0 48180.0 61640.0 ;
      RECT  47475.0 62985.0 48180.0 61640.0 ;
      RECT  47475.0 62985.0 48180.0 64330.0 ;
      RECT  47475.0 65675.0 48180.0 64330.0 ;
      RECT  47475.0 65675.0 48180.0 67020.0 ;
      RECT  47475.0 68365.0 48180.0 67020.0 ;
      RECT  47475.0 68365.0 48180.0 69710.0 ;
      RECT  47475.0 71055.0 48180.0 69710.0 ;
      RECT  47475.0 71055.0 48180.0 72400.0 ;
      RECT  47475.0 73745.0 48180.0 72400.0 ;
      RECT  47475.0 73745.0 48180.0 75090.0 ;
      RECT  47475.0 76435.0 48180.0 75090.0 ;
      RECT  47475.0 76435.0 48180.0 77780.0 ;
      RECT  47475.0 79125.0 48180.0 77780.0 ;
      RECT  47475.0 79125.0 48180.0 80470.0 ;
      RECT  47475.0 81815.0 48180.0 80470.0 ;
      RECT  47475.0 81815.0 48180.0 83160.0 ;
      RECT  47475.0 84505.0 48180.0 83160.0 ;
      RECT  47475.0 84505.0 48180.0 85850.0 ;
      RECT  47475.0 87195.0 48180.0 85850.0 ;
      RECT  47475.0 87195.0 48180.0 88540.0 ;
      RECT  47475.0 89885.0 48180.0 88540.0 ;
      RECT  47475.0 89885.0 48180.0 91230.0 ;
      RECT  47475.0 92575.0 48180.0 91230.0 ;
      RECT  47475.0 92575.0 48180.0 93920.0 ;
      RECT  47475.0 95265.0 48180.0 93920.0 ;
      RECT  47475.0 95265.0 48180.0 96610.0 ;
      RECT  47475.0 97955.0 48180.0 96610.0 ;
      RECT  47475.0 97955.0 48180.0 99300.0 ;
      RECT  47475.0 100645.0 48180.0 99300.0 ;
      RECT  47475.0 100645.0 48180.0 101990.0 ;
      RECT  47475.0 103335.0 48180.0 101990.0 ;
      RECT  47475.0 103335.0 48180.0 104680.0 ;
      RECT  47475.0 106025.0 48180.0 104680.0 ;
      RECT  47475.0 106025.0 48180.0 107370.0 ;
      RECT  47475.0 108715.0 48180.0 107370.0 ;
      RECT  47475.0 108715.0 48180.0 110060.0 ;
      RECT  47475.0 111405.0 48180.0 110060.0 ;
      RECT  47475.0 111405.0 48180.0 112750.0 ;
      RECT  47475.0 114095.0 48180.0 112750.0 ;
      RECT  48180.0 28015.0 48885.0 29360.0 ;
      RECT  48180.0 30705.0 48885.0 29360.0 ;
      RECT  48180.0 30705.0 48885.0 32050.0 ;
      RECT  48180.0 33395.0 48885.0 32050.0 ;
      RECT  48180.0 33395.0 48885.0 34740.0 ;
      RECT  48180.0 36085.0 48885.0 34740.0 ;
      RECT  48180.0 36085.0 48885.0 37430.0 ;
      RECT  48180.0 38775.0 48885.0 37430.0 ;
      RECT  48180.0 38775.0 48885.0 40120.0 ;
      RECT  48180.0 41465.0 48885.0 40120.0 ;
      RECT  48180.0 41465.0 48885.0 42810.0 ;
      RECT  48180.0 44155.0 48885.0 42810.0 ;
      RECT  48180.0 44155.0 48885.0 45500.0 ;
      RECT  48180.0 46845.0 48885.0 45500.0 ;
      RECT  48180.0 46845.0 48885.0 48190.0 ;
      RECT  48180.0 49535.0 48885.0 48190.0 ;
      RECT  48180.0 49535.0 48885.0 50880.0 ;
      RECT  48180.0 52225.0 48885.0 50880.0 ;
      RECT  48180.0 52225.0 48885.0 53570.0 ;
      RECT  48180.0 54915.0 48885.0 53570.0 ;
      RECT  48180.0 54915.0 48885.0 56260.0 ;
      RECT  48180.0 57605.0 48885.0 56260.0 ;
      RECT  48180.0 57605.0 48885.0 58950.0 ;
      RECT  48180.0 60295.0 48885.0 58950.0 ;
      RECT  48180.0 60295.0 48885.0 61640.0 ;
      RECT  48180.0 62985.0 48885.0 61640.0 ;
      RECT  48180.0 62985.0 48885.0 64330.0 ;
      RECT  48180.0 65675.0 48885.0 64330.0 ;
      RECT  48180.0 65675.0 48885.0 67020.0 ;
      RECT  48180.0 68365.0 48885.0 67020.0 ;
      RECT  48180.0 68365.0 48885.0 69710.0 ;
      RECT  48180.0 71055.0 48885.0 69710.0 ;
      RECT  48180.0 71055.0 48885.0 72400.0 ;
      RECT  48180.0 73745.0 48885.0 72400.0 ;
      RECT  48180.0 73745.0 48885.0 75090.0 ;
      RECT  48180.0 76435.0 48885.0 75090.0 ;
      RECT  48180.0 76435.0 48885.0 77780.0 ;
      RECT  48180.0 79125.0 48885.0 77780.0 ;
      RECT  48180.0 79125.0 48885.0 80470.0 ;
      RECT  48180.0 81815.0 48885.0 80470.0 ;
      RECT  48180.0 81815.0 48885.0 83160.0 ;
      RECT  48180.0 84505.0 48885.0 83160.0 ;
      RECT  48180.0 84505.0 48885.0 85850.0 ;
      RECT  48180.0 87195.0 48885.0 85850.0 ;
      RECT  48180.0 87195.0 48885.0 88540.0 ;
      RECT  48180.0 89885.0 48885.0 88540.0 ;
      RECT  48180.0 89885.0 48885.0 91230.0 ;
      RECT  48180.0 92575.0 48885.0 91230.0 ;
      RECT  48180.0 92575.0 48885.0 93920.0 ;
      RECT  48180.0 95265.0 48885.0 93920.0 ;
      RECT  48180.0 95265.0 48885.0 96610.0 ;
      RECT  48180.0 97955.0 48885.0 96610.0 ;
      RECT  48180.0 97955.0 48885.0 99300.0 ;
      RECT  48180.0 100645.0 48885.0 99300.0 ;
      RECT  48180.0 100645.0 48885.0 101990.0 ;
      RECT  48180.0 103335.0 48885.0 101990.0 ;
      RECT  48180.0 103335.0 48885.0 104680.0 ;
      RECT  48180.0 106025.0 48885.0 104680.0 ;
      RECT  48180.0 106025.0 48885.0 107370.0 ;
      RECT  48180.0 108715.0 48885.0 107370.0 ;
      RECT  48180.0 108715.0 48885.0 110060.0 ;
      RECT  48180.0 111405.0 48885.0 110060.0 ;
      RECT  48180.0 111405.0 48885.0 112750.0 ;
      RECT  48180.0 114095.0 48885.0 112750.0 ;
      RECT  48885.0 28015.0 49590.0 29360.0 ;
      RECT  48885.0 30705.0 49590.0 29360.0 ;
      RECT  48885.0 30705.0 49590.0 32050.0 ;
      RECT  48885.0 33395.0 49590.0 32050.0 ;
      RECT  48885.0 33395.0 49590.0 34740.0 ;
      RECT  48885.0 36085.0 49590.0 34740.0 ;
      RECT  48885.0 36085.0 49590.0 37430.0 ;
      RECT  48885.0 38775.0 49590.0 37430.0 ;
      RECT  48885.0 38775.0 49590.0 40120.0 ;
      RECT  48885.0 41465.0 49590.0 40120.0 ;
      RECT  48885.0 41465.0 49590.0 42810.0 ;
      RECT  48885.0 44155.0 49590.0 42810.0 ;
      RECT  48885.0 44155.0 49590.0 45500.0 ;
      RECT  48885.0 46845.0 49590.0 45500.0 ;
      RECT  48885.0 46845.0 49590.0 48190.0 ;
      RECT  48885.0 49535.0 49590.0 48190.0 ;
      RECT  48885.0 49535.0 49590.0 50880.0 ;
      RECT  48885.0 52225.0 49590.0 50880.0 ;
      RECT  48885.0 52225.0 49590.0 53570.0 ;
      RECT  48885.0 54915.0 49590.0 53570.0 ;
      RECT  48885.0 54915.0 49590.0 56260.0 ;
      RECT  48885.0 57605.0 49590.0 56260.0 ;
      RECT  48885.0 57605.0 49590.0 58950.0 ;
      RECT  48885.0 60295.0 49590.0 58950.0 ;
      RECT  48885.0 60295.0 49590.0 61640.0 ;
      RECT  48885.0 62985.0 49590.0 61640.0 ;
      RECT  48885.0 62985.0 49590.0 64330.0 ;
      RECT  48885.0 65675.0 49590.0 64330.0 ;
      RECT  48885.0 65675.0 49590.0 67020.0 ;
      RECT  48885.0 68365.0 49590.0 67020.0 ;
      RECT  48885.0 68365.0 49590.0 69710.0 ;
      RECT  48885.0 71055.0 49590.0 69710.0 ;
      RECT  48885.0 71055.0 49590.0 72400.0 ;
      RECT  48885.0 73745.0 49590.0 72400.0 ;
      RECT  48885.0 73745.0 49590.0 75090.0 ;
      RECT  48885.0 76435.0 49590.0 75090.0 ;
      RECT  48885.0 76435.0 49590.0 77780.0 ;
      RECT  48885.0 79125.0 49590.0 77780.0 ;
      RECT  48885.0 79125.0 49590.0 80470.0 ;
      RECT  48885.0 81815.0 49590.0 80470.0 ;
      RECT  48885.0 81815.0 49590.0 83160.0 ;
      RECT  48885.0 84505.0 49590.0 83160.0 ;
      RECT  48885.0 84505.0 49590.0 85850.0 ;
      RECT  48885.0 87195.0 49590.0 85850.0 ;
      RECT  48885.0 87195.0 49590.0 88540.0 ;
      RECT  48885.0 89885.0 49590.0 88540.0 ;
      RECT  48885.0 89885.0 49590.0 91230.0 ;
      RECT  48885.0 92575.0 49590.0 91230.0 ;
      RECT  48885.0 92575.0 49590.0 93920.0 ;
      RECT  48885.0 95265.0 49590.0 93920.0 ;
      RECT  48885.0 95265.0 49590.0 96610.0 ;
      RECT  48885.0 97955.0 49590.0 96610.0 ;
      RECT  48885.0 97955.0 49590.0 99300.0 ;
      RECT  48885.0 100645.0 49590.0 99300.0 ;
      RECT  48885.0 100645.0 49590.0 101990.0 ;
      RECT  48885.0 103335.0 49590.0 101990.0 ;
      RECT  48885.0 103335.0 49590.0 104680.0 ;
      RECT  48885.0 106025.0 49590.0 104680.0 ;
      RECT  48885.0 106025.0 49590.0 107370.0 ;
      RECT  48885.0 108715.0 49590.0 107370.0 ;
      RECT  48885.0 108715.0 49590.0 110060.0 ;
      RECT  48885.0 111405.0 49590.0 110060.0 ;
      RECT  48885.0 111405.0 49590.0 112750.0 ;
      RECT  48885.0 114095.0 49590.0 112750.0 ;
      RECT  49590.0 28015.0 50295.0 29360.0 ;
      RECT  49590.0 30705.0 50295.0 29360.0 ;
      RECT  49590.0 30705.0 50295.0 32050.0 ;
      RECT  49590.0 33395.0 50295.0 32050.0 ;
      RECT  49590.0 33395.0 50295.0 34740.0 ;
      RECT  49590.0 36085.0 50295.0 34740.0 ;
      RECT  49590.0 36085.0 50295.0 37430.0 ;
      RECT  49590.0 38775.0 50295.0 37430.0 ;
      RECT  49590.0 38775.0 50295.0 40120.0 ;
      RECT  49590.0 41465.0 50295.0 40120.0 ;
      RECT  49590.0 41465.0 50295.0 42810.0 ;
      RECT  49590.0 44155.0 50295.0 42810.0 ;
      RECT  49590.0 44155.0 50295.0 45500.0 ;
      RECT  49590.0 46845.0 50295.0 45500.0 ;
      RECT  49590.0 46845.0 50295.0 48190.0 ;
      RECT  49590.0 49535.0 50295.0 48190.0 ;
      RECT  49590.0 49535.0 50295.0 50880.0 ;
      RECT  49590.0 52225.0 50295.0 50880.0 ;
      RECT  49590.0 52225.0 50295.0 53570.0 ;
      RECT  49590.0 54915.0 50295.0 53570.0 ;
      RECT  49590.0 54915.0 50295.0 56260.0 ;
      RECT  49590.0 57605.0 50295.0 56260.0 ;
      RECT  49590.0 57605.0 50295.0 58950.0 ;
      RECT  49590.0 60295.0 50295.0 58950.0 ;
      RECT  49590.0 60295.0 50295.0 61640.0 ;
      RECT  49590.0 62985.0 50295.0 61640.0 ;
      RECT  49590.0 62985.0 50295.0 64330.0 ;
      RECT  49590.0 65675.0 50295.0 64330.0 ;
      RECT  49590.0 65675.0 50295.0 67020.0 ;
      RECT  49590.0 68365.0 50295.0 67020.0 ;
      RECT  49590.0 68365.0 50295.0 69710.0 ;
      RECT  49590.0 71055.0 50295.0 69710.0 ;
      RECT  49590.0 71055.0 50295.0 72400.0 ;
      RECT  49590.0 73745.0 50295.0 72400.0 ;
      RECT  49590.0 73745.0 50295.0 75090.0 ;
      RECT  49590.0 76435.0 50295.0 75090.0 ;
      RECT  49590.0 76435.0 50295.0 77780.0 ;
      RECT  49590.0 79125.0 50295.0 77780.0 ;
      RECT  49590.0 79125.0 50295.0 80470.0 ;
      RECT  49590.0 81815.0 50295.0 80470.0 ;
      RECT  49590.0 81815.0 50295.0 83160.0 ;
      RECT  49590.0 84505.0 50295.0 83160.0 ;
      RECT  49590.0 84505.0 50295.0 85850.0 ;
      RECT  49590.0 87195.0 50295.0 85850.0 ;
      RECT  49590.0 87195.0 50295.0 88540.0 ;
      RECT  49590.0 89885.0 50295.0 88540.0 ;
      RECT  49590.0 89885.0 50295.0 91230.0 ;
      RECT  49590.0 92575.0 50295.0 91230.0 ;
      RECT  49590.0 92575.0 50295.0 93920.0 ;
      RECT  49590.0 95265.0 50295.0 93920.0 ;
      RECT  49590.0 95265.0 50295.0 96610.0 ;
      RECT  49590.0 97955.0 50295.0 96610.0 ;
      RECT  49590.0 97955.0 50295.0 99300.0 ;
      RECT  49590.0 100645.0 50295.0 99300.0 ;
      RECT  49590.0 100645.0 50295.0 101990.0 ;
      RECT  49590.0 103335.0 50295.0 101990.0 ;
      RECT  49590.0 103335.0 50295.0 104680.0 ;
      RECT  49590.0 106025.0 50295.0 104680.0 ;
      RECT  49590.0 106025.0 50295.0 107370.0 ;
      RECT  49590.0 108715.0 50295.0 107370.0 ;
      RECT  49590.0 108715.0 50295.0 110060.0 ;
      RECT  49590.0 111405.0 50295.0 110060.0 ;
      RECT  49590.0 111405.0 50295.0 112750.0 ;
      RECT  49590.0 114095.0 50295.0 112750.0 ;
      RECT  50295.0 28015.0 51000.0 29360.0 ;
      RECT  50295.0 30705.0 51000.0 29360.0 ;
      RECT  50295.0 30705.0 51000.0 32050.0 ;
      RECT  50295.0 33395.0 51000.0 32050.0 ;
      RECT  50295.0 33395.0 51000.0 34740.0 ;
      RECT  50295.0 36085.0 51000.0 34740.0 ;
      RECT  50295.0 36085.0 51000.0 37430.0 ;
      RECT  50295.0 38775.0 51000.0 37430.0 ;
      RECT  50295.0 38775.0 51000.0 40120.0 ;
      RECT  50295.0 41465.0 51000.0 40120.0 ;
      RECT  50295.0 41465.0 51000.0 42810.0 ;
      RECT  50295.0 44155.0 51000.0 42810.0 ;
      RECT  50295.0 44155.0 51000.0 45500.0 ;
      RECT  50295.0 46845.0 51000.0 45500.0 ;
      RECT  50295.0 46845.0 51000.0 48190.0 ;
      RECT  50295.0 49535.0 51000.0 48190.0 ;
      RECT  50295.0 49535.0 51000.0 50880.0 ;
      RECT  50295.0 52225.0 51000.0 50880.0 ;
      RECT  50295.0 52225.0 51000.0 53570.0 ;
      RECT  50295.0 54915.0 51000.0 53570.0 ;
      RECT  50295.0 54915.0 51000.0 56260.0 ;
      RECT  50295.0 57605.0 51000.0 56260.0 ;
      RECT  50295.0 57605.0 51000.0 58950.0 ;
      RECT  50295.0 60295.0 51000.0 58950.0 ;
      RECT  50295.0 60295.0 51000.0 61640.0 ;
      RECT  50295.0 62985.0 51000.0 61640.0 ;
      RECT  50295.0 62985.0 51000.0 64330.0 ;
      RECT  50295.0 65675.0 51000.0 64330.0 ;
      RECT  50295.0 65675.0 51000.0 67020.0 ;
      RECT  50295.0 68365.0 51000.0 67020.0 ;
      RECT  50295.0 68365.0 51000.0 69710.0 ;
      RECT  50295.0 71055.0 51000.0 69710.0 ;
      RECT  50295.0 71055.0 51000.0 72400.0 ;
      RECT  50295.0 73745.0 51000.0 72400.0 ;
      RECT  50295.0 73745.0 51000.0 75090.0 ;
      RECT  50295.0 76435.0 51000.0 75090.0 ;
      RECT  50295.0 76435.0 51000.0 77780.0 ;
      RECT  50295.0 79125.0 51000.0 77780.0 ;
      RECT  50295.0 79125.0 51000.0 80470.0 ;
      RECT  50295.0 81815.0 51000.0 80470.0 ;
      RECT  50295.0 81815.0 51000.0 83160.0 ;
      RECT  50295.0 84505.0 51000.0 83160.0 ;
      RECT  50295.0 84505.0 51000.0 85850.0 ;
      RECT  50295.0 87195.0 51000.0 85850.0 ;
      RECT  50295.0 87195.0 51000.0 88540.0 ;
      RECT  50295.0 89885.0 51000.0 88540.0 ;
      RECT  50295.0 89885.0 51000.0 91230.0 ;
      RECT  50295.0 92575.0 51000.0 91230.0 ;
      RECT  50295.0 92575.0 51000.0 93920.0 ;
      RECT  50295.0 95265.0 51000.0 93920.0 ;
      RECT  50295.0 95265.0 51000.0 96610.0 ;
      RECT  50295.0 97955.0 51000.0 96610.0 ;
      RECT  50295.0 97955.0 51000.0 99300.0 ;
      RECT  50295.0 100645.0 51000.0 99300.0 ;
      RECT  50295.0 100645.0 51000.0 101990.0 ;
      RECT  50295.0 103335.0 51000.0 101990.0 ;
      RECT  50295.0 103335.0 51000.0 104680.0 ;
      RECT  50295.0 106025.0 51000.0 104680.0 ;
      RECT  50295.0 106025.0 51000.0 107370.0 ;
      RECT  50295.0 108715.0 51000.0 107370.0 ;
      RECT  50295.0 108715.0 51000.0 110060.0 ;
      RECT  50295.0 111405.0 51000.0 110060.0 ;
      RECT  50295.0 111405.0 51000.0 112750.0 ;
      RECT  50295.0 114095.0 51000.0 112750.0 ;
      RECT  51000.0 28015.0 51705.0 29360.0 ;
      RECT  51000.0 30705.0 51705.0 29360.0 ;
      RECT  51000.0 30705.0 51705.0 32050.0 ;
      RECT  51000.0 33395.0 51705.0 32050.0 ;
      RECT  51000.0 33395.0 51705.0 34740.0 ;
      RECT  51000.0 36085.0 51705.0 34740.0 ;
      RECT  51000.0 36085.0 51705.0 37430.0 ;
      RECT  51000.0 38775.0 51705.0 37430.0 ;
      RECT  51000.0 38775.0 51705.0 40120.0 ;
      RECT  51000.0 41465.0 51705.0 40120.0 ;
      RECT  51000.0 41465.0 51705.0 42810.0 ;
      RECT  51000.0 44155.0 51705.0 42810.0 ;
      RECT  51000.0 44155.0 51705.0 45500.0 ;
      RECT  51000.0 46845.0 51705.0 45500.0 ;
      RECT  51000.0 46845.0 51705.0 48190.0 ;
      RECT  51000.0 49535.0 51705.0 48190.0 ;
      RECT  51000.0 49535.0 51705.0 50880.0 ;
      RECT  51000.0 52225.0 51705.0 50880.0 ;
      RECT  51000.0 52225.0 51705.0 53570.0 ;
      RECT  51000.0 54915.0 51705.0 53570.0 ;
      RECT  51000.0 54915.0 51705.0 56260.0 ;
      RECT  51000.0 57605.0 51705.0 56260.0 ;
      RECT  51000.0 57605.0 51705.0 58950.0 ;
      RECT  51000.0 60295.0 51705.0 58950.0 ;
      RECT  51000.0 60295.0 51705.0 61640.0 ;
      RECT  51000.0 62985.0 51705.0 61640.0 ;
      RECT  51000.0 62985.0 51705.0 64330.0 ;
      RECT  51000.0 65675.0 51705.0 64330.0 ;
      RECT  51000.0 65675.0 51705.0 67020.0 ;
      RECT  51000.0 68365.0 51705.0 67020.0 ;
      RECT  51000.0 68365.0 51705.0 69710.0 ;
      RECT  51000.0 71055.0 51705.0 69710.0 ;
      RECT  51000.0 71055.0 51705.0 72400.0 ;
      RECT  51000.0 73745.0 51705.0 72400.0 ;
      RECT  51000.0 73745.0 51705.0 75090.0 ;
      RECT  51000.0 76435.0 51705.0 75090.0 ;
      RECT  51000.0 76435.0 51705.0 77780.0 ;
      RECT  51000.0 79125.0 51705.0 77780.0 ;
      RECT  51000.0 79125.0 51705.0 80470.0 ;
      RECT  51000.0 81815.0 51705.0 80470.0 ;
      RECT  51000.0 81815.0 51705.0 83160.0 ;
      RECT  51000.0 84505.0 51705.0 83160.0 ;
      RECT  51000.0 84505.0 51705.0 85850.0 ;
      RECT  51000.0 87195.0 51705.0 85850.0 ;
      RECT  51000.0 87195.0 51705.0 88540.0 ;
      RECT  51000.0 89885.0 51705.0 88540.0 ;
      RECT  51000.0 89885.0 51705.0 91230.0 ;
      RECT  51000.0 92575.0 51705.0 91230.0 ;
      RECT  51000.0 92575.0 51705.0 93920.0 ;
      RECT  51000.0 95265.0 51705.0 93920.0 ;
      RECT  51000.0 95265.0 51705.0 96610.0 ;
      RECT  51000.0 97955.0 51705.0 96610.0 ;
      RECT  51000.0 97955.0 51705.0 99300.0 ;
      RECT  51000.0 100645.0 51705.0 99300.0 ;
      RECT  51000.0 100645.0 51705.0 101990.0 ;
      RECT  51000.0 103335.0 51705.0 101990.0 ;
      RECT  51000.0 103335.0 51705.0 104680.0 ;
      RECT  51000.0 106025.0 51705.0 104680.0 ;
      RECT  51000.0 106025.0 51705.0 107370.0 ;
      RECT  51000.0 108715.0 51705.0 107370.0 ;
      RECT  51000.0 108715.0 51705.0 110060.0 ;
      RECT  51000.0 111405.0 51705.0 110060.0 ;
      RECT  51000.0 111405.0 51705.0 112750.0 ;
      RECT  51000.0 114095.0 51705.0 112750.0 ;
      RECT  51705.0 28015.0 52410.0 29360.0 ;
      RECT  51705.0 30705.0 52410.0 29360.0 ;
      RECT  51705.0 30705.0 52410.0 32050.0 ;
      RECT  51705.0 33395.0 52410.0 32050.0 ;
      RECT  51705.0 33395.0 52410.0 34740.0 ;
      RECT  51705.0 36085.0 52410.0 34740.0 ;
      RECT  51705.0 36085.0 52410.0 37430.0 ;
      RECT  51705.0 38775.0 52410.0 37430.0 ;
      RECT  51705.0 38775.0 52410.0 40120.0 ;
      RECT  51705.0 41465.0 52410.0 40120.0 ;
      RECT  51705.0 41465.0 52410.0 42810.0 ;
      RECT  51705.0 44155.0 52410.0 42810.0 ;
      RECT  51705.0 44155.0 52410.0 45500.0 ;
      RECT  51705.0 46845.0 52410.0 45500.0 ;
      RECT  51705.0 46845.0 52410.0 48190.0 ;
      RECT  51705.0 49535.0 52410.0 48190.0 ;
      RECT  51705.0 49535.0 52410.0 50880.0 ;
      RECT  51705.0 52225.0 52410.0 50880.0 ;
      RECT  51705.0 52225.0 52410.0 53570.0 ;
      RECT  51705.0 54915.0 52410.0 53570.0 ;
      RECT  51705.0 54915.0 52410.0 56260.0 ;
      RECT  51705.0 57605.0 52410.0 56260.0 ;
      RECT  51705.0 57605.0 52410.0 58950.0 ;
      RECT  51705.0 60295.0 52410.0 58950.0 ;
      RECT  51705.0 60295.0 52410.0 61640.0 ;
      RECT  51705.0 62985.0 52410.0 61640.0 ;
      RECT  51705.0 62985.0 52410.0 64330.0 ;
      RECT  51705.0 65675.0 52410.0 64330.0 ;
      RECT  51705.0 65675.0 52410.0 67020.0 ;
      RECT  51705.0 68365.0 52410.0 67020.0 ;
      RECT  51705.0 68365.0 52410.0 69710.0 ;
      RECT  51705.0 71055.0 52410.0 69710.0 ;
      RECT  51705.0 71055.0 52410.0 72400.0 ;
      RECT  51705.0 73745.0 52410.0 72400.0 ;
      RECT  51705.0 73745.0 52410.0 75090.0 ;
      RECT  51705.0 76435.0 52410.0 75090.0 ;
      RECT  51705.0 76435.0 52410.0 77780.0 ;
      RECT  51705.0 79125.0 52410.0 77780.0 ;
      RECT  51705.0 79125.0 52410.0 80470.0 ;
      RECT  51705.0 81815.0 52410.0 80470.0 ;
      RECT  51705.0 81815.0 52410.0 83160.0 ;
      RECT  51705.0 84505.0 52410.0 83160.0 ;
      RECT  51705.0 84505.0 52410.0 85850.0 ;
      RECT  51705.0 87195.0 52410.0 85850.0 ;
      RECT  51705.0 87195.0 52410.0 88540.0 ;
      RECT  51705.0 89885.0 52410.0 88540.0 ;
      RECT  51705.0 89885.0 52410.0 91230.0 ;
      RECT  51705.0 92575.0 52410.0 91230.0 ;
      RECT  51705.0 92575.0 52410.0 93920.0 ;
      RECT  51705.0 95265.0 52410.0 93920.0 ;
      RECT  51705.0 95265.0 52410.0 96610.0 ;
      RECT  51705.0 97955.0 52410.0 96610.0 ;
      RECT  51705.0 97955.0 52410.0 99300.0 ;
      RECT  51705.0 100645.0 52410.0 99300.0 ;
      RECT  51705.0 100645.0 52410.0 101990.0 ;
      RECT  51705.0 103335.0 52410.0 101990.0 ;
      RECT  51705.0 103335.0 52410.0 104680.0 ;
      RECT  51705.0 106025.0 52410.0 104680.0 ;
      RECT  51705.0 106025.0 52410.0 107370.0 ;
      RECT  51705.0 108715.0 52410.0 107370.0 ;
      RECT  51705.0 108715.0 52410.0 110060.0 ;
      RECT  51705.0 111405.0 52410.0 110060.0 ;
      RECT  51705.0 111405.0 52410.0 112750.0 ;
      RECT  51705.0 114095.0 52410.0 112750.0 ;
      RECT  52410.0 28015.0 53115.0 29360.0 ;
      RECT  52410.0 30705.0 53115.0 29360.0 ;
      RECT  52410.0 30705.0 53115.0 32050.0 ;
      RECT  52410.0 33395.0 53115.0 32050.0 ;
      RECT  52410.0 33395.0 53115.0 34740.0 ;
      RECT  52410.0 36085.0 53115.0 34740.0 ;
      RECT  52410.0 36085.0 53115.0 37430.0 ;
      RECT  52410.0 38775.0 53115.0 37430.0 ;
      RECT  52410.0 38775.0 53115.0 40120.0 ;
      RECT  52410.0 41465.0 53115.0 40120.0 ;
      RECT  52410.0 41465.0 53115.0 42810.0 ;
      RECT  52410.0 44155.0 53115.0 42810.0 ;
      RECT  52410.0 44155.0 53115.0 45500.0 ;
      RECT  52410.0 46845.0 53115.0 45500.0 ;
      RECT  52410.0 46845.0 53115.0 48190.0 ;
      RECT  52410.0 49535.0 53115.0 48190.0 ;
      RECT  52410.0 49535.0 53115.0 50880.0 ;
      RECT  52410.0 52225.0 53115.0 50880.0 ;
      RECT  52410.0 52225.0 53115.0 53570.0 ;
      RECT  52410.0 54915.0 53115.0 53570.0 ;
      RECT  52410.0 54915.0 53115.0 56260.0 ;
      RECT  52410.0 57605.0 53115.0 56260.0 ;
      RECT  52410.0 57605.0 53115.0 58950.0 ;
      RECT  52410.0 60295.0 53115.0 58950.0 ;
      RECT  52410.0 60295.0 53115.0 61640.0 ;
      RECT  52410.0 62985.0 53115.0 61640.0 ;
      RECT  52410.0 62985.0 53115.0 64330.0 ;
      RECT  52410.0 65675.0 53115.0 64330.0 ;
      RECT  52410.0 65675.0 53115.0 67020.0 ;
      RECT  52410.0 68365.0 53115.0 67020.0 ;
      RECT  52410.0 68365.0 53115.0 69710.0 ;
      RECT  52410.0 71055.0 53115.0 69710.0 ;
      RECT  52410.0 71055.0 53115.0 72400.0 ;
      RECT  52410.0 73745.0 53115.0 72400.0 ;
      RECT  52410.0 73745.0 53115.0 75090.0 ;
      RECT  52410.0 76435.0 53115.0 75090.0 ;
      RECT  52410.0 76435.0 53115.0 77780.0 ;
      RECT  52410.0 79125.0 53115.0 77780.0 ;
      RECT  52410.0 79125.0 53115.0 80470.0 ;
      RECT  52410.0 81815.0 53115.0 80470.0 ;
      RECT  52410.0 81815.0 53115.0 83160.0 ;
      RECT  52410.0 84505.0 53115.0 83160.0 ;
      RECT  52410.0 84505.0 53115.0 85850.0 ;
      RECT  52410.0 87195.0 53115.0 85850.0 ;
      RECT  52410.0 87195.0 53115.0 88540.0 ;
      RECT  52410.0 89885.0 53115.0 88540.0 ;
      RECT  52410.0 89885.0 53115.0 91230.0 ;
      RECT  52410.0 92575.0 53115.0 91230.0 ;
      RECT  52410.0 92575.0 53115.0 93920.0 ;
      RECT  52410.0 95265.0 53115.0 93920.0 ;
      RECT  52410.0 95265.0 53115.0 96610.0 ;
      RECT  52410.0 97955.0 53115.0 96610.0 ;
      RECT  52410.0 97955.0 53115.0 99300.0 ;
      RECT  52410.0 100645.0 53115.0 99300.0 ;
      RECT  52410.0 100645.0 53115.0 101990.0 ;
      RECT  52410.0 103335.0 53115.0 101990.0 ;
      RECT  52410.0 103335.0 53115.0 104680.0 ;
      RECT  52410.0 106025.0 53115.0 104680.0 ;
      RECT  52410.0 106025.0 53115.0 107370.0 ;
      RECT  52410.0 108715.0 53115.0 107370.0 ;
      RECT  52410.0 108715.0 53115.0 110060.0 ;
      RECT  52410.0 111405.0 53115.0 110060.0 ;
      RECT  52410.0 111405.0 53115.0 112750.0 ;
      RECT  52410.0 114095.0 53115.0 112750.0 ;
      RECT  53115.0 28015.0 53820.0 29360.0 ;
      RECT  53115.0 30705.0 53820.0 29360.0 ;
      RECT  53115.0 30705.0 53820.0 32050.0 ;
      RECT  53115.0 33395.0 53820.0 32050.0 ;
      RECT  53115.0 33395.0 53820.0 34740.0 ;
      RECT  53115.0 36085.0 53820.0 34740.0 ;
      RECT  53115.0 36085.0 53820.0 37430.0 ;
      RECT  53115.0 38775.0 53820.0 37430.0 ;
      RECT  53115.0 38775.0 53820.0 40120.0 ;
      RECT  53115.0 41465.0 53820.0 40120.0 ;
      RECT  53115.0 41465.0 53820.0 42810.0 ;
      RECT  53115.0 44155.0 53820.0 42810.0 ;
      RECT  53115.0 44155.0 53820.0 45500.0 ;
      RECT  53115.0 46845.0 53820.0 45500.0 ;
      RECT  53115.0 46845.0 53820.0 48190.0 ;
      RECT  53115.0 49535.0 53820.0 48190.0 ;
      RECT  53115.0 49535.0 53820.0 50880.0 ;
      RECT  53115.0 52225.0 53820.0 50880.0 ;
      RECT  53115.0 52225.0 53820.0 53570.0 ;
      RECT  53115.0 54915.0 53820.0 53570.0 ;
      RECT  53115.0 54915.0 53820.0 56260.0 ;
      RECT  53115.0 57605.0 53820.0 56260.0 ;
      RECT  53115.0 57605.0 53820.0 58950.0 ;
      RECT  53115.0 60295.0 53820.0 58950.0 ;
      RECT  53115.0 60295.0 53820.0 61640.0 ;
      RECT  53115.0 62985.0 53820.0 61640.0 ;
      RECT  53115.0 62985.0 53820.0 64330.0 ;
      RECT  53115.0 65675.0 53820.0 64330.0 ;
      RECT  53115.0 65675.0 53820.0 67020.0 ;
      RECT  53115.0 68365.0 53820.0 67020.0 ;
      RECT  53115.0 68365.0 53820.0 69710.0 ;
      RECT  53115.0 71055.0 53820.0 69710.0 ;
      RECT  53115.0 71055.0 53820.0 72400.0 ;
      RECT  53115.0 73745.0 53820.0 72400.0 ;
      RECT  53115.0 73745.0 53820.0 75090.0 ;
      RECT  53115.0 76435.0 53820.0 75090.0 ;
      RECT  53115.0 76435.0 53820.0 77780.0 ;
      RECT  53115.0 79125.0 53820.0 77780.0 ;
      RECT  53115.0 79125.0 53820.0 80470.0 ;
      RECT  53115.0 81815.0 53820.0 80470.0 ;
      RECT  53115.0 81815.0 53820.0 83160.0 ;
      RECT  53115.0 84505.0 53820.0 83160.0 ;
      RECT  53115.0 84505.0 53820.0 85850.0 ;
      RECT  53115.0 87195.0 53820.0 85850.0 ;
      RECT  53115.0 87195.0 53820.0 88540.0 ;
      RECT  53115.0 89885.0 53820.0 88540.0 ;
      RECT  53115.0 89885.0 53820.0 91230.0 ;
      RECT  53115.0 92575.0 53820.0 91230.0 ;
      RECT  53115.0 92575.0 53820.0 93920.0 ;
      RECT  53115.0 95265.0 53820.0 93920.0 ;
      RECT  53115.0 95265.0 53820.0 96610.0 ;
      RECT  53115.0 97955.0 53820.0 96610.0 ;
      RECT  53115.0 97955.0 53820.0 99300.0 ;
      RECT  53115.0 100645.0 53820.0 99300.0 ;
      RECT  53115.0 100645.0 53820.0 101990.0 ;
      RECT  53115.0 103335.0 53820.0 101990.0 ;
      RECT  53115.0 103335.0 53820.0 104680.0 ;
      RECT  53115.0 106025.0 53820.0 104680.0 ;
      RECT  53115.0 106025.0 53820.0 107370.0 ;
      RECT  53115.0 108715.0 53820.0 107370.0 ;
      RECT  53115.0 108715.0 53820.0 110060.0 ;
      RECT  53115.0 111405.0 53820.0 110060.0 ;
      RECT  53115.0 111405.0 53820.0 112750.0 ;
      RECT  53115.0 114095.0 53820.0 112750.0 ;
      RECT  53820.0 28015.0 54525.0 29360.0 ;
      RECT  53820.0 30705.0 54525.0 29360.0 ;
      RECT  53820.0 30705.0 54525.0 32050.0 ;
      RECT  53820.0 33395.0 54525.0 32050.0 ;
      RECT  53820.0 33395.0 54525.0 34740.0 ;
      RECT  53820.0 36085.0 54525.0 34740.0 ;
      RECT  53820.0 36085.0 54525.0 37430.0 ;
      RECT  53820.0 38775.0 54525.0 37430.0 ;
      RECT  53820.0 38775.0 54525.0 40120.0 ;
      RECT  53820.0 41465.0 54525.0 40120.0 ;
      RECT  53820.0 41465.0 54525.0 42810.0 ;
      RECT  53820.0 44155.0 54525.0 42810.0 ;
      RECT  53820.0 44155.0 54525.0 45500.0 ;
      RECT  53820.0 46845.0 54525.0 45500.0 ;
      RECT  53820.0 46845.0 54525.0 48190.0 ;
      RECT  53820.0 49535.0 54525.0 48190.0 ;
      RECT  53820.0 49535.0 54525.0 50880.0 ;
      RECT  53820.0 52225.0 54525.0 50880.0 ;
      RECT  53820.0 52225.0 54525.0 53570.0 ;
      RECT  53820.0 54915.0 54525.0 53570.0 ;
      RECT  53820.0 54915.0 54525.0 56260.0 ;
      RECT  53820.0 57605.0 54525.0 56260.0 ;
      RECT  53820.0 57605.0 54525.0 58950.0 ;
      RECT  53820.0 60295.0 54525.0 58950.0 ;
      RECT  53820.0 60295.0 54525.0 61640.0 ;
      RECT  53820.0 62985.0 54525.0 61640.0 ;
      RECT  53820.0 62985.0 54525.0 64330.0 ;
      RECT  53820.0 65675.0 54525.0 64330.0 ;
      RECT  53820.0 65675.0 54525.0 67020.0 ;
      RECT  53820.0 68365.0 54525.0 67020.0 ;
      RECT  53820.0 68365.0 54525.0 69710.0 ;
      RECT  53820.0 71055.0 54525.0 69710.0 ;
      RECT  53820.0 71055.0 54525.0 72400.0 ;
      RECT  53820.0 73745.0 54525.0 72400.0 ;
      RECT  53820.0 73745.0 54525.0 75090.0 ;
      RECT  53820.0 76435.0 54525.0 75090.0 ;
      RECT  53820.0 76435.0 54525.0 77780.0 ;
      RECT  53820.0 79125.0 54525.0 77780.0 ;
      RECT  53820.0 79125.0 54525.0 80470.0 ;
      RECT  53820.0 81815.0 54525.0 80470.0 ;
      RECT  53820.0 81815.0 54525.0 83160.0 ;
      RECT  53820.0 84505.0 54525.0 83160.0 ;
      RECT  53820.0 84505.0 54525.0 85850.0 ;
      RECT  53820.0 87195.0 54525.0 85850.0 ;
      RECT  53820.0 87195.0 54525.0 88540.0 ;
      RECT  53820.0 89885.0 54525.0 88540.0 ;
      RECT  53820.0 89885.0 54525.0 91230.0 ;
      RECT  53820.0 92575.0 54525.0 91230.0 ;
      RECT  53820.0 92575.0 54525.0 93920.0 ;
      RECT  53820.0 95265.0 54525.0 93920.0 ;
      RECT  53820.0 95265.0 54525.0 96610.0 ;
      RECT  53820.0 97955.0 54525.0 96610.0 ;
      RECT  53820.0 97955.0 54525.0 99300.0 ;
      RECT  53820.0 100645.0 54525.0 99300.0 ;
      RECT  53820.0 100645.0 54525.0 101990.0 ;
      RECT  53820.0 103335.0 54525.0 101990.0 ;
      RECT  53820.0 103335.0 54525.0 104680.0 ;
      RECT  53820.0 106025.0 54525.0 104680.0 ;
      RECT  53820.0 106025.0 54525.0 107370.0 ;
      RECT  53820.0 108715.0 54525.0 107370.0 ;
      RECT  53820.0 108715.0 54525.0 110060.0 ;
      RECT  53820.0 111405.0 54525.0 110060.0 ;
      RECT  53820.0 111405.0 54525.0 112750.0 ;
      RECT  53820.0 114095.0 54525.0 112750.0 ;
      RECT  54525.0 28015.0 55230.0 29360.0 ;
      RECT  54525.0 30705.0 55230.0 29360.0 ;
      RECT  54525.0 30705.0 55230.0 32050.0 ;
      RECT  54525.0 33395.0 55230.0 32050.0 ;
      RECT  54525.0 33395.0 55230.0 34740.0 ;
      RECT  54525.0 36085.0 55230.0 34740.0 ;
      RECT  54525.0 36085.0 55230.0 37430.0 ;
      RECT  54525.0 38775.0 55230.0 37430.0 ;
      RECT  54525.0 38775.0 55230.0 40120.0 ;
      RECT  54525.0 41465.0 55230.0 40120.0 ;
      RECT  54525.0 41465.0 55230.0 42810.0 ;
      RECT  54525.0 44155.0 55230.0 42810.0 ;
      RECT  54525.0 44155.0 55230.0 45500.0 ;
      RECT  54525.0 46845.0 55230.0 45500.0 ;
      RECT  54525.0 46845.0 55230.0 48190.0 ;
      RECT  54525.0 49535.0 55230.0 48190.0 ;
      RECT  54525.0 49535.0 55230.0 50880.0 ;
      RECT  54525.0 52225.0 55230.0 50880.0 ;
      RECT  54525.0 52225.0 55230.0 53570.0 ;
      RECT  54525.0 54915.0 55230.0 53570.0 ;
      RECT  54525.0 54915.0 55230.0 56260.0 ;
      RECT  54525.0 57605.0 55230.0 56260.0 ;
      RECT  54525.0 57605.0 55230.0 58950.0 ;
      RECT  54525.0 60295.0 55230.0 58950.0 ;
      RECT  54525.0 60295.0 55230.0 61640.0 ;
      RECT  54525.0 62985.0 55230.0 61640.0 ;
      RECT  54525.0 62985.0 55230.0 64330.0 ;
      RECT  54525.0 65675.0 55230.0 64330.0 ;
      RECT  54525.0 65675.0 55230.0 67020.0 ;
      RECT  54525.0 68365.0 55230.0 67020.0 ;
      RECT  54525.0 68365.0 55230.0 69710.0 ;
      RECT  54525.0 71055.0 55230.0 69710.0 ;
      RECT  54525.0 71055.0 55230.0 72400.0 ;
      RECT  54525.0 73745.0 55230.0 72400.0 ;
      RECT  54525.0 73745.0 55230.0 75090.0 ;
      RECT  54525.0 76435.0 55230.0 75090.0 ;
      RECT  54525.0 76435.0 55230.0 77780.0 ;
      RECT  54525.0 79125.0 55230.0 77780.0 ;
      RECT  54525.0 79125.0 55230.0 80470.0 ;
      RECT  54525.0 81815.0 55230.0 80470.0 ;
      RECT  54525.0 81815.0 55230.0 83160.0 ;
      RECT  54525.0 84505.0 55230.0 83160.0 ;
      RECT  54525.0 84505.0 55230.0 85850.0 ;
      RECT  54525.0 87195.0 55230.0 85850.0 ;
      RECT  54525.0 87195.0 55230.0 88540.0 ;
      RECT  54525.0 89885.0 55230.0 88540.0 ;
      RECT  54525.0 89885.0 55230.0 91230.0 ;
      RECT  54525.0 92575.0 55230.0 91230.0 ;
      RECT  54525.0 92575.0 55230.0 93920.0 ;
      RECT  54525.0 95265.0 55230.0 93920.0 ;
      RECT  54525.0 95265.0 55230.0 96610.0 ;
      RECT  54525.0 97955.0 55230.0 96610.0 ;
      RECT  54525.0 97955.0 55230.0 99300.0 ;
      RECT  54525.0 100645.0 55230.0 99300.0 ;
      RECT  54525.0 100645.0 55230.0 101990.0 ;
      RECT  54525.0 103335.0 55230.0 101990.0 ;
      RECT  54525.0 103335.0 55230.0 104680.0 ;
      RECT  54525.0 106025.0 55230.0 104680.0 ;
      RECT  54525.0 106025.0 55230.0 107370.0 ;
      RECT  54525.0 108715.0 55230.0 107370.0 ;
      RECT  54525.0 108715.0 55230.0 110060.0 ;
      RECT  54525.0 111405.0 55230.0 110060.0 ;
      RECT  54525.0 111405.0 55230.0 112750.0 ;
      RECT  54525.0 114095.0 55230.0 112750.0 ;
      RECT  55230.0 28015.0 55935.0 29360.0 ;
      RECT  55230.0 30705.0 55935.0 29360.0 ;
      RECT  55230.0 30705.0 55935.0 32050.0 ;
      RECT  55230.0 33395.0 55935.0 32050.0 ;
      RECT  55230.0 33395.0 55935.0 34740.0 ;
      RECT  55230.0 36085.0 55935.0 34740.0 ;
      RECT  55230.0 36085.0 55935.0 37430.0 ;
      RECT  55230.0 38775.0 55935.0 37430.0 ;
      RECT  55230.0 38775.0 55935.0 40120.0 ;
      RECT  55230.0 41465.0 55935.0 40120.0 ;
      RECT  55230.0 41465.0 55935.0 42810.0 ;
      RECT  55230.0 44155.0 55935.0 42810.0 ;
      RECT  55230.0 44155.0 55935.0 45500.0 ;
      RECT  55230.0 46845.0 55935.0 45500.0 ;
      RECT  55230.0 46845.0 55935.0 48190.0 ;
      RECT  55230.0 49535.0 55935.0 48190.0 ;
      RECT  55230.0 49535.0 55935.0 50880.0 ;
      RECT  55230.0 52225.0 55935.0 50880.0 ;
      RECT  55230.0 52225.0 55935.0 53570.0 ;
      RECT  55230.0 54915.0 55935.0 53570.0 ;
      RECT  55230.0 54915.0 55935.0 56260.0 ;
      RECT  55230.0 57605.0 55935.0 56260.0 ;
      RECT  55230.0 57605.0 55935.0 58950.0 ;
      RECT  55230.0 60295.0 55935.0 58950.0 ;
      RECT  55230.0 60295.0 55935.0 61640.0 ;
      RECT  55230.0 62985.0 55935.0 61640.0 ;
      RECT  55230.0 62985.0 55935.0 64330.0 ;
      RECT  55230.0 65675.0 55935.0 64330.0 ;
      RECT  55230.0 65675.0 55935.0 67020.0 ;
      RECT  55230.0 68365.0 55935.0 67020.0 ;
      RECT  55230.0 68365.0 55935.0 69710.0 ;
      RECT  55230.0 71055.0 55935.0 69710.0 ;
      RECT  55230.0 71055.0 55935.0 72400.0 ;
      RECT  55230.0 73745.0 55935.0 72400.0 ;
      RECT  55230.0 73745.0 55935.0 75090.0 ;
      RECT  55230.0 76435.0 55935.0 75090.0 ;
      RECT  55230.0 76435.0 55935.0 77780.0 ;
      RECT  55230.0 79125.0 55935.0 77780.0 ;
      RECT  55230.0 79125.0 55935.0 80470.0 ;
      RECT  55230.0 81815.0 55935.0 80470.0 ;
      RECT  55230.0 81815.0 55935.0 83160.0 ;
      RECT  55230.0 84505.0 55935.0 83160.0 ;
      RECT  55230.0 84505.0 55935.0 85850.0 ;
      RECT  55230.0 87195.0 55935.0 85850.0 ;
      RECT  55230.0 87195.0 55935.0 88540.0 ;
      RECT  55230.0 89885.0 55935.0 88540.0 ;
      RECT  55230.0 89885.0 55935.0 91230.0 ;
      RECT  55230.0 92575.0 55935.0 91230.0 ;
      RECT  55230.0 92575.0 55935.0 93920.0 ;
      RECT  55230.0 95265.0 55935.0 93920.0 ;
      RECT  55230.0 95265.0 55935.0 96610.0 ;
      RECT  55230.0 97955.0 55935.0 96610.0 ;
      RECT  55230.0 97955.0 55935.0 99300.0 ;
      RECT  55230.0 100645.0 55935.0 99300.0 ;
      RECT  55230.0 100645.0 55935.0 101990.0 ;
      RECT  55230.0 103335.0 55935.0 101990.0 ;
      RECT  55230.0 103335.0 55935.0 104680.0 ;
      RECT  55230.0 106025.0 55935.0 104680.0 ;
      RECT  55230.0 106025.0 55935.0 107370.0 ;
      RECT  55230.0 108715.0 55935.0 107370.0 ;
      RECT  55230.0 108715.0 55935.0 110060.0 ;
      RECT  55230.0 111405.0 55935.0 110060.0 ;
      RECT  55230.0 111405.0 55935.0 112750.0 ;
      RECT  55230.0 114095.0 55935.0 112750.0 ;
      RECT  55935.0 28015.0 56640.0 29360.0 ;
      RECT  55935.0 30705.0 56640.0 29360.0 ;
      RECT  55935.0 30705.0 56640.0 32050.0 ;
      RECT  55935.0 33395.0 56640.0 32050.0 ;
      RECT  55935.0 33395.0 56640.0 34740.0 ;
      RECT  55935.0 36085.0 56640.0 34740.0 ;
      RECT  55935.0 36085.0 56640.0 37430.0 ;
      RECT  55935.0 38775.0 56640.0 37430.0 ;
      RECT  55935.0 38775.0 56640.0 40120.0 ;
      RECT  55935.0 41465.0 56640.0 40120.0 ;
      RECT  55935.0 41465.0 56640.0 42810.0 ;
      RECT  55935.0 44155.0 56640.0 42810.0 ;
      RECT  55935.0 44155.0 56640.0 45500.0 ;
      RECT  55935.0 46845.0 56640.0 45500.0 ;
      RECT  55935.0 46845.0 56640.0 48190.0 ;
      RECT  55935.0 49535.0 56640.0 48190.0 ;
      RECT  55935.0 49535.0 56640.0 50880.0 ;
      RECT  55935.0 52225.0 56640.0 50880.0 ;
      RECT  55935.0 52225.0 56640.0 53570.0 ;
      RECT  55935.0 54915.0 56640.0 53570.0 ;
      RECT  55935.0 54915.0 56640.0 56260.0 ;
      RECT  55935.0 57605.0 56640.0 56260.0 ;
      RECT  55935.0 57605.0 56640.0 58950.0 ;
      RECT  55935.0 60295.0 56640.0 58950.0 ;
      RECT  55935.0 60295.0 56640.0 61640.0 ;
      RECT  55935.0 62985.0 56640.0 61640.0 ;
      RECT  55935.0 62985.0 56640.0 64330.0 ;
      RECT  55935.0 65675.0 56640.0 64330.0 ;
      RECT  55935.0 65675.0 56640.0 67020.0 ;
      RECT  55935.0 68365.0 56640.0 67020.0 ;
      RECT  55935.0 68365.0 56640.0 69710.0 ;
      RECT  55935.0 71055.0 56640.0 69710.0 ;
      RECT  55935.0 71055.0 56640.0 72400.0 ;
      RECT  55935.0 73745.0 56640.0 72400.0 ;
      RECT  55935.0 73745.0 56640.0 75090.0 ;
      RECT  55935.0 76435.0 56640.0 75090.0 ;
      RECT  55935.0 76435.0 56640.0 77780.0 ;
      RECT  55935.0 79125.0 56640.0 77780.0 ;
      RECT  55935.0 79125.0 56640.0 80470.0 ;
      RECT  55935.0 81815.0 56640.0 80470.0 ;
      RECT  55935.0 81815.0 56640.0 83160.0 ;
      RECT  55935.0 84505.0 56640.0 83160.0 ;
      RECT  55935.0 84505.0 56640.0 85850.0 ;
      RECT  55935.0 87195.0 56640.0 85850.0 ;
      RECT  55935.0 87195.0 56640.0 88540.0 ;
      RECT  55935.0 89885.0 56640.0 88540.0 ;
      RECT  55935.0 89885.0 56640.0 91230.0 ;
      RECT  55935.0 92575.0 56640.0 91230.0 ;
      RECT  55935.0 92575.0 56640.0 93920.0 ;
      RECT  55935.0 95265.0 56640.0 93920.0 ;
      RECT  55935.0 95265.0 56640.0 96610.0 ;
      RECT  55935.0 97955.0 56640.0 96610.0 ;
      RECT  55935.0 97955.0 56640.0 99300.0 ;
      RECT  55935.0 100645.0 56640.0 99300.0 ;
      RECT  55935.0 100645.0 56640.0 101990.0 ;
      RECT  55935.0 103335.0 56640.0 101990.0 ;
      RECT  55935.0 103335.0 56640.0 104680.0 ;
      RECT  55935.0 106025.0 56640.0 104680.0 ;
      RECT  55935.0 106025.0 56640.0 107370.0 ;
      RECT  55935.0 108715.0 56640.0 107370.0 ;
      RECT  55935.0 108715.0 56640.0 110060.0 ;
      RECT  55935.0 111405.0 56640.0 110060.0 ;
      RECT  55935.0 111405.0 56640.0 112750.0 ;
      RECT  55935.0 114095.0 56640.0 112750.0 ;
      RECT  56640.0 28015.0 57345.0 29360.0 ;
      RECT  56640.0 30705.0 57345.0 29360.0 ;
      RECT  56640.0 30705.0 57345.0 32050.0 ;
      RECT  56640.0 33395.0 57345.0 32050.0 ;
      RECT  56640.0 33395.0 57345.0 34740.0 ;
      RECT  56640.0 36085.0 57345.0 34740.0 ;
      RECT  56640.0 36085.0 57345.0 37430.0 ;
      RECT  56640.0 38775.0 57345.0 37430.0 ;
      RECT  56640.0 38775.0 57345.0 40120.0 ;
      RECT  56640.0 41465.0 57345.0 40120.0 ;
      RECT  56640.0 41465.0 57345.0 42810.0 ;
      RECT  56640.0 44155.0 57345.0 42810.0 ;
      RECT  56640.0 44155.0 57345.0 45500.0 ;
      RECT  56640.0 46845.0 57345.0 45500.0 ;
      RECT  56640.0 46845.0 57345.0 48190.0 ;
      RECT  56640.0 49535.0 57345.0 48190.0 ;
      RECT  56640.0 49535.0 57345.0 50880.0 ;
      RECT  56640.0 52225.0 57345.0 50880.0 ;
      RECT  56640.0 52225.0 57345.0 53570.0 ;
      RECT  56640.0 54915.0 57345.0 53570.0 ;
      RECT  56640.0 54915.0 57345.0 56260.0 ;
      RECT  56640.0 57605.0 57345.0 56260.0 ;
      RECT  56640.0 57605.0 57345.0 58950.0 ;
      RECT  56640.0 60295.0 57345.0 58950.0 ;
      RECT  56640.0 60295.0 57345.0 61640.0 ;
      RECT  56640.0 62985.0 57345.0 61640.0 ;
      RECT  56640.0 62985.0 57345.0 64330.0 ;
      RECT  56640.0 65675.0 57345.0 64330.0 ;
      RECT  56640.0 65675.0 57345.0 67020.0 ;
      RECT  56640.0 68365.0 57345.0 67020.0 ;
      RECT  56640.0 68365.0 57345.0 69710.0 ;
      RECT  56640.0 71055.0 57345.0 69710.0 ;
      RECT  56640.0 71055.0 57345.0 72400.0 ;
      RECT  56640.0 73745.0 57345.0 72400.0 ;
      RECT  56640.0 73745.0 57345.0 75090.0 ;
      RECT  56640.0 76435.0 57345.0 75090.0 ;
      RECT  56640.0 76435.0 57345.0 77780.0 ;
      RECT  56640.0 79125.0 57345.0 77780.0 ;
      RECT  56640.0 79125.0 57345.0 80470.0 ;
      RECT  56640.0 81815.0 57345.0 80470.0 ;
      RECT  56640.0 81815.0 57345.0 83160.0 ;
      RECT  56640.0 84505.0 57345.0 83160.0 ;
      RECT  56640.0 84505.0 57345.0 85850.0 ;
      RECT  56640.0 87195.0 57345.0 85850.0 ;
      RECT  56640.0 87195.0 57345.0 88540.0 ;
      RECT  56640.0 89885.0 57345.0 88540.0 ;
      RECT  56640.0 89885.0 57345.0 91230.0 ;
      RECT  56640.0 92575.0 57345.0 91230.0 ;
      RECT  56640.0 92575.0 57345.0 93920.0 ;
      RECT  56640.0 95265.0 57345.0 93920.0 ;
      RECT  56640.0 95265.0 57345.0 96610.0 ;
      RECT  56640.0 97955.0 57345.0 96610.0 ;
      RECT  56640.0 97955.0 57345.0 99300.0 ;
      RECT  56640.0 100645.0 57345.0 99300.0 ;
      RECT  56640.0 100645.0 57345.0 101990.0 ;
      RECT  56640.0 103335.0 57345.0 101990.0 ;
      RECT  56640.0 103335.0 57345.0 104680.0 ;
      RECT  56640.0 106025.0 57345.0 104680.0 ;
      RECT  56640.0 106025.0 57345.0 107370.0 ;
      RECT  56640.0 108715.0 57345.0 107370.0 ;
      RECT  56640.0 108715.0 57345.0 110060.0 ;
      RECT  56640.0 111405.0 57345.0 110060.0 ;
      RECT  56640.0 111405.0 57345.0 112750.0 ;
      RECT  56640.0 114095.0 57345.0 112750.0 ;
      RECT  57345.0 28015.0 58050.0 29360.0 ;
      RECT  57345.0 30705.0 58050.0 29360.0 ;
      RECT  57345.0 30705.0 58050.0 32050.0 ;
      RECT  57345.0 33395.0 58050.0 32050.0 ;
      RECT  57345.0 33395.0 58050.0 34740.0 ;
      RECT  57345.0 36085.0 58050.0 34740.0 ;
      RECT  57345.0 36085.0 58050.0 37430.0 ;
      RECT  57345.0 38775.0 58050.0 37430.0 ;
      RECT  57345.0 38775.0 58050.0 40120.0 ;
      RECT  57345.0 41465.0 58050.0 40120.0 ;
      RECT  57345.0 41465.0 58050.0 42810.0 ;
      RECT  57345.0 44155.0 58050.0 42810.0 ;
      RECT  57345.0 44155.0 58050.0 45500.0 ;
      RECT  57345.0 46845.0 58050.0 45500.0 ;
      RECT  57345.0 46845.0 58050.0 48190.0 ;
      RECT  57345.0 49535.0 58050.0 48190.0 ;
      RECT  57345.0 49535.0 58050.0 50880.0 ;
      RECT  57345.0 52225.0 58050.0 50880.0 ;
      RECT  57345.0 52225.0 58050.0 53570.0 ;
      RECT  57345.0 54915.0 58050.0 53570.0 ;
      RECT  57345.0 54915.0 58050.0 56260.0 ;
      RECT  57345.0 57605.0 58050.0 56260.0 ;
      RECT  57345.0 57605.0 58050.0 58950.0 ;
      RECT  57345.0 60295.0 58050.0 58950.0 ;
      RECT  57345.0 60295.0 58050.0 61640.0 ;
      RECT  57345.0 62985.0 58050.0 61640.0 ;
      RECT  57345.0 62985.0 58050.0 64330.0 ;
      RECT  57345.0 65675.0 58050.0 64330.0 ;
      RECT  57345.0 65675.0 58050.0 67020.0 ;
      RECT  57345.0 68365.0 58050.0 67020.0 ;
      RECT  57345.0 68365.0 58050.0 69710.0 ;
      RECT  57345.0 71055.0 58050.0 69710.0 ;
      RECT  57345.0 71055.0 58050.0 72400.0 ;
      RECT  57345.0 73745.0 58050.0 72400.0 ;
      RECT  57345.0 73745.0 58050.0 75090.0 ;
      RECT  57345.0 76435.0 58050.0 75090.0 ;
      RECT  57345.0 76435.0 58050.0 77780.0 ;
      RECT  57345.0 79125.0 58050.0 77780.0 ;
      RECT  57345.0 79125.0 58050.0 80470.0 ;
      RECT  57345.0 81815.0 58050.0 80470.0 ;
      RECT  57345.0 81815.0 58050.0 83160.0 ;
      RECT  57345.0 84505.0 58050.0 83160.0 ;
      RECT  57345.0 84505.0 58050.0 85850.0 ;
      RECT  57345.0 87195.0 58050.0 85850.0 ;
      RECT  57345.0 87195.0 58050.0 88540.0 ;
      RECT  57345.0 89885.0 58050.0 88540.0 ;
      RECT  57345.0 89885.0 58050.0 91230.0 ;
      RECT  57345.0 92575.0 58050.0 91230.0 ;
      RECT  57345.0 92575.0 58050.0 93920.0 ;
      RECT  57345.0 95265.0 58050.0 93920.0 ;
      RECT  57345.0 95265.0 58050.0 96610.0 ;
      RECT  57345.0 97955.0 58050.0 96610.0 ;
      RECT  57345.0 97955.0 58050.0 99300.0 ;
      RECT  57345.0 100645.0 58050.0 99300.0 ;
      RECT  57345.0 100645.0 58050.0 101990.0 ;
      RECT  57345.0 103335.0 58050.0 101990.0 ;
      RECT  57345.0 103335.0 58050.0 104680.0 ;
      RECT  57345.0 106025.0 58050.0 104680.0 ;
      RECT  57345.0 106025.0 58050.0 107370.0 ;
      RECT  57345.0 108715.0 58050.0 107370.0 ;
      RECT  57345.0 108715.0 58050.0 110060.0 ;
      RECT  57345.0 111405.0 58050.0 110060.0 ;
      RECT  57345.0 111405.0 58050.0 112750.0 ;
      RECT  57345.0 114095.0 58050.0 112750.0 ;
      RECT  58050.0 28015.0 58755.0 29360.0 ;
      RECT  58050.0 30705.0 58755.0 29360.0 ;
      RECT  58050.0 30705.0 58755.0 32050.0 ;
      RECT  58050.0 33395.0 58755.0 32050.0 ;
      RECT  58050.0 33395.0 58755.0 34740.0 ;
      RECT  58050.0 36085.0 58755.0 34740.0 ;
      RECT  58050.0 36085.0 58755.0 37430.0 ;
      RECT  58050.0 38775.0 58755.0 37430.0 ;
      RECT  58050.0 38775.0 58755.0 40120.0 ;
      RECT  58050.0 41465.0 58755.0 40120.0 ;
      RECT  58050.0 41465.0 58755.0 42810.0 ;
      RECT  58050.0 44155.0 58755.0 42810.0 ;
      RECT  58050.0 44155.0 58755.0 45500.0 ;
      RECT  58050.0 46845.0 58755.0 45500.0 ;
      RECT  58050.0 46845.0 58755.0 48190.0 ;
      RECT  58050.0 49535.0 58755.0 48190.0 ;
      RECT  58050.0 49535.0 58755.0 50880.0 ;
      RECT  58050.0 52225.0 58755.0 50880.0 ;
      RECT  58050.0 52225.0 58755.0 53570.0 ;
      RECT  58050.0 54915.0 58755.0 53570.0 ;
      RECT  58050.0 54915.0 58755.0 56260.0 ;
      RECT  58050.0 57605.0 58755.0 56260.0 ;
      RECT  58050.0 57605.0 58755.0 58950.0 ;
      RECT  58050.0 60295.0 58755.0 58950.0 ;
      RECT  58050.0 60295.0 58755.0 61640.0 ;
      RECT  58050.0 62985.0 58755.0 61640.0 ;
      RECT  58050.0 62985.0 58755.0 64330.0 ;
      RECT  58050.0 65675.0 58755.0 64330.0 ;
      RECT  58050.0 65675.0 58755.0 67020.0 ;
      RECT  58050.0 68365.0 58755.0 67020.0 ;
      RECT  58050.0 68365.0 58755.0 69710.0 ;
      RECT  58050.0 71055.0 58755.0 69710.0 ;
      RECT  58050.0 71055.0 58755.0 72400.0 ;
      RECT  58050.0 73745.0 58755.0 72400.0 ;
      RECT  58050.0 73745.0 58755.0 75090.0 ;
      RECT  58050.0 76435.0 58755.0 75090.0 ;
      RECT  58050.0 76435.0 58755.0 77780.0 ;
      RECT  58050.0 79125.0 58755.0 77780.0 ;
      RECT  58050.0 79125.0 58755.0 80470.0 ;
      RECT  58050.0 81815.0 58755.0 80470.0 ;
      RECT  58050.0 81815.0 58755.0 83160.0 ;
      RECT  58050.0 84505.0 58755.0 83160.0 ;
      RECT  58050.0 84505.0 58755.0 85850.0 ;
      RECT  58050.0 87195.0 58755.0 85850.0 ;
      RECT  58050.0 87195.0 58755.0 88540.0 ;
      RECT  58050.0 89885.0 58755.0 88540.0 ;
      RECT  58050.0 89885.0 58755.0 91230.0 ;
      RECT  58050.0 92575.0 58755.0 91230.0 ;
      RECT  58050.0 92575.0 58755.0 93920.0 ;
      RECT  58050.0 95265.0 58755.0 93920.0 ;
      RECT  58050.0 95265.0 58755.0 96610.0 ;
      RECT  58050.0 97955.0 58755.0 96610.0 ;
      RECT  58050.0 97955.0 58755.0 99300.0 ;
      RECT  58050.0 100645.0 58755.0 99300.0 ;
      RECT  58050.0 100645.0 58755.0 101990.0 ;
      RECT  58050.0 103335.0 58755.0 101990.0 ;
      RECT  58050.0 103335.0 58755.0 104680.0 ;
      RECT  58050.0 106025.0 58755.0 104680.0 ;
      RECT  58050.0 106025.0 58755.0 107370.0 ;
      RECT  58050.0 108715.0 58755.0 107370.0 ;
      RECT  58050.0 108715.0 58755.0 110060.0 ;
      RECT  58050.0 111405.0 58755.0 110060.0 ;
      RECT  58050.0 111405.0 58755.0 112750.0 ;
      RECT  58050.0 114095.0 58755.0 112750.0 ;
      RECT  58755.0 28015.0 59460.0 29360.0 ;
      RECT  58755.0 30705.0 59460.0 29360.0 ;
      RECT  58755.0 30705.0 59460.0 32050.0 ;
      RECT  58755.0 33395.0 59460.0 32050.0 ;
      RECT  58755.0 33395.0 59460.0 34740.0 ;
      RECT  58755.0 36085.0 59460.0 34740.0 ;
      RECT  58755.0 36085.0 59460.0 37430.0 ;
      RECT  58755.0 38775.0 59460.0 37430.0 ;
      RECT  58755.0 38775.0 59460.0 40120.0 ;
      RECT  58755.0 41465.0 59460.0 40120.0 ;
      RECT  58755.0 41465.0 59460.0 42810.0 ;
      RECT  58755.0 44155.0 59460.0 42810.0 ;
      RECT  58755.0 44155.0 59460.0 45500.0 ;
      RECT  58755.0 46845.0 59460.0 45500.0 ;
      RECT  58755.0 46845.0 59460.0 48190.0 ;
      RECT  58755.0 49535.0 59460.0 48190.0 ;
      RECT  58755.0 49535.0 59460.0 50880.0 ;
      RECT  58755.0 52225.0 59460.0 50880.0 ;
      RECT  58755.0 52225.0 59460.0 53570.0 ;
      RECT  58755.0 54915.0 59460.0 53570.0 ;
      RECT  58755.0 54915.0 59460.0 56260.0 ;
      RECT  58755.0 57605.0 59460.0 56260.0 ;
      RECT  58755.0 57605.0 59460.0 58950.0 ;
      RECT  58755.0 60295.0 59460.0 58950.0 ;
      RECT  58755.0 60295.0 59460.0 61640.0 ;
      RECT  58755.0 62985.0 59460.0 61640.0 ;
      RECT  58755.0 62985.0 59460.0 64330.0 ;
      RECT  58755.0 65675.0 59460.0 64330.0 ;
      RECT  58755.0 65675.0 59460.0 67020.0 ;
      RECT  58755.0 68365.0 59460.0 67020.0 ;
      RECT  58755.0 68365.0 59460.0 69710.0 ;
      RECT  58755.0 71055.0 59460.0 69710.0 ;
      RECT  58755.0 71055.0 59460.0 72400.0 ;
      RECT  58755.0 73745.0 59460.0 72400.0 ;
      RECT  58755.0 73745.0 59460.0 75090.0 ;
      RECT  58755.0 76435.0 59460.0 75090.0 ;
      RECT  58755.0 76435.0 59460.0 77780.0 ;
      RECT  58755.0 79125.0 59460.0 77780.0 ;
      RECT  58755.0 79125.0 59460.0 80470.0 ;
      RECT  58755.0 81815.0 59460.0 80470.0 ;
      RECT  58755.0 81815.0 59460.0 83160.0 ;
      RECT  58755.0 84505.0 59460.0 83160.0 ;
      RECT  58755.0 84505.0 59460.0 85850.0 ;
      RECT  58755.0 87195.0 59460.0 85850.0 ;
      RECT  58755.0 87195.0 59460.0 88540.0 ;
      RECT  58755.0 89885.0 59460.0 88540.0 ;
      RECT  58755.0 89885.0 59460.0 91230.0 ;
      RECT  58755.0 92575.0 59460.0 91230.0 ;
      RECT  58755.0 92575.0 59460.0 93920.0 ;
      RECT  58755.0 95265.0 59460.0 93920.0 ;
      RECT  58755.0 95265.0 59460.0 96610.0 ;
      RECT  58755.0 97955.0 59460.0 96610.0 ;
      RECT  58755.0 97955.0 59460.0 99300.0 ;
      RECT  58755.0 100645.0 59460.0 99300.0 ;
      RECT  58755.0 100645.0 59460.0 101990.0 ;
      RECT  58755.0 103335.0 59460.0 101990.0 ;
      RECT  58755.0 103335.0 59460.0 104680.0 ;
      RECT  58755.0 106025.0 59460.0 104680.0 ;
      RECT  58755.0 106025.0 59460.0 107370.0 ;
      RECT  58755.0 108715.0 59460.0 107370.0 ;
      RECT  58755.0 108715.0 59460.0 110060.0 ;
      RECT  58755.0 111405.0 59460.0 110060.0 ;
      RECT  58755.0 111405.0 59460.0 112750.0 ;
      RECT  58755.0 114095.0 59460.0 112750.0 ;
      RECT  59460.0 28015.0 60165.0 29360.0 ;
      RECT  59460.0 30705.0 60165.0 29360.0 ;
      RECT  59460.0 30705.0 60165.0 32050.0 ;
      RECT  59460.0 33395.0 60165.0 32050.0 ;
      RECT  59460.0 33395.0 60165.0 34740.0 ;
      RECT  59460.0 36085.0 60165.0 34740.0 ;
      RECT  59460.0 36085.0 60165.0 37430.0 ;
      RECT  59460.0 38775.0 60165.0 37430.0 ;
      RECT  59460.0 38775.0 60165.0 40120.0 ;
      RECT  59460.0 41465.0 60165.0 40120.0 ;
      RECT  59460.0 41465.0 60165.0 42810.0 ;
      RECT  59460.0 44155.0 60165.0 42810.0 ;
      RECT  59460.0 44155.0 60165.0 45500.0 ;
      RECT  59460.0 46845.0 60165.0 45500.0 ;
      RECT  59460.0 46845.0 60165.0 48190.0 ;
      RECT  59460.0 49535.0 60165.0 48190.0 ;
      RECT  59460.0 49535.0 60165.0 50880.0 ;
      RECT  59460.0 52225.0 60165.0 50880.0 ;
      RECT  59460.0 52225.0 60165.0 53570.0 ;
      RECT  59460.0 54915.0 60165.0 53570.0 ;
      RECT  59460.0 54915.0 60165.0 56260.0 ;
      RECT  59460.0 57605.0 60165.0 56260.0 ;
      RECT  59460.0 57605.0 60165.0 58950.0 ;
      RECT  59460.0 60295.0 60165.0 58950.0 ;
      RECT  59460.0 60295.0 60165.0 61640.0 ;
      RECT  59460.0 62985.0 60165.0 61640.0 ;
      RECT  59460.0 62985.0 60165.0 64330.0 ;
      RECT  59460.0 65675.0 60165.0 64330.0 ;
      RECT  59460.0 65675.0 60165.0 67020.0 ;
      RECT  59460.0 68365.0 60165.0 67020.0 ;
      RECT  59460.0 68365.0 60165.0 69710.0 ;
      RECT  59460.0 71055.0 60165.0 69710.0 ;
      RECT  59460.0 71055.0 60165.0 72400.0 ;
      RECT  59460.0 73745.0 60165.0 72400.0 ;
      RECT  59460.0 73745.0 60165.0 75090.0 ;
      RECT  59460.0 76435.0 60165.0 75090.0 ;
      RECT  59460.0 76435.0 60165.0 77780.0 ;
      RECT  59460.0 79125.0 60165.0 77780.0 ;
      RECT  59460.0 79125.0 60165.0 80470.0 ;
      RECT  59460.0 81815.0 60165.0 80470.0 ;
      RECT  59460.0 81815.0 60165.0 83160.0 ;
      RECT  59460.0 84505.0 60165.0 83160.0 ;
      RECT  59460.0 84505.0 60165.0 85850.0 ;
      RECT  59460.0 87195.0 60165.0 85850.0 ;
      RECT  59460.0 87195.0 60165.0 88540.0 ;
      RECT  59460.0 89885.0 60165.0 88540.0 ;
      RECT  59460.0 89885.0 60165.0 91230.0 ;
      RECT  59460.0 92575.0 60165.0 91230.0 ;
      RECT  59460.0 92575.0 60165.0 93920.0 ;
      RECT  59460.0 95265.0 60165.0 93920.0 ;
      RECT  59460.0 95265.0 60165.0 96610.0 ;
      RECT  59460.0 97955.0 60165.0 96610.0 ;
      RECT  59460.0 97955.0 60165.0 99300.0 ;
      RECT  59460.0 100645.0 60165.0 99300.0 ;
      RECT  59460.0 100645.0 60165.0 101990.0 ;
      RECT  59460.0 103335.0 60165.0 101990.0 ;
      RECT  59460.0 103335.0 60165.0 104680.0 ;
      RECT  59460.0 106025.0 60165.0 104680.0 ;
      RECT  59460.0 106025.0 60165.0 107370.0 ;
      RECT  59460.0 108715.0 60165.0 107370.0 ;
      RECT  59460.0 108715.0 60165.0 110060.0 ;
      RECT  59460.0 111405.0 60165.0 110060.0 ;
      RECT  59460.0 111405.0 60165.0 112750.0 ;
      RECT  59460.0 114095.0 60165.0 112750.0 ;
      RECT  60165.0 28015.0 60870.0 29360.0 ;
      RECT  60165.0 30705.0 60870.0 29360.0 ;
      RECT  60165.0 30705.0 60870.0 32050.0 ;
      RECT  60165.0 33395.0 60870.0 32050.0 ;
      RECT  60165.0 33395.0 60870.0 34740.0 ;
      RECT  60165.0 36085.0 60870.0 34740.0 ;
      RECT  60165.0 36085.0 60870.0 37430.0 ;
      RECT  60165.0 38775.0 60870.0 37430.0 ;
      RECT  60165.0 38775.0 60870.0 40120.0 ;
      RECT  60165.0 41465.0 60870.0 40120.0 ;
      RECT  60165.0 41465.0 60870.0 42810.0 ;
      RECT  60165.0 44155.0 60870.0 42810.0 ;
      RECT  60165.0 44155.0 60870.0 45500.0 ;
      RECT  60165.0 46845.0 60870.0 45500.0 ;
      RECT  60165.0 46845.0 60870.0 48190.0 ;
      RECT  60165.0 49535.0 60870.0 48190.0 ;
      RECT  60165.0 49535.0 60870.0 50880.0 ;
      RECT  60165.0 52225.0 60870.0 50880.0 ;
      RECT  60165.0 52225.0 60870.0 53570.0 ;
      RECT  60165.0 54915.0 60870.0 53570.0 ;
      RECT  60165.0 54915.0 60870.0 56260.0 ;
      RECT  60165.0 57605.0 60870.0 56260.0 ;
      RECT  60165.0 57605.0 60870.0 58950.0 ;
      RECT  60165.0 60295.0 60870.0 58950.0 ;
      RECT  60165.0 60295.0 60870.0 61640.0 ;
      RECT  60165.0 62985.0 60870.0 61640.0 ;
      RECT  60165.0 62985.0 60870.0 64330.0 ;
      RECT  60165.0 65675.0 60870.0 64330.0 ;
      RECT  60165.0 65675.0 60870.0 67020.0 ;
      RECT  60165.0 68365.0 60870.0 67020.0 ;
      RECT  60165.0 68365.0 60870.0 69710.0 ;
      RECT  60165.0 71055.0 60870.0 69710.0 ;
      RECT  60165.0 71055.0 60870.0 72400.0 ;
      RECT  60165.0 73745.0 60870.0 72400.0 ;
      RECT  60165.0 73745.0 60870.0 75090.0 ;
      RECT  60165.0 76435.0 60870.0 75090.0 ;
      RECT  60165.0 76435.0 60870.0 77780.0 ;
      RECT  60165.0 79125.0 60870.0 77780.0 ;
      RECT  60165.0 79125.0 60870.0 80470.0 ;
      RECT  60165.0 81815.0 60870.0 80470.0 ;
      RECT  60165.0 81815.0 60870.0 83160.0 ;
      RECT  60165.0 84505.0 60870.0 83160.0 ;
      RECT  60165.0 84505.0 60870.0 85850.0 ;
      RECT  60165.0 87195.0 60870.0 85850.0 ;
      RECT  60165.0 87195.0 60870.0 88540.0 ;
      RECT  60165.0 89885.0 60870.0 88540.0 ;
      RECT  60165.0 89885.0 60870.0 91230.0 ;
      RECT  60165.0 92575.0 60870.0 91230.0 ;
      RECT  60165.0 92575.0 60870.0 93920.0 ;
      RECT  60165.0 95265.0 60870.0 93920.0 ;
      RECT  60165.0 95265.0 60870.0 96610.0 ;
      RECT  60165.0 97955.0 60870.0 96610.0 ;
      RECT  60165.0 97955.0 60870.0 99300.0 ;
      RECT  60165.0 100645.0 60870.0 99300.0 ;
      RECT  60165.0 100645.0 60870.0 101990.0 ;
      RECT  60165.0 103335.0 60870.0 101990.0 ;
      RECT  60165.0 103335.0 60870.0 104680.0 ;
      RECT  60165.0 106025.0 60870.0 104680.0 ;
      RECT  60165.0 106025.0 60870.0 107370.0 ;
      RECT  60165.0 108715.0 60870.0 107370.0 ;
      RECT  60165.0 108715.0 60870.0 110060.0 ;
      RECT  60165.0 111405.0 60870.0 110060.0 ;
      RECT  60165.0 111405.0 60870.0 112750.0 ;
      RECT  60165.0 114095.0 60870.0 112750.0 ;
      RECT  60870.0 28015.0 61575.0 29360.0 ;
      RECT  60870.0 30705.0 61575.0 29360.0 ;
      RECT  60870.0 30705.0 61575.0 32050.0 ;
      RECT  60870.0 33395.0 61575.0 32050.0 ;
      RECT  60870.0 33395.0 61575.0 34740.0 ;
      RECT  60870.0 36085.0 61575.0 34740.0 ;
      RECT  60870.0 36085.0 61575.0 37430.0 ;
      RECT  60870.0 38775.0 61575.0 37430.0 ;
      RECT  60870.0 38775.0 61575.0 40120.0 ;
      RECT  60870.0 41465.0 61575.0 40120.0 ;
      RECT  60870.0 41465.0 61575.0 42810.0 ;
      RECT  60870.0 44155.0 61575.0 42810.0 ;
      RECT  60870.0 44155.0 61575.0 45500.0 ;
      RECT  60870.0 46845.0 61575.0 45500.0 ;
      RECT  60870.0 46845.0 61575.0 48190.0 ;
      RECT  60870.0 49535.0 61575.0 48190.0 ;
      RECT  60870.0 49535.0 61575.0 50880.0 ;
      RECT  60870.0 52225.0 61575.0 50880.0 ;
      RECT  60870.0 52225.0 61575.0 53570.0 ;
      RECT  60870.0 54915.0 61575.0 53570.0 ;
      RECT  60870.0 54915.0 61575.0 56260.0 ;
      RECT  60870.0 57605.0 61575.0 56260.0 ;
      RECT  60870.0 57605.0 61575.0 58950.0 ;
      RECT  60870.0 60295.0 61575.0 58950.0 ;
      RECT  60870.0 60295.0 61575.0 61640.0 ;
      RECT  60870.0 62985.0 61575.0 61640.0 ;
      RECT  60870.0 62985.0 61575.0 64330.0 ;
      RECT  60870.0 65675.0 61575.0 64330.0 ;
      RECT  60870.0 65675.0 61575.0 67020.0 ;
      RECT  60870.0 68365.0 61575.0 67020.0 ;
      RECT  60870.0 68365.0 61575.0 69710.0 ;
      RECT  60870.0 71055.0 61575.0 69710.0 ;
      RECT  60870.0 71055.0 61575.0 72400.0 ;
      RECT  60870.0 73745.0 61575.0 72400.0 ;
      RECT  60870.0 73745.0 61575.0 75090.0 ;
      RECT  60870.0 76435.0 61575.0 75090.0 ;
      RECT  60870.0 76435.0 61575.0 77780.0 ;
      RECT  60870.0 79125.0 61575.0 77780.0 ;
      RECT  60870.0 79125.0 61575.0 80470.0 ;
      RECT  60870.0 81815.0 61575.0 80470.0 ;
      RECT  60870.0 81815.0 61575.0 83160.0 ;
      RECT  60870.0 84505.0 61575.0 83160.0 ;
      RECT  60870.0 84505.0 61575.0 85850.0 ;
      RECT  60870.0 87195.0 61575.0 85850.0 ;
      RECT  60870.0 87195.0 61575.0 88540.0 ;
      RECT  60870.0 89885.0 61575.0 88540.0 ;
      RECT  60870.0 89885.0 61575.0 91230.0 ;
      RECT  60870.0 92575.0 61575.0 91230.0 ;
      RECT  60870.0 92575.0 61575.0 93920.0 ;
      RECT  60870.0 95265.0 61575.0 93920.0 ;
      RECT  60870.0 95265.0 61575.0 96610.0 ;
      RECT  60870.0 97955.0 61575.0 96610.0 ;
      RECT  60870.0 97955.0 61575.0 99300.0 ;
      RECT  60870.0 100645.0 61575.0 99300.0 ;
      RECT  60870.0 100645.0 61575.0 101990.0 ;
      RECT  60870.0 103335.0 61575.0 101990.0 ;
      RECT  60870.0 103335.0 61575.0 104680.0 ;
      RECT  60870.0 106025.0 61575.0 104680.0 ;
      RECT  60870.0 106025.0 61575.0 107370.0 ;
      RECT  60870.0 108715.0 61575.0 107370.0 ;
      RECT  60870.0 108715.0 61575.0 110060.0 ;
      RECT  60870.0 111405.0 61575.0 110060.0 ;
      RECT  60870.0 111405.0 61575.0 112750.0 ;
      RECT  60870.0 114095.0 61575.0 112750.0 ;
      RECT  61575.0 28015.0 62280.0 29360.0 ;
      RECT  61575.0 30705.0 62280.0 29360.0 ;
      RECT  61575.0 30705.0 62280.0 32050.0 ;
      RECT  61575.0 33395.0 62280.0 32050.0 ;
      RECT  61575.0 33395.0 62280.0 34740.0 ;
      RECT  61575.0 36085.0 62280.0 34740.0 ;
      RECT  61575.0 36085.0 62280.0 37430.0 ;
      RECT  61575.0 38775.0 62280.0 37430.0 ;
      RECT  61575.0 38775.0 62280.0 40120.0 ;
      RECT  61575.0 41465.0 62280.0 40120.0 ;
      RECT  61575.0 41465.0 62280.0 42810.0 ;
      RECT  61575.0 44155.0 62280.0 42810.0 ;
      RECT  61575.0 44155.0 62280.0 45500.0 ;
      RECT  61575.0 46845.0 62280.0 45500.0 ;
      RECT  61575.0 46845.0 62280.0 48190.0 ;
      RECT  61575.0 49535.0 62280.0 48190.0 ;
      RECT  61575.0 49535.0 62280.0 50880.0 ;
      RECT  61575.0 52225.0 62280.0 50880.0 ;
      RECT  61575.0 52225.0 62280.0 53570.0 ;
      RECT  61575.0 54915.0 62280.0 53570.0 ;
      RECT  61575.0 54915.0 62280.0 56260.0 ;
      RECT  61575.0 57605.0 62280.0 56260.0 ;
      RECT  61575.0 57605.0 62280.0 58950.0 ;
      RECT  61575.0 60295.0 62280.0 58950.0 ;
      RECT  61575.0 60295.0 62280.0 61640.0 ;
      RECT  61575.0 62985.0 62280.0 61640.0 ;
      RECT  61575.0 62985.0 62280.0 64330.0 ;
      RECT  61575.0 65675.0 62280.0 64330.0 ;
      RECT  61575.0 65675.0 62280.0 67020.0 ;
      RECT  61575.0 68365.0 62280.0 67020.0 ;
      RECT  61575.0 68365.0 62280.0 69710.0 ;
      RECT  61575.0 71055.0 62280.0 69710.0 ;
      RECT  61575.0 71055.0 62280.0 72400.0 ;
      RECT  61575.0 73745.0 62280.0 72400.0 ;
      RECT  61575.0 73745.0 62280.0 75090.0 ;
      RECT  61575.0 76435.0 62280.0 75090.0 ;
      RECT  61575.0 76435.0 62280.0 77780.0 ;
      RECT  61575.0 79125.0 62280.0 77780.0 ;
      RECT  61575.0 79125.0 62280.0 80470.0 ;
      RECT  61575.0 81815.0 62280.0 80470.0 ;
      RECT  61575.0 81815.0 62280.0 83160.0 ;
      RECT  61575.0 84505.0 62280.0 83160.0 ;
      RECT  61575.0 84505.0 62280.0 85850.0 ;
      RECT  61575.0 87195.0 62280.0 85850.0 ;
      RECT  61575.0 87195.0 62280.0 88540.0 ;
      RECT  61575.0 89885.0 62280.0 88540.0 ;
      RECT  61575.0 89885.0 62280.0 91230.0 ;
      RECT  61575.0 92575.0 62280.0 91230.0 ;
      RECT  61575.0 92575.0 62280.0 93920.0 ;
      RECT  61575.0 95265.0 62280.0 93920.0 ;
      RECT  61575.0 95265.0 62280.0 96610.0 ;
      RECT  61575.0 97955.0 62280.0 96610.0 ;
      RECT  61575.0 97955.0 62280.0 99300.0 ;
      RECT  61575.0 100645.0 62280.0 99300.0 ;
      RECT  61575.0 100645.0 62280.0 101990.0 ;
      RECT  61575.0 103335.0 62280.0 101990.0 ;
      RECT  61575.0 103335.0 62280.0 104680.0 ;
      RECT  61575.0 106025.0 62280.0 104680.0 ;
      RECT  61575.0 106025.0 62280.0 107370.0 ;
      RECT  61575.0 108715.0 62280.0 107370.0 ;
      RECT  61575.0 108715.0 62280.0 110060.0 ;
      RECT  61575.0 111405.0 62280.0 110060.0 ;
      RECT  61575.0 111405.0 62280.0 112750.0 ;
      RECT  61575.0 114095.0 62280.0 112750.0 ;
      RECT  62280.0 28015.0 62985.0 29360.0 ;
      RECT  62280.0 30705.0 62985.0 29360.0 ;
      RECT  62280.0 30705.0 62985.0 32050.0 ;
      RECT  62280.0 33395.0 62985.0 32050.0 ;
      RECT  62280.0 33395.0 62985.0 34740.0 ;
      RECT  62280.0 36085.0 62985.0 34740.0 ;
      RECT  62280.0 36085.0 62985.0 37430.0 ;
      RECT  62280.0 38775.0 62985.0 37430.0 ;
      RECT  62280.0 38775.0 62985.0 40120.0 ;
      RECT  62280.0 41465.0 62985.0 40120.0 ;
      RECT  62280.0 41465.0 62985.0 42810.0 ;
      RECT  62280.0 44155.0 62985.0 42810.0 ;
      RECT  62280.0 44155.0 62985.0 45500.0 ;
      RECT  62280.0 46845.0 62985.0 45500.0 ;
      RECT  62280.0 46845.0 62985.0 48190.0 ;
      RECT  62280.0 49535.0 62985.0 48190.0 ;
      RECT  62280.0 49535.0 62985.0 50880.0 ;
      RECT  62280.0 52225.0 62985.0 50880.0 ;
      RECT  62280.0 52225.0 62985.0 53570.0 ;
      RECT  62280.0 54915.0 62985.0 53570.0 ;
      RECT  62280.0 54915.0 62985.0 56260.0 ;
      RECT  62280.0 57605.0 62985.0 56260.0 ;
      RECT  62280.0 57605.0 62985.0 58950.0 ;
      RECT  62280.0 60295.0 62985.0 58950.0 ;
      RECT  62280.0 60295.0 62985.0 61640.0 ;
      RECT  62280.0 62985.0 62985.0 61640.0 ;
      RECT  62280.0 62985.0 62985.0 64330.0 ;
      RECT  62280.0 65675.0 62985.0 64330.0 ;
      RECT  62280.0 65675.0 62985.0 67020.0 ;
      RECT  62280.0 68365.0 62985.0 67020.0 ;
      RECT  62280.0 68365.0 62985.0 69710.0 ;
      RECT  62280.0 71055.0 62985.0 69710.0 ;
      RECT  62280.0 71055.0 62985.0 72400.0 ;
      RECT  62280.0 73745.0 62985.0 72400.0 ;
      RECT  62280.0 73745.0 62985.0 75090.0 ;
      RECT  62280.0 76435.0 62985.0 75090.0 ;
      RECT  62280.0 76435.0 62985.0 77780.0 ;
      RECT  62280.0 79125.0 62985.0 77780.0 ;
      RECT  62280.0 79125.0 62985.0 80470.0 ;
      RECT  62280.0 81815.0 62985.0 80470.0 ;
      RECT  62280.0 81815.0 62985.0 83160.0 ;
      RECT  62280.0 84505.0 62985.0 83160.0 ;
      RECT  62280.0 84505.0 62985.0 85850.0 ;
      RECT  62280.0 87195.0 62985.0 85850.0 ;
      RECT  62280.0 87195.0 62985.0 88540.0 ;
      RECT  62280.0 89885.0 62985.0 88540.0 ;
      RECT  62280.0 89885.0 62985.0 91230.0 ;
      RECT  62280.0 92575.0 62985.0 91230.0 ;
      RECT  62280.0 92575.0 62985.0 93920.0 ;
      RECT  62280.0 95265.0 62985.0 93920.0 ;
      RECT  62280.0 95265.0 62985.0 96610.0 ;
      RECT  62280.0 97955.0 62985.0 96610.0 ;
      RECT  62280.0 97955.0 62985.0 99300.0 ;
      RECT  62280.0 100645.0 62985.0 99300.0 ;
      RECT  62280.0 100645.0 62985.0 101990.0 ;
      RECT  62280.0 103335.0 62985.0 101990.0 ;
      RECT  62280.0 103335.0 62985.0 104680.0 ;
      RECT  62280.0 106025.0 62985.0 104680.0 ;
      RECT  62280.0 106025.0 62985.0 107370.0 ;
      RECT  62280.0 108715.0 62985.0 107370.0 ;
      RECT  62280.0 108715.0 62985.0 110060.0 ;
      RECT  62280.0 111405.0 62985.0 110060.0 ;
      RECT  62280.0 111405.0 62985.0 112750.0 ;
      RECT  62280.0 114095.0 62985.0 112750.0 ;
      RECT  62985.0 28015.0 63690.0 29360.0 ;
      RECT  62985.0 30705.0 63690.0 29360.0 ;
      RECT  62985.0 30705.0 63690.0 32050.0 ;
      RECT  62985.0 33395.0 63690.0 32050.0 ;
      RECT  62985.0 33395.0 63690.0 34740.0 ;
      RECT  62985.0 36085.0 63690.0 34740.0 ;
      RECT  62985.0 36085.0 63690.0 37430.0 ;
      RECT  62985.0 38775.0 63690.0 37430.0 ;
      RECT  62985.0 38775.0 63690.0 40120.0 ;
      RECT  62985.0 41465.0 63690.0 40120.0 ;
      RECT  62985.0 41465.0 63690.0 42810.0 ;
      RECT  62985.0 44155.0 63690.0 42810.0 ;
      RECT  62985.0 44155.0 63690.0 45500.0 ;
      RECT  62985.0 46845.0 63690.0 45500.0 ;
      RECT  62985.0 46845.0 63690.0 48190.0 ;
      RECT  62985.0 49535.0 63690.0 48190.0 ;
      RECT  62985.0 49535.0 63690.0 50880.0 ;
      RECT  62985.0 52225.0 63690.0 50880.0 ;
      RECT  62985.0 52225.0 63690.0 53570.0 ;
      RECT  62985.0 54915.0 63690.0 53570.0 ;
      RECT  62985.0 54915.0 63690.0 56260.0 ;
      RECT  62985.0 57605.0 63690.0 56260.0 ;
      RECT  62985.0 57605.0 63690.0 58950.0 ;
      RECT  62985.0 60295.0 63690.0 58950.0 ;
      RECT  62985.0 60295.0 63690.0 61640.0 ;
      RECT  62985.0 62985.0 63690.0 61640.0 ;
      RECT  62985.0 62985.0 63690.0 64330.0 ;
      RECT  62985.0 65675.0 63690.0 64330.0 ;
      RECT  62985.0 65675.0 63690.0 67020.0 ;
      RECT  62985.0 68365.0 63690.0 67020.0 ;
      RECT  62985.0 68365.0 63690.0 69710.0 ;
      RECT  62985.0 71055.0 63690.0 69710.0 ;
      RECT  62985.0 71055.0 63690.0 72400.0 ;
      RECT  62985.0 73745.0 63690.0 72400.0 ;
      RECT  62985.0 73745.0 63690.0 75090.0 ;
      RECT  62985.0 76435.0 63690.0 75090.0 ;
      RECT  62985.0 76435.0 63690.0 77780.0 ;
      RECT  62985.0 79125.0 63690.0 77780.0 ;
      RECT  62985.0 79125.0 63690.0 80470.0 ;
      RECT  62985.0 81815.0 63690.0 80470.0 ;
      RECT  62985.0 81815.0 63690.0 83160.0 ;
      RECT  62985.0 84505.0 63690.0 83160.0 ;
      RECT  62985.0 84505.0 63690.0 85850.0 ;
      RECT  62985.0 87195.0 63690.0 85850.0 ;
      RECT  62985.0 87195.0 63690.0 88540.0 ;
      RECT  62985.0 89885.0 63690.0 88540.0 ;
      RECT  62985.0 89885.0 63690.0 91230.0 ;
      RECT  62985.0 92575.0 63690.0 91230.0 ;
      RECT  62985.0 92575.0 63690.0 93920.0 ;
      RECT  62985.0 95265.0 63690.0 93920.0 ;
      RECT  62985.0 95265.0 63690.0 96610.0 ;
      RECT  62985.0 97955.0 63690.0 96610.0 ;
      RECT  62985.0 97955.0 63690.0 99300.0 ;
      RECT  62985.0 100645.0 63690.0 99300.0 ;
      RECT  62985.0 100645.0 63690.0 101990.0 ;
      RECT  62985.0 103335.0 63690.0 101990.0 ;
      RECT  62985.0 103335.0 63690.0 104680.0 ;
      RECT  62985.0 106025.0 63690.0 104680.0 ;
      RECT  62985.0 106025.0 63690.0 107370.0 ;
      RECT  62985.0 108715.0 63690.0 107370.0 ;
      RECT  62985.0 108715.0 63690.0 110060.0 ;
      RECT  62985.0 111405.0 63690.0 110060.0 ;
      RECT  62985.0 111405.0 63690.0 112750.0 ;
      RECT  62985.0 114095.0 63690.0 112750.0 ;
      RECT  63690.0 28015.0 64395.0 29360.0 ;
      RECT  63690.0 30705.0 64395.0 29360.0 ;
      RECT  63690.0 30705.0 64395.0 32050.0 ;
      RECT  63690.0 33395.0 64395.0 32050.0 ;
      RECT  63690.0 33395.0 64395.0 34740.0 ;
      RECT  63690.0 36085.0 64395.0 34740.0 ;
      RECT  63690.0 36085.0 64395.0 37430.0 ;
      RECT  63690.0 38775.0 64395.0 37430.0 ;
      RECT  63690.0 38775.0 64395.0 40120.0 ;
      RECT  63690.0 41465.0 64395.0 40120.0 ;
      RECT  63690.0 41465.0 64395.0 42810.0 ;
      RECT  63690.0 44155.0 64395.0 42810.0 ;
      RECT  63690.0 44155.0 64395.0 45500.0 ;
      RECT  63690.0 46845.0 64395.0 45500.0 ;
      RECT  63690.0 46845.0 64395.0 48190.0 ;
      RECT  63690.0 49535.0 64395.0 48190.0 ;
      RECT  63690.0 49535.0 64395.0 50880.0 ;
      RECT  63690.0 52225.0 64395.0 50880.0 ;
      RECT  63690.0 52225.0 64395.0 53570.0 ;
      RECT  63690.0 54915.0 64395.0 53570.0 ;
      RECT  63690.0 54915.0 64395.0 56260.0 ;
      RECT  63690.0 57605.0 64395.0 56260.0 ;
      RECT  63690.0 57605.0 64395.0 58950.0 ;
      RECT  63690.0 60295.0 64395.0 58950.0 ;
      RECT  63690.0 60295.0 64395.0 61640.0 ;
      RECT  63690.0 62985.0 64395.0 61640.0 ;
      RECT  63690.0 62985.0 64395.0 64330.0 ;
      RECT  63690.0 65675.0 64395.0 64330.0 ;
      RECT  63690.0 65675.0 64395.0 67020.0 ;
      RECT  63690.0 68365.0 64395.0 67020.0 ;
      RECT  63690.0 68365.0 64395.0 69710.0 ;
      RECT  63690.0 71055.0 64395.0 69710.0 ;
      RECT  63690.0 71055.0 64395.0 72400.0 ;
      RECT  63690.0 73745.0 64395.0 72400.0 ;
      RECT  63690.0 73745.0 64395.0 75090.0 ;
      RECT  63690.0 76435.0 64395.0 75090.0 ;
      RECT  63690.0 76435.0 64395.0 77780.0 ;
      RECT  63690.0 79125.0 64395.0 77780.0 ;
      RECT  63690.0 79125.0 64395.0 80470.0 ;
      RECT  63690.0 81815.0 64395.0 80470.0 ;
      RECT  63690.0 81815.0 64395.0 83160.0 ;
      RECT  63690.0 84505.0 64395.0 83160.0 ;
      RECT  63690.0 84505.0 64395.0 85850.0 ;
      RECT  63690.0 87195.0 64395.0 85850.0 ;
      RECT  63690.0 87195.0 64395.0 88540.0 ;
      RECT  63690.0 89885.0 64395.0 88540.0 ;
      RECT  63690.0 89885.0 64395.0 91230.0 ;
      RECT  63690.0 92575.0 64395.0 91230.0 ;
      RECT  63690.0 92575.0 64395.0 93920.0 ;
      RECT  63690.0 95265.0 64395.0 93920.0 ;
      RECT  63690.0 95265.0 64395.0 96610.0 ;
      RECT  63690.0 97955.0 64395.0 96610.0 ;
      RECT  63690.0 97955.0 64395.0 99300.0 ;
      RECT  63690.0 100645.0 64395.0 99300.0 ;
      RECT  63690.0 100645.0 64395.0 101990.0 ;
      RECT  63690.0 103335.0 64395.0 101990.0 ;
      RECT  63690.0 103335.0 64395.0 104680.0 ;
      RECT  63690.0 106025.0 64395.0 104680.0 ;
      RECT  63690.0 106025.0 64395.0 107370.0 ;
      RECT  63690.0 108715.0 64395.0 107370.0 ;
      RECT  63690.0 108715.0 64395.0 110060.0 ;
      RECT  63690.0 111405.0 64395.0 110060.0 ;
      RECT  63690.0 111405.0 64395.0 112750.0 ;
      RECT  63690.0 114095.0 64395.0 112750.0 ;
      RECT  64395.0 28015.0 65100.0 29360.0 ;
      RECT  64395.0 30705.0 65100.0 29360.0 ;
      RECT  64395.0 30705.0 65100.0 32050.0 ;
      RECT  64395.0 33395.0 65100.0 32050.0 ;
      RECT  64395.0 33395.0 65100.0 34740.0 ;
      RECT  64395.0 36085.0 65100.0 34740.0 ;
      RECT  64395.0 36085.0 65100.0 37430.0 ;
      RECT  64395.0 38775.0 65100.0 37430.0 ;
      RECT  64395.0 38775.0 65100.0 40120.0 ;
      RECT  64395.0 41465.0 65100.0 40120.0 ;
      RECT  64395.0 41465.0 65100.0 42810.0 ;
      RECT  64395.0 44155.0 65100.0 42810.0 ;
      RECT  64395.0 44155.0 65100.0 45500.0 ;
      RECT  64395.0 46845.0 65100.0 45500.0 ;
      RECT  64395.0 46845.0 65100.0 48190.0 ;
      RECT  64395.0 49535.0 65100.0 48190.0 ;
      RECT  64395.0 49535.0 65100.0 50880.0 ;
      RECT  64395.0 52225.0 65100.0 50880.0 ;
      RECT  64395.0 52225.0 65100.0 53570.0 ;
      RECT  64395.0 54915.0 65100.0 53570.0 ;
      RECT  64395.0 54915.0 65100.0 56260.0 ;
      RECT  64395.0 57605.0 65100.0 56260.0 ;
      RECT  64395.0 57605.0 65100.0 58950.0 ;
      RECT  64395.0 60295.0 65100.0 58950.0 ;
      RECT  64395.0 60295.0 65100.0 61640.0 ;
      RECT  64395.0 62985.0 65100.0 61640.0 ;
      RECT  64395.0 62985.0 65100.0 64330.0 ;
      RECT  64395.0 65675.0 65100.0 64330.0 ;
      RECT  64395.0 65675.0 65100.0 67020.0 ;
      RECT  64395.0 68365.0 65100.0 67020.0 ;
      RECT  64395.0 68365.0 65100.0 69710.0 ;
      RECT  64395.0 71055.0 65100.0 69710.0 ;
      RECT  64395.0 71055.0 65100.0 72400.0 ;
      RECT  64395.0 73745.0 65100.0 72400.0 ;
      RECT  64395.0 73745.0 65100.0 75090.0 ;
      RECT  64395.0 76435.0 65100.0 75090.0 ;
      RECT  64395.0 76435.0 65100.0 77780.0 ;
      RECT  64395.0 79125.0 65100.0 77780.0 ;
      RECT  64395.0 79125.0 65100.0 80470.0 ;
      RECT  64395.0 81815.0 65100.0 80470.0 ;
      RECT  64395.0 81815.0 65100.0 83160.0 ;
      RECT  64395.0 84505.0 65100.0 83160.0 ;
      RECT  64395.0 84505.0 65100.0 85850.0 ;
      RECT  64395.0 87195.0 65100.0 85850.0 ;
      RECT  64395.0 87195.0 65100.0 88540.0 ;
      RECT  64395.0 89885.0 65100.0 88540.0 ;
      RECT  64395.0 89885.0 65100.0 91230.0 ;
      RECT  64395.0 92575.0 65100.0 91230.0 ;
      RECT  64395.0 92575.0 65100.0 93920.0 ;
      RECT  64395.0 95265.0 65100.0 93920.0 ;
      RECT  64395.0 95265.0 65100.0 96610.0 ;
      RECT  64395.0 97955.0 65100.0 96610.0 ;
      RECT  64395.0 97955.0 65100.0 99300.0 ;
      RECT  64395.0 100645.0 65100.0 99300.0 ;
      RECT  64395.0 100645.0 65100.0 101990.0 ;
      RECT  64395.0 103335.0 65100.0 101990.0 ;
      RECT  64395.0 103335.0 65100.0 104680.0 ;
      RECT  64395.0 106025.0 65100.0 104680.0 ;
      RECT  64395.0 106025.0 65100.0 107370.0 ;
      RECT  64395.0 108715.0 65100.0 107370.0 ;
      RECT  64395.0 108715.0 65100.0 110060.0 ;
      RECT  64395.0 111405.0 65100.0 110060.0 ;
      RECT  64395.0 111405.0 65100.0 112750.0 ;
      RECT  64395.0 114095.0 65100.0 112750.0 ;
      RECT  65100.0 28015.0 65805.0 29360.0 ;
      RECT  65100.0 30705.0 65805.0 29360.0 ;
      RECT  65100.0 30705.0 65805.0 32050.0 ;
      RECT  65100.0 33395.0 65805.0 32050.0 ;
      RECT  65100.0 33395.0 65805.0 34740.0 ;
      RECT  65100.0 36085.0 65805.0 34740.0 ;
      RECT  65100.0 36085.0 65805.0 37430.0 ;
      RECT  65100.0 38775.0 65805.0 37430.0 ;
      RECT  65100.0 38775.0 65805.0 40120.0 ;
      RECT  65100.0 41465.0 65805.0 40120.0 ;
      RECT  65100.0 41465.0 65805.0 42810.0 ;
      RECT  65100.0 44155.0 65805.0 42810.0 ;
      RECT  65100.0 44155.0 65805.0 45500.0 ;
      RECT  65100.0 46845.0 65805.0 45500.0 ;
      RECT  65100.0 46845.0 65805.0 48190.0 ;
      RECT  65100.0 49535.0 65805.0 48190.0 ;
      RECT  65100.0 49535.0 65805.0 50880.0 ;
      RECT  65100.0 52225.0 65805.0 50880.0 ;
      RECT  65100.0 52225.0 65805.0 53570.0 ;
      RECT  65100.0 54915.0 65805.0 53570.0 ;
      RECT  65100.0 54915.0 65805.0 56260.0 ;
      RECT  65100.0 57605.0 65805.0 56260.0 ;
      RECT  65100.0 57605.0 65805.0 58950.0 ;
      RECT  65100.0 60295.0 65805.0 58950.0 ;
      RECT  65100.0 60295.0 65805.0 61640.0 ;
      RECT  65100.0 62985.0 65805.0 61640.0 ;
      RECT  65100.0 62985.0 65805.0 64330.0 ;
      RECT  65100.0 65675.0 65805.0 64330.0 ;
      RECT  65100.0 65675.0 65805.0 67020.0 ;
      RECT  65100.0 68365.0 65805.0 67020.0 ;
      RECT  65100.0 68365.0 65805.0 69710.0 ;
      RECT  65100.0 71055.0 65805.0 69710.0 ;
      RECT  65100.0 71055.0 65805.0 72400.0 ;
      RECT  65100.0 73745.0 65805.0 72400.0 ;
      RECT  65100.0 73745.0 65805.0 75090.0 ;
      RECT  65100.0 76435.0 65805.0 75090.0 ;
      RECT  65100.0 76435.0 65805.0 77780.0 ;
      RECT  65100.0 79125.0 65805.0 77780.0 ;
      RECT  65100.0 79125.0 65805.0 80470.0 ;
      RECT  65100.0 81815.0 65805.0 80470.0 ;
      RECT  65100.0 81815.0 65805.0 83160.0 ;
      RECT  65100.0 84505.0 65805.0 83160.0 ;
      RECT  65100.0 84505.0 65805.0 85850.0 ;
      RECT  65100.0 87195.0 65805.0 85850.0 ;
      RECT  65100.0 87195.0 65805.0 88540.0 ;
      RECT  65100.0 89885.0 65805.0 88540.0 ;
      RECT  65100.0 89885.0 65805.0 91230.0 ;
      RECT  65100.0 92575.0 65805.0 91230.0 ;
      RECT  65100.0 92575.0 65805.0 93920.0 ;
      RECT  65100.0 95265.0 65805.0 93920.0 ;
      RECT  65100.0 95265.0 65805.0 96610.0 ;
      RECT  65100.0 97955.0 65805.0 96610.0 ;
      RECT  65100.0 97955.0 65805.0 99300.0 ;
      RECT  65100.0 100645.0 65805.0 99300.0 ;
      RECT  65100.0 100645.0 65805.0 101990.0 ;
      RECT  65100.0 103335.0 65805.0 101990.0 ;
      RECT  65100.0 103335.0 65805.0 104680.0 ;
      RECT  65100.0 106025.0 65805.0 104680.0 ;
      RECT  65100.0 106025.0 65805.0 107370.0 ;
      RECT  65100.0 108715.0 65805.0 107370.0 ;
      RECT  65100.0 108715.0 65805.0 110060.0 ;
      RECT  65100.0 111405.0 65805.0 110060.0 ;
      RECT  65100.0 111405.0 65805.0 112750.0 ;
      RECT  65100.0 114095.0 65805.0 112750.0 ;
      RECT  65805.0 28015.0 66510.0 29360.0 ;
      RECT  65805.0 30705.0 66510.0 29360.0 ;
      RECT  65805.0 30705.0 66510.0 32050.0 ;
      RECT  65805.0 33395.0 66510.0 32050.0 ;
      RECT  65805.0 33395.0 66510.0 34740.0 ;
      RECT  65805.0 36085.0 66510.0 34740.0 ;
      RECT  65805.0 36085.0 66510.0 37430.0 ;
      RECT  65805.0 38775.0 66510.0 37430.0 ;
      RECT  65805.0 38775.0 66510.0 40120.0 ;
      RECT  65805.0 41465.0 66510.0 40120.0 ;
      RECT  65805.0 41465.0 66510.0 42810.0 ;
      RECT  65805.0 44155.0 66510.0 42810.0 ;
      RECT  65805.0 44155.0 66510.0 45500.0 ;
      RECT  65805.0 46845.0 66510.0 45500.0 ;
      RECT  65805.0 46845.0 66510.0 48190.0 ;
      RECT  65805.0 49535.0 66510.0 48190.0 ;
      RECT  65805.0 49535.0 66510.0 50880.0 ;
      RECT  65805.0 52225.0 66510.0 50880.0 ;
      RECT  65805.0 52225.0 66510.0 53570.0 ;
      RECT  65805.0 54915.0 66510.0 53570.0 ;
      RECT  65805.0 54915.0 66510.0 56260.0 ;
      RECT  65805.0 57605.0 66510.0 56260.0 ;
      RECT  65805.0 57605.0 66510.0 58950.0 ;
      RECT  65805.0 60295.0 66510.0 58950.0 ;
      RECT  65805.0 60295.0 66510.0 61640.0 ;
      RECT  65805.0 62985.0 66510.0 61640.0 ;
      RECT  65805.0 62985.0 66510.0 64330.0 ;
      RECT  65805.0 65675.0 66510.0 64330.0 ;
      RECT  65805.0 65675.0 66510.0 67020.0 ;
      RECT  65805.0 68365.0 66510.0 67020.0 ;
      RECT  65805.0 68365.0 66510.0 69710.0 ;
      RECT  65805.0 71055.0 66510.0 69710.0 ;
      RECT  65805.0 71055.0 66510.0 72400.0 ;
      RECT  65805.0 73745.0 66510.0 72400.0 ;
      RECT  65805.0 73745.0 66510.0 75090.0 ;
      RECT  65805.0 76435.0 66510.0 75090.0 ;
      RECT  65805.0 76435.0 66510.0 77780.0 ;
      RECT  65805.0 79125.0 66510.0 77780.0 ;
      RECT  65805.0 79125.0 66510.0 80470.0 ;
      RECT  65805.0 81815.0 66510.0 80470.0 ;
      RECT  65805.0 81815.0 66510.0 83160.0 ;
      RECT  65805.0 84505.0 66510.0 83160.0 ;
      RECT  65805.0 84505.0 66510.0 85850.0 ;
      RECT  65805.0 87195.0 66510.0 85850.0 ;
      RECT  65805.0 87195.0 66510.0 88540.0 ;
      RECT  65805.0 89885.0 66510.0 88540.0 ;
      RECT  65805.0 89885.0 66510.0 91230.0 ;
      RECT  65805.0 92575.0 66510.0 91230.0 ;
      RECT  65805.0 92575.0 66510.0 93920.0 ;
      RECT  65805.0 95265.0 66510.0 93920.0 ;
      RECT  65805.0 95265.0 66510.0 96610.0 ;
      RECT  65805.0 97955.0 66510.0 96610.0 ;
      RECT  65805.0 97955.0 66510.0 99300.0 ;
      RECT  65805.0 100645.0 66510.0 99300.0 ;
      RECT  65805.0 100645.0 66510.0 101990.0 ;
      RECT  65805.0 103335.0 66510.0 101990.0 ;
      RECT  65805.0 103335.0 66510.0 104680.0 ;
      RECT  65805.0 106025.0 66510.0 104680.0 ;
      RECT  65805.0 106025.0 66510.0 107370.0 ;
      RECT  65805.0 108715.0 66510.0 107370.0 ;
      RECT  65805.0 108715.0 66510.0 110060.0 ;
      RECT  65805.0 111405.0 66510.0 110060.0 ;
      RECT  65805.0 111405.0 66510.0 112750.0 ;
      RECT  65805.0 114095.0 66510.0 112750.0 ;
      RECT  66510.0 28015.0 67215.0 29360.0 ;
      RECT  66510.0 30705.0 67215.0 29360.0 ;
      RECT  66510.0 30705.0 67215.0 32050.0 ;
      RECT  66510.0 33395.0 67215.0 32050.0 ;
      RECT  66510.0 33395.0 67215.0 34740.0 ;
      RECT  66510.0 36085.0 67215.0 34740.0 ;
      RECT  66510.0 36085.0 67215.0 37430.0 ;
      RECT  66510.0 38775.0 67215.0 37430.0 ;
      RECT  66510.0 38775.0 67215.0 40120.0 ;
      RECT  66510.0 41465.0 67215.0 40120.0 ;
      RECT  66510.0 41465.0 67215.0 42810.0 ;
      RECT  66510.0 44155.0 67215.0 42810.0 ;
      RECT  66510.0 44155.0 67215.0 45500.0 ;
      RECT  66510.0 46845.0 67215.0 45500.0 ;
      RECT  66510.0 46845.0 67215.0 48190.0 ;
      RECT  66510.0 49535.0 67215.0 48190.0 ;
      RECT  66510.0 49535.0 67215.0 50880.0 ;
      RECT  66510.0 52225.0 67215.0 50880.0 ;
      RECT  66510.0 52225.0 67215.0 53570.0 ;
      RECT  66510.0 54915.0 67215.0 53570.0 ;
      RECT  66510.0 54915.0 67215.0 56260.0 ;
      RECT  66510.0 57605.0 67215.0 56260.0 ;
      RECT  66510.0 57605.0 67215.0 58950.0 ;
      RECT  66510.0 60295.0 67215.0 58950.0 ;
      RECT  66510.0 60295.0 67215.0 61640.0 ;
      RECT  66510.0 62985.0 67215.0 61640.0 ;
      RECT  66510.0 62985.0 67215.0 64330.0 ;
      RECT  66510.0 65675.0 67215.0 64330.0 ;
      RECT  66510.0 65675.0 67215.0 67020.0 ;
      RECT  66510.0 68365.0 67215.0 67020.0 ;
      RECT  66510.0 68365.0 67215.0 69710.0 ;
      RECT  66510.0 71055.0 67215.0 69710.0 ;
      RECT  66510.0 71055.0 67215.0 72400.0 ;
      RECT  66510.0 73745.0 67215.0 72400.0 ;
      RECT  66510.0 73745.0 67215.0 75090.0 ;
      RECT  66510.0 76435.0 67215.0 75090.0 ;
      RECT  66510.0 76435.0 67215.0 77780.0 ;
      RECT  66510.0 79125.0 67215.0 77780.0 ;
      RECT  66510.0 79125.0 67215.0 80470.0 ;
      RECT  66510.0 81815.0 67215.0 80470.0 ;
      RECT  66510.0 81815.0 67215.0 83160.0 ;
      RECT  66510.0 84505.0 67215.0 83160.0 ;
      RECT  66510.0 84505.0 67215.0 85850.0 ;
      RECT  66510.0 87195.0 67215.0 85850.0 ;
      RECT  66510.0 87195.0 67215.0 88540.0 ;
      RECT  66510.0 89885.0 67215.0 88540.0 ;
      RECT  66510.0 89885.0 67215.0 91230.0 ;
      RECT  66510.0 92575.0 67215.0 91230.0 ;
      RECT  66510.0 92575.0 67215.0 93920.0 ;
      RECT  66510.0 95265.0 67215.0 93920.0 ;
      RECT  66510.0 95265.0 67215.0 96610.0 ;
      RECT  66510.0 97955.0 67215.0 96610.0 ;
      RECT  66510.0 97955.0 67215.0 99300.0 ;
      RECT  66510.0 100645.0 67215.0 99300.0 ;
      RECT  66510.0 100645.0 67215.0 101990.0 ;
      RECT  66510.0 103335.0 67215.0 101990.0 ;
      RECT  66510.0 103335.0 67215.0 104680.0 ;
      RECT  66510.0 106025.0 67215.0 104680.0 ;
      RECT  66510.0 106025.0 67215.0 107370.0 ;
      RECT  66510.0 108715.0 67215.0 107370.0 ;
      RECT  66510.0 108715.0 67215.0 110060.0 ;
      RECT  66510.0 111405.0 67215.0 110060.0 ;
      RECT  66510.0 111405.0 67215.0 112750.0 ;
      RECT  66510.0 114095.0 67215.0 112750.0 ;
      RECT  67215.0 28015.0 67920.0 29360.0 ;
      RECT  67215.0 30705.0 67920.0 29360.0 ;
      RECT  67215.0 30705.0 67920.0 32050.0 ;
      RECT  67215.0 33395.0 67920.0 32050.0 ;
      RECT  67215.0 33395.0 67920.0 34740.0 ;
      RECT  67215.0 36085.0 67920.0 34740.0 ;
      RECT  67215.0 36085.0 67920.0 37430.0 ;
      RECT  67215.0 38775.0 67920.0 37430.0 ;
      RECT  67215.0 38775.0 67920.0 40120.0 ;
      RECT  67215.0 41465.0 67920.0 40120.0 ;
      RECT  67215.0 41465.0 67920.0 42810.0 ;
      RECT  67215.0 44155.0 67920.0 42810.0 ;
      RECT  67215.0 44155.0 67920.0 45500.0 ;
      RECT  67215.0 46845.0 67920.0 45500.0 ;
      RECT  67215.0 46845.0 67920.0 48190.0 ;
      RECT  67215.0 49535.0 67920.0 48190.0 ;
      RECT  67215.0 49535.0 67920.0 50880.0 ;
      RECT  67215.0 52225.0 67920.0 50880.0 ;
      RECT  67215.0 52225.0 67920.0 53570.0 ;
      RECT  67215.0 54915.0 67920.0 53570.0 ;
      RECT  67215.0 54915.0 67920.0 56260.0 ;
      RECT  67215.0 57605.0 67920.0 56260.0 ;
      RECT  67215.0 57605.0 67920.0 58950.0 ;
      RECT  67215.0 60295.0 67920.0 58950.0 ;
      RECT  67215.0 60295.0 67920.0 61640.0 ;
      RECT  67215.0 62985.0 67920.0 61640.0 ;
      RECT  67215.0 62985.0 67920.0 64330.0 ;
      RECT  67215.0 65675.0 67920.0 64330.0 ;
      RECT  67215.0 65675.0 67920.0 67020.0 ;
      RECT  67215.0 68365.0 67920.0 67020.0 ;
      RECT  67215.0 68365.0 67920.0 69710.0 ;
      RECT  67215.0 71055.0 67920.0 69710.0 ;
      RECT  67215.0 71055.0 67920.0 72400.0 ;
      RECT  67215.0 73745.0 67920.0 72400.0 ;
      RECT  67215.0 73745.0 67920.0 75090.0 ;
      RECT  67215.0 76435.0 67920.0 75090.0 ;
      RECT  67215.0 76435.0 67920.0 77780.0 ;
      RECT  67215.0 79125.0 67920.0 77780.0 ;
      RECT  67215.0 79125.0 67920.0 80470.0 ;
      RECT  67215.0 81815.0 67920.0 80470.0 ;
      RECT  67215.0 81815.0 67920.0 83160.0 ;
      RECT  67215.0 84505.0 67920.0 83160.0 ;
      RECT  67215.0 84505.0 67920.0 85850.0 ;
      RECT  67215.0 87195.0 67920.0 85850.0 ;
      RECT  67215.0 87195.0 67920.0 88540.0 ;
      RECT  67215.0 89885.0 67920.0 88540.0 ;
      RECT  67215.0 89885.0 67920.0 91230.0 ;
      RECT  67215.0 92575.0 67920.0 91230.0 ;
      RECT  67215.0 92575.0 67920.0 93920.0 ;
      RECT  67215.0 95265.0 67920.0 93920.0 ;
      RECT  67215.0 95265.0 67920.0 96610.0 ;
      RECT  67215.0 97955.0 67920.0 96610.0 ;
      RECT  67215.0 97955.0 67920.0 99300.0 ;
      RECT  67215.0 100645.0 67920.0 99300.0 ;
      RECT  67215.0 100645.0 67920.0 101990.0 ;
      RECT  67215.0 103335.0 67920.0 101990.0 ;
      RECT  67215.0 103335.0 67920.0 104680.0 ;
      RECT  67215.0 106025.0 67920.0 104680.0 ;
      RECT  67215.0 106025.0 67920.0 107370.0 ;
      RECT  67215.0 108715.0 67920.0 107370.0 ;
      RECT  67215.0 108715.0 67920.0 110060.0 ;
      RECT  67215.0 111405.0 67920.0 110060.0 ;
      RECT  67215.0 111405.0 67920.0 112750.0 ;
      RECT  67215.0 114095.0 67920.0 112750.0 ;
      RECT  67920.0 28015.0 68625.0 29360.0 ;
      RECT  67920.0 30705.0 68625.0 29360.0 ;
      RECT  67920.0 30705.0 68625.0 32050.0 ;
      RECT  67920.0 33395.0 68625.0 32050.0 ;
      RECT  67920.0 33395.0 68625.0 34740.0 ;
      RECT  67920.0 36085.0 68625.0 34740.0 ;
      RECT  67920.0 36085.0 68625.0 37430.0 ;
      RECT  67920.0 38775.0 68625.0 37430.0 ;
      RECT  67920.0 38775.0 68625.0 40120.0 ;
      RECT  67920.0 41465.0 68625.0 40120.0 ;
      RECT  67920.0 41465.0 68625.0 42810.0 ;
      RECT  67920.0 44155.0 68625.0 42810.0 ;
      RECT  67920.0 44155.0 68625.0 45500.0 ;
      RECT  67920.0 46845.0 68625.0 45500.0 ;
      RECT  67920.0 46845.0 68625.0 48190.0 ;
      RECT  67920.0 49535.0 68625.0 48190.0 ;
      RECT  67920.0 49535.0 68625.0 50880.0 ;
      RECT  67920.0 52225.0 68625.0 50880.0 ;
      RECT  67920.0 52225.0 68625.0 53570.0 ;
      RECT  67920.0 54915.0 68625.0 53570.0 ;
      RECT  67920.0 54915.0 68625.0 56260.0 ;
      RECT  67920.0 57605.0 68625.0 56260.0 ;
      RECT  67920.0 57605.0 68625.0 58950.0 ;
      RECT  67920.0 60295.0 68625.0 58950.0 ;
      RECT  67920.0 60295.0 68625.0 61640.0 ;
      RECT  67920.0 62985.0 68625.0 61640.0 ;
      RECT  67920.0 62985.0 68625.0 64330.0 ;
      RECT  67920.0 65675.0 68625.0 64330.0 ;
      RECT  67920.0 65675.0 68625.0 67020.0 ;
      RECT  67920.0 68365.0 68625.0 67020.0 ;
      RECT  67920.0 68365.0 68625.0 69710.0 ;
      RECT  67920.0 71055.0 68625.0 69710.0 ;
      RECT  67920.0 71055.0 68625.0 72400.0 ;
      RECT  67920.0 73745.0 68625.0 72400.0 ;
      RECT  67920.0 73745.0 68625.0 75090.0 ;
      RECT  67920.0 76435.0 68625.0 75090.0 ;
      RECT  67920.0 76435.0 68625.0 77780.0 ;
      RECT  67920.0 79125.0 68625.0 77780.0 ;
      RECT  67920.0 79125.0 68625.0 80470.0 ;
      RECT  67920.0 81815.0 68625.0 80470.0 ;
      RECT  67920.0 81815.0 68625.0 83160.0 ;
      RECT  67920.0 84505.0 68625.0 83160.0 ;
      RECT  67920.0 84505.0 68625.0 85850.0 ;
      RECT  67920.0 87195.0 68625.0 85850.0 ;
      RECT  67920.0 87195.0 68625.0 88540.0 ;
      RECT  67920.0 89885.0 68625.0 88540.0 ;
      RECT  67920.0 89885.0 68625.0 91230.0 ;
      RECT  67920.0 92575.0 68625.0 91230.0 ;
      RECT  67920.0 92575.0 68625.0 93920.0 ;
      RECT  67920.0 95265.0 68625.0 93920.0 ;
      RECT  67920.0 95265.0 68625.0 96610.0 ;
      RECT  67920.0 97955.0 68625.0 96610.0 ;
      RECT  67920.0 97955.0 68625.0 99300.0 ;
      RECT  67920.0 100645.0 68625.0 99300.0 ;
      RECT  67920.0 100645.0 68625.0 101990.0 ;
      RECT  67920.0 103335.0 68625.0 101990.0 ;
      RECT  67920.0 103335.0 68625.0 104680.0 ;
      RECT  67920.0 106025.0 68625.0 104680.0 ;
      RECT  67920.0 106025.0 68625.0 107370.0 ;
      RECT  67920.0 108715.0 68625.0 107370.0 ;
      RECT  67920.0 108715.0 68625.0 110060.0 ;
      RECT  67920.0 111405.0 68625.0 110060.0 ;
      RECT  67920.0 111405.0 68625.0 112750.0 ;
      RECT  67920.0 114095.0 68625.0 112750.0 ;
      RECT  68625.0 28015.0 69330.0 29360.0 ;
      RECT  68625.0 30705.0 69330.0 29360.0 ;
      RECT  68625.0 30705.0 69330.0 32050.0 ;
      RECT  68625.0 33395.0 69330.0 32050.0 ;
      RECT  68625.0 33395.0 69330.0 34740.0 ;
      RECT  68625.0 36085.0 69330.0 34740.0 ;
      RECT  68625.0 36085.0 69330.0 37430.0 ;
      RECT  68625.0 38775.0 69330.0 37430.0 ;
      RECT  68625.0 38775.0 69330.0 40120.0 ;
      RECT  68625.0 41465.0 69330.0 40120.0 ;
      RECT  68625.0 41465.0 69330.0 42810.0 ;
      RECT  68625.0 44155.0 69330.0 42810.0 ;
      RECT  68625.0 44155.0 69330.0 45500.0 ;
      RECT  68625.0 46845.0 69330.0 45500.0 ;
      RECT  68625.0 46845.0 69330.0 48190.0 ;
      RECT  68625.0 49535.0 69330.0 48190.0 ;
      RECT  68625.0 49535.0 69330.0 50880.0 ;
      RECT  68625.0 52225.0 69330.0 50880.0 ;
      RECT  68625.0 52225.0 69330.0 53570.0 ;
      RECT  68625.0 54915.0 69330.0 53570.0 ;
      RECT  68625.0 54915.0 69330.0 56260.0 ;
      RECT  68625.0 57605.0 69330.0 56260.0 ;
      RECT  68625.0 57605.0 69330.0 58950.0 ;
      RECT  68625.0 60295.0 69330.0 58950.0 ;
      RECT  68625.0 60295.0 69330.0 61640.0 ;
      RECT  68625.0 62985.0 69330.0 61640.0 ;
      RECT  68625.0 62985.0 69330.0 64330.0 ;
      RECT  68625.0 65675.0 69330.0 64330.0 ;
      RECT  68625.0 65675.0 69330.0 67020.0 ;
      RECT  68625.0 68365.0 69330.0 67020.0 ;
      RECT  68625.0 68365.0 69330.0 69710.0 ;
      RECT  68625.0 71055.0 69330.0 69710.0 ;
      RECT  68625.0 71055.0 69330.0 72400.0 ;
      RECT  68625.0 73745.0 69330.0 72400.0 ;
      RECT  68625.0 73745.0 69330.0 75090.0 ;
      RECT  68625.0 76435.0 69330.0 75090.0 ;
      RECT  68625.0 76435.0 69330.0 77780.0 ;
      RECT  68625.0 79125.0 69330.0 77780.0 ;
      RECT  68625.0 79125.0 69330.0 80470.0 ;
      RECT  68625.0 81815.0 69330.0 80470.0 ;
      RECT  68625.0 81815.0 69330.0 83160.0 ;
      RECT  68625.0 84505.0 69330.0 83160.0 ;
      RECT  68625.0 84505.0 69330.0 85850.0 ;
      RECT  68625.0 87195.0 69330.0 85850.0 ;
      RECT  68625.0 87195.0 69330.0 88540.0 ;
      RECT  68625.0 89885.0 69330.0 88540.0 ;
      RECT  68625.0 89885.0 69330.0 91230.0 ;
      RECT  68625.0 92575.0 69330.0 91230.0 ;
      RECT  68625.0 92575.0 69330.0 93920.0 ;
      RECT  68625.0 95265.0 69330.0 93920.0 ;
      RECT  68625.0 95265.0 69330.0 96610.0 ;
      RECT  68625.0 97955.0 69330.0 96610.0 ;
      RECT  68625.0 97955.0 69330.0 99300.0 ;
      RECT  68625.0 100645.0 69330.0 99300.0 ;
      RECT  68625.0 100645.0 69330.0 101990.0 ;
      RECT  68625.0 103335.0 69330.0 101990.0 ;
      RECT  68625.0 103335.0 69330.0 104680.0 ;
      RECT  68625.0 106025.0 69330.0 104680.0 ;
      RECT  68625.0 106025.0 69330.0 107370.0 ;
      RECT  68625.0 108715.0 69330.0 107370.0 ;
      RECT  68625.0 108715.0 69330.0 110060.0 ;
      RECT  68625.0 111405.0 69330.0 110060.0 ;
      RECT  68625.0 111405.0 69330.0 112750.0 ;
      RECT  68625.0 114095.0 69330.0 112750.0 ;
      RECT  69330.0 28015.0 70035.0 29360.0 ;
      RECT  69330.0 30705.0 70035.0 29360.0 ;
      RECT  69330.0 30705.0 70035.0 32050.0 ;
      RECT  69330.0 33395.0 70035.0 32050.0 ;
      RECT  69330.0 33395.0 70035.0 34740.0 ;
      RECT  69330.0 36085.0 70035.0 34740.0 ;
      RECT  69330.0 36085.0 70035.0 37430.0 ;
      RECT  69330.0 38775.0 70035.0 37430.0 ;
      RECT  69330.0 38775.0 70035.0 40120.0 ;
      RECT  69330.0 41465.0 70035.0 40120.0 ;
      RECT  69330.0 41465.0 70035.0 42810.0 ;
      RECT  69330.0 44155.0 70035.0 42810.0 ;
      RECT  69330.0 44155.0 70035.0 45500.0 ;
      RECT  69330.0 46845.0 70035.0 45500.0 ;
      RECT  69330.0 46845.0 70035.0 48190.0 ;
      RECT  69330.0 49535.0 70035.0 48190.0 ;
      RECT  69330.0 49535.0 70035.0 50880.0 ;
      RECT  69330.0 52225.0 70035.0 50880.0 ;
      RECT  69330.0 52225.0 70035.0 53570.0 ;
      RECT  69330.0 54915.0 70035.0 53570.0 ;
      RECT  69330.0 54915.0 70035.0 56260.0 ;
      RECT  69330.0 57605.0 70035.0 56260.0 ;
      RECT  69330.0 57605.0 70035.0 58950.0 ;
      RECT  69330.0 60295.0 70035.0 58950.0 ;
      RECT  69330.0 60295.0 70035.0 61640.0 ;
      RECT  69330.0 62985.0 70035.0 61640.0 ;
      RECT  69330.0 62985.0 70035.0 64330.0 ;
      RECT  69330.0 65675.0 70035.0 64330.0 ;
      RECT  69330.0 65675.0 70035.0 67020.0 ;
      RECT  69330.0 68365.0 70035.0 67020.0 ;
      RECT  69330.0 68365.0 70035.0 69710.0 ;
      RECT  69330.0 71055.0 70035.0 69710.0 ;
      RECT  69330.0 71055.0 70035.0 72400.0 ;
      RECT  69330.0 73745.0 70035.0 72400.0 ;
      RECT  69330.0 73745.0 70035.0 75090.0 ;
      RECT  69330.0 76435.0 70035.0 75090.0 ;
      RECT  69330.0 76435.0 70035.0 77780.0 ;
      RECT  69330.0 79125.0 70035.0 77780.0 ;
      RECT  69330.0 79125.0 70035.0 80470.0 ;
      RECT  69330.0 81815.0 70035.0 80470.0 ;
      RECT  69330.0 81815.0 70035.0 83160.0 ;
      RECT  69330.0 84505.0 70035.0 83160.0 ;
      RECT  69330.0 84505.0 70035.0 85850.0 ;
      RECT  69330.0 87195.0 70035.0 85850.0 ;
      RECT  69330.0 87195.0 70035.0 88540.0 ;
      RECT  69330.0 89885.0 70035.0 88540.0 ;
      RECT  69330.0 89885.0 70035.0 91230.0 ;
      RECT  69330.0 92575.0 70035.0 91230.0 ;
      RECT  69330.0 92575.0 70035.0 93920.0 ;
      RECT  69330.0 95265.0 70035.0 93920.0 ;
      RECT  69330.0 95265.0 70035.0 96610.0 ;
      RECT  69330.0 97955.0 70035.0 96610.0 ;
      RECT  69330.0 97955.0 70035.0 99300.0 ;
      RECT  69330.0 100645.0 70035.0 99300.0 ;
      RECT  69330.0 100645.0 70035.0 101990.0 ;
      RECT  69330.0 103335.0 70035.0 101990.0 ;
      RECT  69330.0 103335.0 70035.0 104680.0 ;
      RECT  69330.0 106025.0 70035.0 104680.0 ;
      RECT  69330.0 106025.0 70035.0 107370.0 ;
      RECT  69330.0 108715.0 70035.0 107370.0 ;
      RECT  69330.0 108715.0 70035.0 110060.0 ;
      RECT  69330.0 111405.0 70035.0 110060.0 ;
      RECT  69330.0 111405.0 70035.0 112750.0 ;
      RECT  69330.0 114095.0 70035.0 112750.0 ;
      RECT  70035.0 28015.0 70740.0 29360.0 ;
      RECT  70035.0 30705.0 70740.0 29360.0 ;
      RECT  70035.0 30705.0 70740.0 32050.0 ;
      RECT  70035.0 33395.0 70740.0 32050.0 ;
      RECT  70035.0 33395.0 70740.0 34740.0 ;
      RECT  70035.0 36085.0 70740.0 34740.0 ;
      RECT  70035.0 36085.0 70740.0 37430.0 ;
      RECT  70035.0 38775.0 70740.0 37430.0 ;
      RECT  70035.0 38775.0 70740.0 40120.0 ;
      RECT  70035.0 41465.0 70740.0 40120.0 ;
      RECT  70035.0 41465.0 70740.0 42810.0 ;
      RECT  70035.0 44155.0 70740.0 42810.0 ;
      RECT  70035.0 44155.0 70740.0 45500.0 ;
      RECT  70035.0 46845.0 70740.0 45500.0 ;
      RECT  70035.0 46845.0 70740.0 48190.0 ;
      RECT  70035.0 49535.0 70740.0 48190.0 ;
      RECT  70035.0 49535.0 70740.0 50880.0 ;
      RECT  70035.0 52225.0 70740.0 50880.0 ;
      RECT  70035.0 52225.0 70740.0 53570.0 ;
      RECT  70035.0 54915.0 70740.0 53570.0 ;
      RECT  70035.0 54915.0 70740.0 56260.0 ;
      RECT  70035.0 57605.0 70740.0 56260.0 ;
      RECT  70035.0 57605.0 70740.0 58950.0 ;
      RECT  70035.0 60295.0 70740.0 58950.0 ;
      RECT  70035.0 60295.0 70740.0 61640.0 ;
      RECT  70035.0 62985.0 70740.0 61640.0 ;
      RECT  70035.0 62985.0 70740.0 64330.0 ;
      RECT  70035.0 65675.0 70740.0 64330.0 ;
      RECT  70035.0 65675.0 70740.0 67020.0 ;
      RECT  70035.0 68365.0 70740.0 67020.0 ;
      RECT  70035.0 68365.0 70740.0 69710.0 ;
      RECT  70035.0 71055.0 70740.0 69710.0 ;
      RECT  70035.0 71055.0 70740.0 72400.0 ;
      RECT  70035.0 73745.0 70740.0 72400.0 ;
      RECT  70035.0 73745.0 70740.0 75090.0 ;
      RECT  70035.0 76435.0 70740.0 75090.0 ;
      RECT  70035.0 76435.0 70740.0 77780.0 ;
      RECT  70035.0 79125.0 70740.0 77780.0 ;
      RECT  70035.0 79125.0 70740.0 80470.0 ;
      RECT  70035.0 81815.0 70740.0 80470.0 ;
      RECT  70035.0 81815.0 70740.0 83160.0 ;
      RECT  70035.0 84505.0 70740.0 83160.0 ;
      RECT  70035.0 84505.0 70740.0 85850.0 ;
      RECT  70035.0 87195.0 70740.0 85850.0 ;
      RECT  70035.0 87195.0 70740.0 88540.0 ;
      RECT  70035.0 89885.0 70740.0 88540.0 ;
      RECT  70035.0 89885.0 70740.0 91230.0 ;
      RECT  70035.0 92575.0 70740.0 91230.0 ;
      RECT  70035.0 92575.0 70740.0 93920.0 ;
      RECT  70035.0 95265.0 70740.0 93920.0 ;
      RECT  70035.0 95265.0 70740.0 96610.0 ;
      RECT  70035.0 97955.0 70740.0 96610.0 ;
      RECT  70035.0 97955.0 70740.0 99300.0 ;
      RECT  70035.0 100645.0 70740.0 99300.0 ;
      RECT  70035.0 100645.0 70740.0 101990.0 ;
      RECT  70035.0 103335.0 70740.0 101990.0 ;
      RECT  70035.0 103335.0 70740.0 104680.0 ;
      RECT  70035.0 106025.0 70740.0 104680.0 ;
      RECT  70035.0 106025.0 70740.0 107370.0 ;
      RECT  70035.0 108715.0 70740.0 107370.0 ;
      RECT  70035.0 108715.0 70740.0 110060.0 ;
      RECT  70035.0 111405.0 70740.0 110060.0 ;
      RECT  70035.0 111405.0 70740.0 112750.0 ;
      RECT  70035.0 114095.0 70740.0 112750.0 ;
      RECT  70740.0 28015.0 71445.0 29360.0 ;
      RECT  70740.0 30705.0 71445.0 29360.0 ;
      RECT  70740.0 30705.0 71445.0 32050.0 ;
      RECT  70740.0 33395.0 71445.0 32050.0 ;
      RECT  70740.0 33395.0 71445.0 34740.0 ;
      RECT  70740.0 36085.0 71445.0 34740.0 ;
      RECT  70740.0 36085.0 71445.0 37430.0 ;
      RECT  70740.0 38775.0 71445.0 37430.0 ;
      RECT  70740.0 38775.0 71445.0 40120.0 ;
      RECT  70740.0 41465.0 71445.0 40120.0 ;
      RECT  70740.0 41465.0 71445.0 42810.0 ;
      RECT  70740.0 44155.0 71445.0 42810.0 ;
      RECT  70740.0 44155.0 71445.0 45500.0 ;
      RECT  70740.0 46845.0 71445.0 45500.0 ;
      RECT  70740.0 46845.0 71445.0 48190.0 ;
      RECT  70740.0 49535.0 71445.0 48190.0 ;
      RECT  70740.0 49535.0 71445.0 50880.0 ;
      RECT  70740.0 52225.0 71445.0 50880.0 ;
      RECT  70740.0 52225.0 71445.0 53570.0 ;
      RECT  70740.0 54915.0 71445.0 53570.0 ;
      RECT  70740.0 54915.0 71445.0 56260.0 ;
      RECT  70740.0 57605.0 71445.0 56260.0 ;
      RECT  70740.0 57605.0 71445.0 58950.0 ;
      RECT  70740.0 60295.0 71445.0 58950.0 ;
      RECT  70740.0 60295.0 71445.0 61640.0 ;
      RECT  70740.0 62985.0 71445.0 61640.0 ;
      RECT  70740.0 62985.0 71445.0 64330.0 ;
      RECT  70740.0 65675.0 71445.0 64330.0 ;
      RECT  70740.0 65675.0 71445.0 67020.0 ;
      RECT  70740.0 68365.0 71445.0 67020.0 ;
      RECT  70740.0 68365.0 71445.0 69710.0 ;
      RECT  70740.0 71055.0 71445.0 69710.0 ;
      RECT  70740.0 71055.0 71445.0 72400.0 ;
      RECT  70740.0 73745.0 71445.0 72400.0 ;
      RECT  70740.0 73745.0 71445.0 75090.0 ;
      RECT  70740.0 76435.0 71445.0 75090.0 ;
      RECT  70740.0 76435.0 71445.0 77780.0 ;
      RECT  70740.0 79125.0 71445.0 77780.0 ;
      RECT  70740.0 79125.0 71445.0 80470.0 ;
      RECT  70740.0 81815.0 71445.0 80470.0 ;
      RECT  70740.0 81815.0 71445.0 83160.0 ;
      RECT  70740.0 84505.0 71445.0 83160.0 ;
      RECT  70740.0 84505.0 71445.0 85850.0 ;
      RECT  70740.0 87195.0 71445.0 85850.0 ;
      RECT  70740.0 87195.0 71445.0 88540.0 ;
      RECT  70740.0 89885.0 71445.0 88540.0 ;
      RECT  70740.0 89885.0 71445.0 91230.0 ;
      RECT  70740.0 92575.0 71445.0 91230.0 ;
      RECT  70740.0 92575.0 71445.0 93920.0 ;
      RECT  70740.0 95265.0 71445.0 93920.0 ;
      RECT  70740.0 95265.0 71445.0 96610.0 ;
      RECT  70740.0 97955.0 71445.0 96610.0 ;
      RECT  70740.0 97955.0 71445.0 99300.0 ;
      RECT  70740.0 100645.0 71445.0 99300.0 ;
      RECT  70740.0 100645.0 71445.0 101990.0 ;
      RECT  70740.0 103335.0 71445.0 101990.0 ;
      RECT  70740.0 103335.0 71445.0 104680.0 ;
      RECT  70740.0 106025.0 71445.0 104680.0 ;
      RECT  70740.0 106025.0 71445.0 107370.0 ;
      RECT  70740.0 108715.0 71445.0 107370.0 ;
      RECT  70740.0 108715.0 71445.0 110060.0 ;
      RECT  70740.0 111405.0 71445.0 110060.0 ;
      RECT  70740.0 111405.0 71445.0 112750.0 ;
      RECT  70740.0 114095.0 71445.0 112750.0 ;
      RECT  71445.0 28015.0 72150.0 29360.0 ;
      RECT  71445.0 30705.0 72150.0 29360.0 ;
      RECT  71445.0 30705.0 72150.0 32050.0 ;
      RECT  71445.0 33395.0 72150.0 32050.0 ;
      RECT  71445.0 33395.0 72150.0 34740.0 ;
      RECT  71445.0 36085.0 72150.0 34740.0 ;
      RECT  71445.0 36085.0 72150.0 37430.0 ;
      RECT  71445.0 38775.0 72150.0 37430.0 ;
      RECT  71445.0 38775.0 72150.0 40120.0 ;
      RECT  71445.0 41465.0 72150.0 40120.0 ;
      RECT  71445.0 41465.0 72150.0 42810.0 ;
      RECT  71445.0 44155.0 72150.0 42810.0 ;
      RECT  71445.0 44155.0 72150.0 45500.0 ;
      RECT  71445.0 46845.0 72150.0 45500.0 ;
      RECT  71445.0 46845.0 72150.0 48190.0 ;
      RECT  71445.0 49535.0 72150.0 48190.0 ;
      RECT  71445.0 49535.0 72150.0 50880.0 ;
      RECT  71445.0 52225.0 72150.0 50880.0 ;
      RECT  71445.0 52225.0 72150.0 53570.0 ;
      RECT  71445.0 54915.0 72150.0 53570.0 ;
      RECT  71445.0 54915.0 72150.0 56260.0 ;
      RECT  71445.0 57605.0 72150.0 56260.0 ;
      RECT  71445.0 57605.0 72150.0 58950.0 ;
      RECT  71445.0 60295.0 72150.0 58950.0 ;
      RECT  71445.0 60295.0 72150.0 61640.0 ;
      RECT  71445.0 62985.0 72150.0 61640.0 ;
      RECT  71445.0 62985.0 72150.0 64330.0 ;
      RECT  71445.0 65675.0 72150.0 64330.0 ;
      RECT  71445.0 65675.0 72150.0 67020.0 ;
      RECT  71445.0 68365.0 72150.0 67020.0 ;
      RECT  71445.0 68365.0 72150.0 69710.0 ;
      RECT  71445.0 71055.0 72150.0 69710.0 ;
      RECT  71445.0 71055.0 72150.0 72400.0 ;
      RECT  71445.0 73745.0 72150.0 72400.0 ;
      RECT  71445.0 73745.0 72150.0 75090.0 ;
      RECT  71445.0 76435.0 72150.0 75090.0 ;
      RECT  71445.0 76435.0 72150.0 77780.0 ;
      RECT  71445.0 79125.0 72150.0 77780.0 ;
      RECT  71445.0 79125.0 72150.0 80470.0 ;
      RECT  71445.0 81815.0 72150.0 80470.0 ;
      RECT  71445.0 81815.0 72150.0 83160.0 ;
      RECT  71445.0 84505.0 72150.0 83160.0 ;
      RECT  71445.0 84505.0 72150.0 85850.0 ;
      RECT  71445.0 87195.0 72150.0 85850.0 ;
      RECT  71445.0 87195.0 72150.0 88540.0 ;
      RECT  71445.0 89885.0 72150.0 88540.0 ;
      RECT  71445.0 89885.0 72150.0 91230.0 ;
      RECT  71445.0 92575.0 72150.0 91230.0 ;
      RECT  71445.0 92575.0 72150.0 93920.0 ;
      RECT  71445.0 95265.0 72150.0 93920.0 ;
      RECT  71445.0 95265.0 72150.0 96610.0 ;
      RECT  71445.0 97955.0 72150.0 96610.0 ;
      RECT  71445.0 97955.0 72150.0 99300.0 ;
      RECT  71445.0 100645.0 72150.0 99300.0 ;
      RECT  71445.0 100645.0 72150.0 101990.0 ;
      RECT  71445.0 103335.0 72150.0 101990.0 ;
      RECT  71445.0 103335.0 72150.0 104680.0 ;
      RECT  71445.0 106025.0 72150.0 104680.0 ;
      RECT  71445.0 106025.0 72150.0 107370.0 ;
      RECT  71445.0 108715.0 72150.0 107370.0 ;
      RECT  71445.0 108715.0 72150.0 110060.0 ;
      RECT  71445.0 111405.0 72150.0 110060.0 ;
      RECT  71445.0 111405.0 72150.0 112750.0 ;
      RECT  71445.0 114095.0 72150.0 112750.0 ;
      RECT  72150.0 28015.0 72855.0 29360.0 ;
      RECT  72150.0 30705.0 72855.0 29360.0 ;
      RECT  72150.0 30705.0 72855.0 32050.0 ;
      RECT  72150.0 33395.0 72855.0 32050.0 ;
      RECT  72150.0 33395.0 72855.0 34740.0 ;
      RECT  72150.0 36085.0 72855.0 34740.0 ;
      RECT  72150.0 36085.0 72855.0 37430.0 ;
      RECT  72150.0 38775.0 72855.0 37430.0 ;
      RECT  72150.0 38775.0 72855.0 40120.0 ;
      RECT  72150.0 41465.0 72855.0 40120.0 ;
      RECT  72150.0 41465.0 72855.0 42810.0 ;
      RECT  72150.0 44155.0 72855.0 42810.0 ;
      RECT  72150.0 44155.0 72855.0 45500.0 ;
      RECT  72150.0 46845.0 72855.0 45500.0 ;
      RECT  72150.0 46845.0 72855.0 48190.0 ;
      RECT  72150.0 49535.0 72855.0 48190.0 ;
      RECT  72150.0 49535.0 72855.0 50880.0 ;
      RECT  72150.0 52225.0 72855.0 50880.0 ;
      RECT  72150.0 52225.0 72855.0 53570.0 ;
      RECT  72150.0 54915.0 72855.0 53570.0 ;
      RECT  72150.0 54915.0 72855.0 56260.0 ;
      RECT  72150.0 57605.0 72855.0 56260.0 ;
      RECT  72150.0 57605.0 72855.0 58950.0 ;
      RECT  72150.0 60295.0 72855.0 58950.0 ;
      RECT  72150.0 60295.0 72855.0 61640.0 ;
      RECT  72150.0 62985.0 72855.0 61640.0 ;
      RECT  72150.0 62985.0 72855.0 64330.0 ;
      RECT  72150.0 65675.0 72855.0 64330.0 ;
      RECT  72150.0 65675.0 72855.0 67020.0 ;
      RECT  72150.0 68365.0 72855.0 67020.0 ;
      RECT  72150.0 68365.0 72855.0 69710.0 ;
      RECT  72150.0 71055.0 72855.0 69710.0 ;
      RECT  72150.0 71055.0 72855.0 72400.0 ;
      RECT  72150.0 73745.0 72855.0 72400.0 ;
      RECT  72150.0 73745.0 72855.0 75090.0 ;
      RECT  72150.0 76435.0 72855.0 75090.0 ;
      RECT  72150.0 76435.0 72855.0 77780.0 ;
      RECT  72150.0 79125.0 72855.0 77780.0 ;
      RECT  72150.0 79125.0 72855.0 80470.0 ;
      RECT  72150.0 81815.0 72855.0 80470.0 ;
      RECT  72150.0 81815.0 72855.0 83160.0 ;
      RECT  72150.0 84505.0 72855.0 83160.0 ;
      RECT  72150.0 84505.0 72855.0 85850.0 ;
      RECT  72150.0 87195.0 72855.0 85850.0 ;
      RECT  72150.0 87195.0 72855.0 88540.0 ;
      RECT  72150.0 89885.0 72855.0 88540.0 ;
      RECT  72150.0 89885.0 72855.0 91230.0 ;
      RECT  72150.0 92575.0 72855.0 91230.0 ;
      RECT  72150.0 92575.0 72855.0 93920.0 ;
      RECT  72150.0 95265.0 72855.0 93920.0 ;
      RECT  72150.0 95265.0 72855.0 96610.0 ;
      RECT  72150.0 97955.0 72855.0 96610.0 ;
      RECT  72150.0 97955.0 72855.0 99300.0 ;
      RECT  72150.0 100645.0 72855.0 99300.0 ;
      RECT  72150.0 100645.0 72855.0 101990.0 ;
      RECT  72150.0 103335.0 72855.0 101990.0 ;
      RECT  72150.0 103335.0 72855.0 104680.0 ;
      RECT  72150.0 106025.0 72855.0 104680.0 ;
      RECT  72150.0 106025.0 72855.0 107370.0 ;
      RECT  72150.0 108715.0 72855.0 107370.0 ;
      RECT  72150.0 108715.0 72855.0 110060.0 ;
      RECT  72150.0 111405.0 72855.0 110060.0 ;
      RECT  72150.0 111405.0 72855.0 112750.0 ;
      RECT  72150.0 114095.0 72855.0 112750.0 ;
      RECT  72855.0 28015.0 73560.0 29360.0 ;
      RECT  72855.0 30705.0 73560.0 29360.0 ;
      RECT  72855.0 30705.0 73560.0 32050.0 ;
      RECT  72855.0 33395.0 73560.0 32050.0 ;
      RECT  72855.0 33395.0 73560.0 34740.0 ;
      RECT  72855.0 36085.0 73560.0 34740.0 ;
      RECT  72855.0 36085.0 73560.0 37430.0 ;
      RECT  72855.0 38775.0 73560.0 37430.0 ;
      RECT  72855.0 38775.0 73560.0 40120.0 ;
      RECT  72855.0 41465.0 73560.0 40120.0 ;
      RECT  72855.0 41465.0 73560.0 42810.0 ;
      RECT  72855.0 44155.0 73560.0 42810.0 ;
      RECT  72855.0 44155.0 73560.0 45500.0 ;
      RECT  72855.0 46845.0 73560.0 45500.0 ;
      RECT  72855.0 46845.0 73560.0 48190.0 ;
      RECT  72855.0 49535.0 73560.0 48190.0 ;
      RECT  72855.0 49535.0 73560.0 50880.0 ;
      RECT  72855.0 52225.0 73560.0 50880.0 ;
      RECT  72855.0 52225.0 73560.0 53570.0 ;
      RECT  72855.0 54915.0 73560.0 53570.0 ;
      RECT  72855.0 54915.0 73560.0 56260.0 ;
      RECT  72855.0 57605.0 73560.0 56260.0 ;
      RECT  72855.0 57605.0 73560.0 58950.0 ;
      RECT  72855.0 60295.0 73560.0 58950.0 ;
      RECT  72855.0 60295.0 73560.0 61640.0 ;
      RECT  72855.0 62985.0 73560.0 61640.0 ;
      RECT  72855.0 62985.0 73560.0 64330.0 ;
      RECT  72855.0 65675.0 73560.0 64330.0 ;
      RECT  72855.0 65675.0 73560.0 67020.0 ;
      RECT  72855.0 68365.0 73560.0 67020.0 ;
      RECT  72855.0 68365.0 73560.0 69710.0 ;
      RECT  72855.0 71055.0 73560.0 69710.0 ;
      RECT  72855.0 71055.0 73560.0 72400.0 ;
      RECT  72855.0 73745.0 73560.0 72400.0 ;
      RECT  72855.0 73745.0 73560.0 75090.0 ;
      RECT  72855.0 76435.0 73560.0 75090.0 ;
      RECT  72855.0 76435.0 73560.0 77780.0 ;
      RECT  72855.0 79125.0 73560.0 77780.0 ;
      RECT  72855.0 79125.0 73560.0 80470.0 ;
      RECT  72855.0 81815.0 73560.0 80470.0 ;
      RECT  72855.0 81815.0 73560.0 83160.0 ;
      RECT  72855.0 84505.0 73560.0 83160.0 ;
      RECT  72855.0 84505.0 73560.0 85850.0 ;
      RECT  72855.0 87195.0 73560.0 85850.0 ;
      RECT  72855.0 87195.0 73560.0 88540.0 ;
      RECT  72855.0 89885.0 73560.0 88540.0 ;
      RECT  72855.0 89885.0 73560.0 91230.0 ;
      RECT  72855.0 92575.0 73560.0 91230.0 ;
      RECT  72855.0 92575.0 73560.0 93920.0 ;
      RECT  72855.0 95265.0 73560.0 93920.0 ;
      RECT  72855.0 95265.0 73560.0 96610.0 ;
      RECT  72855.0 97955.0 73560.0 96610.0 ;
      RECT  72855.0 97955.0 73560.0 99300.0 ;
      RECT  72855.0 100645.0 73560.0 99300.0 ;
      RECT  72855.0 100645.0 73560.0 101990.0 ;
      RECT  72855.0 103335.0 73560.0 101990.0 ;
      RECT  72855.0 103335.0 73560.0 104680.0 ;
      RECT  72855.0 106025.0 73560.0 104680.0 ;
      RECT  72855.0 106025.0 73560.0 107370.0 ;
      RECT  72855.0 108715.0 73560.0 107370.0 ;
      RECT  72855.0 108715.0 73560.0 110060.0 ;
      RECT  72855.0 111405.0 73560.0 110060.0 ;
      RECT  72855.0 111405.0 73560.0 112750.0 ;
      RECT  72855.0 114095.0 73560.0 112750.0 ;
      RECT  73560.0 28015.0 74265.0 29360.0 ;
      RECT  73560.0 30705.0 74265.0 29360.0 ;
      RECT  73560.0 30705.0 74265.0 32050.0 ;
      RECT  73560.0 33395.0 74265.0 32050.0 ;
      RECT  73560.0 33395.0 74265.0 34740.0 ;
      RECT  73560.0 36085.0 74265.0 34740.0 ;
      RECT  73560.0 36085.0 74265.0 37430.0 ;
      RECT  73560.0 38775.0 74265.0 37430.0 ;
      RECT  73560.0 38775.0 74265.0 40120.0 ;
      RECT  73560.0 41465.0 74265.0 40120.0 ;
      RECT  73560.0 41465.0 74265.0 42810.0 ;
      RECT  73560.0 44155.0 74265.0 42810.0 ;
      RECT  73560.0 44155.0 74265.0 45500.0 ;
      RECT  73560.0 46845.0 74265.0 45500.0 ;
      RECT  73560.0 46845.0 74265.0 48190.0 ;
      RECT  73560.0 49535.0 74265.0 48190.0 ;
      RECT  73560.0 49535.0 74265.0 50880.0 ;
      RECT  73560.0 52225.0 74265.0 50880.0 ;
      RECT  73560.0 52225.0 74265.0 53570.0 ;
      RECT  73560.0 54915.0 74265.0 53570.0 ;
      RECT  73560.0 54915.0 74265.0 56260.0 ;
      RECT  73560.0 57605.0 74265.0 56260.0 ;
      RECT  73560.0 57605.0 74265.0 58950.0 ;
      RECT  73560.0 60295.0 74265.0 58950.0 ;
      RECT  73560.0 60295.0 74265.0 61640.0 ;
      RECT  73560.0 62985.0 74265.0 61640.0 ;
      RECT  73560.0 62985.0 74265.0 64330.0 ;
      RECT  73560.0 65675.0 74265.0 64330.0 ;
      RECT  73560.0 65675.0 74265.0 67020.0 ;
      RECT  73560.0 68365.0 74265.0 67020.0 ;
      RECT  73560.0 68365.0 74265.0 69710.0 ;
      RECT  73560.0 71055.0 74265.0 69710.0 ;
      RECT  73560.0 71055.0 74265.0 72400.0 ;
      RECT  73560.0 73745.0 74265.0 72400.0 ;
      RECT  73560.0 73745.0 74265.0 75090.0 ;
      RECT  73560.0 76435.0 74265.0 75090.0 ;
      RECT  73560.0 76435.0 74265.0 77780.0 ;
      RECT  73560.0 79125.0 74265.0 77780.0 ;
      RECT  73560.0 79125.0 74265.0 80470.0 ;
      RECT  73560.0 81815.0 74265.0 80470.0 ;
      RECT  73560.0 81815.0 74265.0 83160.0 ;
      RECT  73560.0 84505.0 74265.0 83160.0 ;
      RECT  73560.0 84505.0 74265.0 85850.0 ;
      RECT  73560.0 87195.0 74265.0 85850.0 ;
      RECT  73560.0 87195.0 74265.0 88540.0 ;
      RECT  73560.0 89885.0 74265.0 88540.0 ;
      RECT  73560.0 89885.0 74265.0 91230.0 ;
      RECT  73560.0 92575.0 74265.0 91230.0 ;
      RECT  73560.0 92575.0 74265.0 93920.0 ;
      RECT  73560.0 95265.0 74265.0 93920.0 ;
      RECT  73560.0 95265.0 74265.0 96610.0 ;
      RECT  73560.0 97955.0 74265.0 96610.0 ;
      RECT  73560.0 97955.0 74265.0 99300.0 ;
      RECT  73560.0 100645.0 74265.0 99300.0 ;
      RECT  73560.0 100645.0 74265.0 101990.0 ;
      RECT  73560.0 103335.0 74265.0 101990.0 ;
      RECT  73560.0 103335.0 74265.0 104680.0 ;
      RECT  73560.0 106025.0 74265.0 104680.0 ;
      RECT  73560.0 106025.0 74265.0 107370.0 ;
      RECT  73560.0 108715.0 74265.0 107370.0 ;
      RECT  73560.0 108715.0 74265.0 110060.0 ;
      RECT  73560.0 111405.0 74265.0 110060.0 ;
      RECT  73560.0 111405.0 74265.0 112750.0 ;
      RECT  73560.0 114095.0 74265.0 112750.0 ;
      RECT  74265.0 28015.0 74970.0 29360.0 ;
      RECT  74265.0 30705.0 74970.0 29360.0 ;
      RECT  74265.0 30705.0 74970.0 32050.0 ;
      RECT  74265.0 33395.0 74970.0 32050.0 ;
      RECT  74265.0 33395.0 74970.0 34740.0 ;
      RECT  74265.0 36085.0 74970.0 34740.0 ;
      RECT  74265.0 36085.0 74970.0 37430.0 ;
      RECT  74265.0 38775.0 74970.0 37430.0 ;
      RECT  74265.0 38775.0 74970.0 40120.0 ;
      RECT  74265.0 41465.0 74970.0 40120.0 ;
      RECT  74265.0 41465.0 74970.0 42810.0 ;
      RECT  74265.0 44155.0 74970.0 42810.0 ;
      RECT  74265.0 44155.0 74970.0 45500.0 ;
      RECT  74265.0 46845.0 74970.0 45500.0 ;
      RECT  74265.0 46845.0 74970.0 48190.0 ;
      RECT  74265.0 49535.0 74970.0 48190.0 ;
      RECT  74265.0 49535.0 74970.0 50880.0 ;
      RECT  74265.0 52225.0 74970.0 50880.0 ;
      RECT  74265.0 52225.0 74970.0 53570.0 ;
      RECT  74265.0 54915.0 74970.0 53570.0 ;
      RECT  74265.0 54915.0 74970.0 56260.0 ;
      RECT  74265.0 57605.0 74970.0 56260.0 ;
      RECT  74265.0 57605.0 74970.0 58950.0 ;
      RECT  74265.0 60295.0 74970.0 58950.0 ;
      RECT  74265.0 60295.0 74970.0 61640.0 ;
      RECT  74265.0 62985.0 74970.0 61640.0 ;
      RECT  74265.0 62985.0 74970.0 64330.0 ;
      RECT  74265.0 65675.0 74970.0 64330.0 ;
      RECT  74265.0 65675.0 74970.0 67020.0 ;
      RECT  74265.0 68365.0 74970.0 67020.0 ;
      RECT  74265.0 68365.0 74970.0 69710.0 ;
      RECT  74265.0 71055.0 74970.0 69710.0 ;
      RECT  74265.0 71055.0 74970.0 72400.0 ;
      RECT  74265.0 73745.0 74970.0 72400.0 ;
      RECT  74265.0 73745.0 74970.0 75090.0 ;
      RECT  74265.0 76435.0 74970.0 75090.0 ;
      RECT  74265.0 76435.0 74970.0 77780.0 ;
      RECT  74265.0 79125.0 74970.0 77780.0 ;
      RECT  74265.0 79125.0 74970.0 80470.0 ;
      RECT  74265.0 81815.0 74970.0 80470.0 ;
      RECT  74265.0 81815.0 74970.0 83160.0 ;
      RECT  74265.0 84505.0 74970.0 83160.0 ;
      RECT  74265.0 84505.0 74970.0 85850.0 ;
      RECT  74265.0 87195.0 74970.0 85850.0 ;
      RECT  74265.0 87195.0 74970.0 88540.0 ;
      RECT  74265.0 89885.0 74970.0 88540.0 ;
      RECT  74265.0 89885.0 74970.0 91230.0 ;
      RECT  74265.0 92575.0 74970.0 91230.0 ;
      RECT  74265.0 92575.0 74970.0 93920.0 ;
      RECT  74265.0 95265.0 74970.0 93920.0 ;
      RECT  74265.0 95265.0 74970.0 96610.0 ;
      RECT  74265.0 97955.0 74970.0 96610.0 ;
      RECT  74265.0 97955.0 74970.0 99300.0 ;
      RECT  74265.0 100645.0 74970.0 99300.0 ;
      RECT  74265.0 100645.0 74970.0 101990.0 ;
      RECT  74265.0 103335.0 74970.0 101990.0 ;
      RECT  74265.0 103335.0 74970.0 104680.0 ;
      RECT  74265.0 106025.0 74970.0 104680.0 ;
      RECT  74265.0 106025.0 74970.0 107370.0 ;
      RECT  74265.0 108715.0 74970.0 107370.0 ;
      RECT  74265.0 108715.0 74970.0 110060.0 ;
      RECT  74265.0 111405.0 74970.0 110060.0 ;
      RECT  74265.0 111405.0 74970.0 112750.0 ;
      RECT  74265.0 114095.0 74970.0 112750.0 ;
      RECT  74970.0 28015.0 75675.0 29360.0 ;
      RECT  74970.0 30705.0 75675.0 29360.0 ;
      RECT  74970.0 30705.0 75675.0 32050.0 ;
      RECT  74970.0 33395.0 75675.0 32050.0 ;
      RECT  74970.0 33395.0 75675.0 34740.0 ;
      RECT  74970.0 36085.0 75675.0 34740.0 ;
      RECT  74970.0 36085.0 75675.0 37430.0 ;
      RECT  74970.0 38775.0 75675.0 37430.0 ;
      RECT  74970.0 38775.0 75675.0 40120.0 ;
      RECT  74970.0 41465.0 75675.0 40120.0 ;
      RECT  74970.0 41465.0 75675.0 42810.0 ;
      RECT  74970.0 44155.0 75675.0 42810.0 ;
      RECT  74970.0 44155.0 75675.0 45500.0 ;
      RECT  74970.0 46845.0 75675.0 45500.0 ;
      RECT  74970.0 46845.0 75675.0 48190.0 ;
      RECT  74970.0 49535.0 75675.0 48190.0 ;
      RECT  74970.0 49535.0 75675.0 50880.0 ;
      RECT  74970.0 52225.0 75675.0 50880.0 ;
      RECT  74970.0 52225.0 75675.0 53570.0 ;
      RECT  74970.0 54915.0 75675.0 53570.0 ;
      RECT  74970.0 54915.0 75675.0 56260.0 ;
      RECT  74970.0 57605.0 75675.0 56260.0 ;
      RECT  74970.0 57605.0 75675.0 58950.0 ;
      RECT  74970.0 60295.0 75675.0 58950.0 ;
      RECT  74970.0 60295.0 75675.0 61640.0 ;
      RECT  74970.0 62985.0 75675.0 61640.0 ;
      RECT  74970.0 62985.0 75675.0 64330.0 ;
      RECT  74970.0 65675.0 75675.0 64330.0 ;
      RECT  74970.0 65675.0 75675.0 67020.0 ;
      RECT  74970.0 68365.0 75675.0 67020.0 ;
      RECT  74970.0 68365.0 75675.0 69710.0 ;
      RECT  74970.0 71055.0 75675.0 69710.0 ;
      RECT  74970.0 71055.0 75675.0 72400.0 ;
      RECT  74970.0 73745.0 75675.0 72400.0 ;
      RECT  74970.0 73745.0 75675.0 75090.0 ;
      RECT  74970.0 76435.0 75675.0 75090.0 ;
      RECT  74970.0 76435.0 75675.0 77780.0 ;
      RECT  74970.0 79125.0 75675.0 77780.0 ;
      RECT  74970.0 79125.0 75675.0 80470.0 ;
      RECT  74970.0 81815.0 75675.0 80470.0 ;
      RECT  74970.0 81815.0 75675.0 83160.0 ;
      RECT  74970.0 84505.0 75675.0 83160.0 ;
      RECT  74970.0 84505.0 75675.0 85850.0 ;
      RECT  74970.0 87195.0 75675.0 85850.0 ;
      RECT  74970.0 87195.0 75675.0 88540.0 ;
      RECT  74970.0 89885.0 75675.0 88540.0 ;
      RECT  74970.0 89885.0 75675.0 91230.0 ;
      RECT  74970.0 92575.0 75675.0 91230.0 ;
      RECT  74970.0 92575.0 75675.0 93920.0 ;
      RECT  74970.0 95265.0 75675.0 93920.0 ;
      RECT  74970.0 95265.0 75675.0 96610.0 ;
      RECT  74970.0 97955.0 75675.0 96610.0 ;
      RECT  74970.0 97955.0 75675.0 99300.0 ;
      RECT  74970.0 100645.0 75675.0 99300.0 ;
      RECT  74970.0 100645.0 75675.0 101990.0 ;
      RECT  74970.0 103335.0 75675.0 101990.0 ;
      RECT  74970.0 103335.0 75675.0 104680.0 ;
      RECT  74970.0 106025.0 75675.0 104680.0 ;
      RECT  74970.0 106025.0 75675.0 107370.0 ;
      RECT  74970.0 108715.0 75675.0 107370.0 ;
      RECT  74970.0 108715.0 75675.0 110060.0 ;
      RECT  74970.0 111405.0 75675.0 110060.0 ;
      RECT  74970.0 111405.0 75675.0 112750.0 ;
      RECT  74970.0 114095.0 75675.0 112750.0 ;
      RECT  75675.0 28015.0 76380.0 29360.0 ;
      RECT  75675.0 30705.0 76380.0 29360.0 ;
      RECT  75675.0 30705.0 76380.0 32050.0 ;
      RECT  75675.0 33395.0 76380.0 32050.0 ;
      RECT  75675.0 33395.0 76380.0 34740.0 ;
      RECT  75675.0 36085.0 76380.0 34740.0 ;
      RECT  75675.0 36085.0 76380.0 37430.0 ;
      RECT  75675.0 38775.0 76380.0 37430.0 ;
      RECT  75675.0 38775.0 76380.0 40120.0 ;
      RECT  75675.0 41465.0 76380.0 40120.0 ;
      RECT  75675.0 41465.0 76380.0 42810.0 ;
      RECT  75675.0 44155.0 76380.0 42810.0 ;
      RECT  75675.0 44155.0 76380.0 45500.0 ;
      RECT  75675.0 46845.0 76380.0 45500.0 ;
      RECT  75675.0 46845.0 76380.0 48190.0 ;
      RECT  75675.0 49535.0 76380.0 48190.0 ;
      RECT  75675.0 49535.0 76380.0 50880.0 ;
      RECT  75675.0 52225.0 76380.0 50880.0 ;
      RECT  75675.0 52225.0 76380.0 53570.0 ;
      RECT  75675.0 54915.0 76380.0 53570.0 ;
      RECT  75675.0 54915.0 76380.0 56260.0 ;
      RECT  75675.0 57605.0 76380.0 56260.0 ;
      RECT  75675.0 57605.0 76380.0 58950.0 ;
      RECT  75675.0 60295.0 76380.0 58950.0 ;
      RECT  75675.0 60295.0 76380.0 61640.0 ;
      RECT  75675.0 62985.0 76380.0 61640.0 ;
      RECT  75675.0 62985.0 76380.0 64330.0 ;
      RECT  75675.0 65675.0 76380.0 64330.0 ;
      RECT  75675.0 65675.0 76380.0 67020.0 ;
      RECT  75675.0 68365.0 76380.0 67020.0 ;
      RECT  75675.0 68365.0 76380.0 69710.0 ;
      RECT  75675.0 71055.0 76380.0 69710.0 ;
      RECT  75675.0 71055.0 76380.0 72400.0 ;
      RECT  75675.0 73745.0 76380.0 72400.0 ;
      RECT  75675.0 73745.0 76380.0 75090.0 ;
      RECT  75675.0 76435.0 76380.0 75090.0 ;
      RECT  75675.0 76435.0 76380.0 77780.0 ;
      RECT  75675.0 79125.0 76380.0 77780.0 ;
      RECT  75675.0 79125.0 76380.0 80470.0 ;
      RECT  75675.0 81815.0 76380.0 80470.0 ;
      RECT  75675.0 81815.0 76380.0 83160.0 ;
      RECT  75675.0 84505.0 76380.0 83160.0 ;
      RECT  75675.0 84505.0 76380.0 85850.0 ;
      RECT  75675.0 87195.0 76380.0 85850.0 ;
      RECT  75675.0 87195.0 76380.0 88540.0 ;
      RECT  75675.0 89885.0 76380.0 88540.0 ;
      RECT  75675.0 89885.0 76380.0 91230.0 ;
      RECT  75675.0 92575.0 76380.0 91230.0 ;
      RECT  75675.0 92575.0 76380.0 93920.0 ;
      RECT  75675.0 95265.0 76380.0 93920.0 ;
      RECT  75675.0 95265.0 76380.0 96610.0 ;
      RECT  75675.0 97955.0 76380.0 96610.0 ;
      RECT  75675.0 97955.0 76380.0 99300.0 ;
      RECT  75675.0 100645.0 76380.0 99300.0 ;
      RECT  75675.0 100645.0 76380.0 101990.0 ;
      RECT  75675.0 103335.0 76380.0 101990.0 ;
      RECT  75675.0 103335.0 76380.0 104680.0 ;
      RECT  75675.0 106025.0 76380.0 104680.0 ;
      RECT  75675.0 106025.0 76380.0 107370.0 ;
      RECT  75675.0 108715.0 76380.0 107370.0 ;
      RECT  75675.0 108715.0 76380.0 110060.0 ;
      RECT  75675.0 111405.0 76380.0 110060.0 ;
      RECT  75675.0 111405.0 76380.0 112750.0 ;
      RECT  75675.0 114095.0 76380.0 112750.0 ;
      RECT  76380.0 28015.0 77085.0 29360.0 ;
      RECT  76380.0 30705.0 77085.0 29360.0 ;
      RECT  76380.0 30705.0 77085.0 32050.0 ;
      RECT  76380.0 33395.0 77085.0 32050.0 ;
      RECT  76380.0 33395.0 77085.0 34740.0 ;
      RECT  76380.0 36085.0 77085.0 34740.0 ;
      RECT  76380.0 36085.0 77085.0 37430.0 ;
      RECT  76380.0 38775.0 77085.0 37430.0 ;
      RECT  76380.0 38775.0 77085.0 40120.0 ;
      RECT  76380.0 41465.0 77085.0 40120.0 ;
      RECT  76380.0 41465.0 77085.0 42810.0 ;
      RECT  76380.0 44155.0 77085.0 42810.0 ;
      RECT  76380.0 44155.0 77085.0 45500.0 ;
      RECT  76380.0 46845.0 77085.0 45500.0 ;
      RECT  76380.0 46845.0 77085.0 48190.0 ;
      RECT  76380.0 49535.0 77085.0 48190.0 ;
      RECT  76380.0 49535.0 77085.0 50880.0 ;
      RECT  76380.0 52225.0 77085.0 50880.0 ;
      RECT  76380.0 52225.0 77085.0 53570.0 ;
      RECT  76380.0 54915.0 77085.0 53570.0 ;
      RECT  76380.0 54915.0 77085.0 56260.0 ;
      RECT  76380.0 57605.0 77085.0 56260.0 ;
      RECT  76380.0 57605.0 77085.0 58950.0 ;
      RECT  76380.0 60295.0 77085.0 58950.0 ;
      RECT  76380.0 60295.0 77085.0 61640.0 ;
      RECT  76380.0 62985.0 77085.0 61640.0 ;
      RECT  76380.0 62985.0 77085.0 64330.0 ;
      RECT  76380.0 65675.0 77085.0 64330.0 ;
      RECT  76380.0 65675.0 77085.0 67020.0 ;
      RECT  76380.0 68365.0 77085.0 67020.0 ;
      RECT  76380.0 68365.0 77085.0 69710.0 ;
      RECT  76380.0 71055.0 77085.0 69710.0 ;
      RECT  76380.0 71055.0 77085.0 72400.0 ;
      RECT  76380.0 73745.0 77085.0 72400.0 ;
      RECT  76380.0 73745.0 77085.0 75090.0 ;
      RECT  76380.0 76435.0 77085.0 75090.0 ;
      RECT  76380.0 76435.0 77085.0 77780.0 ;
      RECT  76380.0 79125.0 77085.0 77780.0 ;
      RECT  76380.0 79125.0 77085.0 80470.0 ;
      RECT  76380.0 81815.0 77085.0 80470.0 ;
      RECT  76380.0 81815.0 77085.0 83160.0 ;
      RECT  76380.0 84505.0 77085.0 83160.0 ;
      RECT  76380.0 84505.0 77085.0 85850.0 ;
      RECT  76380.0 87195.0 77085.0 85850.0 ;
      RECT  76380.0 87195.0 77085.0 88540.0 ;
      RECT  76380.0 89885.0 77085.0 88540.0 ;
      RECT  76380.0 89885.0 77085.0 91230.0 ;
      RECT  76380.0 92575.0 77085.0 91230.0 ;
      RECT  76380.0 92575.0 77085.0 93920.0 ;
      RECT  76380.0 95265.0 77085.0 93920.0 ;
      RECT  76380.0 95265.0 77085.0 96610.0 ;
      RECT  76380.0 97955.0 77085.0 96610.0 ;
      RECT  76380.0 97955.0 77085.0 99300.0 ;
      RECT  76380.0 100645.0 77085.0 99300.0 ;
      RECT  76380.0 100645.0 77085.0 101990.0 ;
      RECT  76380.0 103335.0 77085.0 101990.0 ;
      RECT  76380.0 103335.0 77085.0 104680.0 ;
      RECT  76380.0 106025.0 77085.0 104680.0 ;
      RECT  76380.0 106025.0 77085.0 107370.0 ;
      RECT  76380.0 108715.0 77085.0 107370.0 ;
      RECT  76380.0 108715.0 77085.0 110060.0 ;
      RECT  76380.0 111405.0 77085.0 110060.0 ;
      RECT  76380.0 111405.0 77085.0 112750.0 ;
      RECT  76380.0 114095.0 77085.0 112750.0 ;
      RECT  77085.0 28015.0 77790.0 29360.0 ;
      RECT  77085.0 30705.0 77790.0 29360.0 ;
      RECT  77085.0 30705.0 77790.0 32050.0 ;
      RECT  77085.0 33395.0 77790.0 32050.0 ;
      RECT  77085.0 33395.0 77790.0 34740.0 ;
      RECT  77085.0 36085.0 77790.0 34740.0 ;
      RECT  77085.0 36085.0 77790.0 37430.0 ;
      RECT  77085.0 38775.0 77790.0 37430.0 ;
      RECT  77085.0 38775.0 77790.0 40120.0 ;
      RECT  77085.0 41465.0 77790.0 40120.0 ;
      RECT  77085.0 41465.0 77790.0 42810.0 ;
      RECT  77085.0 44155.0 77790.0 42810.0 ;
      RECT  77085.0 44155.0 77790.0 45500.0 ;
      RECT  77085.0 46845.0 77790.0 45500.0 ;
      RECT  77085.0 46845.0 77790.0 48190.0 ;
      RECT  77085.0 49535.0 77790.0 48190.0 ;
      RECT  77085.0 49535.0 77790.0 50880.0 ;
      RECT  77085.0 52225.0 77790.0 50880.0 ;
      RECT  77085.0 52225.0 77790.0 53570.0 ;
      RECT  77085.0 54915.0 77790.0 53570.0 ;
      RECT  77085.0 54915.0 77790.0 56260.0 ;
      RECT  77085.0 57605.0 77790.0 56260.0 ;
      RECT  77085.0 57605.0 77790.0 58950.0 ;
      RECT  77085.0 60295.0 77790.0 58950.0 ;
      RECT  77085.0 60295.0 77790.0 61640.0 ;
      RECT  77085.0 62985.0 77790.0 61640.0 ;
      RECT  77085.0 62985.0 77790.0 64330.0 ;
      RECT  77085.0 65675.0 77790.0 64330.0 ;
      RECT  77085.0 65675.0 77790.0 67020.0 ;
      RECT  77085.0 68365.0 77790.0 67020.0 ;
      RECT  77085.0 68365.0 77790.0 69710.0 ;
      RECT  77085.0 71055.0 77790.0 69710.0 ;
      RECT  77085.0 71055.0 77790.0 72400.0 ;
      RECT  77085.0 73745.0 77790.0 72400.0 ;
      RECT  77085.0 73745.0 77790.0 75090.0 ;
      RECT  77085.0 76435.0 77790.0 75090.0 ;
      RECT  77085.0 76435.0 77790.0 77780.0 ;
      RECT  77085.0 79125.0 77790.0 77780.0 ;
      RECT  77085.0 79125.0 77790.0 80470.0 ;
      RECT  77085.0 81815.0 77790.0 80470.0 ;
      RECT  77085.0 81815.0 77790.0 83160.0 ;
      RECT  77085.0 84505.0 77790.0 83160.0 ;
      RECT  77085.0 84505.0 77790.0 85850.0 ;
      RECT  77085.0 87195.0 77790.0 85850.0 ;
      RECT  77085.0 87195.0 77790.0 88540.0 ;
      RECT  77085.0 89885.0 77790.0 88540.0 ;
      RECT  77085.0 89885.0 77790.0 91230.0 ;
      RECT  77085.0 92575.0 77790.0 91230.0 ;
      RECT  77085.0 92575.0 77790.0 93920.0 ;
      RECT  77085.0 95265.0 77790.0 93920.0 ;
      RECT  77085.0 95265.0 77790.0 96610.0 ;
      RECT  77085.0 97955.0 77790.0 96610.0 ;
      RECT  77085.0 97955.0 77790.0 99300.0 ;
      RECT  77085.0 100645.0 77790.0 99300.0 ;
      RECT  77085.0 100645.0 77790.0 101990.0 ;
      RECT  77085.0 103335.0 77790.0 101990.0 ;
      RECT  77085.0 103335.0 77790.0 104680.0 ;
      RECT  77085.0 106025.0 77790.0 104680.0 ;
      RECT  77085.0 106025.0 77790.0 107370.0 ;
      RECT  77085.0 108715.0 77790.0 107370.0 ;
      RECT  77085.0 108715.0 77790.0 110060.0 ;
      RECT  77085.0 111405.0 77790.0 110060.0 ;
      RECT  77085.0 111405.0 77790.0 112750.0 ;
      RECT  77085.0 114095.0 77790.0 112750.0 ;
      RECT  77790.0 28015.0 78495.0 29360.0 ;
      RECT  77790.0 30705.0 78495.0 29360.0 ;
      RECT  77790.0 30705.0 78495.0 32050.0 ;
      RECT  77790.0 33395.0 78495.0 32050.0 ;
      RECT  77790.0 33395.0 78495.0 34740.0 ;
      RECT  77790.0 36085.0 78495.0 34740.0 ;
      RECT  77790.0 36085.0 78495.0 37430.0 ;
      RECT  77790.0 38775.0 78495.0 37430.0 ;
      RECT  77790.0 38775.0 78495.0 40120.0 ;
      RECT  77790.0 41465.0 78495.0 40120.0 ;
      RECT  77790.0 41465.0 78495.0 42810.0 ;
      RECT  77790.0 44155.0 78495.0 42810.0 ;
      RECT  77790.0 44155.0 78495.0 45500.0 ;
      RECT  77790.0 46845.0 78495.0 45500.0 ;
      RECT  77790.0 46845.0 78495.0 48190.0 ;
      RECT  77790.0 49535.0 78495.0 48190.0 ;
      RECT  77790.0 49535.0 78495.0 50880.0 ;
      RECT  77790.0 52225.0 78495.0 50880.0 ;
      RECT  77790.0 52225.0 78495.0 53570.0 ;
      RECT  77790.0 54915.0 78495.0 53570.0 ;
      RECT  77790.0 54915.0 78495.0 56260.0 ;
      RECT  77790.0 57605.0 78495.0 56260.0 ;
      RECT  77790.0 57605.0 78495.0 58950.0 ;
      RECT  77790.0 60295.0 78495.0 58950.0 ;
      RECT  77790.0 60295.0 78495.0 61640.0 ;
      RECT  77790.0 62985.0 78495.0 61640.0 ;
      RECT  77790.0 62985.0 78495.0 64330.0 ;
      RECT  77790.0 65675.0 78495.0 64330.0 ;
      RECT  77790.0 65675.0 78495.0 67020.0 ;
      RECT  77790.0 68365.0 78495.0 67020.0 ;
      RECT  77790.0 68365.0 78495.0 69710.0 ;
      RECT  77790.0 71055.0 78495.0 69710.0 ;
      RECT  77790.0 71055.0 78495.0 72400.0 ;
      RECT  77790.0 73745.0 78495.0 72400.0 ;
      RECT  77790.0 73745.0 78495.0 75090.0 ;
      RECT  77790.0 76435.0 78495.0 75090.0 ;
      RECT  77790.0 76435.0 78495.0 77780.0 ;
      RECT  77790.0 79125.0 78495.0 77780.0 ;
      RECT  77790.0 79125.0 78495.0 80470.0 ;
      RECT  77790.0 81815.0 78495.0 80470.0 ;
      RECT  77790.0 81815.0 78495.0 83160.0 ;
      RECT  77790.0 84505.0 78495.0 83160.0 ;
      RECT  77790.0 84505.0 78495.0 85850.0 ;
      RECT  77790.0 87195.0 78495.0 85850.0 ;
      RECT  77790.0 87195.0 78495.0 88540.0 ;
      RECT  77790.0 89885.0 78495.0 88540.0 ;
      RECT  77790.0 89885.0 78495.0 91230.0 ;
      RECT  77790.0 92575.0 78495.0 91230.0 ;
      RECT  77790.0 92575.0 78495.0 93920.0 ;
      RECT  77790.0 95265.0 78495.0 93920.0 ;
      RECT  77790.0 95265.0 78495.0 96610.0 ;
      RECT  77790.0 97955.0 78495.0 96610.0 ;
      RECT  77790.0 97955.0 78495.0 99300.0 ;
      RECT  77790.0 100645.0 78495.0 99300.0 ;
      RECT  77790.0 100645.0 78495.0 101990.0 ;
      RECT  77790.0 103335.0 78495.0 101990.0 ;
      RECT  77790.0 103335.0 78495.0 104680.0 ;
      RECT  77790.0 106025.0 78495.0 104680.0 ;
      RECT  77790.0 106025.0 78495.0 107370.0 ;
      RECT  77790.0 108715.0 78495.0 107370.0 ;
      RECT  77790.0 108715.0 78495.0 110060.0 ;
      RECT  77790.0 111405.0 78495.0 110060.0 ;
      RECT  77790.0 111405.0 78495.0 112750.0 ;
      RECT  77790.0 114095.0 78495.0 112750.0 ;
      RECT  78495.0 28015.0 79200.0 29360.0 ;
      RECT  78495.0 30705.0 79200.0 29360.0 ;
      RECT  78495.0 30705.0 79200.0 32050.0 ;
      RECT  78495.0 33395.0 79200.0 32050.0 ;
      RECT  78495.0 33395.0 79200.0 34740.0 ;
      RECT  78495.0 36085.0 79200.0 34740.0 ;
      RECT  78495.0 36085.0 79200.0 37430.0 ;
      RECT  78495.0 38775.0 79200.0 37430.0 ;
      RECT  78495.0 38775.0 79200.0 40120.0 ;
      RECT  78495.0 41465.0 79200.0 40120.0 ;
      RECT  78495.0 41465.0 79200.0 42810.0 ;
      RECT  78495.0 44155.0 79200.0 42810.0 ;
      RECT  78495.0 44155.0 79200.0 45500.0 ;
      RECT  78495.0 46845.0 79200.0 45500.0 ;
      RECT  78495.0 46845.0 79200.0 48190.0 ;
      RECT  78495.0 49535.0 79200.0 48190.0 ;
      RECT  78495.0 49535.0 79200.0 50880.0 ;
      RECT  78495.0 52225.0 79200.0 50880.0 ;
      RECT  78495.0 52225.0 79200.0 53570.0 ;
      RECT  78495.0 54915.0 79200.0 53570.0 ;
      RECT  78495.0 54915.0 79200.0 56260.0 ;
      RECT  78495.0 57605.0 79200.0 56260.0 ;
      RECT  78495.0 57605.0 79200.0 58950.0 ;
      RECT  78495.0 60295.0 79200.0 58950.0 ;
      RECT  78495.0 60295.0 79200.0 61640.0 ;
      RECT  78495.0 62985.0 79200.0 61640.0 ;
      RECT  78495.0 62985.0 79200.0 64330.0 ;
      RECT  78495.0 65675.0 79200.0 64330.0 ;
      RECT  78495.0 65675.0 79200.0 67020.0 ;
      RECT  78495.0 68365.0 79200.0 67020.0 ;
      RECT  78495.0 68365.0 79200.0 69710.0 ;
      RECT  78495.0 71055.0 79200.0 69710.0 ;
      RECT  78495.0 71055.0 79200.0 72400.0 ;
      RECT  78495.0 73745.0 79200.0 72400.0 ;
      RECT  78495.0 73745.0 79200.0 75090.0 ;
      RECT  78495.0 76435.0 79200.0 75090.0 ;
      RECT  78495.0 76435.0 79200.0 77780.0 ;
      RECT  78495.0 79125.0 79200.0 77780.0 ;
      RECT  78495.0 79125.0 79200.0 80470.0 ;
      RECT  78495.0 81815.0 79200.0 80470.0 ;
      RECT  78495.0 81815.0 79200.0 83160.0 ;
      RECT  78495.0 84505.0 79200.0 83160.0 ;
      RECT  78495.0 84505.0 79200.0 85850.0 ;
      RECT  78495.0 87195.0 79200.0 85850.0 ;
      RECT  78495.0 87195.0 79200.0 88540.0 ;
      RECT  78495.0 89885.0 79200.0 88540.0 ;
      RECT  78495.0 89885.0 79200.0 91230.0 ;
      RECT  78495.0 92575.0 79200.0 91230.0 ;
      RECT  78495.0 92575.0 79200.0 93920.0 ;
      RECT  78495.0 95265.0 79200.0 93920.0 ;
      RECT  78495.0 95265.0 79200.0 96610.0 ;
      RECT  78495.0 97955.0 79200.0 96610.0 ;
      RECT  78495.0 97955.0 79200.0 99300.0 ;
      RECT  78495.0 100645.0 79200.0 99300.0 ;
      RECT  78495.0 100645.0 79200.0 101990.0 ;
      RECT  78495.0 103335.0 79200.0 101990.0 ;
      RECT  78495.0 103335.0 79200.0 104680.0 ;
      RECT  78495.0 106025.0 79200.0 104680.0 ;
      RECT  78495.0 106025.0 79200.0 107370.0 ;
      RECT  78495.0 108715.0 79200.0 107370.0 ;
      RECT  78495.0 108715.0 79200.0 110060.0 ;
      RECT  78495.0 111405.0 79200.0 110060.0 ;
      RECT  78495.0 111405.0 79200.0 112750.0 ;
      RECT  78495.0 114095.0 79200.0 112750.0 ;
      RECT  79200.0 28015.0 79905.0 29360.0 ;
      RECT  79200.0 30705.0 79905.0 29360.0 ;
      RECT  79200.0 30705.0 79905.0 32050.0 ;
      RECT  79200.0 33395.0 79905.0 32050.0 ;
      RECT  79200.0 33395.0 79905.0 34740.0 ;
      RECT  79200.0 36085.0 79905.0 34740.0 ;
      RECT  79200.0 36085.0 79905.0 37430.0 ;
      RECT  79200.0 38775.0 79905.0 37430.0 ;
      RECT  79200.0 38775.0 79905.0 40120.0 ;
      RECT  79200.0 41465.0 79905.0 40120.0 ;
      RECT  79200.0 41465.0 79905.0 42810.0 ;
      RECT  79200.0 44155.0 79905.0 42810.0 ;
      RECT  79200.0 44155.0 79905.0 45500.0 ;
      RECT  79200.0 46845.0 79905.0 45500.0 ;
      RECT  79200.0 46845.0 79905.0 48190.0 ;
      RECT  79200.0 49535.0 79905.0 48190.0 ;
      RECT  79200.0 49535.0 79905.0 50880.0 ;
      RECT  79200.0 52225.0 79905.0 50880.0 ;
      RECT  79200.0 52225.0 79905.0 53570.0 ;
      RECT  79200.0 54915.0 79905.0 53570.0 ;
      RECT  79200.0 54915.0 79905.0 56260.0 ;
      RECT  79200.0 57605.0 79905.0 56260.0 ;
      RECT  79200.0 57605.0 79905.0 58950.0 ;
      RECT  79200.0 60295.0 79905.0 58950.0 ;
      RECT  79200.0 60295.0 79905.0 61640.0 ;
      RECT  79200.0 62985.0 79905.0 61640.0 ;
      RECT  79200.0 62985.0 79905.0 64330.0 ;
      RECT  79200.0 65675.0 79905.0 64330.0 ;
      RECT  79200.0 65675.0 79905.0 67020.0 ;
      RECT  79200.0 68365.0 79905.0 67020.0 ;
      RECT  79200.0 68365.0 79905.0 69710.0 ;
      RECT  79200.0 71055.0 79905.0 69710.0 ;
      RECT  79200.0 71055.0 79905.0 72400.0 ;
      RECT  79200.0 73745.0 79905.0 72400.0 ;
      RECT  79200.0 73745.0 79905.0 75090.0 ;
      RECT  79200.0 76435.0 79905.0 75090.0 ;
      RECT  79200.0 76435.0 79905.0 77780.0 ;
      RECT  79200.0 79125.0 79905.0 77780.0 ;
      RECT  79200.0 79125.0 79905.0 80470.0 ;
      RECT  79200.0 81815.0 79905.0 80470.0 ;
      RECT  79200.0 81815.0 79905.0 83160.0 ;
      RECT  79200.0 84505.0 79905.0 83160.0 ;
      RECT  79200.0 84505.0 79905.0 85850.0 ;
      RECT  79200.0 87195.0 79905.0 85850.0 ;
      RECT  79200.0 87195.0 79905.0 88540.0 ;
      RECT  79200.0 89885.0 79905.0 88540.0 ;
      RECT  79200.0 89885.0 79905.0 91230.0 ;
      RECT  79200.0 92575.0 79905.0 91230.0 ;
      RECT  79200.0 92575.0 79905.0 93920.0 ;
      RECT  79200.0 95265.0 79905.0 93920.0 ;
      RECT  79200.0 95265.0 79905.0 96610.0 ;
      RECT  79200.0 97955.0 79905.0 96610.0 ;
      RECT  79200.0 97955.0 79905.0 99300.0 ;
      RECT  79200.0 100645.0 79905.0 99300.0 ;
      RECT  79200.0 100645.0 79905.0 101990.0 ;
      RECT  79200.0 103335.0 79905.0 101990.0 ;
      RECT  79200.0 103335.0 79905.0 104680.0 ;
      RECT  79200.0 106025.0 79905.0 104680.0 ;
      RECT  79200.0 106025.0 79905.0 107370.0 ;
      RECT  79200.0 108715.0 79905.0 107370.0 ;
      RECT  79200.0 108715.0 79905.0 110060.0 ;
      RECT  79200.0 111405.0 79905.0 110060.0 ;
      RECT  79200.0 111405.0 79905.0 112750.0 ;
      RECT  79200.0 114095.0 79905.0 112750.0 ;
      RECT  79905.0 28015.0 80610.0 29360.0 ;
      RECT  79905.0 30705.0 80610.0 29360.0 ;
      RECT  79905.0 30705.0 80610.0 32050.0 ;
      RECT  79905.0 33395.0 80610.0 32050.0 ;
      RECT  79905.0 33395.0 80610.0 34740.0 ;
      RECT  79905.0 36085.0 80610.0 34740.0 ;
      RECT  79905.0 36085.0 80610.0 37430.0 ;
      RECT  79905.0 38775.0 80610.0 37430.0 ;
      RECT  79905.0 38775.0 80610.0 40120.0 ;
      RECT  79905.0 41465.0 80610.0 40120.0 ;
      RECT  79905.0 41465.0 80610.0 42810.0 ;
      RECT  79905.0 44155.0 80610.0 42810.0 ;
      RECT  79905.0 44155.0 80610.0 45500.0 ;
      RECT  79905.0 46845.0 80610.0 45500.0 ;
      RECT  79905.0 46845.0 80610.0 48190.0 ;
      RECT  79905.0 49535.0 80610.0 48190.0 ;
      RECT  79905.0 49535.0 80610.0 50880.0 ;
      RECT  79905.0 52225.0 80610.0 50880.0 ;
      RECT  79905.0 52225.0 80610.0 53570.0 ;
      RECT  79905.0 54915.0 80610.0 53570.0 ;
      RECT  79905.0 54915.0 80610.0 56260.0 ;
      RECT  79905.0 57605.0 80610.0 56260.0 ;
      RECT  79905.0 57605.0 80610.0 58950.0 ;
      RECT  79905.0 60295.0 80610.0 58950.0 ;
      RECT  79905.0 60295.0 80610.0 61640.0 ;
      RECT  79905.0 62985.0 80610.0 61640.0 ;
      RECT  79905.0 62985.0 80610.0 64330.0 ;
      RECT  79905.0 65675.0 80610.0 64330.0 ;
      RECT  79905.0 65675.0 80610.0 67020.0 ;
      RECT  79905.0 68365.0 80610.0 67020.0 ;
      RECT  79905.0 68365.0 80610.0 69710.0 ;
      RECT  79905.0 71055.0 80610.0 69710.0 ;
      RECT  79905.0 71055.0 80610.0 72400.0 ;
      RECT  79905.0 73745.0 80610.0 72400.0 ;
      RECT  79905.0 73745.0 80610.0 75090.0 ;
      RECT  79905.0 76435.0 80610.0 75090.0 ;
      RECT  79905.0 76435.0 80610.0 77780.0 ;
      RECT  79905.0 79125.0 80610.0 77780.0 ;
      RECT  79905.0 79125.0 80610.0 80470.0 ;
      RECT  79905.0 81815.0 80610.0 80470.0 ;
      RECT  79905.0 81815.0 80610.0 83160.0 ;
      RECT  79905.0 84505.0 80610.0 83160.0 ;
      RECT  79905.0 84505.0 80610.0 85850.0 ;
      RECT  79905.0 87195.0 80610.0 85850.0 ;
      RECT  79905.0 87195.0 80610.0 88540.0 ;
      RECT  79905.0 89885.0 80610.0 88540.0 ;
      RECT  79905.0 89885.0 80610.0 91230.0 ;
      RECT  79905.0 92575.0 80610.0 91230.0 ;
      RECT  79905.0 92575.0 80610.0 93920.0 ;
      RECT  79905.0 95265.0 80610.0 93920.0 ;
      RECT  79905.0 95265.0 80610.0 96610.0 ;
      RECT  79905.0 97955.0 80610.0 96610.0 ;
      RECT  79905.0 97955.0 80610.0 99300.0 ;
      RECT  79905.0 100645.0 80610.0 99300.0 ;
      RECT  79905.0 100645.0 80610.0 101990.0 ;
      RECT  79905.0 103335.0 80610.0 101990.0 ;
      RECT  79905.0 103335.0 80610.0 104680.0 ;
      RECT  79905.0 106025.0 80610.0 104680.0 ;
      RECT  79905.0 106025.0 80610.0 107370.0 ;
      RECT  79905.0 108715.0 80610.0 107370.0 ;
      RECT  79905.0 108715.0 80610.0 110060.0 ;
      RECT  79905.0 111405.0 80610.0 110060.0 ;
      RECT  79905.0 111405.0 80610.0 112750.0 ;
      RECT  79905.0 114095.0 80610.0 112750.0 ;
      RECT  80610.0 28015.0 81315.0 29360.0 ;
      RECT  80610.0 30705.0 81315.0 29360.0 ;
      RECT  80610.0 30705.0 81315.0 32050.0 ;
      RECT  80610.0 33395.0 81315.0 32050.0 ;
      RECT  80610.0 33395.0 81315.0 34740.0 ;
      RECT  80610.0 36085.0 81315.0 34740.0 ;
      RECT  80610.0 36085.0 81315.0 37430.0 ;
      RECT  80610.0 38775.0 81315.0 37430.0 ;
      RECT  80610.0 38775.0 81315.0 40120.0 ;
      RECT  80610.0 41465.0 81315.0 40120.0 ;
      RECT  80610.0 41465.0 81315.0 42810.0 ;
      RECT  80610.0 44155.0 81315.0 42810.0 ;
      RECT  80610.0 44155.0 81315.0 45500.0 ;
      RECT  80610.0 46845.0 81315.0 45500.0 ;
      RECT  80610.0 46845.0 81315.0 48190.0 ;
      RECT  80610.0 49535.0 81315.0 48190.0 ;
      RECT  80610.0 49535.0 81315.0 50880.0 ;
      RECT  80610.0 52225.0 81315.0 50880.0 ;
      RECT  80610.0 52225.0 81315.0 53570.0 ;
      RECT  80610.0 54915.0 81315.0 53570.0 ;
      RECT  80610.0 54915.0 81315.0 56260.0 ;
      RECT  80610.0 57605.0 81315.0 56260.0 ;
      RECT  80610.0 57605.0 81315.0 58950.0 ;
      RECT  80610.0 60295.0 81315.0 58950.0 ;
      RECT  80610.0 60295.0 81315.0 61640.0 ;
      RECT  80610.0 62985.0 81315.0 61640.0 ;
      RECT  80610.0 62985.0 81315.0 64330.0 ;
      RECT  80610.0 65675.0 81315.0 64330.0 ;
      RECT  80610.0 65675.0 81315.0 67020.0 ;
      RECT  80610.0 68365.0 81315.0 67020.0 ;
      RECT  80610.0 68365.0 81315.0 69710.0 ;
      RECT  80610.0 71055.0 81315.0 69710.0 ;
      RECT  80610.0 71055.0 81315.0 72400.0 ;
      RECT  80610.0 73745.0 81315.0 72400.0 ;
      RECT  80610.0 73745.0 81315.0 75090.0 ;
      RECT  80610.0 76435.0 81315.0 75090.0 ;
      RECT  80610.0 76435.0 81315.0 77780.0 ;
      RECT  80610.0 79125.0 81315.0 77780.0 ;
      RECT  80610.0 79125.0 81315.0 80470.0 ;
      RECT  80610.0 81815.0 81315.0 80470.0 ;
      RECT  80610.0 81815.0 81315.0 83160.0 ;
      RECT  80610.0 84505.0 81315.0 83160.0 ;
      RECT  80610.0 84505.0 81315.0 85850.0 ;
      RECT  80610.0 87195.0 81315.0 85850.0 ;
      RECT  80610.0 87195.0 81315.0 88540.0 ;
      RECT  80610.0 89885.0 81315.0 88540.0 ;
      RECT  80610.0 89885.0 81315.0 91230.0 ;
      RECT  80610.0 92575.0 81315.0 91230.0 ;
      RECT  80610.0 92575.0 81315.0 93920.0 ;
      RECT  80610.0 95265.0 81315.0 93920.0 ;
      RECT  80610.0 95265.0 81315.0 96610.0 ;
      RECT  80610.0 97955.0 81315.0 96610.0 ;
      RECT  80610.0 97955.0 81315.0 99300.0 ;
      RECT  80610.0 100645.0 81315.0 99300.0 ;
      RECT  80610.0 100645.0 81315.0 101990.0 ;
      RECT  80610.0 103335.0 81315.0 101990.0 ;
      RECT  80610.0 103335.0 81315.0 104680.0 ;
      RECT  80610.0 106025.0 81315.0 104680.0 ;
      RECT  80610.0 106025.0 81315.0 107370.0 ;
      RECT  80610.0 108715.0 81315.0 107370.0 ;
      RECT  80610.0 108715.0 81315.0 110060.0 ;
      RECT  80610.0 111405.0 81315.0 110060.0 ;
      RECT  80610.0 111405.0 81315.0 112750.0 ;
      RECT  80610.0 114095.0 81315.0 112750.0 ;
      RECT  81315.0 28015.0 82020.0 29360.0 ;
      RECT  81315.0 30705.0 82020.0 29360.0 ;
      RECT  81315.0 30705.0 82020.0 32050.0 ;
      RECT  81315.0 33395.0 82020.0 32050.0 ;
      RECT  81315.0 33395.0 82020.0 34740.0 ;
      RECT  81315.0 36085.0 82020.0 34740.0 ;
      RECT  81315.0 36085.0 82020.0 37430.0 ;
      RECT  81315.0 38775.0 82020.0 37430.0 ;
      RECT  81315.0 38775.0 82020.0 40120.0 ;
      RECT  81315.0 41465.0 82020.0 40120.0 ;
      RECT  81315.0 41465.0 82020.0 42810.0 ;
      RECT  81315.0 44155.0 82020.0 42810.0 ;
      RECT  81315.0 44155.0 82020.0 45500.0 ;
      RECT  81315.0 46845.0 82020.0 45500.0 ;
      RECT  81315.0 46845.0 82020.0 48190.0 ;
      RECT  81315.0 49535.0 82020.0 48190.0 ;
      RECT  81315.0 49535.0 82020.0 50880.0 ;
      RECT  81315.0 52225.0 82020.0 50880.0 ;
      RECT  81315.0 52225.0 82020.0 53570.0 ;
      RECT  81315.0 54915.0 82020.0 53570.0 ;
      RECT  81315.0 54915.0 82020.0 56260.0 ;
      RECT  81315.0 57605.0 82020.0 56260.0 ;
      RECT  81315.0 57605.0 82020.0 58950.0 ;
      RECT  81315.0 60295.0 82020.0 58950.0 ;
      RECT  81315.0 60295.0 82020.0 61640.0 ;
      RECT  81315.0 62985.0 82020.0 61640.0 ;
      RECT  81315.0 62985.0 82020.0 64330.0 ;
      RECT  81315.0 65675.0 82020.0 64330.0 ;
      RECT  81315.0 65675.0 82020.0 67020.0 ;
      RECT  81315.0 68365.0 82020.0 67020.0 ;
      RECT  81315.0 68365.0 82020.0 69710.0 ;
      RECT  81315.0 71055.0 82020.0 69710.0 ;
      RECT  81315.0 71055.0 82020.0 72400.0 ;
      RECT  81315.0 73745.0 82020.0 72400.0 ;
      RECT  81315.0 73745.0 82020.0 75090.0 ;
      RECT  81315.0 76435.0 82020.0 75090.0 ;
      RECT  81315.0 76435.0 82020.0 77780.0 ;
      RECT  81315.0 79125.0 82020.0 77780.0 ;
      RECT  81315.0 79125.0 82020.0 80470.0 ;
      RECT  81315.0 81815.0 82020.0 80470.0 ;
      RECT  81315.0 81815.0 82020.0 83160.0 ;
      RECT  81315.0 84505.0 82020.0 83160.0 ;
      RECT  81315.0 84505.0 82020.0 85850.0 ;
      RECT  81315.0 87195.0 82020.0 85850.0 ;
      RECT  81315.0 87195.0 82020.0 88540.0 ;
      RECT  81315.0 89885.0 82020.0 88540.0 ;
      RECT  81315.0 89885.0 82020.0 91230.0 ;
      RECT  81315.0 92575.0 82020.0 91230.0 ;
      RECT  81315.0 92575.0 82020.0 93920.0 ;
      RECT  81315.0 95265.0 82020.0 93920.0 ;
      RECT  81315.0 95265.0 82020.0 96610.0 ;
      RECT  81315.0 97955.0 82020.0 96610.0 ;
      RECT  81315.0 97955.0 82020.0 99300.0 ;
      RECT  81315.0 100645.0 82020.0 99300.0 ;
      RECT  81315.0 100645.0 82020.0 101990.0 ;
      RECT  81315.0 103335.0 82020.0 101990.0 ;
      RECT  81315.0 103335.0 82020.0 104680.0 ;
      RECT  81315.0 106025.0 82020.0 104680.0 ;
      RECT  81315.0 106025.0 82020.0 107370.0 ;
      RECT  81315.0 108715.0 82020.0 107370.0 ;
      RECT  81315.0 108715.0 82020.0 110060.0 ;
      RECT  81315.0 111405.0 82020.0 110060.0 ;
      RECT  81315.0 111405.0 82020.0 112750.0 ;
      RECT  81315.0 114095.0 82020.0 112750.0 ;
      RECT  82020.0 28015.0 82725.0 29360.0 ;
      RECT  82020.0 30705.0 82725.0 29360.0 ;
      RECT  82020.0 30705.0 82725.0 32050.0 ;
      RECT  82020.0 33395.0 82725.0 32050.0 ;
      RECT  82020.0 33395.0 82725.0 34740.0 ;
      RECT  82020.0 36085.0 82725.0 34740.0 ;
      RECT  82020.0 36085.0 82725.0 37430.0 ;
      RECT  82020.0 38775.0 82725.0 37430.0 ;
      RECT  82020.0 38775.0 82725.0 40120.0 ;
      RECT  82020.0 41465.0 82725.0 40120.0 ;
      RECT  82020.0 41465.0 82725.0 42810.0 ;
      RECT  82020.0 44155.0 82725.0 42810.0 ;
      RECT  82020.0 44155.0 82725.0 45500.0 ;
      RECT  82020.0 46845.0 82725.0 45500.0 ;
      RECT  82020.0 46845.0 82725.0 48190.0 ;
      RECT  82020.0 49535.0 82725.0 48190.0 ;
      RECT  82020.0 49535.0 82725.0 50880.0 ;
      RECT  82020.0 52225.0 82725.0 50880.0 ;
      RECT  82020.0 52225.0 82725.0 53570.0 ;
      RECT  82020.0 54915.0 82725.0 53570.0 ;
      RECT  82020.0 54915.0 82725.0 56260.0 ;
      RECT  82020.0 57605.0 82725.0 56260.0 ;
      RECT  82020.0 57605.0 82725.0 58950.0 ;
      RECT  82020.0 60295.0 82725.0 58950.0 ;
      RECT  82020.0 60295.0 82725.0 61640.0 ;
      RECT  82020.0 62985.0 82725.0 61640.0 ;
      RECT  82020.0 62985.0 82725.0 64330.0 ;
      RECT  82020.0 65675.0 82725.0 64330.0 ;
      RECT  82020.0 65675.0 82725.0 67020.0 ;
      RECT  82020.0 68365.0 82725.0 67020.0 ;
      RECT  82020.0 68365.0 82725.0 69710.0 ;
      RECT  82020.0 71055.0 82725.0 69710.0 ;
      RECT  82020.0 71055.0 82725.0 72400.0 ;
      RECT  82020.0 73745.0 82725.0 72400.0 ;
      RECT  82020.0 73745.0 82725.0 75090.0 ;
      RECT  82020.0 76435.0 82725.0 75090.0 ;
      RECT  82020.0 76435.0 82725.0 77780.0 ;
      RECT  82020.0 79125.0 82725.0 77780.0 ;
      RECT  82020.0 79125.0 82725.0 80470.0 ;
      RECT  82020.0 81815.0 82725.0 80470.0 ;
      RECT  82020.0 81815.0 82725.0 83160.0 ;
      RECT  82020.0 84505.0 82725.0 83160.0 ;
      RECT  82020.0 84505.0 82725.0 85850.0 ;
      RECT  82020.0 87195.0 82725.0 85850.0 ;
      RECT  82020.0 87195.0 82725.0 88540.0 ;
      RECT  82020.0 89885.0 82725.0 88540.0 ;
      RECT  82020.0 89885.0 82725.0 91230.0 ;
      RECT  82020.0 92575.0 82725.0 91230.0 ;
      RECT  82020.0 92575.0 82725.0 93920.0 ;
      RECT  82020.0 95265.0 82725.0 93920.0 ;
      RECT  82020.0 95265.0 82725.0 96610.0 ;
      RECT  82020.0 97955.0 82725.0 96610.0 ;
      RECT  82020.0 97955.0 82725.0 99300.0 ;
      RECT  82020.0 100645.0 82725.0 99300.0 ;
      RECT  82020.0 100645.0 82725.0 101990.0 ;
      RECT  82020.0 103335.0 82725.0 101990.0 ;
      RECT  82020.0 103335.0 82725.0 104680.0 ;
      RECT  82020.0 106025.0 82725.0 104680.0 ;
      RECT  82020.0 106025.0 82725.0 107370.0 ;
      RECT  82020.0 108715.0 82725.0 107370.0 ;
      RECT  82020.0 108715.0 82725.0 110060.0 ;
      RECT  82020.0 111405.0 82725.0 110060.0 ;
      RECT  82020.0 111405.0 82725.0 112750.0 ;
      RECT  82020.0 114095.0 82725.0 112750.0 ;
      RECT  82725.0 28015.0 83430.0 29360.0 ;
      RECT  82725.0 30705.0 83430.0 29360.0 ;
      RECT  82725.0 30705.0 83430.0 32050.0 ;
      RECT  82725.0 33395.0 83430.0 32050.0 ;
      RECT  82725.0 33395.0 83430.0 34740.0 ;
      RECT  82725.0 36085.0 83430.0 34740.0 ;
      RECT  82725.0 36085.0 83430.0 37430.0 ;
      RECT  82725.0 38775.0 83430.0 37430.0 ;
      RECT  82725.0 38775.0 83430.0 40120.0 ;
      RECT  82725.0 41465.0 83430.0 40120.0 ;
      RECT  82725.0 41465.0 83430.0 42810.0 ;
      RECT  82725.0 44155.0 83430.0 42810.0 ;
      RECT  82725.0 44155.0 83430.0 45500.0 ;
      RECT  82725.0 46845.0 83430.0 45500.0 ;
      RECT  82725.0 46845.0 83430.0 48190.0 ;
      RECT  82725.0 49535.0 83430.0 48190.0 ;
      RECT  82725.0 49535.0 83430.0 50880.0 ;
      RECT  82725.0 52225.0 83430.0 50880.0 ;
      RECT  82725.0 52225.0 83430.0 53570.0 ;
      RECT  82725.0 54915.0 83430.0 53570.0 ;
      RECT  82725.0 54915.0 83430.0 56260.0 ;
      RECT  82725.0 57605.0 83430.0 56260.0 ;
      RECT  82725.0 57605.0 83430.0 58950.0 ;
      RECT  82725.0 60295.0 83430.0 58950.0 ;
      RECT  82725.0 60295.0 83430.0 61640.0 ;
      RECT  82725.0 62985.0 83430.0 61640.0 ;
      RECT  82725.0 62985.0 83430.0 64330.0 ;
      RECT  82725.0 65675.0 83430.0 64330.0 ;
      RECT  82725.0 65675.0 83430.0 67020.0 ;
      RECT  82725.0 68365.0 83430.0 67020.0 ;
      RECT  82725.0 68365.0 83430.0 69710.0 ;
      RECT  82725.0 71055.0 83430.0 69710.0 ;
      RECT  82725.0 71055.0 83430.0 72400.0 ;
      RECT  82725.0 73745.0 83430.0 72400.0 ;
      RECT  82725.0 73745.0 83430.0 75090.0 ;
      RECT  82725.0 76435.0 83430.0 75090.0 ;
      RECT  82725.0 76435.0 83430.0 77780.0 ;
      RECT  82725.0 79125.0 83430.0 77780.0 ;
      RECT  82725.0 79125.0 83430.0 80470.0 ;
      RECT  82725.0 81815.0 83430.0 80470.0 ;
      RECT  82725.0 81815.0 83430.0 83160.0 ;
      RECT  82725.0 84505.0 83430.0 83160.0 ;
      RECT  82725.0 84505.0 83430.0 85850.0 ;
      RECT  82725.0 87195.0 83430.0 85850.0 ;
      RECT  82725.0 87195.0 83430.0 88540.0 ;
      RECT  82725.0 89885.0 83430.0 88540.0 ;
      RECT  82725.0 89885.0 83430.0 91230.0 ;
      RECT  82725.0 92575.0 83430.0 91230.0 ;
      RECT  82725.0 92575.0 83430.0 93920.0 ;
      RECT  82725.0 95265.0 83430.0 93920.0 ;
      RECT  82725.0 95265.0 83430.0 96610.0 ;
      RECT  82725.0 97955.0 83430.0 96610.0 ;
      RECT  82725.0 97955.0 83430.0 99300.0 ;
      RECT  82725.0 100645.0 83430.0 99300.0 ;
      RECT  82725.0 100645.0 83430.0 101990.0 ;
      RECT  82725.0 103335.0 83430.0 101990.0 ;
      RECT  82725.0 103335.0 83430.0 104680.0 ;
      RECT  82725.0 106025.0 83430.0 104680.0 ;
      RECT  82725.0 106025.0 83430.0 107370.0 ;
      RECT  82725.0 108715.0 83430.0 107370.0 ;
      RECT  82725.0 108715.0 83430.0 110060.0 ;
      RECT  82725.0 111405.0 83430.0 110060.0 ;
      RECT  82725.0 111405.0 83430.0 112750.0 ;
      RECT  82725.0 114095.0 83430.0 112750.0 ;
      RECT  83430.0 28015.0 84135.0 29360.0 ;
      RECT  83430.0 30705.0 84135.0 29360.0 ;
      RECT  83430.0 30705.0 84135.0 32050.0 ;
      RECT  83430.0 33395.0 84135.0 32050.0 ;
      RECT  83430.0 33395.0 84135.0 34740.0 ;
      RECT  83430.0 36085.0 84135.0 34740.0 ;
      RECT  83430.0 36085.0 84135.0 37430.0 ;
      RECT  83430.0 38775.0 84135.0 37430.0 ;
      RECT  83430.0 38775.0 84135.0 40120.0 ;
      RECT  83430.0 41465.0 84135.0 40120.0 ;
      RECT  83430.0 41465.0 84135.0 42810.0 ;
      RECT  83430.0 44155.0 84135.0 42810.0 ;
      RECT  83430.0 44155.0 84135.0 45500.0 ;
      RECT  83430.0 46845.0 84135.0 45500.0 ;
      RECT  83430.0 46845.0 84135.0 48190.0 ;
      RECT  83430.0 49535.0 84135.0 48190.0 ;
      RECT  83430.0 49535.0 84135.0 50880.0 ;
      RECT  83430.0 52225.0 84135.0 50880.0 ;
      RECT  83430.0 52225.0 84135.0 53570.0 ;
      RECT  83430.0 54915.0 84135.0 53570.0 ;
      RECT  83430.0 54915.0 84135.0 56260.0 ;
      RECT  83430.0 57605.0 84135.0 56260.0 ;
      RECT  83430.0 57605.0 84135.0 58950.0 ;
      RECT  83430.0 60295.0 84135.0 58950.0 ;
      RECT  83430.0 60295.0 84135.0 61640.0 ;
      RECT  83430.0 62985.0 84135.0 61640.0 ;
      RECT  83430.0 62985.0 84135.0 64330.0 ;
      RECT  83430.0 65675.0 84135.0 64330.0 ;
      RECT  83430.0 65675.0 84135.0 67020.0 ;
      RECT  83430.0 68365.0 84135.0 67020.0 ;
      RECT  83430.0 68365.0 84135.0 69710.0 ;
      RECT  83430.0 71055.0 84135.0 69710.0 ;
      RECT  83430.0 71055.0 84135.0 72400.0 ;
      RECT  83430.0 73745.0 84135.0 72400.0 ;
      RECT  83430.0 73745.0 84135.0 75090.0 ;
      RECT  83430.0 76435.0 84135.0 75090.0 ;
      RECT  83430.0 76435.0 84135.0 77780.0 ;
      RECT  83430.0 79125.0 84135.0 77780.0 ;
      RECT  83430.0 79125.0 84135.0 80470.0 ;
      RECT  83430.0 81815.0 84135.0 80470.0 ;
      RECT  83430.0 81815.0 84135.0 83160.0 ;
      RECT  83430.0 84505.0 84135.0 83160.0 ;
      RECT  83430.0 84505.0 84135.0 85850.0 ;
      RECT  83430.0 87195.0 84135.0 85850.0 ;
      RECT  83430.0 87195.0 84135.0 88540.0 ;
      RECT  83430.0 89885.0 84135.0 88540.0 ;
      RECT  83430.0 89885.0 84135.0 91230.0 ;
      RECT  83430.0 92575.0 84135.0 91230.0 ;
      RECT  83430.0 92575.0 84135.0 93920.0 ;
      RECT  83430.0 95265.0 84135.0 93920.0 ;
      RECT  83430.0 95265.0 84135.0 96610.0 ;
      RECT  83430.0 97955.0 84135.0 96610.0 ;
      RECT  83430.0 97955.0 84135.0 99300.0 ;
      RECT  83430.0 100645.0 84135.0 99300.0 ;
      RECT  83430.0 100645.0 84135.0 101990.0 ;
      RECT  83430.0 103335.0 84135.0 101990.0 ;
      RECT  83430.0 103335.0 84135.0 104680.0 ;
      RECT  83430.0 106025.0 84135.0 104680.0 ;
      RECT  83430.0 106025.0 84135.0 107370.0 ;
      RECT  83430.0 108715.0 84135.0 107370.0 ;
      RECT  83430.0 108715.0 84135.0 110060.0 ;
      RECT  83430.0 111405.0 84135.0 110060.0 ;
      RECT  83430.0 111405.0 84135.0 112750.0 ;
      RECT  83430.0 114095.0 84135.0 112750.0 ;
      RECT  84135.0 28015.0 84840.0 29360.0 ;
      RECT  84135.0 30705.0 84840.0 29360.0 ;
      RECT  84135.0 30705.0 84840.0 32050.0 ;
      RECT  84135.0 33395.0 84840.0 32050.0 ;
      RECT  84135.0 33395.0 84840.0 34740.0 ;
      RECT  84135.0 36085.0 84840.0 34740.0 ;
      RECT  84135.0 36085.0 84840.0 37430.0 ;
      RECT  84135.0 38775.0 84840.0 37430.0 ;
      RECT  84135.0 38775.0 84840.0 40120.0 ;
      RECT  84135.0 41465.0 84840.0 40120.0 ;
      RECT  84135.0 41465.0 84840.0 42810.0 ;
      RECT  84135.0 44155.0 84840.0 42810.0 ;
      RECT  84135.0 44155.0 84840.0 45500.0 ;
      RECT  84135.0 46845.0 84840.0 45500.0 ;
      RECT  84135.0 46845.0 84840.0 48190.0 ;
      RECT  84135.0 49535.0 84840.0 48190.0 ;
      RECT  84135.0 49535.0 84840.0 50880.0 ;
      RECT  84135.0 52225.0 84840.0 50880.0 ;
      RECT  84135.0 52225.0 84840.0 53570.0 ;
      RECT  84135.0 54915.0 84840.0 53570.0 ;
      RECT  84135.0 54915.0 84840.0 56260.0 ;
      RECT  84135.0 57605.0 84840.0 56260.0 ;
      RECT  84135.0 57605.0 84840.0 58950.0 ;
      RECT  84135.0 60295.0 84840.0 58950.0 ;
      RECT  84135.0 60295.0 84840.0 61640.0 ;
      RECT  84135.0 62985.0 84840.0 61640.0 ;
      RECT  84135.0 62985.0 84840.0 64330.0 ;
      RECT  84135.0 65675.0 84840.0 64330.0 ;
      RECT  84135.0 65675.0 84840.0 67020.0 ;
      RECT  84135.0 68365.0 84840.0 67020.0 ;
      RECT  84135.0 68365.0 84840.0 69710.0 ;
      RECT  84135.0 71055.0 84840.0 69710.0 ;
      RECT  84135.0 71055.0 84840.0 72400.0 ;
      RECT  84135.0 73745.0 84840.0 72400.0 ;
      RECT  84135.0 73745.0 84840.0 75090.0 ;
      RECT  84135.0 76435.0 84840.0 75090.0 ;
      RECT  84135.0 76435.0 84840.0 77780.0 ;
      RECT  84135.0 79125.0 84840.0 77780.0 ;
      RECT  84135.0 79125.0 84840.0 80470.0 ;
      RECT  84135.0 81815.0 84840.0 80470.0 ;
      RECT  84135.0 81815.0 84840.0 83160.0 ;
      RECT  84135.0 84505.0 84840.0 83160.0 ;
      RECT  84135.0 84505.0 84840.0 85850.0 ;
      RECT  84135.0 87195.0 84840.0 85850.0 ;
      RECT  84135.0 87195.0 84840.0 88540.0 ;
      RECT  84135.0 89885.0 84840.0 88540.0 ;
      RECT  84135.0 89885.0 84840.0 91230.0 ;
      RECT  84135.0 92575.0 84840.0 91230.0 ;
      RECT  84135.0 92575.0 84840.0 93920.0 ;
      RECT  84135.0 95265.0 84840.0 93920.0 ;
      RECT  84135.0 95265.0 84840.0 96610.0 ;
      RECT  84135.0 97955.0 84840.0 96610.0 ;
      RECT  84135.0 97955.0 84840.0 99300.0 ;
      RECT  84135.0 100645.0 84840.0 99300.0 ;
      RECT  84135.0 100645.0 84840.0 101990.0 ;
      RECT  84135.0 103335.0 84840.0 101990.0 ;
      RECT  84135.0 103335.0 84840.0 104680.0 ;
      RECT  84135.0 106025.0 84840.0 104680.0 ;
      RECT  84135.0 106025.0 84840.0 107370.0 ;
      RECT  84135.0 108715.0 84840.0 107370.0 ;
      RECT  84135.0 108715.0 84840.0 110060.0 ;
      RECT  84135.0 111405.0 84840.0 110060.0 ;
      RECT  84135.0 111405.0 84840.0 112750.0 ;
      RECT  84135.0 114095.0 84840.0 112750.0 ;
      RECT  84840.0 28015.0 85545.0 29360.0 ;
      RECT  84840.0 30705.0 85545.0 29360.0 ;
      RECT  84840.0 30705.0 85545.0 32050.0 ;
      RECT  84840.0 33395.0 85545.0 32050.0 ;
      RECT  84840.0 33395.0 85545.0 34740.0 ;
      RECT  84840.0 36085.0 85545.0 34740.0 ;
      RECT  84840.0 36085.0 85545.0 37430.0 ;
      RECT  84840.0 38775.0 85545.0 37430.0 ;
      RECT  84840.0 38775.0 85545.0 40120.0 ;
      RECT  84840.0 41465.0 85545.0 40120.0 ;
      RECT  84840.0 41465.0 85545.0 42810.0 ;
      RECT  84840.0 44155.0 85545.0 42810.0 ;
      RECT  84840.0 44155.0 85545.0 45500.0 ;
      RECT  84840.0 46845.0 85545.0 45500.0 ;
      RECT  84840.0 46845.0 85545.0 48190.0 ;
      RECT  84840.0 49535.0 85545.0 48190.0 ;
      RECT  84840.0 49535.0 85545.0 50880.0 ;
      RECT  84840.0 52225.0 85545.0 50880.0 ;
      RECT  84840.0 52225.0 85545.0 53570.0 ;
      RECT  84840.0 54915.0 85545.0 53570.0 ;
      RECT  84840.0 54915.0 85545.0 56260.0 ;
      RECT  84840.0 57605.0 85545.0 56260.0 ;
      RECT  84840.0 57605.0 85545.0 58950.0 ;
      RECT  84840.0 60295.0 85545.0 58950.0 ;
      RECT  84840.0 60295.0 85545.0 61640.0 ;
      RECT  84840.0 62985.0 85545.0 61640.0 ;
      RECT  84840.0 62985.0 85545.0 64330.0 ;
      RECT  84840.0 65675.0 85545.0 64330.0 ;
      RECT  84840.0 65675.0 85545.0 67020.0 ;
      RECT  84840.0 68365.0 85545.0 67020.0 ;
      RECT  84840.0 68365.0 85545.0 69710.0 ;
      RECT  84840.0 71055.0 85545.0 69710.0 ;
      RECT  84840.0 71055.0 85545.0 72400.0 ;
      RECT  84840.0 73745.0 85545.0 72400.0 ;
      RECT  84840.0 73745.0 85545.0 75090.0 ;
      RECT  84840.0 76435.0 85545.0 75090.0 ;
      RECT  84840.0 76435.0 85545.0 77780.0 ;
      RECT  84840.0 79125.0 85545.0 77780.0 ;
      RECT  84840.0 79125.0 85545.0 80470.0 ;
      RECT  84840.0 81815.0 85545.0 80470.0 ;
      RECT  84840.0 81815.0 85545.0 83160.0 ;
      RECT  84840.0 84505.0 85545.0 83160.0 ;
      RECT  84840.0 84505.0 85545.0 85850.0 ;
      RECT  84840.0 87195.0 85545.0 85850.0 ;
      RECT  84840.0 87195.0 85545.0 88540.0 ;
      RECT  84840.0 89885.0 85545.0 88540.0 ;
      RECT  84840.0 89885.0 85545.0 91230.0 ;
      RECT  84840.0 92575.0 85545.0 91230.0 ;
      RECT  84840.0 92575.0 85545.0 93920.0 ;
      RECT  84840.0 95265.0 85545.0 93920.0 ;
      RECT  84840.0 95265.0 85545.0 96610.0 ;
      RECT  84840.0 97955.0 85545.0 96610.0 ;
      RECT  84840.0 97955.0 85545.0 99300.0 ;
      RECT  84840.0 100645.0 85545.0 99300.0 ;
      RECT  84840.0 100645.0 85545.0 101990.0 ;
      RECT  84840.0 103335.0 85545.0 101990.0 ;
      RECT  84840.0 103335.0 85545.0 104680.0 ;
      RECT  84840.0 106025.0 85545.0 104680.0 ;
      RECT  84840.0 106025.0 85545.0 107370.0 ;
      RECT  84840.0 108715.0 85545.0 107370.0 ;
      RECT  84840.0 108715.0 85545.0 110060.0 ;
      RECT  84840.0 111405.0 85545.0 110060.0 ;
      RECT  84840.0 111405.0 85545.0 112750.0 ;
      RECT  84840.0 114095.0 85545.0 112750.0 ;
      RECT  85545.0 28015.0 86250.0 29360.0 ;
      RECT  85545.0 30705.0 86250.0 29360.0 ;
      RECT  85545.0 30705.0 86250.0 32050.0 ;
      RECT  85545.0 33395.0 86250.0 32050.0 ;
      RECT  85545.0 33395.0 86250.0 34740.0 ;
      RECT  85545.0 36085.0 86250.0 34740.0 ;
      RECT  85545.0 36085.0 86250.0 37430.0 ;
      RECT  85545.0 38775.0 86250.0 37430.0 ;
      RECT  85545.0 38775.0 86250.0 40120.0 ;
      RECT  85545.0 41465.0 86250.0 40120.0 ;
      RECT  85545.0 41465.0 86250.0 42810.0 ;
      RECT  85545.0 44155.0 86250.0 42810.0 ;
      RECT  85545.0 44155.0 86250.0 45500.0 ;
      RECT  85545.0 46845.0 86250.0 45500.0 ;
      RECT  85545.0 46845.0 86250.0 48190.0 ;
      RECT  85545.0 49535.0 86250.0 48190.0 ;
      RECT  85545.0 49535.0 86250.0 50880.0 ;
      RECT  85545.0 52225.0 86250.0 50880.0 ;
      RECT  85545.0 52225.0 86250.0 53570.0 ;
      RECT  85545.0 54915.0 86250.0 53570.0 ;
      RECT  85545.0 54915.0 86250.0 56260.0 ;
      RECT  85545.0 57605.0 86250.0 56260.0 ;
      RECT  85545.0 57605.0 86250.0 58950.0 ;
      RECT  85545.0 60295.0 86250.0 58950.0 ;
      RECT  85545.0 60295.0 86250.0 61640.0 ;
      RECT  85545.0 62985.0 86250.0 61640.0 ;
      RECT  85545.0 62985.0 86250.0 64330.0 ;
      RECT  85545.0 65675.0 86250.0 64330.0 ;
      RECT  85545.0 65675.0 86250.0 67020.0 ;
      RECT  85545.0 68365.0 86250.0 67020.0 ;
      RECT  85545.0 68365.0 86250.0 69710.0 ;
      RECT  85545.0 71055.0 86250.0 69710.0 ;
      RECT  85545.0 71055.0 86250.0 72400.0 ;
      RECT  85545.0 73745.0 86250.0 72400.0 ;
      RECT  85545.0 73745.0 86250.0 75090.0 ;
      RECT  85545.0 76435.0 86250.0 75090.0 ;
      RECT  85545.0 76435.0 86250.0 77780.0 ;
      RECT  85545.0 79125.0 86250.0 77780.0 ;
      RECT  85545.0 79125.0 86250.0 80470.0 ;
      RECT  85545.0 81815.0 86250.0 80470.0 ;
      RECT  85545.0 81815.0 86250.0 83160.0 ;
      RECT  85545.0 84505.0 86250.0 83160.0 ;
      RECT  85545.0 84505.0 86250.0 85850.0 ;
      RECT  85545.0 87195.0 86250.0 85850.0 ;
      RECT  85545.0 87195.0 86250.0 88540.0 ;
      RECT  85545.0 89885.0 86250.0 88540.0 ;
      RECT  85545.0 89885.0 86250.0 91230.0 ;
      RECT  85545.0 92575.0 86250.0 91230.0 ;
      RECT  85545.0 92575.0 86250.0 93920.0 ;
      RECT  85545.0 95265.0 86250.0 93920.0 ;
      RECT  85545.0 95265.0 86250.0 96610.0 ;
      RECT  85545.0 97955.0 86250.0 96610.0 ;
      RECT  85545.0 97955.0 86250.0 99300.0 ;
      RECT  85545.0 100645.0 86250.0 99300.0 ;
      RECT  85545.0 100645.0 86250.0 101990.0 ;
      RECT  85545.0 103335.0 86250.0 101990.0 ;
      RECT  85545.0 103335.0 86250.0 104680.0 ;
      RECT  85545.0 106025.0 86250.0 104680.0 ;
      RECT  85545.0 106025.0 86250.0 107370.0 ;
      RECT  85545.0 108715.0 86250.0 107370.0 ;
      RECT  85545.0 108715.0 86250.0 110060.0 ;
      RECT  85545.0 111405.0 86250.0 110060.0 ;
      RECT  85545.0 111405.0 86250.0 112750.0 ;
      RECT  85545.0 114095.0 86250.0 112750.0 ;
      RECT  86250.0 28015.0 86955.0 29360.0 ;
      RECT  86250.0 30705.0 86955.0 29360.0 ;
      RECT  86250.0 30705.0 86955.0 32050.0 ;
      RECT  86250.0 33395.0 86955.0 32050.0 ;
      RECT  86250.0 33395.0 86955.0 34740.0 ;
      RECT  86250.0 36085.0 86955.0 34740.0 ;
      RECT  86250.0 36085.0 86955.0 37430.0 ;
      RECT  86250.0 38775.0 86955.0 37430.0 ;
      RECT  86250.0 38775.0 86955.0 40120.0 ;
      RECT  86250.0 41465.0 86955.0 40120.0 ;
      RECT  86250.0 41465.0 86955.0 42810.0 ;
      RECT  86250.0 44155.0 86955.0 42810.0 ;
      RECT  86250.0 44155.0 86955.0 45500.0 ;
      RECT  86250.0 46845.0 86955.0 45500.0 ;
      RECT  86250.0 46845.0 86955.0 48190.0 ;
      RECT  86250.0 49535.0 86955.0 48190.0 ;
      RECT  86250.0 49535.0 86955.0 50880.0 ;
      RECT  86250.0 52225.0 86955.0 50880.0 ;
      RECT  86250.0 52225.0 86955.0 53570.0 ;
      RECT  86250.0 54915.0 86955.0 53570.0 ;
      RECT  86250.0 54915.0 86955.0 56260.0 ;
      RECT  86250.0 57605.0 86955.0 56260.0 ;
      RECT  86250.0 57605.0 86955.0 58950.0 ;
      RECT  86250.0 60295.0 86955.0 58950.0 ;
      RECT  86250.0 60295.0 86955.0 61640.0 ;
      RECT  86250.0 62985.0 86955.0 61640.0 ;
      RECT  86250.0 62985.0 86955.0 64330.0 ;
      RECT  86250.0 65675.0 86955.0 64330.0 ;
      RECT  86250.0 65675.0 86955.0 67020.0 ;
      RECT  86250.0 68365.0 86955.0 67020.0 ;
      RECT  86250.0 68365.0 86955.0 69710.0 ;
      RECT  86250.0 71055.0 86955.0 69710.0 ;
      RECT  86250.0 71055.0 86955.0 72400.0 ;
      RECT  86250.0 73745.0 86955.0 72400.0 ;
      RECT  86250.0 73745.0 86955.0 75090.0 ;
      RECT  86250.0 76435.0 86955.0 75090.0 ;
      RECT  86250.0 76435.0 86955.0 77780.0 ;
      RECT  86250.0 79125.0 86955.0 77780.0 ;
      RECT  86250.0 79125.0 86955.0 80470.0 ;
      RECT  86250.0 81815.0 86955.0 80470.0 ;
      RECT  86250.0 81815.0 86955.0 83160.0 ;
      RECT  86250.0 84505.0 86955.0 83160.0 ;
      RECT  86250.0 84505.0 86955.0 85850.0 ;
      RECT  86250.0 87195.0 86955.0 85850.0 ;
      RECT  86250.0 87195.0 86955.0 88540.0 ;
      RECT  86250.0 89885.0 86955.0 88540.0 ;
      RECT  86250.0 89885.0 86955.0 91230.0 ;
      RECT  86250.0 92575.0 86955.0 91230.0 ;
      RECT  86250.0 92575.0 86955.0 93920.0 ;
      RECT  86250.0 95265.0 86955.0 93920.0 ;
      RECT  86250.0 95265.0 86955.0 96610.0 ;
      RECT  86250.0 97955.0 86955.0 96610.0 ;
      RECT  86250.0 97955.0 86955.0 99300.0 ;
      RECT  86250.0 100645.0 86955.0 99300.0 ;
      RECT  86250.0 100645.0 86955.0 101990.0 ;
      RECT  86250.0 103335.0 86955.0 101990.0 ;
      RECT  86250.0 103335.0 86955.0 104680.0 ;
      RECT  86250.0 106025.0 86955.0 104680.0 ;
      RECT  86250.0 106025.0 86955.0 107370.0 ;
      RECT  86250.0 108715.0 86955.0 107370.0 ;
      RECT  86250.0 108715.0 86955.0 110060.0 ;
      RECT  86250.0 111405.0 86955.0 110060.0 ;
      RECT  86250.0 111405.0 86955.0 112750.0 ;
      RECT  86250.0 114095.0 86955.0 112750.0 ;
      RECT  86955.0 28015.0 87660.0 29360.0 ;
      RECT  86955.0 30705.0 87660.0 29360.0 ;
      RECT  86955.0 30705.0 87660.0 32050.0 ;
      RECT  86955.0 33395.0 87660.0 32050.0 ;
      RECT  86955.0 33395.0 87660.0 34740.0 ;
      RECT  86955.0 36085.0 87660.0 34740.0 ;
      RECT  86955.0 36085.0 87660.0 37430.0 ;
      RECT  86955.0 38775.0 87660.0 37430.0 ;
      RECT  86955.0 38775.0 87660.0 40120.0 ;
      RECT  86955.0 41465.0 87660.0 40120.0 ;
      RECT  86955.0 41465.0 87660.0 42810.0 ;
      RECT  86955.0 44155.0 87660.0 42810.0 ;
      RECT  86955.0 44155.0 87660.0 45500.0 ;
      RECT  86955.0 46845.0 87660.0 45500.0 ;
      RECT  86955.0 46845.0 87660.0 48190.0 ;
      RECT  86955.0 49535.0 87660.0 48190.0 ;
      RECT  86955.0 49535.0 87660.0 50880.0 ;
      RECT  86955.0 52225.0 87660.0 50880.0 ;
      RECT  86955.0 52225.0 87660.0 53570.0 ;
      RECT  86955.0 54915.0 87660.0 53570.0 ;
      RECT  86955.0 54915.0 87660.0 56260.0 ;
      RECT  86955.0 57605.0 87660.0 56260.0 ;
      RECT  86955.0 57605.0 87660.0 58950.0 ;
      RECT  86955.0 60295.0 87660.0 58950.0 ;
      RECT  86955.0 60295.0 87660.0 61640.0 ;
      RECT  86955.0 62985.0 87660.0 61640.0 ;
      RECT  86955.0 62985.0 87660.0 64330.0 ;
      RECT  86955.0 65675.0 87660.0 64330.0 ;
      RECT  86955.0 65675.0 87660.0 67020.0 ;
      RECT  86955.0 68365.0 87660.0 67020.0 ;
      RECT  86955.0 68365.0 87660.0 69710.0 ;
      RECT  86955.0 71055.0 87660.0 69710.0 ;
      RECT  86955.0 71055.0 87660.0 72400.0 ;
      RECT  86955.0 73745.0 87660.0 72400.0 ;
      RECT  86955.0 73745.0 87660.0 75090.0 ;
      RECT  86955.0 76435.0 87660.0 75090.0 ;
      RECT  86955.0 76435.0 87660.0 77780.0 ;
      RECT  86955.0 79125.0 87660.0 77780.0 ;
      RECT  86955.0 79125.0 87660.0 80470.0 ;
      RECT  86955.0 81815.0 87660.0 80470.0 ;
      RECT  86955.0 81815.0 87660.0 83160.0 ;
      RECT  86955.0 84505.0 87660.0 83160.0 ;
      RECT  86955.0 84505.0 87660.0 85850.0 ;
      RECT  86955.0 87195.0 87660.0 85850.0 ;
      RECT  86955.0 87195.0 87660.0 88540.0 ;
      RECT  86955.0 89885.0 87660.0 88540.0 ;
      RECT  86955.0 89885.0 87660.0 91230.0 ;
      RECT  86955.0 92575.0 87660.0 91230.0 ;
      RECT  86955.0 92575.0 87660.0 93920.0 ;
      RECT  86955.0 95265.0 87660.0 93920.0 ;
      RECT  86955.0 95265.0 87660.0 96610.0 ;
      RECT  86955.0 97955.0 87660.0 96610.0 ;
      RECT  86955.0 97955.0 87660.0 99300.0 ;
      RECT  86955.0 100645.0 87660.0 99300.0 ;
      RECT  86955.0 100645.0 87660.0 101990.0 ;
      RECT  86955.0 103335.0 87660.0 101990.0 ;
      RECT  86955.0 103335.0 87660.0 104680.0 ;
      RECT  86955.0 106025.0 87660.0 104680.0 ;
      RECT  86955.0 106025.0 87660.0 107370.0 ;
      RECT  86955.0 108715.0 87660.0 107370.0 ;
      RECT  86955.0 108715.0 87660.0 110060.0 ;
      RECT  86955.0 111405.0 87660.0 110060.0 ;
      RECT  86955.0 111405.0 87660.0 112750.0 ;
      RECT  86955.0 114095.0 87660.0 112750.0 ;
      RECT  87660.0 28015.0 88365.0 29360.0 ;
      RECT  87660.0 30705.0 88365.0 29360.0 ;
      RECT  87660.0 30705.0 88365.0 32050.0 ;
      RECT  87660.0 33395.0 88365.0 32050.0 ;
      RECT  87660.0 33395.0 88365.0 34740.0 ;
      RECT  87660.0 36085.0 88365.0 34740.0 ;
      RECT  87660.0 36085.0 88365.0 37430.0 ;
      RECT  87660.0 38775.0 88365.0 37430.0 ;
      RECT  87660.0 38775.0 88365.0 40120.0 ;
      RECT  87660.0 41465.0 88365.0 40120.0 ;
      RECT  87660.0 41465.0 88365.0 42810.0 ;
      RECT  87660.0 44155.0 88365.0 42810.0 ;
      RECT  87660.0 44155.0 88365.0 45500.0 ;
      RECT  87660.0 46845.0 88365.0 45500.0 ;
      RECT  87660.0 46845.0 88365.0 48190.0 ;
      RECT  87660.0 49535.0 88365.0 48190.0 ;
      RECT  87660.0 49535.0 88365.0 50880.0 ;
      RECT  87660.0 52225.0 88365.0 50880.0 ;
      RECT  87660.0 52225.0 88365.0 53570.0 ;
      RECT  87660.0 54915.0 88365.0 53570.0 ;
      RECT  87660.0 54915.0 88365.0 56260.0 ;
      RECT  87660.0 57605.0 88365.0 56260.0 ;
      RECT  87660.0 57605.0 88365.0 58950.0 ;
      RECT  87660.0 60295.0 88365.0 58950.0 ;
      RECT  87660.0 60295.0 88365.0 61640.0 ;
      RECT  87660.0 62985.0 88365.0 61640.0 ;
      RECT  87660.0 62985.0 88365.0 64330.0 ;
      RECT  87660.0 65675.0 88365.0 64330.0 ;
      RECT  87660.0 65675.0 88365.0 67020.0 ;
      RECT  87660.0 68365.0 88365.0 67020.0 ;
      RECT  87660.0 68365.0 88365.0 69710.0 ;
      RECT  87660.0 71055.0 88365.0 69710.0 ;
      RECT  87660.0 71055.0 88365.0 72400.0 ;
      RECT  87660.0 73745.0 88365.0 72400.0 ;
      RECT  87660.0 73745.0 88365.0 75090.0 ;
      RECT  87660.0 76435.0 88365.0 75090.0 ;
      RECT  87660.0 76435.0 88365.0 77780.0 ;
      RECT  87660.0 79125.0 88365.0 77780.0 ;
      RECT  87660.0 79125.0 88365.0 80470.0 ;
      RECT  87660.0 81815.0 88365.0 80470.0 ;
      RECT  87660.0 81815.0 88365.0 83160.0 ;
      RECT  87660.0 84505.0 88365.0 83160.0 ;
      RECT  87660.0 84505.0 88365.0 85850.0 ;
      RECT  87660.0 87195.0 88365.0 85850.0 ;
      RECT  87660.0 87195.0 88365.0 88540.0 ;
      RECT  87660.0 89885.0 88365.0 88540.0 ;
      RECT  87660.0 89885.0 88365.0 91230.0 ;
      RECT  87660.0 92575.0 88365.0 91230.0 ;
      RECT  87660.0 92575.0 88365.0 93920.0 ;
      RECT  87660.0 95265.0 88365.0 93920.0 ;
      RECT  87660.0 95265.0 88365.0 96610.0 ;
      RECT  87660.0 97955.0 88365.0 96610.0 ;
      RECT  87660.0 97955.0 88365.0 99300.0 ;
      RECT  87660.0 100645.0 88365.0 99300.0 ;
      RECT  87660.0 100645.0 88365.0 101990.0 ;
      RECT  87660.0 103335.0 88365.0 101990.0 ;
      RECT  87660.0 103335.0 88365.0 104680.0 ;
      RECT  87660.0 106025.0 88365.0 104680.0 ;
      RECT  87660.0 106025.0 88365.0 107370.0 ;
      RECT  87660.0 108715.0 88365.0 107370.0 ;
      RECT  87660.0 108715.0 88365.0 110060.0 ;
      RECT  87660.0 111405.0 88365.0 110060.0 ;
      RECT  87660.0 111405.0 88365.0 112750.0 ;
      RECT  87660.0 114095.0 88365.0 112750.0 ;
      RECT  88365.0 28015.0 89070.0 29360.0 ;
      RECT  88365.0 30705.0 89070.0 29360.0 ;
      RECT  88365.0 30705.0 89070.0 32050.0 ;
      RECT  88365.0 33395.0 89070.0 32050.0 ;
      RECT  88365.0 33395.0 89070.0 34740.0 ;
      RECT  88365.0 36085.0 89070.0 34740.0 ;
      RECT  88365.0 36085.0 89070.0 37430.0 ;
      RECT  88365.0 38775.0 89070.0 37430.0 ;
      RECT  88365.0 38775.0 89070.0 40120.0 ;
      RECT  88365.0 41465.0 89070.0 40120.0 ;
      RECT  88365.0 41465.0 89070.0 42810.0 ;
      RECT  88365.0 44155.0 89070.0 42810.0 ;
      RECT  88365.0 44155.0 89070.0 45500.0 ;
      RECT  88365.0 46845.0 89070.0 45500.0 ;
      RECT  88365.0 46845.0 89070.0 48190.0 ;
      RECT  88365.0 49535.0 89070.0 48190.0 ;
      RECT  88365.0 49535.0 89070.0 50880.0 ;
      RECT  88365.0 52225.0 89070.0 50880.0 ;
      RECT  88365.0 52225.0 89070.0 53570.0 ;
      RECT  88365.0 54915.0 89070.0 53570.0 ;
      RECT  88365.0 54915.0 89070.0 56260.0 ;
      RECT  88365.0 57605.0 89070.0 56260.0 ;
      RECT  88365.0 57605.0 89070.0 58950.0 ;
      RECT  88365.0 60295.0 89070.0 58950.0 ;
      RECT  88365.0 60295.0 89070.0 61640.0 ;
      RECT  88365.0 62985.0 89070.0 61640.0 ;
      RECT  88365.0 62985.0 89070.0 64330.0 ;
      RECT  88365.0 65675.0 89070.0 64330.0 ;
      RECT  88365.0 65675.0 89070.0 67020.0 ;
      RECT  88365.0 68365.0 89070.0 67020.0 ;
      RECT  88365.0 68365.0 89070.0 69710.0 ;
      RECT  88365.0 71055.0 89070.0 69710.0 ;
      RECT  88365.0 71055.0 89070.0 72400.0 ;
      RECT  88365.0 73745.0 89070.0 72400.0 ;
      RECT  88365.0 73745.0 89070.0 75090.0 ;
      RECT  88365.0 76435.0 89070.0 75090.0 ;
      RECT  88365.0 76435.0 89070.0 77780.0 ;
      RECT  88365.0 79125.0 89070.0 77780.0 ;
      RECT  88365.0 79125.0 89070.0 80470.0 ;
      RECT  88365.0 81815.0 89070.0 80470.0 ;
      RECT  88365.0 81815.0 89070.0 83160.0 ;
      RECT  88365.0 84505.0 89070.0 83160.0 ;
      RECT  88365.0 84505.0 89070.0 85850.0 ;
      RECT  88365.0 87195.0 89070.0 85850.0 ;
      RECT  88365.0 87195.0 89070.0 88540.0 ;
      RECT  88365.0 89885.0 89070.0 88540.0 ;
      RECT  88365.0 89885.0 89070.0 91230.0 ;
      RECT  88365.0 92575.0 89070.0 91230.0 ;
      RECT  88365.0 92575.0 89070.0 93920.0 ;
      RECT  88365.0 95265.0 89070.0 93920.0 ;
      RECT  88365.0 95265.0 89070.0 96610.0 ;
      RECT  88365.0 97955.0 89070.0 96610.0 ;
      RECT  88365.0 97955.0 89070.0 99300.0 ;
      RECT  88365.0 100645.0 89070.0 99300.0 ;
      RECT  88365.0 100645.0 89070.0 101990.0 ;
      RECT  88365.0 103335.0 89070.0 101990.0 ;
      RECT  88365.0 103335.0 89070.0 104680.0 ;
      RECT  88365.0 106025.0 89070.0 104680.0 ;
      RECT  88365.0 106025.0 89070.0 107370.0 ;
      RECT  88365.0 108715.0 89070.0 107370.0 ;
      RECT  88365.0 108715.0 89070.0 110060.0 ;
      RECT  88365.0 111405.0 89070.0 110060.0 ;
      RECT  88365.0 111405.0 89070.0 112750.0 ;
      RECT  88365.0 114095.0 89070.0 112750.0 ;
      RECT  89070.0 28015.0 89775.0 29360.0 ;
      RECT  89070.0 30705.0 89775.0 29360.0 ;
      RECT  89070.0 30705.0 89775.0 32050.0 ;
      RECT  89070.0 33395.0 89775.0 32050.0 ;
      RECT  89070.0 33395.0 89775.0 34740.0 ;
      RECT  89070.0 36085.0 89775.0 34740.0 ;
      RECT  89070.0 36085.0 89775.0 37430.0 ;
      RECT  89070.0 38775.0 89775.0 37430.0 ;
      RECT  89070.0 38775.0 89775.0 40120.0 ;
      RECT  89070.0 41465.0 89775.0 40120.0 ;
      RECT  89070.0 41465.0 89775.0 42810.0 ;
      RECT  89070.0 44155.0 89775.0 42810.0 ;
      RECT  89070.0 44155.0 89775.0 45500.0 ;
      RECT  89070.0 46845.0 89775.0 45500.0 ;
      RECT  89070.0 46845.0 89775.0 48190.0 ;
      RECT  89070.0 49535.0 89775.0 48190.0 ;
      RECT  89070.0 49535.0 89775.0 50880.0 ;
      RECT  89070.0 52225.0 89775.0 50880.0 ;
      RECT  89070.0 52225.0 89775.0 53570.0 ;
      RECT  89070.0 54915.0 89775.0 53570.0 ;
      RECT  89070.0 54915.0 89775.0 56260.0 ;
      RECT  89070.0 57605.0 89775.0 56260.0 ;
      RECT  89070.0 57605.0 89775.0 58950.0 ;
      RECT  89070.0 60295.0 89775.0 58950.0 ;
      RECT  89070.0 60295.0 89775.0 61640.0 ;
      RECT  89070.0 62985.0 89775.0 61640.0 ;
      RECT  89070.0 62985.0 89775.0 64330.0 ;
      RECT  89070.0 65675.0 89775.0 64330.0 ;
      RECT  89070.0 65675.0 89775.0 67020.0 ;
      RECT  89070.0 68365.0 89775.0 67020.0 ;
      RECT  89070.0 68365.0 89775.0 69710.0 ;
      RECT  89070.0 71055.0 89775.0 69710.0 ;
      RECT  89070.0 71055.0 89775.0 72400.0 ;
      RECT  89070.0 73745.0 89775.0 72400.0 ;
      RECT  89070.0 73745.0 89775.0 75090.0 ;
      RECT  89070.0 76435.0 89775.0 75090.0 ;
      RECT  89070.0 76435.0 89775.0 77780.0 ;
      RECT  89070.0 79125.0 89775.0 77780.0 ;
      RECT  89070.0 79125.0 89775.0 80470.0 ;
      RECT  89070.0 81815.0 89775.0 80470.0 ;
      RECT  89070.0 81815.0 89775.0 83160.0 ;
      RECT  89070.0 84505.0 89775.0 83160.0 ;
      RECT  89070.0 84505.0 89775.0 85850.0 ;
      RECT  89070.0 87195.0 89775.0 85850.0 ;
      RECT  89070.0 87195.0 89775.0 88540.0 ;
      RECT  89070.0 89885.0 89775.0 88540.0 ;
      RECT  89070.0 89885.0 89775.0 91230.0 ;
      RECT  89070.0 92575.0 89775.0 91230.0 ;
      RECT  89070.0 92575.0 89775.0 93920.0 ;
      RECT  89070.0 95265.0 89775.0 93920.0 ;
      RECT  89070.0 95265.0 89775.0 96610.0 ;
      RECT  89070.0 97955.0 89775.0 96610.0 ;
      RECT  89070.0 97955.0 89775.0 99300.0 ;
      RECT  89070.0 100645.0 89775.0 99300.0 ;
      RECT  89070.0 100645.0 89775.0 101990.0 ;
      RECT  89070.0 103335.0 89775.0 101990.0 ;
      RECT  89070.0 103335.0 89775.0 104680.0 ;
      RECT  89070.0 106025.0 89775.0 104680.0 ;
      RECT  89070.0 106025.0 89775.0 107370.0 ;
      RECT  89070.0 108715.0 89775.0 107370.0 ;
      RECT  89070.0 108715.0 89775.0 110060.0 ;
      RECT  89070.0 111405.0 89775.0 110060.0 ;
      RECT  89070.0 111405.0 89775.0 112750.0 ;
      RECT  89070.0 114095.0 89775.0 112750.0 ;
      RECT  89775.0 28015.0 90480.0 29360.0 ;
      RECT  89775.0 30705.0 90480.0 29360.0 ;
      RECT  89775.0 30705.0 90480.0 32050.0 ;
      RECT  89775.0 33395.0 90480.0 32050.0 ;
      RECT  89775.0 33395.0 90480.0 34740.0 ;
      RECT  89775.0 36085.0 90480.0 34740.0 ;
      RECT  89775.0 36085.0 90480.0 37430.0 ;
      RECT  89775.0 38775.0 90480.0 37430.0 ;
      RECT  89775.0 38775.0 90480.0 40120.0 ;
      RECT  89775.0 41465.0 90480.0 40120.0 ;
      RECT  89775.0 41465.0 90480.0 42810.0 ;
      RECT  89775.0 44155.0 90480.0 42810.0 ;
      RECT  89775.0 44155.0 90480.0 45500.0 ;
      RECT  89775.0 46845.0 90480.0 45500.0 ;
      RECT  89775.0 46845.0 90480.0 48190.0 ;
      RECT  89775.0 49535.0 90480.0 48190.0 ;
      RECT  89775.0 49535.0 90480.0 50880.0 ;
      RECT  89775.0 52225.0 90480.0 50880.0 ;
      RECT  89775.0 52225.0 90480.0 53570.0 ;
      RECT  89775.0 54915.0 90480.0 53570.0 ;
      RECT  89775.0 54915.0 90480.0 56260.0 ;
      RECT  89775.0 57605.0 90480.0 56260.0 ;
      RECT  89775.0 57605.0 90480.0 58950.0 ;
      RECT  89775.0 60295.0 90480.0 58950.0 ;
      RECT  89775.0 60295.0 90480.0 61640.0 ;
      RECT  89775.0 62985.0 90480.0 61640.0 ;
      RECT  89775.0 62985.0 90480.0 64330.0 ;
      RECT  89775.0 65675.0 90480.0 64330.0 ;
      RECT  89775.0 65675.0 90480.0 67020.0 ;
      RECT  89775.0 68365.0 90480.0 67020.0 ;
      RECT  89775.0 68365.0 90480.0 69710.0 ;
      RECT  89775.0 71055.0 90480.0 69710.0 ;
      RECT  89775.0 71055.0 90480.0 72400.0 ;
      RECT  89775.0 73745.0 90480.0 72400.0 ;
      RECT  89775.0 73745.0 90480.0 75090.0 ;
      RECT  89775.0 76435.0 90480.0 75090.0 ;
      RECT  89775.0 76435.0 90480.0 77780.0 ;
      RECT  89775.0 79125.0 90480.0 77780.0 ;
      RECT  89775.0 79125.0 90480.0 80470.0 ;
      RECT  89775.0 81815.0 90480.0 80470.0 ;
      RECT  89775.0 81815.0 90480.0 83160.0 ;
      RECT  89775.0 84505.0 90480.0 83160.0 ;
      RECT  89775.0 84505.0 90480.0 85850.0 ;
      RECT  89775.0 87195.0 90480.0 85850.0 ;
      RECT  89775.0 87195.0 90480.0 88540.0 ;
      RECT  89775.0 89885.0 90480.0 88540.0 ;
      RECT  89775.0 89885.0 90480.0 91230.0 ;
      RECT  89775.0 92575.0 90480.0 91230.0 ;
      RECT  89775.0 92575.0 90480.0 93920.0 ;
      RECT  89775.0 95265.0 90480.0 93920.0 ;
      RECT  89775.0 95265.0 90480.0 96610.0 ;
      RECT  89775.0 97955.0 90480.0 96610.0 ;
      RECT  89775.0 97955.0 90480.0 99300.0 ;
      RECT  89775.0 100645.0 90480.0 99300.0 ;
      RECT  89775.0 100645.0 90480.0 101990.0 ;
      RECT  89775.0 103335.0 90480.0 101990.0 ;
      RECT  89775.0 103335.0 90480.0 104680.0 ;
      RECT  89775.0 106025.0 90480.0 104680.0 ;
      RECT  89775.0 106025.0 90480.0 107370.0 ;
      RECT  89775.0 108715.0 90480.0 107370.0 ;
      RECT  89775.0 108715.0 90480.0 110060.0 ;
      RECT  89775.0 111405.0 90480.0 110060.0 ;
      RECT  89775.0 111405.0 90480.0 112750.0 ;
      RECT  89775.0 114095.0 90480.0 112750.0 ;
      RECT  90480.0 28015.0 91185.0 29360.0 ;
      RECT  90480.0 30705.0 91185.0 29360.0 ;
      RECT  90480.0 30705.0 91185.0 32050.0 ;
      RECT  90480.0 33395.0 91185.0 32050.0 ;
      RECT  90480.0 33395.0 91185.0 34740.0 ;
      RECT  90480.0 36085.0 91185.0 34740.0 ;
      RECT  90480.0 36085.0 91185.0 37430.0 ;
      RECT  90480.0 38775.0 91185.0 37430.0 ;
      RECT  90480.0 38775.0 91185.0 40120.0 ;
      RECT  90480.0 41465.0 91185.0 40120.0 ;
      RECT  90480.0 41465.0 91185.0 42810.0 ;
      RECT  90480.0 44155.0 91185.0 42810.0 ;
      RECT  90480.0 44155.0 91185.0 45500.0 ;
      RECT  90480.0 46845.0 91185.0 45500.0 ;
      RECT  90480.0 46845.0 91185.0 48190.0 ;
      RECT  90480.0 49535.0 91185.0 48190.0 ;
      RECT  90480.0 49535.0 91185.0 50880.0 ;
      RECT  90480.0 52225.0 91185.0 50880.0 ;
      RECT  90480.0 52225.0 91185.0 53570.0 ;
      RECT  90480.0 54915.0 91185.0 53570.0 ;
      RECT  90480.0 54915.0 91185.0 56260.0 ;
      RECT  90480.0 57605.0 91185.0 56260.0 ;
      RECT  90480.0 57605.0 91185.0 58950.0 ;
      RECT  90480.0 60295.0 91185.0 58950.0 ;
      RECT  90480.0 60295.0 91185.0 61640.0 ;
      RECT  90480.0 62985.0 91185.0 61640.0 ;
      RECT  90480.0 62985.0 91185.0 64330.0 ;
      RECT  90480.0 65675.0 91185.0 64330.0 ;
      RECT  90480.0 65675.0 91185.0 67020.0 ;
      RECT  90480.0 68365.0 91185.0 67020.0 ;
      RECT  90480.0 68365.0 91185.0 69710.0 ;
      RECT  90480.0 71055.0 91185.0 69710.0 ;
      RECT  90480.0 71055.0 91185.0 72400.0 ;
      RECT  90480.0 73745.0 91185.0 72400.0 ;
      RECT  90480.0 73745.0 91185.0 75090.0 ;
      RECT  90480.0 76435.0 91185.0 75090.0 ;
      RECT  90480.0 76435.0 91185.0 77780.0 ;
      RECT  90480.0 79125.0 91185.0 77780.0 ;
      RECT  90480.0 79125.0 91185.0 80470.0 ;
      RECT  90480.0 81815.0 91185.0 80470.0 ;
      RECT  90480.0 81815.0 91185.0 83160.0 ;
      RECT  90480.0 84505.0 91185.0 83160.0 ;
      RECT  90480.0 84505.0 91185.0 85850.0 ;
      RECT  90480.0 87195.0 91185.0 85850.0 ;
      RECT  90480.0 87195.0 91185.0 88540.0 ;
      RECT  90480.0 89885.0 91185.0 88540.0 ;
      RECT  90480.0 89885.0 91185.0 91230.0 ;
      RECT  90480.0 92575.0 91185.0 91230.0 ;
      RECT  90480.0 92575.0 91185.0 93920.0 ;
      RECT  90480.0 95265.0 91185.0 93920.0 ;
      RECT  90480.0 95265.0 91185.0 96610.0 ;
      RECT  90480.0 97955.0 91185.0 96610.0 ;
      RECT  90480.0 97955.0 91185.0 99300.0 ;
      RECT  90480.0 100645.0 91185.0 99300.0 ;
      RECT  90480.0 100645.0 91185.0 101990.0 ;
      RECT  90480.0 103335.0 91185.0 101990.0 ;
      RECT  90480.0 103335.0 91185.0 104680.0 ;
      RECT  90480.0 106025.0 91185.0 104680.0 ;
      RECT  90480.0 106025.0 91185.0 107370.0 ;
      RECT  90480.0 108715.0 91185.0 107370.0 ;
      RECT  90480.0 108715.0 91185.0 110060.0 ;
      RECT  90480.0 111405.0 91185.0 110060.0 ;
      RECT  90480.0 111405.0 91185.0 112750.0 ;
      RECT  90480.0 114095.0 91185.0 112750.0 ;
      RECT  91185.0 28015.0 91890.0 29360.0 ;
      RECT  91185.0 30705.0 91890.0 29360.0 ;
      RECT  91185.0 30705.0 91890.0 32050.0 ;
      RECT  91185.0 33395.0 91890.0 32050.0 ;
      RECT  91185.0 33395.0 91890.0 34740.0 ;
      RECT  91185.0 36085.0 91890.0 34740.0 ;
      RECT  91185.0 36085.0 91890.0 37430.0 ;
      RECT  91185.0 38775.0 91890.0 37430.0 ;
      RECT  91185.0 38775.0 91890.0 40120.0 ;
      RECT  91185.0 41465.0 91890.0 40120.0 ;
      RECT  91185.0 41465.0 91890.0 42810.0 ;
      RECT  91185.0 44155.0 91890.0 42810.0 ;
      RECT  91185.0 44155.0 91890.0 45500.0 ;
      RECT  91185.0 46845.0 91890.0 45500.0 ;
      RECT  91185.0 46845.0 91890.0 48190.0 ;
      RECT  91185.0 49535.0 91890.0 48190.0 ;
      RECT  91185.0 49535.0 91890.0 50880.0 ;
      RECT  91185.0 52225.0 91890.0 50880.0 ;
      RECT  91185.0 52225.0 91890.0 53570.0 ;
      RECT  91185.0 54915.0 91890.0 53570.0 ;
      RECT  91185.0 54915.0 91890.0 56260.0 ;
      RECT  91185.0 57605.0 91890.0 56260.0 ;
      RECT  91185.0 57605.0 91890.0 58950.0 ;
      RECT  91185.0 60295.0 91890.0 58950.0 ;
      RECT  91185.0 60295.0 91890.0 61640.0 ;
      RECT  91185.0 62985.0 91890.0 61640.0 ;
      RECT  91185.0 62985.0 91890.0 64330.0 ;
      RECT  91185.0 65675.0 91890.0 64330.0 ;
      RECT  91185.0 65675.0 91890.0 67020.0 ;
      RECT  91185.0 68365.0 91890.0 67020.0 ;
      RECT  91185.0 68365.0 91890.0 69710.0 ;
      RECT  91185.0 71055.0 91890.0 69710.0 ;
      RECT  91185.0 71055.0 91890.0 72400.0 ;
      RECT  91185.0 73745.0 91890.0 72400.0 ;
      RECT  91185.0 73745.0 91890.0 75090.0 ;
      RECT  91185.0 76435.0 91890.0 75090.0 ;
      RECT  91185.0 76435.0 91890.0 77780.0 ;
      RECT  91185.0 79125.0 91890.0 77780.0 ;
      RECT  91185.0 79125.0 91890.0 80470.0 ;
      RECT  91185.0 81815.0 91890.0 80470.0 ;
      RECT  91185.0 81815.0 91890.0 83160.0 ;
      RECT  91185.0 84505.0 91890.0 83160.0 ;
      RECT  91185.0 84505.0 91890.0 85850.0 ;
      RECT  91185.0 87195.0 91890.0 85850.0 ;
      RECT  91185.0 87195.0 91890.0 88540.0 ;
      RECT  91185.0 89885.0 91890.0 88540.0 ;
      RECT  91185.0 89885.0 91890.0 91230.0 ;
      RECT  91185.0 92575.0 91890.0 91230.0 ;
      RECT  91185.0 92575.0 91890.0 93920.0 ;
      RECT  91185.0 95265.0 91890.0 93920.0 ;
      RECT  91185.0 95265.0 91890.0 96610.0 ;
      RECT  91185.0 97955.0 91890.0 96610.0 ;
      RECT  91185.0 97955.0 91890.0 99300.0 ;
      RECT  91185.0 100645.0 91890.0 99300.0 ;
      RECT  91185.0 100645.0 91890.0 101990.0 ;
      RECT  91185.0 103335.0 91890.0 101990.0 ;
      RECT  91185.0 103335.0 91890.0 104680.0 ;
      RECT  91185.0 106025.0 91890.0 104680.0 ;
      RECT  91185.0 106025.0 91890.0 107370.0 ;
      RECT  91185.0 108715.0 91890.0 107370.0 ;
      RECT  91185.0 108715.0 91890.0 110060.0 ;
      RECT  91185.0 111405.0 91890.0 110060.0 ;
      RECT  91185.0 111405.0 91890.0 112750.0 ;
      RECT  91185.0 114095.0 91890.0 112750.0 ;
      RECT  91890.0 28015.0 92595.0 29360.0 ;
      RECT  91890.0 30705.0 92595.0 29360.0 ;
      RECT  91890.0 30705.0 92595.0 32050.0 ;
      RECT  91890.0 33395.0 92595.0 32050.0 ;
      RECT  91890.0 33395.0 92595.0 34740.0 ;
      RECT  91890.0 36085.0 92595.0 34740.0 ;
      RECT  91890.0 36085.0 92595.0 37430.0 ;
      RECT  91890.0 38775.0 92595.0 37430.0 ;
      RECT  91890.0 38775.0 92595.0 40120.0 ;
      RECT  91890.0 41465.0 92595.0 40120.0 ;
      RECT  91890.0 41465.0 92595.0 42810.0 ;
      RECT  91890.0 44155.0 92595.0 42810.0 ;
      RECT  91890.0 44155.0 92595.0 45500.0 ;
      RECT  91890.0 46845.0 92595.0 45500.0 ;
      RECT  91890.0 46845.0 92595.0 48190.0 ;
      RECT  91890.0 49535.0 92595.0 48190.0 ;
      RECT  91890.0 49535.0 92595.0 50880.0 ;
      RECT  91890.0 52225.0 92595.0 50880.0 ;
      RECT  91890.0 52225.0 92595.0 53570.0 ;
      RECT  91890.0 54915.0 92595.0 53570.0 ;
      RECT  91890.0 54915.0 92595.0 56260.0 ;
      RECT  91890.0 57605.0 92595.0 56260.0 ;
      RECT  91890.0 57605.0 92595.0 58950.0 ;
      RECT  91890.0 60295.0 92595.0 58950.0 ;
      RECT  91890.0 60295.0 92595.0 61640.0 ;
      RECT  91890.0 62985.0 92595.0 61640.0 ;
      RECT  91890.0 62985.0 92595.0 64330.0 ;
      RECT  91890.0 65675.0 92595.0 64330.0 ;
      RECT  91890.0 65675.0 92595.0 67020.0 ;
      RECT  91890.0 68365.0 92595.0 67020.0 ;
      RECT  91890.0 68365.0 92595.0 69710.0 ;
      RECT  91890.0 71055.0 92595.0 69710.0 ;
      RECT  91890.0 71055.0 92595.0 72400.0 ;
      RECT  91890.0 73745.0 92595.0 72400.0 ;
      RECT  91890.0 73745.0 92595.0 75090.0 ;
      RECT  91890.0 76435.0 92595.0 75090.0 ;
      RECT  91890.0 76435.0 92595.0 77780.0 ;
      RECT  91890.0 79125.0 92595.0 77780.0 ;
      RECT  91890.0 79125.0 92595.0 80470.0 ;
      RECT  91890.0 81815.0 92595.0 80470.0 ;
      RECT  91890.0 81815.0 92595.0 83160.0 ;
      RECT  91890.0 84505.0 92595.0 83160.0 ;
      RECT  91890.0 84505.0 92595.0 85850.0 ;
      RECT  91890.0 87195.0 92595.0 85850.0 ;
      RECT  91890.0 87195.0 92595.0 88540.0 ;
      RECT  91890.0 89885.0 92595.0 88540.0 ;
      RECT  91890.0 89885.0 92595.0 91230.0 ;
      RECT  91890.0 92575.0 92595.0 91230.0 ;
      RECT  91890.0 92575.0 92595.0 93920.0 ;
      RECT  91890.0 95265.0 92595.0 93920.0 ;
      RECT  91890.0 95265.0 92595.0 96610.0 ;
      RECT  91890.0 97955.0 92595.0 96610.0 ;
      RECT  91890.0 97955.0 92595.0 99300.0 ;
      RECT  91890.0 100645.0 92595.0 99300.0 ;
      RECT  91890.0 100645.0 92595.0 101990.0 ;
      RECT  91890.0 103335.0 92595.0 101990.0 ;
      RECT  91890.0 103335.0 92595.0 104680.0 ;
      RECT  91890.0 106025.0 92595.0 104680.0 ;
      RECT  91890.0 106025.0 92595.0 107370.0 ;
      RECT  91890.0 108715.0 92595.0 107370.0 ;
      RECT  91890.0 108715.0 92595.0 110060.0 ;
      RECT  91890.0 111405.0 92595.0 110060.0 ;
      RECT  91890.0 111405.0 92595.0 112750.0 ;
      RECT  91890.0 114095.0 92595.0 112750.0 ;
      RECT  92595.0 28015.0 93300.0 29360.0 ;
      RECT  92595.0 30705.0 93300.0 29360.0 ;
      RECT  92595.0 30705.0 93300.0 32050.0 ;
      RECT  92595.0 33395.0 93300.0 32050.0 ;
      RECT  92595.0 33395.0 93300.0 34740.0 ;
      RECT  92595.0 36085.0 93300.0 34740.0 ;
      RECT  92595.0 36085.0 93300.0 37430.0 ;
      RECT  92595.0 38775.0 93300.0 37430.0 ;
      RECT  92595.0 38775.0 93300.0 40120.0 ;
      RECT  92595.0 41465.0 93300.0 40120.0 ;
      RECT  92595.0 41465.0 93300.0 42810.0 ;
      RECT  92595.0 44155.0 93300.0 42810.0 ;
      RECT  92595.0 44155.0 93300.0 45500.0 ;
      RECT  92595.0 46845.0 93300.0 45500.0 ;
      RECT  92595.0 46845.0 93300.0 48190.0 ;
      RECT  92595.0 49535.0 93300.0 48190.0 ;
      RECT  92595.0 49535.0 93300.0 50880.0 ;
      RECT  92595.0 52225.0 93300.0 50880.0 ;
      RECT  92595.0 52225.0 93300.0 53570.0 ;
      RECT  92595.0 54915.0 93300.0 53570.0 ;
      RECT  92595.0 54915.0 93300.0 56260.0 ;
      RECT  92595.0 57605.0 93300.0 56260.0 ;
      RECT  92595.0 57605.0 93300.0 58950.0 ;
      RECT  92595.0 60295.0 93300.0 58950.0 ;
      RECT  92595.0 60295.0 93300.0 61640.0 ;
      RECT  92595.0 62985.0 93300.0 61640.0 ;
      RECT  92595.0 62985.0 93300.0 64330.0 ;
      RECT  92595.0 65675.0 93300.0 64330.0 ;
      RECT  92595.0 65675.0 93300.0 67020.0 ;
      RECT  92595.0 68365.0 93300.0 67020.0 ;
      RECT  92595.0 68365.0 93300.0 69710.0 ;
      RECT  92595.0 71055.0 93300.0 69710.0 ;
      RECT  92595.0 71055.0 93300.0 72400.0 ;
      RECT  92595.0 73745.0 93300.0 72400.0 ;
      RECT  92595.0 73745.0 93300.0 75090.0 ;
      RECT  92595.0 76435.0 93300.0 75090.0 ;
      RECT  92595.0 76435.0 93300.0 77780.0 ;
      RECT  92595.0 79125.0 93300.0 77780.0 ;
      RECT  92595.0 79125.0 93300.0 80470.0 ;
      RECT  92595.0 81815.0 93300.0 80470.0 ;
      RECT  92595.0 81815.0 93300.0 83160.0 ;
      RECT  92595.0 84505.0 93300.0 83160.0 ;
      RECT  92595.0 84505.0 93300.0 85850.0 ;
      RECT  92595.0 87195.0 93300.0 85850.0 ;
      RECT  92595.0 87195.0 93300.0 88540.0 ;
      RECT  92595.0 89885.0 93300.0 88540.0 ;
      RECT  92595.0 89885.0 93300.0 91230.0 ;
      RECT  92595.0 92575.0 93300.0 91230.0 ;
      RECT  92595.0 92575.0 93300.0 93920.0 ;
      RECT  92595.0 95265.0 93300.0 93920.0 ;
      RECT  92595.0 95265.0 93300.0 96610.0 ;
      RECT  92595.0 97955.0 93300.0 96610.0 ;
      RECT  92595.0 97955.0 93300.0 99300.0 ;
      RECT  92595.0 100645.0 93300.0 99300.0 ;
      RECT  92595.0 100645.0 93300.0 101990.0 ;
      RECT  92595.0 103335.0 93300.0 101990.0 ;
      RECT  92595.0 103335.0 93300.0 104680.0 ;
      RECT  92595.0 106025.0 93300.0 104680.0 ;
      RECT  92595.0 106025.0 93300.0 107370.0 ;
      RECT  92595.0 108715.0 93300.0 107370.0 ;
      RECT  92595.0 108715.0 93300.0 110060.0 ;
      RECT  92595.0 111405.0 93300.0 110060.0 ;
      RECT  92595.0 111405.0 93300.0 112750.0 ;
      RECT  92595.0 114095.0 93300.0 112750.0 ;
      RECT  93300.0 28015.0 94005.0 29360.0 ;
      RECT  93300.0 30705.0 94005.0 29360.0 ;
      RECT  93300.0 30705.0 94005.0 32050.0 ;
      RECT  93300.0 33395.0 94005.0 32050.0 ;
      RECT  93300.0 33395.0 94005.0 34740.0 ;
      RECT  93300.0 36085.0 94005.0 34740.0 ;
      RECT  93300.0 36085.0 94005.0 37430.0 ;
      RECT  93300.0 38775.0 94005.0 37430.0 ;
      RECT  93300.0 38775.0 94005.0 40120.0 ;
      RECT  93300.0 41465.0 94005.0 40120.0 ;
      RECT  93300.0 41465.0 94005.0 42810.0 ;
      RECT  93300.0 44155.0 94005.0 42810.0 ;
      RECT  93300.0 44155.0 94005.0 45500.0 ;
      RECT  93300.0 46845.0 94005.0 45500.0 ;
      RECT  93300.0 46845.0 94005.0 48190.0 ;
      RECT  93300.0 49535.0 94005.0 48190.0 ;
      RECT  93300.0 49535.0 94005.0 50880.0 ;
      RECT  93300.0 52225.0 94005.0 50880.0 ;
      RECT  93300.0 52225.0 94005.0 53570.0 ;
      RECT  93300.0 54915.0 94005.0 53570.0 ;
      RECT  93300.0 54915.0 94005.0 56260.0 ;
      RECT  93300.0 57605.0 94005.0 56260.0 ;
      RECT  93300.0 57605.0 94005.0 58950.0 ;
      RECT  93300.0 60295.0 94005.0 58950.0 ;
      RECT  93300.0 60295.0 94005.0 61640.0 ;
      RECT  93300.0 62985.0 94005.0 61640.0 ;
      RECT  93300.0 62985.0 94005.0 64330.0 ;
      RECT  93300.0 65675.0 94005.0 64330.0 ;
      RECT  93300.0 65675.0 94005.0 67020.0 ;
      RECT  93300.0 68365.0 94005.0 67020.0 ;
      RECT  93300.0 68365.0 94005.0 69710.0 ;
      RECT  93300.0 71055.0 94005.0 69710.0 ;
      RECT  93300.0 71055.0 94005.0 72400.0 ;
      RECT  93300.0 73745.0 94005.0 72400.0 ;
      RECT  93300.0 73745.0 94005.0 75090.0 ;
      RECT  93300.0 76435.0 94005.0 75090.0 ;
      RECT  93300.0 76435.0 94005.0 77780.0 ;
      RECT  93300.0 79125.0 94005.0 77780.0 ;
      RECT  93300.0 79125.0 94005.0 80470.0 ;
      RECT  93300.0 81815.0 94005.0 80470.0 ;
      RECT  93300.0 81815.0 94005.0 83160.0 ;
      RECT  93300.0 84505.0 94005.0 83160.0 ;
      RECT  93300.0 84505.0 94005.0 85850.0 ;
      RECT  93300.0 87195.0 94005.0 85850.0 ;
      RECT  93300.0 87195.0 94005.0 88540.0 ;
      RECT  93300.0 89885.0 94005.0 88540.0 ;
      RECT  93300.0 89885.0 94005.0 91230.0 ;
      RECT  93300.0 92575.0 94005.0 91230.0 ;
      RECT  93300.0 92575.0 94005.0 93920.0 ;
      RECT  93300.0 95265.0 94005.0 93920.0 ;
      RECT  93300.0 95265.0 94005.0 96610.0 ;
      RECT  93300.0 97955.0 94005.0 96610.0 ;
      RECT  93300.0 97955.0 94005.0 99300.0 ;
      RECT  93300.0 100645.0 94005.0 99300.0 ;
      RECT  93300.0 100645.0 94005.0 101990.0 ;
      RECT  93300.0 103335.0 94005.0 101990.0 ;
      RECT  93300.0 103335.0 94005.0 104680.0 ;
      RECT  93300.0 106025.0 94005.0 104680.0 ;
      RECT  93300.0 106025.0 94005.0 107370.0 ;
      RECT  93300.0 108715.0 94005.0 107370.0 ;
      RECT  93300.0 108715.0 94005.0 110060.0 ;
      RECT  93300.0 111405.0 94005.0 110060.0 ;
      RECT  93300.0 111405.0 94005.0 112750.0 ;
      RECT  93300.0 114095.0 94005.0 112750.0 ;
      RECT  94005.0 28015.0 94710.0 29360.0 ;
      RECT  94005.0 30705.0 94710.0 29360.0 ;
      RECT  94005.0 30705.0 94710.0 32050.0 ;
      RECT  94005.0 33395.0 94710.0 32050.0 ;
      RECT  94005.0 33395.0 94710.0 34740.0 ;
      RECT  94005.0 36085.0 94710.0 34740.0 ;
      RECT  94005.0 36085.0 94710.0 37430.0 ;
      RECT  94005.0 38775.0 94710.0 37430.0 ;
      RECT  94005.0 38775.0 94710.0 40120.0 ;
      RECT  94005.0 41465.0 94710.0 40120.0 ;
      RECT  94005.0 41465.0 94710.0 42810.0 ;
      RECT  94005.0 44155.0 94710.0 42810.0 ;
      RECT  94005.0 44155.0 94710.0 45500.0 ;
      RECT  94005.0 46845.0 94710.0 45500.0 ;
      RECT  94005.0 46845.0 94710.0 48190.0 ;
      RECT  94005.0 49535.0 94710.0 48190.0 ;
      RECT  94005.0 49535.0 94710.0 50880.0 ;
      RECT  94005.0 52225.0 94710.0 50880.0 ;
      RECT  94005.0 52225.0 94710.0 53570.0 ;
      RECT  94005.0 54915.0 94710.0 53570.0 ;
      RECT  94005.0 54915.0 94710.0 56260.0 ;
      RECT  94005.0 57605.0 94710.0 56260.0 ;
      RECT  94005.0 57605.0 94710.0 58950.0 ;
      RECT  94005.0 60295.0 94710.0 58950.0 ;
      RECT  94005.0 60295.0 94710.0 61640.0 ;
      RECT  94005.0 62985.0 94710.0 61640.0 ;
      RECT  94005.0 62985.0 94710.0 64330.0 ;
      RECT  94005.0 65675.0 94710.0 64330.0 ;
      RECT  94005.0 65675.0 94710.0 67020.0 ;
      RECT  94005.0 68365.0 94710.0 67020.0 ;
      RECT  94005.0 68365.0 94710.0 69710.0 ;
      RECT  94005.0 71055.0 94710.0 69710.0 ;
      RECT  94005.0 71055.0 94710.0 72400.0 ;
      RECT  94005.0 73745.0 94710.0 72400.0 ;
      RECT  94005.0 73745.0 94710.0 75090.0 ;
      RECT  94005.0 76435.0 94710.0 75090.0 ;
      RECT  94005.0 76435.0 94710.0 77780.0 ;
      RECT  94005.0 79125.0 94710.0 77780.0 ;
      RECT  94005.0 79125.0 94710.0 80470.0 ;
      RECT  94005.0 81815.0 94710.0 80470.0 ;
      RECT  94005.0 81815.0 94710.0 83160.0 ;
      RECT  94005.0 84505.0 94710.0 83160.0 ;
      RECT  94005.0 84505.0 94710.0 85850.0 ;
      RECT  94005.0 87195.0 94710.0 85850.0 ;
      RECT  94005.0 87195.0 94710.0 88540.0 ;
      RECT  94005.0 89885.0 94710.0 88540.0 ;
      RECT  94005.0 89885.0 94710.0 91230.0 ;
      RECT  94005.0 92575.0 94710.0 91230.0 ;
      RECT  94005.0 92575.0 94710.0 93920.0 ;
      RECT  94005.0 95265.0 94710.0 93920.0 ;
      RECT  94005.0 95265.0 94710.0 96610.0 ;
      RECT  94005.0 97955.0 94710.0 96610.0 ;
      RECT  94005.0 97955.0 94710.0 99300.0 ;
      RECT  94005.0 100645.0 94710.0 99300.0 ;
      RECT  94005.0 100645.0 94710.0 101990.0 ;
      RECT  94005.0 103335.0 94710.0 101990.0 ;
      RECT  94005.0 103335.0 94710.0 104680.0 ;
      RECT  94005.0 106025.0 94710.0 104680.0 ;
      RECT  94005.0 106025.0 94710.0 107370.0 ;
      RECT  94005.0 108715.0 94710.0 107370.0 ;
      RECT  94005.0 108715.0 94710.0 110060.0 ;
      RECT  94005.0 111405.0 94710.0 110060.0 ;
      RECT  94005.0 111405.0 94710.0 112750.0 ;
      RECT  94005.0 114095.0 94710.0 112750.0 ;
      RECT  94710.0 28015.0 95415.0 29360.0 ;
      RECT  94710.0 30705.0 95415.0 29360.0 ;
      RECT  94710.0 30705.0 95415.0 32050.0 ;
      RECT  94710.0 33395.0 95415.0 32050.0 ;
      RECT  94710.0 33395.0 95415.0 34740.0 ;
      RECT  94710.0 36085.0 95415.0 34740.0 ;
      RECT  94710.0 36085.0 95415.0 37430.0 ;
      RECT  94710.0 38775.0 95415.0 37430.0 ;
      RECT  94710.0 38775.0 95415.0 40120.0 ;
      RECT  94710.0 41465.0 95415.0 40120.0 ;
      RECT  94710.0 41465.0 95415.0 42810.0 ;
      RECT  94710.0 44155.0 95415.0 42810.0 ;
      RECT  94710.0 44155.0 95415.0 45500.0 ;
      RECT  94710.0 46845.0 95415.0 45500.0 ;
      RECT  94710.0 46845.0 95415.0 48190.0 ;
      RECT  94710.0 49535.0 95415.0 48190.0 ;
      RECT  94710.0 49535.0 95415.0 50880.0 ;
      RECT  94710.0 52225.0 95415.0 50880.0 ;
      RECT  94710.0 52225.0 95415.0 53570.0 ;
      RECT  94710.0 54915.0 95415.0 53570.0 ;
      RECT  94710.0 54915.0 95415.0 56260.0 ;
      RECT  94710.0 57605.0 95415.0 56260.0 ;
      RECT  94710.0 57605.0 95415.0 58950.0 ;
      RECT  94710.0 60295.0 95415.0 58950.0 ;
      RECT  94710.0 60295.0 95415.0 61640.0 ;
      RECT  94710.0 62985.0 95415.0 61640.0 ;
      RECT  94710.0 62985.0 95415.0 64330.0 ;
      RECT  94710.0 65675.0 95415.0 64330.0 ;
      RECT  94710.0 65675.0 95415.0 67020.0 ;
      RECT  94710.0 68365.0 95415.0 67020.0 ;
      RECT  94710.0 68365.0 95415.0 69710.0 ;
      RECT  94710.0 71055.0 95415.0 69710.0 ;
      RECT  94710.0 71055.0 95415.0 72400.0 ;
      RECT  94710.0 73745.0 95415.0 72400.0 ;
      RECT  94710.0 73745.0 95415.0 75090.0 ;
      RECT  94710.0 76435.0 95415.0 75090.0 ;
      RECT  94710.0 76435.0 95415.0 77780.0 ;
      RECT  94710.0 79125.0 95415.0 77780.0 ;
      RECT  94710.0 79125.0 95415.0 80470.0 ;
      RECT  94710.0 81815.0 95415.0 80470.0 ;
      RECT  94710.0 81815.0 95415.0 83160.0 ;
      RECT  94710.0 84505.0 95415.0 83160.0 ;
      RECT  94710.0 84505.0 95415.0 85850.0 ;
      RECT  94710.0 87195.0 95415.0 85850.0 ;
      RECT  94710.0 87195.0 95415.0 88540.0 ;
      RECT  94710.0 89885.0 95415.0 88540.0 ;
      RECT  94710.0 89885.0 95415.0 91230.0 ;
      RECT  94710.0 92575.0 95415.0 91230.0 ;
      RECT  94710.0 92575.0 95415.0 93920.0 ;
      RECT  94710.0 95265.0 95415.0 93920.0 ;
      RECT  94710.0 95265.0 95415.0 96610.0 ;
      RECT  94710.0 97955.0 95415.0 96610.0 ;
      RECT  94710.0 97955.0 95415.0 99300.0 ;
      RECT  94710.0 100645.0 95415.0 99300.0 ;
      RECT  94710.0 100645.0 95415.0 101990.0 ;
      RECT  94710.0 103335.0 95415.0 101990.0 ;
      RECT  94710.0 103335.0 95415.0 104680.0 ;
      RECT  94710.0 106025.0 95415.0 104680.0 ;
      RECT  94710.0 106025.0 95415.0 107370.0 ;
      RECT  94710.0 108715.0 95415.0 107370.0 ;
      RECT  94710.0 108715.0 95415.0 110060.0 ;
      RECT  94710.0 111405.0 95415.0 110060.0 ;
      RECT  94710.0 111405.0 95415.0 112750.0 ;
      RECT  94710.0 114095.0 95415.0 112750.0 ;
      RECT  95415.0 28015.0 96120.0 29360.0 ;
      RECT  95415.0 30705.0 96120.0 29360.0 ;
      RECT  95415.0 30705.0 96120.0 32050.0 ;
      RECT  95415.0 33395.0 96120.0 32050.0 ;
      RECT  95415.0 33395.0 96120.0 34740.0 ;
      RECT  95415.0 36085.0 96120.0 34740.0 ;
      RECT  95415.0 36085.0 96120.0 37430.0 ;
      RECT  95415.0 38775.0 96120.0 37430.0 ;
      RECT  95415.0 38775.0 96120.0 40120.0 ;
      RECT  95415.0 41465.0 96120.0 40120.0 ;
      RECT  95415.0 41465.0 96120.0 42810.0 ;
      RECT  95415.0 44155.0 96120.0 42810.0 ;
      RECT  95415.0 44155.0 96120.0 45500.0 ;
      RECT  95415.0 46845.0 96120.0 45500.0 ;
      RECT  95415.0 46845.0 96120.0 48190.0 ;
      RECT  95415.0 49535.0 96120.0 48190.0 ;
      RECT  95415.0 49535.0 96120.0 50880.0 ;
      RECT  95415.0 52225.0 96120.0 50880.0 ;
      RECT  95415.0 52225.0 96120.0 53570.0 ;
      RECT  95415.0 54915.0 96120.0 53570.0 ;
      RECT  95415.0 54915.0 96120.0 56260.0 ;
      RECT  95415.0 57605.0 96120.0 56260.0 ;
      RECT  95415.0 57605.0 96120.0 58950.0 ;
      RECT  95415.0 60295.0 96120.0 58950.0 ;
      RECT  95415.0 60295.0 96120.0 61640.0 ;
      RECT  95415.0 62985.0 96120.0 61640.0 ;
      RECT  95415.0 62985.0 96120.0 64330.0 ;
      RECT  95415.0 65675.0 96120.0 64330.0 ;
      RECT  95415.0 65675.0 96120.0 67020.0 ;
      RECT  95415.0 68365.0 96120.0 67020.0 ;
      RECT  95415.0 68365.0 96120.0 69710.0 ;
      RECT  95415.0 71055.0 96120.0 69710.0 ;
      RECT  95415.0 71055.0 96120.0 72400.0 ;
      RECT  95415.0 73745.0 96120.0 72400.0 ;
      RECT  95415.0 73745.0 96120.0 75090.0 ;
      RECT  95415.0 76435.0 96120.0 75090.0 ;
      RECT  95415.0 76435.0 96120.0 77780.0 ;
      RECT  95415.0 79125.0 96120.0 77780.0 ;
      RECT  95415.0 79125.0 96120.0 80470.0 ;
      RECT  95415.0 81815.0 96120.0 80470.0 ;
      RECT  95415.0 81815.0 96120.0 83160.0 ;
      RECT  95415.0 84505.0 96120.0 83160.0 ;
      RECT  95415.0 84505.0 96120.0 85850.0 ;
      RECT  95415.0 87195.0 96120.0 85850.0 ;
      RECT  95415.0 87195.0 96120.0 88540.0 ;
      RECT  95415.0 89885.0 96120.0 88540.0 ;
      RECT  95415.0 89885.0 96120.0 91230.0 ;
      RECT  95415.0 92575.0 96120.0 91230.0 ;
      RECT  95415.0 92575.0 96120.0 93920.0 ;
      RECT  95415.0 95265.0 96120.0 93920.0 ;
      RECT  95415.0 95265.0 96120.0 96610.0 ;
      RECT  95415.0 97955.0 96120.0 96610.0 ;
      RECT  95415.0 97955.0 96120.0 99300.0 ;
      RECT  95415.0 100645.0 96120.0 99300.0 ;
      RECT  95415.0 100645.0 96120.0 101990.0 ;
      RECT  95415.0 103335.0 96120.0 101990.0 ;
      RECT  95415.0 103335.0 96120.0 104680.0 ;
      RECT  95415.0 106025.0 96120.0 104680.0 ;
      RECT  95415.0 106025.0 96120.0 107370.0 ;
      RECT  95415.0 108715.0 96120.0 107370.0 ;
      RECT  95415.0 108715.0 96120.0 110060.0 ;
      RECT  95415.0 111405.0 96120.0 110060.0 ;
      RECT  95415.0 111405.0 96120.0 112750.0 ;
      RECT  95415.0 114095.0 96120.0 112750.0 ;
      RECT  96120.0 28015.0 96825.0 29360.0 ;
      RECT  96120.0 30705.0 96825.0 29360.0 ;
      RECT  96120.0 30705.0 96825.0 32050.0 ;
      RECT  96120.0 33395.0 96825.0 32050.0 ;
      RECT  96120.0 33395.0 96825.0 34740.0 ;
      RECT  96120.0 36085.0 96825.0 34740.0 ;
      RECT  96120.0 36085.0 96825.0 37430.0 ;
      RECT  96120.0 38775.0 96825.0 37430.0 ;
      RECT  96120.0 38775.0 96825.0 40120.0 ;
      RECT  96120.0 41465.0 96825.0 40120.0 ;
      RECT  96120.0 41465.0 96825.0 42810.0 ;
      RECT  96120.0 44155.0 96825.0 42810.0 ;
      RECT  96120.0 44155.0 96825.0 45500.0 ;
      RECT  96120.0 46845.0 96825.0 45500.0 ;
      RECT  96120.0 46845.0 96825.0 48190.0 ;
      RECT  96120.0 49535.0 96825.0 48190.0 ;
      RECT  96120.0 49535.0 96825.0 50880.0 ;
      RECT  96120.0 52225.0 96825.0 50880.0 ;
      RECT  96120.0 52225.0 96825.0 53570.0 ;
      RECT  96120.0 54915.0 96825.0 53570.0 ;
      RECT  96120.0 54915.0 96825.0 56260.0 ;
      RECT  96120.0 57605.0 96825.0 56260.0 ;
      RECT  96120.0 57605.0 96825.0 58950.0 ;
      RECT  96120.0 60295.0 96825.0 58950.0 ;
      RECT  96120.0 60295.0 96825.0 61640.0 ;
      RECT  96120.0 62985.0 96825.0 61640.0 ;
      RECT  96120.0 62985.0 96825.0 64330.0 ;
      RECT  96120.0 65675.0 96825.0 64330.0 ;
      RECT  96120.0 65675.0 96825.0 67020.0 ;
      RECT  96120.0 68365.0 96825.0 67020.0 ;
      RECT  96120.0 68365.0 96825.0 69710.0 ;
      RECT  96120.0 71055.0 96825.0 69710.0 ;
      RECT  96120.0 71055.0 96825.0 72400.0 ;
      RECT  96120.0 73745.0 96825.0 72400.0 ;
      RECT  96120.0 73745.0 96825.0 75090.0 ;
      RECT  96120.0 76435.0 96825.0 75090.0 ;
      RECT  96120.0 76435.0 96825.0 77780.0 ;
      RECT  96120.0 79125.0 96825.0 77780.0 ;
      RECT  96120.0 79125.0 96825.0 80470.0 ;
      RECT  96120.0 81815.0 96825.0 80470.0 ;
      RECT  96120.0 81815.0 96825.0 83160.0 ;
      RECT  96120.0 84505.0 96825.0 83160.0 ;
      RECT  96120.0 84505.0 96825.0 85850.0 ;
      RECT  96120.0 87195.0 96825.0 85850.0 ;
      RECT  96120.0 87195.0 96825.0 88540.0 ;
      RECT  96120.0 89885.0 96825.0 88540.0 ;
      RECT  96120.0 89885.0 96825.0 91230.0 ;
      RECT  96120.0 92575.0 96825.0 91230.0 ;
      RECT  96120.0 92575.0 96825.0 93920.0 ;
      RECT  96120.0 95265.0 96825.0 93920.0 ;
      RECT  96120.0 95265.0 96825.0 96610.0 ;
      RECT  96120.0 97955.0 96825.0 96610.0 ;
      RECT  96120.0 97955.0 96825.0 99300.0 ;
      RECT  96120.0 100645.0 96825.0 99300.0 ;
      RECT  96120.0 100645.0 96825.0 101990.0 ;
      RECT  96120.0 103335.0 96825.0 101990.0 ;
      RECT  96120.0 103335.0 96825.0 104680.0 ;
      RECT  96120.0 106025.0 96825.0 104680.0 ;
      RECT  96120.0 106025.0 96825.0 107370.0 ;
      RECT  96120.0 108715.0 96825.0 107370.0 ;
      RECT  96120.0 108715.0 96825.0 110060.0 ;
      RECT  96120.0 111405.0 96825.0 110060.0 ;
      RECT  96120.0 111405.0 96825.0 112750.0 ;
      RECT  96120.0 114095.0 96825.0 112750.0 ;
      RECT  96825.0 28015.0 97530.0 29360.0 ;
      RECT  96825.0 30705.0 97530.0 29360.0 ;
      RECT  96825.0 30705.0 97530.0 32050.0 ;
      RECT  96825.0 33395.0 97530.0 32050.0 ;
      RECT  96825.0 33395.0 97530.0 34740.0 ;
      RECT  96825.0 36085.0 97530.0 34740.0 ;
      RECT  96825.0 36085.0 97530.0 37430.0 ;
      RECT  96825.0 38775.0 97530.0 37430.0 ;
      RECT  96825.0 38775.0 97530.0 40120.0 ;
      RECT  96825.0 41465.0 97530.0 40120.0 ;
      RECT  96825.0 41465.0 97530.0 42810.0 ;
      RECT  96825.0 44155.0 97530.0 42810.0 ;
      RECT  96825.0 44155.0 97530.0 45500.0 ;
      RECT  96825.0 46845.0 97530.0 45500.0 ;
      RECT  96825.0 46845.0 97530.0 48190.0 ;
      RECT  96825.0 49535.0 97530.0 48190.0 ;
      RECT  96825.0 49535.0 97530.0 50880.0 ;
      RECT  96825.0 52225.0 97530.0 50880.0 ;
      RECT  96825.0 52225.0 97530.0 53570.0 ;
      RECT  96825.0 54915.0 97530.0 53570.0 ;
      RECT  96825.0 54915.0 97530.0 56260.0 ;
      RECT  96825.0 57605.0 97530.0 56260.0 ;
      RECT  96825.0 57605.0 97530.0 58950.0 ;
      RECT  96825.0 60295.0 97530.0 58950.0 ;
      RECT  96825.0 60295.0 97530.0 61640.0 ;
      RECT  96825.0 62985.0 97530.0 61640.0 ;
      RECT  96825.0 62985.0 97530.0 64330.0 ;
      RECT  96825.0 65675.0 97530.0 64330.0 ;
      RECT  96825.0 65675.0 97530.0 67020.0 ;
      RECT  96825.0 68365.0 97530.0 67020.0 ;
      RECT  96825.0 68365.0 97530.0 69710.0 ;
      RECT  96825.0 71055.0 97530.0 69710.0 ;
      RECT  96825.0 71055.0 97530.0 72400.0 ;
      RECT  96825.0 73745.0 97530.0 72400.0 ;
      RECT  96825.0 73745.0 97530.0 75090.0 ;
      RECT  96825.0 76435.0 97530.0 75090.0 ;
      RECT  96825.0 76435.0 97530.0 77780.0 ;
      RECT  96825.0 79125.0 97530.0 77780.0 ;
      RECT  96825.0 79125.0 97530.0 80470.0 ;
      RECT  96825.0 81815.0 97530.0 80470.0 ;
      RECT  96825.0 81815.0 97530.0 83160.0 ;
      RECT  96825.0 84505.0 97530.0 83160.0 ;
      RECT  96825.0 84505.0 97530.0 85850.0 ;
      RECT  96825.0 87195.0 97530.0 85850.0 ;
      RECT  96825.0 87195.0 97530.0 88540.0 ;
      RECT  96825.0 89885.0 97530.0 88540.0 ;
      RECT  96825.0 89885.0 97530.0 91230.0 ;
      RECT  96825.0 92575.0 97530.0 91230.0 ;
      RECT  96825.0 92575.0 97530.0 93920.0 ;
      RECT  96825.0 95265.0 97530.0 93920.0 ;
      RECT  96825.0 95265.0 97530.0 96610.0 ;
      RECT  96825.0 97955.0 97530.0 96610.0 ;
      RECT  96825.0 97955.0 97530.0 99300.0 ;
      RECT  96825.0 100645.0 97530.0 99300.0 ;
      RECT  96825.0 100645.0 97530.0 101990.0 ;
      RECT  96825.0 103335.0 97530.0 101990.0 ;
      RECT  96825.0 103335.0 97530.0 104680.0 ;
      RECT  96825.0 106025.0 97530.0 104680.0 ;
      RECT  96825.0 106025.0 97530.0 107370.0 ;
      RECT  96825.0 108715.0 97530.0 107370.0 ;
      RECT  96825.0 108715.0 97530.0 110060.0 ;
      RECT  96825.0 111405.0 97530.0 110060.0 ;
      RECT  96825.0 111405.0 97530.0 112750.0 ;
      RECT  96825.0 114095.0 97530.0 112750.0 ;
      RECT  97530.0 28015.0 98235.0 29360.0 ;
      RECT  97530.0 30705.0 98235.0 29360.0 ;
      RECT  97530.0 30705.0 98235.0 32050.0 ;
      RECT  97530.0 33395.0 98235.0 32050.0 ;
      RECT  97530.0 33395.0 98235.0 34740.0 ;
      RECT  97530.0 36085.0 98235.0 34740.0 ;
      RECT  97530.0 36085.0 98235.0 37430.0 ;
      RECT  97530.0 38775.0 98235.0 37430.0 ;
      RECT  97530.0 38775.0 98235.0 40120.0 ;
      RECT  97530.0 41465.0 98235.0 40120.0 ;
      RECT  97530.0 41465.0 98235.0 42810.0 ;
      RECT  97530.0 44155.0 98235.0 42810.0 ;
      RECT  97530.0 44155.0 98235.0 45500.0 ;
      RECT  97530.0 46845.0 98235.0 45500.0 ;
      RECT  97530.0 46845.0 98235.0 48190.0 ;
      RECT  97530.0 49535.0 98235.0 48190.0 ;
      RECT  97530.0 49535.0 98235.0 50880.0 ;
      RECT  97530.0 52225.0 98235.0 50880.0 ;
      RECT  97530.0 52225.0 98235.0 53570.0 ;
      RECT  97530.0 54915.0 98235.0 53570.0 ;
      RECT  97530.0 54915.0 98235.0 56260.0 ;
      RECT  97530.0 57605.0 98235.0 56260.0 ;
      RECT  97530.0 57605.0 98235.0 58950.0 ;
      RECT  97530.0 60295.0 98235.0 58950.0 ;
      RECT  97530.0 60295.0 98235.0 61640.0 ;
      RECT  97530.0 62985.0 98235.0 61640.0 ;
      RECT  97530.0 62985.0 98235.0 64330.0 ;
      RECT  97530.0 65675.0 98235.0 64330.0 ;
      RECT  97530.0 65675.0 98235.0 67020.0 ;
      RECT  97530.0 68365.0 98235.0 67020.0 ;
      RECT  97530.0 68365.0 98235.0 69710.0 ;
      RECT  97530.0 71055.0 98235.0 69710.0 ;
      RECT  97530.0 71055.0 98235.0 72400.0 ;
      RECT  97530.0 73745.0 98235.0 72400.0 ;
      RECT  97530.0 73745.0 98235.0 75090.0 ;
      RECT  97530.0 76435.0 98235.0 75090.0 ;
      RECT  97530.0 76435.0 98235.0 77780.0 ;
      RECT  97530.0 79125.0 98235.0 77780.0 ;
      RECT  97530.0 79125.0 98235.0 80470.0 ;
      RECT  97530.0 81815.0 98235.0 80470.0 ;
      RECT  97530.0 81815.0 98235.0 83160.0 ;
      RECT  97530.0 84505.0 98235.0 83160.0 ;
      RECT  97530.0 84505.0 98235.0 85850.0 ;
      RECT  97530.0 87195.0 98235.0 85850.0 ;
      RECT  97530.0 87195.0 98235.0 88540.0 ;
      RECT  97530.0 89885.0 98235.0 88540.0 ;
      RECT  97530.0 89885.0 98235.0 91230.0 ;
      RECT  97530.0 92575.0 98235.0 91230.0 ;
      RECT  97530.0 92575.0 98235.0 93920.0 ;
      RECT  97530.0 95265.0 98235.0 93920.0 ;
      RECT  97530.0 95265.0 98235.0 96610.0 ;
      RECT  97530.0 97955.0 98235.0 96610.0 ;
      RECT  97530.0 97955.0 98235.0 99300.0 ;
      RECT  97530.0 100645.0 98235.0 99300.0 ;
      RECT  97530.0 100645.0 98235.0 101990.0 ;
      RECT  97530.0 103335.0 98235.0 101990.0 ;
      RECT  97530.0 103335.0 98235.0 104680.0 ;
      RECT  97530.0 106025.0 98235.0 104680.0 ;
      RECT  97530.0 106025.0 98235.0 107370.0 ;
      RECT  97530.0 108715.0 98235.0 107370.0 ;
      RECT  97530.0 108715.0 98235.0 110060.0 ;
      RECT  97530.0 111405.0 98235.0 110060.0 ;
      RECT  97530.0 111405.0 98235.0 112750.0 ;
      RECT  97530.0 114095.0 98235.0 112750.0 ;
      RECT  98235.0 28015.0 98940.0 29360.0 ;
      RECT  98235.0 30705.0 98940.0 29360.0 ;
      RECT  98235.0 30705.0 98940.0 32050.0 ;
      RECT  98235.0 33395.0 98940.0 32050.0 ;
      RECT  98235.0 33395.0 98940.0 34740.0 ;
      RECT  98235.0 36085.0 98940.0 34740.0 ;
      RECT  98235.0 36085.0 98940.0 37430.0 ;
      RECT  98235.0 38775.0 98940.0 37430.0 ;
      RECT  98235.0 38775.0 98940.0 40120.0 ;
      RECT  98235.0 41465.0 98940.0 40120.0 ;
      RECT  98235.0 41465.0 98940.0 42810.0 ;
      RECT  98235.0 44155.0 98940.0 42810.0 ;
      RECT  98235.0 44155.0 98940.0 45500.0 ;
      RECT  98235.0 46845.0 98940.0 45500.0 ;
      RECT  98235.0 46845.0 98940.0 48190.0 ;
      RECT  98235.0 49535.0 98940.0 48190.0 ;
      RECT  98235.0 49535.0 98940.0 50880.0 ;
      RECT  98235.0 52225.0 98940.0 50880.0 ;
      RECT  98235.0 52225.0 98940.0 53570.0 ;
      RECT  98235.0 54915.0 98940.0 53570.0 ;
      RECT  98235.0 54915.0 98940.0 56260.0 ;
      RECT  98235.0 57605.0 98940.0 56260.0 ;
      RECT  98235.0 57605.0 98940.0 58950.0 ;
      RECT  98235.0 60295.0 98940.0 58950.0 ;
      RECT  98235.0 60295.0 98940.0 61640.0 ;
      RECT  98235.0 62985.0 98940.0 61640.0 ;
      RECT  98235.0 62985.0 98940.0 64330.0 ;
      RECT  98235.0 65675.0 98940.0 64330.0 ;
      RECT  98235.0 65675.0 98940.0 67020.0 ;
      RECT  98235.0 68365.0 98940.0 67020.0 ;
      RECT  98235.0 68365.0 98940.0 69710.0 ;
      RECT  98235.0 71055.0 98940.0 69710.0 ;
      RECT  98235.0 71055.0 98940.0 72400.0 ;
      RECT  98235.0 73745.0 98940.0 72400.0 ;
      RECT  98235.0 73745.0 98940.0 75090.0 ;
      RECT  98235.0 76435.0 98940.0 75090.0 ;
      RECT  98235.0 76435.0 98940.0 77780.0 ;
      RECT  98235.0 79125.0 98940.0 77780.0 ;
      RECT  98235.0 79125.0 98940.0 80470.0 ;
      RECT  98235.0 81815.0 98940.0 80470.0 ;
      RECT  98235.0 81815.0 98940.0 83160.0 ;
      RECT  98235.0 84505.0 98940.0 83160.0 ;
      RECT  98235.0 84505.0 98940.0 85850.0 ;
      RECT  98235.0 87195.0 98940.0 85850.0 ;
      RECT  98235.0 87195.0 98940.0 88540.0 ;
      RECT  98235.0 89885.0 98940.0 88540.0 ;
      RECT  98235.0 89885.0 98940.0 91230.0 ;
      RECT  98235.0 92575.0 98940.0 91230.0 ;
      RECT  98235.0 92575.0 98940.0 93920.0 ;
      RECT  98235.0 95265.0 98940.0 93920.0 ;
      RECT  98235.0 95265.0 98940.0 96610.0 ;
      RECT  98235.0 97955.0 98940.0 96610.0 ;
      RECT  98235.0 97955.0 98940.0 99300.0 ;
      RECT  98235.0 100645.0 98940.0 99300.0 ;
      RECT  98235.0 100645.0 98940.0 101990.0 ;
      RECT  98235.0 103335.0 98940.0 101990.0 ;
      RECT  98235.0 103335.0 98940.0 104680.0 ;
      RECT  98235.0 106025.0 98940.0 104680.0 ;
      RECT  98235.0 106025.0 98940.0 107370.0 ;
      RECT  98235.0 108715.0 98940.0 107370.0 ;
      RECT  98235.0 108715.0 98940.0 110060.0 ;
      RECT  98235.0 111405.0 98940.0 110060.0 ;
      RECT  98235.0 111405.0 98940.0 112750.0 ;
      RECT  98235.0 114095.0 98940.0 112750.0 ;
      RECT  98940.0 28015.0 99645.0 29360.0 ;
      RECT  98940.0 30705.0 99645.0 29360.0 ;
      RECT  98940.0 30705.0 99645.0 32050.0 ;
      RECT  98940.0 33395.0 99645.0 32050.0 ;
      RECT  98940.0 33395.0 99645.0 34740.0 ;
      RECT  98940.0 36085.0 99645.0 34740.0 ;
      RECT  98940.0 36085.0 99645.0 37430.0 ;
      RECT  98940.0 38775.0 99645.0 37430.0 ;
      RECT  98940.0 38775.0 99645.0 40120.0 ;
      RECT  98940.0 41465.0 99645.0 40120.0 ;
      RECT  98940.0 41465.0 99645.0 42810.0 ;
      RECT  98940.0 44155.0 99645.0 42810.0 ;
      RECT  98940.0 44155.0 99645.0 45500.0 ;
      RECT  98940.0 46845.0 99645.0 45500.0 ;
      RECT  98940.0 46845.0 99645.0 48190.0 ;
      RECT  98940.0 49535.0 99645.0 48190.0 ;
      RECT  98940.0 49535.0 99645.0 50880.0 ;
      RECT  98940.0 52225.0 99645.0 50880.0 ;
      RECT  98940.0 52225.0 99645.0 53570.0 ;
      RECT  98940.0 54915.0 99645.0 53570.0 ;
      RECT  98940.0 54915.0 99645.0 56260.0 ;
      RECT  98940.0 57605.0 99645.0 56260.0 ;
      RECT  98940.0 57605.0 99645.0 58950.0 ;
      RECT  98940.0 60295.0 99645.0 58950.0 ;
      RECT  98940.0 60295.0 99645.0 61640.0 ;
      RECT  98940.0 62985.0 99645.0 61640.0 ;
      RECT  98940.0 62985.0 99645.0 64330.0 ;
      RECT  98940.0 65675.0 99645.0 64330.0 ;
      RECT  98940.0 65675.0 99645.0 67020.0 ;
      RECT  98940.0 68365.0 99645.0 67020.0 ;
      RECT  98940.0 68365.0 99645.0 69710.0 ;
      RECT  98940.0 71055.0 99645.0 69710.0 ;
      RECT  98940.0 71055.0 99645.0 72400.0 ;
      RECT  98940.0 73745.0 99645.0 72400.0 ;
      RECT  98940.0 73745.0 99645.0 75090.0 ;
      RECT  98940.0 76435.0 99645.0 75090.0 ;
      RECT  98940.0 76435.0 99645.0 77780.0 ;
      RECT  98940.0 79125.0 99645.0 77780.0 ;
      RECT  98940.0 79125.0 99645.0 80470.0 ;
      RECT  98940.0 81815.0 99645.0 80470.0 ;
      RECT  98940.0 81815.0 99645.0 83160.0 ;
      RECT  98940.0 84505.0 99645.0 83160.0 ;
      RECT  98940.0 84505.0 99645.0 85850.0 ;
      RECT  98940.0 87195.0 99645.0 85850.0 ;
      RECT  98940.0 87195.0 99645.0 88540.0 ;
      RECT  98940.0 89885.0 99645.0 88540.0 ;
      RECT  98940.0 89885.0 99645.0 91230.0 ;
      RECT  98940.0 92575.0 99645.0 91230.0 ;
      RECT  98940.0 92575.0 99645.0 93920.0 ;
      RECT  98940.0 95265.0 99645.0 93920.0 ;
      RECT  98940.0 95265.0 99645.0 96610.0 ;
      RECT  98940.0 97955.0 99645.0 96610.0 ;
      RECT  98940.0 97955.0 99645.0 99300.0 ;
      RECT  98940.0 100645.0 99645.0 99300.0 ;
      RECT  98940.0 100645.0 99645.0 101990.0 ;
      RECT  98940.0 103335.0 99645.0 101990.0 ;
      RECT  98940.0 103335.0 99645.0 104680.0 ;
      RECT  98940.0 106025.0 99645.0 104680.0 ;
      RECT  98940.0 106025.0 99645.0 107370.0 ;
      RECT  98940.0 108715.0 99645.0 107370.0 ;
      RECT  98940.0 108715.0 99645.0 110060.0 ;
      RECT  98940.0 111405.0 99645.0 110060.0 ;
      RECT  98940.0 111405.0 99645.0 112750.0 ;
      RECT  98940.0 114095.0 99645.0 112750.0 ;
      RECT  99645.0 28015.0 100350.0 29360.0 ;
      RECT  99645.0 30705.0 100350.0 29360.0 ;
      RECT  99645.0 30705.0 100350.0 32050.0 ;
      RECT  99645.0 33395.0 100350.0 32050.0 ;
      RECT  99645.0 33395.0 100350.0 34740.0 ;
      RECT  99645.0 36085.0 100350.0 34740.0 ;
      RECT  99645.0 36085.0 100350.0 37430.0 ;
      RECT  99645.0 38775.0 100350.0 37430.0 ;
      RECT  99645.0 38775.0 100350.0 40120.0 ;
      RECT  99645.0 41465.0 100350.0 40120.0 ;
      RECT  99645.0 41465.0 100350.0 42810.0 ;
      RECT  99645.0 44155.0 100350.0 42810.0 ;
      RECT  99645.0 44155.0 100350.0 45500.0 ;
      RECT  99645.0 46845.0 100350.0 45500.0 ;
      RECT  99645.0 46845.0 100350.0 48190.0 ;
      RECT  99645.0 49535.0 100350.0 48190.0 ;
      RECT  99645.0 49535.0 100350.0 50880.0 ;
      RECT  99645.0 52225.0 100350.0 50880.0 ;
      RECT  99645.0 52225.0 100350.0 53570.0 ;
      RECT  99645.0 54915.0 100350.0 53570.0 ;
      RECT  99645.0 54915.0 100350.0 56260.0 ;
      RECT  99645.0 57605.0 100350.0 56260.0 ;
      RECT  99645.0 57605.0 100350.0 58950.0 ;
      RECT  99645.0 60295.0 100350.0 58950.0 ;
      RECT  99645.0 60295.0 100350.0 61640.0 ;
      RECT  99645.0 62985.0 100350.0 61640.0 ;
      RECT  99645.0 62985.0 100350.0 64330.0 ;
      RECT  99645.0 65675.0 100350.0 64330.0 ;
      RECT  99645.0 65675.0 100350.0 67020.0 ;
      RECT  99645.0 68365.0 100350.0 67020.0 ;
      RECT  99645.0 68365.0 100350.0 69710.0 ;
      RECT  99645.0 71055.0 100350.0 69710.0 ;
      RECT  99645.0 71055.0 100350.0 72400.0 ;
      RECT  99645.0 73745.0 100350.0 72400.0 ;
      RECT  99645.0 73745.0 100350.0 75090.0 ;
      RECT  99645.0 76435.0 100350.0 75090.0 ;
      RECT  99645.0 76435.0 100350.0 77780.0 ;
      RECT  99645.0 79125.0 100350.0 77780.0 ;
      RECT  99645.0 79125.0 100350.0 80470.0 ;
      RECT  99645.0 81815.0 100350.0 80470.0 ;
      RECT  99645.0 81815.0 100350.0 83160.0 ;
      RECT  99645.0 84505.0 100350.0 83160.0 ;
      RECT  99645.0 84505.0 100350.0 85850.0 ;
      RECT  99645.0 87195.0 100350.0 85850.0 ;
      RECT  99645.0 87195.0 100350.0 88540.0 ;
      RECT  99645.0 89885.0 100350.0 88540.0 ;
      RECT  99645.0 89885.0 100350.0 91230.0 ;
      RECT  99645.0 92575.0 100350.0 91230.0 ;
      RECT  99645.0 92575.0 100350.0 93920.0 ;
      RECT  99645.0 95265.0 100350.0 93920.0 ;
      RECT  99645.0 95265.0 100350.0 96610.0 ;
      RECT  99645.0 97955.0 100350.0 96610.0 ;
      RECT  99645.0 97955.0 100350.0 99300.0 ;
      RECT  99645.0 100645.0 100350.0 99300.0 ;
      RECT  99645.0 100645.0 100350.0 101990.0 ;
      RECT  99645.0 103335.0 100350.0 101990.0 ;
      RECT  99645.0 103335.0 100350.0 104680.0 ;
      RECT  99645.0 106025.0 100350.0 104680.0 ;
      RECT  99645.0 106025.0 100350.0 107370.0 ;
      RECT  99645.0 108715.0 100350.0 107370.0 ;
      RECT  99645.0 108715.0 100350.0 110060.0 ;
      RECT  99645.0 111405.0 100350.0 110060.0 ;
      RECT  99645.0 111405.0 100350.0 112750.0 ;
      RECT  99645.0 114095.0 100350.0 112750.0 ;
      RECT  100350.0 28015.0 101055.0 29360.0 ;
      RECT  100350.0 30705.0 101055.0 29360.0 ;
      RECT  100350.0 30705.0 101055.0 32050.0 ;
      RECT  100350.0 33395.0 101055.0 32050.0 ;
      RECT  100350.0 33395.0 101055.0 34740.0 ;
      RECT  100350.0 36085.0 101055.0 34740.0 ;
      RECT  100350.0 36085.0 101055.0 37430.0 ;
      RECT  100350.0 38775.0 101055.0 37430.0 ;
      RECT  100350.0 38775.0 101055.0 40120.0 ;
      RECT  100350.0 41465.0 101055.0 40120.0 ;
      RECT  100350.0 41465.0 101055.0 42810.0 ;
      RECT  100350.0 44155.0 101055.0 42810.0 ;
      RECT  100350.0 44155.0 101055.0 45500.0 ;
      RECT  100350.0 46845.0 101055.0 45500.0 ;
      RECT  100350.0 46845.0 101055.0 48190.0 ;
      RECT  100350.0 49535.0 101055.0 48190.0 ;
      RECT  100350.0 49535.0 101055.0 50880.0 ;
      RECT  100350.0 52225.0 101055.0 50880.0 ;
      RECT  100350.0 52225.0 101055.0 53570.0 ;
      RECT  100350.0 54915.0 101055.0 53570.0 ;
      RECT  100350.0 54915.0 101055.0 56260.0 ;
      RECT  100350.0 57605.0 101055.0 56260.0 ;
      RECT  100350.0 57605.0 101055.0 58950.0 ;
      RECT  100350.0 60295.0 101055.0 58950.0 ;
      RECT  100350.0 60295.0 101055.0 61640.0 ;
      RECT  100350.0 62985.0 101055.0 61640.0 ;
      RECT  100350.0 62985.0 101055.0 64330.0 ;
      RECT  100350.0 65675.0 101055.0 64330.0 ;
      RECT  100350.0 65675.0 101055.0 67020.0 ;
      RECT  100350.0 68365.0 101055.0 67020.0 ;
      RECT  100350.0 68365.0 101055.0 69710.0 ;
      RECT  100350.0 71055.0 101055.0 69710.0 ;
      RECT  100350.0 71055.0 101055.0 72400.0 ;
      RECT  100350.0 73745.0 101055.0 72400.0 ;
      RECT  100350.0 73745.0 101055.0 75090.0 ;
      RECT  100350.0 76435.0 101055.0 75090.0 ;
      RECT  100350.0 76435.0 101055.0 77780.0 ;
      RECT  100350.0 79125.0 101055.0 77780.0 ;
      RECT  100350.0 79125.0 101055.0 80470.0 ;
      RECT  100350.0 81815.0 101055.0 80470.0 ;
      RECT  100350.0 81815.0 101055.0 83160.0 ;
      RECT  100350.0 84505.0 101055.0 83160.0 ;
      RECT  100350.0 84505.0 101055.0 85850.0 ;
      RECT  100350.0 87195.0 101055.0 85850.0 ;
      RECT  100350.0 87195.0 101055.0 88540.0 ;
      RECT  100350.0 89885.0 101055.0 88540.0 ;
      RECT  100350.0 89885.0 101055.0 91230.0 ;
      RECT  100350.0 92575.0 101055.0 91230.0 ;
      RECT  100350.0 92575.0 101055.0 93920.0 ;
      RECT  100350.0 95265.0 101055.0 93920.0 ;
      RECT  100350.0 95265.0 101055.0 96610.0 ;
      RECT  100350.0 97955.0 101055.0 96610.0 ;
      RECT  100350.0 97955.0 101055.0 99300.0 ;
      RECT  100350.0 100645.0 101055.0 99300.0 ;
      RECT  100350.0 100645.0 101055.0 101990.0 ;
      RECT  100350.0 103335.0 101055.0 101990.0 ;
      RECT  100350.0 103335.0 101055.0 104680.0 ;
      RECT  100350.0 106025.0 101055.0 104680.0 ;
      RECT  100350.0 106025.0 101055.0 107370.0 ;
      RECT  100350.0 108715.0 101055.0 107370.0 ;
      RECT  100350.0 108715.0 101055.0 110060.0 ;
      RECT  100350.0 111405.0 101055.0 110060.0 ;
      RECT  100350.0 111405.0 101055.0 112750.0 ;
      RECT  100350.0 114095.0 101055.0 112750.0 ;
      RECT  101055.0 28015.0 101760.0 29360.0 ;
      RECT  101055.0 30705.0 101760.0 29360.0 ;
      RECT  101055.0 30705.0 101760.0 32050.0 ;
      RECT  101055.0 33395.0 101760.0 32050.0 ;
      RECT  101055.0 33395.0 101760.0 34740.0 ;
      RECT  101055.0 36085.0 101760.0 34740.0 ;
      RECT  101055.0 36085.0 101760.0 37430.0 ;
      RECT  101055.0 38775.0 101760.0 37430.0 ;
      RECT  101055.0 38775.0 101760.0 40120.0 ;
      RECT  101055.0 41465.0 101760.0 40120.0 ;
      RECT  101055.0 41465.0 101760.0 42810.0 ;
      RECT  101055.0 44155.0 101760.0 42810.0 ;
      RECT  101055.0 44155.0 101760.0 45500.0 ;
      RECT  101055.0 46845.0 101760.0 45500.0 ;
      RECT  101055.0 46845.0 101760.0 48190.0 ;
      RECT  101055.0 49535.0 101760.0 48190.0 ;
      RECT  101055.0 49535.0 101760.0 50880.0 ;
      RECT  101055.0 52225.0 101760.0 50880.0 ;
      RECT  101055.0 52225.0 101760.0 53570.0 ;
      RECT  101055.0 54915.0 101760.0 53570.0 ;
      RECT  101055.0 54915.0 101760.0 56260.0 ;
      RECT  101055.0 57605.0 101760.0 56260.0 ;
      RECT  101055.0 57605.0 101760.0 58950.0 ;
      RECT  101055.0 60295.0 101760.0 58950.0 ;
      RECT  101055.0 60295.0 101760.0 61640.0 ;
      RECT  101055.0 62985.0 101760.0 61640.0 ;
      RECT  101055.0 62985.0 101760.0 64330.0 ;
      RECT  101055.0 65675.0 101760.0 64330.0 ;
      RECT  101055.0 65675.0 101760.0 67020.0 ;
      RECT  101055.0 68365.0 101760.0 67020.0 ;
      RECT  101055.0 68365.0 101760.0 69710.0 ;
      RECT  101055.0 71055.0 101760.0 69710.0 ;
      RECT  101055.0 71055.0 101760.0 72400.0 ;
      RECT  101055.0 73745.0 101760.0 72400.0 ;
      RECT  101055.0 73745.0 101760.0 75090.0 ;
      RECT  101055.0 76435.0 101760.0 75090.0 ;
      RECT  101055.0 76435.0 101760.0 77780.0 ;
      RECT  101055.0 79125.0 101760.0 77780.0 ;
      RECT  101055.0 79125.0 101760.0 80470.0 ;
      RECT  101055.0 81815.0 101760.0 80470.0 ;
      RECT  101055.0 81815.0 101760.0 83160.0 ;
      RECT  101055.0 84505.0 101760.0 83160.0 ;
      RECT  101055.0 84505.0 101760.0 85850.0 ;
      RECT  101055.0 87195.0 101760.0 85850.0 ;
      RECT  101055.0 87195.0 101760.0 88540.0 ;
      RECT  101055.0 89885.0 101760.0 88540.0 ;
      RECT  101055.0 89885.0 101760.0 91230.0 ;
      RECT  101055.0 92575.0 101760.0 91230.0 ;
      RECT  101055.0 92575.0 101760.0 93920.0 ;
      RECT  101055.0 95265.0 101760.0 93920.0 ;
      RECT  101055.0 95265.0 101760.0 96610.0 ;
      RECT  101055.0 97955.0 101760.0 96610.0 ;
      RECT  101055.0 97955.0 101760.0 99300.0 ;
      RECT  101055.0 100645.0 101760.0 99300.0 ;
      RECT  101055.0 100645.0 101760.0 101990.0 ;
      RECT  101055.0 103335.0 101760.0 101990.0 ;
      RECT  101055.0 103335.0 101760.0 104680.0 ;
      RECT  101055.0 106025.0 101760.0 104680.0 ;
      RECT  101055.0 106025.0 101760.0 107370.0 ;
      RECT  101055.0 108715.0 101760.0 107370.0 ;
      RECT  101055.0 108715.0 101760.0 110060.0 ;
      RECT  101055.0 111405.0 101760.0 110060.0 ;
      RECT  101055.0 111405.0 101760.0 112750.0 ;
      RECT  101055.0 114095.0 101760.0 112750.0 ;
      RECT  101760.0 28015.0 102465.0 29360.0 ;
      RECT  101760.0 30705.0 102465.0 29360.0 ;
      RECT  101760.0 30705.0 102465.0 32050.0 ;
      RECT  101760.0 33395.0 102465.0 32050.0 ;
      RECT  101760.0 33395.0 102465.0 34740.0 ;
      RECT  101760.0 36085.0 102465.0 34740.0 ;
      RECT  101760.0 36085.0 102465.0 37430.0 ;
      RECT  101760.0 38775.0 102465.0 37430.0 ;
      RECT  101760.0 38775.0 102465.0 40120.0 ;
      RECT  101760.0 41465.0 102465.0 40120.0 ;
      RECT  101760.0 41465.0 102465.0 42810.0 ;
      RECT  101760.0 44155.0 102465.0 42810.0 ;
      RECT  101760.0 44155.0 102465.0 45500.0 ;
      RECT  101760.0 46845.0 102465.0 45500.0 ;
      RECT  101760.0 46845.0 102465.0 48190.0 ;
      RECT  101760.0 49535.0 102465.0 48190.0 ;
      RECT  101760.0 49535.0 102465.0 50880.0 ;
      RECT  101760.0 52225.0 102465.0 50880.0 ;
      RECT  101760.0 52225.0 102465.0 53570.0 ;
      RECT  101760.0 54915.0 102465.0 53570.0 ;
      RECT  101760.0 54915.0 102465.0 56260.0 ;
      RECT  101760.0 57605.0 102465.0 56260.0 ;
      RECT  101760.0 57605.0 102465.0 58950.0 ;
      RECT  101760.0 60295.0 102465.0 58950.0 ;
      RECT  101760.0 60295.0 102465.0 61640.0 ;
      RECT  101760.0 62985.0 102465.0 61640.0 ;
      RECT  101760.0 62985.0 102465.0 64330.0 ;
      RECT  101760.0 65675.0 102465.0 64330.0 ;
      RECT  101760.0 65675.0 102465.0 67020.0 ;
      RECT  101760.0 68365.0 102465.0 67020.0 ;
      RECT  101760.0 68365.0 102465.0 69710.0 ;
      RECT  101760.0 71055.0 102465.0 69710.0 ;
      RECT  101760.0 71055.0 102465.0 72400.0 ;
      RECT  101760.0 73745.0 102465.0 72400.0 ;
      RECT  101760.0 73745.0 102465.0 75090.0 ;
      RECT  101760.0 76435.0 102465.0 75090.0 ;
      RECT  101760.0 76435.0 102465.0 77780.0 ;
      RECT  101760.0 79125.0 102465.0 77780.0 ;
      RECT  101760.0 79125.0 102465.0 80470.0 ;
      RECT  101760.0 81815.0 102465.0 80470.0 ;
      RECT  101760.0 81815.0 102465.0 83160.0 ;
      RECT  101760.0 84505.0 102465.0 83160.0 ;
      RECT  101760.0 84505.0 102465.0 85850.0 ;
      RECT  101760.0 87195.0 102465.0 85850.0 ;
      RECT  101760.0 87195.0 102465.0 88540.0 ;
      RECT  101760.0 89885.0 102465.0 88540.0 ;
      RECT  101760.0 89885.0 102465.0 91230.0 ;
      RECT  101760.0 92575.0 102465.0 91230.0 ;
      RECT  101760.0 92575.0 102465.0 93920.0 ;
      RECT  101760.0 95265.0 102465.0 93920.0 ;
      RECT  101760.0 95265.0 102465.0 96610.0 ;
      RECT  101760.0 97955.0 102465.0 96610.0 ;
      RECT  101760.0 97955.0 102465.0 99300.0 ;
      RECT  101760.0 100645.0 102465.0 99300.0 ;
      RECT  101760.0 100645.0 102465.0 101990.0 ;
      RECT  101760.0 103335.0 102465.0 101990.0 ;
      RECT  101760.0 103335.0 102465.0 104680.0 ;
      RECT  101760.0 106025.0 102465.0 104680.0 ;
      RECT  101760.0 106025.0 102465.0 107370.0 ;
      RECT  101760.0 108715.0 102465.0 107370.0 ;
      RECT  101760.0 108715.0 102465.0 110060.0 ;
      RECT  101760.0 111405.0 102465.0 110060.0 ;
      RECT  101760.0 111405.0 102465.0 112750.0 ;
      RECT  101760.0 114095.0 102465.0 112750.0 ;
      RECT  102465.0 28015.0 103170.0 29360.0 ;
      RECT  102465.0 30705.0 103170.0 29360.0 ;
      RECT  102465.0 30705.0 103170.0 32050.0 ;
      RECT  102465.0 33395.0 103170.0 32050.0 ;
      RECT  102465.0 33395.0 103170.0 34740.0 ;
      RECT  102465.0 36085.0 103170.0 34740.0 ;
      RECT  102465.0 36085.0 103170.0 37430.0 ;
      RECT  102465.0 38775.0 103170.0 37430.0 ;
      RECT  102465.0 38775.0 103170.0 40120.0 ;
      RECT  102465.0 41465.0 103170.0 40120.0 ;
      RECT  102465.0 41465.0 103170.0 42810.0 ;
      RECT  102465.0 44155.0 103170.0 42810.0 ;
      RECT  102465.0 44155.0 103170.0 45500.0 ;
      RECT  102465.0 46845.0 103170.0 45500.0 ;
      RECT  102465.0 46845.0 103170.0 48190.0 ;
      RECT  102465.0 49535.0 103170.0 48190.0 ;
      RECT  102465.0 49535.0 103170.0 50880.0 ;
      RECT  102465.0 52225.0 103170.0 50880.0 ;
      RECT  102465.0 52225.0 103170.0 53570.0 ;
      RECT  102465.0 54915.0 103170.0 53570.0 ;
      RECT  102465.0 54915.0 103170.0 56260.0 ;
      RECT  102465.0 57605.0 103170.0 56260.0 ;
      RECT  102465.0 57605.0 103170.0 58950.0 ;
      RECT  102465.0 60295.0 103170.0 58950.0 ;
      RECT  102465.0 60295.0 103170.0 61640.0 ;
      RECT  102465.0 62985.0 103170.0 61640.0 ;
      RECT  102465.0 62985.0 103170.0 64330.0 ;
      RECT  102465.0 65675.0 103170.0 64330.0 ;
      RECT  102465.0 65675.0 103170.0 67020.0 ;
      RECT  102465.0 68365.0 103170.0 67020.0 ;
      RECT  102465.0 68365.0 103170.0 69710.0 ;
      RECT  102465.0 71055.0 103170.0 69710.0 ;
      RECT  102465.0 71055.0 103170.0 72400.0 ;
      RECT  102465.0 73745.0 103170.0 72400.0 ;
      RECT  102465.0 73745.0 103170.0 75090.0 ;
      RECT  102465.0 76435.0 103170.0 75090.0 ;
      RECT  102465.0 76435.0 103170.0 77780.0 ;
      RECT  102465.0 79125.0 103170.0 77780.0 ;
      RECT  102465.0 79125.0 103170.0 80470.0 ;
      RECT  102465.0 81815.0 103170.0 80470.0 ;
      RECT  102465.0 81815.0 103170.0 83160.0 ;
      RECT  102465.0 84505.0 103170.0 83160.0 ;
      RECT  102465.0 84505.0 103170.0 85850.0 ;
      RECT  102465.0 87195.0 103170.0 85850.0 ;
      RECT  102465.0 87195.0 103170.0 88540.0 ;
      RECT  102465.0 89885.0 103170.0 88540.0 ;
      RECT  102465.0 89885.0 103170.0 91230.0 ;
      RECT  102465.0 92575.0 103170.0 91230.0 ;
      RECT  102465.0 92575.0 103170.0 93920.0 ;
      RECT  102465.0 95265.0 103170.0 93920.0 ;
      RECT  102465.0 95265.0 103170.0 96610.0 ;
      RECT  102465.0 97955.0 103170.0 96610.0 ;
      RECT  102465.0 97955.0 103170.0 99300.0 ;
      RECT  102465.0 100645.0 103170.0 99300.0 ;
      RECT  102465.0 100645.0 103170.0 101990.0 ;
      RECT  102465.0 103335.0 103170.0 101990.0 ;
      RECT  102465.0 103335.0 103170.0 104680.0 ;
      RECT  102465.0 106025.0 103170.0 104680.0 ;
      RECT  102465.0 106025.0 103170.0 107370.0 ;
      RECT  102465.0 108715.0 103170.0 107370.0 ;
      RECT  102465.0 108715.0 103170.0 110060.0 ;
      RECT  102465.0 111405.0 103170.0 110060.0 ;
      RECT  102465.0 111405.0 103170.0 112750.0 ;
      RECT  102465.0 114095.0 103170.0 112750.0 ;
      RECT  103170.0 28015.0 103875.0 29360.0 ;
      RECT  103170.0 30705.0 103875.0 29360.0 ;
      RECT  103170.0 30705.0 103875.0 32050.0 ;
      RECT  103170.0 33395.0 103875.0 32050.0 ;
      RECT  103170.0 33395.0 103875.0 34740.0 ;
      RECT  103170.0 36085.0 103875.0 34740.0 ;
      RECT  103170.0 36085.0 103875.0 37430.0 ;
      RECT  103170.0 38775.0 103875.0 37430.0 ;
      RECT  103170.0 38775.0 103875.0 40120.0 ;
      RECT  103170.0 41465.0 103875.0 40120.0 ;
      RECT  103170.0 41465.0 103875.0 42810.0 ;
      RECT  103170.0 44155.0 103875.0 42810.0 ;
      RECT  103170.0 44155.0 103875.0 45500.0 ;
      RECT  103170.0 46845.0 103875.0 45500.0 ;
      RECT  103170.0 46845.0 103875.0 48190.0 ;
      RECT  103170.0 49535.0 103875.0 48190.0 ;
      RECT  103170.0 49535.0 103875.0 50880.0 ;
      RECT  103170.0 52225.0 103875.0 50880.0 ;
      RECT  103170.0 52225.0 103875.0 53570.0 ;
      RECT  103170.0 54915.0 103875.0 53570.0 ;
      RECT  103170.0 54915.0 103875.0 56260.0 ;
      RECT  103170.0 57605.0 103875.0 56260.0 ;
      RECT  103170.0 57605.0 103875.0 58950.0 ;
      RECT  103170.0 60295.0 103875.0 58950.0 ;
      RECT  103170.0 60295.0 103875.0 61640.0 ;
      RECT  103170.0 62985.0 103875.0 61640.0 ;
      RECT  103170.0 62985.0 103875.0 64330.0 ;
      RECT  103170.0 65675.0 103875.0 64330.0 ;
      RECT  103170.0 65675.0 103875.0 67020.0 ;
      RECT  103170.0 68365.0 103875.0 67020.0 ;
      RECT  103170.0 68365.0 103875.0 69710.0 ;
      RECT  103170.0 71055.0 103875.0 69710.0 ;
      RECT  103170.0 71055.0 103875.0 72400.0 ;
      RECT  103170.0 73745.0 103875.0 72400.0 ;
      RECT  103170.0 73745.0 103875.0 75090.0 ;
      RECT  103170.0 76435.0 103875.0 75090.0 ;
      RECT  103170.0 76435.0 103875.0 77780.0 ;
      RECT  103170.0 79125.0 103875.0 77780.0 ;
      RECT  103170.0 79125.0 103875.0 80470.0 ;
      RECT  103170.0 81815.0 103875.0 80470.0 ;
      RECT  103170.0 81815.0 103875.0 83160.0 ;
      RECT  103170.0 84505.0 103875.0 83160.0 ;
      RECT  103170.0 84505.0 103875.0 85850.0 ;
      RECT  103170.0 87195.0 103875.0 85850.0 ;
      RECT  103170.0 87195.0 103875.0 88540.0 ;
      RECT  103170.0 89885.0 103875.0 88540.0 ;
      RECT  103170.0 89885.0 103875.0 91230.0 ;
      RECT  103170.0 92575.0 103875.0 91230.0 ;
      RECT  103170.0 92575.0 103875.0 93920.0 ;
      RECT  103170.0 95265.0 103875.0 93920.0 ;
      RECT  103170.0 95265.0 103875.0 96610.0 ;
      RECT  103170.0 97955.0 103875.0 96610.0 ;
      RECT  103170.0 97955.0 103875.0 99300.0 ;
      RECT  103170.0 100645.0 103875.0 99300.0 ;
      RECT  103170.0 100645.0 103875.0 101990.0 ;
      RECT  103170.0 103335.0 103875.0 101990.0 ;
      RECT  103170.0 103335.0 103875.0 104680.0 ;
      RECT  103170.0 106025.0 103875.0 104680.0 ;
      RECT  103170.0 106025.0 103875.0 107370.0 ;
      RECT  103170.0 108715.0 103875.0 107370.0 ;
      RECT  103170.0 108715.0 103875.0 110060.0 ;
      RECT  103170.0 111405.0 103875.0 110060.0 ;
      RECT  103170.0 111405.0 103875.0 112750.0 ;
      RECT  103170.0 114095.0 103875.0 112750.0 ;
      RECT  103875.0 28015.0 104580.0 29360.0 ;
      RECT  103875.0 30705.0 104580.0 29360.0 ;
      RECT  103875.0 30705.0 104580.0 32050.0 ;
      RECT  103875.0 33395.0 104580.0 32050.0 ;
      RECT  103875.0 33395.0 104580.0 34740.0 ;
      RECT  103875.0 36085.0 104580.0 34740.0 ;
      RECT  103875.0 36085.0 104580.0 37430.0 ;
      RECT  103875.0 38775.0 104580.0 37430.0 ;
      RECT  103875.0 38775.0 104580.0 40120.0 ;
      RECT  103875.0 41465.0 104580.0 40120.0 ;
      RECT  103875.0 41465.0 104580.0 42810.0 ;
      RECT  103875.0 44155.0 104580.0 42810.0 ;
      RECT  103875.0 44155.0 104580.0 45500.0 ;
      RECT  103875.0 46845.0 104580.0 45500.0 ;
      RECT  103875.0 46845.0 104580.0 48190.0 ;
      RECT  103875.0 49535.0 104580.0 48190.0 ;
      RECT  103875.0 49535.0 104580.0 50880.0 ;
      RECT  103875.0 52225.0 104580.0 50880.0 ;
      RECT  103875.0 52225.0 104580.0 53570.0 ;
      RECT  103875.0 54915.0 104580.0 53570.0 ;
      RECT  103875.0 54915.0 104580.0 56260.0 ;
      RECT  103875.0 57605.0 104580.0 56260.0 ;
      RECT  103875.0 57605.0 104580.0 58950.0 ;
      RECT  103875.0 60295.0 104580.0 58950.0 ;
      RECT  103875.0 60295.0 104580.0 61640.0 ;
      RECT  103875.0 62985.0 104580.0 61640.0 ;
      RECT  103875.0 62985.0 104580.0 64330.0 ;
      RECT  103875.0 65675.0 104580.0 64330.0 ;
      RECT  103875.0 65675.0 104580.0 67020.0 ;
      RECT  103875.0 68365.0 104580.0 67020.0 ;
      RECT  103875.0 68365.0 104580.0 69710.0 ;
      RECT  103875.0 71055.0 104580.0 69710.0 ;
      RECT  103875.0 71055.0 104580.0 72400.0 ;
      RECT  103875.0 73745.0 104580.0 72400.0 ;
      RECT  103875.0 73745.0 104580.0 75090.0 ;
      RECT  103875.0 76435.0 104580.0 75090.0 ;
      RECT  103875.0 76435.0 104580.0 77780.0 ;
      RECT  103875.0 79125.0 104580.0 77780.0 ;
      RECT  103875.0 79125.0 104580.0 80470.0 ;
      RECT  103875.0 81815.0 104580.0 80470.0 ;
      RECT  103875.0 81815.0 104580.0 83160.0 ;
      RECT  103875.0 84505.0 104580.0 83160.0 ;
      RECT  103875.0 84505.0 104580.0 85850.0 ;
      RECT  103875.0 87195.0 104580.0 85850.0 ;
      RECT  103875.0 87195.0 104580.0 88540.0 ;
      RECT  103875.0 89885.0 104580.0 88540.0 ;
      RECT  103875.0 89885.0 104580.0 91230.0 ;
      RECT  103875.0 92575.0 104580.0 91230.0 ;
      RECT  103875.0 92575.0 104580.0 93920.0 ;
      RECT  103875.0 95265.0 104580.0 93920.0 ;
      RECT  103875.0 95265.0 104580.0 96610.0 ;
      RECT  103875.0 97955.0 104580.0 96610.0 ;
      RECT  103875.0 97955.0 104580.0 99300.0 ;
      RECT  103875.0 100645.0 104580.0 99300.0 ;
      RECT  103875.0 100645.0 104580.0 101990.0 ;
      RECT  103875.0 103335.0 104580.0 101990.0 ;
      RECT  103875.0 103335.0 104580.0 104680.0 ;
      RECT  103875.0 106025.0 104580.0 104680.0 ;
      RECT  103875.0 106025.0 104580.0 107370.0 ;
      RECT  103875.0 108715.0 104580.0 107370.0 ;
      RECT  103875.0 108715.0 104580.0 110060.0 ;
      RECT  103875.0 111405.0 104580.0 110060.0 ;
      RECT  103875.0 111405.0 104580.0 112750.0 ;
      RECT  103875.0 114095.0 104580.0 112750.0 ;
      RECT  104580.0 28015.0 105285.0 29360.0 ;
      RECT  104580.0 30705.0 105285.0 29360.0 ;
      RECT  104580.0 30705.0 105285.0 32050.0 ;
      RECT  104580.0 33395.0 105285.0 32050.0 ;
      RECT  104580.0 33395.0 105285.0 34740.0 ;
      RECT  104580.0 36085.0 105285.0 34740.0 ;
      RECT  104580.0 36085.0 105285.0 37430.0 ;
      RECT  104580.0 38775.0 105285.0 37430.0 ;
      RECT  104580.0 38775.0 105285.0 40120.0 ;
      RECT  104580.0 41465.0 105285.0 40120.0 ;
      RECT  104580.0 41465.0 105285.0 42810.0 ;
      RECT  104580.0 44155.0 105285.0 42810.0 ;
      RECT  104580.0 44155.0 105285.0 45500.0 ;
      RECT  104580.0 46845.0 105285.0 45500.0 ;
      RECT  104580.0 46845.0 105285.0 48190.0 ;
      RECT  104580.0 49535.0 105285.0 48190.0 ;
      RECT  104580.0 49535.0 105285.0 50880.0 ;
      RECT  104580.0 52225.0 105285.0 50880.0 ;
      RECT  104580.0 52225.0 105285.0 53570.0 ;
      RECT  104580.0 54915.0 105285.0 53570.0 ;
      RECT  104580.0 54915.0 105285.0 56260.0 ;
      RECT  104580.0 57605.0 105285.0 56260.0 ;
      RECT  104580.0 57605.0 105285.0 58950.0 ;
      RECT  104580.0 60295.0 105285.0 58950.0 ;
      RECT  104580.0 60295.0 105285.0 61640.0 ;
      RECT  104580.0 62985.0 105285.0 61640.0 ;
      RECT  104580.0 62985.0 105285.0 64330.0 ;
      RECT  104580.0 65675.0 105285.0 64330.0 ;
      RECT  104580.0 65675.0 105285.0 67020.0 ;
      RECT  104580.0 68365.0 105285.0 67020.0 ;
      RECT  104580.0 68365.0 105285.0 69710.0 ;
      RECT  104580.0 71055.0 105285.0 69710.0 ;
      RECT  104580.0 71055.0 105285.0 72400.0 ;
      RECT  104580.0 73745.0 105285.0 72400.0 ;
      RECT  104580.0 73745.0 105285.0 75090.0 ;
      RECT  104580.0 76435.0 105285.0 75090.0 ;
      RECT  104580.0 76435.0 105285.0 77780.0 ;
      RECT  104580.0 79125.0 105285.0 77780.0 ;
      RECT  104580.0 79125.0 105285.0 80470.0 ;
      RECT  104580.0 81815.0 105285.0 80470.0 ;
      RECT  104580.0 81815.0 105285.0 83160.0 ;
      RECT  104580.0 84505.0 105285.0 83160.0 ;
      RECT  104580.0 84505.0 105285.0 85850.0 ;
      RECT  104580.0 87195.0 105285.0 85850.0 ;
      RECT  104580.0 87195.0 105285.0 88540.0 ;
      RECT  104580.0 89885.0 105285.0 88540.0 ;
      RECT  104580.0 89885.0 105285.0 91230.0 ;
      RECT  104580.0 92575.0 105285.0 91230.0 ;
      RECT  104580.0 92575.0 105285.0 93920.0 ;
      RECT  104580.0 95265.0 105285.0 93920.0 ;
      RECT  104580.0 95265.0 105285.0 96610.0 ;
      RECT  104580.0 97955.0 105285.0 96610.0 ;
      RECT  104580.0 97955.0 105285.0 99300.0 ;
      RECT  104580.0 100645.0 105285.0 99300.0 ;
      RECT  104580.0 100645.0 105285.0 101990.0 ;
      RECT  104580.0 103335.0 105285.0 101990.0 ;
      RECT  104580.0 103335.0 105285.0 104680.0 ;
      RECT  104580.0 106025.0 105285.0 104680.0 ;
      RECT  104580.0 106025.0 105285.0 107370.0 ;
      RECT  104580.0 108715.0 105285.0 107370.0 ;
      RECT  104580.0 108715.0 105285.0 110060.0 ;
      RECT  104580.0 111405.0 105285.0 110060.0 ;
      RECT  104580.0 111405.0 105285.0 112750.0 ;
      RECT  104580.0 114095.0 105285.0 112750.0 ;
      RECT  105285.0 28015.0 105990.0 29360.0 ;
      RECT  105285.0 30705.0 105990.0 29360.0 ;
      RECT  105285.0 30705.0 105990.0 32050.0 ;
      RECT  105285.0 33395.0 105990.0 32050.0 ;
      RECT  105285.0 33395.0 105990.0 34740.0 ;
      RECT  105285.0 36085.0 105990.0 34740.0 ;
      RECT  105285.0 36085.0 105990.0 37430.0 ;
      RECT  105285.0 38775.0 105990.0 37430.0 ;
      RECT  105285.0 38775.0 105990.0 40120.0 ;
      RECT  105285.0 41465.0 105990.0 40120.0 ;
      RECT  105285.0 41465.0 105990.0 42810.0 ;
      RECT  105285.0 44155.0 105990.0 42810.0 ;
      RECT  105285.0 44155.0 105990.0 45500.0 ;
      RECT  105285.0 46845.0 105990.0 45500.0 ;
      RECT  105285.0 46845.0 105990.0 48190.0 ;
      RECT  105285.0 49535.0 105990.0 48190.0 ;
      RECT  105285.0 49535.0 105990.0 50880.0 ;
      RECT  105285.0 52225.0 105990.0 50880.0 ;
      RECT  105285.0 52225.0 105990.0 53570.0 ;
      RECT  105285.0 54915.0 105990.0 53570.0 ;
      RECT  105285.0 54915.0 105990.0 56260.0 ;
      RECT  105285.0 57605.0 105990.0 56260.0 ;
      RECT  105285.0 57605.0 105990.0 58950.0 ;
      RECT  105285.0 60295.0 105990.0 58950.0 ;
      RECT  105285.0 60295.0 105990.0 61640.0 ;
      RECT  105285.0 62985.0 105990.0 61640.0 ;
      RECT  105285.0 62985.0 105990.0 64330.0 ;
      RECT  105285.0 65675.0 105990.0 64330.0 ;
      RECT  105285.0 65675.0 105990.0 67020.0 ;
      RECT  105285.0 68365.0 105990.0 67020.0 ;
      RECT  105285.0 68365.0 105990.0 69710.0 ;
      RECT  105285.0 71055.0 105990.0 69710.0 ;
      RECT  105285.0 71055.0 105990.0 72400.0 ;
      RECT  105285.0 73745.0 105990.0 72400.0 ;
      RECT  105285.0 73745.0 105990.0 75090.0 ;
      RECT  105285.0 76435.0 105990.0 75090.0 ;
      RECT  105285.0 76435.0 105990.0 77780.0 ;
      RECT  105285.0 79125.0 105990.0 77780.0 ;
      RECT  105285.0 79125.0 105990.0 80470.0 ;
      RECT  105285.0 81815.0 105990.0 80470.0 ;
      RECT  105285.0 81815.0 105990.0 83160.0 ;
      RECT  105285.0 84505.0 105990.0 83160.0 ;
      RECT  105285.0 84505.0 105990.0 85850.0 ;
      RECT  105285.0 87195.0 105990.0 85850.0 ;
      RECT  105285.0 87195.0 105990.0 88540.0 ;
      RECT  105285.0 89885.0 105990.0 88540.0 ;
      RECT  105285.0 89885.0 105990.0 91230.0 ;
      RECT  105285.0 92575.0 105990.0 91230.0 ;
      RECT  105285.0 92575.0 105990.0 93920.0 ;
      RECT  105285.0 95265.0 105990.0 93920.0 ;
      RECT  105285.0 95265.0 105990.0 96610.0 ;
      RECT  105285.0 97955.0 105990.0 96610.0 ;
      RECT  105285.0 97955.0 105990.0 99300.0 ;
      RECT  105285.0 100645.0 105990.0 99300.0 ;
      RECT  105285.0 100645.0 105990.0 101990.0 ;
      RECT  105285.0 103335.0 105990.0 101990.0 ;
      RECT  105285.0 103335.0 105990.0 104680.0 ;
      RECT  105285.0 106025.0 105990.0 104680.0 ;
      RECT  105285.0 106025.0 105990.0 107370.0 ;
      RECT  105285.0 108715.0 105990.0 107370.0 ;
      RECT  105285.0 108715.0 105990.0 110060.0 ;
      RECT  105285.0 111405.0 105990.0 110060.0 ;
      RECT  105285.0 111405.0 105990.0 112750.0 ;
      RECT  105285.0 114095.0 105990.0 112750.0 ;
      RECT  15900.0 27915.0 15970.0 114250.0 ;
      RECT  16235.0 27915.0 16305.0 114250.0 ;
      RECT  16605.0 27915.0 16675.0 114250.0 ;
      RECT  16940.0 27915.0 17010.0 114250.0 ;
      RECT  17310.0 27915.0 17380.0 114250.0 ;
      RECT  17645.0 27915.0 17715.0 114250.0 ;
      RECT  18015.0 27915.0 18085.0 114250.0 ;
      RECT  18350.0 27915.0 18420.0 114250.0 ;
      RECT  18720.0 27915.0 18790.0 114250.0 ;
      RECT  19055.0 27915.0 19125.0 114250.0 ;
      RECT  19425.0 27915.0 19495.0 114250.0 ;
      RECT  19760.0 27915.0 19830.0 114250.0 ;
      RECT  20130.0 27915.0 20200.0 114250.0 ;
      RECT  20465.0 27915.0 20535.0 114250.0 ;
      RECT  20835.0 27915.0 20905.0 114250.0 ;
      RECT  21170.0 27915.0 21240.0 114250.0 ;
      RECT  21540.0 27915.0 21610.0 114250.0 ;
      RECT  21875.0 27915.0 21945.0 114250.0 ;
      RECT  22245.0 27915.0 22315.0 114250.0 ;
      RECT  22580.0 27915.0 22650.0 114250.0 ;
      RECT  22950.0 27915.0 23020.0 114250.0 ;
      RECT  23285.0 27915.0 23355.0 114250.0 ;
      RECT  23655.0 27915.0 23725.0 114250.0 ;
      RECT  23990.0 27915.0 24060.0 114250.0 ;
      RECT  24360.0 27915.0 24430.0 114250.0 ;
      RECT  24695.0 27915.0 24765.0 114250.0 ;
      RECT  25065.0 27915.0 25135.0 114250.0 ;
      RECT  25400.0 27915.0 25470.0 114250.0 ;
      RECT  25770.0 27915.0 25840.0 114250.0 ;
      RECT  26105.0 27915.0 26175.0 114250.0 ;
      RECT  26475.0 27915.0 26545.0 114250.0 ;
      RECT  26810.0 27915.0 26880.0 114250.0 ;
      RECT  27180.0 27915.0 27250.0 114250.0 ;
      RECT  27515.0 27915.0 27585.0 114250.0 ;
      RECT  27885.0 27915.0 27955.0 114250.0 ;
      RECT  28220.0 27915.0 28290.0 114250.0 ;
      RECT  28590.0 27915.0 28660.0 114250.0 ;
      RECT  28925.0 27915.0 28995.0 114250.0 ;
      RECT  29295.0 27915.0 29365.0 114250.0 ;
      RECT  29630.0 27915.0 29700.0 114250.0 ;
      RECT  30000.0 27915.0 30070.0 114250.0 ;
      RECT  30335.0 27915.0 30405.0 114250.0 ;
      RECT  30705.0 27915.0 30775.0 114250.0 ;
      RECT  31040.0 27915.0 31110.0 114250.0 ;
      RECT  31410.0 27915.0 31480.0 114250.0 ;
      RECT  31745.0 27915.0 31815.0 114250.0 ;
      RECT  32115.0 27915.0 32185.0 114250.0 ;
      RECT  32450.0 27915.0 32520.0 114250.0 ;
      RECT  32820.0 27915.0 32890.0 114250.0 ;
      RECT  33155.0 27915.0 33225.0 114250.0 ;
      RECT  33525.0 27915.0 33595.0 114250.0 ;
      RECT  33860.0 27915.0 33930.0 114250.0 ;
      RECT  34230.0 27915.0 34300.0 114250.0 ;
      RECT  34565.0 27915.0 34635.0 114250.0 ;
      RECT  34935.0 27915.0 35005.0 114250.0 ;
      RECT  35270.0 27915.0 35340.0 114250.0 ;
      RECT  35640.0 27915.0 35710.0 114250.0 ;
      RECT  35975.0 27915.0 36045.0 114250.0 ;
      RECT  36345.0 27915.0 36415.0 114250.0 ;
      RECT  36680.0 27915.0 36750.0 114250.0 ;
      RECT  37050.0 27915.0 37120.0 114250.0 ;
      RECT  37385.0 27915.0 37455.0 114250.0 ;
      RECT  37755.0 27915.0 37825.0 114250.0 ;
      RECT  38090.0 27915.0 38160.0 114250.0 ;
      RECT  38460.0 27915.0 38530.0 114250.0 ;
      RECT  38795.0 27915.0 38865.0 114250.0 ;
      RECT  39165.0 27915.0 39235.0 114250.0 ;
      RECT  39500.0 27915.0 39570.0 114250.0 ;
      RECT  39870.0 27915.0 39940.0 114250.0 ;
      RECT  40205.0 27915.0 40275.0 114250.0 ;
      RECT  40575.0 27915.0 40645.0 114250.0 ;
      RECT  40910.0 27915.0 40980.0 114250.0 ;
      RECT  41280.0 27915.0 41350.0 114250.0 ;
      RECT  41615.0 27915.0 41685.0 114250.0 ;
      RECT  41985.0 27915.0 42055.0 114250.0 ;
      RECT  42320.0 27915.0 42390.0 114250.0 ;
      RECT  42690.0 27915.0 42760.0 114250.0 ;
      RECT  43025.0 27915.0 43095.0 114250.0 ;
      RECT  43395.0 27915.0 43465.0 114250.0 ;
      RECT  43730.0 27915.0 43800.0 114250.0 ;
      RECT  44100.0 27915.0 44170.0 114250.0 ;
      RECT  44435.0 27915.0 44505.0 114250.0 ;
      RECT  44805.0 27915.0 44875.0 114250.0 ;
      RECT  45140.0 27915.0 45210.0 114250.0 ;
      RECT  45510.0 27915.0 45580.0 114250.0 ;
      RECT  45845.0 27915.0 45915.0 114250.0 ;
      RECT  46215.0 27915.0 46285.0 114250.0 ;
      RECT  46550.0 27915.0 46620.0 114250.0 ;
      RECT  46920.0 27915.0 46990.0 114250.0 ;
      RECT  47255.0 27915.0 47325.0 114250.0 ;
      RECT  47625.0 27915.0 47695.0 114250.0 ;
      RECT  47960.0 27915.0 48030.0 114250.0 ;
      RECT  48330.0 27915.0 48400.0 114250.0 ;
      RECT  48665.0 27915.0 48735.0 114250.0 ;
      RECT  49035.0 27915.0 49105.0 114250.0 ;
      RECT  49370.0 27915.0 49440.0 114250.0 ;
      RECT  49740.0 27915.0 49810.0 114250.0 ;
      RECT  50075.0 27915.0 50145.0 114250.0 ;
      RECT  50445.0 27915.0 50515.0 114250.0 ;
      RECT  50780.0 27915.0 50850.0 114250.0 ;
      RECT  51150.0 27915.0 51220.0 114250.0 ;
      RECT  51485.0 27915.0 51555.0 114250.0 ;
      RECT  51855.0 27915.0 51925.0 114250.0 ;
      RECT  52190.0 27915.0 52260.0 114250.0 ;
      RECT  52560.0 27915.0 52630.0 114250.0 ;
      RECT  52895.0 27915.0 52965.0 114250.0 ;
      RECT  53265.0 27915.0 53335.0 114250.0 ;
      RECT  53600.0 27915.0 53670.0 114250.0 ;
      RECT  53970.0 27915.0 54040.0 114250.0 ;
      RECT  54305.0 27915.0 54375.0 114250.0 ;
      RECT  54675.0 27915.0 54745.0 114250.0 ;
      RECT  55010.0 27915.0 55080.0 114250.0 ;
      RECT  55380.0 27915.0 55450.0 114250.0 ;
      RECT  55715.0 27915.0 55785.0 114250.0 ;
      RECT  56085.0 27915.0 56155.0 114250.0 ;
      RECT  56420.0 27915.0 56490.0 114250.0 ;
      RECT  56790.0 27915.0 56860.0 114250.0 ;
      RECT  57125.0 27915.0 57195.0 114250.0 ;
      RECT  57495.0 27915.0 57565.0 114250.0 ;
      RECT  57830.0 27915.0 57900.0 114250.0 ;
      RECT  58200.0 27915.0 58270.0 114250.0 ;
      RECT  58535.0 27915.0 58605.0 114250.0 ;
      RECT  58905.0 27915.0 58975.0 114250.0 ;
      RECT  59240.0 27915.0 59310.0 114250.0 ;
      RECT  59610.0 27915.0 59680.0 114250.0 ;
      RECT  59945.0 27915.0 60015.0 114250.0 ;
      RECT  60315.0 27915.0 60385.0 114250.0 ;
      RECT  60650.0 27915.0 60720.0 114250.0 ;
      RECT  61020.0 27915.0 61090.0 114250.0 ;
      RECT  61355.0 27915.0 61425.0 114250.0 ;
      RECT  61725.0 27915.0 61795.0 114250.0 ;
      RECT  62060.0 27915.0 62130.0 114250.0 ;
      RECT  62430.0 27915.0 62500.0 114250.0 ;
      RECT  62765.0 27915.0 62835.0 114250.0 ;
      RECT  63135.0 27915.0 63205.0 114250.0 ;
      RECT  63470.0 27915.0 63540.0 114250.0 ;
      RECT  63840.0 27915.0 63910.0 114250.0 ;
      RECT  64175.0 27915.0 64245.0 114250.0 ;
      RECT  64545.0 27915.0 64615.0 114250.0 ;
      RECT  64880.0 27915.0 64950.0 114250.0 ;
      RECT  65250.0 27915.0 65320.0 114250.0 ;
      RECT  65585.0 27915.0 65655.0 114250.0 ;
      RECT  65955.0 27915.0 66025.0 114250.0 ;
      RECT  66290.0 27915.0 66360.0 114250.0 ;
      RECT  66660.0 27915.0 66730.0 114250.0 ;
      RECT  66995.0 27915.0 67065.0 114250.0 ;
      RECT  67365.0 27915.0 67435.0 114250.0 ;
      RECT  67700.0 27915.0 67770.0 114250.0 ;
      RECT  68070.0 27915.0 68140.0 114250.0 ;
      RECT  68405.0 27915.0 68475.0 114250.0 ;
      RECT  68775.0 27915.0 68845.0 114250.0 ;
      RECT  69110.0 27915.0 69180.0 114250.0 ;
      RECT  69480.0 27915.0 69550.0 114250.0 ;
      RECT  69815.0 27915.0 69885.0 114250.0 ;
      RECT  70185.0 27915.0 70255.0 114250.0 ;
      RECT  70520.0 27915.0 70590.0 114250.0 ;
      RECT  70890.0 27915.0 70960.0 114250.0 ;
      RECT  71225.0 27915.0 71295.0 114250.0 ;
      RECT  71595.0 27915.0 71665.0 114250.0 ;
      RECT  71930.0 27915.0 72000.0 114250.0 ;
      RECT  72300.0 27915.0 72370.0 114250.0 ;
      RECT  72635.0 27915.0 72705.0 114250.0 ;
      RECT  73005.0 27915.0 73075.0 114250.0 ;
      RECT  73340.0 27915.0 73410.0 114250.0 ;
      RECT  73710.0 27915.0 73780.0 114250.0 ;
      RECT  74045.0 27915.0 74115.0 114250.0 ;
      RECT  74415.0 27915.0 74485.0 114250.0 ;
      RECT  74750.0 27915.0 74820.0 114250.0 ;
      RECT  75120.0 27915.0 75190.0 114250.0 ;
      RECT  75455.0 27915.0 75525.0 114250.0 ;
      RECT  75825.0 27915.0 75895.0 114250.0 ;
      RECT  76160.0 27915.0 76230.0 114250.0 ;
      RECT  76530.0 27915.0 76600.0 114250.0 ;
      RECT  76865.0 27915.0 76935.0 114250.0 ;
      RECT  77235.0 27915.0 77305.0 114250.0 ;
      RECT  77570.0 27915.0 77640.0 114250.0 ;
      RECT  77940.0 27915.0 78010.0 114250.0 ;
      RECT  78275.0 27915.0 78345.0 114250.0 ;
      RECT  78645.0 27915.0 78715.0 114250.0 ;
      RECT  78980.0 27915.0 79050.0 114250.0 ;
      RECT  79350.0 27915.0 79420.0 114250.0 ;
      RECT  79685.0 27915.0 79755.0 114250.0 ;
      RECT  80055.0 27915.0 80125.0 114250.0 ;
      RECT  80390.0 27915.0 80460.0 114250.0 ;
      RECT  80760.0 27915.0 80830.0 114250.0 ;
      RECT  81095.0 27915.0 81165.0 114250.0 ;
      RECT  81465.0 27915.0 81535.0 114250.0 ;
      RECT  81800.0 27915.0 81870.0 114250.0 ;
      RECT  82170.0 27915.0 82240.0 114250.0 ;
      RECT  82505.0 27915.0 82575.0 114250.0 ;
      RECT  82875.0 27915.0 82945.0 114250.0 ;
      RECT  83210.0 27915.0 83280.0 114250.0 ;
      RECT  83580.0 27915.0 83650.0 114250.0 ;
      RECT  83915.0 27915.0 83985.0 114250.0 ;
      RECT  84285.0 27915.0 84355.0 114250.0 ;
      RECT  84620.0 27915.0 84690.0 114250.0 ;
      RECT  84990.0 27915.0 85060.0 114250.0 ;
      RECT  85325.0 27915.0 85395.0 114250.0 ;
      RECT  85695.0 27915.0 85765.0 114250.0 ;
      RECT  86030.0 27915.0 86100.0 114250.0 ;
      RECT  86400.0 27915.0 86470.0 114250.0 ;
      RECT  86735.0 27915.0 86805.0 114250.0 ;
      RECT  87105.0 27915.0 87175.0 114250.0 ;
      RECT  87440.0 27915.0 87510.0 114250.0 ;
      RECT  87810.0 27915.0 87880.0 114250.0 ;
      RECT  88145.0 27915.0 88215.0 114250.0 ;
      RECT  88515.0 27915.0 88585.0 114250.0 ;
      RECT  88850.0 27915.0 88920.0 114250.0 ;
      RECT  89220.0 27915.0 89290.0 114250.0 ;
      RECT  89555.0 27915.0 89625.0 114250.0 ;
      RECT  89925.0 27915.0 89995.0 114250.0 ;
      RECT  90260.0 27915.0 90330.0 114250.0 ;
      RECT  90630.0 27915.0 90700.0 114250.0 ;
      RECT  90965.0 27915.0 91035.0 114250.0 ;
      RECT  91335.0 27915.0 91405.0 114250.0 ;
      RECT  91670.0 27915.0 91740.0 114250.0 ;
      RECT  92040.0 27915.0 92110.0 114250.0 ;
      RECT  92375.0 27915.0 92445.0 114250.0 ;
      RECT  92745.0 27915.0 92815.0 114250.0 ;
      RECT  93080.0 27915.0 93150.0 114250.0 ;
      RECT  93450.0 27915.0 93520.0 114250.0 ;
      RECT  93785.0 27915.0 93855.0 114250.0 ;
      RECT  94155.0 27915.0 94225.0 114250.0 ;
      RECT  94490.0 27915.0 94560.0 114250.0 ;
      RECT  94860.0 27915.0 94930.0 114250.0 ;
      RECT  95195.0 27915.0 95265.0 114250.0 ;
      RECT  95565.0 27915.0 95635.0 114250.0 ;
      RECT  95900.0 27915.0 95970.0 114250.0 ;
      RECT  96270.0 27915.0 96340.0 114250.0 ;
      RECT  96605.0 27915.0 96675.0 114250.0 ;
      RECT  96975.0 27915.0 97045.0 114250.0 ;
      RECT  97310.0 27915.0 97380.0 114250.0 ;
      RECT  97680.0 27915.0 97750.0 114250.0 ;
      RECT  98015.0 27915.0 98085.0 114250.0 ;
      RECT  98385.0 27915.0 98455.0 114250.0 ;
      RECT  98720.0 27915.0 98790.0 114250.0 ;
      RECT  99090.0 27915.0 99160.0 114250.0 ;
      RECT  99425.0 27915.0 99495.0 114250.0 ;
      RECT  99795.0 27915.0 99865.0 114250.0 ;
      RECT  100130.0 27915.0 100200.0 114250.0 ;
      RECT  100500.0 27915.0 100570.0 114250.0 ;
      RECT  100835.0 27915.0 100905.0 114250.0 ;
      RECT  101205.0 27915.0 101275.0 114250.0 ;
      RECT  101540.0 27915.0 101610.0 114250.0 ;
      RECT  101910.0 27915.0 101980.0 114250.0 ;
      RECT  102245.0 27915.0 102315.0 114250.0 ;
      RECT  102615.0 27915.0 102685.0 114250.0 ;
      RECT  102950.0 27915.0 103020.0 114250.0 ;
      RECT  103320.0 27915.0 103390.0 114250.0 ;
      RECT  103655.0 27915.0 103725.0 114250.0 ;
      RECT  104025.0 27915.0 104095.0 114250.0 ;
      RECT  104360.0 27915.0 104430.0 114250.0 ;
      RECT  104730.0 27915.0 104800.0 114250.0 ;
      RECT  105065.0 27915.0 105135.0 114250.0 ;
      RECT  105435.0 27915.0 105505.0 114250.0 ;
      RECT  105770.0 27915.0 105840.0 114250.0 ;
      RECT  15715.0 27915.0 15785.0 114250.0 ;
      RECT  16420.0 27915.0 16490.0 114250.0 ;
      RECT  17125.0 27915.0 17195.0 114250.0 ;
      RECT  17830.0 27915.0 17900.0 114250.0 ;
      RECT  18535.0 27915.0 18605.0 114250.0 ;
      RECT  19240.0 27915.0 19310.0 114250.0 ;
      RECT  19945.0 27915.0 20015.0 114250.0 ;
      RECT  20650.0 27915.0 20720.0 114250.0 ;
      RECT  21355.0 27915.0 21425.0 114250.0 ;
      RECT  22060.0 27915.0 22130.0 114250.0 ;
      RECT  22765.0 27915.0 22835.0 114250.0 ;
      RECT  23470.0 27915.0 23540.0 114250.0 ;
      RECT  24175.0 27915.0 24245.0 114250.0 ;
      RECT  24880.0 27915.0 24950.0 114250.0 ;
      RECT  25585.0 27915.0 25655.0 114250.0 ;
      RECT  26290.0 27915.0 26360.0 114250.0 ;
      RECT  26995.0 27915.0 27065.0 114250.0 ;
      RECT  27700.0 27915.0 27770.0 114250.0 ;
      RECT  28405.0 27915.0 28475.0 114250.0 ;
      RECT  29110.0 27915.0 29180.0 114250.0 ;
      RECT  29815.0 27915.0 29885.0 114250.0 ;
      RECT  30520.0 27915.0 30590.0 114250.0 ;
      RECT  31225.0 27915.0 31295.0 114250.0 ;
      RECT  31930.0 27915.0 32000.0 114250.0 ;
      RECT  32635.0 27915.0 32705.0 114250.0 ;
      RECT  33340.0 27915.0 33410.0 114250.0 ;
      RECT  34045.0 27915.0 34115.0 114250.0 ;
      RECT  34750.0 27915.0 34820.0 114250.0 ;
      RECT  35455.0 27915.0 35525.0 114250.0 ;
      RECT  36160.0 27915.0 36230.0 114250.0 ;
      RECT  36865.0 27915.0 36935.0 114250.0 ;
      RECT  37570.0 27915.0 37640.0 114250.0 ;
      RECT  38275.0 27915.0 38345.0 114250.0 ;
      RECT  38980.0 27915.0 39050.0 114250.0 ;
      RECT  39685.0 27915.0 39755.0 114250.0 ;
      RECT  40390.0 27915.0 40460.0 114250.0 ;
      RECT  41095.0 27915.0 41165.0 114250.0 ;
      RECT  41800.0 27915.0 41870.0 114250.0 ;
      RECT  42505.0 27915.0 42575.0 114250.0 ;
      RECT  43210.0 27915.0 43280.0 114250.0 ;
      RECT  43915.0 27915.0 43985.0 114250.0 ;
      RECT  44620.0 27915.0 44690.0 114250.0 ;
      RECT  45325.0 27915.0 45395.0 114250.0 ;
      RECT  46030.0 27915.0 46100.0 114250.0 ;
      RECT  46735.0 27915.0 46805.0 114250.0 ;
      RECT  47440.0 27915.0 47510.0 114250.0 ;
      RECT  48145.0 27915.0 48215.0 114250.0 ;
      RECT  48850.0 27915.0 48920.0 114250.0 ;
      RECT  49555.0 27915.0 49625.0 114250.0 ;
      RECT  50260.0 27915.0 50330.0 114250.0 ;
      RECT  50965.0 27915.0 51035.0 114250.0 ;
      RECT  51670.0 27915.0 51740.0 114250.0 ;
      RECT  52375.0 27915.0 52445.0 114250.0 ;
      RECT  53080.0 27915.0 53150.0 114250.0 ;
      RECT  53785.0 27915.0 53855.0 114250.0 ;
      RECT  54490.0 27915.0 54560.0 114250.0 ;
      RECT  55195.0 27915.0 55265.0 114250.0 ;
      RECT  55900.0 27915.0 55970.0 114250.0 ;
      RECT  56605.0 27915.0 56675.0 114250.0 ;
      RECT  57310.0 27915.0 57380.0 114250.0 ;
      RECT  58015.0 27915.0 58085.0 114250.0 ;
      RECT  58720.0 27915.0 58790.0 114250.0 ;
      RECT  59425.0 27915.0 59495.0 114250.0 ;
      RECT  60130.0 27915.0 60200.0 114250.0 ;
      RECT  60835.0 27915.0 60905.0 114250.0 ;
      RECT  61540.0 27915.0 61610.0 114250.0 ;
      RECT  62245.0 27915.0 62315.0 114250.0 ;
      RECT  62950.0 27915.0 63020.0 114250.0 ;
      RECT  63655.0 27915.0 63725.0 114250.0 ;
      RECT  64360.0 27915.0 64430.0 114250.0 ;
      RECT  65065.0 27915.0 65135.0 114250.0 ;
      RECT  65770.0 27915.0 65840.0 114250.0 ;
      RECT  66475.0 27915.0 66545.0 114250.0 ;
      RECT  67180.0 27915.0 67250.0 114250.0 ;
      RECT  67885.0 27915.0 67955.0 114250.0 ;
      RECT  68590.0 27915.0 68660.0 114250.0 ;
      RECT  69295.0 27915.0 69365.0 114250.0 ;
      RECT  70000.0 27915.0 70070.0 114250.0 ;
      RECT  70705.0 27915.0 70775.0 114250.0 ;
      RECT  71410.0 27915.0 71480.0 114250.0 ;
      RECT  72115.0 27915.0 72185.0 114250.0 ;
      RECT  72820.0 27915.0 72890.0 114250.0 ;
      RECT  73525.0 27915.0 73595.0 114250.0 ;
      RECT  74230.0 27915.0 74300.0 114250.0 ;
      RECT  74935.0 27915.0 75005.0 114250.0 ;
      RECT  75640.0 27915.0 75710.0 114250.0 ;
      RECT  76345.0 27915.0 76415.0 114250.0 ;
      RECT  77050.0 27915.0 77120.0 114250.0 ;
      RECT  77755.0 27915.0 77825.0 114250.0 ;
      RECT  78460.0 27915.0 78530.0 114250.0 ;
      RECT  79165.0 27915.0 79235.0 114250.0 ;
      RECT  79870.0 27915.0 79940.0 114250.0 ;
      RECT  80575.0 27915.0 80645.0 114250.0 ;
      RECT  81280.0 27915.0 81350.0 114250.0 ;
      RECT  81985.0 27915.0 82055.0 114250.0 ;
      RECT  82690.0 27915.0 82760.0 114250.0 ;
      RECT  83395.0 27915.0 83465.0 114250.0 ;
      RECT  84100.0 27915.0 84170.0 114250.0 ;
      RECT  84805.0 27915.0 84875.0 114250.0 ;
      RECT  85510.0 27915.0 85580.0 114250.0 ;
      RECT  86215.0 27915.0 86285.0 114250.0 ;
      RECT  86920.0 27915.0 86990.0 114250.0 ;
      RECT  87625.0 27915.0 87695.0 114250.0 ;
      RECT  88330.0 27915.0 88400.0 114250.0 ;
      RECT  89035.0 27915.0 89105.0 114250.0 ;
      RECT  89740.0 27915.0 89810.0 114250.0 ;
      RECT  90445.0 27915.0 90515.0 114250.0 ;
      RECT  91150.0 27915.0 91220.0 114250.0 ;
      RECT  91855.0 27915.0 91925.0 114250.0 ;
      RECT  92560.0 27915.0 92630.0 114250.0 ;
      RECT  93265.0 27915.0 93335.0 114250.0 ;
      RECT  93970.0 27915.0 94040.0 114250.0 ;
      RECT  94675.0 27915.0 94745.0 114250.0 ;
      RECT  95380.0 27915.0 95450.0 114250.0 ;
      RECT  96085.0 27915.0 96155.0 114250.0 ;
      RECT  96790.0 27915.0 96860.0 114250.0 ;
      RECT  97495.0 27915.0 97565.0 114250.0 ;
      RECT  98200.0 27915.0 98270.0 114250.0 ;
      RECT  98905.0 27915.0 98975.0 114250.0 ;
      RECT  99610.0 27915.0 99680.0 114250.0 ;
      RECT  100315.0 27915.0 100385.0 114250.0 ;
      RECT  101020.0 27915.0 101090.0 114250.0 ;
      RECT  101725.0 27915.0 101795.0 114250.0 ;
      RECT  102430.0 27915.0 102500.0 114250.0 ;
      RECT  103135.0 27915.0 103205.0 114250.0 ;
      RECT  103840.0 27915.0 103910.0 114250.0 ;
      RECT  104545.0 27915.0 104615.0 114250.0 ;
      RECT  105250.0 27915.0 105320.0 114250.0 ;
      RECT  105955.0 27915.0 106025.0 114250.0 ;
      RECT  15900.0 114777.5 15977.5 114912.5 ;
      RECT  16102.5 114777.5 16305.0 114912.5 ;
      RECT  15900.0 115307.5 15977.5 115442.5 ;
      RECT  16235.0 115307.5 16357.5 115442.5 ;
      RECT  15910.0 114777.5 15980.0 114912.5 ;
      RECT  16100.0 114777.5 16170.0 114912.5 ;
      RECT  15910.0 115307.5 15980.0 115442.5 ;
      RECT  16290.0 115307.5 16360.0 115442.5 ;
      RECT  15900.0 114655.0 15970.0 115822.5 ;
      RECT  16235.0 114655.0 16305.0 115822.5 ;
      RECT  16605.0 114777.5 16682.5 114912.5 ;
      RECT  16807.5 114777.5 17010.0 114912.5 ;
      RECT  16605.0 115307.5 16682.5 115442.5 ;
      RECT  16940.0 115307.5 17062.5 115442.5 ;
      RECT  16615.0 114777.5 16685.0 114912.5 ;
      RECT  16805.0 114777.5 16875.0 114912.5 ;
      RECT  16615.0 115307.5 16685.0 115442.5 ;
      RECT  16995.0 115307.5 17065.0 115442.5 ;
      RECT  16605.0 114655.0 16675.0 115822.5 ;
      RECT  16940.0 114655.0 17010.0 115822.5 ;
      RECT  17310.0 114777.5 17387.5 114912.5 ;
      RECT  17512.5 114777.5 17715.0 114912.5 ;
      RECT  17310.0 115307.5 17387.5 115442.5 ;
      RECT  17645.0 115307.5 17767.5 115442.5 ;
      RECT  17320.0 114777.5 17390.0 114912.5 ;
      RECT  17510.0 114777.5 17580.0 114912.5 ;
      RECT  17320.0 115307.5 17390.0 115442.5 ;
      RECT  17700.0 115307.5 17770.0 115442.5 ;
      RECT  17310.0 114655.0 17380.0 115822.5 ;
      RECT  17645.0 114655.0 17715.0 115822.5 ;
      RECT  18015.0 114777.5 18092.5 114912.5 ;
      RECT  18217.5 114777.5 18420.0 114912.5 ;
      RECT  18015.0 115307.5 18092.5 115442.5 ;
      RECT  18350.0 115307.5 18472.5 115442.5 ;
      RECT  18025.0 114777.5 18095.0 114912.5 ;
      RECT  18215.0 114777.5 18285.0 114912.5 ;
      RECT  18025.0 115307.5 18095.0 115442.5 ;
      RECT  18405.0 115307.5 18475.0 115442.5 ;
      RECT  18015.0 114655.0 18085.0 115822.5 ;
      RECT  18350.0 114655.0 18420.0 115822.5 ;
      RECT  18720.0 114777.5 18797.5 114912.5 ;
      RECT  18922.5 114777.5 19125.0 114912.5 ;
      RECT  18720.0 115307.5 18797.5 115442.5 ;
      RECT  19055.0 115307.5 19177.5 115442.5 ;
      RECT  18730.0 114777.5 18800.0 114912.5 ;
      RECT  18920.0 114777.5 18990.0 114912.5 ;
      RECT  18730.0 115307.5 18800.0 115442.5 ;
      RECT  19110.0 115307.5 19180.0 115442.5 ;
      RECT  18720.0 114655.0 18790.0 115822.5 ;
      RECT  19055.0 114655.0 19125.0 115822.5 ;
      RECT  19425.0 114777.5 19502.5 114912.5 ;
      RECT  19627.5 114777.5 19830.0 114912.5 ;
      RECT  19425.0 115307.5 19502.5 115442.5 ;
      RECT  19760.0 115307.5 19882.5 115442.5 ;
      RECT  19435.0 114777.5 19505.0 114912.5 ;
      RECT  19625.0 114777.5 19695.0 114912.5 ;
      RECT  19435.0 115307.5 19505.0 115442.5 ;
      RECT  19815.0 115307.5 19885.0 115442.5 ;
      RECT  19425.0 114655.0 19495.0 115822.5 ;
      RECT  19760.0 114655.0 19830.0 115822.5 ;
      RECT  20130.0 114777.5 20207.5 114912.5 ;
      RECT  20332.5 114777.5 20535.0 114912.5 ;
      RECT  20130.0 115307.5 20207.5 115442.5 ;
      RECT  20465.0 115307.5 20587.5 115442.5 ;
      RECT  20140.0 114777.5 20210.0 114912.5 ;
      RECT  20330.0 114777.5 20400.0 114912.5 ;
      RECT  20140.0 115307.5 20210.0 115442.5 ;
      RECT  20520.0 115307.5 20590.0 115442.5 ;
      RECT  20130.0 114655.0 20200.0 115822.5 ;
      RECT  20465.0 114655.0 20535.0 115822.5 ;
      RECT  20835.0 114777.5 20912.5 114912.5 ;
      RECT  21037.5 114777.5 21240.0 114912.5 ;
      RECT  20835.0 115307.5 20912.5 115442.5 ;
      RECT  21170.0 115307.5 21292.5 115442.5 ;
      RECT  20845.0 114777.5 20915.0 114912.5 ;
      RECT  21035.0 114777.5 21105.0 114912.5 ;
      RECT  20845.0 115307.5 20915.0 115442.5 ;
      RECT  21225.0 115307.5 21295.0 115442.5 ;
      RECT  20835.0 114655.0 20905.0 115822.5 ;
      RECT  21170.0 114655.0 21240.0 115822.5 ;
      RECT  21540.0 114777.5 21617.5 114912.5 ;
      RECT  21742.5 114777.5 21945.0 114912.5 ;
      RECT  21540.0 115307.5 21617.5 115442.5 ;
      RECT  21875.0 115307.5 21997.5 115442.5 ;
      RECT  21550.0 114777.5 21620.0 114912.5 ;
      RECT  21740.0 114777.5 21810.0 114912.5 ;
      RECT  21550.0 115307.5 21620.0 115442.5 ;
      RECT  21930.0 115307.5 22000.0 115442.5 ;
      RECT  21540.0 114655.0 21610.0 115822.5 ;
      RECT  21875.0 114655.0 21945.0 115822.5 ;
      RECT  22245.0 114777.5 22322.5 114912.5 ;
      RECT  22447.5 114777.5 22650.0 114912.5 ;
      RECT  22245.0 115307.5 22322.5 115442.5 ;
      RECT  22580.0 115307.5 22702.5 115442.5 ;
      RECT  22255.0 114777.5 22325.0 114912.5 ;
      RECT  22445.0 114777.5 22515.0 114912.5 ;
      RECT  22255.0 115307.5 22325.0 115442.5 ;
      RECT  22635.0 115307.5 22705.0 115442.5 ;
      RECT  22245.0 114655.0 22315.0 115822.5 ;
      RECT  22580.0 114655.0 22650.0 115822.5 ;
      RECT  22950.0 114777.5 23027.5 114912.5 ;
      RECT  23152.5 114777.5 23355.0 114912.5 ;
      RECT  22950.0 115307.5 23027.5 115442.5 ;
      RECT  23285.0 115307.5 23407.5 115442.5 ;
      RECT  22960.0 114777.5 23030.0 114912.5 ;
      RECT  23150.0 114777.5 23220.0 114912.5 ;
      RECT  22960.0 115307.5 23030.0 115442.5 ;
      RECT  23340.0 115307.5 23410.0 115442.5 ;
      RECT  22950.0 114655.0 23020.0 115822.5 ;
      RECT  23285.0 114655.0 23355.0 115822.5 ;
      RECT  23655.0 114777.5 23732.5 114912.5 ;
      RECT  23857.5 114777.5 24060.0 114912.5 ;
      RECT  23655.0 115307.5 23732.5 115442.5 ;
      RECT  23990.0 115307.5 24112.5 115442.5 ;
      RECT  23665.0 114777.5 23735.0 114912.5 ;
      RECT  23855.0 114777.5 23925.0 114912.5 ;
      RECT  23665.0 115307.5 23735.0 115442.5 ;
      RECT  24045.0 115307.5 24115.0 115442.5 ;
      RECT  23655.0 114655.0 23725.0 115822.5 ;
      RECT  23990.0 114655.0 24060.0 115822.5 ;
      RECT  24360.0 114777.5 24437.5 114912.5 ;
      RECT  24562.5 114777.5 24765.0 114912.5 ;
      RECT  24360.0 115307.5 24437.5 115442.5 ;
      RECT  24695.0 115307.5 24817.5 115442.5 ;
      RECT  24370.0 114777.5 24440.0 114912.5 ;
      RECT  24560.0 114777.5 24630.0 114912.5 ;
      RECT  24370.0 115307.5 24440.0 115442.5 ;
      RECT  24750.0 115307.5 24820.0 115442.5 ;
      RECT  24360.0 114655.0 24430.0 115822.5 ;
      RECT  24695.0 114655.0 24765.0 115822.5 ;
      RECT  25065.0 114777.5 25142.5 114912.5 ;
      RECT  25267.5 114777.5 25470.0 114912.5 ;
      RECT  25065.0 115307.5 25142.5 115442.5 ;
      RECT  25400.0 115307.5 25522.5 115442.5 ;
      RECT  25075.0 114777.5 25145.0 114912.5 ;
      RECT  25265.0 114777.5 25335.0 114912.5 ;
      RECT  25075.0 115307.5 25145.0 115442.5 ;
      RECT  25455.0 115307.5 25525.0 115442.5 ;
      RECT  25065.0 114655.0 25135.0 115822.5 ;
      RECT  25400.0 114655.0 25470.0 115822.5 ;
      RECT  25770.0 114777.5 25847.5 114912.5 ;
      RECT  25972.5 114777.5 26175.0 114912.5 ;
      RECT  25770.0 115307.5 25847.5 115442.5 ;
      RECT  26105.0 115307.5 26227.5 115442.5 ;
      RECT  25780.0 114777.5 25850.0 114912.5 ;
      RECT  25970.0 114777.5 26040.0 114912.5 ;
      RECT  25780.0 115307.5 25850.0 115442.5 ;
      RECT  26160.0 115307.5 26230.0 115442.5 ;
      RECT  25770.0 114655.0 25840.0 115822.5 ;
      RECT  26105.0 114655.0 26175.0 115822.5 ;
      RECT  26475.0 114777.5 26552.5 114912.5 ;
      RECT  26677.5 114777.5 26880.0 114912.5 ;
      RECT  26475.0 115307.5 26552.5 115442.5 ;
      RECT  26810.0 115307.5 26932.5 115442.5 ;
      RECT  26485.0 114777.5 26555.0 114912.5 ;
      RECT  26675.0 114777.5 26745.0 114912.5 ;
      RECT  26485.0 115307.5 26555.0 115442.5 ;
      RECT  26865.0 115307.5 26935.0 115442.5 ;
      RECT  26475.0 114655.0 26545.0 115822.5 ;
      RECT  26810.0 114655.0 26880.0 115822.5 ;
      RECT  27180.0 114777.5 27257.5 114912.5 ;
      RECT  27382.5 114777.5 27585.0 114912.5 ;
      RECT  27180.0 115307.5 27257.5 115442.5 ;
      RECT  27515.0 115307.5 27637.5 115442.5 ;
      RECT  27190.0 114777.5 27260.0 114912.5 ;
      RECT  27380.0 114777.5 27450.0 114912.5 ;
      RECT  27190.0 115307.5 27260.0 115442.5 ;
      RECT  27570.0 115307.5 27640.0 115442.5 ;
      RECT  27180.0 114655.0 27250.0 115822.5 ;
      RECT  27515.0 114655.0 27585.0 115822.5 ;
      RECT  27885.0 114777.5 27962.5 114912.5 ;
      RECT  28087.5 114777.5 28290.0 114912.5 ;
      RECT  27885.0 115307.5 27962.5 115442.5 ;
      RECT  28220.0 115307.5 28342.5 115442.5 ;
      RECT  27895.0 114777.5 27965.0 114912.5 ;
      RECT  28085.0 114777.5 28155.0 114912.5 ;
      RECT  27895.0 115307.5 27965.0 115442.5 ;
      RECT  28275.0 115307.5 28345.0 115442.5 ;
      RECT  27885.0 114655.0 27955.0 115822.5 ;
      RECT  28220.0 114655.0 28290.0 115822.5 ;
      RECT  28590.0 114777.5 28667.5 114912.5 ;
      RECT  28792.5 114777.5 28995.0 114912.5 ;
      RECT  28590.0 115307.5 28667.5 115442.5 ;
      RECT  28925.0 115307.5 29047.5 115442.5 ;
      RECT  28600.0 114777.5 28670.0 114912.5 ;
      RECT  28790.0 114777.5 28860.0 114912.5 ;
      RECT  28600.0 115307.5 28670.0 115442.5 ;
      RECT  28980.0 115307.5 29050.0 115442.5 ;
      RECT  28590.0 114655.0 28660.0 115822.5 ;
      RECT  28925.0 114655.0 28995.0 115822.5 ;
      RECT  29295.0 114777.5 29372.5 114912.5 ;
      RECT  29497.5 114777.5 29700.0 114912.5 ;
      RECT  29295.0 115307.5 29372.5 115442.5 ;
      RECT  29630.0 115307.5 29752.5 115442.5 ;
      RECT  29305.0 114777.5 29375.0 114912.5 ;
      RECT  29495.0 114777.5 29565.0 114912.5 ;
      RECT  29305.0 115307.5 29375.0 115442.5 ;
      RECT  29685.0 115307.5 29755.0 115442.5 ;
      RECT  29295.0 114655.0 29365.0 115822.5 ;
      RECT  29630.0 114655.0 29700.0 115822.5 ;
      RECT  30000.0 114777.5 30077.5 114912.5 ;
      RECT  30202.5 114777.5 30405.0 114912.5 ;
      RECT  30000.0 115307.5 30077.5 115442.5 ;
      RECT  30335.0 115307.5 30457.5 115442.5 ;
      RECT  30010.0 114777.5 30080.0 114912.5 ;
      RECT  30200.0 114777.5 30270.0 114912.5 ;
      RECT  30010.0 115307.5 30080.0 115442.5 ;
      RECT  30390.0 115307.5 30460.0 115442.5 ;
      RECT  30000.0 114655.0 30070.0 115822.5 ;
      RECT  30335.0 114655.0 30405.0 115822.5 ;
      RECT  30705.0 114777.5 30782.5 114912.5 ;
      RECT  30907.5 114777.5 31110.0 114912.5 ;
      RECT  30705.0 115307.5 30782.5 115442.5 ;
      RECT  31040.0 115307.5 31162.5 115442.5 ;
      RECT  30715.0 114777.5 30785.0 114912.5 ;
      RECT  30905.0 114777.5 30975.0 114912.5 ;
      RECT  30715.0 115307.5 30785.0 115442.5 ;
      RECT  31095.0 115307.5 31165.0 115442.5 ;
      RECT  30705.0 114655.0 30775.0 115822.5 ;
      RECT  31040.0 114655.0 31110.0 115822.5 ;
      RECT  31410.0 114777.5 31487.5 114912.5 ;
      RECT  31612.5 114777.5 31815.0 114912.5 ;
      RECT  31410.0 115307.5 31487.5 115442.5 ;
      RECT  31745.0 115307.5 31867.5 115442.5 ;
      RECT  31420.0 114777.5 31490.0 114912.5 ;
      RECT  31610.0 114777.5 31680.0 114912.5 ;
      RECT  31420.0 115307.5 31490.0 115442.5 ;
      RECT  31800.0 115307.5 31870.0 115442.5 ;
      RECT  31410.0 114655.0 31480.0 115822.5 ;
      RECT  31745.0 114655.0 31815.0 115822.5 ;
      RECT  32115.0 114777.5 32192.5 114912.5 ;
      RECT  32317.5 114777.5 32520.0 114912.5 ;
      RECT  32115.0 115307.5 32192.5 115442.5 ;
      RECT  32450.0 115307.5 32572.5 115442.5 ;
      RECT  32125.0 114777.5 32195.0 114912.5 ;
      RECT  32315.0 114777.5 32385.0 114912.5 ;
      RECT  32125.0 115307.5 32195.0 115442.5 ;
      RECT  32505.0 115307.5 32575.0 115442.5 ;
      RECT  32115.0 114655.0 32185.0 115822.5 ;
      RECT  32450.0 114655.0 32520.0 115822.5 ;
      RECT  32820.0 114777.5 32897.5 114912.5 ;
      RECT  33022.5 114777.5 33225.0 114912.5 ;
      RECT  32820.0 115307.5 32897.5 115442.5 ;
      RECT  33155.0 115307.5 33277.5 115442.5 ;
      RECT  32830.0 114777.5 32900.0 114912.5 ;
      RECT  33020.0 114777.5 33090.0 114912.5 ;
      RECT  32830.0 115307.5 32900.0 115442.5 ;
      RECT  33210.0 115307.5 33280.0 115442.5 ;
      RECT  32820.0 114655.0 32890.0 115822.5 ;
      RECT  33155.0 114655.0 33225.0 115822.5 ;
      RECT  33525.0 114777.5 33602.5 114912.5 ;
      RECT  33727.5 114777.5 33930.0 114912.5 ;
      RECT  33525.0 115307.5 33602.5 115442.5 ;
      RECT  33860.0 115307.5 33982.5 115442.5 ;
      RECT  33535.0 114777.5 33605.0 114912.5 ;
      RECT  33725.0 114777.5 33795.0 114912.5 ;
      RECT  33535.0 115307.5 33605.0 115442.5 ;
      RECT  33915.0 115307.5 33985.0 115442.5 ;
      RECT  33525.0 114655.0 33595.0 115822.5 ;
      RECT  33860.0 114655.0 33930.0 115822.5 ;
      RECT  34230.0 114777.5 34307.5 114912.5 ;
      RECT  34432.5 114777.5 34635.0 114912.5 ;
      RECT  34230.0 115307.5 34307.5 115442.5 ;
      RECT  34565.0 115307.5 34687.5 115442.5 ;
      RECT  34240.0 114777.5 34310.0 114912.5 ;
      RECT  34430.0 114777.5 34500.0 114912.5 ;
      RECT  34240.0 115307.5 34310.0 115442.5 ;
      RECT  34620.0 115307.5 34690.0 115442.5 ;
      RECT  34230.0 114655.0 34300.0 115822.5 ;
      RECT  34565.0 114655.0 34635.0 115822.5 ;
      RECT  34935.0 114777.5 35012.5 114912.5 ;
      RECT  35137.5 114777.5 35340.0 114912.5 ;
      RECT  34935.0 115307.5 35012.5 115442.5 ;
      RECT  35270.0 115307.5 35392.5 115442.5 ;
      RECT  34945.0 114777.5 35015.0 114912.5 ;
      RECT  35135.0 114777.5 35205.0 114912.5 ;
      RECT  34945.0 115307.5 35015.0 115442.5 ;
      RECT  35325.0 115307.5 35395.0 115442.5 ;
      RECT  34935.0 114655.0 35005.0 115822.5 ;
      RECT  35270.0 114655.0 35340.0 115822.5 ;
      RECT  35640.0 114777.5 35717.5 114912.5 ;
      RECT  35842.5 114777.5 36045.0 114912.5 ;
      RECT  35640.0 115307.5 35717.5 115442.5 ;
      RECT  35975.0 115307.5 36097.5 115442.5 ;
      RECT  35650.0 114777.5 35720.0 114912.5 ;
      RECT  35840.0 114777.5 35910.0 114912.5 ;
      RECT  35650.0 115307.5 35720.0 115442.5 ;
      RECT  36030.0 115307.5 36100.0 115442.5 ;
      RECT  35640.0 114655.0 35710.0 115822.5 ;
      RECT  35975.0 114655.0 36045.0 115822.5 ;
      RECT  36345.0 114777.5 36422.5 114912.5 ;
      RECT  36547.5 114777.5 36750.0 114912.5 ;
      RECT  36345.0 115307.5 36422.5 115442.5 ;
      RECT  36680.0 115307.5 36802.5 115442.5 ;
      RECT  36355.0 114777.5 36425.0 114912.5 ;
      RECT  36545.0 114777.5 36615.0 114912.5 ;
      RECT  36355.0 115307.5 36425.0 115442.5 ;
      RECT  36735.0 115307.5 36805.0 115442.5 ;
      RECT  36345.0 114655.0 36415.0 115822.5 ;
      RECT  36680.0 114655.0 36750.0 115822.5 ;
      RECT  37050.0 114777.5 37127.5 114912.5 ;
      RECT  37252.5 114777.5 37455.0 114912.5 ;
      RECT  37050.0 115307.5 37127.5 115442.5 ;
      RECT  37385.0 115307.5 37507.5 115442.5 ;
      RECT  37060.0 114777.5 37130.0 114912.5 ;
      RECT  37250.0 114777.5 37320.0 114912.5 ;
      RECT  37060.0 115307.5 37130.0 115442.5 ;
      RECT  37440.0 115307.5 37510.0 115442.5 ;
      RECT  37050.0 114655.0 37120.0 115822.5 ;
      RECT  37385.0 114655.0 37455.0 115822.5 ;
      RECT  37755.0 114777.5 37832.5 114912.5 ;
      RECT  37957.5 114777.5 38160.0 114912.5 ;
      RECT  37755.0 115307.5 37832.5 115442.5 ;
      RECT  38090.0 115307.5 38212.5 115442.5 ;
      RECT  37765.0 114777.5 37835.0 114912.5 ;
      RECT  37955.0 114777.5 38025.0 114912.5 ;
      RECT  37765.0 115307.5 37835.0 115442.5 ;
      RECT  38145.0 115307.5 38215.0 115442.5 ;
      RECT  37755.0 114655.0 37825.0 115822.5 ;
      RECT  38090.0 114655.0 38160.0 115822.5 ;
      RECT  38460.0 114777.5 38537.5 114912.5 ;
      RECT  38662.5 114777.5 38865.0 114912.5 ;
      RECT  38460.0 115307.5 38537.5 115442.5 ;
      RECT  38795.0 115307.5 38917.5 115442.5 ;
      RECT  38470.0 114777.5 38540.0 114912.5 ;
      RECT  38660.0 114777.5 38730.0 114912.5 ;
      RECT  38470.0 115307.5 38540.0 115442.5 ;
      RECT  38850.0 115307.5 38920.0 115442.5 ;
      RECT  38460.0 114655.0 38530.0 115822.5 ;
      RECT  38795.0 114655.0 38865.0 115822.5 ;
      RECT  39165.0 114777.5 39242.5 114912.5 ;
      RECT  39367.5 114777.5 39570.0 114912.5 ;
      RECT  39165.0 115307.5 39242.5 115442.5 ;
      RECT  39500.0 115307.5 39622.5 115442.5 ;
      RECT  39175.0 114777.5 39245.0 114912.5 ;
      RECT  39365.0 114777.5 39435.0 114912.5 ;
      RECT  39175.0 115307.5 39245.0 115442.5 ;
      RECT  39555.0 115307.5 39625.0 115442.5 ;
      RECT  39165.0 114655.0 39235.0 115822.5 ;
      RECT  39500.0 114655.0 39570.0 115822.5 ;
      RECT  39870.0 114777.5 39947.5 114912.5 ;
      RECT  40072.5 114777.5 40275.0 114912.5 ;
      RECT  39870.0 115307.5 39947.5 115442.5 ;
      RECT  40205.0 115307.5 40327.5 115442.5 ;
      RECT  39880.0 114777.5 39950.0 114912.5 ;
      RECT  40070.0 114777.5 40140.0 114912.5 ;
      RECT  39880.0 115307.5 39950.0 115442.5 ;
      RECT  40260.0 115307.5 40330.0 115442.5 ;
      RECT  39870.0 114655.0 39940.0 115822.5 ;
      RECT  40205.0 114655.0 40275.0 115822.5 ;
      RECT  40575.0 114777.5 40652.5 114912.5 ;
      RECT  40777.5 114777.5 40980.0 114912.5 ;
      RECT  40575.0 115307.5 40652.5 115442.5 ;
      RECT  40910.0 115307.5 41032.5 115442.5 ;
      RECT  40585.0 114777.5 40655.0 114912.5 ;
      RECT  40775.0 114777.5 40845.0 114912.5 ;
      RECT  40585.0 115307.5 40655.0 115442.5 ;
      RECT  40965.0 115307.5 41035.0 115442.5 ;
      RECT  40575.0 114655.0 40645.0 115822.5 ;
      RECT  40910.0 114655.0 40980.0 115822.5 ;
      RECT  41280.0 114777.5 41357.5 114912.5 ;
      RECT  41482.5 114777.5 41685.0 114912.5 ;
      RECT  41280.0 115307.5 41357.5 115442.5 ;
      RECT  41615.0 115307.5 41737.5 115442.5 ;
      RECT  41290.0 114777.5 41360.0 114912.5 ;
      RECT  41480.0 114777.5 41550.0 114912.5 ;
      RECT  41290.0 115307.5 41360.0 115442.5 ;
      RECT  41670.0 115307.5 41740.0 115442.5 ;
      RECT  41280.0 114655.0 41350.0 115822.5 ;
      RECT  41615.0 114655.0 41685.0 115822.5 ;
      RECT  41985.0 114777.5 42062.5 114912.5 ;
      RECT  42187.5 114777.5 42390.0 114912.5 ;
      RECT  41985.0 115307.5 42062.5 115442.5 ;
      RECT  42320.0 115307.5 42442.5 115442.5 ;
      RECT  41995.0 114777.5 42065.0 114912.5 ;
      RECT  42185.0 114777.5 42255.0 114912.5 ;
      RECT  41995.0 115307.5 42065.0 115442.5 ;
      RECT  42375.0 115307.5 42445.0 115442.5 ;
      RECT  41985.0 114655.0 42055.0 115822.5 ;
      RECT  42320.0 114655.0 42390.0 115822.5 ;
      RECT  42690.0 114777.5 42767.5 114912.5 ;
      RECT  42892.5 114777.5 43095.0 114912.5 ;
      RECT  42690.0 115307.5 42767.5 115442.5 ;
      RECT  43025.0 115307.5 43147.5 115442.5 ;
      RECT  42700.0 114777.5 42770.0 114912.5 ;
      RECT  42890.0 114777.5 42960.0 114912.5 ;
      RECT  42700.0 115307.5 42770.0 115442.5 ;
      RECT  43080.0 115307.5 43150.0 115442.5 ;
      RECT  42690.0 114655.0 42760.0 115822.5 ;
      RECT  43025.0 114655.0 43095.0 115822.5 ;
      RECT  43395.0 114777.5 43472.5 114912.5 ;
      RECT  43597.5 114777.5 43800.0 114912.5 ;
      RECT  43395.0 115307.5 43472.5 115442.5 ;
      RECT  43730.0 115307.5 43852.5 115442.5 ;
      RECT  43405.0 114777.5 43475.0 114912.5 ;
      RECT  43595.0 114777.5 43665.0 114912.5 ;
      RECT  43405.0 115307.5 43475.0 115442.5 ;
      RECT  43785.0 115307.5 43855.0 115442.5 ;
      RECT  43395.0 114655.0 43465.0 115822.5 ;
      RECT  43730.0 114655.0 43800.0 115822.5 ;
      RECT  44100.0 114777.5 44177.5 114912.5 ;
      RECT  44302.5 114777.5 44505.0 114912.5 ;
      RECT  44100.0 115307.5 44177.5 115442.5 ;
      RECT  44435.0 115307.5 44557.5 115442.5 ;
      RECT  44110.0 114777.5 44180.0 114912.5 ;
      RECT  44300.0 114777.5 44370.0 114912.5 ;
      RECT  44110.0 115307.5 44180.0 115442.5 ;
      RECT  44490.0 115307.5 44560.0 115442.5 ;
      RECT  44100.0 114655.0 44170.0 115822.5 ;
      RECT  44435.0 114655.0 44505.0 115822.5 ;
      RECT  44805.0 114777.5 44882.5 114912.5 ;
      RECT  45007.5 114777.5 45210.0 114912.5 ;
      RECT  44805.0 115307.5 44882.5 115442.5 ;
      RECT  45140.0 115307.5 45262.5 115442.5 ;
      RECT  44815.0 114777.5 44885.0 114912.5 ;
      RECT  45005.0 114777.5 45075.0 114912.5 ;
      RECT  44815.0 115307.5 44885.0 115442.5 ;
      RECT  45195.0 115307.5 45265.0 115442.5 ;
      RECT  44805.0 114655.0 44875.0 115822.5 ;
      RECT  45140.0 114655.0 45210.0 115822.5 ;
      RECT  45510.0 114777.5 45587.5 114912.5 ;
      RECT  45712.5 114777.5 45915.0 114912.5 ;
      RECT  45510.0 115307.5 45587.5 115442.5 ;
      RECT  45845.0 115307.5 45967.5 115442.5 ;
      RECT  45520.0 114777.5 45590.0 114912.5 ;
      RECT  45710.0 114777.5 45780.0 114912.5 ;
      RECT  45520.0 115307.5 45590.0 115442.5 ;
      RECT  45900.0 115307.5 45970.0 115442.5 ;
      RECT  45510.0 114655.0 45580.0 115822.5 ;
      RECT  45845.0 114655.0 45915.0 115822.5 ;
      RECT  46215.0 114777.5 46292.5 114912.5 ;
      RECT  46417.5 114777.5 46620.0 114912.5 ;
      RECT  46215.0 115307.5 46292.5 115442.5 ;
      RECT  46550.0 115307.5 46672.5 115442.5 ;
      RECT  46225.0 114777.5 46295.0 114912.5 ;
      RECT  46415.0 114777.5 46485.0 114912.5 ;
      RECT  46225.0 115307.5 46295.0 115442.5 ;
      RECT  46605.0 115307.5 46675.0 115442.5 ;
      RECT  46215.0 114655.0 46285.0 115822.5 ;
      RECT  46550.0 114655.0 46620.0 115822.5 ;
      RECT  46920.0 114777.5 46997.5 114912.5 ;
      RECT  47122.5 114777.5 47325.0 114912.5 ;
      RECT  46920.0 115307.5 46997.5 115442.5 ;
      RECT  47255.0 115307.5 47377.5 115442.5 ;
      RECT  46930.0 114777.5 47000.0 114912.5 ;
      RECT  47120.0 114777.5 47190.0 114912.5 ;
      RECT  46930.0 115307.5 47000.0 115442.5 ;
      RECT  47310.0 115307.5 47380.0 115442.5 ;
      RECT  46920.0 114655.0 46990.0 115822.5 ;
      RECT  47255.0 114655.0 47325.0 115822.5 ;
      RECT  47625.0 114777.5 47702.5 114912.5 ;
      RECT  47827.5 114777.5 48030.0 114912.5 ;
      RECT  47625.0 115307.5 47702.5 115442.5 ;
      RECT  47960.0 115307.5 48082.5 115442.5 ;
      RECT  47635.0 114777.5 47705.0 114912.5 ;
      RECT  47825.0 114777.5 47895.0 114912.5 ;
      RECT  47635.0 115307.5 47705.0 115442.5 ;
      RECT  48015.0 115307.5 48085.0 115442.5 ;
      RECT  47625.0 114655.0 47695.0 115822.5 ;
      RECT  47960.0 114655.0 48030.0 115822.5 ;
      RECT  48330.0 114777.5 48407.5 114912.5 ;
      RECT  48532.5 114777.5 48735.0 114912.5 ;
      RECT  48330.0 115307.5 48407.5 115442.5 ;
      RECT  48665.0 115307.5 48787.5 115442.5 ;
      RECT  48340.0 114777.5 48410.0 114912.5 ;
      RECT  48530.0 114777.5 48600.0 114912.5 ;
      RECT  48340.0 115307.5 48410.0 115442.5 ;
      RECT  48720.0 115307.5 48790.0 115442.5 ;
      RECT  48330.0 114655.0 48400.0 115822.5 ;
      RECT  48665.0 114655.0 48735.0 115822.5 ;
      RECT  49035.0 114777.5 49112.5 114912.5 ;
      RECT  49237.5 114777.5 49440.0 114912.5 ;
      RECT  49035.0 115307.5 49112.5 115442.5 ;
      RECT  49370.0 115307.5 49492.5 115442.5 ;
      RECT  49045.0 114777.5 49115.0 114912.5 ;
      RECT  49235.0 114777.5 49305.0 114912.5 ;
      RECT  49045.0 115307.5 49115.0 115442.5 ;
      RECT  49425.0 115307.5 49495.0 115442.5 ;
      RECT  49035.0 114655.0 49105.0 115822.5 ;
      RECT  49370.0 114655.0 49440.0 115822.5 ;
      RECT  49740.0 114777.5 49817.5 114912.5 ;
      RECT  49942.5 114777.5 50145.0 114912.5 ;
      RECT  49740.0 115307.5 49817.5 115442.5 ;
      RECT  50075.0 115307.5 50197.5 115442.5 ;
      RECT  49750.0 114777.5 49820.0 114912.5 ;
      RECT  49940.0 114777.5 50010.0 114912.5 ;
      RECT  49750.0 115307.5 49820.0 115442.5 ;
      RECT  50130.0 115307.5 50200.0 115442.5 ;
      RECT  49740.0 114655.0 49810.0 115822.5 ;
      RECT  50075.0 114655.0 50145.0 115822.5 ;
      RECT  50445.0 114777.5 50522.5 114912.5 ;
      RECT  50647.5 114777.5 50850.0 114912.5 ;
      RECT  50445.0 115307.5 50522.5 115442.5 ;
      RECT  50780.0 115307.5 50902.5 115442.5 ;
      RECT  50455.0 114777.5 50525.0 114912.5 ;
      RECT  50645.0 114777.5 50715.0 114912.5 ;
      RECT  50455.0 115307.5 50525.0 115442.5 ;
      RECT  50835.0 115307.5 50905.0 115442.5 ;
      RECT  50445.0 114655.0 50515.0 115822.5 ;
      RECT  50780.0 114655.0 50850.0 115822.5 ;
      RECT  51150.0 114777.5 51227.5 114912.5 ;
      RECT  51352.5 114777.5 51555.0 114912.5 ;
      RECT  51150.0 115307.5 51227.5 115442.5 ;
      RECT  51485.0 115307.5 51607.5 115442.5 ;
      RECT  51160.0 114777.5 51230.0 114912.5 ;
      RECT  51350.0 114777.5 51420.0 114912.5 ;
      RECT  51160.0 115307.5 51230.0 115442.5 ;
      RECT  51540.0 115307.5 51610.0 115442.5 ;
      RECT  51150.0 114655.0 51220.0 115822.5 ;
      RECT  51485.0 114655.0 51555.0 115822.5 ;
      RECT  51855.0 114777.5 51932.5 114912.5 ;
      RECT  52057.5 114777.5 52260.0 114912.5 ;
      RECT  51855.0 115307.5 51932.5 115442.5 ;
      RECT  52190.0 115307.5 52312.5 115442.5 ;
      RECT  51865.0 114777.5 51935.0 114912.5 ;
      RECT  52055.0 114777.5 52125.0 114912.5 ;
      RECT  51865.0 115307.5 51935.0 115442.5 ;
      RECT  52245.0 115307.5 52315.0 115442.5 ;
      RECT  51855.0 114655.0 51925.0 115822.5 ;
      RECT  52190.0 114655.0 52260.0 115822.5 ;
      RECT  52560.0 114777.5 52637.5 114912.5 ;
      RECT  52762.5 114777.5 52965.0 114912.5 ;
      RECT  52560.0 115307.5 52637.5 115442.5 ;
      RECT  52895.0 115307.5 53017.5 115442.5 ;
      RECT  52570.0 114777.5 52640.0 114912.5 ;
      RECT  52760.0 114777.5 52830.0 114912.5 ;
      RECT  52570.0 115307.5 52640.0 115442.5 ;
      RECT  52950.0 115307.5 53020.0 115442.5 ;
      RECT  52560.0 114655.0 52630.0 115822.5 ;
      RECT  52895.0 114655.0 52965.0 115822.5 ;
      RECT  53265.0 114777.5 53342.5 114912.5 ;
      RECT  53467.5 114777.5 53670.0 114912.5 ;
      RECT  53265.0 115307.5 53342.5 115442.5 ;
      RECT  53600.0 115307.5 53722.5 115442.5 ;
      RECT  53275.0 114777.5 53345.0 114912.5 ;
      RECT  53465.0 114777.5 53535.0 114912.5 ;
      RECT  53275.0 115307.5 53345.0 115442.5 ;
      RECT  53655.0 115307.5 53725.0 115442.5 ;
      RECT  53265.0 114655.0 53335.0 115822.5 ;
      RECT  53600.0 114655.0 53670.0 115822.5 ;
      RECT  53970.0 114777.5 54047.5 114912.5 ;
      RECT  54172.5 114777.5 54375.0 114912.5 ;
      RECT  53970.0 115307.5 54047.5 115442.5 ;
      RECT  54305.0 115307.5 54427.5 115442.5 ;
      RECT  53980.0 114777.5 54050.0 114912.5 ;
      RECT  54170.0 114777.5 54240.0 114912.5 ;
      RECT  53980.0 115307.5 54050.0 115442.5 ;
      RECT  54360.0 115307.5 54430.0 115442.5 ;
      RECT  53970.0 114655.0 54040.0 115822.5 ;
      RECT  54305.0 114655.0 54375.0 115822.5 ;
      RECT  54675.0 114777.5 54752.5 114912.5 ;
      RECT  54877.5 114777.5 55080.0 114912.5 ;
      RECT  54675.0 115307.5 54752.5 115442.5 ;
      RECT  55010.0 115307.5 55132.5 115442.5 ;
      RECT  54685.0 114777.5 54755.0 114912.5 ;
      RECT  54875.0 114777.5 54945.0 114912.5 ;
      RECT  54685.0 115307.5 54755.0 115442.5 ;
      RECT  55065.0 115307.5 55135.0 115442.5 ;
      RECT  54675.0 114655.0 54745.0 115822.5 ;
      RECT  55010.0 114655.0 55080.0 115822.5 ;
      RECT  55380.0 114777.5 55457.5 114912.5 ;
      RECT  55582.5 114777.5 55785.0 114912.5 ;
      RECT  55380.0 115307.5 55457.5 115442.5 ;
      RECT  55715.0 115307.5 55837.5 115442.5 ;
      RECT  55390.0 114777.5 55460.0 114912.5 ;
      RECT  55580.0 114777.5 55650.0 114912.5 ;
      RECT  55390.0 115307.5 55460.0 115442.5 ;
      RECT  55770.0 115307.5 55840.0 115442.5 ;
      RECT  55380.0 114655.0 55450.0 115822.5 ;
      RECT  55715.0 114655.0 55785.0 115822.5 ;
      RECT  56085.0 114777.5 56162.5 114912.5 ;
      RECT  56287.5 114777.5 56490.0 114912.5 ;
      RECT  56085.0 115307.5 56162.5 115442.5 ;
      RECT  56420.0 115307.5 56542.5 115442.5 ;
      RECT  56095.0 114777.5 56165.0 114912.5 ;
      RECT  56285.0 114777.5 56355.0 114912.5 ;
      RECT  56095.0 115307.5 56165.0 115442.5 ;
      RECT  56475.0 115307.5 56545.0 115442.5 ;
      RECT  56085.0 114655.0 56155.0 115822.5 ;
      RECT  56420.0 114655.0 56490.0 115822.5 ;
      RECT  56790.0 114777.5 56867.5 114912.5 ;
      RECT  56992.5 114777.5 57195.0 114912.5 ;
      RECT  56790.0 115307.5 56867.5 115442.5 ;
      RECT  57125.0 115307.5 57247.5 115442.5 ;
      RECT  56800.0 114777.5 56870.0 114912.5 ;
      RECT  56990.0 114777.5 57060.0 114912.5 ;
      RECT  56800.0 115307.5 56870.0 115442.5 ;
      RECT  57180.0 115307.5 57250.0 115442.5 ;
      RECT  56790.0 114655.0 56860.0 115822.5 ;
      RECT  57125.0 114655.0 57195.0 115822.5 ;
      RECT  57495.0 114777.5 57572.5 114912.5 ;
      RECT  57697.5 114777.5 57900.0 114912.5 ;
      RECT  57495.0 115307.5 57572.5 115442.5 ;
      RECT  57830.0 115307.5 57952.5 115442.5 ;
      RECT  57505.0 114777.5 57575.0 114912.5 ;
      RECT  57695.0 114777.5 57765.0 114912.5 ;
      RECT  57505.0 115307.5 57575.0 115442.5 ;
      RECT  57885.0 115307.5 57955.0 115442.5 ;
      RECT  57495.0 114655.0 57565.0 115822.5 ;
      RECT  57830.0 114655.0 57900.0 115822.5 ;
      RECT  58200.0 114777.5 58277.5 114912.5 ;
      RECT  58402.5 114777.5 58605.0 114912.5 ;
      RECT  58200.0 115307.5 58277.5 115442.5 ;
      RECT  58535.0 115307.5 58657.5 115442.5 ;
      RECT  58210.0 114777.5 58280.0 114912.5 ;
      RECT  58400.0 114777.5 58470.0 114912.5 ;
      RECT  58210.0 115307.5 58280.0 115442.5 ;
      RECT  58590.0 115307.5 58660.0 115442.5 ;
      RECT  58200.0 114655.0 58270.0 115822.5 ;
      RECT  58535.0 114655.0 58605.0 115822.5 ;
      RECT  58905.0 114777.5 58982.5 114912.5 ;
      RECT  59107.5 114777.5 59310.0 114912.5 ;
      RECT  58905.0 115307.5 58982.5 115442.5 ;
      RECT  59240.0 115307.5 59362.5 115442.5 ;
      RECT  58915.0 114777.5 58985.0 114912.5 ;
      RECT  59105.0 114777.5 59175.0 114912.5 ;
      RECT  58915.0 115307.5 58985.0 115442.5 ;
      RECT  59295.0 115307.5 59365.0 115442.5 ;
      RECT  58905.0 114655.0 58975.0 115822.5 ;
      RECT  59240.0 114655.0 59310.0 115822.5 ;
      RECT  59610.0 114777.5 59687.5 114912.5 ;
      RECT  59812.5 114777.5 60015.0 114912.5 ;
      RECT  59610.0 115307.5 59687.5 115442.5 ;
      RECT  59945.0 115307.5 60067.5 115442.5 ;
      RECT  59620.0 114777.5 59690.0 114912.5 ;
      RECT  59810.0 114777.5 59880.0 114912.5 ;
      RECT  59620.0 115307.5 59690.0 115442.5 ;
      RECT  60000.0 115307.5 60070.0 115442.5 ;
      RECT  59610.0 114655.0 59680.0 115822.5 ;
      RECT  59945.0 114655.0 60015.0 115822.5 ;
      RECT  60315.0 114777.5 60392.5 114912.5 ;
      RECT  60517.5 114777.5 60720.0 114912.5 ;
      RECT  60315.0 115307.5 60392.5 115442.5 ;
      RECT  60650.0 115307.5 60772.5 115442.5 ;
      RECT  60325.0 114777.5 60395.0 114912.5 ;
      RECT  60515.0 114777.5 60585.0 114912.5 ;
      RECT  60325.0 115307.5 60395.0 115442.5 ;
      RECT  60705.0 115307.5 60775.0 115442.5 ;
      RECT  60315.0 114655.0 60385.0 115822.5 ;
      RECT  60650.0 114655.0 60720.0 115822.5 ;
      RECT  61020.0 114777.5 61097.5 114912.5 ;
      RECT  61222.5 114777.5 61425.0 114912.5 ;
      RECT  61020.0 115307.5 61097.5 115442.5 ;
      RECT  61355.0 115307.5 61477.5 115442.5 ;
      RECT  61030.0 114777.5 61100.0 114912.5 ;
      RECT  61220.0 114777.5 61290.0 114912.5 ;
      RECT  61030.0 115307.5 61100.0 115442.5 ;
      RECT  61410.0 115307.5 61480.0 115442.5 ;
      RECT  61020.0 114655.0 61090.0 115822.5 ;
      RECT  61355.0 114655.0 61425.0 115822.5 ;
      RECT  61725.0 114777.5 61802.5 114912.5 ;
      RECT  61927.5 114777.5 62130.0 114912.5 ;
      RECT  61725.0 115307.5 61802.5 115442.5 ;
      RECT  62060.0 115307.5 62182.5 115442.5 ;
      RECT  61735.0 114777.5 61805.0 114912.5 ;
      RECT  61925.0 114777.5 61995.0 114912.5 ;
      RECT  61735.0 115307.5 61805.0 115442.5 ;
      RECT  62115.0 115307.5 62185.0 115442.5 ;
      RECT  61725.0 114655.0 61795.0 115822.5 ;
      RECT  62060.0 114655.0 62130.0 115822.5 ;
      RECT  62430.0 114777.5 62507.5 114912.5 ;
      RECT  62632.5 114777.5 62835.0 114912.5 ;
      RECT  62430.0 115307.5 62507.5 115442.5 ;
      RECT  62765.0 115307.5 62887.5 115442.5 ;
      RECT  62440.0 114777.5 62510.0 114912.5 ;
      RECT  62630.0 114777.5 62700.0 114912.5 ;
      RECT  62440.0 115307.5 62510.0 115442.5 ;
      RECT  62820.0 115307.5 62890.0 115442.5 ;
      RECT  62430.0 114655.0 62500.0 115822.5 ;
      RECT  62765.0 114655.0 62835.0 115822.5 ;
      RECT  63135.0 114777.5 63212.5 114912.5 ;
      RECT  63337.5 114777.5 63540.0 114912.5 ;
      RECT  63135.0 115307.5 63212.5 115442.5 ;
      RECT  63470.0 115307.5 63592.5 115442.5 ;
      RECT  63145.0 114777.5 63215.0 114912.5 ;
      RECT  63335.0 114777.5 63405.0 114912.5 ;
      RECT  63145.0 115307.5 63215.0 115442.5 ;
      RECT  63525.0 115307.5 63595.0 115442.5 ;
      RECT  63135.0 114655.0 63205.0 115822.5 ;
      RECT  63470.0 114655.0 63540.0 115822.5 ;
      RECT  63840.0 114777.5 63917.5 114912.5 ;
      RECT  64042.5 114777.5 64245.0 114912.5 ;
      RECT  63840.0 115307.5 63917.5 115442.5 ;
      RECT  64175.0 115307.5 64297.5 115442.5 ;
      RECT  63850.0 114777.5 63920.0 114912.5 ;
      RECT  64040.0 114777.5 64110.0 114912.5 ;
      RECT  63850.0 115307.5 63920.0 115442.5 ;
      RECT  64230.0 115307.5 64300.0 115442.5 ;
      RECT  63840.0 114655.0 63910.0 115822.5 ;
      RECT  64175.0 114655.0 64245.0 115822.5 ;
      RECT  64545.0 114777.5 64622.5 114912.5 ;
      RECT  64747.5 114777.5 64950.0 114912.5 ;
      RECT  64545.0 115307.5 64622.5 115442.5 ;
      RECT  64880.0 115307.5 65002.5 115442.5 ;
      RECT  64555.0 114777.5 64625.0 114912.5 ;
      RECT  64745.0 114777.5 64815.0 114912.5 ;
      RECT  64555.0 115307.5 64625.0 115442.5 ;
      RECT  64935.0 115307.5 65005.0 115442.5 ;
      RECT  64545.0 114655.0 64615.0 115822.5 ;
      RECT  64880.0 114655.0 64950.0 115822.5 ;
      RECT  65250.0 114777.5 65327.5 114912.5 ;
      RECT  65452.5 114777.5 65655.0 114912.5 ;
      RECT  65250.0 115307.5 65327.5 115442.5 ;
      RECT  65585.0 115307.5 65707.5 115442.5 ;
      RECT  65260.0 114777.5 65330.0 114912.5 ;
      RECT  65450.0 114777.5 65520.0 114912.5 ;
      RECT  65260.0 115307.5 65330.0 115442.5 ;
      RECT  65640.0 115307.5 65710.0 115442.5 ;
      RECT  65250.0 114655.0 65320.0 115822.5 ;
      RECT  65585.0 114655.0 65655.0 115822.5 ;
      RECT  65955.0 114777.5 66032.5 114912.5 ;
      RECT  66157.5 114777.5 66360.0 114912.5 ;
      RECT  65955.0 115307.5 66032.5 115442.5 ;
      RECT  66290.0 115307.5 66412.5 115442.5 ;
      RECT  65965.0 114777.5 66035.0 114912.5 ;
      RECT  66155.0 114777.5 66225.0 114912.5 ;
      RECT  65965.0 115307.5 66035.0 115442.5 ;
      RECT  66345.0 115307.5 66415.0 115442.5 ;
      RECT  65955.0 114655.0 66025.0 115822.5 ;
      RECT  66290.0 114655.0 66360.0 115822.5 ;
      RECT  66660.0 114777.5 66737.5 114912.5 ;
      RECT  66862.5 114777.5 67065.0 114912.5 ;
      RECT  66660.0 115307.5 66737.5 115442.5 ;
      RECT  66995.0 115307.5 67117.5 115442.5 ;
      RECT  66670.0 114777.5 66740.0 114912.5 ;
      RECT  66860.0 114777.5 66930.0 114912.5 ;
      RECT  66670.0 115307.5 66740.0 115442.5 ;
      RECT  67050.0 115307.5 67120.0 115442.5 ;
      RECT  66660.0 114655.0 66730.0 115822.5 ;
      RECT  66995.0 114655.0 67065.0 115822.5 ;
      RECT  67365.0 114777.5 67442.5 114912.5 ;
      RECT  67567.5 114777.5 67770.0 114912.5 ;
      RECT  67365.0 115307.5 67442.5 115442.5 ;
      RECT  67700.0 115307.5 67822.5 115442.5 ;
      RECT  67375.0 114777.5 67445.0 114912.5 ;
      RECT  67565.0 114777.5 67635.0 114912.5 ;
      RECT  67375.0 115307.5 67445.0 115442.5 ;
      RECT  67755.0 115307.5 67825.0 115442.5 ;
      RECT  67365.0 114655.0 67435.0 115822.5 ;
      RECT  67700.0 114655.0 67770.0 115822.5 ;
      RECT  68070.0 114777.5 68147.5 114912.5 ;
      RECT  68272.5 114777.5 68475.0 114912.5 ;
      RECT  68070.0 115307.5 68147.5 115442.5 ;
      RECT  68405.0 115307.5 68527.5 115442.5 ;
      RECT  68080.0 114777.5 68150.0 114912.5 ;
      RECT  68270.0 114777.5 68340.0 114912.5 ;
      RECT  68080.0 115307.5 68150.0 115442.5 ;
      RECT  68460.0 115307.5 68530.0 115442.5 ;
      RECT  68070.0 114655.0 68140.0 115822.5 ;
      RECT  68405.0 114655.0 68475.0 115822.5 ;
      RECT  68775.0 114777.5 68852.5 114912.5 ;
      RECT  68977.5 114777.5 69180.0 114912.5 ;
      RECT  68775.0 115307.5 68852.5 115442.5 ;
      RECT  69110.0 115307.5 69232.5 115442.5 ;
      RECT  68785.0 114777.5 68855.0 114912.5 ;
      RECT  68975.0 114777.5 69045.0 114912.5 ;
      RECT  68785.0 115307.5 68855.0 115442.5 ;
      RECT  69165.0 115307.5 69235.0 115442.5 ;
      RECT  68775.0 114655.0 68845.0 115822.5 ;
      RECT  69110.0 114655.0 69180.0 115822.5 ;
      RECT  69480.0 114777.5 69557.5 114912.5 ;
      RECT  69682.5 114777.5 69885.0 114912.5 ;
      RECT  69480.0 115307.5 69557.5 115442.5 ;
      RECT  69815.0 115307.5 69937.5 115442.5 ;
      RECT  69490.0 114777.5 69560.0 114912.5 ;
      RECT  69680.0 114777.5 69750.0 114912.5 ;
      RECT  69490.0 115307.5 69560.0 115442.5 ;
      RECT  69870.0 115307.5 69940.0 115442.5 ;
      RECT  69480.0 114655.0 69550.0 115822.5 ;
      RECT  69815.0 114655.0 69885.0 115822.5 ;
      RECT  70185.0 114777.5 70262.5 114912.5 ;
      RECT  70387.5 114777.5 70590.0 114912.5 ;
      RECT  70185.0 115307.5 70262.5 115442.5 ;
      RECT  70520.0 115307.5 70642.5 115442.5 ;
      RECT  70195.0 114777.5 70265.0 114912.5 ;
      RECT  70385.0 114777.5 70455.0 114912.5 ;
      RECT  70195.0 115307.5 70265.0 115442.5 ;
      RECT  70575.0 115307.5 70645.0 115442.5 ;
      RECT  70185.0 114655.0 70255.0 115822.5 ;
      RECT  70520.0 114655.0 70590.0 115822.5 ;
      RECT  70890.0 114777.5 70967.5 114912.5 ;
      RECT  71092.5 114777.5 71295.0 114912.5 ;
      RECT  70890.0 115307.5 70967.5 115442.5 ;
      RECT  71225.0 115307.5 71347.5 115442.5 ;
      RECT  70900.0 114777.5 70970.0 114912.5 ;
      RECT  71090.0 114777.5 71160.0 114912.5 ;
      RECT  70900.0 115307.5 70970.0 115442.5 ;
      RECT  71280.0 115307.5 71350.0 115442.5 ;
      RECT  70890.0 114655.0 70960.0 115822.5 ;
      RECT  71225.0 114655.0 71295.0 115822.5 ;
      RECT  71595.0 114777.5 71672.5 114912.5 ;
      RECT  71797.5 114777.5 72000.0 114912.5 ;
      RECT  71595.0 115307.5 71672.5 115442.5 ;
      RECT  71930.0 115307.5 72052.5 115442.5 ;
      RECT  71605.0 114777.5 71675.0 114912.5 ;
      RECT  71795.0 114777.5 71865.0 114912.5 ;
      RECT  71605.0 115307.5 71675.0 115442.5 ;
      RECT  71985.0 115307.5 72055.0 115442.5 ;
      RECT  71595.0 114655.0 71665.0 115822.5 ;
      RECT  71930.0 114655.0 72000.0 115822.5 ;
      RECT  72300.0 114777.5 72377.5 114912.5 ;
      RECT  72502.5 114777.5 72705.0 114912.5 ;
      RECT  72300.0 115307.5 72377.5 115442.5 ;
      RECT  72635.0 115307.5 72757.5 115442.5 ;
      RECT  72310.0 114777.5 72380.0 114912.5 ;
      RECT  72500.0 114777.5 72570.0 114912.5 ;
      RECT  72310.0 115307.5 72380.0 115442.5 ;
      RECT  72690.0 115307.5 72760.0 115442.5 ;
      RECT  72300.0 114655.0 72370.0 115822.5 ;
      RECT  72635.0 114655.0 72705.0 115822.5 ;
      RECT  73005.0 114777.5 73082.5 114912.5 ;
      RECT  73207.5 114777.5 73410.0 114912.5 ;
      RECT  73005.0 115307.5 73082.5 115442.5 ;
      RECT  73340.0 115307.5 73462.5 115442.5 ;
      RECT  73015.0 114777.5 73085.0 114912.5 ;
      RECT  73205.0 114777.5 73275.0 114912.5 ;
      RECT  73015.0 115307.5 73085.0 115442.5 ;
      RECT  73395.0 115307.5 73465.0 115442.5 ;
      RECT  73005.0 114655.0 73075.0 115822.5 ;
      RECT  73340.0 114655.0 73410.0 115822.5 ;
      RECT  73710.0 114777.5 73787.5 114912.5 ;
      RECT  73912.5 114777.5 74115.0 114912.5 ;
      RECT  73710.0 115307.5 73787.5 115442.5 ;
      RECT  74045.0 115307.5 74167.5 115442.5 ;
      RECT  73720.0 114777.5 73790.0 114912.5 ;
      RECT  73910.0 114777.5 73980.0 114912.5 ;
      RECT  73720.0 115307.5 73790.0 115442.5 ;
      RECT  74100.0 115307.5 74170.0 115442.5 ;
      RECT  73710.0 114655.0 73780.0 115822.5 ;
      RECT  74045.0 114655.0 74115.0 115822.5 ;
      RECT  74415.0 114777.5 74492.5 114912.5 ;
      RECT  74617.5 114777.5 74820.0 114912.5 ;
      RECT  74415.0 115307.5 74492.5 115442.5 ;
      RECT  74750.0 115307.5 74872.5 115442.5 ;
      RECT  74425.0 114777.5 74495.0 114912.5 ;
      RECT  74615.0 114777.5 74685.0 114912.5 ;
      RECT  74425.0 115307.5 74495.0 115442.5 ;
      RECT  74805.0 115307.5 74875.0 115442.5 ;
      RECT  74415.0 114655.0 74485.0 115822.5 ;
      RECT  74750.0 114655.0 74820.0 115822.5 ;
      RECT  75120.0 114777.5 75197.5 114912.5 ;
      RECT  75322.5 114777.5 75525.0 114912.5 ;
      RECT  75120.0 115307.5 75197.5 115442.5 ;
      RECT  75455.0 115307.5 75577.5 115442.5 ;
      RECT  75130.0 114777.5 75200.0 114912.5 ;
      RECT  75320.0 114777.5 75390.0 114912.5 ;
      RECT  75130.0 115307.5 75200.0 115442.5 ;
      RECT  75510.0 115307.5 75580.0 115442.5 ;
      RECT  75120.0 114655.0 75190.0 115822.5 ;
      RECT  75455.0 114655.0 75525.0 115822.5 ;
      RECT  75825.0 114777.5 75902.5 114912.5 ;
      RECT  76027.5 114777.5 76230.0 114912.5 ;
      RECT  75825.0 115307.5 75902.5 115442.5 ;
      RECT  76160.0 115307.5 76282.5 115442.5 ;
      RECT  75835.0 114777.5 75905.0 114912.5 ;
      RECT  76025.0 114777.5 76095.0 114912.5 ;
      RECT  75835.0 115307.5 75905.0 115442.5 ;
      RECT  76215.0 115307.5 76285.0 115442.5 ;
      RECT  75825.0 114655.0 75895.0 115822.5 ;
      RECT  76160.0 114655.0 76230.0 115822.5 ;
      RECT  76530.0 114777.5 76607.5 114912.5 ;
      RECT  76732.5 114777.5 76935.0 114912.5 ;
      RECT  76530.0 115307.5 76607.5 115442.5 ;
      RECT  76865.0 115307.5 76987.5 115442.5 ;
      RECT  76540.0 114777.5 76610.0 114912.5 ;
      RECT  76730.0 114777.5 76800.0 114912.5 ;
      RECT  76540.0 115307.5 76610.0 115442.5 ;
      RECT  76920.0 115307.5 76990.0 115442.5 ;
      RECT  76530.0 114655.0 76600.0 115822.5 ;
      RECT  76865.0 114655.0 76935.0 115822.5 ;
      RECT  77235.0 114777.5 77312.5 114912.5 ;
      RECT  77437.5 114777.5 77640.0 114912.5 ;
      RECT  77235.0 115307.5 77312.5 115442.5 ;
      RECT  77570.0 115307.5 77692.5 115442.5 ;
      RECT  77245.0 114777.5 77315.0 114912.5 ;
      RECT  77435.0 114777.5 77505.0 114912.5 ;
      RECT  77245.0 115307.5 77315.0 115442.5 ;
      RECT  77625.0 115307.5 77695.0 115442.5 ;
      RECT  77235.0 114655.0 77305.0 115822.5 ;
      RECT  77570.0 114655.0 77640.0 115822.5 ;
      RECT  77940.0 114777.5 78017.5 114912.5 ;
      RECT  78142.5 114777.5 78345.0 114912.5 ;
      RECT  77940.0 115307.5 78017.5 115442.5 ;
      RECT  78275.0 115307.5 78397.5 115442.5 ;
      RECT  77950.0 114777.5 78020.0 114912.5 ;
      RECT  78140.0 114777.5 78210.0 114912.5 ;
      RECT  77950.0 115307.5 78020.0 115442.5 ;
      RECT  78330.0 115307.5 78400.0 115442.5 ;
      RECT  77940.0 114655.0 78010.0 115822.5 ;
      RECT  78275.0 114655.0 78345.0 115822.5 ;
      RECT  78645.0 114777.5 78722.5 114912.5 ;
      RECT  78847.5 114777.5 79050.0 114912.5 ;
      RECT  78645.0 115307.5 78722.5 115442.5 ;
      RECT  78980.0 115307.5 79102.5 115442.5 ;
      RECT  78655.0 114777.5 78725.0 114912.5 ;
      RECT  78845.0 114777.5 78915.0 114912.5 ;
      RECT  78655.0 115307.5 78725.0 115442.5 ;
      RECT  79035.0 115307.5 79105.0 115442.5 ;
      RECT  78645.0 114655.0 78715.0 115822.5 ;
      RECT  78980.0 114655.0 79050.0 115822.5 ;
      RECT  79350.0 114777.5 79427.5 114912.5 ;
      RECT  79552.5 114777.5 79755.0 114912.5 ;
      RECT  79350.0 115307.5 79427.5 115442.5 ;
      RECT  79685.0 115307.5 79807.5 115442.5 ;
      RECT  79360.0 114777.5 79430.0 114912.5 ;
      RECT  79550.0 114777.5 79620.0 114912.5 ;
      RECT  79360.0 115307.5 79430.0 115442.5 ;
      RECT  79740.0 115307.5 79810.0 115442.5 ;
      RECT  79350.0 114655.0 79420.0 115822.5 ;
      RECT  79685.0 114655.0 79755.0 115822.5 ;
      RECT  80055.0 114777.5 80132.5 114912.5 ;
      RECT  80257.5 114777.5 80460.0 114912.5 ;
      RECT  80055.0 115307.5 80132.5 115442.5 ;
      RECT  80390.0 115307.5 80512.5 115442.5 ;
      RECT  80065.0 114777.5 80135.0 114912.5 ;
      RECT  80255.0 114777.5 80325.0 114912.5 ;
      RECT  80065.0 115307.5 80135.0 115442.5 ;
      RECT  80445.0 115307.5 80515.0 115442.5 ;
      RECT  80055.0 114655.0 80125.0 115822.5 ;
      RECT  80390.0 114655.0 80460.0 115822.5 ;
      RECT  80760.0 114777.5 80837.5 114912.5 ;
      RECT  80962.5 114777.5 81165.0 114912.5 ;
      RECT  80760.0 115307.5 80837.5 115442.5 ;
      RECT  81095.0 115307.5 81217.5 115442.5 ;
      RECT  80770.0 114777.5 80840.0 114912.5 ;
      RECT  80960.0 114777.5 81030.0 114912.5 ;
      RECT  80770.0 115307.5 80840.0 115442.5 ;
      RECT  81150.0 115307.5 81220.0 115442.5 ;
      RECT  80760.0 114655.0 80830.0 115822.5 ;
      RECT  81095.0 114655.0 81165.0 115822.5 ;
      RECT  81465.0 114777.5 81542.5 114912.5 ;
      RECT  81667.5 114777.5 81870.0 114912.5 ;
      RECT  81465.0 115307.5 81542.5 115442.5 ;
      RECT  81800.0 115307.5 81922.5 115442.5 ;
      RECT  81475.0 114777.5 81545.0 114912.5 ;
      RECT  81665.0 114777.5 81735.0 114912.5 ;
      RECT  81475.0 115307.5 81545.0 115442.5 ;
      RECT  81855.0 115307.5 81925.0 115442.5 ;
      RECT  81465.0 114655.0 81535.0 115822.5 ;
      RECT  81800.0 114655.0 81870.0 115822.5 ;
      RECT  82170.0 114777.5 82247.5 114912.5 ;
      RECT  82372.5 114777.5 82575.0 114912.5 ;
      RECT  82170.0 115307.5 82247.5 115442.5 ;
      RECT  82505.0 115307.5 82627.5 115442.5 ;
      RECT  82180.0 114777.5 82250.0 114912.5 ;
      RECT  82370.0 114777.5 82440.0 114912.5 ;
      RECT  82180.0 115307.5 82250.0 115442.5 ;
      RECT  82560.0 115307.5 82630.0 115442.5 ;
      RECT  82170.0 114655.0 82240.0 115822.5 ;
      RECT  82505.0 114655.0 82575.0 115822.5 ;
      RECT  82875.0 114777.5 82952.5 114912.5 ;
      RECT  83077.5 114777.5 83280.0 114912.5 ;
      RECT  82875.0 115307.5 82952.5 115442.5 ;
      RECT  83210.0 115307.5 83332.5 115442.5 ;
      RECT  82885.0 114777.5 82955.0 114912.5 ;
      RECT  83075.0 114777.5 83145.0 114912.5 ;
      RECT  82885.0 115307.5 82955.0 115442.5 ;
      RECT  83265.0 115307.5 83335.0 115442.5 ;
      RECT  82875.0 114655.0 82945.0 115822.5 ;
      RECT  83210.0 114655.0 83280.0 115822.5 ;
      RECT  83580.0 114777.5 83657.5 114912.5 ;
      RECT  83782.5 114777.5 83985.0 114912.5 ;
      RECT  83580.0 115307.5 83657.5 115442.5 ;
      RECT  83915.0 115307.5 84037.5 115442.5 ;
      RECT  83590.0 114777.5 83660.0 114912.5 ;
      RECT  83780.0 114777.5 83850.0 114912.5 ;
      RECT  83590.0 115307.5 83660.0 115442.5 ;
      RECT  83970.0 115307.5 84040.0 115442.5 ;
      RECT  83580.0 114655.0 83650.0 115822.5 ;
      RECT  83915.0 114655.0 83985.0 115822.5 ;
      RECT  84285.0 114777.5 84362.5 114912.5 ;
      RECT  84487.5 114777.5 84690.0 114912.5 ;
      RECT  84285.0 115307.5 84362.5 115442.5 ;
      RECT  84620.0 115307.5 84742.5 115442.5 ;
      RECT  84295.0 114777.5 84365.0 114912.5 ;
      RECT  84485.0 114777.5 84555.0 114912.5 ;
      RECT  84295.0 115307.5 84365.0 115442.5 ;
      RECT  84675.0 115307.5 84745.0 115442.5 ;
      RECT  84285.0 114655.0 84355.0 115822.5 ;
      RECT  84620.0 114655.0 84690.0 115822.5 ;
      RECT  84990.0 114777.5 85067.5 114912.5 ;
      RECT  85192.5 114777.5 85395.0 114912.5 ;
      RECT  84990.0 115307.5 85067.5 115442.5 ;
      RECT  85325.0 115307.5 85447.5 115442.5 ;
      RECT  85000.0 114777.5 85070.0 114912.5 ;
      RECT  85190.0 114777.5 85260.0 114912.5 ;
      RECT  85000.0 115307.5 85070.0 115442.5 ;
      RECT  85380.0 115307.5 85450.0 115442.5 ;
      RECT  84990.0 114655.0 85060.0 115822.5 ;
      RECT  85325.0 114655.0 85395.0 115822.5 ;
      RECT  85695.0 114777.5 85772.5 114912.5 ;
      RECT  85897.5 114777.5 86100.0 114912.5 ;
      RECT  85695.0 115307.5 85772.5 115442.5 ;
      RECT  86030.0 115307.5 86152.5 115442.5 ;
      RECT  85705.0 114777.5 85775.0 114912.5 ;
      RECT  85895.0 114777.5 85965.0 114912.5 ;
      RECT  85705.0 115307.5 85775.0 115442.5 ;
      RECT  86085.0 115307.5 86155.0 115442.5 ;
      RECT  85695.0 114655.0 85765.0 115822.5 ;
      RECT  86030.0 114655.0 86100.0 115822.5 ;
      RECT  86400.0 114777.5 86477.5 114912.5 ;
      RECT  86602.5 114777.5 86805.0 114912.5 ;
      RECT  86400.0 115307.5 86477.5 115442.5 ;
      RECT  86735.0 115307.5 86857.5 115442.5 ;
      RECT  86410.0 114777.5 86480.0 114912.5 ;
      RECT  86600.0 114777.5 86670.0 114912.5 ;
      RECT  86410.0 115307.5 86480.0 115442.5 ;
      RECT  86790.0 115307.5 86860.0 115442.5 ;
      RECT  86400.0 114655.0 86470.0 115822.5 ;
      RECT  86735.0 114655.0 86805.0 115822.5 ;
      RECT  87105.0 114777.5 87182.5 114912.5 ;
      RECT  87307.5 114777.5 87510.0 114912.5 ;
      RECT  87105.0 115307.5 87182.5 115442.5 ;
      RECT  87440.0 115307.5 87562.5 115442.5 ;
      RECT  87115.0 114777.5 87185.0 114912.5 ;
      RECT  87305.0 114777.5 87375.0 114912.5 ;
      RECT  87115.0 115307.5 87185.0 115442.5 ;
      RECT  87495.0 115307.5 87565.0 115442.5 ;
      RECT  87105.0 114655.0 87175.0 115822.5 ;
      RECT  87440.0 114655.0 87510.0 115822.5 ;
      RECT  87810.0 114777.5 87887.5 114912.5 ;
      RECT  88012.5 114777.5 88215.0 114912.5 ;
      RECT  87810.0 115307.5 87887.5 115442.5 ;
      RECT  88145.0 115307.5 88267.5 115442.5 ;
      RECT  87820.0 114777.5 87890.0 114912.5 ;
      RECT  88010.0 114777.5 88080.0 114912.5 ;
      RECT  87820.0 115307.5 87890.0 115442.5 ;
      RECT  88200.0 115307.5 88270.0 115442.5 ;
      RECT  87810.0 114655.0 87880.0 115822.5 ;
      RECT  88145.0 114655.0 88215.0 115822.5 ;
      RECT  88515.0 114777.5 88592.5 114912.5 ;
      RECT  88717.5 114777.5 88920.0 114912.5 ;
      RECT  88515.0 115307.5 88592.5 115442.5 ;
      RECT  88850.0 115307.5 88972.5 115442.5 ;
      RECT  88525.0 114777.5 88595.0 114912.5 ;
      RECT  88715.0 114777.5 88785.0 114912.5 ;
      RECT  88525.0 115307.5 88595.0 115442.5 ;
      RECT  88905.0 115307.5 88975.0 115442.5 ;
      RECT  88515.0 114655.0 88585.0 115822.5 ;
      RECT  88850.0 114655.0 88920.0 115822.5 ;
      RECT  89220.0 114777.5 89297.5 114912.5 ;
      RECT  89422.5 114777.5 89625.0 114912.5 ;
      RECT  89220.0 115307.5 89297.5 115442.5 ;
      RECT  89555.0 115307.5 89677.5 115442.5 ;
      RECT  89230.0 114777.5 89300.0 114912.5 ;
      RECT  89420.0 114777.5 89490.0 114912.5 ;
      RECT  89230.0 115307.5 89300.0 115442.5 ;
      RECT  89610.0 115307.5 89680.0 115442.5 ;
      RECT  89220.0 114655.0 89290.0 115822.5 ;
      RECT  89555.0 114655.0 89625.0 115822.5 ;
      RECT  89925.0 114777.5 90002.5 114912.5 ;
      RECT  90127.5 114777.5 90330.0 114912.5 ;
      RECT  89925.0 115307.5 90002.5 115442.5 ;
      RECT  90260.0 115307.5 90382.5 115442.5 ;
      RECT  89935.0 114777.5 90005.0 114912.5 ;
      RECT  90125.0 114777.5 90195.0 114912.5 ;
      RECT  89935.0 115307.5 90005.0 115442.5 ;
      RECT  90315.0 115307.5 90385.0 115442.5 ;
      RECT  89925.0 114655.0 89995.0 115822.5 ;
      RECT  90260.0 114655.0 90330.0 115822.5 ;
      RECT  90630.0 114777.5 90707.5 114912.5 ;
      RECT  90832.5 114777.5 91035.0 114912.5 ;
      RECT  90630.0 115307.5 90707.5 115442.5 ;
      RECT  90965.0 115307.5 91087.5 115442.5 ;
      RECT  90640.0 114777.5 90710.0 114912.5 ;
      RECT  90830.0 114777.5 90900.0 114912.5 ;
      RECT  90640.0 115307.5 90710.0 115442.5 ;
      RECT  91020.0 115307.5 91090.0 115442.5 ;
      RECT  90630.0 114655.0 90700.0 115822.5 ;
      RECT  90965.0 114655.0 91035.0 115822.5 ;
      RECT  91335.0 114777.5 91412.5 114912.5 ;
      RECT  91537.5 114777.5 91740.0 114912.5 ;
      RECT  91335.0 115307.5 91412.5 115442.5 ;
      RECT  91670.0 115307.5 91792.5 115442.5 ;
      RECT  91345.0 114777.5 91415.0 114912.5 ;
      RECT  91535.0 114777.5 91605.0 114912.5 ;
      RECT  91345.0 115307.5 91415.0 115442.5 ;
      RECT  91725.0 115307.5 91795.0 115442.5 ;
      RECT  91335.0 114655.0 91405.0 115822.5 ;
      RECT  91670.0 114655.0 91740.0 115822.5 ;
      RECT  92040.0 114777.5 92117.5 114912.5 ;
      RECT  92242.5 114777.5 92445.0 114912.5 ;
      RECT  92040.0 115307.5 92117.5 115442.5 ;
      RECT  92375.0 115307.5 92497.5 115442.5 ;
      RECT  92050.0 114777.5 92120.0 114912.5 ;
      RECT  92240.0 114777.5 92310.0 114912.5 ;
      RECT  92050.0 115307.5 92120.0 115442.5 ;
      RECT  92430.0 115307.5 92500.0 115442.5 ;
      RECT  92040.0 114655.0 92110.0 115822.5 ;
      RECT  92375.0 114655.0 92445.0 115822.5 ;
      RECT  92745.0 114777.5 92822.5 114912.5 ;
      RECT  92947.5 114777.5 93150.0 114912.5 ;
      RECT  92745.0 115307.5 92822.5 115442.5 ;
      RECT  93080.0 115307.5 93202.5 115442.5 ;
      RECT  92755.0 114777.5 92825.0 114912.5 ;
      RECT  92945.0 114777.5 93015.0 114912.5 ;
      RECT  92755.0 115307.5 92825.0 115442.5 ;
      RECT  93135.0 115307.5 93205.0 115442.5 ;
      RECT  92745.0 114655.0 92815.0 115822.5 ;
      RECT  93080.0 114655.0 93150.0 115822.5 ;
      RECT  93450.0 114777.5 93527.5 114912.5 ;
      RECT  93652.5 114777.5 93855.0 114912.5 ;
      RECT  93450.0 115307.5 93527.5 115442.5 ;
      RECT  93785.0 115307.5 93907.5 115442.5 ;
      RECT  93460.0 114777.5 93530.0 114912.5 ;
      RECT  93650.0 114777.5 93720.0 114912.5 ;
      RECT  93460.0 115307.5 93530.0 115442.5 ;
      RECT  93840.0 115307.5 93910.0 115442.5 ;
      RECT  93450.0 114655.0 93520.0 115822.5 ;
      RECT  93785.0 114655.0 93855.0 115822.5 ;
      RECT  94155.0 114777.5 94232.5 114912.5 ;
      RECT  94357.5 114777.5 94560.0 114912.5 ;
      RECT  94155.0 115307.5 94232.5 115442.5 ;
      RECT  94490.0 115307.5 94612.5 115442.5 ;
      RECT  94165.0 114777.5 94235.0 114912.5 ;
      RECT  94355.0 114777.5 94425.0 114912.5 ;
      RECT  94165.0 115307.5 94235.0 115442.5 ;
      RECT  94545.0 115307.5 94615.0 115442.5 ;
      RECT  94155.0 114655.0 94225.0 115822.5 ;
      RECT  94490.0 114655.0 94560.0 115822.5 ;
      RECT  94860.0 114777.5 94937.5 114912.5 ;
      RECT  95062.5 114777.5 95265.0 114912.5 ;
      RECT  94860.0 115307.5 94937.5 115442.5 ;
      RECT  95195.0 115307.5 95317.5 115442.5 ;
      RECT  94870.0 114777.5 94940.0 114912.5 ;
      RECT  95060.0 114777.5 95130.0 114912.5 ;
      RECT  94870.0 115307.5 94940.0 115442.5 ;
      RECT  95250.0 115307.5 95320.0 115442.5 ;
      RECT  94860.0 114655.0 94930.0 115822.5 ;
      RECT  95195.0 114655.0 95265.0 115822.5 ;
      RECT  95565.0 114777.5 95642.5 114912.5 ;
      RECT  95767.5 114777.5 95970.0 114912.5 ;
      RECT  95565.0 115307.5 95642.5 115442.5 ;
      RECT  95900.0 115307.5 96022.5 115442.5 ;
      RECT  95575.0 114777.5 95645.0 114912.5 ;
      RECT  95765.0 114777.5 95835.0 114912.5 ;
      RECT  95575.0 115307.5 95645.0 115442.5 ;
      RECT  95955.0 115307.5 96025.0 115442.5 ;
      RECT  95565.0 114655.0 95635.0 115822.5 ;
      RECT  95900.0 114655.0 95970.0 115822.5 ;
      RECT  96270.0 114777.5 96347.5 114912.5 ;
      RECT  96472.5 114777.5 96675.0 114912.5 ;
      RECT  96270.0 115307.5 96347.5 115442.5 ;
      RECT  96605.0 115307.5 96727.5 115442.5 ;
      RECT  96280.0 114777.5 96350.0 114912.5 ;
      RECT  96470.0 114777.5 96540.0 114912.5 ;
      RECT  96280.0 115307.5 96350.0 115442.5 ;
      RECT  96660.0 115307.5 96730.0 115442.5 ;
      RECT  96270.0 114655.0 96340.0 115822.5 ;
      RECT  96605.0 114655.0 96675.0 115822.5 ;
      RECT  96975.0 114777.5 97052.5 114912.5 ;
      RECT  97177.5 114777.5 97380.0 114912.5 ;
      RECT  96975.0 115307.5 97052.5 115442.5 ;
      RECT  97310.0 115307.5 97432.5 115442.5 ;
      RECT  96985.0 114777.5 97055.0 114912.5 ;
      RECT  97175.0 114777.5 97245.0 114912.5 ;
      RECT  96985.0 115307.5 97055.0 115442.5 ;
      RECT  97365.0 115307.5 97435.0 115442.5 ;
      RECT  96975.0 114655.0 97045.0 115822.5 ;
      RECT  97310.0 114655.0 97380.0 115822.5 ;
      RECT  97680.0 114777.5 97757.5 114912.5 ;
      RECT  97882.5 114777.5 98085.0 114912.5 ;
      RECT  97680.0 115307.5 97757.5 115442.5 ;
      RECT  98015.0 115307.5 98137.5 115442.5 ;
      RECT  97690.0 114777.5 97760.0 114912.5 ;
      RECT  97880.0 114777.5 97950.0 114912.5 ;
      RECT  97690.0 115307.5 97760.0 115442.5 ;
      RECT  98070.0 115307.5 98140.0 115442.5 ;
      RECT  97680.0 114655.0 97750.0 115822.5 ;
      RECT  98015.0 114655.0 98085.0 115822.5 ;
      RECT  98385.0 114777.5 98462.5 114912.5 ;
      RECT  98587.5 114777.5 98790.0 114912.5 ;
      RECT  98385.0 115307.5 98462.5 115442.5 ;
      RECT  98720.0 115307.5 98842.5 115442.5 ;
      RECT  98395.0 114777.5 98465.0 114912.5 ;
      RECT  98585.0 114777.5 98655.0 114912.5 ;
      RECT  98395.0 115307.5 98465.0 115442.5 ;
      RECT  98775.0 115307.5 98845.0 115442.5 ;
      RECT  98385.0 114655.0 98455.0 115822.5 ;
      RECT  98720.0 114655.0 98790.0 115822.5 ;
      RECT  99090.0 114777.5 99167.5 114912.5 ;
      RECT  99292.5 114777.5 99495.0 114912.5 ;
      RECT  99090.0 115307.5 99167.5 115442.5 ;
      RECT  99425.0 115307.5 99547.5 115442.5 ;
      RECT  99100.0 114777.5 99170.0 114912.5 ;
      RECT  99290.0 114777.5 99360.0 114912.5 ;
      RECT  99100.0 115307.5 99170.0 115442.5 ;
      RECT  99480.0 115307.5 99550.0 115442.5 ;
      RECT  99090.0 114655.0 99160.0 115822.5 ;
      RECT  99425.0 114655.0 99495.0 115822.5 ;
      RECT  99795.0 114777.5 99872.5 114912.5 ;
      RECT  99997.5 114777.5 100200.0 114912.5 ;
      RECT  99795.0 115307.5 99872.5 115442.5 ;
      RECT  100130.0 115307.5 100252.5 115442.5 ;
      RECT  99805.0 114777.5 99875.0 114912.5 ;
      RECT  99995.0 114777.5 100065.0 114912.5 ;
      RECT  99805.0 115307.5 99875.0 115442.5 ;
      RECT  100185.0 115307.5 100255.0 115442.5 ;
      RECT  99795.0 114655.0 99865.0 115822.5 ;
      RECT  100130.0 114655.0 100200.0 115822.5 ;
      RECT  100500.0 114777.5 100577.5 114912.5 ;
      RECT  100702.5 114777.5 100905.0 114912.5 ;
      RECT  100500.0 115307.5 100577.5 115442.5 ;
      RECT  100835.0 115307.5 100957.5 115442.5 ;
      RECT  100510.0 114777.5 100580.0 114912.5 ;
      RECT  100700.0 114777.5 100770.0 114912.5 ;
      RECT  100510.0 115307.5 100580.0 115442.5 ;
      RECT  100890.0 115307.5 100960.0 115442.5 ;
      RECT  100500.0 114655.0 100570.0 115822.5 ;
      RECT  100835.0 114655.0 100905.0 115822.5 ;
      RECT  101205.0 114777.5 101282.5 114912.5 ;
      RECT  101407.5 114777.5 101610.0 114912.5 ;
      RECT  101205.0 115307.5 101282.5 115442.5 ;
      RECT  101540.0 115307.5 101662.5 115442.5 ;
      RECT  101215.0 114777.5 101285.0 114912.5 ;
      RECT  101405.0 114777.5 101475.0 114912.5 ;
      RECT  101215.0 115307.5 101285.0 115442.5 ;
      RECT  101595.0 115307.5 101665.0 115442.5 ;
      RECT  101205.0 114655.0 101275.0 115822.5 ;
      RECT  101540.0 114655.0 101610.0 115822.5 ;
      RECT  101910.0 114777.5 101987.5 114912.5 ;
      RECT  102112.5 114777.5 102315.0 114912.5 ;
      RECT  101910.0 115307.5 101987.5 115442.5 ;
      RECT  102245.0 115307.5 102367.5 115442.5 ;
      RECT  101920.0 114777.5 101990.0 114912.5 ;
      RECT  102110.0 114777.5 102180.0 114912.5 ;
      RECT  101920.0 115307.5 101990.0 115442.5 ;
      RECT  102300.0 115307.5 102370.0 115442.5 ;
      RECT  101910.0 114655.0 101980.0 115822.5 ;
      RECT  102245.0 114655.0 102315.0 115822.5 ;
      RECT  102615.0 114777.5 102692.5 114912.5 ;
      RECT  102817.5 114777.5 103020.0 114912.5 ;
      RECT  102615.0 115307.5 102692.5 115442.5 ;
      RECT  102950.0 115307.5 103072.5 115442.5 ;
      RECT  102625.0 114777.5 102695.0 114912.5 ;
      RECT  102815.0 114777.5 102885.0 114912.5 ;
      RECT  102625.0 115307.5 102695.0 115442.5 ;
      RECT  103005.0 115307.5 103075.0 115442.5 ;
      RECT  102615.0 114655.0 102685.0 115822.5 ;
      RECT  102950.0 114655.0 103020.0 115822.5 ;
      RECT  103320.0 114777.5 103397.5 114912.5 ;
      RECT  103522.5 114777.5 103725.0 114912.5 ;
      RECT  103320.0 115307.5 103397.5 115442.5 ;
      RECT  103655.0 115307.5 103777.5 115442.5 ;
      RECT  103330.0 114777.5 103400.0 114912.5 ;
      RECT  103520.0 114777.5 103590.0 114912.5 ;
      RECT  103330.0 115307.5 103400.0 115442.5 ;
      RECT  103710.0 115307.5 103780.0 115442.5 ;
      RECT  103320.0 114655.0 103390.0 115822.5 ;
      RECT  103655.0 114655.0 103725.0 115822.5 ;
      RECT  104025.0 114777.5 104102.5 114912.5 ;
      RECT  104227.5 114777.5 104430.0 114912.5 ;
      RECT  104025.0 115307.5 104102.5 115442.5 ;
      RECT  104360.0 115307.5 104482.5 115442.5 ;
      RECT  104035.0 114777.5 104105.0 114912.5 ;
      RECT  104225.0 114777.5 104295.0 114912.5 ;
      RECT  104035.0 115307.5 104105.0 115442.5 ;
      RECT  104415.0 115307.5 104485.0 115442.5 ;
      RECT  104025.0 114655.0 104095.0 115822.5 ;
      RECT  104360.0 114655.0 104430.0 115822.5 ;
      RECT  104730.0 114777.5 104807.5 114912.5 ;
      RECT  104932.5 114777.5 105135.0 114912.5 ;
      RECT  104730.0 115307.5 104807.5 115442.5 ;
      RECT  105065.0 115307.5 105187.5 115442.5 ;
      RECT  104740.0 114777.5 104810.0 114912.5 ;
      RECT  104930.0 114777.5 105000.0 114912.5 ;
      RECT  104740.0 115307.5 104810.0 115442.5 ;
      RECT  105120.0 115307.5 105190.0 115442.5 ;
      RECT  104730.0 114655.0 104800.0 115822.5 ;
      RECT  105065.0 114655.0 105135.0 115822.5 ;
      RECT  105435.0 114777.5 105512.5 114912.5 ;
      RECT  105637.5 114777.5 105840.0 114912.5 ;
      RECT  105435.0 115307.5 105512.5 115442.5 ;
      RECT  105770.0 115307.5 105892.5 115442.5 ;
      RECT  105445.0 114777.5 105515.0 114912.5 ;
      RECT  105635.0 114777.5 105705.0 114912.5 ;
      RECT  105445.0 115307.5 105515.0 115442.5 ;
      RECT  105825.0 115307.5 105895.0 115442.5 ;
      RECT  105435.0 114655.0 105505.0 115822.5 ;
      RECT  105770.0 114655.0 105840.0 115822.5 ;
      RECT  15900.0 114655.0 15970.0 115822.5 ;
      RECT  16235.0 114655.0 16305.0 115822.5 ;
      RECT  16605.0 114655.0 16675.0 115822.5 ;
      RECT  16940.0 114655.0 17010.0 115822.5 ;
      RECT  17310.0 114655.0 17380.0 115822.5 ;
      RECT  17645.0 114655.0 17715.0 115822.5 ;
      RECT  18015.0 114655.0 18085.0 115822.5 ;
      RECT  18350.0 114655.0 18420.0 115822.5 ;
      RECT  18720.0 114655.0 18790.0 115822.5 ;
      RECT  19055.0 114655.0 19125.0 115822.5 ;
      RECT  19425.0 114655.0 19495.0 115822.5 ;
      RECT  19760.0 114655.0 19830.0 115822.5 ;
      RECT  20130.0 114655.0 20200.0 115822.5 ;
      RECT  20465.0 114655.0 20535.0 115822.5 ;
      RECT  20835.0 114655.0 20905.0 115822.5 ;
      RECT  21170.0 114655.0 21240.0 115822.5 ;
      RECT  21540.0 114655.0 21610.0 115822.5 ;
      RECT  21875.0 114655.0 21945.0 115822.5 ;
      RECT  22245.0 114655.0 22315.0 115822.5 ;
      RECT  22580.0 114655.0 22650.0 115822.5 ;
      RECT  22950.0 114655.0 23020.0 115822.5 ;
      RECT  23285.0 114655.0 23355.0 115822.5 ;
      RECT  23655.0 114655.0 23725.0 115822.5 ;
      RECT  23990.0 114655.0 24060.0 115822.5 ;
      RECT  24360.0 114655.0 24430.0 115822.5 ;
      RECT  24695.0 114655.0 24765.0 115822.5 ;
      RECT  25065.0 114655.0 25135.0 115822.5 ;
      RECT  25400.0 114655.0 25470.0 115822.5 ;
      RECT  25770.0 114655.0 25840.0 115822.5 ;
      RECT  26105.0 114655.0 26175.0 115822.5 ;
      RECT  26475.0 114655.0 26545.0 115822.5 ;
      RECT  26810.0 114655.0 26880.0 115822.5 ;
      RECT  27180.0 114655.0 27250.0 115822.5 ;
      RECT  27515.0 114655.0 27585.0 115822.5 ;
      RECT  27885.0 114655.0 27955.0 115822.5 ;
      RECT  28220.0 114655.0 28290.0 115822.5 ;
      RECT  28590.0 114655.0 28660.0 115822.5 ;
      RECT  28925.0 114655.0 28995.0 115822.5 ;
      RECT  29295.0 114655.0 29365.0 115822.5 ;
      RECT  29630.0 114655.0 29700.0 115822.5 ;
      RECT  30000.0 114655.0 30070.0 115822.5 ;
      RECT  30335.0 114655.0 30405.0 115822.5 ;
      RECT  30705.0 114655.0 30775.0 115822.5 ;
      RECT  31040.0 114655.0 31110.0 115822.5 ;
      RECT  31410.0 114655.0 31480.0 115822.5 ;
      RECT  31745.0 114655.0 31815.0 115822.5 ;
      RECT  32115.0 114655.0 32185.0 115822.5 ;
      RECT  32450.0 114655.0 32520.0 115822.5 ;
      RECT  32820.0 114655.0 32890.0 115822.5 ;
      RECT  33155.0 114655.0 33225.0 115822.5 ;
      RECT  33525.0 114655.0 33595.0 115822.5 ;
      RECT  33860.0 114655.0 33930.0 115822.5 ;
      RECT  34230.0 114655.0 34300.0 115822.5 ;
      RECT  34565.0 114655.0 34635.0 115822.5 ;
      RECT  34935.0 114655.0 35005.0 115822.5 ;
      RECT  35270.0 114655.0 35340.0 115822.5 ;
      RECT  35640.0 114655.0 35710.0 115822.5 ;
      RECT  35975.0 114655.0 36045.0 115822.5 ;
      RECT  36345.0 114655.0 36415.0 115822.5 ;
      RECT  36680.0 114655.0 36750.0 115822.5 ;
      RECT  37050.0 114655.0 37120.0 115822.5 ;
      RECT  37385.0 114655.0 37455.0 115822.5 ;
      RECT  37755.0 114655.0 37825.0 115822.5 ;
      RECT  38090.0 114655.0 38160.0 115822.5 ;
      RECT  38460.0 114655.0 38530.0 115822.5 ;
      RECT  38795.0 114655.0 38865.0 115822.5 ;
      RECT  39165.0 114655.0 39235.0 115822.5 ;
      RECT  39500.0 114655.0 39570.0 115822.5 ;
      RECT  39870.0 114655.0 39940.0 115822.5 ;
      RECT  40205.0 114655.0 40275.0 115822.5 ;
      RECT  40575.0 114655.0 40645.0 115822.5 ;
      RECT  40910.0 114655.0 40980.0 115822.5 ;
      RECT  41280.0 114655.0 41350.0 115822.5 ;
      RECT  41615.0 114655.0 41685.0 115822.5 ;
      RECT  41985.0 114655.0 42055.0 115822.5 ;
      RECT  42320.0 114655.0 42390.0 115822.5 ;
      RECT  42690.0 114655.0 42760.0 115822.5 ;
      RECT  43025.0 114655.0 43095.0 115822.5 ;
      RECT  43395.0 114655.0 43465.0 115822.5 ;
      RECT  43730.0 114655.0 43800.0 115822.5 ;
      RECT  44100.0 114655.0 44170.0 115822.5 ;
      RECT  44435.0 114655.0 44505.0 115822.5 ;
      RECT  44805.0 114655.0 44875.0 115822.5 ;
      RECT  45140.0 114655.0 45210.0 115822.5 ;
      RECT  45510.0 114655.0 45580.0 115822.5 ;
      RECT  45845.0 114655.0 45915.0 115822.5 ;
      RECT  46215.0 114655.0 46285.0 115822.5 ;
      RECT  46550.0 114655.0 46620.0 115822.5 ;
      RECT  46920.0 114655.0 46990.0 115822.5 ;
      RECT  47255.0 114655.0 47325.0 115822.5 ;
      RECT  47625.0 114655.0 47695.0 115822.5 ;
      RECT  47960.0 114655.0 48030.0 115822.5 ;
      RECT  48330.0 114655.0 48400.0 115822.5 ;
      RECT  48665.0 114655.0 48735.0 115822.5 ;
      RECT  49035.0 114655.0 49105.0 115822.5 ;
      RECT  49370.0 114655.0 49440.0 115822.5 ;
      RECT  49740.0 114655.0 49810.0 115822.5 ;
      RECT  50075.0 114655.0 50145.0 115822.5 ;
      RECT  50445.0 114655.0 50515.0 115822.5 ;
      RECT  50780.0 114655.0 50850.0 115822.5 ;
      RECT  51150.0 114655.0 51220.0 115822.5 ;
      RECT  51485.0 114655.0 51555.0 115822.5 ;
      RECT  51855.0 114655.0 51925.0 115822.5 ;
      RECT  52190.0 114655.0 52260.0 115822.5 ;
      RECT  52560.0 114655.0 52630.0 115822.5 ;
      RECT  52895.0 114655.0 52965.0 115822.5 ;
      RECT  53265.0 114655.0 53335.0 115822.5 ;
      RECT  53600.0 114655.0 53670.0 115822.5 ;
      RECT  53970.0 114655.0 54040.0 115822.5 ;
      RECT  54305.0 114655.0 54375.0 115822.5 ;
      RECT  54675.0 114655.0 54745.0 115822.5 ;
      RECT  55010.0 114655.0 55080.0 115822.5 ;
      RECT  55380.0 114655.0 55450.0 115822.5 ;
      RECT  55715.0 114655.0 55785.0 115822.5 ;
      RECT  56085.0 114655.0 56155.0 115822.5 ;
      RECT  56420.0 114655.0 56490.0 115822.5 ;
      RECT  56790.0 114655.0 56860.0 115822.5 ;
      RECT  57125.0 114655.0 57195.0 115822.5 ;
      RECT  57495.0 114655.0 57565.0 115822.5 ;
      RECT  57830.0 114655.0 57900.0 115822.5 ;
      RECT  58200.0 114655.0 58270.0 115822.5 ;
      RECT  58535.0 114655.0 58605.0 115822.5 ;
      RECT  58905.0 114655.0 58975.0 115822.5 ;
      RECT  59240.0 114655.0 59310.0 115822.5 ;
      RECT  59610.0 114655.0 59680.0 115822.5 ;
      RECT  59945.0 114655.0 60015.0 115822.5 ;
      RECT  60315.0 114655.0 60385.0 115822.5 ;
      RECT  60650.0 114655.0 60720.0 115822.5 ;
      RECT  61020.0 114655.0 61090.0 115822.5 ;
      RECT  61355.0 114655.0 61425.0 115822.5 ;
      RECT  61725.0 114655.0 61795.0 115822.5 ;
      RECT  62060.0 114655.0 62130.0 115822.5 ;
      RECT  62430.0 114655.0 62500.0 115822.5 ;
      RECT  62765.0 114655.0 62835.0 115822.5 ;
      RECT  63135.0 114655.0 63205.0 115822.5 ;
      RECT  63470.0 114655.0 63540.0 115822.5 ;
      RECT  63840.0 114655.0 63910.0 115822.5 ;
      RECT  64175.0 114655.0 64245.0 115822.5 ;
      RECT  64545.0 114655.0 64615.0 115822.5 ;
      RECT  64880.0 114655.0 64950.0 115822.5 ;
      RECT  65250.0 114655.0 65320.0 115822.5 ;
      RECT  65585.0 114655.0 65655.0 115822.5 ;
      RECT  65955.0 114655.0 66025.0 115822.5 ;
      RECT  66290.0 114655.0 66360.0 115822.5 ;
      RECT  66660.0 114655.0 66730.0 115822.5 ;
      RECT  66995.0 114655.0 67065.0 115822.5 ;
      RECT  67365.0 114655.0 67435.0 115822.5 ;
      RECT  67700.0 114655.0 67770.0 115822.5 ;
      RECT  68070.0 114655.0 68140.0 115822.5 ;
      RECT  68405.0 114655.0 68475.0 115822.5 ;
      RECT  68775.0 114655.0 68845.0 115822.5 ;
      RECT  69110.0 114655.0 69180.0 115822.5 ;
      RECT  69480.0 114655.0 69550.0 115822.5 ;
      RECT  69815.0 114655.0 69885.0 115822.5 ;
      RECT  70185.0 114655.0 70255.0 115822.5 ;
      RECT  70520.0 114655.0 70590.0 115822.5 ;
      RECT  70890.0 114655.0 70960.0 115822.5 ;
      RECT  71225.0 114655.0 71295.0 115822.5 ;
      RECT  71595.0 114655.0 71665.0 115822.5 ;
      RECT  71930.0 114655.0 72000.0 115822.5 ;
      RECT  72300.0 114655.0 72370.0 115822.5 ;
      RECT  72635.0 114655.0 72705.0 115822.5 ;
      RECT  73005.0 114655.0 73075.0 115822.5 ;
      RECT  73340.0 114655.0 73410.0 115822.5 ;
      RECT  73710.0 114655.0 73780.0 115822.5 ;
      RECT  74045.0 114655.0 74115.0 115822.5 ;
      RECT  74415.0 114655.0 74485.0 115822.5 ;
      RECT  74750.0 114655.0 74820.0 115822.5 ;
      RECT  75120.0 114655.0 75190.0 115822.5 ;
      RECT  75455.0 114655.0 75525.0 115822.5 ;
      RECT  75825.0 114655.0 75895.0 115822.5 ;
      RECT  76160.0 114655.0 76230.0 115822.5 ;
      RECT  76530.0 114655.0 76600.0 115822.5 ;
      RECT  76865.0 114655.0 76935.0 115822.5 ;
      RECT  77235.0 114655.0 77305.0 115822.5 ;
      RECT  77570.0 114655.0 77640.0 115822.5 ;
      RECT  77940.0 114655.0 78010.0 115822.5 ;
      RECT  78275.0 114655.0 78345.0 115822.5 ;
      RECT  78645.0 114655.0 78715.0 115822.5 ;
      RECT  78980.0 114655.0 79050.0 115822.5 ;
      RECT  79350.0 114655.0 79420.0 115822.5 ;
      RECT  79685.0 114655.0 79755.0 115822.5 ;
      RECT  80055.0 114655.0 80125.0 115822.5 ;
      RECT  80390.0 114655.0 80460.0 115822.5 ;
      RECT  80760.0 114655.0 80830.0 115822.5 ;
      RECT  81095.0 114655.0 81165.0 115822.5 ;
      RECT  81465.0 114655.0 81535.0 115822.5 ;
      RECT  81800.0 114655.0 81870.0 115822.5 ;
      RECT  82170.0 114655.0 82240.0 115822.5 ;
      RECT  82505.0 114655.0 82575.0 115822.5 ;
      RECT  82875.0 114655.0 82945.0 115822.5 ;
      RECT  83210.0 114655.0 83280.0 115822.5 ;
      RECT  83580.0 114655.0 83650.0 115822.5 ;
      RECT  83915.0 114655.0 83985.0 115822.5 ;
      RECT  84285.0 114655.0 84355.0 115822.5 ;
      RECT  84620.0 114655.0 84690.0 115822.5 ;
      RECT  84990.0 114655.0 85060.0 115822.5 ;
      RECT  85325.0 114655.0 85395.0 115822.5 ;
      RECT  85695.0 114655.0 85765.0 115822.5 ;
      RECT  86030.0 114655.0 86100.0 115822.5 ;
      RECT  86400.0 114655.0 86470.0 115822.5 ;
      RECT  86735.0 114655.0 86805.0 115822.5 ;
      RECT  87105.0 114655.0 87175.0 115822.5 ;
      RECT  87440.0 114655.0 87510.0 115822.5 ;
      RECT  87810.0 114655.0 87880.0 115822.5 ;
      RECT  88145.0 114655.0 88215.0 115822.5 ;
      RECT  88515.0 114655.0 88585.0 115822.5 ;
      RECT  88850.0 114655.0 88920.0 115822.5 ;
      RECT  89220.0 114655.0 89290.0 115822.5 ;
      RECT  89555.0 114655.0 89625.0 115822.5 ;
      RECT  89925.0 114655.0 89995.0 115822.5 ;
      RECT  90260.0 114655.0 90330.0 115822.5 ;
      RECT  90630.0 114655.0 90700.0 115822.5 ;
      RECT  90965.0 114655.0 91035.0 115822.5 ;
      RECT  91335.0 114655.0 91405.0 115822.5 ;
      RECT  91670.0 114655.0 91740.0 115822.5 ;
      RECT  92040.0 114655.0 92110.0 115822.5 ;
      RECT  92375.0 114655.0 92445.0 115822.5 ;
      RECT  92745.0 114655.0 92815.0 115822.5 ;
      RECT  93080.0 114655.0 93150.0 115822.5 ;
      RECT  93450.0 114655.0 93520.0 115822.5 ;
      RECT  93785.0 114655.0 93855.0 115822.5 ;
      RECT  94155.0 114655.0 94225.0 115822.5 ;
      RECT  94490.0 114655.0 94560.0 115822.5 ;
      RECT  94860.0 114655.0 94930.0 115822.5 ;
      RECT  95195.0 114655.0 95265.0 115822.5 ;
      RECT  95565.0 114655.0 95635.0 115822.5 ;
      RECT  95900.0 114655.0 95970.0 115822.5 ;
      RECT  96270.0 114655.0 96340.0 115822.5 ;
      RECT  96605.0 114655.0 96675.0 115822.5 ;
      RECT  96975.0 114655.0 97045.0 115822.5 ;
      RECT  97310.0 114655.0 97380.0 115822.5 ;
      RECT  97680.0 114655.0 97750.0 115822.5 ;
      RECT  98015.0 114655.0 98085.0 115822.5 ;
      RECT  98385.0 114655.0 98455.0 115822.5 ;
      RECT  98720.0 114655.0 98790.0 115822.5 ;
      RECT  99090.0 114655.0 99160.0 115822.5 ;
      RECT  99425.0 114655.0 99495.0 115822.5 ;
      RECT  99795.0 114655.0 99865.0 115822.5 ;
      RECT  100130.0 114655.0 100200.0 115822.5 ;
      RECT  100500.0 114655.0 100570.0 115822.5 ;
      RECT  100835.0 114655.0 100905.0 115822.5 ;
      RECT  101205.0 114655.0 101275.0 115822.5 ;
      RECT  101540.0 114655.0 101610.0 115822.5 ;
      RECT  101910.0 114655.0 101980.0 115822.5 ;
      RECT  102245.0 114655.0 102315.0 115822.5 ;
      RECT  102615.0 114655.0 102685.0 115822.5 ;
      RECT  102950.0 114655.0 103020.0 115822.5 ;
      RECT  103320.0 114655.0 103390.0 115822.5 ;
      RECT  103655.0 114655.0 103725.0 115822.5 ;
      RECT  104025.0 114655.0 104095.0 115822.5 ;
      RECT  104360.0 114655.0 104430.0 115822.5 ;
      RECT  104730.0 114655.0 104800.0 115822.5 ;
      RECT  105065.0 114655.0 105135.0 115822.5 ;
      RECT  105435.0 114655.0 105505.0 115822.5 ;
      RECT  105770.0 114655.0 105840.0 115822.5 ;
      RECT  16605.0 25450.0 16675.0 26150.0 ;
      RECT  16940.0 25310.0 17010.0 26150.0 ;
      RECT  17310.0 25450.0 17380.0 26150.0 ;
      RECT  17645.0 25310.0 17715.0 26150.0 ;
      RECT  18015.0 25450.0 18085.0 26150.0 ;
      RECT  18350.0 25310.0 18420.0 26150.0 ;
      RECT  19425.0 25450.0 19495.0 26150.0 ;
      RECT  19760.0 25310.0 19830.0 26150.0 ;
      RECT  20130.0 25450.0 20200.0 26150.0 ;
      RECT  20465.0 25310.0 20535.0 26150.0 ;
      RECT  20835.0 25450.0 20905.0 26150.0 ;
      RECT  21170.0 25310.0 21240.0 26150.0 ;
      RECT  22245.0 25450.0 22315.0 26150.0 ;
      RECT  22580.0 25310.0 22650.0 26150.0 ;
      RECT  22950.0 25450.0 23020.0 26150.0 ;
      RECT  23285.0 25310.0 23355.0 26150.0 ;
      RECT  23655.0 25450.0 23725.0 26150.0 ;
      RECT  23990.0 25310.0 24060.0 26150.0 ;
      RECT  25065.0 25450.0 25135.0 26150.0 ;
      RECT  25400.0 25310.0 25470.0 26150.0 ;
      RECT  25770.0 25450.0 25840.0 26150.0 ;
      RECT  26105.0 25310.0 26175.0 26150.0 ;
      RECT  26475.0 25450.0 26545.0 26150.0 ;
      RECT  26810.0 25310.0 26880.0 26150.0 ;
      RECT  27885.0 25450.0 27955.0 26150.0 ;
      RECT  28220.0 25310.0 28290.0 26150.0 ;
      RECT  28590.0 25450.0 28660.0 26150.0 ;
      RECT  28925.0 25310.0 28995.0 26150.0 ;
      RECT  29295.0 25450.0 29365.0 26150.0 ;
      RECT  29630.0 25310.0 29700.0 26150.0 ;
      RECT  30705.0 25450.0 30775.0 26150.0 ;
      RECT  31040.0 25310.0 31110.0 26150.0 ;
      RECT  31410.0 25450.0 31480.0 26150.0 ;
      RECT  31745.0 25310.0 31815.0 26150.0 ;
      RECT  32115.0 25450.0 32185.0 26150.0 ;
      RECT  32450.0 25310.0 32520.0 26150.0 ;
      RECT  33525.0 25450.0 33595.0 26150.0 ;
      RECT  33860.0 25310.0 33930.0 26150.0 ;
      RECT  34230.0 25450.0 34300.0 26150.0 ;
      RECT  34565.0 25310.0 34635.0 26150.0 ;
      RECT  34935.0 25450.0 35005.0 26150.0 ;
      RECT  35270.0 25310.0 35340.0 26150.0 ;
      RECT  36345.0 25450.0 36415.0 26150.0 ;
      RECT  36680.0 25310.0 36750.0 26150.0 ;
      RECT  37050.0 25450.0 37120.0 26150.0 ;
      RECT  37385.0 25310.0 37455.0 26150.0 ;
      RECT  37755.0 25450.0 37825.0 26150.0 ;
      RECT  38090.0 25310.0 38160.0 26150.0 ;
      RECT  39165.0 25450.0 39235.0 26150.0 ;
      RECT  39500.0 25310.0 39570.0 26150.0 ;
      RECT  39870.0 25450.0 39940.0 26150.0 ;
      RECT  40205.0 25310.0 40275.0 26150.0 ;
      RECT  40575.0 25450.0 40645.0 26150.0 ;
      RECT  40910.0 25310.0 40980.0 26150.0 ;
      RECT  41985.0 25450.0 42055.0 26150.0 ;
      RECT  42320.0 25310.0 42390.0 26150.0 ;
      RECT  42690.0 25450.0 42760.0 26150.0 ;
      RECT  43025.0 25310.0 43095.0 26150.0 ;
      RECT  43395.0 25450.0 43465.0 26150.0 ;
      RECT  43730.0 25310.0 43800.0 26150.0 ;
      RECT  44805.0 25450.0 44875.0 26150.0 ;
      RECT  45140.0 25310.0 45210.0 26150.0 ;
      RECT  45510.0 25450.0 45580.0 26150.0 ;
      RECT  45845.0 25310.0 45915.0 26150.0 ;
      RECT  46215.0 25450.0 46285.0 26150.0 ;
      RECT  46550.0 25310.0 46620.0 26150.0 ;
      RECT  47625.0 25450.0 47695.0 26150.0 ;
      RECT  47960.0 25310.0 48030.0 26150.0 ;
      RECT  48330.0 25450.0 48400.0 26150.0 ;
      RECT  48665.0 25310.0 48735.0 26150.0 ;
      RECT  49035.0 25450.0 49105.0 26150.0 ;
      RECT  49370.0 25310.0 49440.0 26150.0 ;
      RECT  50445.0 25450.0 50515.0 26150.0 ;
      RECT  50780.0 25310.0 50850.0 26150.0 ;
      RECT  51150.0 25450.0 51220.0 26150.0 ;
      RECT  51485.0 25310.0 51555.0 26150.0 ;
      RECT  51855.0 25450.0 51925.0 26150.0 ;
      RECT  52190.0 25310.0 52260.0 26150.0 ;
      RECT  53265.0 25450.0 53335.0 26150.0 ;
      RECT  53600.0 25310.0 53670.0 26150.0 ;
      RECT  53970.0 25450.0 54040.0 26150.0 ;
      RECT  54305.0 25310.0 54375.0 26150.0 ;
      RECT  54675.0 25450.0 54745.0 26150.0 ;
      RECT  55010.0 25310.0 55080.0 26150.0 ;
      RECT  56085.0 25450.0 56155.0 26150.0 ;
      RECT  56420.0 25310.0 56490.0 26150.0 ;
      RECT  56790.0 25450.0 56860.0 26150.0 ;
      RECT  57125.0 25310.0 57195.0 26150.0 ;
      RECT  57495.0 25450.0 57565.0 26150.0 ;
      RECT  57830.0 25310.0 57900.0 26150.0 ;
      RECT  58905.0 25450.0 58975.0 26150.0 ;
      RECT  59240.0 25310.0 59310.0 26150.0 ;
      RECT  59610.0 25450.0 59680.0 26150.0 ;
      RECT  59945.0 25310.0 60015.0 26150.0 ;
      RECT  60315.0 25450.0 60385.0 26150.0 ;
      RECT  60650.0 25310.0 60720.0 26150.0 ;
      RECT  61725.0 25450.0 61795.0 26150.0 ;
      RECT  62060.0 25310.0 62130.0 26150.0 ;
      RECT  62430.0 25450.0 62500.0 26150.0 ;
      RECT  62765.0 25310.0 62835.0 26150.0 ;
      RECT  63135.0 25450.0 63205.0 26150.0 ;
      RECT  63470.0 25310.0 63540.0 26150.0 ;
      RECT  64545.0 25450.0 64615.0 26150.0 ;
      RECT  64880.0 25310.0 64950.0 26150.0 ;
      RECT  65250.0 25450.0 65320.0 26150.0 ;
      RECT  65585.0 25310.0 65655.0 26150.0 ;
      RECT  65955.0 25450.0 66025.0 26150.0 ;
      RECT  66290.0 25310.0 66360.0 26150.0 ;
      RECT  67365.0 25450.0 67435.0 26150.0 ;
      RECT  67700.0 25310.0 67770.0 26150.0 ;
      RECT  68070.0 25450.0 68140.0 26150.0 ;
      RECT  68405.0 25310.0 68475.0 26150.0 ;
      RECT  68775.0 25450.0 68845.0 26150.0 ;
      RECT  69110.0 25310.0 69180.0 26150.0 ;
      RECT  70185.0 25450.0 70255.0 26150.0 ;
      RECT  70520.0 25310.0 70590.0 26150.0 ;
      RECT  70890.0 25450.0 70960.0 26150.0 ;
      RECT  71225.0 25310.0 71295.0 26150.0 ;
      RECT  71595.0 25450.0 71665.0 26150.0 ;
      RECT  71930.0 25310.0 72000.0 26150.0 ;
      RECT  73005.0 25450.0 73075.0 26150.0 ;
      RECT  73340.0 25310.0 73410.0 26150.0 ;
      RECT  73710.0 25450.0 73780.0 26150.0 ;
      RECT  74045.0 25310.0 74115.0 26150.0 ;
      RECT  74415.0 25450.0 74485.0 26150.0 ;
      RECT  74750.0 25310.0 74820.0 26150.0 ;
      RECT  75825.0 25450.0 75895.0 26150.0 ;
      RECT  76160.0 25310.0 76230.0 26150.0 ;
      RECT  76530.0 25450.0 76600.0 26150.0 ;
      RECT  76865.0 25310.0 76935.0 26150.0 ;
      RECT  77235.0 25450.0 77305.0 26150.0 ;
      RECT  77570.0 25310.0 77640.0 26150.0 ;
      RECT  78645.0 25450.0 78715.0 26150.0 ;
      RECT  78980.0 25310.0 79050.0 26150.0 ;
      RECT  79350.0 25450.0 79420.0 26150.0 ;
      RECT  79685.0 25310.0 79755.0 26150.0 ;
      RECT  80055.0 25450.0 80125.0 26150.0 ;
      RECT  80390.0 25310.0 80460.0 26150.0 ;
      RECT  81465.0 25450.0 81535.0 26150.0 ;
      RECT  81800.0 25310.0 81870.0 26150.0 ;
      RECT  82170.0 25450.0 82240.0 26150.0 ;
      RECT  82505.0 25310.0 82575.0 26150.0 ;
      RECT  82875.0 25450.0 82945.0 26150.0 ;
      RECT  83210.0 25310.0 83280.0 26150.0 ;
      RECT  84285.0 25450.0 84355.0 26150.0 ;
      RECT  84620.0 25310.0 84690.0 26150.0 ;
      RECT  84990.0 25450.0 85060.0 26150.0 ;
      RECT  85325.0 25310.0 85395.0 26150.0 ;
      RECT  85695.0 25450.0 85765.0 26150.0 ;
      RECT  86030.0 25310.0 86100.0 26150.0 ;
      RECT  87105.0 25450.0 87175.0 26150.0 ;
      RECT  87440.0 25310.0 87510.0 26150.0 ;
      RECT  87810.0 25450.0 87880.0 26150.0 ;
      RECT  88145.0 25310.0 88215.0 26150.0 ;
      RECT  88515.0 25450.0 88585.0 26150.0 ;
      RECT  88850.0 25310.0 88920.0 26150.0 ;
      RECT  89925.0 25450.0 89995.0 26150.0 ;
      RECT  90260.0 25310.0 90330.0 26150.0 ;
      RECT  90630.0 25450.0 90700.0 26150.0 ;
      RECT  90965.0 25310.0 91035.0 26150.0 ;
      RECT  91335.0 25450.0 91405.0 26150.0 ;
      RECT  91670.0 25310.0 91740.0 26150.0 ;
      RECT  92745.0 25450.0 92815.0 26150.0 ;
      RECT  93080.0 25310.0 93150.0 26150.0 ;
      RECT  93450.0 25450.0 93520.0 26150.0 ;
      RECT  93785.0 25310.0 93855.0 26150.0 ;
      RECT  94155.0 25450.0 94225.0 26150.0 ;
      RECT  94490.0 25310.0 94560.0 26150.0 ;
      RECT  95565.0 25450.0 95635.0 26150.0 ;
      RECT  95900.0 25310.0 95970.0 26150.0 ;
      RECT  96270.0 25450.0 96340.0 26150.0 ;
      RECT  96605.0 25310.0 96675.0 26150.0 ;
      RECT  96975.0 25450.0 97045.0 26150.0 ;
      RECT  97310.0 25310.0 97380.0 26150.0 ;
      RECT  98385.0 25450.0 98455.0 26150.0 ;
      RECT  98720.0 25310.0 98790.0 26150.0 ;
      RECT  99090.0 25450.0 99160.0 26150.0 ;
      RECT  99425.0 25310.0 99495.0 26150.0 ;
      RECT  99795.0 25450.0 99865.0 26150.0 ;
      RECT  100130.0 25310.0 100200.0 26150.0 ;
      RECT  101205.0 25450.0 101275.0 26150.0 ;
      RECT  101540.0 25310.0 101610.0 26150.0 ;
      RECT  101910.0 25450.0 101980.0 26150.0 ;
      RECT  102245.0 25310.0 102315.0 26150.0 ;
      RECT  102615.0 25450.0 102685.0 26150.0 ;
      RECT  102950.0 25310.0 103020.0 26150.0 ;
      RECT  104025.0 25450.0 104095.0 26150.0 ;
      RECT  104360.0 25310.0 104430.0 26150.0 ;
      RECT  104730.0 25450.0 104800.0 26150.0 ;
      RECT  105065.0 25310.0 105135.0 26150.0 ;
      RECT  105435.0 25450.0 105505.0 26150.0 ;
      RECT  105770.0 25310.0 105840.0 26150.0 ;
      RECT  15900.0 26790.0 15970.0 26860.0 ;
      RECT  15972.5 26790.0 16042.5 26860.0 ;
      RECT  15900.0 26290.0 15970.0 26825.0 ;
      RECT  15935.0 26790.0 16007.5 26860.0 ;
      RECT  15972.5 26825.0 16042.5 27357.5 ;
      RECT  16235.0 27202.5 16305.0 27272.5 ;
      RECT  16162.5 27202.5 16232.5 27272.5 ;
      RECT  16235.0 27237.5 16305.0 27840.0 ;
      RECT  16197.5 27202.5 16270.0 27272.5 ;
      RECT  16162.5 26632.5 16232.5 27237.5 ;
      RECT  15900.0 27772.5 15970.0 27907.5 ;
      RECT  16235.0 26222.5 16305.0 26357.5 ;
      RECT  15972.5 27357.5 16042.5 27492.5 ;
      RECT  16162.5 26497.5 16232.5 26632.5 ;
      RECT  16420.0 26397.5 16490.0 26532.5 ;
      RECT  15900.0 27840.0 15970.0 27980.0 ;
      RECT  16235.0 27840.0 16305.0 27980.0 ;
      RECT  15900.0 26150.0 15970.0 26290.0 ;
      RECT  16235.0 26150.0 16305.0 26290.0 ;
      RECT  15715.0 26150.0 15785.0 27980.0 ;
      RECT  16420.0 26150.0 16490.0 27980.0 ;
      RECT  16605.0 26790.0 16675.0 26860.0 ;
      RECT  16677.5 26790.0 16747.5 26860.0 ;
      RECT  16605.0 26290.0 16675.0 26825.0 ;
      RECT  16640.0 26790.0 16712.5 26860.0 ;
      RECT  16677.5 26825.0 16747.5 27357.5 ;
      RECT  16940.0 27202.5 17010.0 27272.5 ;
      RECT  16867.5 27202.5 16937.5 27272.5 ;
      RECT  16940.0 27237.5 17010.0 27840.0 ;
      RECT  16902.5 27202.5 16975.0 27272.5 ;
      RECT  16867.5 26632.5 16937.5 27237.5 ;
      RECT  16605.0 27772.5 16675.0 27907.5 ;
      RECT  16940.0 26222.5 17010.0 26357.5 ;
      RECT  16677.5 27357.5 16747.5 27492.5 ;
      RECT  16867.5 26497.5 16937.5 26632.5 ;
      RECT  17125.0 26397.5 17195.0 26532.5 ;
      RECT  16605.0 27840.0 16675.0 27980.0 ;
      RECT  16940.0 27840.0 17010.0 27980.0 ;
      RECT  16605.0 26150.0 16675.0 26290.0 ;
      RECT  16940.0 26150.0 17010.0 26290.0 ;
      RECT  16420.0 26150.0 16490.0 27980.0 ;
      RECT  17125.0 26150.0 17195.0 27980.0 ;
      RECT  17310.0 26790.0 17380.0 26860.0 ;
      RECT  17382.5 26790.0 17452.5 26860.0 ;
      RECT  17310.0 26290.0 17380.0 26825.0 ;
      RECT  17345.0 26790.0 17417.5 26860.0 ;
      RECT  17382.5 26825.0 17452.5 27357.5 ;
      RECT  17645.0 27202.5 17715.0 27272.5 ;
      RECT  17572.5 27202.5 17642.5 27272.5 ;
      RECT  17645.0 27237.5 17715.0 27840.0 ;
      RECT  17607.5 27202.5 17680.0 27272.5 ;
      RECT  17572.5 26632.5 17642.5 27237.5 ;
      RECT  17310.0 27772.5 17380.0 27907.5 ;
      RECT  17645.0 26222.5 17715.0 26357.5 ;
      RECT  17382.5 27357.5 17452.5 27492.5 ;
      RECT  17572.5 26497.5 17642.5 26632.5 ;
      RECT  17830.0 26397.5 17900.0 26532.5 ;
      RECT  17310.0 27840.0 17380.0 27980.0 ;
      RECT  17645.0 27840.0 17715.0 27980.0 ;
      RECT  17310.0 26150.0 17380.0 26290.0 ;
      RECT  17645.0 26150.0 17715.0 26290.0 ;
      RECT  17125.0 26150.0 17195.0 27980.0 ;
      RECT  17830.0 26150.0 17900.0 27980.0 ;
      RECT  18015.0 26790.0 18085.0 26860.0 ;
      RECT  18087.5 26790.0 18157.5 26860.0 ;
      RECT  18015.0 26290.0 18085.0 26825.0 ;
      RECT  18050.0 26790.0 18122.5 26860.0 ;
      RECT  18087.5 26825.0 18157.5 27357.5 ;
      RECT  18350.0 27202.5 18420.0 27272.5 ;
      RECT  18277.5 27202.5 18347.5 27272.5 ;
      RECT  18350.0 27237.5 18420.0 27840.0 ;
      RECT  18312.5 27202.5 18385.0 27272.5 ;
      RECT  18277.5 26632.5 18347.5 27237.5 ;
      RECT  18015.0 27772.5 18085.0 27907.5 ;
      RECT  18350.0 26222.5 18420.0 26357.5 ;
      RECT  18087.5 27357.5 18157.5 27492.5 ;
      RECT  18277.5 26497.5 18347.5 26632.5 ;
      RECT  18535.0 26397.5 18605.0 26532.5 ;
      RECT  18015.0 27840.0 18085.0 27980.0 ;
      RECT  18350.0 27840.0 18420.0 27980.0 ;
      RECT  18015.0 26150.0 18085.0 26290.0 ;
      RECT  18350.0 26150.0 18420.0 26290.0 ;
      RECT  17830.0 26150.0 17900.0 27980.0 ;
      RECT  18535.0 26150.0 18605.0 27980.0 ;
      RECT  18720.0 26790.0 18790.0 26860.0 ;
      RECT  18792.5 26790.0 18862.5 26860.0 ;
      RECT  18720.0 26290.0 18790.0 26825.0 ;
      RECT  18755.0 26790.0 18827.5 26860.0 ;
      RECT  18792.5 26825.0 18862.5 27357.5 ;
      RECT  19055.0 27202.5 19125.0 27272.5 ;
      RECT  18982.5 27202.5 19052.5 27272.5 ;
      RECT  19055.0 27237.5 19125.0 27840.0 ;
      RECT  19017.5 27202.5 19090.0 27272.5 ;
      RECT  18982.5 26632.5 19052.5 27237.5 ;
      RECT  18720.0 27772.5 18790.0 27907.5 ;
      RECT  19055.0 26222.5 19125.0 26357.5 ;
      RECT  18792.5 27357.5 18862.5 27492.5 ;
      RECT  18982.5 26497.5 19052.5 26632.5 ;
      RECT  19240.0 26397.5 19310.0 26532.5 ;
      RECT  18720.0 27840.0 18790.0 27980.0 ;
      RECT  19055.0 27840.0 19125.0 27980.0 ;
      RECT  18720.0 26150.0 18790.0 26290.0 ;
      RECT  19055.0 26150.0 19125.0 26290.0 ;
      RECT  18535.0 26150.0 18605.0 27980.0 ;
      RECT  19240.0 26150.0 19310.0 27980.0 ;
      RECT  19425.0 26790.0 19495.0 26860.0 ;
      RECT  19497.5 26790.0 19567.5 26860.0 ;
      RECT  19425.0 26290.0 19495.0 26825.0 ;
      RECT  19460.0 26790.0 19532.5 26860.0 ;
      RECT  19497.5 26825.0 19567.5 27357.5 ;
      RECT  19760.0 27202.5 19830.0 27272.5 ;
      RECT  19687.5 27202.5 19757.5 27272.5 ;
      RECT  19760.0 27237.5 19830.0 27840.0 ;
      RECT  19722.5 27202.5 19795.0 27272.5 ;
      RECT  19687.5 26632.5 19757.5 27237.5 ;
      RECT  19425.0 27772.5 19495.0 27907.5 ;
      RECT  19760.0 26222.5 19830.0 26357.5 ;
      RECT  19497.5 27357.5 19567.5 27492.5 ;
      RECT  19687.5 26497.5 19757.5 26632.5 ;
      RECT  19945.0 26397.5 20015.0 26532.5 ;
      RECT  19425.0 27840.0 19495.0 27980.0 ;
      RECT  19760.0 27840.0 19830.0 27980.0 ;
      RECT  19425.0 26150.0 19495.0 26290.0 ;
      RECT  19760.0 26150.0 19830.0 26290.0 ;
      RECT  19240.0 26150.0 19310.0 27980.0 ;
      RECT  19945.0 26150.0 20015.0 27980.0 ;
      RECT  20130.0 26790.0 20200.0 26860.0 ;
      RECT  20202.5 26790.0 20272.5 26860.0 ;
      RECT  20130.0 26290.0 20200.0 26825.0 ;
      RECT  20165.0 26790.0 20237.5 26860.0 ;
      RECT  20202.5 26825.0 20272.5 27357.5 ;
      RECT  20465.0 27202.5 20535.0 27272.5 ;
      RECT  20392.5 27202.5 20462.5 27272.5 ;
      RECT  20465.0 27237.5 20535.0 27840.0 ;
      RECT  20427.5 27202.5 20500.0 27272.5 ;
      RECT  20392.5 26632.5 20462.5 27237.5 ;
      RECT  20130.0 27772.5 20200.0 27907.5 ;
      RECT  20465.0 26222.5 20535.0 26357.5 ;
      RECT  20202.5 27357.5 20272.5 27492.5 ;
      RECT  20392.5 26497.5 20462.5 26632.5 ;
      RECT  20650.0 26397.5 20720.0 26532.5 ;
      RECT  20130.0 27840.0 20200.0 27980.0 ;
      RECT  20465.0 27840.0 20535.0 27980.0 ;
      RECT  20130.0 26150.0 20200.0 26290.0 ;
      RECT  20465.0 26150.0 20535.0 26290.0 ;
      RECT  19945.0 26150.0 20015.0 27980.0 ;
      RECT  20650.0 26150.0 20720.0 27980.0 ;
      RECT  20835.0 26790.0 20905.0 26860.0 ;
      RECT  20907.5 26790.0 20977.5 26860.0 ;
      RECT  20835.0 26290.0 20905.0 26825.0 ;
      RECT  20870.0 26790.0 20942.5 26860.0 ;
      RECT  20907.5 26825.0 20977.5 27357.5 ;
      RECT  21170.0 27202.5 21240.0 27272.5 ;
      RECT  21097.5 27202.5 21167.5 27272.5 ;
      RECT  21170.0 27237.5 21240.0 27840.0 ;
      RECT  21132.5 27202.5 21205.0 27272.5 ;
      RECT  21097.5 26632.5 21167.5 27237.5 ;
      RECT  20835.0 27772.5 20905.0 27907.5 ;
      RECT  21170.0 26222.5 21240.0 26357.5 ;
      RECT  20907.5 27357.5 20977.5 27492.5 ;
      RECT  21097.5 26497.5 21167.5 26632.5 ;
      RECT  21355.0 26397.5 21425.0 26532.5 ;
      RECT  20835.0 27840.0 20905.0 27980.0 ;
      RECT  21170.0 27840.0 21240.0 27980.0 ;
      RECT  20835.0 26150.0 20905.0 26290.0 ;
      RECT  21170.0 26150.0 21240.0 26290.0 ;
      RECT  20650.0 26150.0 20720.0 27980.0 ;
      RECT  21355.0 26150.0 21425.0 27980.0 ;
      RECT  21540.0 26790.0 21610.0 26860.0 ;
      RECT  21612.5 26790.0 21682.5 26860.0 ;
      RECT  21540.0 26290.0 21610.0 26825.0 ;
      RECT  21575.0 26790.0 21647.5 26860.0 ;
      RECT  21612.5 26825.0 21682.5 27357.5 ;
      RECT  21875.0 27202.5 21945.0 27272.5 ;
      RECT  21802.5 27202.5 21872.5 27272.5 ;
      RECT  21875.0 27237.5 21945.0 27840.0 ;
      RECT  21837.5 27202.5 21910.0 27272.5 ;
      RECT  21802.5 26632.5 21872.5 27237.5 ;
      RECT  21540.0 27772.5 21610.0 27907.5 ;
      RECT  21875.0 26222.5 21945.0 26357.5 ;
      RECT  21612.5 27357.5 21682.5 27492.5 ;
      RECT  21802.5 26497.5 21872.5 26632.5 ;
      RECT  22060.0 26397.5 22130.0 26532.5 ;
      RECT  21540.0 27840.0 21610.0 27980.0 ;
      RECT  21875.0 27840.0 21945.0 27980.0 ;
      RECT  21540.0 26150.0 21610.0 26290.0 ;
      RECT  21875.0 26150.0 21945.0 26290.0 ;
      RECT  21355.0 26150.0 21425.0 27980.0 ;
      RECT  22060.0 26150.0 22130.0 27980.0 ;
      RECT  22245.0 26790.0 22315.0 26860.0 ;
      RECT  22317.5 26790.0 22387.5 26860.0 ;
      RECT  22245.0 26290.0 22315.0 26825.0 ;
      RECT  22280.0 26790.0 22352.5 26860.0 ;
      RECT  22317.5 26825.0 22387.5 27357.5 ;
      RECT  22580.0 27202.5 22650.0 27272.5 ;
      RECT  22507.5 27202.5 22577.5 27272.5 ;
      RECT  22580.0 27237.5 22650.0 27840.0 ;
      RECT  22542.5 27202.5 22615.0 27272.5 ;
      RECT  22507.5 26632.5 22577.5 27237.5 ;
      RECT  22245.0 27772.5 22315.0 27907.5 ;
      RECT  22580.0 26222.5 22650.0 26357.5 ;
      RECT  22317.5 27357.5 22387.5 27492.5 ;
      RECT  22507.5 26497.5 22577.5 26632.5 ;
      RECT  22765.0 26397.5 22835.0 26532.5 ;
      RECT  22245.0 27840.0 22315.0 27980.0 ;
      RECT  22580.0 27840.0 22650.0 27980.0 ;
      RECT  22245.0 26150.0 22315.0 26290.0 ;
      RECT  22580.0 26150.0 22650.0 26290.0 ;
      RECT  22060.0 26150.0 22130.0 27980.0 ;
      RECT  22765.0 26150.0 22835.0 27980.0 ;
      RECT  22950.0 26790.0 23020.0 26860.0 ;
      RECT  23022.5 26790.0 23092.5 26860.0 ;
      RECT  22950.0 26290.0 23020.0 26825.0 ;
      RECT  22985.0 26790.0 23057.5 26860.0 ;
      RECT  23022.5 26825.0 23092.5 27357.5 ;
      RECT  23285.0 27202.5 23355.0 27272.5 ;
      RECT  23212.5 27202.5 23282.5 27272.5 ;
      RECT  23285.0 27237.5 23355.0 27840.0 ;
      RECT  23247.5 27202.5 23320.0 27272.5 ;
      RECT  23212.5 26632.5 23282.5 27237.5 ;
      RECT  22950.0 27772.5 23020.0 27907.5 ;
      RECT  23285.0 26222.5 23355.0 26357.5 ;
      RECT  23022.5 27357.5 23092.5 27492.5 ;
      RECT  23212.5 26497.5 23282.5 26632.5 ;
      RECT  23470.0 26397.5 23540.0 26532.5 ;
      RECT  22950.0 27840.0 23020.0 27980.0 ;
      RECT  23285.0 27840.0 23355.0 27980.0 ;
      RECT  22950.0 26150.0 23020.0 26290.0 ;
      RECT  23285.0 26150.0 23355.0 26290.0 ;
      RECT  22765.0 26150.0 22835.0 27980.0 ;
      RECT  23470.0 26150.0 23540.0 27980.0 ;
      RECT  23655.0 26790.0 23725.0 26860.0 ;
      RECT  23727.5 26790.0 23797.5 26860.0 ;
      RECT  23655.0 26290.0 23725.0 26825.0 ;
      RECT  23690.0 26790.0 23762.5 26860.0 ;
      RECT  23727.5 26825.0 23797.5 27357.5 ;
      RECT  23990.0 27202.5 24060.0 27272.5 ;
      RECT  23917.5 27202.5 23987.5 27272.5 ;
      RECT  23990.0 27237.5 24060.0 27840.0 ;
      RECT  23952.5 27202.5 24025.0 27272.5 ;
      RECT  23917.5 26632.5 23987.5 27237.5 ;
      RECT  23655.0 27772.5 23725.0 27907.5 ;
      RECT  23990.0 26222.5 24060.0 26357.5 ;
      RECT  23727.5 27357.5 23797.5 27492.5 ;
      RECT  23917.5 26497.5 23987.5 26632.5 ;
      RECT  24175.0 26397.5 24245.0 26532.5 ;
      RECT  23655.0 27840.0 23725.0 27980.0 ;
      RECT  23990.0 27840.0 24060.0 27980.0 ;
      RECT  23655.0 26150.0 23725.0 26290.0 ;
      RECT  23990.0 26150.0 24060.0 26290.0 ;
      RECT  23470.0 26150.0 23540.0 27980.0 ;
      RECT  24175.0 26150.0 24245.0 27980.0 ;
      RECT  24360.0 26790.0 24430.0 26860.0 ;
      RECT  24432.5 26790.0 24502.5 26860.0 ;
      RECT  24360.0 26290.0 24430.0 26825.0 ;
      RECT  24395.0 26790.0 24467.5 26860.0 ;
      RECT  24432.5 26825.0 24502.5 27357.5 ;
      RECT  24695.0 27202.5 24765.0 27272.5 ;
      RECT  24622.5 27202.5 24692.5 27272.5 ;
      RECT  24695.0 27237.5 24765.0 27840.0 ;
      RECT  24657.5 27202.5 24730.0 27272.5 ;
      RECT  24622.5 26632.5 24692.5 27237.5 ;
      RECT  24360.0 27772.5 24430.0 27907.5 ;
      RECT  24695.0 26222.5 24765.0 26357.5 ;
      RECT  24432.5 27357.5 24502.5 27492.5 ;
      RECT  24622.5 26497.5 24692.5 26632.5 ;
      RECT  24880.0 26397.5 24950.0 26532.5 ;
      RECT  24360.0 27840.0 24430.0 27980.0 ;
      RECT  24695.0 27840.0 24765.0 27980.0 ;
      RECT  24360.0 26150.0 24430.0 26290.0 ;
      RECT  24695.0 26150.0 24765.0 26290.0 ;
      RECT  24175.0 26150.0 24245.0 27980.0 ;
      RECT  24880.0 26150.0 24950.0 27980.0 ;
      RECT  25065.0 26790.0 25135.0 26860.0 ;
      RECT  25137.5 26790.0 25207.5 26860.0 ;
      RECT  25065.0 26290.0 25135.0 26825.0 ;
      RECT  25100.0 26790.0 25172.5 26860.0 ;
      RECT  25137.5 26825.0 25207.5 27357.5 ;
      RECT  25400.0 27202.5 25470.0 27272.5 ;
      RECT  25327.5 27202.5 25397.5 27272.5 ;
      RECT  25400.0 27237.5 25470.0 27840.0 ;
      RECT  25362.5 27202.5 25435.0 27272.5 ;
      RECT  25327.5 26632.5 25397.5 27237.5 ;
      RECT  25065.0 27772.5 25135.0 27907.5 ;
      RECT  25400.0 26222.5 25470.0 26357.5 ;
      RECT  25137.5 27357.5 25207.5 27492.5 ;
      RECT  25327.5 26497.5 25397.5 26632.5 ;
      RECT  25585.0 26397.5 25655.0 26532.5 ;
      RECT  25065.0 27840.0 25135.0 27980.0 ;
      RECT  25400.0 27840.0 25470.0 27980.0 ;
      RECT  25065.0 26150.0 25135.0 26290.0 ;
      RECT  25400.0 26150.0 25470.0 26290.0 ;
      RECT  24880.0 26150.0 24950.0 27980.0 ;
      RECT  25585.0 26150.0 25655.0 27980.0 ;
      RECT  25770.0 26790.0 25840.0 26860.0 ;
      RECT  25842.5 26790.0 25912.5 26860.0 ;
      RECT  25770.0 26290.0 25840.0 26825.0 ;
      RECT  25805.0 26790.0 25877.5 26860.0 ;
      RECT  25842.5 26825.0 25912.5 27357.5 ;
      RECT  26105.0 27202.5 26175.0 27272.5 ;
      RECT  26032.5 27202.5 26102.5 27272.5 ;
      RECT  26105.0 27237.5 26175.0 27840.0 ;
      RECT  26067.5 27202.5 26140.0 27272.5 ;
      RECT  26032.5 26632.5 26102.5 27237.5 ;
      RECT  25770.0 27772.5 25840.0 27907.5 ;
      RECT  26105.0 26222.5 26175.0 26357.5 ;
      RECT  25842.5 27357.5 25912.5 27492.5 ;
      RECT  26032.5 26497.5 26102.5 26632.5 ;
      RECT  26290.0 26397.5 26360.0 26532.5 ;
      RECT  25770.0 27840.0 25840.0 27980.0 ;
      RECT  26105.0 27840.0 26175.0 27980.0 ;
      RECT  25770.0 26150.0 25840.0 26290.0 ;
      RECT  26105.0 26150.0 26175.0 26290.0 ;
      RECT  25585.0 26150.0 25655.0 27980.0 ;
      RECT  26290.0 26150.0 26360.0 27980.0 ;
      RECT  26475.0 26790.0 26545.0 26860.0 ;
      RECT  26547.5 26790.0 26617.5 26860.0 ;
      RECT  26475.0 26290.0 26545.0 26825.0 ;
      RECT  26510.0 26790.0 26582.5 26860.0 ;
      RECT  26547.5 26825.0 26617.5 27357.5 ;
      RECT  26810.0 27202.5 26880.0 27272.5 ;
      RECT  26737.5 27202.5 26807.5 27272.5 ;
      RECT  26810.0 27237.5 26880.0 27840.0 ;
      RECT  26772.5 27202.5 26845.0 27272.5 ;
      RECT  26737.5 26632.5 26807.5 27237.5 ;
      RECT  26475.0 27772.5 26545.0 27907.5 ;
      RECT  26810.0 26222.5 26880.0 26357.5 ;
      RECT  26547.5 27357.5 26617.5 27492.5 ;
      RECT  26737.5 26497.5 26807.5 26632.5 ;
      RECT  26995.0 26397.5 27065.0 26532.5 ;
      RECT  26475.0 27840.0 26545.0 27980.0 ;
      RECT  26810.0 27840.0 26880.0 27980.0 ;
      RECT  26475.0 26150.0 26545.0 26290.0 ;
      RECT  26810.0 26150.0 26880.0 26290.0 ;
      RECT  26290.0 26150.0 26360.0 27980.0 ;
      RECT  26995.0 26150.0 27065.0 27980.0 ;
      RECT  27180.0 26790.0 27250.0 26860.0 ;
      RECT  27252.5 26790.0 27322.5 26860.0 ;
      RECT  27180.0 26290.0 27250.0 26825.0 ;
      RECT  27215.0 26790.0 27287.5 26860.0 ;
      RECT  27252.5 26825.0 27322.5 27357.5 ;
      RECT  27515.0 27202.5 27585.0 27272.5 ;
      RECT  27442.5 27202.5 27512.5 27272.5 ;
      RECT  27515.0 27237.5 27585.0 27840.0 ;
      RECT  27477.5 27202.5 27550.0 27272.5 ;
      RECT  27442.5 26632.5 27512.5 27237.5 ;
      RECT  27180.0 27772.5 27250.0 27907.5 ;
      RECT  27515.0 26222.5 27585.0 26357.5 ;
      RECT  27252.5 27357.5 27322.5 27492.5 ;
      RECT  27442.5 26497.5 27512.5 26632.5 ;
      RECT  27700.0 26397.5 27770.0 26532.5 ;
      RECT  27180.0 27840.0 27250.0 27980.0 ;
      RECT  27515.0 27840.0 27585.0 27980.0 ;
      RECT  27180.0 26150.0 27250.0 26290.0 ;
      RECT  27515.0 26150.0 27585.0 26290.0 ;
      RECT  26995.0 26150.0 27065.0 27980.0 ;
      RECT  27700.0 26150.0 27770.0 27980.0 ;
      RECT  27885.0 26790.0 27955.0 26860.0 ;
      RECT  27957.5 26790.0 28027.5 26860.0 ;
      RECT  27885.0 26290.0 27955.0 26825.0 ;
      RECT  27920.0 26790.0 27992.5 26860.0 ;
      RECT  27957.5 26825.0 28027.5 27357.5 ;
      RECT  28220.0 27202.5 28290.0 27272.5 ;
      RECT  28147.5 27202.5 28217.5 27272.5 ;
      RECT  28220.0 27237.5 28290.0 27840.0 ;
      RECT  28182.5 27202.5 28255.0 27272.5 ;
      RECT  28147.5 26632.5 28217.5 27237.5 ;
      RECT  27885.0 27772.5 27955.0 27907.5 ;
      RECT  28220.0 26222.5 28290.0 26357.5 ;
      RECT  27957.5 27357.5 28027.5 27492.5 ;
      RECT  28147.5 26497.5 28217.5 26632.5 ;
      RECT  28405.0 26397.5 28475.0 26532.5 ;
      RECT  27885.0 27840.0 27955.0 27980.0 ;
      RECT  28220.0 27840.0 28290.0 27980.0 ;
      RECT  27885.0 26150.0 27955.0 26290.0 ;
      RECT  28220.0 26150.0 28290.0 26290.0 ;
      RECT  27700.0 26150.0 27770.0 27980.0 ;
      RECT  28405.0 26150.0 28475.0 27980.0 ;
      RECT  28590.0 26790.0 28660.0 26860.0 ;
      RECT  28662.5 26790.0 28732.5 26860.0 ;
      RECT  28590.0 26290.0 28660.0 26825.0 ;
      RECT  28625.0 26790.0 28697.5 26860.0 ;
      RECT  28662.5 26825.0 28732.5 27357.5 ;
      RECT  28925.0 27202.5 28995.0 27272.5 ;
      RECT  28852.5 27202.5 28922.5 27272.5 ;
      RECT  28925.0 27237.5 28995.0 27840.0 ;
      RECT  28887.5 27202.5 28960.0 27272.5 ;
      RECT  28852.5 26632.5 28922.5 27237.5 ;
      RECT  28590.0 27772.5 28660.0 27907.5 ;
      RECT  28925.0 26222.5 28995.0 26357.5 ;
      RECT  28662.5 27357.5 28732.5 27492.5 ;
      RECT  28852.5 26497.5 28922.5 26632.5 ;
      RECT  29110.0 26397.5 29180.0 26532.5 ;
      RECT  28590.0 27840.0 28660.0 27980.0 ;
      RECT  28925.0 27840.0 28995.0 27980.0 ;
      RECT  28590.0 26150.0 28660.0 26290.0 ;
      RECT  28925.0 26150.0 28995.0 26290.0 ;
      RECT  28405.0 26150.0 28475.0 27980.0 ;
      RECT  29110.0 26150.0 29180.0 27980.0 ;
      RECT  29295.0 26790.0 29365.0 26860.0 ;
      RECT  29367.5 26790.0 29437.5 26860.0 ;
      RECT  29295.0 26290.0 29365.0 26825.0 ;
      RECT  29330.0 26790.0 29402.5 26860.0 ;
      RECT  29367.5 26825.0 29437.5 27357.5 ;
      RECT  29630.0 27202.5 29700.0 27272.5 ;
      RECT  29557.5 27202.5 29627.5 27272.5 ;
      RECT  29630.0 27237.5 29700.0 27840.0 ;
      RECT  29592.5 27202.5 29665.0 27272.5 ;
      RECT  29557.5 26632.5 29627.5 27237.5 ;
      RECT  29295.0 27772.5 29365.0 27907.5 ;
      RECT  29630.0 26222.5 29700.0 26357.5 ;
      RECT  29367.5 27357.5 29437.5 27492.5 ;
      RECT  29557.5 26497.5 29627.5 26632.5 ;
      RECT  29815.0 26397.5 29885.0 26532.5 ;
      RECT  29295.0 27840.0 29365.0 27980.0 ;
      RECT  29630.0 27840.0 29700.0 27980.0 ;
      RECT  29295.0 26150.0 29365.0 26290.0 ;
      RECT  29630.0 26150.0 29700.0 26290.0 ;
      RECT  29110.0 26150.0 29180.0 27980.0 ;
      RECT  29815.0 26150.0 29885.0 27980.0 ;
      RECT  30000.0 26790.0 30070.0 26860.0 ;
      RECT  30072.5 26790.0 30142.5 26860.0 ;
      RECT  30000.0 26290.0 30070.0 26825.0 ;
      RECT  30035.0 26790.0 30107.5 26860.0 ;
      RECT  30072.5 26825.0 30142.5 27357.5 ;
      RECT  30335.0 27202.5 30405.0 27272.5 ;
      RECT  30262.5 27202.5 30332.5 27272.5 ;
      RECT  30335.0 27237.5 30405.0 27840.0 ;
      RECT  30297.5 27202.5 30370.0 27272.5 ;
      RECT  30262.5 26632.5 30332.5 27237.5 ;
      RECT  30000.0 27772.5 30070.0 27907.5 ;
      RECT  30335.0 26222.5 30405.0 26357.5 ;
      RECT  30072.5 27357.5 30142.5 27492.5 ;
      RECT  30262.5 26497.5 30332.5 26632.5 ;
      RECT  30520.0 26397.5 30590.0 26532.5 ;
      RECT  30000.0 27840.0 30070.0 27980.0 ;
      RECT  30335.0 27840.0 30405.0 27980.0 ;
      RECT  30000.0 26150.0 30070.0 26290.0 ;
      RECT  30335.0 26150.0 30405.0 26290.0 ;
      RECT  29815.0 26150.0 29885.0 27980.0 ;
      RECT  30520.0 26150.0 30590.0 27980.0 ;
      RECT  30705.0 26790.0 30775.0 26860.0 ;
      RECT  30777.5 26790.0 30847.5 26860.0 ;
      RECT  30705.0 26290.0 30775.0 26825.0 ;
      RECT  30740.0 26790.0 30812.5 26860.0 ;
      RECT  30777.5 26825.0 30847.5 27357.5 ;
      RECT  31040.0 27202.5 31110.0 27272.5 ;
      RECT  30967.5 27202.5 31037.5 27272.5 ;
      RECT  31040.0 27237.5 31110.0 27840.0 ;
      RECT  31002.5 27202.5 31075.0 27272.5 ;
      RECT  30967.5 26632.5 31037.5 27237.5 ;
      RECT  30705.0 27772.5 30775.0 27907.5 ;
      RECT  31040.0 26222.5 31110.0 26357.5 ;
      RECT  30777.5 27357.5 30847.5 27492.5 ;
      RECT  30967.5 26497.5 31037.5 26632.5 ;
      RECT  31225.0 26397.5 31295.0 26532.5 ;
      RECT  30705.0 27840.0 30775.0 27980.0 ;
      RECT  31040.0 27840.0 31110.0 27980.0 ;
      RECT  30705.0 26150.0 30775.0 26290.0 ;
      RECT  31040.0 26150.0 31110.0 26290.0 ;
      RECT  30520.0 26150.0 30590.0 27980.0 ;
      RECT  31225.0 26150.0 31295.0 27980.0 ;
      RECT  31410.0 26790.0 31480.0 26860.0 ;
      RECT  31482.5 26790.0 31552.5 26860.0 ;
      RECT  31410.0 26290.0 31480.0 26825.0 ;
      RECT  31445.0 26790.0 31517.5 26860.0 ;
      RECT  31482.5 26825.0 31552.5 27357.5 ;
      RECT  31745.0 27202.5 31815.0 27272.5 ;
      RECT  31672.5 27202.5 31742.5 27272.5 ;
      RECT  31745.0 27237.5 31815.0 27840.0 ;
      RECT  31707.5 27202.5 31780.0 27272.5 ;
      RECT  31672.5 26632.5 31742.5 27237.5 ;
      RECT  31410.0 27772.5 31480.0 27907.5 ;
      RECT  31745.0 26222.5 31815.0 26357.5 ;
      RECT  31482.5 27357.5 31552.5 27492.5 ;
      RECT  31672.5 26497.5 31742.5 26632.5 ;
      RECT  31930.0 26397.5 32000.0 26532.5 ;
      RECT  31410.0 27840.0 31480.0 27980.0 ;
      RECT  31745.0 27840.0 31815.0 27980.0 ;
      RECT  31410.0 26150.0 31480.0 26290.0 ;
      RECT  31745.0 26150.0 31815.0 26290.0 ;
      RECT  31225.0 26150.0 31295.0 27980.0 ;
      RECT  31930.0 26150.0 32000.0 27980.0 ;
      RECT  32115.0 26790.0 32185.0 26860.0 ;
      RECT  32187.5 26790.0 32257.5 26860.0 ;
      RECT  32115.0 26290.0 32185.0 26825.0 ;
      RECT  32150.0 26790.0 32222.5 26860.0 ;
      RECT  32187.5 26825.0 32257.5 27357.5 ;
      RECT  32450.0 27202.5 32520.0 27272.5 ;
      RECT  32377.5 27202.5 32447.5 27272.5 ;
      RECT  32450.0 27237.5 32520.0 27840.0 ;
      RECT  32412.5 27202.5 32485.0 27272.5 ;
      RECT  32377.5 26632.5 32447.5 27237.5 ;
      RECT  32115.0 27772.5 32185.0 27907.5 ;
      RECT  32450.0 26222.5 32520.0 26357.5 ;
      RECT  32187.5 27357.5 32257.5 27492.5 ;
      RECT  32377.5 26497.5 32447.5 26632.5 ;
      RECT  32635.0 26397.5 32705.0 26532.5 ;
      RECT  32115.0 27840.0 32185.0 27980.0 ;
      RECT  32450.0 27840.0 32520.0 27980.0 ;
      RECT  32115.0 26150.0 32185.0 26290.0 ;
      RECT  32450.0 26150.0 32520.0 26290.0 ;
      RECT  31930.0 26150.0 32000.0 27980.0 ;
      RECT  32635.0 26150.0 32705.0 27980.0 ;
      RECT  32820.0 26790.0 32890.0 26860.0 ;
      RECT  32892.5 26790.0 32962.5 26860.0 ;
      RECT  32820.0 26290.0 32890.0 26825.0 ;
      RECT  32855.0 26790.0 32927.5 26860.0 ;
      RECT  32892.5 26825.0 32962.5 27357.5 ;
      RECT  33155.0 27202.5 33225.0 27272.5 ;
      RECT  33082.5 27202.5 33152.5 27272.5 ;
      RECT  33155.0 27237.5 33225.0 27840.0 ;
      RECT  33117.5 27202.5 33190.0 27272.5 ;
      RECT  33082.5 26632.5 33152.5 27237.5 ;
      RECT  32820.0 27772.5 32890.0 27907.5 ;
      RECT  33155.0 26222.5 33225.0 26357.5 ;
      RECT  32892.5 27357.5 32962.5 27492.5 ;
      RECT  33082.5 26497.5 33152.5 26632.5 ;
      RECT  33340.0 26397.5 33410.0 26532.5 ;
      RECT  32820.0 27840.0 32890.0 27980.0 ;
      RECT  33155.0 27840.0 33225.0 27980.0 ;
      RECT  32820.0 26150.0 32890.0 26290.0 ;
      RECT  33155.0 26150.0 33225.0 26290.0 ;
      RECT  32635.0 26150.0 32705.0 27980.0 ;
      RECT  33340.0 26150.0 33410.0 27980.0 ;
      RECT  33525.0 26790.0 33595.0 26860.0 ;
      RECT  33597.5 26790.0 33667.5 26860.0 ;
      RECT  33525.0 26290.0 33595.0 26825.0 ;
      RECT  33560.0 26790.0 33632.5 26860.0 ;
      RECT  33597.5 26825.0 33667.5 27357.5 ;
      RECT  33860.0 27202.5 33930.0 27272.5 ;
      RECT  33787.5 27202.5 33857.5 27272.5 ;
      RECT  33860.0 27237.5 33930.0 27840.0 ;
      RECT  33822.5 27202.5 33895.0 27272.5 ;
      RECT  33787.5 26632.5 33857.5 27237.5 ;
      RECT  33525.0 27772.5 33595.0 27907.5 ;
      RECT  33860.0 26222.5 33930.0 26357.5 ;
      RECT  33597.5 27357.5 33667.5 27492.5 ;
      RECT  33787.5 26497.5 33857.5 26632.5 ;
      RECT  34045.0 26397.5 34115.0 26532.5 ;
      RECT  33525.0 27840.0 33595.0 27980.0 ;
      RECT  33860.0 27840.0 33930.0 27980.0 ;
      RECT  33525.0 26150.0 33595.0 26290.0 ;
      RECT  33860.0 26150.0 33930.0 26290.0 ;
      RECT  33340.0 26150.0 33410.0 27980.0 ;
      RECT  34045.0 26150.0 34115.0 27980.0 ;
      RECT  34230.0 26790.0 34300.0 26860.0 ;
      RECT  34302.5 26790.0 34372.5 26860.0 ;
      RECT  34230.0 26290.0 34300.0 26825.0 ;
      RECT  34265.0 26790.0 34337.5 26860.0 ;
      RECT  34302.5 26825.0 34372.5 27357.5 ;
      RECT  34565.0 27202.5 34635.0 27272.5 ;
      RECT  34492.5 27202.5 34562.5 27272.5 ;
      RECT  34565.0 27237.5 34635.0 27840.0 ;
      RECT  34527.5 27202.5 34600.0 27272.5 ;
      RECT  34492.5 26632.5 34562.5 27237.5 ;
      RECT  34230.0 27772.5 34300.0 27907.5 ;
      RECT  34565.0 26222.5 34635.0 26357.5 ;
      RECT  34302.5 27357.5 34372.5 27492.5 ;
      RECT  34492.5 26497.5 34562.5 26632.5 ;
      RECT  34750.0 26397.5 34820.0 26532.5 ;
      RECT  34230.0 27840.0 34300.0 27980.0 ;
      RECT  34565.0 27840.0 34635.0 27980.0 ;
      RECT  34230.0 26150.0 34300.0 26290.0 ;
      RECT  34565.0 26150.0 34635.0 26290.0 ;
      RECT  34045.0 26150.0 34115.0 27980.0 ;
      RECT  34750.0 26150.0 34820.0 27980.0 ;
      RECT  34935.0 26790.0 35005.0 26860.0 ;
      RECT  35007.5 26790.0 35077.5 26860.0 ;
      RECT  34935.0 26290.0 35005.0 26825.0 ;
      RECT  34970.0 26790.0 35042.5 26860.0 ;
      RECT  35007.5 26825.0 35077.5 27357.5 ;
      RECT  35270.0 27202.5 35340.0 27272.5 ;
      RECT  35197.5 27202.5 35267.5 27272.5 ;
      RECT  35270.0 27237.5 35340.0 27840.0 ;
      RECT  35232.5 27202.5 35305.0 27272.5 ;
      RECT  35197.5 26632.5 35267.5 27237.5 ;
      RECT  34935.0 27772.5 35005.0 27907.5 ;
      RECT  35270.0 26222.5 35340.0 26357.5 ;
      RECT  35007.5 27357.5 35077.5 27492.5 ;
      RECT  35197.5 26497.5 35267.5 26632.5 ;
      RECT  35455.0 26397.5 35525.0 26532.5 ;
      RECT  34935.0 27840.0 35005.0 27980.0 ;
      RECT  35270.0 27840.0 35340.0 27980.0 ;
      RECT  34935.0 26150.0 35005.0 26290.0 ;
      RECT  35270.0 26150.0 35340.0 26290.0 ;
      RECT  34750.0 26150.0 34820.0 27980.0 ;
      RECT  35455.0 26150.0 35525.0 27980.0 ;
      RECT  35640.0 26790.0 35710.0 26860.0 ;
      RECT  35712.5 26790.0 35782.5 26860.0 ;
      RECT  35640.0 26290.0 35710.0 26825.0 ;
      RECT  35675.0 26790.0 35747.5 26860.0 ;
      RECT  35712.5 26825.0 35782.5 27357.5 ;
      RECT  35975.0 27202.5 36045.0 27272.5 ;
      RECT  35902.5 27202.5 35972.5 27272.5 ;
      RECT  35975.0 27237.5 36045.0 27840.0 ;
      RECT  35937.5 27202.5 36010.0 27272.5 ;
      RECT  35902.5 26632.5 35972.5 27237.5 ;
      RECT  35640.0 27772.5 35710.0 27907.5 ;
      RECT  35975.0 26222.5 36045.0 26357.5 ;
      RECT  35712.5 27357.5 35782.5 27492.5 ;
      RECT  35902.5 26497.5 35972.5 26632.5 ;
      RECT  36160.0 26397.5 36230.0 26532.5 ;
      RECT  35640.0 27840.0 35710.0 27980.0 ;
      RECT  35975.0 27840.0 36045.0 27980.0 ;
      RECT  35640.0 26150.0 35710.0 26290.0 ;
      RECT  35975.0 26150.0 36045.0 26290.0 ;
      RECT  35455.0 26150.0 35525.0 27980.0 ;
      RECT  36160.0 26150.0 36230.0 27980.0 ;
      RECT  36345.0 26790.0 36415.0 26860.0 ;
      RECT  36417.5 26790.0 36487.5 26860.0 ;
      RECT  36345.0 26290.0 36415.0 26825.0 ;
      RECT  36380.0 26790.0 36452.5 26860.0 ;
      RECT  36417.5 26825.0 36487.5 27357.5 ;
      RECT  36680.0 27202.5 36750.0 27272.5 ;
      RECT  36607.5 27202.5 36677.5 27272.5 ;
      RECT  36680.0 27237.5 36750.0 27840.0 ;
      RECT  36642.5 27202.5 36715.0 27272.5 ;
      RECT  36607.5 26632.5 36677.5 27237.5 ;
      RECT  36345.0 27772.5 36415.0 27907.5 ;
      RECT  36680.0 26222.5 36750.0 26357.5 ;
      RECT  36417.5 27357.5 36487.5 27492.5 ;
      RECT  36607.5 26497.5 36677.5 26632.5 ;
      RECT  36865.0 26397.5 36935.0 26532.5 ;
      RECT  36345.0 27840.0 36415.0 27980.0 ;
      RECT  36680.0 27840.0 36750.0 27980.0 ;
      RECT  36345.0 26150.0 36415.0 26290.0 ;
      RECT  36680.0 26150.0 36750.0 26290.0 ;
      RECT  36160.0 26150.0 36230.0 27980.0 ;
      RECT  36865.0 26150.0 36935.0 27980.0 ;
      RECT  37050.0 26790.0 37120.0 26860.0 ;
      RECT  37122.5 26790.0 37192.5 26860.0 ;
      RECT  37050.0 26290.0 37120.0 26825.0 ;
      RECT  37085.0 26790.0 37157.5 26860.0 ;
      RECT  37122.5 26825.0 37192.5 27357.5 ;
      RECT  37385.0 27202.5 37455.0 27272.5 ;
      RECT  37312.5 27202.5 37382.5 27272.5 ;
      RECT  37385.0 27237.5 37455.0 27840.0 ;
      RECT  37347.5 27202.5 37420.0 27272.5 ;
      RECT  37312.5 26632.5 37382.5 27237.5 ;
      RECT  37050.0 27772.5 37120.0 27907.5 ;
      RECT  37385.0 26222.5 37455.0 26357.5 ;
      RECT  37122.5 27357.5 37192.5 27492.5 ;
      RECT  37312.5 26497.5 37382.5 26632.5 ;
      RECT  37570.0 26397.5 37640.0 26532.5 ;
      RECT  37050.0 27840.0 37120.0 27980.0 ;
      RECT  37385.0 27840.0 37455.0 27980.0 ;
      RECT  37050.0 26150.0 37120.0 26290.0 ;
      RECT  37385.0 26150.0 37455.0 26290.0 ;
      RECT  36865.0 26150.0 36935.0 27980.0 ;
      RECT  37570.0 26150.0 37640.0 27980.0 ;
      RECT  37755.0 26790.0 37825.0 26860.0 ;
      RECT  37827.5 26790.0 37897.5 26860.0 ;
      RECT  37755.0 26290.0 37825.0 26825.0 ;
      RECT  37790.0 26790.0 37862.5 26860.0 ;
      RECT  37827.5 26825.0 37897.5 27357.5 ;
      RECT  38090.0 27202.5 38160.0 27272.5 ;
      RECT  38017.5 27202.5 38087.5 27272.5 ;
      RECT  38090.0 27237.5 38160.0 27840.0 ;
      RECT  38052.5 27202.5 38125.0 27272.5 ;
      RECT  38017.5 26632.5 38087.5 27237.5 ;
      RECT  37755.0 27772.5 37825.0 27907.5 ;
      RECT  38090.0 26222.5 38160.0 26357.5 ;
      RECT  37827.5 27357.5 37897.5 27492.5 ;
      RECT  38017.5 26497.5 38087.5 26632.5 ;
      RECT  38275.0 26397.5 38345.0 26532.5 ;
      RECT  37755.0 27840.0 37825.0 27980.0 ;
      RECT  38090.0 27840.0 38160.0 27980.0 ;
      RECT  37755.0 26150.0 37825.0 26290.0 ;
      RECT  38090.0 26150.0 38160.0 26290.0 ;
      RECT  37570.0 26150.0 37640.0 27980.0 ;
      RECT  38275.0 26150.0 38345.0 27980.0 ;
      RECT  38460.0 26790.0 38530.0 26860.0 ;
      RECT  38532.5 26790.0 38602.5 26860.0 ;
      RECT  38460.0 26290.0 38530.0 26825.0 ;
      RECT  38495.0 26790.0 38567.5 26860.0 ;
      RECT  38532.5 26825.0 38602.5 27357.5 ;
      RECT  38795.0 27202.5 38865.0 27272.5 ;
      RECT  38722.5 27202.5 38792.5 27272.5 ;
      RECT  38795.0 27237.5 38865.0 27840.0 ;
      RECT  38757.5 27202.5 38830.0 27272.5 ;
      RECT  38722.5 26632.5 38792.5 27237.5 ;
      RECT  38460.0 27772.5 38530.0 27907.5 ;
      RECT  38795.0 26222.5 38865.0 26357.5 ;
      RECT  38532.5 27357.5 38602.5 27492.5 ;
      RECT  38722.5 26497.5 38792.5 26632.5 ;
      RECT  38980.0 26397.5 39050.0 26532.5 ;
      RECT  38460.0 27840.0 38530.0 27980.0 ;
      RECT  38795.0 27840.0 38865.0 27980.0 ;
      RECT  38460.0 26150.0 38530.0 26290.0 ;
      RECT  38795.0 26150.0 38865.0 26290.0 ;
      RECT  38275.0 26150.0 38345.0 27980.0 ;
      RECT  38980.0 26150.0 39050.0 27980.0 ;
      RECT  39165.0 26790.0 39235.0 26860.0 ;
      RECT  39237.5 26790.0 39307.5 26860.0 ;
      RECT  39165.0 26290.0 39235.0 26825.0 ;
      RECT  39200.0 26790.0 39272.5 26860.0 ;
      RECT  39237.5 26825.0 39307.5 27357.5 ;
      RECT  39500.0 27202.5 39570.0 27272.5 ;
      RECT  39427.5 27202.5 39497.5 27272.5 ;
      RECT  39500.0 27237.5 39570.0 27840.0 ;
      RECT  39462.5 27202.5 39535.0 27272.5 ;
      RECT  39427.5 26632.5 39497.5 27237.5 ;
      RECT  39165.0 27772.5 39235.0 27907.5 ;
      RECT  39500.0 26222.5 39570.0 26357.5 ;
      RECT  39237.5 27357.5 39307.5 27492.5 ;
      RECT  39427.5 26497.5 39497.5 26632.5 ;
      RECT  39685.0 26397.5 39755.0 26532.5 ;
      RECT  39165.0 27840.0 39235.0 27980.0 ;
      RECT  39500.0 27840.0 39570.0 27980.0 ;
      RECT  39165.0 26150.0 39235.0 26290.0 ;
      RECT  39500.0 26150.0 39570.0 26290.0 ;
      RECT  38980.0 26150.0 39050.0 27980.0 ;
      RECT  39685.0 26150.0 39755.0 27980.0 ;
      RECT  39870.0 26790.0 39940.0 26860.0 ;
      RECT  39942.5 26790.0 40012.5 26860.0 ;
      RECT  39870.0 26290.0 39940.0 26825.0 ;
      RECT  39905.0 26790.0 39977.5 26860.0 ;
      RECT  39942.5 26825.0 40012.5 27357.5 ;
      RECT  40205.0 27202.5 40275.0 27272.5 ;
      RECT  40132.5 27202.5 40202.5 27272.5 ;
      RECT  40205.0 27237.5 40275.0 27840.0 ;
      RECT  40167.5 27202.5 40240.0 27272.5 ;
      RECT  40132.5 26632.5 40202.5 27237.5 ;
      RECT  39870.0 27772.5 39940.0 27907.5 ;
      RECT  40205.0 26222.5 40275.0 26357.5 ;
      RECT  39942.5 27357.5 40012.5 27492.5 ;
      RECT  40132.5 26497.5 40202.5 26632.5 ;
      RECT  40390.0 26397.5 40460.0 26532.5 ;
      RECT  39870.0 27840.0 39940.0 27980.0 ;
      RECT  40205.0 27840.0 40275.0 27980.0 ;
      RECT  39870.0 26150.0 39940.0 26290.0 ;
      RECT  40205.0 26150.0 40275.0 26290.0 ;
      RECT  39685.0 26150.0 39755.0 27980.0 ;
      RECT  40390.0 26150.0 40460.0 27980.0 ;
      RECT  40575.0 26790.0 40645.0 26860.0 ;
      RECT  40647.5 26790.0 40717.5 26860.0 ;
      RECT  40575.0 26290.0 40645.0 26825.0 ;
      RECT  40610.0 26790.0 40682.5 26860.0 ;
      RECT  40647.5 26825.0 40717.5 27357.5 ;
      RECT  40910.0 27202.5 40980.0 27272.5 ;
      RECT  40837.5 27202.5 40907.5 27272.5 ;
      RECT  40910.0 27237.5 40980.0 27840.0 ;
      RECT  40872.5 27202.5 40945.0 27272.5 ;
      RECT  40837.5 26632.5 40907.5 27237.5 ;
      RECT  40575.0 27772.5 40645.0 27907.5 ;
      RECT  40910.0 26222.5 40980.0 26357.5 ;
      RECT  40647.5 27357.5 40717.5 27492.5 ;
      RECT  40837.5 26497.5 40907.5 26632.5 ;
      RECT  41095.0 26397.5 41165.0 26532.5 ;
      RECT  40575.0 27840.0 40645.0 27980.0 ;
      RECT  40910.0 27840.0 40980.0 27980.0 ;
      RECT  40575.0 26150.0 40645.0 26290.0 ;
      RECT  40910.0 26150.0 40980.0 26290.0 ;
      RECT  40390.0 26150.0 40460.0 27980.0 ;
      RECT  41095.0 26150.0 41165.0 27980.0 ;
      RECT  41280.0 26790.0 41350.0 26860.0 ;
      RECT  41352.5 26790.0 41422.5 26860.0 ;
      RECT  41280.0 26290.0 41350.0 26825.0 ;
      RECT  41315.0 26790.0 41387.5 26860.0 ;
      RECT  41352.5 26825.0 41422.5 27357.5 ;
      RECT  41615.0 27202.5 41685.0 27272.5 ;
      RECT  41542.5 27202.5 41612.5 27272.5 ;
      RECT  41615.0 27237.5 41685.0 27840.0 ;
      RECT  41577.5 27202.5 41650.0 27272.5 ;
      RECT  41542.5 26632.5 41612.5 27237.5 ;
      RECT  41280.0 27772.5 41350.0 27907.5 ;
      RECT  41615.0 26222.5 41685.0 26357.5 ;
      RECT  41352.5 27357.5 41422.5 27492.5 ;
      RECT  41542.5 26497.5 41612.5 26632.5 ;
      RECT  41800.0 26397.5 41870.0 26532.5 ;
      RECT  41280.0 27840.0 41350.0 27980.0 ;
      RECT  41615.0 27840.0 41685.0 27980.0 ;
      RECT  41280.0 26150.0 41350.0 26290.0 ;
      RECT  41615.0 26150.0 41685.0 26290.0 ;
      RECT  41095.0 26150.0 41165.0 27980.0 ;
      RECT  41800.0 26150.0 41870.0 27980.0 ;
      RECT  41985.0 26790.0 42055.0 26860.0 ;
      RECT  42057.5 26790.0 42127.5 26860.0 ;
      RECT  41985.0 26290.0 42055.0 26825.0 ;
      RECT  42020.0 26790.0 42092.5 26860.0 ;
      RECT  42057.5 26825.0 42127.5 27357.5 ;
      RECT  42320.0 27202.5 42390.0 27272.5 ;
      RECT  42247.5 27202.5 42317.5 27272.5 ;
      RECT  42320.0 27237.5 42390.0 27840.0 ;
      RECT  42282.5 27202.5 42355.0 27272.5 ;
      RECT  42247.5 26632.5 42317.5 27237.5 ;
      RECT  41985.0 27772.5 42055.0 27907.5 ;
      RECT  42320.0 26222.5 42390.0 26357.5 ;
      RECT  42057.5 27357.5 42127.5 27492.5 ;
      RECT  42247.5 26497.5 42317.5 26632.5 ;
      RECT  42505.0 26397.5 42575.0 26532.5 ;
      RECT  41985.0 27840.0 42055.0 27980.0 ;
      RECT  42320.0 27840.0 42390.0 27980.0 ;
      RECT  41985.0 26150.0 42055.0 26290.0 ;
      RECT  42320.0 26150.0 42390.0 26290.0 ;
      RECT  41800.0 26150.0 41870.0 27980.0 ;
      RECT  42505.0 26150.0 42575.0 27980.0 ;
      RECT  42690.0 26790.0 42760.0 26860.0 ;
      RECT  42762.5 26790.0 42832.5 26860.0 ;
      RECT  42690.0 26290.0 42760.0 26825.0 ;
      RECT  42725.0 26790.0 42797.5 26860.0 ;
      RECT  42762.5 26825.0 42832.5 27357.5 ;
      RECT  43025.0 27202.5 43095.0 27272.5 ;
      RECT  42952.5 27202.5 43022.5 27272.5 ;
      RECT  43025.0 27237.5 43095.0 27840.0 ;
      RECT  42987.5 27202.5 43060.0 27272.5 ;
      RECT  42952.5 26632.5 43022.5 27237.5 ;
      RECT  42690.0 27772.5 42760.0 27907.5 ;
      RECT  43025.0 26222.5 43095.0 26357.5 ;
      RECT  42762.5 27357.5 42832.5 27492.5 ;
      RECT  42952.5 26497.5 43022.5 26632.5 ;
      RECT  43210.0 26397.5 43280.0 26532.5 ;
      RECT  42690.0 27840.0 42760.0 27980.0 ;
      RECT  43025.0 27840.0 43095.0 27980.0 ;
      RECT  42690.0 26150.0 42760.0 26290.0 ;
      RECT  43025.0 26150.0 43095.0 26290.0 ;
      RECT  42505.0 26150.0 42575.0 27980.0 ;
      RECT  43210.0 26150.0 43280.0 27980.0 ;
      RECT  43395.0 26790.0 43465.0 26860.0 ;
      RECT  43467.5 26790.0 43537.5 26860.0 ;
      RECT  43395.0 26290.0 43465.0 26825.0 ;
      RECT  43430.0 26790.0 43502.5 26860.0 ;
      RECT  43467.5 26825.0 43537.5 27357.5 ;
      RECT  43730.0 27202.5 43800.0 27272.5 ;
      RECT  43657.5 27202.5 43727.5 27272.5 ;
      RECT  43730.0 27237.5 43800.0 27840.0 ;
      RECT  43692.5 27202.5 43765.0 27272.5 ;
      RECT  43657.5 26632.5 43727.5 27237.5 ;
      RECT  43395.0 27772.5 43465.0 27907.5 ;
      RECT  43730.0 26222.5 43800.0 26357.5 ;
      RECT  43467.5 27357.5 43537.5 27492.5 ;
      RECT  43657.5 26497.5 43727.5 26632.5 ;
      RECT  43915.0 26397.5 43985.0 26532.5 ;
      RECT  43395.0 27840.0 43465.0 27980.0 ;
      RECT  43730.0 27840.0 43800.0 27980.0 ;
      RECT  43395.0 26150.0 43465.0 26290.0 ;
      RECT  43730.0 26150.0 43800.0 26290.0 ;
      RECT  43210.0 26150.0 43280.0 27980.0 ;
      RECT  43915.0 26150.0 43985.0 27980.0 ;
      RECT  44100.0 26790.0 44170.0 26860.0 ;
      RECT  44172.5 26790.0 44242.5 26860.0 ;
      RECT  44100.0 26290.0 44170.0 26825.0 ;
      RECT  44135.0 26790.0 44207.5 26860.0 ;
      RECT  44172.5 26825.0 44242.5 27357.5 ;
      RECT  44435.0 27202.5 44505.0 27272.5 ;
      RECT  44362.5 27202.5 44432.5 27272.5 ;
      RECT  44435.0 27237.5 44505.0 27840.0 ;
      RECT  44397.5 27202.5 44470.0 27272.5 ;
      RECT  44362.5 26632.5 44432.5 27237.5 ;
      RECT  44100.0 27772.5 44170.0 27907.5 ;
      RECT  44435.0 26222.5 44505.0 26357.5 ;
      RECT  44172.5 27357.5 44242.5 27492.5 ;
      RECT  44362.5 26497.5 44432.5 26632.5 ;
      RECT  44620.0 26397.5 44690.0 26532.5 ;
      RECT  44100.0 27840.0 44170.0 27980.0 ;
      RECT  44435.0 27840.0 44505.0 27980.0 ;
      RECT  44100.0 26150.0 44170.0 26290.0 ;
      RECT  44435.0 26150.0 44505.0 26290.0 ;
      RECT  43915.0 26150.0 43985.0 27980.0 ;
      RECT  44620.0 26150.0 44690.0 27980.0 ;
      RECT  44805.0 26790.0 44875.0 26860.0 ;
      RECT  44877.5 26790.0 44947.5 26860.0 ;
      RECT  44805.0 26290.0 44875.0 26825.0 ;
      RECT  44840.0 26790.0 44912.5 26860.0 ;
      RECT  44877.5 26825.0 44947.5 27357.5 ;
      RECT  45140.0 27202.5 45210.0 27272.5 ;
      RECT  45067.5 27202.5 45137.5 27272.5 ;
      RECT  45140.0 27237.5 45210.0 27840.0 ;
      RECT  45102.5 27202.5 45175.0 27272.5 ;
      RECT  45067.5 26632.5 45137.5 27237.5 ;
      RECT  44805.0 27772.5 44875.0 27907.5 ;
      RECT  45140.0 26222.5 45210.0 26357.5 ;
      RECT  44877.5 27357.5 44947.5 27492.5 ;
      RECT  45067.5 26497.5 45137.5 26632.5 ;
      RECT  45325.0 26397.5 45395.0 26532.5 ;
      RECT  44805.0 27840.0 44875.0 27980.0 ;
      RECT  45140.0 27840.0 45210.0 27980.0 ;
      RECT  44805.0 26150.0 44875.0 26290.0 ;
      RECT  45140.0 26150.0 45210.0 26290.0 ;
      RECT  44620.0 26150.0 44690.0 27980.0 ;
      RECT  45325.0 26150.0 45395.0 27980.0 ;
      RECT  45510.0 26790.0 45580.0 26860.0 ;
      RECT  45582.5 26790.0 45652.5 26860.0 ;
      RECT  45510.0 26290.0 45580.0 26825.0 ;
      RECT  45545.0 26790.0 45617.5 26860.0 ;
      RECT  45582.5 26825.0 45652.5 27357.5 ;
      RECT  45845.0 27202.5 45915.0 27272.5 ;
      RECT  45772.5 27202.5 45842.5 27272.5 ;
      RECT  45845.0 27237.5 45915.0 27840.0 ;
      RECT  45807.5 27202.5 45880.0 27272.5 ;
      RECT  45772.5 26632.5 45842.5 27237.5 ;
      RECT  45510.0 27772.5 45580.0 27907.5 ;
      RECT  45845.0 26222.5 45915.0 26357.5 ;
      RECT  45582.5 27357.5 45652.5 27492.5 ;
      RECT  45772.5 26497.5 45842.5 26632.5 ;
      RECT  46030.0 26397.5 46100.0 26532.5 ;
      RECT  45510.0 27840.0 45580.0 27980.0 ;
      RECT  45845.0 27840.0 45915.0 27980.0 ;
      RECT  45510.0 26150.0 45580.0 26290.0 ;
      RECT  45845.0 26150.0 45915.0 26290.0 ;
      RECT  45325.0 26150.0 45395.0 27980.0 ;
      RECT  46030.0 26150.0 46100.0 27980.0 ;
      RECT  46215.0 26790.0 46285.0 26860.0 ;
      RECT  46287.5 26790.0 46357.5 26860.0 ;
      RECT  46215.0 26290.0 46285.0 26825.0 ;
      RECT  46250.0 26790.0 46322.5 26860.0 ;
      RECT  46287.5 26825.0 46357.5 27357.5 ;
      RECT  46550.0 27202.5 46620.0 27272.5 ;
      RECT  46477.5 27202.5 46547.5 27272.5 ;
      RECT  46550.0 27237.5 46620.0 27840.0 ;
      RECT  46512.5 27202.5 46585.0 27272.5 ;
      RECT  46477.5 26632.5 46547.5 27237.5 ;
      RECT  46215.0 27772.5 46285.0 27907.5 ;
      RECT  46550.0 26222.5 46620.0 26357.5 ;
      RECT  46287.5 27357.5 46357.5 27492.5 ;
      RECT  46477.5 26497.5 46547.5 26632.5 ;
      RECT  46735.0 26397.5 46805.0 26532.5 ;
      RECT  46215.0 27840.0 46285.0 27980.0 ;
      RECT  46550.0 27840.0 46620.0 27980.0 ;
      RECT  46215.0 26150.0 46285.0 26290.0 ;
      RECT  46550.0 26150.0 46620.0 26290.0 ;
      RECT  46030.0 26150.0 46100.0 27980.0 ;
      RECT  46735.0 26150.0 46805.0 27980.0 ;
      RECT  46920.0 26790.0 46990.0 26860.0 ;
      RECT  46992.5 26790.0 47062.5 26860.0 ;
      RECT  46920.0 26290.0 46990.0 26825.0 ;
      RECT  46955.0 26790.0 47027.5 26860.0 ;
      RECT  46992.5 26825.0 47062.5 27357.5 ;
      RECT  47255.0 27202.5 47325.0 27272.5 ;
      RECT  47182.5 27202.5 47252.5 27272.5 ;
      RECT  47255.0 27237.5 47325.0 27840.0 ;
      RECT  47217.5 27202.5 47290.0 27272.5 ;
      RECT  47182.5 26632.5 47252.5 27237.5 ;
      RECT  46920.0 27772.5 46990.0 27907.5 ;
      RECT  47255.0 26222.5 47325.0 26357.5 ;
      RECT  46992.5 27357.5 47062.5 27492.5 ;
      RECT  47182.5 26497.5 47252.5 26632.5 ;
      RECT  47440.0 26397.5 47510.0 26532.5 ;
      RECT  46920.0 27840.0 46990.0 27980.0 ;
      RECT  47255.0 27840.0 47325.0 27980.0 ;
      RECT  46920.0 26150.0 46990.0 26290.0 ;
      RECT  47255.0 26150.0 47325.0 26290.0 ;
      RECT  46735.0 26150.0 46805.0 27980.0 ;
      RECT  47440.0 26150.0 47510.0 27980.0 ;
      RECT  47625.0 26790.0 47695.0 26860.0 ;
      RECT  47697.5 26790.0 47767.5 26860.0 ;
      RECT  47625.0 26290.0 47695.0 26825.0 ;
      RECT  47660.0 26790.0 47732.5 26860.0 ;
      RECT  47697.5 26825.0 47767.5 27357.5 ;
      RECT  47960.0 27202.5 48030.0 27272.5 ;
      RECT  47887.5 27202.5 47957.5 27272.5 ;
      RECT  47960.0 27237.5 48030.0 27840.0 ;
      RECT  47922.5 27202.5 47995.0 27272.5 ;
      RECT  47887.5 26632.5 47957.5 27237.5 ;
      RECT  47625.0 27772.5 47695.0 27907.5 ;
      RECT  47960.0 26222.5 48030.0 26357.5 ;
      RECT  47697.5 27357.5 47767.5 27492.5 ;
      RECT  47887.5 26497.5 47957.5 26632.5 ;
      RECT  48145.0 26397.5 48215.0 26532.5 ;
      RECT  47625.0 27840.0 47695.0 27980.0 ;
      RECT  47960.0 27840.0 48030.0 27980.0 ;
      RECT  47625.0 26150.0 47695.0 26290.0 ;
      RECT  47960.0 26150.0 48030.0 26290.0 ;
      RECT  47440.0 26150.0 47510.0 27980.0 ;
      RECT  48145.0 26150.0 48215.0 27980.0 ;
      RECT  48330.0 26790.0 48400.0 26860.0 ;
      RECT  48402.5 26790.0 48472.5 26860.0 ;
      RECT  48330.0 26290.0 48400.0 26825.0 ;
      RECT  48365.0 26790.0 48437.5 26860.0 ;
      RECT  48402.5 26825.0 48472.5 27357.5 ;
      RECT  48665.0 27202.5 48735.0 27272.5 ;
      RECT  48592.5 27202.5 48662.5 27272.5 ;
      RECT  48665.0 27237.5 48735.0 27840.0 ;
      RECT  48627.5 27202.5 48700.0 27272.5 ;
      RECT  48592.5 26632.5 48662.5 27237.5 ;
      RECT  48330.0 27772.5 48400.0 27907.5 ;
      RECT  48665.0 26222.5 48735.0 26357.5 ;
      RECT  48402.5 27357.5 48472.5 27492.5 ;
      RECT  48592.5 26497.5 48662.5 26632.5 ;
      RECT  48850.0 26397.5 48920.0 26532.5 ;
      RECT  48330.0 27840.0 48400.0 27980.0 ;
      RECT  48665.0 27840.0 48735.0 27980.0 ;
      RECT  48330.0 26150.0 48400.0 26290.0 ;
      RECT  48665.0 26150.0 48735.0 26290.0 ;
      RECT  48145.0 26150.0 48215.0 27980.0 ;
      RECT  48850.0 26150.0 48920.0 27980.0 ;
      RECT  49035.0 26790.0 49105.0 26860.0 ;
      RECT  49107.5 26790.0 49177.5 26860.0 ;
      RECT  49035.0 26290.0 49105.0 26825.0 ;
      RECT  49070.0 26790.0 49142.5 26860.0 ;
      RECT  49107.5 26825.0 49177.5 27357.5 ;
      RECT  49370.0 27202.5 49440.0 27272.5 ;
      RECT  49297.5 27202.5 49367.5 27272.5 ;
      RECT  49370.0 27237.5 49440.0 27840.0 ;
      RECT  49332.5 27202.5 49405.0 27272.5 ;
      RECT  49297.5 26632.5 49367.5 27237.5 ;
      RECT  49035.0 27772.5 49105.0 27907.5 ;
      RECT  49370.0 26222.5 49440.0 26357.5 ;
      RECT  49107.5 27357.5 49177.5 27492.5 ;
      RECT  49297.5 26497.5 49367.5 26632.5 ;
      RECT  49555.0 26397.5 49625.0 26532.5 ;
      RECT  49035.0 27840.0 49105.0 27980.0 ;
      RECT  49370.0 27840.0 49440.0 27980.0 ;
      RECT  49035.0 26150.0 49105.0 26290.0 ;
      RECT  49370.0 26150.0 49440.0 26290.0 ;
      RECT  48850.0 26150.0 48920.0 27980.0 ;
      RECT  49555.0 26150.0 49625.0 27980.0 ;
      RECT  49740.0 26790.0 49810.0 26860.0 ;
      RECT  49812.5 26790.0 49882.5 26860.0 ;
      RECT  49740.0 26290.0 49810.0 26825.0 ;
      RECT  49775.0 26790.0 49847.5 26860.0 ;
      RECT  49812.5 26825.0 49882.5 27357.5 ;
      RECT  50075.0 27202.5 50145.0 27272.5 ;
      RECT  50002.5 27202.5 50072.5 27272.5 ;
      RECT  50075.0 27237.5 50145.0 27840.0 ;
      RECT  50037.5 27202.5 50110.0 27272.5 ;
      RECT  50002.5 26632.5 50072.5 27237.5 ;
      RECT  49740.0 27772.5 49810.0 27907.5 ;
      RECT  50075.0 26222.5 50145.0 26357.5 ;
      RECT  49812.5 27357.5 49882.5 27492.5 ;
      RECT  50002.5 26497.5 50072.5 26632.5 ;
      RECT  50260.0 26397.5 50330.0 26532.5 ;
      RECT  49740.0 27840.0 49810.0 27980.0 ;
      RECT  50075.0 27840.0 50145.0 27980.0 ;
      RECT  49740.0 26150.0 49810.0 26290.0 ;
      RECT  50075.0 26150.0 50145.0 26290.0 ;
      RECT  49555.0 26150.0 49625.0 27980.0 ;
      RECT  50260.0 26150.0 50330.0 27980.0 ;
      RECT  50445.0 26790.0 50515.0 26860.0 ;
      RECT  50517.5 26790.0 50587.5 26860.0 ;
      RECT  50445.0 26290.0 50515.0 26825.0 ;
      RECT  50480.0 26790.0 50552.5 26860.0 ;
      RECT  50517.5 26825.0 50587.5 27357.5 ;
      RECT  50780.0 27202.5 50850.0 27272.5 ;
      RECT  50707.5 27202.5 50777.5 27272.5 ;
      RECT  50780.0 27237.5 50850.0 27840.0 ;
      RECT  50742.5 27202.5 50815.0 27272.5 ;
      RECT  50707.5 26632.5 50777.5 27237.5 ;
      RECT  50445.0 27772.5 50515.0 27907.5 ;
      RECT  50780.0 26222.5 50850.0 26357.5 ;
      RECT  50517.5 27357.5 50587.5 27492.5 ;
      RECT  50707.5 26497.5 50777.5 26632.5 ;
      RECT  50965.0 26397.5 51035.0 26532.5 ;
      RECT  50445.0 27840.0 50515.0 27980.0 ;
      RECT  50780.0 27840.0 50850.0 27980.0 ;
      RECT  50445.0 26150.0 50515.0 26290.0 ;
      RECT  50780.0 26150.0 50850.0 26290.0 ;
      RECT  50260.0 26150.0 50330.0 27980.0 ;
      RECT  50965.0 26150.0 51035.0 27980.0 ;
      RECT  51150.0 26790.0 51220.0 26860.0 ;
      RECT  51222.5 26790.0 51292.5 26860.0 ;
      RECT  51150.0 26290.0 51220.0 26825.0 ;
      RECT  51185.0 26790.0 51257.5 26860.0 ;
      RECT  51222.5 26825.0 51292.5 27357.5 ;
      RECT  51485.0 27202.5 51555.0 27272.5 ;
      RECT  51412.5 27202.5 51482.5 27272.5 ;
      RECT  51485.0 27237.5 51555.0 27840.0 ;
      RECT  51447.5 27202.5 51520.0 27272.5 ;
      RECT  51412.5 26632.5 51482.5 27237.5 ;
      RECT  51150.0 27772.5 51220.0 27907.5 ;
      RECT  51485.0 26222.5 51555.0 26357.5 ;
      RECT  51222.5 27357.5 51292.5 27492.5 ;
      RECT  51412.5 26497.5 51482.5 26632.5 ;
      RECT  51670.0 26397.5 51740.0 26532.5 ;
      RECT  51150.0 27840.0 51220.0 27980.0 ;
      RECT  51485.0 27840.0 51555.0 27980.0 ;
      RECT  51150.0 26150.0 51220.0 26290.0 ;
      RECT  51485.0 26150.0 51555.0 26290.0 ;
      RECT  50965.0 26150.0 51035.0 27980.0 ;
      RECT  51670.0 26150.0 51740.0 27980.0 ;
      RECT  51855.0 26790.0 51925.0 26860.0 ;
      RECT  51927.5 26790.0 51997.5 26860.0 ;
      RECT  51855.0 26290.0 51925.0 26825.0 ;
      RECT  51890.0 26790.0 51962.5 26860.0 ;
      RECT  51927.5 26825.0 51997.5 27357.5 ;
      RECT  52190.0 27202.5 52260.0 27272.5 ;
      RECT  52117.5 27202.5 52187.5 27272.5 ;
      RECT  52190.0 27237.5 52260.0 27840.0 ;
      RECT  52152.5 27202.5 52225.0 27272.5 ;
      RECT  52117.5 26632.5 52187.5 27237.5 ;
      RECT  51855.0 27772.5 51925.0 27907.5 ;
      RECT  52190.0 26222.5 52260.0 26357.5 ;
      RECT  51927.5 27357.5 51997.5 27492.5 ;
      RECT  52117.5 26497.5 52187.5 26632.5 ;
      RECT  52375.0 26397.5 52445.0 26532.5 ;
      RECT  51855.0 27840.0 51925.0 27980.0 ;
      RECT  52190.0 27840.0 52260.0 27980.0 ;
      RECT  51855.0 26150.0 51925.0 26290.0 ;
      RECT  52190.0 26150.0 52260.0 26290.0 ;
      RECT  51670.0 26150.0 51740.0 27980.0 ;
      RECT  52375.0 26150.0 52445.0 27980.0 ;
      RECT  52560.0 26790.0 52630.0 26860.0 ;
      RECT  52632.5 26790.0 52702.5 26860.0 ;
      RECT  52560.0 26290.0 52630.0 26825.0 ;
      RECT  52595.0 26790.0 52667.5 26860.0 ;
      RECT  52632.5 26825.0 52702.5 27357.5 ;
      RECT  52895.0 27202.5 52965.0 27272.5 ;
      RECT  52822.5 27202.5 52892.5 27272.5 ;
      RECT  52895.0 27237.5 52965.0 27840.0 ;
      RECT  52857.5 27202.5 52930.0 27272.5 ;
      RECT  52822.5 26632.5 52892.5 27237.5 ;
      RECT  52560.0 27772.5 52630.0 27907.5 ;
      RECT  52895.0 26222.5 52965.0 26357.5 ;
      RECT  52632.5 27357.5 52702.5 27492.5 ;
      RECT  52822.5 26497.5 52892.5 26632.5 ;
      RECT  53080.0 26397.5 53150.0 26532.5 ;
      RECT  52560.0 27840.0 52630.0 27980.0 ;
      RECT  52895.0 27840.0 52965.0 27980.0 ;
      RECT  52560.0 26150.0 52630.0 26290.0 ;
      RECT  52895.0 26150.0 52965.0 26290.0 ;
      RECT  52375.0 26150.0 52445.0 27980.0 ;
      RECT  53080.0 26150.0 53150.0 27980.0 ;
      RECT  53265.0 26790.0 53335.0 26860.0 ;
      RECT  53337.5 26790.0 53407.5 26860.0 ;
      RECT  53265.0 26290.0 53335.0 26825.0 ;
      RECT  53300.0 26790.0 53372.5 26860.0 ;
      RECT  53337.5 26825.0 53407.5 27357.5 ;
      RECT  53600.0 27202.5 53670.0 27272.5 ;
      RECT  53527.5 27202.5 53597.5 27272.5 ;
      RECT  53600.0 27237.5 53670.0 27840.0 ;
      RECT  53562.5 27202.5 53635.0 27272.5 ;
      RECT  53527.5 26632.5 53597.5 27237.5 ;
      RECT  53265.0 27772.5 53335.0 27907.5 ;
      RECT  53600.0 26222.5 53670.0 26357.5 ;
      RECT  53337.5 27357.5 53407.5 27492.5 ;
      RECT  53527.5 26497.5 53597.5 26632.5 ;
      RECT  53785.0 26397.5 53855.0 26532.5 ;
      RECT  53265.0 27840.0 53335.0 27980.0 ;
      RECT  53600.0 27840.0 53670.0 27980.0 ;
      RECT  53265.0 26150.0 53335.0 26290.0 ;
      RECT  53600.0 26150.0 53670.0 26290.0 ;
      RECT  53080.0 26150.0 53150.0 27980.0 ;
      RECT  53785.0 26150.0 53855.0 27980.0 ;
      RECT  53970.0 26790.0 54040.0 26860.0 ;
      RECT  54042.5 26790.0 54112.5 26860.0 ;
      RECT  53970.0 26290.0 54040.0 26825.0 ;
      RECT  54005.0 26790.0 54077.5 26860.0 ;
      RECT  54042.5 26825.0 54112.5 27357.5 ;
      RECT  54305.0 27202.5 54375.0 27272.5 ;
      RECT  54232.5 27202.5 54302.5 27272.5 ;
      RECT  54305.0 27237.5 54375.0 27840.0 ;
      RECT  54267.5 27202.5 54340.0 27272.5 ;
      RECT  54232.5 26632.5 54302.5 27237.5 ;
      RECT  53970.0 27772.5 54040.0 27907.5 ;
      RECT  54305.0 26222.5 54375.0 26357.5 ;
      RECT  54042.5 27357.5 54112.5 27492.5 ;
      RECT  54232.5 26497.5 54302.5 26632.5 ;
      RECT  54490.0 26397.5 54560.0 26532.5 ;
      RECT  53970.0 27840.0 54040.0 27980.0 ;
      RECT  54305.0 27840.0 54375.0 27980.0 ;
      RECT  53970.0 26150.0 54040.0 26290.0 ;
      RECT  54305.0 26150.0 54375.0 26290.0 ;
      RECT  53785.0 26150.0 53855.0 27980.0 ;
      RECT  54490.0 26150.0 54560.0 27980.0 ;
      RECT  54675.0 26790.0 54745.0 26860.0 ;
      RECT  54747.5 26790.0 54817.5 26860.0 ;
      RECT  54675.0 26290.0 54745.0 26825.0 ;
      RECT  54710.0 26790.0 54782.5 26860.0 ;
      RECT  54747.5 26825.0 54817.5 27357.5 ;
      RECT  55010.0 27202.5 55080.0 27272.5 ;
      RECT  54937.5 27202.5 55007.5 27272.5 ;
      RECT  55010.0 27237.5 55080.0 27840.0 ;
      RECT  54972.5 27202.5 55045.0 27272.5 ;
      RECT  54937.5 26632.5 55007.5 27237.5 ;
      RECT  54675.0 27772.5 54745.0 27907.5 ;
      RECT  55010.0 26222.5 55080.0 26357.5 ;
      RECT  54747.5 27357.5 54817.5 27492.5 ;
      RECT  54937.5 26497.5 55007.5 26632.5 ;
      RECT  55195.0 26397.5 55265.0 26532.5 ;
      RECT  54675.0 27840.0 54745.0 27980.0 ;
      RECT  55010.0 27840.0 55080.0 27980.0 ;
      RECT  54675.0 26150.0 54745.0 26290.0 ;
      RECT  55010.0 26150.0 55080.0 26290.0 ;
      RECT  54490.0 26150.0 54560.0 27980.0 ;
      RECT  55195.0 26150.0 55265.0 27980.0 ;
      RECT  55380.0 26790.0 55450.0 26860.0 ;
      RECT  55452.5 26790.0 55522.5 26860.0 ;
      RECT  55380.0 26290.0 55450.0 26825.0 ;
      RECT  55415.0 26790.0 55487.5 26860.0 ;
      RECT  55452.5 26825.0 55522.5 27357.5 ;
      RECT  55715.0 27202.5 55785.0 27272.5 ;
      RECT  55642.5 27202.5 55712.5 27272.5 ;
      RECT  55715.0 27237.5 55785.0 27840.0 ;
      RECT  55677.5 27202.5 55750.0 27272.5 ;
      RECT  55642.5 26632.5 55712.5 27237.5 ;
      RECT  55380.0 27772.5 55450.0 27907.5 ;
      RECT  55715.0 26222.5 55785.0 26357.5 ;
      RECT  55452.5 27357.5 55522.5 27492.5 ;
      RECT  55642.5 26497.5 55712.5 26632.5 ;
      RECT  55900.0 26397.5 55970.0 26532.5 ;
      RECT  55380.0 27840.0 55450.0 27980.0 ;
      RECT  55715.0 27840.0 55785.0 27980.0 ;
      RECT  55380.0 26150.0 55450.0 26290.0 ;
      RECT  55715.0 26150.0 55785.0 26290.0 ;
      RECT  55195.0 26150.0 55265.0 27980.0 ;
      RECT  55900.0 26150.0 55970.0 27980.0 ;
      RECT  56085.0 26790.0 56155.0 26860.0 ;
      RECT  56157.5 26790.0 56227.5 26860.0 ;
      RECT  56085.0 26290.0 56155.0 26825.0 ;
      RECT  56120.0 26790.0 56192.5 26860.0 ;
      RECT  56157.5 26825.0 56227.5 27357.5 ;
      RECT  56420.0 27202.5 56490.0 27272.5 ;
      RECT  56347.5 27202.5 56417.5 27272.5 ;
      RECT  56420.0 27237.5 56490.0 27840.0 ;
      RECT  56382.5 27202.5 56455.0 27272.5 ;
      RECT  56347.5 26632.5 56417.5 27237.5 ;
      RECT  56085.0 27772.5 56155.0 27907.5 ;
      RECT  56420.0 26222.5 56490.0 26357.5 ;
      RECT  56157.5 27357.5 56227.5 27492.5 ;
      RECT  56347.5 26497.5 56417.5 26632.5 ;
      RECT  56605.0 26397.5 56675.0 26532.5 ;
      RECT  56085.0 27840.0 56155.0 27980.0 ;
      RECT  56420.0 27840.0 56490.0 27980.0 ;
      RECT  56085.0 26150.0 56155.0 26290.0 ;
      RECT  56420.0 26150.0 56490.0 26290.0 ;
      RECT  55900.0 26150.0 55970.0 27980.0 ;
      RECT  56605.0 26150.0 56675.0 27980.0 ;
      RECT  56790.0 26790.0 56860.0 26860.0 ;
      RECT  56862.5 26790.0 56932.5 26860.0 ;
      RECT  56790.0 26290.0 56860.0 26825.0 ;
      RECT  56825.0 26790.0 56897.5 26860.0 ;
      RECT  56862.5 26825.0 56932.5 27357.5 ;
      RECT  57125.0 27202.5 57195.0 27272.5 ;
      RECT  57052.5 27202.5 57122.5 27272.5 ;
      RECT  57125.0 27237.5 57195.0 27840.0 ;
      RECT  57087.5 27202.5 57160.0 27272.5 ;
      RECT  57052.5 26632.5 57122.5 27237.5 ;
      RECT  56790.0 27772.5 56860.0 27907.5 ;
      RECT  57125.0 26222.5 57195.0 26357.5 ;
      RECT  56862.5 27357.5 56932.5 27492.5 ;
      RECT  57052.5 26497.5 57122.5 26632.5 ;
      RECT  57310.0 26397.5 57380.0 26532.5 ;
      RECT  56790.0 27840.0 56860.0 27980.0 ;
      RECT  57125.0 27840.0 57195.0 27980.0 ;
      RECT  56790.0 26150.0 56860.0 26290.0 ;
      RECT  57125.0 26150.0 57195.0 26290.0 ;
      RECT  56605.0 26150.0 56675.0 27980.0 ;
      RECT  57310.0 26150.0 57380.0 27980.0 ;
      RECT  57495.0 26790.0 57565.0 26860.0 ;
      RECT  57567.5 26790.0 57637.5 26860.0 ;
      RECT  57495.0 26290.0 57565.0 26825.0 ;
      RECT  57530.0 26790.0 57602.5 26860.0 ;
      RECT  57567.5 26825.0 57637.5 27357.5 ;
      RECT  57830.0 27202.5 57900.0 27272.5 ;
      RECT  57757.5 27202.5 57827.5 27272.5 ;
      RECT  57830.0 27237.5 57900.0 27840.0 ;
      RECT  57792.5 27202.5 57865.0 27272.5 ;
      RECT  57757.5 26632.5 57827.5 27237.5 ;
      RECT  57495.0 27772.5 57565.0 27907.5 ;
      RECT  57830.0 26222.5 57900.0 26357.5 ;
      RECT  57567.5 27357.5 57637.5 27492.5 ;
      RECT  57757.5 26497.5 57827.5 26632.5 ;
      RECT  58015.0 26397.5 58085.0 26532.5 ;
      RECT  57495.0 27840.0 57565.0 27980.0 ;
      RECT  57830.0 27840.0 57900.0 27980.0 ;
      RECT  57495.0 26150.0 57565.0 26290.0 ;
      RECT  57830.0 26150.0 57900.0 26290.0 ;
      RECT  57310.0 26150.0 57380.0 27980.0 ;
      RECT  58015.0 26150.0 58085.0 27980.0 ;
      RECT  58200.0 26790.0 58270.0 26860.0 ;
      RECT  58272.5 26790.0 58342.5 26860.0 ;
      RECT  58200.0 26290.0 58270.0 26825.0 ;
      RECT  58235.0 26790.0 58307.5 26860.0 ;
      RECT  58272.5 26825.0 58342.5 27357.5 ;
      RECT  58535.0 27202.5 58605.0 27272.5 ;
      RECT  58462.5 27202.5 58532.5 27272.5 ;
      RECT  58535.0 27237.5 58605.0 27840.0 ;
      RECT  58497.5 27202.5 58570.0 27272.5 ;
      RECT  58462.5 26632.5 58532.5 27237.5 ;
      RECT  58200.0 27772.5 58270.0 27907.5 ;
      RECT  58535.0 26222.5 58605.0 26357.5 ;
      RECT  58272.5 27357.5 58342.5 27492.5 ;
      RECT  58462.5 26497.5 58532.5 26632.5 ;
      RECT  58720.0 26397.5 58790.0 26532.5 ;
      RECT  58200.0 27840.0 58270.0 27980.0 ;
      RECT  58535.0 27840.0 58605.0 27980.0 ;
      RECT  58200.0 26150.0 58270.0 26290.0 ;
      RECT  58535.0 26150.0 58605.0 26290.0 ;
      RECT  58015.0 26150.0 58085.0 27980.0 ;
      RECT  58720.0 26150.0 58790.0 27980.0 ;
      RECT  58905.0 26790.0 58975.0 26860.0 ;
      RECT  58977.5 26790.0 59047.5 26860.0 ;
      RECT  58905.0 26290.0 58975.0 26825.0 ;
      RECT  58940.0 26790.0 59012.5 26860.0 ;
      RECT  58977.5 26825.0 59047.5 27357.5 ;
      RECT  59240.0 27202.5 59310.0 27272.5 ;
      RECT  59167.5 27202.5 59237.5 27272.5 ;
      RECT  59240.0 27237.5 59310.0 27840.0 ;
      RECT  59202.5 27202.5 59275.0 27272.5 ;
      RECT  59167.5 26632.5 59237.5 27237.5 ;
      RECT  58905.0 27772.5 58975.0 27907.5 ;
      RECT  59240.0 26222.5 59310.0 26357.5 ;
      RECT  58977.5 27357.5 59047.5 27492.5 ;
      RECT  59167.5 26497.5 59237.5 26632.5 ;
      RECT  59425.0 26397.5 59495.0 26532.5 ;
      RECT  58905.0 27840.0 58975.0 27980.0 ;
      RECT  59240.0 27840.0 59310.0 27980.0 ;
      RECT  58905.0 26150.0 58975.0 26290.0 ;
      RECT  59240.0 26150.0 59310.0 26290.0 ;
      RECT  58720.0 26150.0 58790.0 27980.0 ;
      RECT  59425.0 26150.0 59495.0 27980.0 ;
      RECT  59610.0 26790.0 59680.0 26860.0 ;
      RECT  59682.5 26790.0 59752.5 26860.0 ;
      RECT  59610.0 26290.0 59680.0 26825.0 ;
      RECT  59645.0 26790.0 59717.5 26860.0 ;
      RECT  59682.5 26825.0 59752.5 27357.5 ;
      RECT  59945.0 27202.5 60015.0 27272.5 ;
      RECT  59872.5 27202.5 59942.5 27272.5 ;
      RECT  59945.0 27237.5 60015.0 27840.0 ;
      RECT  59907.5 27202.5 59980.0 27272.5 ;
      RECT  59872.5 26632.5 59942.5 27237.5 ;
      RECT  59610.0 27772.5 59680.0 27907.5 ;
      RECT  59945.0 26222.5 60015.0 26357.5 ;
      RECT  59682.5 27357.5 59752.5 27492.5 ;
      RECT  59872.5 26497.5 59942.5 26632.5 ;
      RECT  60130.0 26397.5 60200.0 26532.5 ;
      RECT  59610.0 27840.0 59680.0 27980.0 ;
      RECT  59945.0 27840.0 60015.0 27980.0 ;
      RECT  59610.0 26150.0 59680.0 26290.0 ;
      RECT  59945.0 26150.0 60015.0 26290.0 ;
      RECT  59425.0 26150.0 59495.0 27980.0 ;
      RECT  60130.0 26150.0 60200.0 27980.0 ;
      RECT  60315.0 26790.0 60385.0 26860.0 ;
      RECT  60387.5 26790.0 60457.5 26860.0 ;
      RECT  60315.0 26290.0 60385.0 26825.0 ;
      RECT  60350.0 26790.0 60422.5 26860.0 ;
      RECT  60387.5 26825.0 60457.5 27357.5 ;
      RECT  60650.0 27202.5 60720.0 27272.5 ;
      RECT  60577.5 27202.5 60647.5 27272.5 ;
      RECT  60650.0 27237.5 60720.0 27840.0 ;
      RECT  60612.5 27202.5 60685.0 27272.5 ;
      RECT  60577.5 26632.5 60647.5 27237.5 ;
      RECT  60315.0 27772.5 60385.0 27907.5 ;
      RECT  60650.0 26222.5 60720.0 26357.5 ;
      RECT  60387.5 27357.5 60457.5 27492.5 ;
      RECT  60577.5 26497.5 60647.5 26632.5 ;
      RECT  60835.0 26397.5 60905.0 26532.5 ;
      RECT  60315.0 27840.0 60385.0 27980.0 ;
      RECT  60650.0 27840.0 60720.0 27980.0 ;
      RECT  60315.0 26150.0 60385.0 26290.0 ;
      RECT  60650.0 26150.0 60720.0 26290.0 ;
      RECT  60130.0 26150.0 60200.0 27980.0 ;
      RECT  60835.0 26150.0 60905.0 27980.0 ;
      RECT  61020.0 26790.0 61090.0 26860.0 ;
      RECT  61092.5 26790.0 61162.5 26860.0 ;
      RECT  61020.0 26290.0 61090.0 26825.0 ;
      RECT  61055.0 26790.0 61127.5 26860.0 ;
      RECT  61092.5 26825.0 61162.5 27357.5 ;
      RECT  61355.0 27202.5 61425.0 27272.5 ;
      RECT  61282.5 27202.5 61352.5 27272.5 ;
      RECT  61355.0 27237.5 61425.0 27840.0 ;
      RECT  61317.5 27202.5 61390.0 27272.5 ;
      RECT  61282.5 26632.5 61352.5 27237.5 ;
      RECT  61020.0 27772.5 61090.0 27907.5 ;
      RECT  61355.0 26222.5 61425.0 26357.5 ;
      RECT  61092.5 27357.5 61162.5 27492.5 ;
      RECT  61282.5 26497.5 61352.5 26632.5 ;
      RECT  61540.0 26397.5 61610.0 26532.5 ;
      RECT  61020.0 27840.0 61090.0 27980.0 ;
      RECT  61355.0 27840.0 61425.0 27980.0 ;
      RECT  61020.0 26150.0 61090.0 26290.0 ;
      RECT  61355.0 26150.0 61425.0 26290.0 ;
      RECT  60835.0 26150.0 60905.0 27980.0 ;
      RECT  61540.0 26150.0 61610.0 27980.0 ;
      RECT  61725.0 26790.0 61795.0 26860.0 ;
      RECT  61797.5 26790.0 61867.5 26860.0 ;
      RECT  61725.0 26290.0 61795.0 26825.0 ;
      RECT  61760.0 26790.0 61832.5 26860.0 ;
      RECT  61797.5 26825.0 61867.5 27357.5 ;
      RECT  62060.0 27202.5 62130.0 27272.5 ;
      RECT  61987.5 27202.5 62057.5 27272.5 ;
      RECT  62060.0 27237.5 62130.0 27840.0 ;
      RECT  62022.5 27202.5 62095.0 27272.5 ;
      RECT  61987.5 26632.5 62057.5 27237.5 ;
      RECT  61725.0 27772.5 61795.0 27907.5 ;
      RECT  62060.0 26222.5 62130.0 26357.5 ;
      RECT  61797.5 27357.5 61867.5 27492.5 ;
      RECT  61987.5 26497.5 62057.5 26632.5 ;
      RECT  62245.0 26397.5 62315.0 26532.5 ;
      RECT  61725.0 27840.0 61795.0 27980.0 ;
      RECT  62060.0 27840.0 62130.0 27980.0 ;
      RECT  61725.0 26150.0 61795.0 26290.0 ;
      RECT  62060.0 26150.0 62130.0 26290.0 ;
      RECT  61540.0 26150.0 61610.0 27980.0 ;
      RECT  62245.0 26150.0 62315.0 27980.0 ;
      RECT  62430.0 26790.0 62500.0 26860.0 ;
      RECT  62502.5 26790.0 62572.5 26860.0 ;
      RECT  62430.0 26290.0 62500.0 26825.0 ;
      RECT  62465.0 26790.0 62537.5 26860.0 ;
      RECT  62502.5 26825.0 62572.5 27357.5 ;
      RECT  62765.0 27202.5 62835.0 27272.5 ;
      RECT  62692.5 27202.5 62762.5 27272.5 ;
      RECT  62765.0 27237.5 62835.0 27840.0 ;
      RECT  62727.5 27202.5 62800.0 27272.5 ;
      RECT  62692.5 26632.5 62762.5 27237.5 ;
      RECT  62430.0 27772.5 62500.0 27907.5 ;
      RECT  62765.0 26222.5 62835.0 26357.5 ;
      RECT  62502.5 27357.5 62572.5 27492.5 ;
      RECT  62692.5 26497.5 62762.5 26632.5 ;
      RECT  62950.0 26397.5 63020.0 26532.5 ;
      RECT  62430.0 27840.0 62500.0 27980.0 ;
      RECT  62765.0 27840.0 62835.0 27980.0 ;
      RECT  62430.0 26150.0 62500.0 26290.0 ;
      RECT  62765.0 26150.0 62835.0 26290.0 ;
      RECT  62245.0 26150.0 62315.0 27980.0 ;
      RECT  62950.0 26150.0 63020.0 27980.0 ;
      RECT  63135.0 26790.0 63205.0 26860.0 ;
      RECT  63207.5 26790.0 63277.5 26860.0 ;
      RECT  63135.0 26290.0 63205.0 26825.0 ;
      RECT  63170.0 26790.0 63242.5 26860.0 ;
      RECT  63207.5 26825.0 63277.5 27357.5 ;
      RECT  63470.0 27202.5 63540.0 27272.5 ;
      RECT  63397.5 27202.5 63467.5 27272.5 ;
      RECT  63470.0 27237.5 63540.0 27840.0 ;
      RECT  63432.5 27202.5 63505.0 27272.5 ;
      RECT  63397.5 26632.5 63467.5 27237.5 ;
      RECT  63135.0 27772.5 63205.0 27907.5 ;
      RECT  63470.0 26222.5 63540.0 26357.5 ;
      RECT  63207.5 27357.5 63277.5 27492.5 ;
      RECT  63397.5 26497.5 63467.5 26632.5 ;
      RECT  63655.0 26397.5 63725.0 26532.5 ;
      RECT  63135.0 27840.0 63205.0 27980.0 ;
      RECT  63470.0 27840.0 63540.0 27980.0 ;
      RECT  63135.0 26150.0 63205.0 26290.0 ;
      RECT  63470.0 26150.0 63540.0 26290.0 ;
      RECT  62950.0 26150.0 63020.0 27980.0 ;
      RECT  63655.0 26150.0 63725.0 27980.0 ;
      RECT  63840.0 26790.0 63910.0 26860.0 ;
      RECT  63912.5 26790.0 63982.5 26860.0 ;
      RECT  63840.0 26290.0 63910.0 26825.0 ;
      RECT  63875.0 26790.0 63947.5 26860.0 ;
      RECT  63912.5 26825.0 63982.5 27357.5 ;
      RECT  64175.0 27202.5 64245.0 27272.5 ;
      RECT  64102.5 27202.5 64172.5 27272.5 ;
      RECT  64175.0 27237.5 64245.0 27840.0 ;
      RECT  64137.5 27202.5 64210.0 27272.5 ;
      RECT  64102.5 26632.5 64172.5 27237.5 ;
      RECT  63840.0 27772.5 63910.0 27907.5 ;
      RECT  64175.0 26222.5 64245.0 26357.5 ;
      RECT  63912.5 27357.5 63982.5 27492.5 ;
      RECT  64102.5 26497.5 64172.5 26632.5 ;
      RECT  64360.0 26397.5 64430.0 26532.5 ;
      RECT  63840.0 27840.0 63910.0 27980.0 ;
      RECT  64175.0 27840.0 64245.0 27980.0 ;
      RECT  63840.0 26150.0 63910.0 26290.0 ;
      RECT  64175.0 26150.0 64245.0 26290.0 ;
      RECT  63655.0 26150.0 63725.0 27980.0 ;
      RECT  64360.0 26150.0 64430.0 27980.0 ;
      RECT  64545.0 26790.0 64615.0 26860.0 ;
      RECT  64617.5 26790.0 64687.5 26860.0 ;
      RECT  64545.0 26290.0 64615.0 26825.0 ;
      RECT  64580.0 26790.0 64652.5 26860.0 ;
      RECT  64617.5 26825.0 64687.5 27357.5 ;
      RECT  64880.0 27202.5 64950.0 27272.5 ;
      RECT  64807.5 27202.5 64877.5 27272.5 ;
      RECT  64880.0 27237.5 64950.0 27840.0 ;
      RECT  64842.5 27202.5 64915.0 27272.5 ;
      RECT  64807.5 26632.5 64877.5 27237.5 ;
      RECT  64545.0 27772.5 64615.0 27907.5 ;
      RECT  64880.0 26222.5 64950.0 26357.5 ;
      RECT  64617.5 27357.5 64687.5 27492.5 ;
      RECT  64807.5 26497.5 64877.5 26632.5 ;
      RECT  65065.0 26397.5 65135.0 26532.5 ;
      RECT  64545.0 27840.0 64615.0 27980.0 ;
      RECT  64880.0 27840.0 64950.0 27980.0 ;
      RECT  64545.0 26150.0 64615.0 26290.0 ;
      RECT  64880.0 26150.0 64950.0 26290.0 ;
      RECT  64360.0 26150.0 64430.0 27980.0 ;
      RECT  65065.0 26150.0 65135.0 27980.0 ;
      RECT  65250.0 26790.0 65320.0 26860.0 ;
      RECT  65322.5 26790.0 65392.5 26860.0 ;
      RECT  65250.0 26290.0 65320.0 26825.0 ;
      RECT  65285.0 26790.0 65357.5 26860.0 ;
      RECT  65322.5 26825.0 65392.5 27357.5 ;
      RECT  65585.0 27202.5 65655.0 27272.5 ;
      RECT  65512.5 27202.5 65582.5 27272.5 ;
      RECT  65585.0 27237.5 65655.0 27840.0 ;
      RECT  65547.5 27202.5 65620.0 27272.5 ;
      RECT  65512.5 26632.5 65582.5 27237.5 ;
      RECT  65250.0 27772.5 65320.0 27907.5 ;
      RECT  65585.0 26222.5 65655.0 26357.5 ;
      RECT  65322.5 27357.5 65392.5 27492.5 ;
      RECT  65512.5 26497.5 65582.5 26632.5 ;
      RECT  65770.0 26397.5 65840.0 26532.5 ;
      RECT  65250.0 27840.0 65320.0 27980.0 ;
      RECT  65585.0 27840.0 65655.0 27980.0 ;
      RECT  65250.0 26150.0 65320.0 26290.0 ;
      RECT  65585.0 26150.0 65655.0 26290.0 ;
      RECT  65065.0 26150.0 65135.0 27980.0 ;
      RECT  65770.0 26150.0 65840.0 27980.0 ;
      RECT  65955.0 26790.0 66025.0 26860.0 ;
      RECT  66027.5 26790.0 66097.5 26860.0 ;
      RECT  65955.0 26290.0 66025.0 26825.0 ;
      RECT  65990.0 26790.0 66062.5 26860.0 ;
      RECT  66027.5 26825.0 66097.5 27357.5 ;
      RECT  66290.0 27202.5 66360.0 27272.5 ;
      RECT  66217.5 27202.5 66287.5 27272.5 ;
      RECT  66290.0 27237.5 66360.0 27840.0 ;
      RECT  66252.5 27202.5 66325.0 27272.5 ;
      RECT  66217.5 26632.5 66287.5 27237.5 ;
      RECT  65955.0 27772.5 66025.0 27907.5 ;
      RECT  66290.0 26222.5 66360.0 26357.5 ;
      RECT  66027.5 27357.5 66097.5 27492.5 ;
      RECT  66217.5 26497.5 66287.5 26632.5 ;
      RECT  66475.0 26397.5 66545.0 26532.5 ;
      RECT  65955.0 27840.0 66025.0 27980.0 ;
      RECT  66290.0 27840.0 66360.0 27980.0 ;
      RECT  65955.0 26150.0 66025.0 26290.0 ;
      RECT  66290.0 26150.0 66360.0 26290.0 ;
      RECT  65770.0 26150.0 65840.0 27980.0 ;
      RECT  66475.0 26150.0 66545.0 27980.0 ;
      RECT  66660.0 26790.0 66730.0 26860.0 ;
      RECT  66732.5 26790.0 66802.5 26860.0 ;
      RECT  66660.0 26290.0 66730.0 26825.0 ;
      RECT  66695.0 26790.0 66767.5 26860.0 ;
      RECT  66732.5 26825.0 66802.5 27357.5 ;
      RECT  66995.0 27202.5 67065.0 27272.5 ;
      RECT  66922.5 27202.5 66992.5 27272.5 ;
      RECT  66995.0 27237.5 67065.0 27840.0 ;
      RECT  66957.5 27202.5 67030.0 27272.5 ;
      RECT  66922.5 26632.5 66992.5 27237.5 ;
      RECT  66660.0 27772.5 66730.0 27907.5 ;
      RECT  66995.0 26222.5 67065.0 26357.5 ;
      RECT  66732.5 27357.5 66802.5 27492.5 ;
      RECT  66922.5 26497.5 66992.5 26632.5 ;
      RECT  67180.0 26397.5 67250.0 26532.5 ;
      RECT  66660.0 27840.0 66730.0 27980.0 ;
      RECT  66995.0 27840.0 67065.0 27980.0 ;
      RECT  66660.0 26150.0 66730.0 26290.0 ;
      RECT  66995.0 26150.0 67065.0 26290.0 ;
      RECT  66475.0 26150.0 66545.0 27980.0 ;
      RECT  67180.0 26150.0 67250.0 27980.0 ;
      RECT  67365.0 26790.0 67435.0 26860.0 ;
      RECT  67437.5 26790.0 67507.5 26860.0 ;
      RECT  67365.0 26290.0 67435.0 26825.0 ;
      RECT  67400.0 26790.0 67472.5 26860.0 ;
      RECT  67437.5 26825.0 67507.5 27357.5 ;
      RECT  67700.0 27202.5 67770.0 27272.5 ;
      RECT  67627.5 27202.5 67697.5 27272.5 ;
      RECT  67700.0 27237.5 67770.0 27840.0 ;
      RECT  67662.5 27202.5 67735.0 27272.5 ;
      RECT  67627.5 26632.5 67697.5 27237.5 ;
      RECT  67365.0 27772.5 67435.0 27907.5 ;
      RECT  67700.0 26222.5 67770.0 26357.5 ;
      RECT  67437.5 27357.5 67507.5 27492.5 ;
      RECT  67627.5 26497.5 67697.5 26632.5 ;
      RECT  67885.0 26397.5 67955.0 26532.5 ;
      RECT  67365.0 27840.0 67435.0 27980.0 ;
      RECT  67700.0 27840.0 67770.0 27980.0 ;
      RECT  67365.0 26150.0 67435.0 26290.0 ;
      RECT  67700.0 26150.0 67770.0 26290.0 ;
      RECT  67180.0 26150.0 67250.0 27980.0 ;
      RECT  67885.0 26150.0 67955.0 27980.0 ;
      RECT  68070.0 26790.0 68140.0 26860.0 ;
      RECT  68142.5 26790.0 68212.5 26860.0 ;
      RECT  68070.0 26290.0 68140.0 26825.0 ;
      RECT  68105.0 26790.0 68177.5 26860.0 ;
      RECT  68142.5 26825.0 68212.5 27357.5 ;
      RECT  68405.0 27202.5 68475.0 27272.5 ;
      RECT  68332.5 27202.5 68402.5 27272.5 ;
      RECT  68405.0 27237.5 68475.0 27840.0 ;
      RECT  68367.5 27202.5 68440.0 27272.5 ;
      RECT  68332.5 26632.5 68402.5 27237.5 ;
      RECT  68070.0 27772.5 68140.0 27907.5 ;
      RECT  68405.0 26222.5 68475.0 26357.5 ;
      RECT  68142.5 27357.5 68212.5 27492.5 ;
      RECT  68332.5 26497.5 68402.5 26632.5 ;
      RECT  68590.0 26397.5 68660.0 26532.5 ;
      RECT  68070.0 27840.0 68140.0 27980.0 ;
      RECT  68405.0 27840.0 68475.0 27980.0 ;
      RECT  68070.0 26150.0 68140.0 26290.0 ;
      RECT  68405.0 26150.0 68475.0 26290.0 ;
      RECT  67885.0 26150.0 67955.0 27980.0 ;
      RECT  68590.0 26150.0 68660.0 27980.0 ;
      RECT  68775.0 26790.0 68845.0 26860.0 ;
      RECT  68847.5 26790.0 68917.5 26860.0 ;
      RECT  68775.0 26290.0 68845.0 26825.0 ;
      RECT  68810.0 26790.0 68882.5 26860.0 ;
      RECT  68847.5 26825.0 68917.5 27357.5 ;
      RECT  69110.0 27202.5 69180.0 27272.5 ;
      RECT  69037.5 27202.5 69107.5 27272.5 ;
      RECT  69110.0 27237.5 69180.0 27840.0 ;
      RECT  69072.5 27202.5 69145.0 27272.5 ;
      RECT  69037.5 26632.5 69107.5 27237.5 ;
      RECT  68775.0 27772.5 68845.0 27907.5 ;
      RECT  69110.0 26222.5 69180.0 26357.5 ;
      RECT  68847.5 27357.5 68917.5 27492.5 ;
      RECT  69037.5 26497.5 69107.5 26632.5 ;
      RECT  69295.0 26397.5 69365.0 26532.5 ;
      RECT  68775.0 27840.0 68845.0 27980.0 ;
      RECT  69110.0 27840.0 69180.0 27980.0 ;
      RECT  68775.0 26150.0 68845.0 26290.0 ;
      RECT  69110.0 26150.0 69180.0 26290.0 ;
      RECT  68590.0 26150.0 68660.0 27980.0 ;
      RECT  69295.0 26150.0 69365.0 27980.0 ;
      RECT  69480.0 26790.0 69550.0 26860.0 ;
      RECT  69552.5 26790.0 69622.5 26860.0 ;
      RECT  69480.0 26290.0 69550.0 26825.0 ;
      RECT  69515.0 26790.0 69587.5 26860.0 ;
      RECT  69552.5 26825.0 69622.5 27357.5 ;
      RECT  69815.0 27202.5 69885.0 27272.5 ;
      RECT  69742.5 27202.5 69812.5 27272.5 ;
      RECT  69815.0 27237.5 69885.0 27840.0 ;
      RECT  69777.5 27202.5 69850.0 27272.5 ;
      RECT  69742.5 26632.5 69812.5 27237.5 ;
      RECT  69480.0 27772.5 69550.0 27907.5 ;
      RECT  69815.0 26222.5 69885.0 26357.5 ;
      RECT  69552.5 27357.5 69622.5 27492.5 ;
      RECT  69742.5 26497.5 69812.5 26632.5 ;
      RECT  70000.0 26397.5 70070.0 26532.5 ;
      RECT  69480.0 27840.0 69550.0 27980.0 ;
      RECT  69815.0 27840.0 69885.0 27980.0 ;
      RECT  69480.0 26150.0 69550.0 26290.0 ;
      RECT  69815.0 26150.0 69885.0 26290.0 ;
      RECT  69295.0 26150.0 69365.0 27980.0 ;
      RECT  70000.0 26150.0 70070.0 27980.0 ;
      RECT  70185.0 26790.0 70255.0 26860.0 ;
      RECT  70257.5 26790.0 70327.5 26860.0 ;
      RECT  70185.0 26290.0 70255.0 26825.0 ;
      RECT  70220.0 26790.0 70292.5 26860.0 ;
      RECT  70257.5 26825.0 70327.5 27357.5 ;
      RECT  70520.0 27202.5 70590.0 27272.5 ;
      RECT  70447.5 27202.5 70517.5 27272.5 ;
      RECT  70520.0 27237.5 70590.0 27840.0 ;
      RECT  70482.5 27202.5 70555.0 27272.5 ;
      RECT  70447.5 26632.5 70517.5 27237.5 ;
      RECT  70185.0 27772.5 70255.0 27907.5 ;
      RECT  70520.0 26222.5 70590.0 26357.5 ;
      RECT  70257.5 27357.5 70327.5 27492.5 ;
      RECT  70447.5 26497.5 70517.5 26632.5 ;
      RECT  70705.0 26397.5 70775.0 26532.5 ;
      RECT  70185.0 27840.0 70255.0 27980.0 ;
      RECT  70520.0 27840.0 70590.0 27980.0 ;
      RECT  70185.0 26150.0 70255.0 26290.0 ;
      RECT  70520.0 26150.0 70590.0 26290.0 ;
      RECT  70000.0 26150.0 70070.0 27980.0 ;
      RECT  70705.0 26150.0 70775.0 27980.0 ;
      RECT  70890.0 26790.0 70960.0 26860.0 ;
      RECT  70962.5 26790.0 71032.5 26860.0 ;
      RECT  70890.0 26290.0 70960.0 26825.0 ;
      RECT  70925.0 26790.0 70997.5 26860.0 ;
      RECT  70962.5 26825.0 71032.5 27357.5 ;
      RECT  71225.0 27202.5 71295.0 27272.5 ;
      RECT  71152.5 27202.5 71222.5 27272.5 ;
      RECT  71225.0 27237.5 71295.0 27840.0 ;
      RECT  71187.5 27202.5 71260.0 27272.5 ;
      RECT  71152.5 26632.5 71222.5 27237.5 ;
      RECT  70890.0 27772.5 70960.0 27907.5 ;
      RECT  71225.0 26222.5 71295.0 26357.5 ;
      RECT  70962.5 27357.5 71032.5 27492.5 ;
      RECT  71152.5 26497.5 71222.5 26632.5 ;
      RECT  71410.0 26397.5 71480.0 26532.5 ;
      RECT  70890.0 27840.0 70960.0 27980.0 ;
      RECT  71225.0 27840.0 71295.0 27980.0 ;
      RECT  70890.0 26150.0 70960.0 26290.0 ;
      RECT  71225.0 26150.0 71295.0 26290.0 ;
      RECT  70705.0 26150.0 70775.0 27980.0 ;
      RECT  71410.0 26150.0 71480.0 27980.0 ;
      RECT  71595.0 26790.0 71665.0 26860.0 ;
      RECT  71667.5 26790.0 71737.5 26860.0 ;
      RECT  71595.0 26290.0 71665.0 26825.0 ;
      RECT  71630.0 26790.0 71702.5 26860.0 ;
      RECT  71667.5 26825.0 71737.5 27357.5 ;
      RECT  71930.0 27202.5 72000.0 27272.5 ;
      RECT  71857.5 27202.5 71927.5 27272.5 ;
      RECT  71930.0 27237.5 72000.0 27840.0 ;
      RECT  71892.5 27202.5 71965.0 27272.5 ;
      RECT  71857.5 26632.5 71927.5 27237.5 ;
      RECT  71595.0 27772.5 71665.0 27907.5 ;
      RECT  71930.0 26222.5 72000.0 26357.5 ;
      RECT  71667.5 27357.5 71737.5 27492.5 ;
      RECT  71857.5 26497.5 71927.5 26632.5 ;
      RECT  72115.0 26397.5 72185.0 26532.5 ;
      RECT  71595.0 27840.0 71665.0 27980.0 ;
      RECT  71930.0 27840.0 72000.0 27980.0 ;
      RECT  71595.0 26150.0 71665.0 26290.0 ;
      RECT  71930.0 26150.0 72000.0 26290.0 ;
      RECT  71410.0 26150.0 71480.0 27980.0 ;
      RECT  72115.0 26150.0 72185.0 27980.0 ;
      RECT  72300.0 26790.0 72370.0 26860.0 ;
      RECT  72372.5 26790.0 72442.5 26860.0 ;
      RECT  72300.0 26290.0 72370.0 26825.0 ;
      RECT  72335.0 26790.0 72407.5 26860.0 ;
      RECT  72372.5 26825.0 72442.5 27357.5 ;
      RECT  72635.0 27202.5 72705.0 27272.5 ;
      RECT  72562.5 27202.5 72632.5 27272.5 ;
      RECT  72635.0 27237.5 72705.0 27840.0 ;
      RECT  72597.5 27202.5 72670.0 27272.5 ;
      RECT  72562.5 26632.5 72632.5 27237.5 ;
      RECT  72300.0 27772.5 72370.0 27907.5 ;
      RECT  72635.0 26222.5 72705.0 26357.5 ;
      RECT  72372.5 27357.5 72442.5 27492.5 ;
      RECT  72562.5 26497.5 72632.5 26632.5 ;
      RECT  72820.0 26397.5 72890.0 26532.5 ;
      RECT  72300.0 27840.0 72370.0 27980.0 ;
      RECT  72635.0 27840.0 72705.0 27980.0 ;
      RECT  72300.0 26150.0 72370.0 26290.0 ;
      RECT  72635.0 26150.0 72705.0 26290.0 ;
      RECT  72115.0 26150.0 72185.0 27980.0 ;
      RECT  72820.0 26150.0 72890.0 27980.0 ;
      RECT  73005.0 26790.0 73075.0 26860.0 ;
      RECT  73077.5 26790.0 73147.5 26860.0 ;
      RECT  73005.0 26290.0 73075.0 26825.0 ;
      RECT  73040.0 26790.0 73112.5 26860.0 ;
      RECT  73077.5 26825.0 73147.5 27357.5 ;
      RECT  73340.0 27202.5 73410.0 27272.5 ;
      RECT  73267.5 27202.5 73337.5 27272.5 ;
      RECT  73340.0 27237.5 73410.0 27840.0 ;
      RECT  73302.5 27202.5 73375.0 27272.5 ;
      RECT  73267.5 26632.5 73337.5 27237.5 ;
      RECT  73005.0 27772.5 73075.0 27907.5 ;
      RECT  73340.0 26222.5 73410.0 26357.5 ;
      RECT  73077.5 27357.5 73147.5 27492.5 ;
      RECT  73267.5 26497.5 73337.5 26632.5 ;
      RECT  73525.0 26397.5 73595.0 26532.5 ;
      RECT  73005.0 27840.0 73075.0 27980.0 ;
      RECT  73340.0 27840.0 73410.0 27980.0 ;
      RECT  73005.0 26150.0 73075.0 26290.0 ;
      RECT  73340.0 26150.0 73410.0 26290.0 ;
      RECT  72820.0 26150.0 72890.0 27980.0 ;
      RECT  73525.0 26150.0 73595.0 27980.0 ;
      RECT  73710.0 26790.0 73780.0 26860.0 ;
      RECT  73782.5 26790.0 73852.5 26860.0 ;
      RECT  73710.0 26290.0 73780.0 26825.0 ;
      RECT  73745.0 26790.0 73817.5 26860.0 ;
      RECT  73782.5 26825.0 73852.5 27357.5 ;
      RECT  74045.0 27202.5 74115.0 27272.5 ;
      RECT  73972.5 27202.5 74042.5 27272.5 ;
      RECT  74045.0 27237.5 74115.0 27840.0 ;
      RECT  74007.5 27202.5 74080.0 27272.5 ;
      RECT  73972.5 26632.5 74042.5 27237.5 ;
      RECT  73710.0 27772.5 73780.0 27907.5 ;
      RECT  74045.0 26222.5 74115.0 26357.5 ;
      RECT  73782.5 27357.5 73852.5 27492.5 ;
      RECT  73972.5 26497.5 74042.5 26632.5 ;
      RECT  74230.0 26397.5 74300.0 26532.5 ;
      RECT  73710.0 27840.0 73780.0 27980.0 ;
      RECT  74045.0 27840.0 74115.0 27980.0 ;
      RECT  73710.0 26150.0 73780.0 26290.0 ;
      RECT  74045.0 26150.0 74115.0 26290.0 ;
      RECT  73525.0 26150.0 73595.0 27980.0 ;
      RECT  74230.0 26150.0 74300.0 27980.0 ;
      RECT  74415.0 26790.0 74485.0 26860.0 ;
      RECT  74487.5 26790.0 74557.5 26860.0 ;
      RECT  74415.0 26290.0 74485.0 26825.0 ;
      RECT  74450.0 26790.0 74522.5 26860.0 ;
      RECT  74487.5 26825.0 74557.5 27357.5 ;
      RECT  74750.0 27202.5 74820.0 27272.5 ;
      RECT  74677.5 27202.5 74747.5 27272.5 ;
      RECT  74750.0 27237.5 74820.0 27840.0 ;
      RECT  74712.5 27202.5 74785.0 27272.5 ;
      RECT  74677.5 26632.5 74747.5 27237.5 ;
      RECT  74415.0 27772.5 74485.0 27907.5 ;
      RECT  74750.0 26222.5 74820.0 26357.5 ;
      RECT  74487.5 27357.5 74557.5 27492.5 ;
      RECT  74677.5 26497.5 74747.5 26632.5 ;
      RECT  74935.0 26397.5 75005.0 26532.5 ;
      RECT  74415.0 27840.0 74485.0 27980.0 ;
      RECT  74750.0 27840.0 74820.0 27980.0 ;
      RECT  74415.0 26150.0 74485.0 26290.0 ;
      RECT  74750.0 26150.0 74820.0 26290.0 ;
      RECT  74230.0 26150.0 74300.0 27980.0 ;
      RECT  74935.0 26150.0 75005.0 27980.0 ;
      RECT  75120.0 26790.0 75190.0 26860.0 ;
      RECT  75192.5 26790.0 75262.5 26860.0 ;
      RECT  75120.0 26290.0 75190.0 26825.0 ;
      RECT  75155.0 26790.0 75227.5 26860.0 ;
      RECT  75192.5 26825.0 75262.5 27357.5 ;
      RECT  75455.0 27202.5 75525.0 27272.5 ;
      RECT  75382.5 27202.5 75452.5 27272.5 ;
      RECT  75455.0 27237.5 75525.0 27840.0 ;
      RECT  75417.5 27202.5 75490.0 27272.5 ;
      RECT  75382.5 26632.5 75452.5 27237.5 ;
      RECT  75120.0 27772.5 75190.0 27907.5 ;
      RECT  75455.0 26222.5 75525.0 26357.5 ;
      RECT  75192.5 27357.5 75262.5 27492.5 ;
      RECT  75382.5 26497.5 75452.5 26632.5 ;
      RECT  75640.0 26397.5 75710.0 26532.5 ;
      RECT  75120.0 27840.0 75190.0 27980.0 ;
      RECT  75455.0 27840.0 75525.0 27980.0 ;
      RECT  75120.0 26150.0 75190.0 26290.0 ;
      RECT  75455.0 26150.0 75525.0 26290.0 ;
      RECT  74935.0 26150.0 75005.0 27980.0 ;
      RECT  75640.0 26150.0 75710.0 27980.0 ;
      RECT  75825.0 26790.0 75895.0 26860.0 ;
      RECT  75897.5 26790.0 75967.5 26860.0 ;
      RECT  75825.0 26290.0 75895.0 26825.0 ;
      RECT  75860.0 26790.0 75932.5 26860.0 ;
      RECT  75897.5 26825.0 75967.5 27357.5 ;
      RECT  76160.0 27202.5 76230.0 27272.5 ;
      RECT  76087.5 27202.5 76157.5 27272.5 ;
      RECT  76160.0 27237.5 76230.0 27840.0 ;
      RECT  76122.5 27202.5 76195.0 27272.5 ;
      RECT  76087.5 26632.5 76157.5 27237.5 ;
      RECT  75825.0 27772.5 75895.0 27907.5 ;
      RECT  76160.0 26222.5 76230.0 26357.5 ;
      RECT  75897.5 27357.5 75967.5 27492.5 ;
      RECT  76087.5 26497.5 76157.5 26632.5 ;
      RECT  76345.0 26397.5 76415.0 26532.5 ;
      RECT  75825.0 27840.0 75895.0 27980.0 ;
      RECT  76160.0 27840.0 76230.0 27980.0 ;
      RECT  75825.0 26150.0 75895.0 26290.0 ;
      RECT  76160.0 26150.0 76230.0 26290.0 ;
      RECT  75640.0 26150.0 75710.0 27980.0 ;
      RECT  76345.0 26150.0 76415.0 27980.0 ;
      RECT  76530.0 26790.0 76600.0 26860.0 ;
      RECT  76602.5 26790.0 76672.5 26860.0 ;
      RECT  76530.0 26290.0 76600.0 26825.0 ;
      RECT  76565.0 26790.0 76637.5 26860.0 ;
      RECT  76602.5 26825.0 76672.5 27357.5 ;
      RECT  76865.0 27202.5 76935.0 27272.5 ;
      RECT  76792.5 27202.5 76862.5 27272.5 ;
      RECT  76865.0 27237.5 76935.0 27840.0 ;
      RECT  76827.5 27202.5 76900.0 27272.5 ;
      RECT  76792.5 26632.5 76862.5 27237.5 ;
      RECT  76530.0 27772.5 76600.0 27907.5 ;
      RECT  76865.0 26222.5 76935.0 26357.5 ;
      RECT  76602.5 27357.5 76672.5 27492.5 ;
      RECT  76792.5 26497.5 76862.5 26632.5 ;
      RECT  77050.0 26397.5 77120.0 26532.5 ;
      RECT  76530.0 27840.0 76600.0 27980.0 ;
      RECT  76865.0 27840.0 76935.0 27980.0 ;
      RECT  76530.0 26150.0 76600.0 26290.0 ;
      RECT  76865.0 26150.0 76935.0 26290.0 ;
      RECT  76345.0 26150.0 76415.0 27980.0 ;
      RECT  77050.0 26150.0 77120.0 27980.0 ;
      RECT  77235.0 26790.0 77305.0 26860.0 ;
      RECT  77307.5 26790.0 77377.5 26860.0 ;
      RECT  77235.0 26290.0 77305.0 26825.0 ;
      RECT  77270.0 26790.0 77342.5 26860.0 ;
      RECT  77307.5 26825.0 77377.5 27357.5 ;
      RECT  77570.0 27202.5 77640.0 27272.5 ;
      RECT  77497.5 27202.5 77567.5 27272.5 ;
      RECT  77570.0 27237.5 77640.0 27840.0 ;
      RECT  77532.5 27202.5 77605.0 27272.5 ;
      RECT  77497.5 26632.5 77567.5 27237.5 ;
      RECT  77235.0 27772.5 77305.0 27907.5 ;
      RECT  77570.0 26222.5 77640.0 26357.5 ;
      RECT  77307.5 27357.5 77377.5 27492.5 ;
      RECT  77497.5 26497.5 77567.5 26632.5 ;
      RECT  77755.0 26397.5 77825.0 26532.5 ;
      RECT  77235.0 27840.0 77305.0 27980.0 ;
      RECT  77570.0 27840.0 77640.0 27980.0 ;
      RECT  77235.0 26150.0 77305.0 26290.0 ;
      RECT  77570.0 26150.0 77640.0 26290.0 ;
      RECT  77050.0 26150.0 77120.0 27980.0 ;
      RECT  77755.0 26150.0 77825.0 27980.0 ;
      RECT  77940.0 26790.0 78010.0 26860.0 ;
      RECT  78012.5 26790.0 78082.5 26860.0 ;
      RECT  77940.0 26290.0 78010.0 26825.0 ;
      RECT  77975.0 26790.0 78047.5 26860.0 ;
      RECT  78012.5 26825.0 78082.5 27357.5 ;
      RECT  78275.0 27202.5 78345.0 27272.5 ;
      RECT  78202.5 27202.5 78272.5 27272.5 ;
      RECT  78275.0 27237.5 78345.0 27840.0 ;
      RECT  78237.5 27202.5 78310.0 27272.5 ;
      RECT  78202.5 26632.5 78272.5 27237.5 ;
      RECT  77940.0 27772.5 78010.0 27907.5 ;
      RECT  78275.0 26222.5 78345.0 26357.5 ;
      RECT  78012.5 27357.5 78082.5 27492.5 ;
      RECT  78202.5 26497.5 78272.5 26632.5 ;
      RECT  78460.0 26397.5 78530.0 26532.5 ;
      RECT  77940.0 27840.0 78010.0 27980.0 ;
      RECT  78275.0 27840.0 78345.0 27980.0 ;
      RECT  77940.0 26150.0 78010.0 26290.0 ;
      RECT  78275.0 26150.0 78345.0 26290.0 ;
      RECT  77755.0 26150.0 77825.0 27980.0 ;
      RECT  78460.0 26150.0 78530.0 27980.0 ;
      RECT  78645.0 26790.0 78715.0 26860.0 ;
      RECT  78717.5 26790.0 78787.5 26860.0 ;
      RECT  78645.0 26290.0 78715.0 26825.0 ;
      RECT  78680.0 26790.0 78752.5 26860.0 ;
      RECT  78717.5 26825.0 78787.5 27357.5 ;
      RECT  78980.0 27202.5 79050.0 27272.5 ;
      RECT  78907.5 27202.5 78977.5 27272.5 ;
      RECT  78980.0 27237.5 79050.0 27840.0 ;
      RECT  78942.5 27202.5 79015.0 27272.5 ;
      RECT  78907.5 26632.5 78977.5 27237.5 ;
      RECT  78645.0 27772.5 78715.0 27907.5 ;
      RECT  78980.0 26222.5 79050.0 26357.5 ;
      RECT  78717.5 27357.5 78787.5 27492.5 ;
      RECT  78907.5 26497.5 78977.5 26632.5 ;
      RECT  79165.0 26397.5 79235.0 26532.5 ;
      RECT  78645.0 27840.0 78715.0 27980.0 ;
      RECT  78980.0 27840.0 79050.0 27980.0 ;
      RECT  78645.0 26150.0 78715.0 26290.0 ;
      RECT  78980.0 26150.0 79050.0 26290.0 ;
      RECT  78460.0 26150.0 78530.0 27980.0 ;
      RECT  79165.0 26150.0 79235.0 27980.0 ;
      RECT  79350.0 26790.0 79420.0 26860.0 ;
      RECT  79422.5 26790.0 79492.5 26860.0 ;
      RECT  79350.0 26290.0 79420.0 26825.0 ;
      RECT  79385.0 26790.0 79457.5 26860.0 ;
      RECT  79422.5 26825.0 79492.5 27357.5 ;
      RECT  79685.0 27202.5 79755.0 27272.5 ;
      RECT  79612.5 27202.5 79682.5 27272.5 ;
      RECT  79685.0 27237.5 79755.0 27840.0 ;
      RECT  79647.5 27202.5 79720.0 27272.5 ;
      RECT  79612.5 26632.5 79682.5 27237.5 ;
      RECT  79350.0 27772.5 79420.0 27907.5 ;
      RECT  79685.0 26222.5 79755.0 26357.5 ;
      RECT  79422.5 27357.5 79492.5 27492.5 ;
      RECT  79612.5 26497.5 79682.5 26632.5 ;
      RECT  79870.0 26397.5 79940.0 26532.5 ;
      RECT  79350.0 27840.0 79420.0 27980.0 ;
      RECT  79685.0 27840.0 79755.0 27980.0 ;
      RECT  79350.0 26150.0 79420.0 26290.0 ;
      RECT  79685.0 26150.0 79755.0 26290.0 ;
      RECT  79165.0 26150.0 79235.0 27980.0 ;
      RECT  79870.0 26150.0 79940.0 27980.0 ;
      RECT  80055.0 26790.0 80125.0 26860.0 ;
      RECT  80127.5 26790.0 80197.5 26860.0 ;
      RECT  80055.0 26290.0 80125.0 26825.0 ;
      RECT  80090.0 26790.0 80162.5 26860.0 ;
      RECT  80127.5 26825.0 80197.5 27357.5 ;
      RECT  80390.0 27202.5 80460.0 27272.5 ;
      RECT  80317.5 27202.5 80387.5 27272.5 ;
      RECT  80390.0 27237.5 80460.0 27840.0 ;
      RECT  80352.5 27202.5 80425.0 27272.5 ;
      RECT  80317.5 26632.5 80387.5 27237.5 ;
      RECT  80055.0 27772.5 80125.0 27907.5 ;
      RECT  80390.0 26222.5 80460.0 26357.5 ;
      RECT  80127.5 27357.5 80197.5 27492.5 ;
      RECT  80317.5 26497.5 80387.5 26632.5 ;
      RECT  80575.0 26397.5 80645.0 26532.5 ;
      RECT  80055.0 27840.0 80125.0 27980.0 ;
      RECT  80390.0 27840.0 80460.0 27980.0 ;
      RECT  80055.0 26150.0 80125.0 26290.0 ;
      RECT  80390.0 26150.0 80460.0 26290.0 ;
      RECT  79870.0 26150.0 79940.0 27980.0 ;
      RECT  80575.0 26150.0 80645.0 27980.0 ;
      RECT  80760.0 26790.0 80830.0 26860.0 ;
      RECT  80832.5 26790.0 80902.5 26860.0 ;
      RECT  80760.0 26290.0 80830.0 26825.0 ;
      RECT  80795.0 26790.0 80867.5 26860.0 ;
      RECT  80832.5 26825.0 80902.5 27357.5 ;
      RECT  81095.0 27202.5 81165.0 27272.5 ;
      RECT  81022.5 27202.5 81092.5 27272.5 ;
      RECT  81095.0 27237.5 81165.0 27840.0 ;
      RECT  81057.5 27202.5 81130.0 27272.5 ;
      RECT  81022.5 26632.5 81092.5 27237.5 ;
      RECT  80760.0 27772.5 80830.0 27907.5 ;
      RECT  81095.0 26222.5 81165.0 26357.5 ;
      RECT  80832.5 27357.5 80902.5 27492.5 ;
      RECT  81022.5 26497.5 81092.5 26632.5 ;
      RECT  81280.0 26397.5 81350.0 26532.5 ;
      RECT  80760.0 27840.0 80830.0 27980.0 ;
      RECT  81095.0 27840.0 81165.0 27980.0 ;
      RECT  80760.0 26150.0 80830.0 26290.0 ;
      RECT  81095.0 26150.0 81165.0 26290.0 ;
      RECT  80575.0 26150.0 80645.0 27980.0 ;
      RECT  81280.0 26150.0 81350.0 27980.0 ;
      RECT  81465.0 26790.0 81535.0 26860.0 ;
      RECT  81537.5 26790.0 81607.5 26860.0 ;
      RECT  81465.0 26290.0 81535.0 26825.0 ;
      RECT  81500.0 26790.0 81572.5 26860.0 ;
      RECT  81537.5 26825.0 81607.5 27357.5 ;
      RECT  81800.0 27202.5 81870.0 27272.5 ;
      RECT  81727.5 27202.5 81797.5 27272.5 ;
      RECT  81800.0 27237.5 81870.0 27840.0 ;
      RECT  81762.5 27202.5 81835.0 27272.5 ;
      RECT  81727.5 26632.5 81797.5 27237.5 ;
      RECT  81465.0 27772.5 81535.0 27907.5 ;
      RECT  81800.0 26222.5 81870.0 26357.5 ;
      RECT  81537.5 27357.5 81607.5 27492.5 ;
      RECT  81727.5 26497.5 81797.5 26632.5 ;
      RECT  81985.0 26397.5 82055.0 26532.5 ;
      RECT  81465.0 27840.0 81535.0 27980.0 ;
      RECT  81800.0 27840.0 81870.0 27980.0 ;
      RECT  81465.0 26150.0 81535.0 26290.0 ;
      RECT  81800.0 26150.0 81870.0 26290.0 ;
      RECT  81280.0 26150.0 81350.0 27980.0 ;
      RECT  81985.0 26150.0 82055.0 27980.0 ;
      RECT  82170.0 26790.0 82240.0 26860.0 ;
      RECT  82242.5 26790.0 82312.5 26860.0 ;
      RECT  82170.0 26290.0 82240.0 26825.0 ;
      RECT  82205.0 26790.0 82277.5 26860.0 ;
      RECT  82242.5 26825.0 82312.5 27357.5 ;
      RECT  82505.0 27202.5 82575.0 27272.5 ;
      RECT  82432.5 27202.5 82502.5 27272.5 ;
      RECT  82505.0 27237.5 82575.0 27840.0 ;
      RECT  82467.5 27202.5 82540.0 27272.5 ;
      RECT  82432.5 26632.5 82502.5 27237.5 ;
      RECT  82170.0 27772.5 82240.0 27907.5 ;
      RECT  82505.0 26222.5 82575.0 26357.5 ;
      RECT  82242.5 27357.5 82312.5 27492.5 ;
      RECT  82432.5 26497.5 82502.5 26632.5 ;
      RECT  82690.0 26397.5 82760.0 26532.5 ;
      RECT  82170.0 27840.0 82240.0 27980.0 ;
      RECT  82505.0 27840.0 82575.0 27980.0 ;
      RECT  82170.0 26150.0 82240.0 26290.0 ;
      RECT  82505.0 26150.0 82575.0 26290.0 ;
      RECT  81985.0 26150.0 82055.0 27980.0 ;
      RECT  82690.0 26150.0 82760.0 27980.0 ;
      RECT  82875.0 26790.0 82945.0 26860.0 ;
      RECT  82947.5 26790.0 83017.5 26860.0 ;
      RECT  82875.0 26290.0 82945.0 26825.0 ;
      RECT  82910.0 26790.0 82982.5 26860.0 ;
      RECT  82947.5 26825.0 83017.5 27357.5 ;
      RECT  83210.0 27202.5 83280.0 27272.5 ;
      RECT  83137.5 27202.5 83207.5 27272.5 ;
      RECT  83210.0 27237.5 83280.0 27840.0 ;
      RECT  83172.5 27202.5 83245.0 27272.5 ;
      RECT  83137.5 26632.5 83207.5 27237.5 ;
      RECT  82875.0 27772.5 82945.0 27907.5 ;
      RECT  83210.0 26222.5 83280.0 26357.5 ;
      RECT  82947.5 27357.5 83017.5 27492.5 ;
      RECT  83137.5 26497.5 83207.5 26632.5 ;
      RECT  83395.0 26397.5 83465.0 26532.5 ;
      RECT  82875.0 27840.0 82945.0 27980.0 ;
      RECT  83210.0 27840.0 83280.0 27980.0 ;
      RECT  82875.0 26150.0 82945.0 26290.0 ;
      RECT  83210.0 26150.0 83280.0 26290.0 ;
      RECT  82690.0 26150.0 82760.0 27980.0 ;
      RECT  83395.0 26150.0 83465.0 27980.0 ;
      RECT  83580.0 26790.0 83650.0 26860.0 ;
      RECT  83652.5 26790.0 83722.5 26860.0 ;
      RECT  83580.0 26290.0 83650.0 26825.0 ;
      RECT  83615.0 26790.0 83687.5 26860.0 ;
      RECT  83652.5 26825.0 83722.5 27357.5 ;
      RECT  83915.0 27202.5 83985.0 27272.5 ;
      RECT  83842.5 27202.5 83912.5 27272.5 ;
      RECT  83915.0 27237.5 83985.0 27840.0 ;
      RECT  83877.5 27202.5 83950.0 27272.5 ;
      RECT  83842.5 26632.5 83912.5 27237.5 ;
      RECT  83580.0 27772.5 83650.0 27907.5 ;
      RECT  83915.0 26222.5 83985.0 26357.5 ;
      RECT  83652.5 27357.5 83722.5 27492.5 ;
      RECT  83842.5 26497.5 83912.5 26632.5 ;
      RECT  84100.0 26397.5 84170.0 26532.5 ;
      RECT  83580.0 27840.0 83650.0 27980.0 ;
      RECT  83915.0 27840.0 83985.0 27980.0 ;
      RECT  83580.0 26150.0 83650.0 26290.0 ;
      RECT  83915.0 26150.0 83985.0 26290.0 ;
      RECT  83395.0 26150.0 83465.0 27980.0 ;
      RECT  84100.0 26150.0 84170.0 27980.0 ;
      RECT  84285.0 26790.0 84355.0 26860.0 ;
      RECT  84357.5 26790.0 84427.5 26860.0 ;
      RECT  84285.0 26290.0 84355.0 26825.0 ;
      RECT  84320.0 26790.0 84392.5 26860.0 ;
      RECT  84357.5 26825.0 84427.5 27357.5 ;
      RECT  84620.0 27202.5 84690.0 27272.5 ;
      RECT  84547.5 27202.5 84617.5 27272.5 ;
      RECT  84620.0 27237.5 84690.0 27840.0 ;
      RECT  84582.5 27202.5 84655.0 27272.5 ;
      RECT  84547.5 26632.5 84617.5 27237.5 ;
      RECT  84285.0 27772.5 84355.0 27907.5 ;
      RECT  84620.0 26222.5 84690.0 26357.5 ;
      RECT  84357.5 27357.5 84427.5 27492.5 ;
      RECT  84547.5 26497.5 84617.5 26632.5 ;
      RECT  84805.0 26397.5 84875.0 26532.5 ;
      RECT  84285.0 27840.0 84355.0 27980.0 ;
      RECT  84620.0 27840.0 84690.0 27980.0 ;
      RECT  84285.0 26150.0 84355.0 26290.0 ;
      RECT  84620.0 26150.0 84690.0 26290.0 ;
      RECT  84100.0 26150.0 84170.0 27980.0 ;
      RECT  84805.0 26150.0 84875.0 27980.0 ;
      RECT  84990.0 26790.0 85060.0 26860.0 ;
      RECT  85062.5 26790.0 85132.5 26860.0 ;
      RECT  84990.0 26290.0 85060.0 26825.0 ;
      RECT  85025.0 26790.0 85097.5 26860.0 ;
      RECT  85062.5 26825.0 85132.5 27357.5 ;
      RECT  85325.0 27202.5 85395.0 27272.5 ;
      RECT  85252.5 27202.5 85322.5 27272.5 ;
      RECT  85325.0 27237.5 85395.0 27840.0 ;
      RECT  85287.5 27202.5 85360.0 27272.5 ;
      RECT  85252.5 26632.5 85322.5 27237.5 ;
      RECT  84990.0 27772.5 85060.0 27907.5 ;
      RECT  85325.0 26222.5 85395.0 26357.5 ;
      RECT  85062.5 27357.5 85132.5 27492.5 ;
      RECT  85252.5 26497.5 85322.5 26632.5 ;
      RECT  85510.0 26397.5 85580.0 26532.5 ;
      RECT  84990.0 27840.0 85060.0 27980.0 ;
      RECT  85325.0 27840.0 85395.0 27980.0 ;
      RECT  84990.0 26150.0 85060.0 26290.0 ;
      RECT  85325.0 26150.0 85395.0 26290.0 ;
      RECT  84805.0 26150.0 84875.0 27980.0 ;
      RECT  85510.0 26150.0 85580.0 27980.0 ;
      RECT  85695.0 26790.0 85765.0 26860.0 ;
      RECT  85767.5 26790.0 85837.5 26860.0 ;
      RECT  85695.0 26290.0 85765.0 26825.0 ;
      RECT  85730.0 26790.0 85802.5 26860.0 ;
      RECT  85767.5 26825.0 85837.5 27357.5 ;
      RECT  86030.0 27202.5 86100.0 27272.5 ;
      RECT  85957.5 27202.5 86027.5 27272.5 ;
      RECT  86030.0 27237.5 86100.0 27840.0 ;
      RECT  85992.5 27202.5 86065.0 27272.5 ;
      RECT  85957.5 26632.5 86027.5 27237.5 ;
      RECT  85695.0 27772.5 85765.0 27907.5 ;
      RECT  86030.0 26222.5 86100.0 26357.5 ;
      RECT  85767.5 27357.5 85837.5 27492.5 ;
      RECT  85957.5 26497.5 86027.5 26632.5 ;
      RECT  86215.0 26397.5 86285.0 26532.5 ;
      RECT  85695.0 27840.0 85765.0 27980.0 ;
      RECT  86030.0 27840.0 86100.0 27980.0 ;
      RECT  85695.0 26150.0 85765.0 26290.0 ;
      RECT  86030.0 26150.0 86100.0 26290.0 ;
      RECT  85510.0 26150.0 85580.0 27980.0 ;
      RECT  86215.0 26150.0 86285.0 27980.0 ;
      RECT  86400.0 26790.0 86470.0 26860.0 ;
      RECT  86472.5 26790.0 86542.5 26860.0 ;
      RECT  86400.0 26290.0 86470.0 26825.0 ;
      RECT  86435.0 26790.0 86507.5 26860.0 ;
      RECT  86472.5 26825.0 86542.5 27357.5 ;
      RECT  86735.0 27202.5 86805.0 27272.5 ;
      RECT  86662.5 27202.5 86732.5 27272.5 ;
      RECT  86735.0 27237.5 86805.0 27840.0 ;
      RECT  86697.5 27202.5 86770.0 27272.5 ;
      RECT  86662.5 26632.5 86732.5 27237.5 ;
      RECT  86400.0 27772.5 86470.0 27907.5 ;
      RECT  86735.0 26222.5 86805.0 26357.5 ;
      RECT  86472.5 27357.5 86542.5 27492.5 ;
      RECT  86662.5 26497.5 86732.5 26632.5 ;
      RECT  86920.0 26397.5 86990.0 26532.5 ;
      RECT  86400.0 27840.0 86470.0 27980.0 ;
      RECT  86735.0 27840.0 86805.0 27980.0 ;
      RECT  86400.0 26150.0 86470.0 26290.0 ;
      RECT  86735.0 26150.0 86805.0 26290.0 ;
      RECT  86215.0 26150.0 86285.0 27980.0 ;
      RECT  86920.0 26150.0 86990.0 27980.0 ;
      RECT  87105.0 26790.0 87175.0 26860.0 ;
      RECT  87177.5 26790.0 87247.5 26860.0 ;
      RECT  87105.0 26290.0 87175.0 26825.0 ;
      RECT  87140.0 26790.0 87212.5 26860.0 ;
      RECT  87177.5 26825.0 87247.5 27357.5 ;
      RECT  87440.0 27202.5 87510.0 27272.5 ;
      RECT  87367.5 27202.5 87437.5 27272.5 ;
      RECT  87440.0 27237.5 87510.0 27840.0 ;
      RECT  87402.5 27202.5 87475.0 27272.5 ;
      RECT  87367.5 26632.5 87437.5 27237.5 ;
      RECT  87105.0 27772.5 87175.0 27907.5 ;
      RECT  87440.0 26222.5 87510.0 26357.5 ;
      RECT  87177.5 27357.5 87247.5 27492.5 ;
      RECT  87367.5 26497.5 87437.5 26632.5 ;
      RECT  87625.0 26397.5 87695.0 26532.5 ;
      RECT  87105.0 27840.0 87175.0 27980.0 ;
      RECT  87440.0 27840.0 87510.0 27980.0 ;
      RECT  87105.0 26150.0 87175.0 26290.0 ;
      RECT  87440.0 26150.0 87510.0 26290.0 ;
      RECT  86920.0 26150.0 86990.0 27980.0 ;
      RECT  87625.0 26150.0 87695.0 27980.0 ;
      RECT  87810.0 26790.0 87880.0 26860.0 ;
      RECT  87882.5 26790.0 87952.5 26860.0 ;
      RECT  87810.0 26290.0 87880.0 26825.0 ;
      RECT  87845.0 26790.0 87917.5 26860.0 ;
      RECT  87882.5 26825.0 87952.5 27357.5 ;
      RECT  88145.0 27202.5 88215.0 27272.5 ;
      RECT  88072.5 27202.5 88142.5 27272.5 ;
      RECT  88145.0 27237.5 88215.0 27840.0 ;
      RECT  88107.5 27202.5 88180.0 27272.5 ;
      RECT  88072.5 26632.5 88142.5 27237.5 ;
      RECT  87810.0 27772.5 87880.0 27907.5 ;
      RECT  88145.0 26222.5 88215.0 26357.5 ;
      RECT  87882.5 27357.5 87952.5 27492.5 ;
      RECT  88072.5 26497.5 88142.5 26632.5 ;
      RECT  88330.0 26397.5 88400.0 26532.5 ;
      RECT  87810.0 27840.0 87880.0 27980.0 ;
      RECT  88145.0 27840.0 88215.0 27980.0 ;
      RECT  87810.0 26150.0 87880.0 26290.0 ;
      RECT  88145.0 26150.0 88215.0 26290.0 ;
      RECT  87625.0 26150.0 87695.0 27980.0 ;
      RECT  88330.0 26150.0 88400.0 27980.0 ;
      RECT  88515.0 26790.0 88585.0 26860.0 ;
      RECT  88587.5 26790.0 88657.5 26860.0 ;
      RECT  88515.0 26290.0 88585.0 26825.0 ;
      RECT  88550.0 26790.0 88622.5 26860.0 ;
      RECT  88587.5 26825.0 88657.5 27357.5 ;
      RECT  88850.0 27202.5 88920.0 27272.5 ;
      RECT  88777.5 27202.5 88847.5 27272.5 ;
      RECT  88850.0 27237.5 88920.0 27840.0 ;
      RECT  88812.5 27202.5 88885.0 27272.5 ;
      RECT  88777.5 26632.5 88847.5 27237.5 ;
      RECT  88515.0 27772.5 88585.0 27907.5 ;
      RECT  88850.0 26222.5 88920.0 26357.5 ;
      RECT  88587.5 27357.5 88657.5 27492.5 ;
      RECT  88777.5 26497.5 88847.5 26632.5 ;
      RECT  89035.0 26397.5 89105.0 26532.5 ;
      RECT  88515.0 27840.0 88585.0 27980.0 ;
      RECT  88850.0 27840.0 88920.0 27980.0 ;
      RECT  88515.0 26150.0 88585.0 26290.0 ;
      RECT  88850.0 26150.0 88920.0 26290.0 ;
      RECT  88330.0 26150.0 88400.0 27980.0 ;
      RECT  89035.0 26150.0 89105.0 27980.0 ;
      RECT  89220.0 26790.0 89290.0 26860.0 ;
      RECT  89292.5 26790.0 89362.5 26860.0 ;
      RECT  89220.0 26290.0 89290.0 26825.0 ;
      RECT  89255.0 26790.0 89327.5 26860.0 ;
      RECT  89292.5 26825.0 89362.5 27357.5 ;
      RECT  89555.0 27202.5 89625.0 27272.5 ;
      RECT  89482.5 27202.5 89552.5 27272.5 ;
      RECT  89555.0 27237.5 89625.0 27840.0 ;
      RECT  89517.5 27202.5 89590.0 27272.5 ;
      RECT  89482.5 26632.5 89552.5 27237.5 ;
      RECT  89220.0 27772.5 89290.0 27907.5 ;
      RECT  89555.0 26222.5 89625.0 26357.5 ;
      RECT  89292.5 27357.5 89362.5 27492.5 ;
      RECT  89482.5 26497.5 89552.5 26632.5 ;
      RECT  89740.0 26397.5 89810.0 26532.5 ;
      RECT  89220.0 27840.0 89290.0 27980.0 ;
      RECT  89555.0 27840.0 89625.0 27980.0 ;
      RECT  89220.0 26150.0 89290.0 26290.0 ;
      RECT  89555.0 26150.0 89625.0 26290.0 ;
      RECT  89035.0 26150.0 89105.0 27980.0 ;
      RECT  89740.0 26150.0 89810.0 27980.0 ;
      RECT  89925.0 26790.0 89995.0 26860.0 ;
      RECT  89997.5 26790.0 90067.5 26860.0 ;
      RECT  89925.0 26290.0 89995.0 26825.0 ;
      RECT  89960.0 26790.0 90032.5 26860.0 ;
      RECT  89997.5 26825.0 90067.5 27357.5 ;
      RECT  90260.0 27202.5 90330.0 27272.5 ;
      RECT  90187.5 27202.5 90257.5 27272.5 ;
      RECT  90260.0 27237.5 90330.0 27840.0 ;
      RECT  90222.5 27202.5 90295.0 27272.5 ;
      RECT  90187.5 26632.5 90257.5 27237.5 ;
      RECT  89925.0 27772.5 89995.0 27907.5 ;
      RECT  90260.0 26222.5 90330.0 26357.5 ;
      RECT  89997.5 27357.5 90067.5 27492.5 ;
      RECT  90187.5 26497.5 90257.5 26632.5 ;
      RECT  90445.0 26397.5 90515.0 26532.5 ;
      RECT  89925.0 27840.0 89995.0 27980.0 ;
      RECT  90260.0 27840.0 90330.0 27980.0 ;
      RECT  89925.0 26150.0 89995.0 26290.0 ;
      RECT  90260.0 26150.0 90330.0 26290.0 ;
      RECT  89740.0 26150.0 89810.0 27980.0 ;
      RECT  90445.0 26150.0 90515.0 27980.0 ;
      RECT  90630.0 26790.0 90700.0 26860.0 ;
      RECT  90702.5 26790.0 90772.5 26860.0 ;
      RECT  90630.0 26290.0 90700.0 26825.0 ;
      RECT  90665.0 26790.0 90737.5 26860.0 ;
      RECT  90702.5 26825.0 90772.5 27357.5 ;
      RECT  90965.0 27202.5 91035.0 27272.5 ;
      RECT  90892.5 27202.5 90962.5 27272.5 ;
      RECT  90965.0 27237.5 91035.0 27840.0 ;
      RECT  90927.5 27202.5 91000.0 27272.5 ;
      RECT  90892.5 26632.5 90962.5 27237.5 ;
      RECT  90630.0 27772.5 90700.0 27907.5 ;
      RECT  90965.0 26222.5 91035.0 26357.5 ;
      RECT  90702.5 27357.5 90772.5 27492.5 ;
      RECT  90892.5 26497.5 90962.5 26632.5 ;
      RECT  91150.0 26397.5 91220.0 26532.5 ;
      RECT  90630.0 27840.0 90700.0 27980.0 ;
      RECT  90965.0 27840.0 91035.0 27980.0 ;
      RECT  90630.0 26150.0 90700.0 26290.0 ;
      RECT  90965.0 26150.0 91035.0 26290.0 ;
      RECT  90445.0 26150.0 90515.0 27980.0 ;
      RECT  91150.0 26150.0 91220.0 27980.0 ;
      RECT  91335.0 26790.0 91405.0 26860.0 ;
      RECT  91407.5 26790.0 91477.5 26860.0 ;
      RECT  91335.0 26290.0 91405.0 26825.0 ;
      RECT  91370.0 26790.0 91442.5 26860.0 ;
      RECT  91407.5 26825.0 91477.5 27357.5 ;
      RECT  91670.0 27202.5 91740.0 27272.5 ;
      RECT  91597.5 27202.5 91667.5 27272.5 ;
      RECT  91670.0 27237.5 91740.0 27840.0 ;
      RECT  91632.5 27202.5 91705.0 27272.5 ;
      RECT  91597.5 26632.5 91667.5 27237.5 ;
      RECT  91335.0 27772.5 91405.0 27907.5 ;
      RECT  91670.0 26222.5 91740.0 26357.5 ;
      RECT  91407.5 27357.5 91477.5 27492.5 ;
      RECT  91597.5 26497.5 91667.5 26632.5 ;
      RECT  91855.0 26397.5 91925.0 26532.5 ;
      RECT  91335.0 27840.0 91405.0 27980.0 ;
      RECT  91670.0 27840.0 91740.0 27980.0 ;
      RECT  91335.0 26150.0 91405.0 26290.0 ;
      RECT  91670.0 26150.0 91740.0 26290.0 ;
      RECT  91150.0 26150.0 91220.0 27980.0 ;
      RECT  91855.0 26150.0 91925.0 27980.0 ;
      RECT  92040.0 26790.0 92110.0 26860.0 ;
      RECT  92112.5 26790.0 92182.5 26860.0 ;
      RECT  92040.0 26290.0 92110.0 26825.0 ;
      RECT  92075.0 26790.0 92147.5 26860.0 ;
      RECT  92112.5 26825.0 92182.5 27357.5 ;
      RECT  92375.0 27202.5 92445.0 27272.5 ;
      RECT  92302.5 27202.5 92372.5 27272.5 ;
      RECT  92375.0 27237.5 92445.0 27840.0 ;
      RECT  92337.5 27202.5 92410.0 27272.5 ;
      RECT  92302.5 26632.5 92372.5 27237.5 ;
      RECT  92040.0 27772.5 92110.0 27907.5 ;
      RECT  92375.0 26222.5 92445.0 26357.5 ;
      RECT  92112.5 27357.5 92182.5 27492.5 ;
      RECT  92302.5 26497.5 92372.5 26632.5 ;
      RECT  92560.0 26397.5 92630.0 26532.5 ;
      RECT  92040.0 27840.0 92110.0 27980.0 ;
      RECT  92375.0 27840.0 92445.0 27980.0 ;
      RECT  92040.0 26150.0 92110.0 26290.0 ;
      RECT  92375.0 26150.0 92445.0 26290.0 ;
      RECT  91855.0 26150.0 91925.0 27980.0 ;
      RECT  92560.0 26150.0 92630.0 27980.0 ;
      RECT  92745.0 26790.0 92815.0 26860.0 ;
      RECT  92817.5 26790.0 92887.5 26860.0 ;
      RECT  92745.0 26290.0 92815.0 26825.0 ;
      RECT  92780.0 26790.0 92852.5 26860.0 ;
      RECT  92817.5 26825.0 92887.5 27357.5 ;
      RECT  93080.0 27202.5 93150.0 27272.5 ;
      RECT  93007.5 27202.5 93077.5 27272.5 ;
      RECT  93080.0 27237.5 93150.0 27840.0 ;
      RECT  93042.5 27202.5 93115.0 27272.5 ;
      RECT  93007.5 26632.5 93077.5 27237.5 ;
      RECT  92745.0 27772.5 92815.0 27907.5 ;
      RECT  93080.0 26222.5 93150.0 26357.5 ;
      RECT  92817.5 27357.5 92887.5 27492.5 ;
      RECT  93007.5 26497.5 93077.5 26632.5 ;
      RECT  93265.0 26397.5 93335.0 26532.5 ;
      RECT  92745.0 27840.0 92815.0 27980.0 ;
      RECT  93080.0 27840.0 93150.0 27980.0 ;
      RECT  92745.0 26150.0 92815.0 26290.0 ;
      RECT  93080.0 26150.0 93150.0 26290.0 ;
      RECT  92560.0 26150.0 92630.0 27980.0 ;
      RECT  93265.0 26150.0 93335.0 27980.0 ;
      RECT  93450.0 26790.0 93520.0 26860.0 ;
      RECT  93522.5 26790.0 93592.5 26860.0 ;
      RECT  93450.0 26290.0 93520.0 26825.0 ;
      RECT  93485.0 26790.0 93557.5 26860.0 ;
      RECT  93522.5 26825.0 93592.5 27357.5 ;
      RECT  93785.0 27202.5 93855.0 27272.5 ;
      RECT  93712.5 27202.5 93782.5 27272.5 ;
      RECT  93785.0 27237.5 93855.0 27840.0 ;
      RECT  93747.5 27202.5 93820.0 27272.5 ;
      RECT  93712.5 26632.5 93782.5 27237.5 ;
      RECT  93450.0 27772.5 93520.0 27907.5 ;
      RECT  93785.0 26222.5 93855.0 26357.5 ;
      RECT  93522.5 27357.5 93592.5 27492.5 ;
      RECT  93712.5 26497.5 93782.5 26632.5 ;
      RECT  93970.0 26397.5 94040.0 26532.5 ;
      RECT  93450.0 27840.0 93520.0 27980.0 ;
      RECT  93785.0 27840.0 93855.0 27980.0 ;
      RECT  93450.0 26150.0 93520.0 26290.0 ;
      RECT  93785.0 26150.0 93855.0 26290.0 ;
      RECT  93265.0 26150.0 93335.0 27980.0 ;
      RECT  93970.0 26150.0 94040.0 27980.0 ;
      RECT  94155.0 26790.0 94225.0 26860.0 ;
      RECT  94227.5 26790.0 94297.5 26860.0 ;
      RECT  94155.0 26290.0 94225.0 26825.0 ;
      RECT  94190.0 26790.0 94262.5 26860.0 ;
      RECT  94227.5 26825.0 94297.5 27357.5 ;
      RECT  94490.0 27202.5 94560.0 27272.5 ;
      RECT  94417.5 27202.5 94487.5 27272.5 ;
      RECT  94490.0 27237.5 94560.0 27840.0 ;
      RECT  94452.5 27202.5 94525.0 27272.5 ;
      RECT  94417.5 26632.5 94487.5 27237.5 ;
      RECT  94155.0 27772.5 94225.0 27907.5 ;
      RECT  94490.0 26222.5 94560.0 26357.5 ;
      RECT  94227.5 27357.5 94297.5 27492.5 ;
      RECT  94417.5 26497.5 94487.5 26632.5 ;
      RECT  94675.0 26397.5 94745.0 26532.5 ;
      RECT  94155.0 27840.0 94225.0 27980.0 ;
      RECT  94490.0 27840.0 94560.0 27980.0 ;
      RECT  94155.0 26150.0 94225.0 26290.0 ;
      RECT  94490.0 26150.0 94560.0 26290.0 ;
      RECT  93970.0 26150.0 94040.0 27980.0 ;
      RECT  94675.0 26150.0 94745.0 27980.0 ;
      RECT  94860.0 26790.0 94930.0 26860.0 ;
      RECT  94932.5 26790.0 95002.5 26860.0 ;
      RECT  94860.0 26290.0 94930.0 26825.0 ;
      RECT  94895.0 26790.0 94967.5 26860.0 ;
      RECT  94932.5 26825.0 95002.5 27357.5 ;
      RECT  95195.0 27202.5 95265.0 27272.5 ;
      RECT  95122.5 27202.5 95192.5 27272.5 ;
      RECT  95195.0 27237.5 95265.0 27840.0 ;
      RECT  95157.5 27202.5 95230.0 27272.5 ;
      RECT  95122.5 26632.5 95192.5 27237.5 ;
      RECT  94860.0 27772.5 94930.0 27907.5 ;
      RECT  95195.0 26222.5 95265.0 26357.5 ;
      RECT  94932.5 27357.5 95002.5 27492.5 ;
      RECT  95122.5 26497.5 95192.5 26632.5 ;
      RECT  95380.0 26397.5 95450.0 26532.5 ;
      RECT  94860.0 27840.0 94930.0 27980.0 ;
      RECT  95195.0 27840.0 95265.0 27980.0 ;
      RECT  94860.0 26150.0 94930.0 26290.0 ;
      RECT  95195.0 26150.0 95265.0 26290.0 ;
      RECT  94675.0 26150.0 94745.0 27980.0 ;
      RECT  95380.0 26150.0 95450.0 27980.0 ;
      RECT  95565.0 26790.0 95635.0 26860.0 ;
      RECT  95637.5 26790.0 95707.5 26860.0 ;
      RECT  95565.0 26290.0 95635.0 26825.0 ;
      RECT  95600.0 26790.0 95672.5 26860.0 ;
      RECT  95637.5 26825.0 95707.5 27357.5 ;
      RECT  95900.0 27202.5 95970.0 27272.5 ;
      RECT  95827.5 27202.5 95897.5 27272.5 ;
      RECT  95900.0 27237.5 95970.0 27840.0 ;
      RECT  95862.5 27202.5 95935.0 27272.5 ;
      RECT  95827.5 26632.5 95897.5 27237.5 ;
      RECT  95565.0 27772.5 95635.0 27907.5 ;
      RECT  95900.0 26222.5 95970.0 26357.5 ;
      RECT  95637.5 27357.5 95707.5 27492.5 ;
      RECT  95827.5 26497.5 95897.5 26632.5 ;
      RECT  96085.0 26397.5 96155.0 26532.5 ;
      RECT  95565.0 27840.0 95635.0 27980.0 ;
      RECT  95900.0 27840.0 95970.0 27980.0 ;
      RECT  95565.0 26150.0 95635.0 26290.0 ;
      RECT  95900.0 26150.0 95970.0 26290.0 ;
      RECT  95380.0 26150.0 95450.0 27980.0 ;
      RECT  96085.0 26150.0 96155.0 27980.0 ;
      RECT  96270.0 26790.0 96340.0 26860.0 ;
      RECT  96342.5 26790.0 96412.5 26860.0 ;
      RECT  96270.0 26290.0 96340.0 26825.0 ;
      RECT  96305.0 26790.0 96377.5 26860.0 ;
      RECT  96342.5 26825.0 96412.5 27357.5 ;
      RECT  96605.0 27202.5 96675.0 27272.5 ;
      RECT  96532.5 27202.5 96602.5 27272.5 ;
      RECT  96605.0 27237.5 96675.0 27840.0 ;
      RECT  96567.5 27202.5 96640.0 27272.5 ;
      RECT  96532.5 26632.5 96602.5 27237.5 ;
      RECT  96270.0 27772.5 96340.0 27907.5 ;
      RECT  96605.0 26222.5 96675.0 26357.5 ;
      RECT  96342.5 27357.5 96412.5 27492.5 ;
      RECT  96532.5 26497.5 96602.5 26632.5 ;
      RECT  96790.0 26397.5 96860.0 26532.5 ;
      RECT  96270.0 27840.0 96340.0 27980.0 ;
      RECT  96605.0 27840.0 96675.0 27980.0 ;
      RECT  96270.0 26150.0 96340.0 26290.0 ;
      RECT  96605.0 26150.0 96675.0 26290.0 ;
      RECT  96085.0 26150.0 96155.0 27980.0 ;
      RECT  96790.0 26150.0 96860.0 27980.0 ;
      RECT  96975.0 26790.0 97045.0 26860.0 ;
      RECT  97047.5 26790.0 97117.5 26860.0 ;
      RECT  96975.0 26290.0 97045.0 26825.0 ;
      RECT  97010.0 26790.0 97082.5 26860.0 ;
      RECT  97047.5 26825.0 97117.5 27357.5 ;
      RECT  97310.0 27202.5 97380.0 27272.5 ;
      RECT  97237.5 27202.5 97307.5 27272.5 ;
      RECT  97310.0 27237.5 97380.0 27840.0 ;
      RECT  97272.5 27202.5 97345.0 27272.5 ;
      RECT  97237.5 26632.5 97307.5 27237.5 ;
      RECT  96975.0 27772.5 97045.0 27907.5 ;
      RECT  97310.0 26222.5 97380.0 26357.5 ;
      RECT  97047.5 27357.5 97117.5 27492.5 ;
      RECT  97237.5 26497.5 97307.5 26632.5 ;
      RECT  97495.0 26397.5 97565.0 26532.5 ;
      RECT  96975.0 27840.0 97045.0 27980.0 ;
      RECT  97310.0 27840.0 97380.0 27980.0 ;
      RECT  96975.0 26150.0 97045.0 26290.0 ;
      RECT  97310.0 26150.0 97380.0 26290.0 ;
      RECT  96790.0 26150.0 96860.0 27980.0 ;
      RECT  97495.0 26150.0 97565.0 27980.0 ;
      RECT  97680.0 26790.0 97750.0 26860.0 ;
      RECT  97752.5 26790.0 97822.5 26860.0 ;
      RECT  97680.0 26290.0 97750.0 26825.0 ;
      RECT  97715.0 26790.0 97787.5 26860.0 ;
      RECT  97752.5 26825.0 97822.5 27357.5 ;
      RECT  98015.0 27202.5 98085.0 27272.5 ;
      RECT  97942.5 27202.5 98012.5 27272.5 ;
      RECT  98015.0 27237.5 98085.0 27840.0 ;
      RECT  97977.5 27202.5 98050.0 27272.5 ;
      RECT  97942.5 26632.5 98012.5 27237.5 ;
      RECT  97680.0 27772.5 97750.0 27907.5 ;
      RECT  98015.0 26222.5 98085.0 26357.5 ;
      RECT  97752.5 27357.5 97822.5 27492.5 ;
      RECT  97942.5 26497.5 98012.5 26632.5 ;
      RECT  98200.0 26397.5 98270.0 26532.5 ;
      RECT  97680.0 27840.0 97750.0 27980.0 ;
      RECT  98015.0 27840.0 98085.0 27980.0 ;
      RECT  97680.0 26150.0 97750.0 26290.0 ;
      RECT  98015.0 26150.0 98085.0 26290.0 ;
      RECT  97495.0 26150.0 97565.0 27980.0 ;
      RECT  98200.0 26150.0 98270.0 27980.0 ;
      RECT  98385.0 26790.0 98455.0 26860.0 ;
      RECT  98457.5 26790.0 98527.5 26860.0 ;
      RECT  98385.0 26290.0 98455.0 26825.0 ;
      RECT  98420.0 26790.0 98492.5 26860.0 ;
      RECT  98457.5 26825.0 98527.5 27357.5 ;
      RECT  98720.0 27202.5 98790.0 27272.5 ;
      RECT  98647.5 27202.5 98717.5 27272.5 ;
      RECT  98720.0 27237.5 98790.0 27840.0 ;
      RECT  98682.5 27202.5 98755.0 27272.5 ;
      RECT  98647.5 26632.5 98717.5 27237.5 ;
      RECT  98385.0 27772.5 98455.0 27907.5 ;
      RECT  98720.0 26222.5 98790.0 26357.5 ;
      RECT  98457.5 27357.5 98527.5 27492.5 ;
      RECT  98647.5 26497.5 98717.5 26632.5 ;
      RECT  98905.0 26397.5 98975.0 26532.5 ;
      RECT  98385.0 27840.0 98455.0 27980.0 ;
      RECT  98720.0 27840.0 98790.0 27980.0 ;
      RECT  98385.0 26150.0 98455.0 26290.0 ;
      RECT  98720.0 26150.0 98790.0 26290.0 ;
      RECT  98200.0 26150.0 98270.0 27980.0 ;
      RECT  98905.0 26150.0 98975.0 27980.0 ;
      RECT  99090.0 26790.0 99160.0 26860.0 ;
      RECT  99162.5 26790.0 99232.5 26860.0 ;
      RECT  99090.0 26290.0 99160.0 26825.0 ;
      RECT  99125.0 26790.0 99197.5 26860.0 ;
      RECT  99162.5 26825.0 99232.5 27357.5 ;
      RECT  99425.0 27202.5 99495.0 27272.5 ;
      RECT  99352.5 27202.5 99422.5 27272.5 ;
      RECT  99425.0 27237.5 99495.0 27840.0 ;
      RECT  99387.5 27202.5 99460.0 27272.5 ;
      RECT  99352.5 26632.5 99422.5 27237.5 ;
      RECT  99090.0 27772.5 99160.0 27907.5 ;
      RECT  99425.0 26222.5 99495.0 26357.5 ;
      RECT  99162.5 27357.5 99232.5 27492.5 ;
      RECT  99352.5 26497.5 99422.5 26632.5 ;
      RECT  99610.0 26397.5 99680.0 26532.5 ;
      RECT  99090.0 27840.0 99160.0 27980.0 ;
      RECT  99425.0 27840.0 99495.0 27980.0 ;
      RECT  99090.0 26150.0 99160.0 26290.0 ;
      RECT  99425.0 26150.0 99495.0 26290.0 ;
      RECT  98905.0 26150.0 98975.0 27980.0 ;
      RECT  99610.0 26150.0 99680.0 27980.0 ;
      RECT  99795.0 26790.0 99865.0 26860.0 ;
      RECT  99867.5 26790.0 99937.5 26860.0 ;
      RECT  99795.0 26290.0 99865.0 26825.0 ;
      RECT  99830.0 26790.0 99902.5 26860.0 ;
      RECT  99867.5 26825.0 99937.5 27357.5 ;
      RECT  100130.0 27202.5 100200.0 27272.5 ;
      RECT  100057.5 27202.5 100127.5 27272.5 ;
      RECT  100130.0 27237.5 100200.0 27840.0 ;
      RECT  100092.5 27202.5 100165.0 27272.5 ;
      RECT  100057.5 26632.5 100127.5 27237.5 ;
      RECT  99795.0 27772.5 99865.0 27907.5 ;
      RECT  100130.0 26222.5 100200.0 26357.5 ;
      RECT  99867.5 27357.5 99937.5 27492.5 ;
      RECT  100057.5 26497.5 100127.5 26632.5 ;
      RECT  100315.0 26397.5 100385.0 26532.5 ;
      RECT  99795.0 27840.0 99865.0 27980.0 ;
      RECT  100130.0 27840.0 100200.0 27980.0 ;
      RECT  99795.0 26150.0 99865.0 26290.0 ;
      RECT  100130.0 26150.0 100200.0 26290.0 ;
      RECT  99610.0 26150.0 99680.0 27980.0 ;
      RECT  100315.0 26150.0 100385.0 27980.0 ;
      RECT  100500.0 26790.0 100570.0 26860.0 ;
      RECT  100572.5 26790.0 100642.5 26860.0 ;
      RECT  100500.0 26290.0 100570.0 26825.0 ;
      RECT  100535.0 26790.0 100607.5 26860.0 ;
      RECT  100572.5 26825.0 100642.5 27357.5 ;
      RECT  100835.0 27202.5 100905.0 27272.5 ;
      RECT  100762.5 27202.5 100832.5 27272.5 ;
      RECT  100835.0 27237.5 100905.0 27840.0 ;
      RECT  100797.5 27202.5 100870.0 27272.5 ;
      RECT  100762.5 26632.5 100832.5 27237.5 ;
      RECT  100500.0 27772.5 100570.0 27907.5 ;
      RECT  100835.0 26222.5 100905.0 26357.5 ;
      RECT  100572.5 27357.5 100642.5 27492.5 ;
      RECT  100762.5 26497.5 100832.5 26632.5 ;
      RECT  101020.0 26397.5 101090.0 26532.5 ;
      RECT  100500.0 27840.0 100570.0 27980.0 ;
      RECT  100835.0 27840.0 100905.0 27980.0 ;
      RECT  100500.0 26150.0 100570.0 26290.0 ;
      RECT  100835.0 26150.0 100905.0 26290.0 ;
      RECT  100315.0 26150.0 100385.0 27980.0 ;
      RECT  101020.0 26150.0 101090.0 27980.0 ;
      RECT  101205.0 26790.0 101275.0 26860.0 ;
      RECT  101277.5 26790.0 101347.5 26860.0 ;
      RECT  101205.0 26290.0 101275.0 26825.0 ;
      RECT  101240.0 26790.0 101312.5 26860.0 ;
      RECT  101277.5 26825.0 101347.5 27357.5 ;
      RECT  101540.0 27202.5 101610.0 27272.5 ;
      RECT  101467.5 27202.5 101537.5 27272.5 ;
      RECT  101540.0 27237.5 101610.0 27840.0 ;
      RECT  101502.5 27202.5 101575.0 27272.5 ;
      RECT  101467.5 26632.5 101537.5 27237.5 ;
      RECT  101205.0 27772.5 101275.0 27907.5 ;
      RECT  101540.0 26222.5 101610.0 26357.5 ;
      RECT  101277.5 27357.5 101347.5 27492.5 ;
      RECT  101467.5 26497.5 101537.5 26632.5 ;
      RECT  101725.0 26397.5 101795.0 26532.5 ;
      RECT  101205.0 27840.0 101275.0 27980.0 ;
      RECT  101540.0 27840.0 101610.0 27980.0 ;
      RECT  101205.0 26150.0 101275.0 26290.0 ;
      RECT  101540.0 26150.0 101610.0 26290.0 ;
      RECT  101020.0 26150.0 101090.0 27980.0 ;
      RECT  101725.0 26150.0 101795.0 27980.0 ;
      RECT  101910.0 26790.0 101980.0 26860.0 ;
      RECT  101982.5 26790.0 102052.5 26860.0 ;
      RECT  101910.0 26290.0 101980.0 26825.0 ;
      RECT  101945.0 26790.0 102017.5 26860.0 ;
      RECT  101982.5 26825.0 102052.5 27357.5 ;
      RECT  102245.0 27202.5 102315.0 27272.5 ;
      RECT  102172.5 27202.5 102242.5 27272.5 ;
      RECT  102245.0 27237.5 102315.0 27840.0 ;
      RECT  102207.5 27202.5 102280.0 27272.5 ;
      RECT  102172.5 26632.5 102242.5 27237.5 ;
      RECT  101910.0 27772.5 101980.0 27907.5 ;
      RECT  102245.0 26222.5 102315.0 26357.5 ;
      RECT  101982.5 27357.5 102052.5 27492.5 ;
      RECT  102172.5 26497.5 102242.5 26632.5 ;
      RECT  102430.0 26397.5 102500.0 26532.5 ;
      RECT  101910.0 27840.0 101980.0 27980.0 ;
      RECT  102245.0 27840.0 102315.0 27980.0 ;
      RECT  101910.0 26150.0 101980.0 26290.0 ;
      RECT  102245.0 26150.0 102315.0 26290.0 ;
      RECT  101725.0 26150.0 101795.0 27980.0 ;
      RECT  102430.0 26150.0 102500.0 27980.0 ;
      RECT  102615.0 26790.0 102685.0 26860.0 ;
      RECT  102687.5 26790.0 102757.5 26860.0 ;
      RECT  102615.0 26290.0 102685.0 26825.0 ;
      RECT  102650.0 26790.0 102722.5 26860.0 ;
      RECT  102687.5 26825.0 102757.5 27357.5 ;
      RECT  102950.0 27202.5 103020.0 27272.5 ;
      RECT  102877.5 27202.5 102947.5 27272.5 ;
      RECT  102950.0 27237.5 103020.0 27840.0 ;
      RECT  102912.5 27202.5 102985.0 27272.5 ;
      RECT  102877.5 26632.5 102947.5 27237.5 ;
      RECT  102615.0 27772.5 102685.0 27907.5 ;
      RECT  102950.0 26222.5 103020.0 26357.5 ;
      RECT  102687.5 27357.5 102757.5 27492.5 ;
      RECT  102877.5 26497.5 102947.5 26632.5 ;
      RECT  103135.0 26397.5 103205.0 26532.5 ;
      RECT  102615.0 27840.0 102685.0 27980.0 ;
      RECT  102950.0 27840.0 103020.0 27980.0 ;
      RECT  102615.0 26150.0 102685.0 26290.0 ;
      RECT  102950.0 26150.0 103020.0 26290.0 ;
      RECT  102430.0 26150.0 102500.0 27980.0 ;
      RECT  103135.0 26150.0 103205.0 27980.0 ;
      RECT  103320.0 26790.0 103390.0 26860.0 ;
      RECT  103392.5 26790.0 103462.5 26860.0 ;
      RECT  103320.0 26290.0 103390.0 26825.0 ;
      RECT  103355.0 26790.0 103427.5 26860.0 ;
      RECT  103392.5 26825.0 103462.5 27357.5 ;
      RECT  103655.0 27202.5 103725.0 27272.5 ;
      RECT  103582.5 27202.5 103652.5 27272.5 ;
      RECT  103655.0 27237.5 103725.0 27840.0 ;
      RECT  103617.5 27202.5 103690.0 27272.5 ;
      RECT  103582.5 26632.5 103652.5 27237.5 ;
      RECT  103320.0 27772.5 103390.0 27907.5 ;
      RECT  103655.0 26222.5 103725.0 26357.5 ;
      RECT  103392.5 27357.5 103462.5 27492.5 ;
      RECT  103582.5 26497.5 103652.5 26632.5 ;
      RECT  103840.0 26397.5 103910.0 26532.5 ;
      RECT  103320.0 27840.0 103390.0 27980.0 ;
      RECT  103655.0 27840.0 103725.0 27980.0 ;
      RECT  103320.0 26150.0 103390.0 26290.0 ;
      RECT  103655.0 26150.0 103725.0 26290.0 ;
      RECT  103135.0 26150.0 103205.0 27980.0 ;
      RECT  103840.0 26150.0 103910.0 27980.0 ;
      RECT  104025.0 26790.0 104095.0 26860.0 ;
      RECT  104097.5 26790.0 104167.5 26860.0 ;
      RECT  104025.0 26290.0 104095.0 26825.0 ;
      RECT  104060.0 26790.0 104132.5 26860.0 ;
      RECT  104097.5 26825.0 104167.5 27357.5 ;
      RECT  104360.0 27202.5 104430.0 27272.5 ;
      RECT  104287.5 27202.5 104357.5 27272.5 ;
      RECT  104360.0 27237.5 104430.0 27840.0 ;
      RECT  104322.5 27202.5 104395.0 27272.5 ;
      RECT  104287.5 26632.5 104357.5 27237.5 ;
      RECT  104025.0 27772.5 104095.0 27907.5 ;
      RECT  104360.0 26222.5 104430.0 26357.5 ;
      RECT  104097.5 27357.5 104167.5 27492.5 ;
      RECT  104287.5 26497.5 104357.5 26632.5 ;
      RECT  104545.0 26397.5 104615.0 26532.5 ;
      RECT  104025.0 27840.0 104095.0 27980.0 ;
      RECT  104360.0 27840.0 104430.0 27980.0 ;
      RECT  104025.0 26150.0 104095.0 26290.0 ;
      RECT  104360.0 26150.0 104430.0 26290.0 ;
      RECT  103840.0 26150.0 103910.0 27980.0 ;
      RECT  104545.0 26150.0 104615.0 27980.0 ;
      RECT  104730.0 26790.0 104800.0 26860.0 ;
      RECT  104802.5 26790.0 104872.5 26860.0 ;
      RECT  104730.0 26290.0 104800.0 26825.0 ;
      RECT  104765.0 26790.0 104837.5 26860.0 ;
      RECT  104802.5 26825.0 104872.5 27357.5 ;
      RECT  105065.0 27202.5 105135.0 27272.5 ;
      RECT  104992.5 27202.5 105062.5 27272.5 ;
      RECT  105065.0 27237.5 105135.0 27840.0 ;
      RECT  105027.5 27202.5 105100.0 27272.5 ;
      RECT  104992.5 26632.5 105062.5 27237.5 ;
      RECT  104730.0 27772.5 104800.0 27907.5 ;
      RECT  105065.0 26222.5 105135.0 26357.5 ;
      RECT  104802.5 27357.5 104872.5 27492.5 ;
      RECT  104992.5 26497.5 105062.5 26632.5 ;
      RECT  105250.0 26397.5 105320.0 26532.5 ;
      RECT  104730.0 27840.0 104800.0 27980.0 ;
      RECT  105065.0 27840.0 105135.0 27980.0 ;
      RECT  104730.0 26150.0 104800.0 26290.0 ;
      RECT  105065.0 26150.0 105135.0 26290.0 ;
      RECT  104545.0 26150.0 104615.0 27980.0 ;
      RECT  105250.0 26150.0 105320.0 27980.0 ;
      RECT  105435.0 26790.0 105505.0 26860.0 ;
      RECT  105507.5 26790.0 105577.5 26860.0 ;
      RECT  105435.0 26290.0 105505.0 26825.0 ;
      RECT  105470.0 26790.0 105542.5 26860.0 ;
      RECT  105507.5 26825.0 105577.5 27357.5 ;
      RECT  105770.0 27202.5 105840.0 27272.5 ;
      RECT  105697.5 27202.5 105767.5 27272.5 ;
      RECT  105770.0 27237.5 105840.0 27840.0 ;
      RECT  105732.5 27202.5 105805.0 27272.5 ;
      RECT  105697.5 26632.5 105767.5 27237.5 ;
      RECT  105435.0 27772.5 105505.0 27907.5 ;
      RECT  105770.0 26222.5 105840.0 26357.5 ;
      RECT  105507.5 27357.5 105577.5 27492.5 ;
      RECT  105697.5 26497.5 105767.5 26632.5 ;
      RECT  105955.0 26397.5 106025.0 26532.5 ;
      RECT  105435.0 27840.0 105505.0 27980.0 ;
      RECT  105770.0 27840.0 105840.0 27980.0 ;
      RECT  105435.0 26150.0 105505.0 26290.0 ;
      RECT  105770.0 26150.0 105840.0 26290.0 ;
      RECT  105250.0 26150.0 105320.0 27980.0 ;
      RECT  105955.0 26150.0 106025.0 27980.0 ;
      RECT  16035.0 25450.0 15900.0 25520.0 ;
      RECT  16235.0 25310.0 16100.0 25380.0 ;
      RECT  16740.0 25450.0 16605.0 25520.0 ;
      RECT  16940.0 25310.0 16805.0 25380.0 ;
      RECT  17445.0 25450.0 17310.0 25520.0 ;
      RECT  17645.0 25310.0 17510.0 25380.0 ;
      RECT  18150.0 25450.0 18015.0 25520.0 ;
      RECT  18350.0 25310.0 18215.0 25380.0 ;
      RECT  18855.0 25450.0 18720.0 25520.0 ;
      RECT  19055.0 25310.0 18920.0 25380.0 ;
      RECT  19560.0 25450.0 19425.0 25520.0 ;
      RECT  19760.0 25310.0 19625.0 25380.0 ;
      RECT  20265.0 25450.0 20130.0 25520.0 ;
      RECT  20465.0 25310.0 20330.0 25380.0 ;
      RECT  20970.0 25450.0 20835.0 25520.0 ;
      RECT  21170.0 25310.0 21035.0 25380.0 ;
      RECT  21675.0 25450.0 21540.0 25520.0 ;
      RECT  21875.0 25310.0 21740.0 25380.0 ;
      RECT  22380.0 25450.0 22245.0 25520.0 ;
      RECT  22580.0 25310.0 22445.0 25380.0 ;
      RECT  23085.0 25450.0 22950.0 25520.0 ;
      RECT  23285.0 25310.0 23150.0 25380.0 ;
      RECT  23790.0 25450.0 23655.0 25520.0 ;
      RECT  23990.0 25310.0 23855.0 25380.0 ;
      RECT  24495.0 25450.0 24360.0 25520.0 ;
      RECT  24695.0 25310.0 24560.0 25380.0 ;
      RECT  25200.0 25450.0 25065.0 25520.0 ;
      RECT  25400.0 25310.0 25265.0 25380.0 ;
      RECT  25905.0 25450.0 25770.0 25520.0 ;
      RECT  26105.0 25310.0 25970.0 25380.0 ;
      RECT  26610.0 25450.0 26475.0 25520.0 ;
      RECT  26810.0 25310.0 26675.0 25380.0 ;
      RECT  27315.0 25450.0 27180.0 25520.0 ;
      RECT  27515.0 25310.0 27380.0 25380.0 ;
      RECT  28020.0 25450.0 27885.0 25520.0 ;
      RECT  28220.0 25310.0 28085.0 25380.0 ;
      RECT  28725.0 25450.0 28590.0 25520.0 ;
      RECT  28925.0 25310.0 28790.0 25380.0 ;
      RECT  29430.0 25450.0 29295.0 25520.0 ;
      RECT  29630.0 25310.0 29495.0 25380.0 ;
      RECT  30135.0 25450.0 30000.0 25520.0 ;
      RECT  30335.0 25310.0 30200.0 25380.0 ;
      RECT  30840.0 25450.0 30705.0 25520.0 ;
      RECT  31040.0 25310.0 30905.0 25380.0 ;
      RECT  31545.0 25450.0 31410.0 25520.0 ;
      RECT  31745.0 25310.0 31610.0 25380.0 ;
      RECT  32250.0 25450.0 32115.0 25520.0 ;
      RECT  32450.0 25310.0 32315.0 25380.0 ;
      RECT  32955.0 25450.0 32820.0 25520.0 ;
      RECT  33155.0 25310.0 33020.0 25380.0 ;
      RECT  33660.0 25450.0 33525.0 25520.0 ;
      RECT  33860.0 25310.0 33725.0 25380.0 ;
      RECT  34365.0 25450.0 34230.0 25520.0 ;
      RECT  34565.0 25310.0 34430.0 25380.0 ;
      RECT  35070.0 25450.0 34935.0 25520.0 ;
      RECT  35270.0 25310.0 35135.0 25380.0 ;
      RECT  35775.0 25450.0 35640.0 25520.0 ;
      RECT  35975.0 25310.0 35840.0 25380.0 ;
      RECT  36480.0 25450.0 36345.0 25520.0 ;
      RECT  36680.0 25310.0 36545.0 25380.0 ;
      RECT  37185.0 25450.0 37050.0 25520.0 ;
      RECT  37385.0 25310.0 37250.0 25380.0 ;
      RECT  37890.0 25450.0 37755.0 25520.0 ;
      RECT  38090.0 25310.0 37955.0 25380.0 ;
      RECT  38595.0 25450.0 38460.0 25520.0 ;
      RECT  38795.0 25310.0 38660.0 25380.0 ;
      RECT  39300.0 25450.0 39165.0 25520.0 ;
      RECT  39500.0 25310.0 39365.0 25380.0 ;
      RECT  40005.0 25450.0 39870.0 25520.0 ;
      RECT  40205.0 25310.0 40070.0 25380.0 ;
      RECT  40710.0 25450.0 40575.0 25520.0 ;
      RECT  40910.0 25310.0 40775.0 25380.0 ;
      RECT  41415.0 25450.0 41280.0 25520.0 ;
      RECT  41615.0 25310.0 41480.0 25380.0 ;
      RECT  42120.0 25450.0 41985.0 25520.0 ;
      RECT  42320.0 25310.0 42185.0 25380.0 ;
      RECT  42825.0 25450.0 42690.0 25520.0 ;
      RECT  43025.0 25310.0 42890.0 25380.0 ;
      RECT  43530.0 25450.0 43395.0 25520.0 ;
      RECT  43730.0 25310.0 43595.0 25380.0 ;
      RECT  44235.0 25450.0 44100.0 25520.0 ;
      RECT  44435.0 25310.0 44300.0 25380.0 ;
      RECT  44940.0 25450.0 44805.0 25520.0 ;
      RECT  45140.0 25310.0 45005.0 25380.0 ;
      RECT  45645.0 25450.0 45510.0 25520.0 ;
      RECT  45845.0 25310.0 45710.0 25380.0 ;
      RECT  46350.0 25450.0 46215.0 25520.0 ;
      RECT  46550.0 25310.0 46415.0 25380.0 ;
      RECT  47055.0 25450.0 46920.0 25520.0 ;
      RECT  47255.0 25310.0 47120.0 25380.0 ;
      RECT  47760.0 25450.0 47625.0 25520.0 ;
      RECT  47960.0 25310.0 47825.0 25380.0 ;
      RECT  48465.0 25450.0 48330.0 25520.0 ;
      RECT  48665.0 25310.0 48530.0 25380.0 ;
      RECT  49170.0 25450.0 49035.0 25520.0 ;
      RECT  49370.0 25310.0 49235.0 25380.0 ;
      RECT  49875.0 25450.0 49740.0 25520.0 ;
      RECT  50075.0 25310.0 49940.0 25380.0 ;
      RECT  50580.0 25450.0 50445.0 25520.0 ;
      RECT  50780.0 25310.0 50645.0 25380.0 ;
      RECT  51285.0 25450.0 51150.0 25520.0 ;
      RECT  51485.0 25310.0 51350.0 25380.0 ;
      RECT  51990.0 25450.0 51855.0 25520.0 ;
      RECT  52190.0 25310.0 52055.0 25380.0 ;
      RECT  52695.0 25450.0 52560.0 25520.0 ;
      RECT  52895.0 25310.0 52760.0 25380.0 ;
      RECT  53400.0 25450.0 53265.0 25520.0 ;
      RECT  53600.0 25310.0 53465.0 25380.0 ;
      RECT  54105.0 25450.0 53970.0 25520.0 ;
      RECT  54305.0 25310.0 54170.0 25380.0 ;
      RECT  54810.0 25450.0 54675.0 25520.0 ;
      RECT  55010.0 25310.0 54875.0 25380.0 ;
      RECT  55515.0 25450.0 55380.0 25520.0 ;
      RECT  55715.0 25310.0 55580.0 25380.0 ;
      RECT  56220.0 25450.0 56085.0 25520.0 ;
      RECT  56420.0 25310.0 56285.0 25380.0 ;
      RECT  56925.0 25450.0 56790.0 25520.0 ;
      RECT  57125.0 25310.0 56990.0 25380.0 ;
      RECT  57630.0 25450.0 57495.0 25520.0 ;
      RECT  57830.0 25310.0 57695.0 25380.0 ;
      RECT  58335.0 25450.0 58200.0 25520.0 ;
      RECT  58535.0 25310.0 58400.0 25380.0 ;
      RECT  59040.0 25450.0 58905.0 25520.0 ;
      RECT  59240.0 25310.0 59105.0 25380.0 ;
      RECT  59745.0 25450.0 59610.0 25520.0 ;
      RECT  59945.0 25310.0 59810.0 25380.0 ;
      RECT  60450.0 25450.0 60315.0 25520.0 ;
      RECT  60650.0 25310.0 60515.0 25380.0 ;
      RECT  61155.0 25450.0 61020.0 25520.0 ;
      RECT  61355.0 25310.0 61220.0 25380.0 ;
      RECT  61860.0 25450.0 61725.0 25520.0 ;
      RECT  62060.0 25310.0 61925.0 25380.0 ;
      RECT  62565.0 25450.0 62430.0 25520.0 ;
      RECT  62765.0 25310.0 62630.0 25380.0 ;
      RECT  63270.0 25450.0 63135.0 25520.0 ;
      RECT  63470.0 25310.0 63335.0 25380.0 ;
      RECT  63975.0 25450.0 63840.0 25520.0 ;
      RECT  64175.0 25310.0 64040.0 25380.0 ;
      RECT  64680.0 25450.0 64545.0 25520.0 ;
      RECT  64880.0 25310.0 64745.0 25380.0 ;
      RECT  65385.0 25450.0 65250.0 25520.0 ;
      RECT  65585.0 25310.0 65450.0 25380.0 ;
      RECT  66090.0 25450.0 65955.0 25520.0 ;
      RECT  66290.0 25310.0 66155.0 25380.0 ;
      RECT  66795.0 25450.0 66660.0 25520.0 ;
      RECT  66995.0 25310.0 66860.0 25380.0 ;
      RECT  67500.0 25450.0 67365.0 25520.0 ;
      RECT  67700.0 25310.0 67565.0 25380.0 ;
      RECT  68205.0 25450.0 68070.0 25520.0 ;
      RECT  68405.0 25310.0 68270.0 25380.0 ;
      RECT  68910.0 25450.0 68775.0 25520.0 ;
      RECT  69110.0 25310.0 68975.0 25380.0 ;
      RECT  69615.0 25450.0 69480.0 25520.0 ;
      RECT  69815.0 25310.0 69680.0 25380.0 ;
      RECT  70320.0 25450.0 70185.0 25520.0 ;
      RECT  70520.0 25310.0 70385.0 25380.0 ;
      RECT  71025.0 25450.0 70890.0 25520.0 ;
      RECT  71225.0 25310.0 71090.0 25380.0 ;
      RECT  71730.0 25450.0 71595.0 25520.0 ;
      RECT  71930.0 25310.0 71795.0 25380.0 ;
      RECT  72435.0 25450.0 72300.0 25520.0 ;
      RECT  72635.0 25310.0 72500.0 25380.0 ;
      RECT  73140.0 25450.0 73005.0 25520.0 ;
      RECT  73340.0 25310.0 73205.0 25380.0 ;
      RECT  73845.0 25450.0 73710.0 25520.0 ;
      RECT  74045.0 25310.0 73910.0 25380.0 ;
      RECT  74550.0 25450.0 74415.0 25520.0 ;
      RECT  74750.0 25310.0 74615.0 25380.0 ;
      RECT  75255.0 25450.0 75120.0 25520.0 ;
      RECT  75455.0 25310.0 75320.0 25380.0 ;
      RECT  75960.0 25450.0 75825.0 25520.0 ;
      RECT  76160.0 25310.0 76025.0 25380.0 ;
      RECT  76665.0 25450.0 76530.0 25520.0 ;
      RECT  76865.0 25310.0 76730.0 25380.0 ;
      RECT  77370.0 25450.0 77235.0 25520.0 ;
      RECT  77570.0 25310.0 77435.0 25380.0 ;
      RECT  78075.0 25450.0 77940.0 25520.0 ;
      RECT  78275.0 25310.0 78140.0 25380.0 ;
      RECT  78780.0 25450.0 78645.0 25520.0 ;
      RECT  78980.0 25310.0 78845.0 25380.0 ;
      RECT  79485.0 25450.0 79350.0 25520.0 ;
      RECT  79685.0 25310.0 79550.0 25380.0 ;
      RECT  80190.0 25450.0 80055.0 25520.0 ;
      RECT  80390.0 25310.0 80255.0 25380.0 ;
      RECT  80895.0 25450.0 80760.0 25520.0 ;
      RECT  81095.0 25310.0 80960.0 25380.0 ;
      RECT  81600.0 25450.0 81465.0 25520.0 ;
      RECT  81800.0 25310.0 81665.0 25380.0 ;
      RECT  82305.0 25450.0 82170.0 25520.0 ;
      RECT  82505.0 25310.0 82370.0 25380.0 ;
      RECT  83010.0 25450.0 82875.0 25520.0 ;
      RECT  83210.0 25310.0 83075.0 25380.0 ;
      RECT  83715.0 25450.0 83580.0 25520.0 ;
      RECT  83915.0 25310.0 83780.0 25380.0 ;
      RECT  84420.0 25450.0 84285.0 25520.0 ;
      RECT  84620.0 25310.0 84485.0 25380.0 ;
      RECT  85125.0 25450.0 84990.0 25520.0 ;
      RECT  85325.0 25310.0 85190.0 25380.0 ;
      RECT  85830.0 25450.0 85695.0 25520.0 ;
      RECT  86030.0 25310.0 85895.0 25380.0 ;
      RECT  86535.0 25450.0 86400.0 25520.0 ;
      RECT  86735.0 25310.0 86600.0 25380.0 ;
      RECT  87240.0 25450.0 87105.0 25520.0 ;
      RECT  87440.0 25310.0 87305.0 25380.0 ;
      RECT  87945.0 25450.0 87810.0 25520.0 ;
      RECT  88145.0 25310.0 88010.0 25380.0 ;
      RECT  88650.0 25450.0 88515.0 25520.0 ;
      RECT  88850.0 25310.0 88715.0 25380.0 ;
      RECT  89355.0 25450.0 89220.0 25520.0 ;
      RECT  89555.0 25310.0 89420.0 25380.0 ;
      RECT  90060.0 25450.0 89925.0 25520.0 ;
      RECT  90260.0 25310.0 90125.0 25380.0 ;
      RECT  90765.0 25450.0 90630.0 25520.0 ;
      RECT  90965.0 25310.0 90830.0 25380.0 ;
      RECT  91470.0 25450.0 91335.0 25520.0 ;
      RECT  91670.0 25310.0 91535.0 25380.0 ;
      RECT  92175.0 25450.0 92040.0 25520.0 ;
      RECT  92375.0 25310.0 92240.0 25380.0 ;
      RECT  92880.0 25450.0 92745.0 25520.0 ;
      RECT  93080.0 25310.0 92945.0 25380.0 ;
      RECT  93585.0 25450.0 93450.0 25520.0 ;
      RECT  93785.0 25310.0 93650.0 25380.0 ;
      RECT  94290.0 25450.0 94155.0 25520.0 ;
      RECT  94490.0 25310.0 94355.0 25380.0 ;
      RECT  94995.0 25450.0 94860.0 25520.0 ;
      RECT  95195.0 25310.0 95060.0 25380.0 ;
      RECT  95700.0 25450.0 95565.0 25520.0 ;
      RECT  95900.0 25310.0 95765.0 25380.0 ;
      RECT  96405.0 25450.0 96270.0 25520.0 ;
      RECT  96605.0 25310.0 96470.0 25380.0 ;
      RECT  97110.0 25450.0 96975.0 25520.0 ;
      RECT  97310.0 25310.0 97175.0 25380.0 ;
      RECT  97815.0 25450.0 97680.0 25520.0 ;
      RECT  98015.0 25310.0 97880.0 25380.0 ;
      RECT  98520.0 25450.0 98385.0 25520.0 ;
      RECT  98720.0 25310.0 98585.0 25380.0 ;
      RECT  99225.0 25450.0 99090.0 25520.0 ;
      RECT  99425.0 25310.0 99290.0 25380.0 ;
      RECT  99930.0 25450.0 99795.0 25520.0 ;
      RECT  100130.0 25310.0 99995.0 25380.0 ;
      RECT  100635.0 25450.0 100500.0 25520.0 ;
      RECT  100835.0 25310.0 100700.0 25380.0 ;
      RECT  101340.0 25450.0 101205.0 25520.0 ;
      RECT  101540.0 25310.0 101405.0 25380.0 ;
      RECT  102045.0 25450.0 101910.0 25520.0 ;
      RECT  102245.0 25310.0 102110.0 25380.0 ;
      RECT  102750.0 25450.0 102615.0 25520.0 ;
      RECT  102950.0 25310.0 102815.0 25380.0 ;
      RECT  103455.0 25450.0 103320.0 25520.0 ;
      RECT  103655.0 25310.0 103520.0 25380.0 ;
      RECT  104160.0 25450.0 104025.0 25520.0 ;
      RECT  104360.0 25310.0 104225.0 25380.0 ;
      RECT  104865.0 25450.0 104730.0 25520.0 ;
      RECT  105065.0 25310.0 104930.0 25380.0 ;
      RECT  105570.0 25450.0 105435.0 25520.0 ;
      RECT  105770.0 25310.0 105635.0 25380.0 ;
      RECT  15900.0 27840.0 15970.0 27980.0 ;
      RECT  16235.0 27840.0 16305.0 27980.0 ;
      RECT  16605.0 27840.0 16675.0 27980.0 ;
      RECT  16940.0 27840.0 17010.0 27980.0 ;
      RECT  17310.0 27840.0 17380.0 27980.0 ;
      RECT  17645.0 27840.0 17715.0 27980.0 ;
      RECT  18015.0 27840.0 18085.0 27980.0 ;
      RECT  18350.0 27840.0 18420.0 27980.0 ;
      RECT  18720.0 27840.0 18790.0 27980.0 ;
      RECT  19055.0 27840.0 19125.0 27980.0 ;
      RECT  19425.0 27840.0 19495.0 27980.0 ;
      RECT  19760.0 27840.0 19830.0 27980.0 ;
      RECT  20130.0 27840.0 20200.0 27980.0 ;
      RECT  20465.0 27840.0 20535.0 27980.0 ;
      RECT  20835.0 27840.0 20905.0 27980.0 ;
      RECT  21170.0 27840.0 21240.0 27980.0 ;
      RECT  21540.0 27840.0 21610.0 27980.0 ;
      RECT  21875.0 27840.0 21945.0 27980.0 ;
      RECT  22245.0 27840.0 22315.0 27980.0 ;
      RECT  22580.0 27840.0 22650.0 27980.0 ;
      RECT  22950.0 27840.0 23020.0 27980.0 ;
      RECT  23285.0 27840.0 23355.0 27980.0 ;
      RECT  23655.0 27840.0 23725.0 27980.0 ;
      RECT  23990.0 27840.0 24060.0 27980.0 ;
      RECT  24360.0 27840.0 24430.0 27980.0 ;
      RECT  24695.0 27840.0 24765.0 27980.0 ;
      RECT  25065.0 27840.0 25135.0 27980.0 ;
      RECT  25400.0 27840.0 25470.0 27980.0 ;
      RECT  25770.0 27840.0 25840.0 27980.0 ;
      RECT  26105.0 27840.0 26175.0 27980.0 ;
      RECT  26475.0 27840.0 26545.0 27980.0 ;
      RECT  26810.0 27840.0 26880.0 27980.0 ;
      RECT  27180.0 27840.0 27250.0 27980.0 ;
      RECT  27515.0 27840.0 27585.0 27980.0 ;
      RECT  27885.0 27840.0 27955.0 27980.0 ;
      RECT  28220.0 27840.0 28290.0 27980.0 ;
      RECT  28590.0 27840.0 28660.0 27980.0 ;
      RECT  28925.0 27840.0 28995.0 27980.0 ;
      RECT  29295.0 27840.0 29365.0 27980.0 ;
      RECT  29630.0 27840.0 29700.0 27980.0 ;
      RECT  30000.0 27840.0 30070.0 27980.0 ;
      RECT  30335.0 27840.0 30405.0 27980.0 ;
      RECT  30705.0 27840.0 30775.0 27980.0 ;
      RECT  31040.0 27840.0 31110.0 27980.0 ;
      RECT  31410.0 27840.0 31480.0 27980.0 ;
      RECT  31745.0 27840.0 31815.0 27980.0 ;
      RECT  32115.0 27840.0 32185.0 27980.0 ;
      RECT  32450.0 27840.0 32520.0 27980.0 ;
      RECT  32820.0 27840.0 32890.0 27980.0 ;
      RECT  33155.0 27840.0 33225.0 27980.0 ;
      RECT  33525.0 27840.0 33595.0 27980.0 ;
      RECT  33860.0 27840.0 33930.0 27980.0 ;
      RECT  34230.0 27840.0 34300.0 27980.0 ;
      RECT  34565.0 27840.0 34635.0 27980.0 ;
      RECT  34935.0 27840.0 35005.0 27980.0 ;
      RECT  35270.0 27840.0 35340.0 27980.0 ;
      RECT  35640.0 27840.0 35710.0 27980.0 ;
      RECT  35975.0 27840.0 36045.0 27980.0 ;
      RECT  36345.0 27840.0 36415.0 27980.0 ;
      RECT  36680.0 27840.0 36750.0 27980.0 ;
      RECT  37050.0 27840.0 37120.0 27980.0 ;
      RECT  37385.0 27840.0 37455.0 27980.0 ;
      RECT  37755.0 27840.0 37825.0 27980.0 ;
      RECT  38090.0 27840.0 38160.0 27980.0 ;
      RECT  38460.0 27840.0 38530.0 27980.0 ;
      RECT  38795.0 27840.0 38865.0 27980.0 ;
      RECT  39165.0 27840.0 39235.0 27980.0 ;
      RECT  39500.0 27840.0 39570.0 27980.0 ;
      RECT  39870.0 27840.0 39940.0 27980.0 ;
      RECT  40205.0 27840.0 40275.0 27980.0 ;
      RECT  40575.0 27840.0 40645.0 27980.0 ;
      RECT  40910.0 27840.0 40980.0 27980.0 ;
      RECT  41280.0 27840.0 41350.0 27980.0 ;
      RECT  41615.0 27840.0 41685.0 27980.0 ;
      RECT  41985.0 27840.0 42055.0 27980.0 ;
      RECT  42320.0 27840.0 42390.0 27980.0 ;
      RECT  42690.0 27840.0 42760.0 27980.0 ;
      RECT  43025.0 27840.0 43095.0 27980.0 ;
      RECT  43395.0 27840.0 43465.0 27980.0 ;
      RECT  43730.0 27840.0 43800.0 27980.0 ;
      RECT  44100.0 27840.0 44170.0 27980.0 ;
      RECT  44435.0 27840.0 44505.0 27980.0 ;
      RECT  44805.0 27840.0 44875.0 27980.0 ;
      RECT  45140.0 27840.0 45210.0 27980.0 ;
      RECT  45510.0 27840.0 45580.0 27980.0 ;
      RECT  45845.0 27840.0 45915.0 27980.0 ;
      RECT  46215.0 27840.0 46285.0 27980.0 ;
      RECT  46550.0 27840.0 46620.0 27980.0 ;
      RECT  46920.0 27840.0 46990.0 27980.0 ;
      RECT  47255.0 27840.0 47325.0 27980.0 ;
      RECT  47625.0 27840.0 47695.0 27980.0 ;
      RECT  47960.0 27840.0 48030.0 27980.0 ;
      RECT  48330.0 27840.0 48400.0 27980.0 ;
      RECT  48665.0 27840.0 48735.0 27980.0 ;
      RECT  49035.0 27840.0 49105.0 27980.0 ;
      RECT  49370.0 27840.0 49440.0 27980.0 ;
      RECT  49740.0 27840.0 49810.0 27980.0 ;
      RECT  50075.0 27840.0 50145.0 27980.0 ;
      RECT  50445.0 27840.0 50515.0 27980.0 ;
      RECT  50780.0 27840.0 50850.0 27980.0 ;
      RECT  51150.0 27840.0 51220.0 27980.0 ;
      RECT  51485.0 27840.0 51555.0 27980.0 ;
      RECT  51855.0 27840.0 51925.0 27980.0 ;
      RECT  52190.0 27840.0 52260.0 27980.0 ;
      RECT  52560.0 27840.0 52630.0 27980.0 ;
      RECT  52895.0 27840.0 52965.0 27980.0 ;
      RECT  53265.0 27840.0 53335.0 27980.0 ;
      RECT  53600.0 27840.0 53670.0 27980.0 ;
      RECT  53970.0 27840.0 54040.0 27980.0 ;
      RECT  54305.0 27840.0 54375.0 27980.0 ;
      RECT  54675.0 27840.0 54745.0 27980.0 ;
      RECT  55010.0 27840.0 55080.0 27980.0 ;
      RECT  55380.0 27840.0 55450.0 27980.0 ;
      RECT  55715.0 27840.0 55785.0 27980.0 ;
      RECT  56085.0 27840.0 56155.0 27980.0 ;
      RECT  56420.0 27840.0 56490.0 27980.0 ;
      RECT  56790.0 27840.0 56860.0 27980.0 ;
      RECT  57125.0 27840.0 57195.0 27980.0 ;
      RECT  57495.0 27840.0 57565.0 27980.0 ;
      RECT  57830.0 27840.0 57900.0 27980.0 ;
      RECT  58200.0 27840.0 58270.0 27980.0 ;
      RECT  58535.0 27840.0 58605.0 27980.0 ;
      RECT  58905.0 27840.0 58975.0 27980.0 ;
      RECT  59240.0 27840.0 59310.0 27980.0 ;
      RECT  59610.0 27840.0 59680.0 27980.0 ;
      RECT  59945.0 27840.0 60015.0 27980.0 ;
      RECT  60315.0 27840.0 60385.0 27980.0 ;
      RECT  60650.0 27840.0 60720.0 27980.0 ;
      RECT  61020.0 27840.0 61090.0 27980.0 ;
      RECT  61355.0 27840.0 61425.0 27980.0 ;
      RECT  61725.0 27840.0 61795.0 27980.0 ;
      RECT  62060.0 27840.0 62130.0 27980.0 ;
      RECT  62430.0 27840.0 62500.0 27980.0 ;
      RECT  62765.0 27840.0 62835.0 27980.0 ;
      RECT  63135.0 27840.0 63205.0 27980.0 ;
      RECT  63470.0 27840.0 63540.0 27980.0 ;
      RECT  63840.0 27840.0 63910.0 27980.0 ;
      RECT  64175.0 27840.0 64245.0 27980.0 ;
      RECT  64545.0 27840.0 64615.0 27980.0 ;
      RECT  64880.0 27840.0 64950.0 27980.0 ;
      RECT  65250.0 27840.0 65320.0 27980.0 ;
      RECT  65585.0 27840.0 65655.0 27980.0 ;
      RECT  65955.0 27840.0 66025.0 27980.0 ;
      RECT  66290.0 27840.0 66360.0 27980.0 ;
      RECT  66660.0 27840.0 66730.0 27980.0 ;
      RECT  66995.0 27840.0 67065.0 27980.0 ;
      RECT  67365.0 27840.0 67435.0 27980.0 ;
      RECT  67700.0 27840.0 67770.0 27980.0 ;
      RECT  68070.0 27840.0 68140.0 27980.0 ;
      RECT  68405.0 27840.0 68475.0 27980.0 ;
      RECT  68775.0 27840.0 68845.0 27980.0 ;
      RECT  69110.0 27840.0 69180.0 27980.0 ;
      RECT  69480.0 27840.0 69550.0 27980.0 ;
      RECT  69815.0 27840.0 69885.0 27980.0 ;
      RECT  70185.0 27840.0 70255.0 27980.0 ;
      RECT  70520.0 27840.0 70590.0 27980.0 ;
      RECT  70890.0 27840.0 70960.0 27980.0 ;
      RECT  71225.0 27840.0 71295.0 27980.0 ;
      RECT  71595.0 27840.0 71665.0 27980.0 ;
      RECT  71930.0 27840.0 72000.0 27980.0 ;
      RECT  72300.0 27840.0 72370.0 27980.0 ;
      RECT  72635.0 27840.0 72705.0 27980.0 ;
      RECT  73005.0 27840.0 73075.0 27980.0 ;
      RECT  73340.0 27840.0 73410.0 27980.0 ;
      RECT  73710.0 27840.0 73780.0 27980.0 ;
      RECT  74045.0 27840.0 74115.0 27980.0 ;
      RECT  74415.0 27840.0 74485.0 27980.0 ;
      RECT  74750.0 27840.0 74820.0 27980.0 ;
      RECT  75120.0 27840.0 75190.0 27980.0 ;
      RECT  75455.0 27840.0 75525.0 27980.0 ;
      RECT  75825.0 27840.0 75895.0 27980.0 ;
      RECT  76160.0 27840.0 76230.0 27980.0 ;
      RECT  76530.0 27840.0 76600.0 27980.0 ;
      RECT  76865.0 27840.0 76935.0 27980.0 ;
      RECT  77235.0 27840.0 77305.0 27980.0 ;
      RECT  77570.0 27840.0 77640.0 27980.0 ;
      RECT  77940.0 27840.0 78010.0 27980.0 ;
      RECT  78275.0 27840.0 78345.0 27980.0 ;
      RECT  78645.0 27840.0 78715.0 27980.0 ;
      RECT  78980.0 27840.0 79050.0 27980.0 ;
      RECT  79350.0 27840.0 79420.0 27980.0 ;
      RECT  79685.0 27840.0 79755.0 27980.0 ;
      RECT  80055.0 27840.0 80125.0 27980.0 ;
      RECT  80390.0 27840.0 80460.0 27980.0 ;
      RECT  80760.0 27840.0 80830.0 27980.0 ;
      RECT  81095.0 27840.0 81165.0 27980.0 ;
      RECT  81465.0 27840.0 81535.0 27980.0 ;
      RECT  81800.0 27840.0 81870.0 27980.0 ;
      RECT  82170.0 27840.0 82240.0 27980.0 ;
      RECT  82505.0 27840.0 82575.0 27980.0 ;
      RECT  82875.0 27840.0 82945.0 27980.0 ;
      RECT  83210.0 27840.0 83280.0 27980.0 ;
      RECT  83580.0 27840.0 83650.0 27980.0 ;
      RECT  83915.0 27840.0 83985.0 27980.0 ;
      RECT  84285.0 27840.0 84355.0 27980.0 ;
      RECT  84620.0 27840.0 84690.0 27980.0 ;
      RECT  84990.0 27840.0 85060.0 27980.0 ;
      RECT  85325.0 27840.0 85395.0 27980.0 ;
      RECT  85695.0 27840.0 85765.0 27980.0 ;
      RECT  86030.0 27840.0 86100.0 27980.0 ;
      RECT  86400.0 27840.0 86470.0 27980.0 ;
      RECT  86735.0 27840.0 86805.0 27980.0 ;
      RECT  87105.0 27840.0 87175.0 27980.0 ;
      RECT  87440.0 27840.0 87510.0 27980.0 ;
      RECT  87810.0 27840.0 87880.0 27980.0 ;
      RECT  88145.0 27840.0 88215.0 27980.0 ;
      RECT  88515.0 27840.0 88585.0 27980.0 ;
      RECT  88850.0 27840.0 88920.0 27980.0 ;
      RECT  89220.0 27840.0 89290.0 27980.0 ;
      RECT  89555.0 27840.0 89625.0 27980.0 ;
      RECT  89925.0 27840.0 89995.0 27980.0 ;
      RECT  90260.0 27840.0 90330.0 27980.0 ;
      RECT  90630.0 27840.0 90700.0 27980.0 ;
      RECT  90965.0 27840.0 91035.0 27980.0 ;
      RECT  91335.0 27840.0 91405.0 27980.0 ;
      RECT  91670.0 27840.0 91740.0 27980.0 ;
      RECT  92040.0 27840.0 92110.0 27980.0 ;
      RECT  92375.0 27840.0 92445.0 27980.0 ;
      RECT  92745.0 27840.0 92815.0 27980.0 ;
      RECT  93080.0 27840.0 93150.0 27980.0 ;
      RECT  93450.0 27840.0 93520.0 27980.0 ;
      RECT  93785.0 27840.0 93855.0 27980.0 ;
      RECT  94155.0 27840.0 94225.0 27980.0 ;
      RECT  94490.0 27840.0 94560.0 27980.0 ;
      RECT  94860.0 27840.0 94930.0 27980.0 ;
      RECT  95195.0 27840.0 95265.0 27980.0 ;
      RECT  95565.0 27840.0 95635.0 27980.0 ;
      RECT  95900.0 27840.0 95970.0 27980.0 ;
      RECT  96270.0 27840.0 96340.0 27980.0 ;
      RECT  96605.0 27840.0 96675.0 27980.0 ;
      RECT  96975.0 27840.0 97045.0 27980.0 ;
      RECT  97310.0 27840.0 97380.0 27980.0 ;
      RECT  97680.0 27840.0 97750.0 27980.0 ;
      RECT  98015.0 27840.0 98085.0 27980.0 ;
      RECT  98385.0 27840.0 98455.0 27980.0 ;
      RECT  98720.0 27840.0 98790.0 27980.0 ;
      RECT  99090.0 27840.0 99160.0 27980.0 ;
      RECT  99425.0 27840.0 99495.0 27980.0 ;
      RECT  99795.0 27840.0 99865.0 27980.0 ;
      RECT  100130.0 27840.0 100200.0 27980.0 ;
      RECT  100500.0 27840.0 100570.0 27980.0 ;
      RECT  100835.0 27840.0 100905.0 27980.0 ;
      RECT  101205.0 27840.0 101275.0 27980.0 ;
      RECT  101540.0 27840.0 101610.0 27980.0 ;
      RECT  101910.0 27840.0 101980.0 27980.0 ;
      RECT  102245.0 27840.0 102315.0 27980.0 ;
      RECT  102615.0 27840.0 102685.0 27980.0 ;
      RECT  102950.0 27840.0 103020.0 27980.0 ;
      RECT  103320.0 27840.0 103390.0 27980.0 ;
      RECT  103655.0 27840.0 103725.0 27980.0 ;
      RECT  104025.0 27840.0 104095.0 27980.0 ;
      RECT  104360.0 27840.0 104430.0 27980.0 ;
      RECT  104730.0 27840.0 104800.0 27980.0 ;
      RECT  105065.0 27840.0 105135.0 27980.0 ;
      RECT  105435.0 27840.0 105505.0 27980.0 ;
      RECT  105770.0 27840.0 105840.0 27980.0 ;
      RECT  15900.0 25170.0 15970.0 26150.0 ;
      RECT  16235.0 25170.0 16305.0 26150.0 ;
      RECT  18720.0 25170.0 18790.0 26150.0 ;
      RECT  19055.0 25170.0 19125.0 26150.0 ;
      RECT  21540.0 25170.0 21610.0 26150.0 ;
      RECT  21875.0 25170.0 21945.0 26150.0 ;
      RECT  24360.0 25170.0 24430.0 26150.0 ;
      RECT  24695.0 25170.0 24765.0 26150.0 ;
      RECT  27180.0 25170.0 27250.0 26150.0 ;
      RECT  27515.0 25170.0 27585.0 26150.0 ;
      RECT  30000.0 25170.0 30070.0 26150.0 ;
      RECT  30335.0 25170.0 30405.0 26150.0 ;
      RECT  32820.0 25170.0 32890.0 26150.0 ;
      RECT  33155.0 25170.0 33225.0 26150.0 ;
      RECT  35640.0 25170.0 35710.0 26150.0 ;
      RECT  35975.0 25170.0 36045.0 26150.0 ;
      RECT  38460.0 25170.0 38530.0 26150.0 ;
      RECT  38795.0 25170.0 38865.0 26150.0 ;
      RECT  41280.0 25170.0 41350.0 26150.0 ;
      RECT  41615.0 25170.0 41685.0 26150.0 ;
      RECT  44100.0 25170.0 44170.0 26150.0 ;
      RECT  44435.0 25170.0 44505.0 26150.0 ;
      RECT  46920.0 25170.0 46990.0 26150.0 ;
      RECT  47255.0 25170.0 47325.0 26150.0 ;
      RECT  49740.0 25170.0 49810.0 26150.0 ;
      RECT  50075.0 25170.0 50145.0 26150.0 ;
      RECT  52560.0 25170.0 52630.0 26150.0 ;
      RECT  52895.0 25170.0 52965.0 26150.0 ;
      RECT  55380.0 25170.0 55450.0 26150.0 ;
      RECT  55715.0 25170.0 55785.0 26150.0 ;
      RECT  58200.0 25170.0 58270.0 26150.0 ;
      RECT  58535.0 25170.0 58605.0 26150.0 ;
      RECT  61020.0 25170.0 61090.0 26150.0 ;
      RECT  61355.0 25170.0 61425.0 26150.0 ;
      RECT  63840.0 25170.0 63910.0 26150.0 ;
      RECT  64175.0 25170.0 64245.0 26150.0 ;
      RECT  66660.0 25170.0 66730.0 26150.0 ;
      RECT  66995.0 25170.0 67065.0 26150.0 ;
      RECT  69480.0 25170.0 69550.0 26150.0 ;
      RECT  69815.0 25170.0 69885.0 26150.0 ;
      RECT  72300.0 25170.0 72370.0 26150.0 ;
      RECT  72635.0 25170.0 72705.0 26150.0 ;
      RECT  75120.0 25170.0 75190.0 26150.0 ;
      RECT  75455.0 25170.0 75525.0 26150.0 ;
      RECT  77940.0 25170.0 78010.0 26150.0 ;
      RECT  78275.0 25170.0 78345.0 26150.0 ;
      RECT  80760.0 25170.0 80830.0 26150.0 ;
      RECT  81095.0 25170.0 81165.0 26150.0 ;
      RECT  83580.0 25170.0 83650.0 26150.0 ;
      RECT  83915.0 25170.0 83985.0 26150.0 ;
      RECT  86400.0 25170.0 86470.0 26150.0 ;
      RECT  86735.0 25170.0 86805.0 26150.0 ;
      RECT  89220.0 25170.0 89290.0 26150.0 ;
      RECT  89555.0 25170.0 89625.0 26150.0 ;
      RECT  92040.0 25170.0 92110.0 26150.0 ;
      RECT  92375.0 25170.0 92445.0 26150.0 ;
      RECT  94860.0 25170.0 94930.0 26150.0 ;
      RECT  95195.0 25170.0 95265.0 26150.0 ;
      RECT  97680.0 25170.0 97750.0 26150.0 ;
      RECT  98015.0 25170.0 98085.0 26150.0 ;
      RECT  100500.0 25170.0 100570.0 26150.0 ;
      RECT  100835.0 25170.0 100905.0 26150.0 ;
      RECT  103320.0 25170.0 103390.0 26150.0 ;
      RECT  103655.0 25170.0 103725.0 26150.0 ;
      RECT  15715.0 25170.0 15785.0 27980.0 ;
      RECT  16420.0 25170.0 16490.0 27980.0 ;
      RECT  17125.0 25170.0 17195.0 27980.0 ;
      RECT  17830.0 25170.0 17900.0 27980.0 ;
      RECT  18535.0 25170.0 18605.0 27980.0 ;
      RECT  19240.0 25170.0 19310.0 27980.0 ;
      RECT  19945.0 25170.0 20015.0 27980.0 ;
      RECT  20650.0 25170.0 20720.0 27980.0 ;
      RECT  21355.0 25170.0 21425.0 27980.0 ;
      RECT  22060.0 25170.0 22130.0 27980.0 ;
      RECT  22765.0 25170.0 22835.0 27980.0 ;
      RECT  23470.0 25170.0 23540.0 27980.0 ;
      RECT  24175.0 25170.0 24245.0 27980.0 ;
      RECT  24880.0 25170.0 24950.0 27980.0 ;
      RECT  25585.0 25170.0 25655.0 27980.0 ;
      RECT  26290.0 25170.0 26360.0 27980.0 ;
      RECT  26995.0 25170.0 27065.0 27980.0 ;
      RECT  27700.0 25170.0 27770.0 27980.0 ;
      RECT  28405.0 25170.0 28475.0 27980.0 ;
      RECT  29110.0 25170.0 29180.0 27980.0 ;
      RECT  29815.0 25170.0 29885.0 27980.0 ;
      RECT  30520.0 25170.0 30590.0 27980.0 ;
      RECT  31225.0 25170.0 31295.0 27980.0 ;
      RECT  31930.0 25170.0 32000.0 27980.0 ;
      RECT  32635.0 25170.0 32705.0 27980.0 ;
      RECT  33340.0 25170.0 33410.0 27980.0 ;
      RECT  34045.0 25170.0 34115.0 27980.0 ;
      RECT  34750.0 25170.0 34820.0 27980.0 ;
      RECT  35455.0 25170.0 35525.0 27980.0 ;
      RECT  36160.0 25170.0 36230.0 27980.0 ;
      RECT  36865.0 25170.0 36935.0 27980.0 ;
      RECT  37570.0 25170.0 37640.0 27980.0 ;
      RECT  38275.0 25170.0 38345.0 27980.0 ;
      RECT  38980.0 25170.0 39050.0 27980.0 ;
      RECT  39685.0 25170.0 39755.0 27980.0 ;
      RECT  40390.0 25170.0 40460.0 27980.0 ;
      RECT  41095.0 25170.0 41165.0 27980.0 ;
      RECT  41800.0 25170.0 41870.0 27980.0 ;
      RECT  42505.0 25170.0 42575.0 27980.0 ;
      RECT  43210.0 25170.0 43280.0 27980.0 ;
      RECT  43915.0 25170.0 43985.0 27980.0 ;
      RECT  44620.0 25170.0 44690.0 27980.0 ;
      RECT  45325.0 25170.0 45395.0 27980.0 ;
      RECT  46030.0 25170.0 46100.0 27980.0 ;
      RECT  46735.0 25170.0 46805.0 27980.0 ;
      RECT  47440.0 25170.0 47510.0 27980.0 ;
      RECT  48145.0 25170.0 48215.0 27980.0 ;
      RECT  48850.0 25170.0 48920.0 27980.0 ;
      RECT  49555.0 25170.0 49625.0 27980.0 ;
      RECT  50260.0 25170.0 50330.0 27980.0 ;
      RECT  50965.0 25170.0 51035.0 27980.0 ;
      RECT  51670.0 25170.0 51740.0 27980.0 ;
      RECT  52375.0 25170.0 52445.0 27980.0 ;
      RECT  53080.0 25170.0 53150.0 27980.0 ;
      RECT  53785.0 25170.0 53855.0 27980.0 ;
      RECT  54490.0 25170.0 54560.0 27980.0 ;
      RECT  55195.0 25170.0 55265.0 27980.0 ;
      RECT  55900.0 25170.0 55970.0 27980.0 ;
      RECT  56605.0 25170.0 56675.0 27980.0 ;
      RECT  57310.0 25170.0 57380.0 27980.0 ;
      RECT  58015.0 25170.0 58085.0 27980.0 ;
      RECT  58720.0 25170.0 58790.0 27980.0 ;
      RECT  59425.0 25170.0 59495.0 27980.0 ;
      RECT  60130.0 25170.0 60200.0 27980.0 ;
      RECT  60835.0 25170.0 60905.0 27980.0 ;
      RECT  61540.0 25170.0 61610.0 27980.0 ;
      RECT  62245.0 25170.0 62315.0 27980.0 ;
      RECT  62950.0 25170.0 63020.0 27980.0 ;
      RECT  63655.0 25170.0 63725.0 27980.0 ;
      RECT  64360.0 25170.0 64430.0 27980.0 ;
      RECT  65065.0 25170.0 65135.0 27980.0 ;
      RECT  65770.0 25170.0 65840.0 27980.0 ;
      RECT  66475.0 25170.0 66545.0 27980.0 ;
      RECT  67180.0 25170.0 67250.0 27980.0 ;
      RECT  67885.0 25170.0 67955.0 27980.0 ;
      RECT  68590.0 25170.0 68660.0 27980.0 ;
      RECT  69295.0 25170.0 69365.0 27980.0 ;
      RECT  70000.0 25170.0 70070.0 27980.0 ;
      RECT  70705.0 25170.0 70775.0 27980.0 ;
      RECT  71410.0 25170.0 71480.0 27980.0 ;
      RECT  72115.0 25170.0 72185.0 27980.0 ;
      RECT  72820.0 25170.0 72890.0 27980.0 ;
      RECT  73525.0 25170.0 73595.0 27980.0 ;
      RECT  74230.0 25170.0 74300.0 27980.0 ;
      RECT  74935.0 25170.0 75005.0 27980.0 ;
      RECT  75640.0 25170.0 75710.0 27980.0 ;
      RECT  76345.0 25170.0 76415.0 27980.0 ;
      RECT  77050.0 25170.0 77120.0 27980.0 ;
      RECT  77755.0 25170.0 77825.0 27980.0 ;
      RECT  78460.0 25170.0 78530.0 27980.0 ;
      RECT  79165.0 25170.0 79235.0 27980.0 ;
      RECT  79870.0 25170.0 79940.0 27980.0 ;
      RECT  80575.0 25170.0 80645.0 27980.0 ;
      RECT  81280.0 25170.0 81350.0 27980.0 ;
      RECT  81985.0 25170.0 82055.0 27980.0 ;
      RECT  82690.0 25170.0 82760.0 27980.0 ;
      RECT  83395.0 25170.0 83465.0 27980.0 ;
      RECT  84100.0 25170.0 84170.0 27980.0 ;
      RECT  84805.0 25170.0 84875.0 27980.0 ;
      RECT  85510.0 25170.0 85580.0 27980.0 ;
      RECT  86215.0 25170.0 86285.0 27980.0 ;
      RECT  86920.0 25170.0 86990.0 27980.0 ;
      RECT  87625.0 25170.0 87695.0 27980.0 ;
      RECT  88330.0 25170.0 88400.0 27980.0 ;
      RECT  89035.0 25170.0 89105.0 27980.0 ;
      RECT  89740.0 25170.0 89810.0 27980.0 ;
      RECT  90445.0 25170.0 90515.0 27980.0 ;
      RECT  91150.0 25170.0 91220.0 27980.0 ;
      RECT  91855.0 25170.0 91925.0 27980.0 ;
      RECT  92560.0 25170.0 92630.0 27980.0 ;
      RECT  93265.0 25170.0 93335.0 27980.0 ;
      RECT  93970.0 25170.0 94040.0 27980.0 ;
      RECT  94675.0 25170.0 94745.0 27980.0 ;
      RECT  95380.0 25170.0 95450.0 27980.0 ;
      RECT  96085.0 25170.0 96155.0 27980.0 ;
      RECT  96790.0 25170.0 96860.0 27980.0 ;
      RECT  97495.0 25170.0 97565.0 27980.0 ;
      RECT  98200.0 25170.0 98270.0 27980.0 ;
      RECT  98905.0 25170.0 98975.0 27980.0 ;
      RECT  99610.0 25170.0 99680.0 27980.0 ;
      RECT  100315.0 25170.0 100385.0 27980.0 ;
      RECT  101020.0 25170.0 101090.0 27980.0 ;
      RECT  101725.0 25170.0 101795.0 27980.0 ;
      RECT  102430.0 25170.0 102500.0 27980.0 ;
      RECT  103135.0 25170.0 103205.0 27980.0 ;
      RECT  103840.0 25170.0 103910.0 27980.0 ;
      RECT  104545.0 25170.0 104615.0 27980.0 ;
      RECT  105250.0 25170.0 105320.0 27980.0 ;
      RECT  8655.0 35.0 8725.0 5275.0 ;
      RECT  8930.0 35.0 9000.0 5275.0 ;
      RECT  8105.0 35.0 8175.0 5275.0 ;
      RECT  8380.0 35.0 8450.0 5275.0 ;
      RECT  9460.0 640.0 9530.0 710.0 ;
      RECT  9650.0 640.0 9720.0 710.0 ;
      RECT  9460.0 675.0 9530.0 1037.5 ;
      RECT  9495.0 640.0 9685.0 710.0 ;
      RECT  9650.0 332.5 9720.0 675.0 ;
      RECT  9460.0 1037.5 9530.0 1172.5 ;
      RECT  9650.0 197.5 9720.0 332.5 ;
      RECT  9752.5 640.0 9617.5 710.0 ;
      RECT  9460.0 2120.0 9530.0 2050.0 ;
      RECT  9650.0 2120.0 9720.0 2050.0 ;
      RECT  9460.0 2085.0 9530.0 1722.5 ;
      RECT  9495.0 2120.0 9685.0 2050.0 ;
      RECT  9650.0 2427.5 9720.0 2085.0 ;
      RECT  9460.0 1722.5 9530.0 1587.5 ;
      RECT  9650.0 2562.5 9720.0 2427.5 ;
      RECT  9752.5 2120.0 9617.5 2050.0 ;
      RECT  9460.0 3330.0 9530.0 3400.0 ;
      RECT  9650.0 3330.0 9720.0 3400.0 ;
      RECT  9460.0 3365.0 9530.0 3727.5 ;
      RECT  9495.0 3330.0 9685.0 3400.0 ;
      RECT  9650.0 3022.5 9720.0 3365.0 ;
      RECT  9460.0 3727.5 9530.0 3862.5 ;
      RECT  9650.0 2887.5 9720.0 3022.5 ;
      RECT  9752.5 3330.0 9617.5 3400.0 ;
      RECT  9460.0 4810.0 9530.0 4740.0 ;
      RECT  9650.0 4810.0 9720.0 4740.0 ;
      RECT  9460.0 4775.0 9530.0 4412.5 ;
      RECT  9495.0 4810.0 9685.0 4740.0 ;
      RECT  9650.0 5117.5 9720.0 4775.0 ;
      RECT  9460.0 4412.5 9530.0 4277.5 ;
      RECT  9650.0 5252.5 9720.0 5117.5 ;
      RECT  9752.5 4810.0 9617.5 4740.0 ;
      RECT  8207.5 1150.0 8072.5 1220.0 ;
      RECT  6822.5 627.5 6687.5 697.5 ;
      RECT  8482.5 2495.0 8347.5 2565.0 ;
      RECT  7097.5 2062.5 6962.5 2132.5 ;
      RECT  6822.5 2825.0 6687.5 2895.0 ;
      RECT  8757.5 2825.0 8622.5 2895.0 ;
      RECT  7097.5 4170.0 6962.5 4240.0 ;
      RECT  9032.5 4170.0 8897.5 4240.0 ;
      RECT  8207.5 640.0 8072.5 710.0 ;
      RECT  8482.5 425.0 8347.5 495.0 ;
      RECT  8757.5 2050.0 8622.5 2120.0 ;
      RECT  8482.5 2265.0 8347.5 2335.0 ;
      RECT  8207.5 3330.0 8072.5 3400.0 ;
      RECT  9032.5 3115.0 8897.5 3185.0 ;
      RECT  8757.5 4740.0 8622.5 4810.0 ;
      RECT  9032.5 4955.0 8897.5 5025.0 ;
      RECT  6720.0 35.0 6790.0 5275.0 ;
      RECT  6995.0 35.0 7065.0 5275.0 ;
      RECT  15750.0 20285.0 16455.0 25170.0 ;
      RECT  18570.0 20285.0 19275.0 25170.0 ;
      RECT  21390.0 20285.0 22095.0 25170.0 ;
      RECT  24210.0 20285.0 24915.0 25170.0 ;
      RECT  27030.0 20285.0 27735.0 25170.0 ;
      RECT  29850.0 20285.0 30555.0 25170.0 ;
      RECT  32670.0 20285.0 33375.0 25170.0 ;
      RECT  35490.0 20285.0 36195.0 25170.0 ;
      RECT  38310.0 20285.0 39015.0 25170.0 ;
      RECT  41130.0 20285.0 41835.0 25170.0 ;
      RECT  43950.0 20285.0 44655.0 25170.0 ;
      RECT  46770.0 20285.0 47475.0 25170.0 ;
      RECT  49590.0 20285.0 50295.0 25170.0 ;
      RECT  52410.0 20285.0 53115.0 25170.0 ;
      RECT  55230.0 20285.0 55935.0 25170.0 ;
      RECT  58050.0 20285.0 58755.0 25170.0 ;
      RECT  60870.0 20285.0 61575.0 25170.0 ;
      RECT  63690.0 20285.0 64395.0 25170.0 ;
      RECT  66510.0 20285.0 67215.0 25170.0 ;
      RECT  69330.0 20285.0 70035.0 25170.0 ;
      RECT  72150.0 20285.0 72855.0 25170.0 ;
      RECT  74970.0 20285.0 75675.0 25170.0 ;
      RECT  77790.0 20285.0 78495.0 25170.0 ;
      RECT  80610.0 20285.0 81315.0 25170.0 ;
      RECT  83430.0 20285.0 84135.0 25170.0 ;
      RECT  86250.0 20285.0 86955.0 25170.0 ;
      RECT  89070.0 20285.0 89775.0 25170.0 ;
      RECT  91890.0 20285.0 92595.0 25170.0 ;
      RECT  94710.0 20285.0 95415.0 25170.0 ;
      RECT  97530.0 20285.0 98235.0 25170.0 ;
      RECT  100350.0 20285.0 101055.0 25170.0 ;
      RECT  103170.0 20285.0 103875.0 25170.0 ;
      RECT  15900.0 20285.0 15970.0 25170.0 ;
      RECT  16235.0 20285.0 16305.0 24370.0 ;
      RECT  18720.0 20285.0 18790.0 25170.0 ;
      RECT  19055.0 20285.0 19125.0 24370.0 ;
      RECT  21540.0 20285.0 21610.0 25170.0 ;
      RECT  21875.0 20285.0 21945.0 24370.0 ;
      RECT  24360.0 20285.0 24430.0 25170.0 ;
      RECT  24695.0 20285.0 24765.0 24370.0 ;
      RECT  27180.0 20285.0 27250.0 25170.0 ;
      RECT  27515.0 20285.0 27585.0 24370.0 ;
      RECT  30000.0 20285.0 30070.0 25170.0 ;
      RECT  30335.0 20285.0 30405.0 24370.0 ;
      RECT  32820.0 20285.0 32890.0 25170.0 ;
      RECT  33155.0 20285.0 33225.0 24370.0 ;
      RECT  35640.0 20285.0 35710.0 25170.0 ;
      RECT  35975.0 20285.0 36045.0 24370.0 ;
      RECT  38460.0 20285.0 38530.0 25170.0 ;
      RECT  38795.0 20285.0 38865.0 24370.0 ;
      RECT  41280.0 20285.0 41350.0 25170.0 ;
      RECT  41615.0 20285.0 41685.0 24370.0 ;
      RECT  44100.0 20285.0 44170.0 25170.0 ;
      RECT  44435.0 20285.0 44505.0 24370.0 ;
      RECT  46920.0 20285.0 46990.0 25170.0 ;
      RECT  47255.0 20285.0 47325.0 24370.0 ;
      RECT  49740.0 20285.0 49810.0 25170.0 ;
      RECT  50075.0 20285.0 50145.0 24370.0 ;
      RECT  52560.0 20285.0 52630.0 25170.0 ;
      RECT  52895.0 20285.0 52965.0 24370.0 ;
      RECT  55380.0 20285.0 55450.0 25170.0 ;
      RECT  55715.0 20285.0 55785.0 24370.0 ;
      RECT  58200.0 20285.0 58270.0 25170.0 ;
      RECT  58535.0 20285.0 58605.0 24370.0 ;
      RECT  61020.0 20285.0 61090.0 25170.0 ;
      RECT  61355.0 20285.0 61425.0 24370.0 ;
      RECT  63840.0 20285.0 63910.0 25170.0 ;
      RECT  64175.0 20285.0 64245.0 24370.0 ;
      RECT  66660.0 20285.0 66730.0 25170.0 ;
      RECT  66995.0 20285.0 67065.0 24370.0 ;
      RECT  69480.0 20285.0 69550.0 25170.0 ;
      RECT  69815.0 20285.0 69885.0 24370.0 ;
      RECT  72300.0 20285.0 72370.0 25170.0 ;
      RECT  72635.0 20285.0 72705.0 24370.0 ;
      RECT  75120.0 20285.0 75190.0 25170.0 ;
      RECT  75455.0 20285.0 75525.0 24370.0 ;
      RECT  77940.0 20285.0 78010.0 25170.0 ;
      RECT  78275.0 20285.0 78345.0 24370.0 ;
      RECT  80760.0 20285.0 80830.0 25170.0 ;
      RECT  81095.0 20285.0 81165.0 24370.0 ;
      RECT  83580.0 20285.0 83650.0 25170.0 ;
      RECT  83915.0 20285.0 83985.0 24370.0 ;
      RECT  86400.0 20285.0 86470.0 25170.0 ;
      RECT  86735.0 20285.0 86805.0 24370.0 ;
      RECT  89220.0 20285.0 89290.0 25170.0 ;
      RECT  89555.0 20285.0 89625.0 24370.0 ;
      RECT  92040.0 20285.0 92110.0 25170.0 ;
      RECT  92375.0 20285.0 92445.0 24370.0 ;
      RECT  94860.0 20285.0 94930.0 25170.0 ;
      RECT  95195.0 20285.0 95265.0 24370.0 ;
      RECT  97680.0 20285.0 97750.0 25170.0 ;
      RECT  98015.0 20285.0 98085.0 24370.0 ;
      RECT  100500.0 20285.0 100570.0 25170.0 ;
      RECT  100835.0 20285.0 100905.0 24370.0 ;
      RECT  103320.0 20285.0 103390.0 25170.0 ;
      RECT  103655.0 20285.0 103725.0 24370.0 ;
      RECT  15750.0 16110.0 16455.0 20285.0 ;
      RECT  18570.0 16110.0 19275.0 20285.0 ;
      RECT  21390.0 16110.0 22095.0 20285.0 ;
      RECT  24210.0 16110.0 24915.0 20285.0 ;
      RECT  27030.0 16110.0 27735.0 20285.0 ;
      RECT  29850.0 16110.0 30555.0 20285.0 ;
      RECT  32670.0 16110.0 33375.0 20285.0 ;
      RECT  35490.0 16110.0 36195.0 20285.0 ;
      RECT  38310.0 16110.0 39015.0 20285.0 ;
      RECT  41130.0 16110.0 41835.0 20285.0 ;
      RECT  43950.0 16110.0 44655.0 20285.0 ;
      RECT  46770.0 16110.0 47475.0 20285.0 ;
      RECT  49590.0 16110.0 50295.0 20285.0 ;
      RECT  52410.0 16110.0 53115.0 20285.0 ;
      RECT  55230.0 16110.0 55935.0 20285.0 ;
      RECT  58050.0 16110.0 58755.0 20285.0 ;
      RECT  60870.0 16110.0 61575.0 20285.0 ;
      RECT  63690.0 16110.0 64395.0 20285.0 ;
      RECT  66510.0 16110.0 67215.0 20285.0 ;
      RECT  69330.0 16110.0 70035.0 20285.0 ;
      RECT  72150.0 16110.0 72855.0 20285.0 ;
      RECT  74970.0 16110.0 75675.0 20285.0 ;
      RECT  77790.0 16110.0 78495.0 20285.0 ;
      RECT  80610.0 16110.0 81315.0 20285.0 ;
      RECT  83430.0 16110.0 84135.0 20285.0 ;
      RECT  86250.0 16110.0 86955.0 20285.0 ;
      RECT  89070.0 16110.0 89775.0 20285.0 ;
      RECT  91890.0 16110.0 92595.0 20285.0 ;
      RECT  94710.0 16110.0 95415.0 20285.0 ;
      RECT  97530.0 16110.0 98235.0 20285.0 ;
      RECT  100350.0 16110.0 101055.0 20285.0 ;
      RECT  103170.0 16110.0 103875.0 20285.0 ;
      RECT  16067.5 16110.0 16137.5 16250.0 ;
      RECT  18887.5 16110.0 18957.5 16250.0 ;
      RECT  21707.5 16110.0 21777.5 16250.0 ;
      RECT  24527.5 16110.0 24597.5 16250.0 ;
      RECT  27347.5 16110.0 27417.5 16250.0 ;
      RECT  30167.5 16110.0 30237.5 16250.0 ;
      RECT  32987.5 16110.0 33057.5 16250.0 ;
      RECT  35807.5 16110.0 35877.5 16250.0 ;
      RECT  38627.5 16110.0 38697.5 16250.0 ;
      RECT  41447.5 16110.0 41517.5 16250.0 ;
      RECT  44267.5 16110.0 44337.5 16250.0 ;
      RECT  47087.5 16110.0 47157.5 16250.0 ;
      RECT  49907.5 16110.0 49977.5 16250.0 ;
      RECT  52727.5 16110.0 52797.5 16250.0 ;
      RECT  55547.5 16110.0 55617.5 16250.0 ;
      RECT  58367.5 16110.0 58437.5 16250.0 ;
      RECT  61187.5 16110.0 61257.5 16250.0 ;
      RECT  64007.5 16110.0 64077.5 16250.0 ;
      RECT  66827.5 16110.0 66897.5 16250.0 ;
      RECT  69647.5 16110.0 69717.5 16250.0 ;
      RECT  72467.5 16110.0 72537.5 16250.0 ;
      RECT  75287.5 16110.0 75357.5 16250.0 ;
      RECT  78107.5 16110.0 78177.5 16250.0 ;
      RECT  80927.5 16110.0 80997.5 16250.0 ;
      RECT  83747.5 16110.0 83817.5 16250.0 ;
      RECT  86567.5 16110.0 86637.5 16250.0 ;
      RECT  89387.5 16110.0 89457.5 16250.0 ;
      RECT  92207.5 16110.0 92277.5 16250.0 ;
      RECT  95027.5 16110.0 95097.5 16250.0 ;
      RECT  97847.5 16110.0 97917.5 16250.0 ;
      RECT  100667.5 16110.0 100737.5 16250.0 ;
      RECT  103487.5 16110.0 103557.5 16250.0 ;
      RECT  15900.0 19985.0 15970.0 20285.0 ;
      RECT  16235.0 17845.0 16305.0 20285.0 ;
      RECT  18720.0 19985.0 18790.0 20285.0 ;
      RECT  19055.0 17845.0 19125.0 20285.0 ;
      RECT  21540.0 19985.0 21610.0 20285.0 ;
      RECT  21875.0 17845.0 21945.0 20285.0 ;
      RECT  24360.0 19985.0 24430.0 20285.0 ;
      RECT  24695.0 17845.0 24765.0 20285.0 ;
      RECT  27180.0 19985.0 27250.0 20285.0 ;
      RECT  27515.0 17845.0 27585.0 20285.0 ;
      RECT  30000.0 19985.0 30070.0 20285.0 ;
      RECT  30335.0 17845.0 30405.0 20285.0 ;
      RECT  32820.0 19985.0 32890.0 20285.0 ;
      RECT  33155.0 17845.0 33225.0 20285.0 ;
      RECT  35640.0 19985.0 35710.0 20285.0 ;
      RECT  35975.0 17845.0 36045.0 20285.0 ;
      RECT  38460.0 19985.0 38530.0 20285.0 ;
      RECT  38795.0 17845.0 38865.0 20285.0 ;
      RECT  41280.0 19985.0 41350.0 20285.0 ;
      RECT  41615.0 17845.0 41685.0 20285.0 ;
      RECT  44100.0 19985.0 44170.0 20285.0 ;
      RECT  44435.0 17845.0 44505.0 20285.0 ;
      RECT  46920.0 19985.0 46990.0 20285.0 ;
      RECT  47255.0 17845.0 47325.0 20285.0 ;
      RECT  49740.0 19985.0 49810.0 20285.0 ;
      RECT  50075.0 17845.0 50145.0 20285.0 ;
      RECT  52560.0 19985.0 52630.0 20285.0 ;
      RECT  52895.0 17845.0 52965.0 20285.0 ;
      RECT  55380.0 19985.0 55450.0 20285.0 ;
      RECT  55715.0 17845.0 55785.0 20285.0 ;
      RECT  58200.0 19985.0 58270.0 20285.0 ;
      RECT  58535.0 17845.0 58605.0 20285.0 ;
      RECT  61020.0 19985.0 61090.0 20285.0 ;
      RECT  61355.0 17845.0 61425.0 20285.0 ;
      RECT  63840.0 19985.0 63910.0 20285.0 ;
      RECT  64175.0 17845.0 64245.0 20285.0 ;
      RECT  66660.0 19985.0 66730.0 20285.0 ;
      RECT  66995.0 17845.0 67065.0 20285.0 ;
      RECT  69480.0 19985.0 69550.0 20285.0 ;
      RECT  69815.0 17845.0 69885.0 20285.0 ;
      RECT  72300.0 19985.0 72370.0 20285.0 ;
      RECT  72635.0 17845.0 72705.0 20285.0 ;
      RECT  75120.0 19985.0 75190.0 20285.0 ;
      RECT  75455.0 17845.0 75525.0 20285.0 ;
      RECT  77940.0 19985.0 78010.0 20285.0 ;
      RECT  78275.0 17845.0 78345.0 20285.0 ;
      RECT  80760.0 19985.0 80830.0 20285.0 ;
      RECT  81095.0 17845.0 81165.0 20285.0 ;
      RECT  83580.0 19985.0 83650.0 20285.0 ;
      RECT  83915.0 17845.0 83985.0 20285.0 ;
      RECT  86400.0 19985.0 86470.0 20285.0 ;
      RECT  86735.0 17845.0 86805.0 20285.0 ;
      RECT  89220.0 19985.0 89290.0 20285.0 ;
      RECT  89555.0 17845.0 89625.0 20285.0 ;
      RECT  92040.0 19985.0 92110.0 20285.0 ;
      RECT  92375.0 17845.0 92445.0 20285.0 ;
      RECT  94860.0 19985.0 94930.0 20285.0 ;
      RECT  95195.0 17845.0 95265.0 20285.0 ;
      RECT  97680.0 19985.0 97750.0 20285.0 ;
      RECT  98015.0 17845.0 98085.0 20285.0 ;
      RECT  100500.0 19985.0 100570.0 20285.0 ;
      RECT  100835.0 17845.0 100905.0 20285.0 ;
      RECT  103320.0 19985.0 103390.0 20285.0 ;
      RECT  103655.0 17845.0 103725.0 20285.0 ;
      RECT  15750.0 9670.0 16455.0 16110.0 ;
      RECT  18570.0 9670.0 19275.0 16110.0 ;
      RECT  21390.0 9670.0 22095.0 16110.0 ;
      RECT  24210.0 9670.0 24915.0 16110.0 ;
      RECT  27030.0 9670.0 27735.0 16110.0 ;
      RECT  29850.0 9670.0 30555.0 16110.0 ;
      RECT  32670.0 9670.0 33375.0 16110.0 ;
      RECT  35490.0 9670.0 36195.0 16110.0 ;
      RECT  38310.0 9670.0 39015.0 16110.0 ;
      RECT  41130.0 9670.0 41835.0 16110.0 ;
      RECT  43950.0 9670.0 44655.0 16110.0 ;
      RECT  46770.0 9670.0 47475.0 16110.0 ;
      RECT  49590.0 9670.0 50295.0 16110.0 ;
      RECT  52410.0 9670.0 53115.0 16110.0 ;
      RECT  55230.0 9670.0 55935.0 16110.0 ;
      RECT  58050.0 9670.0 58755.0 16110.0 ;
      RECT  60870.0 9670.0 61575.0 16110.0 ;
      RECT  63690.0 9670.0 64395.0 16110.0 ;
      RECT  66510.0 9670.0 67215.0 16110.0 ;
      RECT  69330.0 9670.0 70035.0 16110.0 ;
      RECT  72150.0 9670.0 72855.0 16110.0 ;
      RECT  74970.0 9670.0 75675.0 16110.0 ;
      RECT  77790.0 9670.0 78495.0 16110.0 ;
      RECT  80610.0 9670.0 81315.0 16110.0 ;
      RECT  83430.0 9670.0 84135.0 16110.0 ;
      RECT  86250.0 9670.0 86955.0 16110.0 ;
      RECT  89070.0 9670.0 89775.0 16110.0 ;
      RECT  91890.0 9670.0 92595.0 16110.0 ;
      RECT  94710.0 9670.0 95415.0 16110.0 ;
      RECT  97530.0 9670.0 98235.0 16110.0 ;
      RECT  100350.0 9670.0 101055.0 16110.0 ;
      RECT  103170.0 9670.0 103875.0 16110.0 ;
      RECT  16067.5 9670.0 16137.5 9815.0 ;
      RECT  18887.5 9670.0 18957.5 9815.0 ;
      RECT  21707.5 9670.0 21777.5 9815.0 ;
      RECT  24527.5 9670.0 24597.5 9815.0 ;
      RECT  27347.5 9670.0 27417.5 9815.0 ;
      RECT  30167.5 9670.0 30237.5 9815.0 ;
      RECT  32987.5 9670.0 33057.5 9815.0 ;
      RECT  35807.5 9670.0 35877.5 9815.0 ;
      RECT  38627.5 9670.0 38697.5 9815.0 ;
      RECT  41447.5 9670.0 41517.5 9815.0 ;
      RECT  44267.5 9670.0 44337.5 9815.0 ;
      RECT  47087.5 9670.0 47157.5 9815.0 ;
      RECT  49907.5 9670.0 49977.5 9815.0 ;
      RECT  52727.5 9670.0 52797.5 9815.0 ;
      RECT  55547.5 9670.0 55617.5 9815.0 ;
      RECT  58367.5 9670.0 58437.5 9815.0 ;
      RECT  61187.5 9670.0 61257.5 9815.0 ;
      RECT  64007.5 9670.0 64077.5 9815.0 ;
      RECT  66827.5 9670.0 66897.5 9815.0 ;
      RECT  69647.5 9670.0 69717.5 9815.0 ;
      RECT  72467.5 9670.0 72537.5 9815.0 ;
      RECT  75287.5 9670.0 75357.5 9815.0 ;
      RECT  78107.5 9670.0 78177.5 9815.0 ;
      RECT  80927.5 9670.0 80997.5 9815.0 ;
      RECT  83747.5 9670.0 83817.5 9815.0 ;
      RECT  86567.5 9670.0 86637.5 9815.0 ;
      RECT  89387.5 9670.0 89457.5 9815.0 ;
      RECT  92207.5 9670.0 92277.5 9815.0 ;
      RECT  95027.5 9670.0 95097.5 9815.0 ;
      RECT  97847.5 9670.0 97917.5 9815.0 ;
      RECT  100667.5 9670.0 100737.5 9815.0 ;
      RECT  103487.5 9670.0 103557.5 9815.0 ;
      RECT  16067.5 15840.0 16137.5 16110.0 ;
      RECT  15912.5 15422.5 15982.5 16110.0 ;
      RECT  18887.5 15840.0 18957.5 16110.0 ;
      RECT  18732.5 15422.5 18802.5 16110.0 ;
      RECT  21707.5 15840.0 21777.5 16110.0 ;
      RECT  21552.5 15422.5 21622.5 16110.0 ;
      RECT  24527.5 15840.0 24597.5 16110.0 ;
      RECT  24372.5 15422.5 24442.5 16110.0 ;
      RECT  27347.5 15840.0 27417.5 16110.0 ;
      RECT  27192.5 15422.5 27262.5 16110.0 ;
      RECT  30167.5 15840.0 30237.5 16110.0 ;
      RECT  30012.5 15422.5 30082.5 16110.0 ;
      RECT  32987.5 15840.0 33057.5 16110.0 ;
      RECT  32832.5 15422.5 32902.5 16110.0 ;
      RECT  35807.5 15840.0 35877.5 16110.0 ;
      RECT  35652.5 15422.5 35722.5 16110.0 ;
      RECT  38627.5 15840.0 38697.5 16110.0 ;
      RECT  38472.5 15422.5 38542.5 16110.0 ;
      RECT  41447.5 15840.0 41517.5 16110.0 ;
      RECT  41292.5 15422.5 41362.5 16110.0 ;
      RECT  44267.5 15840.0 44337.5 16110.0 ;
      RECT  44112.5 15422.5 44182.5 16110.0 ;
      RECT  47087.5 15840.0 47157.5 16110.0 ;
      RECT  46932.5 15422.5 47002.5 16110.0 ;
      RECT  49907.5 15840.0 49977.5 16110.0 ;
      RECT  49752.5 15422.5 49822.5 16110.0 ;
      RECT  52727.5 15840.0 52797.5 16110.0 ;
      RECT  52572.5 15422.5 52642.5 16110.0 ;
      RECT  55547.5 15840.0 55617.5 16110.0 ;
      RECT  55392.5 15422.5 55462.5 16110.0 ;
      RECT  58367.5 15840.0 58437.5 16110.0 ;
      RECT  58212.5 15422.5 58282.5 16110.0 ;
      RECT  61187.5 15840.0 61257.5 16110.0 ;
      RECT  61032.5 15422.5 61102.5 16110.0 ;
      RECT  64007.5 15840.0 64077.5 16110.0 ;
      RECT  63852.5 15422.5 63922.5 16110.0 ;
      RECT  66827.5 15840.0 66897.5 16110.0 ;
      RECT  66672.5 15422.5 66742.5 16110.0 ;
      RECT  69647.5 15840.0 69717.5 16110.0 ;
      RECT  69492.5 15422.5 69562.5 16110.0 ;
      RECT  72467.5 15840.0 72537.5 16110.0 ;
      RECT  72312.5 15422.5 72382.5 16110.0 ;
      RECT  75287.5 15840.0 75357.5 16110.0 ;
      RECT  75132.5 15422.5 75202.5 16110.0 ;
      RECT  78107.5 15840.0 78177.5 16110.0 ;
      RECT  77952.5 15422.5 78022.5 16110.0 ;
      RECT  80927.5 15840.0 80997.5 16110.0 ;
      RECT  80772.5 15422.5 80842.5 16110.0 ;
      RECT  83747.5 15840.0 83817.5 16110.0 ;
      RECT  83592.5 15422.5 83662.5 16110.0 ;
      RECT  86567.5 15840.0 86637.5 16110.0 ;
      RECT  86412.5 15422.5 86482.5 16110.0 ;
      RECT  89387.5 15840.0 89457.5 16110.0 ;
      RECT  89232.5 15422.5 89302.5 16110.0 ;
      RECT  92207.5 15840.0 92277.5 16110.0 ;
      RECT  92052.5 15422.5 92122.5 16110.0 ;
      RECT  95027.5 15840.0 95097.5 16110.0 ;
      RECT  94872.5 15422.5 94942.5 16110.0 ;
      RECT  97847.5 15840.0 97917.5 16110.0 ;
      RECT  97692.5 15422.5 97762.5 16110.0 ;
      RECT  100667.5 15840.0 100737.5 16110.0 ;
      RECT  100512.5 15422.5 100582.5 16110.0 ;
      RECT  103487.5 15840.0 103557.5 16110.0 ;
      RECT  103332.5 15422.5 103402.5 16110.0 ;
      RECT  15715.0 9670.0 15785.0 16110.0 ;
      RECT  16420.0 9670.0 16490.0 16110.0 ;
      RECT  18535.0 9670.0 18605.0 16110.0 ;
      RECT  19240.0 9670.0 19310.0 16110.0 ;
      RECT  21355.0 9670.0 21425.0 16110.0 ;
      RECT  22060.0 9670.0 22130.0 16110.0 ;
      RECT  24175.0 9670.0 24245.0 16110.0 ;
      RECT  24880.0 9670.0 24950.0 16110.0 ;
      RECT  26995.0 9670.0 27065.0 16110.0 ;
      RECT  27700.0 9670.0 27770.0 16110.0 ;
      RECT  29815.0 9670.0 29885.0 16110.0 ;
      RECT  30520.0 9670.0 30590.0 16110.0 ;
      RECT  32635.0 9670.0 32705.0 16110.0 ;
      RECT  33340.0 9670.0 33410.0 16110.0 ;
      RECT  35455.0 9670.0 35525.0 16110.0 ;
      RECT  36160.0 9670.0 36230.0 16110.0 ;
      RECT  38275.0 9670.0 38345.0 16110.0 ;
      RECT  38980.0 9670.0 39050.0 16110.0 ;
      RECT  41095.0 9670.0 41165.0 16110.0 ;
      RECT  41800.0 9670.0 41870.0 16110.0 ;
      RECT  43915.0 9670.0 43985.0 16110.0 ;
      RECT  44620.0 9670.0 44690.0 16110.0 ;
      RECT  46735.0 9670.0 46805.0 16110.0 ;
      RECT  47440.0 9670.0 47510.0 16110.0 ;
      RECT  49555.0 9670.0 49625.0 16110.0 ;
      RECT  50260.0 9670.0 50330.0 16110.0 ;
      RECT  52375.0 9670.0 52445.0 16110.0 ;
      RECT  53080.0 9670.0 53150.0 16110.0 ;
      RECT  55195.0 9670.0 55265.0 16110.0 ;
      RECT  55900.0 9670.0 55970.0 16110.0 ;
      RECT  58015.0 9670.0 58085.0 16110.0 ;
      RECT  58720.0 9670.0 58790.0 16110.0 ;
      RECT  60835.0 9670.0 60905.0 16110.0 ;
      RECT  61540.0 9670.0 61610.0 16110.0 ;
      RECT  63655.0 9670.0 63725.0 16110.0 ;
      RECT  64360.0 9670.0 64430.0 16110.0 ;
      RECT  66475.0 9670.0 66545.0 16110.0 ;
      RECT  67180.0 9670.0 67250.0 16110.0 ;
      RECT  69295.0 9670.0 69365.0 16110.0 ;
      RECT  70000.0 9670.0 70070.0 16110.0 ;
      RECT  72115.0 9670.0 72185.0 16110.0 ;
      RECT  72820.0 9670.0 72890.0 16110.0 ;
      RECT  74935.0 9670.0 75005.0 16110.0 ;
      RECT  75640.0 9670.0 75710.0 16110.0 ;
      RECT  77755.0 9670.0 77825.0 16110.0 ;
      RECT  78460.0 9670.0 78530.0 16110.0 ;
      RECT  80575.0 9670.0 80645.0 16110.0 ;
      RECT  81280.0 9670.0 81350.0 16110.0 ;
      RECT  83395.0 9670.0 83465.0 16110.0 ;
      RECT  84100.0 9670.0 84170.0 16110.0 ;
      RECT  86215.0 9670.0 86285.0 16110.0 ;
      RECT  86920.0 9670.0 86990.0 16110.0 ;
      RECT  89035.0 9670.0 89105.0 16110.0 ;
      RECT  89740.0 9670.0 89810.0 16110.0 ;
      RECT  91855.0 9670.0 91925.0 16110.0 ;
      RECT  92560.0 9670.0 92630.0 16110.0 ;
      RECT  94675.0 9670.0 94745.0 16110.0 ;
      RECT  95380.0 9670.0 95450.0 16110.0 ;
      RECT  97495.0 9670.0 97565.0 16110.0 ;
      RECT  98200.0 9670.0 98270.0 16110.0 ;
      RECT  100315.0 9670.0 100385.0 16110.0 ;
      RECT  101020.0 9670.0 101090.0 16110.0 ;
      RECT  103135.0 9670.0 103205.0 16110.0 ;
      RECT  103840.0 9670.0 103910.0 16110.0 ;
      RECT  15750.0 9670.0 16455.0 6695.0 ;
      RECT  18570.0 9670.0 19275.0 6695.0 ;
      RECT  21390.0 9670.0 22095.0 6695.0 ;
      RECT  24210.0 9670.0 24915.0 6695.0 ;
      RECT  27030.0 9670.0 27735.0 6695.0 ;
      RECT  29850.0 9670.0 30555.0 6695.0 ;
      RECT  32670.0 9670.0 33375.0 6695.0 ;
      RECT  35490.0 9670.0 36195.0 6695.0 ;
      RECT  38310.0 9670.0 39015.0 6695.0 ;
      RECT  41130.0 9670.0 41835.0 6695.0 ;
      RECT  43950.0 9670.0 44655.0 6695.0 ;
      RECT  46770.0 9670.0 47475.0 6695.0 ;
      RECT  49590.0 9670.0 50295.0 6695.0 ;
      RECT  52410.0 9670.0 53115.0 6695.0 ;
      RECT  55230.0 9670.0 55935.0 6695.0 ;
      RECT  58050.0 9670.0 58755.0 6695.0 ;
      RECT  60870.0 9670.0 61575.0 6695.0 ;
      RECT  63690.0 9670.0 64395.0 6695.0 ;
      RECT  66510.0 9670.0 67215.0 6695.0 ;
      RECT  69330.0 9670.0 70035.0 6695.0 ;
      RECT  72150.0 9670.0 72855.0 6695.0 ;
      RECT  74970.0 9670.0 75675.0 6695.0 ;
      RECT  77790.0 9670.0 78495.0 6695.0 ;
      RECT  80610.0 9670.0 81315.0 6695.0 ;
      RECT  83430.0 9670.0 84135.0 6695.0 ;
      RECT  86250.0 9670.0 86955.0 6695.0 ;
      RECT  89070.0 9670.0 89775.0 6695.0 ;
      RECT  91890.0 9670.0 92595.0 6695.0 ;
      RECT  94710.0 9670.0 95415.0 6695.0 ;
      RECT  97530.0 9670.0 98235.0 6695.0 ;
      RECT  100350.0 9670.0 101055.0 6695.0 ;
      RECT  103170.0 9670.0 103875.0 6695.0 ;
      RECT  16067.5 6935.0 16137.5 6695.0 ;
      RECT  18887.5 6935.0 18957.5 6695.0 ;
      RECT  21707.5 6935.0 21777.5 6695.0 ;
      RECT  24527.5 6935.0 24597.5 6695.0 ;
      RECT  27347.5 6935.0 27417.5 6695.0 ;
      RECT  30167.5 6935.0 30237.5 6695.0 ;
      RECT  32987.5 6935.0 33057.5 6695.0 ;
      RECT  35807.5 6935.0 35877.5 6695.0 ;
      RECT  38627.5 6935.0 38697.5 6695.0 ;
      RECT  41447.5 6935.0 41517.5 6695.0 ;
      RECT  44267.5 6935.0 44337.5 6695.0 ;
      RECT  47087.5 6935.0 47157.5 6695.0 ;
      RECT  49907.5 6935.0 49977.5 6695.0 ;
      RECT  52727.5 6935.0 52797.5 6695.0 ;
      RECT  55547.5 6935.0 55617.5 6695.0 ;
      RECT  58367.5 6935.0 58437.5 6695.0 ;
      RECT  61187.5 6935.0 61257.5 6695.0 ;
      RECT  64007.5 6935.0 64077.5 6695.0 ;
      RECT  66827.5 6935.0 66897.5 6695.0 ;
      RECT  69647.5 6935.0 69717.5 6695.0 ;
      RECT  72467.5 6935.0 72537.5 6695.0 ;
      RECT  75287.5 6935.0 75357.5 6695.0 ;
      RECT  78107.5 6935.0 78177.5 6695.0 ;
      RECT  80927.5 6935.0 80997.5 6695.0 ;
      RECT  83747.5 6935.0 83817.5 6695.0 ;
      RECT  86567.5 6935.0 86637.5 6695.0 ;
      RECT  89387.5 6935.0 89457.5 6695.0 ;
      RECT  92207.5 6935.0 92277.5 6695.0 ;
      RECT  95027.5 6935.0 95097.5 6695.0 ;
      RECT  97847.5 6935.0 97917.5 6695.0 ;
      RECT  100667.5 6935.0 100737.5 6695.0 ;
      RECT  103487.5 6935.0 103557.5 6695.0 ;
      RECT  16067.5 9670.0 16137.5 9320.0 ;
      RECT  18887.5 9670.0 18957.5 9320.0 ;
      RECT  21707.5 9670.0 21777.5 9320.0 ;
      RECT  24527.5 9670.0 24597.5 9320.0 ;
      RECT  27347.5 9670.0 27417.5 9320.0 ;
      RECT  30167.5 9670.0 30237.5 9320.0 ;
      RECT  32987.5 9670.0 33057.5 9320.0 ;
      RECT  35807.5 9670.0 35877.5 9320.0 ;
      RECT  38627.5 9670.0 38697.5 9320.0 ;
      RECT  41447.5 9670.0 41517.5 9320.0 ;
      RECT  44267.5 9670.0 44337.5 9320.0 ;
      RECT  47087.5 9670.0 47157.5 9320.0 ;
      RECT  49907.5 9670.0 49977.5 9320.0 ;
      RECT  52727.5 9670.0 52797.5 9320.0 ;
      RECT  55547.5 9670.0 55617.5 9320.0 ;
      RECT  58367.5 9670.0 58437.5 9320.0 ;
      RECT  61187.5 9670.0 61257.5 9320.0 ;
      RECT  64007.5 9670.0 64077.5 9320.0 ;
      RECT  66827.5 9670.0 66897.5 9320.0 ;
      RECT  69647.5 9670.0 69717.5 9320.0 ;
      RECT  72467.5 9670.0 72537.5 9320.0 ;
      RECT  75287.5 9670.0 75357.5 9320.0 ;
      RECT  78107.5 9670.0 78177.5 9320.0 ;
      RECT  80927.5 9670.0 80997.5 9320.0 ;
      RECT  83747.5 9670.0 83817.5 9320.0 ;
      RECT  86567.5 9670.0 86637.5 9320.0 ;
      RECT  89387.5 9670.0 89457.5 9320.0 ;
      RECT  92207.5 9670.0 92277.5 9320.0 ;
      RECT  95027.5 9670.0 95097.5 9320.0 ;
      RECT  97847.5 9670.0 97917.5 9320.0 ;
      RECT  100667.5 9670.0 100737.5 9320.0 ;
      RECT  103487.5 9670.0 103557.5 9320.0 ;
      RECT  5030.0 11875.0 5100.0 114095.0 ;
      RECT  5205.0 11875.0 5275.0 114095.0 ;
      RECT  5380.0 11875.0 5450.0 114095.0 ;
      RECT  5555.0 11875.0 5625.0 114095.0 ;
      RECT  5730.0 11875.0 5800.0 114095.0 ;
      RECT  5905.0 11875.0 5975.0 114095.0 ;
      RECT  6080.0 11875.0 6150.0 114095.0 ;
      RECT  6255.0 11875.0 6325.0 114095.0 ;
      RECT  6430.0 11875.0 6500.0 114095.0 ;
      RECT  6605.0 11875.0 6675.0 114095.0 ;
      RECT  6780.0 11875.0 6850.0 114095.0 ;
      RECT  6955.0 11875.0 7025.0 114095.0 ;
      RECT  9160.0 11875.0 9090.0 17115.0 ;
      RECT  8885.0 11875.0 8815.0 17115.0 ;
      RECT  9710.0 11875.0 9640.0 17115.0 ;
      RECT  9435.0 11875.0 9365.0 17115.0 ;
      RECT  8355.0 12480.0 8285.0 12550.0 ;
      RECT  8165.0 12480.0 8095.0 12550.0 ;
      RECT  8355.0 12515.0 8285.0 12877.5 ;
      RECT  8320.0 12480.0 8130.0 12550.0 ;
      RECT  8165.0 12172.5 8095.0 12515.0 ;
      RECT  8355.0 12877.5 8285.0 13012.5 ;
      RECT  8165.0 12037.5 8095.0 12172.5 ;
      RECT  8062.5 12480.0 8197.5 12550.0 ;
      RECT  8355.0 13960.0 8285.0 13890.0 ;
      RECT  8165.0 13960.0 8095.0 13890.0 ;
      RECT  8355.0 13925.0 8285.0 13562.5 ;
      RECT  8320.0 13960.0 8130.0 13890.0 ;
      RECT  8165.0 14267.5 8095.0 13925.0 ;
      RECT  8355.0 13562.5 8285.0 13427.5 ;
      RECT  8165.0 14402.5 8095.0 14267.5 ;
      RECT  8062.5 13960.0 8197.5 13890.0 ;
      RECT  8355.0 15170.0 8285.0 15240.0 ;
      RECT  8165.0 15170.0 8095.0 15240.0 ;
      RECT  8355.0 15205.0 8285.0 15567.5 ;
      RECT  8320.0 15170.0 8130.0 15240.0 ;
      RECT  8165.0 14862.5 8095.0 15205.0 ;
      RECT  8355.0 15567.5 8285.0 15702.5 ;
      RECT  8165.0 14727.5 8095.0 14862.5 ;
      RECT  8062.5 15170.0 8197.5 15240.0 ;
      RECT  8355.0 16650.0 8285.0 16580.0 ;
      RECT  8165.0 16650.0 8095.0 16580.0 ;
      RECT  8355.0 16615.0 8285.0 16252.5 ;
      RECT  8320.0 16650.0 8130.0 16580.0 ;
      RECT  8165.0 16957.5 8095.0 16615.0 ;
      RECT  8355.0 16252.5 8285.0 16117.5 ;
      RECT  8165.0 17092.5 8095.0 16957.5 ;
      RECT  8062.5 16650.0 8197.5 16580.0 ;
      RECT  9607.5 12990.0 9742.5 13060.0 ;
      RECT  10992.5 12467.5 11127.5 12537.5 ;
      RECT  9332.5 14335.0 9467.5 14405.0 ;
      RECT  10717.5 13902.5 10852.5 13972.5 ;
      RECT  10992.5 14665.0 11127.5 14735.0 ;
      RECT  9057.5 14665.0 9192.5 14735.0 ;
      RECT  10717.5 16010.0 10852.5 16080.0 ;
      RECT  8782.5 16010.0 8917.5 16080.0 ;
      RECT  9607.5 12480.0 9742.5 12550.0 ;
      RECT  9332.5 12265.0 9467.5 12335.0 ;
      RECT  9057.5 13890.0 9192.5 13960.0 ;
      RECT  9332.5 14105.0 9467.5 14175.0 ;
      RECT  9607.5 15170.0 9742.5 15240.0 ;
      RECT  8782.5 14955.0 8917.5 15025.0 ;
      RECT  9057.5 16580.0 9192.5 16650.0 ;
      RECT  8782.5 16795.0 8917.5 16865.0 ;
      RECT  11095.0 11875.0 11025.0 17115.0 ;
      RECT  10820.0 11875.0 10750.0 17115.0 ;
      RECT  9160.0 17255.0 9090.0 22495.0 ;
      RECT  8885.0 17255.0 8815.0 22495.0 ;
      RECT  9710.0 17255.0 9640.0 22495.0 ;
      RECT  9435.0 17255.0 9365.0 22495.0 ;
      RECT  8355.0 17860.0 8285.0 17930.0 ;
      RECT  8165.0 17860.0 8095.0 17930.0 ;
      RECT  8355.0 17895.0 8285.0 18257.5 ;
      RECT  8320.0 17860.0 8130.0 17930.0 ;
      RECT  8165.0 17552.5 8095.0 17895.0 ;
      RECT  8355.0 18257.5 8285.0 18392.5 ;
      RECT  8165.0 17417.5 8095.0 17552.5 ;
      RECT  8062.5 17860.0 8197.5 17930.0 ;
      RECT  8355.0 19340.0 8285.0 19270.0 ;
      RECT  8165.0 19340.0 8095.0 19270.0 ;
      RECT  8355.0 19305.0 8285.0 18942.5 ;
      RECT  8320.0 19340.0 8130.0 19270.0 ;
      RECT  8165.0 19647.5 8095.0 19305.0 ;
      RECT  8355.0 18942.5 8285.0 18807.5 ;
      RECT  8165.0 19782.5 8095.0 19647.5 ;
      RECT  8062.5 19340.0 8197.5 19270.0 ;
      RECT  8355.0 20550.0 8285.0 20620.0 ;
      RECT  8165.0 20550.0 8095.0 20620.0 ;
      RECT  8355.0 20585.0 8285.0 20947.5 ;
      RECT  8320.0 20550.0 8130.0 20620.0 ;
      RECT  8165.0 20242.5 8095.0 20585.0 ;
      RECT  8355.0 20947.5 8285.0 21082.5 ;
      RECT  8165.0 20107.5 8095.0 20242.5 ;
      RECT  8062.5 20550.0 8197.5 20620.0 ;
      RECT  8355.0 22030.0 8285.0 21960.0 ;
      RECT  8165.0 22030.0 8095.0 21960.0 ;
      RECT  8355.0 21995.0 8285.0 21632.5 ;
      RECT  8320.0 22030.0 8130.0 21960.0 ;
      RECT  8165.0 22337.5 8095.0 21995.0 ;
      RECT  8355.0 21632.5 8285.0 21497.5 ;
      RECT  8165.0 22472.5 8095.0 22337.5 ;
      RECT  8062.5 22030.0 8197.5 21960.0 ;
      RECT  9607.5 18370.0 9742.5 18440.0 ;
      RECT  10992.5 17847.5 11127.5 17917.5 ;
      RECT  9332.5 19715.0 9467.5 19785.0 ;
      RECT  10717.5 19282.5 10852.5 19352.5 ;
      RECT  10992.5 20045.0 11127.5 20115.0 ;
      RECT  9057.5 20045.0 9192.5 20115.0 ;
      RECT  10717.5 21390.0 10852.5 21460.0 ;
      RECT  8782.5 21390.0 8917.5 21460.0 ;
      RECT  9607.5 17860.0 9742.5 17930.0 ;
      RECT  9332.5 17645.0 9467.5 17715.0 ;
      RECT  9057.5 19270.0 9192.5 19340.0 ;
      RECT  9332.5 19485.0 9467.5 19555.0 ;
      RECT  9607.5 20550.0 9742.5 20620.0 ;
      RECT  8782.5 20335.0 8917.5 20405.0 ;
      RECT  9057.5 21960.0 9192.5 22030.0 ;
      RECT  8782.5 22175.0 8917.5 22245.0 ;
      RECT  11095.0 17255.0 11025.0 22495.0 ;
      RECT  10820.0 17255.0 10750.0 22495.0 ;
      RECT  9160.0 22635.0 9090.0 27875.0 ;
      RECT  8885.0 22635.0 8815.0 27875.0 ;
      RECT  9710.0 22635.0 9640.0 27875.0 ;
      RECT  9435.0 22635.0 9365.0 27875.0 ;
      RECT  8355.0 23240.0 8285.0 23310.0 ;
      RECT  8165.0 23240.0 8095.0 23310.0 ;
      RECT  8355.0 23275.0 8285.0 23637.5 ;
      RECT  8320.0 23240.0 8130.0 23310.0 ;
      RECT  8165.0 22932.5 8095.0 23275.0 ;
      RECT  8355.0 23637.5 8285.0 23772.5 ;
      RECT  8165.0 22797.5 8095.0 22932.5 ;
      RECT  8062.5 23240.0 8197.5 23310.0 ;
      RECT  8355.0 24720.0 8285.0 24650.0 ;
      RECT  8165.0 24720.0 8095.0 24650.0 ;
      RECT  8355.0 24685.0 8285.0 24322.5 ;
      RECT  8320.0 24720.0 8130.0 24650.0 ;
      RECT  8165.0 25027.5 8095.0 24685.0 ;
      RECT  8355.0 24322.5 8285.0 24187.5 ;
      RECT  8165.0 25162.5 8095.0 25027.5 ;
      RECT  8062.5 24720.0 8197.5 24650.0 ;
      RECT  8355.0 25930.0 8285.0 26000.0 ;
      RECT  8165.0 25930.0 8095.0 26000.0 ;
      RECT  8355.0 25965.0 8285.0 26327.5 ;
      RECT  8320.0 25930.0 8130.0 26000.0 ;
      RECT  8165.0 25622.5 8095.0 25965.0 ;
      RECT  8355.0 26327.5 8285.0 26462.5 ;
      RECT  8165.0 25487.5 8095.0 25622.5 ;
      RECT  8062.5 25930.0 8197.5 26000.0 ;
      RECT  8355.0 27410.0 8285.0 27340.0 ;
      RECT  8165.0 27410.0 8095.0 27340.0 ;
      RECT  8355.0 27375.0 8285.0 27012.5 ;
      RECT  8320.0 27410.0 8130.0 27340.0 ;
      RECT  8165.0 27717.5 8095.0 27375.0 ;
      RECT  8355.0 27012.5 8285.0 26877.5 ;
      RECT  8165.0 27852.5 8095.0 27717.5 ;
      RECT  8062.5 27410.0 8197.5 27340.0 ;
      RECT  9607.5 23750.0 9742.5 23820.0 ;
      RECT  10992.5 23227.5 11127.5 23297.5 ;
      RECT  9332.5 25095.0 9467.5 25165.0 ;
      RECT  10717.5 24662.5 10852.5 24732.5 ;
      RECT  10992.5 25425.0 11127.5 25495.0 ;
      RECT  9057.5 25425.0 9192.5 25495.0 ;
      RECT  10717.5 26770.0 10852.5 26840.0 ;
      RECT  8782.5 26770.0 8917.5 26840.0 ;
      RECT  9607.5 23240.0 9742.5 23310.0 ;
      RECT  9332.5 23025.0 9467.5 23095.0 ;
      RECT  9057.5 24650.0 9192.5 24720.0 ;
      RECT  9332.5 24865.0 9467.5 24935.0 ;
      RECT  9607.5 25930.0 9742.5 26000.0 ;
      RECT  8782.5 25715.0 8917.5 25785.0 ;
      RECT  9057.5 27340.0 9192.5 27410.0 ;
      RECT  8782.5 27555.0 8917.5 27625.0 ;
      RECT  11095.0 22635.0 11025.0 27875.0 ;
      RECT  10820.0 22635.0 10750.0 27875.0 ;
      RECT  7765.0 28312.5 7835.0 29017.5 ;
      RECT  7385.0 28667.5 7455.0 28737.5 ;
      RECT  7765.0 28667.5 7835.0 28737.5 ;
      RECT  7385.0 28702.5 7455.0 29017.5 ;
      RECT  7420.0 28667.5 7800.0 28737.5 ;
      RECT  7765.0 28312.5 7835.0 28702.5 ;
      RECT  7385.0 29017.5 7455.0 29152.5 ;
      RECT  7765.0 29017.5 7835.0 29152.5 ;
      RECT  7765.0 28177.5 7835.0 28312.5 ;
      RECT  7765.0 28635.0 7835.0 28770.0 ;
      RECT  7765.0 30407.5 7835.0 29702.5 ;
      RECT  7385.0 30052.5 7455.0 29982.5 ;
      RECT  7765.0 30052.5 7835.0 29982.5 ;
      RECT  7385.0 30017.5 7455.0 29702.5 ;
      RECT  7420.0 30052.5 7800.0 29982.5 ;
      RECT  7765.0 30407.5 7835.0 30017.5 ;
      RECT  7385.0 29702.5 7455.0 29567.5 ;
      RECT  7765.0 29702.5 7835.0 29567.5 ;
      RECT  7765.0 30542.5 7835.0 30407.5 ;
      RECT  7765.0 30085.0 7835.0 29950.0 ;
      RECT  7765.0 31002.5 7835.0 31707.5 ;
      RECT  7385.0 31357.5 7455.0 31427.5 ;
      RECT  7765.0 31357.5 7835.0 31427.5 ;
      RECT  7385.0 31392.5 7455.0 31707.5 ;
      RECT  7420.0 31357.5 7800.0 31427.5 ;
      RECT  7765.0 31002.5 7835.0 31392.5 ;
      RECT  7385.0 31707.5 7455.0 31842.5 ;
      RECT  7765.0 31707.5 7835.0 31842.5 ;
      RECT  7765.0 30867.5 7835.0 31002.5 ;
      RECT  7765.0 31325.0 7835.0 31460.0 ;
      RECT  7765.0 33097.5 7835.0 32392.5 ;
      RECT  7385.0 32742.5 7455.0 32672.5 ;
      RECT  7765.0 32742.5 7835.0 32672.5 ;
      RECT  7385.0 32707.5 7455.0 32392.5 ;
      RECT  7420.0 32742.5 7800.0 32672.5 ;
      RECT  7765.0 33097.5 7835.0 32707.5 ;
      RECT  7385.0 32392.5 7455.0 32257.5 ;
      RECT  7765.0 32392.5 7835.0 32257.5 ;
      RECT  7765.0 33232.5 7835.0 33097.5 ;
      RECT  7765.0 32775.0 7835.0 32640.0 ;
      RECT  7765.0 33692.5 7835.0 34397.5 ;
      RECT  7385.0 34047.5 7455.0 34117.5 ;
      RECT  7765.0 34047.5 7835.0 34117.5 ;
      RECT  7385.0 34082.5 7455.0 34397.5 ;
      RECT  7420.0 34047.5 7800.0 34117.5 ;
      RECT  7765.0 33692.5 7835.0 34082.5 ;
      RECT  7385.0 34397.5 7455.0 34532.5 ;
      RECT  7765.0 34397.5 7835.0 34532.5 ;
      RECT  7765.0 33557.5 7835.0 33692.5 ;
      RECT  7765.0 34015.0 7835.0 34150.0 ;
      RECT  7765.0 35787.5 7835.0 35082.5 ;
      RECT  7385.0 35432.5 7455.0 35362.5 ;
      RECT  7765.0 35432.5 7835.0 35362.5 ;
      RECT  7385.0 35397.5 7455.0 35082.5 ;
      RECT  7420.0 35432.5 7800.0 35362.5 ;
      RECT  7765.0 35787.5 7835.0 35397.5 ;
      RECT  7385.0 35082.5 7455.0 34947.5 ;
      RECT  7765.0 35082.5 7835.0 34947.5 ;
      RECT  7765.0 35922.5 7835.0 35787.5 ;
      RECT  7765.0 35465.0 7835.0 35330.0 ;
      RECT  7765.0 36382.5 7835.0 37087.5 ;
      RECT  7385.0 36737.5 7455.0 36807.5 ;
      RECT  7765.0 36737.5 7835.0 36807.5 ;
      RECT  7385.0 36772.5 7455.0 37087.5 ;
      RECT  7420.0 36737.5 7800.0 36807.5 ;
      RECT  7765.0 36382.5 7835.0 36772.5 ;
      RECT  7385.0 37087.5 7455.0 37222.5 ;
      RECT  7765.0 37087.5 7835.0 37222.5 ;
      RECT  7765.0 36247.5 7835.0 36382.5 ;
      RECT  7765.0 36705.0 7835.0 36840.0 ;
      RECT  7765.0 38477.5 7835.0 37772.5 ;
      RECT  7385.0 38122.5 7455.0 38052.5 ;
      RECT  7765.0 38122.5 7835.0 38052.5 ;
      RECT  7385.0 38087.5 7455.0 37772.5 ;
      RECT  7420.0 38122.5 7800.0 38052.5 ;
      RECT  7765.0 38477.5 7835.0 38087.5 ;
      RECT  7385.0 37772.5 7455.0 37637.5 ;
      RECT  7765.0 37772.5 7835.0 37637.5 ;
      RECT  7765.0 38612.5 7835.0 38477.5 ;
      RECT  7765.0 38155.0 7835.0 38020.0 ;
      RECT  7765.0 39072.5 7835.0 39777.5 ;
      RECT  7385.0 39427.5 7455.0 39497.5 ;
      RECT  7765.0 39427.5 7835.0 39497.5 ;
      RECT  7385.0 39462.5 7455.0 39777.5 ;
      RECT  7420.0 39427.5 7800.0 39497.5 ;
      RECT  7765.0 39072.5 7835.0 39462.5 ;
      RECT  7385.0 39777.5 7455.0 39912.5 ;
      RECT  7765.0 39777.5 7835.0 39912.5 ;
      RECT  7765.0 38937.5 7835.0 39072.5 ;
      RECT  7765.0 39395.0 7835.0 39530.0 ;
      RECT  7765.0 41167.5 7835.0 40462.5 ;
      RECT  7385.0 40812.5 7455.0 40742.5 ;
      RECT  7765.0 40812.5 7835.0 40742.5 ;
      RECT  7385.0 40777.5 7455.0 40462.5 ;
      RECT  7420.0 40812.5 7800.0 40742.5 ;
      RECT  7765.0 41167.5 7835.0 40777.5 ;
      RECT  7385.0 40462.5 7455.0 40327.5 ;
      RECT  7765.0 40462.5 7835.0 40327.5 ;
      RECT  7765.0 41302.5 7835.0 41167.5 ;
      RECT  7765.0 40845.0 7835.0 40710.0 ;
      RECT  7765.0 41762.5 7835.0 42467.5 ;
      RECT  7385.0 42117.5 7455.0 42187.5 ;
      RECT  7765.0 42117.5 7835.0 42187.5 ;
      RECT  7385.0 42152.5 7455.0 42467.5 ;
      RECT  7420.0 42117.5 7800.0 42187.5 ;
      RECT  7765.0 41762.5 7835.0 42152.5 ;
      RECT  7385.0 42467.5 7455.0 42602.5 ;
      RECT  7765.0 42467.5 7835.0 42602.5 ;
      RECT  7765.0 41627.5 7835.0 41762.5 ;
      RECT  7765.0 42085.0 7835.0 42220.0 ;
      RECT  7765.0 43857.5 7835.0 43152.5 ;
      RECT  7385.0 43502.5 7455.0 43432.5 ;
      RECT  7765.0 43502.5 7835.0 43432.5 ;
      RECT  7385.0 43467.5 7455.0 43152.5 ;
      RECT  7420.0 43502.5 7800.0 43432.5 ;
      RECT  7765.0 43857.5 7835.0 43467.5 ;
      RECT  7385.0 43152.5 7455.0 43017.5 ;
      RECT  7765.0 43152.5 7835.0 43017.5 ;
      RECT  7765.0 43992.5 7835.0 43857.5 ;
      RECT  7765.0 43535.0 7835.0 43400.0 ;
      RECT  7765.0 44452.5 7835.0 45157.5 ;
      RECT  7385.0 44807.5 7455.0 44877.5 ;
      RECT  7765.0 44807.5 7835.0 44877.5 ;
      RECT  7385.0 44842.5 7455.0 45157.5 ;
      RECT  7420.0 44807.5 7800.0 44877.5 ;
      RECT  7765.0 44452.5 7835.0 44842.5 ;
      RECT  7385.0 45157.5 7455.0 45292.5 ;
      RECT  7765.0 45157.5 7835.0 45292.5 ;
      RECT  7765.0 44317.5 7835.0 44452.5 ;
      RECT  7765.0 44775.0 7835.0 44910.0 ;
      RECT  7765.0 46547.5 7835.0 45842.5 ;
      RECT  7385.0 46192.5 7455.0 46122.5 ;
      RECT  7765.0 46192.5 7835.0 46122.5 ;
      RECT  7385.0 46157.5 7455.0 45842.5 ;
      RECT  7420.0 46192.5 7800.0 46122.5 ;
      RECT  7765.0 46547.5 7835.0 46157.5 ;
      RECT  7385.0 45842.5 7455.0 45707.5 ;
      RECT  7765.0 45842.5 7835.0 45707.5 ;
      RECT  7765.0 46682.5 7835.0 46547.5 ;
      RECT  7765.0 46225.0 7835.0 46090.0 ;
      RECT  7765.0 47142.5 7835.0 47847.5 ;
      RECT  7385.0 47497.5 7455.0 47567.5 ;
      RECT  7765.0 47497.5 7835.0 47567.5 ;
      RECT  7385.0 47532.5 7455.0 47847.5 ;
      RECT  7420.0 47497.5 7800.0 47567.5 ;
      RECT  7765.0 47142.5 7835.0 47532.5 ;
      RECT  7385.0 47847.5 7455.0 47982.5 ;
      RECT  7765.0 47847.5 7835.0 47982.5 ;
      RECT  7765.0 47007.5 7835.0 47142.5 ;
      RECT  7765.0 47465.0 7835.0 47600.0 ;
      RECT  7765.0 49237.5 7835.0 48532.5 ;
      RECT  7385.0 48882.5 7455.0 48812.5 ;
      RECT  7765.0 48882.5 7835.0 48812.5 ;
      RECT  7385.0 48847.5 7455.0 48532.5 ;
      RECT  7420.0 48882.5 7800.0 48812.5 ;
      RECT  7765.0 49237.5 7835.0 48847.5 ;
      RECT  7385.0 48532.5 7455.0 48397.5 ;
      RECT  7765.0 48532.5 7835.0 48397.5 ;
      RECT  7765.0 49372.5 7835.0 49237.5 ;
      RECT  7765.0 48915.0 7835.0 48780.0 ;
      RECT  7765.0 49832.5 7835.0 50537.5 ;
      RECT  7385.0 50187.5 7455.0 50257.5 ;
      RECT  7765.0 50187.5 7835.0 50257.5 ;
      RECT  7385.0 50222.5 7455.0 50537.5 ;
      RECT  7420.0 50187.5 7800.0 50257.5 ;
      RECT  7765.0 49832.5 7835.0 50222.5 ;
      RECT  7385.0 50537.5 7455.0 50672.5 ;
      RECT  7765.0 50537.5 7835.0 50672.5 ;
      RECT  7765.0 49697.5 7835.0 49832.5 ;
      RECT  7765.0 50155.0 7835.0 50290.0 ;
      RECT  7765.0 51927.5 7835.0 51222.5 ;
      RECT  7385.0 51572.5 7455.0 51502.5 ;
      RECT  7765.0 51572.5 7835.0 51502.5 ;
      RECT  7385.0 51537.5 7455.0 51222.5 ;
      RECT  7420.0 51572.5 7800.0 51502.5 ;
      RECT  7765.0 51927.5 7835.0 51537.5 ;
      RECT  7385.0 51222.5 7455.0 51087.5 ;
      RECT  7765.0 51222.5 7835.0 51087.5 ;
      RECT  7765.0 52062.5 7835.0 51927.5 ;
      RECT  7765.0 51605.0 7835.0 51470.0 ;
      RECT  7765.0 52522.5 7835.0 53227.5 ;
      RECT  7385.0 52877.5 7455.0 52947.5 ;
      RECT  7765.0 52877.5 7835.0 52947.5 ;
      RECT  7385.0 52912.5 7455.0 53227.5 ;
      RECT  7420.0 52877.5 7800.0 52947.5 ;
      RECT  7765.0 52522.5 7835.0 52912.5 ;
      RECT  7385.0 53227.5 7455.0 53362.5 ;
      RECT  7765.0 53227.5 7835.0 53362.5 ;
      RECT  7765.0 52387.5 7835.0 52522.5 ;
      RECT  7765.0 52845.0 7835.0 52980.0 ;
      RECT  7765.0 54617.5 7835.0 53912.5 ;
      RECT  7385.0 54262.5 7455.0 54192.5 ;
      RECT  7765.0 54262.5 7835.0 54192.5 ;
      RECT  7385.0 54227.5 7455.0 53912.5 ;
      RECT  7420.0 54262.5 7800.0 54192.5 ;
      RECT  7765.0 54617.5 7835.0 54227.5 ;
      RECT  7385.0 53912.5 7455.0 53777.5 ;
      RECT  7765.0 53912.5 7835.0 53777.5 ;
      RECT  7765.0 54752.5 7835.0 54617.5 ;
      RECT  7765.0 54295.0 7835.0 54160.0 ;
      RECT  7765.0 55212.5 7835.0 55917.5 ;
      RECT  7385.0 55567.5 7455.0 55637.5 ;
      RECT  7765.0 55567.5 7835.0 55637.5 ;
      RECT  7385.0 55602.5 7455.0 55917.5 ;
      RECT  7420.0 55567.5 7800.0 55637.5 ;
      RECT  7765.0 55212.5 7835.0 55602.5 ;
      RECT  7385.0 55917.5 7455.0 56052.5 ;
      RECT  7765.0 55917.5 7835.0 56052.5 ;
      RECT  7765.0 55077.5 7835.0 55212.5 ;
      RECT  7765.0 55535.0 7835.0 55670.0 ;
      RECT  7765.0 57307.5 7835.0 56602.5 ;
      RECT  7385.0 56952.5 7455.0 56882.5 ;
      RECT  7765.0 56952.5 7835.0 56882.5 ;
      RECT  7385.0 56917.5 7455.0 56602.5 ;
      RECT  7420.0 56952.5 7800.0 56882.5 ;
      RECT  7765.0 57307.5 7835.0 56917.5 ;
      RECT  7385.0 56602.5 7455.0 56467.5 ;
      RECT  7765.0 56602.5 7835.0 56467.5 ;
      RECT  7765.0 57442.5 7835.0 57307.5 ;
      RECT  7765.0 56985.0 7835.0 56850.0 ;
      RECT  7765.0 57902.5 7835.0 58607.5 ;
      RECT  7385.0 58257.5 7455.0 58327.5 ;
      RECT  7765.0 58257.5 7835.0 58327.5 ;
      RECT  7385.0 58292.5 7455.0 58607.5 ;
      RECT  7420.0 58257.5 7800.0 58327.5 ;
      RECT  7765.0 57902.5 7835.0 58292.5 ;
      RECT  7385.0 58607.5 7455.0 58742.5 ;
      RECT  7765.0 58607.5 7835.0 58742.5 ;
      RECT  7765.0 57767.5 7835.0 57902.5 ;
      RECT  7765.0 58225.0 7835.0 58360.0 ;
      RECT  7765.0 59997.5 7835.0 59292.5 ;
      RECT  7385.0 59642.5 7455.0 59572.5 ;
      RECT  7765.0 59642.5 7835.0 59572.5 ;
      RECT  7385.0 59607.5 7455.0 59292.5 ;
      RECT  7420.0 59642.5 7800.0 59572.5 ;
      RECT  7765.0 59997.5 7835.0 59607.5 ;
      RECT  7385.0 59292.5 7455.0 59157.5 ;
      RECT  7765.0 59292.5 7835.0 59157.5 ;
      RECT  7765.0 60132.5 7835.0 59997.5 ;
      RECT  7765.0 59675.0 7835.0 59540.0 ;
      RECT  7765.0 60592.5 7835.0 61297.5 ;
      RECT  7385.0 60947.5 7455.0 61017.5 ;
      RECT  7765.0 60947.5 7835.0 61017.5 ;
      RECT  7385.0 60982.5 7455.0 61297.5 ;
      RECT  7420.0 60947.5 7800.0 61017.5 ;
      RECT  7765.0 60592.5 7835.0 60982.5 ;
      RECT  7385.0 61297.5 7455.0 61432.5 ;
      RECT  7765.0 61297.5 7835.0 61432.5 ;
      RECT  7765.0 60457.5 7835.0 60592.5 ;
      RECT  7765.0 60915.0 7835.0 61050.0 ;
      RECT  7765.0 62687.5 7835.0 61982.5 ;
      RECT  7385.0 62332.5 7455.0 62262.5 ;
      RECT  7765.0 62332.5 7835.0 62262.5 ;
      RECT  7385.0 62297.5 7455.0 61982.5 ;
      RECT  7420.0 62332.5 7800.0 62262.5 ;
      RECT  7765.0 62687.5 7835.0 62297.5 ;
      RECT  7385.0 61982.5 7455.0 61847.5 ;
      RECT  7765.0 61982.5 7835.0 61847.5 ;
      RECT  7765.0 62822.5 7835.0 62687.5 ;
      RECT  7765.0 62365.0 7835.0 62230.0 ;
      RECT  7765.0 63282.5 7835.0 63987.5 ;
      RECT  7385.0 63637.5 7455.0 63707.5 ;
      RECT  7765.0 63637.5 7835.0 63707.5 ;
      RECT  7385.0 63672.5 7455.0 63987.5 ;
      RECT  7420.0 63637.5 7800.0 63707.5 ;
      RECT  7765.0 63282.5 7835.0 63672.5 ;
      RECT  7385.0 63987.5 7455.0 64122.5 ;
      RECT  7765.0 63987.5 7835.0 64122.5 ;
      RECT  7765.0 63147.5 7835.0 63282.5 ;
      RECT  7765.0 63605.0 7835.0 63740.0 ;
      RECT  7765.0 65377.5 7835.0 64672.5 ;
      RECT  7385.0 65022.5 7455.0 64952.5 ;
      RECT  7765.0 65022.5 7835.0 64952.5 ;
      RECT  7385.0 64987.5 7455.0 64672.5 ;
      RECT  7420.0 65022.5 7800.0 64952.5 ;
      RECT  7765.0 65377.5 7835.0 64987.5 ;
      RECT  7385.0 64672.5 7455.0 64537.5 ;
      RECT  7765.0 64672.5 7835.0 64537.5 ;
      RECT  7765.0 65512.5 7835.0 65377.5 ;
      RECT  7765.0 65055.0 7835.0 64920.0 ;
      RECT  7765.0 65972.5 7835.0 66677.5 ;
      RECT  7385.0 66327.5 7455.0 66397.5 ;
      RECT  7765.0 66327.5 7835.0 66397.5 ;
      RECT  7385.0 66362.5 7455.0 66677.5 ;
      RECT  7420.0 66327.5 7800.0 66397.5 ;
      RECT  7765.0 65972.5 7835.0 66362.5 ;
      RECT  7385.0 66677.5 7455.0 66812.5 ;
      RECT  7765.0 66677.5 7835.0 66812.5 ;
      RECT  7765.0 65837.5 7835.0 65972.5 ;
      RECT  7765.0 66295.0 7835.0 66430.0 ;
      RECT  7765.0 68067.5 7835.0 67362.5 ;
      RECT  7385.0 67712.5 7455.0 67642.5 ;
      RECT  7765.0 67712.5 7835.0 67642.5 ;
      RECT  7385.0 67677.5 7455.0 67362.5 ;
      RECT  7420.0 67712.5 7800.0 67642.5 ;
      RECT  7765.0 68067.5 7835.0 67677.5 ;
      RECT  7385.0 67362.5 7455.0 67227.5 ;
      RECT  7765.0 67362.5 7835.0 67227.5 ;
      RECT  7765.0 68202.5 7835.0 68067.5 ;
      RECT  7765.0 67745.0 7835.0 67610.0 ;
      RECT  7765.0 68662.5 7835.0 69367.5 ;
      RECT  7385.0 69017.5 7455.0 69087.5 ;
      RECT  7765.0 69017.5 7835.0 69087.5 ;
      RECT  7385.0 69052.5 7455.0 69367.5 ;
      RECT  7420.0 69017.5 7800.0 69087.5 ;
      RECT  7765.0 68662.5 7835.0 69052.5 ;
      RECT  7385.0 69367.5 7455.0 69502.5 ;
      RECT  7765.0 69367.5 7835.0 69502.5 ;
      RECT  7765.0 68527.5 7835.0 68662.5 ;
      RECT  7765.0 68985.0 7835.0 69120.0 ;
      RECT  7765.0 70757.5 7835.0 70052.5 ;
      RECT  7385.0 70402.5 7455.0 70332.5 ;
      RECT  7765.0 70402.5 7835.0 70332.5 ;
      RECT  7385.0 70367.5 7455.0 70052.5 ;
      RECT  7420.0 70402.5 7800.0 70332.5 ;
      RECT  7765.0 70757.5 7835.0 70367.5 ;
      RECT  7385.0 70052.5 7455.0 69917.5 ;
      RECT  7765.0 70052.5 7835.0 69917.5 ;
      RECT  7765.0 70892.5 7835.0 70757.5 ;
      RECT  7765.0 70435.0 7835.0 70300.0 ;
      RECT  7765.0 71352.5 7835.0 72057.5 ;
      RECT  7385.0 71707.5 7455.0 71777.5 ;
      RECT  7765.0 71707.5 7835.0 71777.5 ;
      RECT  7385.0 71742.5 7455.0 72057.5 ;
      RECT  7420.0 71707.5 7800.0 71777.5 ;
      RECT  7765.0 71352.5 7835.0 71742.5 ;
      RECT  7385.0 72057.5 7455.0 72192.5 ;
      RECT  7765.0 72057.5 7835.0 72192.5 ;
      RECT  7765.0 71217.5 7835.0 71352.5 ;
      RECT  7765.0 71675.0 7835.0 71810.0 ;
      RECT  7765.0 73447.5 7835.0 72742.5 ;
      RECT  7385.0 73092.5 7455.0 73022.5 ;
      RECT  7765.0 73092.5 7835.0 73022.5 ;
      RECT  7385.0 73057.5 7455.0 72742.5 ;
      RECT  7420.0 73092.5 7800.0 73022.5 ;
      RECT  7765.0 73447.5 7835.0 73057.5 ;
      RECT  7385.0 72742.5 7455.0 72607.5 ;
      RECT  7765.0 72742.5 7835.0 72607.5 ;
      RECT  7765.0 73582.5 7835.0 73447.5 ;
      RECT  7765.0 73125.0 7835.0 72990.0 ;
      RECT  7765.0 74042.5 7835.0 74747.5 ;
      RECT  7385.0 74397.5 7455.0 74467.5 ;
      RECT  7765.0 74397.5 7835.0 74467.5 ;
      RECT  7385.0 74432.5 7455.0 74747.5 ;
      RECT  7420.0 74397.5 7800.0 74467.5 ;
      RECT  7765.0 74042.5 7835.0 74432.5 ;
      RECT  7385.0 74747.5 7455.0 74882.5 ;
      RECT  7765.0 74747.5 7835.0 74882.5 ;
      RECT  7765.0 73907.5 7835.0 74042.5 ;
      RECT  7765.0 74365.0 7835.0 74500.0 ;
      RECT  7765.0 76137.5 7835.0 75432.5 ;
      RECT  7385.0 75782.5 7455.0 75712.5 ;
      RECT  7765.0 75782.5 7835.0 75712.5 ;
      RECT  7385.0 75747.5 7455.0 75432.5 ;
      RECT  7420.0 75782.5 7800.0 75712.5 ;
      RECT  7765.0 76137.5 7835.0 75747.5 ;
      RECT  7385.0 75432.5 7455.0 75297.5 ;
      RECT  7765.0 75432.5 7835.0 75297.5 ;
      RECT  7765.0 76272.5 7835.0 76137.5 ;
      RECT  7765.0 75815.0 7835.0 75680.0 ;
      RECT  7765.0 76732.5 7835.0 77437.5 ;
      RECT  7385.0 77087.5 7455.0 77157.5 ;
      RECT  7765.0 77087.5 7835.0 77157.5 ;
      RECT  7385.0 77122.5 7455.0 77437.5 ;
      RECT  7420.0 77087.5 7800.0 77157.5 ;
      RECT  7765.0 76732.5 7835.0 77122.5 ;
      RECT  7385.0 77437.5 7455.0 77572.5 ;
      RECT  7765.0 77437.5 7835.0 77572.5 ;
      RECT  7765.0 76597.5 7835.0 76732.5 ;
      RECT  7765.0 77055.0 7835.0 77190.0 ;
      RECT  7765.0 78827.5 7835.0 78122.5 ;
      RECT  7385.0 78472.5 7455.0 78402.5 ;
      RECT  7765.0 78472.5 7835.0 78402.5 ;
      RECT  7385.0 78437.5 7455.0 78122.5 ;
      RECT  7420.0 78472.5 7800.0 78402.5 ;
      RECT  7765.0 78827.5 7835.0 78437.5 ;
      RECT  7385.0 78122.5 7455.0 77987.5 ;
      RECT  7765.0 78122.5 7835.0 77987.5 ;
      RECT  7765.0 78962.5 7835.0 78827.5 ;
      RECT  7765.0 78505.0 7835.0 78370.0 ;
      RECT  7765.0 79422.5 7835.0 80127.5 ;
      RECT  7385.0 79777.5 7455.0 79847.5 ;
      RECT  7765.0 79777.5 7835.0 79847.5 ;
      RECT  7385.0 79812.5 7455.0 80127.5 ;
      RECT  7420.0 79777.5 7800.0 79847.5 ;
      RECT  7765.0 79422.5 7835.0 79812.5 ;
      RECT  7385.0 80127.5 7455.0 80262.5 ;
      RECT  7765.0 80127.5 7835.0 80262.5 ;
      RECT  7765.0 79287.5 7835.0 79422.5 ;
      RECT  7765.0 79745.0 7835.0 79880.0 ;
      RECT  7765.0 81517.5 7835.0 80812.5 ;
      RECT  7385.0 81162.5 7455.0 81092.5 ;
      RECT  7765.0 81162.5 7835.0 81092.5 ;
      RECT  7385.0 81127.5 7455.0 80812.5 ;
      RECT  7420.0 81162.5 7800.0 81092.5 ;
      RECT  7765.0 81517.5 7835.0 81127.5 ;
      RECT  7385.0 80812.5 7455.0 80677.5 ;
      RECT  7765.0 80812.5 7835.0 80677.5 ;
      RECT  7765.0 81652.5 7835.0 81517.5 ;
      RECT  7765.0 81195.0 7835.0 81060.0 ;
      RECT  7765.0 82112.5 7835.0 82817.5 ;
      RECT  7385.0 82467.5 7455.0 82537.5 ;
      RECT  7765.0 82467.5 7835.0 82537.5 ;
      RECT  7385.0 82502.5 7455.0 82817.5 ;
      RECT  7420.0 82467.5 7800.0 82537.5 ;
      RECT  7765.0 82112.5 7835.0 82502.5 ;
      RECT  7385.0 82817.5 7455.0 82952.5 ;
      RECT  7765.0 82817.5 7835.0 82952.5 ;
      RECT  7765.0 81977.5 7835.0 82112.5 ;
      RECT  7765.0 82435.0 7835.0 82570.0 ;
      RECT  7765.0 84207.5 7835.0 83502.5 ;
      RECT  7385.0 83852.5 7455.0 83782.5 ;
      RECT  7765.0 83852.5 7835.0 83782.5 ;
      RECT  7385.0 83817.5 7455.0 83502.5 ;
      RECT  7420.0 83852.5 7800.0 83782.5 ;
      RECT  7765.0 84207.5 7835.0 83817.5 ;
      RECT  7385.0 83502.5 7455.0 83367.5 ;
      RECT  7765.0 83502.5 7835.0 83367.5 ;
      RECT  7765.0 84342.5 7835.0 84207.5 ;
      RECT  7765.0 83885.0 7835.0 83750.0 ;
      RECT  7765.0 84802.5 7835.0 85507.5 ;
      RECT  7385.0 85157.5 7455.0 85227.5 ;
      RECT  7765.0 85157.5 7835.0 85227.5 ;
      RECT  7385.0 85192.5 7455.0 85507.5 ;
      RECT  7420.0 85157.5 7800.0 85227.5 ;
      RECT  7765.0 84802.5 7835.0 85192.5 ;
      RECT  7385.0 85507.5 7455.0 85642.5 ;
      RECT  7765.0 85507.5 7835.0 85642.5 ;
      RECT  7765.0 84667.5 7835.0 84802.5 ;
      RECT  7765.0 85125.0 7835.0 85260.0 ;
      RECT  7765.0 86897.5 7835.0 86192.5 ;
      RECT  7385.0 86542.5 7455.0 86472.5 ;
      RECT  7765.0 86542.5 7835.0 86472.5 ;
      RECT  7385.0 86507.5 7455.0 86192.5 ;
      RECT  7420.0 86542.5 7800.0 86472.5 ;
      RECT  7765.0 86897.5 7835.0 86507.5 ;
      RECT  7385.0 86192.5 7455.0 86057.5 ;
      RECT  7765.0 86192.5 7835.0 86057.5 ;
      RECT  7765.0 87032.5 7835.0 86897.5 ;
      RECT  7765.0 86575.0 7835.0 86440.0 ;
      RECT  7765.0 87492.5 7835.0 88197.5 ;
      RECT  7385.0 87847.5 7455.0 87917.5 ;
      RECT  7765.0 87847.5 7835.0 87917.5 ;
      RECT  7385.0 87882.5 7455.0 88197.5 ;
      RECT  7420.0 87847.5 7800.0 87917.5 ;
      RECT  7765.0 87492.5 7835.0 87882.5 ;
      RECT  7385.0 88197.5 7455.0 88332.5 ;
      RECT  7765.0 88197.5 7835.0 88332.5 ;
      RECT  7765.0 87357.5 7835.0 87492.5 ;
      RECT  7765.0 87815.0 7835.0 87950.0 ;
      RECT  7765.0 89587.5 7835.0 88882.5 ;
      RECT  7385.0 89232.5 7455.0 89162.5 ;
      RECT  7765.0 89232.5 7835.0 89162.5 ;
      RECT  7385.0 89197.5 7455.0 88882.5 ;
      RECT  7420.0 89232.5 7800.0 89162.5 ;
      RECT  7765.0 89587.5 7835.0 89197.5 ;
      RECT  7385.0 88882.5 7455.0 88747.5 ;
      RECT  7765.0 88882.5 7835.0 88747.5 ;
      RECT  7765.0 89722.5 7835.0 89587.5 ;
      RECT  7765.0 89265.0 7835.0 89130.0 ;
      RECT  7765.0 90182.5 7835.0 90887.5 ;
      RECT  7385.0 90537.5 7455.0 90607.5 ;
      RECT  7765.0 90537.5 7835.0 90607.5 ;
      RECT  7385.0 90572.5 7455.0 90887.5 ;
      RECT  7420.0 90537.5 7800.0 90607.5 ;
      RECT  7765.0 90182.5 7835.0 90572.5 ;
      RECT  7385.0 90887.5 7455.0 91022.5 ;
      RECT  7765.0 90887.5 7835.0 91022.5 ;
      RECT  7765.0 90047.5 7835.0 90182.5 ;
      RECT  7765.0 90505.0 7835.0 90640.0 ;
      RECT  7765.0 92277.5 7835.0 91572.5 ;
      RECT  7385.0 91922.5 7455.0 91852.5 ;
      RECT  7765.0 91922.5 7835.0 91852.5 ;
      RECT  7385.0 91887.5 7455.0 91572.5 ;
      RECT  7420.0 91922.5 7800.0 91852.5 ;
      RECT  7765.0 92277.5 7835.0 91887.5 ;
      RECT  7385.0 91572.5 7455.0 91437.5 ;
      RECT  7765.0 91572.5 7835.0 91437.5 ;
      RECT  7765.0 92412.5 7835.0 92277.5 ;
      RECT  7765.0 91955.0 7835.0 91820.0 ;
      RECT  7765.0 92872.5 7835.0 93577.5 ;
      RECT  7385.0 93227.5 7455.0 93297.5 ;
      RECT  7765.0 93227.5 7835.0 93297.5 ;
      RECT  7385.0 93262.5 7455.0 93577.5 ;
      RECT  7420.0 93227.5 7800.0 93297.5 ;
      RECT  7765.0 92872.5 7835.0 93262.5 ;
      RECT  7385.0 93577.5 7455.0 93712.5 ;
      RECT  7765.0 93577.5 7835.0 93712.5 ;
      RECT  7765.0 92737.5 7835.0 92872.5 ;
      RECT  7765.0 93195.0 7835.0 93330.0 ;
      RECT  7765.0 94967.5 7835.0 94262.5 ;
      RECT  7385.0 94612.5 7455.0 94542.5 ;
      RECT  7765.0 94612.5 7835.0 94542.5 ;
      RECT  7385.0 94577.5 7455.0 94262.5 ;
      RECT  7420.0 94612.5 7800.0 94542.5 ;
      RECT  7765.0 94967.5 7835.0 94577.5 ;
      RECT  7385.0 94262.5 7455.0 94127.5 ;
      RECT  7765.0 94262.5 7835.0 94127.5 ;
      RECT  7765.0 95102.5 7835.0 94967.5 ;
      RECT  7765.0 94645.0 7835.0 94510.0 ;
      RECT  7765.0 95562.5 7835.0 96267.5 ;
      RECT  7385.0 95917.5 7455.0 95987.5 ;
      RECT  7765.0 95917.5 7835.0 95987.5 ;
      RECT  7385.0 95952.5 7455.0 96267.5 ;
      RECT  7420.0 95917.5 7800.0 95987.5 ;
      RECT  7765.0 95562.5 7835.0 95952.5 ;
      RECT  7385.0 96267.5 7455.0 96402.5 ;
      RECT  7765.0 96267.5 7835.0 96402.5 ;
      RECT  7765.0 95427.5 7835.0 95562.5 ;
      RECT  7765.0 95885.0 7835.0 96020.0 ;
      RECT  7765.0 97657.5 7835.0 96952.5 ;
      RECT  7385.0 97302.5 7455.0 97232.5 ;
      RECT  7765.0 97302.5 7835.0 97232.5 ;
      RECT  7385.0 97267.5 7455.0 96952.5 ;
      RECT  7420.0 97302.5 7800.0 97232.5 ;
      RECT  7765.0 97657.5 7835.0 97267.5 ;
      RECT  7385.0 96952.5 7455.0 96817.5 ;
      RECT  7765.0 96952.5 7835.0 96817.5 ;
      RECT  7765.0 97792.5 7835.0 97657.5 ;
      RECT  7765.0 97335.0 7835.0 97200.0 ;
      RECT  7765.0 98252.5 7835.0 98957.5 ;
      RECT  7385.0 98607.5 7455.0 98677.5 ;
      RECT  7765.0 98607.5 7835.0 98677.5 ;
      RECT  7385.0 98642.5 7455.0 98957.5 ;
      RECT  7420.0 98607.5 7800.0 98677.5 ;
      RECT  7765.0 98252.5 7835.0 98642.5 ;
      RECT  7385.0 98957.5 7455.0 99092.5 ;
      RECT  7765.0 98957.5 7835.0 99092.5 ;
      RECT  7765.0 98117.5 7835.0 98252.5 ;
      RECT  7765.0 98575.0 7835.0 98710.0 ;
      RECT  7765.0 100347.5 7835.0 99642.5 ;
      RECT  7385.0 99992.5 7455.0 99922.5 ;
      RECT  7765.0 99992.5 7835.0 99922.5 ;
      RECT  7385.0 99957.5 7455.0 99642.5 ;
      RECT  7420.0 99992.5 7800.0 99922.5 ;
      RECT  7765.0 100347.5 7835.0 99957.5 ;
      RECT  7385.0 99642.5 7455.0 99507.5 ;
      RECT  7765.0 99642.5 7835.0 99507.5 ;
      RECT  7765.0 100482.5 7835.0 100347.5 ;
      RECT  7765.0 100025.0 7835.0 99890.0 ;
      RECT  7765.0 100942.5 7835.0 101647.5 ;
      RECT  7385.0 101297.5 7455.0 101367.5 ;
      RECT  7765.0 101297.5 7835.0 101367.5 ;
      RECT  7385.0 101332.5 7455.0 101647.5 ;
      RECT  7420.0 101297.5 7800.0 101367.5 ;
      RECT  7765.0 100942.5 7835.0 101332.5 ;
      RECT  7385.0 101647.5 7455.0 101782.5 ;
      RECT  7765.0 101647.5 7835.0 101782.5 ;
      RECT  7765.0 100807.5 7835.0 100942.5 ;
      RECT  7765.0 101265.0 7835.0 101400.0 ;
      RECT  7765.0 103037.5 7835.0 102332.5 ;
      RECT  7385.0 102682.5 7455.0 102612.5 ;
      RECT  7765.0 102682.5 7835.0 102612.5 ;
      RECT  7385.0 102647.5 7455.0 102332.5 ;
      RECT  7420.0 102682.5 7800.0 102612.5 ;
      RECT  7765.0 103037.5 7835.0 102647.5 ;
      RECT  7385.0 102332.5 7455.0 102197.5 ;
      RECT  7765.0 102332.5 7835.0 102197.5 ;
      RECT  7765.0 103172.5 7835.0 103037.5 ;
      RECT  7765.0 102715.0 7835.0 102580.0 ;
      RECT  7765.0 103632.5 7835.0 104337.5 ;
      RECT  7385.0 103987.5 7455.0 104057.5 ;
      RECT  7765.0 103987.5 7835.0 104057.5 ;
      RECT  7385.0 104022.5 7455.0 104337.5 ;
      RECT  7420.0 103987.5 7800.0 104057.5 ;
      RECT  7765.0 103632.5 7835.0 104022.5 ;
      RECT  7385.0 104337.5 7455.0 104472.5 ;
      RECT  7765.0 104337.5 7835.0 104472.5 ;
      RECT  7765.0 103497.5 7835.0 103632.5 ;
      RECT  7765.0 103955.0 7835.0 104090.0 ;
      RECT  7765.0 105727.5 7835.0 105022.5 ;
      RECT  7385.0 105372.5 7455.0 105302.5 ;
      RECT  7765.0 105372.5 7835.0 105302.5 ;
      RECT  7385.0 105337.5 7455.0 105022.5 ;
      RECT  7420.0 105372.5 7800.0 105302.5 ;
      RECT  7765.0 105727.5 7835.0 105337.5 ;
      RECT  7385.0 105022.5 7455.0 104887.5 ;
      RECT  7765.0 105022.5 7835.0 104887.5 ;
      RECT  7765.0 105862.5 7835.0 105727.5 ;
      RECT  7765.0 105405.0 7835.0 105270.0 ;
      RECT  7765.0 106322.5 7835.0 107027.5 ;
      RECT  7385.0 106677.5 7455.0 106747.5 ;
      RECT  7765.0 106677.5 7835.0 106747.5 ;
      RECT  7385.0 106712.5 7455.0 107027.5 ;
      RECT  7420.0 106677.5 7800.0 106747.5 ;
      RECT  7765.0 106322.5 7835.0 106712.5 ;
      RECT  7385.0 107027.5 7455.0 107162.5 ;
      RECT  7765.0 107027.5 7835.0 107162.5 ;
      RECT  7765.0 106187.5 7835.0 106322.5 ;
      RECT  7765.0 106645.0 7835.0 106780.0 ;
      RECT  7765.0 108417.5 7835.0 107712.5 ;
      RECT  7385.0 108062.5 7455.0 107992.5 ;
      RECT  7765.0 108062.5 7835.0 107992.5 ;
      RECT  7385.0 108027.5 7455.0 107712.5 ;
      RECT  7420.0 108062.5 7800.0 107992.5 ;
      RECT  7765.0 108417.5 7835.0 108027.5 ;
      RECT  7385.0 107712.5 7455.0 107577.5 ;
      RECT  7765.0 107712.5 7835.0 107577.5 ;
      RECT  7765.0 108552.5 7835.0 108417.5 ;
      RECT  7765.0 108095.0 7835.0 107960.0 ;
      RECT  7765.0 109012.5 7835.0 109717.5 ;
      RECT  7385.0 109367.5 7455.0 109437.5 ;
      RECT  7765.0 109367.5 7835.0 109437.5 ;
      RECT  7385.0 109402.5 7455.0 109717.5 ;
      RECT  7420.0 109367.5 7800.0 109437.5 ;
      RECT  7765.0 109012.5 7835.0 109402.5 ;
      RECT  7385.0 109717.5 7455.0 109852.5 ;
      RECT  7765.0 109717.5 7835.0 109852.5 ;
      RECT  7765.0 108877.5 7835.0 109012.5 ;
      RECT  7765.0 109335.0 7835.0 109470.0 ;
      RECT  7765.0 111107.5 7835.0 110402.5 ;
      RECT  7385.0 110752.5 7455.0 110682.5 ;
      RECT  7765.0 110752.5 7835.0 110682.5 ;
      RECT  7385.0 110717.5 7455.0 110402.5 ;
      RECT  7420.0 110752.5 7800.0 110682.5 ;
      RECT  7765.0 111107.5 7835.0 110717.5 ;
      RECT  7385.0 110402.5 7455.0 110267.5 ;
      RECT  7765.0 110402.5 7835.0 110267.5 ;
      RECT  7765.0 111242.5 7835.0 111107.5 ;
      RECT  7765.0 110785.0 7835.0 110650.0 ;
      RECT  7765.0 111702.5 7835.0 112407.5 ;
      RECT  7385.0 112057.5 7455.0 112127.5 ;
      RECT  7765.0 112057.5 7835.0 112127.5 ;
      RECT  7385.0 112092.5 7455.0 112407.5 ;
      RECT  7420.0 112057.5 7800.0 112127.5 ;
      RECT  7765.0 111702.5 7835.0 112092.5 ;
      RECT  7385.0 112407.5 7455.0 112542.5 ;
      RECT  7765.0 112407.5 7835.0 112542.5 ;
      RECT  7765.0 111567.5 7835.0 111702.5 ;
      RECT  7765.0 112025.0 7835.0 112160.0 ;
      RECT  7765.0 113797.5 7835.0 113092.5 ;
      RECT  7385.0 113442.5 7455.0 113372.5 ;
      RECT  7765.0 113442.5 7835.0 113372.5 ;
      RECT  7385.0 113407.5 7455.0 113092.5 ;
      RECT  7420.0 113442.5 7800.0 113372.5 ;
      RECT  7765.0 113797.5 7835.0 113407.5 ;
      RECT  7385.0 113092.5 7455.0 112957.5 ;
      RECT  7765.0 113092.5 7835.0 112957.5 ;
      RECT  7765.0 113932.5 7835.0 113797.5 ;
      RECT  7765.0 113475.0 7835.0 113340.0 ;
      RECT  5132.5 12467.5 4997.5 12537.5 ;
      RECT  5307.5 13902.5 5172.5 13972.5 ;
      RECT  5482.5 15157.5 5347.5 15227.5 ;
      RECT  5657.5 16592.5 5522.5 16662.5 ;
      RECT  5832.5 17847.5 5697.5 17917.5 ;
      RECT  6007.5 19282.5 5872.5 19352.5 ;
      RECT  6182.5 20537.5 6047.5 20607.5 ;
      RECT  6357.5 21972.5 6222.5 22042.5 ;
      RECT  6532.5 23227.5 6397.5 23297.5 ;
      RECT  6707.5 24662.5 6572.5 24732.5 ;
      RECT  6882.5 25917.5 6747.5 25987.5 ;
      RECT  7057.5 27352.5 6922.5 27422.5 ;
      RECT  5132.5 28667.5 4997.5 28737.5 ;
      RECT  5832.5 28527.5 5697.5 28597.5 ;
      RECT  6532.5 28387.5 6397.5 28457.5 ;
      RECT  5132.5 29982.5 4997.5 30052.5 ;
      RECT  5832.5 30122.5 5697.5 30192.5 ;
      RECT  6707.5 30262.5 6572.5 30332.5 ;
      RECT  5132.5 31357.5 4997.5 31427.5 ;
      RECT  5832.5 31217.5 5697.5 31287.5 ;
      RECT  6882.5 31077.5 6747.5 31147.5 ;
      RECT  5132.5 32672.5 4997.5 32742.5 ;
      RECT  5832.5 32812.5 5697.5 32882.5 ;
      RECT  7057.5 32952.5 6922.5 33022.5 ;
      RECT  5132.5 34047.5 4997.5 34117.5 ;
      RECT  6007.5 33907.5 5872.5 33977.5 ;
      RECT  6532.5 33767.5 6397.5 33837.5 ;
      RECT  5132.5 35362.5 4997.5 35432.5 ;
      RECT  6007.5 35502.5 5872.5 35572.5 ;
      RECT  6707.5 35642.5 6572.5 35712.5 ;
      RECT  5132.5 36737.5 4997.5 36807.5 ;
      RECT  6007.5 36597.5 5872.5 36667.5 ;
      RECT  6882.5 36457.5 6747.5 36527.5 ;
      RECT  5132.5 38052.5 4997.5 38122.5 ;
      RECT  6007.5 38192.5 5872.5 38262.5 ;
      RECT  7057.5 38332.5 6922.5 38402.5 ;
      RECT  5132.5 39427.5 4997.5 39497.5 ;
      RECT  6182.5 39287.5 6047.5 39357.5 ;
      RECT  6532.5 39147.5 6397.5 39217.5 ;
      RECT  5132.5 40742.5 4997.5 40812.5 ;
      RECT  6182.5 40882.5 6047.5 40952.5 ;
      RECT  6707.5 41022.5 6572.5 41092.5 ;
      RECT  5132.5 42117.5 4997.5 42187.5 ;
      RECT  6182.5 41977.5 6047.5 42047.5 ;
      RECT  6882.5 41837.5 6747.5 41907.5 ;
      RECT  5132.5 43432.5 4997.5 43502.5 ;
      RECT  6182.5 43572.5 6047.5 43642.5 ;
      RECT  7057.5 43712.5 6922.5 43782.5 ;
      RECT  5132.5 44807.5 4997.5 44877.5 ;
      RECT  6357.5 44667.5 6222.5 44737.5 ;
      RECT  6532.5 44527.5 6397.5 44597.5 ;
      RECT  5132.5 46122.5 4997.5 46192.5 ;
      RECT  6357.5 46262.5 6222.5 46332.5 ;
      RECT  6707.5 46402.5 6572.5 46472.5 ;
      RECT  5132.5 47497.5 4997.5 47567.5 ;
      RECT  6357.5 47357.5 6222.5 47427.5 ;
      RECT  6882.5 47217.5 6747.5 47287.5 ;
      RECT  5132.5 48812.5 4997.5 48882.5 ;
      RECT  6357.5 48952.5 6222.5 49022.5 ;
      RECT  7057.5 49092.5 6922.5 49162.5 ;
      RECT  5307.5 50187.5 5172.5 50257.5 ;
      RECT  5832.5 50047.5 5697.5 50117.5 ;
      RECT  6532.5 49907.5 6397.5 49977.5 ;
      RECT  5307.5 51502.5 5172.5 51572.5 ;
      RECT  5832.5 51642.5 5697.5 51712.5 ;
      RECT  6707.5 51782.5 6572.5 51852.5 ;
      RECT  5307.5 52877.5 5172.5 52947.5 ;
      RECT  5832.5 52737.5 5697.5 52807.5 ;
      RECT  6882.5 52597.5 6747.5 52667.5 ;
      RECT  5307.5 54192.5 5172.5 54262.5 ;
      RECT  5832.5 54332.5 5697.5 54402.5 ;
      RECT  7057.5 54472.5 6922.5 54542.5 ;
      RECT  5307.5 55567.5 5172.5 55637.5 ;
      RECT  6007.5 55427.5 5872.5 55497.5 ;
      RECT  6532.5 55287.5 6397.5 55357.5 ;
      RECT  5307.5 56882.5 5172.5 56952.5 ;
      RECT  6007.5 57022.5 5872.5 57092.5 ;
      RECT  6707.5 57162.5 6572.5 57232.5 ;
      RECT  5307.5 58257.5 5172.5 58327.5 ;
      RECT  6007.5 58117.5 5872.5 58187.5 ;
      RECT  6882.5 57977.5 6747.5 58047.5 ;
      RECT  5307.5 59572.5 5172.5 59642.5 ;
      RECT  6007.5 59712.5 5872.5 59782.5 ;
      RECT  7057.5 59852.5 6922.5 59922.5 ;
      RECT  5307.5 60947.5 5172.5 61017.5 ;
      RECT  6182.5 60807.5 6047.5 60877.5 ;
      RECT  6532.5 60667.5 6397.5 60737.5 ;
      RECT  5307.5 62262.5 5172.5 62332.5 ;
      RECT  6182.5 62402.5 6047.5 62472.5 ;
      RECT  6707.5 62542.5 6572.5 62612.5 ;
      RECT  5307.5 63637.5 5172.5 63707.5 ;
      RECT  6182.5 63497.5 6047.5 63567.5 ;
      RECT  6882.5 63357.5 6747.5 63427.5 ;
      RECT  5307.5 64952.5 5172.5 65022.5 ;
      RECT  6182.5 65092.5 6047.5 65162.5 ;
      RECT  7057.5 65232.5 6922.5 65302.5 ;
      RECT  5307.5 66327.5 5172.5 66397.5 ;
      RECT  6357.5 66187.5 6222.5 66257.5 ;
      RECT  6532.5 66047.5 6397.5 66117.5 ;
      RECT  5307.5 67642.5 5172.5 67712.5 ;
      RECT  6357.5 67782.5 6222.5 67852.5 ;
      RECT  6707.5 67922.5 6572.5 67992.5 ;
      RECT  5307.5 69017.5 5172.5 69087.5 ;
      RECT  6357.5 68877.5 6222.5 68947.5 ;
      RECT  6882.5 68737.5 6747.5 68807.5 ;
      RECT  5307.5 70332.5 5172.5 70402.5 ;
      RECT  6357.5 70472.5 6222.5 70542.5 ;
      RECT  7057.5 70612.5 6922.5 70682.5 ;
      RECT  5482.5 71707.5 5347.5 71777.5 ;
      RECT  5832.5 71567.5 5697.5 71637.5 ;
      RECT  6532.5 71427.5 6397.5 71497.5 ;
      RECT  5482.5 73022.5 5347.5 73092.5 ;
      RECT  5832.5 73162.5 5697.5 73232.5 ;
      RECT  6707.5 73302.5 6572.5 73372.5 ;
      RECT  5482.5 74397.5 5347.5 74467.5 ;
      RECT  5832.5 74257.5 5697.5 74327.5 ;
      RECT  6882.5 74117.5 6747.5 74187.5 ;
      RECT  5482.5 75712.5 5347.5 75782.5 ;
      RECT  5832.5 75852.5 5697.5 75922.5 ;
      RECT  7057.5 75992.5 6922.5 76062.5 ;
      RECT  5482.5 77087.5 5347.5 77157.5 ;
      RECT  6007.5 76947.5 5872.5 77017.5 ;
      RECT  6532.5 76807.5 6397.5 76877.5 ;
      RECT  5482.5 78402.5 5347.5 78472.5 ;
      RECT  6007.5 78542.5 5872.5 78612.5 ;
      RECT  6707.5 78682.5 6572.5 78752.5 ;
      RECT  5482.5 79777.5 5347.5 79847.5 ;
      RECT  6007.5 79637.5 5872.5 79707.5 ;
      RECT  6882.5 79497.5 6747.5 79567.5 ;
      RECT  5482.5 81092.5 5347.5 81162.5 ;
      RECT  6007.5 81232.5 5872.5 81302.5 ;
      RECT  7057.5 81372.5 6922.5 81442.5 ;
      RECT  5482.5 82467.5 5347.5 82537.5 ;
      RECT  6182.5 82327.5 6047.5 82397.5 ;
      RECT  6532.5 82187.5 6397.5 82257.5 ;
      RECT  5482.5 83782.5 5347.5 83852.5 ;
      RECT  6182.5 83922.5 6047.5 83992.5 ;
      RECT  6707.5 84062.5 6572.5 84132.5 ;
      RECT  5482.5 85157.5 5347.5 85227.5 ;
      RECT  6182.5 85017.5 6047.5 85087.5 ;
      RECT  6882.5 84877.5 6747.5 84947.5 ;
      RECT  5482.5 86472.5 5347.5 86542.5 ;
      RECT  6182.5 86612.5 6047.5 86682.5 ;
      RECT  7057.5 86752.5 6922.5 86822.5 ;
      RECT  5482.5 87847.5 5347.5 87917.5 ;
      RECT  6357.5 87707.5 6222.5 87777.5 ;
      RECT  6532.5 87567.5 6397.5 87637.5 ;
      RECT  5482.5 89162.5 5347.5 89232.5 ;
      RECT  6357.5 89302.5 6222.5 89372.5 ;
      RECT  6707.5 89442.5 6572.5 89512.5 ;
      RECT  5482.5 90537.5 5347.5 90607.5 ;
      RECT  6357.5 90397.5 6222.5 90467.5 ;
      RECT  6882.5 90257.5 6747.5 90327.5 ;
      RECT  5482.5 91852.5 5347.5 91922.5 ;
      RECT  6357.5 91992.5 6222.5 92062.5 ;
      RECT  7057.5 92132.5 6922.5 92202.5 ;
      RECT  5657.5 93227.5 5522.5 93297.5 ;
      RECT  5832.5 93087.5 5697.5 93157.5 ;
      RECT  6532.5 92947.5 6397.5 93017.5 ;
      RECT  5657.5 94542.5 5522.5 94612.5 ;
      RECT  5832.5 94682.5 5697.5 94752.5 ;
      RECT  6707.5 94822.5 6572.5 94892.5 ;
      RECT  5657.5 95917.5 5522.5 95987.5 ;
      RECT  5832.5 95777.5 5697.5 95847.5 ;
      RECT  6882.5 95637.5 6747.5 95707.5 ;
      RECT  5657.5 97232.5 5522.5 97302.5 ;
      RECT  5832.5 97372.5 5697.5 97442.5 ;
      RECT  7057.5 97512.5 6922.5 97582.5 ;
      RECT  5657.5 98607.5 5522.5 98677.5 ;
      RECT  6007.5 98467.5 5872.5 98537.5 ;
      RECT  6532.5 98327.5 6397.5 98397.5 ;
      RECT  5657.5 99922.5 5522.5 99992.5 ;
      RECT  6007.5 100062.5 5872.5 100132.5 ;
      RECT  6707.5 100202.5 6572.5 100272.5 ;
      RECT  5657.5 101297.5 5522.5 101367.5 ;
      RECT  6007.5 101157.5 5872.5 101227.5 ;
      RECT  6882.5 101017.5 6747.5 101087.5 ;
      RECT  5657.5 102612.5 5522.5 102682.5 ;
      RECT  6007.5 102752.5 5872.5 102822.5 ;
      RECT  7057.5 102892.5 6922.5 102962.5 ;
      RECT  5657.5 103987.5 5522.5 104057.5 ;
      RECT  6182.5 103847.5 6047.5 103917.5 ;
      RECT  6532.5 103707.5 6397.5 103777.5 ;
      RECT  5657.5 105302.5 5522.5 105372.5 ;
      RECT  6182.5 105442.5 6047.5 105512.5 ;
      RECT  6707.5 105582.5 6572.5 105652.5 ;
      RECT  5657.5 106677.5 5522.5 106747.5 ;
      RECT  6182.5 106537.5 6047.5 106607.5 ;
      RECT  6882.5 106397.5 6747.5 106467.5 ;
      RECT  5657.5 107992.5 5522.5 108062.5 ;
      RECT  6182.5 108132.5 6047.5 108202.5 ;
      RECT  7057.5 108272.5 6922.5 108342.5 ;
      RECT  5657.5 109367.5 5522.5 109437.5 ;
      RECT  6357.5 109227.5 6222.5 109297.5 ;
      RECT  6532.5 109087.5 6397.5 109157.5 ;
      RECT  5657.5 110682.5 5522.5 110752.5 ;
      RECT  6357.5 110822.5 6222.5 110892.5 ;
      RECT  6707.5 110962.5 6572.5 111032.5 ;
      RECT  5657.5 112057.5 5522.5 112127.5 ;
      RECT  6357.5 111917.5 6222.5 111987.5 ;
      RECT  6882.5 111777.5 6747.5 111847.5 ;
      RECT  5657.5 113372.5 5522.5 113442.5 ;
      RECT  6357.5 113512.5 6222.5 113582.5 ;
      RECT  7057.5 113652.5 6922.5 113722.5 ;
      RECT  11025.0 11875.0 11095.0 17115.0 ;
      RECT  10750.0 11875.0 10820.0 17115.0 ;
      RECT  11025.0 17255.0 11095.0 22495.0 ;
      RECT  10750.0 17255.0 10820.0 22495.0 ;
      RECT  11025.0 22635.0 11095.0 27875.0 ;
      RECT  10750.0 22635.0 10820.0 27875.0 ;
      RECT  9035.0 28405.0 9105.0 28475.0 ;
      RECT  9035.0 28370.0 9105.0 28440.0 ;
      RECT  9070.0 28405.0 10032.5 28475.0 ;
      RECT  9035.0 30245.0 9105.0 30315.0 ;
      RECT  9035.0 30280.0 9105.0 30350.0 ;
      RECT  9070.0 30245.0 10032.5 30315.0 ;
      RECT  9035.0 31095.0 9105.0 31165.0 ;
      RECT  9035.0 31060.0 9105.0 31130.0 ;
      RECT  9070.0 31095.0 10032.5 31165.0 ;
      RECT  9035.0 32935.0 9105.0 33005.0 ;
      RECT  9035.0 32970.0 9105.0 33040.0 ;
      RECT  9070.0 32935.0 10032.5 33005.0 ;
      RECT  9035.0 33785.0 9105.0 33855.0 ;
      RECT  9035.0 33750.0 9105.0 33820.0 ;
      RECT  9070.0 33785.0 10032.5 33855.0 ;
      RECT  9035.0 35625.0 9105.0 35695.0 ;
      RECT  9035.0 35660.0 9105.0 35730.0 ;
      RECT  9070.0 35625.0 10032.5 35695.0 ;
      RECT  9035.0 36475.0 9105.0 36545.0 ;
      RECT  9035.0 36440.0 9105.0 36510.0 ;
      RECT  9070.0 36475.0 10032.5 36545.0 ;
      RECT  9035.0 38315.0 9105.0 38385.0 ;
      RECT  9035.0 38350.0 9105.0 38420.0 ;
      RECT  9070.0 38315.0 10032.5 38385.0 ;
      RECT  9035.0 39165.0 9105.0 39235.0 ;
      RECT  9035.0 39130.0 9105.0 39200.0 ;
      RECT  9070.0 39165.0 10032.5 39235.0 ;
      RECT  9035.0 41005.0 9105.0 41075.0 ;
      RECT  9035.0 41040.0 9105.0 41110.0 ;
      RECT  9070.0 41005.0 10032.5 41075.0 ;
      RECT  9035.0 41855.0 9105.0 41925.0 ;
      RECT  9035.0 41820.0 9105.0 41890.0 ;
      RECT  9070.0 41855.0 10032.5 41925.0 ;
      RECT  9035.0 43695.0 9105.0 43765.0 ;
      RECT  9035.0 43730.0 9105.0 43800.0 ;
      RECT  9070.0 43695.0 10032.5 43765.0 ;
      RECT  9035.0 44545.0 9105.0 44615.0 ;
      RECT  9035.0 44510.0 9105.0 44580.0 ;
      RECT  9070.0 44545.0 10032.5 44615.0 ;
      RECT  9035.0 46385.0 9105.0 46455.0 ;
      RECT  9035.0 46420.0 9105.0 46490.0 ;
      RECT  9070.0 46385.0 10032.5 46455.0 ;
      RECT  9035.0 47235.0 9105.0 47305.0 ;
      RECT  9035.0 47200.0 9105.0 47270.0 ;
      RECT  9070.0 47235.0 10032.5 47305.0 ;
      RECT  9035.0 49075.0 9105.0 49145.0 ;
      RECT  9035.0 49110.0 9105.0 49180.0 ;
      RECT  9070.0 49075.0 10032.5 49145.0 ;
      RECT  9035.0 49925.0 9105.0 49995.0 ;
      RECT  9035.0 49890.0 9105.0 49960.0 ;
      RECT  9070.0 49925.0 10032.5 49995.0 ;
      RECT  9035.0 51765.0 9105.0 51835.0 ;
      RECT  9035.0 51800.0 9105.0 51870.0 ;
      RECT  9070.0 51765.0 10032.5 51835.0 ;
      RECT  9035.0 52615.0 9105.0 52685.0 ;
      RECT  9035.0 52580.0 9105.0 52650.0 ;
      RECT  9070.0 52615.0 10032.5 52685.0 ;
      RECT  9035.0 54455.0 9105.0 54525.0 ;
      RECT  9035.0 54490.0 9105.0 54560.0 ;
      RECT  9070.0 54455.0 10032.5 54525.0 ;
      RECT  9035.0 55305.0 9105.0 55375.0 ;
      RECT  9035.0 55270.0 9105.0 55340.0 ;
      RECT  9070.0 55305.0 10032.5 55375.0 ;
      RECT  9035.0 57145.0 9105.0 57215.0 ;
      RECT  9035.0 57180.0 9105.0 57250.0 ;
      RECT  9070.0 57145.0 10032.5 57215.0 ;
      RECT  9035.0 57995.0 9105.0 58065.0 ;
      RECT  9035.0 57960.0 9105.0 58030.0 ;
      RECT  9070.0 57995.0 10032.5 58065.0 ;
      RECT  9035.0 59835.0 9105.0 59905.0 ;
      RECT  9035.0 59870.0 9105.0 59940.0 ;
      RECT  9070.0 59835.0 10032.5 59905.0 ;
      RECT  9035.0 60685.0 9105.0 60755.0 ;
      RECT  9035.0 60650.0 9105.0 60720.0 ;
      RECT  9070.0 60685.0 10032.5 60755.0 ;
      RECT  9035.0 62525.0 9105.0 62595.0 ;
      RECT  9035.0 62560.0 9105.0 62630.0 ;
      RECT  9070.0 62525.0 10032.5 62595.0 ;
      RECT  9035.0 63375.0 9105.0 63445.0 ;
      RECT  9035.0 63340.0 9105.0 63410.0 ;
      RECT  9070.0 63375.0 10032.5 63445.0 ;
      RECT  9035.0 65215.0 9105.0 65285.0 ;
      RECT  9035.0 65250.0 9105.0 65320.0 ;
      RECT  9070.0 65215.0 10032.5 65285.0 ;
      RECT  9035.0 66065.0 9105.0 66135.0 ;
      RECT  9035.0 66030.0 9105.0 66100.0 ;
      RECT  9070.0 66065.0 10032.5 66135.0 ;
      RECT  9035.0 67905.0 9105.0 67975.0 ;
      RECT  9035.0 67940.0 9105.0 68010.0 ;
      RECT  9070.0 67905.0 10032.5 67975.0 ;
      RECT  9035.0 68755.0 9105.0 68825.0 ;
      RECT  9035.0 68720.0 9105.0 68790.0 ;
      RECT  9070.0 68755.0 10032.5 68825.0 ;
      RECT  9035.0 70595.0 9105.0 70665.0 ;
      RECT  9035.0 70630.0 9105.0 70700.0 ;
      RECT  9070.0 70595.0 10032.5 70665.0 ;
      RECT  9035.0 71445.0 9105.0 71515.0 ;
      RECT  9035.0 71410.0 9105.0 71480.0 ;
      RECT  9070.0 71445.0 10032.5 71515.0 ;
      RECT  9035.0 73285.0 9105.0 73355.0 ;
      RECT  9035.0 73320.0 9105.0 73390.0 ;
      RECT  9070.0 73285.0 10032.5 73355.0 ;
      RECT  9035.0 74135.0 9105.0 74205.0 ;
      RECT  9035.0 74100.0 9105.0 74170.0 ;
      RECT  9070.0 74135.0 10032.5 74205.0 ;
      RECT  9035.0 75975.0 9105.0 76045.0 ;
      RECT  9035.0 76010.0 9105.0 76080.0 ;
      RECT  9070.0 75975.0 10032.5 76045.0 ;
      RECT  9035.0 76825.0 9105.0 76895.0 ;
      RECT  9035.0 76790.0 9105.0 76860.0 ;
      RECT  9070.0 76825.0 10032.5 76895.0 ;
      RECT  9035.0 78665.0 9105.0 78735.0 ;
      RECT  9035.0 78700.0 9105.0 78770.0 ;
      RECT  9070.0 78665.0 10032.5 78735.0 ;
      RECT  9035.0 79515.0 9105.0 79585.0 ;
      RECT  9035.0 79480.0 9105.0 79550.0 ;
      RECT  9070.0 79515.0 10032.5 79585.0 ;
      RECT  9035.0 81355.0 9105.0 81425.0 ;
      RECT  9035.0 81390.0 9105.0 81460.0 ;
      RECT  9070.0 81355.0 10032.5 81425.0 ;
      RECT  9035.0 82205.0 9105.0 82275.0 ;
      RECT  9035.0 82170.0 9105.0 82240.0 ;
      RECT  9070.0 82205.0 10032.5 82275.0 ;
      RECT  9035.0 84045.0 9105.0 84115.0 ;
      RECT  9035.0 84080.0 9105.0 84150.0 ;
      RECT  9070.0 84045.0 10032.5 84115.0 ;
      RECT  9035.0 84895.0 9105.0 84965.0 ;
      RECT  9035.0 84860.0 9105.0 84930.0 ;
      RECT  9070.0 84895.0 10032.5 84965.0 ;
      RECT  9035.0 86735.0 9105.0 86805.0 ;
      RECT  9035.0 86770.0 9105.0 86840.0 ;
      RECT  9070.0 86735.0 10032.5 86805.0 ;
      RECT  9035.0 87585.0 9105.0 87655.0 ;
      RECT  9035.0 87550.0 9105.0 87620.0 ;
      RECT  9070.0 87585.0 10032.5 87655.0 ;
      RECT  9035.0 89425.0 9105.0 89495.0 ;
      RECT  9035.0 89460.0 9105.0 89530.0 ;
      RECT  9070.0 89425.0 10032.5 89495.0 ;
      RECT  9035.0 90275.0 9105.0 90345.0 ;
      RECT  9035.0 90240.0 9105.0 90310.0 ;
      RECT  9070.0 90275.0 10032.5 90345.0 ;
      RECT  9035.0 92115.0 9105.0 92185.0 ;
      RECT  9035.0 92150.0 9105.0 92220.0 ;
      RECT  9070.0 92115.0 10032.5 92185.0 ;
      RECT  9035.0 92965.0 9105.0 93035.0 ;
      RECT  9035.0 92930.0 9105.0 93000.0 ;
      RECT  9070.0 92965.0 10032.5 93035.0 ;
      RECT  9035.0 94805.0 9105.0 94875.0 ;
      RECT  9035.0 94840.0 9105.0 94910.0 ;
      RECT  9070.0 94805.0 10032.5 94875.0 ;
      RECT  9035.0 95655.0 9105.0 95725.0 ;
      RECT  9035.0 95620.0 9105.0 95690.0 ;
      RECT  9070.0 95655.0 10032.5 95725.0 ;
      RECT  9035.0 97495.0 9105.0 97565.0 ;
      RECT  9035.0 97530.0 9105.0 97600.0 ;
      RECT  9070.0 97495.0 10032.5 97565.0 ;
      RECT  9035.0 98345.0 9105.0 98415.0 ;
      RECT  9035.0 98310.0 9105.0 98380.0 ;
      RECT  9070.0 98345.0 10032.5 98415.0 ;
      RECT  9035.0 100185.0 9105.0 100255.0 ;
      RECT  9035.0 100220.0 9105.0 100290.0 ;
      RECT  9070.0 100185.0 10032.5 100255.0 ;
      RECT  9035.0 101035.0 9105.0 101105.0 ;
      RECT  9035.0 101000.0 9105.0 101070.0 ;
      RECT  9070.0 101035.0 10032.5 101105.0 ;
      RECT  9035.0 102875.0 9105.0 102945.0 ;
      RECT  9035.0 102910.0 9105.0 102980.0 ;
      RECT  9070.0 102875.0 10032.5 102945.0 ;
      RECT  9035.0 103725.0 9105.0 103795.0 ;
      RECT  9035.0 103690.0 9105.0 103760.0 ;
      RECT  9070.0 103725.0 10032.5 103795.0 ;
      RECT  9035.0 105565.0 9105.0 105635.0 ;
      RECT  9035.0 105600.0 9105.0 105670.0 ;
      RECT  9070.0 105565.0 10032.5 105635.0 ;
      RECT  9035.0 106415.0 9105.0 106485.0 ;
      RECT  9035.0 106380.0 9105.0 106450.0 ;
      RECT  9070.0 106415.0 10032.5 106485.0 ;
      RECT  9035.0 108255.0 9105.0 108325.0 ;
      RECT  9035.0 108290.0 9105.0 108360.0 ;
      RECT  9070.0 108255.0 10032.5 108325.0 ;
      RECT  9035.0 109105.0 9105.0 109175.0 ;
      RECT  9035.0 109070.0 9105.0 109140.0 ;
      RECT  9070.0 109105.0 10032.5 109175.0 ;
      RECT  9035.0 110945.0 9105.0 111015.0 ;
      RECT  9035.0 110980.0 9105.0 111050.0 ;
      RECT  9070.0 110945.0 10032.5 111015.0 ;
      RECT  9035.0 111795.0 9105.0 111865.0 ;
      RECT  9035.0 111760.0 9105.0 111830.0 ;
      RECT  9070.0 111795.0 10032.5 111865.0 ;
      RECT  9035.0 113635.0 9105.0 113705.0 ;
      RECT  9035.0 113670.0 9105.0 113740.0 ;
      RECT  9070.0 113635.0 10032.5 113705.0 ;
      RECT  9970.0 28620.0 10040.0 28690.0 ;
      RECT  10160.0 28620.0 10230.0 28690.0 ;
      RECT  9970.0 28655.0 10040.0 29017.5 ;
      RECT  10005.0 28620.0 10195.0 28690.0 ;
      RECT  10160.0 28312.5 10230.0 28655.0 ;
      RECT  9970.0 29017.5 10040.0 29152.5 ;
      RECT  10160.0 28177.5 10230.0 28312.5 ;
      RECT  10262.5 28620.0 10127.5 28690.0 ;
      RECT  8895.0 28575.0 8965.0 28710.0 ;
      RECT  9035.0 28302.5 9105.0 28437.5 ;
      RECT  10032.5 28405.0 9897.5 28475.0 ;
      RECT  9970.0 30100.0 10040.0 30030.0 ;
      RECT  10160.0 30100.0 10230.0 30030.0 ;
      RECT  9970.0 30065.0 10040.0 29702.5 ;
      RECT  10005.0 30100.0 10195.0 30030.0 ;
      RECT  10160.0 30407.5 10230.0 30065.0 ;
      RECT  9970.0 29702.5 10040.0 29567.5 ;
      RECT  10160.0 30542.5 10230.0 30407.5 ;
      RECT  10262.5 30100.0 10127.5 30030.0 ;
      RECT  8895.0 30010.0 8965.0 30145.0 ;
      RECT  9035.0 30282.5 9105.0 30417.5 ;
      RECT  10032.5 30245.0 9897.5 30315.0 ;
      RECT  9970.0 31310.0 10040.0 31380.0 ;
      RECT  10160.0 31310.0 10230.0 31380.0 ;
      RECT  9970.0 31345.0 10040.0 31707.5 ;
      RECT  10005.0 31310.0 10195.0 31380.0 ;
      RECT  10160.0 31002.5 10230.0 31345.0 ;
      RECT  9970.0 31707.5 10040.0 31842.5 ;
      RECT  10160.0 30867.5 10230.0 31002.5 ;
      RECT  10262.5 31310.0 10127.5 31380.0 ;
      RECT  8895.0 31265.0 8965.0 31400.0 ;
      RECT  9035.0 30992.5 9105.0 31127.5 ;
      RECT  10032.5 31095.0 9897.5 31165.0 ;
      RECT  9970.0 32790.0 10040.0 32720.0 ;
      RECT  10160.0 32790.0 10230.0 32720.0 ;
      RECT  9970.0 32755.0 10040.0 32392.5 ;
      RECT  10005.0 32790.0 10195.0 32720.0 ;
      RECT  10160.0 33097.5 10230.0 32755.0 ;
      RECT  9970.0 32392.5 10040.0 32257.5 ;
      RECT  10160.0 33232.5 10230.0 33097.5 ;
      RECT  10262.5 32790.0 10127.5 32720.0 ;
      RECT  8895.0 32700.0 8965.0 32835.0 ;
      RECT  9035.0 32972.5 9105.0 33107.5 ;
      RECT  10032.5 32935.0 9897.5 33005.0 ;
      RECT  9970.0 34000.0 10040.0 34070.0 ;
      RECT  10160.0 34000.0 10230.0 34070.0 ;
      RECT  9970.0 34035.0 10040.0 34397.5 ;
      RECT  10005.0 34000.0 10195.0 34070.0 ;
      RECT  10160.0 33692.5 10230.0 34035.0 ;
      RECT  9970.0 34397.5 10040.0 34532.5 ;
      RECT  10160.0 33557.5 10230.0 33692.5 ;
      RECT  10262.5 34000.0 10127.5 34070.0 ;
      RECT  8895.0 33955.0 8965.0 34090.0 ;
      RECT  9035.0 33682.5 9105.0 33817.5 ;
      RECT  10032.5 33785.0 9897.5 33855.0 ;
      RECT  9970.0 35480.0 10040.0 35410.0 ;
      RECT  10160.0 35480.0 10230.0 35410.0 ;
      RECT  9970.0 35445.0 10040.0 35082.5 ;
      RECT  10005.0 35480.0 10195.0 35410.0 ;
      RECT  10160.0 35787.5 10230.0 35445.0 ;
      RECT  9970.0 35082.5 10040.0 34947.5 ;
      RECT  10160.0 35922.5 10230.0 35787.5 ;
      RECT  10262.5 35480.0 10127.5 35410.0 ;
      RECT  8895.0 35390.0 8965.0 35525.0 ;
      RECT  9035.0 35662.5 9105.0 35797.5 ;
      RECT  10032.5 35625.0 9897.5 35695.0 ;
      RECT  9970.0 36690.0 10040.0 36760.0 ;
      RECT  10160.0 36690.0 10230.0 36760.0 ;
      RECT  9970.0 36725.0 10040.0 37087.5 ;
      RECT  10005.0 36690.0 10195.0 36760.0 ;
      RECT  10160.0 36382.5 10230.0 36725.0 ;
      RECT  9970.0 37087.5 10040.0 37222.5 ;
      RECT  10160.0 36247.5 10230.0 36382.5 ;
      RECT  10262.5 36690.0 10127.5 36760.0 ;
      RECT  8895.0 36645.0 8965.0 36780.0 ;
      RECT  9035.0 36372.5 9105.0 36507.5 ;
      RECT  10032.5 36475.0 9897.5 36545.0 ;
      RECT  9970.0 38170.0 10040.0 38100.0 ;
      RECT  10160.0 38170.0 10230.0 38100.0 ;
      RECT  9970.0 38135.0 10040.0 37772.5 ;
      RECT  10005.0 38170.0 10195.0 38100.0 ;
      RECT  10160.0 38477.5 10230.0 38135.0 ;
      RECT  9970.0 37772.5 10040.0 37637.5 ;
      RECT  10160.0 38612.5 10230.0 38477.5 ;
      RECT  10262.5 38170.0 10127.5 38100.0 ;
      RECT  8895.0 38080.0 8965.0 38215.0 ;
      RECT  9035.0 38352.5 9105.0 38487.5 ;
      RECT  10032.5 38315.0 9897.5 38385.0 ;
      RECT  9970.0 39380.0 10040.0 39450.0 ;
      RECT  10160.0 39380.0 10230.0 39450.0 ;
      RECT  9970.0 39415.0 10040.0 39777.5 ;
      RECT  10005.0 39380.0 10195.0 39450.0 ;
      RECT  10160.0 39072.5 10230.0 39415.0 ;
      RECT  9970.0 39777.5 10040.0 39912.5 ;
      RECT  10160.0 38937.5 10230.0 39072.5 ;
      RECT  10262.5 39380.0 10127.5 39450.0 ;
      RECT  8895.0 39335.0 8965.0 39470.0 ;
      RECT  9035.0 39062.5 9105.0 39197.5 ;
      RECT  10032.5 39165.0 9897.5 39235.0 ;
      RECT  9970.0 40860.0 10040.0 40790.0 ;
      RECT  10160.0 40860.0 10230.0 40790.0 ;
      RECT  9970.0 40825.0 10040.0 40462.5 ;
      RECT  10005.0 40860.0 10195.0 40790.0 ;
      RECT  10160.0 41167.5 10230.0 40825.0 ;
      RECT  9970.0 40462.5 10040.0 40327.5 ;
      RECT  10160.0 41302.5 10230.0 41167.5 ;
      RECT  10262.5 40860.0 10127.5 40790.0 ;
      RECT  8895.0 40770.0 8965.0 40905.0 ;
      RECT  9035.0 41042.5 9105.0 41177.5 ;
      RECT  10032.5 41005.0 9897.5 41075.0 ;
      RECT  9970.0 42070.0 10040.0 42140.0 ;
      RECT  10160.0 42070.0 10230.0 42140.0 ;
      RECT  9970.0 42105.0 10040.0 42467.5 ;
      RECT  10005.0 42070.0 10195.0 42140.0 ;
      RECT  10160.0 41762.5 10230.0 42105.0 ;
      RECT  9970.0 42467.5 10040.0 42602.5 ;
      RECT  10160.0 41627.5 10230.0 41762.5 ;
      RECT  10262.5 42070.0 10127.5 42140.0 ;
      RECT  8895.0 42025.0 8965.0 42160.0 ;
      RECT  9035.0 41752.5 9105.0 41887.5 ;
      RECT  10032.5 41855.0 9897.5 41925.0 ;
      RECT  9970.0 43550.0 10040.0 43480.0 ;
      RECT  10160.0 43550.0 10230.0 43480.0 ;
      RECT  9970.0 43515.0 10040.0 43152.5 ;
      RECT  10005.0 43550.0 10195.0 43480.0 ;
      RECT  10160.0 43857.5 10230.0 43515.0 ;
      RECT  9970.0 43152.5 10040.0 43017.5 ;
      RECT  10160.0 43992.5 10230.0 43857.5 ;
      RECT  10262.5 43550.0 10127.5 43480.0 ;
      RECT  8895.0 43460.0 8965.0 43595.0 ;
      RECT  9035.0 43732.5 9105.0 43867.5 ;
      RECT  10032.5 43695.0 9897.5 43765.0 ;
      RECT  9970.0 44760.0 10040.0 44830.0 ;
      RECT  10160.0 44760.0 10230.0 44830.0 ;
      RECT  9970.0 44795.0 10040.0 45157.5 ;
      RECT  10005.0 44760.0 10195.0 44830.0 ;
      RECT  10160.0 44452.5 10230.0 44795.0 ;
      RECT  9970.0 45157.5 10040.0 45292.5 ;
      RECT  10160.0 44317.5 10230.0 44452.5 ;
      RECT  10262.5 44760.0 10127.5 44830.0 ;
      RECT  8895.0 44715.0 8965.0 44850.0 ;
      RECT  9035.0 44442.5 9105.0 44577.5 ;
      RECT  10032.5 44545.0 9897.5 44615.0 ;
      RECT  9970.0 46240.0 10040.0 46170.0 ;
      RECT  10160.0 46240.0 10230.0 46170.0 ;
      RECT  9970.0 46205.0 10040.0 45842.5 ;
      RECT  10005.0 46240.0 10195.0 46170.0 ;
      RECT  10160.0 46547.5 10230.0 46205.0 ;
      RECT  9970.0 45842.5 10040.0 45707.5 ;
      RECT  10160.0 46682.5 10230.0 46547.5 ;
      RECT  10262.5 46240.0 10127.5 46170.0 ;
      RECT  8895.0 46150.0 8965.0 46285.0 ;
      RECT  9035.0 46422.5 9105.0 46557.5 ;
      RECT  10032.5 46385.0 9897.5 46455.0 ;
      RECT  9970.0 47450.0 10040.0 47520.0 ;
      RECT  10160.0 47450.0 10230.0 47520.0 ;
      RECT  9970.0 47485.0 10040.0 47847.5 ;
      RECT  10005.0 47450.0 10195.0 47520.0 ;
      RECT  10160.0 47142.5 10230.0 47485.0 ;
      RECT  9970.0 47847.5 10040.0 47982.5 ;
      RECT  10160.0 47007.5 10230.0 47142.5 ;
      RECT  10262.5 47450.0 10127.5 47520.0 ;
      RECT  8895.0 47405.0 8965.0 47540.0 ;
      RECT  9035.0 47132.5 9105.0 47267.5 ;
      RECT  10032.5 47235.0 9897.5 47305.0 ;
      RECT  9970.0 48930.0 10040.0 48860.0 ;
      RECT  10160.0 48930.0 10230.0 48860.0 ;
      RECT  9970.0 48895.0 10040.0 48532.5 ;
      RECT  10005.0 48930.0 10195.0 48860.0 ;
      RECT  10160.0 49237.5 10230.0 48895.0 ;
      RECT  9970.0 48532.5 10040.0 48397.5 ;
      RECT  10160.0 49372.5 10230.0 49237.5 ;
      RECT  10262.5 48930.0 10127.5 48860.0 ;
      RECT  8895.0 48840.0 8965.0 48975.0 ;
      RECT  9035.0 49112.5 9105.0 49247.5 ;
      RECT  10032.5 49075.0 9897.5 49145.0 ;
      RECT  9970.0 50140.0 10040.0 50210.0 ;
      RECT  10160.0 50140.0 10230.0 50210.0 ;
      RECT  9970.0 50175.0 10040.0 50537.5 ;
      RECT  10005.0 50140.0 10195.0 50210.0 ;
      RECT  10160.0 49832.5 10230.0 50175.0 ;
      RECT  9970.0 50537.5 10040.0 50672.5 ;
      RECT  10160.0 49697.5 10230.0 49832.5 ;
      RECT  10262.5 50140.0 10127.5 50210.0 ;
      RECT  8895.0 50095.0 8965.0 50230.0 ;
      RECT  9035.0 49822.5 9105.0 49957.5 ;
      RECT  10032.5 49925.0 9897.5 49995.0 ;
      RECT  9970.0 51620.0 10040.0 51550.0 ;
      RECT  10160.0 51620.0 10230.0 51550.0 ;
      RECT  9970.0 51585.0 10040.0 51222.5 ;
      RECT  10005.0 51620.0 10195.0 51550.0 ;
      RECT  10160.0 51927.5 10230.0 51585.0 ;
      RECT  9970.0 51222.5 10040.0 51087.5 ;
      RECT  10160.0 52062.5 10230.0 51927.5 ;
      RECT  10262.5 51620.0 10127.5 51550.0 ;
      RECT  8895.0 51530.0 8965.0 51665.0 ;
      RECT  9035.0 51802.5 9105.0 51937.5 ;
      RECT  10032.5 51765.0 9897.5 51835.0 ;
      RECT  9970.0 52830.0 10040.0 52900.0 ;
      RECT  10160.0 52830.0 10230.0 52900.0 ;
      RECT  9970.0 52865.0 10040.0 53227.5 ;
      RECT  10005.0 52830.0 10195.0 52900.0 ;
      RECT  10160.0 52522.5 10230.0 52865.0 ;
      RECT  9970.0 53227.5 10040.0 53362.5 ;
      RECT  10160.0 52387.5 10230.0 52522.5 ;
      RECT  10262.5 52830.0 10127.5 52900.0 ;
      RECT  8895.0 52785.0 8965.0 52920.0 ;
      RECT  9035.0 52512.5 9105.0 52647.5 ;
      RECT  10032.5 52615.0 9897.5 52685.0 ;
      RECT  9970.0 54310.0 10040.0 54240.0 ;
      RECT  10160.0 54310.0 10230.0 54240.0 ;
      RECT  9970.0 54275.0 10040.0 53912.5 ;
      RECT  10005.0 54310.0 10195.0 54240.0 ;
      RECT  10160.0 54617.5 10230.0 54275.0 ;
      RECT  9970.0 53912.5 10040.0 53777.5 ;
      RECT  10160.0 54752.5 10230.0 54617.5 ;
      RECT  10262.5 54310.0 10127.5 54240.0 ;
      RECT  8895.0 54220.0 8965.0 54355.0 ;
      RECT  9035.0 54492.5 9105.0 54627.5 ;
      RECT  10032.5 54455.0 9897.5 54525.0 ;
      RECT  9970.0 55520.0 10040.0 55590.0 ;
      RECT  10160.0 55520.0 10230.0 55590.0 ;
      RECT  9970.0 55555.0 10040.0 55917.5 ;
      RECT  10005.0 55520.0 10195.0 55590.0 ;
      RECT  10160.0 55212.5 10230.0 55555.0 ;
      RECT  9970.0 55917.5 10040.0 56052.5 ;
      RECT  10160.0 55077.5 10230.0 55212.5 ;
      RECT  10262.5 55520.0 10127.5 55590.0 ;
      RECT  8895.0 55475.0 8965.0 55610.0 ;
      RECT  9035.0 55202.5 9105.0 55337.5 ;
      RECT  10032.5 55305.0 9897.5 55375.0 ;
      RECT  9970.0 57000.0 10040.0 56930.0 ;
      RECT  10160.0 57000.0 10230.0 56930.0 ;
      RECT  9970.0 56965.0 10040.0 56602.5 ;
      RECT  10005.0 57000.0 10195.0 56930.0 ;
      RECT  10160.0 57307.5 10230.0 56965.0 ;
      RECT  9970.0 56602.5 10040.0 56467.5 ;
      RECT  10160.0 57442.5 10230.0 57307.5 ;
      RECT  10262.5 57000.0 10127.5 56930.0 ;
      RECT  8895.0 56910.0 8965.0 57045.0 ;
      RECT  9035.0 57182.5 9105.0 57317.5 ;
      RECT  10032.5 57145.0 9897.5 57215.0 ;
      RECT  9970.0 58210.0 10040.0 58280.0 ;
      RECT  10160.0 58210.0 10230.0 58280.0 ;
      RECT  9970.0 58245.0 10040.0 58607.5 ;
      RECT  10005.0 58210.0 10195.0 58280.0 ;
      RECT  10160.0 57902.5 10230.0 58245.0 ;
      RECT  9970.0 58607.5 10040.0 58742.5 ;
      RECT  10160.0 57767.5 10230.0 57902.5 ;
      RECT  10262.5 58210.0 10127.5 58280.0 ;
      RECT  8895.0 58165.0 8965.0 58300.0 ;
      RECT  9035.0 57892.5 9105.0 58027.5 ;
      RECT  10032.5 57995.0 9897.5 58065.0 ;
      RECT  9970.0 59690.0 10040.0 59620.0 ;
      RECT  10160.0 59690.0 10230.0 59620.0 ;
      RECT  9970.0 59655.0 10040.0 59292.5 ;
      RECT  10005.0 59690.0 10195.0 59620.0 ;
      RECT  10160.0 59997.5 10230.0 59655.0 ;
      RECT  9970.0 59292.5 10040.0 59157.5 ;
      RECT  10160.0 60132.5 10230.0 59997.5 ;
      RECT  10262.5 59690.0 10127.5 59620.0 ;
      RECT  8895.0 59600.0 8965.0 59735.0 ;
      RECT  9035.0 59872.5 9105.0 60007.5 ;
      RECT  10032.5 59835.0 9897.5 59905.0 ;
      RECT  9970.0 60900.0 10040.0 60970.0 ;
      RECT  10160.0 60900.0 10230.0 60970.0 ;
      RECT  9970.0 60935.0 10040.0 61297.5 ;
      RECT  10005.0 60900.0 10195.0 60970.0 ;
      RECT  10160.0 60592.5 10230.0 60935.0 ;
      RECT  9970.0 61297.5 10040.0 61432.5 ;
      RECT  10160.0 60457.5 10230.0 60592.5 ;
      RECT  10262.5 60900.0 10127.5 60970.0 ;
      RECT  8895.0 60855.0 8965.0 60990.0 ;
      RECT  9035.0 60582.5 9105.0 60717.5 ;
      RECT  10032.5 60685.0 9897.5 60755.0 ;
      RECT  9970.0 62380.0 10040.0 62310.0 ;
      RECT  10160.0 62380.0 10230.0 62310.0 ;
      RECT  9970.0 62345.0 10040.0 61982.5 ;
      RECT  10005.0 62380.0 10195.0 62310.0 ;
      RECT  10160.0 62687.5 10230.0 62345.0 ;
      RECT  9970.0 61982.5 10040.0 61847.5 ;
      RECT  10160.0 62822.5 10230.0 62687.5 ;
      RECT  10262.5 62380.0 10127.5 62310.0 ;
      RECT  8895.0 62290.0 8965.0 62425.0 ;
      RECT  9035.0 62562.5 9105.0 62697.5 ;
      RECT  10032.5 62525.0 9897.5 62595.0 ;
      RECT  9970.0 63590.0 10040.0 63660.0 ;
      RECT  10160.0 63590.0 10230.0 63660.0 ;
      RECT  9970.0 63625.0 10040.0 63987.5 ;
      RECT  10005.0 63590.0 10195.0 63660.0 ;
      RECT  10160.0 63282.5 10230.0 63625.0 ;
      RECT  9970.0 63987.5 10040.0 64122.5 ;
      RECT  10160.0 63147.5 10230.0 63282.5 ;
      RECT  10262.5 63590.0 10127.5 63660.0 ;
      RECT  8895.0 63545.0 8965.0 63680.0 ;
      RECT  9035.0 63272.5 9105.0 63407.5 ;
      RECT  10032.5 63375.0 9897.5 63445.0 ;
      RECT  9970.0 65070.0 10040.0 65000.0 ;
      RECT  10160.0 65070.0 10230.0 65000.0 ;
      RECT  9970.0 65035.0 10040.0 64672.5 ;
      RECT  10005.0 65070.0 10195.0 65000.0 ;
      RECT  10160.0 65377.5 10230.0 65035.0 ;
      RECT  9970.0 64672.5 10040.0 64537.5 ;
      RECT  10160.0 65512.5 10230.0 65377.5 ;
      RECT  10262.5 65070.0 10127.5 65000.0 ;
      RECT  8895.0 64980.0 8965.0 65115.0 ;
      RECT  9035.0 65252.5 9105.0 65387.5 ;
      RECT  10032.5 65215.0 9897.5 65285.0 ;
      RECT  9970.0 66280.0 10040.0 66350.0 ;
      RECT  10160.0 66280.0 10230.0 66350.0 ;
      RECT  9970.0 66315.0 10040.0 66677.5 ;
      RECT  10005.0 66280.0 10195.0 66350.0 ;
      RECT  10160.0 65972.5 10230.0 66315.0 ;
      RECT  9970.0 66677.5 10040.0 66812.5 ;
      RECT  10160.0 65837.5 10230.0 65972.5 ;
      RECT  10262.5 66280.0 10127.5 66350.0 ;
      RECT  8895.0 66235.0 8965.0 66370.0 ;
      RECT  9035.0 65962.5 9105.0 66097.5 ;
      RECT  10032.5 66065.0 9897.5 66135.0 ;
      RECT  9970.0 67760.0 10040.0 67690.0 ;
      RECT  10160.0 67760.0 10230.0 67690.0 ;
      RECT  9970.0 67725.0 10040.0 67362.5 ;
      RECT  10005.0 67760.0 10195.0 67690.0 ;
      RECT  10160.0 68067.5 10230.0 67725.0 ;
      RECT  9970.0 67362.5 10040.0 67227.5 ;
      RECT  10160.0 68202.5 10230.0 68067.5 ;
      RECT  10262.5 67760.0 10127.5 67690.0 ;
      RECT  8895.0 67670.0 8965.0 67805.0 ;
      RECT  9035.0 67942.5 9105.0 68077.5 ;
      RECT  10032.5 67905.0 9897.5 67975.0 ;
      RECT  9970.0 68970.0 10040.0 69040.0 ;
      RECT  10160.0 68970.0 10230.0 69040.0 ;
      RECT  9970.0 69005.0 10040.0 69367.5 ;
      RECT  10005.0 68970.0 10195.0 69040.0 ;
      RECT  10160.0 68662.5 10230.0 69005.0 ;
      RECT  9970.0 69367.5 10040.0 69502.5 ;
      RECT  10160.0 68527.5 10230.0 68662.5 ;
      RECT  10262.5 68970.0 10127.5 69040.0 ;
      RECT  8895.0 68925.0 8965.0 69060.0 ;
      RECT  9035.0 68652.5 9105.0 68787.5 ;
      RECT  10032.5 68755.0 9897.5 68825.0 ;
      RECT  9970.0 70450.0 10040.0 70380.0 ;
      RECT  10160.0 70450.0 10230.0 70380.0 ;
      RECT  9970.0 70415.0 10040.0 70052.5 ;
      RECT  10005.0 70450.0 10195.0 70380.0 ;
      RECT  10160.0 70757.5 10230.0 70415.0 ;
      RECT  9970.0 70052.5 10040.0 69917.5 ;
      RECT  10160.0 70892.5 10230.0 70757.5 ;
      RECT  10262.5 70450.0 10127.5 70380.0 ;
      RECT  8895.0 70360.0 8965.0 70495.0 ;
      RECT  9035.0 70632.5 9105.0 70767.5 ;
      RECT  10032.5 70595.0 9897.5 70665.0 ;
      RECT  9970.0 71660.0 10040.0 71730.0 ;
      RECT  10160.0 71660.0 10230.0 71730.0 ;
      RECT  9970.0 71695.0 10040.0 72057.5 ;
      RECT  10005.0 71660.0 10195.0 71730.0 ;
      RECT  10160.0 71352.5 10230.0 71695.0 ;
      RECT  9970.0 72057.5 10040.0 72192.5 ;
      RECT  10160.0 71217.5 10230.0 71352.5 ;
      RECT  10262.5 71660.0 10127.5 71730.0 ;
      RECT  8895.0 71615.0 8965.0 71750.0 ;
      RECT  9035.0 71342.5 9105.0 71477.5 ;
      RECT  10032.5 71445.0 9897.5 71515.0 ;
      RECT  9970.0 73140.0 10040.0 73070.0 ;
      RECT  10160.0 73140.0 10230.0 73070.0 ;
      RECT  9970.0 73105.0 10040.0 72742.5 ;
      RECT  10005.0 73140.0 10195.0 73070.0 ;
      RECT  10160.0 73447.5 10230.0 73105.0 ;
      RECT  9970.0 72742.5 10040.0 72607.5 ;
      RECT  10160.0 73582.5 10230.0 73447.5 ;
      RECT  10262.5 73140.0 10127.5 73070.0 ;
      RECT  8895.0 73050.0 8965.0 73185.0 ;
      RECT  9035.0 73322.5 9105.0 73457.5 ;
      RECT  10032.5 73285.0 9897.5 73355.0 ;
      RECT  9970.0 74350.0 10040.0 74420.0 ;
      RECT  10160.0 74350.0 10230.0 74420.0 ;
      RECT  9970.0 74385.0 10040.0 74747.5 ;
      RECT  10005.0 74350.0 10195.0 74420.0 ;
      RECT  10160.0 74042.5 10230.0 74385.0 ;
      RECT  9970.0 74747.5 10040.0 74882.5 ;
      RECT  10160.0 73907.5 10230.0 74042.5 ;
      RECT  10262.5 74350.0 10127.5 74420.0 ;
      RECT  8895.0 74305.0 8965.0 74440.0 ;
      RECT  9035.0 74032.5 9105.0 74167.5 ;
      RECT  10032.5 74135.0 9897.5 74205.0 ;
      RECT  9970.0 75830.0 10040.0 75760.0 ;
      RECT  10160.0 75830.0 10230.0 75760.0 ;
      RECT  9970.0 75795.0 10040.0 75432.5 ;
      RECT  10005.0 75830.0 10195.0 75760.0 ;
      RECT  10160.0 76137.5 10230.0 75795.0 ;
      RECT  9970.0 75432.5 10040.0 75297.5 ;
      RECT  10160.0 76272.5 10230.0 76137.5 ;
      RECT  10262.5 75830.0 10127.5 75760.0 ;
      RECT  8895.0 75740.0 8965.0 75875.0 ;
      RECT  9035.0 76012.5 9105.0 76147.5 ;
      RECT  10032.5 75975.0 9897.5 76045.0 ;
      RECT  9970.0 77040.0 10040.0 77110.0 ;
      RECT  10160.0 77040.0 10230.0 77110.0 ;
      RECT  9970.0 77075.0 10040.0 77437.5 ;
      RECT  10005.0 77040.0 10195.0 77110.0 ;
      RECT  10160.0 76732.5 10230.0 77075.0 ;
      RECT  9970.0 77437.5 10040.0 77572.5 ;
      RECT  10160.0 76597.5 10230.0 76732.5 ;
      RECT  10262.5 77040.0 10127.5 77110.0 ;
      RECT  8895.0 76995.0 8965.0 77130.0 ;
      RECT  9035.0 76722.5 9105.0 76857.5 ;
      RECT  10032.5 76825.0 9897.5 76895.0 ;
      RECT  9970.0 78520.0 10040.0 78450.0 ;
      RECT  10160.0 78520.0 10230.0 78450.0 ;
      RECT  9970.0 78485.0 10040.0 78122.5 ;
      RECT  10005.0 78520.0 10195.0 78450.0 ;
      RECT  10160.0 78827.5 10230.0 78485.0 ;
      RECT  9970.0 78122.5 10040.0 77987.5 ;
      RECT  10160.0 78962.5 10230.0 78827.5 ;
      RECT  10262.5 78520.0 10127.5 78450.0 ;
      RECT  8895.0 78430.0 8965.0 78565.0 ;
      RECT  9035.0 78702.5 9105.0 78837.5 ;
      RECT  10032.5 78665.0 9897.5 78735.0 ;
      RECT  9970.0 79730.0 10040.0 79800.0 ;
      RECT  10160.0 79730.0 10230.0 79800.0 ;
      RECT  9970.0 79765.0 10040.0 80127.5 ;
      RECT  10005.0 79730.0 10195.0 79800.0 ;
      RECT  10160.0 79422.5 10230.0 79765.0 ;
      RECT  9970.0 80127.5 10040.0 80262.5 ;
      RECT  10160.0 79287.5 10230.0 79422.5 ;
      RECT  10262.5 79730.0 10127.5 79800.0 ;
      RECT  8895.0 79685.0 8965.0 79820.0 ;
      RECT  9035.0 79412.5 9105.0 79547.5 ;
      RECT  10032.5 79515.0 9897.5 79585.0 ;
      RECT  9970.0 81210.0 10040.0 81140.0 ;
      RECT  10160.0 81210.0 10230.0 81140.0 ;
      RECT  9970.0 81175.0 10040.0 80812.5 ;
      RECT  10005.0 81210.0 10195.0 81140.0 ;
      RECT  10160.0 81517.5 10230.0 81175.0 ;
      RECT  9970.0 80812.5 10040.0 80677.5 ;
      RECT  10160.0 81652.5 10230.0 81517.5 ;
      RECT  10262.5 81210.0 10127.5 81140.0 ;
      RECT  8895.0 81120.0 8965.0 81255.0 ;
      RECT  9035.0 81392.5 9105.0 81527.5 ;
      RECT  10032.5 81355.0 9897.5 81425.0 ;
      RECT  9970.0 82420.0 10040.0 82490.0 ;
      RECT  10160.0 82420.0 10230.0 82490.0 ;
      RECT  9970.0 82455.0 10040.0 82817.5 ;
      RECT  10005.0 82420.0 10195.0 82490.0 ;
      RECT  10160.0 82112.5 10230.0 82455.0 ;
      RECT  9970.0 82817.5 10040.0 82952.5 ;
      RECT  10160.0 81977.5 10230.0 82112.5 ;
      RECT  10262.5 82420.0 10127.5 82490.0 ;
      RECT  8895.0 82375.0 8965.0 82510.0 ;
      RECT  9035.0 82102.5 9105.0 82237.5 ;
      RECT  10032.5 82205.0 9897.5 82275.0 ;
      RECT  9970.0 83900.0 10040.0 83830.0 ;
      RECT  10160.0 83900.0 10230.0 83830.0 ;
      RECT  9970.0 83865.0 10040.0 83502.5 ;
      RECT  10005.0 83900.0 10195.0 83830.0 ;
      RECT  10160.0 84207.5 10230.0 83865.0 ;
      RECT  9970.0 83502.5 10040.0 83367.5 ;
      RECT  10160.0 84342.5 10230.0 84207.5 ;
      RECT  10262.5 83900.0 10127.5 83830.0 ;
      RECT  8895.0 83810.0 8965.0 83945.0 ;
      RECT  9035.0 84082.5 9105.0 84217.5 ;
      RECT  10032.5 84045.0 9897.5 84115.0 ;
      RECT  9970.0 85110.0 10040.0 85180.0 ;
      RECT  10160.0 85110.0 10230.0 85180.0 ;
      RECT  9970.0 85145.0 10040.0 85507.5 ;
      RECT  10005.0 85110.0 10195.0 85180.0 ;
      RECT  10160.0 84802.5 10230.0 85145.0 ;
      RECT  9970.0 85507.5 10040.0 85642.5 ;
      RECT  10160.0 84667.5 10230.0 84802.5 ;
      RECT  10262.5 85110.0 10127.5 85180.0 ;
      RECT  8895.0 85065.0 8965.0 85200.0 ;
      RECT  9035.0 84792.5 9105.0 84927.5 ;
      RECT  10032.5 84895.0 9897.5 84965.0 ;
      RECT  9970.0 86590.0 10040.0 86520.0 ;
      RECT  10160.0 86590.0 10230.0 86520.0 ;
      RECT  9970.0 86555.0 10040.0 86192.5 ;
      RECT  10005.0 86590.0 10195.0 86520.0 ;
      RECT  10160.0 86897.5 10230.0 86555.0 ;
      RECT  9970.0 86192.5 10040.0 86057.5 ;
      RECT  10160.0 87032.5 10230.0 86897.5 ;
      RECT  10262.5 86590.0 10127.5 86520.0 ;
      RECT  8895.0 86500.0 8965.0 86635.0 ;
      RECT  9035.0 86772.5 9105.0 86907.5 ;
      RECT  10032.5 86735.0 9897.5 86805.0 ;
      RECT  9970.0 87800.0 10040.0 87870.0 ;
      RECT  10160.0 87800.0 10230.0 87870.0 ;
      RECT  9970.0 87835.0 10040.0 88197.5 ;
      RECT  10005.0 87800.0 10195.0 87870.0 ;
      RECT  10160.0 87492.5 10230.0 87835.0 ;
      RECT  9970.0 88197.5 10040.0 88332.5 ;
      RECT  10160.0 87357.5 10230.0 87492.5 ;
      RECT  10262.5 87800.0 10127.5 87870.0 ;
      RECT  8895.0 87755.0 8965.0 87890.0 ;
      RECT  9035.0 87482.5 9105.0 87617.5 ;
      RECT  10032.5 87585.0 9897.5 87655.0 ;
      RECT  9970.0 89280.0 10040.0 89210.0 ;
      RECT  10160.0 89280.0 10230.0 89210.0 ;
      RECT  9970.0 89245.0 10040.0 88882.5 ;
      RECT  10005.0 89280.0 10195.0 89210.0 ;
      RECT  10160.0 89587.5 10230.0 89245.0 ;
      RECT  9970.0 88882.5 10040.0 88747.5 ;
      RECT  10160.0 89722.5 10230.0 89587.5 ;
      RECT  10262.5 89280.0 10127.5 89210.0 ;
      RECT  8895.0 89190.0 8965.0 89325.0 ;
      RECT  9035.0 89462.5 9105.0 89597.5 ;
      RECT  10032.5 89425.0 9897.5 89495.0 ;
      RECT  9970.0 90490.0 10040.0 90560.0 ;
      RECT  10160.0 90490.0 10230.0 90560.0 ;
      RECT  9970.0 90525.0 10040.0 90887.5 ;
      RECT  10005.0 90490.0 10195.0 90560.0 ;
      RECT  10160.0 90182.5 10230.0 90525.0 ;
      RECT  9970.0 90887.5 10040.0 91022.5 ;
      RECT  10160.0 90047.5 10230.0 90182.5 ;
      RECT  10262.5 90490.0 10127.5 90560.0 ;
      RECT  8895.0 90445.0 8965.0 90580.0 ;
      RECT  9035.0 90172.5 9105.0 90307.5 ;
      RECT  10032.5 90275.0 9897.5 90345.0 ;
      RECT  9970.0 91970.0 10040.0 91900.0 ;
      RECT  10160.0 91970.0 10230.0 91900.0 ;
      RECT  9970.0 91935.0 10040.0 91572.5 ;
      RECT  10005.0 91970.0 10195.0 91900.0 ;
      RECT  10160.0 92277.5 10230.0 91935.0 ;
      RECT  9970.0 91572.5 10040.0 91437.5 ;
      RECT  10160.0 92412.5 10230.0 92277.5 ;
      RECT  10262.5 91970.0 10127.5 91900.0 ;
      RECT  8895.0 91880.0 8965.0 92015.0 ;
      RECT  9035.0 92152.5 9105.0 92287.5 ;
      RECT  10032.5 92115.0 9897.5 92185.0 ;
      RECT  9970.0 93180.0 10040.0 93250.0 ;
      RECT  10160.0 93180.0 10230.0 93250.0 ;
      RECT  9970.0 93215.0 10040.0 93577.5 ;
      RECT  10005.0 93180.0 10195.0 93250.0 ;
      RECT  10160.0 92872.5 10230.0 93215.0 ;
      RECT  9970.0 93577.5 10040.0 93712.5 ;
      RECT  10160.0 92737.5 10230.0 92872.5 ;
      RECT  10262.5 93180.0 10127.5 93250.0 ;
      RECT  8895.0 93135.0 8965.0 93270.0 ;
      RECT  9035.0 92862.5 9105.0 92997.5 ;
      RECT  10032.5 92965.0 9897.5 93035.0 ;
      RECT  9970.0 94660.0 10040.0 94590.0 ;
      RECT  10160.0 94660.0 10230.0 94590.0 ;
      RECT  9970.0 94625.0 10040.0 94262.5 ;
      RECT  10005.0 94660.0 10195.0 94590.0 ;
      RECT  10160.0 94967.5 10230.0 94625.0 ;
      RECT  9970.0 94262.5 10040.0 94127.5 ;
      RECT  10160.0 95102.5 10230.0 94967.5 ;
      RECT  10262.5 94660.0 10127.5 94590.0 ;
      RECT  8895.0 94570.0 8965.0 94705.0 ;
      RECT  9035.0 94842.5 9105.0 94977.5 ;
      RECT  10032.5 94805.0 9897.5 94875.0 ;
      RECT  9970.0 95870.0 10040.0 95940.0 ;
      RECT  10160.0 95870.0 10230.0 95940.0 ;
      RECT  9970.0 95905.0 10040.0 96267.5 ;
      RECT  10005.0 95870.0 10195.0 95940.0 ;
      RECT  10160.0 95562.5 10230.0 95905.0 ;
      RECT  9970.0 96267.5 10040.0 96402.5 ;
      RECT  10160.0 95427.5 10230.0 95562.5 ;
      RECT  10262.5 95870.0 10127.5 95940.0 ;
      RECT  8895.0 95825.0 8965.0 95960.0 ;
      RECT  9035.0 95552.5 9105.0 95687.5 ;
      RECT  10032.5 95655.0 9897.5 95725.0 ;
      RECT  9970.0 97350.0 10040.0 97280.0 ;
      RECT  10160.0 97350.0 10230.0 97280.0 ;
      RECT  9970.0 97315.0 10040.0 96952.5 ;
      RECT  10005.0 97350.0 10195.0 97280.0 ;
      RECT  10160.0 97657.5 10230.0 97315.0 ;
      RECT  9970.0 96952.5 10040.0 96817.5 ;
      RECT  10160.0 97792.5 10230.0 97657.5 ;
      RECT  10262.5 97350.0 10127.5 97280.0 ;
      RECT  8895.0 97260.0 8965.0 97395.0 ;
      RECT  9035.0 97532.5 9105.0 97667.5 ;
      RECT  10032.5 97495.0 9897.5 97565.0 ;
      RECT  9970.0 98560.0 10040.0 98630.0 ;
      RECT  10160.0 98560.0 10230.0 98630.0 ;
      RECT  9970.0 98595.0 10040.0 98957.5 ;
      RECT  10005.0 98560.0 10195.0 98630.0 ;
      RECT  10160.0 98252.5 10230.0 98595.0 ;
      RECT  9970.0 98957.5 10040.0 99092.5 ;
      RECT  10160.0 98117.5 10230.0 98252.5 ;
      RECT  10262.5 98560.0 10127.5 98630.0 ;
      RECT  8895.0 98515.0 8965.0 98650.0 ;
      RECT  9035.0 98242.5 9105.0 98377.5 ;
      RECT  10032.5 98345.0 9897.5 98415.0 ;
      RECT  9970.0 100040.0 10040.0 99970.0 ;
      RECT  10160.0 100040.0 10230.0 99970.0 ;
      RECT  9970.0 100005.0 10040.0 99642.5 ;
      RECT  10005.0 100040.0 10195.0 99970.0 ;
      RECT  10160.0 100347.5 10230.0 100005.0 ;
      RECT  9970.0 99642.5 10040.0 99507.5 ;
      RECT  10160.0 100482.5 10230.0 100347.5 ;
      RECT  10262.5 100040.0 10127.5 99970.0 ;
      RECT  8895.0 99950.0 8965.0 100085.0 ;
      RECT  9035.0 100222.5 9105.0 100357.5 ;
      RECT  10032.5 100185.0 9897.5 100255.0 ;
      RECT  9970.0 101250.0 10040.0 101320.0 ;
      RECT  10160.0 101250.0 10230.0 101320.0 ;
      RECT  9970.0 101285.0 10040.0 101647.5 ;
      RECT  10005.0 101250.0 10195.0 101320.0 ;
      RECT  10160.0 100942.5 10230.0 101285.0 ;
      RECT  9970.0 101647.5 10040.0 101782.5 ;
      RECT  10160.0 100807.5 10230.0 100942.5 ;
      RECT  10262.5 101250.0 10127.5 101320.0 ;
      RECT  8895.0 101205.0 8965.0 101340.0 ;
      RECT  9035.0 100932.5 9105.0 101067.5 ;
      RECT  10032.5 101035.0 9897.5 101105.0 ;
      RECT  9970.0 102730.0 10040.0 102660.0 ;
      RECT  10160.0 102730.0 10230.0 102660.0 ;
      RECT  9970.0 102695.0 10040.0 102332.5 ;
      RECT  10005.0 102730.0 10195.0 102660.0 ;
      RECT  10160.0 103037.5 10230.0 102695.0 ;
      RECT  9970.0 102332.5 10040.0 102197.5 ;
      RECT  10160.0 103172.5 10230.0 103037.5 ;
      RECT  10262.5 102730.0 10127.5 102660.0 ;
      RECT  8895.0 102640.0 8965.0 102775.0 ;
      RECT  9035.0 102912.5 9105.0 103047.5 ;
      RECT  10032.5 102875.0 9897.5 102945.0 ;
      RECT  9970.0 103940.0 10040.0 104010.0 ;
      RECT  10160.0 103940.0 10230.0 104010.0 ;
      RECT  9970.0 103975.0 10040.0 104337.5 ;
      RECT  10005.0 103940.0 10195.0 104010.0 ;
      RECT  10160.0 103632.5 10230.0 103975.0 ;
      RECT  9970.0 104337.5 10040.0 104472.5 ;
      RECT  10160.0 103497.5 10230.0 103632.5 ;
      RECT  10262.5 103940.0 10127.5 104010.0 ;
      RECT  8895.0 103895.0 8965.0 104030.0 ;
      RECT  9035.0 103622.5 9105.0 103757.5 ;
      RECT  10032.5 103725.0 9897.5 103795.0 ;
      RECT  9970.0 105420.0 10040.0 105350.0 ;
      RECT  10160.0 105420.0 10230.0 105350.0 ;
      RECT  9970.0 105385.0 10040.0 105022.5 ;
      RECT  10005.0 105420.0 10195.0 105350.0 ;
      RECT  10160.0 105727.5 10230.0 105385.0 ;
      RECT  9970.0 105022.5 10040.0 104887.5 ;
      RECT  10160.0 105862.5 10230.0 105727.5 ;
      RECT  10262.5 105420.0 10127.5 105350.0 ;
      RECT  8895.0 105330.0 8965.0 105465.0 ;
      RECT  9035.0 105602.5 9105.0 105737.5 ;
      RECT  10032.5 105565.0 9897.5 105635.0 ;
      RECT  9970.0 106630.0 10040.0 106700.0 ;
      RECT  10160.0 106630.0 10230.0 106700.0 ;
      RECT  9970.0 106665.0 10040.0 107027.5 ;
      RECT  10005.0 106630.0 10195.0 106700.0 ;
      RECT  10160.0 106322.5 10230.0 106665.0 ;
      RECT  9970.0 107027.5 10040.0 107162.5 ;
      RECT  10160.0 106187.5 10230.0 106322.5 ;
      RECT  10262.5 106630.0 10127.5 106700.0 ;
      RECT  8895.0 106585.0 8965.0 106720.0 ;
      RECT  9035.0 106312.5 9105.0 106447.5 ;
      RECT  10032.5 106415.0 9897.5 106485.0 ;
      RECT  9970.0 108110.0 10040.0 108040.0 ;
      RECT  10160.0 108110.0 10230.0 108040.0 ;
      RECT  9970.0 108075.0 10040.0 107712.5 ;
      RECT  10005.0 108110.0 10195.0 108040.0 ;
      RECT  10160.0 108417.5 10230.0 108075.0 ;
      RECT  9970.0 107712.5 10040.0 107577.5 ;
      RECT  10160.0 108552.5 10230.0 108417.5 ;
      RECT  10262.5 108110.0 10127.5 108040.0 ;
      RECT  8895.0 108020.0 8965.0 108155.0 ;
      RECT  9035.0 108292.5 9105.0 108427.5 ;
      RECT  10032.5 108255.0 9897.5 108325.0 ;
      RECT  9970.0 109320.0 10040.0 109390.0 ;
      RECT  10160.0 109320.0 10230.0 109390.0 ;
      RECT  9970.0 109355.0 10040.0 109717.5 ;
      RECT  10005.0 109320.0 10195.0 109390.0 ;
      RECT  10160.0 109012.5 10230.0 109355.0 ;
      RECT  9970.0 109717.5 10040.0 109852.5 ;
      RECT  10160.0 108877.5 10230.0 109012.5 ;
      RECT  10262.5 109320.0 10127.5 109390.0 ;
      RECT  8895.0 109275.0 8965.0 109410.0 ;
      RECT  9035.0 109002.5 9105.0 109137.5 ;
      RECT  10032.5 109105.0 9897.5 109175.0 ;
      RECT  9970.0 110800.0 10040.0 110730.0 ;
      RECT  10160.0 110800.0 10230.0 110730.0 ;
      RECT  9970.0 110765.0 10040.0 110402.5 ;
      RECT  10005.0 110800.0 10195.0 110730.0 ;
      RECT  10160.0 111107.5 10230.0 110765.0 ;
      RECT  9970.0 110402.5 10040.0 110267.5 ;
      RECT  10160.0 111242.5 10230.0 111107.5 ;
      RECT  10262.5 110800.0 10127.5 110730.0 ;
      RECT  8895.0 110710.0 8965.0 110845.0 ;
      RECT  9035.0 110982.5 9105.0 111117.5 ;
      RECT  10032.5 110945.0 9897.5 111015.0 ;
      RECT  9970.0 112010.0 10040.0 112080.0 ;
      RECT  10160.0 112010.0 10230.0 112080.0 ;
      RECT  9970.0 112045.0 10040.0 112407.5 ;
      RECT  10005.0 112010.0 10195.0 112080.0 ;
      RECT  10160.0 111702.5 10230.0 112045.0 ;
      RECT  9970.0 112407.5 10040.0 112542.5 ;
      RECT  10160.0 111567.5 10230.0 111702.5 ;
      RECT  10262.5 112010.0 10127.5 112080.0 ;
      RECT  8895.0 111965.0 8965.0 112100.0 ;
      RECT  9035.0 111692.5 9105.0 111827.5 ;
      RECT  10032.5 111795.0 9897.5 111865.0 ;
      RECT  9970.0 113490.0 10040.0 113420.0 ;
      RECT  10160.0 113490.0 10230.0 113420.0 ;
      RECT  9970.0 113455.0 10040.0 113092.5 ;
      RECT  10005.0 113490.0 10195.0 113420.0 ;
      RECT  10160.0 113797.5 10230.0 113455.0 ;
      RECT  9970.0 113092.5 10040.0 112957.5 ;
      RECT  10160.0 113932.5 10230.0 113797.5 ;
      RECT  10262.5 113490.0 10127.5 113420.0 ;
      RECT  8895.0 113400.0 8965.0 113535.0 ;
      RECT  9035.0 113672.5 9105.0 113807.5 ;
      RECT  10032.5 113635.0 9897.5 113705.0 ;
      RECT  8895.0 28015.0 8965.0 114095.0 ;
      RECT  4655.0 11465.0 11095.0 10760.0 ;
      RECT  4655.0 10055.0 11095.0 10760.0 ;
      RECT  4655.0 10055.0 11095.0 9350.0 ;
      RECT  4655.0 8645.0 11095.0 9350.0 ;
      RECT  4655.0 8645.0 11095.0 7940.0 ;
      RECT  4655.0 7235.0 11095.0 7940.0 ;
      RECT  4655.0 7235.0 11095.0 6530.0 ;
      RECT  4655.0 5825.0 11095.0 6530.0 ;
      RECT  4655.0 11147.5 4800.0 11077.5 ;
      RECT  4655.0 10442.5 4800.0 10372.5 ;
      RECT  4655.0 9737.5 4800.0 9667.5 ;
      RECT  4655.0 9032.5 4800.0 8962.5 ;
      RECT  4655.0 8327.5 4800.0 8257.5 ;
      RECT  4655.0 7622.5 4800.0 7552.5 ;
      RECT  4655.0 6917.5 4800.0 6847.5 ;
      RECT  4655.0 6212.5 4800.0 6142.5 ;
      RECT  10825.0 11147.5 11095.0 11077.5 ;
      RECT  10407.5 11302.5 11095.0 11232.5 ;
      RECT  10825.0 10442.5 11095.0 10372.5 ;
      RECT  10407.5 10287.5 11095.0 10217.5 ;
      RECT  10825.0 9737.5 11095.0 9667.5 ;
      RECT  10407.5 9892.5 11095.0 9822.5 ;
      RECT  10825.0 9032.5 11095.0 8962.5 ;
      RECT  10407.5 8877.5 11095.0 8807.5 ;
      RECT  10825.0 8327.5 11095.0 8257.5 ;
      RECT  10407.5 8482.5 11095.0 8412.5 ;
      RECT  10825.0 7622.5 11095.0 7552.5 ;
      RECT  10407.5 7467.5 11095.0 7397.5 ;
      RECT  10825.0 6917.5 11095.0 6847.5 ;
      RECT  10407.5 7072.5 11095.0 7002.5 ;
      RECT  10825.0 6212.5 11095.0 6142.5 ;
      RECT  10407.5 6057.5 11095.0 5987.5 ;
      RECT  4655.0 11500.0 11095.0 11430.0 ;
      RECT  4655.0 10795.0 11095.0 10725.0 ;
      RECT  4655.0 10090.0 11095.0 10020.0 ;
      RECT  4655.0 9385.0 11095.0 9315.0 ;
      RECT  4655.0 8680.0 11095.0 8610.0 ;
      RECT  4655.0 7975.0 11095.0 7905.0 ;
      RECT  4655.0 7270.0 11095.0 7200.0 ;
      RECT  4655.0 6565.0 11095.0 6495.0 ;
      RECT  4655.0 5860.0 11095.0 5790.0 ;
      RECT  15857.5 6520.0 15927.5 6655.0 ;
      RECT  18677.5 6520.0 18747.5 6655.0 ;
      RECT  21497.5 6520.0 21567.5 6655.0 ;
      RECT  24317.5 6520.0 24387.5 6655.0 ;
      RECT  27137.5 6520.0 27207.5 6655.0 ;
      RECT  29957.5 6520.0 30027.5 6655.0 ;
      RECT  32777.5 6520.0 32847.5 6655.0 ;
      RECT  35597.5 6520.0 35667.5 6655.0 ;
      RECT  38417.5 6520.0 38487.5 6655.0 ;
      RECT  41237.5 6520.0 41307.5 6655.0 ;
      RECT  44057.5 6520.0 44127.5 6655.0 ;
      RECT  46877.5 6520.0 46947.5 6655.0 ;
      RECT  49697.5 6520.0 49767.5 6655.0 ;
      RECT  52517.5 6520.0 52587.5 6655.0 ;
      RECT  55337.5 6520.0 55407.5 6655.0 ;
      RECT  58157.5 6520.0 58227.5 6655.0 ;
      RECT  60977.5 6520.0 61047.5 6655.0 ;
      RECT  63797.5 6520.0 63867.5 6655.0 ;
      RECT  66617.5 6520.0 66687.5 6655.0 ;
      RECT  69437.5 6520.0 69507.5 6655.0 ;
      RECT  72257.5 6520.0 72327.5 6655.0 ;
      RECT  75077.5 6520.0 75147.5 6655.0 ;
      RECT  77897.5 6520.0 77967.5 6655.0 ;
      RECT  80717.5 6520.0 80787.5 6655.0 ;
      RECT  83537.5 6520.0 83607.5 6655.0 ;
      RECT  86357.5 6520.0 86427.5 6655.0 ;
      RECT  89177.5 6520.0 89247.5 6655.0 ;
      RECT  91997.5 6520.0 92067.5 6655.0 ;
      RECT  94817.5 6520.0 94887.5 6655.0 ;
      RECT  97637.5 6520.0 97707.5 6655.0 ;
      RECT  100457.5 6520.0 100527.5 6655.0 ;
      RECT  103277.5 6520.0 103347.5 6655.0 ;
      RECT  16067.5 35.0 16137.5 170.0 ;
      RECT  18887.5 35.0 18957.5 170.0 ;
      RECT  21707.5 35.0 21777.5 170.0 ;
      RECT  24527.5 35.0 24597.5 170.0 ;
      RECT  27347.5 35.0 27417.5 170.0 ;
      RECT  30167.5 35.0 30237.5 170.0 ;
      RECT  32987.5 35.0 33057.5 170.0 ;
      RECT  35807.5 35.0 35877.5 170.0 ;
      RECT  38627.5 35.0 38697.5 170.0 ;
      RECT  41447.5 35.0 41517.5 170.0 ;
      RECT  44267.5 35.0 44337.5 170.0 ;
      RECT  47087.5 35.0 47157.5 170.0 ;
      RECT  49907.5 35.0 49977.5 170.0 ;
      RECT  52727.5 35.0 52797.5 170.0 ;
      RECT  55547.5 35.0 55617.5 170.0 ;
      RECT  58367.5 35.0 58437.5 170.0 ;
      RECT  61187.5 35.0 61257.5 170.0 ;
      RECT  64007.5 35.0 64077.5 170.0 ;
      RECT  66827.5 35.0 66897.5 170.0 ;
      RECT  69647.5 35.0 69717.5 170.0 ;
      RECT  72467.5 35.0 72537.5 170.0 ;
      RECT  75287.5 35.0 75357.5 170.0 ;
      RECT  78107.5 35.0 78177.5 170.0 ;
      RECT  80927.5 35.0 80997.5 170.0 ;
      RECT  83747.5 35.0 83817.5 170.0 ;
      RECT  86567.5 35.0 86637.5 170.0 ;
      RECT  89387.5 35.0 89457.5 170.0 ;
      RECT  92207.5 35.0 92277.5 170.0 ;
      RECT  95027.5 35.0 95097.5 170.0 ;
      RECT  97847.5 35.0 97917.5 170.0 ;
      RECT  100667.5 35.0 100737.5 170.0 ;
      RECT  103487.5 35.0 103557.5 170.0 ;
      RECT  13657.5 28050.0 13792.5 27980.0 ;
      RECT  13657.5 30740.0 13792.5 30670.0 ;
      RECT  13657.5 33430.0 13792.5 33360.0 ;
      RECT  13657.5 36120.0 13792.5 36050.0 ;
      RECT  13657.5 38810.0 13792.5 38740.0 ;
      RECT  13657.5 41500.0 13792.5 41430.0 ;
      RECT  13657.5 44190.0 13792.5 44120.0 ;
      RECT  13657.5 46880.0 13792.5 46810.0 ;
      RECT  13657.5 49570.0 13792.5 49500.0 ;
      RECT  13657.5 52260.0 13792.5 52190.0 ;
      RECT  13657.5 54950.0 13792.5 54880.0 ;
      RECT  13657.5 57640.0 13792.5 57570.0 ;
      RECT  13657.5 60330.0 13792.5 60260.0 ;
      RECT  13657.5 63020.0 13792.5 62950.0 ;
      RECT  13657.5 65710.0 13792.5 65640.0 ;
      RECT  13657.5 68400.0 13792.5 68330.0 ;
      RECT  13657.5 71090.0 13792.5 71020.0 ;
      RECT  13657.5 73780.0 13792.5 73710.0 ;
      RECT  13657.5 76470.0 13792.5 76400.0 ;
      RECT  13657.5 79160.0 13792.5 79090.0 ;
      RECT  13657.5 81850.0 13792.5 81780.0 ;
      RECT  13657.5 84540.0 13792.5 84470.0 ;
      RECT  13657.5 87230.0 13792.5 87160.0 ;
      RECT  13657.5 89920.0 13792.5 89850.0 ;
      RECT  13657.5 92610.0 13792.5 92540.0 ;
      RECT  13657.5 95300.0 13792.5 95230.0 ;
      RECT  13657.5 97990.0 13792.5 97920.0 ;
      RECT  13657.5 100680.0 13792.5 100610.0 ;
      RECT  13657.5 103370.0 13792.5 103300.0 ;
      RECT  13657.5 106060.0 13792.5 105990.0 ;
      RECT  13657.5 108750.0 13792.5 108680.0 ;
      RECT  13657.5 111440.0 13792.5 111370.0 ;
      RECT  13657.5 114130.0 13792.5 114060.0 ;
      RECT  11095.0 12045.0 10960.0 12115.0 ;
      RECT  11505.0 12045.0 11370.0 12115.0 ;
      RECT  10820.0 13390.0 10685.0 13460.0 ;
      RECT  11710.0 13390.0 11575.0 13460.0 ;
      RECT  11095.0 17425.0 10960.0 17495.0 ;
      RECT  11915.0 17425.0 11780.0 17495.0 ;
      RECT  10820.0 18770.0 10685.0 18840.0 ;
      RECT  12120.0 18770.0 11985.0 18840.0 ;
      RECT  11095.0 22805.0 10960.0 22875.0 ;
      RECT  12325.0 22805.0 12190.0 22875.0 ;
      RECT  10820.0 24150.0 10685.0 24220.0 ;
      RECT  12530.0 24150.0 12395.0 24220.0 ;
      RECT  11300.0 11840.0 11165.0 11910.0 ;
      RECT  11300.0 11840.0 11165.0 11910.0 ;
      RECT  13590.0 11910.0 13725.0 11840.0 ;
      RECT  11300.0 14530.0 11165.0 14600.0 ;
      RECT  11300.0 14530.0 11165.0 14600.0 ;
      RECT  13590.0 14600.0 13725.0 14530.0 ;
      RECT  11300.0 17220.0 11165.0 17290.0 ;
      RECT  11300.0 17220.0 11165.0 17290.0 ;
      RECT  13590.0 17290.0 13725.0 17220.0 ;
      RECT  11300.0 19910.0 11165.0 19980.0 ;
      RECT  11300.0 19910.0 11165.0 19980.0 ;
      RECT  13590.0 19980.0 13725.0 19910.0 ;
      RECT  11300.0 22600.0 11165.0 22670.0 ;
      RECT  11300.0 22600.0 11165.0 22670.0 ;
      RECT  13590.0 22670.0 13725.0 22600.0 ;
      RECT  11300.0 25290.0 11165.0 25360.0 ;
      RECT  11300.0 25290.0 11165.0 25360.0 ;
      RECT  13590.0 25360.0 13725.0 25290.0 ;
      RECT  12735.0 26010.0 12600.0 26080.0 ;
      RECT  12940.0 25870.0 12805.0 25940.0 ;
      RECT  13145.0 25730.0 13010.0 25800.0 ;
      RECT  13350.0 25590.0 13215.0 25660.0 ;
      RECT  12735.0 627.5 12600.0 697.5 ;
      RECT  12940.0 2062.5 12805.0 2132.5 ;
      RECT  13145.0 3317.5 13010.0 3387.5 ;
      RECT  13350.0 4752.5 13215.0 4822.5 ;
      RECT  13657.5 70.0 13792.5 2.49800180541e-13 ;
      RECT  13657.5 2760.0 13792.5 2690.0 ;
      RECT  13657.5 5450.0 13792.5 5380.0 ;
      RECT  11162.5 6847.5 11027.5 6917.5 ;
      RECT  6720.0 5207.5 6790.0 5342.5 ;
      RECT  11162.5 6142.5 11027.5 6212.5 ;
      RECT  6995.0 5207.5 7065.0 5342.5 ;
      RECT  11162.5 11077.5 11027.5 11147.5 ;
      RECT  11505.0 11077.5 11370.0 11147.5 ;
      RECT  11162.5 10372.5 11027.5 10442.5 ;
      RECT  11710.0 10372.5 11575.0 10442.5 ;
      RECT  11162.5 9667.5 11027.5 9737.5 ;
      RECT  11915.0 9667.5 11780.0 9737.5 ;
      RECT  11162.5 8962.5 11027.5 9032.5 ;
      RECT  12120.0 8962.5 11985.0 9032.5 ;
      RECT  11162.5 8257.5 11027.5 8327.5 ;
      RECT  12325.0 8257.5 12190.0 8327.5 ;
      RECT  11162.5 7552.5 11027.5 7622.5 ;
      RECT  12530.0 7552.5 12395.0 7622.5 ;
      RECT  11230.0 11430.0 11095.0 11500.0 ;
      RECT  13792.5 11430.0 13657.5 11500.0 ;
      RECT  11230.0 10725.0 11095.0 10795.0 ;
      RECT  13792.5 10725.0 13657.5 10795.0 ;
      RECT  11230.0 10020.0 11095.0 10090.0 ;
      RECT  13792.5 10020.0 13657.5 10090.0 ;
      RECT  11230.0 9315.0 11095.0 9385.0 ;
      RECT  13792.5 9315.0 13657.5 9385.0 ;
      RECT  11230.0 8610.0 11095.0 8680.0 ;
      RECT  13792.5 8610.0 13657.5 8680.0 ;
      RECT  11230.0 7905.0 11095.0 7975.0 ;
      RECT  13792.5 7905.0 13657.5 7975.0 ;
      RECT  11230.0 7200.0 11095.0 7270.0 ;
      RECT  13792.5 7200.0 13657.5 7270.0 ;
      RECT  11230.0 6495.0 11095.0 6565.0 ;
      RECT  13792.5 6495.0 13657.5 6565.0 ;
      RECT  11230.0 5790.0 11095.0 5860.0 ;
      RECT  13792.5 5790.0 13657.5 5860.0 ;
      RECT  14930.0 9872.5 14795.0 9942.5 ;
      RECT  14520.0 7687.5 14385.0 7757.5 ;
      RECT  14725.0 9235.0 14590.0 9305.0 ;
      RECT  14930.0 115070.0 14795.0 115140.0 ;
      RECT  15135.0 16375.0 15000.0 16445.0 ;
      RECT  15340.0 20400.0 15205.0 20470.0 ;
      RECT  14315.0 11635.0 14180.0 11705.0 ;
      RECT  8997.5 114265.0 8862.5 114335.0 ;
      RECT  14315.0 114265.0 14180.0 114335.0 ;
      RECT  14007.5 9105.0 13872.5 9175.0 ;
      RECT  14007.5 20530.0 13872.5 20600.0 ;
      RECT  14007.5 10032.5 13872.5 10102.5 ;
      RECT  14007.5 17307.5 13872.5 17377.5 ;
      RECT  16067.5 35.0 16137.5 175.0 ;
      RECT  18887.5 35.0 18957.5 175.0 ;
      RECT  21707.5 35.0 21777.5 175.0 ;
      RECT  24527.5 35.0 24597.5 175.0 ;
      RECT  27347.5 35.0 27417.5 175.0 ;
      RECT  30167.5 35.0 30237.5 175.0 ;
      RECT  32987.5 35.0 33057.5 175.0 ;
      RECT  35807.5 35.0 35877.5 175.0 ;
      RECT  38627.5 35.0 38697.5 175.0 ;
      RECT  41447.5 35.0 41517.5 175.0 ;
      RECT  44267.5 35.0 44337.5 175.0 ;
      RECT  47087.5 35.0 47157.5 175.0 ;
      RECT  49907.5 35.0 49977.5 175.0 ;
      RECT  52727.5 35.0 52797.5 175.0 ;
      RECT  55547.5 35.0 55617.5 175.0 ;
      RECT  58367.5 35.0 58437.5 175.0 ;
      RECT  61187.5 35.0 61257.5 175.0 ;
      RECT  64007.5 35.0 64077.5 175.0 ;
      RECT  66827.5 35.0 66897.5 175.0 ;
      RECT  69647.5 35.0 69717.5 175.0 ;
      RECT  72467.5 35.0 72537.5 175.0 ;
      RECT  75287.5 35.0 75357.5 175.0 ;
      RECT  78107.5 35.0 78177.5 175.0 ;
      RECT  80927.5 35.0 80997.5 175.0 ;
      RECT  83747.5 35.0 83817.5 175.0 ;
      RECT  86567.5 35.0 86637.5 175.0 ;
      RECT  89387.5 35.0 89457.5 175.0 ;
      RECT  92207.5 35.0 92277.5 175.0 ;
      RECT  95027.5 35.0 95097.5 175.0 ;
      RECT  97847.5 35.0 97917.5 175.0 ;
      RECT  100667.5 35.0 100737.5 175.0 ;
      RECT  103487.5 35.0 103557.5 175.0 ;
      RECT  15237.5 35.0 15307.5 115822.5 ;
      RECT  15032.5 35.0 15102.5 115822.5 ;
      RECT  14417.5 35.0 14487.5 115822.5 ;
      RECT  14622.5 35.0 14692.5 115822.5 ;
      RECT  14827.5 35.0 14897.5 115822.5 ;
      RECT  14212.5 35.0 14282.5 115822.5 ;
      RECT  13657.5 35.0 14007.5 115822.5 ;
      RECT  4035.0 35415.0 8.881784197e-13 35485.0 ;
      RECT  4035.0 35620.0 8.881784197e-13 35690.0 ;
      RECT  4035.0 35825.0 8.881784197e-13 35895.0 ;
      RECT  4035.0 36235.0 8.881784197e-13 36305.0 ;
      RECT  3422.5 30925.0 2690.0 30995.0 ;
      RECT  2520.0 28392.5 2450.0 35040.0 ;
      RECT  4035.0 35210.0 3830.0 35280.0 ;
      RECT  2895.0 36030.0 2690.0 36100.0 ;
      RECT  1550.0 35210.0 1345.0 35280.0 ;
      RECT  205.0 36030.0 8.881784197e-13 36100.0 ;
      RECT  165.0 28155.0 870.0 34595.0 ;
      RECT  1575.0 28155.0 870.0 34595.0 ;
      RECT  1575.0 28155.0 2280.0 34595.0 ;
      RECT  482.5 28155.0 552.5 28300.0 ;
      RECT  1187.5 28155.0 1257.5 28300.0 ;
      RECT  1892.5 28155.0 1962.5 28300.0 ;
      RECT  482.5 34325.0 552.5 34595.0 ;
      RECT  327.5 33907.5 397.5 34595.0 ;
      RECT  1187.5 34325.0 1257.5 34595.0 ;
      RECT  1342.5 33907.5 1412.5 34595.0 ;
      RECT  1892.5 34325.0 1962.5 34595.0 ;
      RECT  1737.5 33907.5 1807.5 34595.0 ;
      RECT  130.0 28155.0 200.0 34595.0 ;
      RECT  835.0 28155.0 905.0 34595.0 ;
      RECT  1540.0 28155.0 1610.0 34595.0 ;
      RECT  2245.0 28155.0 2315.0 34595.0 ;
      RECT  3737.5 37485.0 3032.5 37555.0 ;
      RECT  3382.5 37105.0 3312.5 37175.0 ;
      RECT  3382.5 37485.0 3312.5 37555.0 ;
      RECT  3347.5 37105.0 3032.5 37175.0 ;
      RECT  3382.5 37140.0 3312.5 37520.0 ;
      RECT  3737.5 37485.0 3347.5 37555.0 ;
      RECT  3032.5 37105.0 2897.5 37175.0 ;
      RECT  3032.5 37485.0 2897.5 37555.0 ;
      RECT  3872.5 37485.0 3737.5 37555.0 ;
      RECT  3415.0 37485.0 3280.0 37555.0 ;
      RECT  1895.0 37295.0 1965.0 37365.0 ;
      RECT  1930.0 37295.0 2280.0 37365.0 ;
      RECT  1895.0 37330.0 1965.0 37400.0 ;
      RECT  1495.0 37295.0 1565.0 37365.0 ;
      RECT  1495.0 37172.5 1565.0 37330.0 ;
      RECT  1530.0 37295.0 1930.0 37365.0 ;
      RECT  2280.0 37295.0 2415.0 37365.0 ;
      RECT  1495.0 37207.5 1565.0 37072.5 ;
      RECT  1895.0 37467.5 1965.0 37332.5 ;
      RECT  1950.0 38250.0 2020.0 38320.0 ;
      RECT  1950.0 38440.0 2020.0 38510.0 ;
      RECT  1985.0 38250.0 2347.5 38320.0 ;
      RECT  1950.0 38285.0 2020.0 38475.0 ;
      RECT  1642.5 38440.0 1985.0 38510.0 ;
      RECT  2347.5 38250.0 2482.5 38320.0 ;
      RECT  1507.5 38440.0 1642.5 38510.0 ;
      RECT  1950.0 38542.5 2020.0 38407.5 ;
      RECT  1047.5 38045.0 342.5 38115.0 ;
      RECT  692.5 37665.0 622.5 37735.0 ;
      RECT  692.5 38045.0 622.5 38115.0 ;
      RECT  657.5 37665.0 342.5 37735.0 ;
      RECT  692.5 37700.0 622.5 38080.0 ;
      RECT  1047.5 38045.0 657.5 38115.0 ;
      RECT  342.5 37665.0 207.5 37735.0 ;
      RECT  342.5 38045.0 207.5 38115.0 ;
      RECT  1182.5 38045.0 1047.5 38115.0 ;
      RECT  725.0 38045.0 590.0 38115.0 ;
      RECT  397.5 34662.5 327.5 34527.5 ;
      RECT  397.5 36337.5 327.5 36202.5 ;
      RECT  552.5 34662.5 482.5 34527.5 ;
      RECT  552.5 35517.5 482.5 35382.5 ;
      RECT  1412.5 34662.5 1342.5 34527.5 ;
      RECT  1412.5 35722.5 1342.5 35587.5 ;
      RECT  1807.5 34662.5 1737.5 34527.5 ;
      RECT  1807.5 35927.5 1737.5 35792.5 ;
      RECT  200.0 34662.5 130.0 34527.5 ;
      RECT  200.0 35312.5 130.0 35177.5 ;
      RECT  905.0 34662.5 835.0 34527.5 ;
      RECT  905.0 35312.5 835.0 35177.5 ;
      RECT  1610.0 34662.5 1540.0 34527.5 ;
      RECT  1610.0 35312.5 1540.0 35177.5 ;
      RECT  2315.0 34662.5 2245.0 34527.5 ;
      RECT  2315.0 35312.5 2245.0 35177.5 ;
      RECT  1380.0 40820.0 1310.0 60675.0 ;
      RECT  970.0 40820.0 900.0 60365.0 ;
      RECT  265.0 40820.0 195.0 60365.0 ;
      RECT  1207.5 40987.5 1137.5 41585.0 ;
      RECT  785.0 40987.5 715.0 41267.5 ;
      RECT  3372.5 43382.5 3442.5 43777.5 ;
      RECT  3372.5 43777.5 3442.5 44337.5 ;
      RECT  3372.5 44337.5 3442.5 44897.5 ;
      RECT  3372.5 45062.5 3442.5 45457.5 ;
      RECT  3372.5 45457.5 3442.5 46017.5 ;
      RECT  3372.5 46017.5 3442.5 46577.5 ;
      RECT  2655.0 46707.5 2725.0 46777.5 ;
      RECT  2655.0 46227.5 2725.0 46297.5 ;
      RECT  2690.0 46707.5 3407.5 46777.5 ;
      RECT  2655.0 46262.5 2725.0 46742.5 ;
      RECT  1972.5 46227.5 2690.0 46297.5 ;
      RECT  1937.5 45702.5 2007.5 46262.5 ;
      RECT  1937.5 45142.5 2007.5 45702.5 ;
      RECT  1937.5 44582.5 2007.5 44977.5 ;
      RECT  1937.5 44022.5 2007.5 44582.5 ;
      RECT  1937.5 43462.5 2007.5 44022.5 ;
      RECT  3340.0 43742.5 3475.0 43812.5 ;
      RECT  3340.0 44302.5 3475.0 44372.5 ;
      RECT  3340.0 44862.5 3475.0 44932.5 ;
      RECT  3340.0 45422.5 3475.0 45492.5 ;
      RECT  3340.0 45982.5 3475.0 46052.5 ;
      RECT  3340.0 46542.5 3475.0 46612.5 ;
      RECT  1905.0 46227.5 2040.0 46297.5 ;
      RECT  1905.0 45667.5 2040.0 45737.5 ;
      RECT  1905.0 45107.5 2040.0 45177.5 ;
      RECT  1905.0 44547.5 2040.0 44617.5 ;
      RECT  1905.0 43987.5 2040.0 44057.5 ;
      RECT  1905.0 43427.5 2040.0 43497.5 ;
      RECT  3340.0 43347.5 3475.0 43417.5 ;
      RECT  3340.0 45027.5 3475.0 45097.5 ;
      RECT  3340.0 46707.5 3475.0 46777.5 ;
      RECT  1905.0 44942.5 2040.0 45012.5 ;
      RECT  935.0 42725.0 225.0 41380.0 ;
      RECT  935.0 42725.0 230.0 44070.0 ;
      RECT  935.0 45415.0 230.0 44070.0 ;
      RECT  935.0 45415.0 230.0 46760.0 ;
      RECT  935.0 48105.0 230.0 46760.0 ;
      RECT  935.0 48105.0 230.0 49450.0 ;
      RECT  935.0 50795.0 230.0 49450.0 ;
      RECT  935.0 50795.0 230.0 52140.0 ;
      RECT  935.0 53485.0 230.0 52140.0 ;
      RECT  935.0 53485.0 230.0 54830.0 ;
      RECT  935.0 56175.0 230.0 54830.0 ;
      RECT  935.0 56175.0 230.0 57520.0 ;
      RECT  935.0 58865.0 230.0 57520.0 ;
      RECT  935.0 58865.0 230.0 60210.0 ;
      RECT  785.0 42625.0 715.0 60365.0 ;
      RECT  450.0 42625.0 380.0 60365.0 ;
      RECT  970.0 42625.0 900.0 60365.0 ;
      RECT  265.0 42625.0 195.0 60365.0 ;
      RECT  1347.5 42797.5 1277.5 42932.5 ;
      RECT  1347.5 45207.5 1277.5 45342.5 ;
      RECT  1347.5 45487.5 1277.5 45622.5 ;
      RECT  1347.5 47897.5 1277.5 48032.5 ;
      RECT  1347.5 48177.5 1277.5 48312.5 ;
      RECT  1347.5 50587.5 1277.5 50722.5 ;
      RECT  1347.5 50867.5 1277.5 51002.5 ;
      RECT  1347.5 53277.5 1277.5 53412.5 ;
      RECT  1347.5 53557.5 1277.5 53692.5 ;
      RECT  1347.5 55967.5 1277.5 56102.5 ;
      RECT  1347.5 56247.5 1277.5 56382.5 ;
      RECT  1347.5 58657.5 1277.5 58792.5 ;
      RECT  1347.5 58937.5 1277.5 59072.5 ;
      RECT  1345.0 43060.0 1275.0 43195.0 ;
      RECT  1380.0 40685.0 1310.0 40820.0 ;
      RECT  867.5 40785.0 1002.5 40855.0 ;
      RECT  162.5 40785.0 297.5 40855.0 ;
      RECT  1105.0 41550.0 1240.0 41620.0 ;
      RECT  1105.0 40952.5 1240.0 41022.5 ;
      RECT  682.5 40952.5 817.5 41022.5 ;
      RECT  3457.5 35107.5 3387.5 34972.5 ;
      RECT  3457.5 31027.5 3387.5 30892.5 ;
      RECT  2725.0 31027.5 2655.0 30892.5 ;
      RECT  2725.0 36542.5 2655.0 36407.5 ;
      RECT  2520.0 28460.0 2450.0 28325.0 ;
      RECT  1965.0 35107.5 1895.0 34972.5 ;
      RECT  1750.0 35517.5 1680.0 35382.5 ;
      RECT  2020.0 38055.0 1950.0 37920.0 ;
      RECT  2020.0 38055.0 1950.0 37920.0 ;
      RECT  2020.0 36542.5 1950.0 36407.5 ;
      RECT  1805.0 38312.5 1735.0 38177.5 ;
      RECT  1805.0 38312.5 1735.0 38177.5 ;
      RECT  1805.0 36337.5 1735.0 36202.5 ;
      RECT  3382.5 36542.5 3312.5 36407.5 ;
      RECT  3522.5 36337.5 3452.5 36202.5 ;
      RECT  3662.5 35722.5 3592.5 35587.5 ;
      RECT  692.5 36542.5 622.5 36407.5 ;
      RECT  832.5 35722.5 762.5 35587.5 ;
      RECT  972.5 35927.5 902.5 35792.5 ;
      RECT  1997.5 37735.0 1862.5 37805.0 ;
      RECT  2052.5 38880.0 1917.5 38950.0 ;
      RECT  785.0 40065.0 650.0 40135.0 ;
      RECT  2040.0 39105.0 1905.0 39175.0 ;
      RECT  4070.0 35312.5 4000.0 35177.5 ;
      RECT  2725.0 36132.5 2655.0 35997.5 ;
      RECT  1380.0 35312.5 1310.0 35177.5 ;
      RECT  35.0 36132.5 -35.0 35997.5 ;
      RECT  4035.0 39105.0 1972.5 39175.0 ;
      RECT  4035.0 40065.0 717.5 40135.0 ;
      RECT  4035.0 37735.0 1930.0 37805.0 ;
      RECT  4035.0 38880.0 1985.0 38950.0 ;
      RECT  4035.0 36440.0 8.881784197e-13 36510.0 ;
      RECT  4035.0 35005.0 0.0 35075.0 ;
      RECT  4035.0 36030.0 8.881784197e-13 36100.0 ;
      RECT  4035.0 35210.0 0.0 35280.0 ;
      RECT  15340.0 39105.0 15205.0 39175.0 ;
      RECT  4035.0 39105.0 3900.0 39175.0 ;
      RECT  15135.0 40065.0 15000.0 40135.0 ;
      RECT  4035.0 40065.0 3900.0 40135.0 ;
      RECT  14725.0 37735.0 14590.0 37805.0 ;
      RECT  4035.0 37735.0 3900.0 37805.0 ;
      RECT  14520.0 38880.0 14385.0 38950.0 ;
      RECT  4035.0 38880.0 3900.0 38950.0 ;
      RECT  14930.0 36440.0 14795.0 36510.0 ;
      RECT  4035.0 36440.0 3900.0 36510.0 ;
      RECT  14315.0 35005.0 14180.0 35075.0 ;
      RECT  4035.0 35005.0 3900.0 35075.0 ;
      RECT  4417.5 36030.0 4282.5 36100.0 ;
      RECT  13900.0 35210.0 13765.0 35280.0 ;
      RECT  4035.0 35210.0 3900.0 35280.0 ;
   LAYER  metal3 ;
      RECT  4035.0 39105.0 15272.5 39175.0 ;
      RECT  4035.0 40065.0 15067.5 40135.0 ;
      RECT  4035.0 37735.0 14657.5 37805.0 ;
      RECT  4035.0 38880.0 14452.5 38950.0 ;
      RECT  4035.0 36440.0 14862.5 36510.0 ;
      RECT  4035.0 35005.0 14247.5 35075.0 ;
      RECT  4035.0 35210.0 13832.5 35280.0 ;
      RECT  15857.5 25065.0 15927.5 25135.0 ;
      RECT  15857.5 6555.0 15927.5 25100.0 ;
      RECT  15892.5 25065.0 16062.5 25135.0 ;
      RECT  18677.5 25065.0 18747.5 25135.0 ;
      RECT  18677.5 6555.0 18747.5 25100.0 ;
      RECT  18712.5 25065.0 18882.5 25135.0 ;
      RECT  21497.5 25065.0 21567.5 25135.0 ;
      RECT  21497.5 6555.0 21567.5 25100.0 ;
      RECT  21532.5 25065.0 21702.5 25135.0 ;
      RECT  24317.5 25065.0 24387.5 25135.0 ;
      RECT  24317.5 6555.0 24387.5 25100.0 ;
      RECT  24352.5 25065.0 24522.5 25135.0 ;
      RECT  27137.5 25065.0 27207.5 25135.0 ;
      RECT  27137.5 6555.0 27207.5 25100.0 ;
      RECT  27172.5 25065.0 27342.5 25135.0 ;
      RECT  29957.5 25065.0 30027.5 25135.0 ;
      RECT  29957.5 6555.0 30027.5 25100.0 ;
      RECT  29992.5 25065.0 30162.5 25135.0 ;
      RECT  32777.5 25065.0 32847.5 25135.0 ;
      RECT  32777.5 6555.0 32847.5 25100.0 ;
      RECT  32812.5 25065.0 32982.5 25135.0 ;
      RECT  35597.5 25065.0 35667.5 25135.0 ;
      RECT  35597.5 6555.0 35667.5 25100.0 ;
      RECT  35632.5 25065.0 35802.5 25135.0 ;
      RECT  38417.5 25065.0 38487.5 25135.0 ;
      RECT  38417.5 6555.0 38487.5 25100.0 ;
      RECT  38452.5 25065.0 38622.5 25135.0 ;
      RECT  41237.5 25065.0 41307.5 25135.0 ;
      RECT  41237.5 6555.0 41307.5 25100.0 ;
      RECT  41272.5 25065.0 41442.5 25135.0 ;
      RECT  44057.5 25065.0 44127.5 25135.0 ;
      RECT  44057.5 6555.0 44127.5 25100.0 ;
      RECT  44092.5 25065.0 44262.5 25135.0 ;
      RECT  46877.5 25065.0 46947.5 25135.0 ;
      RECT  46877.5 6555.0 46947.5 25100.0 ;
      RECT  46912.5 25065.0 47082.5 25135.0 ;
      RECT  49697.5 25065.0 49767.5 25135.0 ;
      RECT  49697.5 6555.0 49767.5 25100.0 ;
      RECT  49732.5 25065.0 49902.5 25135.0 ;
      RECT  52517.5 25065.0 52587.5 25135.0 ;
      RECT  52517.5 6555.0 52587.5 25100.0 ;
      RECT  52552.5 25065.0 52722.5 25135.0 ;
      RECT  55337.5 25065.0 55407.5 25135.0 ;
      RECT  55337.5 6555.0 55407.5 25100.0 ;
      RECT  55372.5 25065.0 55542.5 25135.0 ;
      RECT  58157.5 25065.0 58227.5 25135.0 ;
      RECT  58157.5 6555.0 58227.5 25100.0 ;
      RECT  58192.5 25065.0 58362.5 25135.0 ;
      RECT  60977.5 25065.0 61047.5 25135.0 ;
      RECT  60977.5 6555.0 61047.5 25100.0 ;
      RECT  61012.5 25065.0 61182.5 25135.0 ;
      RECT  63797.5 25065.0 63867.5 25135.0 ;
      RECT  63797.5 6555.0 63867.5 25100.0 ;
      RECT  63832.5 25065.0 64002.5 25135.0 ;
      RECT  66617.5 25065.0 66687.5 25135.0 ;
      RECT  66617.5 6555.0 66687.5 25100.0 ;
      RECT  66652.5 25065.0 66822.5 25135.0 ;
      RECT  69437.5 25065.0 69507.5 25135.0 ;
      RECT  69437.5 6555.0 69507.5 25100.0 ;
      RECT  69472.5 25065.0 69642.5 25135.0 ;
      RECT  72257.5 25065.0 72327.5 25135.0 ;
      RECT  72257.5 6555.0 72327.5 25100.0 ;
      RECT  72292.5 25065.0 72462.5 25135.0 ;
      RECT  75077.5 25065.0 75147.5 25135.0 ;
      RECT  75077.5 6555.0 75147.5 25100.0 ;
      RECT  75112.5 25065.0 75282.5 25135.0 ;
      RECT  77897.5 25065.0 77967.5 25135.0 ;
      RECT  77897.5 6555.0 77967.5 25100.0 ;
      RECT  77932.5 25065.0 78102.5 25135.0 ;
      RECT  80717.5 25065.0 80787.5 25135.0 ;
      RECT  80717.5 6555.0 80787.5 25100.0 ;
      RECT  80752.5 25065.0 80922.5 25135.0 ;
      RECT  83537.5 25065.0 83607.5 25135.0 ;
      RECT  83537.5 6555.0 83607.5 25100.0 ;
      RECT  83572.5 25065.0 83742.5 25135.0 ;
      RECT  86357.5 25065.0 86427.5 25135.0 ;
      RECT  86357.5 6555.0 86427.5 25100.0 ;
      RECT  86392.5 25065.0 86562.5 25135.0 ;
      RECT  89177.5 25065.0 89247.5 25135.0 ;
      RECT  89177.5 6555.0 89247.5 25100.0 ;
      RECT  89212.5 25065.0 89382.5 25135.0 ;
      RECT  91997.5 25065.0 92067.5 25135.0 ;
      RECT  91997.5 6555.0 92067.5 25100.0 ;
      RECT  92032.5 25065.0 92202.5 25135.0 ;
      RECT  94817.5 25065.0 94887.5 25135.0 ;
      RECT  94817.5 6555.0 94887.5 25100.0 ;
      RECT  94852.5 25065.0 95022.5 25135.0 ;
      RECT  97637.5 25065.0 97707.5 25135.0 ;
      RECT  97637.5 6555.0 97707.5 25100.0 ;
      RECT  97672.5 25065.0 97842.5 25135.0 ;
      RECT  100457.5 25065.0 100527.5 25135.0 ;
      RECT  100457.5 6555.0 100527.5 25100.0 ;
      RECT  100492.5 25065.0 100662.5 25135.0 ;
      RECT  103277.5 25065.0 103347.5 25135.0 ;
      RECT  103277.5 6555.0 103347.5 25100.0 ;
      RECT  103312.5 25065.0 103482.5 25135.0 ;
      RECT  16067.5 35.0 16137.5 9670.0 ;
      RECT  18887.5 35.0 18957.5 9670.0 ;
      RECT  21707.5 35.0 21777.5 9670.0 ;
      RECT  24527.5 35.0 24597.5 9670.0 ;
      RECT  27347.5 35.0 27417.5 9670.0 ;
      RECT  30167.5 35.0 30237.5 9670.0 ;
      RECT  32987.5 35.0 33057.5 9670.0 ;
      RECT  35807.5 35.0 35877.5 9670.0 ;
      RECT  38627.5 35.0 38697.5 9670.0 ;
      RECT  41447.5 35.0 41517.5 9670.0 ;
      RECT  44267.5 35.0 44337.5 9670.0 ;
      RECT  47087.5 35.0 47157.5 9670.0 ;
      RECT  49907.5 35.0 49977.5 9670.0 ;
      RECT  52727.5 35.0 52797.5 9670.0 ;
      RECT  55547.5 35.0 55617.5 9670.0 ;
      RECT  58367.5 35.0 58437.5 9670.0 ;
      RECT  61187.5 35.0 61257.5 9670.0 ;
      RECT  64007.5 35.0 64077.5 9670.0 ;
      RECT  66827.5 35.0 66897.5 9670.0 ;
      RECT  69647.5 35.0 69717.5 9670.0 ;
      RECT  72467.5 35.0 72537.5 9670.0 ;
      RECT  75287.5 35.0 75357.5 9670.0 ;
      RECT  78107.5 35.0 78177.5 9670.0 ;
      RECT  80927.5 35.0 80997.5 9670.0 ;
      RECT  83747.5 35.0 83817.5 9670.0 ;
      RECT  86567.5 35.0 86637.5 9670.0 ;
      RECT  89387.5 35.0 89457.5 9670.0 ;
      RECT  92207.5 35.0 92277.5 9670.0 ;
      RECT  95027.5 35.0 95097.5 9670.0 ;
      RECT  97847.5 35.0 97917.5 9670.0 ;
      RECT  100667.5 35.0 100737.5 9670.0 ;
      RECT  103487.5 35.0 103557.5 9670.0 ;
      RECT  11232.5 11840.0 13657.5 11910.0 ;
      RECT  11232.5 14530.0 13657.5 14600.0 ;
      RECT  11232.5 17220.0 13657.5 17290.0 ;
      RECT  11232.5 19910.0 13657.5 19980.0 ;
      RECT  11232.5 22600.0 13657.5 22670.0 ;
      RECT  11232.5 25290.0 13657.5 25360.0 ;
      RECT  6720.0 6847.5 6790.0 6917.5 ;
      RECT  6755.0 6847.5 11095.0 6917.5 ;
      RECT  6720.0 5275.0 6790.0 6882.5 ;
      RECT  6995.0 6142.5 7065.0 6212.5 ;
      RECT  7030.0 6142.5 11095.0 6212.5 ;
      RECT  6995.0 5275.0 7065.0 6177.5 ;
      RECT  16062.5 25030.0 16132.5 25170.0 ;
      RECT  18882.5 25030.0 18952.5 25170.0 ;
      RECT  21702.5 25030.0 21772.5 25170.0 ;
      RECT  24522.5 25030.0 24592.5 25170.0 ;
      RECT  27342.5 25030.0 27412.5 25170.0 ;
      RECT  30162.5 25030.0 30232.5 25170.0 ;
      RECT  32982.5 25030.0 33052.5 25170.0 ;
      RECT  35802.5 25030.0 35872.5 25170.0 ;
      RECT  38622.5 25030.0 38692.5 25170.0 ;
      RECT  41442.5 25030.0 41512.5 25170.0 ;
      RECT  44262.5 25030.0 44332.5 25170.0 ;
      RECT  47082.5 25030.0 47152.5 25170.0 ;
      RECT  49902.5 25030.0 49972.5 25170.0 ;
      RECT  52722.5 25030.0 52792.5 25170.0 ;
      RECT  55542.5 25030.0 55612.5 25170.0 ;
      RECT  58362.5 25030.0 58432.5 25170.0 ;
      RECT  61182.5 25030.0 61252.5 25170.0 ;
      RECT  64002.5 25030.0 64072.5 25170.0 ;
      RECT  66822.5 25030.0 66892.5 25170.0 ;
      RECT  69642.5 25030.0 69712.5 25170.0 ;
      RECT  72462.5 25030.0 72532.5 25170.0 ;
      RECT  75282.5 25030.0 75352.5 25170.0 ;
      RECT  78102.5 25030.0 78172.5 25170.0 ;
      RECT  80922.5 25030.0 80992.5 25170.0 ;
      RECT  83742.5 25030.0 83812.5 25170.0 ;
      RECT  86562.5 25030.0 86632.5 25170.0 ;
      RECT  89382.5 25030.0 89452.5 25170.0 ;
      RECT  92202.5 25030.0 92272.5 25170.0 ;
      RECT  95022.5 25030.0 95092.5 25170.0 ;
      RECT  97842.5 25030.0 97912.5 25170.0 ;
      RECT  100662.5 25030.0 100732.5 25170.0 ;
      RECT  103482.5 25030.0 103552.5 25170.0 ;
      RECT  16067.5 9670.0 16137.5 9810.0 ;
      RECT  18887.5 9670.0 18957.5 9810.0 ;
      RECT  21707.5 9670.0 21777.5 9810.0 ;
      RECT  24527.5 9670.0 24597.5 9810.0 ;
      RECT  27347.5 9670.0 27417.5 9810.0 ;
      RECT  30167.5 9670.0 30237.5 9810.0 ;
      RECT  32987.5 9670.0 33057.5 9810.0 ;
      RECT  35807.5 9670.0 35877.5 9810.0 ;
      RECT  38627.5 9670.0 38697.5 9810.0 ;
      RECT  41447.5 9670.0 41517.5 9810.0 ;
      RECT  44267.5 9670.0 44337.5 9810.0 ;
      RECT  47087.5 9670.0 47157.5 9810.0 ;
      RECT  49907.5 9670.0 49977.5 9810.0 ;
      RECT  52727.5 9670.0 52797.5 9810.0 ;
      RECT  55547.5 9670.0 55617.5 9810.0 ;
      RECT  58367.5 9670.0 58437.5 9810.0 ;
      RECT  61187.5 9670.0 61257.5 9810.0 ;
      RECT  64007.5 9670.0 64077.5 9810.0 ;
      RECT  66827.5 9670.0 66897.5 9810.0 ;
      RECT  69647.5 9670.0 69717.5 9810.0 ;
      RECT  72467.5 9670.0 72537.5 9810.0 ;
      RECT  75287.5 9670.0 75357.5 9810.0 ;
      RECT  78107.5 9670.0 78177.5 9810.0 ;
      RECT  80927.5 9670.0 80997.5 9810.0 ;
      RECT  83747.5 9670.0 83817.5 9810.0 ;
      RECT  86567.5 9670.0 86637.5 9810.0 ;
      RECT  89387.5 9670.0 89457.5 9810.0 ;
      RECT  92207.5 9670.0 92277.5 9810.0 ;
      RECT  95027.5 9670.0 95097.5 9810.0 ;
      RECT  97847.5 9670.0 97917.5 9810.0 ;
      RECT  100667.5 9670.0 100737.5 9810.0 ;
      RECT  103487.5 9670.0 103557.5 9810.0 ;
      RECT  4655.0 11147.5 4795.0 11077.5 ;
      RECT  4655.0 10442.5 4795.0 10372.5 ;
      RECT  4655.0 9737.5 4795.0 9667.5 ;
      RECT  4655.0 9032.5 4795.0 8962.5 ;
      RECT  4655.0 8327.5 4795.0 8257.5 ;
      RECT  4655.0 7622.5 4795.0 7552.5 ;
      RECT  4655.0 6917.5 4795.0 6847.5 ;
      RECT  4655.0 6212.5 4795.0 6142.5 ;
      RECT  15857.5 6520.0 15927.5 6655.0 ;
      RECT  18677.5 6520.0 18747.5 6655.0 ;
      RECT  21497.5 6520.0 21567.5 6655.0 ;
      RECT  24317.5 6520.0 24387.5 6655.0 ;
      RECT  27137.5 6520.0 27207.5 6655.0 ;
      RECT  29957.5 6520.0 30027.5 6655.0 ;
      RECT  32777.5 6520.0 32847.5 6655.0 ;
      RECT  35597.5 6520.0 35667.5 6655.0 ;
      RECT  38417.5 6520.0 38487.5 6655.0 ;
      RECT  41237.5 6520.0 41307.5 6655.0 ;
      RECT  44057.5 6520.0 44127.5 6655.0 ;
      RECT  46877.5 6520.0 46947.5 6655.0 ;
      RECT  49697.5 6520.0 49767.5 6655.0 ;
      RECT  52517.5 6520.0 52587.5 6655.0 ;
      RECT  55337.5 6520.0 55407.5 6655.0 ;
      RECT  58157.5 6520.0 58227.5 6655.0 ;
      RECT  60977.5 6520.0 61047.5 6655.0 ;
      RECT  63797.5 6520.0 63867.5 6655.0 ;
      RECT  66617.5 6520.0 66687.5 6655.0 ;
      RECT  69437.5 6520.0 69507.5 6655.0 ;
      RECT  72257.5 6520.0 72327.5 6655.0 ;
      RECT  75077.5 6520.0 75147.5 6655.0 ;
      RECT  77897.5 6520.0 77967.5 6655.0 ;
      RECT  80717.5 6520.0 80787.5 6655.0 ;
      RECT  83537.5 6520.0 83607.5 6655.0 ;
      RECT  86357.5 6520.0 86427.5 6655.0 ;
      RECT  89177.5 6520.0 89247.5 6655.0 ;
      RECT  91997.5 6520.0 92067.5 6655.0 ;
      RECT  94817.5 6520.0 94887.5 6655.0 ;
      RECT  97637.5 6520.0 97707.5 6655.0 ;
      RECT  100457.5 6520.0 100527.5 6655.0 ;
      RECT  103277.5 6520.0 103347.5 6655.0 ;
      RECT  16067.5 35.0 16137.5 170.0 ;
      RECT  18887.5 35.0 18957.5 170.0 ;
      RECT  21707.5 35.0 21777.5 170.0 ;
      RECT  24527.5 35.0 24597.5 170.0 ;
      RECT  27347.5 35.0 27417.5 170.0 ;
      RECT  30167.5 35.0 30237.5 170.0 ;
      RECT  32987.5 35.0 33057.5 170.0 ;
      RECT  35807.5 35.0 35877.5 170.0 ;
      RECT  38627.5 35.0 38697.5 170.0 ;
      RECT  41447.5 35.0 41517.5 170.0 ;
      RECT  44267.5 35.0 44337.5 170.0 ;
      RECT  47087.5 35.0 47157.5 170.0 ;
      RECT  49907.5 35.0 49977.5 170.0 ;
      RECT  52727.5 35.0 52797.5 170.0 ;
      RECT  55547.5 35.0 55617.5 170.0 ;
      RECT  58367.5 35.0 58437.5 170.0 ;
      RECT  61187.5 35.0 61257.5 170.0 ;
      RECT  64007.5 35.0 64077.5 170.0 ;
      RECT  66827.5 35.0 66897.5 170.0 ;
      RECT  69647.5 35.0 69717.5 170.0 ;
      RECT  72467.5 35.0 72537.5 170.0 ;
      RECT  75287.5 35.0 75357.5 170.0 ;
      RECT  78107.5 35.0 78177.5 170.0 ;
      RECT  80927.5 35.0 80997.5 170.0 ;
      RECT  83747.5 35.0 83817.5 170.0 ;
      RECT  86567.5 35.0 86637.5 170.0 ;
      RECT  89387.5 35.0 89457.5 170.0 ;
      RECT  92207.5 35.0 92277.5 170.0 ;
      RECT  95027.5 35.0 95097.5 170.0 ;
      RECT  97847.5 35.0 97917.5 170.0 ;
      RECT  100667.5 35.0 100737.5 170.0 ;
      RECT  103487.5 35.0 103557.5 170.0 ;
      RECT  11300.0 11840.0 11165.0 11910.0 ;
      RECT  13590.0 11910.0 13725.0 11840.0 ;
      RECT  11300.0 14530.0 11165.0 14600.0 ;
      RECT  13590.0 14600.0 13725.0 14530.0 ;
      RECT  11300.0 17220.0 11165.0 17290.0 ;
      RECT  13590.0 17290.0 13725.0 17220.0 ;
      RECT  11300.0 19910.0 11165.0 19980.0 ;
      RECT  13590.0 19980.0 13725.0 19910.0 ;
      RECT  11300.0 22600.0 11165.0 22670.0 ;
      RECT  13590.0 22670.0 13725.0 22600.0 ;
      RECT  11300.0 25290.0 11165.0 25360.0 ;
      RECT  13590.0 25360.0 13725.0 25290.0 ;
      RECT  11162.5 6847.5 11027.5 6917.5 ;
      RECT  6720.0 5207.5 6790.0 5342.5 ;
      RECT  11162.5 6142.5 11027.5 6212.5 ;
      RECT  6995.0 5207.5 7065.0 5342.5 ;
      RECT  4175.0 11077.5 4655.0 11147.5 ;
      RECT  4175.0 10372.5 4655.0 10442.5 ;
      RECT  4175.0 9667.5 4655.0 9737.5 ;
      RECT  4175.0 8962.5 4655.0 9032.5 ;
      RECT  4175.0 8257.5 4655.0 8327.5 ;
      RECT  4175.0 7552.5 4655.0 7622.5 ;
      RECT  4175.0 6847.5 4655.0 6917.5 ;
      RECT  4175.0 6142.5 4655.0 6212.5 ;
      RECT  397.5 34595.0 327.5 36270.0 ;
      RECT  552.5 34595.0 482.5 35450.0 ;
      RECT  1412.5 34595.0 1342.5 35655.0 ;
      RECT  1807.5 34595.0 1737.5 35860.0 ;
      RECT  200.0 34595.0 130.0 35245.0 ;
      RECT  905.0 34595.0 835.0 35245.0 ;
      RECT  1610.0 34595.0 1540.0 35245.0 ;
      RECT  2315.0 34595.0 2245.0 35245.0 ;
      RECT  2725.0 30960.0 2655.0 36475.0 ;
      RECT  2020.0 36475.0 1950.0 37987.5 ;
      RECT  1805.0 36270.0 1735.0 38245.0 ;
      RECT  482.5 28155.0 552.5 28295.0 ;
      RECT  1187.5 28155.0 1257.5 28295.0 ;
      RECT  1892.5 28155.0 1962.5 28295.0 ;
      RECT  397.5 34662.5 327.5 34527.5 ;
      RECT  397.5 36337.5 327.5 36202.5 ;
      RECT  552.5 34662.5 482.5 34527.5 ;
      RECT  552.5 35517.5 482.5 35382.5 ;
      RECT  1412.5 34662.5 1342.5 34527.5 ;
      RECT  1412.5 35722.5 1342.5 35587.5 ;
      RECT  1807.5 34662.5 1737.5 34527.5 ;
      RECT  1807.5 35927.5 1737.5 35792.5 ;
      RECT  200.0 34662.5 130.0 34527.5 ;
      RECT  200.0 35312.5 130.0 35177.5 ;
      RECT  905.0 34662.5 835.0 34527.5 ;
      RECT  905.0 35312.5 835.0 35177.5 ;
      RECT  1610.0 34662.5 1540.0 34527.5 ;
      RECT  1610.0 35312.5 1540.0 35177.5 ;
      RECT  2315.0 34662.5 2245.0 34527.5 ;
      RECT  2315.0 35312.5 2245.0 35177.5 ;
      RECT  2725.0 31027.5 2655.0 30892.5 ;
      RECT  2725.0 36542.5 2655.0 36407.5 ;
      RECT  2020.0 38055.0 1950.0 37920.0 ;
      RECT  2020.0 36542.5 1950.0 36407.5 ;
      RECT  1805.0 38312.5 1735.0 38177.5 ;
      RECT  1805.0 36337.5 1735.0 36202.5 ;
      RECT  1257.5 28155.0 1187.5 28295.0 ;
      RECT  1962.5 28155.0 1892.5 28295.0 ;
      RECT  552.5 28155.0 482.5 28295.0 ;
      RECT  15340.0 39105.0 15205.0 39175.0 ;
      RECT  4035.0 39105.0 3900.0 39175.0 ;
      RECT  15135.0 40065.0 15000.0 40135.0 ;
      RECT  4035.0 40065.0 3900.0 40135.0 ;
      RECT  14725.0 37735.0 14590.0 37805.0 ;
      RECT  4035.0 37735.0 3900.0 37805.0 ;
      RECT  14520.0 38880.0 14385.0 38950.0 ;
      RECT  4035.0 38880.0 3900.0 38950.0 ;
      RECT  14930.0 36440.0 14795.0 36510.0 ;
      RECT  4035.0 36440.0 3900.0 36510.0 ;
      RECT  14315.0 35005.0 14180.0 35075.0 ;
      RECT  4035.0 35005.0 3900.0 35075.0 ;
      RECT  13900.0 35210.0 13765.0 35280.0 ;
      RECT  4035.0 35210.0 3900.0 35280.0 ;
   END
   END    sram_1rw_32b_256w_1bank_freepdk45
END    LIBRARY
