magic
tech scmos
timestamp 1523654621
<< nwell >>
rect 12 43 44 102
rect 12 -17 52 7
<< pwell >>
rect 12 102 44 131
rect 12 7 52 43
<< ntransistor >>
rect 23 119 25 125
rect 28 119 30 125
rect 23 29 25 35
rect 28 29 30 35
rect 23 13 25 17
rect 39 13 41 17
<< ptransistor >>
rect 23 84 25 96
rect 28 84 30 96
rect 23 50 25 62
rect 28 50 30 62
rect 23 -6 25 1
rect 39 -6 41 1
<< ndiffusion >>
rect 22 119 23 125
rect 25 119 28 125
rect 30 119 31 125
rect 22 29 23 35
rect 25 29 28 35
rect 30 29 31 35
rect 22 13 23 17
rect 25 13 26 17
rect 38 13 39 17
rect 41 13 42 17
<< pdiffusion >>
rect 22 84 23 96
rect 25 84 28 96
rect 30 84 31 96
rect 22 50 23 62
rect 25 50 28 62
rect 30 50 31 62
rect 22 -6 23 1
rect 25 -6 26 1
rect 38 -6 39 1
rect 41 -6 42 1
<< ndcontact >>
rect 18 119 22 125
rect 31 119 35 125
rect 18 29 22 35
rect 31 29 35 35
rect 18 13 22 17
rect 26 13 30 17
rect 34 13 38 17
rect 42 13 46 17
<< pdcontact >>
rect 18 84 22 96
rect 31 84 35 96
rect 18 50 22 62
rect 31 50 35 62
rect 18 -6 22 1
rect 26 -6 30 1
rect 34 -6 38 1
rect 42 -6 46 1
<< psubstratepcontact >>
rect 18 111 22 115
rect 26 21 30 25
rect 34 21 38 25
<< nsubstratencontact >>
rect 18 76 22 80
rect 18 66 22 70
rect 18 -14 22 -10
<< polysilicon >>
rect 23 125 25 127
rect 28 125 30 127
rect 23 107 25 119
rect 28 117 30 119
rect 28 115 40 117
rect 23 96 25 103
rect 28 96 30 98
rect 23 81 25 84
rect 23 62 25 64
rect 28 62 30 84
rect 23 35 25 50
rect 28 42 30 50
rect 38 38 40 115
rect 28 36 40 38
rect 28 35 30 36
rect 23 17 25 29
rect 28 28 30 29
rect 28 26 41 28
rect 39 17 41 26
rect 23 1 25 13
rect 39 1 41 13
rect 23 -8 25 -6
rect 23 -10 32 -8
rect 30 -25 32 -10
rect 39 -9 41 -6
rect 39 -11 43 -9
rect 41 -17 43 -11
<< polycontact >>
rect 22 103 26 107
rect 30 42 34 46
rect 41 -21 45 -17
rect 30 -29 34 -25
<< metal1 >>
rect 25 134 29 138
rect 25 130 35 134
rect 31 125 35 130
rect 18 110 22 111
rect 35 91 39 125
rect 42 84 46 125
rect 18 80 22 84
rect 18 70 22 72
rect 18 62 22 66
rect 41 80 46 84
rect 41 62 45 80
rect 35 58 45 62
rect 41 35 45 58
rect 35 31 45 35
rect 18 25 22 29
rect 18 21 26 25
rect 30 21 34 25
rect 38 21 47 25
rect 18 17 22 21
rect 26 8 30 13
rect 26 1 30 4
rect 46 13 47 17
rect 34 8 38 13
rect 34 1 38 4
rect 18 -10 22 -6
rect 42 -10 46 -6
rect 26 -14 46 -10
rect 16 -21 41 -17
rect 45 -21 49 -17
<< m2contact >>
rect 25 138 29 142
rect 42 125 46 129
rect 18 115 22 119
rect 26 103 30 107
rect 18 72 22 76
rect 34 41 38 45
rect 47 21 51 25
rect 26 4 30 8
rect 47 13 51 17
rect 34 4 38 8
rect 22 -14 26 -10
rect 30 -33 34 -29
<< metal2 >>
rect 25 142 29 162
rect 35 142 39 162
rect 35 138 46 142
rect 42 129 46 138
rect 18 114 22 115
rect 18 110 51 114
rect 18 -6 22 72
rect 26 8 30 103
rect 34 8 38 41
rect 47 25 51 110
rect 47 17 51 21
rect 18 -10 26 -6
rect 30 -40 34 -33
<< m3p >>
rect 15 -40 49 162
<< labels >>
rlabel metal1 19 -19 19 -19 1 en
rlabel metal2 27 161 27 161 5 bl
rlabel metal2 37 161 37 161 5 br
rlabel metal2 32 -38 32 -38 1 din
rlabel metal2 50 101 50 101 7 gnd
rlabel metal2 20 41 20 41 1 vdd
<< end >>
