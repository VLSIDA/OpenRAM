VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO sram_2_16_scn4m_subm
   CLASS BLOCK ;
   SIZE 209.1 BY 424.8 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  108.8 11.4 109.6 12.2 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  130.6 11.4 131.4 12.2 ;
      END
   END din0[1]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  65.2 353.4 66.0 354.2 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  65.2 375.4 66.0 376.2 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  65.2 393.4 66.0 394.2 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  65.2 415.4 66.0 416.2 ;
      END
   END addr0[3]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  10.0 11.4 10.8 12.2 ;
      END
   END csb0
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  10.0 33.4 10.8 34.2 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  54.1 12.3 54.7 12.9 ;
      END
   END clk0
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER m2 ;
         RECT  187.5 112.6 188.3 115.6 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER m2 ;
         RECT  194.3 112.6 195.1 115.6 ;
      END
   END dout0[1]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER m3 ;
         RECT  81.6 163.2 207.6 164.4 ;
         LAYER m3 ;
         RECT  0.0 67.2 207.6 68.4 ;
         LAYER m3 ;
         RECT  72.0 422.4 207.6 423.6 ;
         LAYER m3 ;
         RECT  0.0 153.6 75.6 154.8 ;
         LAYER m3 ;
         RECT  0.0 417.6 207.6 418.8 ;
         LAYER m3 ;
         RECT  0.0 230.4 207.6 231.6 ;
         LAYER m3 ;
         RECT  0.0 28.8 27.6 30.0 ;
         LAYER m4 ;
         RECT  141.6 2.4 142.8 423.6 ;
         LAYER m3 ;
         RECT  183.6 159.6 184.4 160.4 ;
         LAYER m3 ;
         RECT  167.5 342.4 168.3 343.2 ;
         LAYER m4 ;
         RECT  98.4 2.4 99.6 423.6 ;
         LAYER m3 ;
         RECT  23.2 263.2 24.0 264.0 ;
         LAYER m3 ;
         RECT  0.0 225.6 87.6 226.8 ;
         LAYER m3 ;
         RECT  0.0 19.2 207.6 20.4 ;
         LAYER m3 ;
         RECT  176.3 217.2 177.1 218.0 ;
         LAYER m3 ;
         RECT  197.2 159.6 198.0 160.4 ;
         LAYER m3 ;
         RECT  0.0 24.0 37.2 25.2 ;
         LAYER m3 ;
         RECT  111.7 22.4 112.5 23.2 ;
         LAYER m3 ;
         RECT  167.5 259.2 168.3 260.0 ;
         LAYER m3 ;
         RECT  129.6 201.6 169.2 202.8 ;
         LAYER m3 ;
         RECT  0.0 240.0 207.6 241.2 ;
         LAYER m4 ;
         RECT  79.2 2.4 80.4 423.6 ;
         LAYER m3 ;
         RECT  86.4 355.2 166.8 356.4 ;
         LAYER m4 ;
         RECT  55.2 2.4 56.4 423.6 ;
         LAYER m3 ;
         RECT  112.8 225.6 147.6 226.8 ;
         LAYER m3 ;
         RECT  176.3 258.8 177.1 259.6 ;
         LAYER m3 ;
         RECT  172.8 331.2 207.6 332.4 ;
         LAYER m3 ;
         RECT  190.1 91.4 190.9 92.2 ;
         LAYER m3 ;
         RECT  72.0 345.6 169.2 346.8 ;
         LAYER m3 ;
         RECT  177.6 355.2 205.2 356.4 ;
         LAYER m3 ;
         RECT  0.0 144.0 207.6 145.2 ;
         LAYER m3 ;
         RECT  0.0 350.4 147.6 351.6 ;
         LAYER m4 ;
         RECT  21.6 2.4 22.8 423.6 ;
         LAYER m3 ;
         RECT  0.0 86.4 188.4 87.6 ;
         LAYER m4 ;
         RECT  189.6 2.4 190.8 423.6 ;
         LAYER m3 ;
         RECT  0.0 211.2 116.4 212.4 ;
         LAYER m4 ;
         RECT  184.8 2.4 186.0 423.6 ;
         LAYER m4 ;
         RECT  175.2 2.4 176.4 423.6 ;
         LAYER m3 ;
         RECT  93.1 259.2 93.9 260.0 ;
         LAYER m3 ;
         RECT  203.5 175.6 204.3 176.4 ;
         LAYER m3 ;
         RECT  68.1 364.4 68.9 365.2 ;
         LAYER m4 ;
         RECT  74.4 2.4 75.6 423.6 ;
         LAYER m3 ;
         RECT  33.6 235.2 207.6 236.4 ;
         LAYER m4 ;
         RECT  16.8 2.4 18.0 423.6 ;
         LAYER m4 ;
         RECT  194.4 2.4 195.6 423.6 ;
         LAYER m3 ;
         RECT  33.6 254.4 116.4 255.6 ;
         LAYER m3 ;
         RECT  129.6 264.0 169.2 265.2 ;
         LAYER m3 ;
         RECT  129.6 273.6 169.2 274.8 ;
         LAYER m3 ;
         RECT  170.4 91.2 207.6 92.4 ;
         LAYER m3 ;
         RECT  0.0 110.4 207.6 111.6 ;
         LAYER m3 ;
         RECT  10.0 224.0 10.8 224.8 ;
         LAYER m3 ;
         RECT  129.6 220.8 169.2 222.0 ;
         LAYER m4 ;
         RECT  60.0 2.4 61.2 423.6 ;
         LAYER m4 ;
         RECT  112.8 2.4 114.0 423.6 ;
         LAYER m3 ;
         RECT  23.2 224.0 24.0 224.8 ;
         LAYER m3 ;
         RECT  26.4 206.4 87.6 207.6 ;
         LAYER m3 ;
         RECT  0.0 278.4 121.2 279.6 ;
         LAYER m3 ;
         RECT  0.0 48.0 207.6 49.2 ;
         LAYER m3 ;
         RECT  152.0 321.6 152.8 322.4 ;
         LAYER m3 ;
         RECT  189.9 175.6 190.7 176.4 ;
         LAYER m3 ;
         RECT  108.1 196.8 108.9 197.6 ;
         LAYER m3 ;
         RECT  176.3 279.6 177.1 280.4 ;
         LAYER m3 ;
         RECT  23.2 184.8 24.0 185.6 ;
         LAYER m3 ;
         RECT  0.0 9.6 207.6 10.8 ;
         LAYER m3 ;
         RECT  203.5 217.2 204.3 218.0 ;
         LAYER m3 ;
         RECT  152.0 300.8 152.8 301.6 ;
         LAYER m4 ;
         RECT  7.2 2.4 8.4 423.6 ;
         LAYER m3 ;
         RECT  152.0 259.2 152.8 260.0 ;
         LAYER m3 ;
         RECT  67.2 52.8 207.6 54.0 ;
         LAYER m3 ;
         RECT  203.5 321.2 204.3 322.0 ;
         LAYER m3 ;
         RECT  129.6 192.0 169.2 193.2 ;
         LAYER m3 ;
         RECT  167.5 238.4 168.3 239.2 ;
         LAYER m3 ;
         RECT  0.0 120.0 73.2 121.2 ;
         LAYER m3 ;
         RECT  176.3 362.8 177.1 363.6 ;
         LAYER m3 ;
         RECT  0.0 316.8 169.2 318.0 ;
         LAYER m4 ;
         RECT  40.8 2.4 42.0 423.6 ;
         LAYER m3 ;
         RECT  33.6 273.6 116.4 274.8 ;
         LAYER m3 ;
         RECT  177.6 168.0 205.2 169.2 ;
         LAYER m4 ;
         RECT  69.6 2.4 70.8 423.6 ;
         LAYER m3 ;
         RECT  196.7 175.6 197.5 176.4 ;
         LAYER m3 ;
         RECT  68.1 404.4 68.9 405.2 ;
         LAYER m3 ;
         RECT  91.2 393.6 207.6 394.8 ;
         LAYER m3 ;
         RECT  0.0 216.0 121.2 217.2 ;
         LAYER m4 ;
         RECT  103.2 2.4 104.4 423.6 ;
         LAYER m3 ;
         RECT  203.5 300.4 204.3 301.2 ;
         LAYER m3 ;
         RECT  0.0 259.2 121.2 260.4 ;
         LAYER m3 ;
         RECT  152.0 280.0 152.8 280.8 ;
         LAYER m3 ;
         RECT  93.1 280.0 93.9 280.8 ;
         LAYER m3 ;
         RECT  176.3 196.4 177.1 197.2 ;
         LAYER m3 ;
         RECT  0.0 72.0 75.6 73.2 ;
         LAYER m3 ;
         RECT  108.1 259.2 108.9 260.0 ;
         LAYER m3 ;
         RECT  77.6 142.4 78.4 143.2 ;
         LAYER m3 ;
         RECT  175.2 72.0 207.6 73.2 ;
         LAYER m3 ;
         RECT  23.2 341.6 24.0 342.4 ;
         LAYER m3 ;
         RECT  93.1 217.6 93.9 218.4 ;
         LAYER m4 ;
         RECT  64.8 2.4 66.0 423.6 ;
         LAYER m4 ;
         RECT  136.8 2.4 138.0 423.6 ;
         LAYER m4 ;
         RECT  132.0 2.4 133.2 423.6 ;
         LAYER m3 ;
         RECT  129.6 283.2 169.2 284.4 ;
         LAYER m3 ;
         RECT  172.8 249.6 207.6 250.8 ;
         LAYER m3 ;
         RECT  172.8 350.4 207.6 351.6 ;
         LAYER m3 ;
         RECT  196.9 91.4 197.7 92.2 ;
         LAYER m3 ;
         RECT  167.5 217.6 168.3 218.4 ;
         LAYER m3 ;
         RECT  77.6 102.4 78.4 103.2 ;
         LAYER m3 ;
         RECT  152.0 238.4 152.8 239.2 ;
         LAYER m3 ;
         RECT  0.0 38.4 207.6 39.6 ;
         LAYER m3 ;
         RECT  0.0 187.2 87.6 188.4 ;
         LAYER m3 ;
         RECT  172.8 187.2 207.6 188.4 ;
         LAYER m3 ;
         RECT  196.7 362.8 197.5 363.6 ;
         LAYER m3 ;
         RECT  0.0 369.6 207.6 370.8 ;
         LAYER m3 ;
         RECT  112.8 288.0 147.6 289.2 ;
         LAYER m3 ;
         RECT  0.0 192.0 116.4 193.2 ;
         LAYER m3 ;
         RECT  172.8 268.8 207.6 270.0 ;
         LAYER m3 ;
         RECT  0.0 345.6 63.6 346.8 ;
         LAYER m3 ;
         RECT  0.0 422.4 63.6 423.6 ;
         LAYER m3 ;
         RECT  0.0 336.0 169.2 337.2 ;
         LAYER m4 ;
         RECT  204.0 2.4 205.2 423.6 ;
         LAYER m3 ;
         RECT  167.5 300.8 168.3 301.6 ;
         LAYER m3 ;
         RECT  183.1 362.8 183.9 363.6 ;
         LAYER m3 ;
         RECT  108.1 217.6 108.9 218.4 ;
         LAYER m3 ;
         RECT  10.0 302.4 10.8 303.2 ;
         LAYER m3 ;
         RECT  81.6 81.6 186.0 82.8 ;
         LAYER m3 ;
         RECT  0.0 57.6 207.6 58.8 ;
         LAYER m3 ;
         RECT  33.6 331.2 147.6 332.4 ;
         LAYER m3 ;
         RECT  77.6 22.4 78.4 23.2 ;
         LAYER m3 ;
         RECT  0.0 326.4 169.2 327.6 ;
         LAYER m3 ;
         RECT  0.0 360.0 207.6 361.2 ;
         LAYER m3 ;
         RECT  4.8 43.2 73.2 44.4 ;
         LAYER m3 ;
         RECT  132.0 196.8 207.6 198.0 ;
         LAYER m3 ;
         RECT  0.0 403.2 207.6 404.4 ;
         LAYER m3 ;
         RECT  203.5 258.8 204.3 259.6 ;
         LAYER m4 ;
         RECT  199.2 2.4 200.4 423.6 ;
         LAYER m3 ;
         RECT  26.4 321.6 207.6 322.8 ;
         LAYER m3 ;
         RECT  0.0 196.8 121.2 198.0 ;
         LAYER m4 ;
         RECT  180.0 2.4 181.2 423.6 ;
         LAYER m3 ;
         RECT  183.1 175.6 183.9 176.4 ;
         LAYER m3 ;
         RECT  176.3 321.2 177.1 322.0 ;
         LAYER m3 ;
         RECT  190.4 159.6 191.2 160.4 ;
         LAYER m3 ;
         RECT  0.0 33.6 207.6 34.8 ;
         LAYER m3 ;
         RECT  0.0 96.0 207.6 97.2 ;
         LAYER m3 ;
         RECT  172.8 288.0 207.6 289.2 ;
         LAYER m3 ;
         RECT  0.0 302.4 207.6 303.6 ;
         LAYER m3 ;
         RECT  81.6 43.2 207.6 44.4 ;
         LAYER m3 ;
         RECT  2.0 22.4 2.8 23.2 ;
         LAYER m3 ;
         RECT  141.6 278.4 207.6 279.6 ;
         LAYER m3 ;
         RECT  152.0 196.8 152.8 197.6 ;
         LAYER m3 ;
         RECT  192.3 125.4 193.1 126.2 ;
         LAYER m3 ;
         RECT  203.5 362.8 204.3 363.6 ;
         LAYER m3 ;
         RECT  176.3 300.4 177.1 301.2 ;
         LAYER m4 ;
         RECT  31.2 2.4 32.4 423.6 ;
         LAYER m3 ;
         RECT  108.1 280.0 108.9 280.8 ;
         LAYER m3 ;
         RECT  176.3 342.0 177.1 342.8 ;
         LAYER m3 ;
         RECT  33.6 312.0 147.6 313.2 ;
         LAYER m3 ;
         RECT  148.8 4.8 207.6 6.0 ;
         LAYER m3 ;
         RECT  10.0 341.6 10.8 342.4 ;
         LAYER m3 ;
         RECT  0.0 182.4 169.2 183.6 ;
         LAYER m3 ;
         RECT  203.5 196.4 204.3 197.2 ;
         LAYER m3 ;
         RECT  0.0 374.4 70.8 375.6 ;
         LAYER m3 ;
         RECT  0.0 220.8 121.2 222.0 ;
         LAYER m3 ;
         RECT  170.4 153.6 207.6 154.8 ;
         LAYER m3 ;
         RECT  0.0 129.6 207.6 130.8 ;
         LAYER m3 ;
         RECT  199.1 125.4 199.9 126.2 ;
         LAYER m3 ;
         RECT  0.0 398.4 207.6 399.6 ;
         LAYER m4 ;
         RECT  88.8 2.4 90.0 423.6 ;
         LAYER m4 ;
         RECT  146.4 2.4 147.6 423.6 ;
         LAYER m3 ;
         RECT  0.0 14.4 27.6 15.6 ;
         LAYER m3 ;
         RECT  93.1 196.8 93.9 197.6 ;
         LAYER m3 ;
         RECT  0.0 91.2 75.6 92.4 ;
         LAYER m3 ;
         RECT  60.0 124.8 207.6 126.0 ;
         LAYER m3 ;
         RECT  26.4 283.2 121.2 284.4 ;
         LAYER m3 ;
         RECT  0.0 393.6 70.8 394.8 ;
         LAYER m3 ;
         RECT  0.0 168.0 166.8 169.2 ;
         LAYER m3 ;
         RECT  0.0 76.8 207.6 78.0 ;
         LAYER m3 ;
         RECT  33.6 292.8 207.6 294.0 ;
         LAYER m4 ;
         RECT  156.0 2.4 157.2 423.6 ;
         LAYER m3 ;
         RECT  0.0 379.2 207.6 380.4 ;
         LAYER m4 ;
         RECT  50.4 2.4 51.6 423.6 ;
         LAYER m4 ;
         RECT  93.6 2.4 94.8 423.6 ;
         LAYER m3 ;
         RECT  0.0 134.4 207.6 135.6 ;
         LAYER m3 ;
         RECT  0.0 139.2 188.4 140.4 ;
         LAYER m3 ;
         RECT  134.4 216.0 207.6 217.2 ;
         LAYER m4 ;
         RECT  108.0 2.4 109.2 423.6 ;
         LAYER m3 ;
         RECT  26.4 163.2 73.2 164.4 ;
         LAYER m4 ;
         RECT  160.8 2.4 162.0 423.6 ;
         LAYER m3 ;
         RECT  0.0 4.8 44.4 6.0 ;
         LAYER m3 ;
         RECT  0.0 81.6 73.2 82.8 ;
         LAYER m4 ;
         RECT  36.0 2.4 37.2 423.6 ;
         LAYER m3 ;
         RECT  203.5 342.0 204.3 342.8 ;
         LAYER m4 ;
         RECT  84.0 2.4 85.2 423.6 ;
         LAYER m4 ;
         RECT  45.6 2.4 46.8 423.6 ;
         LAYER m3 ;
         RECT  0.0 307.2 169.2 308.4 ;
         LAYER m3 ;
         RECT  77.6 62.4 78.4 63.2 ;
         LAYER m3 ;
         RECT  167.5 321.6 168.3 322.4 ;
         LAYER m3 ;
         RECT  10.0 263.2 10.8 264.0 ;
         LAYER m3 ;
         RECT  69.6 384.0 207.6 385.2 ;
         LAYER m3 ;
         RECT  176.3 238.0 177.1 238.8 ;
         LAYER m3 ;
         RECT  10.0 184.8 10.8 185.6 ;
         LAYER m3 ;
         RECT  203.5 279.6 204.3 280.4 ;
         LAYER m3 ;
         RECT  0.0 52.8 39.6 54.0 ;
         LAYER m4 ;
         RECT  122.4 2.4 123.6 423.6 ;
         LAYER m3 ;
         RECT  0.0 62.4 207.6 63.6 ;
         LAYER m3 ;
         RECT  0.0 177.6 207.6 178.8 ;
         LAYER m3 ;
         RECT  0.0 340.8 207.6 342.0 ;
         LAYER m4 ;
         RECT  165.6 2.4 166.8 423.6 ;
         LAYER m3 ;
         RECT  0.0 264.0 116.4 265.2 ;
         LAYER m4 ;
         RECT  170.4 2.4 171.6 423.6 ;
         LAYER m3 ;
         RECT  197.5 74.0 198.3 74.8 ;
         LAYER m3 ;
         RECT  91.2 412.8 207.6 414.0 ;
         LAYER m3 ;
         RECT  0.0 412.8 70.8 414.0 ;
         LAYER m4 ;
         RECT  151.2 2.4 152.4 423.6 ;
         LAYER m3 ;
         RECT  0.0 148.8 27.6 150.0 ;
         LAYER m3 ;
         RECT  0.0 268.8 87.6 270.0 ;
         LAYER m3 ;
         RECT  74.4 24.0 207.6 25.2 ;
         LAYER m3 ;
         RECT  0.0 158.4 207.6 159.6 ;
         LAYER m3 ;
         RECT  52.8 14.4 207.6 15.6 ;
         LAYER m3 ;
         RECT  129.6 211.2 169.2 212.4 ;
         LAYER m3 ;
         RECT  136.8 259.2 207.6 260.4 ;
         LAYER m3 ;
         RECT  0.0 384.0 63.6 385.2 ;
         LAYER m3 ;
         RECT  26.4 244.8 169.2 246.0 ;
         LAYER m4 ;
         RECT  26.4 2.4 27.6 423.6 ;
         LAYER m4 ;
         RECT  127.2 2.4 128.4 423.6 ;
         LAYER m3 ;
         RECT  203.5 238.0 204.3 238.8 ;
         LAYER m4 ;
         RECT  2.4 2.4 3.6 423.6 ;
         LAYER m3 ;
         RECT  152.0 217.6 152.8 218.4 ;
         LAYER m3 ;
         RECT  172.8 225.6 207.6 226.8 ;
         LAYER m3 ;
         RECT  0.0 100.8 183.6 102.0 ;
         LAYER m3 ;
         RECT  0.0 201.6 116.4 202.8 ;
         LAYER m3 ;
         RECT  0.0 297.6 207.6 298.8 ;
         LAYER m3 ;
         RECT  0.0 355.2 70.8 356.4 ;
         LAYER m3 ;
         RECT  167.5 196.8 168.3 197.6 ;
         LAYER m3 ;
         RECT  88.8 374.4 207.6 375.6 ;
         LAYER m3 ;
         RECT  0.0 288.0 87.6 289.2 ;
         LAYER m4 ;
         RECT  117.6 2.4 118.8 423.6 ;
         LAYER m3 ;
         RECT  176.3 175.6 177.1 176.4 ;
         LAYER m3 ;
         RECT  0.0 408.0 207.6 409.2 ;
         LAYER m4 ;
         RECT  12.0 2.4 13.2 423.6 ;
         LAYER m3 ;
         RECT  172.8 206.4 207.6 207.6 ;
         LAYER m3 ;
         RECT  133.5 22.4 134.3 23.2 ;
         LAYER m3 ;
         RECT  152.0 342.4 152.8 343.2 ;
         LAYER m3 ;
         RECT  129.6 254.4 169.2 255.6 ;
         LAYER m3 ;
         RECT  190.7 74.0 191.5 74.8 ;
         LAYER m3 ;
         RECT  48.0 28.8 207.6 30.0 ;
         LAYER m3 ;
         RECT  0.0 115.2 207.6 116.4 ;
         LAYER m3 ;
         RECT  0.0 388.8 207.6 390.0 ;
         LAYER m3 ;
         RECT  0.0 124.8 34.8 126.0 ;
         LAYER m3 ;
         RECT  0.0 249.6 87.6 250.8 ;
         LAYER m3 ;
         RECT  167.5 280.0 168.3 280.8 ;
         LAYER m3 ;
         RECT  189.9 362.8 190.7 363.6 ;
         LAYER m3 ;
         RECT  172.8 312.0 207.6 313.2 ;
         LAYER m3 ;
         RECT  33.6 172.8 207.6 174.0 ;
         LAYER m3 ;
         RECT  23.2 302.4 24.0 303.2 ;
         LAYER m3 ;
         RECT  0.0 105.6 207.6 106.8 ;
         LAYER m3 ;
         RECT  0.0 364.8 207.6 366.0 ;
         LAYER m3 ;
         RECT  81.6 120.0 207.6 121.2 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER m3 ;
         RECT  179.7 347.0 180.5 347.8 ;
         LAYER m3 ;
         RECT  0.0 74.4 75.6 75.6 ;
         LAYER m3 ;
         RECT  172.9 337.0 173.7 337.8 ;
         LAYER m3 ;
         RECT  200.1 295.4 200.9 296.2 ;
         LAYER m4 ;
         RECT  96.0 2.4 97.2 423.6 ;
         LAYER m3 ;
         RECT  179.7 284.6 180.5 285.4 ;
         LAYER m3 ;
         RECT  0.0 266.4 207.6 267.6 ;
         LAYER m3 ;
         RECT  186.5 170.6 187.3 171.4 ;
         LAYER m3 ;
         RECT  72.0 362.4 171.6 363.6 ;
         LAYER m3 ;
         RECT  172.9 191.4 173.7 192.2 ;
         LAYER m3 ;
         RECT  172.8 112.8 207.6 114.0 ;
         LAYER m4 ;
         RECT  182.4 2.4 183.6 423.6 ;
         LAYER m3 ;
         RECT  179.7 191.4 180.5 192.2 ;
         LAYER m3 ;
         RECT  179.7 212.2 180.5 213.0 ;
         LAYER m3 ;
         RECT  0.0 204.0 207.6 205.2 ;
         LAYER m3 ;
         RECT  172.9 274.6 173.7 275.4 ;
         LAYER m3 ;
         RECT  172.9 170.6 173.7 171.4 ;
         LAYER m3 ;
         RECT  77.6 122.4 78.4 123.2 ;
         LAYER m4 ;
         RECT  196.8 2.4 198.0 423.6 ;
         LAYER m3 ;
         RECT  0.0 218.4 87.6 219.6 ;
         LAYER m3 ;
         RECT  0.0 391.2 207.6 392.4 ;
         LAYER m4 ;
         RECT  192.0 2.4 193.2 423.6 ;
         LAYER m3 ;
         RECT  167.5 207.2 168.3 208.0 ;
         LAYER m3 ;
         RECT  129.6 276.0 207.6 277.2 ;
         LAYER m4 ;
         RECT  9.6 2.4 10.8 423.6 ;
         LAYER m3 ;
         RECT  206.9 201.4 207.7 202.2 ;
         LAYER m3 ;
         RECT  0.0 228.0 207.6 229.2 ;
         LAYER m3 ;
         RECT  0.0 93.6 207.6 94.8 ;
         LAYER m3 ;
         RECT  0.0 127.2 188.4 128.4 ;
         LAYER m4 ;
         RECT  124.8 2.4 126.0 423.6 ;
         LAYER m3 ;
         RECT  179.7 274.6 180.5 275.4 ;
         LAYER m3 ;
         RECT  0.0 7.2 75.6 8.4 ;
         LAYER m3 ;
         RECT  2.0 42.4 2.8 43.2 ;
         LAYER m3 ;
         RECT  200.1 316.2 200.9 317.0 ;
         LAYER m3 ;
         RECT  0.0 112.8 75.6 114.0 ;
         LAYER m3 ;
         RECT  23.2 204.4 24.0 205.2 ;
         LAYER m3 ;
         RECT  206.9 316.2 207.7 317.0 ;
         LAYER m3 ;
         RECT  33.6 232.8 207.6 234.0 ;
         LAYER m3 ;
         RECT  206.9 191.4 207.7 192.2 ;
         LAYER m3 ;
         RECT  172.9 180.6 173.7 181.4 ;
         LAYER m3 ;
         RECT  172.9 316.2 173.7 317.0 ;
         LAYER m3 ;
         RECT  0.0 26.4 37.2 27.6 ;
         LAYER m3 ;
         RECT  0.0 348.0 54.0 349.2 ;
         LAYER m3 ;
         RECT  0.0 40.8 207.6 42.0 ;
         LAYER m3 ;
         RECT  0.0 242.4 207.6 243.6 ;
         LAYER m3 ;
         RECT  0.0 386.4 207.6 387.6 ;
         LAYER m4 ;
         RECT  144.0 2.4 145.2 423.6 ;
         LAYER m3 ;
         RECT  206.9 357.8 207.7 358.6 ;
         LAYER m4 ;
         RECT  28.8 2.4 30.0 423.6 ;
         LAYER m3 ;
         RECT  68.1 344.4 68.9 345.2 ;
         LAYER m3 ;
         RECT  179.7 337.0 180.5 337.8 ;
         LAYER m3 ;
         RECT  152.0 207.2 152.8 208.0 ;
         LAYER m3 ;
         RECT  0.0 108.0 207.6 109.2 ;
         LAYER m3 ;
         RECT  0.0 367.2 207.6 368.4 ;
         LAYER m3 ;
         RECT  60.0 122.4 207.6 123.6 ;
         LAYER m3 ;
         RECT  132.0 184.8 207.6 186.0 ;
         LAYER m3 ;
         RECT  111.7 2.4 112.5 3.2 ;
         LAYER m4 ;
         RECT  148.8 2.4 150.0 423.6 ;
         LAYER m3 ;
         RECT  129.6 252.0 207.6 253.2 ;
         LAYER m3 ;
         RECT  0.0 165.6 207.6 166.8 ;
         LAYER m3 ;
         RECT  0.0 362.4 63.6 363.6 ;
         LAYER m3 ;
         RECT  167.5 332.0 168.3 332.8 ;
         LAYER m3 ;
         RECT  0.0 79.2 207.6 80.4 ;
         LAYER m4 ;
         RECT  76.8 2.4 78.0 423.6 ;
         LAYER m3 ;
         RECT  0.0 84.0 207.6 85.2 ;
         LAYER m3 ;
         RECT  179.7 253.8 180.5 254.6 ;
         LAYER m3 ;
         RECT  129.6 261.6 207.6 262.8 ;
         LAYER m3 ;
         RECT  0.0 160.8 178.8 162.0 ;
         LAYER m4 ;
         RECT  163.2 2.4 164.4 423.6 ;
         LAYER m3 ;
         RECT  209.0 167.8 209.8 168.6 ;
         LAYER m3 ;
         RECT  172.9 357.8 173.7 358.6 ;
         LAYER m3 ;
         RECT  0.0 319.2 147.6 320.4 ;
         LAYER m4 ;
         RECT  105.6 2.4 106.8 423.6 ;
         LAYER m3 ;
         RECT  206.9 284.6 207.7 285.4 ;
         LAYER m3 ;
         RECT  148.8 7.2 207.6 8.4 ;
         LAYER m3 ;
         RECT  93.1 207.2 93.9 208.0 ;
         LAYER m3 ;
         RECT  81.6 103.2 207.6 104.4 ;
         LAYER m3 ;
         RECT  93.1 186.4 93.9 187.2 ;
         LAYER m3 ;
         RECT  167.5 186.4 168.3 187.2 ;
         LAYER m3 ;
         RECT  206.9 295.4 207.7 296.2 ;
         LAYER m3 ;
         RECT  26.4 343.2 147.6 344.4 ;
         LAYER m3 ;
         RECT  200.1 357.8 200.9 358.6 ;
         LAYER m3 ;
         RECT  112.8 256.8 147.6 258.0 ;
         LAYER m3 ;
         RECT  179.7 233.0 180.5 233.8 ;
         LAYER m3 ;
         RECT  0.0 98.4 207.6 99.6 ;
         LAYER m3 ;
         RECT  206.9 233.0 207.7 233.8 ;
         LAYER m3 ;
         RECT  172.9 263.8 173.7 264.6 ;
         LAYER m3 ;
         RECT  206.9 347.0 207.7 347.8 ;
         LAYER m3 ;
         RECT  200.1 253.8 200.9 254.6 ;
         LAYER m3 ;
         RECT  93.1 228.0 93.9 228.8 ;
         LAYER m3 ;
         RECT  0.0 64.8 207.6 66.0 ;
         LAYER m3 ;
         RECT  0.0 88.8 207.6 90.0 ;
         LAYER m3 ;
         RECT  112.8 194.4 147.6 195.6 ;
         LAYER m3 ;
         RECT  179.7 170.6 180.5 171.4 ;
         LAYER m3 ;
         RECT  0.0 50.4 39.6 51.6 ;
         LAYER m3 ;
         RECT  152.0 186.4 152.8 187.2 ;
         LAYER m3 ;
         RECT  172.9 295.4 173.7 296.2 ;
         LAYER m3 ;
         RECT  108.1 207.2 108.9 208.0 ;
         LAYER m3 ;
         RECT  129.6 223.2 207.6 224.4 ;
         LAYER m3 ;
         RECT  108.1 269.6 108.9 270.4 ;
         LAYER m3 ;
         RECT  172.9 243.0 173.7 243.8 ;
         LAYER m3 ;
         RECT  33.6 194.4 87.6 195.6 ;
         LAYER m3 ;
         RECT  23.2 243.6 24.0 244.4 ;
         LAYER m3 ;
         RECT  200.1 138.8 200.9 139.6 ;
         LAYER m3 ;
         RECT  0.0 189.6 116.4 190.8 ;
         LAYER m4 ;
         RECT  67.2 2.4 68.4 423.6 ;
         LAYER m3 ;
         RECT  152.0 352.8 152.8 353.6 ;
         LAYER m3 ;
         RECT  0.0 280.8 87.6 282.0 ;
         LAYER m3 ;
         RECT  0.0 36.0 34.8 37.2 ;
         LAYER m3 ;
         RECT  26.4 300.0 147.6 301.2 ;
         LAYER m3 ;
         RECT  0.0 276.0 116.4 277.2 ;
         LAYER m4 ;
         RECT  33.6 2.4 34.8 423.6 ;
         LAYER m3 ;
         RECT  0.0 180.0 207.6 181.2 ;
         LAYER m3 ;
         RECT  0.0 16.8 207.6 18.0 ;
         LAYER m3 ;
         RECT  0.0 357.6 207.6 358.8 ;
         LAYER m3 ;
         RECT  0.0 122.4 34.8 123.6 ;
         LAYER m3 ;
         RECT  0.0 55.2 207.6 56.4 ;
         LAYER m3 ;
         RECT  0.0 117.6 207.6 118.8 ;
         LAYER m3 ;
         RECT  0.0 314.4 207.6 315.6 ;
         LAYER m3 ;
         RECT  139.2 21.6 207.6 22.8 ;
         LAYER m3 ;
         RECT  33.6 290.4 207.6 291.6 ;
         LAYER m3 ;
         RECT  68.1 424.4 68.9 425.2 ;
         LAYER m3 ;
         RECT  179.7 305.4 180.5 306.2 ;
         LAYER m3 ;
         RECT  68.1 384.4 68.9 385.2 ;
         LAYER m3 ;
         RECT  179.7 180.6 180.5 181.4 ;
         LAYER m3 ;
         RECT  2.0 2.4 2.8 3.2 ;
         LAYER m3 ;
         RECT  23.2 322.0 24.0 322.8 ;
         LAYER m3 ;
         RECT  0.0 208.8 121.2 210.0 ;
         LAYER m3 ;
         RECT  152.0 228.0 152.8 228.8 ;
         LAYER m3 ;
         RECT  200.1 263.8 200.9 264.6 ;
         LAYER m3 ;
         RECT  0.0 376.8 207.6 378.0 ;
         LAYER m3 ;
         RECT  0.0 304.8 207.6 306.0 ;
         LAYER m3 ;
         RECT  206.9 212.2 207.7 213.0 ;
         LAYER m3 ;
         RECT  133.5 2.4 134.3 3.2 ;
         LAYER m4 ;
         RECT  129.6 2.4 130.8 423.6 ;
         LAYER m4 ;
         RECT  134.4 2.4 135.6 423.6 ;
         LAYER m3 ;
         RECT  0.0 136.8 207.6 138.0 ;
         LAYER m3 ;
         RECT  26.4 223.2 116.4 224.4 ;
         LAYER m3 ;
         RECT  206.9 170.6 207.7 171.4 ;
         LAYER m3 ;
         RECT  26.4 184.8 121.2 186.0 ;
         LAYER m3 ;
         RECT  179.7 263.8 180.5 264.6 ;
         LAYER m3 ;
         RECT  172.9 326.2 173.7 327.0 ;
         LAYER m4 ;
         RECT  0.0 2.4 1.2 423.6 ;
         LAYER m3 ;
         RECT  0.0 60.0 73.2 61.2 ;
         LAYER m3 ;
         RECT  33.6 271.2 121.2 272.4 ;
         LAYER m3 ;
         RECT  152.0 332.0 152.8 332.8 ;
         LAYER m3 ;
         RECT  0.0 405.6 63.6 406.8 ;
         LAYER m3 ;
         RECT  167.5 311.2 168.3 312.0 ;
         LAYER m4 ;
         RECT  168.0 2.4 169.2 423.6 ;
         LAYER m3 ;
         RECT  0.0 2.4 44.4 3.6 ;
         LAYER m4 ;
         RECT  62.4 2.4 63.6 423.6 ;
         LAYER m3 ;
         RECT  72.0 405.6 207.6 406.8 ;
         LAYER m3 ;
         RECT  179.7 316.2 180.5 317.0 ;
         LAYER m3 ;
         RECT  167.5 228.0 168.3 228.8 ;
         LAYER m3 ;
         RECT  206.9 243.0 207.7 243.8 ;
         LAYER m3 ;
         RECT  172.9 212.2 173.7 213.0 ;
         LAYER m3 ;
         RECT  179.7 357.8 180.5 358.6 ;
         LAYER m3 ;
         RECT  0.0 328.8 207.6 330.0 ;
         LAYER m3 ;
         RECT  200.1 201.4 200.9 202.2 ;
         LAYER m3 ;
         RECT  0.0 352.8 70.8 354.0 ;
         LAYER m3 ;
         RECT  0.0 396.0 207.6 397.2 ;
         LAYER m3 ;
         RECT  134.4 208.8 207.6 210.0 ;
         LAYER m3 ;
         RECT  0.0 415.2 70.8 416.4 ;
         LAYER m3 ;
         RECT  152.0 269.6 152.8 270.4 ;
         LAYER m3 ;
         RECT  0.0 237.6 147.6 238.8 ;
         LAYER m3 ;
         RECT  4.8 21.6 73.2 22.8 ;
         LAYER m3 ;
         RECT  86.4 348.0 207.6 349.2 ;
         LAYER m3 ;
         RECT  93.1 290.4 93.9 291.2 ;
         LAYER m3 ;
         RECT  67.2 36.0 207.6 37.2 ;
         LAYER m3 ;
         RECT  200.1 170.6 200.9 171.4 ;
         LAYER m3 ;
         RECT  167.5 269.6 168.3 270.4 ;
         LAYER m3 ;
         RECT  170.4 151.2 207.6 152.4 ;
         LAYER m3 ;
         RECT  200.1 274.6 200.9 275.4 ;
         LAYER m3 ;
         RECT  86.4 352.8 207.6 354.0 ;
         LAYER m3 ;
         RECT  81.6 60.0 207.6 61.2 ;
         LAYER m3 ;
         RECT  172.9 305.4 173.7 306.2 ;
         LAYER m3 ;
         RECT  0.0 69.6 207.6 70.8 ;
         LAYER m3 ;
         RECT  200.1 243.0 200.9 243.8 ;
         LAYER m3 ;
         RECT  152.0 290.4 152.8 291.2 ;
         LAYER m3 ;
         RECT  129.6 189.6 207.6 190.8 ;
         LAYER m4 ;
         RECT  158.4 2.4 159.6 423.6 ;
         LAYER m3 ;
         RECT  172.9 253.8 173.7 254.6 ;
         LAYER m3 ;
         RECT  192.1 85.0 192.9 85.8 ;
         LAYER m3 ;
         RECT  0.0 156.0 207.6 157.2 ;
         LAYER m3 ;
         RECT  179.7 222.2 180.5 223.0 ;
         LAYER m3 ;
         RECT  206.9 326.2 207.7 327.0 ;
         LAYER m4 ;
         RECT  38.4 2.4 39.6 423.6 ;
         LAYER m3 ;
         RECT  0.0 132.0 207.6 133.2 ;
         LAYER m3 ;
         RECT  77.6 2.4 78.4 3.2 ;
         LAYER m4 ;
         RECT  4.8 2.4 6.0 423.6 ;
         LAYER m3 ;
         RECT  167.5 290.4 168.3 291.2 ;
         LAYER m3 ;
         RECT  33.6 175.2 171.6 176.4 ;
         LAYER m3 ;
         RECT  206.9 253.8 207.7 254.6 ;
         LAYER m3 ;
         RECT  10.0 165.2 10.8 166.0 ;
         LAYER m3 ;
         RECT  179.7 201.4 180.5 202.2 ;
         LAYER m3 ;
         RECT  200.1 180.6 200.9 181.4 ;
         LAYER m4 ;
         RECT  57.6 2.4 58.8 423.6 ;
         LAYER m4 ;
         RECT  72.0 2.4 73.2 423.6 ;
         LAYER m4 ;
         RECT  201.6 2.4 202.8 423.6 ;
         LAYER m3 ;
         RECT  0.0 400.8 207.6 402.0 ;
         LAYER m3 ;
         RECT  172.9 201.4 173.7 202.2 ;
         LAYER m3 ;
         RECT  0.0 420.0 207.6 421.2 ;
         LAYER m3 ;
         RECT  172.9 284.6 173.7 285.4 ;
         LAYER m3 ;
         RECT  10.0 243.6 10.8 244.4 ;
         LAYER m3 ;
         RECT  0.0 256.8 87.6 258.0 ;
         LAYER m3 ;
         RECT  0.0 151.2 75.6 152.4 ;
         LAYER m3 ;
         RECT  200.1 212.2 200.9 213.0 ;
         LAYER m4 ;
         RECT  19.2 2.4 20.4 423.6 ;
         LAYER m3 ;
         RECT  200.1 284.6 200.9 285.4 ;
         LAYER m3 ;
         RECT  0.0 285.6 116.4 286.8 ;
         LAYER m3 ;
         RECT  172.9 222.2 173.7 223.0 ;
         LAYER m3 ;
         RECT  108.1 248.8 108.9 249.6 ;
         LAYER m3 ;
         RECT  206.9 180.6 207.7 181.4 ;
         LAYER m4 ;
         RECT  153.6 2.4 154.8 423.6 ;
         LAYER m3 ;
         RECT  197.5 80.6 198.3 81.4 ;
         LAYER m3 ;
         RECT  10.0 322.0 10.8 322.8 ;
         LAYER m3 ;
         RECT  76.8 2.4 207.6 3.6 ;
         LAYER m3 ;
         RECT  0.0 410.4 207.6 411.6 ;
         LAYER m3 ;
         RECT  200.1 337.0 200.9 337.8 ;
         LAYER m3 ;
         RECT  139.2 271.2 207.6 272.4 ;
         LAYER m3 ;
         RECT  77.6 82.4 78.4 83.2 ;
         LAYER m3 ;
         RECT  172.9 233.0 173.7 233.8 ;
         LAYER m3 ;
         RECT  167.5 352.8 168.3 353.6 ;
         LAYER m3 ;
         RECT  200.1 233.0 200.9 233.8 ;
         LAYER m3 ;
         RECT  200.1 191.4 200.9 192.2 ;
         LAYER m4 ;
         RECT  81.6 2.4 82.8 423.6 ;
         LAYER m3 ;
         RECT  190.7 80.6 191.5 81.4 ;
         LAYER m3 ;
         RECT  170.8 355.0 171.6 355.8 ;
         LAYER m3 ;
         RECT  0.0 324.0 207.6 325.2 ;
         LAYER m3 ;
         RECT  200.1 222.2 200.9 223.0 ;
         LAYER m3 ;
         RECT  77.6 162.4 78.4 163.2 ;
         LAYER m3 ;
         RECT  129.6 199.2 207.6 200.4 ;
         LAYER m4 ;
         RECT  91.2 2.4 92.4 423.6 ;
         LAYER m4 ;
         RECT  139.2 2.4 140.4 423.6 ;
         LAYER m3 ;
         RECT  193.3 170.6 194.1 171.4 ;
         LAYER m3 ;
         RECT  196.1 99.6 196.9 100.4 ;
         LAYER m4 ;
         RECT  120.0 2.4 121.2 423.6 ;
         LAYER m3 ;
         RECT  206.9 263.8 207.7 264.6 ;
         LAYER m3 ;
         RECT  0.0 170.4 207.6 171.6 ;
         LAYER m3 ;
         RECT  193.3 357.8 194.1 358.6 ;
         LAYER m3 ;
         RECT  152.0 248.8 152.8 249.6 ;
         LAYER m3 ;
         RECT  0.0 247.2 121.2 248.4 ;
         LAYER m3 ;
         RECT  179.7 243.0 180.5 243.8 ;
         LAYER m3 ;
         RECT  206.9 337.0 207.7 337.8 ;
         LAYER m3 ;
         RECT  93.1 269.6 93.9 270.4 ;
         LAYER m4 ;
         RECT  206.4 2.4 207.6 423.6 ;
         LAYER m3 ;
         RECT  108.1 290.4 108.9 291.2 ;
         LAYER m3 ;
         RECT  0.0 199.2 121.2 200.4 ;
         LAYER m3 ;
         RECT  129.6 285.6 207.6 286.8 ;
         LAYER m4 ;
         RECT  177.6 2.4 178.8 423.6 ;
         LAYER m3 ;
         RECT  209.0 355.0 209.8 355.8 ;
         LAYER m3 ;
         RECT  193.3 138.8 194.1 139.6 ;
         LAYER m4 ;
         RECT  48.0 2.4 49.2 423.6 ;
         LAYER m3 ;
         RECT  108.1 186.4 108.9 187.2 ;
         LAYER m3 ;
         RECT  206.9 274.6 207.7 275.4 ;
         LAYER m3 ;
         RECT  0.0 146.4 27.6 147.6 ;
         LAYER m3 ;
         RECT  0.0 372.0 207.6 373.2 ;
         LAYER m3 ;
         RECT  198.9 85.0 199.7 85.8 ;
         LAYER m3 ;
         RECT  136.8 247.2 207.6 248.4 ;
         LAYER m4 ;
         RECT  14.4 2.4 15.6 423.6 ;
         LAYER m3 ;
         RECT  74.4 26.4 207.6 27.6 ;
         LAYER m3 ;
         RECT  33.6 213.6 116.4 214.8 ;
         LAYER m3 ;
         RECT  206.9 222.2 207.7 223.0 ;
         LAYER m3 ;
         RECT  81.6 141.6 207.6 142.8 ;
         LAYER m3 ;
         RECT  91.2 415.2 207.6 416.4 ;
         LAYER m4 ;
         RECT  110.4 2.4 111.6 423.6 ;
         LAYER m3 ;
         RECT  0.0 141.6 73.2 142.8 ;
         LAYER m3 ;
         RECT  200.1 326.2 200.9 327.0 ;
         LAYER m3 ;
         RECT  0.0 31.2 27.6 32.4 ;
         LAYER m4 ;
         RECT  100.8 2.4 102.0 423.6 ;
         LAYER m3 ;
         RECT  152.0 311.2 152.8 312.0 ;
         LAYER m3 ;
         RECT  33.6 252.0 116.4 253.2 ;
         LAYER m3 ;
         RECT  108.1 228.0 108.9 228.8 ;
         LAYER m3 ;
         RECT  172.9 347.0 173.7 347.8 ;
         LAYER m3 ;
         RECT  129.6 213.6 207.6 214.8 ;
         LAYER m3 ;
         RECT  200.1 305.4 200.9 306.2 ;
         LAYER m3 ;
         RECT  186.5 357.8 187.3 358.6 ;
         LAYER m3 ;
         RECT  10.0 282.8 10.8 283.6 ;
         LAYER m3 ;
         RECT  67.2 50.4 207.6 51.6 ;
         LAYER m3 ;
         RECT  0.0 295.2 207.6 296.4 ;
         LAYER m3 ;
         RECT  206.9 305.4 207.7 306.2 ;
         LAYER m3 ;
         RECT  0.0 309.6 207.6 310.8 ;
         LAYER m3 ;
         RECT  170.8 167.8 171.6 168.6 ;
         LAYER m3 ;
         RECT  23.2 282.8 24.0 283.6 ;
         LAYER m4 ;
         RECT  187.2 2.4 188.4 423.6 ;
         LAYER m3 ;
         RECT  23.2 165.2 24.0 166.0 ;
         LAYER m3 ;
         RECT  0.0 333.6 207.6 334.8 ;
         LAYER m3 ;
         RECT  0.0 103.2 73.2 104.4 ;
         LAYER m4 ;
         RECT  43.2 2.4 44.4 423.6 ;
         LAYER m3 ;
         RECT  0.0 12.0 207.6 13.2 ;
         LAYER m4 ;
         RECT  115.2 2.4 116.4 423.6 ;
         LAYER m4 ;
         RECT  86.4 2.4 87.6 423.6 ;
         LAYER m3 ;
         RECT  179.7 295.4 180.5 296.2 ;
         LAYER m3 ;
         RECT  0.0 45.6 207.6 46.8 ;
         LAYER m3 ;
         RECT  200.1 347.0 200.9 347.8 ;
         LAYER m3 ;
         RECT  48.0 31.2 207.6 32.4 ;
         LAYER m3 ;
         RECT  77.6 42.4 78.4 43.2 ;
         LAYER m3 ;
         RECT  0.0 381.6 207.6 382.8 ;
         LAYER m3 ;
         RECT  26.4 261.6 121.2 262.8 ;
         LAYER m4 ;
         RECT  52.8 2.4 54.0 423.6 ;
         LAYER m3 ;
         RECT  10.0 204.4 10.8 205.2 ;
         LAYER m4 ;
         RECT  172.8 2.4 174.0 423.6 ;
         LAYER m4 ;
         RECT  24.0 2.4 25.2 423.6 ;
         LAYER m3 ;
         RECT  0.0 338.4 207.6 339.6 ;
         LAYER m3 ;
         RECT  179.7 326.2 180.5 327.0 ;
         LAYER m3 ;
         RECT  189.3 99.6 190.1 100.4 ;
         LAYER m3 ;
         RECT  167.5 248.8 168.3 249.6 ;
         LAYER m3 ;
         RECT  93.1 248.8 93.9 249.6 ;
      END
   END gnd
   OBS
   LAYER  m1 ;
      RECT  188.9 190.4 189.9 191.2 ;
      RECT  191.3 194.8 192.3 195.6 ;
      RECT  191.5 191.2 192.3 191.6 ;
      RECT  190.3 189.4 191.1 189.6 ;
      RECT  193.3 190.0 194.1 194.2 ;
      RECT  189.1 193.4 190.7 194.2 ;
      RECT  191.5 190.4 192.5 191.2 ;
      RECT  186.5 196.4 194.1 197.2 ;
      RECT  186.5 194.8 187.3 196.4 ;
      RECT  189.1 194.8 190.1 195.6 ;
      RECT  189.1 194.2 189.9 194.8 ;
      RECT  191.5 192.4 192.3 194.8 ;
      RECT  191.1 191.6 192.3 192.4 ;
      RECT  186.5 188.6 194.1 189.4 ;
      RECT  186.5 190.0 187.3 194.2 ;
      RECT  189.1 191.2 189.9 193.4 ;
      RECT  190.9 187.2 192.5 188.0 ;
      RECT  193.3 194.8 194.1 196.4 ;
      RECT  188.1 187.2 189.7 188.0 ;
      RECT  188.9 203.2 189.9 202.4 ;
      RECT  191.3 198.8 192.3 198.0 ;
      RECT  191.5 202.4 192.3 202.0 ;
      RECT  190.3 204.2 191.1 204.0 ;
      RECT  193.3 203.6 194.1 199.4 ;
      RECT  189.1 200.2 190.7 199.4 ;
      RECT  191.5 203.2 192.5 202.4 ;
      RECT  186.5 197.2 194.1 196.4 ;
      RECT  186.5 198.8 187.3 197.2 ;
      RECT  189.1 198.8 190.1 198.0 ;
      RECT  189.1 199.4 189.9 198.8 ;
      RECT  191.5 201.2 192.3 198.8 ;
      RECT  191.1 202.0 192.3 201.2 ;
      RECT  186.5 205.0 194.1 204.2 ;
      RECT  186.5 203.6 187.3 199.4 ;
      RECT  189.1 202.4 189.9 200.2 ;
      RECT  190.9 206.4 192.5 205.6 ;
      RECT  193.3 198.8 194.1 197.2 ;
      RECT  188.1 206.4 189.7 205.6 ;
      RECT  188.9 211.2 189.9 212.0 ;
      RECT  191.3 215.6 192.3 216.4 ;
      RECT  191.5 212.0 192.3 212.4 ;
      RECT  190.3 210.2 191.1 210.4 ;
      RECT  193.3 210.8 194.1 215.0 ;
      RECT  189.1 214.2 190.7 215.0 ;
      RECT  191.5 211.2 192.5 212.0 ;
      RECT  186.5 217.2 194.1 218.0 ;
      RECT  186.5 215.6 187.3 217.2 ;
      RECT  189.1 215.6 190.1 216.4 ;
      RECT  189.1 215.0 189.9 215.6 ;
      RECT  191.5 213.2 192.3 215.6 ;
      RECT  191.1 212.4 192.3 213.2 ;
      RECT  186.5 209.4 194.1 210.2 ;
      RECT  186.5 210.8 187.3 215.0 ;
      RECT  189.1 212.0 189.9 214.2 ;
      RECT  190.9 208.0 192.5 208.8 ;
      RECT  193.3 215.6 194.1 217.2 ;
      RECT  188.1 208.0 189.7 208.8 ;
      RECT  188.9 224.0 189.9 223.2 ;
      RECT  191.3 219.6 192.3 218.8 ;
      RECT  191.5 223.2 192.3 222.8 ;
      RECT  190.3 225.0 191.1 224.8 ;
      RECT  193.3 224.4 194.1 220.2 ;
      RECT  189.1 221.0 190.7 220.2 ;
      RECT  191.5 224.0 192.5 223.2 ;
      RECT  186.5 218.0 194.1 217.2 ;
      RECT  186.5 219.6 187.3 218.0 ;
      RECT  189.1 219.6 190.1 218.8 ;
      RECT  189.1 220.2 189.9 219.6 ;
      RECT  191.5 222.0 192.3 219.6 ;
      RECT  191.1 222.8 192.3 222.0 ;
      RECT  186.5 225.8 194.1 225.0 ;
      RECT  186.5 224.4 187.3 220.2 ;
      RECT  189.1 223.2 189.9 221.0 ;
      RECT  190.9 227.2 192.5 226.4 ;
      RECT  193.3 219.6 194.1 218.0 ;
      RECT  188.1 227.2 189.7 226.4 ;
      RECT  188.9 232.0 189.9 232.8 ;
      RECT  191.3 236.4 192.3 237.2 ;
      RECT  191.5 232.8 192.3 233.2 ;
      RECT  190.3 231.0 191.1 231.2 ;
      RECT  193.3 231.6 194.1 235.8 ;
      RECT  189.1 235.0 190.7 235.8 ;
      RECT  191.5 232.0 192.5 232.8 ;
      RECT  186.5 238.0 194.1 238.8 ;
      RECT  186.5 236.4 187.3 238.0 ;
      RECT  189.1 236.4 190.1 237.2 ;
      RECT  189.1 235.8 189.9 236.4 ;
      RECT  191.5 234.0 192.3 236.4 ;
      RECT  191.1 233.2 192.3 234.0 ;
      RECT  186.5 230.2 194.1 231.0 ;
      RECT  186.5 231.6 187.3 235.8 ;
      RECT  189.1 232.8 189.9 235.0 ;
      RECT  190.9 228.8 192.5 229.6 ;
      RECT  193.3 236.4 194.1 238.0 ;
      RECT  188.1 228.8 189.7 229.6 ;
      RECT  188.9 244.8 189.9 244.0 ;
      RECT  191.3 240.4 192.3 239.6 ;
      RECT  191.5 244.0 192.3 243.6 ;
      RECT  190.3 245.8 191.1 245.6 ;
      RECT  193.3 245.2 194.1 241.0 ;
      RECT  189.1 241.8 190.7 241.0 ;
      RECT  191.5 244.8 192.5 244.0 ;
      RECT  186.5 238.8 194.1 238.0 ;
      RECT  186.5 240.4 187.3 238.8 ;
      RECT  189.1 240.4 190.1 239.6 ;
      RECT  189.1 241.0 189.9 240.4 ;
      RECT  191.5 242.8 192.3 240.4 ;
      RECT  191.1 243.6 192.3 242.8 ;
      RECT  186.5 246.6 194.1 245.8 ;
      RECT  186.5 245.2 187.3 241.0 ;
      RECT  189.1 244.0 189.9 241.8 ;
      RECT  190.9 248.0 192.5 247.2 ;
      RECT  193.3 240.4 194.1 238.8 ;
      RECT  188.1 248.0 189.7 247.2 ;
      RECT  188.9 252.8 189.9 253.6 ;
      RECT  191.3 257.2 192.3 258.0 ;
      RECT  191.5 253.6 192.3 254.0 ;
      RECT  190.3 251.8 191.1 252.0 ;
      RECT  193.3 252.4 194.1 256.6 ;
      RECT  189.1 255.8 190.7 256.6 ;
      RECT  191.5 252.8 192.5 253.6 ;
      RECT  186.5 258.8 194.1 259.6 ;
      RECT  186.5 257.2 187.3 258.8 ;
      RECT  189.1 257.2 190.1 258.0 ;
      RECT  189.1 256.6 189.9 257.2 ;
      RECT  191.5 254.8 192.3 257.2 ;
      RECT  191.1 254.0 192.3 254.8 ;
      RECT  186.5 251.0 194.1 251.8 ;
      RECT  186.5 252.4 187.3 256.6 ;
      RECT  189.1 253.6 189.9 255.8 ;
      RECT  190.9 249.6 192.5 250.4 ;
      RECT  193.3 257.2 194.1 258.8 ;
      RECT  188.1 249.6 189.7 250.4 ;
      RECT  188.9 265.6 189.9 264.8 ;
      RECT  191.3 261.2 192.3 260.4 ;
      RECT  191.5 264.8 192.3 264.4 ;
      RECT  190.3 266.6 191.1 266.4 ;
      RECT  193.3 266.0 194.1 261.8 ;
      RECT  189.1 262.6 190.7 261.8 ;
      RECT  191.5 265.6 192.5 264.8 ;
      RECT  186.5 259.6 194.1 258.8 ;
      RECT  186.5 261.2 187.3 259.6 ;
      RECT  189.1 261.2 190.1 260.4 ;
      RECT  189.1 261.8 189.9 261.2 ;
      RECT  191.5 263.6 192.3 261.2 ;
      RECT  191.1 264.4 192.3 263.6 ;
      RECT  186.5 267.4 194.1 266.6 ;
      RECT  186.5 266.0 187.3 261.8 ;
      RECT  189.1 264.8 189.9 262.6 ;
      RECT  190.9 268.8 192.5 268.0 ;
      RECT  193.3 261.2 194.1 259.6 ;
      RECT  188.1 268.8 189.7 268.0 ;
      RECT  188.9 273.6 189.9 274.4 ;
      RECT  191.3 278.0 192.3 278.8 ;
      RECT  191.5 274.4 192.3 274.8 ;
      RECT  190.3 272.6 191.1 272.8 ;
      RECT  193.3 273.2 194.1 277.4 ;
      RECT  189.1 276.6 190.7 277.4 ;
      RECT  191.5 273.6 192.5 274.4 ;
      RECT  186.5 279.6 194.1 280.4 ;
      RECT  186.5 278.0 187.3 279.6 ;
      RECT  189.1 278.0 190.1 278.8 ;
      RECT  189.1 277.4 189.9 278.0 ;
      RECT  191.5 275.6 192.3 278.0 ;
      RECT  191.1 274.8 192.3 275.6 ;
      RECT  186.5 271.8 194.1 272.6 ;
      RECT  186.5 273.2 187.3 277.4 ;
      RECT  189.1 274.4 189.9 276.6 ;
      RECT  190.9 270.4 192.5 271.2 ;
      RECT  193.3 278.0 194.1 279.6 ;
      RECT  188.1 270.4 189.7 271.2 ;
      RECT  188.9 286.4 189.9 285.6 ;
      RECT  191.3 282.0 192.3 281.2 ;
      RECT  191.5 285.6 192.3 285.2 ;
      RECT  190.3 287.4 191.1 287.2 ;
      RECT  193.3 286.8 194.1 282.6 ;
      RECT  189.1 283.4 190.7 282.6 ;
      RECT  191.5 286.4 192.5 285.6 ;
      RECT  186.5 280.4 194.1 279.6 ;
      RECT  186.5 282.0 187.3 280.4 ;
      RECT  189.1 282.0 190.1 281.2 ;
      RECT  189.1 282.6 189.9 282.0 ;
      RECT  191.5 284.4 192.3 282.0 ;
      RECT  191.1 285.2 192.3 284.4 ;
      RECT  186.5 288.2 194.1 287.4 ;
      RECT  186.5 286.8 187.3 282.6 ;
      RECT  189.1 285.6 189.9 283.4 ;
      RECT  190.9 289.6 192.5 288.8 ;
      RECT  193.3 282.0 194.1 280.4 ;
      RECT  188.1 289.6 189.7 288.8 ;
      RECT  188.9 294.4 189.9 295.2 ;
      RECT  191.3 298.8 192.3 299.6 ;
      RECT  191.5 295.2 192.3 295.6 ;
      RECT  190.3 293.4 191.1 293.6 ;
      RECT  193.3 294.0 194.1 298.2 ;
      RECT  189.1 297.4 190.7 298.2 ;
      RECT  191.5 294.4 192.5 295.2 ;
      RECT  186.5 300.4 194.1 301.2 ;
      RECT  186.5 298.8 187.3 300.4 ;
      RECT  189.1 298.8 190.1 299.6 ;
      RECT  189.1 298.2 189.9 298.8 ;
      RECT  191.5 296.4 192.3 298.8 ;
      RECT  191.1 295.6 192.3 296.4 ;
      RECT  186.5 292.6 194.1 293.4 ;
      RECT  186.5 294.0 187.3 298.2 ;
      RECT  189.1 295.2 189.9 297.4 ;
      RECT  190.9 291.2 192.5 292.0 ;
      RECT  193.3 298.8 194.1 300.4 ;
      RECT  188.1 291.2 189.7 292.0 ;
      RECT  188.9 307.2 189.9 306.4 ;
      RECT  191.3 302.8 192.3 302.0 ;
      RECT  191.5 306.4 192.3 306.0 ;
      RECT  190.3 308.2 191.1 308.0 ;
      RECT  193.3 307.6 194.1 303.4 ;
      RECT  189.1 304.2 190.7 303.4 ;
      RECT  191.5 307.2 192.5 306.4 ;
      RECT  186.5 301.2 194.1 300.4 ;
      RECT  186.5 302.8 187.3 301.2 ;
      RECT  189.1 302.8 190.1 302.0 ;
      RECT  189.1 303.4 189.9 302.8 ;
      RECT  191.5 305.2 192.3 302.8 ;
      RECT  191.1 306.0 192.3 305.2 ;
      RECT  186.5 309.0 194.1 308.2 ;
      RECT  186.5 307.6 187.3 303.4 ;
      RECT  189.1 306.4 189.9 304.2 ;
      RECT  190.9 310.4 192.5 309.6 ;
      RECT  193.3 302.8 194.1 301.2 ;
      RECT  188.1 310.4 189.7 309.6 ;
      RECT  188.9 315.2 189.9 316.0 ;
      RECT  191.3 319.6 192.3 320.4 ;
      RECT  191.5 316.0 192.3 316.4 ;
      RECT  190.3 314.2 191.1 314.4 ;
      RECT  193.3 314.8 194.1 319.0 ;
      RECT  189.1 318.2 190.7 319.0 ;
      RECT  191.5 315.2 192.5 316.0 ;
      RECT  186.5 321.2 194.1 322.0 ;
      RECT  186.5 319.6 187.3 321.2 ;
      RECT  189.1 319.6 190.1 320.4 ;
      RECT  189.1 319.0 189.9 319.6 ;
      RECT  191.5 317.2 192.3 319.6 ;
      RECT  191.1 316.4 192.3 317.2 ;
      RECT  186.5 313.4 194.1 314.2 ;
      RECT  186.5 314.8 187.3 319.0 ;
      RECT  189.1 316.0 189.9 318.2 ;
      RECT  190.9 312.0 192.5 312.8 ;
      RECT  193.3 319.6 194.1 321.2 ;
      RECT  188.1 312.0 189.7 312.8 ;
      RECT  188.9 328.0 189.9 327.2 ;
      RECT  191.3 323.6 192.3 322.8 ;
      RECT  191.5 327.2 192.3 326.8 ;
      RECT  190.3 329.0 191.1 328.8 ;
      RECT  193.3 328.4 194.1 324.2 ;
      RECT  189.1 325.0 190.7 324.2 ;
      RECT  191.5 328.0 192.5 327.2 ;
      RECT  186.5 322.0 194.1 321.2 ;
      RECT  186.5 323.6 187.3 322.0 ;
      RECT  189.1 323.6 190.1 322.8 ;
      RECT  189.1 324.2 189.9 323.6 ;
      RECT  191.5 326.0 192.3 323.6 ;
      RECT  191.1 326.8 192.3 326.0 ;
      RECT  186.5 329.8 194.1 329.0 ;
      RECT  186.5 328.4 187.3 324.2 ;
      RECT  189.1 327.2 189.9 325.0 ;
      RECT  190.9 331.2 192.5 330.4 ;
      RECT  193.3 323.6 194.1 322.0 ;
      RECT  188.1 331.2 189.7 330.4 ;
      RECT  188.9 336.0 189.9 336.8 ;
      RECT  191.3 340.4 192.3 341.2 ;
      RECT  191.5 336.8 192.3 337.2 ;
      RECT  190.3 335.0 191.1 335.2 ;
      RECT  193.3 335.6 194.1 339.8 ;
      RECT  189.1 339.0 190.7 339.8 ;
      RECT  191.5 336.0 192.5 336.8 ;
      RECT  186.5 342.0 194.1 342.8 ;
      RECT  186.5 340.4 187.3 342.0 ;
      RECT  189.1 340.4 190.1 341.2 ;
      RECT  189.1 339.8 189.9 340.4 ;
      RECT  191.5 338.0 192.3 340.4 ;
      RECT  191.1 337.2 192.3 338.0 ;
      RECT  186.5 334.2 194.1 335.0 ;
      RECT  186.5 335.6 187.3 339.8 ;
      RECT  189.1 336.8 189.9 339.0 ;
      RECT  190.9 332.8 192.5 333.6 ;
      RECT  193.3 340.4 194.1 342.0 ;
      RECT  188.1 332.8 189.7 333.6 ;
      RECT  188.9 348.8 189.9 348.0 ;
      RECT  191.3 344.4 192.3 343.6 ;
      RECT  191.5 348.0 192.3 347.6 ;
      RECT  190.3 349.8 191.1 349.6 ;
      RECT  193.3 349.2 194.1 345.0 ;
      RECT  189.1 345.8 190.7 345.0 ;
      RECT  191.5 348.8 192.5 348.0 ;
      RECT  186.5 342.8 194.1 342.0 ;
      RECT  186.5 344.4 187.3 342.8 ;
      RECT  189.1 344.4 190.1 343.6 ;
      RECT  189.1 345.0 189.9 344.4 ;
      RECT  191.5 346.8 192.3 344.4 ;
      RECT  191.1 347.6 192.3 346.8 ;
      RECT  186.5 350.6 194.1 349.8 ;
      RECT  186.5 349.2 187.3 345.0 ;
      RECT  189.1 348.0 189.9 345.8 ;
      RECT  190.9 352.0 192.5 351.2 ;
      RECT  193.3 344.4 194.1 342.8 ;
      RECT  188.1 352.0 189.7 351.2 ;
      RECT  195.7 190.4 196.7 191.2 ;
      RECT  198.1 194.8 199.1 195.6 ;
      RECT  198.3 191.2 199.1 191.6 ;
      RECT  197.1 189.4 197.9 189.6 ;
      RECT  200.1 190.0 200.9 194.2 ;
      RECT  195.9 193.4 197.5 194.2 ;
      RECT  198.3 190.4 199.3 191.2 ;
      RECT  193.3 196.4 200.9 197.2 ;
      RECT  193.3 194.8 194.1 196.4 ;
      RECT  195.9 194.8 196.9 195.6 ;
      RECT  195.9 194.2 196.7 194.8 ;
      RECT  198.3 192.4 199.1 194.8 ;
      RECT  197.9 191.6 199.1 192.4 ;
      RECT  193.3 188.6 200.9 189.4 ;
      RECT  193.3 190.0 194.1 194.2 ;
      RECT  195.9 191.2 196.7 193.4 ;
      RECT  197.7 187.2 199.3 188.0 ;
      RECT  200.1 194.8 200.9 196.4 ;
      RECT  194.9 187.2 196.5 188.0 ;
      RECT  195.7 203.2 196.7 202.4 ;
      RECT  198.1 198.8 199.1 198.0 ;
      RECT  198.3 202.4 199.1 202.0 ;
      RECT  197.1 204.2 197.9 204.0 ;
      RECT  200.1 203.6 200.9 199.4 ;
      RECT  195.9 200.2 197.5 199.4 ;
      RECT  198.3 203.2 199.3 202.4 ;
      RECT  193.3 197.2 200.9 196.4 ;
      RECT  193.3 198.8 194.1 197.2 ;
      RECT  195.9 198.8 196.9 198.0 ;
      RECT  195.9 199.4 196.7 198.8 ;
      RECT  198.3 201.2 199.1 198.8 ;
      RECT  197.9 202.0 199.1 201.2 ;
      RECT  193.3 205.0 200.9 204.2 ;
      RECT  193.3 203.6 194.1 199.4 ;
      RECT  195.9 202.4 196.7 200.2 ;
      RECT  197.7 206.4 199.3 205.6 ;
      RECT  200.1 198.8 200.9 197.2 ;
      RECT  194.9 206.4 196.5 205.6 ;
      RECT  195.7 211.2 196.7 212.0 ;
      RECT  198.1 215.6 199.1 216.4 ;
      RECT  198.3 212.0 199.1 212.4 ;
      RECT  197.1 210.2 197.9 210.4 ;
      RECT  200.1 210.8 200.9 215.0 ;
      RECT  195.9 214.2 197.5 215.0 ;
      RECT  198.3 211.2 199.3 212.0 ;
      RECT  193.3 217.2 200.9 218.0 ;
      RECT  193.3 215.6 194.1 217.2 ;
      RECT  195.9 215.6 196.9 216.4 ;
      RECT  195.9 215.0 196.7 215.6 ;
      RECT  198.3 213.2 199.1 215.6 ;
      RECT  197.9 212.4 199.1 213.2 ;
      RECT  193.3 209.4 200.9 210.2 ;
      RECT  193.3 210.8 194.1 215.0 ;
      RECT  195.9 212.0 196.7 214.2 ;
      RECT  197.7 208.0 199.3 208.8 ;
      RECT  200.1 215.6 200.9 217.2 ;
      RECT  194.9 208.0 196.5 208.8 ;
      RECT  195.7 224.0 196.7 223.2 ;
      RECT  198.1 219.6 199.1 218.8 ;
      RECT  198.3 223.2 199.1 222.8 ;
      RECT  197.1 225.0 197.9 224.8 ;
      RECT  200.1 224.4 200.9 220.2 ;
      RECT  195.9 221.0 197.5 220.2 ;
      RECT  198.3 224.0 199.3 223.2 ;
      RECT  193.3 218.0 200.9 217.2 ;
      RECT  193.3 219.6 194.1 218.0 ;
      RECT  195.9 219.6 196.9 218.8 ;
      RECT  195.9 220.2 196.7 219.6 ;
      RECT  198.3 222.0 199.1 219.6 ;
      RECT  197.9 222.8 199.1 222.0 ;
      RECT  193.3 225.8 200.9 225.0 ;
      RECT  193.3 224.4 194.1 220.2 ;
      RECT  195.9 223.2 196.7 221.0 ;
      RECT  197.7 227.2 199.3 226.4 ;
      RECT  200.1 219.6 200.9 218.0 ;
      RECT  194.9 227.2 196.5 226.4 ;
      RECT  195.7 232.0 196.7 232.8 ;
      RECT  198.1 236.4 199.1 237.2 ;
      RECT  198.3 232.8 199.1 233.2 ;
      RECT  197.1 231.0 197.9 231.2 ;
      RECT  200.1 231.6 200.9 235.8 ;
      RECT  195.9 235.0 197.5 235.8 ;
      RECT  198.3 232.0 199.3 232.8 ;
      RECT  193.3 238.0 200.9 238.8 ;
      RECT  193.3 236.4 194.1 238.0 ;
      RECT  195.9 236.4 196.9 237.2 ;
      RECT  195.9 235.8 196.7 236.4 ;
      RECT  198.3 234.0 199.1 236.4 ;
      RECT  197.9 233.2 199.1 234.0 ;
      RECT  193.3 230.2 200.9 231.0 ;
      RECT  193.3 231.6 194.1 235.8 ;
      RECT  195.9 232.8 196.7 235.0 ;
      RECT  197.7 228.8 199.3 229.6 ;
      RECT  200.1 236.4 200.9 238.0 ;
      RECT  194.9 228.8 196.5 229.6 ;
      RECT  195.7 244.8 196.7 244.0 ;
      RECT  198.1 240.4 199.1 239.6 ;
      RECT  198.3 244.0 199.1 243.6 ;
      RECT  197.1 245.8 197.9 245.6 ;
      RECT  200.1 245.2 200.9 241.0 ;
      RECT  195.9 241.8 197.5 241.0 ;
      RECT  198.3 244.8 199.3 244.0 ;
      RECT  193.3 238.8 200.9 238.0 ;
      RECT  193.3 240.4 194.1 238.8 ;
      RECT  195.9 240.4 196.9 239.6 ;
      RECT  195.9 241.0 196.7 240.4 ;
      RECT  198.3 242.8 199.1 240.4 ;
      RECT  197.9 243.6 199.1 242.8 ;
      RECT  193.3 246.6 200.9 245.8 ;
      RECT  193.3 245.2 194.1 241.0 ;
      RECT  195.9 244.0 196.7 241.8 ;
      RECT  197.7 248.0 199.3 247.2 ;
      RECT  200.1 240.4 200.9 238.8 ;
      RECT  194.9 248.0 196.5 247.2 ;
      RECT  195.7 252.8 196.7 253.6 ;
      RECT  198.1 257.2 199.1 258.0 ;
      RECT  198.3 253.6 199.1 254.0 ;
      RECT  197.1 251.8 197.9 252.0 ;
      RECT  200.1 252.4 200.9 256.6 ;
      RECT  195.9 255.8 197.5 256.6 ;
      RECT  198.3 252.8 199.3 253.6 ;
      RECT  193.3 258.8 200.9 259.6 ;
      RECT  193.3 257.2 194.1 258.8 ;
      RECT  195.9 257.2 196.9 258.0 ;
      RECT  195.9 256.6 196.7 257.2 ;
      RECT  198.3 254.8 199.1 257.2 ;
      RECT  197.9 254.0 199.1 254.8 ;
      RECT  193.3 251.0 200.9 251.8 ;
      RECT  193.3 252.4 194.1 256.6 ;
      RECT  195.9 253.6 196.7 255.8 ;
      RECT  197.7 249.6 199.3 250.4 ;
      RECT  200.1 257.2 200.9 258.8 ;
      RECT  194.9 249.6 196.5 250.4 ;
      RECT  195.7 265.6 196.7 264.8 ;
      RECT  198.1 261.2 199.1 260.4 ;
      RECT  198.3 264.8 199.1 264.4 ;
      RECT  197.1 266.6 197.9 266.4 ;
      RECT  200.1 266.0 200.9 261.8 ;
      RECT  195.9 262.6 197.5 261.8 ;
      RECT  198.3 265.6 199.3 264.8 ;
      RECT  193.3 259.6 200.9 258.8 ;
      RECT  193.3 261.2 194.1 259.6 ;
      RECT  195.9 261.2 196.9 260.4 ;
      RECT  195.9 261.8 196.7 261.2 ;
      RECT  198.3 263.6 199.1 261.2 ;
      RECT  197.9 264.4 199.1 263.6 ;
      RECT  193.3 267.4 200.9 266.6 ;
      RECT  193.3 266.0 194.1 261.8 ;
      RECT  195.9 264.8 196.7 262.6 ;
      RECT  197.7 268.8 199.3 268.0 ;
      RECT  200.1 261.2 200.9 259.6 ;
      RECT  194.9 268.8 196.5 268.0 ;
      RECT  195.7 273.6 196.7 274.4 ;
      RECT  198.1 278.0 199.1 278.8 ;
      RECT  198.3 274.4 199.1 274.8 ;
      RECT  197.1 272.6 197.9 272.8 ;
      RECT  200.1 273.2 200.9 277.4 ;
      RECT  195.9 276.6 197.5 277.4 ;
      RECT  198.3 273.6 199.3 274.4 ;
      RECT  193.3 279.6 200.9 280.4 ;
      RECT  193.3 278.0 194.1 279.6 ;
      RECT  195.9 278.0 196.9 278.8 ;
      RECT  195.9 277.4 196.7 278.0 ;
      RECT  198.3 275.6 199.1 278.0 ;
      RECT  197.9 274.8 199.1 275.6 ;
      RECT  193.3 271.8 200.9 272.6 ;
      RECT  193.3 273.2 194.1 277.4 ;
      RECT  195.9 274.4 196.7 276.6 ;
      RECT  197.7 270.4 199.3 271.2 ;
      RECT  200.1 278.0 200.9 279.6 ;
      RECT  194.9 270.4 196.5 271.2 ;
      RECT  195.7 286.4 196.7 285.6 ;
      RECT  198.1 282.0 199.1 281.2 ;
      RECT  198.3 285.6 199.1 285.2 ;
      RECT  197.1 287.4 197.9 287.2 ;
      RECT  200.1 286.8 200.9 282.6 ;
      RECT  195.9 283.4 197.5 282.6 ;
      RECT  198.3 286.4 199.3 285.6 ;
      RECT  193.3 280.4 200.9 279.6 ;
      RECT  193.3 282.0 194.1 280.4 ;
      RECT  195.9 282.0 196.9 281.2 ;
      RECT  195.9 282.6 196.7 282.0 ;
      RECT  198.3 284.4 199.1 282.0 ;
      RECT  197.9 285.2 199.1 284.4 ;
      RECT  193.3 288.2 200.9 287.4 ;
      RECT  193.3 286.8 194.1 282.6 ;
      RECT  195.9 285.6 196.7 283.4 ;
      RECT  197.7 289.6 199.3 288.8 ;
      RECT  200.1 282.0 200.9 280.4 ;
      RECT  194.9 289.6 196.5 288.8 ;
      RECT  195.7 294.4 196.7 295.2 ;
      RECT  198.1 298.8 199.1 299.6 ;
      RECT  198.3 295.2 199.1 295.6 ;
      RECT  197.1 293.4 197.9 293.6 ;
      RECT  200.1 294.0 200.9 298.2 ;
      RECT  195.9 297.4 197.5 298.2 ;
      RECT  198.3 294.4 199.3 295.2 ;
      RECT  193.3 300.4 200.9 301.2 ;
      RECT  193.3 298.8 194.1 300.4 ;
      RECT  195.9 298.8 196.9 299.6 ;
      RECT  195.9 298.2 196.7 298.8 ;
      RECT  198.3 296.4 199.1 298.8 ;
      RECT  197.9 295.6 199.1 296.4 ;
      RECT  193.3 292.6 200.9 293.4 ;
      RECT  193.3 294.0 194.1 298.2 ;
      RECT  195.9 295.2 196.7 297.4 ;
      RECT  197.7 291.2 199.3 292.0 ;
      RECT  200.1 298.8 200.9 300.4 ;
      RECT  194.9 291.2 196.5 292.0 ;
      RECT  195.7 307.2 196.7 306.4 ;
      RECT  198.1 302.8 199.1 302.0 ;
      RECT  198.3 306.4 199.1 306.0 ;
      RECT  197.1 308.2 197.9 308.0 ;
      RECT  200.1 307.6 200.9 303.4 ;
      RECT  195.9 304.2 197.5 303.4 ;
      RECT  198.3 307.2 199.3 306.4 ;
      RECT  193.3 301.2 200.9 300.4 ;
      RECT  193.3 302.8 194.1 301.2 ;
      RECT  195.9 302.8 196.9 302.0 ;
      RECT  195.9 303.4 196.7 302.8 ;
      RECT  198.3 305.2 199.1 302.8 ;
      RECT  197.9 306.0 199.1 305.2 ;
      RECT  193.3 309.0 200.9 308.2 ;
      RECT  193.3 307.6 194.1 303.4 ;
      RECT  195.9 306.4 196.7 304.2 ;
      RECT  197.7 310.4 199.3 309.6 ;
      RECT  200.1 302.8 200.9 301.2 ;
      RECT  194.9 310.4 196.5 309.6 ;
      RECT  195.7 315.2 196.7 316.0 ;
      RECT  198.1 319.6 199.1 320.4 ;
      RECT  198.3 316.0 199.1 316.4 ;
      RECT  197.1 314.2 197.9 314.4 ;
      RECT  200.1 314.8 200.9 319.0 ;
      RECT  195.9 318.2 197.5 319.0 ;
      RECT  198.3 315.2 199.3 316.0 ;
      RECT  193.3 321.2 200.9 322.0 ;
      RECT  193.3 319.6 194.1 321.2 ;
      RECT  195.9 319.6 196.9 320.4 ;
      RECT  195.9 319.0 196.7 319.6 ;
      RECT  198.3 317.2 199.1 319.6 ;
      RECT  197.9 316.4 199.1 317.2 ;
      RECT  193.3 313.4 200.9 314.2 ;
      RECT  193.3 314.8 194.1 319.0 ;
      RECT  195.9 316.0 196.7 318.2 ;
      RECT  197.7 312.0 199.3 312.8 ;
      RECT  200.1 319.6 200.9 321.2 ;
      RECT  194.9 312.0 196.5 312.8 ;
      RECT  195.7 328.0 196.7 327.2 ;
      RECT  198.1 323.6 199.1 322.8 ;
      RECT  198.3 327.2 199.1 326.8 ;
      RECT  197.1 329.0 197.9 328.8 ;
      RECT  200.1 328.4 200.9 324.2 ;
      RECT  195.9 325.0 197.5 324.2 ;
      RECT  198.3 328.0 199.3 327.2 ;
      RECT  193.3 322.0 200.9 321.2 ;
      RECT  193.3 323.6 194.1 322.0 ;
      RECT  195.9 323.6 196.9 322.8 ;
      RECT  195.9 324.2 196.7 323.6 ;
      RECT  198.3 326.0 199.1 323.6 ;
      RECT  197.9 326.8 199.1 326.0 ;
      RECT  193.3 329.8 200.9 329.0 ;
      RECT  193.3 328.4 194.1 324.2 ;
      RECT  195.9 327.2 196.7 325.0 ;
      RECT  197.7 331.2 199.3 330.4 ;
      RECT  200.1 323.6 200.9 322.0 ;
      RECT  194.9 331.2 196.5 330.4 ;
      RECT  195.7 336.0 196.7 336.8 ;
      RECT  198.1 340.4 199.1 341.2 ;
      RECT  198.3 336.8 199.1 337.2 ;
      RECT  197.1 335.0 197.9 335.2 ;
      RECT  200.1 335.6 200.9 339.8 ;
      RECT  195.9 339.0 197.5 339.8 ;
      RECT  198.3 336.0 199.3 336.8 ;
      RECT  193.3 342.0 200.9 342.8 ;
      RECT  193.3 340.4 194.1 342.0 ;
      RECT  195.9 340.4 196.9 341.2 ;
      RECT  195.9 339.8 196.7 340.4 ;
      RECT  198.3 338.0 199.1 340.4 ;
      RECT  197.9 337.2 199.1 338.0 ;
      RECT  193.3 334.2 200.9 335.0 ;
      RECT  193.3 335.6 194.1 339.8 ;
      RECT  195.9 336.8 196.7 339.0 ;
      RECT  197.7 332.8 199.3 333.6 ;
      RECT  200.1 340.4 200.9 342.0 ;
      RECT  194.9 332.8 196.5 333.6 ;
      RECT  195.7 348.8 196.7 348.0 ;
      RECT  198.1 344.4 199.1 343.6 ;
      RECT  198.3 348.0 199.1 347.6 ;
      RECT  197.1 349.8 197.9 349.6 ;
      RECT  200.1 349.2 200.9 345.0 ;
      RECT  195.9 345.8 197.5 345.0 ;
      RECT  198.3 348.8 199.3 348.0 ;
      RECT  193.3 342.8 200.9 342.0 ;
      RECT  193.3 344.4 194.1 342.8 ;
      RECT  195.9 344.4 196.9 343.6 ;
      RECT  195.9 345.0 196.7 344.4 ;
      RECT  198.3 346.8 199.1 344.4 ;
      RECT  197.9 347.6 199.1 346.8 ;
      RECT  193.3 350.6 200.9 349.8 ;
      RECT  193.3 349.2 194.1 345.0 ;
      RECT  195.9 348.0 196.7 345.8 ;
      RECT  197.7 352.0 199.3 351.2 ;
      RECT  200.1 344.4 200.9 342.8 ;
      RECT  194.9 352.0 196.5 351.2 ;
      RECT  186.9 188.6 200.5 189.4 ;
      RECT  186.9 204.2 200.5 205.0 ;
      RECT  186.9 209.4 200.5 210.2 ;
      RECT  186.9 225.0 200.5 225.8 ;
      RECT  186.9 230.2 200.5 231.0 ;
      RECT  186.9 245.8 200.5 246.6 ;
      RECT  186.9 251.0 200.5 251.8 ;
      RECT  186.9 266.6 200.5 267.4 ;
      RECT  186.9 271.8 200.5 272.6 ;
      RECT  186.9 287.4 200.5 288.2 ;
      RECT  186.9 292.6 200.5 293.4 ;
      RECT  186.9 308.2 200.5 309.0 ;
      RECT  186.9 313.4 200.5 314.2 ;
      RECT  186.9 329.0 200.5 329.8 ;
      RECT  186.9 334.2 200.5 335.0 ;
      RECT  186.9 349.8 200.5 350.6 ;
      RECT  182.1 169.6 183.1 170.4 ;
      RECT  184.5 174.0 185.5 174.8 ;
      RECT  184.7 170.4 185.5 170.8 ;
      RECT  183.5 168.6 184.3 168.8 ;
      RECT  186.5 169.2 187.3 173.4 ;
      RECT  182.3 172.6 183.9 173.4 ;
      RECT  184.7 169.6 185.7 170.4 ;
      RECT  182.1 166.4 182.9 167.2 ;
      RECT  179.7 175.6 187.3 176.4 ;
      RECT  179.7 174.0 180.5 175.6 ;
      RECT  182.3 174.0 183.3 174.8 ;
      RECT  182.3 173.4 183.1 174.0 ;
      RECT  184.7 171.6 185.5 174.0 ;
      RECT  184.3 170.8 185.5 171.6 ;
      RECT  179.7 167.8 187.3 168.6 ;
      RECT  184.9 166.4 185.7 167.2 ;
      RECT  179.7 169.2 180.5 173.4 ;
      RECT  182.3 170.4 183.1 172.6 ;
      RECT  186.5 174.0 187.3 175.6 ;
      RECT  182.1 182.4 183.1 181.6 ;
      RECT  184.5 178.0 185.5 177.2 ;
      RECT  184.7 181.6 185.5 181.2 ;
      RECT  183.5 183.4 184.3 183.2 ;
      RECT  186.5 182.8 187.3 178.6 ;
      RECT  182.3 179.4 183.9 178.6 ;
      RECT  184.5 177.2 185.3 176.4 ;
      RECT  184.7 182.4 185.7 181.6 ;
      RECT  179.7 176.4 187.3 175.6 ;
      RECT  179.7 178.0 180.5 176.4 ;
      RECT  182.3 178.0 183.3 177.2 ;
      RECT  182.3 178.6 183.1 178.0 ;
      RECT  184.7 180.4 185.5 178.0 ;
      RECT  184.3 181.2 185.5 180.4 ;
      RECT  179.7 184.2 187.3 183.4 ;
      RECT  179.7 182.8 180.5 178.6 ;
      RECT  182.3 181.6 183.1 179.4 ;
      RECT  184.1 185.6 185.7 184.8 ;
      RECT  186.5 178.0 187.3 176.4 ;
      RECT  181.3 185.6 182.9 184.8 ;
      RECT  182.1 190.4 183.1 191.2 ;
      RECT  184.5 194.8 185.5 195.6 ;
      RECT  184.7 191.2 185.5 191.6 ;
      RECT  183.5 189.4 184.3 189.6 ;
      RECT  186.5 190.0 187.3 194.2 ;
      RECT  182.3 193.4 183.9 194.2 ;
      RECT  184.5 195.6 185.3 196.4 ;
      RECT  184.7 190.4 185.7 191.2 ;
      RECT  179.7 196.4 187.3 197.2 ;
      RECT  179.7 194.8 180.5 196.4 ;
      RECT  182.3 194.8 183.3 195.6 ;
      RECT  182.3 194.2 183.1 194.8 ;
      RECT  184.7 192.4 185.5 194.8 ;
      RECT  184.3 191.6 185.5 192.4 ;
      RECT  179.7 188.6 187.3 189.4 ;
      RECT  179.7 190.0 180.5 194.2 ;
      RECT  182.3 191.2 183.1 193.4 ;
      RECT  184.1 187.2 185.7 188.0 ;
      RECT  186.5 194.8 187.3 196.4 ;
      RECT  181.3 187.2 182.9 188.0 ;
      RECT  182.1 203.2 183.1 202.4 ;
      RECT  184.5 198.8 185.5 198.0 ;
      RECT  184.7 202.4 185.5 202.0 ;
      RECT  183.5 204.2 184.3 204.0 ;
      RECT  186.5 203.6 187.3 199.4 ;
      RECT  182.3 200.2 183.9 199.4 ;
      RECT  184.5 198.0 185.3 197.2 ;
      RECT  184.7 203.2 185.7 202.4 ;
      RECT  179.7 197.2 187.3 196.4 ;
      RECT  179.7 198.8 180.5 197.2 ;
      RECT  182.3 198.8 183.3 198.0 ;
      RECT  182.3 199.4 183.1 198.8 ;
      RECT  184.7 201.2 185.5 198.8 ;
      RECT  184.3 202.0 185.5 201.2 ;
      RECT  179.7 205.0 187.3 204.2 ;
      RECT  179.7 203.6 180.5 199.4 ;
      RECT  182.3 202.4 183.1 200.2 ;
      RECT  184.1 206.4 185.7 205.6 ;
      RECT  186.5 198.8 187.3 197.2 ;
      RECT  181.3 206.4 182.9 205.6 ;
      RECT  182.1 211.2 183.1 212.0 ;
      RECT  184.5 215.6 185.5 216.4 ;
      RECT  184.7 212.0 185.5 212.4 ;
      RECT  183.5 210.2 184.3 210.4 ;
      RECT  186.5 210.8 187.3 215.0 ;
      RECT  182.3 214.2 183.9 215.0 ;
      RECT  184.5 216.4 185.3 217.2 ;
      RECT  184.7 211.2 185.7 212.0 ;
      RECT  179.7 217.2 187.3 218.0 ;
      RECT  179.7 215.6 180.5 217.2 ;
      RECT  182.3 215.6 183.3 216.4 ;
      RECT  182.3 215.0 183.1 215.6 ;
      RECT  184.7 213.2 185.5 215.6 ;
      RECT  184.3 212.4 185.5 213.2 ;
      RECT  179.7 209.4 187.3 210.2 ;
      RECT  179.7 210.8 180.5 215.0 ;
      RECT  182.3 212.0 183.1 214.2 ;
      RECT  184.1 208.0 185.7 208.8 ;
      RECT  186.5 215.6 187.3 217.2 ;
      RECT  181.3 208.0 182.9 208.8 ;
      RECT  182.1 224.0 183.1 223.2 ;
      RECT  184.5 219.6 185.5 218.8 ;
      RECT  184.7 223.2 185.5 222.8 ;
      RECT  183.5 225.0 184.3 224.8 ;
      RECT  186.5 224.4 187.3 220.2 ;
      RECT  182.3 221.0 183.9 220.2 ;
      RECT  184.5 218.8 185.3 218.0 ;
      RECT  184.7 224.0 185.7 223.2 ;
      RECT  179.7 218.0 187.3 217.2 ;
      RECT  179.7 219.6 180.5 218.0 ;
      RECT  182.3 219.6 183.3 218.8 ;
      RECT  182.3 220.2 183.1 219.6 ;
      RECT  184.7 222.0 185.5 219.6 ;
      RECT  184.3 222.8 185.5 222.0 ;
      RECT  179.7 225.8 187.3 225.0 ;
      RECT  179.7 224.4 180.5 220.2 ;
      RECT  182.3 223.2 183.1 221.0 ;
      RECT  184.1 227.2 185.7 226.4 ;
      RECT  186.5 219.6 187.3 218.0 ;
      RECT  181.3 227.2 182.9 226.4 ;
      RECT  182.1 232.0 183.1 232.8 ;
      RECT  184.5 236.4 185.5 237.2 ;
      RECT  184.7 232.8 185.5 233.2 ;
      RECT  183.5 231.0 184.3 231.2 ;
      RECT  186.5 231.6 187.3 235.8 ;
      RECT  182.3 235.0 183.9 235.8 ;
      RECT  184.5 237.2 185.3 238.0 ;
      RECT  184.7 232.0 185.7 232.8 ;
      RECT  179.7 238.0 187.3 238.8 ;
      RECT  179.7 236.4 180.5 238.0 ;
      RECT  182.3 236.4 183.3 237.2 ;
      RECT  182.3 235.8 183.1 236.4 ;
      RECT  184.7 234.0 185.5 236.4 ;
      RECT  184.3 233.2 185.5 234.0 ;
      RECT  179.7 230.2 187.3 231.0 ;
      RECT  179.7 231.6 180.5 235.8 ;
      RECT  182.3 232.8 183.1 235.0 ;
      RECT  184.1 228.8 185.7 229.6 ;
      RECT  186.5 236.4 187.3 238.0 ;
      RECT  181.3 228.8 182.9 229.6 ;
      RECT  182.1 244.8 183.1 244.0 ;
      RECT  184.5 240.4 185.5 239.6 ;
      RECT  184.7 244.0 185.5 243.6 ;
      RECT  183.5 245.8 184.3 245.6 ;
      RECT  186.5 245.2 187.3 241.0 ;
      RECT  182.3 241.8 183.9 241.0 ;
      RECT  184.5 239.6 185.3 238.8 ;
      RECT  184.7 244.8 185.7 244.0 ;
      RECT  179.7 238.8 187.3 238.0 ;
      RECT  179.7 240.4 180.5 238.8 ;
      RECT  182.3 240.4 183.3 239.6 ;
      RECT  182.3 241.0 183.1 240.4 ;
      RECT  184.7 242.8 185.5 240.4 ;
      RECT  184.3 243.6 185.5 242.8 ;
      RECT  179.7 246.6 187.3 245.8 ;
      RECT  179.7 245.2 180.5 241.0 ;
      RECT  182.3 244.0 183.1 241.8 ;
      RECT  184.1 248.0 185.7 247.2 ;
      RECT  186.5 240.4 187.3 238.8 ;
      RECT  181.3 248.0 182.9 247.2 ;
      RECT  182.1 252.8 183.1 253.6 ;
      RECT  184.5 257.2 185.5 258.0 ;
      RECT  184.7 253.6 185.5 254.0 ;
      RECT  183.5 251.8 184.3 252.0 ;
      RECT  186.5 252.4 187.3 256.6 ;
      RECT  182.3 255.8 183.9 256.6 ;
      RECT  184.5 258.0 185.3 258.8 ;
      RECT  184.7 252.8 185.7 253.6 ;
      RECT  179.7 258.8 187.3 259.6 ;
      RECT  179.7 257.2 180.5 258.8 ;
      RECT  182.3 257.2 183.3 258.0 ;
      RECT  182.3 256.6 183.1 257.2 ;
      RECT  184.7 254.8 185.5 257.2 ;
      RECT  184.3 254.0 185.5 254.8 ;
      RECT  179.7 251.0 187.3 251.8 ;
      RECT  179.7 252.4 180.5 256.6 ;
      RECT  182.3 253.6 183.1 255.8 ;
      RECT  184.1 249.6 185.7 250.4 ;
      RECT  186.5 257.2 187.3 258.8 ;
      RECT  181.3 249.6 182.9 250.4 ;
      RECT  182.1 265.6 183.1 264.8 ;
      RECT  184.5 261.2 185.5 260.4 ;
      RECT  184.7 264.8 185.5 264.4 ;
      RECT  183.5 266.6 184.3 266.4 ;
      RECT  186.5 266.0 187.3 261.8 ;
      RECT  182.3 262.6 183.9 261.8 ;
      RECT  184.5 260.4 185.3 259.6 ;
      RECT  184.7 265.6 185.7 264.8 ;
      RECT  179.7 259.6 187.3 258.8 ;
      RECT  179.7 261.2 180.5 259.6 ;
      RECT  182.3 261.2 183.3 260.4 ;
      RECT  182.3 261.8 183.1 261.2 ;
      RECT  184.7 263.6 185.5 261.2 ;
      RECT  184.3 264.4 185.5 263.6 ;
      RECT  179.7 267.4 187.3 266.6 ;
      RECT  179.7 266.0 180.5 261.8 ;
      RECT  182.3 264.8 183.1 262.6 ;
      RECT  184.1 268.8 185.7 268.0 ;
      RECT  186.5 261.2 187.3 259.6 ;
      RECT  181.3 268.8 182.9 268.0 ;
      RECT  182.1 273.6 183.1 274.4 ;
      RECT  184.5 278.0 185.5 278.8 ;
      RECT  184.7 274.4 185.5 274.8 ;
      RECT  183.5 272.6 184.3 272.8 ;
      RECT  186.5 273.2 187.3 277.4 ;
      RECT  182.3 276.6 183.9 277.4 ;
      RECT  184.5 278.8 185.3 279.6 ;
      RECT  184.7 273.6 185.7 274.4 ;
      RECT  179.7 279.6 187.3 280.4 ;
      RECT  179.7 278.0 180.5 279.6 ;
      RECT  182.3 278.0 183.3 278.8 ;
      RECT  182.3 277.4 183.1 278.0 ;
      RECT  184.7 275.6 185.5 278.0 ;
      RECT  184.3 274.8 185.5 275.6 ;
      RECT  179.7 271.8 187.3 272.6 ;
      RECT  179.7 273.2 180.5 277.4 ;
      RECT  182.3 274.4 183.1 276.6 ;
      RECT  184.1 270.4 185.7 271.2 ;
      RECT  186.5 278.0 187.3 279.6 ;
      RECT  181.3 270.4 182.9 271.2 ;
      RECT  182.1 286.4 183.1 285.6 ;
      RECT  184.5 282.0 185.5 281.2 ;
      RECT  184.7 285.6 185.5 285.2 ;
      RECT  183.5 287.4 184.3 287.2 ;
      RECT  186.5 286.8 187.3 282.6 ;
      RECT  182.3 283.4 183.9 282.6 ;
      RECT  184.5 281.2 185.3 280.4 ;
      RECT  184.7 286.4 185.7 285.6 ;
      RECT  179.7 280.4 187.3 279.6 ;
      RECT  179.7 282.0 180.5 280.4 ;
      RECT  182.3 282.0 183.3 281.2 ;
      RECT  182.3 282.6 183.1 282.0 ;
      RECT  184.7 284.4 185.5 282.0 ;
      RECT  184.3 285.2 185.5 284.4 ;
      RECT  179.7 288.2 187.3 287.4 ;
      RECT  179.7 286.8 180.5 282.6 ;
      RECT  182.3 285.6 183.1 283.4 ;
      RECT  184.1 289.6 185.7 288.8 ;
      RECT  186.5 282.0 187.3 280.4 ;
      RECT  181.3 289.6 182.9 288.8 ;
      RECT  182.1 294.4 183.1 295.2 ;
      RECT  184.5 298.8 185.5 299.6 ;
      RECT  184.7 295.2 185.5 295.6 ;
      RECT  183.5 293.4 184.3 293.6 ;
      RECT  186.5 294.0 187.3 298.2 ;
      RECT  182.3 297.4 183.9 298.2 ;
      RECT  184.5 299.6 185.3 300.4 ;
      RECT  184.7 294.4 185.7 295.2 ;
      RECT  179.7 300.4 187.3 301.2 ;
      RECT  179.7 298.8 180.5 300.4 ;
      RECT  182.3 298.8 183.3 299.6 ;
      RECT  182.3 298.2 183.1 298.8 ;
      RECT  184.7 296.4 185.5 298.8 ;
      RECT  184.3 295.6 185.5 296.4 ;
      RECT  179.7 292.6 187.3 293.4 ;
      RECT  179.7 294.0 180.5 298.2 ;
      RECT  182.3 295.2 183.1 297.4 ;
      RECT  184.1 291.2 185.7 292.0 ;
      RECT  186.5 298.8 187.3 300.4 ;
      RECT  181.3 291.2 182.9 292.0 ;
      RECT  182.1 307.2 183.1 306.4 ;
      RECT  184.5 302.8 185.5 302.0 ;
      RECT  184.7 306.4 185.5 306.0 ;
      RECT  183.5 308.2 184.3 308.0 ;
      RECT  186.5 307.6 187.3 303.4 ;
      RECT  182.3 304.2 183.9 303.4 ;
      RECT  184.5 302.0 185.3 301.2 ;
      RECT  184.7 307.2 185.7 306.4 ;
      RECT  179.7 301.2 187.3 300.4 ;
      RECT  179.7 302.8 180.5 301.2 ;
      RECT  182.3 302.8 183.3 302.0 ;
      RECT  182.3 303.4 183.1 302.8 ;
      RECT  184.7 305.2 185.5 302.8 ;
      RECT  184.3 306.0 185.5 305.2 ;
      RECT  179.7 309.0 187.3 308.2 ;
      RECT  179.7 307.6 180.5 303.4 ;
      RECT  182.3 306.4 183.1 304.2 ;
      RECT  184.1 310.4 185.7 309.6 ;
      RECT  186.5 302.8 187.3 301.2 ;
      RECT  181.3 310.4 182.9 309.6 ;
      RECT  182.1 315.2 183.1 316.0 ;
      RECT  184.5 319.6 185.5 320.4 ;
      RECT  184.7 316.0 185.5 316.4 ;
      RECT  183.5 314.2 184.3 314.4 ;
      RECT  186.5 314.8 187.3 319.0 ;
      RECT  182.3 318.2 183.9 319.0 ;
      RECT  184.5 320.4 185.3 321.2 ;
      RECT  184.7 315.2 185.7 316.0 ;
      RECT  179.7 321.2 187.3 322.0 ;
      RECT  179.7 319.6 180.5 321.2 ;
      RECT  182.3 319.6 183.3 320.4 ;
      RECT  182.3 319.0 183.1 319.6 ;
      RECT  184.7 317.2 185.5 319.6 ;
      RECT  184.3 316.4 185.5 317.2 ;
      RECT  179.7 313.4 187.3 314.2 ;
      RECT  179.7 314.8 180.5 319.0 ;
      RECT  182.3 316.0 183.1 318.2 ;
      RECT  184.1 312.0 185.7 312.8 ;
      RECT  186.5 319.6 187.3 321.2 ;
      RECT  181.3 312.0 182.9 312.8 ;
      RECT  182.1 328.0 183.1 327.2 ;
      RECT  184.5 323.6 185.5 322.8 ;
      RECT  184.7 327.2 185.5 326.8 ;
      RECT  183.5 329.0 184.3 328.8 ;
      RECT  186.5 328.4 187.3 324.2 ;
      RECT  182.3 325.0 183.9 324.2 ;
      RECT  184.5 322.8 185.3 322.0 ;
      RECT  184.7 328.0 185.7 327.2 ;
      RECT  179.7 322.0 187.3 321.2 ;
      RECT  179.7 323.6 180.5 322.0 ;
      RECT  182.3 323.6 183.3 322.8 ;
      RECT  182.3 324.2 183.1 323.6 ;
      RECT  184.7 326.0 185.5 323.6 ;
      RECT  184.3 326.8 185.5 326.0 ;
      RECT  179.7 329.8 187.3 329.0 ;
      RECT  179.7 328.4 180.5 324.2 ;
      RECT  182.3 327.2 183.1 325.0 ;
      RECT  184.1 331.2 185.7 330.4 ;
      RECT  186.5 323.6 187.3 322.0 ;
      RECT  181.3 331.2 182.9 330.4 ;
      RECT  182.1 336.0 183.1 336.8 ;
      RECT  184.5 340.4 185.5 341.2 ;
      RECT  184.7 336.8 185.5 337.2 ;
      RECT  183.5 335.0 184.3 335.2 ;
      RECT  186.5 335.6 187.3 339.8 ;
      RECT  182.3 339.0 183.9 339.8 ;
      RECT  184.5 341.2 185.3 342.0 ;
      RECT  184.7 336.0 185.7 336.8 ;
      RECT  179.7 342.0 187.3 342.8 ;
      RECT  179.7 340.4 180.5 342.0 ;
      RECT  182.3 340.4 183.3 341.2 ;
      RECT  182.3 339.8 183.1 340.4 ;
      RECT  184.7 338.0 185.5 340.4 ;
      RECT  184.3 337.2 185.5 338.0 ;
      RECT  179.7 334.2 187.3 335.0 ;
      RECT  179.7 335.6 180.5 339.8 ;
      RECT  182.3 336.8 183.1 339.0 ;
      RECT  184.1 332.8 185.7 333.6 ;
      RECT  186.5 340.4 187.3 342.0 ;
      RECT  181.3 332.8 182.9 333.6 ;
      RECT  182.1 348.8 183.1 348.0 ;
      RECT  184.5 344.4 185.5 343.6 ;
      RECT  184.7 348.0 185.5 347.6 ;
      RECT  183.5 349.8 184.3 349.6 ;
      RECT  186.5 349.2 187.3 345.0 ;
      RECT  182.3 345.8 183.9 345.0 ;
      RECT  184.5 343.6 185.3 342.8 ;
      RECT  184.7 348.8 185.7 348.0 ;
      RECT  179.7 342.8 187.3 342.0 ;
      RECT  179.7 344.4 180.5 342.8 ;
      RECT  182.3 344.4 183.3 343.6 ;
      RECT  182.3 345.0 183.1 344.4 ;
      RECT  184.7 346.8 185.5 344.4 ;
      RECT  184.3 347.6 185.5 346.8 ;
      RECT  179.7 350.6 187.3 349.8 ;
      RECT  179.7 349.2 180.5 345.0 ;
      RECT  182.3 348.0 183.1 345.8 ;
      RECT  184.1 352.0 185.7 351.2 ;
      RECT  186.5 344.4 187.3 342.8 ;
      RECT  181.3 352.0 182.9 351.2 ;
      RECT  182.1 356.8 183.1 357.6 ;
      RECT  184.5 361.2 185.5 362.0 ;
      RECT  184.7 357.6 185.5 358.0 ;
      RECT  183.5 355.8 184.3 356.0 ;
      RECT  186.5 356.4 187.3 360.6 ;
      RECT  182.3 359.8 183.9 360.6 ;
      RECT  184.7 356.8 185.7 357.6 ;
      RECT  182.1 353.6 182.9 354.4 ;
      RECT  179.7 362.8 187.3 363.6 ;
      RECT  179.7 361.2 180.5 362.8 ;
      RECT  182.3 361.2 183.3 362.0 ;
      RECT  182.3 360.6 183.1 361.2 ;
      RECT  184.7 358.8 185.5 361.2 ;
      RECT  184.3 358.0 185.5 358.8 ;
      RECT  179.7 355.0 187.3 355.8 ;
      RECT  184.9 353.6 185.7 354.4 ;
      RECT  179.7 356.4 180.5 360.6 ;
      RECT  182.3 357.6 183.1 359.8 ;
      RECT  186.5 361.2 187.3 362.8 ;
      RECT  180.1 167.8 186.9 168.6 ;
      RECT  180.1 183.4 186.9 184.2 ;
      RECT  180.1 188.6 186.9 189.4 ;
      RECT  180.1 204.2 186.9 205.0 ;
      RECT  180.1 209.4 186.9 210.2 ;
      RECT  180.1 225.0 186.9 225.8 ;
      RECT  180.1 230.2 186.9 231.0 ;
      RECT  180.1 245.8 186.9 246.6 ;
      RECT  180.1 251.0 186.9 251.8 ;
      RECT  180.1 266.6 186.9 267.4 ;
      RECT  180.1 271.8 186.9 272.6 ;
      RECT  180.1 287.4 186.9 288.2 ;
      RECT  180.1 292.6 186.9 293.4 ;
      RECT  180.1 308.2 186.9 309.0 ;
      RECT  180.1 313.4 186.9 314.2 ;
      RECT  180.1 329.0 186.9 329.8 ;
      RECT  180.1 334.2 186.9 335.0 ;
      RECT  180.1 349.8 186.9 350.6 ;
      RECT  180.1 355.0 186.9 355.8 ;
      RECT  188.9 182.4 189.9 181.6 ;
      RECT  191.3 178.0 192.3 177.2 ;
      RECT  191.5 181.6 192.3 181.2 ;
      RECT  190.3 183.4 191.1 183.2 ;
      RECT  193.3 182.8 194.1 178.6 ;
      RECT  189.1 179.4 190.7 178.6 ;
      RECT  191.5 182.4 192.5 181.6 ;
      RECT  188.9 185.6 189.7 184.8 ;
      RECT  186.5 176.4 194.1 175.6 ;
      RECT  186.5 178.0 187.3 176.4 ;
      RECT  189.1 178.0 190.1 177.2 ;
      RECT  189.1 178.6 189.9 178.0 ;
      RECT  191.5 180.4 192.3 178.0 ;
      RECT  191.1 181.2 192.3 180.4 ;
      RECT  186.5 184.2 194.1 183.4 ;
      RECT  191.7 185.6 192.5 184.8 ;
      RECT  186.5 182.8 187.3 178.6 ;
      RECT  189.1 181.6 189.9 179.4 ;
      RECT  193.3 178.0 194.1 176.4 ;
      RECT  195.7 182.4 196.7 181.6 ;
      RECT  198.1 178.0 199.1 177.2 ;
      RECT  198.3 181.6 199.1 181.2 ;
      RECT  197.1 183.4 197.9 183.2 ;
      RECT  200.1 182.8 200.9 178.6 ;
      RECT  195.9 179.4 197.5 178.6 ;
      RECT  198.3 182.4 199.3 181.6 ;
      RECT  195.7 185.6 196.5 184.8 ;
      RECT  193.3 176.4 200.9 175.6 ;
      RECT  193.3 178.0 194.1 176.4 ;
      RECT  195.9 178.0 196.9 177.2 ;
      RECT  195.9 178.6 196.7 178.0 ;
      RECT  198.3 180.4 199.1 178.0 ;
      RECT  197.9 181.2 199.1 180.4 ;
      RECT  193.3 184.2 200.9 183.4 ;
      RECT  198.5 185.6 199.3 184.8 ;
      RECT  193.3 182.8 194.1 178.6 ;
      RECT  195.9 181.6 196.7 179.4 ;
      RECT  200.1 178.0 200.9 176.4 ;
      RECT  186.9 184.2 200.5 183.4 ;
      RECT  188.9 169.6 189.9 170.4 ;
      RECT  191.3 174.0 192.3 174.8 ;
      RECT  191.5 170.4 192.3 170.8 ;
      RECT  190.3 168.6 191.1 168.8 ;
      RECT  193.3 169.2 194.1 173.4 ;
      RECT  189.1 172.6 190.7 173.4 ;
      RECT  191.5 169.6 192.5 170.4 ;
      RECT  188.9 166.4 189.7 167.2 ;
      RECT  186.5 175.6 194.1 176.4 ;
      RECT  186.5 174.0 187.3 175.6 ;
      RECT  189.1 174.0 190.1 174.8 ;
      RECT  189.1 173.4 189.9 174.0 ;
      RECT  191.5 171.6 192.3 174.0 ;
      RECT  191.1 170.8 192.3 171.6 ;
      RECT  186.5 167.8 194.1 168.6 ;
      RECT  191.7 166.4 192.5 167.2 ;
      RECT  186.5 169.2 187.3 173.4 ;
      RECT  189.1 170.4 189.9 172.6 ;
      RECT  193.3 174.0 194.1 175.6 ;
      RECT  195.7 169.6 196.7 170.4 ;
      RECT  198.1 174.0 199.1 174.8 ;
      RECT  198.3 170.4 199.1 170.8 ;
      RECT  197.1 168.6 197.9 168.8 ;
      RECT  200.1 169.2 200.9 173.4 ;
      RECT  195.9 172.6 197.5 173.4 ;
      RECT  198.3 169.6 199.3 170.4 ;
      RECT  195.7 166.4 196.5 167.2 ;
      RECT  193.3 175.6 200.9 176.4 ;
      RECT  193.3 174.0 194.1 175.6 ;
      RECT  195.9 174.0 196.9 174.8 ;
      RECT  195.9 173.4 196.7 174.0 ;
      RECT  198.3 171.6 199.1 174.0 ;
      RECT  197.9 170.8 199.1 171.6 ;
      RECT  193.3 167.8 200.9 168.6 ;
      RECT  198.5 166.4 199.3 167.2 ;
      RECT  193.3 169.2 194.1 173.4 ;
      RECT  195.9 170.4 196.7 172.6 ;
      RECT  200.1 174.0 200.9 175.6 ;
      RECT  186.9 167.8 200.5 168.6 ;
      RECT  188.9 356.8 189.9 357.6 ;
      RECT  191.3 361.2 192.3 362.0 ;
      RECT  191.5 357.6 192.3 358.0 ;
      RECT  190.3 355.8 191.1 356.0 ;
      RECT  193.3 356.4 194.1 360.6 ;
      RECT  189.1 359.8 190.7 360.6 ;
      RECT  191.5 356.8 192.5 357.6 ;
      RECT  188.9 353.6 189.7 354.4 ;
      RECT  186.5 362.8 194.1 363.6 ;
      RECT  186.5 361.2 187.3 362.8 ;
      RECT  189.1 361.2 190.1 362.0 ;
      RECT  189.1 360.6 189.9 361.2 ;
      RECT  191.5 358.8 192.3 361.2 ;
      RECT  191.1 358.0 192.3 358.8 ;
      RECT  186.5 355.0 194.1 355.8 ;
      RECT  191.7 353.6 192.5 354.4 ;
      RECT  186.5 356.4 187.3 360.6 ;
      RECT  189.1 357.6 189.9 359.8 ;
      RECT  193.3 361.2 194.1 362.8 ;
      RECT  195.7 356.8 196.7 357.6 ;
      RECT  198.1 361.2 199.1 362.0 ;
      RECT  198.3 357.6 199.1 358.0 ;
      RECT  197.1 355.8 197.9 356.0 ;
      RECT  200.1 356.4 200.9 360.6 ;
      RECT  195.9 359.8 197.5 360.6 ;
      RECT  198.3 356.8 199.3 357.6 ;
      RECT  195.7 353.6 196.5 354.4 ;
      RECT  193.3 362.8 200.9 363.6 ;
      RECT  193.3 361.2 194.1 362.8 ;
      RECT  195.9 361.2 196.9 362.0 ;
      RECT  195.9 360.6 196.7 361.2 ;
      RECT  198.3 358.8 199.1 361.2 ;
      RECT  197.9 358.0 199.1 358.8 ;
      RECT  193.3 355.0 200.9 355.8 ;
      RECT  198.5 353.6 199.3 354.4 ;
      RECT  193.3 356.4 194.1 360.6 ;
      RECT  195.9 357.6 196.7 359.8 ;
      RECT  200.1 361.2 200.9 362.8 ;
      RECT  186.9 355.0 200.5 355.8 ;
      RECT  175.3 169.6 176.3 170.4 ;
      RECT  177.7 174.0 178.7 174.8 ;
      RECT  177.9 170.4 178.7 170.8 ;
      RECT  176.7 168.6 177.5 168.8 ;
      RECT  179.7 169.2 180.5 173.4 ;
      RECT  175.5 172.6 177.1 173.4 ;
      RECT  177.9 169.6 178.9 170.4 ;
      RECT  175.3 166.4 176.1 167.2 ;
      RECT  172.9 175.6 180.5 176.4 ;
      RECT  172.9 174.0 173.7 175.6 ;
      RECT  175.5 174.0 176.5 174.8 ;
      RECT  175.5 173.4 176.3 174.0 ;
      RECT  177.9 171.6 178.7 174.0 ;
      RECT  177.5 170.8 178.7 171.6 ;
      RECT  172.9 167.8 180.5 168.6 ;
      RECT  178.1 166.4 178.9 167.2 ;
      RECT  172.9 169.2 173.7 173.4 ;
      RECT  175.5 170.4 176.3 172.6 ;
      RECT  179.7 174.0 180.5 175.6 ;
      RECT  175.3 182.4 176.3 181.6 ;
      RECT  177.7 178.0 178.7 177.2 ;
      RECT  177.9 181.6 178.7 181.2 ;
      RECT  176.7 183.4 177.5 183.2 ;
      RECT  179.7 182.8 180.5 178.6 ;
      RECT  175.5 179.4 177.1 178.6 ;
      RECT  177.9 182.4 178.9 181.6 ;
      RECT  175.3 185.6 176.1 184.8 ;
      RECT  172.9 176.4 180.5 175.6 ;
      RECT  172.9 178.0 173.7 176.4 ;
      RECT  175.5 178.0 176.5 177.2 ;
      RECT  175.5 178.6 176.3 178.0 ;
      RECT  177.9 180.4 178.7 178.0 ;
      RECT  177.5 181.2 178.7 180.4 ;
      RECT  172.9 184.2 180.5 183.4 ;
      RECT  178.1 185.6 178.9 184.8 ;
      RECT  172.9 182.8 173.7 178.6 ;
      RECT  175.5 181.6 176.3 179.4 ;
      RECT  179.7 178.0 180.5 176.4 ;
      RECT  175.3 190.4 176.3 191.2 ;
      RECT  177.7 194.8 178.7 195.6 ;
      RECT  177.9 191.2 178.7 191.6 ;
      RECT  176.7 189.4 177.5 189.6 ;
      RECT  179.7 190.0 180.5 194.2 ;
      RECT  175.5 193.4 177.1 194.2 ;
      RECT  177.9 190.4 178.9 191.2 ;
      RECT  175.3 187.2 176.1 188.0 ;
      RECT  172.9 196.4 180.5 197.2 ;
      RECT  172.9 194.8 173.7 196.4 ;
      RECT  175.5 194.8 176.5 195.6 ;
      RECT  175.5 194.2 176.3 194.8 ;
      RECT  177.9 192.4 178.7 194.8 ;
      RECT  177.5 191.6 178.7 192.4 ;
      RECT  172.9 188.6 180.5 189.4 ;
      RECT  178.1 187.2 178.9 188.0 ;
      RECT  172.9 190.0 173.7 194.2 ;
      RECT  175.5 191.2 176.3 193.4 ;
      RECT  179.7 194.8 180.5 196.4 ;
      RECT  175.3 203.2 176.3 202.4 ;
      RECT  177.7 198.8 178.7 198.0 ;
      RECT  177.9 202.4 178.7 202.0 ;
      RECT  176.7 204.2 177.5 204.0 ;
      RECT  179.7 203.6 180.5 199.4 ;
      RECT  175.5 200.2 177.1 199.4 ;
      RECT  177.9 203.2 178.9 202.4 ;
      RECT  175.3 206.4 176.1 205.6 ;
      RECT  172.9 197.2 180.5 196.4 ;
      RECT  172.9 198.8 173.7 197.2 ;
      RECT  175.5 198.8 176.5 198.0 ;
      RECT  175.5 199.4 176.3 198.8 ;
      RECT  177.9 201.2 178.7 198.8 ;
      RECT  177.5 202.0 178.7 201.2 ;
      RECT  172.9 205.0 180.5 204.2 ;
      RECT  178.1 206.4 178.9 205.6 ;
      RECT  172.9 203.6 173.7 199.4 ;
      RECT  175.5 202.4 176.3 200.2 ;
      RECT  179.7 198.8 180.5 197.2 ;
      RECT  175.3 211.2 176.3 212.0 ;
      RECT  177.7 215.6 178.7 216.4 ;
      RECT  177.9 212.0 178.7 212.4 ;
      RECT  176.7 210.2 177.5 210.4 ;
      RECT  179.7 210.8 180.5 215.0 ;
      RECT  175.5 214.2 177.1 215.0 ;
      RECT  177.9 211.2 178.9 212.0 ;
      RECT  175.3 208.0 176.1 208.8 ;
      RECT  172.9 217.2 180.5 218.0 ;
      RECT  172.9 215.6 173.7 217.2 ;
      RECT  175.5 215.6 176.5 216.4 ;
      RECT  175.5 215.0 176.3 215.6 ;
      RECT  177.9 213.2 178.7 215.6 ;
      RECT  177.5 212.4 178.7 213.2 ;
      RECT  172.9 209.4 180.5 210.2 ;
      RECT  178.1 208.0 178.9 208.8 ;
      RECT  172.9 210.8 173.7 215.0 ;
      RECT  175.5 212.0 176.3 214.2 ;
      RECT  179.7 215.6 180.5 217.2 ;
      RECT  175.3 224.0 176.3 223.2 ;
      RECT  177.7 219.6 178.7 218.8 ;
      RECT  177.9 223.2 178.7 222.8 ;
      RECT  176.7 225.0 177.5 224.8 ;
      RECT  179.7 224.4 180.5 220.2 ;
      RECT  175.5 221.0 177.1 220.2 ;
      RECT  177.9 224.0 178.9 223.2 ;
      RECT  175.3 227.2 176.1 226.4 ;
      RECT  172.9 218.0 180.5 217.2 ;
      RECT  172.9 219.6 173.7 218.0 ;
      RECT  175.5 219.6 176.5 218.8 ;
      RECT  175.5 220.2 176.3 219.6 ;
      RECT  177.9 222.0 178.7 219.6 ;
      RECT  177.5 222.8 178.7 222.0 ;
      RECT  172.9 225.8 180.5 225.0 ;
      RECT  178.1 227.2 178.9 226.4 ;
      RECT  172.9 224.4 173.7 220.2 ;
      RECT  175.5 223.2 176.3 221.0 ;
      RECT  179.7 219.6 180.5 218.0 ;
      RECT  175.3 232.0 176.3 232.8 ;
      RECT  177.7 236.4 178.7 237.2 ;
      RECT  177.9 232.8 178.7 233.2 ;
      RECT  176.7 231.0 177.5 231.2 ;
      RECT  179.7 231.6 180.5 235.8 ;
      RECT  175.5 235.0 177.1 235.8 ;
      RECT  177.9 232.0 178.9 232.8 ;
      RECT  175.3 228.8 176.1 229.6 ;
      RECT  172.9 238.0 180.5 238.8 ;
      RECT  172.9 236.4 173.7 238.0 ;
      RECT  175.5 236.4 176.5 237.2 ;
      RECT  175.5 235.8 176.3 236.4 ;
      RECT  177.9 234.0 178.7 236.4 ;
      RECT  177.5 233.2 178.7 234.0 ;
      RECT  172.9 230.2 180.5 231.0 ;
      RECT  178.1 228.8 178.9 229.6 ;
      RECT  172.9 231.6 173.7 235.8 ;
      RECT  175.5 232.8 176.3 235.0 ;
      RECT  179.7 236.4 180.5 238.0 ;
      RECT  175.3 244.8 176.3 244.0 ;
      RECT  177.7 240.4 178.7 239.6 ;
      RECT  177.9 244.0 178.7 243.6 ;
      RECT  176.7 245.8 177.5 245.6 ;
      RECT  179.7 245.2 180.5 241.0 ;
      RECT  175.5 241.8 177.1 241.0 ;
      RECT  177.9 244.8 178.9 244.0 ;
      RECT  175.3 248.0 176.1 247.2 ;
      RECT  172.9 238.8 180.5 238.0 ;
      RECT  172.9 240.4 173.7 238.8 ;
      RECT  175.5 240.4 176.5 239.6 ;
      RECT  175.5 241.0 176.3 240.4 ;
      RECT  177.9 242.8 178.7 240.4 ;
      RECT  177.5 243.6 178.7 242.8 ;
      RECT  172.9 246.6 180.5 245.8 ;
      RECT  178.1 248.0 178.9 247.2 ;
      RECT  172.9 245.2 173.7 241.0 ;
      RECT  175.5 244.0 176.3 241.8 ;
      RECT  179.7 240.4 180.5 238.8 ;
      RECT  175.3 252.8 176.3 253.6 ;
      RECT  177.7 257.2 178.7 258.0 ;
      RECT  177.9 253.6 178.7 254.0 ;
      RECT  176.7 251.8 177.5 252.0 ;
      RECT  179.7 252.4 180.5 256.6 ;
      RECT  175.5 255.8 177.1 256.6 ;
      RECT  177.9 252.8 178.9 253.6 ;
      RECT  175.3 249.6 176.1 250.4 ;
      RECT  172.9 258.8 180.5 259.6 ;
      RECT  172.9 257.2 173.7 258.8 ;
      RECT  175.5 257.2 176.5 258.0 ;
      RECT  175.5 256.6 176.3 257.2 ;
      RECT  177.9 254.8 178.7 257.2 ;
      RECT  177.5 254.0 178.7 254.8 ;
      RECT  172.9 251.0 180.5 251.8 ;
      RECT  178.1 249.6 178.9 250.4 ;
      RECT  172.9 252.4 173.7 256.6 ;
      RECT  175.5 253.6 176.3 255.8 ;
      RECT  179.7 257.2 180.5 258.8 ;
      RECT  175.3 265.6 176.3 264.8 ;
      RECT  177.7 261.2 178.7 260.4 ;
      RECT  177.9 264.8 178.7 264.4 ;
      RECT  176.7 266.6 177.5 266.4 ;
      RECT  179.7 266.0 180.5 261.8 ;
      RECT  175.5 262.6 177.1 261.8 ;
      RECT  177.9 265.6 178.9 264.8 ;
      RECT  175.3 268.8 176.1 268.0 ;
      RECT  172.9 259.6 180.5 258.8 ;
      RECT  172.9 261.2 173.7 259.6 ;
      RECT  175.5 261.2 176.5 260.4 ;
      RECT  175.5 261.8 176.3 261.2 ;
      RECT  177.9 263.6 178.7 261.2 ;
      RECT  177.5 264.4 178.7 263.6 ;
      RECT  172.9 267.4 180.5 266.6 ;
      RECT  178.1 268.8 178.9 268.0 ;
      RECT  172.9 266.0 173.7 261.8 ;
      RECT  175.5 264.8 176.3 262.6 ;
      RECT  179.7 261.2 180.5 259.6 ;
      RECT  175.3 273.6 176.3 274.4 ;
      RECT  177.7 278.0 178.7 278.8 ;
      RECT  177.9 274.4 178.7 274.8 ;
      RECT  176.7 272.6 177.5 272.8 ;
      RECT  179.7 273.2 180.5 277.4 ;
      RECT  175.5 276.6 177.1 277.4 ;
      RECT  177.9 273.6 178.9 274.4 ;
      RECT  175.3 270.4 176.1 271.2 ;
      RECT  172.9 279.6 180.5 280.4 ;
      RECT  172.9 278.0 173.7 279.6 ;
      RECT  175.5 278.0 176.5 278.8 ;
      RECT  175.5 277.4 176.3 278.0 ;
      RECT  177.9 275.6 178.7 278.0 ;
      RECT  177.5 274.8 178.7 275.6 ;
      RECT  172.9 271.8 180.5 272.6 ;
      RECT  178.1 270.4 178.9 271.2 ;
      RECT  172.9 273.2 173.7 277.4 ;
      RECT  175.5 274.4 176.3 276.6 ;
      RECT  179.7 278.0 180.5 279.6 ;
      RECT  175.3 286.4 176.3 285.6 ;
      RECT  177.7 282.0 178.7 281.2 ;
      RECT  177.9 285.6 178.7 285.2 ;
      RECT  176.7 287.4 177.5 287.2 ;
      RECT  179.7 286.8 180.5 282.6 ;
      RECT  175.5 283.4 177.1 282.6 ;
      RECT  177.9 286.4 178.9 285.6 ;
      RECT  175.3 289.6 176.1 288.8 ;
      RECT  172.9 280.4 180.5 279.6 ;
      RECT  172.9 282.0 173.7 280.4 ;
      RECT  175.5 282.0 176.5 281.2 ;
      RECT  175.5 282.6 176.3 282.0 ;
      RECT  177.9 284.4 178.7 282.0 ;
      RECT  177.5 285.2 178.7 284.4 ;
      RECT  172.9 288.2 180.5 287.4 ;
      RECT  178.1 289.6 178.9 288.8 ;
      RECT  172.9 286.8 173.7 282.6 ;
      RECT  175.5 285.6 176.3 283.4 ;
      RECT  179.7 282.0 180.5 280.4 ;
      RECT  175.3 294.4 176.3 295.2 ;
      RECT  177.7 298.8 178.7 299.6 ;
      RECT  177.9 295.2 178.7 295.6 ;
      RECT  176.7 293.4 177.5 293.6 ;
      RECT  179.7 294.0 180.5 298.2 ;
      RECT  175.5 297.4 177.1 298.2 ;
      RECT  177.9 294.4 178.9 295.2 ;
      RECT  175.3 291.2 176.1 292.0 ;
      RECT  172.9 300.4 180.5 301.2 ;
      RECT  172.9 298.8 173.7 300.4 ;
      RECT  175.5 298.8 176.5 299.6 ;
      RECT  175.5 298.2 176.3 298.8 ;
      RECT  177.9 296.4 178.7 298.8 ;
      RECT  177.5 295.6 178.7 296.4 ;
      RECT  172.9 292.6 180.5 293.4 ;
      RECT  178.1 291.2 178.9 292.0 ;
      RECT  172.9 294.0 173.7 298.2 ;
      RECT  175.5 295.2 176.3 297.4 ;
      RECT  179.7 298.8 180.5 300.4 ;
      RECT  175.3 307.2 176.3 306.4 ;
      RECT  177.7 302.8 178.7 302.0 ;
      RECT  177.9 306.4 178.7 306.0 ;
      RECT  176.7 308.2 177.5 308.0 ;
      RECT  179.7 307.6 180.5 303.4 ;
      RECT  175.5 304.2 177.1 303.4 ;
      RECT  177.9 307.2 178.9 306.4 ;
      RECT  175.3 310.4 176.1 309.6 ;
      RECT  172.9 301.2 180.5 300.4 ;
      RECT  172.9 302.8 173.7 301.2 ;
      RECT  175.5 302.8 176.5 302.0 ;
      RECT  175.5 303.4 176.3 302.8 ;
      RECT  177.9 305.2 178.7 302.8 ;
      RECT  177.5 306.0 178.7 305.2 ;
      RECT  172.9 309.0 180.5 308.2 ;
      RECT  178.1 310.4 178.9 309.6 ;
      RECT  172.9 307.6 173.7 303.4 ;
      RECT  175.5 306.4 176.3 304.2 ;
      RECT  179.7 302.8 180.5 301.2 ;
      RECT  175.3 315.2 176.3 316.0 ;
      RECT  177.7 319.6 178.7 320.4 ;
      RECT  177.9 316.0 178.7 316.4 ;
      RECT  176.7 314.2 177.5 314.4 ;
      RECT  179.7 314.8 180.5 319.0 ;
      RECT  175.5 318.2 177.1 319.0 ;
      RECT  177.9 315.2 178.9 316.0 ;
      RECT  175.3 312.0 176.1 312.8 ;
      RECT  172.9 321.2 180.5 322.0 ;
      RECT  172.9 319.6 173.7 321.2 ;
      RECT  175.5 319.6 176.5 320.4 ;
      RECT  175.5 319.0 176.3 319.6 ;
      RECT  177.9 317.2 178.7 319.6 ;
      RECT  177.5 316.4 178.7 317.2 ;
      RECT  172.9 313.4 180.5 314.2 ;
      RECT  178.1 312.0 178.9 312.8 ;
      RECT  172.9 314.8 173.7 319.0 ;
      RECT  175.5 316.0 176.3 318.2 ;
      RECT  179.7 319.6 180.5 321.2 ;
      RECT  175.3 328.0 176.3 327.2 ;
      RECT  177.7 323.6 178.7 322.8 ;
      RECT  177.9 327.2 178.7 326.8 ;
      RECT  176.7 329.0 177.5 328.8 ;
      RECT  179.7 328.4 180.5 324.2 ;
      RECT  175.5 325.0 177.1 324.2 ;
      RECT  177.9 328.0 178.9 327.2 ;
      RECT  175.3 331.2 176.1 330.4 ;
      RECT  172.9 322.0 180.5 321.2 ;
      RECT  172.9 323.6 173.7 322.0 ;
      RECT  175.5 323.6 176.5 322.8 ;
      RECT  175.5 324.2 176.3 323.6 ;
      RECT  177.9 326.0 178.7 323.6 ;
      RECT  177.5 326.8 178.7 326.0 ;
      RECT  172.9 329.8 180.5 329.0 ;
      RECT  178.1 331.2 178.9 330.4 ;
      RECT  172.9 328.4 173.7 324.2 ;
      RECT  175.5 327.2 176.3 325.0 ;
      RECT  179.7 323.6 180.5 322.0 ;
      RECT  175.3 336.0 176.3 336.8 ;
      RECT  177.7 340.4 178.7 341.2 ;
      RECT  177.9 336.8 178.7 337.2 ;
      RECT  176.7 335.0 177.5 335.2 ;
      RECT  179.7 335.6 180.5 339.8 ;
      RECT  175.5 339.0 177.1 339.8 ;
      RECT  177.9 336.0 178.9 336.8 ;
      RECT  175.3 332.8 176.1 333.6 ;
      RECT  172.9 342.0 180.5 342.8 ;
      RECT  172.9 340.4 173.7 342.0 ;
      RECT  175.5 340.4 176.5 341.2 ;
      RECT  175.5 339.8 176.3 340.4 ;
      RECT  177.9 338.0 178.7 340.4 ;
      RECT  177.5 337.2 178.7 338.0 ;
      RECT  172.9 334.2 180.5 335.0 ;
      RECT  178.1 332.8 178.9 333.6 ;
      RECT  172.9 335.6 173.7 339.8 ;
      RECT  175.5 336.8 176.3 339.0 ;
      RECT  179.7 340.4 180.5 342.0 ;
      RECT  175.3 348.8 176.3 348.0 ;
      RECT  177.7 344.4 178.7 343.6 ;
      RECT  177.9 348.0 178.7 347.6 ;
      RECT  176.7 349.8 177.5 349.6 ;
      RECT  179.7 349.2 180.5 345.0 ;
      RECT  175.5 345.8 177.1 345.0 ;
      RECT  177.9 348.8 178.9 348.0 ;
      RECT  175.3 352.0 176.1 351.2 ;
      RECT  172.9 342.8 180.5 342.0 ;
      RECT  172.9 344.4 173.7 342.8 ;
      RECT  175.5 344.4 176.5 343.6 ;
      RECT  175.5 345.0 176.3 344.4 ;
      RECT  177.9 346.8 178.7 344.4 ;
      RECT  177.5 347.6 178.7 346.8 ;
      RECT  172.9 350.6 180.5 349.8 ;
      RECT  178.1 352.0 178.9 351.2 ;
      RECT  172.9 349.2 173.7 345.0 ;
      RECT  175.5 348.0 176.3 345.8 ;
      RECT  179.7 344.4 180.5 342.8 ;
      RECT  175.3 356.8 176.3 357.6 ;
      RECT  177.7 361.2 178.7 362.0 ;
      RECT  177.9 357.6 178.7 358.0 ;
      RECT  176.7 355.8 177.5 356.0 ;
      RECT  179.7 356.4 180.5 360.6 ;
      RECT  175.5 359.8 177.1 360.6 ;
      RECT  177.9 356.8 178.9 357.6 ;
      RECT  175.3 353.6 176.1 354.4 ;
      RECT  172.9 362.8 180.5 363.6 ;
      RECT  172.9 361.2 173.7 362.8 ;
      RECT  175.5 361.2 176.5 362.0 ;
      RECT  175.5 360.6 176.3 361.2 ;
      RECT  177.9 358.8 178.7 361.2 ;
      RECT  177.5 358.0 178.7 358.8 ;
      RECT  172.9 355.0 180.5 355.8 ;
      RECT  178.1 353.6 178.9 354.4 ;
      RECT  172.9 356.4 173.7 360.6 ;
      RECT  175.5 357.6 176.3 359.8 ;
      RECT  179.7 361.2 180.5 362.8 ;
      RECT  173.3 167.8 180.1 168.6 ;
      RECT  173.3 183.4 180.1 184.2 ;
      RECT  173.3 188.6 180.1 189.4 ;
      RECT  173.3 204.2 180.1 205.0 ;
      RECT  173.3 209.4 180.1 210.2 ;
      RECT  173.3 225.0 180.1 225.8 ;
      RECT  173.3 230.2 180.1 231.0 ;
      RECT  173.3 245.8 180.1 246.6 ;
      RECT  173.3 251.0 180.1 251.8 ;
      RECT  173.3 266.6 180.1 267.4 ;
      RECT  173.3 271.8 180.1 272.6 ;
      RECT  173.3 287.4 180.1 288.2 ;
      RECT  173.3 292.6 180.1 293.4 ;
      RECT  173.3 308.2 180.1 309.0 ;
      RECT  173.3 313.4 180.1 314.2 ;
      RECT  173.3 329.0 180.1 329.8 ;
      RECT  173.3 334.2 180.1 335.0 ;
      RECT  173.3 349.8 180.1 350.6 ;
      RECT  173.3 355.0 180.1 355.8 ;
      RECT  202.5 169.6 203.5 170.4 ;
      RECT  204.9 174.0 205.9 174.8 ;
      RECT  205.1 170.4 205.9 170.8 ;
      RECT  203.9 168.6 204.7 168.8 ;
      RECT  206.9 169.2 207.7 173.4 ;
      RECT  202.7 172.6 204.3 173.4 ;
      RECT  205.1 169.6 206.1 170.4 ;
      RECT  202.5 166.4 203.3 167.2 ;
      RECT  200.1 175.6 207.7 176.4 ;
      RECT  200.1 174.0 200.9 175.6 ;
      RECT  202.7 174.0 203.7 174.8 ;
      RECT  202.7 173.4 203.5 174.0 ;
      RECT  205.1 171.6 205.9 174.0 ;
      RECT  204.7 170.8 205.9 171.6 ;
      RECT  200.1 167.8 207.7 168.6 ;
      RECT  205.3 166.4 206.1 167.2 ;
      RECT  200.1 169.2 200.9 173.4 ;
      RECT  202.7 170.4 203.5 172.6 ;
      RECT  206.9 174.0 207.7 175.6 ;
      RECT  202.5 182.4 203.5 181.6 ;
      RECT  204.9 178.0 205.9 177.2 ;
      RECT  205.1 181.6 205.9 181.2 ;
      RECT  203.9 183.4 204.7 183.2 ;
      RECT  206.9 182.8 207.7 178.6 ;
      RECT  202.7 179.4 204.3 178.6 ;
      RECT  205.1 182.4 206.1 181.6 ;
      RECT  202.5 185.6 203.3 184.8 ;
      RECT  200.1 176.4 207.7 175.6 ;
      RECT  200.1 178.0 200.9 176.4 ;
      RECT  202.7 178.0 203.7 177.2 ;
      RECT  202.7 178.6 203.5 178.0 ;
      RECT  205.1 180.4 205.9 178.0 ;
      RECT  204.7 181.2 205.9 180.4 ;
      RECT  200.1 184.2 207.7 183.4 ;
      RECT  205.3 185.6 206.1 184.8 ;
      RECT  200.1 182.8 200.9 178.6 ;
      RECT  202.7 181.6 203.5 179.4 ;
      RECT  206.9 178.0 207.7 176.4 ;
      RECT  202.5 190.4 203.5 191.2 ;
      RECT  204.9 194.8 205.9 195.6 ;
      RECT  205.1 191.2 205.9 191.6 ;
      RECT  203.9 189.4 204.7 189.6 ;
      RECT  206.9 190.0 207.7 194.2 ;
      RECT  202.7 193.4 204.3 194.2 ;
      RECT  205.1 190.4 206.1 191.2 ;
      RECT  202.5 187.2 203.3 188.0 ;
      RECT  200.1 196.4 207.7 197.2 ;
      RECT  200.1 194.8 200.9 196.4 ;
      RECT  202.7 194.8 203.7 195.6 ;
      RECT  202.7 194.2 203.5 194.8 ;
      RECT  205.1 192.4 205.9 194.8 ;
      RECT  204.7 191.6 205.9 192.4 ;
      RECT  200.1 188.6 207.7 189.4 ;
      RECT  205.3 187.2 206.1 188.0 ;
      RECT  200.1 190.0 200.9 194.2 ;
      RECT  202.7 191.2 203.5 193.4 ;
      RECT  206.9 194.8 207.7 196.4 ;
      RECT  202.5 203.2 203.5 202.4 ;
      RECT  204.9 198.8 205.9 198.0 ;
      RECT  205.1 202.4 205.9 202.0 ;
      RECT  203.9 204.2 204.7 204.0 ;
      RECT  206.9 203.6 207.7 199.4 ;
      RECT  202.7 200.2 204.3 199.4 ;
      RECT  205.1 203.2 206.1 202.4 ;
      RECT  202.5 206.4 203.3 205.6 ;
      RECT  200.1 197.2 207.7 196.4 ;
      RECT  200.1 198.8 200.9 197.2 ;
      RECT  202.7 198.8 203.7 198.0 ;
      RECT  202.7 199.4 203.5 198.8 ;
      RECT  205.1 201.2 205.9 198.8 ;
      RECT  204.7 202.0 205.9 201.2 ;
      RECT  200.1 205.0 207.7 204.2 ;
      RECT  205.3 206.4 206.1 205.6 ;
      RECT  200.1 203.6 200.9 199.4 ;
      RECT  202.7 202.4 203.5 200.2 ;
      RECT  206.9 198.8 207.7 197.2 ;
      RECT  202.5 211.2 203.5 212.0 ;
      RECT  204.9 215.6 205.9 216.4 ;
      RECT  205.1 212.0 205.9 212.4 ;
      RECT  203.9 210.2 204.7 210.4 ;
      RECT  206.9 210.8 207.7 215.0 ;
      RECT  202.7 214.2 204.3 215.0 ;
      RECT  205.1 211.2 206.1 212.0 ;
      RECT  202.5 208.0 203.3 208.8 ;
      RECT  200.1 217.2 207.7 218.0 ;
      RECT  200.1 215.6 200.9 217.2 ;
      RECT  202.7 215.6 203.7 216.4 ;
      RECT  202.7 215.0 203.5 215.6 ;
      RECT  205.1 213.2 205.9 215.6 ;
      RECT  204.7 212.4 205.9 213.2 ;
      RECT  200.1 209.4 207.7 210.2 ;
      RECT  205.3 208.0 206.1 208.8 ;
      RECT  200.1 210.8 200.9 215.0 ;
      RECT  202.7 212.0 203.5 214.2 ;
      RECT  206.9 215.6 207.7 217.2 ;
      RECT  202.5 224.0 203.5 223.2 ;
      RECT  204.9 219.6 205.9 218.8 ;
      RECT  205.1 223.2 205.9 222.8 ;
      RECT  203.9 225.0 204.7 224.8 ;
      RECT  206.9 224.4 207.7 220.2 ;
      RECT  202.7 221.0 204.3 220.2 ;
      RECT  205.1 224.0 206.1 223.2 ;
      RECT  202.5 227.2 203.3 226.4 ;
      RECT  200.1 218.0 207.7 217.2 ;
      RECT  200.1 219.6 200.9 218.0 ;
      RECT  202.7 219.6 203.7 218.8 ;
      RECT  202.7 220.2 203.5 219.6 ;
      RECT  205.1 222.0 205.9 219.6 ;
      RECT  204.7 222.8 205.9 222.0 ;
      RECT  200.1 225.8 207.7 225.0 ;
      RECT  205.3 227.2 206.1 226.4 ;
      RECT  200.1 224.4 200.9 220.2 ;
      RECT  202.7 223.2 203.5 221.0 ;
      RECT  206.9 219.6 207.7 218.0 ;
      RECT  202.5 232.0 203.5 232.8 ;
      RECT  204.9 236.4 205.9 237.2 ;
      RECT  205.1 232.8 205.9 233.2 ;
      RECT  203.9 231.0 204.7 231.2 ;
      RECT  206.9 231.6 207.7 235.8 ;
      RECT  202.7 235.0 204.3 235.8 ;
      RECT  205.1 232.0 206.1 232.8 ;
      RECT  202.5 228.8 203.3 229.6 ;
      RECT  200.1 238.0 207.7 238.8 ;
      RECT  200.1 236.4 200.9 238.0 ;
      RECT  202.7 236.4 203.7 237.2 ;
      RECT  202.7 235.8 203.5 236.4 ;
      RECT  205.1 234.0 205.9 236.4 ;
      RECT  204.7 233.2 205.9 234.0 ;
      RECT  200.1 230.2 207.7 231.0 ;
      RECT  205.3 228.8 206.1 229.6 ;
      RECT  200.1 231.6 200.9 235.8 ;
      RECT  202.7 232.8 203.5 235.0 ;
      RECT  206.9 236.4 207.7 238.0 ;
      RECT  202.5 244.8 203.5 244.0 ;
      RECT  204.9 240.4 205.9 239.6 ;
      RECT  205.1 244.0 205.9 243.6 ;
      RECT  203.9 245.8 204.7 245.6 ;
      RECT  206.9 245.2 207.7 241.0 ;
      RECT  202.7 241.8 204.3 241.0 ;
      RECT  205.1 244.8 206.1 244.0 ;
      RECT  202.5 248.0 203.3 247.2 ;
      RECT  200.1 238.8 207.7 238.0 ;
      RECT  200.1 240.4 200.9 238.8 ;
      RECT  202.7 240.4 203.7 239.6 ;
      RECT  202.7 241.0 203.5 240.4 ;
      RECT  205.1 242.8 205.9 240.4 ;
      RECT  204.7 243.6 205.9 242.8 ;
      RECT  200.1 246.6 207.7 245.8 ;
      RECT  205.3 248.0 206.1 247.2 ;
      RECT  200.1 245.2 200.9 241.0 ;
      RECT  202.7 244.0 203.5 241.8 ;
      RECT  206.9 240.4 207.7 238.8 ;
      RECT  202.5 252.8 203.5 253.6 ;
      RECT  204.9 257.2 205.9 258.0 ;
      RECT  205.1 253.6 205.9 254.0 ;
      RECT  203.9 251.8 204.7 252.0 ;
      RECT  206.9 252.4 207.7 256.6 ;
      RECT  202.7 255.8 204.3 256.6 ;
      RECT  205.1 252.8 206.1 253.6 ;
      RECT  202.5 249.6 203.3 250.4 ;
      RECT  200.1 258.8 207.7 259.6 ;
      RECT  200.1 257.2 200.9 258.8 ;
      RECT  202.7 257.2 203.7 258.0 ;
      RECT  202.7 256.6 203.5 257.2 ;
      RECT  205.1 254.8 205.9 257.2 ;
      RECT  204.7 254.0 205.9 254.8 ;
      RECT  200.1 251.0 207.7 251.8 ;
      RECT  205.3 249.6 206.1 250.4 ;
      RECT  200.1 252.4 200.9 256.6 ;
      RECT  202.7 253.6 203.5 255.8 ;
      RECT  206.9 257.2 207.7 258.8 ;
      RECT  202.5 265.6 203.5 264.8 ;
      RECT  204.9 261.2 205.9 260.4 ;
      RECT  205.1 264.8 205.9 264.4 ;
      RECT  203.9 266.6 204.7 266.4 ;
      RECT  206.9 266.0 207.7 261.8 ;
      RECT  202.7 262.6 204.3 261.8 ;
      RECT  205.1 265.6 206.1 264.8 ;
      RECT  202.5 268.8 203.3 268.0 ;
      RECT  200.1 259.6 207.7 258.8 ;
      RECT  200.1 261.2 200.9 259.6 ;
      RECT  202.7 261.2 203.7 260.4 ;
      RECT  202.7 261.8 203.5 261.2 ;
      RECT  205.1 263.6 205.9 261.2 ;
      RECT  204.7 264.4 205.9 263.6 ;
      RECT  200.1 267.4 207.7 266.6 ;
      RECT  205.3 268.8 206.1 268.0 ;
      RECT  200.1 266.0 200.9 261.8 ;
      RECT  202.7 264.8 203.5 262.6 ;
      RECT  206.9 261.2 207.7 259.6 ;
      RECT  202.5 273.6 203.5 274.4 ;
      RECT  204.9 278.0 205.9 278.8 ;
      RECT  205.1 274.4 205.9 274.8 ;
      RECT  203.9 272.6 204.7 272.8 ;
      RECT  206.9 273.2 207.7 277.4 ;
      RECT  202.7 276.6 204.3 277.4 ;
      RECT  205.1 273.6 206.1 274.4 ;
      RECT  202.5 270.4 203.3 271.2 ;
      RECT  200.1 279.6 207.7 280.4 ;
      RECT  200.1 278.0 200.9 279.6 ;
      RECT  202.7 278.0 203.7 278.8 ;
      RECT  202.7 277.4 203.5 278.0 ;
      RECT  205.1 275.6 205.9 278.0 ;
      RECT  204.7 274.8 205.9 275.6 ;
      RECT  200.1 271.8 207.7 272.6 ;
      RECT  205.3 270.4 206.1 271.2 ;
      RECT  200.1 273.2 200.9 277.4 ;
      RECT  202.7 274.4 203.5 276.6 ;
      RECT  206.9 278.0 207.7 279.6 ;
      RECT  202.5 286.4 203.5 285.6 ;
      RECT  204.9 282.0 205.9 281.2 ;
      RECT  205.1 285.6 205.9 285.2 ;
      RECT  203.9 287.4 204.7 287.2 ;
      RECT  206.9 286.8 207.7 282.6 ;
      RECT  202.7 283.4 204.3 282.6 ;
      RECT  205.1 286.4 206.1 285.6 ;
      RECT  202.5 289.6 203.3 288.8 ;
      RECT  200.1 280.4 207.7 279.6 ;
      RECT  200.1 282.0 200.9 280.4 ;
      RECT  202.7 282.0 203.7 281.2 ;
      RECT  202.7 282.6 203.5 282.0 ;
      RECT  205.1 284.4 205.9 282.0 ;
      RECT  204.7 285.2 205.9 284.4 ;
      RECT  200.1 288.2 207.7 287.4 ;
      RECT  205.3 289.6 206.1 288.8 ;
      RECT  200.1 286.8 200.9 282.6 ;
      RECT  202.7 285.6 203.5 283.4 ;
      RECT  206.9 282.0 207.7 280.4 ;
      RECT  202.5 294.4 203.5 295.2 ;
      RECT  204.9 298.8 205.9 299.6 ;
      RECT  205.1 295.2 205.9 295.6 ;
      RECT  203.9 293.4 204.7 293.6 ;
      RECT  206.9 294.0 207.7 298.2 ;
      RECT  202.7 297.4 204.3 298.2 ;
      RECT  205.1 294.4 206.1 295.2 ;
      RECT  202.5 291.2 203.3 292.0 ;
      RECT  200.1 300.4 207.7 301.2 ;
      RECT  200.1 298.8 200.9 300.4 ;
      RECT  202.7 298.8 203.7 299.6 ;
      RECT  202.7 298.2 203.5 298.8 ;
      RECT  205.1 296.4 205.9 298.8 ;
      RECT  204.7 295.6 205.9 296.4 ;
      RECT  200.1 292.6 207.7 293.4 ;
      RECT  205.3 291.2 206.1 292.0 ;
      RECT  200.1 294.0 200.9 298.2 ;
      RECT  202.7 295.2 203.5 297.4 ;
      RECT  206.9 298.8 207.7 300.4 ;
      RECT  202.5 307.2 203.5 306.4 ;
      RECT  204.9 302.8 205.9 302.0 ;
      RECT  205.1 306.4 205.9 306.0 ;
      RECT  203.9 308.2 204.7 308.0 ;
      RECT  206.9 307.6 207.7 303.4 ;
      RECT  202.7 304.2 204.3 303.4 ;
      RECT  205.1 307.2 206.1 306.4 ;
      RECT  202.5 310.4 203.3 309.6 ;
      RECT  200.1 301.2 207.7 300.4 ;
      RECT  200.1 302.8 200.9 301.2 ;
      RECT  202.7 302.8 203.7 302.0 ;
      RECT  202.7 303.4 203.5 302.8 ;
      RECT  205.1 305.2 205.9 302.8 ;
      RECT  204.7 306.0 205.9 305.2 ;
      RECT  200.1 309.0 207.7 308.2 ;
      RECT  205.3 310.4 206.1 309.6 ;
      RECT  200.1 307.6 200.9 303.4 ;
      RECT  202.7 306.4 203.5 304.2 ;
      RECT  206.9 302.8 207.7 301.2 ;
      RECT  202.5 315.2 203.5 316.0 ;
      RECT  204.9 319.6 205.9 320.4 ;
      RECT  205.1 316.0 205.9 316.4 ;
      RECT  203.9 314.2 204.7 314.4 ;
      RECT  206.9 314.8 207.7 319.0 ;
      RECT  202.7 318.2 204.3 319.0 ;
      RECT  205.1 315.2 206.1 316.0 ;
      RECT  202.5 312.0 203.3 312.8 ;
      RECT  200.1 321.2 207.7 322.0 ;
      RECT  200.1 319.6 200.9 321.2 ;
      RECT  202.7 319.6 203.7 320.4 ;
      RECT  202.7 319.0 203.5 319.6 ;
      RECT  205.1 317.2 205.9 319.6 ;
      RECT  204.7 316.4 205.9 317.2 ;
      RECT  200.1 313.4 207.7 314.2 ;
      RECT  205.3 312.0 206.1 312.8 ;
      RECT  200.1 314.8 200.9 319.0 ;
      RECT  202.7 316.0 203.5 318.2 ;
      RECT  206.9 319.6 207.7 321.2 ;
      RECT  202.5 328.0 203.5 327.2 ;
      RECT  204.9 323.6 205.9 322.8 ;
      RECT  205.1 327.2 205.9 326.8 ;
      RECT  203.9 329.0 204.7 328.8 ;
      RECT  206.9 328.4 207.7 324.2 ;
      RECT  202.7 325.0 204.3 324.2 ;
      RECT  205.1 328.0 206.1 327.2 ;
      RECT  202.5 331.2 203.3 330.4 ;
      RECT  200.1 322.0 207.7 321.2 ;
      RECT  200.1 323.6 200.9 322.0 ;
      RECT  202.7 323.6 203.7 322.8 ;
      RECT  202.7 324.2 203.5 323.6 ;
      RECT  205.1 326.0 205.9 323.6 ;
      RECT  204.7 326.8 205.9 326.0 ;
      RECT  200.1 329.8 207.7 329.0 ;
      RECT  205.3 331.2 206.1 330.4 ;
      RECT  200.1 328.4 200.9 324.2 ;
      RECT  202.7 327.2 203.5 325.0 ;
      RECT  206.9 323.6 207.7 322.0 ;
      RECT  202.5 336.0 203.5 336.8 ;
      RECT  204.9 340.4 205.9 341.2 ;
      RECT  205.1 336.8 205.9 337.2 ;
      RECT  203.9 335.0 204.7 335.2 ;
      RECT  206.9 335.6 207.7 339.8 ;
      RECT  202.7 339.0 204.3 339.8 ;
      RECT  205.1 336.0 206.1 336.8 ;
      RECT  202.5 332.8 203.3 333.6 ;
      RECT  200.1 342.0 207.7 342.8 ;
      RECT  200.1 340.4 200.9 342.0 ;
      RECT  202.7 340.4 203.7 341.2 ;
      RECT  202.7 339.8 203.5 340.4 ;
      RECT  205.1 338.0 205.9 340.4 ;
      RECT  204.7 337.2 205.9 338.0 ;
      RECT  200.1 334.2 207.7 335.0 ;
      RECT  205.3 332.8 206.1 333.6 ;
      RECT  200.1 335.6 200.9 339.8 ;
      RECT  202.7 336.8 203.5 339.0 ;
      RECT  206.9 340.4 207.7 342.0 ;
      RECT  202.5 348.8 203.5 348.0 ;
      RECT  204.9 344.4 205.9 343.6 ;
      RECT  205.1 348.0 205.9 347.6 ;
      RECT  203.9 349.8 204.7 349.6 ;
      RECT  206.9 349.2 207.7 345.0 ;
      RECT  202.7 345.8 204.3 345.0 ;
      RECT  205.1 348.8 206.1 348.0 ;
      RECT  202.5 352.0 203.3 351.2 ;
      RECT  200.1 342.8 207.7 342.0 ;
      RECT  200.1 344.4 200.9 342.8 ;
      RECT  202.7 344.4 203.7 343.6 ;
      RECT  202.7 345.0 203.5 344.4 ;
      RECT  205.1 346.8 205.9 344.4 ;
      RECT  204.7 347.6 205.9 346.8 ;
      RECT  200.1 350.6 207.7 349.8 ;
      RECT  205.3 352.0 206.1 351.2 ;
      RECT  200.1 349.2 200.9 345.0 ;
      RECT  202.7 348.0 203.5 345.8 ;
      RECT  206.9 344.4 207.7 342.8 ;
      RECT  202.5 356.8 203.5 357.6 ;
      RECT  204.9 361.2 205.9 362.0 ;
      RECT  205.1 357.6 205.9 358.0 ;
      RECT  203.9 355.8 204.7 356.0 ;
      RECT  206.9 356.4 207.7 360.6 ;
      RECT  202.7 359.8 204.3 360.6 ;
      RECT  205.1 356.8 206.1 357.6 ;
      RECT  202.5 353.6 203.3 354.4 ;
      RECT  200.1 362.8 207.7 363.6 ;
      RECT  200.1 361.2 200.9 362.8 ;
      RECT  202.7 361.2 203.7 362.0 ;
      RECT  202.7 360.6 203.5 361.2 ;
      RECT  205.1 358.8 205.9 361.2 ;
      RECT  204.7 358.0 205.9 358.8 ;
      RECT  200.1 355.0 207.7 355.8 ;
      RECT  205.3 353.6 206.1 354.4 ;
      RECT  200.1 356.4 200.9 360.6 ;
      RECT  202.7 357.6 203.5 359.8 ;
      RECT  206.9 361.2 207.7 362.8 ;
      RECT  200.5 167.8 207.3 168.6 ;
      RECT  200.5 183.4 207.3 184.2 ;
      RECT  200.5 188.6 207.3 189.4 ;
      RECT  200.5 204.2 207.3 205.0 ;
      RECT  200.5 209.4 207.3 210.2 ;
      RECT  200.5 225.0 207.3 225.8 ;
      RECT  200.5 230.2 207.3 231.0 ;
      RECT  200.5 245.8 207.3 246.6 ;
      RECT  200.5 251.0 207.3 251.8 ;
      RECT  200.5 266.6 207.3 267.4 ;
      RECT  200.5 271.8 207.3 272.6 ;
      RECT  200.5 287.4 207.3 288.2 ;
      RECT  200.5 292.6 207.3 293.4 ;
      RECT  200.5 308.2 207.3 309.0 ;
      RECT  200.5 313.4 207.3 314.2 ;
      RECT  200.5 329.0 207.3 329.8 ;
      RECT  200.5 334.2 207.3 335.0 ;
      RECT  200.5 349.8 207.3 350.6 ;
      RECT  200.5 355.0 207.3 355.8 ;
      RECT  173.3 167.8 207.3 168.6 ;
      RECT  173.3 183.4 207.3 184.2 ;
      RECT  173.3 188.6 207.3 189.4 ;
      RECT  173.3 204.2 207.3 205.0 ;
      RECT  173.3 209.4 207.3 210.2 ;
      RECT  173.3 225.0 207.3 225.8 ;
      RECT  173.3 230.2 207.3 231.0 ;
      RECT  173.3 245.8 207.3 246.6 ;
      RECT  173.3 251.0 207.3 251.8 ;
      RECT  173.3 266.6 207.3 267.4 ;
      RECT  173.3 271.8 207.3 272.6 ;
      RECT  173.3 287.4 207.3 288.2 ;
      RECT  173.3 292.6 207.3 293.4 ;
      RECT  173.3 308.2 207.3 309.0 ;
      RECT  173.3 313.4 207.3 314.2 ;
      RECT  173.3 329.0 207.3 329.8 ;
      RECT  173.3 334.2 207.3 335.0 ;
      RECT  173.3 349.8 207.3 350.6 ;
      RECT  173.3 355.0 207.3 355.8 ;
      RECT  183.6 152.4 184.4 153.2 ;
      RECT  181.6 152.4 182.4 153.2 ;
      RECT  183.6 156.8 184.4 157.6 ;
      RECT  181.6 156.8 182.4 157.6 ;
      RECT  185.6 156.8 186.4 157.6 ;
      RECT  183.6 156.8 184.4 157.6 ;
      RECT  180.1 150.3 186.9 150.9 ;
      RECT  190.4 152.4 191.2 153.2 ;
      RECT  188.4 152.4 189.2 153.2 ;
      RECT  190.4 156.8 191.2 157.6 ;
      RECT  188.4 156.8 189.2 157.6 ;
      RECT  192.4 156.8 193.2 157.6 ;
      RECT  190.4 156.8 191.2 157.6 ;
      RECT  186.9 150.3 193.7 150.9 ;
      RECT  197.2 152.4 198.0 153.2 ;
      RECT  195.2 152.4 196.0 153.2 ;
      RECT  197.2 156.8 198.0 157.6 ;
      RECT  195.2 156.8 196.0 157.6 ;
      RECT  199.2 156.8 200.0 157.6 ;
      RECT  197.2 156.8 198.0 157.6 ;
      RECT  193.7 150.3 200.5 150.9 ;
      RECT  180.1 150.3 200.5 150.9 ;
      RECT  189.7 116.6 190.5 121.4 ;
      RECT  192.3 125.8 193.1 127.0 ;
      RECT  191.5 133.6 192.3 136.0 ;
      RECT  189.9 134.2 190.7 136.0 ;
      RECT  193.3 140.0 194.1 140.8 ;
      RECT  188.1 117.2 188.9 121.4 ;
      RECT  189.9 127.0 193.1 127.6 ;
      RECT  188.3 126.4 189.1 136.0 ;
      RECT  193.1 121.4 193.7 122.8 ;
      RECT  186.5 142.4 194.1 143.2 ;
      RECT  188.3 125.6 189.5 126.4 ;
      RECT  188.1 122.8 189.5 123.4 ;
      RECT  188.7 123.4 189.5 123.6 ;
      RECT  191.7 140.0 192.5 140.4 ;
      RECT  191.3 116.6 192.1 122.2 ;
      RECT  189.5 121.4 190.3 122.2 ;
      RECT  188.1 121.4 188.7 122.8 ;
      RECT  190.1 136.0 190.7 138.6 ;
      RECT  192.9 116.6 193.7 121.4 ;
      RECT  190.1 138.6 190.9 140.4 ;
      RECT  187.5 114.8 188.3 116.6 ;
      RECT  191.5 128.2 192.3 132.8 ;
      RECT  187.5 116.6 188.9 117.2 ;
      RECT  192.7 122.8 193.7 123.6 ;
      RECT  189.9 128.2 190.7 131.8 ;
      RECT  191.7 139.2 194.1 140.0 ;
      RECT  189.9 127.6 190.5 128.2 ;
      RECT  191.5 132.8 192.9 133.6 ;
      RECT  191.7 138.6 192.5 139.2 ;
      RECT  196.5 116.6 197.3 121.4 ;
      RECT  199.1 125.8 199.9 127.0 ;
      RECT  198.3 133.6 199.1 136.0 ;
      RECT  196.7 134.2 197.5 136.0 ;
      RECT  200.1 140.0 200.9 140.8 ;
      RECT  194.9 117.2 195.7 121.4 ;
      RECT  196.7 127.0 199.9 127.6 ;
      RECT  195.1 126.4 195.9 136.0 ;
      RECT  199.9 121.4 200.5 122.8 ;
      RECT  193.3 142.4 200.9 143.2 ;
      RECT  195.1 125.6 196.3 126.4 ;
      RECT  194.9 122.8 196.3 123.4 ;
      RECT  195.5 123.4 196.3 123.6 ;
      RECT  198.5 140.0 199.3 140.4 ;
      RECT  198.1 116.6 198.9 122.2 ;
      RECT  196.3 121.4 197.1 122.2 ;
      RECT  194.9 121.4 195.5 122.8 ;
      RECT  196.9 136.0 197.5 138.6 ;
      RECT  199.7 116.6 200.5 121.4 ;
      RECT  196.9 138.6 197.7 140.4 ;
      RECT  194.3 114.8 195.1 116.6 ;
      RECT  198.3 128.2 199.1 132.8 ;
      RECT  194.3 116.6 195.7 117.2 ;
      RECT  199.5 122.8 200.5 123.6 ;
      RECT  196.7 128.2 197.5 131.8 ;
      RECT  198.5 139.2 200.9 140.0 ;
      RECT  196.7 127.6 197.3 128.2 ;
      RECT  198.3 132.8 199.7 133.6 ;
      RECT  198.5 138.6 199.3 139.2 ;
      RECT  186.9 142.5 200.5 143.1 ;
      RECT  187.9 84.2 188.7 88.0 ;
      RECT  191.1 87.0 192.3 87.8 ;
      RECT  187.5 72.6 193.1 73.4 ;
      RECT  187.9 106.4 189.7 107.2 ;
      RECT  187.5 74.8 188.3 76.8 ;
      RECT  190.9 92.8 191.7 95.4 ;
      RECT  189.5 89.2 190.3 91.4 ;
      RECT  187.5 74.0 191.5 74.8 ;
      RECT  189.5 84.2 190.3 85.6 ;
      RECT  187.9 88.6 188.7 90.6 ;
      RECT  189.1 75.4 189.9 77.4 ;
      RECT  187.5 78.0 188.3 80.6 ;
      RECT  190.9 96.2 191.7 97.4 ;
      RECT  187.7 92.8 188.5 101.4 ;
      RECT  187.9 88.0 191.9 88.6 ;
      RECT  189.3 91.4 190.9 92.2 ;
      RECT  190.7 74.8 191.5 76.8 ;
      RECT  191.1 88.6 191.9 90.6 ;
      RECT  189.1 79.2 189.9 80.6 ;
      RECT  191.1 87.8 191.9 88.0 ;
      RECT  190.9 103.4 191.7 106.6 ;
      RECT  189.3 92.2 190.1 94.2 ;
      RECT  190.9 95.4 193.5 96.2 ;
      RECT  187.5 82.0 188.3 82.8 ;
      RECT  191.9 85.6 192.9 85.8 ;
      RECT  187.9 105.8 188.5 106.4 ;
      RECT  189.3 96.6 190.1 105.8 ;
      RECT  187.7 103.4 188.5 105.8 ;
      RECT  187.5 77.4 189.9 78.0 ;
      RECT  192.5 104.2 193.5 105.0 ;
      RECT  187.7 80.6 188.3 82.0 ;
      RECT  189.9 69.0 190.7 70.6 ;
      RECT  190.7 79.2 191.5 81.4 ;
      RECT  192.9 96.2 193.5 104.2 ;
      RECT  191.5 82.8 193.1 83.6 ;
      RECT  191.1 84.2 192.9 85.6 ;
      RECT  192.3 75.4 193.1 82.8 ;
      RECT  194.7 84.2 195.5 88.0 ;
      RECT  197.9 87.0 199.1 87.8 ;
      RECT  194.3 72.6 199.9 73.4 ;
      RECT  194.7 106.4 196.5 107.2 ;
      RECT  194.3 74.8 195.1 76.8 ;
      RECT  197.7 92.8 198.5 95.4 ;
      RECT  196.3 89.2 197.1 91.4 ;
      RECT  194.3 74.0 198.3 74.8 ;
      RECT  196.3 84.2 197.1 85.6 ;
      RECT  194.7 88.6 195.5 90.6 ;
      RECT  195.9 75.4 196.7 77.4 ;
      RECT  194.3 78.0 195.1 80.6 ;
      RECT  197.7 96.2 198.5 97.4 ;
      RECT  194.5 92.8 195.3 101.4 ;
      RECT  194.7 88.0 198.7 88.6 ;
      RECT  196.1 91.4 197.7 92.2 ;
      RECT  197.5 74.8 198.3 76.8 ;
      RECT  197.9 88.6 198.7 90.6 ;
      RECT  195.9 79.2 196.7 80.6 ;
      RECT  197.9 87.8 198.7 88.0 ;
      RECT  197.7 103.4 198.5 106.6 ;
      RECT  196.1 92.2 196.9 94.2 ;
      RECT  197.7 95.4 200.3 96.2 ;
      RECT  194.3 82.0 195.1 82.8 ;
      RECT  198.7 85.6 199.7 85.8 ;
      RECT  194.7 105.8 195.3 106.4 ;
      RECT  196.1 96.6 196.9 105.8 ;
      RECT  194.5 103.4 195.3 105.8 ;
      RECT  194.3 77.4 196.7 78.0 ;
      RECT  199.3 104.2 200.3 105.0 ;
      RECT  194.5 80.6 195.1 82.0 ;
      RECT  196.7 69.0 197.5 70.6 ;
      RECT  197.5 79.2 198.3 81.4 ;
      RECT  199.7 96.2 200.3 104.2 ;
      RECT  198.3 82.8 199.9 83.6 ;
      RECT  197.9 84.2 199.7 85.6 ;
      RECT  199.1 75.4 199.9 82.8 ;
      RECT  186.9 72.6 200.5 73.2 ;
      RECT  186.9 143.1 200.5 142.5 ;
      RECT  180.1 150.9 200.5 150.3 ;
      RECT  186.9 73.2 200.5 72.6 ;
      RECT  97.3 195.1 98.1 195.9 ;
      RECT  95.3 195.1 96.1 195.9 ;
      RECT  97.3 187.7 98.1 188.5 ;
      RECT  95.3 187.7 96.1 188.5 ;
      RECT  95.7 191.4 96.5 192.2 ;
      RECT  97.7 191.5 98.3 192.1 ;
      RECT  94.1 196.9 100.7 197.5 ;
      RECT  94.1 186.5 100.7 187.1 ;
      RECT  97.3 199.3 98.1 198.5 ;
      RECT  95.3 199.3 96.1 198.5 ;
      RECT  97.3 206.7 98.1 205.9 ;
      RECT  95.3 206.7 96.1 205.9 ;
      RECT  95.7 203.0 96.5 202.2 ;
      RECT  97.7 202.9 98.3 202.3 ;
      RECT  94.1 197.5 100.7 196.9 ;
      RECT  94.1 207.9 100.7 207.3 ;
      RECT  112.3 195.1 113.1 195.9 ;
      RECT  110.3 195.1 111.1 195.9 ;
      RECT  114.3 195.1 115.1 195.9 ;
      RECT  112.3 195.1 113.1 195.9 ;
      RECT  110.3 188.1 111.1 188.9 ;
      RECT  114.3 188.1 115.1 188.9 ;
      RECT  111.3 189.6 112.1 190.4 ;
      RECT  113.3 192.4 114.1 193.2 ;
      RECT  115.8 193.8 116.4 194.4 ;
      RECT  109.1 196.9 117.7 197.5 ;
      RECT  109.1 186.5 117.7 187.1 ;
      RECT  120.9 195.1 121.7 195.9 ;
      RECT  118.9 195.1 119.7 195.9 ;
      RECT  120.9 187.7 121.7 188.5 ;
      RECT  118.9 187.7 119.7 188.5 ;
      RECT  119.3 191.4 120.1 192.2 ;
      RECT  121.3 191.5 121.9 192.1 ;
      RECT  117.7 196.9 124.3 197.5 ;
      RECT  117.7 186.5 124.3 187.1 ;
      RECT  111.3 189.6 112.1 190.4 ;
      RECT  113.3 192.4 114.1 193.2 ;
      RECT  121.3 191.5 121.9 192.1 ;
      RECT  109.1 196.9 124.3 197.5 ;
      RECT  109.1 186.5 124.3 187.1 ;
      RECT  112.3 199.3 113.1 198.5 ;
      RECT  110.3 199.3 111.1 198.5 ;
      RECT  114.3 199.3 115.1 198.5 ;
      RECT  112.3 199.3 113.1 198.5 ;
      RECT  110.3 206.3 111.1 205.5 ;
      RECT  114.3 206.3 115.1 205.5 ;
      RECT  111.3 204.8 112.1 204.0 ;
      RECT  113.3 202.0 114.1 201.2 ;
      RECT  115.8 200.6 116.4 200.0 ;
      RECT  109.1 197.5 117.7 196.9 ;
      RECT  109.1 207.9 117.7 207.3 ;
      RECT  120.9 199.3 121.7 198.5 ;
      RECT  118.9 199.3 119.7 198.5 ;
      RECT  120.9 206.7 121.7 205.9 ;
      RECT  118.9 206.7 119.7 205.9 ;
      RECT  119.3 203.0 120.1 202.2 ;
      RECT  121.3 202.9 121.9 202.3 ;
      RECT  117.7 197.5 124.3 196.9 ;
      RECT  117.7 207.9 124.3 207.3 ;
      RECT  111.3 204.8 112.1 204.0 ;
      RECT  113.3 202.0 114.1 201.2 ;
      RECT  121.3 202.9 121.9 202.3 ;
      RECT  109.1 197.5 124.3 196.9 ;
      RECT  109.1 207.9 124.3 207.3 ;
      RECT  112.3 215.9 113.1 216.7 ;
      RECT  110.3 215.9 111.1 216.7 ;
      RECT  114.3 215.9 115.1 216.7 ;
      RECT  112.3 215.9 113.1 216.7 ;
      RECT  110.3 208.9 111.1 209.7 ;
      RECT  114.3 208.9 115.1 209.7 ;
      RECT  111.3 210.4 112.1 211.2 ;
      RECT  113.3 213.2 114.1 214.0 ;
      RECT  115.8 214.6 116.4 215.2 ;
      RECT  109.1 217.7 117.7 218.3 ;
      RECT  109.1 207.3 117.7 207.9 ;
      RECT  120.9 215.9 121.7 216.7 ;
      RECT  118.9 215.9 119.7 216.7 ;
      RECT  120.9 208.5 121.7 209.3 ;
      RECT  118.9 208.5 119.7 209.3 ;
      RECT  119.3 212.2 120.1 213.0 ;
      RECT  121.3 212.3 121.9 212.9 ;
      RECT  117.7 217.7 124.3 218.3 ;
      RECT  117.7 207.3 124.3 207.9 ;
      RECT  111.3 210.4 112.1 211.2 ;
      RECT  113.3 213.2 114.1 214.0 ;
      RECT  121.3 212.3 121.9 212.9 ;
      RECT  109.1 217.7 124.3 218.3 ;
      RECT  109.1 207.3 124.3 207.9 ;
      RECT  112.3 220.1 113.1 219.3 ;
      RECT  110.3 220.1 111.1 219.3 ;
      RECT  114.3 220.1 115.1 219.3 ;
      RECT  112.3 220.1 113.1 219.3 ;
      RECT  110.3 227.1 111.1 226.3 ;
      RECT  114.3 227.1 115.1 226.3 ;
      RECT  111.3 225.6 112.1 224.8 ;
      RECT  113.3 222.8 114.1 222.0 ;
      RECT  115.8 221.4 116.4 220.8 ;
      RECT  109.1 218.3 117.7 217.7 ;
      RECT  109.1 228.7 117.7 228.1 ;
      RECT  120.9 220.1 121.7 219.3 ;
      RECT  118.9 220.1 119.7 219.3 ;
      RECT  120.9 227.5 121.7 226.7 ;
      RECT  118.9 227.5 119.7 226.7 ;
      RECT  119.3 223.8 120.1 223.0 ;
      RECT  121.3 223.7 121.9 223.1 ;
      RECT  117.7 218.3 124.3 217.7 ;
      RECT  117.7 228.7 124.3 228.1 ;
      RECT  111.3 225.6 112.1 224.8 ;
      RECT  113.3 222.8 114.1 222.0 ;
      RECT  121.3 223.7 121.9 223.1 ;
      RECT  109.1 218.3 124.3 217.7 ;
      RECT  109.1 228.7 124.3 228.1 ;
      RECT  121.3 191.5 121.9 192.1 ;
      RECT  121.3 202.3 121.9 202.9 ;
      RECT  121.3 212.3 121.9 212.9 ;
      RECT  121.3 223.1 121.9 223.7 ;
      RECT  97.3 257.5 98.1 258.3 ;
      RECT  95.3 257.5 96.1 258.3 ;
      RECT  97.3 250.1 98.1 250.9 ;
      RECT  95.3 250.1 96.1 250.9 ;
      RECT  95.7 253.8 96.5 254.6 ;
      RECT  97.7 253.9 98.3 254.5 ;
      RECT  94.1 259.3 100.7 259.9 ;
      RECT  94.1 248.9 100.7 249.5 ;
      RECT  97.3 261.7 98.1 260.9 ;
      RECT  95.3 261.7 96.1 260.9 ;
      RECT  97.3 269.1 98.1 268.3 ;
      RECT  95.3 269.1 96.1 268.3 ;
      RECT  95.7 265.4 96.5 264.6 ;
      RECT  97.7 265.3 98.3 264.7 ;
      RECT  94.1 259.9 100.7 259.3 ;
      RECT  94.1 270.3 100.7 269.7 ;
      RECT  112.3 257.5 113.1 258.3 ;
      RECT  110.3 257.5 111.1 258.3 ;
      RECT  114.3 257.5 115.1 258.3 ;
      RECT  112.3 257.5 113.1 258.3 ;
      RECT  110.3 250.5 111.1 251.3 ;
      RECT  114.3 250.5 115.1 251.3 ;
      RECT  111.3 252.0 112.1 252.8 ;
      RECT  113.3 254.8 114.1 255.6 ;
      RECT  115.8 256.2 116.4 256.8 ;
      RECT  109.1 259.3 117.7 259.9 ;
      RECT  109.1 248.9 117.7 249.5 ;
      RECT  120.9 257.5 121.7 258.3 ;
      RECT  118.9 257.5 119.7 258.3 ;
      RECT  120.9 250.1 121.7 250.9 ;
      RECT  118.9 250.1 119.7 250.9 ;
      RECT  119.3 253.8 120.1 254.6 ;
      RECT  121.3 253.9 121.9 254.5 ;
      RECT  117.7 259.3 124.3 259.9 ;
      RECT  117.7 248.9 124.3 249.5 ;
      RECT  111.3 252.0 112.1 252.8 ;
      RECT  113.3 254.8 114.1 255.6 ;
      RECT  121.3 253.9 121.9 254.5 ;
      RECT  109.1 259.3 124.3 259.9 ;
      RECT  109.1 248.9 124.3 249.5 ;
      RECT  112.3 261.7 113.1 260.9 ;
      RECT  110.3 261.7 111.1 260.9 ;
      RECT  114.3 261.7 115.1 260.9 ;
      RECT  112.3 261.7 113.1 260.9 ;
      RECT  110.3 268.7 111.1 267.9 ;
      RECT  114.3 268.7 115.1 267.9 ;
      RECT  111.3 267.2 112.1 266.4 ;
      RECT  113.3 264.4 114.1 263.6 ;
      RECT  115.8 263.0 116.4 262.4 ;
      RECT  109.1 259.9 117.7 259.3 ;
      RECT  109.1 270.3 117.7 269.7 ;
      RECT  120.9 261.7 121.7 260.9 ;
      RECT  118.9 261.7 119.7 260.9 ;
      RECT  120.9 269.1 121.7 268.3 ;
      RECT  118.9 269.1 119.7 268.3 ;
      RECT  119.3 265.4 120.1 264.6 ;
      RECT  121.3 265.3 121.9 264.7 ;
      RECT  117.7 259.9 124.3 259.3 ;
      RECT  117.7 270.3 124.3 269.7 ;
      RECT  111.3 267.2 112.1 266.4 ;
      RECT  113.3 264.4 114.1 263.6 ;
      RECT  121.3 265.3 121.9 264.7 ;
      RECT  109.1 259.9 124.3 259.3 ;
      RECT  109.1 270.3 124.3 269.7 ;
      RECT  112.3 278.3 113.1 279.1 ;
      RECT  110.3 278.3 111.1 279.1 ;
      RECT  114.3 278.3 115.1 279.1 ;
      RECT  112.3 278.3 113.1 279.1 ;
      RECT  110.3 271.3 111.1 272.1 ;
      RECT  114.3 271.3 115.1 272.1 ;
      RECT  111.3 272.8 112.1 273.6 ;
      RECT  113.3 275.6 114.1 276.4 ;
      RECT  115.8 277.0 116.4 277.6 ;
      RECT  109.1 280.1 117.7 280.7 ;
      RECT  109.1 269.7 117.7 270.3 ;
      RECT  120.9 278.3 121.7 279.1 ;
      RECT  118.9 278.3 119.7 279.1 ;
      RECT  120.9 270.9 121.7 271.7 ;
      RECT  118.9 270.9 119.7 271.7 ;
      RECT  119.3 274.6 120.1 275.4 ;
      RECT  121.3 274.7 121.9 275.3 ;
      RECT  117.7 280.1 124.3 280.7 ;
      RECT  117.7 269.7 124.3 270.3 ;
      RECT  111.3 272.8 112.1 273.6 ;
      RECT  113.3 275.6 114.1 276.4 ;
      RECT  121.3 274.7 121.9 275.3 ;
      RECT  109.1 280.1 124.3 280.7 ;
      RECT  109.1 269.7 124.3 270.3 ;
      RECT  112.3 282.5 113.1 281.7 ;
      RECT  110.3 282.5 111.1 281.7 ;
      RECT  114.3 282.5 115.1 281.7 ;
      RECT  112.3 282.5 113.1 281.7 ;
      RECT  110.3 289.5 111.1 288.7 ;
      RECT  114.3 289.5 115.1 288.7 ;
      RECT  111.3 288.0 112.1 287.2 ;
      RECT  113.3 285.2 114.1 284.4 ;
      RECT  115.8 283.8 116.4 283.2 ;
      RECT  109.1 280.7 117.7 280.1 ;
      RECT  109.1 291.1 117.7 290.5 ;
      RECT  120.9 282.5 121.7 281.7 ;
      RECT  118.9 282.5 119.7 281.7 ;
      RECT  120.9 289.9 121.7 289.1 ;
      RECT  118.9 289.9 119.7 289.1 ;
      RECT  119.3 286.2 120.1 285.4 ;
      RECT  121.3 286.1 121.9 285.5 ;
      RECT  117.7 280.7 124.3 280.1 ;
      RECT  117.7 291.1 124.3 290.5 ;
      RECT  111.3 288.0 112.1 287.2 ;
      RECT  113.3 285.2 114.1 284.4 ;
      RECT  121.3 286.1 121.9 285.5 ;
      RECT  109.1 280.7 124.3 280.1 ;
      RECT  109.1 291.1 124.3 290.5 ;
      RECT  121.3 253.9 121.9 254.5 ;
      RECT  121.3 264.7 121.9 265.3 ;
      RECT  121.3 274.7 121.9 275.3 ;
      RECT  121.3 285.5 121.9 286.1 ;
      RECT  140.1 195.1 140.9 195.9 ;
      RECT  138.1 195.1 138.9 195.9 ;
      RECT  142.1 195.1 142.9 195.9 ;
      RECT  140.1 195.1 140.9 195.9 ;
      RECT  138.1 188.1 138.9 188.9 ;
      RECT  142.1 188.1 142.9 188.9 ;
      RECT  139.1 189.6 139.9 190.4 ;
      RECT  141.1 192.4 141.9 193.2 ;
      RECT  143.6 193.8 144.2 194.4 ;
      RECT  136.9 196.9 145.5 197.5 ;
      RECT  136.9 186.5 145.5 187.1 ;
      RECT  148.7 195.1 149.5 195.9 ;
      RECT  146.7 195.1 147.5 195.9 ;
      RECT  148.7 187.7 149.5 188.5 ;
      RECT  146.7 187.7 147.5 188.5 ;
      RECT  147.1 191.4 147.9 192.2 ;
      RECT  149.1 191.5 149.7 192.1 ;
      RECT  145.5 196.9 152.1 197.5 ;
      RECT  145.5 186.5 152.1 187.1 ;
      RECT  139.1 189.6 139.9 190.4 ;
      RECT  141.1 192.4 141.9 193.2 ;
      RECT  149.1 191.5 149.7 192.1 ;
      RECT  136.9 196.9 152.1 197.5 ;
      RECT  136.9 186.5 152.1 187.1 ;
      RECT  140.1 199.3 140.9 198.5 ;
      RECT  138.1 199.3 138.9 198.5 ;
      RECT  142.1 199.3 142.9 198.5 ;
      RECT  140.1 199.3 140.9 198.5 ;
      RECT  138.1 206.3 138.9 205.5 ;
      RECT  142.1 206.3 142.9 205.5 ;
      RECT  139.1 204.8 139.9 204.0 ;
      RECT  141.1 202.0 141.9 201.2 ;
      RECT  143.6 200.6 144.2 200.0 ;
      RECT  136.9 197.5 145.5 196.9 ;
      RECT  136.9 207.9 145.5 207.3 ;
      RECT  148.7 199.3 149.5 198.5 ;
      RECT  146.7 199.3 147.5 198.5 ;
      RECT  148.7 206.7 149.5 205.9 ;
      RECT  146.7 206.7 147.5 205.9 ;
      RECT  147.1 203.0 147.9 202.2 ;
      RECT  149.1 202.9 149.7 202.3 ;
      RECT  145.5 197.5 152.1 196.9 ;
      RECT  145.5 207.9 152.1 207.3 ;
      RECT  139.1 204.8 139.9 204.0 ;
      RECT  141.1 202.0 141.9 201.2 ;
      RECT  149.1 202.9 149.7 202.3 ;
      RECT  136.9 197.5 152.1 196.9 ;
      RECT  136.9 207.9 152.1 207.3 ;
      RECT  140.1 215.9 140.9 216.7 ;
      RECT  138.1 215.9 138.9 216.7 ;
      RECT  142.1 215.9 142.9 216.7 ;
      RECT  140.1 215.9 140.9 216.7 ;
      RECT  138.1 208.9 138.9 209.7 ;
      RECT  142.1 208.9 142.9 209.7 ;
      RECT  139.1 210.4 139.9 211.2 ;
      RECT  141.1 213.2 141.9 214.0 ;
      RECT  143.6 214.6 144.2 215.2 ;
      RECT  136.9 217.7 145.5 218.3 ;
      RECT  136.9 207.3 145.5 207.9 ;
      RECT  148.7 215.9 149.5 216.7 ;
      RECT  146.7 215.9 147.5 216.7 ;
      RECT  148.7 208.5 149.5 209.3 ;
      RECT  146.7 208.5 147.5 209.3 ;
      RECT  147.1 212.2 147.9 213.0 ;
      RECT  149.1 212.3 149.7 212.9 ;
      RECT  145.5 217.7 152.1 218.3 ;
      RECT  145.5 207.3 152.1 207.9 ;
      RECT  139.1 210.4 139.9 211.2 ;
      RECT  141.1 213.2 141.9 214.0 ;
      RECT  149.1 212.3 149.7 212.9 ;
      RECT  136.9 217.7 152.1 218.3 ;
      RECT  136.9 207.3 152.1 207.9 ;
      RECT  140.1 220.1 140.9 219.3 ;
      RECT  138.1 220.1 138.9 219.3 ;
      RECT  142.1 220.1 142.9 219.3 ;
      RECT  140.1 220.1 140.9 219.3 ;
      RECT  138.1 227.1 138.9 226.3 ;
      RECT  142.1 227.1 142.9 226.3 ;
      RECT  139.1 225.6 139.9 224.8 ;
      RECT  141.1 222.8 141.9 222.0 ;
      RECT  143.6 221.4 144.2 220.8 ;
      RECT  136.9 218.3 145.5 217.7 ;
      RECT  136.9 228.7 145.5 228.1 ;
      RECT  148.7 220.1 149.5 219.3 ;
      RECT  146.7 220.1 147.5 219.3 ;
      RECT  148.7 227.5 149.5 226.7 ;
      RECT  146.7 227.5 147.5 226.7 ;
      RECT  147.1 223.8 147.9 223.0 ;
      RECT  149.1 223.7 149.7 223.1 ;
      RECT  145.5 218.3 152.1 217.7 ;
      RECT  145.5 228.7 152.1 228.1 ;
      RECT  139.1 225.6 139.9 224.8 ;
      RECT  141.1 222.8 141.9 222.0 ;
      RECT  149.1 223.7 149.7 223.1 ;
      RECT  136.9 218.3 152.1 217.7 ;
      RECT  136.9 228.7 152.1 228.1 ;
      RECT  140.1 236.7 140.9 237.5 ;
      RECT  138.1 236.7 138.9 237.5 ;
      RECT  142.1 236.7 142.9 237.5 ;
      RECT  140.1 236.7 140.9 237.5 ;
      RECT  138.1 229.7 138.9 230.5 ;
      RECT  142.1 229.7 142.9 230.5 ;
      RECT  139.1 231.2 139.9 232.0 ;
      RECT  141.1 234.0 141.9 234.8 ;
      RECT  143.6 235.4 144.2 236.0 ;
      RECT  136.9 238.5 145.5 239.1 ;
      RECT  136.9 228.1 145.5 228.7 ;
      RECT  148.7 236.7 149.5 237.5 ;
      RECT  146.7 236.7 147.5 237.5 ;
      RECT  148.7 229.3 149.5 230.1 ;
      RECT  146.7 229.3 147.5 230.1 ;
      RECT  147.1 233.0 147.9 233.8 ;
      RECT  149.1 233.1 149.7 233.7 ;
      RECT  145.5 238.5 152.1 239.1 ;
      RECT  145.5 228.1 152.1 228.7 ;
      RECT  139.1 231.2 139.9 232.0 ;
      RECT  141.1 234.0 141.9 234.8 ;
      RECT  149.1 233.1 149.7 233.7 ;
      RECT  136.9 238.5 152.1 239.1 ;
      RECT  136.9 228.1 152.1 228.7 ;
      RECT  140.1 240.9 140.9 240.1 ;
      RECT  138.1 240.9 138.9 240.1 ;
      RECT  142.1 240.9 142.9 240.1 ;
      RECT  140.1 240.9 140.9 240.1 ;
      RECT  138.1 247.9 138.9 247.1 ;
      RECT  142.1 247.9 142.9 247.1 ;
      RECT  139.1 246.4 139.9 245.6 ;
      RECT  141.1 243.6 141.9 242.8 ;
      RECT  143.6 242.2 144.2 241.6 ;
      RECT  136.9 239.1 145.5 238.5 ;
      RECT  136.9 249.5 145.5 248.9 ;
      RECT  148.7 240.9 149.5 240.1 ;
      RECT  146.7 240.9 147.5 240.1 ;
      RECT  148.7 248.3 149.5 247.5 ;
      RECT  146.7 248.3 147.5 247.5 ;
      RECT  147.1 244.6 147.9 243.8 ;
      RECT  149.1 244.5 149.7 243.9 ;
      RECT  145.5 239.1 152.1 238.5 ;
      RECT  145.5 249.5 152.1 248.9 ;
      RECT  139.1 246.4 139.9 245.6 ;
      RECT  141.1 243.6 141.9 242.8 ;
      RECT  149.1 244.5 149.7 243.9 ;
      RECT  136.9 239.1 152.1 238.5 ;
      RECT  136.9 249.5 152.1 248.9 ;
      RECT  140.1 257.5 140.9 258.3 ;
      RECT  138.1 257.5 138.9 258.3 ;
      RECT  142.1 257.5 142.9 258.3 ;
      RECT  140.1 257.5 140.9 258.3 ;
      RECT  138.1 250.5 138.9 251.3 ;
      RECT  142.1 250.5 142.9 251.3 ;
      RECT  139.1 252.0 139.9 252.8 ;
      RECT  141.1 254.8 141.9 255.6 ;
      RECT  143.6 256.2 144.2 256.8 ;
      RECT  136.9 259.3 145.5 259.9 ;
      RECT  136.9 248.9 145.5 249.5 ;
      RECT  148.7 257.5 149.5 258.3 ;
      RECT  146.7 257.5 147.5 258.3 ;
      RECT  148.7 250.1 149.5 250.9 ;
      RECT  146.7 250.1 147.5 250.9 ;
      RECT  147.1 253.8 147.9 254.6 ;
      RECT  149.1 253.9 149.7 254.5 ;
      RECT  145.5 259.3 152.1 259.9 ;
      RECT  145.5 248.9 152.1 249.5 ;
      RECT  139.1 252.0 139.9 252.8 ;
      RECT  141.1 254.8 141.9 255.6 ;
      RECT  149.1 253.9 149.7 254.5 ;
      RECT  136.9 259.3 152.1 259.9 ;
      RECT  136.9 248.9 152.1 249.5 ;
      RECT  140.1 261.7 140.9 260.9 ;
      RECT  138.1 261.7 138.9 260.9 ;
      RECT  142.1 261.7 142.9 260.9 ;
      RECT  140.1 261.7 140.9 260.9 ;
      RECT  138.1 268.7 138.9 267.9 ;
      RECT  142.1 268.7 142.9 267.9 ;
      RECT  139.1 267.2 139.9 266.4 ;
      RECT  141.1 264.4 141.9 263.6 ;
      RECT  143.6 263.0 144.2 262.4 ;
      RECT  136.9 259.9 145.5 259.3 ;
      RECT  136.9 270.3 145.5 269.7 ;
      RECT  148.7 261.7 149.5 260.9 ;
      RECT  146.7 261.7 147.5 260.9 ;
      RECT  148.7 269.1 149.5 268.3 ;
      RECT  146.7 269.1 147.5 268.3 ;
      RECT  147.1 265.4 147.9 264.6 ;
      RECT  149.1 265.3 149.7 264.7 ;
      RECT  145.5 259.9 152.1 259.3 ;
      RECT  145.5 270.3 152.1 269.7 ;
      RECT  139.1 267.2 139.9 266.4 ;
      RECT  141.1 264.4 141.9 263.6 ;
      RECT  149.1 265.3 149.7 264.7 ;
      RECT  136.9 259.9 152.1 259.3 ;
      RECT  136.9 270.3 152.1 269.7 ;
      RECT  140.1 278.3 140.9 279.1 ;
      RECT  138.1 278.3 138.9 279.1 ;
      RECT  142.1 278.3 142.9 279.1 ;
      RECT  140.1 278.3 140.9 279.1 ;
      RECT  138.1 271.3 138.9 272.1 ;
      RECT  142.1 271.3 142.9 272.1 ;
      RECT  139.1 272.8 139.9 273.6 ;
      RECT  141.1 275.6 141.9 276.4 ;
      RECT  143.6 277.0 144.2 277.6 ;
      RECT  136.9 280.1 145.5 280.7 ;
      RECT  136.9 269.7 145.5 270.3 ;
      RECT  148.7 278.3 149.5 279.1 ;
      RECT  146.7 278.3 147.5 279.1 ;
      RECT  148.7 270.9 149.5 271.7 ;
      RECT  146.7 270.9 147.5 271.7 ;
      RECT  147.1 274.6 147.9 275.4 ;
      RECT  149.1 274.7 149.7 275.3 ;
      RECT  145.5 280.1 152.1 280.7 ;
      RECT  145.5 269.7 152.1 270.3 ;
      RECT  139.1 272.8 139.9 273.6 ;
      RECT  141.1 275.6 141.9 276.4 ;
      RECT  149.1 274.7 149.7 275.3 ;
      RECT  136.9 280.1 152.1 280.7 ;
      RECT  136.9 269.7 152.1 270.3 ;
      RECT  140.1 282.5 140.9 281.7 ;
      RECT  138.1 282.5 138.9 281.7 ;
      RECT  142.1 282.5 142.9 281.7 ;
      RECT  140.1 282.5 140.9 281.7 ;
      RECT  138.1 289.5 138.9 288.7 ;
      RECT  142.1 289.5 142.9 288.7 ;
      RECT  139.1 288.0 139.9 287.2 ;
      RECT  141.1 285.2 141.9 284.4 ;
      RECT  143.6 283.8 144.2 283.2 ;
      RECT  136.9 280.7 145.5 280.1 ;
      RECT  136.9 291.1 145.5 290.5 ;
      RECT  148.7 282.5 149.5 281.7 ;
      RECT  146.7 282.5 147.5 281.7 ;
      RECT  148.7 289.9 149.5 289.1 ;
      RECT  146.7 289.9 147.5 289.1 ;
      RECT  147.1 286.2 147.9 285.4 ;
      RECT  149.1 286.1 149.7 285.5 ;
      RECT  145.5 280.7 152.1 280.1 ;
      RECT  145.5 291.1 152.1 290.5 ;
      RECT  139.1 288.0 139.9 287.2 ;
      RECT  141.1 285.2 141.9 284.4 ;
      RECT  149.1 286.1 149.7 285.5 ;
      RECT  136.9 280.7 152.1 280.1 ;
      RECT  136.9 291.1 152.1 290.5 ;
      RECT  140.1 299.1 140.9 299.9 ;
      RECT  138.1 299.1 138.9 299.9 ;
      RECT  142.1 299.1 142.9 299.9 ;
      RECT  140.1 299.1 140.9 299.9 ;
      RECT  138.1 292.1 138.9 292.9 ;
      RECT  142.1 292.1 142.9 292.9 ;
      RECT  139.1 293.6 139.9 294.4 ;
      RECT  141.1 296.4 141.9 297.2 ;
      RECT  143.6 297.8 144.2 298.4 ;
      RECT  136.9 300.9 145.5 301.5 ;
      RECT  136.9 290.5 145.5 291.1 ;
      RECT  148.7 299.1 149.5 299.9 ;
      RECT  146.7 299.1 147.5 299.9 ;
      RECT  148.7 291.7 149.5 292.5 ;
      RECT  146.7 291.7 147.5 292.5 ;
      RECT  147.1 295.4 147.9 296.2 ;
      RECT  149.1 295.5 149.7 296.1 ;
      RECT  145.5 300.9 152.1 301.5 ;
      RECT  145.5 290.5 152.1 291.1 ;
      RECT  139.1 293.6 139.9 294.4 ;
      RECT  141.1 296.4 141.9 297.2 ;
      RECT  149.1 295.5 149.7 296.1 ;
      RECT  136.9 300.9 152.1 301.5 ;
      RECT  136.9 290.5 152.1 291.1 ;
      RECT  140.1 303.3 140.9 302.5 ;
      RECT  138.1 303.3 138.9 302.5 ;
      RECT  142.1 303.3 142.9 302.5 ;
      RECT  140.1 303.3 140.9 302.5 ;
      RECT  138.1 310.3 138.9 309.5 ;
      RECT  142.1 310.3 142.9 309.5 ;
      RECT  139.1 308.8 139.9 308.0 ;
      RECT  141.1 306.0 141.9 305.2 ;
      RECT  143.6 304.6 144.2 304.0 ;
      RECT  136.9 301.5 145.5 300.9 ;
      RECT  136.9 311.9 145.5 311.3 ;
      RECT  148.7 303.3 149.5 302.5 ;
      RECT  146.7 303.3 147.5 302.5 ;
      RECT  148.7 310.7 149.5 309.9 ;
      RECT  146.7 310.7 147.5 309.9 ;
      RECT  147.1 307.0 147.9 306.2 ;
      RECT  149.1 306.9 149.7 306.3 ;
      RECT  145.5 301.5 152.1 300.9 ;
      RECT  145.5 311.9 152.1 311.3 ;
      RECT  139.1 308.8 139.9 308.0 ;
      RECT  141.1 306.0 141.9 305.2 ;
      RECT  149.1 306.9 149.7 306.3 ;
      RECT  136.9 301.5 152.1 300.9 ;
      RECT  136.9 311.9 152.1 311.3 ;
      RECT  140.1 319.9 140.9 320.7 ;
      RECT  138.1 319.9 138.9 320.7 ;
      RECT  142.1 319.9 142.9 320.7 ;
      RECT  140.1 319.9 140.9 320.7 ;
      RECT  138.1 312.9 138.9 313.7 ;
      RECT  142.1 312.9 142.9 313.7 ;
      RECT  139.1 314.4 139.9 315.2 ;
      RECT  141.1 317.2 141.9 318.0 ;
      RECT  143.6 318.6 144.2 319.2 ;
      RECT  136.9 321.7 145.5 322.3 ;
      RECT  136.9 311.3 145.5 311.9 ;
      RECT  148.7 319.9 149.5 320.7 ;
      RECT  146.7 319.9 147.5 320.7 ;
      RECT  148.7 312.5 149.5 313.3 ;
      RECT  146.7 312.5 147.5 313.3 ;
      RECT  147.1 316.2 147.9 317.0 ;
      RECT  149.1 316.3 149.7 316.9 ;
      RECT  145.5 321.7 152.1 322.3 ;
      RECT  145.5 311.3 152.1 311.9 ;
      RECT  139.1 314.4 139.9 315.2 ;
      RECT  141.1 317.2 141.9 318.0 ;
      RECT  149.1 316.3 149.7 316.9 ;
      RECT  136.9 321.7 152.1 322.3 ;
      RECT  136.9 311.3 152.1 311.9 ;
      RECT  140.1 324.1 140.9 323.3 ;
      RECT  138.1 324.1 138.9 323.3 ;
      RECT  142.1 324.1 142.9 323.3 ;
      RECT  140.1 324.1 140.9 323.3 ;
      RECT  138.1 331.1 138.9 330.3 ;
      RECT  142.1 331.1 142.9 330.3 ;
      RECT  139.1 329.6 139.9 328.8 ;
      RECT  141.1 326.8 141.9 326.0 ;
      RECT  143.6 325.4 144.2 324.8 ;
      RECT  136.9 322.3 145.5 321.7 ;
      RECT  136.9 332.7 145.5 332.1 ;
      RECT  148.7 324.1 149.5 323.3 ;
      RECT  146.7 324.1 147.5 323.3 ;
      RECT  148.7 331.5 149.5 330.7 ;
      RECT  146.7 331.5 147.5 330.7 ;
      RECT  147.1 327.8 147.9 327.0 ;
      RECT  149.1 327.7 149.7 327.1 ;
      RECT  145.5 322.3 152.1 321.7 ;
      RECT  145.5 332.7 152.1 332.1 ;
      RECT  139.1 329.6 139.9 328.8 ;
      RECT  141.1 326.8 141.9 326.0 ;
      RECT  149.1 327.7 149.7 327.1 ;
      RECT  136.9 322.3 152.1 321.7 ;
      RECT  136.9 332.7 152.1 332.1 ;
      RECT  140.1 340.7 140.9 341.5 ;
      RECT  138.1 340.7 138.9 341.5 ;
      RECT  142.1 340.7 142.9 341.5 ;
      RECT  140.1 340.7 140.9 341.5 ;
      RECT  138.1 333.7 138.9 334.5 ;
      RECT  142.1 333.7 142.9 334.5 ;
      RECT  139.1 335.2 139.9 336.0 ;
      RECT  141.1 338.0 141.9 338.8 ;
      RECT  143.6 339.4 144.2 340.0 ;
      RECT  136.9 342.5 145.5 343.1 ;
      RECT  136.9 332.1 145.5 332.7 ;
      RECT  148.7 340.7 149.5 341.5 ;
      RECT  146.7 340.7 147.5 341.5 ;
      RECT  148.7 333.3 149.5 334.1 ;
      RECT  146.7 333.3 147.5 334.1 ;
      RECT  147.1 337.0 147.9 337.8 ;
      RECT  149.1 337.1 149.7 337.7 ;
      RECT  145.5 342.5 152.1 343.1 ;
      RECT  145.5 332.1 152.1 332.7 ;
      RECT  139.1 335.2 139.9 336.0 ;
      RECT  141.1 338.0 141.9 338.8 ;
      RECT  149.1 337.1 149.7 337.7 ;
      RECT  136.9 342.5 152.1 343.1 ;
      RECT  136.9 332.1 152.1 332.7 ;
      RECT  140.1 344.9 140.9 344.1 ;
      RECT  138.1 344.9 138.9 344.1 ;
      RECT  142.1 344.9 142.9 344.1 ;
      RECT  140.1 344.9 140.9 344.1 ;
      RECT  138.1 351.9 138.9 351.1 ;
      RECT  142.1 351.9 142.9 351.1 ;
      RECT  139.1 350.4 139.9 349.6 ;
      RECT  141.1 347.6 141.9 346.8 ;
      RECT  143.6 346.2 144.2 345.6 ;
      RECT  136.9 343.1 145.5 342.5 ;
      RECT  136.9 353.5 145.5 352.9 ;
      RECT  148.7 344.9 149.5 344.1 ;
      RECT  146.7 344.9 147.5 344.1 ;
      RECT  148.7 352.3 149.5 351.5 ;
      RECT  146.7 352.3 147.5 351.5 ;
      RECT  147.1 348.6 147.9 347.8 ;
      RECT  149.1 348.5 149.7 347.9 ;
      RECT  145.5 343.1 152.1 342.5 ;
      RECT  145.5 353.5 152.1 352.9 ;
      RECT  139.1 350.4 139.9 349.6 ;
      RECT  141.1 347.6 141.9 346.8 ;
      RECT  149.1 348.5 149.7 347.9 ;
      RECT  136.9 343.1 152.1 342.5 ;
      RECT  136.9 353.5 152.1 352.9 ;
      RECT  149.1 191.5 149.7 192.1 ;
      RECT  149.1 202.3 149.7 202.9 ;
      RECT  149.1 212.3 149.7 212.9 ;
      RECT  149.1 223.1 149.7 223.7 ;
      RECT  149.1 233.1 149.7 233.7 ;
      RECT  149.1 243.9 149.7 244.5 ;
      RECT  149.1 253.9 149.7 254.5 ;
      RECT  149.1 264.7 149.7 265.3 ;
      RECT  149.1 274.7 149.7 275.3 ;
      RECT  149.1 285.5 149.7 286.1 ;
      RECT  149.1 295.5 149.7 296.1 ;
      RECT  149.1 306.3 149.7 306.9 ;
      RECT  149.1 316.3 149.7 316.9 ;
      RECT  149.1 327.1 149.7 327.7 ;
      RECT  149.1 337.1 149.7 337.7 ;
      RECT  149.1 347.9 149.7 348.5 ;
      RECT  155.9 195.1 156.7 195.9 ;
      RECT  153.9 195.1 154.7 195.9 ;
      RECT  157.9 195.1 158.7 195.9 ;
      RECT  155.9 195.1 156.7 195.9 ;
      RECT  153.9 188.1 154.7 188.9 ;
      RECT  157.9 188.1 158.7 188.9 ;
      RECT  154.9 189.6 155.7 190.4 ;
      RECT  156.9 192.4 157.7 193.2 ;
      RECT  159.4 193.8 160.0 194.4 ;
      RECT  152.7 196.9 161.3 197.5 ;
      RECT  152.7 186.5 161.3 187.1 ;
      RECT  164.5 194.3 165.3 195.1 ;
      RECT  162.5 194.3 163.3 195.1 ;
      RECT  164.5 188.1 165.3 188.9 ;
      RECT  162.5 188.1 163.3 188.9 ;
      RECT  162.9 191.2 163.7 192.0 ;
      RECT  164.9 191.3 165.5 191.9 ;
      RECT  161.3 196.9 167.9 197.5 ;
      RECT  161.3 186.5 167.9 187.1 ;
      RECT  154.9 189.6 155.7 190.4 ;
      RECT  156.9 192.4 157.7 193.2 ;
      RECT  164.9 191.3 165.5 191.9 ;
      RECT  152.7 196.9 167.9 197.5 ;
      RECT  152.7 186.5 167.9 187.1 ;
      RECT  155.9 199.3 156.7 198.5 ;
      RECT  153.9 199.3 154.7 198.5 ;
      RECT  157.9 199.3 158.7 198.5 ;
      RECT  155.9 199.3 156.7 198.5 ;
      RECT  153.9 206.3 154.7 205.5 ;
      RECT  157.9 206.3 158.7 205.5 ;
      RECT  154.9 204.8 155.7 204.0 ;
      RECT  156.9 202.0 157.7 201.2 ;
      RECT  159.4 200.6 160.0 200.0 ;
      RECT  152.7 197.5 161.3 196.9 ;
      RECT  152.7 207.9 161.3 207.3 ;
      RECT  164.5 200.1 165.3 199.3 ;
      RECT  162.5 200.1 163.3 199.3 ;
      RECT  164.5 206.3 165.3 205.5 ;
      RECT  162.5 206.3 163.3 205.5 ;
      RECT  162.9 203.2 163.7 202.4 ;
      RECT  164.9 203.1 165.5 202.5 ;
      RECT  161.3 197.5 167.9 196.9 ;
      RECT  161.3 207.9 167.9 207.3 ;
      RECT  154.9 204.8 155.7 204.0 ;
      RECT  156.9 202.0 157.7 201.2 ;
      RECT  164.9 203.1 165.5 202.5 ;
      RECT  152.7 197.5 167.9 196.9 ;
      RECT  152.7 207.9 167.9 207.3 ;
      RECT  155.9 215.9 156.7 216.7 ;
      RECT  153.9 215.9 154.7 216.7 ;
      RECT  157.9 215.9 158.7 216.7 ;
      RECT  155.9 215.9 156.7 216.7 ;
      RECT  153.9 208.9 154.7 209.7 ;
      RECT  157.9 208.9 158.7 209.7 ;
      RECT  154.9 210.4 155.7 211.2 ;
      RECT  156.9 213.2 157.7 214.0 ;
      RECT  159.4 214.6 160.0 215.2 ;
      RECT  152.7 217.7 161.3 218.3 ;
      RECT  152.7 207.3 161.3 207.9 ;
      RECT  164.5 215.1 165.3 215.9 ;
      RECT  162.5 215.1 163.3 215.9 ;
      RECT  164.5 208.9 165.3 209.7 ;
      RECT  162.5 208.9 163.3 209.7 ;
      RECT  162.9 212.0 163.7 212.8 ;
      RECT  164.9 212.1 165.5 212.7 ;
      RECT  161.3 217.7 167.9 218.3 ;
      RECT  161.3 207.3 167.9 207.9 ;
      RECT  154.9 210.4 155.7 211.2 ;
      RECT  156.9 213.2 157.7 214.0 ;
      RECT  164.9 212.1 165.5 212.7 ;
      RECT  152.7 217.7 167.9 218.3 ;
      RECT  152.7 207.3 167.9 207.9 ;
      RECT  155.9 220.1 156.7 219.3 ;
      RECT  153.9 220.1 154.7 219.3 ;
      RECT  157.9 220.1 158.7 219.3 ;
      RECT  155.9 220.1 156.7 219.3 ;
      RECT  153.9 227.1 154.7 226.3 ;
      RECT  157.9 227.1 158.7 226.3 ;
      RECT  154.9 225.6 155.7 224.8 ;
      RECT  156.9 222.8 157.7 222.0 ;
      RECT  159.4 221.4 160.0 220.8 ;
      RECT  152.7 218.3 161.3 217.7 ;
      RECT  152.7 228.7 161.3 228.1 ;
      RECT  164.5 220.9 165.3 220.1 ;
      RECT  162.5 220.9 163.3 220.1 ;
      RECT  164.5 227.1 165.3 226.3 ;
      RECT  162.5 227.1 163.3 226.3 ;
      RECT  162.9 224.0 163.7 223.2 ;
      RECT  164.9 223.9 165.5 223.3 ;
      RECT  161.3 218.3 167.9 217.7 ;
      RECT  161.3 228.7 167.9 228.1 ;
      RECT  154.9 225.6 155.7 224.8 ;
      RECT  156.9 222.8 157.7 222.0 ;
      RECT  164.9 223.9 165.5 223.3 ;
      RECT  152.7 218.3 167.9 217.7 ;
      RECT  152.7 228.7 167.9 228.1 ;
      RECT  155.9 236.7 156.7 237.5 ;
      RECT  153.9 236.7 154.7 237.5 ;
      RECT  157.9 236.7 158.7 237.5 ;
      RECT  155.9 236.7 156.7 237.5 ;
      RECT  153.9 229.7 154.7 230.5 ;
      RECT  157.9 229.7 158.7 230.5 ;
      RECT  154.9 231.2 155.7 232.0 ;
      RECT  156.9 234.0 157.7 234.8 ;
      RECT  159.4 235.4 160.0 236.0 ;
      RECT  152.7 238.5 161.3 239.1 ;
      RECT  152.7 228.1 161.3 228.7 ;
      RECT  164.5 235.9 165.3 236.7 ;
      RECT  162.5 235.9 163.3 236.7 ;
      RECT  164.5 229.7 165.3 230.5 ;
      RECT  162.5 229.7 163.3 230.5 ;
      RECT  162.9 232.8 163.7 233.6 ;
      RECT  164.9 232.9 165.5 233.5 ;
      RECT  161.3 238.5 167.9 239.1 ;
      RECT  161.3 228.1 167.9 228.7 ;
      RECT  154.9 231.2 155.7 232.0 ;
      RECT  156.9 234.0 157.7 234.8 ;
      RECT  164.9 232.9 165.5 233.5 ;
      RECT  152.7 238.5 167.9 239.1 ;
      RECT  152.7 228.1 167.9 228.7 ;
      RECT  155.9 240.9 156.7 240.1 ;
      RECT  153.9 240.9 154.7 240.1 ;
      RECT  157.9 240.9 158.7 240.1 ;
      RECT  155.9 240.9 156.7 240.1 ;
      RECT  153.9 247.9 154.7 247.1 ;
      RECT  157.9 247.9 158.7 247.1 ;
      RECT  154.9 246.4 155.7 245.6 ;
      RECT  156.9 243.6 157.7 242.8 ;
      RECT  159.4 242.2 160.0 241.6 ;
      RECT  152.7 239.1 161.3 238.5 ;
      RECT  152.7 249.5 161.3 248.9 ;
      RECT  164.5 241.7 165.3 240.9 ;
      RECT  162.5 241.7 163.3 240.9 ;
      RECT  164.5 247.9 165.3 247.1 ;
      RECT  162.5 247.9 163.3 247.1 ;
      RECT  162.9 244.8 163.7 244.0 ;
      RECT  164.9 244.7 165.5 244.1 ;
      RECT  161.3 239.1 167.9 238.5 ;
      RECT  161.3 249.5 167.9 248.9 ;
      RECT  154.9 246.4 155.7 245.6 ;
      RECT  156.9 243.6 157.7 242.8 ;
      RECT  164.9 244.7 165.5 244.1 ;
      RECT  152.7 239.1 167.9 238.5 ;
      RECT  152.7 249.5 167.9 248.9 ;
      RECT  155.9 257.5 156.7 258.3 ;
      RECT  153.9 257.5 154.7 258.3 ;
      RECT  157.9 257.5 158.7 258.3 ;
      RECT  155.9 257.5 156.7 258.3 ;
      RECT  153.9 250.5 154.7 251.3 ;
      RECT  157.9 250.5 158.7 251.3 ;
      RECT  154.9 252.0 155.7 252.8 ;
      RECT  156.9 254.8 157.7 255.6 ;
      RECT  159.4 256.2 160.0 256.8 ;
      RECT  152.7 259.3 161.3 259.9 ;
      RECT  152.7 248.9 161.3 249.5 ;
      RECT  164.5 256.7 165.3 257.5 ;
      RECT  162.5 256.7 163.3 257.5 ;
      RECT  164.5 250.5 165.3 251.3 ;
      RECT  162.5 250.5 163.3 251.3 ;
      RECT  162.9 253.6 163.7 254.4 ;
      RECT  164.9 253.7 165.5 254.3 ;
      RECT  161.3 259.3 167.9 259.9 ;
      RECT  161.3 248.9 167.9 249.5 ;
      RECT  154.9 252.0 155.7 252.8 ;
      RECT  156.9 254.8 157.7 255.6 ;
      RECT  164.9 253.7 165.5 254.3 ;
      RECT  152.7 259.3 167.9 259.9 ;
      RECT  152.7 248.9 167.9 249.5 ;
      RECT  155.9 261.7 156.7 260.9 ;
      RECT  153.9 261.7 154.7 260.9 ;
      RECT  157.9 261.7 158.7 260.9 ;
      RECT  155.9 261.7 156.7 260.9 ;
      RECT  153.9 268.7 154.7 267.9 ;
      RECT  157.9 268.7 158.7 267.9 ;
      RECT  154.9 267.2 155.7 266.4 ;
      RECT  156.9 264.4 157.7 263.6 ;
      RECT  159.4 263.0 160.0 262.4 ;
      RECT  152.7 259.9 161.3 259.3 ;
      RECT  152.7 270.3 161.3 269.7 ;
      RECT  164.5 262.5 165.3 261.7 ;
      RECT  162.5 262.5 163.3 261.7 ;
      RECT  164.5 268.7 165.3 267.9 ;
      RECT  162.5 268.7 163.3 267.9 ;
      RECT  162.9 265.6 163.7 264.8 ;
      RECT  164.9 265.5 165.5 264.9 ;
      RECT  161.3 259.9 167.9 259.3 ;
      RECT  161.3 270.3 167.9 269.7 ;
      RECT  154.9 267.2 155.7 266.4 ;
      RECT  156.9 264.4 157.7 263.6 ;
      RECT  164.9 265.5 165.5 264.9 ;
      RECT  152.7 259.9 167.9 259.3 ;
      RECT  152.7 270.3 167.9 269.7 ;
      RECT  155.9 278.3 156.7 279.1 ;
      RECT  153.9 278.3 154.7 279.1 ;
      RECT  157.9 278.3 158.7 279.1 ;
      RECT  155.9 278.3 156.7 279.1 ;
      RECT  153.9 271.3 154.7 272.1 ;
      RECT  157.9 271.3 158.7 272.1 ;
      RECT  154.9 272.8 155.7 273.6 ;
      RECT  156.9 275.6 157.7 276.4 ;
      RECT  159.4 277.0 160.0 277.6 ;
      RECT  152.7 280.1 161.3 280.7 ;
      RECT  152.7 269.7 161.3 270.3 ;
      RECT  164.5 277.5 165.3 278.3 ;
      RECT  162.5 277.5 163.3 278.3 ;
      RECT  164.5 271.3 165.3 272.1 ;
      RECT  162.5 271.3 163.3 272.1 ;
      RECT  162.9 274.4 163.7 275.2 ;
      RECT  164.9 274.5 165.5 275.1 ;
      RECT  161.3 280.1 167.9 280.7 ;
      RECT  161.3 269.7 167.9 270.3 ;
      RECT  154.9 272.8 155.7 273.6 ;
      RECT  156.9 275.6 157.7 276.4 ;
      RECT  164.9 274.5 165.5 275.1 ;
      RECT  152.7 280.1 167.9 280.7 ;
      RECT  152.7 269.7 167.9 270.3 ;
      RECT  155.9 282.5 156.7 281.7 ;
      RECT  153.9 282.5 154.7 281.7 ;
      RECT  157.9 282.5 158.7 281.7 ;
      RECT  155.9 282.5 156.7 281.7 ;
      RECT  153.9 289.5 154.7 288.7 ;
      RECT  157.9 289.5 158.7 288.7 ;
      RECT  154.9 288.0 155.7 287.2 ;
      RECT  156.9 285.2 157.7 284.4 ;
      RECT  159.4 283.8 160.0 283.2 ;
      RECT  152.7 280.7 161.3 280.1 ;
      RECT  152.7 291.1 161.3 290.5 ;
      RECT  164.5 283.3 165.3 282.5 ;
      RECT  162.5 283.3 163.3 282.5 ;
      RECT  164.5 289.5 165.3 288.7 ;
      RECT  162.5 289.5 163.3 288.7 ;
      RECT  162.9 286.4 163.7 285.6 ;
      RECT  164.9 286.3 165.5 285.7 ;
      RECT  161.3 280.7 167.9 280.1 ;
      RECT  161.3 291.1 167.9 290.5 ;
      RECT  154.9 288.0 155.7 287.2 ;
      RECT  156.9 285.2 157.7 284.4 ;
      RECT  164.9 286.3 165.5 285.7 ;
      RECT  152.7 280.7 167.9 280.1 ;
      RECT  152.7 291.1 167.9 290.5 ;
      RECT  155.9 299.1 156.7 299.9 ;
      RECT  153.9 299.1 154.7 299.9 ;
      RECT  157.9 299.1 158.7 299.9 ;
      RECT  155.9 299.1 156.7 299.9 ;
      RECT  153.9 292.1 154.7 292.9 ;
      RECT  157.9 292.1 158.7 292.9 ;
      RECT  154.9 293.6 155.7 294.4 ;
      RECT  156.9 296.4 157.7 297.2 ;
      RECT  159.4 297.8 160.0 298.4 ;
      RECT  152.7 300.9 161.3 301.5 ;
      RECT  152.7 290.5 161.3 291.1 ;
      RECT  164.5 298.3 165.3 299.1 ;
      RECT  162.5 298.3 163.3 299.1 ;
      RECT  164.5 292.1 165.3 292.9 ;
      RECT  162.5 292.1 163.3 292.9 ;
      RECT  162.9 295.2 163.7 296.0 ;
      RECT  164.9 295.3 165.5 295.9 ;
      RECT  161.3 300.9 167.9 301.5 ;
      RECT  161.3 290.5 167.9 291.1 ;
      RECT  154.9 293.6 155.7 294.4 ;
      RECT  156.9 296.4 157.7 297.2 ;
      RECT  164.9 295.3 165.5 295.9 ;
      RECT  152.7 300.9 167.9 301.5 ;
      RECT  152.7 290.5 167.9 291.1 ;
      RECT  155.9 303.3 156.7 302.5 ;
      RECT  153.9 303.3 154.7 302.5 ;
      RECT  157.9 303.3 158.7 302.5 ;
      RECT  155.9 303.3 156.7 302.5 ;
      RECT  153.9 310.3 154.7 309.5 ;
      RECT  157.9 310.3 158.7 309.5 ;
      RECT  154.9 308.8 155.7 308.0 ;
      RECT  156.9 306.0 157.7 305.2 ;
      RECT  159.4 304.6 160.0 304.0 ;
      RECT  152.7 301.5 161.3 300.9 ;
      RECT  152.7 311.9 161.3 311.3 ;
      RECT  164.5 304.1 165.3 303.3 ;
      RECT  162.5 304.1 163.3 303.3 ;
      RECT  164.5 310.3 165.3 309.5 ;
      RECT  162.5 310.3 163.3 309.5 ;
      RECT  162.9 307.2 163.7 306.4 ;
      RECT  164.9 307.1 165.5 306.5 ;
      RECT  161.3 301.5 167.9 300.9 ;
      RECT  161.3 311.9 167.9 311.3 ;
      RECT  154.9 308.8 155.7 308.0 ;
      RECT  156.9 306.0 157.7 305.2 ;
      RECT  164.9 307.1 165.5 306.5 ;
      RECT  152.7 301.5 167.9 300.9 ;
      RECT  152.7 311.9 167.9 311.3 ;
      RECT  155.9 319.9 156.7 320.7 ;
      RECT  153.9 319.9 154.7 320.7 ;
      RECT  157.9 319.9 158.7 320.7 ;
      RECT  155.9 319.9 156.7 320.7 ;
      RECT  153.9 312.9 154.7 313.7 ;
      RECT  157.9 312.9 158.7 313.7 ;
      RECT  154.9 314.4 155.7 315.2 ;
      RECT  156.9 317.2 157.7 318.0 ;
      RECT  159.4 318.6 160.0 319.2 ;
      RECT  152.7 321.7 161.3 322.3 ;
      RECT  152.7 311.3 161.3 311.9 ;
      RECT  164.5 319.1 165.3 319.9 ;
      RECT  162.5 319.1 163.3 319.9 ;
      RECT  164.5 312.9 165.3 313.7 ;
      RECT  162.5 312.9 163.3 313.7 ;
      RECT  162.9 316.0 163.7 316.8 ;
      RECT  164.9 316.1 165.5 316.7 ;
      RECT  161.3 321.7 167.9 322.3 ;
      RECT  161.3 311.3 167.9 311.9 ;
      RECT  154.9 314.4 155.7 315.2 ;
      RECT  156.9 317.2 157.7 318.0 ;
      RECT  164.9 316.1 165.5 316.7 ;
      RECT  152.7 321.7 167.9 322.3 ;
      RECT  152.7 311.3 167.9 311.9 ;
      RECT  155.9 324.1 156.7 323.3 ;
      RECT  153.9 324.1 154.7 323.3 ;
      RECT  157.9 324.1 158.7 323.3 ;
      RECT  155.9 324.1 156.7 323.3 ;
      RECT  153.9 331.1 154.7 330.3 ;
      RECT  157.9 331.1 158.7 330.3 ;
      RECT  154.9 329.6 155.7 328.8 ;
      RECT  156.9 326.8 157.7 326.0 ;
      RECT  159.4 325.4 160.0 324.8 ;
      RECT  152.7 322.3 161.3 321.7 ;
      RECT  152.7 332.7 161.3 332.1 ;
      RECT  164.5 324.9 165.3 324.1 ;
      RECT  162.5 324.9 163.3 324.1 ;
      RECT  164.5 331.1 165.3 330.3 ;
      RECT  162.5 331.1 163.3 330.3 ;
      RECT  162.9 328.0 163.7 327.2 ;
      RECT  164.9 327.9 165.5 327.3 ;
      RECT  161.3 322.3 167.9 321.7 ;
      RECT  161.3 332.7 167.9 332.1 ;
      RECT  154.9 329.6 155.7 328.8 ;
      RECT  156.9 326.8 157.7 326.0 ;
      RECT  164.9 327.9 165.5 327.3 ;
      RECT  152.7 322.3 167.9 321.7 ;
      RECT  152.7 332.7 167.9 332.1 ;
      RECT  155.9 340.7 156.7 341.5 ;
      RECT  153.9 340.7 154.7 341.5 ;
      RECT  157.9 340.7 158.7 341.5 ;
      RECT  155.9 340.7 156.7 341.5 ;
      RECT  153.9 333.7 154.7 334.5 ;
      RECT  157.9 333.7 158.7 334.5 ;
      RECT  154.9 335.2 155.7 336.0 ;
      RECT  156.9 338.0 157.7 338.8 ;
      RECT  159.4 339.4 160.0 340.0 ;
      RECT  152.7 342.5 161.3 343.1 ;
      RECT  152.7 332.1 161.3 332.7 ;
      RECT  164.5 339.9 165.3 340.7 ;
      RECT  162.5 339.9 163.3 340.7 ;
      RECT  164.5 333.7 165.3 334.5 ;
      RECT  162.5 333.7 163.3 334.5 ;
      RECT  162.9 336.8 163.7 337.6 ;
      RECT  164.9 336.9 165.5 337.5 ;
      RECT  161.3 342.5 167.9 343.1 ;
      RECT  161.3 332.1 167.9 332.7 ;
      RECT  154.9 335.2 155.7 336.0 ;
      RECT  156.9 338.0 157.7 338.8 ;
      RECT  164.9 336.9 165.5 337.5 ;
      RECT  152.7 342.5 167.9 343.1 ;
      RECT  152.7 332.1 167.9 332.7 ;
      RECT  155.9 344.9 156.7 344.1 ;
      RECT  153.9 344.9 154.7 344.1 ;
      RECT  157.9 344.9 158.7 344.1 ;
      RECT  155.9 344.9 156.7 344.1 ;
      RECT  153.9 351.9 154.7 351.1 ;
      RECT  157.9 351.9 158.7 351.1 ;
      RECT  154.9 350.4 155.7 349.6 ;
      RECT  156.9 347.6 157.7 346.8 ;
      RECT  159.4 346.2 160.0 345.6 ;
      RECT  152.7 343.1 161.3 342.5 ;
      RECT  152.7 353.5 161.3 352.9 ;
      RECT  164.5 345.7 165.3 344.9 ;
      RECT  162.5 345.7 163.3 344.9 ;
      RECT  164.5 351.9 165.3 351.1 ;
      RECT  162.5 351.9 163.3 351.1 ;
      RECT  162.9 348.8 163.7 348.0 ;
      RECT  164.9 348.7 165.5 348.1 ;
      RECT  161.3 343.1 167.9 342.5 ;
      RECT  161.3 353.5 167.9 352.9 ;
      RECT  154.9 350.4 155.7 349.6 ;
      RECT  156.9 347.6 157.7 346.8 ;
      RECT  164.9 348.7 165.5 348.1 ;
      RECT  152.7 343.1 167.9 342.5 ;
      RECT  152.7 353.5 167.9 352.9 ;
      RECT  154.9 189.6 155.7 190.4 ;
      RECT  154.9 204.0 155.7 204.8 ;
      RECT  154.9 210.4 155.7 211.2 ;
      RECT  154.9 224.8 155.7 225.6 ;
      RECT  154.9 231.2 155.7 232.0 ;
      RECT  154.9 245.6 155.7 246.4 ;
      RECT  154.9 252.0 155.7 252.8 ;
      RECT  154.9 266.4 155.7 267.2 ;
      RECT  154.9 272.8 155.7 273.6 ;
      RECT  154.9 287.2 155.7 288.0 ;
      RECT  154.9 293.6 155.7 294.4 ;
      RECT  154.9 308.0 155.7 308.8 ;
      RECT  154.9 314.4 155.7 315.2 ;
      RECT  154.9 328.8 155.7 329.6 ;
      RECT  154.9 335.2 155.7 336.0 ;
      RECT  154.9 349.6 155.7 350.4 ;
      RECT  164.9 191.3 165.5 191.9 ;
      RECT  164.9 202.5 165.5 203.1 ;
      RECT  164.9 212.1 165.5 212.7 ;
      RECT  164.9 223.3 165.5 223.9 ;
      RECT  164.9 232.9 165.5 233.5 ;
      RECT  164.9 244.1 165.5 244.7 ;
      RECT  164.9 253.7 165.5 254.3 ;
      RECT  164.9 264.9 165.5 265.5 ;
      RECT  164.9 274.5 165.5 275.1 ;
      RECT  164.9 285.7 165.5 286.3 ;
      RECT  164.9 295.3 165.5 295.9 ;
      RECT  164.9 306.5 165.5 307.1 ;
      RECT  164.9 316.1 165.5 316.7 ;
      RECT  164.9 327.3 165.5 327.9 ;
      RECT  164.9 336.9 165.5 337.5 ;
      RECT  164.9 348.1 165.5 348.7 ;
      RECT  164.9 191.3 165.5 191.9 ;
      RECT  164.9 202.5 165.5 203.1 ;
      RECT  164.9 212.1 165.5 212.7 ;
      RECT  164.9 223.3 165.5 223.9 ;
      RECT  164.9 232.9 165.5 233.5 ;
      RECT  164.9 244.1 165.5 244.7 ;
      RECT  164.9 253.7 165.5 254.3 ;
      RECT  164.9 264.9 165.5 265.5 ;
      RECT  164.9 274.5 165.5 275.1 ;
      RECT  164.9 285.7 165.5 286.3 ;
      RECT  164.9 295.3 165.5 295.9 ;
      RECT  164.9 306.5 165.5 307.1 ;
      RECT  164.9 316.1 165.5 316.7 ;
      RECT  164.9 327.3 165.5 327.9 ;
      RECT  164.9 336.9 165.5 337.5 ;
      RECT  164.9 348.1 165.5 348.7 ;
      RECT  16.4 10.8 17.2 11.0 ;
      RECT  3.6 4.0 4.4 8.8 ;
      RECT  12.4 17.0 13.0 17.6 ;
      RECT  10.2 16.4 13.8 17.0 ;
      RECT  3.6 12.6 9.2 12.8 ;
      RECT  4.4 9.6 15.4 10.2 ;
      RECT  21.2 13.0 22.0 21.6 ;
      RECT  12.4 6.0 13.0 6.6 ;
      RECT  8.0 4.0 8.8 5.4 ;
      RECT  10.2 16.2 11.0 16.4 ;
      RECT  16.4 16.8 17.2 17.6 ;
      RECT  12.8 13.6 13.4 14.8 ;
      RECT  6.8 17.6 8.8 18.2 ;
      RECT  14.0 3.4 14.8 6.0 ;
      RECT  10.2 6.6 13.0 7.2 ;
      RECT  6.8 5.4 8.8 6.0 ;
      RECT  21.2 9.0 22.0 12.4 ;
      RECT  16.6 17.6 17.8 21.6 ;
      RECT  5.2 13.8 6.0 22.2 ;
      RECT  6.8 14.2 12.2 14.8 ;
      RECT  14.8 10.2 15.4 13.4 ;
      RECT  2.4 22.2 24.2 23.4 ;
      RECT  17.8 12.4 22.0 13.0 ;
      RECT  19.6 13.6 20.4 22.2 ;
      RECT  22.8 3.4 23.6 4.8 ;
      RECT  16.6 14.0 17.2 15.0 ;
      RECT  14.8 13.4 17.2 14.0 ;
      RECT  3.6 13.2 4.4 21.6 ;
      RECT  16.4 5.4 17.8 6.0 ;
      RECT  12.8 14.8 15.0 15.4 ;
      RECT  8.0 18.2 8.8 21.6 ;
      RECT  5.8 11.4 10.8 12.0 ;
      RECT  22.8 20.6 23.6 22.2 ;
      RECT  16.4 11.0 20.2 11.6 ;
      RECT  16.4 6.0 17.2 6.8 ;
      RECT  2.4 2.2 24.2 3.4 ;
      RECT  10.0 12.0 10.8 12.2 ;
      RECT  7.4 10.2 8.2 10.4 ;
      RECT  13.0 16.2 13.8 16.4 ;
      RECT  21.2 4.0 22.0 8.4 ;
      RECT  4.4 9.4 6.0 9.6 ;
      RECT  6.8 16.8 7.6 17.6 ;
      RECT  12.4 4.0 13.2 6.0 ;
      RECT  5.8 11.2 6.6 11.4 ;
      RECT  6.8 14.8 7.6 15.0 ;
      RECT  18.2 8.2 19.0 8.4 ;
      RECT  8.4 6.6 9.2 7.4 ;
      RECT  19.6 3.4 20.4 7.8 ;
      RECT  14.2 14.6 15.0 14.8 ;
      RECT  10.6 3.4 11.6 6.0 ;
      RECT  8.6 7.4 9.2 9.6 ;
      RECT  14.0 17.6 14.8 22.2 ;
      RECT  10.8 17.6 11.6 22.2 ;
      RECT  14.2 9.4 15.0 9.6 ;
      RECT  8.6 13.2 13.4 13.6 ;
      RECT  3.6 12.8 9.4 13.0 ;
      RECT  12.4 17.6 13.2 21.6 ;
      RECT  19.4 11.6 20.2 11.8 ;
      RECT  3.6 13.0 13.4 13.2 ;
      RECT  11.4 14.8 12.2 15.0 ;
      RECT  16.6 4.0 17.8 5.4 ;
      RECT  10.2 7.2 11.0 7.4 ;
      RECT  16.6 15.0 18.0 15.8 ;
      RECT  17.8 12.2 18.6 12.4 ;
      RECT  6.8 6.0 7.6 6.8 ;
      RECT  5.2 3.4 6.0 8.0 ;
      RECT  18.2 8.4 22.0 9.0 ;
      RECT  29.8 19.9 30.6 20.7 ;
      RECT  27.8 19.9 28.6 20.7 ;
      RECT  29.8 4.1 30.6 4.9 ;
      RECT  27.8 4.1 28.6 4.9 ;
      RECT  28.2 12.0 29.0 12.8 ;
      RECT  30.2 12.1 30.8 12.7 ;
      RECT  26.6 22.5 33.2 23.1 ;
      RECT  26.6 2.5 33.2 3.1 ;
      RECT  36.4 18.3 37.2 19.1 ;
      RECT  34.4 18.3 35.2 19.1 ;
      RECT  36.4 4.9 37.2 5.7 ;
      RECT  34.4 4.9 35.2 5.7 ;
      RECT  34.8 11.6 35.6 12.4 ;
      RECT  36.8 11.7 37.4 12.3 ;
      RECT  33.2 22.5 39.8 23.1 ;
      RECT  33.2 2.5 39.8 3.1 ;
      RECT  2.4 22.2 39.8 23.4 ;
      RECT  2.4 2.2 39.8 3.4 ;
      RECT  16.4 34.8 17.2 34.6 ;
      RECT  3.6 41.6 4.4 36.8 ;
      RECT  12.4 28.6 13.0 28.0 ;
      RECT  10.2 29.2 13.8 28.6 ;
      RECT  3.6 33.0 9.2 32.8 ;
      RECT  4.4 36.0 15.4 35.4 ;
      RECT  21.2 32.6 22.0 24.0 ;
      RECT  12.4 39.6 13.0 39.0 ;
      RECT  8.0 41.6 8.8 40.2 ;
      RECT  10.2 29.4 11.0 29.2 ;
      RECT  16.4 28.8 17.2 28.0 ;
      RECT  12.8 32.0 13.4 30.8 ;
      RECT  6.8 28.0 8.8 27.4 ;
      RECT  14.0 42.2 14.8 39.6 ;
      RECT  10.2 39.0 13.0 38.4 ;
      RECT  6.8 40.2 8.8 39.6 ;
      RECT  21.2 36.6 22.0 33.2 ;
      RECT  16.6 28.0 17.8 24.0 ;
      RECT  5.2 31.8 6.0 23.4 ;
      RECT  6.8 31.4 12.2 30.8 ;
      RECT  14.8 35.4 15.4 32.2 ;
      RECT  2.4 23.4 24.2 22.2 ;
      RECT  17.8 33.2 22.0 32.6 ;
      RECT  19.6 32.0 20.4 23.4 ;
      RECT  22.8 42.2 23.6 40.8 ;
      RECT  16.6 31.6 17.2 30.6 ;
      RECT  14.8 32.2 17.2 31.6 ;
      RECT  3.6 32.4 4.4 24.0 ;
      RECT  16.4 40.2 17.8 39.6 ;
      RECT  12.8 30.8 15.0 30.2 ;
      RECT  8.0 27.4 8.8 24.0 ;
      RECT  5.8 34.2 10.8 33.6 ;
      RECT  22.8 25.0 23.6 23.4 ;
      RECT  16.4 34.6 20.2 34.0 ;
      RECT  16.4 39.6 17.2 38.8 ;
      RECT  2.4 43.4 24.2 42.2 ;
      RECT  10.0 33.6 10.8 33.4 ;
      RECT  7.4 35.4 8.2 35.2 ;
      RECT  13.0 29.4 13.8 29.2 ;
      RECT  21.2 41.6 22.0 37.2 ;
      RECT  4.4 36.2 6.0 36.0 ;
      RECT  6.8 28.8 7.6 28.0 ;
      RECT  12.4 41.6 13.2 39.6 ;
      RECT  5.8 34.4 6.6 34.2 ;
      RECT  6.8 30.8 7.6 30.6 ;
      RECT  18.2 37.4 19.0 37.2 ;
      RECT  8.4 39.0 9.2 38.2 ;
      RECT  19.6 42.2 20.4 37.8 ;
      RECT  14.2 31.0 15.0 30.8 ;
      RECT  10.6 42.2 11.6 39.6 ;
      RECT  8.6 38.2 9.2 36.0 ;
      RECT  14.0 28.0 14.8 23.4 ;
      RECT  10.8 28.0 11.6 23.4 ;
      RECT  14.2 36.2 15.0 36.0 ;
      RECT  8.6 32.4 13.4 32.0 ;
      RECT  3.6 32.8 9.4 32.6 ;
      RECT  12.4 28.0 13.2 24.0 ;
      RECT  19.4 34.0 20.2 33.8 ;
      RECT  3.6 32.6 13.4 32.4 ;
      RECT  11.4 30.8 12.2 30.6 ;
      RECT  16.6 41.6 17.8 40.2 ;
      RECT  10.2 38.4 11.0 38.2 ;
      RECT  16.6 30.6 18.0 29.8 ;
      RECT  17.8 33.4 18.6 33.2 ;
      RECT  6.8 39.6 7.6 38.8 ;
      RECT  5.2 42.2 6.0 37.6 ;
      RECT  18.2 37.2 22.0 36.6 ;
      RECT  29.8 25.7 30.6 24.9 ;
      RECT  27.8 25.7 28.6 24.9 ;
      RECT  29.8 41.5 30.6 40.7 ;
      RECT  27.8 41.5 28.6 40.7 ;
      RECT  28.2 33.6 29.0 32.8 ;
      RECT  30.2 33.5 30.8 32.9 ;
      RECT  26.6 23.1 33.2 22.5 ;
      RECT  26.6 43.1 33.2 42.5 ;
      RECT  36.4 27.3 37.2 26.5 ;
      RECT  34.4 27.3 35.2 26.5 ;
      RECT  36.4 40.7 37.2 39.9 ;
      RECT  34.4 40.7 35.2 39.9 ;
      RECT  34.8 34.0 35.6 33.2 ;
      RECT  36.8 33.9 37.4 33.3 ;
      RECT  33.2 23.1 39.8 22.5 ;
      RECT  33.2 43.1 39.8 42.5 ;
      RECT  2.4 23.4 39.8 22.2 ;
      RECT  2.4 43.4 39.8 42.2 ;
      RECT  55.6 20.7 56.4 21.5 ;
      RECT  53.6 20.7 54.4 21.5 ;
      RECT  55.6 3.7 56.4 4.5 ;
      RECT  53.6 3.7 54.4 4.5 ;
      RECT  54.0 12.2 54.8 13.0 ;
      RECT  56.0 12.3 56.6 12.9 ;
      RECT  52.4 22.5 59.0 23.1 ;
      RECT  52.4 2.5 59.0 3.1 ;
      RECT  62.2 19.9 63.0 20.7 ;
      RECT  60.2 19.9 61.0 20.7 ;
      RECT  62.2 4.1 63.0 4.9 ;
      RECT  60.2 4.1 61.0 4.9 ;
      RECT  60.6 12.0 61.4 12.8 ;
      RECT  62.6 12.1 63.2 12.7 ;
      RECT  59.0 22.5 64.2 23.1 ;
      RECT  59.0 2.5 64.2 3.1 ;
      RECT  67.4 17.5 68.2 18.3 ;
      RECT  65.4 17.5 66.2 18.3 ;
      RECT  67.4 5.3 68.2 6.1 ;
      RECT  65.4 5.3 66.2 6.1 ;
      RECT  65.8 11.4 66.6 12.2 ;
      RECT  67.8 11.5 68.4 12.1 ;
      RECT  64.2 22.5 69.4 23.1 ;
      RECT  64.2 2.5 69.4 3.1 ;
      RECT  72.5 16.3 76.5 16.9 ;
      RECT  70.6 17.5 71.4 18.3 ;
      RECT  74.0 17.5 74.8 18.3 ;
      RECT  72.5 6.7 76.5 7.3 ;
      RECT  70.6 5.3 71.4 6.1 ;
      RECT  74.0 5.3 74.8 6.1 ;
      RECT  71.0 11.4 71.8 12.2 ;
      RECT  74.5 11.5 75.1 12.1 ;
      RECT  69.4 22.5 78.0 23.1 ;
      RECT  69.4 2.5 78.0 3.1 ;
      RECT  54.0 12.2 54.8 13.0 ;
      RECT  74.5 11.5 75.1 12.1 ;
      RECT  52.4 22.5 78.0 23.1 ;
      RECT  52.4 2.5 78.0 3.1 ;
      RECT  55.6 24.9 56.4 24.1 ;
      RECT  53.6 24.9 54.4 24.1 ;
      RECT  55.6 41.9 56.4 41.1 ;
      RECT  53.6 41.9 54.4 41.1 ;
      RECT  54.0 33.4 54.8 32.6 ;
      RECT  56.0 33.3 56.6 32.7 ;
      RECT  52.4 23.1 59.0 22.5 ;
      RECT  52.4 43.1 59.0 42.5 ;
      RECT  62.2 24.9 63.0 24.1 ;
      RECT  60.2 24.9 61.0 24.1 ;
      RECT  64.2 24.9 65.0 24.1 ;
      RECT  62.2 24.9 63.0 24.1 ;
      RECT  60.2 41.5 61.0 40.7 ;
      RECT  64.2 41.5 65.0 40.7 ;
      RECT  61.2 40.0 62.0 39.2 ;
      RECT  63.2 37.2 64.0 36.4 ;
      RECT  65.7 26.2 66.3 25.6 ;
      RECT  59.0 23.1 66.6 22.5 ;
      RECT  59.0 43.1 66.6 42.5 ;
      RECT  69.7 28.5 73.7 27.9 ;
      RECT  71.2 27.3 72.0 26.5 ;
      RECT  67.8 27.3 68.6 26.5 ;
      RECT  69.7 39.3 73.7 38.7 ;
      RECT  71.2 40.7 72.0 39.9 ;
      RECT  67.8 40.7 68.6 39.9 ;
      RECT  68.2 34.0 69.0 33.2 ;
      RECT  71.7 33.9 72.3 33.3 ;
      RECT  66.6 23.1 76.4 22.5 ;
      RECT  66.6 43.1 76.4 42.5 ;
      RECT  68.2 34.0 69.0 33.2 ;
      RECT  71.7 33.9 72.3 33.3 ;
      RECT  66.6 23.1 76.4 22.5 ;
      RECT  66.6 43.1 76.4 42.5 ;
      RECT  61.2 40.0 62.0 39.2 ;
      RECT  63.2 37.2 64.0 36.4 ;
      RECT  71.7 33.9 72.3 33.3 ;
      RECT  59.0 23.1 76.4 22.5 ;
      RECT  59.0 43.1 76.4 42.5 ;
      RECT  55.6 60.7 56.4 61.5 ;
      RECT  53.6 60.7 54.4 61.5 ;
      RECT  57.6 60.7 58.4 61.5 ;
      RECT  55.6 60.7 56.4 61.5 ;
      RECT  53.6 44.1 54.4 44.9 ;
      RECT  57.6 44.1 58.4 44.9 ;
      RECT  54.6 45.6 55.4 46.4 ;
      RECT  56.6 48.4 57.4 49.2 ;
      RECT  59.1 59.4 59.7 60.0 ;
      RECT  52.4 62.5 60.0 63.1 ;
      RECT  52.4 42.5 60.0 43.1 ;
      RECT  63.1 57.1 67.1 57.7 ;
      RECT  64.6 58.3 65.4 59.1 ;
      RECT  61.2 58.3 62.0 59.1 ;
      RECT  63.1 46.3 67.1 46.9 ;
      RECT  64.6 44.9 65.4 45.7 ;
      RECT  61.2 44.9 62.0 45.7 ;
      RECT  61.6 51.6 62.4 52.4 ;
      RECT  65.1 51.7 65.7 52.3 ;
      RECT  60.0 62.5 69.8 63.1 ;
      RECT  60.0 42.5 69.8 43.1 ;
      RECT  61.6 51.6 62.4 52.4 ;
      RECT  65.1 51.7 65.7 52.3 ;
      RECT  60.0 62.5 69.8 63.1 ;
      RECT  60.0 42.5 69.8 43.1 ;
      RECT  54.6 45.6 55.4 46.4 ;
      RECT  56.6 48.4 57.4 49.2 ;
      RECT  65.1 51.7 65.7 52.3 ;
      RECT  52.4 62.5 69.8 63.1 ;
      RECT  52.4 42.5 69.8 43.1 ;
      RECT  55.6 64.9 56.4 64.1 ;
      RECT  53.6 64.9 54.4 64.1 ;
      RECT  55.6 81.9 56.4 81.1 ;
      RECT  53.6 81.9 54.4 81.1 ;
      RECT  54.0 73.4 54.8 72.6 ;
      RECT  56.0 73.3 56.6 72.7 ;
      RECT  52.4 63.1 59.0 62.5 ;
      RECT  52.4 83.1 59.0 82.5 ;
      RECT  62.2 64.9 63.0 64.1 ;
      RECT  60.2 64.9 61.0 64.1 ;
      RECT  62.2 81.9 63.0 81.1 ;
      RECT  60.2 81.9 61.0 81.1 ;
      RECT  60.6 73.4 61.4 72.6 ;
      RECT  62.6 73.3 63.2 72.7 ;
      RECT  59.0 63.1 64.2 62.5 ;
      RECT  59.0 83.1 64.2 82.5 ;
      RECT  67.4 65.7 68.2 64.9 ;
      RECT  65.4 65.7 66.2 64.9 ;
      RECT  67.4 81.5 68.2 80.7 ;
      RECT  65.4 81.5 66.2 80.7 ;
      RECT  65.8 73.6 66.6 72.8 ;
      RECT  67.8 73.5 68.4 72.9 ;
      RECT  64.2 63.1 69.4 62.5 ;
      RECT  64.2 83.1 69.4 82.5 ;
      RECT  72.6 68.1 73.4 67.3 ;
      RECT  70.6 68.1 71.4 67.3 ;
      RECT  72.6 80.3 73.4 79.5 ;
      RECT  70.6 80.3 71.4 79.5 ;
      RECT  71.0 74.2 71.8 73.4 ;
      RECT  73.0 74.1 73.6 73.5 ;
      RECT  69.4 63.1 74.6 62.5 ;
      RECT  69.4 83.1 74.6 82.5 ;
      RECT  54.0 73.4 54.8 72.6 ;
      RECT  73.0 74.1 73.6 73.5 ;
      RECT  52.4 63.1 74.6 62.5 ;
      RECT  52.4 83.1 74.6 82.5 ;
      RECT  55.6 140.7 56.4 141.5 ;
      RECT  53.6 140.7 54.4 141.5 ;
      RECT  55.6 123.7 56.4 124.5 ;
      RECT  53.6 123.7 54.4 124.5 ;
      RECT  54.0 132.2 54.8 133.0 ;
      RECT  56.0 132.3 56.6 132.9 ;
      RECT  52.4 142.5 59.0 143.1 ;
      RECT  52.4 122.5 59.0 123.1 ;
      RECT  55.6 100.7 56.4 101.5 ;
      RECT  53.6 100.7 54.4 101.5 ;
      RECT  57.6 100.7 58.4 101.5 ;
      RECT  55.6 100.7 56.4 101.5 ;
      RECT  59.6 100.7 60.4 101.5 ;
      RECT  57.6 100.7 58.4 101.5 ;
      RECT  53.6 84.1 54.4 84.9 ;
      RECT  59.6 84.1 60.4 84.9 ;
      RECT  54.2 85.6 55.0 86.4 ;
      RECT  56.6 87.0 57.4 87.8 ;
      RECT  59.0 88.4 59.8 89.2 ;
      RECT  61.1 99.5 61.7 100.1 ;
      RECT  52.4 102.5 62.0 103.1 ;
      RECT  52.4 82.5 62.0 83.1 ;
      RECT  65.0 97.5 65.8 98.3 ;
      RECT  63.2 97.5 64.0 98.3 ;
      RECT  66.8 97.5 67.6 98.3 ;
      RECT  65.0 85.3 65.8 86.1 ;
      RECT  63.2 85.3 64.0 86.1 ;
      RECT  66.8 85.3 67.6 86.1 ;
      RECT  63.6 91.4 64.4 92.2 ;
      RECT  65.4 91.5 66.0 92.1 ;
      RECT  62.0 102.5 70.2 103.1 ;
      RECT  62.0 82.5 70.2 83.1 ;
      RECT  63.6 91.4 64.4 92.2 ;
      RECT  65.4 91.5 66.0 92.1 ;
      RECT  62.0 102.5 70.2 103.1 ;
      RECT  62.0 82.5 70.2 83.1 ;
      RECT  54.2 85.6 55.0 86.4 ;
      RECT  56.6 87.0 57.4 87.8 ;
      RECT  59.0 88.4 59.8 89.2 ;
      RECT  65.4 91.5 66.0 92.1 ;
      RECT  52.4 102.5 70.2 103.1 ;
      RECT  52.4 82.5 70.2 83.1 ;
      RECT  55.6 144.9 56.4 144.1 ;
      RECT  53.6 144.9 54.4 144.1 ;
      RECT  57.6 144.9 58.4 144.1 ;
      RECT  55.6 144.9 56.4 144.1 ;
      RECT  59.6 144.9 60.4 144.1 ;
      RECT  57.6 144.9 58.4 144.1 ;
      RECT  53.6 161.5 54.4 160.7 ;
      RECT  59.6 161.5 60.4 160.7 ;
      RECT  54.2 160.0 55.0 159.2 ;
      RECT  56.6 158.6 57.4 157.8 ;
      RECT  59.0 157.2 59.8 156.4 ;
      RECT  61.1 146.1 61.7 145.5 ;
      RECT  52.4 143.1 62.0 142.5 ;
      RECT  52.4 163.1 62.0 162.5 ;
      RECT  65.2 145.7 66.0 144.9 ;
      RECT  63.2 145.7 64.0 144.9 ;
      RECT  65.2 161.5 66.0 160.7 ;
      RECT  63.2 161.5 64.0 160.7 ;
      RECT  63.6 153.6 64.4 152.8 ;
      RECT  65.6 153.5 66.2 152.9 ;
      RECT  62.0 143.1 68.6 142.5 ;
      RECT  62.0 163.1 68.6 162.5 ;
      RECT  63.6 153.6 64.4 152.8 ;
      RECT  65.6 153.5 66.2 152.9 ;
      RECT  62.0 143.1 68.6 142.5 ;
      RECT  62.0 163.1 68.6 162.5 ;
      RECT  54.2 160.0 55.0 159.2 ;
      RECT  56.6 158.6 57.4 157.8 ;
      RECT  59.0 157.2 59.8 156.4 ;
      RECT  65.6 153.5 66.2 152.9 ;
      RECT  52.4 143.1 68.6 142.5 ;
      RECT  52.4 163.1 68.6 162.5 ;
      RECT  32.2 183.1 31.4 183.9 ;
      RECT  34.2 183.1 33.4 183.9 ;
      RECT  32.2 166.5 31.4 167.3 ;
      RECT  34.2 166.5 33.4 167.3 ;
      RECT  33.8 174.8 33.0 175.6 ;
      RECT  31.8 174.9 31.2 175.5 ;
      RECT  35.4 184.9 28.8 185.5 ;
      RECT  35.4 165.3 28.8 165.9 ;
      RECT  25.6 183.1 24.8 183.9 ;
      RECT  27.6 183.1 26.8 183.9 ;
      RECT  25.6 166.5 24.8 167.3 ;
      RECT  27.6 166.5 26.8 167.3 ;
      RECT  27.2 174.8 26.4 175.6 ;
      RECT  25.2 174.9 24.6 175.5 ;
      RECT  28.8 184.9 22.2 185.5 ;
      RECT  28.8 165.3 22.2 165.9 ;
      RECT  19.0 183.1 18.2 183.9 ;
      RECT  21.0 183.1 20.2 183.9 ;
      RECT  19.0 166.5 18.2 167.3 ;
      RECT  21.0 166.5 20.2 167.3 ;
      RECT  20.6 174.8 19.8 175.6 ;
      RECT  18.6 174.9 18.0 175.5 ;
      RECT  22.2 184.9 15.6 185.5 ;
      RECT  22.2 165.3 15.6 165.9 ;
      RECT  12.4 183.1 11.6 183.9 ;
      RECT  14.4 183.1 13.6 183.9 ;
      RECT  12.4 166.5 11.6 167.3 ;
      RECT  14.4 166.5 13.6 167.3 ;
      RECT  14.0 174.8 13.2 175.6 ;
      RECT  12.0 174.9 11.4 175.5 ;
      RECT  15.6 184.9 9.0 185.5 ;
      RECT  15.6 165.3 9.0 165.9 ;
      RECT  5.8 183.1 5.0 183.9 ;
      RECT  7.8 183.1 7.0 183.9 ;
      RECT  5.8 166.5 5.0 167.3 ;
      RECT  7.8 166.5 7.0 167.3 ;
      RECT  7.4 174.8 6.6 175.6 ;
      RECT  5.4 174.9 4.8 175.5 ;
      RECT  9.0 184.9 2.4 185.5 ;
      RECT  9.0 165.3 2.4 165.9 ;
      RECT  32.2 187.3 31.4 186.5 ;
      RECT  34.2 187.3 33.4 186.5 ;
      RECT  32.2 203.9 31.4 203.1 ;
      RECT  34.2 203.9 33.4 203.1 ;
      RECT  33.8 195.6 33.0 194.8 ;
      RECT  31.8 195.5 31.2 194.9 ;
      RECT  35.4 185.5 28.8 184.9 ;
      RECT  35.4 205.1 28.8 204.5 ;
      RECT  25.6 187.3 24.8 186.5 ;
      RECT  27.6 187.3 26.8 186.5 ;
      RECT  25.6 203.9 24.8 203.1 ;
      RECT  27.6 203.9 26.8 203.1 ;
      RECT  27.2 195.6 26.4 194.8 ;
      RECT  25.2 195.5 24.6 194.9 ;
      RECT  28.8 185.5 22.2 184.9 ;
      RECT  28.8 205.1 22.2 204.5 ;
      RECT  19.0 187.3 18.2 186.5 ;
      RECT  21.0 187.3 20.2 186.5 ;
      RECT  19.0 203.9 18.2 203.1 ;
      RECT  21.0 203.9 20.2 203.1 ;
      RECT  20.6 195.6 19.8 194.8 ;
      RECT  18.6 195.5 18.0 194.9 ;
      RECT  22.2 185.5 15.6 184.9 ;
      RECT  22.2 205.1 15.6 204.5 ;
      RECT  12.4 187.3 11.6 186.5 ;
      RECT  14.4 187.3 13.6 186.5 ;
      RECT  12.4 203.9 11.6 203.1 ;
      RECT  14.4 203.9 13.6 203.1 ;
      RECT  14.0 195.6 13.2 194.8 ;
      RECT  12.0 195.5 11.4 194.9 ;
      RECT  15.6 185.5 9.0 184.9 ;
      RECT  15.6 205.1 9.0 204.5 ;
      RECT  5.8 187.3 5.0 186.5 ;
      RECT  7.8 187.3 7.0 186.5 ;
      RECT  5.8 203.9 5.0 203.1 ;
      RECT  7.8 203.9 7.0 203.1 ;
      RECT  7.4 195.6 6.6 194.8 ;
      RECT  5.4 195.5 4.8 194.9 ;
      RECT  9.0 185.5 2.4 184.9 ;
      RECT  9.0 205.1 2.4 204.5 ;
      RECT  32.2 222.3 31.4 223.1 ;
      RECT  34.2 222.3 33.4 223.1 ;
      RECT  32.2 205.7 31.4 206.5 ;
      RECT  34.2 205.7 33.4 206.5 ;
      RECT  33.8 214.0 33.0 214.8 ;
      RECT  31.8 214.1 31.2 214.7 ;
      RECT  35.4 224.1 28.8 224.7 ;
      RECT  35.4 204.5 28.8 205.1 ;
      RECT  25.6 222.3 24.8 223.1 ;
      RECT  27.6 222.3 26.8 223.1 ;
      RECT  25.6 205.7 24.8 206.5 ;
      RECT  27.6 205.7 26.8 206.5 ;
      RECT  27.2 214.0 26.4 214.8 ;
      RECT  25.2 214.1 24.6 214.7 ;
      RECT  28.8 224.1 22.2 224.7 ;
      RECT  28.8 204.5 22.2 205.1 ;
      RECT  19.0 222.3 18.2 223.1 ;
      RECT  21.0 222.3 20.2 223.1 ;
      RECT  19.0 205.7 18.2 206.5 ;
      RECT  21.0 205.7 20.2 206.5 ;
      RECT  20.6 214.0 19.8 214.8 ;
      RECT  18.6 214.1 18.0 214.7 ;
      RECT  22.2 224.1 15.6 224.7 ;
      RECT  22.2 204.5 15.6 205.1 ;
      RECT  12.4 222.3 11.6 223.1 ;
      RECT  14.4 222.3 13.6 223.1 ;
      RECT  12.4 205.7 11.6 206.5 ;
      RECT  14.4 205.7 13.6 206.5 ;
      RECT  14.0 214.0 13.2 214.8 ;
      RECT  12.0 214.1 11.4 214.7 ;
      RECT  15.6 224.1 9.0 224.7 ;
      RECT  15.6 204.5 9.0 205.1 ;
      RECT  5.8 222.3 5.0 223.1 ;
      RECT  7.8 222.3 7.0 223.1 ;
      RECT  5.8 205.7 5.0 206.5 ;
      RECT  7.8 205.7 7.0 206.5 ;
      RECT  7.4 214.0 6.6 214.8 ;
      RECT  5.4 214.1 4.8 214.7 ;
      RECT  9.0 224.1 2.4 224.7 ;
      RECT  9.0 204.5 2.4 205.1 ;
      RECT  32.2 226.5 31.4 225.7 ;
      RECT  34.2 226.5 33.4 225.7 ;
      RECT  32.2 243.1 31.4 242.3 ;
      RECT  34.2 243.1 33.4 242.3 ;
      RECT  33.8 234.8 33.0 234.0 ;
      RECT  31.8 234.7 31.2 234.1 ;
      RECT  35.4 224.7 28.8 224.1 ;
      RECT  35.4 244.3 28.8 243.7 ;
      RECT  25.6 226.5 24.8 225.7 ;
      RECT  27.6 226.5 26.8 225.7 ;
      RECT  25.6 243.1 24.8 242.3 ;
      RECT  27.6 243.1 26.8 242.3 ;
      RECT  27.2 234.8 26.4 234.0 ;
      RECT  25.2 234.7 24.6 234.1 ;
      RECT  28.8 224.7 22.2 224.1 ;
      RECT  28.8 244.3 22.2 243.7 ;
      RECT  19.0 226.5 18.2 225.7 ;
      RECT  21.0 226.5 20.2 225.7 ;
      RECT  19.0 243.1 18.2 242.3 ;
      RECT  21.0 243.1 20.2 242.3 ;
      RECT  20.6 234.8 19.8 234.0 ;
      RECT  18.6 234.7 18.0 234.1 ;
      RECT  22.2 224.7 15.6 224.1 ;
      RECT  22.2 244.3 15.6 243.7 ;
      RECT  12.4 226.5 11.6 225.7 ;
      RECT  14.4 226.5 13.6 225.7 ;
      RECT  12.4 243.1 11.6 242.3 ;
      RECT  14.4 243.1 13.6 242.3 ;
      RECT  14.0 234.8 13.2 234.0 ;
      RECT  12.0 234.7 11.4 234.1 ;
      RECT  15.6 224.7 9.0 224.1 ;
      RECT  15.6 244.3 9.0 243.7 ;
      RECT  5.8 226.5 5.0 225.7 ;
      RECT  7.8 226.5 7.0 225.7 ;
      RECT  5.8 243.1 5.0 242.3 ;
      RECT  7.8 243.1 7.0 242.3 ;
      RECT  7.4 234.8 6.6 234.0 ;
      RECT  5.4 234.7 4.8 234.1 ;
      RECT  9.0 224.7 2.4 224.1 ;
      RECT  9.0 244.3 2.4 243.7 ;
      RECT  32.2 261.5 31.4 262.3 ;
      RECT  34.2 261.5 33.4 262.3 ;
      RECT  32.2 244.9 31.4 245.7 ;
      RECT  34.2 244.9 33.4 245.7 ;
      RECT  33.8 253.2 33.0 254.0 ;
      RECT  31.8 253.3 31.2 253.9 ;
      RECT  35.4 263.3 28.8 263.9 ;
      RECT  35.4 243.7 28.8 244.3 ;
      RECT  25.6 261.5 24.8 262.3 ;
      RECT  27.6 261.5 26.8 262.3 ;
      RECT  25.6 244.9 24.8 245.7 ;
      RECT  27.6 244.9 26.8 245.7 ;
      RECT  27.2 253.2 26.4 254.0 ;
      RECT  25.2 253.3 24.6 253.9 ;
      RECT  28.8 263.3 22.2 263.9 ;
      RECT  28.8 243.7 22.2 244.3 ;
      RECT  19.0 261.5 18.2 262.3 ;
      RECT  21.0 261.5 20.2 262.3 ;
      RECT  19.0 244.9 18.2 245.7 ;
      RECT  21.0 244.9 20.2 245.7 ;
      RECT  20.6 253.2 19.8 254.0 ;
      RECT  18.6 253.3 18.0 253.9 ;
      RECT  22.2 263.3 15.6 263.9 ;
      RECT  22.2 243.7 15.6 244.3 ;
      RECT  12.4 261.5 11.6 262.3 ;
      RECT  14.4 261.5 13.6 262.3 ;
      RECT  12.4 244.9 11.6 245.7 ;
      RECT  14.4 244.9 13.6 245.7 ;
      RECT  14.0 253.2 13.2 254.0 ;
      RECT  12.0 253.3 11.4 253.9 ;
      RECT  15.6 263.3 9.0 263.9 ;
      RECT  15.6 243.7 9.0 244.3 ;
      RECT  5.8 261.5 5.0 262.3 ;
      RECT  7.8 261.5 7.0 262.3 ;
      RECT  5.8 244.9 5.0 245.7 ;
      RECT  7.8 244.9 7.0 245.7 ;
      RECT  7.4 253.2 6.6 254.0 ;
      RECT  5.4 253.3 4.8 253.9 ;
      RECT  9.0 263.3 2.4 263.9 ;
      RECT  9.0 243.7 2.4 244.3 ;
      RECT  32.2 265.7 31.4 264.9 ;
      RECT  34.2 265.7 33.4 264.9 ;
      RECT  32.2 282.3 31.4 281.5 ;
      RECT  34.2 282.3 33.4 281.5 ;
      RECT  33.8 274.0 33.0 273.2 ;
      RECT  31.8 273.9 31.2 273.3 ;
      RECT  35.4 263.9 28.8 263.3 ;
      RECT  35.4 283.5 28.8 282.9 ;
      RECT  25.6 265.7 24.8 264.9 ;
      RECT  27.6 265.7 26.8 264.9 ;
      RECT  25.6 282.3 24.8 281.5 ;
      RECT  27.6 282.3 26.8 281.5 ;
      RECT  27.2 274.0 26.4 273.2 ;
      RECT  25.2 273.9 24.6 273.3 ;
      RECT  28.8 263.9 22.2 263.3 ;
      RECT  28.8 283.5 22.2 282.9 ;
      RECT  19.0 265.7 18.2 264.9 ;
      RECT  21.0 265.7 20.2 264.9 ;
      RECT  19.0 282.3 18.2 281.5 ;
      RECT  21.0 282.3 20.2 281.5 ;
      RECT  20.6 274.0 19.8 273.2 ;
      RECT  18.6 273.9 18.0 273.3 ;
      RECT  22.2 263.9 15.6 263.3 ;
      RECT  22.2 283.5 15.6 282.9 ;
      RECT  12.4 265.7 11.6 264.9 ;
      RECT  14.4 265.7 13.6 264.9 ;
      RECT  12.4 282.3 11.6 281.5 ;
      RECT  14.4 282.3 13.6 281.5 ;
      RECT  14.0 274.0 13.2 273.2 ;
      RECT  12.0 273.9 11.4 273.3 ;
      RECT  15.6 263.9 9.0 263.3 ;
      RECT  15.6 283.5 9.0 282.9 ;
      RECT  5.8 265.7 5.0 264.9 ;
      RECT  7.8 265.7 7.0 264.9 ;
      RECT  5.8 282.3 5.0 281.5 ;
      RECT  7.8 282.3 7.0 281.5 ;
      RECT  7.4 274.0 6.6 273.2 ;
      RECT  5.4 273.9 4.8 273.3 ;
      RECT  9.0 263.9 2.4 263.3 ;
      RECT  9.0 283.5 2.4 282.9 ;
      RECT  32.2 300.7 31.4 301.5 ;
      RECT  34.2 300.7 33.4 301.5 ;
      RECT  32.2 284.1 31.4 284.9 ;
      RECT  34.2 284.1 33.4 284.9 ;
      RECT  33.8 292.4 33.0 293.2 ;
      RECT  31.8 292.5 31.2 293.1 ;
      RECT  35.4 302.5 28.8 303.1 ;
      RECT  35.4 282.9 28.8 283.5 ;
      RECT  25.6 300.7 24.8 301.5 ;
      RECT  27.6 300.7 26.8 301.5 ;
      RECT  25.6 284.1 24.8 284.9 ;
      RECT  27.6 284.1 26.8 284.9 ;
      RECT  27.2 292.4 26.4 293.2 ;
      RECT  25.2 292.5 24.6 293.1 ;
      RECT  28.8 302.5 22.2 303.1 ;
      RECT  28.8 282.9 22.2 283.5 ;
      RECT  19.0 300.7 18.2 301.5 ;
      RECT  21.0 300.7 20.2 301.5 ;
      RECT  19.0 284.1 18.2 284.9 ;
      RECT  21.0 284.1 20.2 284.9 ;
      RECT  20.6 292.4 19.8 293.2 ;
      RECT  18.6 292.5 18.0 293.1 ;
      RECT  22.2 302.5 15.6 303.1 ;
      RECT  22.2 282.9 15.6 283.5 ;
      RECT  12.4 300.7 11.6 301.5 ;
      RECT  14.4 300.7 13.6 301.5 ;
      RECT  12.4 284.1 11.6 284.9 ;
      RECT  14.4 284.1 13.6 284.9 ;
      RECT  14.0 292.4 13.2 293.2 ;
      RECT  12.0 292.5 11.4 293.1 ;
      RECT  15.6 302.5 9.0 303.1 ;
      RECT  15.6 282.9 9.0 283.5 ;
      RECT  5.8 300.7 5.0 301.5 ;
      RECT  7.8 300.7 7.0 301.5 ;
      RECT  5.8 284.1 5.0 284.9 ;
      RECT  7.8 284.1 7.0 284.9 ;
      RECT  7.4 292.4 6.6 293.2 ;
      RECT  5.4 292.5 4.8 293.1 ;
      RECT  9.0 302.5 2.4 303.1 ;
      RECT  9.0 282.9 2.4 283.5 ;
      RECT  32.2 304.9 31.4 304.1 ;
      RECT  34.2 304.9 33.4 304.1 ;
      RECT  32.2 321.5 31.4 320.7 ;
      RECT  34.2 321.5 33.4 320.7 ;
      RECT  33.8 313.2 33.0 312.4 ;
      RECT  31.8 313.1 31.2 312.5 ;
      RECT  35.4 303.1 28.8 302.5 ;
      RECT  35.4 322.7 28.8 322.1 ;
      RECT  25.6 304.9 24.8 304.1 ;
      RECT  27.6 304.9 26.8 304.1 ;
      RECT  25.6 321.5 24.8 320.7 ;
      RECT  27.6 321.5 26.8 320.7 ;
      RECT  27.2 313.2 26.4 312.4 ;
      RECT  25.2 313.1 24.6 312.5 ;
      RECT  28.8 303.1 22.2 302.5 ;
      RECT  28.8 322.7 22.2 322.1 ;
      RECT  19.0 304.9 18.2 304.1 ;
      RECT  21.0 304.9 20.2 304.1 ;
      RECT  19.0 321.5 18.2 320.7 ;
      RECT  21.0 321.5 20.2 320.7 ;
      RECT  20.6 313.2 19.8 312.4 ;
      RECT  18.6 313.1 18.0 312.5 ;
      RECT  22.2 303.1 15.6 302.5 ;
      RECT  22.2 322.7 15.6 322.1 ;
      RECT  12.4 304.9 11.6 304.1 ;
      RECT  14.4 304.9 13.6 304.1 ;
      RECT  12.4 321.5 11.6 320.7 ;
      RECT  14.4 321.5 13.6 320.7 ;
      RECT  14.0 313.2 13.2 312.4 ;
      RECT  12.0 313.1 11.4 312.5 ;
      RECT  15.6 303.1 9.0 302.5 ;
      RECT  15.6 322.7 9.0 322.1 ;
      RECT  5.8 304.9 5.0 304.1 ;
      RECT  7.8 304.9 7.0 304.1 ;
      RECT  5.8 321.5 5.0 320.7 ;
      RECT  7.8 321.5 7.0 320.7 ;
      RECT  7.4 313.2 6.6 312.4 ;
      RECT  5.4 313.1 4.8 312.5 ;
      RECT  9.0 303.1 2.4 302.5 ;
      RECT  9.0 322.7 2.4 322.1 ;
      RECT  32.2 339.9 31.4 340.7 ;
      RECT  34.2 339.9 33.4 340.7 ;
      RECT  32.2 323.3 31.4 324.1 ;
      RECT  34.2 323.3 33.4 324.1 ;
      RECT  33.8 331.6 33.0 332.4 ;
      RECT  31.8 331.7 31.2 332.3 ;
      RECT  35.4 341.7 28.8 342.3 ;
      RECT  35.4 322.1 28.8 322.7 ;
      RECT  25.6 339.9 24.8 340.7 ;
      RECT  27.6 339.9 26.8 340.7 ;
      RECT  25.6 323.3 24.8 324.1 ;
      RECT  27.6 323.3 26.8 324.1 ;
      RECT  27.2 331.6 26.4 332.4 ;
      RECT  25.2 331.7 24.6 332.3 ;
      RECT  28.8 341.7 22.2 342.3 ;
      RECT  28.8 322.1 22.2 322.7 ;
      RECT  19.0 339.9 18.2 340.7 ;
      RECT  21.0 339.9 20.2 340.7 ;
      RECT  19.0 323.3 18.2 324.1 ;
      RECT  21.0 323.3 20.2 324.1 ;
      RECT  20.6 331.6 19.8 332.4 ;
      RECT  18.6 331.7 18.0 332.3 ;
      RECT  22.2 341.7 15.6 342.3 ;
      RECT  22.2 322.1 15.6 322.7 ;
      RECT  12.4 339.9 11.6 340.7 ;
      RECT  14.4 339.9 13.6 340.7 ;
      RECT  12.4 323.3 11.6 324.1 ;
      RECT  14.4 323.3 13.6 324.1 ;
      RECT  14.0 331.6 13.2 332.4 ;
      RECT  12.0 331.7 11.4 332.3 ;
      RECT  15.6 341.7 9.0 342.3 ;
      RECT  15.6 322.1 9.0 322.7 ;
      RECT  5.8 339.9 5.0 340.7 ;
      RECT  7.8 339.9 7.0 340.7 ;
      RECT  5.8 323.3 5.0 324.1 ;
      RECT  7.8 323.3 7.0 324.1 ;
      RECT  7.4 331.6 6.6 332.4 ;
      RECT  5.4 331.7 4.8 332.3 ;
      RECT  9.0 341.7 2.4 342.3 ;
      RECT  9.0 322.1 2.4 322.7 ;
      RECT  55.6 104.9 56.4 104.1 ;
      RECT  53.6 104.9 54.4 104.1 ;
      RECT  57.6 104.9 58.4 104.1 ;
      RECT  55.6 104.9 56.4 104.1 ;
      RECT  53.6 121.5 54.4 120.7 ;
      RECT  57.6 121.5 58.4 120.7 ;
      RECT  54.6 120.0 55.4 119.2 ;
      RECT  56.6 117.2 57.4 116.4 ;
      RECT  59.1 106.2 59.7 105.6 ;
      RECT  52.4 103.1 61.0 102.5 ;
      RECT  52.4 123.1 61.0 122.5 ;
      RECT  64.2 104.9 65.0 104.1 ;
      RECT  62.2 104.9 63.0 104.1 ;
      RECT  64.2 121.9 65.0 121.1 ;
      RECT  62.2 121.9 63.0 121.1 ;
      RECT  62.6 113.4 63.4 112.6 ;
      RECT  64.6 113.3 65.2 112.7 ;
      RECT  61.0 103.1 67.6 102.5 ;
      RECT  61.0 123.1 67.6 122.5 ;
      RECT  70.8 104.9 71.6 104.1 ;
      RECT  68.8 104.9 69.6 104.1 ;
      RECT  70.8 121.9 71.6 121.1 ;
      RECT  68.8 121.9 69.6 121.1 ;
      RECT  69.2 113.4 70.0 112.6 ;
      RECT  71.2 113.3 71.8 112.7 ;
      RECT  67.6 103.1 72.8 102.5 ;
      RECT  67.6 123.1 72.8 122.5 ;
      RECT  62.6 113.4 63.4 112.6 ;
      RECT  71.2 113.3 71.8 112.7 ;
      RECT  61.0 103.1 72.8 102.5 ;
      RECT  61.0 123.1 72.8 122.5 ;
      RECT  71.6 352.8 72.4 353.0 ;
      RECT  58.8 346.0 59.6 350.8 ;
      RECT  67.6 359.0 68.2 359.6 ;
      RECT  65.4 358.4 69.0 359.0 ;
      RECT  58.8 354.6 64.4 354.8 ;
      RECT  59.6 351.6 70.6 352.2 ;
      RECT  76.4 355.0 77.2 363.6 ;
      RECT  67.6 348.0 68.2 348.6 ;
      RECT  63.2 346.0 64.0 347.4 ;
      RECT  65.4 358.2 66.2 358.4 ;
      RECT  71.6 358.8 72.4 359.6 ;
      RECT  68.0 355.6 68.6 356.8 ;
      RECT  62.0 359.6 64.0 360.2 ;
      RECT  69.2 345.4 70.0 348.0 ;
      RECT  65.4 348.6 68.2 349.2 ;
      RECT  62.0 347.4 64.0 348.0 ;
      RECT  76.4 351.0 77.2 354.4 ;
      RECT  71.8 359.6 73.0 363.6 ;
      RECT  60.4 355.8 61.2 364.2 ;
      RECT  62.0 356.2 67.4 356.8 ;
      RECT  70.0 352.2 70.6 355.4 ;
      RECT  57.6 364.2 79.4 365.4 ;
      RECT  73.0 354.4 77.2 355.0 ;
      RECT  74.8 355.6 75.6 364.2 ;
      RECT  78.0 345.4 78.8 346.8 ;
      RECT  71.8 356.0 72.4 357.0 ;
      RECT  70.0 355.4 72.4 356.0 ;
      RECT  58.8 355.2 59.6 363.6 ;
      RECT  71.6 347.4 73.0 348.0 ;
      RECT  68.0 356.8 70.2 357.4 ;
      RECT  63.2 360.2 64.0 363.6 ;
      RECT  61.0 353.4 66.0 354.0 ;
      RECT  78.0 362.6 78.8 364.2 ;
      RECT  71.6 353.0 75.4 353.6 ;
      RECT  71.6 348.0 72.4 348.8 ;
      RECT  57.6 344.2 79.4 345.4 ;
      RECT  65.2 354.0 66.0 354.2 ;
      RECT  62.6 352.2 63.4 352.4 ;
      RECT  68.2 358.2 69.0 358.4 ;
      RECT  76.4 346.0 77.2 350.4 ;
      RECT  59.6 351.4 61.2 351.6 ;
      RECT  62.0 358.8 62.8 359.6 ;
      RECT  67.6 346.0 68.4 348.0 ;
      RECT  61.0 353.2 61.8 353.4 ;
      RECT  62.0 356.8 62.8 357.0 ;
      RECT  73.4 350.2 74.2 350.4 ;
      RECT  63.6 348.6 64.4 349.4 ;
      RECT  74.8 345.4 75.6 349.8 ;
      RECT  69.4 356.6 70.2 356.8 ;
      RECT  65.8 345.4 66.8 348.0 ;
      RECT  63.8 349.4 64.4 351.6 ;
      RECT  69.2 359.6 70.0 364.2 ;
      RECT  66.0 359.6 66.8 364.2 ;
      RECT  69.4 351.4 70.2 351.6 ;
      RECT  63.8 355.2 68.6 355.6 ;
      RECT  58.8 354.8 64.6 355.0 ;
      RECT  67.6 359.6 68.4 363.6 ;
      RECT  74.6 353.6 75.4 353.8 ;
      RECT  58.8 355.0 68.6 355.2 ;
      RECT  66.6 356.8 67.4 357.0 ;
      RECT  71.8 346.0 73.0 347.4 ;
      RECT  65.4 349.2 66.2 349.4 ;
      RECT  71.8 357.0 73.2 357.8 ;
      RECT  73.0 354.2 73.8 354.4 ;
      RECT  62.0 348.0 62.8 348.8 ;
      RECT  60.4 345.4 61.2 350.0 ;
      RECT  73.4 350.4 77.2 351.0 ;
      RECT  71.6 376.8 72.4 376.6 ;
      RECT  58.8 383.6 59.6 378.8 ;
      RECT  67.6 370.6 68.2 370.0 ;
      RECT  65.4 371.2 69.0 370.6 ;
      RECT  58.8 375.0 64.4 374.8 ;
      RECT  59.6 378.0 70.6 377.4 ;
      RECT  76.4 374.6 77.2 366.0 ;
      RECT  67.6 381.6 68.2 381.0 ;
      RECT  63.2 383.6 64.0 382.2 ;
      RECT  65.4 371.4 66.2 371.2 ;
      RECT  71.6 370.8 72.4 370.0 ;
      RECT  68.0 374.0 68.6 372.8 ;
      RECT  62.0 370.0 64.0 369.4 ;
      RECT  69.2 384.2 70.0 381.6 ;
      RECT  65.4 381.0 68.2 380.4 ;
      RECT  62.0 382.2 64.0 381.6 ;
      RECT  76.4 378.6 77.2 375.2 ;
      RECT  71.8 370.0 73.0 366.0 ;
      RECT  60.4 373.8 61.2 365.4 ;
      RECT  62.0 373.4 67.4 372.8 ;
      RECT  70.0 377.4 70.6 374.2 ;
      RECT  57.6 365.4 79.4 364.2 ;
      RECT  73.0 375.2 77.2 374.6 ;
      RECT  74.8 374.0 75.6 365.4 ;
      RECT  78.0 384.2 78.8 382.8 ;
      RECT  71.8 373.6 72.4 372.6 ;
      RECT  70.0 374.2 72.4 373.6 ;
      RECT  58.8 374.4 59.6 366.0 ;
      RECT  71.6 382.2 73.0 381.6 ;
      RECT  68.0 372.8 70.2 372.2 ;
      RECT  63.2 369.4 64.0 366.0 ;
      RECT  61.0 376.2 66.0 375.6 ;
      RECT  78.0 367.0 78.8 365.4 ;
      RECT  71.6 376.6 75.4 376.0 ;
      RECT  71.6 381.6 72.4 380.8 ;
      RECT  57.6 385.4 79.4 384.2 ;
      RECT  65.2 375.6 66.0 375.4 ;
      RECT  62.6 377.4 63.4 377.2 ;
      RECT  68.2 371.4 69.0 371.2 ;
      RECT  76.4 383.6 77.2 379.2 ;
      RECT  59.6 378.2 61.2 378.0 ;
      RECT  62.0 370.8 62.8 370.0 ;
      RECT  67.6 383.6 68.4 381.6 ;
      RECT  61.0 376.4 61.8 376.2 ;
      RECT  62.0 372.8 62.8 372.6 ;
      RECT  73.4 379.4 74.2 379.2 ;
      RECT  63.6 381.0 64.4 380.2 ;
      RECT  74.8 384.2 75.6 379.8 ;
      RECT  69.4 373.0 70.2 372.8 ;
      RECT  65.8 384.2 66.8 381.6 ;
      RECT  63.8 380.2 64.4 378.0 ;
      RECT  69.2 370.0 70.0 365.4 ;
      RECT  66.0 370.0 66.8 365.4 ;
      RECT  69.4 378.2 70.2 378.0 ;
      RECT  63.8 374.4 68.6 374.0 ;
      RECT  58.8 374.8 64.6 374.6 ;
      RECT  67.6 370.0 68.4 366.0 ;
      RECT  74.6 376.0 75.4 375.8 ;
      RECT  58.8 374.6 68.6 374.4 ;
      RECT  66.6 372.8 67.4 372.6 ;
      RECT  71.8 383.6 73.0 382.2 ;
      RECT  65.4 380.4 66.2 380.2 ;
      RECT  71.8 372.6 73.2 371.8 ;
      RECT  73.0 375.4 73.8 375.2 ;
      RECT  62.0 381.6 62.8 380.8 ;
      RECT  60.4 384.2 61.2 379.6 ;
      RECT  73.4 379.2 77.2 378.6 ;
      RECT  71.6 392.8 72.4 393.0 ;
      RECT  58.8 386.0 59.6 390.8 ;
      RECT  67.6 399.0 68.2 399.6 ;
      RECT  65.4 398.4 69.0 399.0 ;
      RECT  58.8 394.6 64.4 394.8 ;
      RECT  59.6 391.6 70.6 392.2 ;
      RECT  76.4 395.0 77.2 403.6 ;
      RECT  67.6 388.0 68.2 388.6 ;
      RECT  63.2 386.0 64.0 387.4 ;
      RECT  65.4 398.2 66.2 398.4 ;
      RECT  71.6 398.8 72.4 399.6 ;
      RECT  68.0 395.6 68.6 396.8 ;
      RECT  62.0 399.6 64.0 400.2 ;
      RECT  69.2 385.4 70.0 388.0 ;
      RECT  65.4 388.6 68.2 389.2 ;
      RECT  62.0 387.4 64.0 388.0 ;
      RECT  76.4 391.0 77.2 394.4 ;
      RECT  71.8 399.6 73.0 403.6 ;
      RECT  60.4 395.8 61.2 404.2 ;
      RECT  62.0 396.2 67.4 396.8 ;
      RECT  70.0 392.2 70.6 395.4 ;
      RECT  57.6 404.2 79.4 405.4 ;
      RECT  73.0 394.4 77.2 395.0 ;
      RECT  74.8 395.6 75.6 404.2 ;
      RECT  78.0 385.4 78.8 386.8 ;
      RECT  71.8 396.0 72.4 397.0 ;
      RECT  70.0 395.4 72.4 396.0 ;
      RECT  58.8 395.2 59.6 403.6 ;
      RECT  71.6 387.4 73.0 388.0 ;
      RECT  68.0 396.8 70.2 397.4 ;
      RECT  63.2 400.2 64.0 403.6 ;
      RECT  61.0 393.4 66.0 394.0 ;
      RECT  78.0 402.6 78.8 404.2 ;
      RECT  71.6 393.0 75.4 393.6 ;
      RECT  71.6 388.0 72.4 388.8 ;
      RECT  57.6 384.2 79.4 385.4 ;
      RECT  65.2 394.0 66.0 394.2 ;
      RECT  62.6 392.2 63.4 392.4 ;
      RECT  68.2 398.2 69.0 398.4 ;
      RECT  76.4 386.0 77.2 390.4 ;
      RECT  59.6 391.4 61.2 391.6 ;
      RECT  62.0 398.8 62.8 399.6 ;
      RECT  67.6 386.0 68.4 388.0 ;
      RECT  61.0 393.2 61.8 393.4 ;
      RECT  62.0 396.8 62.8 397.0 ;
      RECT  73.4 390.2 74.2 390.4 ;
      RECT  63.6 388.6 64.4 389.4 ;
      RECT  74.8 385.4 75.6 389.8 ;
      RECT  69.4 396.6 70.2 396.8 ;
      RECT  65.8 385.4 66.8 388.0 ;
      RECT  63.8 389.4 64.4 391.6 ;
      RECT  69.2 399.6 70.0 404.2 ;
      RECT  66.0 399.6 66.8 404.2 ;
      RECT  69.4 391.4 70.2 391.6 ;
      RECT  63.8 395.2 68.6 395.6 ;
      RECT  58.8 394.8 64.6 395.0 ;
      RECT  67.6 399.6 68.4 403.6 ;
      RECT  74.6 393.6 75.4 393.8 ;
      RECT  58.8 395.0 68.6 395.2 ;
      RECT  66.6 396.8 67.4 397.0 ;
      RECT  71.8 386.0 73.0 387.4 ;
      RECT  65.4 389.2 66.2 389.4 ;
      RECT  71.8 397.0 73.2 397.8 ;
      RECT  73.0 394.2 73.8 394.4 ;
      RECT  62.0 388.0 62.8 388.8 ;
      RECT  60.4 385.4 61.2 390.0 ;
      RECT  73.4 390.4 77.2 391.0 ;
      RECT  71.6 416.8 72.4 416.6 ;
      RECT  58.8 423.6 59.6 418.8 ;
      RECT  67.6 410.6 68.2 410.0 ;
      RECT  65.4 411.2 69.0 410.6 ;
      RECT  58.8 415.0 64.4 414.8 ;
      RECT  59.6 418.0 70.6 417.4 ;
      RECT  76.4 414.6 77.2 406.0 ;
      RECT  67.6 421.6 68.2 421.0 ;
      RECT  63.2 423.6 64.0 422.2 ;
      RECT  65.4 411.4 66.2 411.2 ;
      RECT  71.6 410.8 72.4 410.0 ;
      RECT  68.0 414.0 68.6 412.8 ;
      RECT  62.0 410.0 64.0 409.4 ;
      RECT  69.2 424.2 70.0 421.6 ;
      RECT  65.4 421.0 68.2 420.4 ;
      RECT  62.0 422.2 64.0 421.6 ;
      RECT  76.4 418.6 77.2 415.2 ;
      RECT  71.8 410.0 73.0 406.0 ;
      RECT  60.4 413.8 61.2 405.4 ;
      RECT  62.0 413.4 67.4 412.8 ;
      RECT  70.0 417.4 70.6 414.2 ;
      RECT  57.6 405.4 79.4 404.2 ;
      RECT  73.0 415.2 77.2 414.6 ;
      RECT  74.8 414.0 75.6 405.4 ;
      RECT  78.0 424.2 78.8 422.8 ;
      RECT  71.8 413.6 72.4 412.6 ;
      RECT  70.0 414.2 72.4 413.6 ;
      RECT  58.8 414.4 59.6 406.0 ;
      RECT  71.6 422.2 73.0 421.6 ;
      RECT  68.0 412.8 70.2 412.2 ;
      RECT  63.2 409.4 64.0 406.0 ;
      RECT  61.0 416.2 66.0 415.6 ;
      RECT  78.0 407.0 78.8 405.4 ;
      RECT  71.6 416.6 75.4 416.0 ;
      RECT  71.6 421.6 72.4 420.8 ;
      RECT  57.6 425.4 79.4 424.2 ;
      RECT  65.2 415.6 66.0 415.4 ;
      RECT  62.6 417.4 63.4 417.2 ;
      RECT  68.2 411.4 69.0 411.2 ;
      RECT  76.4 423.6 77.2 419.2 ;
      RECT  59.6 418.2 61.2 418.0 ;
      RECT  62.0 410.8 62.8 410.0 ;
      RECT  67.6 423.6 68.4 421.6 ;
      RECT  61.0 416.4 61.8 416.2 ;
      RECT  62.0 412.8 62.8 412.6 ;
      RECT  73.4 419.4 74.2 419.2 ;
      RECT  63.6 421.0 64.4 420.2 ;
      RECT  74.8 424.2 75.6 419.8 ;
      RECT  69.4 413.0 70.2 412.8 ;
      RECT  65.8 424.2 66.8 421.6 ;
      RECT  63.8 420.2 64.4 418.0 ;
      RECT  69.2 410.0 70.0 405.4 ;
      RECT  66.0 410.0 66.8 405.4 ;
      RECT  69.4 418.2 70.2 418.0 ;
      RECT  63.8 414.4 68.6 414.0 ;
      RECT  58.8 414.8 64.6 414.6 ;
      RECT  67.6 410.0 68.4 406.0 ;
      RECT  74.6 416.0 75.4 415.8 ;
      RECT  58.8 414.6 68.6 414.4 ;
      RECT  66.6 412.8 67.4 412.6 ;
      RECT  71.8 423.6 73.0 422.2 ;
      RECT  65.4 420.4 66.2 420.2 ;
      RECT  71.8 412.6 73.2 411.8 ;
      RECT  73.0 415.4 73.8 415.2 ;
      RECT  62.0 421.6 62.8 420.8 ;
      RECT  60.4 424.2 61.2 419.6 ;
      RECT  73.4 419.2 77.2 418.6 ;
      RECT  115.2 10.8 116.0 11.0 ;
      RECT  102.4 4.0 103.2 8.8 ;
      RECT  111.2 17.0 111.8 17.6 ;
      RECT  109.0 16.4 112.6 17.0 ;
      RECT  102.4 12.6 108.0 12.8 ;
      RECT  103.2 9.6 114.2 10.2 ;
      RECT  120.0 13.0 120.8 21.6 ;
      RECT  111.2 6.0 111.8 6.6 ;
      RECT  106.8 4.0 107.6 5.4 ;
      RECT  109.0 16.2 109.8 16.4 ;
      RECT  115.2 16.8 116.0 17.6 ;
      RECT  111.6 13.6 112.2 14.8 ;
      RECT  105.6 17.6 107.6 18.2 ;
      RECT  112.8 3.4 113.6 6.0 ;
      RECT  109.0 6.6 111.8 7.2 ;
      RECT  105.6 5.4 107.6 6.0 ;
      RECT  120.0 9.0 120.8 12.4 ;
      RECT  115.4 17.6 116.6 21.6 ;
      RECT  104.0 13.8 104.8 22.2 ;
      RECT  105.6 14.2 111.0 14.8 ;
      RECT  113.6 10.2 114.2 13.4 ;
      RECT  101.2 22.2 123.0 23.4 ;
      RECT  116.6 12.4 120.8 13.0 ;
      RECT  118.4 13.6 119.2 22.2 ;
      RECT  121.6 3.4 122.4 4.8 ;
      RECT  115.4 14.0 116.0 15.0 ;
      RECT  113.6 13.4 116.0 14.0 ;
      RECT  102.4 13.2 103.2 21.6 ;
      RECT  115.2 5.4 116.6 6.0 ;
      RECT  111.6 14.8 113.8 15.4 ;
      RECT  106.8 18.2 107.6 21.6 ;
      RECT  104.6 11.4 109.6 12.0 ;
      RECT  121.6 20.6 122.4 22.2 ;
      RECT  115.2 11.0 119.0 11.6 ;
      RECT  115.2 6.0 116.0 6.8 ;
      RECT  101.2 2.2 123.0 3.4 ;
      RECT  108.8 12.0 109.6 12.2 ;
      RECT  106.2 10.2 107.0 10.4 ;
      RECT  111.8 16.2 112.6 16.4 ;
      RECT  120.0 4.0 120.8 8.4 ;
      RECT  103.2 9.4 104.8 9.6 ;
      RECT  105.6 16.8 106.4 17.6 ;
      RECT  111.2 4.0 112.0 6.0 ;
      RECT  104.6 11.2 105.4 11.4 ;
      RECT  105.6 14.8 106.4 15.0 ;
      RECT  117.0 8.2 117.8 8.4 ;
      RECT  107.2 6.6 108.0 7.4 ;
      RECT  118.4 3.4 119.2 7.8 ;
      RECT  113.0 14.6 113.8 14.8 ;
      RECT  109.4 3.4 110.4 6.0 ;
      RECT  107.4 7.4 108.0 9.6 ;
      RECT  112.8 17.6 113.6 22.2 ;
      RECT  109.6 17.6 110.4 22.2 ;
      RECT  113.0 9.4 113.8 9.6 ;
      RECT  107.4 13.2 112.2 13.6 ;
      RECT  102.4 12.8 108.2 13.0 ;
      RECT  111.2 17.6 112.0 21.6 ;
      RECT  118.2 11.6 119.0 11.8 ;
      RECT  102.4 13.0 112.2 13.2 ;
      RECT  110.2 14.8 111.0 15.0 ;
      RECT  115.4 4.0 116.6 5.4 ;
      RECT  109.0 7.2 109.8 7.4 ;
      RECT  115.4 15.0 116.8 15.8 ;
      RECT  116.6 12.2 117.4 12.4 ;
      RECT  105.6 6.0 106.4 6.8 ;
      RECT  104.0 3.4 104.8 8.0 ;
      RECT  117.0 8.4 120.8 9.0 ;
      RECT  137.0 10.8 137.8 11.0 ;
      RECT  124.2 4.0 125.0 8.8 ;
      RECT  133.0 17.0 133.6 17.6 ;
      RECT  130.8 16.4 134.4 17.0 ;
      RECT  124.2 12.6 129.8 12.8 ;
      RECT  125.0 9.6 136.0 10.2 ;
      RECT  141.8 13.0 142.6 21.6 ;
      RECT  133.0 6.0 133.6 6.6 ;
      RECT  128.6 4.0 129.4 5.4 ;
      RECT  130.8 16.2 131.6 16.4 ;
      RECT  137.0 16.8 137.8 17.6 ;
      RECT  133.4 13.6 134.0 14.8 ;
      RECT  127.4 17.6 129.4 18.2 ;
      RECT  134.6 3.4 135.4 6.0 ;
      RECT  130.8 6.6 133.6 7.2 ;
      RECT  127.4 5.4 129.4 6.0 ;
      RECT  141.8 9.0 142.6 12.4 ;
      RECT  137.2 17.6 138.4 21.6 ;
      RECT  125.8 13.8 126.6 22.2 ;
      RECT  127.4 14.2 132.8 14.8 ;
      RECT  135.4 10.2 136.0 13.4 ;
      RECT  123.0 22.2 144.8 23.4 ;
      RECT  138.4 12.4 142.6 13.0 ;
      RECT  140.2 13.6 141.0 22.2 ;
      RECT  143.4 3.4 144.2 4.8 ;
      RECT  137.2 14.0 137.8 15.0 ;
      RECT  135.4 13.4 137.8 14.0 ;
      RECT  124.2 13.2 125.0 21.6 ;
      RECT  137.0 5.4 138.4 6.0 ;
      RECT  133.4 14.8 135.6 15.4 ;
      RECT  128.6 18.2 129.4 21.6 ;
      RECT  126.4 11.4 131.4 12.0 ;
      RECT  143.4 20.6 144.2 22.2 ;
      RECT  137.0 11.0 140.8 11.6 ;
      RECT  137.0 6.0 137.8 6.8 ;
      RECT  123.0 2.2 144.8 3.4 ;
      RECT  130.6 12.0 131.4 12.2 ;
      RECT  128.0 10.2 128.8 10.4 ;
      RECT  133.6 16.2 134.4 16.4 ;
      RECT  141.8 4.0 142.6 8.4 ;
      RECT  125.0 9.4 126.6 9.6 ;
      RECT  127.4 16.8 128.2 17.6 ;
      RECT  133.0 4.0 133.8 6.0 ;
      RECT  126.4 11.2 127.2 11.4 ;
      RECT  127.4 14.8 128.2 15.0 ;
      RECT  138.8 8.2 139.6 8.4 ;
      RECT  129.0 6.6 129.8 7.4 ;
      RECT  140.2 3.4 141.0 7.8 ;
      RECT  134.8 14.6 135.6 14.8 ;
      RECT  131.2 3.4 132.2 6.0 ;
      RECT  129.2 7.4 129.8 9.6 ;
      RECT  134.6 17.6 135.4 22.2 ;
      RECT  131.4 17.6 132.2 22.2 ;
      RECT  134.8 9.4 135.6 9.6 ;
      RECT  129.2 13.2 134.0 13.6 ;
      RECT  124.2 12.8 130.0 13.0 ;
      RECT  133.0 17.6 133.8 21.6 ;
      RECT  140.0 11.6 140.8 11.8 ;
      RECT  124.2 13.0 134.0 13.2 ;
      RECT  132.0 14.8 132.8 15.0 ;
      RECT  137.2 4.0 138.4 5.4 ;
      RECT  130.8 7.2 131.6 7.4 ;
      RECT  137.2 15.0 138.6 15.8 ;
      RECT  138.4 12.2 139.2 12.4 ;
      RECT  127.4 6.0 128.2 6.8 ;
      RECT  125.8 3.4 126.6 8.0 ;
      RECT  138.8 8.4 142.6 9.0 ;
   LAYER  m2 ;
      RECT  189.9 196.4 190.7 197.2 ;
      RECT  186.5 186.4 187.3 197.2 ;
      RECT  191.7 188.0 192.5 197.2 ;
      RECT  188.1 186.4 188.9 197.2 ;
      RECT  190.9 187.2 192.5 188.0 ;
      RECT  193.3 186.4 194.1 197.2 ;
      RECT  191.7 186.4 192.5 187.2 ;
      RECT  189.9 197.2 190.7 196.4 ;
      RECT  186.5 207.2 187.3 196.4 ;
      RECT  191.7 205.6 192.5 196.4 ;
      RECT  188.1 207.2 188.9 196.4 ;
      RECT  190.9 206.4 192.5 205.6 ;
      RECT  193.3 207.2 194.1 196.4 ;
      RECT  191.7 207.2 192.5 206.4 ;
      RECT  189.9 217.2 190.7 218.0 ;
      RECT  186.5 207.2 187.3 218.0 ;
      RECT  191.7 208.8 192.5 218.0 ;
      RECT  188.1 207.2 188.9 218.0 ;
      RECT  190.9 208.0 192.5 208.8 ;
      RECT  193.3 207.2 194.1 218.0 ;
      RECT  191.7 207.2 192.5 208.0 ;
      RECT  189.9 218.0 190.7 217.2 ;
      RECT  186.5 228.0 187.3 217.2 ;
      RECT  191.7 226.4 192.5 217.2 ;
      RECT  188.1 228.0 188.9 217.2 ;
      RECT  190.9 227.2 192.5 226.4 ;
      RECT  193.3 228.0 194.1 217.2 ;
      RECT  191.7 228.0 192.5 227.2 ;
      RECT  189.9 238.0 190.7 238.8 ;
      RECT  186.5 228.0 187.3 238.8 ;
      RECT  191.7 229.6 192.5 238.8 ;
      RECT  188.1 228.0 188.9 238.8 ;
      RECT  190.9 228.8 192.5 229.6 ;
      RECT  193.3 228.0 194.1 238.8 ;
      RECT  191.7 228.0 192.5 228.8 ;
      RECT  189.9 238.8 190.7 238.0 ;
      RECT  186.5 248.8 187.3 238.0 ;
      RECT  191.7 247.2 192.5 238.0 ;
      RECT  188.1 248.8 188.9 238.0 ;
      RECT  190.9 248.0 192.5 247.2 ;
      RECT  193.3 248.8 194.1 238.0 ;
      RECT  191.7 248.8 192.5 248.0 ;
      RECT  189.9 258.8 190.7 259.6 ;
      RECT  186.5 248.8 187.3 259.6 ;
      RECT  191.7 250.4 192.5 259.6 ;
      RECT  188.1 248.8 188.9 259.6 ;
      RECT  190.9 249.6 192.5 250.4 ;
      RECT  193.3 248.8 194.1 259.6 ;
      RECT  191.7 248.8 192.5 249.6 ;
      RECT  189.9 259.6 190.7 258.8 ;
      RECT  186.5 269.6 187.3 258.8 ;
      RECT  191.7 268.0 192.5 258.8 ;
      RECT  188.1 269.6 188.9 258.8 ;
      RECT  190.9 268.8 192.5 268.0 ;
      RECT  193.3 269.6 194.1 258.8 ;
      RECT  191.7 269.6 192.5 268.8 ;
      RECT  189.9 279.6 190.7 280.4 ;
      RECT  186.5 269.6 187.3 280.4 ;
      RECT  191.7 271.2 192.5 280.4 ;
      RECT  188.1 269.6 188.9 280.4 ;
      RECT  190.9 270.4 192.5 271.2 ;
      RECT  193.3 269.6 194.1 280.4 ;
      RECT  191.7 269.6 192.5 270.4 ;
      RECT  189.9 280.4 190.7 279.6 ;
      RECT  186.5 290.4 187.3 279.6 ;
      RECT  191.7 288.8 192.5 279.6 ;
      RECT  188.1 290.4 188.9 279.6 ;
      RECT  190.9 289.6 192.5 288.8 ;
      RECT  193.3 290.4 194.1 279.6 ;
      RECT  191.7 290.4 192.5 289.6 ;
      RECT  189.9 300.4 190.7 301.2 ;
      RECT  186.5 290.4 187.3 301.2 ;
      RECT  191.7 292.0 192.5 301.2 ;
      RECT  188.1 290.4 188.9 301.2 ;
      RECT  190.9 291.2 192.5 292.0 ;
      RECT  193.3 290.4 194.1 301.2 ;
      RECT  191.7 290.4 192.5 291.2 ;
      RECT  189.9 301.2 190.7 300.4 ;
      RECT  186.5 311.2 187.3 300.4 ;
      RECT  191.7 309.6 192.5 300.4 ;
      RECT  188.1 311.2 188.9 300.4 ;
      RECT  190.9 310.4 192.5 309.6 ;
      RECT  193.3 311.2 194.1 300.4 ;
      RECT  191.7 311.2 192.5 310.4 ;
      RECT  189.9 321.2 190.7 322.0 ;
      RECT  186.5 311.2 187.3 322.0 ;
      RECT  191.7 312.8 192.5 322.0 ;
      RECT  188.1 311.2 188.9 322.0 ;
      RECT  190.9 312.0 192.5 312.8 ;
      RECT  193.3 311.2 194.1 322.0 ;
      RECT  191.7 311.2 192.5 312.0 ;
      RECT  189.9 322.0 190.7 321.2 ;
      RECT  186.5 332.0 187.3 321.2 ;
      RECT  191.7 330.4 192.5 321.2 ;
      RECT  188.1 332.0 188.9 321.2 ;
      RECT  190.9 331.2 192.5 330.4 ;
      RECT  193.3 332.0 194.1 321.2 ;
      RECT  191.7 332.0 192.5 331.2 ;
      RECT  189.9 342.0 190.7 342.8 ;
      RECT  186.5 332.0 187.3 342.8 ;
      RECT  191.7 333.6 192.5 342.8 ;
      RECT  188.1 332.0 188.9 342.8 ;
      RECT  190.9 332.8 192.5 333.6 ;
      RECT  193.3 332.0 194.1 342.8 ;
      RECT  191.7 332.0 192.5 332.8 ;
      RECT  189.9 342.8 190.7 342.0 ;
      RECT  186.5 352.8 187.3 342.0 ;
      RECT  191.7 351.2 192.5 342.0 ;
      RECT  188.1 352.8 188.9 342.0 ;
      RECT  190.9 352.0 192.5 351.2 ;
      RECT  193.3 352.8 194.1 342.0 ;
      RECT  191.7 352.8 192.5 352.0 ;
      RECT  196.7 196.4 197.5 197.2 ;
      RECT  193.3 186.4 194.1 197.2 ;
      RECT  198.5 188.0 199.3 197.2 ;
      RECT  194.9 186.4 195.7 197.2 ;
      RECT  197.7 187.2 199.3 188.0 ;
      RECT  200.1 186.4 200.9 197.2 ;
      RECT  198.5 186.4 199.3 187.2 ;
      RECT  196.7 197.2 197.5 196.4 ;
      RECT  193.3 207.2 194.1 196.4 ;
      RECT  198.5 205.6 199.3 196.4 ;
      RECT  194.9 207.2 195.7 196.4 ;
      RECT  197.7 206.4 199.3 205.6 ;
      RECT  200.1 207.2 200.9 196.4 ;
      RECT  198.5 207.2 199.3 206.4 ;
      RECT  196.7 217.2 197.5 218.0 ;
      RECT  193.3 207.2 194.1 218.0 ;
      RECT  198.5 208.8 199.3 218.0 ;
      RECT  194.9 207.2 195.7 218.0 ;
      RECT  197.7 208.0 199.3 208.8 ;
      RECT  200.1 207.2 200.9 218.0 ;
      RECT  198.5 207.2 199.3 208.0 ;
      RECT  196.7 218.0 197.5 217.2 ;
      RECT  193.3 228.0 194.1 217.2 ;
      RECT  198.5 226.4 199.3 217.2 ;
      RECT  194.9 228.0 195.7 217.2 ;
      RECT  197.7 227.2 199.3 226.4 ;
      RECT  200.1 228.0 200.9 217.2 ;
      RECT  198.5 228.0 199.3 227.2 ;
      RECT  196.7 238.0 197.5 238.8 ;
      RECT  193.3 228.0 194.1 238.8 ;
      RECT  198.5 229.6 199.3 238.8 ;
      RECT  194.9 228.0 195.7 238.8 ;
      RECT  197.7 228.8 199.3 229.6 ;
      RECT  200.1 228.0 200.9 238.8 ;
      RECT  198.5 228.0 199.3 228.8 ;
      RECT  196.7 238.8 197.5 238.0 ;
      RECT  193.3 248.8 194.1 238.0 ;
      RECT  198.5 247.2 199.3 238.0 ;
      RECT  194.9 248.8 195.7 238.0 ;
      RECT  197.7 248.0 199.3 247.2 ;
      RECT  200.1 248.8 200.9 238.0 ;
      RECT  198.5 248.8 199.3 248.0 ;
      RECT  196.7 258.8 197.5 259.6 ;
      RECT  193.3 248.8 194.1 259.6 ;
      RECT  198.5 250.4 199.3 259.6 ;
      RECT  194.9 248.8 195.7 259.6 ;
      RECT  197.7 249.6 199.3 250.4 ;
      RECT  200.1 248.8 200.9 259.6 ;
      RECT  198.5 248.8 199.3 249.6 ;
      RECT  196.7 259.6 197.5 258.8 ;
      RECT  193.3 269.6 194.1 258.8 ;
      RECT  198.5 268.0 199.3 258.8 ;
      RECT  194.9 269.6 195.7 258.8 ;
      RECT  197.7 268.8 199.3 268.0 ;
      RECT  200.1 269.6 200.9 258.8 ;
      RECT  198.5 269.6 199.3 268.8 ;
      RECT  196.7 279.6 197.5 280.4 ;
      RECT  193.3 269.6 194.1 280.4 ;
      RECT  198.5 271.2 199.3 280.4 ;
      RECT  194.9 269.6 195.7 280.4 ;
      RECT  197.7 270.4 199.3 271.2 ;
      RECT  200.1 269.6 200.9 280.4 ;
      RECT  198.5 269.6 199.3 270.4 ;
      RECT  196.7 280.4 197.5 279.6 ;
      RECT  193.3 290.4 194.1 279.6 ;
      RECT  198.5 288.8 199.3 279.6 ;
      RECT  194.9 290.4 195.7 279.6 ;
      RECT  197.7 289.6 199.3 288.8 ;
      RECT  200.1 290.4 200.9 279.6 ;
      RECT  198.5 290.4 199.3 289.6 ;
      RECT  196.7 300.4 197.5 301.2 ;
      RECT  193.3 290.4 194.1 301.2 ;
      RECT  198.5 292.0 199.3 301.2 ;
      RECT  194.9 290.4 195.7 301.2 ;
      RECT  197.7 291.2 199.3 292.0 ;
      RECT  200.1 290.4 200.9 301.2 ;
      RECT  198.5 290.4 199.3 291.2 ;
      RECT  196.7 301.2 197.5 300.4 ;
      RECT  193.3 311.2 194.1 300.4 ;
      RECT  198.5 309.6 199.3 300.4 ;
      RECT  194.9 311.2 195.7 300.4 ;
      RECT  197.7 310.4 199.3 309.6 ;
      RECT  200.1 311.2 200.9 300.4 ;
      RECT  198.5 311.2 199.3 310.4 ;
      RECT  196.7 321.2 197.5 322.0 ;
      RECT  193.3 311.2 194.1 322.0 ;
      RECT  198.5 312.8 199.3 322.0 ;
      RECT  194.9 311.2 195.7 322.0 ;
      RECT  197.7 312.0 199.3 312.8 ;
      RECT  200.1 311.2 200.9 322.0 ;
      RECT  198.5 311.2 199.3 312.0 ;
      RECT  196.7 322.0 197.5 321.2 ;
      RECT  193.3 332.0 194.1 321.2 ;
      RECT  198.5 330.4 199.3 321.2 ;
      RECT  194.9 332.0 195.7 321.2 ;
      RECT  197.7 331.2 199.3 330.4 ;
      RECT  200.1 332.0 200.9 321.2 ;
      RECT  198.5 332.0 199.3 331.2 ;
      RECT  196.7 342.0 197.5 342.8 ;
      RECT  193.3 332.0 194.1 342.8 ;
      RECT  198.5 333.6 199.3 342.8 ;
      RECT  194.9 332.0 195.7 342.8 ;
      RECT  197.7 332.8 199.3 333.6 ;
      RECT  200.1 332.0 200.9 342.8 ;
      RECT  198.5 332.0 199.3 332.8 ;
      RECT  196.7 342.8 197.5 342.0 ;
      RECT  193.3 352.8 194.1 342.0 ;
      RECT  198.5 351.2 199.3 342.0 ;
      RECT  194.9 352.8 195.7 342.0 ;
      RECT  197.7 352.0 199.3 351.2 ;
      RECT  200.1 352.8 200.9 342.0 ;
      RECT  198.5 352.8 199.3 352.0 ;
      RECT  188.1 186.4 188.9 352.8 ;
      RECT  191.7 186.4 192.5 352.8 ;
      RECT  194.9 186.4 195.7 352.8 ;
      RECT  198.5 186.4 199.3 352.8 ;
      RECT  189.9 321.2 190.7 322.0 ;
      RECT  189.9 321.2 190.7 322.0 ;
      RECT  189.9 342.0 190.7 342.8 ;
      RECT  189.9 258.8 190.7 259.6 ;
      RECT  196.7 196.4 197.5 197.2 ;
      RECT  196.7 300.4 197.5 301.2 ;
      RECT  196.7 300.4 197.5 301.2 ;
      RECT  196.7 342.0 197.5 342.8 ;
      RECT  196.7 238.0 197.5 238.8 ;
      RECT  189.9 300.4 190.7 301.2 ;
      RECT  196.7 238.0 197.5 238.8 ;
      RECT  189.9 300.4 190.7 301.2 ;
      RECT  189.9 196.4 190.7 197.2 ;
      RECT  189.9 238.0 190.7 238.8 ;
      RECT  196.7 217.2 197.5 218.0 ;
      RECT  189.9 279.6 190.7 280.4 ;
      RECT  196.7 258.8 197.5 259.6 ;
      RECT  196.7 321.2 197.5 322.0 ;
      RECT  196.7 321.2 197.5 322.0 ;
      RECT  189.9 217.2 190.7 218.0 ;
      RECT  196.7 279.6 197.5 280.4 ;
      RECT  189.9 238.0 190.7 238.8 ;
      RECT  200.1 207.2 200.9 218.0 ;
      RECT  200.1 279.6 200.9 290.4 ;
      RECT  193.3 290.4 194.1 301.2 ;
      RECT  200.1 342.0 200.9 352.8 ;
      RECT  200.1 321.2 200.9 332.0 ;
      RECT  200.1 258.8 200.9 269.6 ;
      RECT  186.5 258.8 187.3 269.6 ;
      RECT  186.5 196.4 187.3 207.2 ;
      RECT  186.5 228.0 187.3 238.8 ;
      RECT  193.3 238.0 194.1 248.8 ;
      RECT  193.3 238.0 194.1 248.8 ;
      RECT  200.1 228.0 200.9 238.8 ;
      RECT  200.1 186.4 200.9 197.2 ;
      RECT  186.5 269.6 187.3 280.4 ;
      RECT  186.5 238.0 187.3 248.8 ;
      RECT  186.5 290.4 187.3 301.2 ;
      RECT  200.1 311.2 200.9 322.0 ;
      RECT  186.5 342.0 187.3 352.8 ;
      RECT  193.3 300.4 194.1 311.2 ;
      RECT  186.5 248.8 187.3 259.6 ;
      RECT  186.5 217.2 187.3 228.0 ;
      RECT  193.3 342.0 194.1 352.8 ;
      RECT  193.3 186.4 194.1 197.2 ;
      RECT  193.3 186.4 194.1 197.2 ;
      RECT  200.1 290.4 200.9 301.2 ;
      RECT  193.3 342.0 194.1 352.8 ;
      RECT  186.5 279.6 187.3 290.4 ;
      RECT  193.3 207.2 194.1 218.0 ;
      RECT  193.3 207.2 194.1 218.0 ;
      RECT  200.1 332.0 200.9 342.8 ;
      RECT  200.1 217.2 200.9 228.0 ;
      RECT  186.5 186.4 187.3 197.2 ;
      RECT  193.3 228.0 194.1 238.8 ;
      RECT  193.3 228.0 194.1 238.8 ;
      RECT  193.3 258.8 194.1 269.6 ;
      RECT  193.3 258.8 194.1 269.6 ;
      RECT  200.1 238.0 200.9 248.8 ;
      RECT  193.3 332.0 194.1 342.8 ;
      RECT  193.3 332.0 194.1 342.8 ;
      RECT  186.5 311.2 187.3 322.0 ;
      RECT  193.3 217.2 194.1 228.0 ;
      RECT  193.3 217.2 194.1 228.0 ;
      RECT  200.1 248.8 200.9 259.6 ;
      RECT  193.3 196.4 194.1 207.2 ;
      RECT  193.3 196.4 194.1 207.2 ;
      RECT  193.3 269.6 194.1 280.4 ;
      RECT  193.3 269.6 194.1 280.4 ;
      RECT  200.1 300.4 200.9 311.2 ;
      RECT  193.3 248.8 194.1 259.6 ;
      RECT  193.3 248.8 194.1 259.6 ;
      RECT  200.1 269.6 200.9 280.4 ;
      RECT  186.5 321.2 187.3 332.0 ;
      RECT  186.5 207.2 187.3 218.0 ;
      RECT  193.3 279.6 194.1 290.4 ;
      RECT  193.3 279.6 194.1 290.4 ;
      RECT  200.1 196.4 200.9 207.2 ;
      RECT  186.5 300.4 187.3 311.2 ;
      RECT  193.3 311.2 194.1 322.0 ;
      RECT  193.3 311.2 194.1 322.0 ;
      RECT  193.3 321.2 194.1 332.0 ;
      RECT  193.3 321.2 194.1 332.0 ;
      RECT  193.3 290.4 194.1 301.2 ;
      RECT  186.5 332.0 187.3 342.8 ;
      RECT  193.3 300.4 194.1 311.2 ;
      RECT  183.1 175.6 183.9 176.4 ;
      RECT  179.7 165.6 180.5 176.4 ;
      RECT  181.3 165.6 182.1 176.4 ;
      RECT  184.9 165.6 185.7 176.4 ;
      RECT  186.5 165.6 187.3 176.4 ;
      RECT  183.1 176.4 183.9 175.6 ;
      RECT  179.7 186.4 180.5 175.6 ;
      RECT  184.9 184.8 185.7 175.6 ;
      RECT  181.3 186.4 182.1 175.6 ;
      RECT  184.1 185.6 185.7 184.8 ;
      RECT  186.5 186.4 187.3 175.6 ;
      RECT  184.9 186.4 185.7 185.6 ;
      RECT  183.1 196.4 183.9 197.2 ;
      RECT  179.7 186.4 180.5 197.2 ;
      RECT  184.9 188.0 185.7 197.2 ;
      RECT  181.3 186.4 182.1 197.2 ;
      RECT  184.1 187.2 185.7 188.0 ;
      RECT  186.5 186.4 187.3 197.2 ;
      RECT  184.9 186.4 185.7 187.2 ;
      RECT  183.1 197.2 183.9 196.4 ;
      RECT  179.7 207.2 180.5 196.4 ;
      RECT  184.9 205.6 185.7 196.4 ;
      RECT  181.3 207.2 182.1 196.4 ;
      RECT  184.1 206.4 185.7 205.6 ;
      RECT  186.5 207.2 187.3 196.4 ;
      RECT  184.9 207.2 185.7 206.4 ;
      RECT  183.1 217.2 183.9 218.0 ;
      RECT  179.7 207.2 180.5 218.0 ;
      RECT  184.9 208.8 185.7 218.0 ;
      RECT  181.3 207.2 182.1 218.0 ;
      RECT  184.1 208.0 185.7 208.8 ;
      RECT  186.5 207.2 187.3 218.0 ;
      RECT  184.9 207.2 185.7 208.0 ;
      RECT  183.1 218.0 183.9 217.2 ;
      RECT  179.7 228.0 180.5 217.2 ;
      RECT  184.9 226.4 185.7 217.2 ;
      RECT  181.3 228.0 182.1 217.2 ;
      RECT  184.1 227.2 185.7 226.4 ;
      RECT  186.5 228.0 187.3 217.2 ;
      RECT  184.9 228.0 185.7 227.2 ;
      RECT  183.1 238.0 183.9 238.8 ;
      RECT  179.7 228.0 180.5 238.8 ;
      RECT  184.9 229.6 185.7 238.8 ;
      RECT  181.3 228.0 182.1 238.8 ;
      RECT  184.1 228.8 185.7 229.6 ;
      RECT  186.5 228.0 187.3 238.8 ;
      RECT  184.9 228.0 185.7 228.8 ;
      RECT  183.1 238.8 183.9 238.0 ;
      RECT  179.7 248.8 180.5 238.0 ;
      RECT  184.9 247.2 185.7 238.0 ;
      RECT  181.3 248.8 182.1 238.0 ;
      RECT  184.1 248.0 185.7 247.2 ;
      RECT  186.5 248.8 187.3 238.0 ;
      RECT  184.9 248.8 185.7 248.0 ;
      RECT  183.1 258.8 183.9 259.6 ;
      RECT  179.7 248.8 180.5 259.6 ;
      RECT  184.9 250.4 185.7 259.6 ;
      RECT  181.3 248.8 182.1 259.6 ;
      RECT  184.1 249.6 185.7 250.4 ;
      RECT  186.5 248.8 187.3 259.6 ;
      RECT  184.9 248.8 185.7 249.6 ;
      RECT  183.1 259.6 183.9 258.8 ;
      RECT  179.7 269.6 180.5 258.8 ;
      RECT  184.9 268.0 185.7 258.8 ;
      RECT  181.3 269.6 182.1 258.8 ;
      RECT  184.1 268.8 185.7 268.0 ;
      RECT  186.5 269.6 187.3 258.8 ;
      RECT  184.9 269.6 185.7 268.8 ;
      RECT  183.1 279.6 183.9 280.4 ;
      RECT  179.7 269.6 180.5 280.4 ;
      RECT  184.9 271.2 185.7 280.4 ;
      RECT  181.3 269.6 182.1 280.4 ;
      RECT  184.1 270.4 185.7 271.2 ;
      RECT  186.5 269.6 187.3 280.4 ;
      RECT  184.9 269.6 185.7 270.4 ;
      RECT  183.1 280.4 183.9 279.6 ;
      RECT  179.7 290.4 180.5 279.6 ;
      RECT  184.9 288.8 185.7 279.6 ;
      RECT  181.3 290.4 182.1 279.6 ;
      RECT  184.1 289.6 185.7 288.8 ;
      RECT  186.5 290.4 187.3 279.6 ;
      RECT  184.9 290.4 185.7 289.6 ;
      RECT  183.1 300.4 183.9 301.2 ;
      RECT  179.7 290.4 180.5 301.2 ;
      RECT  184.9 292.0 185.7 301.2 ;
      RECT  181.3 290.4 182.1 301.2 ;
      RECT  184.1 291.2 185.7 292.0 ;
      RECT  186.5 290.4 187.3 301.2 ;
      RECT  184.9 290.4 185.7 291.2 ;
      RECT  183.1 301.2 183.9 300.4 ;
      RECT  179.7 311.2 180.5 300.4 ;
      RECT  184.9 309.6 185.7 300.4 ;
      RECT  181.3 311.2 182.1 300.4 ;
      RECT  184.1 310.4 185.7 309.6 ;
      RECT  186.5 311.2 187.3 300.4 ;
      RECT  184.9 311.2 185.7 310.4 ;
      RECT  183.1 321.2 183.9 322.0 ;
      RECT  179.7 311.2 180.5 322.0 ;
      RECT  184.9 312.8 185.7 322.0 ;
      RECT  181.3 311.2 182.1 322.0 ;
      RECT  184.1 312.0 185.7 312.8 ;
      RECT  186.5 311.2 187.3 322.0 ;
      RECT  184.9 311.2 185.7 312.0 ;
      RECT  183.1 322.0 183.9 321.2 ;
      RECT  179.7 332.0 180.5 321.2 ;
      RECT  184.9 330.4 185.7 321.2 ;
      RECT  181.3 332.0 182.1 321.2 ;
      RECT  184.1 331.2 185.7 330.4 ;
      RECT  186.5 332.0 187.3 321.2 ;
      RECT  184.9 332.0 185.7 331.2 ;
      RECT  183.1 342.0 183.9 342.8 ;
      RECT  179.7 332.0 180.5 342.8 ;
      RECT  184.9 333.6 185.7 342.8 ;
      RECT  181.3 332.0 182.1 342.8 ;
      RECT  184.1 332.8 185.7 333.6 ;
      RECT  186.5 332.0 187.3 342.8 ;
      RECT  184.9 332.0 185.7 332.8 ;
      RECT  183.1 342.8 183.9 342.0 ;
      RECT  179.7 352.8 180.5 342.0 ;
      RECT  184.9 351.2 185.7 342.0 ;
      RECT  181.3 352.8 182.1 342.0 ;
      RECT  184.1 352.0 185.7 351.2 ;
      RECT  186.5 352.8 187.3 342.0 ;
      RECT  184.9 352.8 185.7 352.0 ;
      RECT  183.1 362.8 183.9 363.6 ;
      RECT  179.7 352.8 180.5 363.6 ;
      RECT  181.3 352.8 182.1 363.6 ;
      RECT  184.9 352.8 185.7 363.6 ;
      RECT  186.5 352.8 187.3 363.6 ;
      RECT  183.1 300.4 183.9 301.2 ;
      RECT  183.1 279.6 183.9 280.4 ;
      RECT  183.1 300.4 183.9 301.2 ;
      RECT  183.1 321.2 183.9 322.0 ;
      RECT  183.1 238.0 183.9 238.8 ;
      RECT  183.1 196.4 183.9 197.2 ;
      RECT  183.1 258.8 183.9 259.6 ;
      RECT  183.1 342.0 183.9 342.8 ;
      RECT  183.1 217.2 183.9 218.0 ;
      RECT  183.1 175.6 183.9 176.4 ;
      RECT  183.1 217.2 183.9 218.0 ;
      RECT  183.1 279.6 183.9 280.4 ;
      RECT  186.5 269.6 187.3 280.4 ;
      RECT  179.7 342.0 180.5 352.8 ;
      RECT  179.7 238.0 180.5 248.8 ;
      RECT  186.5 342.0 187.3 352.8 ;
      RECT  179.7 207.2 180.5 218.0 ;
      RECT  179.7 175.6 180.5 186.4 ;
      RECT  186.5 217.2 187.3 228.0 ;
      RECT  186.5 332.0 187.3 342.8 ;
      RECT  179.7 248.8 180.5 259.6 ;
      RECT  179.7 332.0 180.5 342.8 ;
      RECT  179.7 217.2 180.5 228.0 ;
      RECT  179.7 269.6 180.5 280.4 ;
      RECT  179.7 321.2 180.5 332.0 ;
      RECT  179.7 228.0 180.5 238.8 ;
      RECT  179.7 196.4 180.5 207.2 ;
      RECT  186.5 321.2 187.3 332.0 ;
      RECT  179.7 258.8 180.5 269.6 ;
      RECT  186.5 186.4 187.3 197.2 ;
      RECT  186.5 207.2 187.3 218.0 ;
      RECT  186.5 311.2 187.3 322.0 ;
      RECT  186.5 238.0 187.3 248.8 ;
      RECT  179.7 290.4 180.5 301.2 ;
      RECT  186.5 196.4 187.3 207.2 ;
      RECT  186.5 175.6 187.3 186.4 ;
      RECT  186.5 248.8 187.3 259.6 ;
      RECT  186.5 228.0 187.3 238.8 ;
      RECT  179.7 300.4 180.5 311.2 ;
      RECT  179.7 186.4 180.5 197.2 ;
      RECT  186.5 258.8 187.3 269.6 ;
      RECT  186.5 290.4 187.3 301.2 ;
      RECT  179.7 279.6 180.5 290.4 ;
      RECT  186.5 300.4 187.3 311.2 ;
      RECT  179.7 311.2 180.5 322.0 ;
      RECT  186.5 279.6 187.3 290.4 ;
      RECT  189.9 176.4 190.7 175.6 ;
      RECT  186.5 186.4 187.3 175.6 ;
      RECT  188.1 186.4 188.9 175.6 ;
      RECT  191.7 186.4 192.5 175.6 ;
      RECT  193.3 186.4 194.1 175.6 ;
      RECT  196.7 176.4 197.5 175.6 ;
      RECT  193.3 186.4 194.1 175.6 ;
      RECT  194.9 186.4 195.7 175.6 ;
      RECT  198.5 186.4 199.3 175.6 ;
      RECT  200.1 186.4 200.9 175.6 ;
      RECT  188.1 186.4 188.9 176.0 ;
      RECT  191.7 186.4 192.5 176.0 ;
      RECT  194.9 186.4 195.7 176.0 ;
      RECT  198.5 186.4 199.3 176.0 ;
      RECT  189.9 176.4 190.7 175.6 ;
      RECT  196.7 176.4 197.5 175.6 ;
      RECT  200.1 186.4 200.9 175.6 ;
      RECT  193.3 186.4 194.1 175.6 ;
      RECT  193.3 186.4 194.1 175.6 ;
      RECT  186.5 186.4 187.3 175.6 ;
      RECT  189.9 175.6 190.7 176.4 ;
      RECT  186.5 165.6 187.3 176.4 ;
      RECT  188.1 165.6 188.9 176.4 ;
      RECT  191.7 165.6 192.5 176.4 ;
      RECT  193.3 165.6 194.1 176.4 ;
      RECT  196.7 175.6 197.5 176.4 ;
      RECT  193.3 165.6 194.1 176.4 ;
      RECT  194.9 165.6 195.7 176.4 ;
      RECT  198.5 165.6 199.3 176.4 ;
      RECT  200.1 165.6 200.9 176.4 ;
      RECT  188.1 165.6 188.9 176.0 ;
      RECT  191.7 165.6 192.5 176.0 ;
      RECT  194.9 165.6 195.7 176.0 ;
      RECT  198.5 165.6 199.3 176.0 ;
      RECT  189.9 175.6 190.7 176.4 ;
      RECT  196.7 175.6 197.5 176.4 ;
      RECT  200.1 165.6 200.9 176.4 ;
      RECT  193.3 165.6 194.1 176.4 ;
      RECT  193.3 165.6 194.1 176.4 ;
      RECT  186.5 165.6 187.3 176.4 ;
      RECT  189.9 362.8 190.7 363.6 ;
      RECT  186.5 352.8 187.3 363.6 ;
      RECT  188.1 352.8 188.9 363.6 ;
      RECT  191.7 352.8 192.5 363.6 ;
      RECT  193.3 352.8 194.1 363.6 ;
      RECT  196.7 362.8 197.5 363.6 ;
      RECT  193.3 352.8 194.1 363.6 ;
      RECT  194.9 352.8 195.7 363.6 ;
      RECT  198.5 352.8 199.3 363.6 ;
      RECT  200.1 352.8 200.9 363.6 ;
      RECT  188.1 352.8 188.9 363.2 ;
      RECT  191.7 352.8 192.5 363.2 ;
      RECT  194.9 352.8 195.7 363.2 ;
      RECT  198.5 352.8 199.3 363.2 ;
      RECT  189.9 362.8 190.7 363.6 ;
      RECT  196.7 362.8 197.5 363.6 ;
      RECT  200.1 352.8 200.9 363.6 ;
      RECT  193.3 352.8 194.1 363.6 ;
      RECT  193.3 352.8 194.1 363.6 ;
      RECT  186.5 352.8 187.3 363.6 ;
      RECT  176.3 175.6 177.1 176.4 ;
      RECT  172.9 165.6 173.7 176.4 ;
      RECT  174.5 165.6 175.3 176.4 ;
      RECT  178.1 165.6 178.9 176.4 ;
      RECT  179.7 165.6 180.5 176.4 ;
      RECT  176.3 176.4 177.1 175.6 ;
      RECT  172.9 186.4 173.7 175.6 ;
      RECT  174.5 186.4 175.3 175.6 ;
      RECT  178.1 186.4 178.9 175.6 ;
      RECT  179.7 186.4 180.5 175.6 ;
      RECT  176.3 196.4 177.1 197.2 ;
      RECT  172.9 186.4 173.7 197.2 ;
      RECT  174.5 186.4 175.3 197.2 ;
      RECT  178.1 186.4 178.9 197.2 ;
      RECT  179.7 186.4 180.5 197.2 ;
      RECT  176.3 197.2 177.1 196.4 ;
      RECT  172.9 207.2 173.7 196.4 ;
      RECT  174.5 207.2 175.3 196.4 ;
      RECT  178.1 207.2 178.9 196.4 ;
      RECT  179.7 207.2 180.5 196.4 ;
      RECT  176.3 217.2 177.1 218.0 ;
      RECT  172.9 207.2 173.7 218.0 ;
      RECT  174.5 207.2 175.3 218.0 ;
      RECT  178.1 207.2 178.9 218.0 ;
      RECT  179.7 207.2 180.5 218.0 ;
      RECT  176.3 218.0 177.1 217.2 ;
      RECT  172.9 228.0 173.7 217.2 ;
      RECT  174.5 228.0 175.3 217.2 ;
      RECT  178.1 228.0 178.9 217.2 ;
      RECT  179.7 228.0 180.5 217.2 ;
      RECT  176.3 238.0 177.1 238.8 ;
      RECT  172.9 228.0 173.7 238.8 ;
      RECT  174.5 228.0 175.3 238.8 ;
      RECT  178.1 228.0 178.9 238.8 ;
      RECT  179.7 228.0 180.5 238.8 ;
      RECT  176.3 238.8 177.1 238.0 ;
      RECT  172.9 248.8 173.7 238.0 ;
      RECT  174.5 248.8 175.3 238.0 ;
      RECT  178.1 248.8 178.9 238.0 ;
      RECT  179.7 248.8 180.5 238.0 ;
      RECT  176.3 258.8 177.1 259.6 ;
      RECT  172.9 248.8 173.7 259.6 ;
      RECT  174.5 248.8 175.3 259.6 ;
      RECT  178.1 248.8 178.9 259.6 ;
      RECT  179.7 248.8 180.5 259.6 ;
      RECT  176.3 259.6 177.1 258.8 ;
      RECT  172.9 269.6 173.7 258.8 ;
      RECT  174.5 269.6 175.3 258.8 ;
      RECT  178.1 269.6 178.9 258.8 ;
      RECT  179.7 269.6 180.5 258.8 ;
      RECT  176.3 279.6 177.1 280.4 ;
      RECT  172.9 269.6 173.7 280.4 ;
      RECT  174.5 269.6 175.3 280.4 ;
      RECT  178.1 269.6 178.9 280.4 ;
      RECT  179.7 269.6 180.5 280.4 ;
      RECT  176.3 280.4 177.1 279.6 ;
      RECT  172.9 290.4 173.7 279.6 ;
      RECT  174.5 290.4 175.3 279.6 ;
      RECT  178.1 290.4 178.9 279.6 ;
      RECT  179.7 290.4 180.5 279.6 ;
      RECT  176.3 300.4 177.1 301.2 ;
      RECT  172.9 290.4 173.7 301.2 ;
      RECT  174.5 290.4 175.3 301.2 ;
      RECT  178.1 290.4 178.9 301.2 ;
      RECT  179.7 290.4 180.5 301.2 ;
      RECT  176.3 301.2 177.1 300.4 ;
      RECT  172.9 311.2 173.7 300.4 ;
      RECT  174.5 311.2 175.3 300.4 ;
      RECT  178.1 311.2 178.9 300.4 ;
      RECT  179.7 311.2 180.5 300.4 ;
      RECT  176.3 321.2 177.1 322.0 ;
      RECT  172.9 311.2 173.7 322.0 ;
      RECT  174.5 311.2 175.3 322.0 ;
      RECT  178.1 311.2 178.9 322.0 ;
      RECT  179.7 311.2 180.5 322.0 ;
      RECT  176.3 322.0 177.1 321.2 ;
      RECT  172.9 332.0 173.7 321.2 ;
      RECT  174.5 332.0 175.3 321.2 ;
      RECT  178.1 332.0 178.9 321.2 ;
      RECT  179.7 332.0 180.5 321.2 ;
      RECT  176.3 342.0 177.1 342.8 ;
      RECT  172.9 332.0 173.7 342.8 ;
      RECT  174.5 332.0 175.3 342.8 ;
      RECT  178.1 332.0 178.9 342.8 ;
      RECT  179.7 332.0 180.5 342.8 ;
      RECT  176.3 342.8 177.1 342.0 ;
      RECT  172.9 352.8 173.7 342.0 ;
      RECT  174.5 352.8 175.3 342.0 ;
      RECT  178.1 352.8 178.9 342.0 ;
      RECT  179.7 352.8 180.5 342.0 ;
      RECT  176.3 362.8 177.1 363.6 ;
      RECT  172.9 352.8 173.7 363.6 ;
      RECT  174.5 352.8 175.3 363.6 ;
      RECT  178.1 352.8 178.9 363.6 ;
      RECT  179.7 352.8 180.5 363.6 ;
      RECT  174.5 165.6 175.3 363.2 ;
      RECT  178.1 165.6 178.9 363.2 ;
      RECT  176.3 300.4 177.1 301.2 ;
      RECT  176.3 279.6 177.1 280.4 ;
      RECT  176.3 300.4 177.1 301.2 ;
      RECT  176.3 321.2 177.1 322.0 ;
      RECT  176.3 362.8 177.1 363.6 ;
      RECT  176.3 238.0 177.1 238.8 ;
      RECT  176.3 196.4 177.1 197.2 ;
      RECT  176.3 258.8 177.1 259.6 ;
      RECT  176.3 342.0 177.1 342.8 ;
      RECT  176.3 217.2 177.1 218.0 ;
      RECT  176.3 175.6 177.1 176.4 ;
      RECT  176.3 217.2 177.1 218.0 ;
      RECT  176.3 279.6 177.1 280.4 ;
      RECT  172.9 342.0 173.7 352.8 ;
      RECT  172.9 238.0 173.7 248.8 ;
      RECT  179.7 342.0 180.5 352.8 ;
      RECT  179.7 352.8 180.5 363.6 ;
      RECT  172.9 175.6 173.7 186.4 ;
      RECT  172.9 207.2 173.7 218.0 ;
      RECT  179.7 217.2 180.5 228.0 ;
      RECT  179.7 332.0 180.5 342.8 ;
      RECT  172.9 248.8 173.7 259.6 ;
      RECT  172.9 352.8 173.7 363.6 ;
      RECT  172.9 332.0 173.7 342.8 ;
      RECT  172.9 217.2 173.7 228.0 ;
      RECT  172.9 269.6 173.7 280.4 ;
      RECT  172.9 321.2 173.7 332.0 ;
      RECT  172.9 228.0 173.7 238.8 ;
      RECT  172.9 196.4 173.7 207.2 ;
      RECT  179.7 321.2 180.5 332.0 ;
      RECT  179.7 165.6 180.5 176.4 ;
      RECT  172.9 258.8 173.7 269.6 ;
      RECT  179.7 186.4 180.5 197.2 ;
      RECT  179.7 207.2 180.5 218.0 ;
      RECT  172.9 165.6 173.7 176.4 ;
      RECT  179.7 238.0 180.5 248.8 ;
      RECT  179.7 311.2 180.5 322.0 ;
      RECT  172.9 290.4 173.7 301.2 ;
      RECT  179.7 196.4 180.5 207.2 ;
      RECT  179.7 175.6 180.5 186.4 ;
      RECT  179.7 248.8 180.5 259.6 ;
      RECT  179.7 228.0 180.5 238.8 ;
      RECT  172.9 300.4 173.7 311.2 ;
      RECT  172.9 186.4 173.7 197.2 ;
      RECT  179.7 258.8 180.5 269.6 ;
      RECT  179.7 290.4 180.5 301.2 ;
      RECT  172.9 279.6 173.7 290.4 ;
      RECT  179.7 300.4 180.5 311.2 ;
      RECT  172.9 311.2 173.7 322.0 ;
      RECT  179.7 269.6 180.5 280.4 ;
      RECT  179.7 279.6 180.5 290.4 ;
      RECT  203.5 175.6 204.3 176.4 ;
      RECT  200.1 165.6 200.9 176.4 ;
      RECT  201.7 165.6 202.5 176.4 ;
      RECT  205.3 165.6 206.1 176.4 ;
      RECT  206.9 165.6 207.7 176.4 ;
      RECT  203.5 176.4 204.3 175.6 ;
      RECT  200.1 186.4 200.9 175.6 ;
      RECT  201.7 186.4 202.5 175.6 ;
      RECT  205.3 186.4 206.1 175.6 ;
      RECT  206.9 186.4 207.7 175.6 ;
      RECT  203.5 196.4 204.3 197.2 ;
      RECT  200.1 186.4 200.9 197.2 ;
      RECT  201.7 186.4 202.5 197.2 ;
      RECT  205.3 186.4 206.1 197.2 ;
      RECT  206.9 186.4 207.7 197.2 ;
      RECT  203.5 197.2 204.3 196.4 ;
      RECT  200.1 207.2 200.9 196.4 ;
      RECT  201.7 207.2 202.5 196.4 ;
      RECT  205.3 207.2 206.1 196.4 ;
      RECT  206.9 207.2 207.7 196.4 ;
      RECT  203.5 217.2 204.3 218.0 ;
      RECT  200.1 207.2 200.9 218.0 ;
      RECT  201.7 207.2 202.5 218.0 ;
      RECT  205.3 207.2 206.1 218.0 ;
      RECT  206.9 207.2 207.7 218.0 ;
      RECT  203.5 218.0 204.3 217.2 ;
      RECT  200.1 228.0 200.9 217.2 ;
      RECT  201.7 228.0 202.5 217.2 ;
      RECT  205.3 228.0 206.1 217.2 ;
      RECT  206.9 228.0 207.7 217.2 ;
      RECT  203.5 238.0 204.3 238.8 ;
      RECT  200.1 228.0 200.9 238.8 ;
      RECT  201.7 228.0 202.5 238.8 ;
      RECT  205.3 228.0 206.1 238.8 ;
      RECT  206.9 228.0 207.7 238.8 ;
      RECT  203.5 238.8 204.3 238.0 ;
      RECT  200.1 248.8 200.9 238.0 ;
      RECT  201.7 248.8 202.5 238.0 ;
      RECT  205.3 248.8 206.1 238.0 ;
      RECT  206.9 248.8 207.7 238.0 ;
      RECT  203.5 258.8 204.3 259.6 ;
      RECT  200.1 248.8 200.9 259.6 ;
      RECT  201.7 248.8 202.5 259.6 ;
      RECT  205.3 248.8 206.1 259.6 ;
      RECT  206.9 248.8 207.7 259.6 ;
      RECT  203.5 259.6 204.3 258.8 ;
      RECT  200.1 269.6 200.9 258.8 ;
      RECT  201.7 269.6 202.5 258.8 ;
      RECT  205.3 269.6 206.1 258.8 ;
      RECT  206.9 269.6 207.7 258.8 ;
      RECT  203.5 279.6 204.3 280.4 ;
      RECT  200.1 269.6 200.9 280.4 ;
      RECT  201.7 269.6 202.5 280.4 ;
      RECT  205.3 269.6 206.1 280.4 ;
      RECT  206.9 269.6 207.7 280.4 ;
      RECT  203.5 280.4 204.3 279.6 ;
      RECT  200.1 290.4 200.9 279.6 ;
      RECT  201.7 290.4 202.5 279.6 ;
      RECT  205.3 290.4 206.1 279.6 ;
      RECT  206.9 290.4 207.7 279.6 ;
      RECT  203.5 300.4 204.3 301.2 ;
      RECT  200.1 290.4 200.9 301.2 ;
      RECT  201.7 290.4 202.5 301.2 ;
      RECT  205.3 290.4 206.1 301.2 ;
      RECT  206.9 290.4 207.7 301.2 ;
      RECT  203.5 301.2 204.3 300.4 ;
      RECT  200.1 311.2 200.9 300.4 ;
      RECT  201.7 311.2 202.5 300.4 ;
      RECT  205.3 311.2 206.1 300.4 ;
      RECT  206.9 311.2 207.7 300.4 ;
      RECT  203.5 321.2 204.3 322.0 ;
      RECT  200.1 311.2 200.9 322.0 ;
      RECT  201.7 311.2 202.5 322.0 ;
      RECT  205.3 311.2 206.1 322.0 ;
      RECT  206.9 311.2 207.7 322.0 ;
      RECT  203.5 322.0 204.3 321.2 ;
      RECT  200.1 332.0 200.9 321.2 ;
      RECT  201.7 332.0 202.5 321.2 ;
      RECT  205.3 332.0 206.1 321.2 ;
      RECT  206.9 332.0 207.7 321.2 ;
      RECT  203.5 342.0 204.3 342.8 ;
      RECT  200.1 332.0 200.9 342.8 ;
      RECT  201.7 332.0 202.5 342.8 ;
      RECT  205.3 332.0 206.1 342.8 ;
      RECT  206.9 332.0 207.7 342.8 ;
      RECT  203.5 342.8 204.3 342.0 ;
      RECT  200.1 352.8 200.9 342.0 ;
      RECT  201.7 352.8 202.5 342.0 ;
      RECT  205.3 352.8 206.1 342.0 ;
      RECT  206.9 352.8 207.7 342.0 ;
      RECT  203.5 362.8 204.3 363.6 ;
      RECT  200.1 352.8 200.9 363.6 ;
      RECT  201.7 352.8 202.5 363.6 ;
      RECT  205.3 352.8 206.1 363.6 ;
      RECT  206.9 352.8 207.7 363.6 ;
      RECT  201.7 165.6 202.5 363.2 ;
      RECT  205.3 165.6 206.1 363.2 ;
      RECT  203.5 300.4 204.3 301.2 ;
      RECT  203.5 279.6 204.3 280.4 ;
      RECT  203.5 300.4 204.3 301.2 ;
      RECT  203.5 321.2 204.3 322.0 ;
      RECT  203.5 362.8 204.3 363.6 ;
      RECT  203.5 238.0 204.3 238.8 ;
      RECT  203.5 196.4 204.3 197.2 ;
      RECT  203.5 258.8 204.3 259.6 ;
      RECT  203.5 342.0 204.3 342.8 ;
      RECT  203.5 217.2 204.3 218.0 ;
      RECT  203.5 175.6 204.3 176.4 ;
      RECT  203.5 217.2 204.3 218.0 ;
      RECT  203.5 279.6 204.3 280.4 ;
      RECT  200.1 342.0 200.9 352.8 ;
      RECT  200.1 238.0 200.9 248.8 ;
      RECT  206.9 342.0 207.7 352.8 ;
      RECT  206.9 352.8 207.7 363.6 ;
      RECT  200.1 175.6 200.9 186.4 ;
      RECT  200.1 207.2 200.9 218.0 ;
      RECT  206.9 217.2 207.7 228.0 ;
      RECT  206.9 332.0 207.7 342.8 ;
      RECT  200.1 248.8 200.9 259.6 ;
      RECT  200.1 352.8 200.9 363.6 ;
      RECT  200.1 332.0 200.9 342.8 ;
      RECT  200.1 217.2 200.9 228.0 ;
      RECT  200.1 269.6 200.9 280.4 ;
      RECT  200.1 321.2 200.9 332.0 ;
      RECT  200.1 228.0 200.9 238.8 ;
      RECT  200.1 196.4 200.9 207.2 ;
      RECT  206.9 321.2 207.7 332.0 ;
      RECT  206.9 165.6 207.7 176.4 ;
      RECT  200.1 258.8 200.9 269.6 ;
      RECT  206.9 186.4 207.7 197.2 ;
      RECT  206.9 207.2 207.7 218.0 ;
      RECT  200.1 165.6 200.9 176.4 ;
      RECT  206.9 238.0 207.7 248.8 ;
      RECT  206.9 311.2 207.7 322.0 ;
      RECT  200.1 290.4 200.9 301.2 ;
      RECT  206.9 196.4 207.7 207.2 ;
      RECT  206.9 175.6 207.7 186.4 ;
      RECT  206.9 248.8 207.7 259.6 ;
      RECT  206.9 228.0 207.7 238.8 ;
      RECT  200.1 300.4 200.9 311.2 ;
      RECT  200.1 186.4 200.9 197.2 ;
      RECT  206.9 258.8 207.7 269.6 ;
      RECT  206.9 290.4 207.7 301.2 ;
      RECT  200.1 279.6 200.9 290.4 ;
      RECT  206.9 300.4 207.7 311.2 ;
      RECT  200.1 311.2 200.9 322.0 ;
      RECT  206.9 269.6 207.7 280.4 ;
      RECT  206.9 279.6 207.7 290.4 ;
      RECT  181.3 165.6 182.1 363.2 ;
      RECT  184.9 165.6 185.7 363.2 ;
      RECT  188.1 165.6 188.9 363.2 ;
      RECT  191.7 165.6 192.5 363.2 ;
      RECT  194.9 165.6 195.7 363.2 ;
      RECT  198.5 165.6 199.3 363.2 ;
      RECT  183.1 175.6 183.9 176.4 ;
      RECT  183.1 279.6 183.9 280.4 ;
      RECT  183.1 321.2 183.9 322.0 ;
      RECT  183.1 217.2 183.9 218.0 ;
      RECT  183.1 342.0 183.9 342.8 ;
      RECT  183.1 196.4 183.9 197.2 ;
      RECT  183.1 238.0 183.9 238.8 ;
      RECT  183.1 300.4 183.9 301.2 ;
      RECT  183.1 258.8 183.9 259.6 ;
      RECT  179.7 342.0 180.5 352.8 ;
      RECT  179.7 217.2 180.5 228.0 ;
      RECT  186.5 207.2 187.3 218.0 ;
      RECT  186.5 311.2 187.3 322.0 ;
      RECT  179.7 238.0 180.5 248.8 ;
      RECT  186.5 196.4 187.3 207.2 ;
      RECT  179.7 196.4 180.5 207.2 ;
      RECT  186.5 279.6 187.3 290.4 ;
      RECT  186.5 248.8 187.3 259.6 ;
      RECT  179.7 290.4 180.5 301.2 ;
      RECT  179.7 269.6 180.5 280.4 ;
      RECT  186.5 332.0 187.3 342.8 ;
      RECT  179.7 186.4 180.5 197.2 ;
      RECT  186.5 217.2 187.3 228.0 ;
      RECT  179.7 175.6 180.5 186.4 ;
      RECT  186.5 342.0 187.3 352.8 ;
      RECT  179.7 228.0 180.5 238.8 ;
      RECT  186.5 300.4 187.3 311.2 ;
      RECT  179.7 258.8 180.5 269.6 ;
      RECT  186.5 186.4 187.3 197.2 ;
      RECT  186.5 258.8 187.3 269.6 ;
      RECT  179.7 332.0 180.5 342.8 ;
      RECT  186.5 290.4 187.3 301.2 ;
      RECT  179.7 248.8 180.5 259.6 ;
      RECT  186.5 321.2 187.3 332.0 ;
      RECT  186.5 238.0 187.3 248.8 ;
      RECT  179.7 321.2 180.5 332.0 ;
      RECT  186.5 269.6 187.3 280.4 ;
      RECT  179.7 207.2 180.5 218.0 ;
      RECT  179.7 311.2 180.5 322.0 ;
      RECT  186.5 228.0 187.3 238.8 ;
      RECT  179.7 300.4 180.5 311.2 ;
      RECT  186.5 175.6 187.3 186.4 ;
      RECT  179.7 279.6 180.5 290.4 ;
      RECT  181.2 149.4 181.8 161.4 ;
      RECT  185.2 149.4 185.8 161.4 ;
      RECT  188.0 149.4 188.6 161.4 ;
      RECT  192.0 149.4 192.6 161.4 ;
      RECT  194.8 149.4 195.4 161.4 ;
      RECT  198.8 149.4 199.4 161.4 ;
      RECT  181.2 149.4 181.8 161.4 ;
      RECT  185.2 149.4 185.8 161.4 ;
      RECT  188.0 149.4 188.6 161.4 ;
      RECT  192.0 149.4 192.6 161.4 ;
      RECT  194.8 149.4 195.4 161.4 ;
      RECT  198.8 149.4 199.4 161.4 ;
      RECT  188.9 122.2 189.7 145.2 ;
      RECT  190.9 122.2 191.7 145.2 ;
      RECT  190.9 112.6 191.7 121.4 ;
      RECT  187.5 112.6 188.3 115.6 ;
      RECT  193.3 138.4 194.1 140.0 ;
      RECT  190.9 121.4 192.1 122.2 ;
      RECT  188.9 112.6 189.7 121.4 ;
      RECT  192.3 125.0 193.1 126.6 ;
      RECT  188.9 121.4 190.3 122.2 ;
      RECT  195.7 122.2 196.5 145.2 ;
      RECT  197.7 122.2 198.5 145.2 ;
      RECT  197.7 112.6 198.5 121.4 ;
      RECT  194.3 112.6 195.1 115.6 ;
      RECT  200.1 138.4 200.9 140.0 ;
      RECT  197.7 121.4 198.9 122.2 ;
      RECT  195.7 112.6 196.5 121.4 ;
      RECT  199.1 125.0 199.9 126.6 ;
      RECT  195.7 121.4 197.1 122.2 ;
      RECT  187.5 112.6 188.3 115.6 ;
      RECT  188.9 122.2 189.7 145.2 ;
      RECT  190.9 122.2 191.7 145.2 ;
      RECT  194.3 112.6 195.1 115.6 ;
      RECT  195.7 122.2 196.5 145.2 ;
      RECT  197.7 122.2 198.5 145.2 ;
      RECT  190.9 103.4 191.7 108.4 ;
      RECT  192.1 85.0 192.9 85.8 ;
      RECT  190.7 80.6 191.5 81.4 ;
      RECT  188.9 106.4 189.7 108.4 ;
      RECT  189.3 99.6 190.1 100.4 ;
      RECT  190.1 91.4 190.9 92.2 ;
      RECT  189.9 67.8 190.7 69.8 ;
      RECT  190.7 74.0 191.5 74.8 ;
      RECT  197.7 103.4 198.5 108.4 ;
      RECT  198.9 85.0 199.7 85.8 ;
      RECT  197.5 80.6 198.3 81.4 ;
      RECT  195.7 106.4 196.5 108.4 ;
      RECT  196.1 99.6 196.9 100.4 ;
      RECT  196.9 91.4 197.7 92.2 ;
      RECT  196.7 67.8 197.5 69.8 ;
      RECT  197.5 74.0 198.3 74.8 ;
      RECT  189.9 67.8 190.7 69.8 ;
      RECT  196.7 67.8 197.5 69.8 ;
      RECT  188.9 106.4 189.7 108.4 ;
      RECT  190.9 103.4 191.7 108.4 ;
      RECT  195.7 106.4 196.5 108.4 ;
      RECT  197.7 103.4 198.5 108.4 ;
      RECT  181.2 161.4 181.8 149.4 ;
      RECT  185.2 161.4 185.8 149.4 ;
      RECT  188.0 161.4 188.6 149.4 ;
      RECT  192.0 161.4 192.6 149.4 ;
      RECT  194.8 161.4 195.4 149.4 ;
      RECT  198.8 161.4 199.4 149.4 ;
      RECT  187.5 115.6 188.3 112.6 ;
      RECT  194.3 115.6 195.1 112.6 ;
      RECT  189.9 69.8 190.7 67.8 ;
      RECT  196.7 69.8 197.5 67.8 ;
      RECT  89.8 191.4 90.6 192.2 ;
      RECT  91.2 202.2 92.0 203.0 ;
      RECT  89.8 253.8 90.6 254.6 ;
      RECT  91.2 264.6 92.0 265.4 ;
      RECT  82.3 186.8 82.9 290.8 ;
      RECT  83.7 186.8 84.3 290.8 ;
      RECT  85.1 186.8 85.7 290.8 ;
      RECT  86.5 186.8 87.1 290.8 ;
      RECT  156.9 186.8 157.5 353.2 ;
      RECT  82.3 186.8 82.9 290.8 ;
      RECT  83.7 186.8 84.3 290.8 ;
      RECT  85.1 186.8 85.7 290.8 ;
      RECT  86.5 186.8 87.1 290.8 ;
      RECT  156.9 186.8 157.5 353.2 ;
      RECT  187.5 112.6 188.3 115.6 ;
      RECT  194.3 112.6 195.1 115.6 ;
      RECT  189.9 67.8 190.7 69.8 ;
      RECT  196.7 67.8 197.5 69.8 ;
      RECT  82.3 186.8 82.9 290.8 ;
      RECT  83.7 186.8 84.3 290.8 ;
      RECT  85.1 186.8 85.7 290.8 ;
      RECT  86.5 186.8 87.1 290.8 ;
      RECT  164.9 67.8 165.5 183.6 ;
      RECT  167.7 67.8 168.3 183.6 ;
      RECT  166.3 67.8 166.9 183.6 ;
      RECT  169.1 67.8 169.7 183.6 ;
      RECT  10.0 11.4 10.8 12.2 ;
      RECT  21.2 12.2 22.0 13.0 ;
      RECT  5.2 9.4 6.0 10.2 ;
      RECT  3.6 8.0 4.4 13.6 ;
      RECT  6.8 6.0 7.6 17.6 ;
      RECT  16.4 6.0 17.2 17.6 ;
      RECT  10.0 11.4 10.8 12.2 ;
      RECT  38.2 8.9 38.8 9.5 ;
      RECT  32.6 14.9 33.2 15.5 ;
      RECT  5.2 9.4 6.0 10.2 ;
      RECT  10.0 34.2 10.8 33.4 ;
      RECT  21.2 33.4 22.0 32.6 ;
      RECT  5.2 36.2 6.0 35.4 ;
      RECT  3.6 37.6 4.4 32.0 ;
      RECT  6.8 39.6 7.6 28.0 ;
      RECT  16.4 39.6 17.2 28.0 ;
      RECT  10.0 34.2 10.8 33.4 ;
      RECT  38.2 36.7 38.8 36.1 ;
      RECT  32.6 30.7 33.2 30.1 ;
      RECT  5.2 36.2 6.0 35.4 ;
      RECT  10.0 11.4 10.8 12.2 ;
      RECT  10.0 33.4 10.8 34.2 ;
      RECT  38.2 8.9 38.8 9.5 ;
      RECT  32.6 14.9 33.2 15.5 ;
      RECT  38.2 36.1 38.8 36.7 ;
      RECT  32.6 30.1 33.2 30.7 ;
      RECT  5.2 2.8 5.8 42.8 ;
      RECT  33.8 165.6 33.2 175.2 ;
      RECT  5.5 165.6 4.9 332.0 ;
      RECT  10.0 11.4 10.8 12.2 ;
      RECT  10.0 33.4 10.8 34.2 ;
      RECT  54.1 12.3 54.7 12.9 ;
      RECT  33.2 165.6 33.8 175.2 ;
      RECT  65.9 152.9 79.4 153.5 ;
      RECT  65.7 91.5 79.4 92.1 ;
      RECT  71.5 112.7 79.4 113.3 ;
      RECT  73.3 73.5 79.4 74.1 ;
      RECT  74.8 11.5 79.4 12.1 ;
      RECT  65.2 353.4 66.0 354.2 ;
      RECT  76.4 354.2 77.2 355.0 ;
      RECT  60.4 351.4 61.2 352.2 ;
      RECT  58.8 350.0 59.6 355.6 ;
      RECT  62.0 348.0 62.8 359.6 ;
      RECT  71.6 348.0 72.4 359.6 ;
      RECT  65.2 376.2 66.0 375.4 ;
      RECT  76.4 375.4 77.2 374.6 ;
      RECT  60.4 378.2 61.2 377.4 ;
      RECT  58.8 379.6 59.6 374.0 ;
      RECT  62.0 381.6 62.8 370.0 ;
      RECT  71.6 381.6 72.4 370.0 ;
      RECT  65.2 393.4 66.0 394.2 ;
      RECT  76.4 394.2 77.2 395.0 ;
      RECT  60.4 391.4 61.2 392.2 ;
      RECT  58.8 390.0 59.6 395.6 ;
      RECT  62.0 388.0 62.8 399.6 ;
      RECT  71.6 388.0 72.4 399.6 ;
      RECT  65.2 416.2 66.0 415.4 ;
      RECT  76.4 415.4 77.2 414.6 ;
      RECT  60.4 418.2 61.2 417.4 ;
      RECT  58.8 419.6 59.6 414.0 ;
      RECT  62.0 421.6 62.8 410.0 ;
      RECT  71.6 421.6 72.4 410.0 ;
      RECT  65.2 353.4 66.0 354.2 ;
      RECT  65.2 375.4 66.0 376.2 ;
      RECT  65.2 393.4 66.0 394.2 ;
      RECT  65.2 415.4 66.0 416.2 ;
      RECT  76.4 354.2 77.2 355.0 ;
      RECT  76.4 374.6 77.2 375.4 ;
      RECT  76.4 394.2 77.2 395.0 ;
      RECT  76.4 414.6 77.2 415.4 ;
      RECT  108.8 11.4 109.6 12.2 ;
      RECT  120.0 12.2 120.8 13.0 ;
      RECT  104.0 9.4 104.8 10.2 ;
      RECT  102.4 8.0 103.2 13.6 ;
      RECT  105.6 6.0 106.4 17.6 ;
      RECT  115.2 6.0 116.0 17.6 ;
      RECT  130.6 11.4 131.4 12.2 ;
      RECT  141.8 12.2 142.6 13.0 ;
      RECT  125.8 9.4 126.6 10.2 ;
      RECT  124.2 8.0 125.0 13.6 ;
      RECT  127.4 6.0 128.2 17.6 ;
      RECT  137.0 6.0 137.8 17.6 ;
      RECT  108.8 11.4 109.6 12.2 ;
      RECT  130.6 11.4 131.4 12.2 ;
      RECT  120.0 12.2 120.8 13.0 ;
      RECT  141.8 12.2 142.6 13.0 ;
   LAYER  m3 ;
      RECT  183.1 175.6 183.9 176.4 ;
      RECT  183.1 362.8 183.9 363.6 ;
      RECT  186.5 357.8 187.3 358.6 ;
      RECT  179.7 357.8 180.5 358.6 ;
      RECT  186.5 170.6 187.3 171.4 ;
      RECT  179.7 170.6 180.5 171.4 ;
      RECT  203.5 279.6 204.3 280.4 ;
      RECT  183.1 175.6 183.9 176.4 ;
      RECT  176.3 238.0 177.1 238.8 ;
      RECT  203.5 342.0 204.3 342.8 ;
      RECT  176.3 217.2 177.1 218.0 ;
      RECT  176.3 175.6 177.1 176.4 ;
      RECT  176.3 362.8 177.1 363.6 ;
      RECT  196.7 175.6 197.5 176.4 ;
      RECT  203.5 300.4 204.3 301.2 ;
      RECT  176.3 321.2 177.1 322.0 ;
      RECT  176.3 279.6 177.1 280.4 ;
      RECT  176.3 258.8 177.1 259.6 ;
      RECT  176.3 196.4 177.1 197.2 ;
      RECT  203.5 362.8 204.3 363.6 ;
      RECT  196.7 362.8 197.5 363.6 ;
      RECT  203.5 258.8 204.3 259.6 ;
      RECT  189.9 362.8 190.7 363.6 ;
      RECT  203.5 321.2 204.3 322.0 ;
      RECT  203.5 175.6 204.3 176.4 ;
      RECT  203.5 196.4 204.3 197.2 ;
      RECT  176.3 342.0 177.1 342.8 ;
      RECT  203.5 238.0 204.3 238.8 ;
      RECT  203.5 217.2 204.3 218.0 ;
      RECT  183.1 362.8 183.9 363.6 ;
      RECT  176.3 300.4 177.1 301.2 ;
      RECT  189.9 175.6 190.7 176.4 ;
      RECT  200.1 305.4 200.9 306.2 ;
      RECT  200.1 274.6 200.9 275.4 ;
      RECT  206.9 284.6 207.7 285.4 ;
      RECT  179.7 326.2 180.5 327.0 ;
      RECT  200.1 263.8 200.9 264.6 ;
      RECT  179.7 337.0 180.5 337.8 ;
      RECT  179.7 191.4 180.5 192.2 ;
      RECT  206.9 263.8 207.7 264.6 ;
      RECT  179.7 274.6 180.5 275.4 ;
      RECT  200.1 284.6 200.9 285.4 ;
      RECT  193.3 170.6 194.1 171.4 ;
      RECT  179.7 347.0 180.5 347.8 ;
      RECT  200.1 191.4 200.9 192.2 ;
      RECT  200.1 295.4 200.9 296.2 ;
      RECT  179.7 233.0 180.5 233.8 ;
      RECT  172.9 253.8 173.7 254.6 ;
      RECT  179.7 316.2 180.5 317.0 ;
      RECT  206.9 357.8 207.7 358.6 ;
      RECT  200.1 243.0 200.9 243.8 ;
      RECT  200.1 326.2 200.9 327.0 ;
      RECT  206.9 347.0 207.7 347.8 ;
      RECT  200.1 347.0 200.9 347.8 ;
      RECT  206.9 295.4 207.7 296.2 ;
      RECT  179.7 201.4 180.5 202.2 ;
      RECT  172.9 212.2 173.7 213.0 ;
      RECT  172.9 326.2 173.7 327.0 ;
      RECT  172.9 305.4 173.7 306.2 ;
      RECT  179.7 263.8 180.5 264.6 ;
      RECT  179.7 357.8 180.5 358.6 ;
      RECT  179.7 357.8 180.5 358.6 ;
      RECT  193.3 357.8 194.1 358.6 ;
      RECT  172.9 295.4 173.7 296.2 ;
      RECT  186.5 357.8 187.3 358.6 ;
      RECT  186.5 357.8 187.3 358.6 ;
      RECT  179.7 212.2 180.5 213.0 ;
      RECT  206.9 191.4 207.7 192.2 ;
      RECT  200.1 201.4 200.9 202.2 ;
      RECT  172.9 284.6 173.7 285.4 ;
      RECT  206.9 337.0 207.7 337.8 ;
      RECT  206.9 222.2 207.7 223.0 ;
      RECT  206.9 243.0 207.7 243.8 ;
      RECT  172.9 201.4 173.7 202.2 ;
      RECT  206.9 274.6 207.7 275.4 ;
      RECT  179.7 295.4 180.5 296.2 ;
      RECT  172.9 337.0 173.7 337.8 ;
      RECT  172.9 263.8 173.7 264.6 ;
      RECT  206.9 180.6 207.7 181.4 ;
      RECT  206.9 201.4 207.7 202.2 ;
      RECT  179.7 180.6 180.5 181.4 ;
      RECT  179.7 253.8 180.5 254.6 ;
      RECT  200.1 180.6 200.9 181.4 ;
      RECT  172.9 180.6 173.7 181.4 ;
      RECT  172.9 274.6 173.7 275.4 ;
      RECT  172.9 357.8 173.7 358.6 ;
      RECT  200.1 357.8 200.9 358.6 ;
      RECT  172.9 233.0 173.7 233.8 ;
      RECT  172.9 191.4 173.7 192.2 ;
      RECT  200.1 212.2 200.9 213.0 ;
      RECT  179.7 222.2 180.5 223.0 ;
      RECT  206.9 326.2 207.7 327.0 ;
      RECT  172.9 347.0 173.7 347.8 ;
      RECT  179.7 243.0 180.5 243.8 ;
      RECT  172.9 316.2 173.7 317.0 ;
      RECT  200.1 170.6 200.9 171.4 ;
      RECT  200.1 253.8 200.9 254.6 ;
      RECT  200.1 337.0 200.9 337.8 ;
      RECT  206.9 305.4 207.7 306.2 ;
      RECT  172.9 222.2 173.7 223.0 ;
      RECT  206.9 253.8 207.7 254.6 ;
      RECT  206.9 316.2 207.7 317.0 ;
      RECT  206.9 212.2 207.7 213.0 ;
      RECT  179.7 284.6 180.5 285.4 ;
      RECT  179.7 305.4 180.5 306.2 ;
      RECT  186.5 170.6 187.3 171.4 ;
      RECT  186.5 170.6 187.3 171.4 ;
      RECT  200.1 233.0 200.9 233.8 ;
      RECT  206.9 170.6 207.7 171.4 ;
      RECT  200.1 316.2 200.9 317.0 ;
      RECT  179.7 170.6 180.5 171.4 ;
      RECT  179.7 170.6 180.5 171.4 ;
      RECT  172.9 243.0 173.7 243.8 ;
      RECT  200.1 222.2 200.9 223.0 ;
      RECT  206.9 233.0 207.7 233.8 ;
      RECT  172.9 170.6 173.7 171.4 ;
      RECT  183.6 159.6 184.4 160.4 ;
      RECT  190.4 159.6 191.2 160.4 ;
      RECT  197.2 159.6 198.0 160.4 ;
      RECT  190.4 159.6 191.2 160.4 ;
      RECT  183.6 159.6 184.4 160.4 ;
      RECT  197.2 159.6 198.0 160.4 ;
      RECT  192.3 125.4 193.1 126.2 ;
      RECT  199.1 125.4 199.9 126.2 ;
      RECT  193.3 138.8 194.1 139.6 ;
      RECT  200.1 138.8 200.9 139.6 ;
      RECT  196.9 91.4 197.7 92.2 ;
      RECT  197.5 74.0 198.3 74.8 ;
      RECT  190.1 91.4 190.9 92.2 ;
      RECT  190.7 74.0 191.5 74.8 ;
      RECT  190.7 80.6 191.5 81.4 ;
      RECT  189.3 99.6 190.1 100.4 ;
      RECT  198.9 85.0 199.7 85.8 ;
      RECT  196.1 99.6 196.9 100.4 ;
      RECT  197.5 80.6 198.3 81.4 ;
      RECT  192.1 85.0 192.9 85.8 ;
      RECT  190.4 160.4 191.2 159.6 ;
      RECT  199.1 126.2 199.9 125.4 ;
      RECT  190.1 92.2 190.9 91.4 ;
      RECT  197.2 160.4 198.0 159.6 ;
      RECT  190.7 74.8 191.5 74.0 ;
      RECT  196.9 92.2 197.7 91.4 ;
      RECT  183.6 160.4 184.4 159.6 ;
      RECT  192.3 126.2 193.1 125.4 ;
      RECT  197.5 74.8 198.3 74.0 ;
      RECT  193.3 139.6 194.1 138.8 ;
      RECT  189.3 100.4 190.1 99.6 ;
      RECT  197.5 81.4 198.3 80.6 ;
      RECT  190.7 81.4 191.5 80.6 ;
      RECT  192.1 85.8 192.9 85.0 ;
      RECT  196.1 100.4 196.9 99.6 ;
      RECT  198.9 85.8 199.7 85.0 ;
      RECT  200.1 139.6 200.9 138.8 ;
      RECT  93.1 217.6 93.9 218.4 ;
      RECT  93.1 217.6 93.9 218.4 ;
      RECT  93.1 196.8 93.9 197.6 ;
      RECT  93.1 196.8 93.9 197.6 ;
      RECT  108.1 217.6 108.9 218.4 ;
      RECT  108.1 196.8 108.9 197.6 ;
      RECT  108.1 196.8 108.9 197.6 ;
      RECT  108.1 217.6 108.9 218.4 ;
      RECT  108.1 228.0 108.9 228.8 ;
      RECT  93.1 186.4 93.9 187.2 ;
      RECT  108.1 207.2 108.9 208.0 ;
      RECT  108.1 186.4 108.9 187.2 ;
      RECT  93.1 228.0 93.9 228.8 ;
      RECT  93.1 207.2 93.9 208.0 ;
      RECT  93.1 280.0 93.9 280.8 ;
      RECT  93.1 280.0 93.9 280.8 ;
      RECT  93.1 259.2 93.9 260.0 ;
      RECT  93.1 259.2 93.9 260.0 ;
      RECT  108.1 280.0 108.9 280.8 ;
      RECT  108.1 259.2 108.9 260.0 ;
      RECT  108.1 259.2 108.9 260.0 ;
      RECT  108.1 280.0 108.9 280.8 ;
      RECT  108.1 290.4 108.9 291.2 ;
      RECT  93.1 248.8 93.9 249.6 ;
      RECT  108.1 269.6 108.9 270.4 ;
      RECT  108.1 248.8 108.9 249.6 ;
      RECT  93.1 290.4 93.9 291.2 ;
      RECT  93.1 269.6 93.9 270.4 ;
      RECT  108.1 259.2 108.9 260.0 ;
      RECT  152.0 321.6 152.8 322.4 ;
      RECT  152.0 280.0 152.8 280.8 ;
      RECT  152.0 280.0 152.8 280.8 ;
      RECT  108.1 217.6 108.9 218.4 ;
      RECT  152.0 238.4 152.8 239.2 ;
      RECT  93.1 259.2 93.9 260.0 ;
      RECT  108.1 280.0 108.9 280.8 ;
      RECT  152.0 259.2 152.8 260.0 ;
      RECT  152.0 259.2 152.8 260.0 ;
      RECT  152.0 300.8 152.8 301.6 ;
      RECT  108.1 196.8 108.9 197.6 ;
      RECT  93.1 280.0 93.9 280.8 ;
      RECT  152.0 196.8 152.8 197.6 ;
      RECT  152.0 196.8 152.8 197.6 ;
      RECT  93.1 217.6 93.9 218.4 ;
      RECT  152.0 217.6 152.8 218.4 ;
      RECT  152.0 217.6 152.8 218.4 ;
      RECT  93.1 196.8 93.9 197.6 ;
      RECT  152.0 342.4 152.8 343.2 ;
      RECT  152.0 269.6 152.8 270.4 ;
      RECT  152.0 311.2 152.8 312.0 ;
      RECT  152.0 228.0 152.8 228.8 ;
      RECT  93.1 207.2 93.9 208.0 ;
      RECT  93.1 248.8 93.9 249.6 ;
      RECT  152.0 352.8 152.8 353.6 ;
      RECT  152.0 290.4 152.8 291.2 ;
      RECT  152.0 332.0 152.8 332.8 ;
      RECT  108.1 248.8 108.9 249.6 ;
      RECT  93.1 290.4 93.9 291.2 ;
      RECT  108.1 228.0 108.9 228.8 ;
      RECT  108.1 207.2 108.9 208.0 ;
      RECT  93.1 269.6 93.9 270.4 ;
      RECT  108.1 186.4 108.9 187.2 ;
      RECT  93.1 186.4 93.9 187.2 ;
      RECT  152.0 207.2 152.8 208.0 ;
      RECT  152.0 186.4 152.8 187.2 ;
      RECT  108.1 269.6 108.9 270.4 ;
      RECT  152.0 248.8 152.8 249.6 ;
      RECT  108.1 290.4 108.9 291.2 ;
      RECT  93.1 228.0 93.9 228.8 ;
      RECT  167.5 217.6 168.3 218.4 ;
      RECT  167.5 196.8 168.3 197.6 ;
      RECT  167.5 217.6 168.3 218.4 ;
      RECT  167.5 196.8 168.3 197.6 ;
      RECT  167.5 321.6 168.3 322.4 ;
      RECT  167.5 342.4 168.3 343.2 ;
      RECT  167.5 280.0 168.3 280.8 ;
      RECT  167.5 280.0 168.3 280.8 ;
      RECT  167.5 259.2 168.3 260.0 ;
      RECT  167.5 259.2 168.3 260.0 ;
      RECT  167.5 300.8 168.3 301.6 ;
      RECT  167.5 238.4 168.3 239.2 ;
      RECT  167.5 269.6 168.3 270.4 ;
      RECT  167.5 332.0 168.3 332.8 ;
      RECT  167.5 207.2 168.3 208.0 ;
      RECT  167.5 248.8 168.3 249.6 ;
      RECT  167.5 186.4 168.3 187.2 ;
      RECT  167.5 352.8 168.3 353.6 ;
      RECT  167.5 290.4 168.3 291.2 ;
      RECT  167.5 311.2 168.3 312.0 ;
      RECT  167.5 228.0 168.3 228.8 ;
      RECT  167.5 321.6 168.3 322.4 ;
      RECT  167.5 342.4 168.3 343.2 ;
      RECT  152.0 217.6 152.8 218.4 ;
      RECT  152.0 259.2 152.8 260.0 ;
      RECT  108.1 280.0 108.9 280.8 ;
      RECT  152.0 342.4 152.8 343.2 ;
      RECT  108.1 196.8 108.9 197.6 ;
      RECT  108.1 217.6 108.9 218.4 ;
      RECT  167.5 300.8 168.3 301.6 ;
      RECT  167.5 238.4 168.3 239.2 ;
      RECT  152.0 196.8 152.8 197.6 ;
      RECT  152.0 238.4 152.8 239.2 ;
      RECT  167.5 196.8 168.3 197.6 ;
      RECT  93.1 280.0 93.9 280.8 ;
      RECT  167.5 217.6 168.3 218.4 ;
      RECT  152.0 280.0 152.8 280.8 ;
      RECT  167.5 259.2 168.3 260.0 ;
      RECT  152.0 300.8 152.8 301.6 ;
      RECT  93.1 196.8 93.9 197.6 ;
      RECT  152.0 321.6 152.8 322.4 ;
      RECT  93.1 259.2 93.9 260.0 ;
      RECT  108.1 259.2 108.9 260.0 ;
      RECT  93.1 217.6 93.9 218.4 ;
      RECT  167.5 280.0 168.3 280.8 ;
      RECT  167.5 311.2 168.3 312.0 ;
      RECT  152.0 207.2 152.8 208.0 ;
      RECT  167.5 269.6 168.3 270.4 ;
      RECT  108.1 207.2 108.9 208.0 ;
      RECT  167.5 207.2 168.3 208.0 ;
      RECT  152.0 186.4 152.8 187.2 ;
      RECT  93.1 248.8 93.9 249.6 ;
      RECT  152.0 228.0 152.8 228.8 ;
      RECT  152.0 290.4 152.8 291.2 ;
      RECT  93.1 207.2 93.9 208.0 ;
      RECT  167.5 228.0 168.3 228.8 ;
      RECT  167.5 290.4 168.3 291.2 ;
      RECT  93.1 290.4 93.9 291.2 ;
      RECT  152.0 352.8 152.8 353.6 ;
      RECT  167.5 332.0 168.3 332.8 ;
      RECT  167.5 248.8 168.3 249.6 ;
      RECT  108.1 186.4 108.9 187.2 ;
      RECT  93.1 269.6 93.9 270.4 ;
      RECT  152.0 311.2 152.8 312.0 ;
      RECT  108.1 248.8 108.9 249.6 ;
      RECT  152.0 248.8 152.8 249.6 ;
      RECT  108.1 290.4 108.9 291.2 ;
      RECT  93.1 186.4 93.9 187.2 ;
      RECT  167.5 186.4 168.3 187.2 ;
      RECT  152.0 269.6 152.8 270.4 ;
      RECT  93.1 228.0 93.9 228.8 ;
      RECT  152.0 332.0 152.8 332.8 ;
      RECT  108.1 269.6 108.9 270.4 ;
      RECT  167.5 352.8 168.3 353.6 ;
      RECT  108.1 228.0 108.9 228.8 ;
      RECT  152.0 342.4 152.8 343.2 ;
      RECT  190.1 91.4 190.9 92.2 ;
      RECT  108.1 196.8 108.9 197.6 ;
      RECT  203.5 279.6 204.3 280.4 ;
      RECT  190.7 74.0 191.5 74.8 ;
      RECT  93.1 259.2 93.9 260.0 ;
      RECT  183.1 175.6 183.9 176.4 ;
      RECT  176.3 238.0 177.1 238.8 ;
      RECT  167.5 196.8 168.3 197.6 ;
      RECT  167.5 280.0 168.3 280.8 ;
      RECT  167.5 259.2 168.3 260.0 ;
      RECT  203.5 342.0 204.3 342.8 ;
      RECT  176.3 217.2 177.1 218.0 ;
      RECT  192.3 125.4 193.1 126.2 ;
      RECT  167.5 321.6 168.3 322.4 ;
      RECT  176.3 175.6 177.1 176.4 ;
      RECT  176.3 362.8 177.1 363.6 ;
      RECT  196.7 175.6 197.5 176.4 ;
      RECT  167.5 342.4 168.3 343.2 ;
      RECT  203.5 300.4 204.3 301.2 ;
      RECT  197.5 74.0 198.3 74.8 ;
      RECT  152.0 238.4 152.8 239.2 ;
      RECT  176.3 321.2 177.1 322.0 ;
      RECT  167.5 300.8 168.3 301.6 ;
      RECT  108.1 217.6 108.9 218.4 ;
      RECT  176.3 279.6 177.1 280.4 ;
      RECT  93.1 196.8 93.9 197.6 ;
      RECT  176.3 258.8 177.1 259.6 ;
      RECT  176.3 196.4 177.1 197.2 ;
      RECT  93.1 280.0 93.9 280.8 ;
      RECT  167.5 217.6 168.3 218.4 ;
      RECT  203.5 362.8 204.3 363.6 ;
      RECT  196.7 362.8 197.5 363.6 ;
      RECT  203.5 258.8 204.3 259.6 ;
      RECT  189.9 362.8 190.7 363.6 ;
      RECT  199.1 125.4 199.9 126.2 ;
      RECT  167.5 238.4 168.3 239.2 ;
      RECT  93.1 217.6 93.9 218.4 ;
      RECT  203.5 321.2 204.3 322.0 ;
      RECT  197.2 159.6 198.0 160.4 ;
      RECT  108.1 280.0 108.9 280.8 ;
      RECT  203.5 175.6 204.3 176.4 ;
      RECT  152.0 196.8 152.8 197.6 ;
      RECT  152.0 300.8 152.8 301.6 ;
      RECT  203.5 196.4 204.3 197.2 ;
      RECT  176.3 342.0 177.1 342.8 ;
      RECT  203.5 238.0 204.3 238.8 ;
      RECT  152.0 259.2 152.8 260.0 ;
      RECT  203.5 217.2 204.3 218.0 ;
      RECT  152.0 217.6 152.8 218.4 ;
      RECT  152.0 321.6 152.8 322.4 ;
      RECT  152.0 280.0 152.8 280.8 ;
      RECT  183.1 362.8 183.9 363.6 ;
      RECT  196.9 91.4 197.7 92.2 ;
      RECT  176.3 300.4 177.1 301.2 ;
      RECT  183.6 159.6 184.4 160.4 ;
      RECT  108.1 259.2 108.9 260.0 ;
      RECT  190.4 159.6 191.2 160.4 ;
      RECT  189.9 175.6 190.7 176.4 ;
      RECT  200.1 305.4 200.9 306.2 ;
      RECT  200.1 138.8 200.9 139.6 ;
      RECT  200.1 274.6 200.9 275.4 ;
      RECT  206.9 284.6 207.7 285.4 ;
      RECT  200.1 263.8 200.9 264.6 ;
      RECT  209.0 355.0 209.8 355.8 ;
      RECT  179.7 326.2 180.5 327.0 ;
      RECT  93.1 207.2 93.9 208.0 ;
      RECT  179.7 337.0 180.5 337.8 ;
      RECT  179.7 191.4 180.5 192.2 ;
      RECT  193.3 138.8 194.1 139.6 ;
      RECT  152.0 269.6 152.8 270.4 ;
      RECT  152.0 311.2 152.8 312.0 ;
      RECT  206.9 263.8 207.7 264.6 ;
      RECT  179.7 274.6 180.5 275.4 ;
      RECT  200.1 284.6 200.9 285.4 ;
      RECT  193.3 170.6 194.1 171.4 ;
      RECT  179.7 347.0 180.5 347.8 ;
      RECT  200.1 191.4 200.9 192.2 ;
      RECT  167.5 228.0 168.3 228.8 ;
      RECT  200.1 295.4 200.9 296.2 ;
      RECT  179.7 233.0 180.5 233.8 ;
      RECT  172.9 253.8 173.7 254.6 ;
      RECT  179.7 316.2 180.5 317.0 ;
      RECT  206.9 357.8 207.7 358.6 ;
      RECT  93.1 248.8 93.9 249.6 ;
      RECT  200.1 243.0 200.9 243.8 ;
      RECT  167.5 290.4 168.3 291.2 ;
      RECT  93.1 269.6 93.9 270.4 ;
      RECT  190.7 80.6 191.5 81.4 ;
      RECT  200.1 326.2 200.9 327.0 ;
      RECT  206.9 347.0 207.7 347.8 ;
      RECT  200.1 347.0 200.9 347.8 ;
      RECT  206.9 295.4 207.7 296.2 ;
      RECT  179.7 201.4 180.5 202.2 ;
      RECT  172.9 212.2 173.7 213.0 ;
      RECT  192.1 85.0 192.9 85.8 ;
      RECT  172.9 326.2 173.7 327.0 ;
      RECT  172.9 305.4 173.7 306.2 ;
      RECT  179.7 263.8 180.5 264.6 ;
      RECT  108.1 290.4 108.9 291.2 ;
      RECT  179.7 357.8 180.5 358.6 ;
      RECT  93.1 228.0 93.9 228.8 ;
      RECT  198.9 85.0 199.7 85.8 ;
      RECT  193.3 357.8 194.1 358.6 ;
      RECT  172.9 295.4 173.7 296.2 ;
      RECT  93.1 186.4 93.9 187.2 ;
      RECT  197.5 80.6 198.3 81.4 ;
      RECT  186.5 357.8 187.3 358.6 ;
      RECT  179.7 212.2 180.5 213.0 ;
      RECT  209.0 167.8 209.8 168.6 ;
      RECT  206.9 191.4 207.7 192.2 ;
      RECT  167.5 332.0 168.3 332.8 ;
      RECT  200.1 201.4 200.9 202.2 ;
      RECT  172.9 284.6 173.7 285.4 ;
      RECT  206.9 337.0 207.7 337.8 ;
      RECT  206.9 222.2 207.7 223.0 ;
      RECT  206.9 243.0 207.7 243.8 ;
      RECT  152.0 207.2 152.8 208.0 ;
      RECT  152.0 248.8 152.8 249.6 ;
      RECT  172.9 201.4 173.7 202.2 ;
      RECT  152.0 228.0 152.8 228.8 ;
      RECT  196.1 99.6 196.9 100.4 ;
      RECT  108.1 207.2 108.9 208.0 ;
      RECT  206.9 274.6 207.7 275.4 ;
      RECT  167.5 248.8 168.3 249.6 ;
      RECT  170.8 167.8 171.6 168.6 ;
      RECT  179.7 295.4 180.5 296.2 ;
      RECT  172.9 337.0 173.7 337.8 ;
      RECT  172.9 263.8 173.7 264.6 ;
      RECT  206.9 180.6 207.7 181.4 ;
      RECT  206.9 201.4 207.7 202.2 ;
      RECT  179.7 180.6 180.5 181.4 ;
      RECT  179.7 253.8 180.5 254.6 ;
      RECT  200.1 180.6 200.9 181.4 ;
      RECT  172.9 180.6 173.7 181.4 ;
      RECT  172.9 274.6 173.7 275.4 ;
      RECT  172.9 357.8 173.7 358.6 ;
      RECT  200.1 357.8 200.9 358.6 ;
      RECT  172.9 233.0 173.7 233.8 ;
      RECT  152.0 352.8 152.8 353.6 ;
      RECT  172.9 191.4 173.7 192.2 ;
      RECT  200.1 212.2 200.9 213.0 ;
      RECT  179.7 222.2 180.5 223.0 ;
      RECT  206.9 326.2 207.7 327.0 ;
      RECT  172.9 347.0 173.7 347.8 ;
      RECT  167.5 352.8 168.3 353.6 ;
      RECT  152.0 332.0 152.8 332.8 ;
      RECT  93.1 290.4 93.9 291.2 ;
      RECT  108.1 248.8 108.9 249.6 ;
      RECT  179.7 243.0 180.5 243.8 ;
      RECT  172.9 316.2 173.7 317.0 ;
      RECT  200.1 170.6 200.9 171.4 ;
      RECT  200.1 253.8 200.9 254.6 ;
      RECT  200.1 337.0 200.9 337.8 ;
      RECT  152.0 290.4 152.8 291.2 ;
      RECT  206.9 305.4 207.7 306.2 ;
      RECT  108.1 228.0 108.9 228.8 ;
      RECT  167.5 269.6 168.3 270.4 ;
      RECT  172.9 222.2 173.7 223.0 ;
      RECT  206.9 253.8 207.7 254.6 ;
      RECT  108.1 186.4 108.9 187.2 ;
      RECT  206.9 316.2 207.7 317.0 ;
      RECT  206.9 212.2 207.7 213.0 ;
      RECT  179.7 284.6 180.5 285.4 ;
      RECT  179.7 305.4 180.5 306.2 ;
      RECT  186.5 170.6 187.3 171.4 ;
      RECT  167.5 207.2 168.3 208.0 ;
      RECT  200.1 233.0 200.9 233.8 ;
      RECT  108.1 269.6 108.9 270.4 ;
      RECT  206.9 170.6 207.7 171.4 ;
      RECT  200.1 316.2 200.9 317.0 ;
      RECT  179.7 170.6 180.5 171.4 ;
      RECT  167.5 186.4 168.3 187.2 ;
      RECT  172.9 243.0 173.7 243.8 ;
      RECT  200.1 222.2 200.9 223.0 ;
      RECT  189.3 99.6 190.1 100.4 ;
      RECT  206.9 233.0 207.7 233.8 ;
      RECT  172.9 170.6 173.7 171.4 ;
      RECT  167.5 311.2 168.3 312.0 ;
      RECT  152.0 186.4 152.8 187.2 ;
      RECT  170.8 355.0 171.6 355.8 ;
      RECT  2.0 22.4 2.8 23.2 ;
      RECT  2.0 2.4 2.8 3.2 ;
      RECT  2.0 42.4 2.8 43.2 ;
      RECT  10.8 224.0 10.0 224.8 ;
      RECT  10.8 341.6 10.0 342.4 ;
      RECT  24.0 341.6 23.2 342.4 ;
      RECT  24.0 263.2 23.2 264.0 ;
      RECT  24.0 184.8 23.2 185.6 ;
      RECT  10.8 263.2 10.0 264.0 ;
      RECT  24.0 302.4 23.2 303.2 ;
      RECT  24.0 224.0 23.2 224.8 ;
      RECT  10.8 302.4 10.0 303.2 ;
      RECT  10.8 184.8 10.0 185.6 ;
      RECT  24.0 243.6 23.2 244.4 ;
      RECT  10.8 322.0 10.0 322.8 ;
      RECT  24.0 204.4 23.2 205.2 ;
      RECT  10.8 243.6 10.0 244.4 ;
      RECT  10.8 204.4 10.0 205.2 ;
      RECT  24.0 322.0 23.2 322.8 ;
      RECT  24.0 282.8 23.2 283.6 ;
      RECT  24.0 165.2 23.2 166.0 ;
      RECT  10.8 165.2 10.0 166.0 ;
      RECT  10.8 282.8 10.0 283.6 ;
      RECT  10.0 302.4 10.8 303.2 ;
      RECT  10.0 341.6 10.8 342.4 ;
      RECT  2.0 22.4 2.8 23.2 ;
      RECT  77.6 22.4 78.4 23.2 ;
      RECT  77.6 102.4 78.4 103.2 ;
      RECT  10.0 224.0 10.8 224.8 ;
      RECT  77.6 142.4 78.4 143.2 ;
      RECT  23.2 184.8 24.0 185.6 ;
      RECT  23.2 302.4 24.0 303.2 ;
      RECT  23.2 224.0 24.0 224.8 ;
      RECT  23.2 341.6 24.0 342.4 ;
      RECT  10.0 263.2 10.8 264.0 ;
      RECT  23.2 263.2 24.0 264.0 ;
      RECT  77.6 62.4 78.4 63.2 ;
      RECT  10.0 184.8 10.8 185.6 ;
      RECT  10.0 204.4 10.8 205.2 ;
      RECT  77.6 2.4 78.4 3.2 ;
      RECT  77.6 42.4 78.4 43.2 ;
      RECT  77.6 162.4 78.4 163.2 ;
      RECT  77.6 82.4 78.4 83.2 ;
      RECT  23.2 243.6 24.0 244.4 ;
      RECT  10.0 243.6 10.8 244.4 ;
      RECT  23.2 282.8 24.0 283.6 ;
      RECT  23.2 322.0 24.0 322.8 ;
      RECT  77.6 122.4 78.4 123.2 ;
      RECT  23.2 204.4 24.0 205.2 ;
      RECT  2.0 2.4 2.8 3.2 ;
      RECT  10.0 282.8 10.8 283.6 ;
      RECT  10.0 165.2 10.8 166.0 ;
      RECT  2.0 42.4 2.8 43.2 ;
      RECT  23.2 165.2 24.0 166.0 ;
      RECT  10.0 322.0 10.8 322.8 ;
      RECT  57.6 347.9 79.4 348.5 ;
      RECT  68.1 404.4 68.9 405.2 ;
      RECT  68.1 364.4 68.9 365.2 ;
      RECT  68.1 424.4 68.9 425.2 ;
      RECT  68.1 344.4 68.9 345.2 ;
      RECT  68.1 384.4 68.9 385.2 ;
      RECT  101.2 5.9 144.8 6.5 ;
      RECT  111.7 22.4 112.5 23.2 ;
      RECT  133.5 22.4 134.3 23.2 ;
      RECT  133.5 2.4 134.3 3.2 ;
      RECT  111.7 2.4 112.5 3.2 ;
   LAYER  m4 ;
   END
   END    sram_2_16_scn4m_subm
END    LIBRARY
